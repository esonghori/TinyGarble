
module sum_N16384_CC16 ( clk, rst, a, b, c );
  input [1023:0] a;
  input [1023:0] b;
  output [1023:0] c;
  input clk, rst;
  wire   carry_on, carry_on_d, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118;

  DFF carry_on_reg ( .D(carry_on_d), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        carry_on) );
  XOR U4 ( .A(n2), .B(n3), .Z(carry_on_d) );
  ANDN U5 ( .B(n4), .A(n5), .Z(n2) );
  XOR U6 ( .A(b[1023]), .B(n3), .Z(n4) );
  XNOR U7 ( .A(b[9]), .B(n6), .Z(c[9]) );
  XNOR U8 ( .A(b[99]), .B(n7), .Z(c[99]) );
  XNOR U9 ( .A(b[999]), .B(n8), .Z(c[999]) );
  XNOR U10 ( .A(b[998]), .B(n9), .Z(c[998]) );
  XNOR U11 ( .A(b[997]), .B(n10), .Z(c[997]) );
  XNOR U12 ( .A(b[996]), .B(n11), .Z(c[996]) );
  XNOR U13 ( .A(b[995]), .B(n12), .Z(c[995]) );
  XNOR U14 ( .A(b[994]), .B(n13), .Z(c[994]) );
  XNOR U15 ( .A(b[993]), .B(n14), .Z(c[993]) );
  XNOR U16 ( .A(b[992]), .B(n15), .Z(c[992]) );
  XNOR U17 ( .A(b[991]), .B(n16), .Z(c[991]) );
  XNOR U18 ( .A(b[990]), .B(n17), .Z(c[990]) );
  XNOR U19 ( .A(b[98]), .B(n18), .Z(c[98]) );
  XNOR U20 ( .A(b[989]), .B(n19), .Z(c[989]) );
  XNOR U21 ( .A(b[988]), .B(n20), .Z(c[988]) );
  XNOR U22 ( .A(b[987]), .B(n21), .Z(c[987]) );
  XNOR U23 ( .A(b[986]), .B(n22), .Z(c[986]) );
  XNOR U24 ( .A(b[985]), .B(n23), .Z(c[985]) );
  XNOR U25 ( .A(b[984]), .B(n24), .Z(c[984]) );
  XNOR U26 ( .A(b[983]), .B(n25), .Z(c[983]) );
  XNOR U27 ( .A(b[982]), .B(n26), .Z(c[982]) );
  XNOR U28 ( .A(b[981]), .B(n27), .Z(c[981]) );
  XNOR U29 ( .A(b[980]), .B(n28), .Z(c[980]) );
  XNOR U30 ( .A(b[97]), .B(n29), .Z(c[97]) );
  XNOR U31 ( .A(b[979]), .B(n30), .Z(c[979]) );
  XNOR U32 ( .A(b[978]), .B(n31), .Z(c[978]) );
  XNOR U33 ( .A(b[977]), .B(n32), .Z(c[977]) );
  XNOR U34 ( .A(b[976]), .B(n33), .Z(c[976]) );
  XNOR U35 ( .A(b[975]), .B(n34), .Z(c[975]) );
  XNOR U36 ( .A(b[974]), .B(n35), .Z(c[974]) );
  XNOR U37 ( .A(b[973]), .B(n36), .Z(c[973]) );
  XNOR U38 ( .A(b[972]), .B(n37), .Z(c[972]) );
  XNOR U39 ( .A(b[971]), .B(n38), .Z(c[971]) );
  XNOR U40 ( .A(b[970]), .B(n39), .Z(c[970]) );
  XNOR U41 ( .A(b[96]), .B(n40), .Z(c[96]) );
  XNOR U42 ( .A(b[969]), .B(n41), .Z(c[969]) );
  XNOR U43 ( .A(b[968]), .B(n42), .Z(c[968]) );
  XNOR U44 ( .A(b[967]), .B(n43), .Z(c[967]) );
  XNOR U45 ( .A(b[966]), .B(n44), .Z(c[966]) );
  XNOR U46 ( .A(b[965]), .B(n45), .Z(c[965]) );
  XNOR U47 ( .A(b[964]), .B(n46), .Z(c[964]) );
  XNOR U48 ( .A(b[963]), .B(n47), .Z(c[963]) );
  XNOR U49 ( .A(b[962]), .B(n48), .Z(c[962]) );
  XNOR U50 ( .A(b[961]), .B(n49), .Z(c[961]) );
  XNOR U51 ( .A(b[960]), .B(n50), .Z(c[960]) );
  XNOR U52 ( .A(b[95]), .B(n51), .Z(c[95]) );
  XNOR U53 ( .A(b[959]), .B(n52), .Z(c[959]) );
  XNOR U54 ( .A(b[958]), .B(n53), .Z(c[958]) );
  XNOR U55 ( .A(b[957]), .B(n54), .Z(c[957]) );
  XNOR U56 ( .A(b[956]), .B(n55), .Z(c[956]) );
  XNOR U57 ( .A(b[955]), .B(n56), .Z(c[955]) );
  XNOR U58 ( .A(b[954]), .B(n57), .Z(c[954]) );
  XNOR U59 ( .A(b[953]), .B(n58), .Z(c[953]) );
  XNOR U60 ( .A(b[952]), .B(n59), .Z(c[952]) );
  XNOR U61 ( .A(b[951]), .B(n60), .Z(c[951]) );
  XNOR U62 ( .A(b[950]), .B(n61), .Z(c[950]) );
  XNOR U63 ( .A(b[94]), .B(n62), .Z(c[94]) );
  XNOR U64 ( .A(b[949]), .B(n63), .Z(c[949]) );
  XNOR U65 ( .A(b[948]), .B(n64), .Z(c[948]) );
  XNOR U66 ( .A(b[947]), .B(n65), .Z(c[947]) );
  XNOR U67 ( .A(b[946]), .B(n66), .Z(c[946]) );
  XNOR U68 ( .A(b[945]), .B(n67), .Z(c[945]) );
  XNOR U69 ( .A(b[944]), .B(n68), .Z(c[944]) );
  XNOR U70 ( .A(b[943]), .B(n69), .Z(c[943]) );
  XNOR U71 ( .A(b[942]), .B(n70), .Z(c[942]) );
  XNOR U72 ( .A(b[941]), .B(n71), .Z(c[941]) );
  XNOR U73 ( .A(b[940]), .B(n72), .Z(c[940]) );
  XNOR U74 ( .A(b[93]), .B(n73), .Z(c[93]) );
  XNOR U75 ( .A(b[939]), .B(n74), .Z(c[939]) );
  XNOR U76 ( .A(b[938]), .B(n75), .Z(c[938]) );
  XNOR U77 ( .A(b[937]), .B(n76), .Z(c[937]) );
  XNOR U78 ( .A(b[936]), .B(n77), .Z(c[936]) );
  XNOR U79 ( .A(b[935]), .B(n78), .Z(c[935]) );
  XNOR U80 ( .A(b[934]), .B(n79), .Z(c[934]) );
  XNOR U81 ( .A(b[933]), .B(n80), .Z(c[933]) );
  XNOR U82 ( .A(b[932]), .B(n81), .Z(c[932]) );
  XNOR U83 ( .A(b[931]), .B(n82), .Z(c[931]) );
  XNOR U84 ( .A(b[930]), .B(n83), .Z(c[930]) );
  XNOR U85 ( .A(b[92]), .B(n84), .Z(c[92]) );
  XNOR U86 ( .A(b[929]), .B(n85), .Z(c[929]) );
  XNOR U87 ( .A(b[928]), .B(n86), .Z(c[928]) );
  XNOR U88 ( .A(b[927]), .B(n87), .Z(c[927]) );
  XNOR U89 ( .A(b[926]), .B(n88), .Z(c[926]) );
  XNOR U90 ( .A(b[925]), .B(n89), .Z(c[925]) );
  XNOR U91 ( .A(b[924]), .B(n90), .Z(c[924]) );
  XNOR U92 ( .A(b[923]), .B(n91), .Z(c[923]) );
  XNOR U93 ( .A(b[922]), .B(n92), .Z(c[922]) );
  XNOR U94 ( .A(b[921]), .B(n93), .Z(c[921]) );
  XNOR U95 ( .A(b[920]), .B(n94), .Z(c[920]) );
  XNOR U96 ( .A(b[91]), .B(n95), .Z(c[91]) );
  XNOR U97 ( .A(b[919]), .B(n96), .Z(c[919]) );
  XNOR U98 ( .A(b[918]), .B(n97), .Z(c[918]) );
  XNOR U99 ( .A(b[917]), .B(n98), .Z(c[917]) );
  XNOR U100 ( .A(b[916]), .B(n99), .Z(c[916]) );
  XNOR U101 ( .A(b[915]), .B(n100), .Z(c[915]) );
  XNOR U102 ( .A(b[914]), .B(n101), .Z(c[914]) );
  XNOR U103 ( .A(b[913]), .B(n102), .Z(c[913]) );
  XNOR U104 ( .A(b[912]), .B(n103), .Z(c[912]) );
  XNOR U105 ( .A(b[911]), .B(n104), .Z(c[911]) );
  XNOR U106 ( .A(b[910]), .B(n105), .Z(c[910]) );
  XNOR U107 ( .A(b[90]), .B(n106), .Z(c[90]) );
  XNOR U108 ( .A(b[909]), .B(n107), .Z(c[909]) );
  XNOR U109 ( .A(b[908]), .B(n108), .Z(c[908]) );
  XNOR U110 ( .A(b[907]), .B(n109), .Z(c[907]) );
  XNOR U111 ( .A(b[906]), .B(n110), .Z(c[906]) );
  XNOR U112 ( .A(b[905]), .B(n111), .Z(c[905]) );
  XNOR U113 ( .A(b[904]), .B(n112), .Z(c[904]) );
  XNOR U114 ( .A(b[903]), .B(n113), .Z(c[903]) );
  XNOR U115 ( .A(b[902]), .B(n114), .Z(c[902]) );
  XNOR U116 ( .A(b[901]), .B(n115), .Z(c[901]) );
  XNOR U117 ( .A(b[900]), .B(n116), .Z(c[900]) );
  XNOR U118 ( .A(b[8]), .B(n117), .Z(c[8]) );
  XNOR U119 ( .A(b[89]), .B(n118), .Z(c[89]) );
  XNOR U120 ( .A(b[899]), .B(n119), .Z(c[899]) );
  XNOR U121 ( .A(b[898]), .B(n120), .Z(c[898]) );
  XNOR U122 ( .A(b[897]), .B(n121), .Z(c[897]) );
  XNOR U123 ( .A(b[896]), .B(n122), .Z(c[896]) );
  XNOR U124 ( .A(b[895]), .B(n123), .Z(c[895]) );
  XNOR U125 ( .A(b[894]), .B(n124), .Z(c[894]) );
  XNOR U126 ( .A(b[893]), .B(n125), .Z(c[893]) );
  XNOR U127 ( .A(b[892]), .B(n126), .Z(c[892]) );
  XNOR U128 ( .A(b[891]), .B(n127), .Z(c[891]) );
  XNOR U129 ( .A(b[890]), .B(n128), .Z(c[890]) );
  XNOR U130 ( .A(b[88]), .B(n129), .Z(c[88]) );
  XNOR U131 ( .A(b[889]), .B(n130), .Z(c[889]) );
  XNOR U132 ( .A(b[888]), .B(n131), .Z(c[888]) );
  XNOR U133 ( .A(b[887]), .B(n132), .Z(c[887]) );
  XNOR U134 ( .A(b[886]), .B(n133), .Z(c[886]) );
  XNOR U135 ( .A(b[885]), .B(n134), .Z(c[885]) );
  XNOR U136 ( .A(b[884]), .B(n135), .Z(c[884]) );
  XNOR U137 ( .A(b[883]), .B(n136), .Z(c[883]) );
  XNOR U138 ( .A(b[882]), .B(n137), .Z(c[882]) );
  XNOR U139 ( .A(b[881]), .B(n138), .Z(c[881]) );
  XNOR U140 ( .A(b[880]), .B(n139), .Z(c[880]) );
  XNOR U141 ( .A(b[87]), .B(n140), .Z(c[87]) );
  XNOR U142 ( .A(b[879]), .B(n141), .Z(c[879]) );
  XNOR U143 ( .A(b[878]), .B(n142), .Z(c[878]) );
  XNOR U144 ( .A(b[877]), .B(n143), .Z(c[877]) );
  XNOR U145 ( .A(b[876]), .B(n144), .Z(c[876]) );
  XNOR U146 ( .A(b[875]), .B(n145), .Z(c[875]) );
  XNOR U147 ( .A(b[874]), .B(n146), .Z(c[874]) );
  XNOR U148 ( .A(b[873]), .B(n147), .Z(c[873]) );
  XNOR U149 ( .A(b[872]), .B(n148), .Z(c[872]) );
  XNOR U150 ( .A(b[871]), .B(n149), .Z(c[871]) );
  XNOR U151 ( .A(b[870]), .B(n150), .Z(c[870]) );
  XNOR U152 ( .A(b[86]), .B(n151), .Z(c[86]) );
  XNOR U153 ( .A(b[869]), .B(n152), .Z(c[869]) );
  XNOR U154 ( .A(b[868]), .B(n153), .Z(c[868]) );
  XNOR U155 ( .A(b[867]), .B(n154), .Z(c[867]) );
  XNOR U156 ( .A(b[866]), .B(n155), .Z(c[866]) );
  XNOR U157 ( .A(b[865]), .B(n156), .Z(c[865]) );
  XNOR U158 ( .A(b[864]), .B(n157), .Z(c[864]) );
  XNOR U159 ( .A(b[863]), .B(n158), .Z(c[863]) );
  XNOR U160 ( .A(b[862]), .B(n159), .Z(c[862]) );
  XNOR U161 ( .A(b[861]), .B(n160), .Z(c[861]) );
  XNOR U162 ( .A(b[860]), .B(n161), .Z(c[860]) );
  XNOR U163 ( .A(b[85]), .B(n162), .Z(c[85]) );
  XNOR U164 ( .A(b[859]), .B(n163), .Z(c[859]) );
  XNOR U165 ( .A(b[858]), .B(n164), .Z(c[858]) );
  XNOR U166 ( .A(b[857]), .B(n165), .Z(c[857]) );
  XNOR U167 ( .A(b[856]), .B(n166), .Z(c[856]) );
  XNOR U168 ( .A(b[855]), .B(n167), .Z(c[855]) );
  XNOR U169 ( .A(b[854]), .B(n168), .Z(c[854]) );
  XNOR U170 ( .A(b[853]), .B(n169), .Z(c[853]) );
  XNOR U171 ( .A(b[852]), .B(n170), .Z(c[852]) );
  XNOR U172 ( .A(b[851]), .B(n171), .Z(c[851]) );
  XNOR U173 ( .A(b[850]), .B(n172), .Z(c[850]) );
  XNOR U174 ( .A(b[84]), .B(n173), .Z(c[84]) );
  XNOR U175 ( .A(b[849]), .B(n174), .Z(c[849]) );
  XNOR U176 ( .A(b[848]), .B(n175), .Z(c[848]) );
  XNOR U177 ( .A(b[847]), .B(n176), .Z(c[847]) );
  XNOR U178 ( .A(b[846]), .B(n177), .Z(c[846]) );
  XNOR U179 ( .A(b[845]), .B(n178), .Z(c[845]) );
  XNOR U180 ( .A(b[844]), .B(n179), .Z(c[844]) );
  XNOR U181 ( .A(b[843]), .B(n180), .Z(c[843]) );
  XNOR U182 ( .A(b[842]), .B(n181), .Z(c[842]) );
  XNOR U183 ( .A(b[841]), .B(n182), .Z(c[841]) );
  XNOR U184 ( .A(b[840]), .B(n183), .Z(c[840]) );
  XNOR U185 ( .A(b[83]), .B(n184), .Z(c[83]) );
  XNOR U186 ( .A(b[839]), .B(n185), .Z(c[839]) );
  XNOR U187 ( .A(b[838]), .B(n186), .Z(c[838]) );
  XNOR U188 ( .A(b[837]), .B(n187), .Z(c[837]) );
  XNOR U189 ( .A(b[836]), .B(n188), .Z(c[836]) );
  XNOR U190 ( .A(b[835]), .B(n189), .Z(c[835]) );
  XNOR U191 ( .A(b[834]), .B(n190), .Z(c[834]) );
  XNOR U192 ( .A(b[833]), .B(n191), .Z(c[833]) );
  XNOR U193 ( .A(b[832]), .B(n192), .Z(c[832]) );
  XNOR U194 ( .A(b[831]), .B(n193), .Z(c[831]) );
  XNOR U195 ( .A(b[830]), .B(n194), .Z(c[830]) );
  XNOR U196 ( .A(b[82]), .B(n195), .Z(c[82]) );
  XNOR U197 ( .A(b[829]), .B(n196), .Z(c[829]) );
  XNOR U198 ( .A(b[828]), .B(n197), .Z(c[828]) );
  XNOR U199 ( .A(b[827]), .B(n198), .Z(c[827]) );
  XNOR U200 ( .A(b[826]), .B(n199), .Z(c[826]) );
  XNOR U201 ( .A(b[825]), .B(n200), .Z(c[825]) );
  XNOR U202 ( .A(b[824]), .B(n201), .Z(c[824]) );
  XNOR U203 ( .A(b[823]), .B(n202), .Z(c[823]) );
  XNOR U204 ( .A(b[822]), .B(n203), .Z(c[822]) );
  XNOR U205 ( .A(b[821]), .B(n204), .Z(c[821]) );
  XNOR U206 ( .A(b[820]), .B(n205), .Z(c[820]) );
  XNOR U207 ( .A(b[81]), .B(n206), .Z(c[81]) );
  XNOR U208 ( .A(b[819]), .B(n207), .Z(c[819]) );
  XNOR U209 ( .A(b[818]), .B(n208), .Z(c[818]) );
  XNOR U210 ( .A(b[817]), .B(n209), .Z(c[817]) );
  XNOR U211 ( .A(b[816]), .B(n210), .Z(c[816]) );
  XNOR U212 ( .A(b[815]), .B(n211), .Z(c[815]) );
  XNOR U213 ( .A(b[814]), .B(n212), .Z(c[814]) );
  XNOR U214 ( .A(b[813]), .B(n213), .Z(c[813]) );
  XNOR U215 ( .A(b[812]), .B(n214), .Z(c[812]) );
  XNOR U216 ( .A(b[811]), .B(n215), .Z(c[811]) );
  XNOR U217 ( .A(b[810]), .B(n216), .Z(c[810]) );
  XNOR U218 ( .A(b[80]), .B(n217), .Z(c[80]) );
  XNOR U219 ( .A(b[809]), .B(n218), .Z(c[809]) );
  XNOR U220 ( .A(b[808]), .B(n219), .Z(c[808]) );
  XNOR U221 ( .A(b[807]), .B(n220), .Z(c[807]) );
  XNOR U222 ( .A(b[806]), .B(n221), .Z(c[806]) );
  XNOR U223 ( .A(b[805]), .B(n222), .Z(c[805]) );
  XNOR U224 ( .A(b[804]), .B(n223), .Z(c[804]) );
  XNOR U225 ( .A(b[803]), .B(n224), .Z(c[803]) );
  XNOR U226 ( .A(b[802]), .B(n225), .Z(c[802]) );
  XNOR U227 ( .A(b[801]), .B(n226), .Z(c[801]) );
  XNOR U228 ( .A(b[800]), .B(n227), .Z(c[800]) );
  XNOR U229 ( .A(b[7]), .B(n228), .Z(c[7]) );
  XNOR U230 ( .A(b[79]), .B(n229), .Z(c[79]) );
  XNOR U231 ( .A(b[799]), .B(n230), .Z(c[799]) );
  XNOR U232 ( .A(b[798]), .B(n231), .Z(c[798]) );
  XNOR U233 ( .A(b[797]), .B(n232), .Z(c[797]) );
  XNOR U234 ( .A(b[796]), .B(n233), .Z(c[796]) );
  XNOR U235 ( .A(b[795]), .B(n234), .Z(c[795]) );
  XNOR U236 ( .A(b[794]), .B(n235), .Z(c[794]) );
  XNOR U237 ( .A(b[793]), .B(n236), .Z(c[793]) );
  XNOR U238 ( .A(b[792]), .B(n237), .Z(c[792]) );
  XNOR U239 ( .A(b[791]), .B(n238), .Z(c[791]) );
  XNOR U240 ( .A(b[790]), .B(n239), .Z(c[790]) );
  XNOR U241 ( .A(b[78]), .B(n240), .Z(c[78]) );
  XNOR U242 ( .A(b[789]), .B(n241), .Z(c[789]) );
  XNOR U243 ( .A(b[788]), .B(n242), .Z(c[788]) );
  XNOR U244 ( .A(b[787]), .B(n243), .Z(c[787]) );
  XNOR U245 ( .A(b[786]), .B(n244), .Z(c[786]) );
  XNOR U246 ( .A(b[785]), .B(n245), .Z(c[785]) );
  XNOR U247 ( .A(b[784]), .B(n246), .Z(c[784]) );
  XNOR U248 ( .A(b[783]), .B(n247), .Z(c[783]) );
  XNOR U249 ( .A(b[782]), .B(n248), .Z(c[782]) );
  XNOR U250 ( .A(b[781]), .B(n249), .Z(c[781]) );
  XNOR U251 ( .A(b[780]), .B(n250), .Z(c[780]) );
  XNOR U252 ( .A(b[77]), .B(n251), .Z(c[77]) );
  XNOR U253 ( .A(b[779]), .B(n252), .Z(c[779]) );
  XNOR U254 ( .A(b[778]), .B(n253), .Z(c[778]) );
  XNOR U255 ( .A(b[777]), .B(n254), .Z(c[777]) );
  XNOR U256 ( .A(b[776]), .B(n255), .Z(c[776]) );
  XNOR U257 ( .A(b[775]), .B(n256), .Z(c[775]) );
  XNOR U258 ( .A(b[774]), .B(n257), .Z(c[774]) );
  XNOR U259 ( .A(b[773]), .B(n258), .Z(c[773]) );
  XNOR U260 ( .A(b[772]), .B(n259), .Z(c[772]) );
  XNOR U261 ( .A(b[771]), .B(n260), .Z(c[771]) );
  XNOR U262 ( .A(b[770]), .B(n261), .Z(c[770]) );
  XNOR U263 ( .A(b[76]), .B(n262), .Z(c[76]) );
  XNOR U264 ( .A(b[769]), .B(n263), .Z(c[769]) );
  XNOR U265 ( .A(b[768]), .B(n264), .Z(c[768]) );
  XNOR U266 ( .A(b[767]), .B(n265), .Z(c[767]) );
  XNOR U267 ( .A(b[766]), .B(n266), .Z(c[766]) );
  XNOR U268 ( .A(b[765]), .B(n267), .Z(c[765]) );
  XNOR U269 ( .A(b[764]), .B(n268), .Z(c[764]) );
  XNOR U270 ( .A(b[763]), .B(n269), .Z(c[763]) );
  XNOR U271 ( .A(b[762]), .B(n270), .Z(c[762]) );
  XNOR U272 ( .A(b[761]), .B(n271), .Z(c[761]) );
  XNOR U273 ( .A(b[760]), .B(n272), .Z(c[760]) );
  XNOR U274 ( .A(b[75]), .B(n273), .Z(c[75]) );
  XNOR U275 ( .A(b[759]), .B(n274), .Z(c[759]) );
  XNOR U276 ( .A(b[758]), .B(n275), .Z(c[758]) );
  XNOR U277 ( .A(b[757]), .B(n276), .Z(c[757]) );
  XNOR U278 ( .A(b[756]), .B(n277), .Z(c[756]) );
  XNOR U279 ( .A(b[755]), .B(n278), .Z(c[755]) );
  XNOR U280 ( .A(b[754]), .B(n279), .Z(c[754]) );
  XNOR U281 ( .A(b[753]), .B(n280), .Z(c[753]) );
  XNOR U282 ( .A(b[752]), .B(n281), .Z(c[752]) );
  XNOR U283 ( .A(b[751]), .B(n282), .Z(c[751]) );
  XNOR U284 ( .A(b[750]), .B(n283), .Z(c[750]) );
  XNOR U285 ( .A(b[74]), .B(n284), .Z(c[74]) );
  XNOR U286 ( .A(b[749]), .B(n285), .Z(c[749]) );
  XNOR U287 ( .A(b[748]), .B(n286), .Z(c[748]) );
  XNOR U288 ( .A(b[747]), .B(n287), .Z(c[747]) );
  XNOR U289 ( .A(b[746]), .B(n288), .Z(c[746]) );
  XNOR U290 ( .A(b[745]), .B(n289), .Z(c[745]) );
  XNOR U291 ( .A(b[744]), .B(n290), .Z(c[744]) );
  XNOR U292 ( .A(b[743]), .B(n291), .Z(c[743]) );
  XNOR U293 ( .A(b[742]), .B(n292), .Z(c[742]) );
  XNOR U294 ( .A(b[741]), .B(n293), .Z(c[741]) );
  XNOR U295 ( .A(b[740]), .B(n294), .Z(c[740]) );
  XNOR U296 ( .A(b[73]), .B(n295), .Z(c[73]) );
  XNOR U297 ( .A(b[739]), .B(n296), .Z(c[739]) );
  XNOR U298 ( .A(b[738]), .B(n297), .Z(c[738]) );
  XNOR U299 ( .A(b[737]), .B(n298), .Z(c[737]) );
  XNOR U300 ( .A(b[736]), .B(n299), .Z(c[736]) );
  XNOR U301 ( .A(b[735]), .B(n300), .Z(c[735]) );
  XNOR U302 ( .A(b[734]), .B(n301), .Z(c[734]) );
  XNOR U303 ( .A(b[733]), .B(n302), .Z(c[733]) );
  XNOR U304 ( .A(b[732]), .B(n303), .Z(c[732]) );
  XNOR U305 ( .A(b[731]), .B(n304), .Z(c[731]) );
  XNOR U306 ( .A(b[730]), .B(n305), .Z(c[730]) );
  XNOR U307 ( .A(b[72]), .B(n306), .Z(c[72]) );
  XNOR U308 ( .A(b[729]), .B(n307), .Z(c[729]) );
  XNOR U309 ( .A(b[728]), .B(n308), .Z(c[728]) );
  XNOR U310 ( .A(b[727]), .B(n309), .Z(c[727]) );
  XNOR U311 ( .A(b[726]), .B(n310), .Z(c[726]) );
  XNOR U312 ( .A(b[725]), .B(n311), .Z(c[725]) );
  XNOR U313 ( .A(b[724]), .B(n312), .Z(c[724]) );
  XNOR U314 ( .A(b[723]), .B(n313), .Z(c[723]) );
  XNOR U315 ( .A(b[722]), .B(n314), .Z(c[722]) );
  XNOR U316 ( .A(b[721]), .B(n315), .Z(c[721]) );
  XNOR U317 ( .A(b[720]), .B(n316), .Z(c[720]) );
  XNOR U318 ( .A(b[71]), .B(n317), .Z(c[71]) );
  XNOR U319 ( .A(b[719]), .B(n318), .Z(c[719]) );
  XNOR U320 ( .A(b[718]), .B(n319), .Z(c[718]) );
  XNOR U321 ( .A(b[717]), .B(n320), .Z(c[717]) );
  XNOR U322 ( .A(b[716]), .B(n321), .Z(c[716]) );
  XNOR U323 ( .A(b[715]), .B(n322), .Z(c[715]) );
  XNOR U324 ( .A(b[714]), .B(n323), .Z(c[714]) );
  XNOR U325 ( .A(b[713]), .B(n324), .Z(c[713]) );
  XNOR U326 ( .A(b[712]), .B(n325), .Z(c[712]) );
  XNOR U327 ( .A(b[711]), .B(n326), .Z(c[711]) );
  XNOR U328 ( .A(b[710]), .B(n327), .Z(c[710]) );
  XNOR U329 ( .A(b[70]), .B(n328), .Z(c[70]) );
  XNOR U330 ( .A(b[709]), .B(n329), .Z(c[709]) );
  XNOR U331 ( .A(b[708]), .B(n330), .Z(c[708]) );
  XNOR U332 ( .A(b[707]), .B(n331), .Z(c[707]) );
  XNOR U333 ( .A(b[706]), .B(n332), .Z(c[706]) );
  XNOR U334 ( .A(b[705]), .B(n333), .Z(c[705]) );
  XNOR U335 ( .A(b[704]), .B(n334), .Z(c[704]) );
  XNOR U336 ( .A(b[703]), .B(n335), .Z(c[703]) );
  XNOR U337 ( .A(b[702]), .B(n336), .Z(c[702]) );
  XNOR U338 ( .A(b[701]), .B(n337), .Z(c[701]) );
  XNOR U339 ( .A(b[700]), .B(n338), .Z(c[700]) );
  XNOR U340 ( .A(b[6]), .B(n339), .Z(c[6]) );
  XNOR U341 ( .A(b[69]), .B(n340), .Z(c[69]) );
  XNOR U342 ( .A(b[699]), .B(n341), .Z(c[699]) );
  XNOR U343 ( .A(b[698]), .B(n342), .Z(c[698]) );
  XNOR U344 ( .A(b[697]), .B(n343), .Z(c[697]) );
  XNOR U345 ( .A(b[696]), .B(n344), .Z(c[696]) );
  XNOR U346 ( .A(b[695]), .B(n345), .Z(c[695]) );
  XNOR U347 ( .A(b[694]), .B(n346), .Z(c[694]) );
  XNOR U348 ( .A(b[693]), .B(n347), .Z(c[693]) );
  XNOR U349 ( .A(b[692]), .B(n348), .Z(c[692]) );
  XNOR U350 ( .A(b[691]), .B(n349), .Z(c[691]) );
  XNOR U351 ( .A(b[690]), .B(n350), .Z(c[690]) );
  XNOR U352 ( .A(b[68]), .B(n351), .Z(c[68]) );
  XNOR U353 ( .A(b[689]), .B(n352), .Z(c[689]) );
  XNOR U354 ( .A(b[688]), .B(n353), .Z(c[688]) );
  XNOR U355 ( .A(b[687]), .B(n354), .Z(c[687]) );
  XNOR U356 ( .A(b[686]), .B(n355), .Z(c[686]) );
  XNOR U357 ( .A(b[685]), .B(n356), .Z(c[685]) );
  XNOR U358 ( .A(b[684]), .B(n357), .Z(c[684]) );
  XNOR U359 ( .A(b[683]), .B(n358), .Z(c[683]) );
  XNOR U360 ( .A(b[682]), .B(n359), .Z(c[682]) );
  XNOR U361 ( .A(b[681]), .B(n360), .Z(c[681]) );
  XNOR U362 ( .A(b[680]), .B(n361), .Z(c[680]) );
  XNOR U363 ( .A(b[67]), .B(n362), .Z(c[67]) );
  XNOR U364 ( .A(b[679]), .B(n363), .Z(c[679]) );
  XNOR U365 ( .A(b[678]), .B(n364), .Z(c[678]) );
  XNOR U366 ( .A(b[677]), .B(n365), .Z(c[677]) );
  XNOR U367 ( .A(b[676]), .B(n366), .Z(c[676]) );
  XNOR U368 ( .A(b[675]), .B(n367), .Z(c[675]) );
  XNOR U369 ( .A(b[674]), .B(n368), .Z(c[674]) );
  XNOR U370 ( .A(b[673]), .B(n369), .Z(c[673]) );
  XNOR U371 ( .A(b[672]), .B(n370), .Z(c[672]) );
  XNOR U372 ( .A(b[671]), .B(n371), .Z(c[671]) );
  XNOR U373 ( .A(b[670]), .B(n372), .Z(c[670]) );
  XNOR U374 ( .A(b[66]), .B(n373), .Z(c[66]) );
  XNOR U375 ( .A(b[669]), .B(n374), .Z(c[669]) );
  XNOR U376 ( .A(b[668]), .B(n375), .Z(c[668]) );
  XNOR U377 ( .A(b[667]), .B(n376), .Z(c[667]) );
  XNOR U378 ( .A(b[666]), .B(n377), .Z(c[666]) );
  XNOR U379 ( .A(b[665]), .B(n378), .Z(c[665]) );
  XNOR U380 ( .A(b[664]), .B(n379), .Z(c[664]) );
  XNOR U381 ( .A(b[663]), .B(n380), .Z(c[663]) );
  XNOR U382 ( .A(b[662]), .B(n381), .Z(c[662]) );
  XNOR U383 ( .A(b[661]), .B(n382), .Z(c[661]) );
  XNOR U384 ( .A(b[660]), .B(n383), .Z(c[660]) );
  XNOR U385 ( .A(b[65]), .B(n384), .Z(c[65]) );
  XNOR U386 ( .A(b[659]), .B(n385), .Z(c[659]) );
  XNOR U387 ( .A(b[658]), .B(n386), .Z(c[658]) );
  XNOR U388 ( .A(b[657]), .B(n387), .Z(c[657]) );
  XNOR U389 ( .A(b[656]), .B(n388), .Z(c[656]) );
  XNOR U390 ( .A(b[655]), .B(n389), .Z(c[655]) );
  XNOR U391 ( .A(b[654]), .B(n390), .Z(c[654]) );
  XNOR U392 ( .A(b[653]), .B(n391), .Z(c[653]) );
  XNOR U393 ( .A(b[652]), .B(n392), .Z(c[652]) );
  XNOR U394 ( .A(b[651]), .B(n393), .Z(c[651]) );
  XNOR U395 ( .A(b[650]), .B(n394), .Z(c[650]) );
  XNOR U396 ( .A(b[64]), .B(n395), .Z(c[64]) );
  XNOR U397 ( .A(b[649]), .B(n396), .Z(c[649]) );
  XNOR U398 ( .A(b[648]), .B(n397), .Z(c[648]) );
  XNOR U399 ( .A(b[647]), .B(n398), .Z(c[647]) );
  XNOR U400 ( .A(b[646]), .B(n399), .Z(c[646]) );
  XNOR U401 ( .A(b[645]), .B(n400), .Z(c[645]) );
  XNOR U402 ( .A(b[644]), .B(n401), .Z(c[644]) );
  XNOR U403 ( .A(b[643]), .B(n402), .Z(c[643]) );
  XNOR U404 ( .A(b[642]), .B(n403), .Z(c[642]) );
  XNOR U405 ( .A(b[641]), .B(n404), .Z(c[641]) );
  XNOR U406 ( .A(b[640]), .B(n405), .Z(c[640]) );
  XNOR U407 ( .A(b[63]), .B(n406), .Z(c[63]) );
  XNOR U408 ( .A(b[639]), .B(n407), .Z(c[639]) );
  XNOR U409 ( .A(b[638]), .B(n408), .Z(c[638]) );
  XNOR U410 ( .A(b[637]), .B(n409), .Z(c[637]) );
  XNOR U411 ( .A(b[636]), .B(n410), .Z(c[636]) );
  XNOR U412 ( .A(b[635]), .B(n411), .Z(c[635]) );
  XNOR U413 ( .A(b[634]), .B(n412), .Z(c[634]) );
  XNOR U414 ( .A(b[633]), .B(n413), .Z(c[633]) );
  XNOR U415 ( .A(b[632]), .B(n414), .Z(c[632]) );
  XNOR U416 ( .A(b[631]), .B(n415), .Z(c[631]) );
  XNOR U417 ( .A(b[630]), .B(n416), .Z(c[630]) );
  XNOR U418 ( .A(b[62]), .B(n417), .Z(c[62]) );
  XNOR U419 ( .A(b[629]), .B(n418), .Z(c[629]) );
  XNOR U420 ( .A(b[628]), .B(n419), .Z(c[628]) );
  XNOR U421 ( .A(b[627]), .B(n420), .Z(c[627]) );
  XNOR U422 ( .A(b[626]), .B(n421), .Z(c[626]) );
  XNOR U423 ( .A(b[625]), .B(n422), .Z(c[625]) );
  XNOR U424 ( .A(b[624]), .B(n423), .Z(c[624]) );
  XNOR U425 ( .A(b[623]), .B(n424), .Z(c[623]) );
  XNOR U426 ( .A(b[622]), .B(n425), .Z(c[622]) );
  XNOR U427 ( .A(b[621]), .B(n426), .Z(c[621]) );
  XNOR U428 ( .A(b[620]), .B(n427), .Z(c[620]) );
  XNOR U429 ( .A(b[61]), .B(n428), .Z(c[61]) );
  XNOR U430 ( .A(b[619]), .B(n429), .Z(c[619]) );
  XNOR U431 ( .A(b[618]), .B(n430), .Z(c[618]) );
  XNOR U432 ( .A(b[617]), .B(n431), .Z(c[617]) );
  XNOR U433 ( .A(b[616]), .B(n432), .Z(c[616]) );
  XNOR U434 ( .A(b[615]), .B(n433), .Z(c[615]) );
  XNOR U435 ( .A(b[614]), .B(n434), .Z(c[614]) );
  XNOR U436 ( .A(b[613]), .B(n435), .Z(c[613]) );
  XNOR U437 ( .A(b[612]), .B(n436), .Z(c[612]) );
  XNOR U438 ( .A(b[611]), .B(n437), .Z(c[611]) );
  XNOR U439 ( .A(b[610]), .B(n438), .Z(c[610]) );
  XNOR U440 ( .A(b[60]), .B(n439), .Z(c[60]) );
  XNOR U441 ( .A(b[609]), .B(n440), .Z(c[609]) );
  XNOR U442 ( .A(b[608]), .B(n441), .Z(c[608]) );
  XNOR U443 ( .A(b[607]), .B(n442), .Z(c[607]) );
  XNOR U444 ( .A(b[606]), .B(n443), .Z(c[606]) );
  XNOR U445 ( .A(b[605]), .B(n444), .Z(c[605]) );
  XNOR U446 ( .A(b[604]), .B(n445), .Z(c[604]) );
  XNOR U447 ( .A(b[603]), .B(n446), .Z(c[603]) );
  XNOR U448 ( .A(b[602]), .B(n447), .Z(c[602]) );
  XNOR U449 ( .A(b[601]), .B(n448), .Z(c[601]) );
  XNOR U450 ( .A(b[600]), .B(n449), .Z(c[600]) );
  XNOR U451 ( .A(b[5]), .B(n450), .Z(c[5]) );
  XNOR U452 ( .A(b[59]), .B(n451), .Z(c[59]) );
  XNOR U453 ( .A(b[599]), .B(n452), .Z(c[599]) );
  XNOR U454 ( .A(b[598]), .B(n453), .Z(c[598]) );
  XNOR U455 ( .A(b[597]), .B(n454), .Z(c[597]) );
  XNOR U456 ( .A(b[596]), .B(n455), .Z(c[596]) );
  XNOR U457 ( .A(b[595]), .B(n456), .Z(c[595]) );
  XNOR U458 ( .A(b[594]), .B(n457), .Z(c[594]) );
  XNOR U459 ( .A(b[593]), .B(n458), .Z(c[593]) );
  XNOR U460 ( .A(b[592]), .B(n459), .Z(c[592]) );
  XNOR U461 ( .A(b[591]), .B(n460), .Z(c[591]) );
  XNOR U462 ( .A(b[590]), .B(n461), .Z(c[590]) );
  XNOR U463 ( .A(b[58]), .B(n462), .Z(c[58]) );
  XNOR U464 ( .A(b[589]), .B(n463), .Z(c[589]) );
  XNOR U465 ( .A(b[588]), .B(n464), .Z(c[588]) );
  XNOR U466 ( .A(b[587]), .B(n465), .Z(c[587]) );
  XNOR U467 ( .A(b[586]), .B(n466), .Z(c[586]) );
  XNOR U468 ( .A(b[585]), .B(n467), .Z(c[585]) );
  XNOR U469 ( .A(b[584]), .B(n468), .Z(c[584]) );
  XNOR U470 ( .A(b[583]), .B(n469), .Z(c[583]) );
  XNOR U471 ( .A(b[582]), .B(n470), .Z(c[582]) );
  XNOR U472 ( .A(b[581]), .B(n471), .Z(c[581]) );
  XNOR U473 ( .A(b[580]), .B(n472), .Z(c[580]) );
  XNOR U474 ( .A(b[57]), .B(n473), .Z(c[57]) );
  XNOR U475 ( .A(b[579]), .B(n474), .Z(c[579]) );
  XNOR U476 ( .A(b[578]), .B(n475), .Z(c[578]) );
  XNOR U477 ( .A(b[577]), .B(n476), .Z(c[577]) );
  XNOR U478 ( .A(b[576]), .B(n477), .Z(c[576]) );
  XNOR U479 ( .A(b[575]), .B(n478), .Z(c[575]) );
  XNOR U480 ( .A(b[574]), .B(n479), .Z(c[574]) );
  XNOR U481 ( .A(b[573]), .B(n480), .Z(c[573]) );
  XNOR U482 ( .A(b[572]), .B(n481), .Z(c[572]) );
  XNOR U483 ( .A(b[571]), .B(n482), .Z(c[571]) );
  XNOR U484 ( .A(b[570]), .B(n483), .Z(c[570]) );
  XNOR U485 ( .A(b[56]), .B(n484), .Z(c[56]) );
  XNOR U486 ( .A(b[569]), .B(n485), .Z(c[569]) );
  XNOR U487 ( .A(b[568]), .B(n486), .Z(c[568]) );
  XNOR U488 ( .A(b[567]), .B(n487), .Z(c[567]) );
  XNOR U489 ( .A(b[566]), .B(n488), .Z(c[566]) );
  XNOR U490 ( .A(b[565]), .B(n489), .Z(c[565]) );
  XNOR U491 ( .A(b[564]), .B(n490), .Z(c[564]) );
  XNOR U492 ( .A(b[563]), .B(n491), .Z(c[563]) );
  XNOR U493 ( .A(b[562]), .B(n492), .Z(c[562]) );
  XNOR U494 ( .A(b[561]), .B(n493), .Z(c[561]) );
  XNOR U495 ( .A(b[560]), .B(n494), .Z(c[560]) );
  XNOR U496 ( .A(b[55]), .B(n495), .Z(c[55]) );
  XNOR U497 ( .A(b[559]), .B(n496), .Z(c[559]) );
  XNOR U498 ( .A(b[558]), .B(n497), .Z(c[558]) );
  XNOR U499 ( .A(b[557]), .B(n498), .Z(c[557]) );
  XNOR U500 ( .A(b[556]), .B(n499), .Z(c[556]) );
  XNOR U501 ( .A(b[555]), .B(n500), .Z(c[555]) );
  XNOR U502 ( .A(b[554]), .B(n501), .Z(c[554]) );
  XNOR U503 ( .A(b[553]), .B(n502), .Z(c[553]) );
  XNOR U504 ( .A(b[552]), .B(n503), .Z(c[552]) );
  XNOR U505 ( .A(b[551]), .B(n504), .Z(c[551]) );
  XNOR U506 ( .A(b[550]), .B(n505), .Z(c[550]) );
  XNOR U507 ( .A(b[54]), .B(n506), .Z(c[54]) );
  XNOR U508 ( .A(b[549]), .B(n507), .Z(c[549]) );
  XNOR U509 ( .A(b[548]), .B(n508), .Z(c[548]) );
  XNOR U510 ( .A(b[547]), .B(n509), .Z(c[547]) );
  XNOR U511 ( .A(b[546]), .B(n510), .Z(c[546]) );
  XNOR U512 ( .A(b[545]), .B(n511), .Z(c[545]) );
  XNOR U513 ( .A(b[544]), .B(n512), .Z(c[544]) );
  XNOR U514 ( .A(b[543]), .B(n513), .Z(c[543]) );
  XNOR U515 ( .A(b[542]), .B(n514), .Z(c[542]) );
  XNOR U516 ( .A(b[541]), .B(n515), .Z(c[541]) );
  XNOR U517 ( .A(b[540]), .B(n516), .Z(c[540]) );
  XNOR U518 ( .A(b[53]), .B(n517), .Z(c[53]) );
  XNOR U519 ( .A(b[539]), .B(n518), .Z(c[539]) );
  XNOR U520 ( .A(b[538]), .B(n519), .Z(c[538]) );
  XNOR U521 ( .A(b[537]), .B(n520), .Z(c[537]) );
  XNOR U522 ( .A(b[536]), .B(n521), .Z(c[536]) );
  XNOR U523 ( .A(b[535]), .B(n522), .Z(c[535]) );
  XNOR U524 ( .A(b[534]), .B(n523), .Z(c[534]) );
  XNOR U525 ( .A(b[533]), .B(n524), .Z(c[533]) );
  XNOR U526 ( .A(b[532]), .B(n525), .Z(c[532]) );
  XNOR U527 ( .A(b[531]), .B(n526), .Z(c[531]) );
  XNOR U528 ( .A(b[530]), .B(n527), .Z(c[530]) );
  XNOR U529 ( .A(b[52]), .B(n528), .Z(c[52]) );
  XNOR U530 ( .A(b[529]), .B(n529), .Z(c[529]) );
  XNOR U531 ( .A(b[528]), .B(n530), .Z(c[528]) );
  XNOR U532 ( .A(b[527]), .B(n531), .Z(c[527]) );
  XNOR U533 ( .A(b[526]), .B(n532), .Z(c[526]) );
  XNOR U534 ( .A(b[525]), .B(n533), .Z(c[525]) );
  XNOR U535 ( .A(b[524]), .B(n534), .Z(c[524]) );
  XNOR U536 ( .A(b[523]), .B(n535), .Z(c[523]) );
  XNOR U537 ( .A(b[522]), .B(n536), .Z(c[522]) );
  XNOR U538 ( .A(b[521]), .B(n537), .Z(c[521]) );
  XNOR U539 ( .A(b[520]), .B(n538), .Z(c[520]) );
  XNOR U540 ( .A(b[51]), .B(n539), .Z(c[51]) );
  XNOR U541 ( .A(b[519]), .B(n540), .Z(c[519]) );
  XNOR U542 ( .A(b[518]), .B(n541), .Z(c[518]) );
  XNOR U543 ( .A(b[517]), .B(n542), .Z(c[517]) );
  XNOR U544 ( .A(b[516]), .B(n543), .Z(c[516]) );
  XNOR U545 ( .A(b[515]), .B(n544), .Z(c[515]) );
  XNOR U546 ( .A(b[514]), .B(n545), .Z(c[514]) );
  XNOR U547 ( .A(b[513]), .B(n546), .Z(c[513]) );
  XNOR U548 ( .A(b[512]), .B(n547), .Z(c[512]) );
  XNOR U549 ( .A(b[511]), .B(n548), .Z(c[511]) );
  XNOR U550 ( .A(b[510]), .B(n549), .Z(c[510]) );
  XNOR U551 ( .A(b[50]), .B(n550), .Z(c[50]) );
  XNOR U552 ( .A(b[509]), .B(n551), .Z(c[509]) );
  XNOR U553 ( .A(b[508]), .B(n552), .Z(c[508]) );
  XNOR U554 ( .A(b[507]), .B(n553), .Z(c[507]) );
  XNOR U555 ( .A(b[506]), .B(n554), .Z(c[506]) );
  XNOR U556 ( .A(b[505]), .B(n555), .Z(c[505]) );
  XNOR U557 ( .A(b[504]), .B(n556), .Z(c[504]) );
  XNOR U558 ( .A(b[503]), .B(n557), .Z(c[503]) );
  XNOR U559 ( .A(b[502]), .B(n558), .Z(c[502]) );
  XNOR U560 ( .A(b[501]), .B(n559), .Z(c[501]) );
  XNOR U561 ( .A(b[500]), .B(n560), .Z(c[500]) );
  XNOR U562 ( .A(b[4]), .B(n561), .Z(c[4]) );
  XNOR U563 ( .A(b[49]), .B(n562), .Z(c[49]) );
  XNOR U564 ( .A(b[499]), .B(n563), .Z(c[499]) );
  XNOR U565 ( .A(b[498]), .B(n564), .Z(c[498]) );
  XNOR U566 ( .A(b[497]), .B(n565), .Z(c[497]) );
  XNOR U567 ( .A(b[496]), .B(n566), .Z(c[496]) );
  XNOR U568 ( .A(b[495]), .B(n567), .Z(c[495]) );
  XNOR U569 ( .A(b[494]), .B(n568), .Z(c[494]) );
  XNOR U570 ( .A(b[493]), .B(n569), .Z(c[493]) );
  XNOR U571 ( .A(b[492]), .B(n570), .Z(c[492]) );
  XNOR U572 ( .A(b[491]), .B(n571), .Z(c[491]) );
  XNOR U573 ( .A(b[490]), .B(n572), .Z(c[490]) );
  XNOR U574 ( .A(b[48]), .B(n573), .Z(c[48]) );
  XNOR U575 ( .A(b[489]), .B(n574), .Z(c[489]) );
  XNOR U576 ( .A(b[488]), .B(n575), .Z(c[488]) );
  XNOR U577 ( .A(b[487]), .B(n576), .Z(c[487]) );
  XNOR U578 ( .A(b[486]), .B(n577), .Z(c[486]) );
  XNOR U579 ( .A(b[485]), .B(n578), .Z(c[485]) );
  XNOR U580 ( .A(b[484]), .B(n579), .Z(c[484]) );
  XNOR U581 ( .A(b[483]), .B(n580), .Z(c[483]) );
  XNOR U582 ( .A(b[482]), .B(n581), .Z(c[482]) );
  XNOR U583 ( .A(b[481]), .B(n582), .Z(c[481]) );
  XNOR U584 ( .A(b[480]), .B(n583), .Z(c[480]) );
  XNOR U585 ( .A(b[47]), .B(n584), .Z(c[47]) );
  XNOR U586 ( .A(b[479]), .B(n585), .Z(c[479]) );
  XNOR U587 ( .A(b[478]), .B(n586), .Z(c[478]) );
  XNOR U588 ( .A(b[477]), .B(n587), .Z(c[477]) );
  XNOR U589 ( .A(b[476]), .B(n588), .Z(c[476]) );
  XNOR U590 ( .A(b[475]), .B(n589), .Z(c[475]) );
  XNOR U591 ( .A(b[474]), .B(n590), .Z(c[474]) );
  XNOR U592 ( .A(b[473]), .B(n591), .Z(c[473]) );
  XNOR U593 ( .A(b[472]), .B(n592), .Z(c[472]) );
  XNOR U594 ( .A(b[471]), .B(n593), .Z(c[471]) );
  XNOR U595 ( .A(b[470]), .B(n594), .Z(c[470]) );
  XNOR U596 ( .A(b[46]), .B(n595), .Z(c[46]) );
  XNOR U597 ( .A(b[469]), .B(n596), .Z(c[469]) );
  XNOR U598 ( .A(b[468]), .B(n597), .Z(c[468]) );
  XNOR U599 ( .A(b[467]), .B(n598), .Z(c[467]) );
  XNOR U600 ( .A(b[466]), .B(n599), .Z(c[466]) );
  XNOR U601 ( .A(b[465]), .B(n600), .Z(c[465]) );
  XNOR U602 ( .A(b[464]), .B(n601), .Z(c[464]) );
  XNOR U603 ( .A(b[463]), .B(n602), .Z(c[463]) );
  XNOR U604 ( .A(b[462]), .B(n603), .Z(c[462]) );
  XNOR U605 ( .A(b[461]), .B(n604), .Z(c[461]) );
  XNOR U606 ( .A(b[460]), .B(n605), .Z(c[460]) );
  XNOR U607 ( .A(b[45]), .B(n606), .Z(c[45]) );
  XNOR U608 ( .A(b[459]), .B(n607), .Z(c[459]) );
  XNOR U609 ( .A(b[458]), .B(n608), .Z(c[458]) );
  XNOR U610 ( .A(b[457]), .B(n609), .Z(c[457]) );
  XNOR U611 ( .A(b[456]), .B(n610), .Z(c[456]) );
  XNOR U612 ( .A(b[455]), .B(n611), .Z(c[455]) );
  XNOR U613 ( .A(b[454]), .B(n612), .Z(c[454]) );
  XNOR U614 ( .A(b[453]), .B(n613), .Z(c[453]) );
  XNOR U615 ( .A(b[452]), .B(n614), .Z(c[452]) );
  XNOR U616 ( .A(b[451]), .B(n615), .Z(c[451]) );
  XNOR U617 ( .A(b[450]), .B(n616), .Z(c[450]) );
  XNOR U618 ( .A(b[44]), .B(n617), .Z(c[44]) );
  XNOR U619 ( .A(b[449]), .B(n618), .Z(c[449]) );
  XNOR U620 ( .A(b[448]), .B(n619), .Z(c[448]) );
  XNOR U621 ( .A(b[447]), .B(n620), .Z(c[447]) );
  XNOR U622 ( .A(b[446]), .B(n621), .Z(c[446]) );
  XNOR U623 ( .A(b[445]), .B(n622), .Z(c[445]) );
  XNOR U624 ( .A(b[444]), .B(n623), .Z(c[444]) );
  XNOR U625 ( .A(b[443]), .B(n624), .Z(c[443]) );
  XNOR U626 ( .A(b[442]), .B(n625), .Z(c[442]) );
  XNOR U627 ( .A(b[441]), .B(n626), .Z(c[441]) );
  XNOR U628 ( .A(b[440]), .B(n627), .Z(c[440]) );
  XNOR U629 ( .A(b[43]), .B(n628), .Z(c[43]) );
  XNOR U630 ( .A(b[439]), .B(n629), .Z(c[439]) );
  XNOR U631 ( .A(b[438]), .B(n630), .Z(c[438]) );
  XNOR U632 ( .A(b[437]), .B(n631), .Z(c[437]) );
  XNOR U633 ( .A(b[436]), .B(n632), .Z(c[436]) );
  XNOR U634 ( .A(b[435]), .B(n633), .Z(c[435]) );
  XNOR U635 ( .A(b[434]), .B(n634), .Z(c[434]) );
  XNOR U636 ( .A(b[433]), .B(n635), .Z(c[433]) );
  XNOR U637 ( .A(b[432]), .B(n636), .Z(c[432]) );
  XNOR U638 ( .A(b[431]), .B(n637), .Z(c[431]) );
  XNOR U639 ( .A(b[430]), .B(n638), .Z(c[430]) );
  XNOR U640 ( .A(b[42]), .B(n639), .Z(c[42]) );
  XNOR U641 ( .A(b[429]), .B(n640), .Z(c[429]) );
  XNOR U642 ( .A(b[428]), .B(n641), .Z(c[428]) );
  XNOR U643 ( .A(b[427]), .B(n642), .Z(c[427]) );
  XNOR U644 ( .A(b[426]), .B(n643), .Z(c[426]) );
  XNOR U645 ( .A(b[425]), .B(n644), .Z(c[425]) );
  XNOR U646 ( .A(b[424]), .B(n645), .Z(c[424]) );
  XNOR U647 ( .A(b[423]), .B(n646), .Z(c[423]) );
  XNOR U648 ( .A(b[422]), .B(n647), .Z(c[422]) );
  XNOR U649 ( .A(b[421]), .B(n648), .Z(c[421]) );
  XNOR U650 ( .A(b[420]), .B(n649), .Z(c[420]) );
  XNOR U651 ( .A(b[41]), .B(n650), .Z(c[41]) );
  XNOR U652 ( .A(b[419]), .B(n651), .Z(c[419]) );
  XNOR U653 ( .A(b[418]), .B(n652), .Z(c[418]) );
  XNOR U654 ( .A(b[417]), .B(n653), .Z(c[417]) );
  XNOR U655 ( .A(b[416]), .B(n654), .Z(c[416]) );
  XNOR U656 ( .A(b[415]), .B(n655), .Z(c[415]) );
  XNOR U657 ( .A(b[414]), .B(n656), .Z(c[414]) );
  XNOR U658 ( .A(b[413]), .B(n657), .Z(c[413]) );
  XNOR U659 ( .A(b[412]), .B(n658), .Z(c[412]) );
  XNOR U660 ( .A(b[411]), .B(n659), .Z(c[411]) );
  XNOR U661 ( .A(b[410]), .B(n660), .Z(c[410]) );
  XNOR U662 ( .A(b[40]), .B(n661), .Z(c[40]) );
  XNOR U663 ( .A(b[409]), .B(n662), .Z(c[409]) );
  XNOR U664 ( .A(b[408]), .B(n663), .Z(c[408]) );
  XNOR U665 ( .A(b[407]), .B(n664), .Z(c[407]) );
  XNOR U666 ( .A(b[406]), .B(n665), .Z(c[406]) );
  XNOR U667 ( .A(b[405]), .B(n666), .Z(c[405]) );
  XNOR U668 ( .A(b[404]), .B(n667), .Z(c[404]) );
  XNOR U669 ( .A(b[403]), .B(n668), .Z(c[403]) );
  XNOR U670 ( .A(b[402]), .B(n669), .Z(c[402]) );
  XNOR U671 ( .A(b[401]), .B(n670), .Z(c[401]) );
  XNOR U672 ( .A(b[400]), .B(n671), .Z(c[400]) );
  XNOR U673 ( .A(b[3]), .B(n672), .Z(c[3]) );
  XNOR U674 ( .A(b[39]), .B(n673), .Z(c[39]) );
  XNOR U675 ( .A(b[399]), .B(n674), .Z(c[399]) );
  XNOR U676 ( .A(b[398]), .B(n675), .Z(c[398]) );
  XNOR U677 ( .A(b[397]), .B(n676), .Z(c[397]) );
  XNOR U678 ( .A(b[396]), .B(n677), .Z(c[396]) );
  XNOR U679 ( .A(b[395]), .B(n678), .Z(c[395]) );
  XNOR U680 ( .A(b[394]), .B(n679), .Z(c[394]) );
  XNOR U681 ( .A(b[393]), .B(n680), .Z(c[393]) );
  XNOR U682 ( .A(b[392]), .B(n681), .Z(c[392]) );
  XNOR U683 ( .A(b[391]), .B(n682), .Z(c[391]) );
  XNOR U684 ( .A(b[390]), .B(n683), .Z(c[390]) );
  XNOR U685 ( .A(b[38]), .B(n684), .Z(c[38]) );
  XNOR U686 ( .A(b[389]), .B(n685), .Z(c[389]) );
  XNOR U687 ( .A(b[388]), .B(n686), .Z(c[388]) );
  XNOR U688 ( .A(b[387]), .B(n687), .Z(c[387]) );
  XNOR U689 ( .A(b[386]), .B(n688), .Z(c[386]) );
  XNOR U690 ( .A(b[385]), .B(n689), .Z(c[385]) );
  XNOR U691 ( .A(b[384]), .B(n690), .Z(c[384]) );
  XNOR U692 ( .A(b[383]), .B(n691), .Z(c[383]) );
  XNOR U693 ( .A(b[382]), .B(n692), .Z(c[382]) );
  XNOR U694 ( .A(b[381]), .B(n693), .Z(c[381]) );
  XNOR U695 ( .A(b[380]), .B(n694), .Z(c[380]) );
  XNOR U696 ( .A(b[37]), .B(n695), .Z(c[37]) );
  XNOR U697 ( .A(b[379]), .B(n696), .Z(c[379]) );
  XNOR U698 ( .A(b[378]), .B(n697), .Z(c[378]) );
  XNOR U699 ( .A(b[377]), .B(n698), .Z(c[377]) );
  XNOR U700 ( .A(b[376]), .B(n699), .Z(c[376]) );
  XNOR U701 ( .A(b[375]), .B(n700), .Z(c[375]) );
  XNOR U702 ( .A(b[374]), .B(n701), .Z(c[374]) );
  XNOR U703 ( .A(b[373]), .B(n702), .Z(c[373]) );
  XNOR U704 ( .A(b[372]), .B(n703), .Z(c[372]) );
  XNOR U705 ( .A(b[371]), .B(n704), .Z(c[371]) );
  XNOR U706 ( .A(b[370]), .B(n705), .Z(c[370]) );
  XNOR U707 ( .A(b[36]), .B(n706), .Z(c[36]) );
  XNOR U708 ( .A(b[369]), .B(n707), .Z(c[369]) );
  XNOR U709 ( .A(b[368]), .B(n708), .Z(c[368]) );
  XNOR U710 ( .A(b[367]), .B(n709), .Z(c[367]) );
  XNOR U711 ( .A(b[366]), .B(n710), .Z(c[366]) );
  XNOR U712 ( .A(b[365]), .B(n711), .Z(c[365]) );
  XNOR U713 ( .A(b[364]), .B(n712), .Z(c[364]) );
  XNOR U714 ( .A(b[363]), .B(n713), .Z(c[363]) );
  XNOR U715 ( .A(b[362]), .B(n714), .Z(c[362]) );
  XNOR U716 ( .A(b[361]), .B(n715), .Z(c[361]) );
  XNOR U717 ( .A(b[360]), .B(n716), .Z(c[360]) );
  XNOR U718 ( .A(b[35]), .B(n717), .Z(c[35]) );
  XNOR U719 ( .A(b[359]), .B(n718), .Z(c[359]) );
  XNOR U720 ( .A(b[358]), .B(n719), .Z(c[358]) );
  XNOR U721 ( .A(b[357]), .B(n720), .Z(c[357]) );
  XNOR U722 ( .A(b[356]), .B(n721), .Z(c[356]) );
  XNOR U723 ( .A(b[355]), .B(n722), .Z(c[355]) );
  XNOR U724 ( .A(b[354]), .B(n723), .Z(c[354]) );
  XNOR U725 ( .A(b[353]), .B(n724), .Z(c[353]) );
  XNOR U726 ( .A(b[352]), .B(n725), .Z(c[352]) );
  XNOR U727 ( .A(b[351]), .B(n726), .Z(c[351]) );
  XNOR U728 ( .A(b[350]), .B(n727), .Z(c[350]) );
  XNOR U729 ( .A(b[34]), .B(n728), .Z(c[34]) );
  XNOR U730 ( .A(b[349]), .B(n729), .Z(c[349]) );
  XNOR U731 ( .A(b[348]), .B(n730), .Z(c[348]) );
  XNOR U732 ( .A(b[347]), .B(n731), .Z(c[347]) );
  XNOR U733 ( .A(b[346]), .B(n732), .Z(c[346]) );
  XNOR U734 ( .A(b[345]), .B(n733), .Z(c[345]) );
  XNOR U735 ( .A(b[344]), .B(n734), .Z(c[344]) );
  XNOR U736 ( .A(b[343]), .B(n735), .Z(c[343]) );
  XNOR U737 ( .A(b[342]), .B(n736), .Z(c[342]) );
  XNOR U738 ( .A(b[341]), .B(n737), .Z(c[341]) );
  XNOR U739 ( .A(b[340]), .B(n738), .Z(c[340]) );
  XNOR U740 ( .A(b[33]), .B(n739), .Z(c[33]) );
  XNOR U741 ( .A(b[339]), .B(n740), .Z(c[339]) );
  XNOR U742 ( .A(b[338]), .B(n741), .Z(c[338]) );
  XNOR U743 ( .A(b[337]), .B(n742), .Z(c[337]) );
  XNOR U744 ( .A(b[336]), .B(n743), .Z(c[336]) );
  XNOR U745 ( .A(b[335]), .B(n744), .Z(c[335]) );
  XNOR U746 ( .A(b[334]), .B(n745), .Z(c[334]) );
  XNOR U747 ( .A(b[333]), .B(n746), .Z(c[333]) );
  XNOR U748 ( .A(b[332]), .B(n747), .Z(c[332]) );
  XNOR U749 ( .A(b[331]), .B(n748), .Z(c[331]) );
  XNOR U750 ( .A(b[330]), .B(n749), .Z(c[330]) );
  XNOR U751 ( .A(b[32]), .B(n750), .Z(c[32]) );
  XNOR U752 ( .A(b[329]), .B(n751), .Z(c[329]) );
  XNOR U753 ( .A(b[328]), .B(n752), .Z(c[328]) );
  XNOR U754 ( .A(b[327]), .B(n753), .Z(c[327]) );
  XNOR U755 ( .A(b[326]), .B(n754), .Z(c[326]) );
  XNOR U756 ( .A(b[325]), .B(n755), .Z(c[325]) );
  XNOR U757 ( .A(b[324]), .B(n756), .Z(c[324]) );
  XNOR U758 ( .A(b[323]), .B(n757), .Z(c[323]) );
  XNOR U759 ( .A(b[322]), .B(n758), .Z(c[322]) );
  XNOR U760 ( .A(b[321]), .B(n759), .Z(c[321]) );
  XNOR U761 ( .A(b[320]), .B(n760), .Z(c[320]) );
  XNOR U762 ( .A(b[31]), .B(n761), .Z(c[31]) );
  XNOR U763 ( .A(b[319]), .B(n762), .Z(c[319]) );
  XNOR U764 ( .A(b[318]), .B(n763), .Z(c[318]) );
  XNOR U765 ( .A(b[317]), .B(n764), .Z(c[317]) );
  XNOR U766 ( .A(b[316]), .B(n765), .Z(c[316]) );
  XNOR U767 ( .A(b[315]), .B(n766), .Z(c[315]) );
  XNOR U768 ( .A(b[314]), .B(n767), .Z(c[314]) );
  XNOR U769 ( .A(b[313]), .B(n768), .Z(c[313]) );
  XNOR U770 ( .A(b[312]), .B(n769), .Z(c[312]) );
  XNOR U771 ( .A(b[311]), .B(n770), .Z(c[311]) );
  XNOR U772 ( .A(b[310]), .B(n771), .Z(c[310]) );
  XNOR U773 ( .A(b[30]), .B(n772), .Z(c[30]) );
  XNOR U774 ( .A(b[309]), .B(n773), .Z(c[309]) );
  XNOR U775 ( .A(b[308]), .B(n774), .Z(c[308]) );
  XNOR U776 ( .A(b[307]), .B(n775), .Z(c[307]) );
  XNOR U777 ( .A(b[306]), .B(n776), .Z(c[306]) );
  XNOR U778 ( .A(b[305]), .B(n777), .Z(c[305]) );
  XNOR U779 ( .A(b[304]), .B(n778), .Z(c[304]) );
  XNOR U780 ( .A(b[303]), .B(n779), .Z(c[303]) );
  XNOR U781 ( .A(b[302]), .B(n780), .Z(c[302]) );
  XNOR U782 ( .A(b[301]), .B(n781), .Z(c[301]) );
  XNOR U783 ( .A(b[300]), .B(n782), .Z(c[300]) );
  XNOR U784 ( .A(b[2]), .B(n783), .Z(c[2]) );
  XNOR U785 ( .A(b[29]), .B(n784), .Z(c[29]) );
  XNOR U786 ( .A(b[299]), .B(n785), .Z(c[299]) );
  XNOR U787 ( .A(b[298]), .B(n786), .Z(c[298]) );
  XNOR U788 ( .A(b[297]), .B(n787), .Z(c[297]) );
  XNOR U789 ( .A(b[296]), .B(n788), .Z(c[296]) );
  XNOR U790 ( .A(b[295]), .B(n789), .Z(c[295]) );
  XNOR U791 ( .A(b[294]), .B(n790), .Z(c[294]) );
  XNOR U792 ( .A(b[293]), .B(n791), .Z(c[293]) );
  XNOR U793 ( .A(b[292]), .B(n792), .Z(c[292]) );
  XNOR U794 ( .A(b[291]), .B(n793), .Z(c[291]) );
  XNOR U795 ( .A(b[290]), .B(n794), .Z(c[290]) );
  XNOR U796 ( .A(b[28]), .B(n795), .Z(c[28]) );
  XNOR U797 ( .A(b[289]), .B(n796), .Z(c[289]) );
  XNOR U798 ( .A(b[288]), .B(n797), .Z(c[288]) );
  XNOR U799 ( .A(b[287]), .B(n798), .Z(c[287]) );
  XNOR U800 ( .A(b[286]), .B(n799), .Z(c[286]) );
  XNOR U801 ( .A(b[285]), .B(n800), .Z(c[285]) );
  XNOR U802 ( .A(b[284]), .B(n801), .Z(c[284]) );
  XNOR U803 ( .A(b[283]), .B(n802), .Z(c[283]) );
  XNOR U804 ( .A(b[282]), .B(n803), .Z(c[282]) );
  XNOR U805 ( .A(b[281]), .B(n804), .Z(c[281]) );
  XNOR U806 ( .A(b[280]), .B(n805), .Z(c[280]) );
  XNOR U807 ( .A(b[27]), .B(n806), .Z(c[27]) );
  XNOR U808 ( .A(b[279]), .B(n807), .Z(c[279]) );
  XNOR U809 ( .A(b[278]), .B(n808), .Z(c[278]) );
  XNOR U810 ( .A(b[277]), .B(n809), .Z(c[277]) );
  XNOR U811 ( .A(b[276]), .B(n810), .Z(c[276]) );
  XNOR U812 ( .A(b[275]), .B(n811), .Z(c[275]) );
  XNOR U813 ( .A(b[274]), .B(n812), .Z(c[274]) );
  XNOR U814 ( .A(b[273]), .B(n813), .Z(c[273]) );
  XNOR U815 ( .A(b[272]), .B(n814), .Z(c[272]) );
  XNOR U816 ( .A(b[271]), .B(n815), .Z(c[271]) );
  XNOR U817 ( .A(b[270]), .B(n816), .Z(c[270]) );
  XNOR U818 ( .A(b[26]), .B(n817), .Z(c[26]) );
  XNOR U819 ( .A(b[269]), .B(n818), .Z(c[269]) );
  XNOR U820 ( .A(b[268]), .B(n819), .Z(c[268]) );
  XNOR U821 ( .A(b[267]), .B(n820), .Z(c[267]) );
  XNOR U822 ( .A(b[266]), .B(n821), .Z(c[266]) );
  XNOR U823 ( .A(b[265]), .B(n822), .Z(c[265]) );
  XNOR U824 ( .A(b[264]), .B(n823), .Z(c[264]) );
  XNOR U825 ( .A(b[263]), .B(n824), .Z(c[263]) );
  XNOR U826 ( .A(b[262]), .B(n825), .Z(c[262]) );
  XNOR U827 ( .A(b[261]), .B(n826), .Z(c[261]) );
  XNOR U828 ( .A(b[260]), .B(n827), .Z(c[260]) );
  XNOR U829 ( .A(b[25]), .B(n828), .Z(c[25]) );
  XNOR U830 ( .A(b[259]), .B(n829), .Z(c[259]) );
  XNOR U831 ( .A(b[258]), .B(n830), .Z(c[258]) );
  XNOR U832 ( .A(b[257]), .B(n831), .Z(c[257]) );
  XNOR U833 ( .A(b[256]), .B(n832), .Z(c[256]) );
  XNOR U834 ( .A(b[255]), .B(n833), .Z(c[255]) );
  XNOR U835 ( .A(b[254]), .B(n834), .Z(c[254]) );
  XNOR U836 ( .A(b[253]), .B(n835), .Z(c[253]) );
  XNOR U837 ( .A(b[252]), .B(n836), .Z(c[252]) );
  XNOR U838 ( .A(b[251]), .B(n837), .Z(c[251]) );
  XNOR U839 ( .A(b[250]), .B(n838), .Z(c[250]) );
  XNOR U840 ( .A(b[24]), .B(n839), .Z(c[24]) );
  XNOR U841 ( .A(b[249]), .B(n840), .Z(c[249]) );
  XNOR U842 ( .A(b[248]), .B(n841), .Z(c[248]) );
  XNOR U843 ( .A(b[247]), .B(n842), .Z(c[247]) );
  XNOR U844 ( .A(b[246]), .B(n843), .Z(c[246]) );
  XNOR U845 ( .A(b[245]), .B(n844), .Z(c[245]) );
  XNOR U846 ( .A(b[244]), .B(n845), .Z(c[244]) );
  XNOR U847 ( .A(b[243]), .B(n846), .Z(c[243]) );
  XNOR U848 ( .A(b[242]), .B(n847), .Z(c[242]) );
  XNOR U849 ( .A(b[241]), .B(n848), .Z(c[241]) );
  XNOR U850 ( .A(b[240]), .B(n849), .Z(c[240]) );
  XNOR U851 ( .A(b[23]), .B(n850), .Z(c[23]) );
  XNOR U852 ( .A(b[239]), .B(n851), .Z(c[239]) );
  XNOR U853 ( .A(b[238]), .B(n852), .Z(c[238]) );
  XNOR U854 ( .A(b[237]), .B(n853), .Z(c[237]) );
  XNOR U855 ( .A(b[236]), .B(n854), .Z(c[236]) );
  XNOR U856 ( .A(b[235]), .B(n855), .Z(c[235]) );
  XNOR U857 ( .A(b[234]), .B(n856), .Z(c[234]) );
  XNOR U858 ( .A(b[233]), .B(n857), .Z(c[233]) );
  XNOR U859 ( .A(b[232]), .B(n858), .Z(c[232]) );
  XNOR U860 ( .A(b[231]), .B(n859), .Z(c[231]) );
  XNOR U861 ( .A(b[230]), .B(n860), .Z(c[230]) );
  XNOR U862 ( .A(b[22]), .B(n861), .Z(c[22]) );
  XNOR U863 ( .A(b[229]), .B(n862), .Z(c[229]) );
  XNOR U864 ( .A(b[228]), .B(n863), .Z(c[228]) );
  XNOR U865 ( .A(b[227]), .B(n864), .Z(c[227]) );
  XNOR U866 ( .A(b[226]), .B(n865), .Z(c[226]) );
  XNOR U867 ( .A(b[225]), .B(n866), .Z(c[225]) );
  XNOR U868 ( .A(b[224]), .B(n867), .Z(c[224]) );
  XNOR U869 ( .A(b[223]), .B(n868), .Z(c[223]) );
  XNOR U870 ( .A(b[222]), .B(n869), .Z(c[222]) );
  XNOR U871 ( .A(b[221]), .B(n870), .Z(c[221]) );
  XNOR U872 ( .A(b[220]), .B(n871), .Z(c[220]) );
  XNOR U873 ( .A(b[21]), .B(n872), .Z(c[21]) );
  XNOR U874 ( .A(b[219]), .B(n873), .Z(c[219]) );
  XNOR U875 ( .A(b[218]), .B(n874), .Z(c[218]) );
  XNOR U876 ( .A(b[217]), .B(n875), .Z(c[217]) );
  XNOR U877 ( .A(b[216]), .B(n876), .Z(c[216]) );
  XNOR U878 ( .A(b[215]), .B(n877), .Z(c[215]) );
  XNOR U879 ( .A(b[214]), .B(n878), .Z(c[214]) );
  XNOR U880 ( .A(b[213]), .B(n879), .Z(c[213]) );
  XNOR U881 ( .A(b[212]), .B(n880), .Z(c[212]) );
  XNOR U882 ( .A(b[211]), .B(n881), .Z(c[211]) );
  XNOR U883 ( .A(b[210]), .B(n882), .Z(c[210]) );
  XNOR U884 ( .A(b[20]), .B(n883), .Z(c[20]) );
  XNOR U885 ( .A(b[209]), .B(n884), .Z(c[209]) );
  XNOR U886 ( .A(b[208]), .B(n885), .Z(c[208]) );
  XNOR U887 ( .A(b[207]), .B(n886), .Z(c[207]) );
  XNOR U888 ( .A(b[206]), .B(n887), .Z(c[206]) );
  XNOR U889 ( .A(b[205]), .B(n888), .Z(c[205]) );
  XNOR U890 ( .A(b[204]), .B(n889), .Z(c[204]) );
  XNOR U891 ( .A(b[203]), .B(n890), .Z(c[203]) );
  XNOR U892 ( .A(b[202]), .B(n891), .Z(c[202]) );
  XNOR U893 ( .A(b[201]), .B(n892), .Z(c[201]) );
  XNOR U894 ( .A(b[200]), .B(n893), .Z(c[200]) );
  XNOR U895 ( .A(b[1]), .B(n894), .Z(c[1]) );
  XNOR U896 ( .A(b[19]), .B(n895), .Z(c[19]) );
  XNOR U897 ( .A(b[199]), .B(n896), .Z(c[199]) );
  XNOR U898 ( .A(b[198]), .B(n897), .Z(c[198]) );
  XNOR U899 ( .A(b[197]), .B(n898), .Z(c[197]) );
  XNOR U900 ( .A(b[196]), .B(n899), .Z(c[196]) );
  XNOR U901 ( .A(b[195]), .B(n900), .Z(c[195]) );
  XNOR U902 ( .A(b[194]), .B(n901), .Z(c[194]) );
  XNOR U903 ( .A(b[193]), .B(n902), .Z(c[193]) );
  XNOR U904 ( .A(b[192]), .B(n903), .Z(c[192]) );
  XNOR U905 ( .A(b[191]), .B(n904), .Z(c[191]) );
  XNOR U906 ( .A(b[190]), .B(n905), .Z(c[190]) );
  XNOR U907 ( .A(b[18]), .B(n906), .Z(c[18]) );
  XNOR U908 ( .A(b[189]), .B(n907), .Z(c[189]) );
  XNOR U909 ( .A(b[188]), .B(n908), .Z(c[188]) );
  XNOR U910 ( .A(b[187]), .B(n909), .Z(c[187]) );
  XNOR U911 ( .A(b[186]), .B(n910), .Z(c[186]) );
  XNOR U912 ( .A(b[185]), .B(n911), .Z(c[185]) );
  XNOR U913 ( .A(b[184]), .B(n912), .Z(c[184]) );
  XNOR U914 ( .A(b[183]), .B(n913), .Z(c[183]) );
  XNOR U915 ( .A(b[182]), .B(n914), .Z(c[182]) );
  XNOR U916 ( .A(b[181]), .B(n915), .Z(c[181]) );
  XNOR U917 ( .A(b[180]), .B(n916), .Z(c[180]) );
  XNOR U918 ( .A(b[17]), .B(n917), .Z(c[17]) );
  XNOR U919 ( .A(b[179]), .B(n918), .Z(c[179]) );
  XNOR U920 ( .A(b[178]), .B(n919), .Z(c[178]) );
  XNOR U921 ( .A(b[177]), .B(n920), .Z(c[177]) );
  XNOR U922 ( .A(b[176]), .B(n921), .Z(c[176]) );
  XNOR U923 ( .A(b[175]), .B(n922), .Z(c[175]) );
  XNOR U924 ( .A(b[174]), .B(n923), .Z(c[174]) );
  XNOR U925 ( .A(b[173]), .B(n924), .Z(c[173]) );
  XNOR U926 ( .A(b[172]), .B(n925), .Z(c[172]) );
  XNOR U927 ( .A(b[171]), .B(n926), .Z(c[171]) );
  XNOR U928 ( .A(b[170]), .B(n927), .Z(c[170]) );
  XNOR U929 ( .A(b[16]), .B(n928), .Z(c[16]) );
  XNOR U930 ( .A(b[169]), .B(n929), .Z(c[169]) );
  XNOR U931 ( .A(b[168]), .B(n930), .Z(c[168]) );
  XNOR U932 ( .A(b[167]), .B(n931), .Z(c[167]) );
  XNOR U933 ( .A(b[166]), .B(n932), .Z(c[166]) );
  XNOR U934 ( .A(b[165]), .B(n933), .Z(c[165]) );
  XNOR U935 ( .A(b[164]), .B(n934), .Z(c[164]) );
  XNOR U936 ( .A(b[163]), .B(n935), .Z(c[163]) );
  XNOR U937 ( .A(b[162]), .B(n936), .Z(c[162]) );
  XNOR U938 ( .A(b[161]), .B(n937), .Z(c[161]) );
  XNOR U939 ( .A(b[160]), .B(n938), .Z(c[160]) );
  XNOR U940 ( .A(b[15]), .B(n939), .Z(c[15]) );
  XNOR U941 ( .A(b[159]), .B(n940), .Z(c[159]) );
  XNOR U942 ( .A(b[158]), .B(n941), .Z(c[158]) );
  XNOR U943 ( .A(b[157]), .B(n942), .Z(c[157]) );
  XNOR U944 ( .A(b[156]), .B(n943), .Z(c[156]) );
  XNOR U945 ( .A(b[155]), .B(n944), .Z(c[155]) );
  XNOR U946 ( .A(b[154]), .B(n945), .Z(c[154]) );
  XNOR U947 ( .A(b[153]), .B(n946), .Z(c[153]) );
  XNOR U948 ( .A(b[152]), .B(n947), .Z(c[152]) );
  XNOR U949 ( .A(b[151]), .B(n948), .Z(c[151]) );
  XNOR U950 ( .A(b[150]), .B(n949), .Z(c[150]) );
  XNOR U951 ( .A(b[14]), .B(n950), .Z(c[14]) );
  XNOR U952 ( .A(b[149]), .B(n951), .Z(c[149]) );
  XNOR U953 ( .A(b[148]), .B(n952), .Z(c[148]) );
  XNOR U954 ( .A(b[147]), .B(n953), .Z(c[147]) );
  XNOR U955 ( .A(b[146]), .B(n954), .Z(c[146]) );
  XNOR U956 ( .A(b[145]), .B(n955), .Z(c[145]) );
  XNOR U957 ( .A(b[144]), .B(n956), .Z(c[144]) );
  XNOR U958 ( .A(b[143]), .B(n957), .Z(c[143]) );
  XNOR U959 ( .A(b[142]), .B(n958), .Z(c[142]) );
  XNOR U960 ( .A(b[141]), .B(n959), .Z(c[141]) );
  XNOR U961 ( .A(b[140]), .B(n960), .Z(c[140]) );
  XNOR U962 ( .A(b[13]), .B(n961), .Z(c[13]) );
  XNOR U963 ( .A(b[139]), .B(n962), .Z(c[139]) );
  XNOR U964 ( .A(b[138]), .B(n963), .Z(c[138]) );
  XNOR U965 ( .A(b[137]), .B(n964), .Z(c[137]) );
  XNOR U966 ( .A(b[136]), .B(n965), .Z(c[136]) );
  XNOR U967 ( .A(b[135]), .B(n966), .Z(c[135]) );
  XNOR U968 ( .A(b[134]), .B(n967), .Z(c[134]) );
  XNOR U969 ( .A(b[133]), .B(n968), .Z(c[133]) );
  XNOR U970 ( .A(b[132]), .B(n969), .Z(c[132]) );
  XNOR U971 ( .A(b[131]), .B(n970), .Z(c[131]) );
  XNOR U972 ( .A(b[130]), .B(n971), .Z(c[130]) );
  XNOR U973 ( .A(b[12]), .B(n972), .Z(c[12]) );
  XNOR U974 ( .A(b[129]), .B(n973), .Z(c[129]) );
  XNOR U975 ( .A(b[128]), .B(n974), .Z(c[128]) );
  XNOR U976 ( .A(b[127]), .B(n975), .Z(c[127]) );
  XNOR U977 ( .A(b[126]), .B(n976), .Z(c[126]) );
  XNOR U978 ( .A(b[125]), .B(n977), .Z(c[125]) );
  XNOR U979 ( .A(b[124]), .B(n978), .Z(c[124]) );
  XNOR U980 ( .A(b[123]), .B(n979), .Z(c[123]) );
  XNOR U981 ( .A(b[122]), .B(n980), .Z(c[122]) );
  XNOR U982 ( .A(b[121]), .B(n981), .Z(c[121]) );
  XNOR U983 ( .A(b[120]), .B(n982), .Z(c[120]) );
  XNOR U984 ( .A(b[11]), .B(n983), .Z(c[11]) );
  XNOR U985 ( .A(b[119]), .B(n984), .Z(c[119]) );
  XNOR U986 ( .A(b[118]), .B(n985), .Z(c[118]) );
  XNOR U987 ( .A(b[117]), .B(n986), .Z(c[117]) );
  XNOR U988 ( .A(b[116]), .B(n987), .Z(c[116]) );
  XNOR U989 ( .A(b[115]), .B(n988), .Z(c[115]) );
  XNOR U990 ( .A(b[114]), .B(n989), .Z(c[114]) );
  XNOR U991 ( .A(b[113]), .B(n990), .Z(c[113]) );
  XNOR U992 ( .A(b[112]), .B(n991), .Z(c[112]) );
  XNOR U993 ( .A(b[111]), .B(n992), .Z(c[111]) );
  XNOR U994 ( .A(b[110]), .B(n993), .Z(c[110]) );
  XNOR U995 ( .A(b[10]), .B(n994), .Z(c[10]) );
  XNOR U996 ( .A(b[109]), .B(n995), .Z(c[109]) );
  XNOR U997 ( .A(b[108]), .B(n996), .Z(c[108]) );
  XNOR U998 ( .A(b[107]), .B(n997), .Z(c[107]) );
  XNOR U999 ( .A(b[106]), .B(n998), .Z(c[106]) );
  XNOR U1000 ( .A(b[105]), .B(n999), .Z(c[105]) );
  XNOR U1001 ( .A(b[104]), .B(n1000), .Z(c[104]) );
  XNOR U1002 ( .A(b[103]), .B(n1001), .Z(c[103]) );
  XNOR U1003 ( .A(b[102]), .B(n1002), .Z(c[102]) );
  XNOR U1004 ( .A(b[1023]), .B(n5), .Z(c[1023]) );
  XNOR U1005 ( .A(a[1023]), .B(n3), .Z(n5) );
  XNOR U1006 ( .A(n1003), .B(n1004), .Z(n3) );
  ANDN U1007 ( .B(n1005), .A(n1006), .Z(n1003) );
  XNOR U1008 ( .A(b[1022]), .B(n1004), .Z(n1005) );
  XNOR U1009 ( .A(b[1022]), .B(n1006), .Z(c[1022]) );
  XNOR U1010 ( .A(a[1022]), .B(n1007), .Z(n1006) );
  IV U1011 ( .A(n1004), .Z(n1007) );
  XOR U1012 ( .A(n1008), .B(n1009), .Z(n1004) );
  ANDN U1013 ( .B(n1010), .A(n1011), .Z(n1008) );
  XNOR U1014 ( .A(b[1021]), .B(n1009), .Z(n1010) );
  XNOR U1015 ( .A(b[1021]), .B(n1011), .Z(c[1021]) );
  XNOR U1016 ( .A(a[1021]), .B(n1012), .Z(n1011) );
  IV U1017 ( .A(n1009), .Z(n1012) );
  XOR U1018 ( .A(n1013), .B(n1014), .Z(n1009) );
  ANDN U1019 ( .B(n1015), .A(n1016), .Z(n1013) );
  XNOR U1020 ( .A(b[1020]), .B(n1014), .Z(n1015) );
  XNOR U1021 ( .A(b[1020]), .B(n1016), .Z(c[1020]) );
  XNOR U1022 ( .A(a[1020]), .B(n1017), .Z(n1016) );
  IV U1023 ( .A(n1014), .Z(n1017) );
  XOR U1024 ( .A(n1018), .B(n1019), .Z(n1014) );
  ANDN U1025 ( .B(n1020), .A(n1021), .Z(n1018) );
  XNOR U1026 ( .A(b[1019]), .B(n1019), .Z(n1020) );
  XNOR U1027 ( .A(b[101]), .B(n1022), .Z(c[101]) );
  XNOR U1028 ( .A(b[1019]), .B(n1021), .Z(c[1019]) );
  XNOR U1029 ( .A(a[1019]), .B(n1023), .Z(n1021) );
  IV U1030 ( .A(n1019), .Z(n1023) );
  XOR U1031 ( .A(n1024), .B(n1025), .Z(n1019) );
  ANDN U1032 ( .B(n1026), .A(n1027), .Z(n1024) );
  XNOR U1033 ( .A(b[1018]), .B(n1025), .Z(n1026) );
  XNOR U1034 ( .A(b[1018]), .B(n1027), .Z(c[1018]) );
  XNOR U1035 ( .A(a[1018]), .B(n1028), .Z(n1027) );
  IV U1036 ( .A(n1025), .Z(n1028) );
  XOR U1037 ( .A(n1029), .B(n1030), .Z(n1025) );
  ANDN U1038 ( .B(n1031), .A(n1032), .Z(n1029) );
  XNOR U1039 ( .A(b[1017]), .B(n1030), .Z(n1031) );
  XNOR U1040 ( .A(b[1017]), .B(n1032), .Z(c[1017]) );
  XNOR U1041 ( .A(a[1017]), .B(n1033), .Z(n1032) );
  IV U1042 ( .A(n1030), .Z(n1033) );
  XOR U1043 ( .A(n1034), .B(n1035), .Z(n1030) );
  ANDN U1044 ( .B(n1036), .A(n1037), .Z(n1034) );
  XNOR U1045 ( .A(b[1016]), .B(n1035), .Z(n1036) );
  XNOR U1046 ( .A(b[1016]), .B(n1037), .Z(c[1016]) );
  XNOR U1047 ( .A(a[1016]), .B(n1038), .Z(n1037) );
  IV U1048 ( .A(n1035), .Z(n1038) );
  XOR U1049 ( .A(n1039), .B(n1040), .Z(n1035) );
  ANDN U1050 ( .B(n1041), .A(n1042), .Z(n1039) );
  XNOR U1051 ( .A(b[1015]), .B(n1040), .Z(n1041) );
  XNOR U1052 ( .A(b[1015]), .B(n1042), .Z(c[1015]) );
  XNOR U1053 ( .A(a[1015]), .B(n1043), .Z(n1042) );
  IV U1054 ( .A(n1040), .Z(n1043) );
  XOR U1055 ( .A(n1044), .B(n1045), .Z(n1040) );
  ANDN U1056 ( .B(n1046), .A(n1047), .Z(n1044) );
  XNOR U1057 ( .A(b[1014]), .B(n1045), .Z(n1046) );
  XNOR U1058 ( .A(b[1014]), .B(n1047), .Z(c[1014]) );
  XNOR U1059 ( .A(a[1014]), .B(n1048), .Z(n1047) );
  IV U1060 ( .A(n1045), .Z(n1048) );
  XOR U1061 ( .A(n1049), .B(n1050), .Z(n1045) );
  ANDN U1062 ( .B(n1051), .A(n1052), .Z(n1049) );
  XNOR U1063 ( .A(b[1013]), .B(n1050), .Z(n1051) );
  XNOR U1064 ( .A(b[1013]), .B(n1052), .Z(c[1013]) );
  XNOR U1065 ( .A(a[1013]), .B(n1053), .Z(n1052) );
  IV U1066 ( .A(n1050), .Z(n1053) );
  XOR U1067 ( .A(n1054), .B(n1055), .Z(n1050) );
  ANDN U1068 ( .B(n1056), .A(n1057), .Z(n1054) );
  XNOR U1069 ( .A(b[1012]), .B(n1055), .Z(n1056) );
  XNOR U1070 ( .A(b[1012]), .B(n1057), .Z(c[1012]) );
  XNOR U1071 ( .A(a[1012]), .B(n1058), .Z(n1057) );
  IV U1072 ( .A(n1055), .Z(n1058) );
  XOR U1073 ( .A(n1059), .B(n1060), .Z(n1055) );
  ANDN U1074 ( .B(n1061), .A(n1062), .Z(n1059) );
  XNOR U1075 ( .A(b[1011]), .B(n1060), .Z(n1061) );
  XNOR U1076 ( .A(b[1011]), .B(n1062), .Z(c[1011]) );
  XNOR U1077 ( .A(a[1011]), .B(n1063), .Z(n1062) );
  IV U1078 ( .A(n1060), .Z(n1063) );
  XOR U1079 ( .A(n1064), .B(n1065), .Z(n1060) );
  ANDN U1080 ( .B(n1066), .A(n1067), .Z(n1064) );
  XNOR U1081 ( .A(b[1010]), .B(n1065), .Z(n1066) );
  XNOR U1082 ( .A(b[1010]), .B(n1067), .Z(c[1010]) );
  XNOR U1083 ( .A(a[1010]), .B(n1068), .Z(n1067) );
  IV U1084 ( .A(n1065), .Z(n1068) );
  XOR U1085 ( .A(n1069), .B(n1070), .Z(n1065) );
  ANDN U1086 ( .B(n1071), .A(n1072), .Z(n1069) );
  XNOR U1087 ( .A(b[1009]), .B(n1070), .Z(n1071) );
  XNOR U1088 ( .A(b[100]), .B(n1073), .Z(c[100]) );
  XNOR U1089 ( .A(b[1009]), .B(n1072), .Z(c[1009]) );
  XNOR U1090 ( .A(a[1009]), .B(n1074), .Z(n1072) );
  IV U1091 ( .A(n1070), .Z(n1074) );
  XOR U1092 ( .A(n1075), .B(n1076), .Z(n1070) );
  ANDN U1093 ( .B(n1077), .A(n1078), .Z(n1075) );
  XNOR U1094 ( .A(b[1008]), .B(n1076), .Z(n1077) );
  XNOR U1095 ( .A(b[1008]), .B(n1078), .Z(c[1008]) );
  XNOR U1096 ( .A(a[1008]), .B(n1079), .Z(n1078) );
  IV U1097 ( .A(n1076), .Z(n1079) );
  XOR U1098 ( .A(n1080), .B(n1081), .Z(n1076) );
  ANDN U1099 ( .B(n1082), .A(n1083), .Z(n1080) );
  XNOR U1100 ( .A(b[1007]), .B(n1081), .Z(n1082) );
  XNOR U1101 ( .A(b[1007]), .B(n1083), .Z(c[1007]) );
  XNOR U1102 ( .A(a[1007]), .B(n1084), .Z(n1083) );
  IV U1103 ( .A(n1081), .Z(n1084) );
  XOR U1104 ( .A(n1085), .B(n1086), .Z(n1081) );
  ANDN U1105 ( .B(n1087), .A(n1088), .Z(n1085) );
  XNOR U1106 ( .A(b[1006]), .B(n1086), .Z(n1087) );
  XNOR U1107 ( .A(b[1006]), .B(n1088), .Z(c[1006]) );
  XNOR U1108 ( .A(a[1006]), .B(n1089), .Z(n1088) );
  IV U1109 ( .A(n1086), .Z(n1089) );
  XOR U1110 ( .A(n1090), .B(n1091), .Z(n1086) );
  ANDN U1111 ( .B(n1092), .A(n1093), .Z(n1090) );
  XNOR U1112 ( .A(b[1005]), .B(n1091), .Z(n1092) );
  XNOR U1113 ( .A(b[1005]), .B(n1093), .Z(c[1005]) );
  XNOR U1114 ( .A(a[1005]), .B(n1094), .Z(n1093) );
  IV U1115 ( .A(n1091), .Z(n1094) );
  XOR U1116 ( .A(n1095), .B(n1096), .Z(n1091) );
  ANDN U1117 ( .B(n1097), .A(n1098), .Z(n1095) );
  XNOR U1118 ( .A(b[1004]), .B(n1096), .Z(n1097) );
  XNOR U1119 ( .A(b[1004]), .B(n1098), .Z(c[1004]) );
  XNOR U1120 ( .A(a[1004]), .B(n1099), .Z(n1098) );
  IV U1121 ( .A(n1096), .Z(n1099) );
  XOR U1122 ( .A(n1100), .B(n1101), .Z(n1096) );
  ANDN U1123 ( .B(n1102), .A(n1103), .Z(n1100) );
  XNOR U1124 ( .A(b[1003]), .B(n1101), .Z(n1102) );
  XNOR U1125 ( .A(b[1003]), .B(n1103), .Z(c[1003]) );
  XNOR U1126 ( .A(a[1003]), .B(n1104), .Z(n1103) );
  IV U1127 ( .A(n1101), .Z(n1104) );
  XOR U1128 ( .A(n1105), .B(n1106), .Z(n1101) );
  ANDN U1129 ( .B(n1107), .A(n1108), .Z(n1105) );
  XNOR U1130 ( .A(b[1002]), .B(n1106), .Z(n1107) );
  XNOR U1131 ( .A(b[1002]), .B(n1108), .Z(c[1002]) );
  XNOR U1132 ( .A(a[1002]), .B(n1109), .Z(n1108) );
  IV U1133 ( .A(n1106), .Z(n1109) );
  XOR U1134 ( .A(n1110), .B(n1111), .Z(n1106) );
  ANDN U1135 ( .B(n1112), .A(n1113), .Z(n1110) );
  XNOR U1136 ( .A(b[1001]), .B(n1111), .Z(n1112) );
  XNOR U1137 ( .A(b[1001]), .B(n1113), .Z(c[1001]) );
  XNOR U1138 ( .A(a[1001]), .B(n1114), .Z(n1113) );
  IV U1139 ( .A(n1111), .Z(n1114) );
  XOR U1140 ( .A(n1115), .B(n1116), .Z(n1111) );
  ANDN U1141 ( .B(n1117), .A(n1118), .Z(n1115) );
  XNOR U1142 ( .A(b[1000]), .B(n1116), .Z(n1117) );
  XNOR U1143 ( .A(b[1000]), .B(n1118), .Z(c[1000]) );
  XNOR U1144 ( .A(a[1000]), .B(n1119), .Z(n1118) );
  IV U1145 ( .A(n1116), .Z(n1119) );
  XOR U1146 ( .A(n1120), .B(n1121), .Z(n1116) );
  ANDN U1147 ( .B(n1122), .A(n8), .Z(n1120) );
  XNOR U1148 ( .A(a[999]), .B(n1123), .Z(n8) );
  IV U1149 ( .A(n1121), .Z(n1123) );
  XNOR U1150 ( .A(b[999]), .B(n1121), .Z(n1122) );
  XOR U1151 ( .A(n1124), .B(n1125), .Z(n1121) );
  ANDN U1152 ( .B(n1126), .A(n9), .Z(n1124) );
  XNOR U1153 ( .A(a[998]), .B(n1127), .Z(n9) );
  IV U1154 ( .A(n1125), .Z(n1127) );
  XNOR U1155 ( .A(b[998]), .B(n1125), .Z(n1126) );
  XOR U1156 ( .A(n1128), .B(n1129), .Z(n1125) );
  ANDN U1157 ( .B(n1130), .A(n10), .Z(n1128) );
  XNOR U1158 ( .A(a[997]), .B(n1131), .Z(n10) );
  IV U1159 ( .A(n1129), .Z(n1131) );
  XNOR U1160 ( .A(b[997]), .B(n1129), .Z(n1130) );
  XOR U1161 ( .A(n1132), .B(n1133), .Z(n1129) );
  ANDN U1162 ( .B(n1134), .A(n11), .Z(n1132) );
  XNOR U1163 ( .A(a[996]), .B(n1135), .Z(n11) );
  IV U1164 ( .A(n1133), .Z(n1135) );
  XNOR U1165 ( .A(b[996]), .B(n1133), .Z(n1134) );
  XOR U1166 ( .A(n1136), .B(n1137), .Z(n1133) );
  ANDN U1167 ( .B(n1138), .A(n12), .Z(n1136) );
  XNOR U1168 ( .A(a[995]), .B(n1139), .Z(n12) );
  IV U1169 ( .A(n1137), .Z(n1139) );
  XNOR U1170 ( .A(b[995]), .B(n1137), .Z(n1138) );
  XOR U1171 ( .A(n1140), .B(n1141), .Z(n1137) );
  ANDN U1172 ( .B(n1142), .A(n13), .Z(n1140) );
  XNOR U1173 ( .A(a[994]), .B(n1143), .Z(n13) );
  IV U1174 ( .A(n1141), .Z(n1143) );
  XNOR U1175 ( .A(b[994]), .B(n1141), .Z(n1142) );
  XOR U1176 ( .A(n1144), .B(n1145), .Z(n1141) );
  ANDN U1177 ( .B(n1146), .A(n14), .Z(n1144) );
  XNOR U1178 ( .A(a[993]), .B(n1147), .Z(n14) );
  IV U1179 ( .A(n1145), .Z(n1147) );
  XNOR U1180 ( .A(b[993]), .B(n1145), .Z(n1146) );
  XOR U1181 ( .A(n1148), .B(n1149), .Z(n1145) );
  ANDN U1182 ( .B(n1150), .A(n15), .Z(n1148) );
  XNOR U1183 ( .A(a[992]), .B(n1151), .Z(n15) );
  IV U1184 ( .A(n1149), .Z(n1151) );
  XNOR U1185 ( .A(b[992]), .B(n1149), .Z(n1150) );
  XOR U1186 ( .A(n1152), .B(n1153), .Z(n1149) );
  ANDN U1187 ( .B(n1154), .A(n16), .Z(n1152) );
  XNOR U1188 ( .A(a[991]), .B(n1155), .Z(n16) );
  IV U1189 ( .A(n1153), .Z(n1155) );
  XNOR U1190 ( .A(b[991]), .B(n1153), .Z(n1154) );
  XOR U1191 ( .A(n1156), .B(n1157), .Z(n1153) );
  ANDN U1192 ( .B(n1158), .A(n17), .Z(n1156) );
  XNOR U1193 ( .A(a[990]), .B(n1159), .Z(n17) );
  IV U1194 ( .A(n1157), .Z(n1159) );
  XNOR U1195 ( .A(b[990]), .B(n1157), .Z(n1158) );
  XOR U1196 ( .A(n1160), .B(n1161), .Z(n1157) );
  ANDN U1197 ( .B(n1162), .A(n19), .Z(n1160) );
  XNOR U1198 ( .A(a[989]), .B(n1163), .Z(n19) );
  IV U1199 ( .A(n1161), .Z(n1163) );
  XNOR U1200 ( .A(b[989]), .B(n1161), .Z(n1162) );
  XOR U1201 ( .A(n1164), .B(n1165), .Z(n1161) );
  ANDN U1202 ( .B(n1166), .A(n20), .Z(n1164) );
  XNOR U1203 ( .A(a[988]), .B(n1167), .Z(n20) );
  IV U1204 ( .A(n1165), .Z(n1167) );
  XNOR U1205 ( .A(b[988]), .B(n1165), .Z(n1166) );
  XOR U1206 ( .A(n1168), .B(n1169), .Z(n1165) );
  ANDN U1207 ( .B(n1170), .A(n21), .Z(n1168) );
  XNOR U1208 ( .A(a[987]), .B(n1171), .Z(n21) );
  IV U1209 ( .A(n1169), .Z(n1171) );
  XNOR U1210 ( .A(b[987]), .B(n1169), .Z(n1170) );
  XOR U1211 ( .A(n1172), .B(n1173), .Z(n1169) );
  ANDN U1212 ( .B(n1174), .A(n22), .Z(n1172) );
  XNOR U1213 ( .A(a[986]), .B(n1175), .Z(n22) );
  IV U1214 ( .A(n1173), .Z(n1175) );
  XNOR U1215 ( .A(b[986]), .B(n1173), .Z(n1174) );
  XOR U1216 ( .A(n1176), .B(n1177), .Z(n1173) );
  ANDN U1217 ( .B(n1178), .A(n23), .Z(n1176) );
  XNOR U1218 ( .A(a[985]), .B(n1179), .Z(n23) );
  IV U1219 ( .A(n1177), .Z(n1179) );
  XNOR U1220 ( .A(b[985]), .B(n1177), .Z(n1178) );
  XOR U1221 ( .A(n1180), .B(n1181), .Z(n1177) );
  ANDN U1222 ( .B(n1182), .A(n24), .Z(n1180) );
  XNOR U1223 ( .A(a[984]), .B(n1183), .Z(n24) );
  IV U1224 ( .A(n1181), .Z(n1183) );
  XNOR U1225 ( .A(b[984]), .B(n1181), .Z(n1182) );
  XOR U1226 ( .A(n1184), .B(n1185), .Z(n1181) );
  ANDN U1227 ( .B(n1186), .A(n25), .Z(n1184) );
  XNOR U1228 ( .A(a[983]), .B(n1187), .Z(n25) );
  IV U1229 ( .A(n1185), .Z(n1187) );
  XNOR U1230 ( .A(b[983]), .B(n1185), .Z(n1186) );
  XOR U1231 ( .A(n1188), .B(n1189), .Z(n1185) );
  ANDN U1232 ( .B(n1190), .A(n26), .Z(n1188) );
  XNOR U1233 ( .A(a[982]), .B(n1191), .Z(n26) );
  IV U1234 ( .A(n1189), .Z(n1191) );
  XNOR U1235 ( .A(b[982]), .B(n1189), .Z(n1190) );
  XOR U1236 ( .A(n1192), .B(n1193), .Z(n1189) );
  ANDN U1237 ( .B(n1194), .A(n27), .Z(n1192) );
  XNOR U1238 ( .A(a[981]), .B(n1195), .Z(n27) );
  IV U1239 ( .A(n1193), .Z(n1195) );
  XNOR U1240 ( .A(b[981]), .B(n1193), .Z(n1194) );
  XOR U1241 ( .A(n1196), .B(n1197), .Z(n1193) );
  ANDN U1242 ( .B(n1198), .A(n28), .Z(n1196) );
  XNOR U1243 ( .A(a[980]), .B(n1199), .Z(n28) );
  IV U1244 ( .A(n1197), .Z(n1199) );
  XNOR U1245 ( .A(b[980]), .B(n1197), .Z(n1198) );
  XOR U1246 ( .A(n1200), .B(n1201), .Z(n1197) );
  ANDN U1247 ( .B(n1202), .A(n30), .Z(n1200) );
  XNOR U1248 ( .A(a[979]), .B(n1203), .Z(n30) );
  IV U1249 ( .A(n1201), .Z(n1203) );
  XNOR U1250 ( .A(b[979]), .B(n1201), .Z(n1202) );
  XOR U1251 ( .A(n1204), .B(n1205), .Z(n1201) );
  ANDN U1252 ( .B(n1206), .A(n31), .Z(n1204) );
  XNOR U1253 ( .A(a[978]), .B(n1207), .Z(n31) );
  IV U1254 ( .A(n1205), .Z(n1207) );
  XNOR U1255 ( .A(b[978]), .B(n1205), .Z(n1206) );
  XOR U1256 ( .A(n1208), .B(n1209), .Z(n1205) );
  ANDN U1257 ( .B(n1210), .A(n32), .Z(n1208) );
  XNOR U1258 ( .A(a[977]), .B(n1211), .Z(n32) );
  IV U1259 ( .A(n1209), .Z(n1211) );
  XNOR U1260 ( .A(b[977]), .B(n1209), .Z(n1210) );
  XOR U1261 ( .A(n1212), .B(n1213), .Z(n1209) );
  ANDN U1262 ( .B(n1214), .A(n33), .Z(n1212) );
  XNOR U1263 ( .A(a[976]), .B(n1215), .Z(n33) );
  IV U1264 ( .A(n1213), .Z(n1215) );
  XNOR U1265 ( .A(b[976]), .B(n1213), .Z(n1214) );
  XOR U1266 ( .A(n1216), .B(n1217), .Z(n1213) );
  ANDN U1267 ( .B(n1218), .A(n34), .Z(n1216) );
  XNOR U1268 ( .A(a[975]), .B(n1219), .Z(n34) );
  IV U1269 ( .A(n1217), .Z(n1219) );
  XNOR U1270 ( .A(b[975]), .B(n1217), .Z(n1218) );
  XOR U1271 ( .A(n1220), .B(n1221), .Z(n1217) );
  ANDN U1272 ( .B(n1222), .A(n35), .Z(n1220) );
  XNOR U1273 ( .A(a[974]), .B(n1223), .Z(n35) );
  IV U1274 ( .A(n1221), .Z(n1223) );
  XNOR U1275 ( .A(b[974]), .B(n1221), .Z(n1222) );
  XOR U1276 ( .A(n1224), .B(n1225), .Z(n1221) );
  ANDN U1277 ( .B(n1226), .A(n36), .Z(n1224) );
  XNOR U1278 ( .A(a[973]), .B(n1227), .Z(n36) );
  IV U1279 ( .A(n1225), .Z(n1227) );
  XNOR U1280 ( .A(b[973]), .B(n1225), .Z(n1226) );
  XOR U1281 ( .A(n1228), .B(n1229), .Z(n1225) );
  ANDN U1282 ( .B(n1230), .A(n37), .Z(n1228) );
  XNOR U1283 ( .A(a[972]), .B(n1231), .Z(n37) );
  IV U1284 ( .A(n1229), .Z(n1231) );
  XNOR U1285 ( .A(b[972]), .B(n1229), .Z(n1230) );
  XOR U1286 ( .A(n1232), .B(n1233), .Z(n1229) );
  ANDN U1287 ( .B(n1234), .A(n38), .Z(n1232) );
  XNOR U1288 ( .A(a[971]), .B(n1235), .Z(n38) );
  IV U1289 ( .A(n1233), .Z(n1235) );
  XNOR U1290 ( .A(b[971]), .B(n1233), .Z(n1234) );
  XOR U1291 ( .A(n1236), .B(n1237), .Z(n1233) );
  ANDN U1292 ( .B(n1238), .A(n39), .Z(n1236) );
  XNOR U1293 ( .A(a[970]), .B(n1239), .Z(n39) );
  IV U1294 ( .A(n1237), .Z(n1239) );
  XNOR U1295 ( .A(b[970]), .B(n1237), .Z(n1238) );
  XOR U1296 ( .A(n1240), .B(n1241), .Z(n1237) );
  ANDN U1297 ( .B(n1242), .A(n41), .Z(n1240) );
  XNOR U1298 ( .A(a[969]), .B(n1243), .Z(n41) );
  IV U1299 ( .A(n1241), .Z(n1243) );
  XNOR U1300 ( .A(b[969]), .B(n1241), .Z(n1242) );
  XOR U1301 ( .A(n1244), .B(n1245), .Z(n1241) );
  ANDN U1302 ( .B(n1246), .A(n42), .Z(n1244) );
  XNOR U1303 ( .A(a[968]), .B(n1247), .Z(n42) );
  IV U1304 ( .A(n1245), .Z(n1247) );
  XNOR U1305 ( .A(b[968]), .B(n1245), .Z(n1246) );
  XOR U1306 ( .A(n1248), .B(n1249), .Z(n1245) );
  ANDN U1307 ( .B(n1250), .A(n43), .Z(n1248) );
  XNOR U1308 ( .A(a[967]), .B(n1251), .Z(n43) );
  IV U1309 ( .A(n1249), .Z(n1251) );
  XNOR U1310 ( .A(b[967]), .B(n1249), .Z(n1250) );
  XOR U1311 ( .A(n1252), .B(n1253), .Z(n1249) );
  ANDN U1312 ( .B(n1254), .A(n44), .Z(n1252) );
  XNOR U1313 ( .A(a[966]), .B(n1255), .Z(n44) );
  IV U1314 ( .A(n1253), .Z(n1255) );
  XNOR U1315 ( .A(b[966]), .B(n1253), .Z(n1254) );
  XOR U1316 ( .A(n1256), .B(n1257), .Z(n1253) );
  ANDN U1317 ( .B(n1258), .A(n45), .Z(n1256) );
  XNOR U1318 ( .A(a[965]), .B(n1259), .Z(n45) );
  IV U1319 ( .A(n1257), .Z(n1259) );
  XNOR U1320 ( .A(b[965]), .B(n1257), .Z(n1258) );
  XOR U1321 ( .A(n1260), .B(n1261), .Z(n1257) );
  ANDN U1322 ( .B(n1262), .A(n46), .Z(n1260) );
  XNOR U1323 ( .A(a[964]), .B(n1263), .Z(n46) );
  IV U1324 ( .A(n1261), .Z(n1263) );
  XNOR U1325 ( .A(b[964]), .B(n1261), .Z(n1262) );
  XOR U1326 ( .A(n1264), .B(n1265), .Z(n1261) );
  ANDN U1327 ( .B(n1266), .A(n47), .Z(n1264) );
  XNOR U1328 ( .A(a[963]), .B(n1267), .Z(n47) );
  IV U1329 ( .A(n1265), .Z(n1267) );
  XNOR U1330 ( .A(b[963]), .B(n1265), .Z(n1266) );
  XOR U1331 ( .A(n1268), .B(n1269), .Z(n1265) );
  ANDN U1332 ( .B(n1270), .A(n48), .Z(n1268) );
  XNOR U1333 ( .A(a[962]), .B(n1271), .Z(n48) );
  IV U1334 ( .A(n1269), .Z(n1271) );
  XNOR U1335 ( .A(b[962]), .B(n1269), .Z(n1270) );
  XOR U1336 ( .A(n1272), .B(n1273), .Z(n1269) );
  ANDN U1337 ( .B(n1274), .A(n49), .Z(n1272) );
  XNOR U1338 ( .A(a[961]), .B(n1275), .Z(n49) );
  IV U1339 ( .A(n1273), .Z(n1275) );
  XNOR U1340 ( .A(b[961]), .B(n1273), .Z(n1274) );
  XOR U1341 ( .A(n1276), .B(n1277), .Z(n1273) );
  ANDN U1342 ( .B(n1278), .A(n50), .Z(n1276) );
  XNOR U1343 ( .A(a[960]), .B(n1279), .Z(n50) );
  IV U1344 ( .A(n1277), .Z(n1279) );
  XNOR U1345 ( .A(b[960]), .B(n1277), .Z(n1278) );
  XOR U1346 ( .A(n1280), .B(n1281), .Z(n1277) );
  ANDN U1347 ( .B(n1282), .A(n52), .Z(n1280) );
  XNOR U1348 ( .A(a[959]), .B(n1283), .Z(n52) );
  IV U1349 ( .A(n1281), .Z(n1283) );
  XNOR U1350 ( .A(b[959]), .B(n1281), .Z(n1282) );
  XOR U1351 ( .A(n1284), .B(n1285), .Z(n1281) );
  ANDN U1352 ( .B(n1286), .A(n53), .Z(n1284) );
  XNOR U1353 ( .A(a[958]), .B(n1287), .Z(n53) );
  IV U1354 ( .A(n1285), .Z(n1287) );
  XNOR U1355 ( .A(b[958]), .B(n1285), .Z(n1286) );
  XOR U1356 ( .A(n1288), .B(n1289), .Z(n1285) );
  ANDN U1357 ( .B(n1290), .A(n54), .Z(n1288) );
  XNOR U1358 ( .A(a[957]), .B(n1291), .Z(n54) );
  IV U1359 ( .A(n1289), .Z(n1291) );
  XNOR U1360 ( .A(b[957]), .B(n1289), .Z(n1290) );
  XOR U1361 ( .A(n1292), .B(n1293), .Z(n1289) );
  ANDN U1362 ( .B(n1294), .A(n55), .Z(n1292) );
  XNOR U1363 ( .A(a[956]), .B(n1295), .Z(n55) );
  IV U1364 ( .A(n1293), .Z(n1295) );
  XNOR U1365 ( .A(b[956]), .B(n1293), .Z(n1294) );
  XOR U1366 ( .A(n1296), .B(n1297), .Z(n1293) );
  ANDN U1367 ( .B(n1298), .A(n56), .Z(n1296) );
  XNOR U1368 ( .A(a[955]), .B(n1299), .Z(n56) );
  IV U1369 ( .A(n1297), .Z(n1299) );
  XNOR U1370 ( .A(b[955]), .B(n1297), .Z(n1298) );
  XOR U1371 ( .A(n1300), .B(n1301), .Z(n1297) );
  ANDN U1372 ( .B(n1302), .A(n57), .Z(n1300) );
  XNOR U1373 ( .A(a[954]), .B(n1303), .Z(n57) );
  IV U1374 ( .A(n1301), .Z(n1303) );
  XNOR U1375 ( .A(b[954]), .B(n1301), .Z(n1302) );
  XOR U1376 ( .A(n1304), .B(n1305), .Z(n1301) );
  ANDN U1377 ( .B(n1306), .A(n58), .Z(n1304) );
  XNOR U1378 ( .A(a[953]), .B(n1307), .Z(n58) );
  IV U1379 ( .A(n1305), .Z(n1307) );
  XNOR U1380 ( .A(b[953]), .B(n1305), .Z(n1306) );
  XOR U1381 ( .A(n1308), .B(n1309), .Z(n1305) );
  ANDN U1382 ( .B(n1310), .A(n59), .Z(n1308) );
  XNOR U1383 ( .A(a[952]), .B(n1311), .Z(n59) );
  IV U1384 ( .A(n1309), .Z(n1311) );
  XNOR U1385 ( .A(b[952]), .B(n1309), .Z(n1310) );
  XOR U1386 ( .A(n1312), .B(n1313), .Z(n1309) );
  ANDN U1387 ( .B(n1314), .A(n60), .Z(n1312) );
  XNOR U1388 ( .A(a[951]), .B(n1315), .Z(n60) );
  IV U1389 ( .A(n1313), .Z(n1315) );
  XNOR U1390 ( .A(b[951]), .B(n1313), .Z(n1314) );
  XOR U1391 ( .A(n1316), .B(n1317), .Z(n1313) );
  ANDN U1392 ( .B(n1318), .A(n61), .Z(n1316) );
  XNOR U1393 ( .A(a[950]), .B(n1319), .Z(n61) );
  IV U1394 ( .A(n1317), .Z(n1319) );
  XNOR U1395 ( .A(b[950]), .B(n1317), .Z(n1318) );
  XOR U1396 ( .A(n1320), .B(n1321), .Z(n1317) );
  ANDN U1397 ( .B(n1322), .A(n63), .Z(n1320) );
  XNOR U1398 ( .A(a[949]), .B(n1323), .Z(n63) );
  IV U1399 ( .A(n1321), .Z(n1323) );
  XNOR U1400 ( .A(b[949]), .B(n1321), .Z(n1322) );
  XOR U1401 ( .A(n1324), .B(n1325), .Z(n1321) );
  ANDN U1402 ( .B(n1326), .A(n64), .Z(n1324) );
  XNOR U1403 ( .A(a[948]), .B(n1327), .Z(n64) );
  IV U1404 ( .A(n1325), .Z(n1327) );
  XNOR U1405 ( .A(b[948]), .B(n1325), .Z(n1326) );
  XOR U1406 ( .A(n1328), .B(n1329), .Z(n1325) );
  ANDN U1407 ( .B(n1330), .A(n65), .Z(n1328) );
  XNOR U1408 ( .A(a[947]), .B(n1331), .Z(n65) );
  IV U1409 ( .A(n1329), .Z(n1331) );
  XNOR U1410 ( .A(b[947]), .B(n1329), .Z(n1330) );
  XOR U1411 ( .A(n1332), .B(n1333), .Z(n1329) );
  ANDN U1412 ( .B(n1334), .A(n66), .Z(n1332) );
  XNOR U1413 ( .A(a[946]), .B(n1335), .Z(n66) );
  IV U1414 ( .A(n1333), .Z(n1335) );
  XNOR U1415 ( .A(b[946]), .B(n1333), .Z(n1334) );
  XOR U1416 ( .A(n1336), .B(n1337), .Z(n1333) );
  ANDN U1417 ( .B(n1338), .A(n67), .Z(n1336) );
  XNOR U1418 ( .A(a[945]), .B(n1339), .Z(n67) );
  IV U1419 ( .A(n1337), .Z(n1339) );
  XNOR U1420 ( .A(b[945]), .B(n1337), .Z(n1338) );
  XOR U1421 ( .A(n1340), .B(n1341), .Z(n1337) );
  ANDN U1422 ( .B(n1342), .A(n68), .Z(n1340) );
  XNOR U1423 ( .A(a[944]), .B(n1343), .Z(n68) );
  IV U1424 ( .A(n1341), .Z(n1343) );
  XNOR U1425 ( .A(b[944]), .B(n1341), .Z(n1342) );
  XOR U1426 ( .A(n1344), .B(n1345), .Z(n1341) );
  ANDN U1427 ( .B(n1346), .A(n69), .Z(n1344) );
  XNOR U1428 ( .A(a[943]), .B(n1347), .Z(n69) );
  IV U1429 ( .A(n1345), .Z(n1347) );
  XNOR U1430 ( .A(b[943]), .B(n1345), .Z(n1346) );
  XOR U1431 ( .A(n1348), .B(n1349), .Z(n1345) );
  ANDN U1432 ( .B(n1350), .A(n70), .Z(n1348) );
  XNOR U1433 ( .A(a[942]), .B(n1351), .Z(n70) );
  IV U1434 ( .A(n1349), .Z(n1351) );
  XNOR U1435 ( .A(b[942]), .B(n1349), .Z(n1350) );
  XOR U1436 ( .A(n1352), .B(n1353), .Z(n1349) );
  ANDN U1437 ( .B(n1354), .A(n71), .Z(n1352) );
  XNOR U1438 ( .A(a[941]), .B(n1355), .Z(n71) );
  IV U1439 ( .A(n1353), .Z(n1355) );
  XNOR U1440 ( .A(b[941]), .B(n1353), .Z(n1354) );
  XOR U1441 ( .A(n1356), .B(n1357), .Z(n1353) );
  ANDN U1442 ( .B(n1358), .A(n72), .Z(n1356) );
  XNOR U1443 ( .A(a[940]), .B(n1359), .Z(n72) );
  IV U1444 ( .A(n1357), .Z(n1359) );
  XNOR U1445 ( .A(b[940]), .B(n1357), .Z(n1358) );
  XOR U1446 ( .A(n1360), .B(n1361), .Z(n1357) );
  ANDN U1447 ( .B(n1362), .A(n74), .Z(n1360) );
  XNOR U1448 ( .A(a[939]), .B(n1363), .Z(n74) );
  IV U1449 ( .A(n1361), .Z(n1363) );
  XNOR U1450 ( .A(b[939]), .B(n1361), .Z(n1362) );
  XOR U1451 ( .A(n1364), .B(n1365), .Z(n1361) );
  ANDN U1452 ( .B(n1366), .A(n75), .Z(n1364) );
  XNOR U1453 ( .A(a[938]), .B(n1367), .Z(n75) );
  IV U1454 ( .A(n1365), .Z(n1367) );
  XNOR U1455 ( .A(b[938]), .B(n1365), .Z(n1366) );
  XOR U1456 ( .A(n1368), .B(n1369), .Z(n1365) );
  ANDN U1457 ( .B(n1370), .A(n76), .Z(n1368) );
  XNOR U1458 ( .A(a[937]), .B(n1371), .Z(n76) );
  IV U1459 ( .A(n1369), .Z(n1371) );
  XNOR U1460 ( .A(b[937]), .B(n1369), .Z(n1370) );
  XOR U1461 ( .A(n1372), .B(n1373), .Z(n1369) );
  ANDN U1462 ( .B(n1374), .A(n77), .Z(n1372) );
  XNOR U1463 ( .A(a[936]), .B(n1375), .Z(n77) );
  IV U1464 ( .A(n1373), .Z(n1375) );
  XNOR U1465 ( .A(b[936]), .B(n1373), .Z(n1374) );
  XOR U1466 ( .A(n1376), .B(n1377), .Z(n1373) );
  ANDN U1467 ( .B(n1378), .A(n78), .Z(n1376) );
  XNOR U1468 ( .A(a[935]), .B(n1379), .Z(n78) );
  IV U1469 ( .A(n1377), .Z(n1379) );
  XNOR U1470 ( .A(b[935]), .B(n1377), .Z(n1378) );
  XOR U1471 ( .A(n1380), .B(n1381), .Z(n1377) );
  ANDN U1472 ( .B(n1382), .A(n79), .Z(n1380) );
  XNOR U1473 ( .A(a[934]), .B(n1383), .Z(n79) );
  IV U1474 ( .A(n1381), .Z(n1383) );
  XNOR U1475 ( .A(b[934]), .B(n1381), .Z(n1382) );
  XOR U1476 ( .A(n1384), .B(n1385), .Z(n1381) );
  ANDN U1477 ( .B(n1386), .A(n80), .Z(n1384) );
  XNOR U1478 ( .A(a[933]), .B(n1387), .Z(n80) );
  IV U1479 ( .A(n1385), .Z(n1387) );
  XNOR U1480 ( .A(b[933]), .B(n1385), .Z(n1386) );
  XOR U1481 ( .A(n1388), .B(n1389), .Z(n1385) );
  ANDN U1482 ( .B(n1390), .A(n81), .Z(n1388) );
  XNOR U1483 ( .A(a[932]), .B(n1391), .Z(n81) );
  IV U1484 ( .A(n1389), .Z(n1391) );
  XNOR U1485 ( .A(b[932]), .B(n1389), .Z(n1390) );
  XOR U1486 ( .A(n1392), .B(n1393), .Z(n1389) );
  ANDN U1487 ( .B(n1394), .A(n82), .Z(n1392) );
  XNOR U1488 ( .A(a[931]), .B(n1395), .Z(n82) );
  IV U1489 ( .A(n1393), .Z(n1395) );
  XNOR U1490 ( .A(b[931]), .B(n1393), .Z(n1394) );
  XOR U1491 ( .A(n1396), .B(n1397), .Z(n1393) );
  ANDN U1492 ( .B(n1398), .A(n83), .Z(n1396) );
  XNOR U1493 ( .A(a[930]), .B(n1399), .Z(n83) );
  IV U1494 ( .A(n1397), .Z(n1399) );
  XNOR U1495 ( .A(b[930]), .B(n1397), .Z(n1398) );
  XOR U1496 ( .A(n1400), .B(n1401), .Z(n1397) );
  ANDN U1497 ( .B(n1402), .A(n85), .Z(n1400) );
  XNOR U1498 ( .A(a[929]), .B(n1403), .Z(n85) );
  IV U1499 ( .A(n1401), .Z(n1403) );
  XNOR U1500 ( .A(b[929]), .B(n1401), .Z(n1402) );
  XOR U1501 ( .A(n1404), .B(n1405), .Z(n1401) );
  ANDN U1502 ( .B(n1406), .A(n86), .Z(n1404) );
  XNOR U1503 ( .A(a[928]), .B(n1407), .Z(n86) );
  IV U1504 ( .A(n1405), .Z(n1407) );
  XNOR U1505 ( .A(b[928]), .B(n1405), .Z(n1406) );
  XOR U1506 ( .A(n1408), .B(n1409), .Z(n1405) );
  ANDN U1507 ( .B(n1410), .A(n87), .Z(n1408) );
  XNOR U1508 ( .A(a[927]), .B(n1411), .Z(n87) );
  IV U1509 ( .A(n1409), .Z(n1411) );
  XNOR U1510 ( .A(b[927]), .B(n1409), .Z(n1410) );
  XOR U1511 ( .A(n1412), .B(n1413), .Z(n1409) );
  ANDN U1512 ( .B(n1414), .A(n88), .Z(n1412) );
  XNOR U1513 ( .A(a[926]), .B(n1415), .Z(n88) );
  IV U1514 ( .A(n1413), .Z(n1415) );
  XNOR U1515 ( .A(b[926]), .B(n1413), .Z(n1414) );
  XOR U1516 ( .A(n1416), .B(n1417), .Z(n1413) );
  ANDN U1517 ( .B(n1418), .A(n89), .Z(n1416) );
  XNOR U1518 ( .A(a[925]), .B(n1419), .Z(n89) );
  IV U1519 ( .A(n1417), .Z(n1419) );
  XNOR U1520 ( .A(b[925]), .B(n1417), .Z(n1418) );
  XOR U1521 ( .A(n1420), .B(n1421), .Z(n1417) );
  ANDN U1522 ( .B(n1422), .A(n90), .Z(n1420) );
  XNOR U1523 ( .A(a[924]), .B(n1423), .Z(n90) );
  IV U1524 ( .A(n1421), .Z(n1423) );
  XNOR U1525 ( .A(b[924]), .B(n1421), .Z(n1422) );
  XOR U1526 ( .A(n1424), .B(n1425), .Z(n1421) );
  ANDN U1527 ( .B(n1426), .A(n91), .Z(n1424) );
  XNOR U1528 ( .A(a[923]), .B(n1427), .Z(n91) );
  IV U1529 ( .A(n1425), .Z(n1427) );
  XNOR U1530 ( .A(b[923]), .B(n1425), .Z(n1426) );
  XOR U1531 ( .A(n1428), .B(n1429), .Z(n1425) );
  ANDN U1532 ( .B(n1430), .A(n92), .Z(n1428) );
  XNOR U1533 ( .A(a[922]), .B(n1431), .Z(n92) );
  IV U1534 ( .A(n1429), .Z(n1431) );
  XNOR U1535 ( .A(b[922]), .B(n1429), .Z(n1430) );
  XOR U1536 ( .A(n1432), .B(n1433), .Z(n1429) );
  ANDN U1537 ( .B(n1434), .A(n93), .Z(n1432) );
  XNOR U1538 ( .A(a[921]), .B(n1435), .Z(n93) );
  IV U1539 ( .A(n1433), .Z(n1435) );
  XNOR U1540 ( .A(b[921]), .B(n1433), .Z(n1434) );
  XOR U1541 ( .A(n1436), .B(n1437), .Z(n1433) );
  ANDN U1542 ( .B(n1438), .A(n94), .Z(n1436) );
  XNOR U1543 ( .A(a[920]), .B(n1439), .Z(n94) );
  IV U1544 ( .A(n1437), .Z(n1439) );
  XNOR U1545 ( .A(b[920]), .B(n1437), .Z(n1438) );
  XOR U1546 ( .A(n1440), .B(n1441), .Z(n1437) );
  ANDN U1547 ( .B(n1442), .A(n96), .Z(n1440) );
  XNOR U1548 ( .A(a[919]), .B(n1443), .Z(n96) );
  IV U1549 ( .A(n1441), .Z(n1443) );
  XNOR U1550 ( .A(b[919]), .B(n1441), .Z(n1442) );
  XOR U1551 ( .A(n1444), .B(n1445), .Z(n1441) );
  ANDN U1552 ( .B(n1446), .A(n97), .Z(n1444) );
  XNOR U1553 ( .A(a[918]), .B(n1447), .Z(n97) );
  IV U1554 ( .A(n1445), .Z(n1447) );
  XNOR U1555 ( .A(b[918]), .B(n1445), .Z(n1446) );
  XOR U1556 ( .A(n1448), .B(n1449), .Z(n1445) );
  ANDN U1557 ( .B(n1450), .A(n98), .Z(n1448) );
  XNOR U1558 ( .A(a[917]), .B(n1451), .Z(n98) );
  IV U1559 ( .A(n1449), .Z(n1451) );
  XNOR U1560 ( .A(b[917]), .B(n1449), .Z(n1450) );
  XOR U1561 ( .A(n1452), .B(n1453), .Z(n1449) );
  ANDN U1562 ( .B(n1454), .A(n99), .Z(n1452) );
  XNOR U1563 ( .A(a[916]), .B(n1455), .Z(n99) );
  IV U1564 ( .A(n1453), .Z(n1455) );
  XNOR U1565 ( .A(b[916]), .B(n1453), .Z(n1454) );
  XOR U1566 ( .A(n1456), .B(n1457), .Z(n1453) );
  ANDN U1567 ( .B(n1458), .A(n100), .Z(n1456) );
  XNOR U1568 ( .A(a[915]), .B(n1459), .Z(n100) );
  IV U1569 ( .A(n1457), .Z(n1459) );
  XNOR U1570 ( .A(b[915]), .B(n1457), .Z(n1458) );
  XOR U1571 ( .A(n1460), .B(n1461), .Z(n1457) );
  ANDN U1572 ( .B(n1462), .A(n101), .Z(n1460) );
  XNOR U1573 ( .A(a[914]), .B(n1463), .Z(n101) );
  IV U1574 ( .A(n1461), .Z(n1463) );
  XNOR U1575 ( .A(b[914]), .B(n1461), .Z(n1462) );
  XOR U1576 ( .A(n1464), .B(n1465), .Z(n1461) );
  ANDN U1577 ( .B(n1466), .A(n102), .Z(n1464) );
  XNOR U1578 ( .A(a[913]), .B(n1467), .Z(n102) );
  IV U1579 ( .A(n1465), .Z(n1467) );
  XNOR U1580 ( .A(b[913]), .B(n1465), .Z(n1466) );
  XOR U1581 ( .A(n1468), .B(n1469), .Z(n1465) );
  ANDN U1582 ( .B(n1470), .A(n103), .Z(n1468) );
  XNOR U1583 ( .A(a[912]), .B(n1471), .Z(n103) );
  IV U1584 ( .A(n1469), .Z(n1471) );
  XNOR U1585 ( .A(b[912]), .B(n1469), .Z(n1470) );
  XOR U1586 ( .A(n1472), .B(n1473), .Z(n1469) );
  ANDN U1587 ( .B(n1474), .A(n104), .Z(n1472) );
  XNOR U1588 ( .A(a[911]), .B(n1475), .Z(n104) );
  IV U1589 ( .A(n1473), .Z(n1475) );
  XNOR U1590 ( .A(b[911]), .B(n1473), .Z(n1474) );
  XOR U1591 ( .A(n1476), .B(n1477), .Z(n1473) );
  ANDN U1592 ( .B(n1478), .A(n105), .Z(n1476) );
  XNOR U1593 ( .A(a[910]), .B(n1479), .Z(n105) );
  IV U1594 ( .A(n1477), .Z(n1479) );
  XNOR U1595 ( .A(b[910]), .B(n1477), .Z(n1478) );
  XOR U1596 ( .A(n1480), .B(n1481), .Z(n1477) );
  ANDN U1597 ( .B(n1482), .A(n107), .Z(n1480) );
  XNOR U1598 ( .A(a[909]), .B(n1483), .Z(n107) );
  IV U1599 ( .A(n1481), .Z(n1483) );
  XNOR U1600 ( .A(b[909]), .B(n1481), .Z(n1482) );
  XOR U1601 ( .A(n1484), .B(n1485), .Z(n1481) );
  ANDN U1602 ( .B(n1486), .A(n108), .Z(n1484) );
  XNOR U1603 ( .A(a[908]), .B(n1487), .Z(n108) );
  IV U1604 ( .A(n1485), .Z(n1487) );
  XNOR U1605 ( .A(b[908]), .B(n1485), .Z(n1486) );
  XOR U1606 ( .A(n1488), .B(n1489), .Z(n1485) );
  ANDN U1607 ( .B(n1490), .A(n109), .Z(n1488) );
  XNOR U1608 ( .A(a[907]), .B(n1491), .Z(n109) );
  IV U1609 ( .A(n1489), .Z(n1491) );
  XNOR U1610 ( .A(b[907]), .B(n1489), .Z(n1490) );
  XOR U1611 ( .A(n1492), .B(n1493), .Z(n1489) );
  ANDN U1612 ( .B(n1494), .A(n110), .Z(n1492) );
  XNOR U1613 ( .A(a[906]), .B(n1495), .Z(n110) );
  IV U1614 ( .A(n1493), .Z(n1495) );
  XNOR U1615 ( .A(b[906]), .B(n1493), .Z(n1494) );
  XOR U1616 ( .A(n1496), .B(n1497), .Z(n1493) );
  ANDN U1617 ( .B(n1498), .A(n111), .Z(n1496) );
  XNOR U1618 ( .A(a[905]), .B(n1499), .Z(n111) );
  IV U1619 ( .A(n1497), .Z(n1499) );
  XNOR U1620 ( .A(b[905]), .B(n1497), .Z(n1498) );
  XOR U1621 ( .A(n1500), .B(n1501), .Z(n1497) );
  ANDN U1622 ( .B(n1502), .A(n112), .Z(n1500) );
  XNOR U1623 ( .A(a[904]), .B(n1503), .Z(n112) );
  IV U1624 ( .A(n1501), .Z(n1503) );
  XNOR U1625 ( .A(b[904]), .B(n1501), .Z(n1502) );
  XOR U1626 ( .A(n1504), .B(n1505), .Z(n1501) );
  ANDN U1627 ( .B(n1506), .A(n113), .Z(n1504) );
  XNOR U1628 ( .A(a[903]), .B(n1507), .Z(n113) );
  IV U1629 ( .A(n1505), .Z(n1507) );
  XNOR U1630 ( .A(b[903]), .B(n1505), .Z(n1506) );
  XOR U1631 ( .A(n1508), .B(n1509), .Z(n1505) );
  ANDN U1632 ( .B(n1510), .A(n114), .Z(n1508) );
  XNOR U1633 ( .A(a[902]), .B(n1511), .Z(n114) );
  IV U1634 ( .A(n1509), .Z(n1511) );
  XNOR U1635 ( .A(b[902]), .B(n1509), .Z(n1510) );
  XOR U1636 ( .A(n1512), .B(n1513), .Z(n1509) );
  ANDN U1637 ( .B(n1514), .A(n115), .Z(n1512) );
  XNOR U1638 ( .A(a[901]), .B(n1515), .Z(n115) );
  IV U1639 ( .A(n1513), .Z(n1515) );
  XNOR U1640 ( .A(b[901]), .B(n1513), .Z(n1514) );
  XOR U1641 ( .A(n1516), .B(n1517), .Z(n1513) );
  ANDN U1642 ( .B(n1518), .A(n116), .Z(n1516) );
  XNOR U1643 ( .A(a[900]), .B(n1519), .Z(n116) );
  IV U1644 ( .A(n1517), .Z(n1519) );
  XNOR U1645 ( .A(b[900]), .B(n1517), .Z(n1518) );
  XOR U1646 ( .A(n1520), .B(n1521), .Z(n1517) );
  ANDN U1647 ( .B(n1522), .A(n119), .Z(n1520) );
  XNOR U1648 ( .A(a[899]), .B(n1523), .Z(n119) );
  IV U1649 ( .A(n1521), .Z(n1523) );
  XNOR U1650 ( .A(b[899]), .B(n1521), .Z(n1522) );
  XOR U1651 ( .A(n1524), .B(n1525), .Z(n1521) );
  ANDN U1652 ( .B(n1526), .A(n120), .Z(n1524) );
  XNOR U1653 ( .A(a[898]), .B(n1527), .Z(n120) );
  IV U1654 ( .A(n1525), .Z(n1527) );
  XNOR U1655 ( .A(b[898]), .B(n1525), .Z(n1526) );
  XOR U1656 ( .A(n1528), .B(n1529), .Z(n1525) );
  ANDN U1657 ( .B(n1530), .A(n121), .Z(n1528) );
  XNOR U1658 ( .A(a[897]), .B(n1531), .Z(n121) );
  IV U1659 ( .A(n1529), .Z(n1531) );
  XNOR U1660 ( .A(b[897]), .B(n1529), .Z(n1530) );
  XOR U1661 ( .A(n1532), .B(n1533), .Z(n1529) );
  ANDN U1662 ( .B(n1534), .A(n122), .Z(n1532) );
  XNOR U1663 ( .A(a[896]), .B(n1535), .Z(n122) );
  IV U1664 ( .A(n1533), .Z(n1535) );
  XNOR U1665 ( .A(b[896]), .B(n1533), .Z(n1534) );
  XOR U1666 ( .A(n1536), .B(n1537), .Z(n1533) );
  ANDN U1667 ( .B(n1538), .A(n123), .Z(n1536) );
  XNOR U1668 ( .A(a[895]), .B(n1539), .Z(n123) );
  IV U1669 ( .A(n1537), .Z(n1539) );
  XNOR U1670 ( .A(b[895]), .B(n1537), .Z(n1538) );
  XOR U1671 ( .A(n1540), .B(n1541), .Z(n1537) );
  ANDN U1672 ( .B(n1542), .A(n124), .Z(n1540) );
  XNOR U1673 ( .A(a[894]), .B(n1543), .Z(n124) );
  IV U1674 ( .A(n1541), .Z(n1543) );
  XNOR U1675 ( .A(b[894]), .B(n1541), .Z(n1542) );
  XOR U1676 ( .A(n1544), .B(n1545), .Z(n1541) );
  ANDN U1677 ( .B(n1546), .A(n125), .Z(n1544) );
  XNOR U1678 ( .A(a[893]), .B(n1547), .Z(n125) );
  IV U1679 ( .A(n1545), .Z(n1547) );
  XNOR U1680 ( .A(b[893]), .B(n1545), .Z(n1546) );
  XOR U1681 ( .A(n1548), .B(n1549), .Z(n1545) );
  ANDN U1682 ( .B(n1550), .A(n126), .Z(n1548) );
  XNOR U1683 ( .A(a[892]), .B(n1551), .Z(n126) );
  IV U1684 ( .A(n1549), .Z(n1551) );
  XNOR U1685 ( .A(b[892]), .B(n1549), .Z(n1550) );
  XOR U1686 ( .A(n1552), .B(n1553), .Z(n1549) );
  ANDN U1687 ( .B(n1554), .A(n127), .Z(n1552) );
  XNOR U1688 ( .A(a[891]), .B(n1555), .Z(n127) );
  IV U1689 ( .A(n1553), .Z(n1555) );
  XNOR U1690 ( .A(b[891]), .B(n1553), .Z(n1554) );
  XOR U1691 ( .A(n1556), .B(n1557), .Z(n1553) );
  ANDN U1692 ( .B(n1558), .A(n128), .Z(n1556) );
  XNOR U1693 ( .A(a[890]), .B(n1559), .Z(n128) );
  IV U1694 ( .A(n1557), .Z(n1559) );
  XNOR U1695 ( .A(b[890]), .B(n1557), .Z(n1558) );
  XOR U1696 ( .A(n1560), .B(n1561), .Z(n1557) );
  ANDN U1697 ( .B(n1562), .A(n130), .Z(n1560) );
  XNOR U1698 ( .A(a[889]), .B(n1563), .Z(n130) );
  IV U1699 ( .A(n1561), .Z(n1563) );
  XNOR U1700 ( .A(b[889]), .B(n1561), .Z(n1562) );
  XOR U1701 ( .A(n1564), .B(n1565), .Z(n1561) );
  ANDN U1702 ( .B(n1566), .A(n131), .Z(n1564) );
  XNOR U1703 ( .A(a[888]), .B(n1567), .Z(n131) );
  IV U1704 ( .A(n1565), .Z(n1567) );
  XNOR U1705 ( .A(b[888]), .B(n1565), .Z(n1566) );
  XOR U1706 ( .A(n1568), .B(n1569), .Z(n1565) );
  ANDN U1707 ( .B(n1570), .A(n132), .Z(n1568) );
  XNOR U1708 ( .A(a[887]), .B(n1571), .Z(n132) );
  IV U1709 ( .A(n1569), .Z(n1571) );
  XNOR U1710 ( .A(b[887]), .B(n1569), .Z(n1570) );
  XOR U1711 ( .A(n1572), .B(n1573), .Z(n1569) );
  ANDN U1712 ( .B(n1574), .A(n133), .Z(n1572) );
  XNOR U1713 ( .A(a[886]), .B(n1575), .Z(n133) );
  IV U1714 ( .A(n1573), .Z(n1575) );
  XNOR U1715 ( .A(b[886]), .B(n1573), .Z(n1574) );
  XOR U1716 ( .A(n1576), .B(n1577), .Z(n1573) );
  ANDN U1717 ( .B(n1578), .A(n134), .Z(n1576) );
  XNOR U1718 ( .A(a[885]), .B(n1579), .Z(n134) );
  IV U1719 ( .A(n1577), .Z(n1579) );
  XNOR U1720 ( .A(b[885]), .B(n1577), .Z(n1578) );
  XOR U1721 ( .A(n1580), .B(n1581), .Z(n1577) );
  ANDN U1722 ( .B(n1582), .A(n135), .Z(n1580) );
  XNOR U1723 ( .A(a[884]), .B(n1583), .Z(n135) );
  IV U1724 ( .A(n1581), .Z(n1583) );
  XNOR U1725 ( .A(b[884]), .B(n1581), .Z(n1582) );
  XOR U1726 ( .A(n1584), .B(n1585), .Z(n1581) );
  ANDN U1727 ( .B(n1586), .A(n136), .Z(n1584) );
  XNOR U1728 ( .A(a[883]), .B(n1587), .Z(n136) );
  IV U1729 ( .A(n1585), .Z(n1587) );
  XNOR U1730 ( .A(b[883]), .B(n1585), .Z(n1586) );
  XOR U1731 ( .A(n1588), .B(n1589), .Z(n1585) );
  ANDN U1732 ( .B(n1590), .A(n137), .Z(n1588) );
  XNOR U1733 ( .A(a[882]), .B(n1591), .Z(n137) );
  IV U1734 ( .A(n1589), .Z(n1591) );
  XNOR U1735 ( .A(b[882]), .B(n1589), .Z(n1590) );
  XOR U1736 ( .A(n1592), .B(n1593), .Z(n1589) );
  ANDN U1737 ( .B(n1594), .A(n138), .Z(n1592) );
  XNOR U1738 ( .A(a[881]), .B(n1595), .Z(n138) );
  IV U1739 ( .A(n1593), .Z(n1595) );
  XNOR U1740 ( .A(b[881]), .B(n1593), .Z(n1594) );
  XOR U1741 ( .A(n1596), .B(n1597), .Z(n1593) );
  ANDN U1742 ( .B(n1598), .A(n139), .Z(n1596) );
  XNOR U1743 ( .A(a[880]), .B(n1599), .Z(n139) );
  IV U1744 ( .A(n1597), .Z(n1599) );
  XNOR U1745 ( .A(b[880]), .B(n1597), .Z(n1598) );
  XOR U1746 ( .A(n1600), .B(n1601), .Z(n1597) );
  ANDN U1747 ( .B(n1602), .A(n141), .Z(n1600) );
  XNOR U1748 ( .A(a[879]), .B(n1603), .Z(n141) );
  IV U1749 ( .A(n1601), .Z(n1603) );
  XNOR U1750 ( .A(b[879]), .B(n1601), .Z(n1602) );
  XOR U1751 ( .A(n1604), .B(n1605), .Z(n1601) );
  ANDN U1752 ( .B(n1606), .A(n142), .Z(n1604) );
  XNOR U1753 ( .A(a[878]), .B(n1607), .Z(n142) );
  IV U1754 ( .A(n1605), .Z(n1607) );
  XNOR U1755 ( .A(b[878]), .B(n1605), .Z(n1606) );
  XOR U1756 ( .A(n1608), .B(n1609), .Z(n1605) );
  ANDN U1757 ( .B(n1610), .A(n143), .Z(n1608) );
  XNOR U1758 ( .A(a[877]), .B(n1611), .Z(n143) );
  IV U1759 ( .A(n1609), .Z(n1611) );
  XNOR U1760 ( .A(b[877]), .B(n1609), .Z(n1610) );
  XOR U1761 ( .A(n1612), .B(n1613), .Z(n1609) );
  ANDN U1762 ( .B(n1614), .A(n144), .Z(n1612) );
  XNOR U1763 ( .A(a[876]), .B(n1615), .Z(n144) );
  IV U1764 ( .A(n1613), .Z(n1615) );
  XNOR U1765 ( .A(b[876]), .B(n1613), .Z(n1614) );
  XOR U1766 ( .A(n1616), .B(n1617), .Z(n1613) );
  ANDN U1767 ( .B(n1618), .A(n145), .Z(n1616) );
  XNOR U1768 ( .A(a[875]), .B(n1619), .Z(n145) );
  IV U1769 ( .A(n1617), .Z(n1619) );
  XNOR U1770 ( .A(b[875]), .B(n1617), .Z(n1618) );
  XOR U1771 ( .A(n1620), .B(n1621), .Z(n1617) );
  ANDN U1772 ( .B(n1622), .A(n146), .Z(n1620) );
  XNOR U1773 ( .A(a[874]), .B(n1623), .Z(n146) );
  IV U1774 ( .A(n1621), .Z(n1623) );
  XNOR U1775 ( .A(b[874]), .B(n1621), .Z(n1622) );
  XOR U1776 ( .A(n1624), .B(n1625), .Z(n1621) );
  ANDN U1777 ( .B(n1626), .A(n147), .Z(n1624) );
  XNOR U1778 ( .A(a[873]), .B(n1627), .Z(n147) );
  IV U1779 ( .A(n1625), .Z(n1627) );
  XNOR U1780 ( .A(b[873]), .B(n1625), .Z(n1626) );
  XOR U1781 ( .A(n1628), .B(n1629), .Z(n1625) );
  ANDN U1782 ( .B(n1630), .A(n148), .Z(n1628) );
  XNOR U1783 ( .A(a[872]), .B(n1631), .Z(n148) );
  IV U1784 ( .A(n1629), .Z(n1631) );
  XNOR U1785 ( .A(b[872]), .B(n1629), .Z(n1630) );
  XOR U1786 ( .A(n1632), .B(n1633), .Z(n1629) );
  ANDN U1787 ( .B(n1634), .A(n149), .Z(n1632) );
  XNOR U1788 ( .A(a[871]), .B(n1635), .Z(n149) );
  IV U1789 ( .A(n1633), .Z(n1635) );
  XNOR U1790 ( .A(b[871]), .B(n1633), .Z(n1634) );
  XOR U1791 ( .A(n1636), .B(n1637), .Z(n1633) );
  ANDN U1792 ( .B(n1638), .A(n150), .Z(n1636) );
  XNOR U1793 ( .A(a[870]), .B(n1639), .Z(n150) );
  IV U1794 ( .A(n1637), .Z(n1639) );
  XNOR U1795 ( .A(b[870]), .B(n1637), .Z(n1638) );
  XOR U1796 ( .A(n1640), .B(n1641), .Z(n1637) );
  ANDN U1797 ( .B(n1642), .A(n152), .Z(n1640) );
  XNOR U1798 ( .A(a[869]), .B(n1643), .Z(n152) );
  IV U1799 ( .A(n1641), .Z(n1643) );
  XNOR U1800 ( .A(b[869]), .B(n1641), .Z(n1642) );
  XOR U1801 ( .A(n1644), .B(n1645), .Z(n1641) );
  ANDN U1802 ( .B(n1646), .A(n153), .Z(n1644) );
  XNOR U1803 ( .A(a[868]), .B(n1647), .Z(n153) );
  IV U1804 ( .A(n1645), .Z(n1647) );
  XNOR U1805 ( .A(b[868]), .B(n1645), .Z(n1646) );
  XOR U1806 ( .A(n1648), .B(n1649), .Z(n1645) );
  ANDN U1807 ( .B(n1650), .A(n154), .Z(n1648) );
  XNOR U1808 ( .A(a[867]), .B(n1651), .Z(n154) );
  IV U1809 ( .A(n1649), .Z(n1651) );
  XNOR U1810 ( .A(b[867]), .B(n1649), .Z(n1650) );
  XOR U1811 ( .A(n1652), .B(n1653), .Z(n1649) );
  ANDN U1812 ( .B(n1654), .A(n155), .Z(n1652) );
  XNOR U1813 ( .A(a[866]), .B(n1655), .Z(n155) );
  IV U1814 ( .A(n1653), .Z(n1655) );
  XNOR U1815 ( .A(b[866]), .B(n1653), .Z(n1654) );
  XOR U1816 ( .A(n1656), .B(n1657), .Z(n1653) );
  ANDN U1817 ( .B(n1658), .A(n156), .Z(n1656) );
  XNOR U1818 ( .A(a[865]), .B(n1659), .Z(n156) );
  IV U1819 ( .A(n1657), .Z(n1659) );
  XNOR U1820 ( .A(b[865]), .B(n1657), .Z(n1658) );
  XOR U1821 ( .A(n1660), .B(n1661), .Z(n1657) );
  ANDN U1822 ( .B(n1662), .A(n157), .Z(n1660) );
  XNOR U1823 ( .A(a[864]), .B(n1663), .Z(n157) );
  IV U1824 ( .A(n1661), .Z(n1663) );
  XNOR U1825 ( .A(b[864]), .B(n1661), .Z(n1662) );
  XOR U1826 ( .A(n1664), .B(n1665), .Z(n1661) );
  ANDN U1827 ( .B(n1666), .A(n158), .Z(n1664) );
  XNOR U1828 ( .A(a[863]), .B(n1667), .Z(n158) );
  IV U1829 ( .A(n1665), .Z(n1667) );
  XNOR U1830 ( .A(b[863]), .B(n1665), .Z(n1666) );
  XOR U1831 ( .A(n1668), .B(n1669), .Z(n1665) );
  ANDN U1832 ( .B(n1670), .A(n159), .Z(n1668) );
  XNOR U1833 ( .A(a[862]), .B(n1671), .Z(n159) );
  IV U1834 ( .A(n1669), .Z(n1671) );
  XNOR U1835 ( .A(b[862]), .B(n1669), .Z(n1670) );
  XOR U1836 ( .A(n1672), .B(n1673), .Z(n1669) );
  ANDN U1837 ( .B(n1674), .A(n160), .Z(n1672) );
  XNOR U1838 ( .A(a[861]), .B(n1675), .Z(n160) );
  IV U1839 ( .A(n1673), .Z(n1675) );
  XNOR U1840 ( .A(b[861]), .B(n1673), .Z(n1674) );
  XOR U1841 ( .A(n1676), .B(n1677), .Z(n1673) );
  ANDN U1842 ( .B(n1678), .A(n161), .Z(n1676) );
  XNOR U1843 ( .A(a[860]), .B(n1679), .Z(n161) );
  IV U1844 ( .A(n1677), .Z(n1679) );
  XNOR U1845 ( .A(b[860]), .B(n1677), .Z(n1678) );
  XOR U1846 ( .A(n1680), .B(n1681), .Z(n1677) );
  ANDN U1847 ( .B(n1682), .A(n163), .Z(n1680) );
  XNOR U1848 ( .A(a[859]), .B(n1683), .Z(n163) );
  IV U1849 ( .A(n1681), .Z(n1683) );
  XNOR U1850 ( .A(b[859]), .B(n1681), .Z(n1682) );
  XOR U1851 ( .A(n1684), .B(n1685), .Z(n1681) );
  ANDN U1852 ( .B(n1686), .A(n164), .Z(n1684) );
  XNOR U1853 ( .A(a[858]), .B(n1687), .Z(n164) );
  IV U1854 ( .A(n1685), .Z(n1687) );
  XNOR U1855 ( .A(b[858]), .B(n1685), .Z(n1686) );
  XOR U1856 ( .A(n1688), .B(n1689), .Z(n1685) );
  ANDN U1857 ( .B(n1690), .A(n165), .Z(n1688) );
  XNOR U1858 ( .A(a[857]), .B(n1691), .Z(n165) );
  IV U1859 ( .A(n1689), .Z(n1691) );
  XNOR U1860 ( .A(b[857]), .B(n1689), .Z(n1690) );
  XOR U1861 ( .A(n1692), .B(n1693), .Z(n1689) );
  ANDN U1862 ( .B(n1694), .A(n166), .Z(n1692) );
  XNOR U1863 ( .A(a[856]), .B(n1695), .Z(n166) );
  IV U1864 ( .A(n1693), .Z(n1695) );
  XNOR U1865 ( .A(b[856]), .B(n1693), .Z(n1694) );
  XOR U1866 ( .A(n1696), .B(n1697), .Z(n1693) );
  ANDN U1867 ( .B(n1698), .A(n167), .Z(n1696) );
  XNOR U1868 ( .A(a[855]), .B(n1699), .Z(n167) );
  IV U1869 ( .A(n1697), .Z(n1699) );
  XNOR U1870 ( .A(b[855]), .B(n1697), .Z(n1698) );
  XOR U1871 ( .A(n1700), .B(n1701), .Z(n1697) );
  ANDN U1872 ( .B(n1702), .A(n168), .Z(n1700) );
  XNOR U1873 ( .A(a[854]), .B(n1703), .Z(n168) );
  IV U1874 ( .A(n1701), .Z(n1703) );
  XNOR U1875 ( .A(b[854]), .B(n1701), .Z(n1702) );
  XOR U1876 ( .A(n1704), .B(n1705), .Z(n1701) );
  ANDN U1877 ( .B(n1706), .A(n169), .Z(n1704) );
  XNOR U1878 ( .A(a[853]), .B(n1707), .Z(n169) );
  IV U1879 ( .A(n1705), .Z(n1707) );
  XNOR U1880 ( .A(b[853]), .B(n1705), .Z(n1706) );
  XOR U1881 ( .A(n1708), .B(n1709), .Z(n1705) );
  ANDN U1882 ( .B(n1710), .A(n170), .Z(n1708) );
  XNOR U1883 ( .A(a[852]), .B(n1711), .Z(n170) );
  IV U1884 ( .A(n1709), .Z(n1711) );
  XNOR U1885 ( .A(b[852]), .B(n1709), .Z(n1710) );
  XOR U1886 ( .A(n1712), .B(n1713), .Z(n1709) );
  ANDN U1887 ( .B(n1714), .A(n171), .Z(n1712) );
  XNOR U1888 ( .A(a[851]), .B(n1715), .Z(n171) );
  IV U1889 ( .A(n1713), .Z(n1715) );
  XNOR U1890 ( .A(b[851]), .B(n1713), .Z(n1714) );
  XOR U1891 ( .A(n1716), .B(n1717), .Z(n1713) );
  ANDN U1892 ( .B(n1718), .A(n172), .Z(n1716) );
  XNOR U1893 ( .A(a[850]), .B(n1719), .Z(n172) );
  IV U1894 ( .A(n1717), .Z(n1719) );
  XNOR U1895 ( .A(b[850]), .B(n1717), .Z(n1718) );
  XOR U1896 ( .A(n1720), .B(n1721), .Z(n1717) );
  ANDN U1897 ( .B(n1722), .A(n174), .Z(n1720) );
  XNOR U1898 ( .A(a[849]), .B(n1723), .Z(n174) );
  IV U1899 ( .A(n1721), .Z(n1723) );
  XNOR U1900 ( .A(b[849]), .B(n1721), .Z(n1722) );
  XOR U1901 ( .A(n1724), .B(n1725), .Z(n1721) );
  ANDN U1902 ( .B(n1726), .A(n175), .Z(n1724) );
  XNOR U1903 ( .A(a[848]), .B(n1727), .Z(n175) );
  IV U1904 ( .A(n1725), .Z(n1727) );
  XNOR U1905 ( .A(b[848]), .B(n1725), .Z(n1726) );
  XOR U1906 ( .A(n1728), .B(n1729), .Z(n1725) );
  ANDN U1907 ( .B(n1730), .A(n176), .Z(n1728) );
  XNOR U1908 ( .A(a[847]), .B(n1731), .Z(n176) );
  IV U1909 ( .A(n1729), .Z(n1731) );
  XNOR U1910 ( .A(b[847]), .B(n1729), .Z(n1730) );
  XOR U1911 ( .A(n1732), .B(n1733), .Z(n1729) );
  ANDN U1912 ( .B(n1734), .A(n177), .Z(n1732) );
  XNOR U1913 ( .A(a[846]), .B(n1735), .Z(n177) );
  IV U1914 ( .A(n1733), .Z(n1735) );
  XNOR U1915 ( .A(b[846]), .B(n1733), .Z(n1734) );
  XOR U1916 ( .A(n1736), .B(n1737), .Z(n1733) );
  ANDN U1917 ( .B(n1738), .A(n178), .Z(n1736) );
  XNOR U1918 ( .A(a[845]), .B(n1739), .Z(n178) );
  IV U1919 ( .A(n1737), .Z(n1739) );
  XNOR U1920 ( .A(b[845]), .B(n1737), .Z(n1738) );
  XOR U1921 ( .A(n1740), .B(n1741), .Z(n1737) );
  ANDN U1922 ( .B(n1742), .A(n179), .Z(n1740) );
  XNOR U1923 ( .A(a[844]), .B(n1743), .Z(n179) );
  IV U1924 ( .A(n1741), .Z(n1743) );
  XNOR U1925 ( .A(b[844]), .B(n1741), .Z(n1742) );
  XOR U1926 ( .A(n1744), .B(n1745), .Z(n1741) );
  ANDN U1927 ( .B(n1746), .A(n180), .Z(n1744) );
  XNOR U1928 ( .A(a[843]), .B(n1747), .Z(n180) );
  IV U1929 ( .A(n1745), .Z(n1747) );
  XNOR U1930 ( .A(b[843]), .B(n1745), .Z(n1746) );
  XOR U1931 ( .A(n1748), .B(n1749), .Z(n1745) );
  ANDN U1932 ( .B(n1750), .A(n181), .Z(n1748) );
  XNOR U1933 ( .A(a[842]), .B(n1751), .Z(n181) );
  IV U1934 ( .A(n1749), .Z(n1751) );
  XNOR U1935 ( .A(b[842]), .B(n1749), .Z(n1750) );
  XOR U1936 ( .A(n1752), .B(n1753), .Z(n1749) );
  ANDN U1937 ( .B(n1754), .A(n182), .Z(n1752) );
  XNOR U1938 ( .A(a[841]), .B(n1755), .Z(n182) );
  IV U1939 ( .A(n1753), .Z(n1755) );
  XNOR U1940 ( .A(b[841]), .B(n1753), .Z(n1754) );
  XOR U1941 ( .A(n1756), .B(n1757), .Z(n1753) );
  ANDN U1942 ( .B(n1758), .A(n183), .Z(n1756) );
  XNOR U1943 ( .A(a[840]), .B(n1759), .Z(n183) );
  IV U1944 ( .A(n1757), .Z(n1759) );
  XNOR U1945 ( .A(b[840]), .B(n1757), .Z(n1758) );
  XOR U1946 ( .A(n1760), .B(n1761), .Z(n1757) );
  ANDN U1947 ( .B(n1762), .A(n185), .Z(n1760) );
  XNOR U1948 ( .A(a[839]), .B(n1763), .Z(n185) );
  IV U1949 ( .A(n1761), .Z(n1763) );
  XNOR U1950 ( .A(b[839]), .B(n1761), .Z(n1762) );
  XOR U1951 ( .A(n1764), .B(n1765), .Z(n1761) );
  ANDN U1952 ( .B(n1766), .A(n186), .Z(n1764) );
  XNOR U1953 ( .A(a[838]), .B(n1767), .Z(n186) );
  IV U1954 ( .A(n1765), .Z(n1767) );
  XNOR U1955 ( .A(b[838]), .B(n1765), .Z(n1766) );
  XOR U1956 ( .A(n1768), .B(n1769), .Z(n1765) );
  ANDN U1957 ( .B(n1770), .A(n187), .Z(n1768) );
  XNOR U1958 ( .A(a[837]), .B(n1771), .Z(n187) );
  IV U1959 ( .A(n1769), .Z(n1771) );
  XNOR U1960 ( .A(b[837]), .B(n1769), .Z(n1770) );
  XOR U1961 ( .A(n1772), .B(n1773), .Z(n1769) );
  ANDN U1962 ( .B(n1774), .A(n188), .Z(n1772) );
  XNOR U1963 ( .A(a[836]), .B(n1775), .Z(n188) );
  IV U1964 ( .A(n1773), .Z(n1775) );
  XNOR U1965 ( .A(b[836]), .B(n1773), .Z(n1774) );
  XOR U1966 ( .A(n1776), .B(n1777), .Z(n1773) );
  ANDN U1967 ( .B(n1778), .A(n189), .Z(n1776) );
  XNOR U1968 ( .A(a[835]), .B(n1779), .Z(n189) );
  IV U1969 ( .A(n1777), .Z(n1779) );
  XNOR U1970 ( .A(b[835]), .B(n1777), .Z(n1778) );
  XOR U1971 ( .A(n1780), .B(n1781), .Z(n1777) );
  ANDN U1972 ( .B(n1782), .A(n190), .Z(n1780) );
  XNOR U1973 ( .A(a[834]), .B(n1783), .Z(n190) );
  IV U1974 ( .A(n1781), .Z(n1783) );
  XNOR U1975 ( .A(b[834]), .B(n1781), .Z(n1782) );
  XOR U1976 ( .A(n1784), .B(n1785), .Z(n1781) );
  ANDN U1977 ( .B(n1786), .A(n191), .Z(n1784) );
  XNOR U1978 ( .A(a[833]), .B(n1787), .Z(n191) );
  IV U1979 ( .A(n1785), .Z(n1787) );
  XNOR U1980 ( .A(b[833]), .B(n1785), .Z(n1786) );
  XOR U1981 ( .A(n1788), .B(n1789), .Z(n1785) );
  ANDN U1982 ( .B(n1790), .A(n192), .Z(n1788) );
  XNOR U1983 ( .A(a[832]), .B(n1791), .Z(n192) );
  IV U1984 ( .A(n1789), .Z(n1791) );
  XNOR U1985 ( .A(b[832]), .B(n1789), .Z(n1790) );
  XOR U1986 ( .A(n1792), .B(n1793), .Z(n1789) );
  ANDN U1987 ( .B(n1794), .A(n193), .Z(n1792) );
  XNOR U1988 ( .A(a[831]), .B(n1795), .Z(n193) );
  IV U1989 ( .A(n1793), .Z(n1795) );
  XNOR U1990 ( .A(b[831]), .B(n1793), .Z(n1794) );
  XOR U1991 ( .A(n1796), .B(n1797), .Z(n1793) );
  ANDN U1992 ( .B(n1798), .A(n194), .Z(n1796) );
  XNOR U1993 ( .A(a[830]), .B(n1799), .Z(n194) );
  IV U1994 ( .A(n1797), .Z(n1799) );
  XNOR U1995 ( .A(b[830]), .B(n1797), .Z(n1798) );
  XOR U1996 ( .A(n1800), .B(n1801), .Z(n1797) );
  ANDN U1997 ( .B(n1802), .A(n196), .Z(n1800) );
  XNOR U1998 ( .A(a[829]), .B(n1803), .Z(n196) );
  IV U1999 ( .A(n1801), .Z(n1803) );
  XNOR U2000 ( .A(b[829]), .B(n1801), .Z(n1802) );
  XOR U2001 ( .A(n1804), .B(n1805), .Z(n1801) );
  ANDN U2002 ( .B(n1806), .A(n197), .Z(n1804) );
  XNOR U2003 ( .A(a[828]), .B(n1807), .Z(n197) );
  IV U2004 ( .A(n1805), .Z(n1807) );
  XNOR U2005 ( .A(b[828]), .B(n1805), .Z(n1806) );
  XOR U2006 ( .A(n1808), .B(n1809), .Z(n1805) );
  ANDN U2007 ( .B(n1810), .A(n198), .Z(n1808) );
  XNOR U2008 ( .A(a[827]), .B(n1811), .Z(n198) );
  IV U2009 ( .A(n1809), .Z(n1811) );
  XNOR U2010 ( .A(b[827]), .B(n1809), .Z(n1810) );
  XOR U2011 ( .A(n1812), .B(n1813), .Z(n1809) );
  ANDN U2012 ( .B(n1814), .A(n199), .Z(n1812) );
  XNOR U2013 ( .A(a[826]), .B(n1815), .Z(n199) );
  IV U2014 ( .A(n1813), .Z(n1815) );
  XNOR U2015 ( .A(b[826]), .B(n1813), .Z(n1814) );
  XOR U2016 ( .A(n1816), .B(n1817), .Z(n1813) );
  ANDN U2017 ( .B(n1818), .A(n200), .Z(n1816) );
  XNOR U2018 ( .A(a[825]), .B(n1819), .Z(n200) );
  IV U2019 ( .A(n1817), .Z(n1819) );
  XNOR U2020 ( .A(b[825]), .B(n1817), .Z(n1818) );
  XOR U2021 ( .A(n1820), .B(n1821), .Z(n1817) );
  ANDN U2022 ( .B(n1822), .A(n201), .Z(n1820) );
  XNOR U2023 ( .A(a[824]), .B(n1823), .Z(n201) );
  IV U2024 ( .A(n1821), .Z(n1823) );
  XNOR U2025 ( .A(b[824]), .B(n1821), .Z(n1822) );
  XOR U2026 ( .A(n1824), .B(n1825), .Z(n1821) );
  ANDN U2027 ( .B(n1826), .A(n202), .Z(n1824) );
  XNOR U2028 ( .A(a[823]), .B(n1827), .Z(n202) );
  IV U2029 ( .A(n1825), .Z(n1827) );
  XNOR U2030 ( .A(b[823]), .B(n1825), .Z(n1826) );
  XOR U2031 ( .A(n1828), .B(n1829), .Z(n1825) );
  ANDN U2032 ( .B(n1830), .A(n203), .Z(n1828) );
  XNOR U2033 ( .A(a[822]), .B(n1831), .Z(n203) );
  IV U2034 ( .A(n1829), .Z(n1831) );
  XNOR U2035 ( .A(b[822]), .B(n1829), .Z(n1830) );
  XOR U2036 ( .A(n1832), .B(n1833), .Z(n1829) );
  ANDN U2037 ( .B(n1834), .A(n204), .Z(n1832) );
  XNOR U2038 ( .A(a[821]), .B(n1835), .Z(n204) );
  IV U2039 ( .A(n1833), .Z(n1835) );
  XNOR U2040 ( .A(b[821]), .B(n1833), .Z(n1834) );
  XOR U2041 ( .A(n1836), .B(n1837), .Z(n1833) );
  ANDN U2042 ( .B(n1838), .A(n205), .Z(n1836) );
  XNOR U2043 ( .A(a[820]), .B(n1839), .Z(n205) );
  IV U2044 ( .A(n1837), .Z(n1839) );
  XNOR U2045 ( .A(b[820]), .B(n1837), .Z(n1838) );
  XOR U2046 ( .A(n1840), .B(n1841), .Z(n1837) );
  ANDN U2047 ( .B(n1842), .A(n207), .Z(n1840) );
  XNOR U2048 ( .A(a[819]), .B(n1843), .Z(n207) );
  IV U2049 ( .A(n1841), .Z(n1843) );
  XNOR U2050 ( .A(b[819]), .B(n1841), .Z(n1842) );
  XOR U2051 ( .A(n1844), .B(n1845), .Z(n1841) );
  ANDN U2052 ( .B(n1846), .A(n208), .Z(n1844) );
  XNOR U2053 ( .A(a[818]), .B(n1847), .Z(n208) );
  IV U2054 ( .A(n1845), .Z(n1847) );
  XNOR U2055 ( .A(b[818]), .B(n1845), .Z(n1846) );
  XOR U2056 ( .A(n1848), .B(n1849), .Z(n1845) );
  ANDN U2057 ( .B(n1850), .A(n209), .Z(n1848) );
  XNOR U2058 ( .A(a[817]), .B(n1851), .Z(n209) );
  IV U2059 ( .A(n1849), .Z(n1851) );
  XNOR U2060 ( .A(b[817]), .B(n1849), .Z(n1850) );
  XOR U2061 ( .A(n1852), .B(n1853), .Z(n1849) );
  ANDN U2062 ( .B(n1854), .A(n210), .Z(n1852) );
  XNOR U2063 ( .A(a[816]), .B(n1855), .Z(n210) );
  IV U2064 ( .A(n1853), .Z(n1855) );
  XNOR U2065 ( .A(b[816]), .B(n1853), .Z(n1854) );
  XOR U2066 ( .A(n1856), .B(n1857), .Z(n1853) );
  ANDN U2067 ( .B(n1858), .A(n211), .Z(n1856) );
  XNOR U2068 ( .A(a[815]), .B(n1859), .Z(n211) );
  IV U2069 ( .A(n1857), .Z(n1859) );
  XNOR U2070 ( .A(b[815]), .B(n1857), .Z(n1858) );
  XOR U2071 ( .A(n1860), .B(n1861), .Z(n1857) );
  ANDN U2072 ( .B(n1862), .A(n212), .Z(n1860) );
  XNOR U2073 ( .A(a[814]), .B(n1863), .Z(n212) );
  IV U2074 ( .A(n1861), .Z(n1863) );
  XNOR U2075 ( .A(b[814]), .B(n1861), .Z(n1862) );
  XOR U2076 ( .A(n1864), .B(n1865), .Z(n1861) );
  ANDN U2077 ( .B(n1866), .A(n213), .Z(n1864) );
  XNOR U2078 ( .A(a[813]), .B(n1867), .Z(n213) );
  IV U2079 ( .A(n1865), .Z(n1867) );
  XNOR U2080 ( .A(b[813]), .B(n1865), .Z(n1866) );
  XOR U2081 ( .A(n1868), .B(n1869), .Z(n1865) );
  ANDN U2082 ( .B(n1870), .A(n214), .Z(n1868) );
  XNOR U2083 ( .A(a[812]), .B(n1871), .Z(n214) );
  IV U2084 ( .A(n1869), .Z(n1871) );
  XNOR U2085 ( .A(b[812]), .B(n1869), .Z(n1870) );
  XOR U2086 ( .A(n1872), .B(n1873), .Z(n1869) );
  ANDN U2087 ( .B(n1874), .A(n215), .Z(n1872) );
  XNOR U2088 ( .A(a[811]), .B(n1875), .Z(n215) );
  IV U2089 ( .A(n1873), .Z(n1875) );
  XNOR U2090 ( .A(b[811]), .B(n1873), .Z(n1874) );
  XOR U2091 ( .A(n1876), .B(n1877), .Z(n1873) );
  ANDN U2092 ( .B(n1878), .A(n216), .Z(n1876) );
  XNOR U2093 ( .A(a[810]), .B(n1879), .Z(n216) );
  IV U2094 ( .A(n1877), .Z(n1879) );
  XNOR U2095 ( .A(b[810]), .B(n1877), .Z(n1878) );
  XOR U2096 ( .A(n1880), .B(n1881), .Z(n1877) );
  ANDN U2097 ( .B(n1882), .A(n218), .Z(n1880) );
  XNOR U2098 ( .A(a[809]), .B(n1883), .Z(n218) );
  IV U2099 ( .A(n1881), .Z(n1883) );
  XNOR U2100 ( .A(b[809]), .B(n1881), .Z(n1882) );
  XOR U2101 ( .A(n1884), .B(n1885), .Z(n1881) );
  ANDN U2102 ( .B(n1886), .A(n219), .Z(n1884) );
  XNOR U2103 ( .A(a[808]), .B(n1887), .Z(n219) );
  IV U2104 ( .A(n1885), .Z(n1887) );
  XNOR U2105 ( .A(b[808]), .B(n1885), .Z(n1886) );
  XOR U2106 ( .A(n1888), .B(n1889), .Z(n1885) );
  ANDN U2107 ( .B(n1890), .A(n220), .Z(n1888) );
  XNOR U2108 ( .A(a[807]), .B(n1891), .Z(n220) );
  IV U2109 ( .A(n1889), .Z(n1891) );
  XNOR U2110 ( .A(b[807]), .B(n1889), .Z(n1890) );
  XOR U2111 ( .A(n1892), .B(n1893), .Z(n1889) );
  ANDN U2112 ( .B(n1894), .A(n221), .Z(n1892) );
  XNOR U2113 ( .A(a[806]), .B(n1895), .Z(n221) );
  IV U2114 ( .A(n1893), .Z(n1895) );
  XNOR U2115 ( .A(b[806]), .B(n1893), .Z(n1894) );
  XOR U2116 ( .A(n1896), .B(n1897), .Z(n1893) );
  ANDN U2117 ( .B(n1898), .A(n222), .Z(n1896) );
  XNOR U2118 ( .A(a[805]), .B(n1899), .Z(n222) );
  IV U2119 ( .A(n1897), .Z(n1899) );
  XNOR U2120 ( .A(b[805]), .B(n1897), .Z(n1898) );
  XOR U2121 ( .A(n1900), .B(n1901), .Z(n1897) );
  ANDN U2122 ( .B(n1902), .A(n223), .Z(n1900) );
  XNOR U2123 ( .A(a[804]), .B(n1903), .Z(n223) );
  IV U2124 ( .A(n1901), .Z(n1903) );
  XNOR U2125 ( .A(b[804]), .B(n1901), .Z(n1902) );
  XOR U2126 ( .A(n1904), .B(n1905), .Z(n1901) );
  ANDN U2127 ( .B(n1906), .A(n224), .Z(n1904) );
  XNOR U2128 ( .A(a[803]), .B(n1907), .Z(n224) );
  IV U2129 ( .A(n1905), .Z(n1907) );
  XNOR U2130 ( .A(b[803]), .B(n1905), .Z(n1906) );
  XOR U2131 ( .A(n1908), .B(n1909), .Z(n1905) );
  ANDN U2132 ( .B(n1910), .A(n225), .Z(n1908) );
  XNOR U2133 ( .A(a[802]), .B(n1911), .Z(n225) );
  IV U2134 ( .A(n1909), .Z(n1911) );
  XNOR U2135 ( .A(b[802]), .B(n1909), .Z(n1910) );
  XOR U2136 ( .A(n1912), .B(n1913), .Z(n1909) );
  ANDN U2137 ( .B(n1914), .A(n226), .Z(n1912) );
  XNOR U2138 ( .A(a[801]), .B(n1915), .Z(n226) );
  IV U2139 ( .A(n1913), .Z(n1915) );
  XNOR U2140 ( .A(b[801]), .B(n1913), .Z(n1914) );
  XOR U2141 ( .A(n1916), .B(n1917), .Z(n1913) );
  ANDN U2142 ( .B(n1918), .A(n227), .Z(n1916) );
  XNOR U2143 ( .A(a[800]), .B(n1919), .Z(n227) );
  IV U2144 ( .A(n1917), .Z(n1919) );
  XNOR U2145 ( .A(b[800]), .B(n1917), .Z(n1918) );
  XOR U2146 ( .A(n1920), .B(n1921), .Z(n1917) );
  ANDN U2147 ( .B(n1922), .A(n230), .Z(n1920) );
  XNOR U2148 ( .A(a[799]), .B(n1923), .Z(n230) );
  IV U2149 ( .A(n1921), .Z(n1923) );
  XNOR U2150 ( .A(b[799]), .B(n1921), .Z(n1922) );
  XOR U2151 ( .A(n1924), .B(n1925), .Z(n1921) );
  ANDN U2152 ( .B(n1926), .A(n231), .Z(n1924) );
  XNOR U2153 ( .A(a[798]), .B(n1927), .Z(n231) );
  IV U2154 ( .A(n1925), .Z(n1927) );
  XNOR U2155 ( .A(b[798]), .B(n1925), .Z(n1926) );
  XOR U2156 ( .A(n1928), .B(n1929), .Z(n1925) );
  ANDN U2157 ( .B(n1930), .A(n232), .Z(n1928) );
  XNOR U2158 ( .A(a[797]), .B(n1931), .Z(n232) );
  IV U2159 ( .A(n1929), .Z(n1931) );
  XNOR U2160 ( .A(b[797]), .B(n1929), .Z(n1930) );
  XOR U2161 ( .A(n1932), .B(n1933), .Z(n1929) );
  ANDN U2162 ( .B(n1934), .A(n233), .Z(n1932) );
  XNOR U2163 ( .A(a[796]), .B(n1935), .Z(n233) );
  IV U2164 ( .A(n1933), .Z(n1935) );
  XNOR U2165 ( .A(b[796]), .B(n1933), .Z(n1934) );
  XOR U2166 ( .A(n1936), .B(n1937), .Z(n1933) );
  ANDN U2167 ( .B(n1938), .A(n234), .Z(n1936) );
  XNOR U2168 ( .A(a[795]), .B(n1939), .Z(n234) );
  IV U2169 ( .A(n1937), .Z(n1939) );
  XNOR U2170 ( .A(b[795]), .B(n1937), .Z(n1938) );
  XOR U2171 ( .A(n1940), .B(n1941), .Z(n1937) );
  ANDN U2172 ( .B(n1942), .A(n235), .Z(n1940) );
  XNOR U2173 ( .A(a[794]), .B(n1943), .Z(n235) );
  IV U2174 ( .A(n1941), .Z(n1943) );
  XNOR U2175 ( .A(b[794]), .B(n1941), .Z(n1942) );
  XOR U2176 ( .A(n1944), .B(n1945), .Z(n1941) );
  ANDN U2177 ( .B(n1946), .A(n236), .Z(n1944) );
  XNOR U2178 ( .A(a[793]), .B(n1947), .Z(n236) );
  IV U2179 ( .A(n1945), .Z(n1947) );
  XNOR U2180 ( .A(b[793]), .B(n1945), .Z(n1946) );
  XOR U2181 ( .A(n1948), .B(n1949), .Z(n1945) );
  ANDN U2182 ( .B(n1950), .A(n237), .Z(n1948) );
  XNOR U2183 ( .A(a[792]), .B(n1951), .Z(n237) );
  IV U2184 ( .A(n1949), .Z(n1951) );
  XNOR U2185 ( .A(b[792]), .B(n1949), .Z(n1950) );
  XOR U2186 ( .A(n1952), .B(n1953), .Z(n1949) );
  ANDN U2187 ( .B(n1954), .A(n238), .Z(n1952) );
  XNOR U2188 ( .A(a[791]), .B(n1955), .Z(n238) );
  IV U2189 ( .A(n1953), .Z(n1955) );
  XNOR U2190 ( .A(b[791]), .B(n1953), .Z(n1954) );
  XOR U2191 ( .A(n1956), .B(n1957), .Z(n1953) );
  ANDN U2192 ( .B(n1958), .A(n239), .Z(n1956) );
  XNOR U2193 ( .A(a[790]), .B(n1959), .Z(n239) );
  IV U2194 ( .A(n1957), .Z(n1959) );
  XNOR U2195 ( .A(b[790]), .B(n1957), .Z(n1958) );
  XOR U2196 ( .A(n1960), .B(n1961), .Z(n1957) );
  ANDN U2197 ( .B(n1962), .A(n241), .Z(n1960) );
  XNOR U2198 ( .A(a[789]), .B(n1963), .Z(n241) );
  IV U2199 ( .A(n1961), .Z(n1963) );
  XNOR U2200 ( .A(b[789]), .B(n1961), .Z(n1962) );
  XOR U2201 ( .A(n1964), .B(n1965), .Z(n1961) );
  ANDN U2202 ( .B(n1966), .A(n242), .Z(n1964) );
  XNOR U2203 ( .A(a[788]), .B(n1967), .Z(n242) );
  IV U2204 ( .A(n1965), .Z(n1967) );
  XNOR U2205 ( .A(b[788]), .B(n1965), .Z(n1966) );
  XOR U2206 ( .A(n1968), .B(n1969), .Z(n1965) );
  ANDN U2207 ( .B(n1970), .A(n243), .Z(n1968) );
  XNOR U2208 ( .A(a[787]), .B(n1971), .Z(n243) );
  IV U2209 ( .A(n1969), .Z(n1971) );
  XNOR U2210 ( .A(b[787]), .B(n1969), .Z(n1970) );
  XOR U2211 ( .A(n1972), .B(n1973), .Z(n1969) );
  ANDN U2212 ( .B(n1974), .A(n244), .Z(n1972) );
  XNOR U2213 ( .A(a[786]), .B(n1975), .Z(n244) );
  IV U2214 ( .A(n1973), .Z(n1975) );
  XNOR U2215 ( .A(b[786]), .B(n1973), .Z(n1974) );
  XOR U2216 ( .A(n1976), .B(n1977), .Z(n1973) );
  ANDN U2217 ( .B(n1978), .A(n245), .Z(n1976) );
  XNOR U2218 ( .A(a[785]), .B(n1979), .Z(n245) );
  IV U2219 ( .A(n1977), .Z(n1979) );
  XNOR U2220 ( .A(b[785]), .B(n1977), .Z(n1978) );
  XOR U2221 ( .A(n1980), .B(n1981), .Z(n1977) );
  ANDN U2222 ( .B(n1982), .A(n246), .Z(n1980) );
  XNOR U2223 ( .A(a[784]), .B(n1983), .Z(n246) );
  IV U2224 ( .A(n1981), .Z(n1983) );
  XNOR U2225 ( .A(b[784]), .B(n1981), .Z(n1982) );
  XOR U2226 ( .A(n1984), .B(n1985), .Z(n1981) );
  ANDN U2227 ( .B(n1986), .A(n247), .Z(n1984) );
  XNOR U2228 ( .A(a[783]), .B(n1987), .Z(n247) );
  IV U2229 ( .A(n1985), .Z(n1987) );
  XNOR U2230 ( .A(b[783]), .B(n1985), .Z(n1986) );
  XOR U2231 ( .A(n1988), .B(n1989), .Z(n1985) );
  ANDN U2232 ( .B(n1990), .A(n248), .Z(n1988) );
  XNOR U2233 ( .A(a[782]), .B(n1991), .Z(n248) );
  IV U2234 ( .A(n1989), .Z(n1991) );
  XNOR U2235 ( .A(b[782]), .B(n1989), .Z(n1990) );
  XOR U2236 ( .A(n1992), .B(n1993), .Z(n1989) );
  ANDN U2237 ( .B(n1994), .A(n249), .Z(n1992) );
  XNOR U2238 ( .A(a[781]), .B(n1995), .Z(n249) );
  IV U2239 ( .A(n1993), .Z(n1995) );
  XNOR U2240 ( .A(b[781]), .B(n1993), .Z(n1994) );
  XOR U2241 ( .A(n1996), .B(n1997), .Z(n1993) );
  ANDN U2242 ( .B(n1998), .A(n250), .Z(n1996) );
  XNOR U2243 ( .A(a[780]), .B(n1999), .Z(n250) );
  IV U2244 ( .A(n1997), .Z(n1999) );
  XNOR U2245 ( .A(b[780]), .B(n1997), .Z(n1998) );
  XOR U2246 ( .A(n2000), .B(n2001), .Z(n1997) );
  ANDN U2247 ( .B(n2002), .A(n252), .Z(n2000) );
  XNOR U2248 ( .A(a[779]), .B(n2003), .Z(n252) );
  IV U2249 ( .A(n2001), .Z(n2003) );
  XNOR U2250 ( .A(b[779]), .B(n2001), .Z(n2002) );
  XOR U2251 ( .A(n2004), .B(n2005), .Z(n2001) );
  ANDN U2252 ( .B(n2006), .A(n253), .Z(n2004) );
  XNOR U2253 ( .A(a[778]), .B(n2007), .Z(n253) );
  IV U2254 ( .A(n2005), .Z(n2007) );
  XNOR U2255 ( .A(b[778]), .B(n2005), .Z(n2006) );
  XOR U2256 ( .A(n2008), .B(n2009), .Z(n2005) );
  ANDN U2257 ( .B(n2010), .A(n254), .Z(n2008) );
  XNOR U2258 ( .A(a[777]), .B(n2011), .Z(n254) );
  IV U2259 ( .A(n2009), .Z(n2011) );
  XNOR U2260 ( .A(b[777]), .B(n2009), .Z(n2010) );
  XOR U2261 ( .A(n2012), .B(n2013), .Z(n2009) );
  ANDN U2262 ( .B(n2014), .A(n255), .Z(n2012) );
  XNOR U2263 ( .A(a[776]), .B(n2015), .Z(n255) );
  IV U2264 ( .A(n2013), .Z(n2015) );
  XNOR U2265 ( .A(b[776]), .B(n2013), .Z(n2014) );
  XOR U2266 ( .A(n2016), .B(n2017), .Z(n2013) );
  ANDN U2267 ( .B(n2018), .A(n256), .Z(n2016) );
  XNOR U2268 ( .A(a[775]), .B(n2019), .Z(n256) );
  IV U2269 ( .A(n2017), .Z(n2019) );
  XNOR U2270 ( .A(b[775]), .B(n2017), .Z(n2018) );
  XOR U2271 ( .A(n2020), .B(n2021), .Z(n2017) );
  ANDN U2272 ( .B(n2022), .A(n257), .Z(n2020) );
  XNOR U2273 ( .A(a[774]), .B(n2023), .Z(n257) );
  IV U2274 ( .A(n2021), .Z(n2023) );
  XNOR U2275 ( .A(b[774]), .B(n2021), .Z(n2022) );
  XOR U2276 ( .A(n2024), .B(n2025), .Z(n2021) );
  ANDN U2277 ( .B(n2026), .A(n258), .Z(n2024) );
  XNOR U2278 ( .A(a[773]), .B(n2027), .Z(n258) );
  IV U2279 ( .A(n2025), .Z(n2027) );
  XNOR U2280 ( .A(b[773]), .B(n2025), .Z(n2026) );
  XOR U2281 ( .A(n2028), .B(n2029), .Z(n2025) );
  ANDN U2282 ( .B(n2030), .A(n259), .Z(n2028) );
  XNOR U2283 ( .A(a[772]), .B(n2031), .Z(n259) );
  IV U2284 ( .A(n2029), .Z(n2031) );
  XNOR U2285 ( .A(b[772]), .B(n2029), .Z(n2030) );
  XOR U2286 ( .A(n2032), .B(n2033), .Z(n2029) );
  ANDN U2287 ( .B(n2034), .A(n260), .Z(n2032) );
  XNOR U2288 ( .A(a[771]), .B(n2035), .Z(n260) );
  IV U2289 ( .A(n2033), .Z(n2035) );
  XNOR U2290 ( .A(b[771]), .B(n2033), .Z(n2034) );
  XOR U2291 ( .A(n2036), .B(n2037), .Z(n2033) );
  ANDN U2292 ( .B(n2038), .A(n261), .Z(n2036) );
  XNOR U2293 ( .A(a[770]), .B(n2039), .Z(n261) );
  IV U2294 ( .A(n2037), .Z(n2039) );
  XNOR U2295 ( .A(b[770]), .B(n2037), .Z(n2038) );
  XOR U2296 ( .A(n2040), .B(n2041), .Z(n2037) );
  ANDN U2297 ( .B(n2042), .A(n263), .Z(n2040) );
  XNOR U2298 ( .A(a[769]), .B(n2043), .Z(n263) );
  IV U2299 ( .A(n2041), .Z(n2043) );
  XNOR U2300 ( .A(b[769]), .B(n2041), .Z(n2042) );
  XOR U2301 ( .A(n2044), .B(n2045), .Z(n2041) );
  ANDN U2302 ( .B(n2046), .A(n264), .Z(n2044) );
  XNOR U2303 ( .A(a[768]), .B(n2047), .Z(n264) );
  IV U2304 ( .A(n2045), .Z(n2047) );
  XNOR U2305 ( .A(b[768]), .B(n2045), .Z(n2046) );
  XOR U2306 ( .A(n2048), .B(n2049), .Z(n2045) );
  ANDN U2307 ( .B(n2050), .A(n265), .Z(n2048) );
  XNOR U2308 ( .A(a[767]), .B(n2051), .Z(n265) );
  IV U2309 ( .A(n2049), .Z(n2051) );
  XNOR U2310 ( .A(b[767]), .B(n2049), .Z(n2050) );
  XOR U2311 ( .A(n2052), .B(n2053), .Z(n2049) );
  ANDN U2312 ( .B(n2054), .A(n266), .Z(n2052) );
  XNOR U2313 ( .A(a[766]), .B(n2055), .Z(n266) );
  IV U2314 ( .A(n2053), .Z(n2055) );
  XNOR U2315 ( .A(b[766]), .B(n2053), .Z(n2054) );
  XOR U2316 ( .A(n2056), .B(n2057), .Z(n2053) );
  ANDN U2317 ( .B(n2058), .A(n267), .Z(n2056) );
  XNOR U2318 ( .A(a[765]), .B(n2059), .Z(n267) );
  IV U2319 ( .A(n2057), .Z(n2059) );
  XNOR U2320 ( .A(b[765]), .B(n2057), .Z(n2058) );
  XOR U2321 ( .A(n2060), .B(n2061), .Z(n2057) );
  ANDN U2322 ( .B(n2062), .A(n268), .Z(n2060) );
  XNOR U2323 ( .A(a[764]), .B(n2063), .Z(n268) );
  IV U2324 ( .A(n2061), .Z(n2063) );
  XNOR U2325 ( .A(b[764]), .B(n2061), .Z(n2062) );
  XOR U2326 ( .A(n2064), .B(n2065), .Z(n2061) );
  ANDN U2327 ( .B(n2066), .A(n269), .Z(n2064) );
  XNOR U2328 ( .A(a[763]), .B(n2067), .Z(n269) );
  IV U2329 ( .A(n2065), .Z(n2067) );
  XNOR U2330 ( .A(b[763]), .B(n2065), .Z(n2066) );
  XOR U2331 ( .A(n2068), .B(n2069), .Z(n2065) );
  ANDN U2332 ( .B(n2070), .A(n270), .Z(n2068) );
  XNOR U2333 ( .A(a[762]), .B(n2071), .Z(n270) );
  IV U2334 ( .A(n2069), .Z(n2071) );
  XNOR U2335 ( .A(b[762]), .B(n2069), .Z(n2070) );
  XOR U2336 ( .A(n2072), .B(n2073), .Z(n2069) );
  ANDN U2337 ( .B(n2074), .A(n271), .Z(n2072) );
  XNOR U2338 ( .A(a[761]), .B(n2075), .Z(n271) );
  IV U2339 ( .A(n2073), .Z(n2075) );
  XNOR U2340 ( .A(b[761]), .B(n2073), .Z(n2074) );
  XOR U2341 ( .A(n2076), .B(n2077), .Z(n2073) );
  ANDN U2342 ( .B(n2078), .A(n272), .Z(n2076) );
  XNOR U2343 ( .A(a[760]), .B(n2079), .Z(n272) );
  IV U2344 ( .A(n2077), .Z(n2079) );
  XNOR U2345 ( .A(b[760]), .B(n2077), .Z(n2078) );
  XOR U2346 ( .A(n2080), .B(n2081), .Z(n2077) );
  ANDN U2347 ( .B(n2082), .A(n274), .Z(n2080) );
  XNOR U2348 ( .A(a[759]), .B(n2083), .Z(n274) );
  IV U2349 ( .A(n2081), .Z(n2083) );
  XNOR U2350 ( .A(b[759]), .B(n2081), .Z(n2082) );
  XOR U2351 ( .A(n2084), .B(n2085), .Z(n2081) );
  ANDN U2352 ( .B(n2086), .A(n275), .Z(n2084) );
  XNOR U2353 ( .A(a[758]), .B(n2087), .Z(n275) );
  IV U2354 ( .A(n2085), .Z(n2087) );
  XNOR U2355 ( .A(b[758]), .B(n2085), .Z(n2086) );
  XOR U2356 ( .A(n2088), .B(n2089), .Z(n2085) );
  ANDN U2357 ( .B(n2090), .A(n276), .Z(n2088) );
  XNOR U2358 ( .A(a[757]), .B(n2091), .Z(n276) );
  IV U2359 ( .A(n2089), .Z(n2091) );
  XNOR U2360 ( .A(b[757]), .B(n2089), .Z(n2090) );
  XOR U2361 ( .A(n2092), .B(n2093), .Z(n2089) );
  ANDN U2362 ( .B(n2094), .A(n277), .Z(n2092) );
  XNOR U2363 ( .A(a[756]), .B(n2095), .Z(n277) );
  IV U2364 ( .A(n2093), .Z(n2095) );
  XNOR U2365 ( .A(b[756]), .B(n2093), .Z(n2094) );
  XOR U2366 ( .A(n2096), .B(n2097), .Z(n2093) );
  ANDN U2367 ( .B(n2098), .A(n278), .Z(n2096) );
  XNOR U2368 ( .A(a[755]), .B(n2099), .Z(n278) );
  IV U2369 ( .A(n2097), .Z(n2099) );
  XNOR U2370 ( .A(b[755]), .B(n2097), .Z(n2098) );
  XOR U2371 ( .A(n2100), .B(n2101), .Z(n2097) );
  ANDN U2372 ( .B(n2102), .A(n279), .Z(n2100) );
  XNOR U2373 ( .A(a[754]), .B(n2103), .Z(n279) );
  IV U2374 ( .A(n2101), .Z(n2103) );
  XNOR U2375 ( .A(b[754]), .B(n2101), .Z(n2102) );
  XOR U2376 ( .A(n2104), .B(n2105), .Z(n2101) );
  ANDN U2377 ( .B(n2106), .A(n280), .Z(n2104) );
  XNOR U2378 ( .A(a[753]), .B(n2107), .Z(n280) );
  IV U2379 ( .A(n2105), .Z(n2107) );
  XNOR U2380 ( .A(b[753]), .B(n2105), .Z(n2106) );
  XOR U2381 ( .A(n2108), .B(n2109), .Z(n2105) );
  ANDN U2382 ( .B(n2110), .A(n281), .Z(n2108) );
  XNOR U2383 ( .A(a[752]), .B(n2111), .Z(n281) );
  IV U2384 ( .A(n2109), .Z(n2111) );
  XNOR U2385 ( .A(b[752]), .B(n2109), .Z(n2110) );
  XOR U2386 ( .A(n2112), .B(n2113), .Z(n2109) );
  ANDN U2387 ( .B(n2114), .A(n282), .Z(n2112) );
  XNOR U2388 ( .A(a[751]), .B(n2115), .Z(n282) );
  IV U2389 ( .A(n2113), .Z(n2115) );
  XNOR U2390 ( .A(b[751]), .B(n2113), .Z(n2114) );
  XOR U2391 ( .A(n2116), .B(n2117), .Z(n2113) );
  ANDN U2392 ( .B(n2118), .A(n283), .Z(n2116) );
  XNOR U2393 ( .A(a[750]), .B(n2119), .Z(n283) );
  IV U2394 ( .A(n2117), .Z(n2119) );
  XNOR U2395 ( .A(b[750]), .B(n2117), .Z(n2118) );
  XOR U2396 ( .A(n2120), .B(n2121), .Z(n2117) );
  ANDN U2397 ( .B(n2122), .A(n285), .Z(n2120) );
  XNOR U2398 ( .A(a[749]), .B(n2123), .Z(n285) );
  IV U2399 ( .A(n2121), .Z(n2123) );
  XNOR U2400 ( .A(b[749]), .B(n2121), .Z(n2122) );
  XOR U2401 ( .A(n2124), .B(n2125), .Z(n2121) );
  ANDN U2402 ( .B(n2126), .A(n286), .Z(n2124) );
  XNOR U2403 ( .A(a[748]), .B(n2127), .Z(n286) );
  IV U2404 ( .A(n2125), .Z(n2127) );
  XNOR U2405 ( .A(b[748]), .B(n2125), .Z(n2126) );
  XOR U2406 ( .A(n2128), .B(n2129), .Z(n2125) );
  ANDN U2407 ( .B(n2130), .A(n287), .Z(n2128) );
  XNOR U2408 ( .A(a[747]), .B(n2131), .Z(n287) );
  IV U2409 ( .A(n2129), .Z(n2131) );
  XNOR U2410 ( .A(b[747]), .B(n2129), .Z(n2130) );
  XOR U2411 ( .A(n2132), .B(n2133), .Z(n2129) );
  ANDN U2412 ( .B(n2134), .A(n288), .Z(n2132) );
  XNOR U2413 ( .A(a[746]), .B(n2135), .Z(n288) );
  IV U2414 ( .A(n2133), .Z(n2135) );
  XNOR U2415 ( .A(b[746]), .B(n2133), .Z(n2134) );
  XOR U2416 ( .A(n2136), .B(n2137), .Z(n2133) );
  ANDN U2417 ( .B(n2138), .A(n289), .Z(n2136) );
  XNOR U2418 ( .A(a[745]), .B(n2139), .Z(n289) );
  IV U2419 ( .A(n2137), .Z(n2139) );
  XNOR U2420 ( .A(b[745]), .B(n2137), .Z(n2138) );
  XOR U2421 ( .A(n2140), .B(n2141), .Z(n2137) );
  ANDN U2422 ( .B(n2142), .A(n290), .Z(n2140) );
  XNOR U2423 ( .A(a[744]), .B(n2143), .Z(n290) );
  IV U2424 ( .A(n2141), .Z(n2143) );
  XNOR U2425 ( .A(b[744]), .B(n2141), .Z(n2142) );
  XOR U2426 ( .A(n2144), .B(n2145), .Z(n2141) );
  ANDN U2427 ( .B(n2146), .A(n291), .Z(n2144) );
  XNOR U2428 ( .A(a[743]), .B(n2147), .Z(n291) );
  IV U2429 ( .A(n2145), .Z(n2147) );
  XNOR U2430 ( .A(b[743]), .B(n2145), .Z(n2146) );
  XOR U2431 ( .A(n2148), .B(n2149), .Z(n2145) );
  ANDN U2432 ( .B(n2150), .A(n292), .Z(n2148) );
  XNOR U2433 ( .A(a[742]), .B(n2151), .Z(n292) );
  IV U2434 ( .A(n2149), .Z(n2151) );
  XNOR U2435 ( .A(b[742]), .B(n2149), .Z(n2150) );
  XOR U2436 ( .A(n2152), .B(n2153), .Z(n2149) );
  ANDN U2437 ( .B(n2154), .A(n293), .Z(n2152) );
  XNOR U2438 ( .A(a[741]), .B(n2155), .Z(n293) );
  IV U2439 ( .A(n2153), .Z(n2155) );
  XNOR U2440 ( .A(b[741]), .B(n2153), .Z(n2154) );
  XOR U2441 ( .A(n2156), .B(n2157), .Z(n2153) );
  ANDN U2442 ( .B(n2158), .A(n294), .Z(n2156) );
  XNOR U2443 ( .A(a[740]), .B(n2159), .Z(n294) );
  IV U2444 ( .A(n2157), .Z(n2159) );
  XNOR U2445 ( .A(b[740]), .B(n2157), .Z(n2158) );
  XOR U2446 ( .A(n2160), .B(n2161), .Z(n2157) );
  ANDN U2447 ( .B(n2162), .A(n296), .Z(n2160) );
  XNOR U2448 ( .A(a[739]), .B(n2163), .Z(n296) );
  IV U2449 ( .A(n2161), .Z(n2163) );
  XNOR U2450 ( .A(b[739]), .B(n2161), .Z(n2162) );
  XOR U2451 ( .A(n2164), .B(n2165), .Z(n2161) );
  ANDN U2452 ( .B(n2166), .A(n297), .Z(n2164) );
  XNOR U2453 ( .A(a[738]), .B(n2167), .Z(n297) );
  IV U2454 ( .A(n2165), .Z(n2167) );
  XNOR U2455 ( .A(b[738]), .B(n2165), .Z(n2166) );
  XOR U2456 ( .A(n2168), .B(n2169), .Z(n2165) );
  ANDN U2457 ( .B(n2170), .A(n298), .Z(n2168) );
  XNOR U2458 ( .A(a[737]), .B(n2171), .Z(n298) );
  IV U2459 ( .A(n2169), .Z(n2171) );
  XNOR U2460 ( .A(b[737]), .B(n2169), .Z(n2170) );
  XOR U2461 ( .A(n2172), .B(n2173), .Z(n2169) );
  ANDN U2462 ( .B(n2174), .A(n299), .Z(n2172) );
  XNOR U2463 ( .A(a[736]), .B(n2175), .Z(n299) );
  IV U2464 ( .A(n2173), .Z(n2175) );
  XNOR U2465 ( .A(b[736]), .B(n2173), .Z(n2174) );
  XOR U2466 ( .A(n2176), .B(n2177), .Z(n2173) );
  ANDN U2467 ( .B(n2178), .A(n300), .Z(n2176) );
  XNOR U2468 ( .A(a[735]), .B(n2179), .Z(n300) );
  IV U2469 ( .A(n2177), .Z(n2179) );
  XNOR U2470 ( .A(b[735]), .B(n2177), .Z(n2178) );
  XOR U2471 ( .A(n2180), .B(n2181), .Z(n2177) );
  ANDN U2472 ( .B(n2182), .A(n301), .Z(n2180) );
  XNOR U2473 ( .A(a[734]), .B(n2183), .Z(n301) );
  IV U2474 ( .A(n2181), .Z(n2183) );
  XNOR U2475 ( .A(b[734]), .B(n2181), .Z(n2182) );
  XOR U2476 ( .A(n2184), .B(n2185), .Z(n2181) );
  ANDN U2477 ( .B(n2186), .A(n302), .Z(n2184) );
  XNOR U2478 ( .A(a[733]), .B(n2187), .Z(n302) );
  IV U2479 ( .A(n2185), .Z(n2187) );
  XNOR U2480 ( .A(b[733]), .B(n2185), .Z(n2186) );
  XOR U2481 ( .A(n2188), .B(n2189), .Z(n2185) );
  ANDN U2482 ( .B(n2190), .A(n303), .Z(n2188) );
  XNOR U2483 ( .A(a[732]), .B(n2191), .Z(n303) );
  IV U2484 ( .A(n2189), .Z(n2191) );
  XNOR U2485 ( .A(b[732]), .B(n2189), .Z(n2190) );
  XOR U2486 ( .A(n2192), .B(n2193), .Z(n2189) );
  ANDN U2487 ( .B(n2194), .A(n304), .Z(n2192) );
  XNOR U2488 ( .A(a[731]), .B(n2195), .Z(n304) );
  IV U2489 ( .A(n2193), .Z(n2195) );
  XNOR U2490 ( .A(b[731]), .B(n2193), .Z(n2194) );
  XOR U2491 ( .A(n2196), .B(n2197), .Z(n2193) );
  ANDN U2492 ( .B(n2198), .A(n305), .Z(n2196) );
  XNOR U2493 ( .A(a[730]), .B(n2199), .Z(n305) );
  IV U2494 ( .A(n2197), .Z(n2199) );
  XNOR U2495 ( .A(b[730]), .B(n2197), .Z(n2198) );
  XOR U2496 ( .A(n2200), .B(n2201), .Z(n2197) );
  ANDN U2497 ( .B(n2202), .A(n307), .Z(n2200) );
  XNOR U2498 ( .A(a[729]), .B(n2203), .Z(n307) );
  IV U2499 ( .A(n2201), .Z(n2203) );
  XNOR U2500 ( .A(b[729]), .B(n2201), .Z(n2202) );
  XOR U2501 ( .A(n2204), .B(n2205), .Z(n2201) );
  ANDN U2502 ( .B(n2206), .A(n308), .Z(n2204) );
  XNOR U2503 ( .A(a[728]), .B(n2207), .Z(n308) );
  IV U2504 ( .A(n2205), .Z(n2207) );
  XNOR U2505 ( .A(b[728]), .B(n2205), .Z(n2206) );
  XOR U2506 ( .A(n2208), .B(n2209), .Z(n2205) );
  ANDN U2507 ( .B(n2210), .A(n309), .Z(n2208) );
  XNOR U2508 ( .A(a[727]), .B(n2211), .Z(n309) );
  IV U2509 ( .A(n2209), .Z(n2211) );
  XNOR U2510 ( .A(b[727]), .B(n2209), .Z(n2210) );
  XOR U2511 ( .A(n2212), .B(n2213), .Z(n2209) );
  ANDN U2512 ( .B(n2214), .A(n310), .Z(n2212) );
  XNOR U2513 ( .A(a[726]), .B(n2215), .Z(n310) );
  IV U2514 ( .A(n2213), .Z(n2215) );
  XNOR U2515 ( .A(b[726]), .B(n2213), .Z(n2214) );
  XOR U2516 ( .A(n2216), .B(n2217), .Z(n2213) );
  ANDN U2517 ( .B(n2218), .A(n311), .Z(n2216) );
  XNOR U2518 ( .A(a[725]), .B(n2219), .Z(n311) );
  IV U2519 ( .A(n2217), .Z(n2219) );
  XNOR U2520 ( .A(b[725]), .B(n2217), .Z(n2218) );
  XOR U2521 ( .A(n2220), .B(n2221), .Z(n2217) );
  ANDN U2522 ( .B(n2222), .A(n312), .Z(n2220) );
  XNOR U2523 ( .A(a[724]), .B(n2223), .Z(n312) );
  IV U2524 ( .A(n2221), .Z(n2223) );
  XNOR U2525 ( .A(b[724]), .B(n2221), .Z(n2222) );
  XOR U2526 ( .A(n2224), .B(n2225), .Z(n2221) );
  ANDN U2527 ( .B(n2226), .A(n313), .Z(n2224) );
  XNOR U2528 ( .A(a[723]), .B(n2227), .Z(n313) );
  IV U2529 ( .A(n2225), .Z(n2227) );
  XNOR U2530 ( .A(b[723]), .B(n2225), .Z(n2226) );
  XOR U2531 ( .A(n2228), .B(n2229), .Z(n2225) );
  ANDN U2532 ( .B(n2230), .A(n314), .Z(n2228) );
  XNOR U2533 ( .A(a[722]), .B(n2231), .Z(n314) );
  IV U2534 ( .A(n2229), .Z(n2231) );
  XNOR U2535 ( .A(b[722]), .B(n2229), .Z(n2230) );
  XOR U2536 ( .A(n2232), .B(n2233), .Z(n2229) );
  ANDN U2537 ( .B(n2234), .A(n315), .Z(n2232) );
  XNOR U2538 ( .A(a[721]), .B(n2235), .Z(n315) );
  IV U2539 ( .A(n2233), .Z(n2235) );
  XNOR U2540 ( .A(b[721]), .B(n2233), .Z(n2234) );
  XOR U2541 ( .A(n2236), .B(n2237), .Z(n2233) );
  ANDN U2542 ( .B(n2238), .A(n316), .Z(n2236) );
  XNOR U2543 ( .A(a[720]), .B(n2239), .Z(n316) );
  IV U2544 ( .A(n2237), .Z(n2239) );
  XNOR U2545 ( .A(b[720]), .B(n2237), .Z(n2238) );
  XOR U2546 ( .A(n2240), .B(n2241), .Z(n2237) );
  ANDN U2547 ( .B(n2242), .A(n318), .Z(n2240) );
  XNOR U2548 ( .A(a[719]), .B(n2243), .Z(n318) );
  IV U2549 ( .A(n2241), .Z(n2243) );
  XNOR U2550 ( .A(b[719]), .B(n2241), .Z(n2242) );
  XOR U2551 ( .A(n2244), .B(n2245), .Z(n2241) );
  ANDN U2552 ( .B(n2246), .A(n319), .Z(n2244) );
  XNOR U2553 ( .A(a[718]), .B(n2247), .Z(n319) );
  IV U2554 ( .A(n2245), .Z(n2247) );
  XNOR U2555 ( .A(b[718]), .B(n2245), .Z(n2246) );
  XOR U2556 ( .A(n2248), .B(n2249), .Z(n2245) );
  ANDN U2557 ( .B(n2250), .A(n320), .Z(n2248) );
  XNOR U2558 ( .A(a[717]), .B(n2251), .Z(n320) );
  IV U2559 ( .A(n2249), .Z(n2251) );
  XNOR U2560 ( .A(b[717]), .B(n2249), .Z(n2250) );
  XOR U2561 ( .A(n2252), .B(n2253), .Z(n2249) );
  ANDN U2562 ( .B(n2254), .A(n321), .Z(n2252) );
  XNOR U2563 ( .A(a[716]), .B(n2255), .Z(n321) );
  IV U2564 ( .A(n2253), .Z(n2255) );
  XNOR U2565 ( .A(b[716]), .B(n2253), .Z(n2254) );
  XOR U2566 ( .A(n2256), .B(n2257), .Z(n2253) );
  ANDN U2567 ( .B(n2258), .A(n322), .Z(n2256) );
  XNOR U2568 ( .A(a[715]), .B(n2259), .Z(n322) );
  IV U2569 ( .A(n2257), .Z(n2259) );
  XNOR U2570 ( .A(b[715]), .B(n2257), .Z(n2258) );
  XOR U2571 ( .A(n2260), .B(n2261), .Z(n2257) );
  ANDN U2572 ( .B(n2262), .A(n323), .Z(n2260) );
  XNOR U2573 ( .A(a[714]), .B(n2263), .Z(n323) );
  IV U2574 ( .A(n2261), .Z(n2263) );
  XNOR U2575 ( .A(b[714]), .B(n2261), .Z(n2262) );
  XOR U2576 ( .A(n2264), .B(n2265), .Z(n2261) );
  ANDN U2577 ( .B(n2266), .A(n324), .Z(n2264) );
  XNOR U2578 ( .A(a[713]), .B(n2267), .Z(n324) );
  IV U2579 ( .A(n2265), .Z(n2267) );
  XNOR U2580 ( .A(b[713]), .B(n2265), .Z(n2266) );
  XOR U2581 ( .A(n2268), .B(n2269), .Z(n2265) );
  ANDN U2582 ( .B(n2270), .A(n325), .Z(n2268) );
  XNOR U2583 ( .A(a[712]), .B(n2271), .Z(n325) );
  IV U2584 ( .A(n2269), .Z(n2271) );
  XNOR U2585 ( .A(b[712]), .B(n2269), .Z(n2270) );
  XOR U2586 ( .A(n2272), .B(n2273), .Z(n2269) );
  ANDN U2587 ( .B(n2274), .A(n326), .Z(n2272) );
  XNOR U2588 ( .A(a[711]), .B(n2275), .Z(n326) );
  IV U2589 ( .A(n2273), .Z(n2275) );
  XNOR U2590 ( .A(b[711]), .B(n2273), .Z(n2274) );
  XOR U2591 ( .A(n2276), .B(n2277), .Z(n2273) );
  ANDN U2592 ( .B(n2278), .A(n327), .Z(n2276) );
  XNOR U2593 ( .A(a[710]), .B(n2279), .Z(n327) );
  IV U2594 ( .A(n2277), .Z(n2279) );
  XNOR U2595 ( .A(b[710]), .B(n2277), .Z(n2278) );
  XOR U2596 ( .A(n2280), .B(n2281), .Z(n2277) );
  ANDN U2597 ( .B(n2282), .A(n329), .Z(n2280) );
  XNOR U2598 ( .A(a[709]), .B(n2283), .Z(n329) );
  IV U2599 ( .A(n2281), .Z(n2283) );
  XNOR U2600 ( .A(b[709]), .B(n2281), .Z(n2282) );
  XOR U2601 ( .A(n2284), .B(n2285), .Z(n2281) );
  ANDN U2602 ( .B(n2286), .A(n330), .Z(n2284) );
  XNOR U2603 ( .A(a[708]), .B(n2287), .Z(n330) );
  IV U2604 ( .A(n2285), .Z(n2287) );
  XNOR U2605 ( .A(b[708]), .B(n2285), .Z(n2286) );
  XOR U2606 ( .A(n2288), .B(n2289), .Z(n2285) );
  ANDN U2607 ( .B(n2290), .A(n331), .Z(n2288) );
  XNOR U2608 ( .A(a[707]), .B(n2291), .Z(n331) );
  IV U2609 ( .A(n2289), .Z(n2291) );
  XNOR U2610 ( .A(b[707]), .B(n2289), .Z(n2290) );
  XOR U2611 ( .A(n2292), .B(n2293), .Z(n2289) );
  ANDN U2612 ( .B(n2294), .A(n332), .Z(n2292) );
  XNOR U2613 ( .A(a[706]), .B(n2295), .Z(n332) );
  IV U2614 ( .A(n2293), .Z(n2295) );
  XNOR U2615 ( .A(b[706]), .B(n2293), .Z(n2294) );
  XOR U2616 ( .A(n2296), .B(n2297), .Z(n2293) );
  ANDN U2617 ( .B(n2298), .A(n333), .Z(n2296) );
  XNOR U2618 ( .A(a[705]), .B(n2299), .Z(n333) );
  IV U2619 ( .A(n2297), .Z(n2299) );
  XNOR U2620 ( .A(b[705]), .B(n2297), .Z(n2298) );
  XOR U2621 ( .A(n2300), .B(n2301), .Z(n2297) );
  ANDN U2622 ( .B(n2302), .A(n334), .Z(n2300) );
  XNOR U2623 ( .A(a[704]), .B(n2303), .Z(n334) );
  IV U2624 ( .A(n2301), .Z(n2303) );
  XNOR U2625 ( .A(b[704]), .B(n2301), .Z(n2302) );
  XOR U2626 ( .A(n2304), .B(n2305), .Z(n2301) );
  ANDN U2627 ( .B(n2306), .A(n335), .Z(n2304) );
  XNOR U2628 ( .A(a[703]), .B(n2307), .Z(n335) );
  IV U2629 ( .A(n2305), .Z(n2307) );
  XNOR U2630 ( .A(b[703]), .B(n2305), .Z(n2306) );
  XOR U2631 ( .A(n2308), .B(n2309), .Z(n2305) );
  ANDN U2632 ( .B(n2310), .A(n336), .Z(n2308) );
  XNOR U2633 ( .A(a[702]), .B(n2311), .Z(n336) );
  IV U2634 ( .A(n2309), .Z(n2311) );
  XNOR U2635 ( .A(b[702]), .B(n2309), .Z(n2310) );
  XOR U2636 ( .A(n2312), .B(n2313), .Z(n2309) );
  ANDN U2637 ( .B(n2314), .A(n337), .Z(n2312) );
  XNOR U2638 ( .A(a[701]), .B(n2315), .Z(n337) );
  IV U2639 ( .A(n2313), .Z(n2315) );
  XNOR U2640 ( .A(b[701]), .B(n2313), .Z(n2314) );
  XOR U2641 ( .A(n2316), .B(n2317), .Z(n2313) );
  ANDN U2642 ( .B(n2318), .A(n338), .Z(n2316) );
  XNOR U2643 ( .A(a[700]), .B(n2319), .Z(n338) );
  IV U2644 ( .A(n2317), .Z(n2319) );
  XNOR U2645 ( .A(b[700]), .B(n2317), .Z(n2318) );
  XOR U2646 ( .A(n2320), .B(n2321), .Z(n2317) );
  ANDN U2647 ( .B(n2322), .A(n341), .Z(n2320) );
  XNOR U2648 ( .A(a[699]), .B(n2323), .Z(n341) );
  IV U2649 ( .A(n2321), .Z(n2323) );
  XNOR U2650 ( .A(b[699]), .B(n2321), .Z(n2322) );
  XOR U2651 ( .A(n2324), .B(n2325), .Z(n2321) );
  ANDN U2652 ( .B(n2326), .A(n342), .Z(n2324) );
  XNOR U2653 ( .A(a[698]), .B(n2327), .Z(n342) );
  IV U2654 ( .A(n2325), .Z(n2327) );
  XNOR U2655 ( .A(b[698]), .B(n2325), .Z(n2326) );
  XOR U2656 ( .A(n2328), .B(n2329), .Z(n2325) );
  ANDN U2657 ( .B(n2330), .A(n343), .Z(n2328) );
  XNOR U2658 ( .A(a[697]), .B(n2331), .Z(n343) );
  IV U2659 ( .A(n2329), .Z(n2331) );
  XNOR U2660 ( .A(b[697]), .B(n2329), .Z(n2330) );
  XOR U2661 ( .A(n2332), .B(n2333), .Z(n2329) );
  ANDN U2662 ( .B(n2334), .A(n344), .Z(n2332) );
  XNOR U2663 ( .A(a[696]), .B(n2335), .Z(n344) );
  IV U2664 ( .A(n2333), .Z(n2335) );
  XNOR U2665 ( .A(b[696]), .B(n2333), .Z(n2334) );
  XOR U2666 ( .A(n2336), .B(n2337), .Z(n2333) );
  ANDN U2667 ( .B(n2338), .A(n345), .Z(n2336) );
  XNOR U2668 ( .A(a[695]), .B(n2339), .Z(n345) );
  IV U2669 ( .A(n2337), .Z(n2339) );
  XNOR U2670 ( .A(b[695]), .B(n2337), .Z(n2338) );
  XOR U2671 ( .A(n2340), .B(n2341), .Z(n2337) );
  ANDN U2672 ( .B(n2342), .A(n346), .Z(n2340) );
  XNOR U2673 ( .A(a[694]), .B(n2343), .Z(n346) );
  IV U2674 ( .A(n2341), .Z(n2343) );
  XNOR U2675 ( .A(b[694]), .B(n2341), .Z(n2342) );
  XOR U2676 ( .A(n2344), .B(n2345), .Z(n2341) );
  ANDN U2677 ( .B(n2346), .A(n347), .Z(n2344) );
  XNOR U2678 ( .A(a[693]), .B(n2347), .Z(n347) );
  IV U2679 ( .A(n2345), .Z(n2347) );
  XNOR U2680 ( .A(b[693]), .B(n2345), .Z(n2346) );
  XOR U2681 ( .A(n2348), .B(n2349), .Z(n2345) );
  ANDN U2682 ( .B(n2350), .A(n348), .Z(n2348) );
  XNOR U2683 ( .A(a[692]), .B(n2351), .Z(n348) );
  IV U2684 ( .A(n2349), .Z(n2351) );
  XNOR U2685 ( .A(b[692]), .B(n2349), .Z(n2350) );
  XOR U2686 ( .A(n2352), .B(n2353), .Z(n2349) );
  ANDN U2687 ( .B(n2354), .A(n349), .Z(n2352) );
  XNOR U2688 ( .A(a[691]), .B(n2355), .Z(n349) );
  IV U2689 ( .A(n2353), .Z(n2355) );
  XNOR U2690 ( .A(b[691]), .B(n2353), .Z(n2354) );
  XOR U2691 ( .A(n2356), .B(n2357), .Z(n2353) );
  ANDN U2692 ( .B(n2358), .A(n350), .Z(n2356) );
  XNOR U2693 ( .A(a[690]), .B(n2359), .Z(n350) );
  IV U2694 ( .A(n2357), .Z(n2359) );
  XNOR U2695 ( .A(b[690]), .B(n2357), .Z(n2358) );
  XOR U2696 ( .A(n2360), .B(n2361), .Z(n2357) );
  ANDN U2697 ( .B(n2362), .A(n352), .Z(n2360) );
  XNOR U2698 ( .A(a[689]), .B(n2363), .Z(n352) );
  IV U2699 ( .A(n2361), .Z(n2363) );
  XNOR U2700 ( .A(b[689]), .B(n2361), .Z(n2362) );
  XOR U2701 ( .A(n2364), .B(n2365), .Z(n2361) );
  ANDN U2702 ( .B(n2366), .A(n353), .Z(n2364) );
  XNOR U2703 ( .A(a[688]), .B(n2367), .Z(n353) );
  IV U2704 ( .A(n2365), .Z(n2367) );
  XNOR U2705 ( .A(b[688]), .B(n2365), .Z(n2366) );
  XOR U2706 ( .A(n2368), .B(n2369), .Z(n2365) );
  ANDN U2707 ( .B(n2370), .A(n354), .Z(n2368) );
  XNOR U2708 ( .A(a[687]), .B(n2371), .Z(n354) );
  IV U2709 ( .A(n2369), .Z(n2371) );
  XNOR U2710 ( .A(b[687]), .B(n2369), .Z(n2370) );
  XOR U2711 ( .A(n2372), .B(n2373), .Z(n2369) );
  ANDN U2712 ( .B(n2374), .A(n355), .Z(n2372) );
  XNOR U2713 ( .A(a[686]), .B(n2375), .Z(n355) );
  IV U2714 ( .A(n2373), .Z(n2375) );
  XNOR U2715 ( .A(b[686]), .B(n2373), .Z(n2374) );
  XOR U2716 ( .A(n2376), .B(n2377), .Z(n2373) );
  ANDN U2717 ( .B(n2378), .A(n356), .Z(n2376) );
  XNOR U2718 ( .A(a[685]), .B(n2379), .Z(n356) );
  IV U2719 ( .A(n2377), .Z(n2379) );
  XNOR U2720 ( .A(b[685]), .B(n2377), .Z(n2378) );
  XOR U2721 ( .A(n2380), .B(n2381), .Z(n2377) );
  ANDN U2722 ( .B(n2382), .A(n357), .Z(n2380) );
  XNOR U2723 ( .A(a[684]), .B(n2383), .Z(n357) );
  IV U2724 ( .A(n2381), .Z(n2383) );
  XNOR U2725 ( .A(b[684]), .B(n2381), .Z(n2382) );
  XOR U2726 ( .A(n2384), .B(n2385), .Z(n2381) );
  ANDN U2727 ( .B(n2386), .A(n358), .Z(n2384) );
  XNOR U2728 ( .A(a[683]), .B(n2387), .Z(n358) );
  IV U2729 ( .A(n2385), .Z(n2387) );
  XNOR U2730 ( .A(b[683]), .B(n2385), .Z(n2386) );
  XOR U2731 ( .A(n2388), .B(n2389), .Z(n2385) );
  ANDN U2732 ( .B(n2390), .A(n359), .Z(n2388) );
  XNOR U2733 ( .A(a[682]), .B(n2391), .Z(n359) );
  IV U2734 ( .A(n2389), .Z(n2391) );
  XNOR U2735 ( .A(b[682]), .B(n2389), .Z(n2390) );
  XOR U2736 ( .A(n2392), .B(n2393), .Z(n2389) );
  ANDN U2737 ( .B(n2394), .A(n360), .Z(n2392) );
  XNOR U2738 ( .A(a[681]), .B(n2395), .Z(n360) );
  IV U2739 ( .A(n2393), .Z(n2395) );
  XNOR U2740 ( .A(b[681]), .B(n2393), .Z(n2394) );
  XOR U2741 ( .A(n2396), .B(n2397), .Z(n2393) );
  ANDN U2742 ( .B(n2398), .A(n361), .Z(n2396) );
  XNOR U2743 ( .A(a[680]), .B(n2399), .Z(n361) );
  IV U2744 ( .A(n2397), .Z(n2399) );
  XNOR U2745 ( .A(b[680]), .B(n2397), .Z(n2398) );
  XOR U2746 ( .A(n2400), .B(n2401), .Z(n2397) );
  ANDN U2747 ( .B(n2402), .A(n363), .Z(n2400) );
  XNOR U2748 ( .A(a[679]), .B(n2403), .Z(n363) );
  IV U2749 ( .A(n2401), .Z(n2403) );
  XNOR U2750 ( .A(b[679]), .B(n2401), .Z(n2402) );
  XOR U2751 ( .A(n2404), .B(n2405), .Z(n2401) );
  ANDN U2752 ( .B(n2406), .A(n364), .Z(n2404) );
  XNOR U2753 ( .A(a[678]), .B(n2407), .Z(n364) );
  IV U2754 ( .A(n2405), .Z(n2407) );
  XNOR U2755 ( .A(b[678]), .B(n2405), .Z(n2406) );
  XOR U2756 ( .A(n2408), .B(n2409), .Z(n2405) );
  ANDN U2757 ( .B(n2410), .A(n365), .Z(n2408) );
  XNOR U2758 ( .A(a[677]), .B(n2411), .Z(n365) );
  IV U2759 ( .A(n2409), .Z(n2411) );
  XNOR U2760 ( .A(b[677]), .B(n2409), .Z(n2410) );
  XOR U2761 ( .A(n2412), .B(n2413), .Z(n2409) );
  ANDN U2762 ( .B(n2414), .A(n366), .Z(n2412) );
  XNOR U2763 ( .A(a[676]), .B(n2415), .Z(n366) );
  IV U2764 ( .A(n2413), .Z(n2415) );
  XNOR U2765 ( .A(b[676]), .B(n2413), .Z(n2414) );
  XOR U2766 ( .A(n2416), .B(n2417), .Z(n2413) );
  ANDN U2767 ( .B(n2418), .A(n367), .Z(n2416) );
  XNOR U2768 ( .A(a[675]), .B(n2419), .Z(n367) );
  IV U2769 ( .A(n2417), .Z(n2419) );
  XNOR U2770 ( .A(b[675]), .B(n2417), .Z(n2418) );
  XOR U2771 ( .A(n2420), .B(n2421), .Z(n2417) );
  ANDN U2772 ( .B(n2422), .A(n368), .Z(n2420) );
  XNOR U2773 ( .A(a[674]), .B(n2423), .Z(n368) );
  IV U2774 ( .A(n2421), .Z(n2423) );
  XNOR U2775 ( .A(b[674]), .B(n2421), .Z(n2422) );
  XOR U2776 ( .A(n2424), .B(n2425), .Z(n2421) );
  ANDN U2777 ( .B(n2426), .A(n369), .Z(n2424) );
  XNOR U2778 ( .A(a[673]), .B(n2427), .Z(n369) );
  IV U2779 ( .A(n2425), .Z(n2427) );
  XNOR U2780 ( .A(b[673]), .B(n2425), .Z(n2426) );
  XOR U2781 ( .A(n2428), .B(n2429), .Z(n2425) );
  ANDN U2782 ( .B(n2430), .A(n370), .Z(n2428) );
  XNOR U2783 ( .A(a[672]), .B(n2431), .Z(n370) );
  IV U2784 ( .A(n2429), .Z(n2431) );
  XNOR U2785 ( .A(b[672]), .B(n2429), .Z(n2430) );
  XOR U2786 ( .A(n2432), .B(n2433), .Z(n2429) );
  ANDN U2787 ( .B(n2434), .A(n371), .Z(n2432) );
  XNOR U2788 ( .A(a[671]), .B(n2435), .Z(n371) );
  IV U2789 ( .A(n2433), .Z(n2435) );
  XNOR U2790 ( .A(b[671]), .B(n2433), .Z(n2434) );
  XOR U2791 ( .A(n2436), .B(n2437), .Z(n2433) );
  ANDN U2792 ( .B(n2438), .A(n372), .Z(n2436) );
  XNOR U2793 ( .A(a[670]), .B(n2439), .Z(n372) );
  IV U2794 ( .A(n2437), .Z(n2439) );
  XNOR U2795 ( .A(b[670]), .B(n2437), .Z(n2438) );
  XOR U2796 ( .A(n2440), .B(n2441), .Z(n2437) );
  ANDN U2797 ( .B(n2442), .A(n374), .Z(n2440) );
  XNOR U2798 ( .A(a[669]), .B(n2443), .Z(n374) );
  IV U2799 ( .A(n2441), .Z(n2443) );
  XNOR U2800 ( .A(b[669]), .B(n2441), .Z(n2442) );
  XOR U2801 ( .A(n2444), .B(n2445), .Z(n2441) );
  ANDN U2802 ( .B(n2446), .A(n375), .Z(n2444) );
  XNOR U2803 ( .A(a[668]), .B(n2447), .Z(n375) );
  IV U2804 ( .A(n2445), .Z(n2447) );
  XNOR U2805 ( .A(b[668]), .B(n2445), .Z(n2446) );
  XOR U2806 ( .A(n2448), .B(n2449), .Z(n2445) );
  ANDN U2807 ( .B(n2450), .A(n376), .Z(n2448) );
  XNOR U2808 ( .A(a[667]), .B(n2451), .Z(n376) );
  IV U2809 ( .A(n2449), .Z(n2451) );
  XNOR U2810 ( .A(b[667]), .B(n2449), .Z(n2450) );
  XOR U2811 ( .A(n2452), .B(n2453), .Z(n2449) );
  ANDN U2812 ( .B(n2454), .A(n377), .Z(n2452) );
  XNOR U2813 ( .A(a[666]), .B(n2455), .Z(n377) );
  IV U2814 ( .A(n2453), .Z(n2455) );
  XNOR U2815 ( .A(b[666]), .B(n2453), .Z(n2454) );
  XOR U2816 ( .A(n2456), .B(n2457), .Z(n2453) );
  ANDN U2817 ( .B(n2458), .A(n378), .Z(n2456) );
  XNOR U2818 ( .A(a[665]), .B(n2459), .Z(n378) );
  IV U2819 ( .A(n2457), .Z(n2459) );
  XNOR U2820 ( .A(b[665]), .B(n2457), .Z(n2458) );
  XOR U2821 ( .A(n2460), .B(n2461), .Z(n2457) );
  ANDN U2822 ( .B(n2462), .A(n379), .Z(n2460) );
  XNOR U2823 ( .A(a[664]), .B(n2463), .Z(n379) );
  IV U2824 ( .A(n2461), .Z(n2463) );
  XNOR U2825 ( .A(b[664]), .B(n2461), .Z(n2462) );
  XOR U2826 ( .A(n2464), .B(n2465), .Z(n2461) );
  ANDN U2827 ( .B(n2466), .A(n380), .Z(n2464) );
  XNOR U2828 ( .A(a[663]), .B(n2467), .Z(n380) );
  IV U2829 ( .A(n2465), .Z(n2467) );
  XNOR U2830 ( .A(b[663]), .B(n2465), .Z(n2466) );
  XOR U2831 ( .A(n2468), .B(n2469), .Z(n2465) );
  ANDN U2832 ( .B(n2470), .A(n381), .Z(n2468) );
  XNOR U2833 ( .A(a[662]), .B(n2471), .Z(n381) );
  IV U2834 ( .A(n2469), .Z(n2471) );
  XNOR U2835 ( .A(b[662]), .B(n2469), .Z(n2470) );
  XOR U2836 ( .A(n2472), .B(n2473), .Z(n2469) );
  ANDN U2837 ( .B(n2474), .A(n382), .Z(n2472) );
  XNOR U2838 ( .A(a[661]), .B(n2475), .Z(n382) );
  IV U2839 ( .A(n2473), .Z(n2475) );
  XNOR U2840 ( .A(b[661]), .B(n2473), .Z(n2474) );
  XOR U2841 ( .A(n2476), .B(n2477), .Z(n2473) );
  ANDN U2842 ( .B(n2478), .A(n383), .Z(n2476) );
  XNOR U2843 ( .A(a[660]), .B(n2479), .Z(n383) );
  IV U2844 ( .A(n2477), .Z(n2479) );
  XNOR U2845 ( .A(b[660]), .B(n2477), .Z(n2478) );
  XOR U2846 ( .A(n2480), .B(n2481), .Z(n2477) );
  ANDN U2847 ( .B(n2482), .A(n385), .Z(n2480) );
  XNOR U2848 ( .A(a[659]), .B(n2483), .Z(n385) );
  IV U2849 ( .A(n2481), .Z(n2483) );
  XNOR U2850 ( .A(b[659]), .B(n2481), .Z(n2482) );
  XOR U2851 ( .A(n2484), .B(n2485), .Z(n2481) );
  ANDN U2852 ( .B(n2486), .A(n386), .Z(n2484) );
  XNOR U2853 ( .A(a[658]), .B(n2487), .Z(n386) );
  IV U2854 ( .A(n2485), .Z(n2487) );
  XNOR U2855 ( .A(b[658]), .B(n2485), .Z(n2486) );
  XOR U2856 ( .A(n2488), .B(n2489), .Z(n2485) );
  ANDN U2857 ( .B(n2490), .A(n387), .Z(n2488) );
  XNOR U2858 ( .A(a[657]), .B(n2491), .Z(n387) );
  IV U2859 ( .A(n2489), .Z(n2491) );
  XNOR U2860 ( .A(b[657]), .B(n2489), .Z(n2490) );
  XOR U2861 ( .A(n2492), .B(n2493), .Z(n2489) );
  ANDN U2862 ( .B(n2494), .A(n388), .Z(n2492) );
  XNOR U2863 ( .A(a[656]), .B(n2495), .Z(n388) );
  IV U2864 ( .A(n2493), .Z(n2495) );
  XNOR U2865 ( .A(b[656]), .B(n2493), .Z(n2494) );
  XOR U2866 ( .A(n2496), .B(n2497), .Z(n2493) );
  ANDN U2867 ( .B(n2498), .A(n389), .Z(n2496) );
  XNOR U2868 ( .A(a[655]), .B(n2499), .Z(n389) );
  IV U2869 ( .A(n2497), .Z(n2499) );
  XNOR U2870 ( .A(b[655]), .B(n2497), .Z(n2498) );
  XOR U2871 ( .A(n2500), .B(n2501), .Z(n2497) );
  ANDN U2872 ( .B(n2502), .A(n390), .Z(n2500) );
  XNOR U2873 ( .A(a[654]), .B(n2503), .Z(n390) );
  IV U2874 ( .A(n2501), .Z(n2503) );
  XNOR U2875 ( .A(b[654]), .B(n2501), .Z(n2502) );
  XOR U2876 ( .A(n2504), .B(n2505), .Z(n2501) );
  ANDN U2877 ( .B(n2506), .A(n391), .Z(n2504) );
  XNOR U2878 ( .A(a[653]), .B(n2507), .Z(n391) );
  IV U2879 ( .A(n2505), .Z(n2507) );
  XNOR U2880 ( .A(b[653]), .B(n2505), .Z(n2506) );
  XOR U2881 ( .A(n2508), .B(n2509), .Z(n2505) );
  ANDN U2882 ( .B(n2510), .A(n392), .Z(n2508) );
  XNOR U2883 ( .A(a[652]), .B(n2511), .Z(n392) );
  IV U2884 ( .A(n2509), .Z(n2511) );
  XNOR U2885 ( .A(b[652]), .B(n2509), .Z(n2510) );
  XOR U2886 ( .A(n2512), .B(n2513), .Z(n2509) );
  ANDN U2887 ( .B(n2514), .A(n393), .Z(n2512) );
  XNOR U2888 ( .A(a[651]), .B(n2515), .Z(n393) );
  IV U2889 ( .A(n2513), .Z(n2515) );
  XNOR U2890 ( .A(b[651]), .B(n2513), .Z(n2514) );
  XOR U2891 ( .A(n2516), .B(n2517), .Z(n2513) );
  ANDN U2892 ( .B(n2518), .A(n394), .Z(n2516) );
  XNOR U2893 ( .A(a[650]), .B(n2519), .Z(n394) );
  IV U2894 ( .A(n2517), .Z(n2519) );
  XNOR U2895 ( .A(b[650]), .B(n2517), .Z(n2518) );
  XOR U2896 ( .A(n2520), .B(n2521), .Z(n2517) );
  ANDN U2897 ( .B(n2522), .A(n396), .Z(n2520) );
  XNOR U2898 ( .A(a[649]), .B(n2523), .Z(n396) );
  IV U2899 ( .A(n2521), .Z(n2523) );
  XNOR U2900 ( .A(b[649]), .B(n2521), .Z(n2522) );
  XOR U2901 ( .A(n2524), .B(n2525), .Z(n2521) );
  ANDN U2902 ( .B(n2526), .A(n397), .Z(n2524) );
  XNOR U2903 ( .A(a[648]), .B(n2527), .Z(n397) );
  IV U2904 ( .A(n2525), .Z(n2527) );
  XNOR U2905 ( .A(b[648]), .B(n2525), .Z(n2526) );
  XOR U2906 ( .A(n2528), .B(n2529), .Z(n2525) );
  ANDN U2907 ( .B(n2530), .A(n398), .Z(n2528) );
  XNOR U2908 ( .A(a[647]), .B(n2531), .Z(n398) );
  IV U2909 ( .A(n2529), .Z(n2531) );
  XNOR U2910 ( .A(b[647]), .B(n2529), .Z(n2530) );
  XOR U2911 ( .A(n2532), .B(n2533), .Z(n2529) );
  ANDN U2912 ( .B(n2534), .A(n399), .Z(n2532) );
  XNOR U2913 ( .A(a[646]), .B(n2535), .Z(n399) );
  IV U2914 ( .A(n2533), .Z(n2535) );
  XNOR U2915 ( .A(b[646]), .B(n2533), .Z(n2534) );
  XOR U2916 ( .A(n2536), .B(n2537), .Z(n2533) );
  ANDN U2917 ( .B(n2538), .A(n400), .Z(n2536) );
  XNOR U2918 ( .A(a[645]), .B(n2539), .Z(n400) );
  IV U2919 ( .A(n2537), .Z(n2539) );
  XNOR U2920 ( .A(b[645]), .B(n2537), .Z(n2538) );
  XOR U2921 ( .A(n2540), .B(n2541), .Z(n2537) );
  ANDN U2922 ( .B(n2542), .A(n401), .Z(n2540) );
  XNOR U2923 ( .A(a[644]), .B(n2543), .Z(n401) );
  IV U2924 ( .A(n2541), .Z(n2543) );
  XNOR U2925 ( .A(b[644]), .B(n2541), .Z(n2542) );
  XOR U2926 ( .A(n2544), .B(n2545), .Z(n2541) );
  ANDN U2927 ( .B(n2546), .A(n402), .Z(n2544) );
  XNOR U2928 ( .A(a[643]), .B(n2547), .Z(n402) );
  IV U2929 ( .A(n2545), .Z(n2547) );
  XNOR U2930 ( .A(b[643]), .B(n2545), .Z(n2546) );
  XOR U2931 ( .A(n2548), .B(n2549), .Z(n2545) );
  ANDN U2932 ( .B(n2550), .A(n403), .Z(n2548) );
  XNOR U2933 ( .A(a[642]), .B(n2551), .Z(n403) );
  IV U2934 ( .A(n2549), .Z(n2551) );
  XNOR U2935 ( .A(b[642]), .B(n2549), .Z(n2550) );
  XOR U2936 ( .A(n2552), .B(n2553), .Z(n2549) );
  ANDN U2937 ( .B(n2554), .A(n404), .Z(n2552) );
  XNOR U2938 ( .A(a[641]), .B(n2555), .Z(n404) );
  IV U2939 ( .A(n2553), .Z(n2555) );
  XNOR U2940 ( .A(b[641]), .B(n2553), .Z(n2554) );
  XOR U2941 ( .A(n2556), .B(n2557), .Z(n2553) );
  ANDN U2942 ( .B(n2558), .A(n405), .Z(n2556) );
  XNOR U2943 ( .A(a[640]), .B(n2559), .Z(n405) );
  IV U2944 ( .A(n2557), .Z(n2559) );
  XNOR U2945 ( .A(b[640]), .B(n2557), .Z(n2558) );
  XOR U2946 ( .A(n2560), .B(n2561), .Z(n2557) );
  ANDN U2947 ( .B(n2562), .A(n407), .Z(n2560) );
  XNOR U2948 ( .A(a[639]), .B(n2563), .Z(n407) );
  IV U2949 ( .A(n2561), .Z(n2563) );
  XNOR U2950 ( .A(b[639]), .B(n2561), .Z(n2562) );
  XOR U2951 ( .A(n2564), .B(n2565), .Z(n2561) );
  ANDN U2952 ( .B(n2566), .A(n408), .Z(n2564) );
  XNOR U2953 ( .A(a[638]), .B(n2567), .Z(n408) );
  IV U2954 ( .A(n2565), .Z(n2567) );
  XNOR U2955 ( .A(b[638]), .B(n2565), .Z(n2566) );
  XOR U2956 ( .A(n2568), .B(n2569), .Z(n2565) );
  ANDN U2957 ( .B(n2570), .A(n409), .Z(n2568) );
  XNOR U2958 ( .A(a[637]), .B(n2571), .Z(n409) );
  IV U2959 ( .A(n2569), .Z(n2571) );
  XNOR U2960 ( .A(b[637]), .B(n2569), .Z(n2570) );
  XOR U2961 ( .A(n2572), .B(n2573), .Z(n2569) );
  ANDN U2962 ( .B(n2574), .A(n410), .Z(n2572) );
  XNOR U2963 ( .A(a[636]), .B(n2575), .Z(n410) );
  IV U2964 ( .A(n2573), .Z(n2575) );
  XNOR U2965 ( .A(b[636]), .B(n2573), .Z(n2574) );
  XOR U2966 ( .A(n2576), .B(n2577), .Z(n2573) );
  ANDN U2967 ( .B(n2578), .A(n411), .Z(n2576) );
  XNOR U2968 ( .A(a[635]), .B(n2579), .Z(n411) );
  IV U2969 ( .A(n2577), .Z(n2579) );
  XNOR U2970 ( .A(b[635]), .B(n2577), .Z(n2578) );
  XOR U2971 ( .A(n2580), .B(n2581), .Z(n2577) );
  ANDN U2972 ( .B(n2582), .A(n412), .Z(n2580) );
  XNOR U2973 ( .A(a[634]), .B(n2583), .Z(n412) );
  IV U2974 ( .A(n2581), .Z(n2583) );
  XNOR U2975 ( .A(b[634]), .B(n2581), .Z(n2582) );
  XOR U2976 ( .A(n2584), .B(n2585), .Z(n2581) );
  ANDN U2977 ( .B(n2586), .A(n413), .Z(n2584) );
  XNOR U2978 ( .A(a[633]), .B(n2587), .Z(n413) );
  IV U2979 ( .A(n2585), .Z(n2587) );
  XNOR U2980 ( .A(b[633]), .B(n2585), .Z(n2586) );
  XOR U2981 ( .A(n2588), .B(n2589), .Z(n2585) );
  ANDN U2982 ( .B(n2590), .A(n414), .Z(n2588) );
  XNOR U2983 ( .A(a[632]), .B(n2591), .Z(n414) );
  IV U2984 ( .A(n2589), .Z(n2591) );
  XNOR U2985 ( .A(b[632]), .B(n2589), .Z(n2590) );
  XOR U2986 ( .A(n2592), .B(n2593), .Z(n2589) );
  ANDN U2987 ( .B(n2594), .A(n415), .Z(n2592) );
  XNOR U2988 ( .A(a[631]), .B(n2595), .Z(n415) );
  IV U2989 ( .A(n2593), .Z(n2595) );
  XNOR U2990 ( .A(b[631]), .B(n2593), .Z(n2594) );
  XOR U2991 ( .A(n2596), .B(n2597), .Z(n2593) );
  ANDN U2992 ( .B(n2598), .A(n416), .Z(n2596) );
  XNOR U2993 ( .A(a[630]), .B(n2599), .Z(n416) );
  IV U2994 ( .A(n2597), .Z(n2599) );
  XNOR U2995 ( .A(b[630]), .B(n2597), .Z(n2598) );
  XOR U2996 ( .A(n2600), .B(n2601), .Z(n2597) );
  ANDN U2997 ( .B(n2602), .A(n418), .Z(n2600) );
  XNOR U2998 ( .A(a[629]), .B(n2603), .Z(n418) );
  IV U2999 ( .A(n2601), .Z(n2603) );
  XNOR U3000 ( .A(b[629]), .B(n2601), .Z(n2602) );
  XOR U3001 ( .A(n2604), .B(n2605), .Z(n2601) );
  ANDN U3002 ( .B(n2606), .A(n419), .Z(n2604) );
  XNOR U3003 ( .A(a[628]), .B(n2607), .Z(n419) );
  IV U3004 ( .A(n2605), .Z(n2607) );
  XNOR U3005 ( .A(b[628]), .B(n2605), .Z(n2606) );
  XOR U3006 ( .A(n2608), .B(n2609), .Z(n2605) );
  ANDN U3007 ( .B(n2610), .A(n420), .Z(n2608) );
  XNOR U3008 ( .A(a[627]), .B(n2611), .Z(n420) );
  IV U3009 ( .A(n2609), .Z(n2611) );
  XNOR U3010 ( .A(b[627]), .B(n2609), .Z(n2610) );
  XOR U3011 ( .A(n2612), .B(n2613), .Z(n2609) );
  ANDN U3012 ( .B(n2614), .A(n421), .Z(n2612) );
  XNOR U3013 ( .A(a[626]), .B(n2615), .Z(n421) );
  IV U3014 ( .A(n2613), .Z(n2615) );
  XNOR U3015 ( .A(b[626]), .B(n2613), .Z(n2614) );
  XOR U3016 ( .A(n2616), .B(n2617), .Z(n2613) );
  ANDN U3017 ( .B(n2618), .A(n422), .Z(n2616) );
  XNOR U3018 ( .A(a[625]), .B(n2619), .Z(n422) );
  IV U3019 ( .A(n2617), .Z(n2619) );
  XNOR U3020 ( .A(b[625]), .B(n2617), .Z(n2618) );
  XOR U3021 ( .A(n2620), .B(n2621), .Z(n2617) );
  ANDN U3022 ( .B(n2622), .A(n423), .Z(n2620) );
  XNOR U3023 ( .A(a[624]), .B(n2623), .Z(n423) );
  IV U3024 ( .A(n2621), .Z(n2623) );
  XNOR U3025 ( .A(b[624]), .B(n2621), .Z(n2622) );
  XOR U3026 ( .A(n2624), .B(n2625), .Z(n2621) );
  ANDN U3027 ( .B(n2626), .A(n424), .Z(n2624) );
  XNOR U3028 ( .A(a[623]), .B(n2627), .Z(n424) );
  IV U3029 ( .A(n2625), .Z(n2627) );
  XNOR U3030 ( .A(b[623]), .B(n2625), .Z(n2626) );
  XOR U3031 ( .A(n2628), .B(n2629), .Z(n2625) );
  ANDN U3032 ( .B(n2630), .A(n425), .Z(n2628) );
  XNOR U3033 ( .A(a[622]), .B(n2631), .Z(n425) );
  IV U3034 ( .A(n2629), .Z(n2631) );
  XNOR U3035 ( .A(b[622]), .B(n2629), .Z(n2630) );
  XOR U3036 ( .A(n2632), .B(n2633), .Z(n2629) );
  ANDN U3037 ( .B(n2634), .A(n426), .Z(n2632) );
  XNOR U3038 ( .A(a[621]), .B(n2635), .Z(n426) );
  IV U3039 ( .A(n2633), .Z(n2635) );
  XNOR U3040 ( .A(b[621]), .B(n2633), .Z(n2634) );
  XOR U3041 ( .A(n2636), .B(n2637), .Z(n2633) );
  ANDN U3042 ( .B(n2638), .A(n427), .Z(n2636) );
  XNOR U3043 ( .A(a[620]), .B(n2639), .Z(n427) );
  IV U3044 ( .A(n2637), .Z(n2639) );
  XNOR U3045 ( .A(b[620]), .B(n2637), .Z(n2638) );
  XOR U3046 ( .A(n2640), .B(n2641), .Z(n2637) );
  ANDN U3047 ( .B(n2642), .A(n429), .Z(n2640) );
  XNOR U3048 ( .A(a[619]), .B(n2643), .Z(n429) );
  IV U3049 ( .A(n2641), .Z(n2643) );
  XNOR U3050 ( .A(b[619]), .B(n2641), .Z(n2642) );
  XOR U3051 ( .A(n2644), .B(n2645), .Z(n2641) );
  ANDN U3052 ( .B(n2646), .A(n430), .Z(n2644) );
  XNOR U3053 ( .A(a[618]), .B(n2647), .Z(n430) );
  IV U3054 ( .A(n2645), .Z(n2647) );
  XNOR U3055 ( .A(b[618]), .B(n2645), .Z(n2646) );
  XOR U3056 ( .A(n2648), .B(n2649), .Z(n2645) );
  ANDN U3057 ( .B(n2650), .A(n431), .Z(n2648) );
  XNOR U3058 ( .A(a[617]), .B(n2651), .Z(n431) );
  IV U3059 ( .A(n2649), .Z(n2651) );
  XNOR U3060 ( .A(b[617]), .B(n2649), .Z(n2650) );
  XOR U3061 ( .A(n2652), .B(n2653), .Z(n2649) );
  ANDN U3062 ( .B(n2654), .A(n432), .Z(n2652) );
  XNOR U3063 ( .A(a[616]), .B(n2655), .Z(n432) );
  IV U3064 ( .A(n2653), .Z(n2655) );
  XNOR U3065 ( .A(b[616]), .B(n2653), .Z(n2654) );
  XOR U3066 ( .A(n2656), .B(n2657), .Z(n2653) );
  ANDN U3067 ( .B(n2658), .A(n433), .Z(n2656) );
  XNOR U3068 ( .A(a[615]), .B(n2659), .Z(n433) );
  IV U3069 ( .A(n2657), .Z(n2659) );
  XNOR U3070 ( .A(b[615]), .B(n2657), .Z(n2658) );
  XOR U3071 ( .A(n2660), .B(n2661), .Z(n2657) );
  ANDN U3072 ( .B(n2662), .A(n434), .Z(n2660) );
  XNOR U3073 ( .A(a[614]), .B(n2663), .Z(n434) );
  IV U3074 ( .A(n2661), .Z(n2663) );
  XNOR U3075 ( .A(b[614]), .B(n2661), .Z(n2662) );
  XOR U3076 ( .A(n2664), .B(n2665), .Z(n2661) );
  ANDN U3077 ( .B(n2666), .A(n435), .Z(n2664) );
  XNOR U3078 ( .A(a[613]), .B(n2667), .Z(n435) );
  IV U3079 ( .A(n2665), .Z(n2667) );
  XNOR U3080 ( .A(b[613]), .B(n2665), .Z(n2666) );
  XOR U3081 ( .A(n2668), .B(n2669), .Z(n2665) );
  ANDN U3082 ( .B(n2670), .A(n436), .Z(n2668) );
  XNOR U3083 ( .A(a[612]), .B(n2671), .Z(n436) );
  IV U3084 ( .A(n2669), .Z(n2671) );
  XNOR U3085 ( .A(b[612]), .B(n2669), .Z(n2670) );
  XOR U3086 ( .A(n2672), .B(n2673), .Z(n2669) );
  ANDN U3087 ( .B(n2674), .A(n437), .Z(n2672) );
  XNOR U3088 ( .A(a[611]), .B(n2675), .Z(n437) );
  IV U3089 ( .A(n2673), .Z(n2675) );
  XNOR U3090 ( .A(b[611]), .B(n2673), .Z(n2674) );
  XOR U3091 ( .A(n2676), .B(n2677), .Z(n2673) );
  ANDN U3092 ( .B(n2678), .A(n438), .Z(n2676) );
  XNOR U3093 ( .A(a[610]), .B(n2679), .Z(n438) );
  IV U3094 ( .A(n2677), .Z(n2679) );
  XNOR U3095 ( .A(b[610]), .B(n2677), .Z(n2678) );
  XOR U3096 ( .A(n2680), .B(n2681), .Z(n2677) );
  ANDN U3097 ( .B(n2682), .A(n440), .Z(n2680) );
  XNOR U3098 ( .A(a[609]), .B(n2683), .Z(n440) );
  IV U3099 ( .A(n2681), .Z(n2683) );
  XNOR U3100 ( .A(b[609]), .B(n2681), .Z(n2682) );
  XOR U3101 ( .A(n2684), .B(n2685), .Z(n2681) );
  ANDN U3102 ( .B(n2686), .A(n441), .Z(n2684) );
  XNOR U3103 ( .A(a[608]), .B(n2687), .Z(n441) );
  IV U3104 ( .A(n2685), .Z(n2687) );
  XNOR U3105 ( .A(b[608]), .B(n2685), .Z(n2686) );
  XOR U3106 ( .A(n2688), .B(n2689), .Z(n2685) );
  ANDN U3107 ( .B(n2690), .A(n442), .Z(n2688) );
  XNOR U3108 ( .A(a[607]), .B(n2691), .Z(n442) );
  IV U3109 ( .A(n2689), .Z(n2691) );
  XNOR U3110 ( .A(b[607]), .B(n2689), .Z(n2690) );
  XOR U3111 ( .A(n2692), .B(n2693), .Z(n2689) );
  ANDN U3112 ( .B(n2694), .A(n443), .Z(n2692) );
  XNOR U3113 ( .A(a[606]), .B(n2695), .Z(n443) );
  IV U3114 ( .A(n2693), .Z(n2695) );
  XNOR U3115 ( .A(b[606]), .B(n2693), .Z(n2694) );
  XOR U3116 ( .A(n2696), .B(n2697), .Z(n2693) );
  ANDN U3117 ( .B(n2698), .A(n444), .Z(n2696) );
  XNOR U3118 ( .A(a[605]), .B(n2699), .Z(n444) );
  IV U3119 ( .A(n2697), .Z(n2699) );
  XNOR U3120 ( .A(b[605]), .B(n2697), .Z(n2698) );
  XOR U3121 ( .A(n2700), .B(n2701), .Z(n2697) );
  ANDN U3122 ( .B(n2702), .A(n445), .Z(n2700) );
  XNOR U3123 ( .A(a[604]), .B(n2703), .Z(n445) );
  IV U3124 ( .A(n2701), .Z(n2703) );
  XNOR U3125 ( .A(b[604]), .B(n2701), .Z(n2702) );
  XOR U3126 ( .A(n2704), .B(n2705), .Z(n2701) );
  ANDN U3127 ( .B(n2706), .A(n446), .Z(n2704) );
  XNOR U3128 ( .A(a[603]), .B(n2707), .Z(n446) );
  IV U3129 ( .A(n2705), .Z(n2707) );
  XNOR U3130 ( .A(b[603]), .B(n2705), .Z(n2706) );
  XOR U3131 ( .A(n2708), .B(n2709), .Z(n2705) );
  ANDN U3132 ( .B(n2710), .A(n447), .Z(n2708) );
  XNOR U3133 ( .A(a[602]), .B(n2711), .Z(n447) );
  IV U3134 ( .A(n2709), .Z(n2711) );
  XNOR U3135 ( .A(b[602]), .B(n2709), .Z(n2710) );
  XOR U3136 ( .A(n2712), .B(n2713), .Z(n2709) );
  ANDN U3137 ( .B(n2714), .A(n448), .Z(n2712) );
  XNOR U3138 ( .A(a[601]), .B(n2715), .Z(n448) );
  IV U3139 ( .A(n2713), .Z(n2715) );
  XNOR U3140 ( .A(b[601]), .B(n2713), .Z(n2714) );
  XOR U3141 ( .A(n2716), .B(n2717), .Z(n2713) );
  ANDN U3142 ( .B(n2718), .A(n449), .Z(n2716) );
  XNOR U3143 ( .A(a[600]), .B(n2719), .Z(n449) );
  IV U3144 ( .A(n2717), .Z(n2719) );
  XNOR U3145 ( .A(b[600]), .B(n2717), .Z(n2718) );
  XOR U3146 ( .A(n2720), .B(n2721), .Z(n2717) );
  ANDN U3147 ( .B(n2722), .A(n452), .Z(n2720) );
  XNOR U3148 ( .A(a[599]), .B(n2723), .Z(n452) );
  IV U3149 ( .A(n2721), .Z(n2723) );
  XNOR U3150 ( .A(b[599]), .B(n2721), .Z(n2722) );
  XOR U3151 ( .A(n2724), .B(n2725), .Z(n2721) );
  ANDN U3152 ( .B(n2726), .A(n453), .Z(n2724) );
  XNOR U3153 ( .A(a[598]), .B(n2727), .Z(n453) );
  IV U3154 ( .A(n2725), .Z(n2727) );
  XNOR U3155 ( .A(b[598]), .B(n2725), .Z(n2726) );
  XOR U3156 ( .A(n2728), .B(n2729), .Z(n2725) );
  ANDN U3157 ( .B(n2730), .A(n454), .Z(n2728) );
  XNOR U3158 ( .A(a[597]), .B(n2731), .Z(n454) );
  IV U3159 ( .A(n2729), .Z(n2731) );
  XNOR U3160 ( .A(b[597]), .B(n2729), .Z(n2730) );
  XOR U3161 ( .A(n2732), .B(n2733), .Z(n2729) );
  ANDN U3162 ( .B(n2734), .A(n455), .Z(n2732) );
  XNOR U3163 ( .A(a[596]), .B(n2735), .Z(n455) );
  IV U3164 ( .A(n2733), .Z(n2735) );
  XNOR U3165 ( .A(b[596]), .B(n2733), .Z(n2734) );
  XOR U3166 ( .A(n2736), .B(n2737), .Z(n2733) );
  ANDN U3167 ( .B(n2738), .A(n456), .Z(n2736) );
  XNOR U3168 ( .A(a[595]), .B(n2739), .Z(n456) );
  IV U3169 ( .A(n2737), .Z(n2739) );
  XNOR U3170 ( .A(b[595]), .B(n2737), .Z(n2738) );
  XOR U3171 ( .A(n2740), .B(n2741), .Z(n2737) );
  ANDN U3172 ( .B(n2742), .A(n457), .Z(n2740) );
  XNOR U3173 ( .A(a[594]), .B(n2743), .Z(n457) );
  IV U3174 ( .A(n2741), .Z(n2743) );
  XNOR U3175 ( .A(b[594]), .B(n2741), .Z(n2742) );
  XOR U3176 ( .A(n2744), .B(n2745), .Z(n2741) );
  ANDN U3177 ( .B(n2746), .A(n458), .Z(n2744) );
  XNOR U3178 ( .A(a[593]), .B(n2747), .Z(n458) );
  IV U3179 ( .A(n2745), .Z(n2747) );
  XNOR U3180 ( .A(b[593]), .B(n2745), .Z(n2746) );
  XOR U3181 ( .A(n2748), .B(n2749), .Z(n2745) );
  ANDN U3182 ( .B(n2750), .A(n459), .Z(n2748) );
  XNOR U3183 ( .A(a[592]), .B(n2751), .Z(n459) );
  IV U3184 ( .A(n2749), .Z(n2751) );
  XNOR U3185 ( .A(b[592]), .B(n2749), .Z(n2750) );
  XOR U3186 ( .A(n2752), .B(n2753), .Z(n2749) );
  ANDN U3187 ( .B(n2754), .A(n460), .Z(n2752) );
  XNOR U3188 ( .A(a[591]), .B(n2755), .Z(n460) );
  IV U3189 ( .A(n2753), .Z(n2755) );
  XNOR U3190 ( .A(b[591]), .B(n2753), .Z(n2754) );
  XOR U3191 ( .A(n2756), .B(n2757), .Z(n2753) );
  ANDN U3192 ( .B(n2758), .A(n461), .Z(n2756) );
  XNOR U3193 ( .A(a[590]), .B(n2759), .Z(n461) );
  IV U3194 ( .A(n2757), .Z(n2759) );
  XNOR U3195 ( .A(b[590]), .B(n2757), .Z(n2758) );
  XOR U3196 ( .A(n2760), .B(n2761), .Z(n2757) );
  ANDN U3197 ( .B(n2762), .A(n463), .Z(n2760) );
  XNOR U3198 ( .A(a[589]), .B(n2763), .Z(n463) );
  IV U3199 ( .A(n2761), .Z(n2763) );
  XNOR U3200 ( .A(b[589]), .B(n2761), .Z(n2762) );
  XOR U3201 ( .A(n2764), .B(n2765), .Z(n2761) );
  ANDN U3202 ( .B(n2766), .A(n464), .Z(n2764) );
  XNOR U3203 ( .A(a[588]), .B(n2767), .Z(n464) );
  IV U3204 ( .A(n2765), .Z(n2767) );
  XNOR U3205 ( .A(b[588]), .B(n2765), .Z(n2766) );
  XOR U3206 ( .A(n2768), .B(n2769), .Z(n2765) );
  ANDN U3207 ( .B(n2770), .A(n465), .Z(n2768) );
  XNOR U3208 ( .A(a[587]), .B(n2771), .Z(n465) );
  IV U3209 ( .A(n2769), .Z(n2771) );
  XNOR U3210 ( .A(b[587]), .B(n2769), .Z(n2770) );
  XOR U3211 ( .A(n2772), .B(n2773), .Z(n2769) );
  ANDN U3212 ( .B(n2774), .A(n466), .Z(n2772) );
  XNOR U3213 ( .A(a[586]), .B(n2775), .Z(n466) );
  IV U3214 ( .A(n2773), .Z(n2775) );
  XNOR U3215 ( .A(b[586]), .B(n2773), .Z(n2774) );
  XOR U3216 ( .A(n2776), .B(n2777), .Z(n2773) );
  ANDN U3217 ( .B(n2778), .A(n467), .Z(n2776) );
  XNOR U3218 ( .A(a[585]), .B(n2779), .Z(n467) );
  IV U3219 ( .A(n2777), .Z(n2779) );
  XNOR U3220 ( .A(b[585]), .B(n2777), .Z(n2778) );
  XOR U3221 ( .A(n2780), .B(n2781), .Z(n2777) );
  ANDN U3222 ( .B(n2782), .A(n468), .Z(n2780) );
  XNOR U3223 ( .A(a[584]), .B(n2783), .Z(n468) );
  IV U3224 ( .A(n2781), .Z(n2783) );
  XNOR U3225 ( .A(b[584]), .B(n2781), .Z(n2782) );
  XOR U3226 ( .A(n2784), .B(n2785), .Z(n2781) );
  ANDN U3227 ( .B(n2786), .A(n469), .Z(n2784) );
  XNOR U3228 ( .A(a[583]), .B(n2787), .Z(n469) );
  IV U3229 ( .A(n2785), .Z(n2787) );
  XNOR U3230 ( .A(b[583]), .B(n2785), .Z(n2786) );
  XOR U3231 ( .A(n2788), .B(n2789), .Z(n2785) );
  ANDN U3232 ( .B(n2790), .A(n470), .Z(n2788) );
  XNOR U3233 ( .A(a[582]), .B(n2791), .Z(n470) );
  IV U3234 ( .A(n2789), .Z(n2791) );
  XNOR U3235 ( .A(b[582]), .B(n2789), .Z(n2790) );
  XOR U3236 ( .A(n2792), .B(n2793), .Z(n2789) );
  ANDN U3237 ( .B(n2794), .A(n471), .Z(n2792) );
  XNOR U3238 ( .A(a[581]), .B(n2795), .Z(n471) );
  IV U3239 ( .A(n2793), .Z(n2795) );
  XNOR U3240 ( .A(b[581]), .B(n2793), .Z(n2794) );
  XOR U3241 ( .A(n2796), .B(n2797), .Z(n2793) );
  ANDN U3242 ( .B(n2798), .A(n472), .Z(n2796) );
  XNOR U3243 ( .A(a[580]), .B(n2799), .Z(n472) );
  IV U3244 ( .A(n2797), .Z(n2799) );
  XNOR U3245 ( .A(b[580]), .B(n2797), .Z(n2798) );
  XOR U3246 ( .A(n2800), .B(n2801), .Z(n2797) );
  ANDN U3247 ( .B(n2802), .A(n474), .Z(n2800) );
  XNOR U3248 ( .A(a[579]), .B(n2803), .Z(n474) );
  IV U3249 ( .A(n2801), .Z(n2803) );
  XNOR U3250 ( .A(b[579]), .B(n2801), .Z(n2802) );
  XOR U3251 ( .A(n2804), .B(n2805), .Z(n2801) );
  ANDN U3252 ( .B(n2806), .A(n475), .Z(n2804) );
  XNOR U3253 ( .A(a[578]), .B(n2807), .Z(n475) );
  IV U3254 ( .A(n2805), .Z(n2807) );
  XNOR U3255 ( .A(b[578]), .B(n2805), .Z(n2806) );
  XOR U3256 ( .A(n2808), .B(n2809), .Z(n2805) );
  ANDN U3257 ( .B(n2810), .A(n476), .Z(n2808) );
  XNOR U3258 ( .A(a[577]), .B(n2811), .Z(n476) );
  IV U3259 ( .A(n2809), .Z(n2811) );
  XNOR U3260 ( .A(b[577]), .B(n2809), .Z(n2810) );
  XOR U3261 ( .A(n2812), .B(n2813), .Z(n2809) );
  ANDN U3262 ( .B(n2814), .A(n477), .Z(n2812) );
  XNOR U3263 ( .A(a[576]), .B(n2815), .Z(n477) );
  IV U3264 ( .A(n2813), .Z(n2815) );
  XNOR U3265 ( .A(b[576]), .B(n2813), .Z(n2814) );
  XOR U3266 ( .A(n2816), .B(n2817), .Z(n2813) );
  ANDN U3267 ( .B(n2818), .A(n478), .Z(n2816) );
  XNOR U3268 ( .A(a[575]), .B(n2819), .Z(n478) );
  IV U3269 ( .A(n2817), .Z(n2819) );
  XNOR U3270 ( .A(b[575]), .B(n2817), .Z(n2818) );
  XOR U3271 ( .A(n2820), .B(n2821), .Z(n2817) );
  ANDN U3272 ( .B(n2822), .A(n479), .Z(n2820) );
  XNOR U3273 ( .A(a[574]), .B(n2823), .Z(n479) );
  IV U3274 ( .A(n2821), .Z(n2823) );
  XNOR U3275 ( .A(b[574]), .B(n2821), .Z(n2822) );
  XOR U3276 ( .A(n2824), .B(n2825), .Z(n2821) );
  ANDN U3277 ( .B(n2826), .A(n480), .Z(n2824) );
  XNOR U3278 ( .A(a[573]), .B(n2827), .Z(n480) );
  IV U3279 ( .A(n2825), .Z(n2827) );
  XNOR U3280 ( .A(b[573]), .B(n2825), .Z(n2826) );
  XOR U3281 ( .A(n2828), .B(n2829), .Z(n2825) );
  ANDN U3282 ( .B(n2830), .A(n481), .Z(n2828) );
  XNOR U3283 ( .A(a[572]), .B(n2831), .Z(n481) );
  IV U3284 ( .A(n2829), .Z(n2831) );
  XNOR U3285 ( .A(b[572]), .B(n2829), .Z(n2830) );
  XOR U3286 ( .A(n2832), .B(n2833), .Z(n2829) );
  ANDN U3287 ( .B(n2834), .A(n482), .Z(n2832) );
  XNOR U3288 ( .A(a[571]), .B(n2835), .Z(n482) );
  IV U3289 ( .A(n2833), .Z(n2835) );
  XNOR U3290 ( .A(b[571]), .B(n2833), .Z(n2834) );
  XOR U3291 ( .A(n2836), .B(n2837), .Z(n2833) );
  ANDN U3292 ( .B(n2838), .A(n483), .Z(n2836) );
  XNOR U3293 ( .A(a[570]), .B(n2839), .Z(n483) );
  IV U3294 ( .A(n2837), .Z(n2839) );
  XNOR U3295 ( .A(b[570]), .B(n2837), .Z(n2838) );
  XOR U3296 ( .A(n2840), .B(n2841), .Z(n2837) );
  ANDN U3297 ( .B(n2842), .A(n485), .Z(n2840) );
  XNOR U3298 ( .A(a[569]), .B(n2843), .Z(n485) );
  IV U3299 ( .A(n2841), .Z(n2843) );
  XNOR U3300 ( .A(b[569]), .B(n2841), .Z(n2842) );
  XOR U3301 ( .A(n2844), .B(n2845), .Z(n2841) );
  ANDN U3302 ( .B(n2846), .A(n486), .Z(n2844) );
  XNOR U3303 ( .A(a[568]), .B(n2847), .Z(n486) );
  IV U3304 ( .A(n2845), .Z(n2847) );
  XNOR U3305 ( .A(b[568]), .B(n2845), .Z(n2846) );
  XOR U3306 ( .A(n2848), .B(n2849), .Z(n2845) );
  ANDN U3307 ( .B(n2850), .A(n487), .Z(n2848) );
  XNOR U3308 ( .A(a[567]), .B(n2851), .Z(n487) );
  IV U3309 ( .A(n2849), .Z(n2851) );
  XNOR U3310 ( .A(b[567]), .B(n2849), .Z(n2850) );
  XOR U3311 ( .A(n2852), .B(n2853), .Z(n2849) );
  ANDN U3312 ( .B(n2854), .A(n488), .Z(n2852) );
  XNOR U3313 ( .A(a[566]), .B(n2855), .Z(n488) );
  IV U3314 ( .A(n2853), .Z(n2855) );
  XNOR U3315 ( .A(b[566]), .B(n2853), .Z(n2854) );
  XOR U3316 ( .A(n2856), .B(n2857), .Z(n2853) );
  ANDN U3317 ( .B(n2858), .A(n489), .Z(n2856) );
  XNOR U3318 ( .A(a[565]), .B(n2859), .Z(n489) );
  IV U3319 ( .A(n2857), .Z(n2859) );
  XNOR U3320 ( .A(b[565]), .B(n2857), .Z(n2858) );
  XOR U3321 ( .A(n2860), .B(n2861), .Z(n2857) );
  ANDN U3322 ( .B(n2862), .A(n490), .Z(n2860) );
  XNOR U3323 ( .A(a[564]), .B(n2863), .Z(n490) );
  IV U3324 ( .A(n2861), .Z(n2863) );
  XNOR U3325 ( .A(b[564]), .B(n2861), .Z(n2862) );
  XOR U3326 ( .A(n2864), .B(n2865), .Z(n2861) );
  ANDN U3327 ( .B(n2866), .A(n491), .Z(n2864) );
  XNOR U3328 ( .A(a[563]), .B(n2867), .Z(n491) );
  IV U3329 ( .A(n2865), .Z(n2867) );
  XNOR U3330 ( .A(b[563]), .B(n2865), .Z(n2866) );
  XOR U3331 ( .A(n2868), .B(n2869), .Z(n2865) );
  ANDN U3332 ( .B(n2870), .A(n492), .Z(n2868) );
  XNOR U3333 ( .A(a[562]), .B(n2871), .Z(n492) );
  IV U3334 ( .A(n2869), .Z(n2871) );
  XNOR U3335 ( .A(b[562]), .B(n2869), .Z(n2870) );
  XOR U3336 ( .A(n2872), .B(n2873), .Z(n2869) );
  ANDN U3337 ( .B(n2874), .A(n493), .Z(n2872) );
  XNOR U3338 ( .A(a[561]), .B(n2875), .Z(n493) );
  IV U3339 ( .A(n2873), .Z(n2875) );
  XNOR U3340 ( .A(b[561]), .B(n2873), .Z(n2874) );
  XOR U3341 ( .A(n2876), .B(n2877), .Z(n2873) );
  ANDN U3342 ( .B(n2878), .A(n494), .Z(n2876) );
  XNOR U3343 ( .A(a[560]), .B(n2879), .Z(n494) );
  IV U3344 ( .A(n2877), .Z(n2879) );
  XNOR U3345 ( .A(b[560]), .B(n2877), .Z(n2878) );
  XOR U3346 ( .A(n2880), .B(n2881), .Z(n2877) );
  ANDN U3347 ( .B(n2882), .A(n496), .Z(n2880) );
  XNOR U3348 ( .A(a[559]), .B(n2883), .Z(n496) );
  IV U3349 ( .A(n2881), .Z(n2883) );
  XNOR U3350 ( .A(b[559]), .B(n2881), .Z(n2882) );
  XOR U3351 ( .A(n2884), .B(n2885), .Z(n2881) );
  ANDN U3352 ( .B(n2886), .A(n497), .Z(n2884) );
  XNOR U3353 ( .A(a[558]), .B(n2887), .Z(n497) );
  IV U3354 ( .A(n2885), .Z(n2887) );
  XNOR U3355 ( .A(b[558]), .B(n2885), .Z(n2886) );
  XOR U3356 ( .A(n2888), .B(n2889), .Z(n2885) );
  ANDN U3357 ( .B(n2890), .A(n498), .Z(n2888) );
  XNOR U3358 ( .A(a[557]), .B(n2891), .Z(n498) );
  IV U3359 ( .A(n2889), .Z(n2891) );
  XNOR U3360 ( .A(b[557]), .B(n2889), .Z(n2890) );
  XOR U3361 ( .A(n2892), .B(n2893), .Z(n2889) );
  ANDN U3362 ( .B(n2894), .A(n499), .Z(n2892) );
  XNOR U3363 ( .A(a[556]), .B(n2895), .Z(n499) );
  IV U3364 ( .A(n2893), .Z(n2895) );
  XNOR U3365 ( .A(b[556]), .B(n2893), .Z(n2894) );
  XOR U3366 ( .A(n2896), .B(n2897), .Z(n2893) );
  ANDN U3367 ( .B(n2898), .A(n500), .Z(n2896) );
  XNOR U3368 ( .A(a[555]), .B(n2899), .Z(n500) );
  IV U3369 ( .A(n2897), .Z(n2899) );
  XNOR U3370 ( .A(b[555]), .B(n2897), .Z(n2898) );
  XOR U3371 ( .A(n2900), .B(n2901), .Z(n2897) );
  ANDN U3372 ( .B(n2902), .A(n501), .Z(n2900) );
  XNOR U3373 ( .A(a[554]), .B(n2903), .Z(n501) );
  IV U3374 ( .A(n2901), .Z(n2903) );
  XNOR U3375 ( .A(b[554]), .B(n2901), .Z(n2902) );
  XOR U3376 ( .A(n2904), .B(n2905), .Z(n2901) );
  ANDN U3377 ( .B(n2906), .A(n502), .Z(n2904) );
  XNOR U3378 ( .A(a[553]), .B(n2907), .Z(n502) );
  IV U3379 ( .A(n2905), .Z(n2907) );
  XNOR U3380 ( .A(b[553]), .B(n2905), .Z(n2906) );
  XOR U3381 ( .A(n2908), .B(n2909), .Z(n2905) );
  ANDN U3382 ( .B(n2910), .A(n503), .Z(n2908) );
  XNOR U3383 ( .A(a[552]), .B(n2911), .Z(n503) );
  IV U3384 ( .A(n2909), .Z(n2911) );
  XNOR U3385 ( .A(b[552]), .B(n2909), .Z(n2910) );
  XOR U3386 ( .A(n2912), .B(n2913), .Z(n2909) );
  ANDN U3387 ( .B(n2914), .A(n504), .Z(n2912) );
  XNOR U3388 ( .A(a[551]), .B(n2915), .Z(n504) );
  IV U3389 ( .A(n2913), .Z(n2915) );
  XNOR U3390 ( .A(b[551]), .B(n2913), .Z(n2914) );
  XOR U3391 ( .A(n2916), .B(n2917), .Z(n2913) );
  ANDN U3392 ( .B(n2918), .A(n505), .Z(n2916) );
  XNOR U3393 ( .A(a[550]), .B(n2919), .Z(n505) );
  IV U3394 ( .A(n2917), .Z(n2919) );
  XNOR U3395 ( .A(b[550]), .B(n2917), .Z(n2918) );
  XOR U3396 ( .A(n2920), .B(n2921), .Z(n2917) );
  ANDN U3397 ( .B(n2922), .A(n507), .Z(n2920) );
  XNOR U3398 ( .A(a[549]), .B(n2923), .Z(n507) );
  IV U3399 ( .A(n2921), .Z(n2923) );
  XNOR U3400 ( .A(b[549]), .B(n2921), .Z(n2922) );
  XOR U3401 ( .A(n2924), .B(n2925), .Z(n2921) );
  ANDN U3402 ( .B(n2926), .A(n508), .Z(n2924) );
  XNOR U3403 ( .A(a[548]), .B(n2927), .Z(n508) );
  IV U3404 ( .A(n2925), .Z(n2927) );
  XNOR U3405 ( .A(b[548]), .B(n2925), .Z(n2926) );
  XOR U3406 ( .A(n2928), .B(n2929), .Z(n2925) );
  ANDN U3407 ( .B(n2930), .A(n509), .Z(n2928) );
  XNOR U3408 ( .A(a[547]), .B(n2931), .Z(n509) );
  IV U3409 ( .A(n2929), .Z(n2931) );
  XNOR U3410 ( .A(b[547]), .B(n2929), .Z(n2930) );
  XOR U3411 ( .A(n2932), .B(n2933), .Z(n2929) );
  ANDN U3412 ( .B(n2934), .A(n510), .Z(n2932) );
  XNOR U3413 ( .A(a[546]), .B(n2935), .Z(n510) );
  IV U3414 ( .A(n2933), .Z(n2935) );
  XNOR U3415 ( .A(b[546]), .B(n2933), .Z(n2934) );
  XOR U3416 ( .A(n2936), .B(n2937), .Z(n2933) );
  ANDN U3417 ( .B(n2938), .A(n511), .Z(n2936) );
  XNOR U3418 ( .A(a[545]), .B(n2939), .Z(n511) );
  IV U3419 ( .A(n2937), .Z(n2939) );
  XNOR U3420 ( .A(b[545]), .B(n2937), .Z(n2938) );
  XOR U3421 ( .A(n2940), .B(n2941), .Z(n2937) );
  ANDN U3422 ( .B(n2942), .A(n512), .Z(n2940) );
  XNOR U3423 ( .A(a[544]), .B(n2943), .Z(n512) );
  IV U3424 ( .A(n2941), .Z(n2943) );
  XNOR U3425 ( .A(b[544]), .B(n2941), .Z(n2942) );
  XOR U3426 ( .A(n2944), .B(n2945), .Z(n2941) );
  ANDN U3427 ( .B(n2946), .A(n513), .Z(n2944) );
  XNOR U3428 ( .A(a[543]), .B(n2947), .Z(n513) );
  IV U3429 ( .A(n2945), .Z(n2947) );
  XNOR U3430 ( .A(b[543]), .B(n2945), .Z(n2946) );
  XOR U3431 ( .A(n2948), .B(n2949), .Z(n2945) );
  ANDN U3432 ( .B(n2950), .A(n514), .Z(n2948) );
  XNOR U3433 ( .A(a[542]), .B(n2951), .Z(n514) );
  IV U3434 ( .A(n2949), .Z(n2951) );
  XNOR U3435 ( .A(b[542]), .B(n2949), .Z(n2950) );
  XOR U3436 ( .A(n2952), .B(n2953), .Z(n2949) );
  ANDN U3437 ( .B(n2954), .A(n515), .Z(n2952) );
  XNOR U3438 ( .A(a[541]), .B(n2955), .Z(n515) );
  IV U3439 ( .A(n2953), .Z(n2955) );
  XNOR U3440 ( .A(b[541]), .B(n2953), .Z(n2954) );
  XOR U3441 ( .A(n2956), .B(n2957), .Z(n2953) );
  ANDN U3442 ( .B(n2958), .A(n516), .Z(n2956) );
  XNOR U3443 ( .A(a[540]), .B(n2959), .Z(n516) );
  IV U3444 ( .A(n2957), .Z(n2959) );
  XNOR U3445 ( .A(b[540]), .B(n2957), .Z(n2958) );
  XOR U3446 ( .A(n2960), .B(n2961), .Z(n2957) );
  ANDN U3447 ( .B(n2962), .A(n518), .Z(n2960) );
  XNOR U3448 ( .A(a[539]), .B(n2963), .Z(n518) );
  IV U3449 ( .A(n2961), .Z(n2963) );
  XNOR U3450 ( .A(b[539]), .B(n2961), .Z(n2962) );
  XOR U3451 ( .A(n2964), .B(n2965), .Z(n2961) );
  ANDN U3452 ( .B(n2966), .A(n519), .Z(n2964) );
  XNOR U3453 ( .A(a[538]), .B(n2967), .Z(n519) );
  IV U3454 ( .A(n2965), .Z(n2967) );
  XNOR U3455 ( .A(b[538]), .B(n2965), .Z(n2966) );
  XOR U3456 ( .A(n2968), .B(n2969), .Z(n2965) );
  ANDN U3457 ( .B(n2970), .A(n520), .Z(n2968) );
  XNOR U3458 ( .A(a[537]), .B(n2971), .Z(n520) );
  IV U3459 ( .A(n2969), .Z(n2971) );
  XNOR U3460 ( .A(b[537]), .B(n2969), .Z(n2970) );
  XOR U3461 ( .A(n2972), .B(n2973), .Z(n2969) );
  ANDN U3462 ( .B(n2974), .A(n521), .Z(n2972) );
  XNOR U3463 ( .A(a[536]), .B(n2975), .Z(n521) );
  IV U3464 ( .A(n2973), .Z(n2975) );
  XNOR U3465 ( .A(b[536]), .B(n2973), .Z(n2974) );
  XOR U3466 ( .A(n2976), .B(n2977), .Z(n2973) );
  ANDN U3467 ( .B(n2978), .A(n522), .Z(n2976) );
  XNOR U3468 ( .A(a[535]), .B(n2979), .Z(n522) );
  IV U3469 ( .A(n2977), .Z(n2979) );
  XNOR U3470 ( .A(b[535]), .B(n2977), .Z(n2978) );
  XOR U3471 ( .A(n2980), .B(n2981), .Z(n2977) );
  ANDN U3472 ( .B(n2982), .A(n523), .Z(n2980) );
  XNOR U3473 ( .A(a[534]), .B(n2983), .Z(n523) );
  IV U3474 ( .A(n2981), .Z(n2983) );
  XNOR U3475 ( .A(b[534]), .B(n2981), .Z(n2982) );
  XOR U3476 ( .A(n2984), .B(n2985), .Z(n2981) );
  ANDN U3477 ( .B(n2986), .A(n524), .Z(n2984) );
  XNOR U3478 ( .A(a[533]), .B(n2987), .Z(n524) );
  IV U3479 ( .A(n2985), .Z(n2987) );
  XNOR U3480 ( .A(b[533]), .B(n2985), .Z(n2986) );
  XOR U3481 ( .A(n2988), .B(n2989), .Z(n2985) );
  ANDN U3482 ( .B(n2990), .A(n525), .Z(n2988) );
  XNOR U3483 ( .A(a[532]), .B(n2991), .Z(n525) );
  IV U3484 ( .A(n2989), .Z(n2991) );
  XNOR U3485 ( .A(b[532]), .B(n2989), .Z(n2990) );
  XOR U3486 ( .A(n2992), .B(n2993), .Z(n2989) );
  ANDN U3487 ( .B(n2994), .A(n526), .Z(n2992) );
  XNOR U3488 ( .A(a[531]), .B(n2995), .Z(n526) );
  IV U3489 ( .A(n2993), .Z(n2995) );
  XNOR U3490 ( .A(b[531]), .B(n2993), .Z(n2994) );
  XOR U3491 ( .A(n2996), .B(n2997), .Z(n2993) );
  ANDN U3492 ( .B(n2998), .A(n527), .Z(n2996) );
  XNOR U3493 ( .A(a[530]), .B(n2999), .Z(n527) );
  IV U3494 ( .A(n2997), .Z(n2999) );
  XNOR U3495 ( .A(b[530]), .B(n2997), .Z(n2998) );
  XOR U3496 ( .A(n3000), .B(n3001), .Z(n2997) );
  ANDN U3497 ( .B(n3002), .A(n529), .Z(n3000) );
  XNOR U3498 ( .A(a[529]), .B(n3003), .Z(n529) );
  IV U3499 ( .A(n3001), .Z(n3003) );
  XNOR U3500 ( .A(b[529]), .B(n3001), .Z(n3002) );
  XOR U3501 ( .A(n3004), .B(n3005), .Z(n3001) );
  ANDN U3502 ( .B(n3006), .A(n530), .Z(n3004) );
  XNOR U3503 ( .A(a[528]), .B(n3007), .Z(n530) );
  IV U3504 ( .A(n3005), .Z(n3007) );
  XNOR U3505 ( .A(b[528]), .B(n3005), .Z(n3006) );
  XOR U3506 ( .A(n3008), .B(n3009), .Z(n3005) );
  ANDN U3507 ( .B(n3010), .A(n531), .Z(n3008) );
  XNOR U3508 ( .A(a[527]), .B(n3011), .Z(n531) );
  IV U3509 ( .A(n3009), .Z(n3011) );
  XNOR U3510 ( .A(b[527]), .B(n3009), .Z(n3010) );
  XOR U3511 ( .A(n3012), .B(n3013), .Z(n3009) );
  ANDN U3512 ( .B(n3014), .A(n532), .Z(n3012) );
  XNOR U3513 ( .A(a[526]), .B(n3015), .Z(n532) );
  IV U3514 ( .A(n3013), .Z(n3015) );
  XNOR U3515 ( .A(b[526]), .B(n3013), .Z(n3014) );
  XOR U3516 ( .A(n3016), .B(n3017), .Z(n3013) );
  ANDN U3517 ( .B(n3018), .A(n533), .Z(n3016) );
  XNOR U3518 ( .A(a[525]), .B(n3019), .Z(n533) );
  IV U3519 ( .A(n3017), .Z(n3019) );
  XNOR U3520 ( .A(b[525]), .B(n3017), .Z(n3018) );
  XOR U3521 ( .A(n3020), .B(n3021), .Z(n3017) );
  ANDN U3522 ( .B(n3022), .A(n534), .Z(n3020) );
  XNOR U3523 ( .A(a[524]), .B(n3023), .Z(n534) );
  IV U3524 ( .A(n3021), .Z(n3023) );
  XNOR U3525 ( .A(b[524]), .B(n3021), .Z(n3022) );
  XOR U3526 ( .A(n3024), .B(n3025), .Z(n3021) );
  ANDN U3527 ( .B(n3026), .A(n535), .Z(n3024) );
  XNOR U3528 ( .A(a[523]), .B(n3027), .Z(n535) );
  IV U3529 ( .A(n3025), .Z(n3027) );
  XNOR U3530 ( .A(b[523]), .B(n3025), .Z(n3026) );
  XOR U3531 ( .A(n3028), .B(n3029), .Z(n3025) );
  ANDN U3532 ( .B(n3030), .A(n536), .Z(n3028) );
  XNOR U3533 ( .A(a[522]), .B(n3031), .Z(n536) );
  IV U3534 ( .A(n3029), .Z(n3031) );
  XNOR U3535 ( .A(b[522]), .B(n3029), .Z(n3030) );
  XOR U3536 ( .A(n3032), .B(n3033), .Z(n3029) );
  ANDN U3537 ( .B(n3034), .A(n537), .Z(n3032) );
  XNOR U3538 ( .A(a[521]), .B(n3035), .Z(n537) );
  IV U3539 ( .A(n3033), .Z(n3035) );
  XNOR U3540 ( .A(b[521]), .B(n3033), .Z(n3034) );
  XOR U3541 ( .A(n3036), .B(n3037), .Z(n3033) );
  ANDN U3542 ( .B(n3038), .A(n538), .Z(n3036) );
  XNOR U3543 ( .A(a[520]), .B(n3039), .Z(n538) );
  IV U3544 ( .A(n3037), .Z(n3039) );
  XNOR U3545 ( .A(b[520]), .B(n3037), .Z(n3038) );
  XOR U3546 ( .A(n3040), .B(n3041), .Z(n3037) );
  ANDN U3547 ( .B(n3042), .A(n540), .Z(n3040) );
  XNOR U3548 ( .A(a[519]), .B(n3043), .Z(n540) );
  IV U3549 ( .A(n3041), .Z(n3043) );
  XNOR U3550 ( .A(b[519]), .B(n3041), .Z(n3042) );
  XOR U3551 ( .A(n3044), .B(n3045), .Z(n3041) );
  ANDN U3552 ( .B(n3046), .A(n541), .Z(n3044) );
  XNOR U3553 ( .A(a[518]), .B(n3047), .Z(n541) );
  IV U3554 ( .A(n3045), .Z(n3047) );
  XNOR U3555 ( .A(b[518]), .B(n3045), .Z(n3046) );
  XOR U3556 ( .A(n3048), .B(n3049), .Z(n3045) );
  ANDN U3557 ( .B(n3050), .A(n542), .Z(n3048) );
  XNOR U3558 ( .A(a[517]), .B(n3051), .Z(n542) );
  IV U3559 ( .A(n3049), .Z(n3051) );
  XNOR U3560 ( .A(b[517]), .B(n3049), .Z(n3050) );
  XOR U3561 ( .A(n3052), .B(n3053), .Z(n3049) );
  ANDN U3562 ( .B(n3054), .A(n543), .Z(n3052) );
  XNOR U3563 ( .A(a[516]), .B(n3055), .Z(n543) );
  IV U3564 ( .A(n3053), .Z(n3055) );
  XNOR U3565 ( .A(b[516]), .B(n3053), .Z(n3054) );
  XOR U3566 ( .A(n3056), .B(n3057), .Z(n3053) );
  ANDN U3567 ( .B(n3058), .A(n544), .Z(n3056) );
  XNOR U3568 ( .A(a[515]), .B(n3059), .Z(n544) );
  IV U3569 ( .A(n3057), .Z(n3059) );
  XNOR U3570 ( .A(b[515]), .B(n3057), .Z(n3058) );
  XOR U3571 ( .A(n3060), .B(n3061), .Z(n3057) );
  ANDN U3572 ( .B(n3062), .A(n545), .Z(n3060) );
  XNOR U3573 ( .A(a[514]), .B(n3063), .Z(n545) );
  IV U3574 ( .A(n3061), .Z(n3063) );
  XNOR U3575 ( .A(b[514]), .B(n3061), .Z(n3062) );
  XOR U3576 ( .A(n3064), .B(n3065), .Z(n3061) );
  ANDN U3577 ( .B(n3066), .A(n546), .Z(n3064) );
  XNOR U3578 ( .A(a[513]), .B(n3067), .Z(n546) );
  IV U3579 ( .A(n3065), .Z(n3067) );
  XNOR U3580 ( .A(b[513]), .B(n3065), .Z(n3066) );
  XOR U3581 ( .A(n3068), .B(n3069), .Z(n3065) );
  ANDN U3582 ( .B(n3070), .A(n547), .Z(n3068) );
  XNOR U3583 ( .A(a[512]), .B(n3071), .Z(n547) );
  IV U3584 ( .A(n3069), .Z(n3071) );
  XNOR U3585 ( .A(b[512]), .B(n3069), .Z(n3070) );
  XOR U3586 ( .A(n3072), .B(n3073), .Z(n3069) );
  ANDN U3587 ( .B(n3074), .A(n548), .Z(n3072) );
  XNOR U3588 ( .A(a[511]), .B(n3075), .Z(n548) );
  IV U3589 ( .A(n3073), .Z(n3075) );
  XNOR U3590 ( .A(b[511]), .B(n3073), .Z(n3074) );
  XOR U3591 ( .A(n3076), .B(n3077), .Z(n3073) );
  ANDN U3592 ( .B(n3078), .A(n549), .Z(n3076) );
  XNOR U3593 ( .A(a[510]), .B(n3079), .Z(n549) );
  IV U3594 ( .A(n3077), .Z(n3079) );
  XNOR U3595 ( .A(b[510]), .B(n3077), .Z(n3078) );
  XOR U3596 ( .A(n3080), .B(n3081), .Z(n3077) );
  ANDN U3597 ( .B(n3082), .A(n551), .Z(n3080) );
  XNOR U3598 ( .A(a[509]), .B(n3083), .Z(n551) );
  IV U3599 ( .A(n3081), .Z(n3083) );
  XNOR U3600 ( .A(b[509]), .B(n3081), .Z(n3082) );
  XOR U3601 ( .A(n3084), .B(n3085), .Z(n3081) );
  ANDN U3602 ( .B(n3086), .A(n552), .Z(n3084) );
  XNOR U3603 ( .A(a[508]), .B(n3087), .Z(n552) );
  IV U3604 ( .A(n3085), .Z(n3087) );
  XNOR U3605 ( .A(b[508]), .B(n3085), .Z(n3086) );
  XOR U3606 ( .A(n3088), .B(n3089), .Z(n3085) );
  ANDN U3607 ( .B(n3090), .A(n553), .Z(n3088) );
  XNOR U3608 ( .A(a[507]), .B(n3091), .Z(n553) );
  IV U3609 ( .A(n3089), .Z(n3091) );
  XNOR U3610 ( .A(b[507]), .B(n3089), .Z(n3090) );
  XOR U3611 ( .A(n3092), .B(n3093), .Z(n3089) );
  ANDN U3612 ( .B(n3094), .A(n554), .Z(n3092) );
  XNOR U3613 ( .A(a[506]), .B(n3095), .Z(n554) );
  IV U3614 ( .A(n3093), .Z(n3095) );
  XNOR U3615 ( .A(b[506]), .B(n3093), .Z(n3094) );
  XOR U3616 ( .A(n3096), .B(n3097), .Z(n3093) );
  ANDN U3617 ( .B(n3098), .A(n555), .Z(n3096) );
  XNOR U3618 ( .A(a[505]), .B(n3099), .Z(n555) );
  IV U3619 ( .A(n3097), .Z(n3099) );
  XNOR U3620 ( .A(b[505]), .B(n3097), .Z(n3098) );
  XOR U3621 ( .A(n3100), .B(n3101), .Z(n3097) );
  ANDN U3622 ( .B(n3102), .A(n556), .Z(n3100) );
  XNOR U3623 ( .A(a[504]), .B(n3103), .Z(n556) );
  IV U3624 ( .A(n3101), .Z(n3103) );
  XNOR U3625 ( .A(b[504]), .B(n3101), .Z(n3102) );
  XOR U3626 ( .A(n3104), .B(n3105), .Z(n3101) );
  ANDN U3627 ( .B(n3106), .A(n557), .Z(n3104) );
  XNOR U3628 ( .A(a[503]), .B(n3107), .Z(n557) );
  IV U3629 ( .A(n3105), .Z(n3107) );
  XNOR U3630 ( .A(b[503]), .B(n3105), .Z(n3106) );
  XOR U3631 ( .A(n3108), .B(n3109), .Z(n3105) );
  ANDN U3632 ( .B(n3110), .A(n558), .Z(n3108) );
  XNOR U3633 ( .A(a[502]), .B(n3111), .Z(n558) );
  IV U3634 ( .A(n3109), .Z(n3111) );
  XNOR U3635 ( .A(b[502]), .B(n3109), .Z(n3110) );
  XOR U3636 ( .A(n3112), .B(n3113), .Z(n3109) );
  ANDN U3637 ( .B(n3114), .A(n559), .Z(n3112) );
  XNOR U3638 ( .A(a[501]), .B(n3115), .Z(n559) );
  IV U3639 ( .A(n3113), .Z(n3115) );
  XNOR U3640 ( .A(b[501]), .B(n3113), .Z(n3114) );
  XOR U3641 ( .A(n3116), .B(n3117), .Z(n3113) );
  ANDN U3642 ( .B(n3118), .A(n560), .Z(n3116) );
  XNOR U3643 ( .A(a[500]), .B(n3119), .Z(n560) );
  IV U3644 ( .A(n3117), .Z(n3119) );
  XNOR U3645 ( .A(b[500]), .B(n3117), .Z(n3118) );
  XOR U3646 ( .A(n3120), .B(n3121), .Z(n3117) );
  ANDN U3647 ( .B(n3122), .A(n563), .Z(n3120) );
  XNOR U3648 ( .A(a[499]), .B(n3123), .Z(n563) );
  IV U3649 ( .A(n3121), .Z(n3123) );
  XNOR U3650 ( .A(b[499]), .B(n3121), .Z(n3122) );
  XOR U3651 ( .A(n3124), .B(n3125), .Z(n3121) );
  ANDN U3652 ( .B(n3126), .A(n564), .Z(n3124) );
  XNOR U3653 ( .A(a[498]), .B(n3127), .Z(n564) );
  IV U3654 ( .A(n3125), .Z(n3127) );
  XNOR U3655 ( .A(b[498]), .B(n3125), .Z(n3126) );
  XOR U3656 ( .A(n3128), .B(n3129), .Z(n3125) );
  ANDN U3657 ( .B(n3130), .A(n565), .Z(n3128) );
  XNOR U3658 ( .A(a[497]), .B(n3131), .Z(n565) );
  IV U3659 ( .A(n3129), .Z(n3131) );
  XNOR U3660 ( .A(b[497]), .B(n3129), .Z(n3130) );
  XOR U3661 ( .A(n3132), .B(n3133), .Z(n3129) );
  ANDN U3662 ( .B(n3134), .A(n566), .Z(n3132) );
  XNOR U3663 ( .A(a[496]), .B(n3135), .Z(n566) );
  IV U3664 ( .A(n3133), .Z(n3135) );
  XNOR U3665 ( .A(b[496]), .B(n3133), .Z(n3134) );
  XOR U3666 ( .A(n3136), .B(n3137), .Z(n3133) );
  ANDN U3667 ( .B(n3138), .A(n567), .Z(n3136) );
  XNOR U3668 ( .A(a[495]), .B(n3139), .Z(n567) );
  IV U3669 ( .A(n3137), .Z(n3139) );
  XNOR U3670 ( .A(b[495]), .B(n3137), .Z(n3138) );
  XOR U3671 ( .A(n3140), .B(n3141), .Z(n3137) );
  ANDN U3672 ( .B(n3142), .A(n568), .Z(n3140) );
  XNOR U3673 ( .A(a[494]), .B(n3143), .Z(n568) );
  IV U3674 ( .A(n3141), .Z(n3143) );
  XNOR U3675 ( .A(b[494]), .B(n3141), .Z(n3142) );
  XOR U3676 ( .A(n3144), .B(n3145), .Z(n3141) );
  ANDN U3677 ( .B(n3146), .A(n569), .Z(n3144) );
  XNOR U3678 ( .A(a[493]), .B(n3147), .Z(n569) );
  IV U3679 ( .A(n3145), .Z(n3147) );
  XNOR U3680 ( .A(b[493]), .B(n3145), .Z(n3146) );
  XOR U3681 ( .A(n3148), .B(n3149), .Z(n3145) );
  ANDN U3682 ( .B(n3150), .A(n570), .Z(n3148) );
  XNOR U3683 ( .A(a[492]), .B(n3151), .Z(n570) );
  IV U3684 ( .A(n3149), .Z(n3151) );
  XNOR U3685 ( .A(b[492]), .B(n3149), .Z(n3150) );
  XOR U3686 ( .A(n3152), .B(n3153), .Z(n3149) );
  ANDN U3687 ( .B(n3154), .A(n571), .Z(n3152) );
  XNOR U3688 ( .A(a[491]), .B(n3155), .Z(n571) );
  IV U3689 ( .A(n3153), .Z(n3155) );
  XNOR U3690 ( .A(b[491]), .B(n3153), .Z(n3154) );
  XOR U3691 ( .A(n3156), .B(n3157), .Z(n3153) );
  ANDN U3692 ( .B(n3158), .A(n572), .Z(n3156) );
  XNOR U3693 ( .A(a[490]), .B(n3159), .Z(n572) );
  IV U3694 ( .A(n3157), .Z(n3159) );
  XNOR U3695 ( .A(b[490]), .B(n3157), .Z(n3158) );
  XOR U3696 ( .A(n3160), .B(n3161), .Z(n3157) );
  ANDN U3697 ( .B(n3162), .A(n574), .Z(n3160) );
  XNOR U3698 ( .A(a[489]), .B(n3163), .Z(n574) );
  IV U3699 ( .A(n3161), .Z(n3163) );
  XNOR U3700 ( .A(b[489]), .B(n3161), .Z(n3162) );
  XOR U3701 ( .A(n3164), .B(n3165), .Z(n3161) );
  ANDN U3702 ( .B(n3166), .A(n575), .Z(n3164) );
  XNOR U3703 ( .A(a[488]), .B(n3167), .Z(n575) );
  IV U3704 ( .A(n3165), .Z(n3167) );
  XNOR U3705 ( .A(b[488]), .B(n3165), .Z(n3166) );
  XOR U3706 ( .A(n3168), .B(n3169), .Z(n3165) );
  ANDN U3707 ( .B(n3170), .A(n576), .Z(n3168) );
  XNOR U3708 ( .A(a[487]), .B(n3171), .Z(n576) );
  IV U3709 ( .A(n3169), .Z(n3171) );
  XNOR U3710 ( .A(b[487]), .B(n3169), .Z(n3170) );
  XOR U3711 ( .A(n3172), .B(n3173), .Z(n3169) );
  ANDN U3712 ( .B(n3174), .A(n577), .Z(n3172) );
  XNOR U3713 ( .A(a[486]), .B(n3175), .Z(n577) );
  IV U3714 ( .A(n3173), .Z(n3175) );
  XNOR U3715 ( .A(b[486]), .B(n3173), .Z(n3174) );
  XOR U3716 ( .A(n3176), .B(n3177), .Z(n3173) );
  ANDN U3717 ( .B(n3178), .A(n578), .Z(n3176) );
  XNOR U3718 ( .A(a[485]), .B(n3179), .Z(n578) );
  IV U3719 ( .A(n3177), .Z(n3179) );
  XNOR U3720 ( .A(b[485]), .B(n3177), .Z(n3178) );
  XOR U3721 ( .A(n3180), .B(n3181), .Z(n3177) );
  ANDN U3722 ( .B(n3182), .A(n579), .Z(n3180) );
  XNOR U3723 ( .A(a[484]), .B(n3183), .Z(n579) );
  IV U3724 ( .A(n3181), .Z(n3183) );
  XNOR U3725 ( .A(b[484]), .B(n3181), .Z(n3182) );
  XOR U3726 ( .A(n3184), .B(n3185), .Z(n3181) );
  ANDN U3727 ( .B(n3186), .A(n580), .Z(n3184) );
  XNOR U3728 ( .A(a[483]), .B(n3187), .Z(n580) );
  IV U3729 ( .A(n3185), .Z(n3187) );
  XNOR U3730 ( .A(b[483]), .B(n3185), .Z(n3186) );
  XOR U3731 ( .A(n3188), .B(n3189), .Z(n3185) );
  ANDN U3732 ( .B(n3190), .A(n581), .Z(n3188) );
  XNOR U3733 ( .A(a[482]), .B(n3191), .Z(n581) );
  IV U3734 ( .A(n3189), .Z(n3191) );
  XNOR U3735 ( .A(b[482]), .B(n3189), .Z(n3190) );
  XOR U3736 ( .A(n3192), .B(n3193), .Z(n3189) );
  ANDN U3737 ( .B(n3194), .A(n582), .Z(n3192) );
  XNOR U3738 ( .A(a[481]), .B(n3195), .Z(n582) );
  IV U3739 ( .A(n3193), .Z(n3195) );
  XNOR U3740 ( .A(b[481]), .B(n3193), .Z(n3194) );
  XOR U3741 ( .A(n3196), .B(n3197), .Z(n3193) );
  ANDN U3742 ( .B(n3198), .A(n583), .Z(n3196) );
  XNOR U3743 ( .A(a[480]), .B(n3199), .Z(n583) );
  IV U3744 ( .A(n3197), .Z(n3199) );
  XNOR U3745 ( .A(b[480]), .B(n3197), .Z(n3198) );
  XOR U3746 ( .A(n3200), .B(n3201), .Z(n3197) );
  ANDN U3747 ( .B(n3202), .A(n585), .Z(n3200) );
  XNOR U3748 ( .A(a[479]), .B(n3203), .Z(n585) );
  IV U3749 ( .A(n3201), .Z(n3203) );
  XNOR U3750 ( .A(b[479]), .B(n3201), .Z(n3202) );
  XOR U3751 ( .A(n3204), .B(n3205), .Z(n3201) );
  ANDN U3752 ( .B(n3206), .A(n586), .Z(n3204) );
  XNOR U3753 ( .A(a[478]), .B(n3207), .Z(n586) );
  IV U3754 ( .A(n3205), .Z(n3207) );
  XNOR U3755 ( .A(b[478]), .B(n3205), .Z(n3206) );
  XOR U3756 ( .A(n3208), .B(n3209), .Z(n3205) );
  ANDN U3757 ( .B(n3210), .A(n587), .Z(n3208) );
  XNOR U3758 ( .A(a[477]), .B(n3211), .Z(n587) );
  IV U3759 ( .A(n3209), .Z(n3211) );
  XNOR U3760 ( .A(b[477]), .B(n3209), .Z(n3210) );
  XOR U3761 ( .A(n3212), .B(n3213), .Z(n3209) );
  ANDN U3762 ( .B(n3214), .A(n588), .Z(n3212) );
  XNOR U3763 ( .A(a[476]), .B(n3215), .Z(n588) );
  IV U3764 ( .A(n3213), .Z(n3215) );
  XNOR U3765 ( .A(b[476]), .B(n3213), .Z(n3214) );
  XOR U3766 ( .A(n3216), .B(n3217), .Z(n3213) );
  ANDN U3767 ( .B(n3218), .A(n589), .Z(n3216) );
  XNOR U3768 ( .A(a[475]), .B(n3219), .Z(n589) );
  IV U3769 ( .A(n3217), .Z(n3219) );
  XNOR U3770 ( .A(b[475]), .B(n3217), .Z(n3218) );
  XOR U3771 ( .A(n3220), .B(n3221), .Z(n3217) );
  ANDN U3772 ( .B(n3222), .A(n590), .Z(n3220) );
  XNOR U3773 ( .A(a[474]), .B(n3223), .Z(n590) );
  IV U3774 ( .A(n3221), .Z(n3223) );
  XNOR U3775 ( .A(b[474]), .B(n3221), .Z(n3222) );
  XOR U3776 ( .A(n3224), .B(n3225), .Z(n3221) );
  ANDN U3777 ( .B(n3226), .A(n591), .Z(n3224) );
  XNOR U3778 ( .A(a[473]), .B(n3227), .Z(n591) );
  IV U3779 ( .A(n3225), .Z(n3227) );
  XNOR U3780 ( .A(b[473]), .B(n3225), .Z(n3226) );
  XOR U3781 ( .A(n3228), .B(n3229), .Z(n3225) );
  ANDN U3782 ( .B(n3230), .A(n592), .Z(n3228) );
  XNOR U3783 ( .A(a[472]), .B(n3231), .Z(n592) );
  IV U3784 ( .A(n3229), .Z(n3231) );
  XNOR U3785 ( .A(b[472]), .B(n3229), .Z(n3230) );
  XOR U3786 ( .A(n3232), .B(n3233), .Z(n3229) );
  ANDN U3787 ( .B(n3234), .A(n593), .Z(n3232) );
  XNOR U3788 ( .A(a[471]), .B(n3235), .Z(n593) );
  IV U3789 ( .A(n3233), .Z(n3235) );
  XNOR U3790 ( .A(b[471]), .B(n3233), .Z(n3234) );
  XOR U3791 ( .A(n3236), .B(n3237), .Z(n3233) );
  ANDN U3792 ( .B(n3238), .A(n594), .Z(n3236) );
  XNOR U3793 ( .A(a[470]), .B(n3239), .Z(n594) );
  IV U3794 ( .A(n3237), .Z(n3239) );
  XNOR U3795 ( .A(b[470]), .B(n3237), .Z(n3238) );
  XOR U3796 ( .A(n3240), .B(n3241), .Z(n3237) );
  ANDN U3797 ( .B(n3242), .A(n596), .Z(n3240) );
  XNOR U3798 ( .A(a[469]), .B(n3243), .Z(n596) );
  IV U3799 ( .A(n3241), .Z(n3243) );
  XNOR U3800 ( .A(b[469]), .B(n3241), .Z(n3242) );
  XOR U3801 ( .A(n3244), .B(n3245), .Z(n3241) );
  ANDN U3802 ( .B(n3246), .A(n597), .Z(n3244) );
  XNOR U3803 ( .A(a[468]), .B(n3247), .Z(n597) );
  IV U3804 ( .A(n3245), .Z(n3247) );
  XNOR U3805 ( .A(b[468]), .B(n3245), .Z(n3246) );
  XOR U3806 ( .A(n3248), .B(n3249), .Z(n3245) );
  ANDN U3807 ( .B(n3250), .A(n598), .Z(n3248) );
  XNOR U3808 ( .A(a[467]), .B(n3251), .Z(n598) );
  IV U3809 ( .A(n3249), .Z(n3251) );
  XNOR U3810 ( .A(b[467]), .B(n3249), .Z(n3250) );
  XOR U3811 ( .A(n3252), .B(n3253), .Z(n3249) );
  ANDN U3812 ( .B(n3254), .A(n599), .Z(n3252) );
  XNOR U3813 ( .A(a[466]), .B(n3255), .Z(n599) );
  IV U3814 ( .A(n3253), .Z(n3255) );
  XNOR U3815 ( .A(b[466]), .B(n3253), .Z(n3254) );
  XOR U3816 ( .A(n3256), .B(n3257), .Z(n3253) );
  ANDN U3817 ( .B(n3258), .A(n600), .Z(n3256) );
  XNOR U3818 ( .A(a[465]), .B(n3259), .Z(n600) );
  IV U3819 ( .A(n3257), .Z(n3259) );
  XNOR U3820 ( .A(b[465]), .B(n3257), .Z(n3258) );
  XOR U3821 ( .A(n3260), .B(n3261), .Z(n3257) );
  ANDN U3822 ( .B(n3262), .A(n601), .Z(n3260) );
  XNOR U3823 ( .A(a[464]), .B(n3263), .Z(n601) );
  IV U3824 ( .A(n3261), .Z(n3263) );
  XNOR U3825 ( .A(b[464]), .B(n3261), .Z(n3262) );
  XOR U3826 ( .A(n3264), .B(n3265), .Z(n3261) );
  ANDN U3827 ( .B(n3266), .A(n602), .Z(n3264) );
  XNOR U3828 ( .A(a[463]), .B(n3267), .Z(n602) );
  IV U3829 ( .A(n3265), .Z(n3267) );
  XNOR U3830 ( .A(b[463]), .B(n3265), .Z(n3266) );
  XOR U3831 ( .A(n3268), .B(n3269), .Z(n3265) );
  ANDN U3832 ( .B(n3270), .A(n603), .Z(n3268) );
  XNOR U3833 ( .A(a[462]), .B(n3271), .Z(n603) );
  IV U3834 ( .A(n3269), .Z(n3271) );
  XNOR U3835 ( .A(b[462]), .B(n3269), .Z(n3270) );
  XOR U3836 ( .A(n3272), .B(n3273), .Z(n3269) );
  ANDN U3837 ( .B(n3274), .A(n604), .Z(n3272) );
  XNOR U3838 ( .A(a[461]), .B(n3275), .Z(n604) );
  IV U3839 ( .A(n3273), .Z(n3275) );
  XNOR U3840 ( .A(b[461]), .B(n3273), .Z(n3274) );
  XOR U3841 ( .A(n3276), .B(n3277), .Z(n3273) );
  ANDN U3842 ( .B(n3278), .A(n605), .Z(n3276) );
  XNOR U3843 ( .A(a[460]), .B(n3279), .Z(n605) );
  IV U3844 ( .A(n3277), .Z(n3279) );
  XNOR U3845 ( .A(b[460]), .B(n3277), .Z(n3278) );
  XOR U3846 ( .A(n3280), .B(n3281), .Z(n3277) );
  ANDN U3847 ( .B(n3282), .A(n607), .Z(n3280) );
  XNOR U3848 ( .A(a[459]), .B(n3283), .Z(n607) );
  IV U3849 ( .A(n3281), .Z(n3283) );
  XNOR U3850 ( .A(b[459]), .B(n3281), .Z(n3282) );
  XOR U3851 ( .A(n3284), .B(n3285), .Z(n3281) );
  ANDN U3852 ( .B(n3286), .A(n608), .Z(n3284) );
  XNOR U3853 ( .A(a[458]), .B(n3287), .Z(n608) );
  IV U3854 ( .A(n3285), .Z(n3287) );
  XNOR U3855 ( .A(b[458]), .B(n3285), .Z(n3286) );
  XOR U3856 ( .A(n3288), .B(n3289), .Z(n3285) );
  ANDN U3857 ( .B(n3290), .A(n609), .Z(n3288) );
  XNOR U3858 ( .A(a[457]), .B(n3291), .Z(n609) );
  IV U3859 ( .A(n3289), .Z(n3291) );
  XNOR U3860 ( .A(b[457]), .B(n3289), .Z(n3290) );
  XOR U3861 ( .A(n3292), .B(n3293), .Z(n3289) );
  ANDN U3862 ( .B(n3294), .A(n610), .Z(n3292) );
  XNOR U3863 ( .A(a[456]), .B(n3295), .Z(n610) );
  IV U3864 ( .A(n3293), .Z(n3295) );
  XNOR U3865 ( .A(b[456]), .B(n3293), .Z(n3294) );
  XOR U3866 ( .A(n3296), .B(n3297), .Z(n3293) );
  ANDN U3867 ( .B(n3298), .A(n611), .Z(n3296) );
  XNOR U3868 ( .A(a[455]), .B(n3299), .Z(n611) );
  IV U3869 ( .A(n3297), .Z(n3299) );
  XNOR U3870 ( .A(b[455]), .B(n3297), .Z(n3298) );
  XOR U3871 ( .A(n3300), .B(n3301), .Z(n3297) );
  ANDN U3872 ( .B(n3302), .A(n612), .Z(n3300) );
  XNOR U3873 ( .A(a[454]), .B(n3303), .Z(n612) );
  IV U3874 ( .A(n3301), .Z(n3303) );
  XNOR U3875 ( .A(b[454]), .B(n3301), .Z(n3302) );
  XOR U3876 ( .A(n3304), .B(n3305), .Z(n3301) );
  ANDN U3877 ( .B(n3306), .A(n613), .Z(n3304) );
  XNOR U3878 ( .A(a[453]), .B(n3307), .Z(n613) );
  IV U3879 ( .A(n3305), .Z(n3307) );
  XNOR U3880 ( .A(b[453]), .B(n3305), .Z(n3306) );
  XOR U3881 ( .A(n3308), .B(n3309), .Z(n3305) );
  ANDN U3882 ( .B(n3310), .A(n614), .Z(n3308) );
  XNOR U3883 ( .A(a[452]), .B(n3311), .Z(n614) );
  IV U3884 ( .A(n3309), .Z(n3311) );
  XNOR U3885 ( .A(b[452]), .B(n3309), .Z(n3310) );
  XOR U3886 ( .A(n3312), .B(n3313), .Z(n3309) );
  ANDN U3887 ( .B(n3314), .A(n615), .Z(n3312) );
  XNOR U3888 ( .A(a[451]), .B(n3315), .Z(n615) );
  IV U3889 ( .A(n3313), .Z(n3315) );
  XNOR U3890 ( .A(b[451]), .B(n3313), .Z(n3314) );
  XOR U3891 ( .A(n3316), .B(n3317), .Z(n3313) );
  ANDN U3892 ( .B(n3318), .A(n616), .Z(n3316) );
  XNOR U3893 ( .A(a[450]), .B(n3319), .Z(n616) );
  IV U3894 ( .A(n3317), .Z(n3319) );
  XNOR U3895 ( .A(b[450]), .B(n3317), .Z(n3318) );
  XOR U3896 ( .A(n3320), .B(n3321), .Z(n3317) );
  ANDN U3897 ( .B(n3322), .A(n618), .Z(n3320) );
  XNOR U3898 ( .A(a[449]), .B(n3323), .Z(n618) );
  IV U3899 ( .A(n3321), .Z(n3323) );
  XNOR U3900 ( .A(b[449]), .B(n3321), .Z(n3322) );
  XOR U3901 ( .A(n3324), .B(n3325), .Z(n3321) );
  ANDN U3902 ( .B(n3326), .A(n619), .Z(n3324) );
  XNOR U3903 ( .A(a[448]), .B(n3327), .Z(n619) );
  IV U3904 ( .A(n3325), .Z(n3327) );
  XNOR U3905 ( .A(b[448]), .B(n3325), .Z(n3326) );
  XOR U3906 ( .A(n3328), .B(n3329), .Z(n3325) );
  ANDN U3907 ( .B(n3330), .A(n620), .Z(n3328) );
  XNOR U3908 ( .A(a[447]), .B(n3331), .Z(n620) );
  IV U3909 ( .A(n3329), .Z(n3331) );
  XNOR U3910 ( .A(b[447]), .B(n3329), .Z(n3330) );
  XOR U3911 ( .A(n3332), .B(n3333), .Z(n3329) );
  ANDN U3912 ( .B(n3334), .A(n621), .Z(n3332) );
  XNOR U3913 ( .A(a[446]), .B(n3335), .Z(n621) );
  IV U3914 ( .A(n3333), .Z(n3335) );
  XNOR U3915 ( .A(b[446]), .B(n3333), .Z(n3334) );
  XOR U3916 ( .A(n3336), .B(n3337), .Z(n3333) );
  ANDN U3917 ( .B(n3338), .A(n622), .Z(n3336) );
  XNOR U3918 ( .A(a[445]), .B(n3339), .Z(n622) );
  IV U3919 ( .A(n3337), .Z(n3339) );
  XNOR U3920 ( .A(b[445]), .B(n3337), .Z(n3338) );
  XOR U3921 ( .A(n3340), .B(n3341), .Z(n3337) );
  ANDN U3922 ( .B(n3342), .A(n623), .Z(n3340) );
  XNOR U3923 ( .A(a[444]), .B(n3343), .Z(n623) );
  IV U3924 ( .A(n3341), .Z(n3343) );
  XNOR U3925 ( .A(b[444]), .B(n3341), .Z(n3342) );
  XOR U3926 ( .A(n3344), .B(n3345), .Z(n3341) );
  ANDN U3927 ( .B(n3346), .A(n624), .Z(n3344) );
  XNOR U3928 ( .A(a[443]), .B(n3347), .Z(n624) );
  IV U3929 ( .A(n3345), .Z(n3347) );
  XNOR U3930 ( .A(b[443]), .B(n3345), .Z(n3346) );
  XOR U3931 ( .A(n3348), .B(n3349), .Z(n3345) );
  ANDN U3932 ( .B(n3350), .A(n625), .Z(n3348) );
  XNOR U3933 ( .A(a[442]), .B(n3351), .Z(n625) );
  IV U3934 ( .A(n3349), .Z(n3351) );
  XNOR U3935 ( .A(b[442]), .B(n3349), .Z(n3350) );
  XOR U3936 ( .A(n3352), .B(n3353), .Z(n3349) );
  ANDN U3937 ( .B(n3354), .A(n626), .Z(n3352) );
  XNOR U3938 ( .A(a[441]), .B(n3355), .Z(n626) );
  IV U3939 ( .A(n3353), .Z(n3355) );
  XNOR U3940 ( .A(b[441]), .B(n3353), .Z(n3354) );
  XOR U3941 ( .A(n3356), .B(n3357), .Z(n3353) );
  ANDN U3942 ( .B(n3358), .A(n627), .Z(n3356) );
  XNOR U3943 ( .A(a[440]), .B(n3359), .Z(n627) );
  IV U3944 ( .A(n3357), .Z(n3359) );
  XNOR U3945 ( .A(b[440]), .B(n3357), .Z(n3358) );
  XOR U3946 ( .A(n3360), .B(n3361), .Z(n3357) );
  ANDN U3947 ( .B(n3362), .A(n629), .Z(n3360) );
  XNOR U3948 ( .A(a[439]), .B(n3363), .Z(n629) );
  IV U3949 ( .A(n3361), .Z(n3363) );
  XNOR U3950 ( .A(b[439]), .B(n3361), .Z(n3362) );
  XOR U3951 ( .A(n3364), .B(n3365), .Z(n3361) );
  ANDN U3952 ( .B(n3366), .A(n630), .Z(n3364) );
  XNOR U3953 ( .A(a[438]), .B(n3367), .Z(n630) );
  IV U3954 ( .A(n3365), .Z(n3367) );
  XNOR U3955 ( .A(b[438]), .B(n3365), .Z(n3366) );
  XOR U3956 ( .A(n3368), .B(n3369), .Z(n3365) );
  ANDN U3957 ( .B(n3370), .A(n631), .Z(n3368) );
  XNOR U3958 ( .A(a[437]), .B(n3371), .Z(n631) );
  IV U3959 ( .A(n3369), .Z(n3371) );
  XNOR U3960 ( .A(b[437]), .B(n3369), .Z(n3370) );
  XOR U3961 ( .A(n3372), .B(n3373), .Z(n3369) );
  ANDN U3962 ( .B(n3374), .A(n632), .Z(n3372) );
  XNOR U3963 ( .A(a[436]), .B(n3375), .Z(n632) );
  IV U3964 ( .A(n3373), .Z(n3375) );
  XNOR U3965 ( .A(b[436]), .B(n3373), .Z(n3374) );
  XOR U3966 ( .A(n3376), .B(n3377), .Z(n3373) );
  ANDN U3967 ( .B(n3378), .A(n633), .Z(n3376) );
  XNOR U3968 ( .A(a[435]), .B(n3379), .Z(n633) );
  IV U3969 ( .A(n3377), .Z(n3379) );
  XNOR U3970 ( .A(b[435]), .B(n3377), .Z(n3378) );
  XOR U3971 ( .A(n3380), .B(n3381), .Z(n3377) );
  ANDN U3972 ( .B(n3382), .A(n634), .Z(n3380) );
  XNOR U3973 ( .A(a[434]), .B(n3383), .Z(n634) );
  IV U3974 ( .A(n3381), .Z(n3383) );
  XNOR U3975 ( .A(b[434]), .B(n3381), .Z(n3382) );
  XOR U3976 ( .A(n3384), .B(n3385), .Z(n3381) );
  ANDN U3977 ( .B(n3386), .A(n635), .Z(n3384) );
  XNOR U3978 ( .A(a[433]), .B(n3387), .Z(n635) );
  IV U3979 ( .A(n3385), .Z(n3387) );
  XNOR U3980 ( .A(b[433]), .B(n3385), .Z(n3386) );
  XOR U3981 ( .A(n3388), .B(n3389), .Z(n3385) );
  ANDN U3982 ( .B(n3390), .A(n636), .Z(n3388) );
  XNOR U3983 ( .A(a[432]), .B(n3391), .Z(n636) );
  IV U3984 ( .A(n3389), .Z(n3391) );
  XNOR U3985 ( .A(b[432]), .B(n3389), .Z(n3390) );
  XOR U3986 ( .A(n3392), .B(n3393), .Z(n3389) );
  ANDN U3987 ( .B(n3394), .A(n637), .Z(n3392) );
  XNOR U3988 ( .A(a[431]), .B(n3395), .Z(n637) );
  IV U3989 ( .A(n3393), .Z(n3395) );
  XNOR U3990 ( .A(b[431]), .B(n3393), .Z(n3394) );
  XOR U3991 ( .A(n3396), .B(n3397), .Z(n3393) );
  ANDN U3992 ( .B(n3398), .A(n638), .Z(n3396) );
  XNOR U3993 ( .A(a[430]), .B(n3399), .Z(n638) );
  IV U3994 ( .A(n3397), .Z(n3399) );
  XNOR U3995 ( .A(b[430]), .B(n3397), .Z(n3398) );
  XOR U3996 ( .A(n3400), .B(n3401), .Z(n3397) );
  ANDN U3997 ( .B(n3402), .A(n640), .Z(n3400) );
  XNOR U3998 ( .A(a[429]), .B(n3403), .Z(n640) );
  IV U3999 ( .A(n3401), .Z(n3403) );
  XNOR U4000 ( .A(b[429]), .B(n3401), .Z(n3402) );
  XOR U4001 ( .A(n3404), .B(n3405), .Z(n3401) );
  ANDN U4002 ( .B(n3406), .A(n641), .Z(n3404) );
  XNOR U4003 ( .A(a[428]), .B(n3407), .Z(n641) );
  IV U4004 ( .A(n3405), .Z(n3407) );
  XNOR U4005 ( .A(b[428]), .B(n3405), .Z(n3406) );
  XOR U4006 ( .A(n3408), .B(n3409), .Z(n3405) );
  ANDN U4007 ( .B(n3410), .A(n642), .Z(n3408) );
  XNOR U4008 ( .A(a[427]), .B(n3411), .Z(n642) );
  IV U4009 ( .A(n3409), .Z(n3411) );
  XNOR U4010 ( .A(b[427]), .B(n3409), .Z(n3410) );
  XOR U4011 ( .A(n3412), .B(n3413), .Z(n3409) );
  ANDN U4012 ( .B(n3414), .A(n643), .Z(n3412) );
  XNOR U4013 ( .A(a[426]), .B(n3415), .Z(n643) );
  IV U4014 ( .A(n3413), .Z(n3415) );
  XNOR U4015 ( .A(b[426]), .B(n3413), .Z(n3414) );
  XOR U4016 ( .A(n3416), .B(n3417), .Z(n3413) );
  ANDN U4017 ( .B(n3418), .A(n644), .Z(n3416) );
  XNOR U4018 ( .A(a[425]), .B(n3419), .Z(n644) );
  IV U4019 ( .A(n3417), .Z(n3419) );
  XNOR U4020 ( .A(b[425]), .B(n3417), .Z(n3418) );
  XOR U4021 ( .A(n3420), .B(n3421), .Z(n3417) );
  ANDN U4022 ( .B(n3422), .A(n645), .Z(n3420) );
  XNOR U4023 ( .A(a[424]), .B(n3423), .Z(n645) );
  IV U4024 ( .A(n3421), .Z(n3423) );
  XNOR U4025 ( .A(b[424]), .B(n3421), .Z(n3422) );
  XOR U4026 ( .A(n3424), .B(n3425), .Z(n3421) );
  ANDN U4027 ( .B(n3426), .A(n646), .Z(n3424) );
  XNOR U4028 ( .A(a[423]), .B(n3427), .Z(n646) );
  IV U4029 ( .A(n3425), .Z(n3427) );
  XNOR U4030 ( .A(b[423]), .B(n3425), .Z(n3426) );
  XOR U4031 ( .A(n3428), .B(n3429), .Z(n3425) );
  ANDN U4032 ( .B(n3430), .A(n647), .Z(n3428) );
  XNOR U4033 ( .A(a[422]), .B(n3431), .Z(n647) );
  IV U4034 ( .A(n3429), .Z(n3431) );
  XNOR U4035 ( .A(b[422]), .B(n3429), .Z(n3430) );
  XOR U4036 ( .A(n3432), .B(n3433), .Z(n3429) );
  ANDN U4037 ( .B(n3434), .A(n648), .Z(n3432) );
  XNOR U4038 ( .A(a[421]), .B(n3435), .Z(n648) );
  IV U4039 ( .A(n3433), .Z(n3435) );
  XNOR U4040 ( .A(b[421]), .B(n3433), .Z(n3434) );
  XOR U4041 ( .A(n3436), .B(n3437), .Z(n3433) );
  ANDN U4042 ( .B(n3438), .A(n649), .Z(n3436) );
  XNOR U4043 ( .A(a[420]), .B(n3439), .Z(n649) );
  IV U4044 ( .A(n3437), .Z(n3439) );
  XNOR U4045 ( .A(b[420]), .B(n3437), .Z(n3438) );
  XOR U4046 ( .A(n3440), .B(n3441), .Z(n3437) );
  ANDN U4047 ( .B(n3442), .A(n651), .Z(n3440) );
  XNOR U4048 ( .A(a[419]), .B(n3443), .Z(n651) );
  IV U4049 ( .A(n3441), .Z(n3443) );
  XNOR U4050 ( .A(b[419]), .B(n3441), .Z(n3442) );
  XOR U4051 ( .A(n3444), .B(n3445), .Z(n3441) );
  ANDN U4052 ( .B(n3446), .A(n652), .Z(n3444) );
  XNOR U4053 ( .A(a[418]), .B(n3447), .Z(n652) );
  IV U4054 ( .A(n3445), .Z(n3447) );
  XNOR U4055 ( .A(b[418]), .B(n3445), .Z(n3446) );
  XOR U4056 ( .A(n3448), .B(n3449), .Z(n3445) );
  ANDN U4057 ( .B(n3450), .A(n653), .Z(n3448) );
  XNOR U4058 ( .A(a[417]), .B(n3451), .Z(n653) );
  IV U4059 ( .A(n3449), .Z(n3451) );
  XNOR U4060 ( .A(b[417]), .B(n3449), .Z(n3450) );
  XOR U4061 ( .A(n3452), .B(n3453), .Z(n3449) );
  ANDN U4062 ( .B(n3454), .A(n654), .Z(n3452) );
  XNOR U4063 ( .A(a[416]), .B(n3455), .Z(n654) );
  IV U4064 ( .A(n3453), .Z(n3455) );
  XNOR U4065 ( .A(b[416]), .B(n3453), .Z(n3454) );
  XOR U4066 ( .A(n3456), .B(n3457), .Z(n3453) );
  ANDN U4067 ( .B(n3458), .A(n655), .Z(n3456) );
  XNOR U4068 ( .A(a[415]), .B(n3459), .Z(n655) );
  IV U4069 ( .A(n3457), .Z(n3459) );
  XNOR U4070 ( .A(b[415]), .B(n3457), .Z(n3458) );
  XOR U4071 ( .A(n3460), .B(n3461), .Z(n3457) );
  ANDN U4072 ( .B(n3462), .A(n656), .Z(n3460) );
  XNOR U4073 ( .A(a[414]), .B(n3463), .Z(n656) );
  IV U4074 ( .A(n3461), .Z(n3463) );
  XNOR U4075 ( .A(b[414]), .B(n3461), .Z(n3462) );
  XOR U4076 ( .A(n3464), .B(n3465), .Z(n3461) );
  ANDN U4077 ( .B(n3466), .A(n657), .Z(n3464) );
  XNOR U4078 ( .A(a[413]), .B(n3467), .Z(n657) );
  IV U4079 ( .A(n3465), .Z(n3467) );
  XNOR U4080 ( .A(b[413]), .B(n3465), .Z(n3466) );
  XOR U4081 ( .A(n3468), .B(n3469), .Z(n3465) );
  ANDN U4082 ( .B(n3470), .A(n658), .Z(n3468) );
  XNOR U4083 ( .A(a[412]), .B(n3471), .Z(n658) );
  IV U4084 ( .A(n3469), .Z(n3471) );
  XNOR U4085 ( .A(b[412]), .B(n3469), .Z(n3470) );
  XOR U4086 ( .A(n3472), .B(n3473), .Z(n3469) );
  ANDN U4087 ( .B(n3474), .A(n659), .Z(n3472) );
  XNOR U4088 ( .A(a[411]), .B(n3475), .Z(n659) );
  IV U4089 ( .A(n3473), .Z(n3475) );
  XNOR U4090 ( .A(b[411]), .B(n3473), .Z(n3474) );
  XOR U4091 ( .A(n3476), .B(n3477), .Z(n3473) );
  ANDN U4092 ( .B(n3478), .A(n660), .Z(n3476) );
  XNOR U4093 ( .A(a[410]), .B(n3479), .Z(n660) );
  IV U4094 ( .A(n3477), .Z(n3479) );
  XNOR U4095 ( .A(b[410]), .B(n3477), .Z(n3478) );
  XOR U4096 ( .A(n3480), .B(n3481), .Z(n3477) );
  ANDN U4097 ( .B(n3482), .A(n662), .Z(n3480) );
  XNOR U4098 ( .A(a[409]), .B(n3483), .Z(n662) );
  IV U4099 ( .A(n3481), .Z(n3483) );
  XNOR U4100 ( .A(b[409]), .B(n3481), .Z(n3482) );
  XOR U4101 ( .A(n3484), .B(n3485), .Z(n3481) );
  ANDN U4102 ( .B(n3486), .A(n663), .Z(n3484) );
  XNOR U4103 ( .A(a[408]), .B(n3487), .Z(n663) );
  IV U4104 ( .A(n3485), .Z(n3487) );
  XNOR U4105 ( .A(b[408]), .B(n3485), .Z(n3486) );
  XOR U4106 ( .A(n3488), .B(n3489), .Z(n3485) );
  ANDN U4107 ( .B(n3490), .A(n664), .Z(n3488) );
  XNOR U4108 ( .A(a[407]), .B(n3491), .Z(n664) );
  IV U4109 ( .A(n3489), .Z(n3491) );
  XNOR U4110 ( .A(b[407]), .B(n3489), .Z(n3490) );
  XOR U4111 ( .A(n3492), .B(n3493), .Z(n3489) );
  ANDN U4112 ( .B(n3494), .A(n665), .Z(n3492) );
  XNOR U4113 ( .A(a[406]), .B(n3495), .Z(n665) );
  IV U4114 ( .A(n3493), .Z(n3495) );
  XNOR U4115 ( .A(b[406]), .B(n3493), .Z(n3494) );
  XOR U4116 ( .A(n3496), .B(n3497), .Z(n3493) );
  ANDN U4117 ( .B(n3498), .A(n666), .Z(n3496) );
  XNOR U4118 ( .A(a[405]), .B(n3499), .Z(n666) );
  IV U4119 ( .A(n3497), .Z(n3499) );
  XNOR U4120 ( .A(b[405]), .B(n3497), .Z(n3498) );
  XOR U4121 ( .A(n3500), .B(n3501), .Z(n3497) );
  ANDN U4122 ( .B(n3502), .A(n667), .Z(n3500) );
  XNOR U4123 ( .A(a[404]), .B(n3503), .Z(n667) );
  IV U4124 ( .A(n3501), .Z(n3503) );
  XNOR U4125 ( .A(b[404]), .B(n3501), .Z(n3502) );
  XOR U4126 ( .A(n3504), .B(n3505), .Z(n3501) );
  ANDN U4127 ( .B(n3506), .A(n668), .Z(n3504) );
  XNOR U4128 ( .A(a[403]), .B(n3507), .Z(n668) );
  IV U4129 ( .A(n3505), .Z(n3507) );
  XNOR U4130 ( .A(b[403]), .B(n3505), .Z(n3506) );
  XOR U4131 ( .A(n3508), .B(n3509), .Z(n3505) );
  ANDN U4132 ( .B(n3510), .A(n669), .Z(n3508) );
  XNOR U4133 ( .A(a[402]), .B(n3511), .Z(n669) );
  IV U4134 ( .A(n3509), .Z(n3511) );
  XNOR U4135 ( .A(b[402]), .B(n3509), .Z(n3510) );
  XOR U4136 ( .A(n3512), .B(n3513), .Z(n3509) );
  ANDN U4137 ( .B(n3514), .A(n670), .Z(n3512) );
  XNOR U4138 ( .A(a[401]), .B(n3515), .Z(n670) );
  IV U4139 ( .A(n3513), .Z(n3515) );
  XNOR U4140 ( .A(b[401]), .B(n3513), .Z(n3514) );
  XOR U4141 ( .A(n3516), .B(n3517), .Z(n3513) );
  ANDN U4142 ( .B(n3518), .A(n671), .Z(n3516) );
  XNOR U4143 ( .A(a[400]), .B(n3519), .Z(n671) );
  IV U4144 ( .A(n3517), .Z(n3519) );
  XNOR U4145 ( .A(b[400]), .B(n3517), .Z(n3518) );
  XOR U4146 ( .A(n3520), .B(n3521), .Z(n3517) );
  ANDN U4147 ( .B(n3522), .A(n674), .Z(n3520) );
  XNOR U4148 ( .A(a[399]), .B(n3523), .Z(n674) );
  IV U4149 ( .A(n3521), .Z(n3523) );
  XNOR U4150 ( .A(b[399]), .B(n3521), .Z(n3522) );
  XOR U4151 ( .A(n3524), .B(n3525), .Z(n3521) );
  ANDN U4152 ( .B(n3526), .A(n675), .Z(n3524) );
  XNOR U4153 ( .A(a[398]), .B(n3527), .Z(n675) );
  IV U4154 ( .A(n3525), .Z(n3527) );
  XNOR U4155 ( .A(b[398]), .B(n3525), .Z(n3526) );
  XOR U4156 ( .A(n3528), .B(n3529), .Z(n3525) );
  ANDN U4157 ( .B(n3530), .A(n676), .Z(n3528) );
  XNOR U4158 ( .A(a[397]), .B(n3531), .Z(n676) );
  IV U4159 ( .A(n3529), .Z(n3531) );
  XNOR U4160 ( .A(b[397]), .B(n3529), .Z(n3530) );
  XOR U4161 ( .A(n3532), .B(n3533), .Z(n3529) );
  ANDN U4162 ( .B(n3534), .A(n677), .Z(n3532) );
  XNOR U4163 ( .A(a[396]), .B(n3535), .Z(n677) );
  IV U4164 ( .A(n3533), .Z(n3535) );
  XNOR U4165 ( .A(b[396]), .B(n3533), .Z(n3534) );
  XOR U4166 ( .A(n3536), .B(n3537), .Z(n3533) );
  ANDN U4167 ( .B(n3538), .A(n678), .Z(n3536) );
  XNOR U4168 ( .A(a[395]), .B(n3539), .Z(n678) );
  IV U4169 ( .A(n3537), .Z(n3539) );
  XNOR U4170 ( .A(b[395]), .B(n3537), .Z(n3538) );
  XOR U4171 ( .A(n3540), .B(n3541), .Z(n3537) );
  ANDN U4172 ( .B(n3542), .A(n679), .Z(n3540) );
  XNOR U4173 ( .A(a[394]), .B(n3543), .Z(n679) );
  IV U4174 ( .A(n3541), .Z(n3543) );
  XNOR U4175 ( .A(b[394]), .B(n3541), .Z(n3542) );
  XOR U4176 ( .A(n3544), .B(n3545), .Z(n3541) );
  ANDN U4177 ( .B(n3546), .A(n680), .Z(n3544) );
  XNOR U4178 ( .A(a[393]), .B(n3547), .Z(n680) );
  IV U4179 ( .A(n3545), .Z(n3547) );
  XNOR U4180 ( .A(b[393]), .B(n3545), .Z(n3546) );
  XOR U4181 ( .A(n3548), .B(n3549), .Z(n3545) );
  ANDN U4182 ( .B(n3550), .A(n681), .Z(n3548) );
  XNOR U4183 ( .A(a[392]), .B(n3551), .Z(n681) );
  IV U4184 ( .A(n3549), .Z(n3551) );
  XNOR U4185 ( .A(b[392]), .B(n3549), .Z(n3550) );
  XOR U4186 ( .A(n3552), .B(n3553), .Z(n3549) );
  ANDN U4187 ( .B(n3554), .A(n682), .Z(n3552) );
  XNOR U4188 ( .A(a[391]), .B(n3555), .Z(n682) );
  IV U4189 ( .A(n3553), .Z(n3555) );
  XNOR U4190 ( .A(b[391]), .B(n3553), .Z(n3554) );
  XOR U4191 ( .A(n3556), .B(n3557), .Z(n3553) );
  ANDN U4192 ( .B(n3558), .A(n683), .Z(n3556) );
  XNOR U4193 ( .A(a[390]), .B(n3559), .Z(n683) );
  IV U4194 ( .A(n3557), .Z(n3559) );
  XNOR U4195 ( .A(b[390]), .B(n3557), .Z(n3558) );
  XOR U4196 ( .A(n3560), .B(n3561), .Z(n3557) );
  ANDN U4197 ( .B(n3562), .A(n685), .Z(n3560) );
  XNOR U4198 ( .A(a[389]), .B(n3563), .Z(n685) );
  IV U4199 ( .A(n3561), .Z(n3563) );
  XNOR U4200 ( .A(b[389]), .B(n3561), .Z(n3562) );
  XOR U4201 ( .A(n3564), .B(n3565), .Z(n3561) );
  ANDN U4202 ( .B(n3566), .A(n686), .Z(n3564) );
  XNOR U4203 ( .A(a[388]), .B(n3567), .Z(n686) );
  IV U4204 ( .A(n3565), .Z(n3567) );
  XNOR U4205 ( .A(b[388]), .B(n3565), .Z(n3566) );
  XOR U4206 ( .A(n3568), .B(n3569), .Z(n3565) );
  ANDN U4207 ( .B(n3570), .A(n687), .Z(n3568) );
  XNOR U4208 ( .A(a[387]), .B(n3571), .Z(n687) );
  IV U4209 ( .A(n3569), .Z(n3571) );
  XNOR U4210 ( .A(b[387]), .B(n3569), .Z(n3570) );
  XOR U4211 ( .A(n3572), .B(n3573), .Z(n3569) );
  ANDN U4212 ( .B(n3574), .A(n688), .Z(n3572) );
  XNOR U4213 ( .A(a[386]), .B(n3575), .Z(n688) );
  IV U4214 ( .A(n3573), .Z(n3575) );
  XNOR U4215 ( .A(b[386]), .B(n3573), .Z(n3574) );
  XOR U4216 ( .A(n3576), .B(n3577), .Z(n3573) );
  ANDN U4217 ( .B(n3578), .A(n689), .Z(n3576) );
  XNOR U4218 ( .A(a[385]), .B(n3579), .Z(n689) );
  IV U4219 ( .A(n3577), .Z(n3579) );
  XNOR U4220 ( .A(b[385]), .B(n3577), .Z(n3578) );
  XOR U4221 ( .A(n3580), .B(n3581), .Z(n3577) );
  ANDN U4222 ( .B(n3582), .A(n690), .Z(n3580) );
  XNOR U4223 ( .A(a[384]), .B(n3583), .Z(n690) );
  IV U4224 ( .A(n3581), .Z(n3583) );
  XNOR U4225 ( .A(b[384]), .B(n3581), .Z(n3582) );
  XOR U4226 ( .A(n3584), .B(n3585), .Z(n3581) );
  ANDN U4227 ( .B(n3586), .A(n691), .Z(n3584) );
  XNOR U4228 ( .A(a[383]), .B(n3587), .Z(n691) );
  IV U4229 ( .A(n3585), .Z(n3587) );
  XNOR U4230 ( .A(b[383]), .B(n3585), .Z(n3586) );
  XOR U4231 ( .A(n3588), .B(n3589), .Z(n3585) );
  ANDN U4232 ( .B(n3590), .A(n692), .Z(n3588) );
  XNOR U4233 ( .A(a[382]), .B(n3591), .Z(n692) );
  IV U4234 ( .A(n3589), .Z(n3591) );
  XNOR U4235 ( .A(b[382]), .B(n3589), .Z(n3590) );
  XOR U4236 ( .A(n3592), .B(n3593), .Z(n3589) );
  ANDN U4237 ( .B(n3594), .A(n693), .Z(n3592) );
  XNOR U4238 ( .A(a[381]), .B(n3595), .Z(n693) );
  IV U4239 ( .A(n3593), .Z(n3595) );
  XNOR U4240 ( .A(b[381]), .B(n3593), .Z(n3594) );
  XOR U4241 ( .A(n3596), .B(n3597), .Z(n3593) );
  ANDN U4242 ( .B(n3598), .A(n694), .Z(n3596) );
  XNOR U4243 ( .A(a[380]), .B(n3599), .Z(n694) );
  IV U4244 ( .A(n3597), .Z(n3599) );
  XNOR U4245 ( .A(b[380]), .B(n3597), .Z(n3598) );
  XOR U4246 ( .A(n3600), .B(n3601), .Z(n3597) );
  ANDN U4247 ( .B(n3602), .A(n696), .Z(n3600) );
  XNOR U4248 ( .A(a[379]), .B(n3603), .Z(n696) );
  IV U4249 ( .A(n3601), .Z(n3603) );
  XNOR U4250 ( .A(b[379]), .B(n3601), .Z(n3602) );
  XOR U4251 ( .A(n3604), .B(n3605), .Z(n3601) );
  ANDN U4252 ( .B(n3606), .A(n697), .Z(n3604) );
  XNOR U4253 ( .A(a[378]), .B(n3607), .Z(n697) );
  IV U4254 ( .A(n3605), .Z(n3607) );
  XNOR U4255 ( .A(b[378]), .B(n3605), .Z(n3606) );
  XOR U4256 ( .A(n3608), .B(n3609), .Z(n3605) );
  ANDN U4257 ( .B(n3610), .A(n698), .Z(n3608) );
  XNOR U4258 ( .A(a[377]), .B(n3611), .Z(n698) );
  IV U4259 ( .A(n3609), .Z(n3611) );
  XNOR U4260 ( .A(b[377]), .B(n3609), .Z(n3610) );
  XOR U4261 ( .A(n3612), .B(n3613), .Z(n3609) );
  ANDN U4262 ( .B(n3614), .A(n699), .Z(n3612) );
  XNOR U4263 ( .A(a[376]), .B(n3615), .Z(n699) );
  IV U4264 ( .A(n3613), .Z(n3615) );
  XNOR U4265 ( .A(b[376]), .B(n3613), .Z(n3614) );
  XOR U4266 ( .A(n3616), .B(n3617), .Z(n3613) );
  ANDN U4267 ( .B(n3618), .A(n700), .Z(n3616) );
  XNOR U4268 ( .A(a[375]), .B(n3619), .Z(n700) );
  IV U4269 ( .A(n3617), .Z(n3619) );
  XNOR U4270 ( .A(b[375]), .B(n3617), .Z(n3618) );
  XOR U4271 ( .A(n3620), .B(n3621), .Z(n3617) );
  ANDN U4272 ( .B(n3622), .A(n701), .Z(n3620) );
  XNOR U4273 ( .A(a[374]), .B(n3623), .Z(n701) );
  IV U4274 ( .A(n3621), .Z(n3623) );
  XNOR U4275 ( .A(b[374]), .B(n3621), .Z(n3622) );
  XOR U4276 ( .A(n3624), .B(n3625), .Z(n3621) );
  ANDN U4277 ( .B(n3626), .A(n702), .Z(n3624) );
  XNOR U4278 ( .A(a[373]), .B(n3627), .Z(n702) );
  IV U4279 ( .A(n3625), .Z(n3627) );
  XNOR U4280 ( .A(b[373]), .B(n3625), .Z(n3626) );
  XOR U4281 ( .A(n3628), .B(n3629), .Z(n3625) );
  ANDN U4282 ( .B(n3630), .A(n703), .Z(n3628) );
  XNOR U4283 ( .A(a[372]), .B(n3631), .Z(n703) );
  IV U4284 ( .A(n3629), .Z(n3631) );
  XNOR U4285 ( .A(b[372]), .B(n3629), .Z(n3630) );
  XOR U4286 ( .A(n3632), .B(n3633), .Z(n3629) );
  ANDN U4287 ( .B(n3634), .A(n704), .Z(n3632) );
  XNOR U4288 ( .A(a[371]), .B(n3635), .Z(n704) );
  IV U4289 ( .A(n3633), .Z(n3635) );
  XNOR U4290 ( .A(b[371]), .B(n3633), .Z(n3634) );
  XOR U4291 ( .A(n3636), .B(n3637), .Z(n3633) );
  ANDN U4292 ( .B(n3638), .A(n705), .Z(n3636) );
  XNOR U4293 ( .A(a[370]), .B(n3639), .Z(n705) );
  IV U4294 ( .A(n3637), .Z(n3639) );
  XNOR U4295 ( .A(b[370]), .B(n3637), .Z(n3638) );
  XOR U4296 ( .A(n3640), .B(n3641), .Z(n3637) );
  ANDN U4297 ( .B(n3642), .A(n707), .Z(n3640) );
  XNOR U4298 ( .A(a[369]), .B(n3643), .Z(n707) );
  IV U4299 ( .A(n3641), .Z(n3643) );
  XNOR U4300 ( .A(b[369]), .B(n3641), .Z(n3642) );
  XOR U4301 ( .A(n3644), .B(n3645), .Z(n3641) );
  ANDN U4302 ( .B(n3646), .A(n708), .Z(n3644) );
  XNOR U4303 ( .A(a[368]), .B(n3647), .Z(n708) );
  IV U4304 ( .A(n3645), .Z(n3647) );
  XNOR U4305 ( .A(b[368]), .B(n3645), .Z(n3646) );
  XOR U4306 ( .A(n3648), .B(n3649), .Z(n3645) );
  ANDN U4307 ( .B(n3650), .A(n709), .Z(n3648) );
  XNOR U4308 ( .A(a[367]), .B(n3651), .Z(n709) );
  IV U4309 ( .A(n3649), .Z(n3651) );
  XNOR U4310 ( .A(b[367]), .B(n3649), .Z(n3650) );
  XOR U4311 ( .A(n3652), .B(n3653), .Z(n3649) );
  ANDN U4312 ( .B(n3654), .A(n710), .Z(n3652) );
  XNOR U4313 ( .A(a[366]), .B(n3655), .Z(n710) );
  IV U4314 ( .A(n3653), .Z(n3655) );
  XNOR U4315 ( .A(b[366]), .B(n3653), .Z(n3654) );
  XOR U4316 ( .A(n3656), .B(n3657), .Z(n3653) );
  ANDN U4317 ( .B(n3658), .A(n711), .Z(n3656) );
  XNOR U4318 ( .A(a[365]), .B(n3659), .Z(n711) );
  IV U4319 ( .A(n3657), .Z(n3659) );
  XNOR U4320 ( .A(b[365]), .B(n3657), .Z(n3658) );
  XOR U4321 ( .A(n3660), .B(n3661), .Z(n3657) );
  ANDN U4322 ( .B(n3662), .A(n712), .Z(n3660) );
  XNOR U4323 ( .A(a[364]), .B(n3663), .Z(n712) );
  IV U4324 ( .A(n3661), .Z(n3663) );
  XNOR U4325 ( .A(b[364]), .B(n3661), .Z(n3662) );
  XOR U4326 ( .A(n3664), .B(n3665), .Z(n3661) );
  ANDN U4327 ( .B(n3666), .A(n713), .Z(n3664) );
  XNOR U4328 ( .A(a[363]), .B(n3667), .Z(n713) );
  IV U4329 ( .A(n3665), .Z(n3667) );
  XNOR U4330 ( .A(b[363]), .B(n3665), .Z(n3666) );
  XOR U4331 ( .A(n3668), .B(n3669), .Z(n3665) );
  ANDN U4332 ( .B(n3670), .A(n714), .Z(n3668) );
  XNOR U4333 ( .A(a[362]), .B(n3671), .Z(n714) );
  IV U4334 ( .A(n3669), .Z(n3671) );
  XNOR U4335 ( .A(b[362]), .B(n3669), .Z(n3670) );
  XOR U4336 ( .A(n3672), .B(n3673), .Z(n3669) );
  ANDN U4337 ( .B(n3674), .A(n715), .Z(n3672) );
  XNOR U4338 ( .A(a[361]), .B(n3675), .Z(n715) );
  IV U4339 ( .A(n3673), .Z(n3675) );
  XNOR U4340 ( .A(b[361]), .B(n3673), .Z(n3674) );
  XOR U4341 ( .A(n3676), .B(n3677), .Z(n3673) );
  ANDN U4342 ( .B(n3678), .A(n716), .Z(n3676) );
  XNOR U4343 ( .A(a[360]), .B(n3679), .Z(n716) );
  IV U4344 ( .A(n3677), .Z(n3679) );
  XNOR U4345 ( .A(b[360]), .B(n3677), .Z(n3678) );
  XOR U4346 ( .A(n3680), .B(n3681), .Z(n3677) );
  ANDN U4347 ( .B(n3682), .A(n718), .Z(n3680) );
  XNOR U4348 ( .A(a[359]), .B(n3683), .Z(n718) );
  IV U4349 ( .A(n3681), .Z(n3683) );
  XNOR U4350 ( .A(b[359]), .B(n3681), .Z(n3682) );
  XOR U4351 ( .A(n3684), .B(n3685), .Z(n3681) );
  ANDN U4352 ( .B(n3686), .A(n719), .Z(n3684) );
  XNOR U4353 ( .A(a[358]), .B(n3687), .Z(n719) );
  IV U4354 ( .A(n3685), .Z(n3687) );
  XNOR U4355 ( .A(b[358]), .B(n3685), .Z(n3686) );
  XOR U4356 ( .A(n3688), .B(n3689), .Z(n3685) );
  ANDN U4357 ( .B(n3690), .A(n720), .Z(n3688) );
  XNOR U4358 ( .A(a[357]), .B(n3691), .Z(n720) );
  IV U4359 ( .A(n3689), .Z(n3691) );
  XNOR U4360 ( .A(b[357]), .B(n3689), .Z(n3690) );
  XOR U4361 ( .A(n3692), .B(n3693), .Z(n3689) );
  ANDN U4362 ( .B(n3694), .A(n721), .Z(n3692) );
  XNOR U4363 ( .A(a[356]), .B(n3695), .Z(n721) );
  IV U4364 ( .A(n3693), .Z(n3695) );
  XNOR U4365 ( .A(b[356]), .B(n3693), .Z(n3694) );
  XOR U4366 ( .A(n3696), .B(n3697), .Z(n3693) );
  ANDN U4367 ( .B(n3698), .A(n722), .Z(n3696) );
  XNOR U4368 ( .A(a[355]), .B(n3699), .Z(n722) );
  IV U4369 ( .A(n3697), .Z(n3699) );
  XNOR U4370 ( .A(b[355]), .B(n3697), .Z(n3698) );
  XOR U4371 ( .A(n3700), .B(n3701), .Z(n3697) );
  ANDN U4372 ( .B(n3702), .A(n723), .Z(n3700) );
  XNOR U4373 ( .A(a[354]), .B(n3703), .Z(n723) );
  IV U4374 ( .A(n3701), .Z(n3703) );
  XNOR U4375 ( .A(b[354]), .B(n3701), .Z(n3702) );
  XOR U4376 ( .A(n3704), .B(n3705), .Z(n3701) );
  ANDN U4377 ( .B(n3706), .A(n724), .Z(n3704) );
  XNOR U4378 ( .A(a[353]), .B(n3707), .Z(n724) );
  IV U4379 ( .A(n3705), .Z(n3707) );
  XNOR U4380 ( .A(b[353]), .B(n3705), .Z(n3706) );
  XOR U4381 ( .A(n3708), .B(n3709), .Z(n3705) );
  ANDN U4382 ( .B(n3710), .A(n725), .Z(n3708) );
  XNOR U4383 ( .A(a[352]), .B(n3711), .Z(n725) );
  IV U4384 ( .A(n3709), .Z(n3711) );
  XNOR U4385 ( .A(b[352]), .B(n3709), .Z(n3710) );
  XOR U4386 ( .A(n3712), .B(n3713), .Z(n3709) );
  ANDN U4387 ( .B(n3714), .A(n726), .Z(n3712) );
  XNOR U4388 ( .A(a[351]), .B(n3715), .Z(n726) );
  IV U4389 ( .A(n3713), .Z(n3715) );
  XNOR U4390 ( .A(b[351]), .B(n3713), .Z(n3714) );
  XOR U4391 ( .A(n3716), .B(n3717), .Z(n3713) );
  ANDN U4392 ( .B(n3718), .A(n727), .Z(n3716) );
  XNOR U4393 ( .A(a[350]), .B(n3719), .Z(n727) );
  IV U4394 ( .A(n3717), .Z(n3719) );
  XNOR U4395 ( .A(b[350]), .B(n3717), .Z(n3718) );
  XOR U4396 ( .A(n3720), .B(n3721), .Z(n3717) );
  ANDN U4397 ( .B(n3722), .A(n729), .Z(n3720) );
  XNOR U4398 ( .A(a[349]), .B(n3723), .Z(n729) );
  IV U4399 ( .A(n3721), .Z(n3723) );
  XNOR U4400 ( .A(b[349]), .B(n3721), .Z(n3722) );
  XOR U4401 ( .A(n3724), .B(n3725), .Z(n3721) );
  ANDN U4402 ( .B(n3726), .A(n730), .Z(n3724) );
  XNOR U4403 ( .A(a[348]), .B(n3727), .Z(n730) );
  IV U4404 ( .A(n3725), .Z(n3727) );
  XNOR U4405 ( .A(b[348]), .B(n3725), .Z(n3726) );
  XOR U4406 ( .A(n3728), .B(n3729), .Z(n3725) );
  ANDN U4407 ( .B(n3730), .A(n731), .Z(n3728) );
  XNOR U4408 ( .A(a[347]), .B(n3731), .Z(n731) );
  IV U4409 ( .A(n3729), .Z(n3731) );
  XNOR U4410 ( .A(b[347]), .B(n3729), .Z(n3730) );
  XOR U4411 ( .A(n3732), .B(n3733), .Z(n3729) );
  ANDN U4412 ( .B(n3734), .A(n732), .Z(n3732) );
  XNOR U4413 ( .A(a[346]), .B(n3735), .Z(n732) );
  IV U4414 ( .A(n3733), .Z(n3735) );
  XNOR U4415 ( .A(b[346]), .B(n3733), .Z(n3734) );
  XOR U4416 ( .A(n3736), .B(n3737), .Z(n3733) );
  ANDN U4417 ( .B(n3738), .A(n733), .Z(n3736) );
  XNOR U4418 ( .A(a[345]), .B(n3739), .Z(n733) );
  IV U4419 ( .A(n3737), .Z(n3739) );
  XNOR U4420 ( .A(b[345]), .B(n3737), .Z(n3738) );
  XOR U4421 ( .A(n3740), .B(n3741), .Z(n3737) );
  ANDN U4422 ( .B(n3742), .A(n734), .Z(n3740) );
  XNOR U4423 ( .A(a[344]), .B(n3743), .Z(n734) );
  IV U4424 ( .A(n3741), .Z(n3743) );
  XNOR U4425 ( .A(b[344]), .B(n3741), .Z(n3742) );
  XOR U4426 ( .A(n3744), .B(n3745), .Z(n3741) );
  ANDN U4427 ( .B(n3746), .A(n735), .Z(n3744) );
  XNOR U4428 ( .A(a[343]), .B(n3747), .Z(n735) );
  IV U4429 ( .A(n3745), .Z(n3747) );
  XNOR U4430 ( .A(b[343]), .B(n3745), .Z(n3746) );
  XOR U4431 ( .A(n3748), .B(n3749), .Z(n3745) );
  ANDN U4432 ( .B(n3750), .A(n736), .Z(n3748) );
  XNOR U4433 ( .A(a[342]), .B(n3751), .Z(n736) );
  IV U4434 ( .A(n3749), .Z(n3751) );
  XNOR U4435 ( .A(b[342]), .B(n3749), .Z(n3750) );
  XOR U4436 ( .A(n3752), .B(n3753), .Z(n3749) );
  ANDN U4437 ( .B(n3754), .A(n737), .Z(n3752) );
  XNOR U4438 ( .A(a[341]), .B(n3755), .Z(n737) );
  IV U4439 ( .A(n3753), .Z(n3755) );
  XNOR U4440 ( .A(b[341]), .B(n3753), .Z(n3754) );
  XOR U4441 ( .A(n3756), .B(n3757), .Z(n3753) );
  ANDN U4442 ( .B(n3758), .A(n738), .Z(n3756) );
  XNOR U4443 ( .A(a[340]), .B(n3759), .Z(n738) );
  IV U4444 ( .A(n3757), .Z(n3759) );
  XNOR U4445 ( .A(b[340]), .B(n3757), .Z(n3758) );
  XOR U4446 ( .A(n3760), .B(n3761), .Z(n3757) );
  ANDN U4447 ( .B(n3762), .A(n740), .Z(n3760) );
  XNOR U4448 ( .A(a[339]), .B(n3763), .Z(n740) );
  IV U4449 ( .A(n3761), .Z(n3763) );
  XNOR U4450 ( .A(b[339]), .B(n3761), .Z(n3762) );
  XOR U4451 ( .A(n3764), .B(n3765), .Z(n3761) );
  ANDN U4452 ( .B(n3766), .A(n741), .Z(n3764) );
  XNOR U4453 ( .A(a[338]), .B(n3767), .Z(n741) );
  IV U4454 ( .A(n3765), .Z(n3767) );
  XNOR U4455 ( .A(b[338]), .B(n3765), .Z(n3766) );
  XOR U4456 ( .A(n3768), .B(n3769), .Z(n3765) );
  ANDN U4457 ( .B(n3770), .A(n742), .Z(n3768) );
  XNOR U4458 ( .A(a[337]), .B(n3771), .Z(n742) );
  IV U4459 ( .A(n3769), .Z(n3771) );
  XNOR U4460 ( .A(b[337]), .B(n3769), .Z(n3770) );
  XOR U4461 ( .A(n3772), .B(n3773), .Z(n3769) );
  ANDN U4462 ( .B(n3774), .A(n743), .Z(n3772) );
  XNOR U4463 ( .A(a[336]), .B(n3775), .Z(n743) );
  IV U4464 ( .A(n3773), .Z(n3775) );
  XNOR U4465 ( .A(b[336]), .B(n3773), .Z(n3774) );
  XOR U4466 ( .A(n3776), .B(n3777), .Z(n3773) );
  ANDN U4467 ( .B(n3778), .A(n744), .Z(n3776) );
  XNOR U4468 ( .A(a[335]), .B(n3779), .Z(n744) );
  IV U4469 ( .A(n3777), .Z(n3779) );
  XNOR U4470 ( .A(b[335]), .B(n3777), .Z(n3778) );
  XOR U4471 ( .A(n3780), .B(n3781), .Z(n3777) );
  ANDN U4472 ( .B(n3782), .A(n745), .Z(n3780) );
  XNOR U4473 ( .A(a[334]), .B(n3783), .Z(n745) );
  IV U4474 ( .A(n3781), .Z(n3783) );
  XNOR U4475 ( .A(b[334]), .B(n3781), .Z(n3782) );
  XOR U4476 ( .A(n3784), .B(n3785), .Z(n3781) );
  ANDN U4477 ( .B(n3786), .A(n746), .Z(n3784) );
  XNOR U4478 ( .A(a[333]), .B(n3787), .Z(n746) );
  IV U4479 ( .A(n3785), .Z(n3787) );
  XNOR U4480 ( .A(b[333]), .B(n3785), .Z(n3786) );
  XOR U4481 ( .A(n3788), .B(n3789), .Z(n3785) );
  ANDN U4482 ( .B(n3790), .A(n747), .Z(n3788) );
  XNOR U4483 ( .A(a[332]), .B(n3791), .Z(n747) );
  IV U4484 ( .A(n3789), .Z(n3791) );
  XNOR U4485 ( .A(b[332]), .B(n3789), .Z(n3790) );
  XOR U4486 ( .A(n3792), .B(n3793), .Z(n3789) );
  ANDN U4487 ( .B(n3794), .A(n748), .Z(n3792) );
  XNOR U4488 ( .A(a[331]), .B(n3795), .Z(n748) );
  IV U4489 ( .A(n3793), .Z(n3795) );
  XNOR U4490 ( .A(b[331]), .B(n3793), .Z(n3794) );
  XOR U4491 ( .A(n3796), .B(n3797), .Z(n3793) );
  ANDN U4492 ( .B(n3798), .A(n749), .Z(n3796) );
  XNOR U4493 ( .A(a[330]), .B(n3799), .Z(n749) );
  IV U4494 ( .A(n3797), .Z(n3799) );
  XNOR U4495 ( .A(b[330]), .B(n3797), .Z(n3798) );
  XOR U4496 ( .A(n3800), .B(n3801), .Z(n3797) );
  ANDN U4497 ( .B(n3802), .A(n751), .Z(n3800) );
  XNOR U4498 ( .A(a[329]), .B(n3803), .Z(n751) );
  IV U4499 ( .A(n3801), .Z(n3803) );
  XNOR U4500 ( .A(b[329]), .B(n3801), .Z(n3802) );
  XOR U4501 ( .A(n3804), .B(n3805), .Z(n3801) );
  ANDN U4502 ( .B(n3806), .A(n752), .Z(n3804) );
  XNOR U4503 ( .A(a[328]), .B(n3807), .Z(n752) );
  IV U4504 ( .A(n3805), .Z(n3807) );
  XNOR U4505 ( .A(b[328]), .B(n3805), .Z(n3806) );
  XOR U4506 ( .A(n3808), .B(n3809), .Z(n3805) );
  ANDN U4507 ( .B(n3810), .A(n753), .Z(n3808) );
  XNOR U4508 ( .A(a[327]), .B(n3811), .Z(n753) );
  IV U4509 ( .A(n3809), .Z(n3811) );
  XNOR U4510 ( .A(b[327]), .B(n3809), .Z(n3810) );
  XOR U4511 ( .A(n3812), .B(n3813), .Z(n3809) );
  ANDN U4512 ( .B(n3814), .A(n754), .Z(n3812) );
  XNOR U4513 ( .A(a[326]), .B(n3815), .Z(n754) );
  IV U4514 ( .A(n3813), .Z(n3815) );
  XNOR U4515 ( .A(b[326]), .B(n3813), .Z(n3814) );
  XOR U4516 ( .A(n3816), .B(n3817), .Z(n3813) );
  ANDN U4517 ( .B(n3818), .A(n755), .Z(n3816) );
  XNOR U4518 ( .A(a[325]), .B(n3819), .Z(n755) );
  IV U4519 ( .A(n3817), .Z(n3819) );
  XNOR U4520 ( .A(b[325]), .B(n3817), .Z(n3818) );
  XOR U4521 ( .A(n3820), .B(n3821), .Z(n3817) );
  ANDN U4522 ( .B(n3822), .A(n756), .Z(n3820) );
  XNOR U4523 ( .A(a[324]), .B(n3823), .Z(n756) );
  IV U4524 ( .A(n3821), .Z(n3823) );
  XNOR U4525 ( .A(b[324]), .B(n3821), .Z(n3822) );
  XOR U4526 ( .A(n3824), .B(n3825), .Z(n3821) );
  ANDN U4527 ( .B(n3826), .A(n757), .Z(n3824) );
  XNOR U4528 ( .A(a[323]), .B(n3827), .Z(n757) );
  IV U4529 ( .A(n3825), .Z(n3827) );
  XNOR U4530 ( .A(b[323]), .B(n3825), .Z(n3826) );
  XOR U4531 ( .A(n3828), .B(n3829), .Z(n3825) );
  ANDN U4532 ( .B(n3830), .A(n758), .Z(n3828) );
  XNOR U4533 ( .A(a[322]), .B(n3831), .Z(n758) );
  IV U4534 ( .A(n3829), .Z(n3831) );
  XNOR U4535 ( .A(b[322]), .B(n3829), .Z(n3830) );
  XOR U4536 ( .A(n3832), .B(n3833), .Z(n3829) );
  ANDN U4537 ( .B(n3834), .A(n759), .Z(n3832) );
  XNOR U4538 ( .A(a[321]), .B(n3835), .Z(n759) );
  IV U4539 ( .A(n3833), .Z(n3835) );
  XNOR U4540 ( .A(b[321]), .B(n3833), .Z(n3834) );
  XOR U4541 ( .A(n3836), .B(n3837), .Z(n3833) );
  ANDN U4542 ( .B(n3838), .A(n760), .Z(n3836) );
  XNOR U4543 ( .A(a[320]), .B(n3839), .Z(n760) );
  IV U4544 ( .A(n3837), .Z(n3839) );
  XNOR U4545 ( .A(b[320]), .B(n3837), .Z(n3838) );
  XOR U4546 ( .A(n3840), .B(n3841), .Z(n3837) );
  ANDN U4547 ( .B(n3842), .A(n762), .Z(n3840) );
  XNOR U4548 ( .A(a[319]), .B(n3843), .Z(n762) );
  IV U4549 ( .A(n3841), .Z(n3843) );
  XNOR U4550 ( .A(b[319]), .B(n3841), .Z(n3842) );
  XOR U4551 ( .A(n3844), .B(n3845), .Z(n3841) );
  ANDN U4552 ( .B(n3846), .A(n763), .Z(n3844) );
  XNOR U4553 ( .A(a[318]), .B(n3847), .Z(n763) );
  IV U4554 ( .A(n3845), .Z(n3847) );
  XNOR U4555 ( .A(b[318]), .B(n3845), .Z(n3846) );
  XOR U4556 ( .A(n3848), .B(n3849), .Z(n3845) );
  ANDN U4557 ( .B(n3850), .A(n764), .Z(n3848) );
  XNOR U4558 ( .A(a[317]), .B(n3851), .Z(n764) );
  IV U4559 ( .A(n3849), .Z(n3851) );
  XNOR U4560 ( .A(b[317]), .B(n3849), .Z(n3850) );
  XOR U4561 ( .A(n3852), .B(n3853), .Z(n3849) );
  ANDN U4562 ( .B(n3854), .A(n765), .Z(n3852) );
  XNOR U4563 ( .A(a[316]), .B(n3855), .Z(n765) );
  IV U4564 ( .A(n3853), .Z(n3855) );
  XNOR U4565 ( .A(b[316]), .B(n3853), .Z(n3854) );
  XOR U4566 ( .A(n3856), .B(n3857), .Z(n3853) );
  ANDN U4567 ( .B(n3858), .A(n766), .Z(n3856) );
  XNOR U4568 ( .A(a[315]), .B(n3859), .Z(n766) );
  IV U4569 ( .A(n3857), .Z(n3859) );
  XNOR U4570 ( .A(b[315]), .B(n3857), .Z(n3858) );
  XOR U4571 ( .A(n3860), .B(n3861), .Z(n3857) );
  ANDN U4572 ( .B(n3862), .A(n767), .Z(n3860) );
  XNOR U4573 ( .A(a[314]), .B(n3863), .Z(n767) );
  IV U4574 ( .A(n3861), .Z(n3863) );
  XNOR U4575 ( .A(b[314]), .B(n3861), .Z(n3862) );
  XOR U4576 ( .A(n3864), .B(n3865), .Z(n3861) );
  ANDN U4577 ( .B(n3866), .A(n768), .Z(n3864) );
  XNOR U4578 ( .A(a[313]), .B(n3867), .Z(n768) );
  IV U4579 ( .A(n3865), .Z(n3867) );
  XNOR U4580 ( .A(b[313]), .B(n3865), .Z(n3866) );
  XOR U4581 ( .A(n3868), .B(n3869), .Z(n3865) );
  ANDN U4582 ( .B(n3870), .A(n769), .Z(n3868) );
  XNOR U4583 ( .A(a[312]), .B(n3871), .Z(n769) );
  IV U4584 ( .A(n3869), .Z(n3871) );
  XNOR U4585 ( .A(b[312]), .B(n3869), .Z(n3870) );
  XOR U4586 ( .A(n3872), .B(n3873), .Z(n3869) );
  ANDN U4587 ( .B(n3874), .A(n770), .Z(n3872) );
  XNOR U4588 ( .A(a[311]), .B(n3875), .Z(n770) );
  IV U4589 ( .A(n3873), .Z(n3875) );
  XNOR U4590 ( .A(b[311]), .B(n3873), .Z(n3874) );
  XOR U4591 ( .A(n3876), .B(n3877), .Z(n3873) );
  ANDN U4592 ( .B(n3878), .A(n771), .Z(n3876) );
  XNOR U4593 ( .A(a[310]), .B(n3879), .Z(n771) );
  IV U4594 ( .A(n3877), .Z(n3879) );
  XNOR U4595 ( .A(b[310]), .B(n3877), .Z(n3878) );
  XOR U4596 ( .A(n3880), .B(n3881), .Z(n3877) );
  ANDN U4597 ( .B(n3882), .A(n773), .Z(n3880) );
  XNOR U4598 ( .A(a[309]), .B(n3883), .Z(n773) );
  IV U4599 ( .A(n3881), .Z(n3883) );
  XNOR U4600 ( .A(b[309]), .B(n3881), .Z(n3882) );
  XOR U4601 ( .A(n3884), .B(n3885), .Z(n3881) );
  ANDN U4602 ( .B(n3886), .A(n774), .Z(n3884) );
  XNOR U4603 ( .A(a[308]), .B(n3887), .Z(n774) );
  IV U4604 ( .A(n3885), .Z(n3887) );
  XNOR U4605 ( .A(b[308]), .B(n3885), .Z(n3886) );
  XOR U4606 ( .A(n3888), .B(n3889), .Z(n3885) );
  ANDN U4607 ( .B(n3890), .A(n775), .Z(n3888) );
  XNOR U4608 ( .A(a[307]), .B(n3891), .Z(n775) );
  IV U4609 ( .A(n3889), .Z(n3891) );
  XNOR U4610 ( .A(b[307]), .B(n3889), .Z(n3890) );
  XOR U4611 ( .A(n3892), .B(n3893), .Z(n3889) );
  ANDN U4612 ( .B(n3894), .A(n776), .Z(n3892) );
  XNOR U4613 ( .A(a[306]), .B(n3895), .Z(n776) );
  IV U4614 ( .A(n3893), .Z(n3895) );
  XNOR U4615 ( .A(b[306]), .B(n3893), .Z(n3894) );
  XOR U4616 ( .A(n3896), .B(n3897), .Z(n3893) );
  ANDN U4617 ( .B(n3898), .A(n777), .Z(n3896) );
  XNOR U4618 ( .A(a[305]), .B(n3899), .Z(n777) );
  IV U4619 ( .A(n3897), .Z(n3899) );
  XNOR U4620 ( .A(b[305]), .B(n3897), .Z(n3898) );
  XOR U4621 ( .A(n3900), .B(n3901), .Z(n3897) );
  ANDN U4622 ( .B(n3902), .A(n778), .Z(n3900) );
  XNOR U4623 ( .A(a[304]), .B(n3903), .Z(n778) );
  IV U4624 ( .A(n3901), .Z(n3903) );
  XNOR U4625 ( .A(b[304]), .B(n3901), .Z(n3902) );
  XOR U4626 ( .A(n3904), .B(n3905), .Z(n3901) );
  ANDN U4627 ( .B(n3906), .A(n779), .Z(n3904) );
  XNOR U4628 ( .A(a[303]), .B(n3907), .Z(n779) );
  IV U4629 ( .A(n3905), .Z(n3907) );
  XNOR U4630 ( .A(b[303]), .B(n3905), .Z(n3906) );
  XOR U4631 ( .A(n3908), .B(n3909), .Z(n3905) );
  ANDN U4632 ( .B(n3910), .A(n780), .Z(n3908) );
  XNOR U4633 ( .A(a[302]), .B(n3911), .Z(n780) );
  IV U4634 ( .A(n3909), .Z(n3911) );
  XNOR U4635 ( .A(b[302]), .B(n3909), .Z(n3910) );
  XOR U4636 ( .A(n3912), .B(n3913), .Z(n3909) );
  ANDN U4637 ( .B(n3914), .A(n781), .Z(n3912) );
  XNOR U4638 ( .A(a[301]), .B(n3915), .Z(n781) );
  IV U4639 ( .A(n3913), .Z(n3915) );
  XNOR U4640 ( .A(b[301]), .B(n3913), .Z(n3914) );
  XOR U4641 ( .A(n3916), .B(n3917), .Z(n3913) );
  ANDN U4642 ( .B(n3918), .A(n782), .Z(n3916) );
  XNOR U4643 ( .A(a[300]), .B(n3919), .Z(n782) );
  IV U4644 ( .A(n3917), .Z(n3919) );
  XNOR U4645 ( .A(b[300]), .B(n3917), .Z(n3918) );
  XOR U4646 ( .A(n3920), .B(n3921), .Z(n3917) );
  ANDN U4647 ( .B(n3922), .A(n785), .Z(n3920) );
  XNOR U4648 ( .A(a[299]), .B(n3923), .Z(n785) );
  IV U4649 ( .A(n3921), .Z(n3923) );
  XNOR U4650 ( .A(b[299]), .B(n3921), .Z(n3922) );
  XOR U4651 ( .A(n3924), .B(n3925), .Z(n3921) );
  ANDN U4652 ( .B(n3926), .A(n786), .Z(n3924) );
  XNOR U4653 ( .A(a[298]), .B(n3927), .Z(n786) );
  IV U4654 ( .A(n3925), .Z(n3927) );
  XNOR U4655 ( .A(b[298]), .B(n3925), .Z(n3926) );
  XOR U4656 ( .A(n3928), .B(n3929), .Z(n3925) );
  ANDN U4657 ( .B(n3930), .A(n787), .Z(n3928) );
  XNOR U4658 ( .A(a[297]), .B(n3931), .Z(n787) );
  IV U4659 ( .A(n3929), .Z(n3931) );
  XNOR U4660 ( .A(b[297]), .B(n3929), .Z(n3930) );
  XOR U4661 ( .A(n3932), .B(n3933), .Z(n3929) );
  ANDN U4662 ( .B(n3934), .A(n788), .Z(n3932) );
  XNOR U4663 ( .A(a[296]), .B(n3935), .Z(n788) );
  IV U4664 ( .A(n3933), .Z(n3935) );
  XNOR U4665 ( .A(b[296]), .B(n3933), .Z(n3934) );
  XOR U4666 ( .A(n3936), .B(n3937), .Z(n3933) );
  ANDN U4667 ( .B(n3938), .A(n789), .Z(n3936) );
  XNOR U4668 ( .A(a[295]), .B(n3939), .Z(n789) );
  IV U4669 ( .A(n3937), .Z(n3939) );
  XNOR U4670 ( .A(b[295]), .B(n3937), .Z(n3938) );
  XOR U4671 ( .A(n3940), .B(n3941), .Z(n3937) );
  ANDN U4672 ( .B(n3942), .A(n790), .Z(n3940) );
  XNOR U4673 ( .A(a[294]), .B(n3943), .Z(n790) );
  IV U4674 ( .A(n3941), .Z(n3943) );
  XNOR U4675 ( .A(b[294]), .B(n3941), .Z(n3942) );
  XOR U4676 ( .A(n3944), .B(n3945), .Z(n3941) );
  ANDN U4677 ( .B(n3946), .A(n791), .Z(n3944) );
  XNOR U4678 ( .A(a[293]), .B(n3947), .Z(n791) );
  IV U4679 ( .A(n3945), .Z(n3947) );
  XNOR U4680 ( .A(b[293]), .B(n3945), .Z(n3946) );
  XOR U4681 ( .A(n3948), .B(n3949), .Z(n3945) );
  ANDN U4682 ( .B(n3950), .A(n792), .Z(n3948) );
  XNOR U4683 ( .A(a[292]), .B(n3951), .Z(n792) );
  IV U4684 ( .A(n3949), .Z(n3951) );
  XNOR U4685 ( .A(b[292]), .B(n3949), .Z(n3950) );
  XOR U4686 ( .A(n3952), .B(n3953), .Z(n3949) );
  ANDN U4687 ( .B(n3954), .A(n793), .Z(n3952) );
  XNOR U4688 ( .A(a[291]), .B(n3955), .Z(n793) );
  IV U4689 ( .A(n3953), .Z(n3955) );
  XNOR U4690 ( .A(b[291]), .B(n3953), .Z(n3954) );
  XOR U4691 ( .A(n3956), .B(n3957), .Z(n3953) );
  ANDN U4692 ( .B(n3958), .A(n794), .Z(n3956) );
  XNOR U4693 ( .A(a[290]), .B(n3959), .Z(n794) );
  IV U4694 ( .A(n3957), .Z(n3959) );
  XNOR U4695 ( .A(b[290]), .B(n3957), .Z(n3958) );
  XOR U4696 ( .A(n3960), .B(n3961), .Z(n3957) );
  ANDN U4697 ( .B(n3962), .A(n796), .Z(n3960) );
  XNOR U4698 ( .A(a[289]), .B(n3963), .Z(n796) );
  IV U4699 ( .A(n3961), .Z(n3963) );
  XNOR U4700 ( .A(b[289]), .B(n3961), .Z(n3962) );
  XOR U4701 ( .A(n3964), .B(n3965), .Z(n3961) );
  ANDN U4702 ( .B(n3966), .A(n797), .Z(n3964) );
  XNOR U4703 ( .A(a[288]), .B(n3967), .Z(n797) );
  IV U4704 ( .A(n3965), .Z(n3967) );
  XNOR U4705 ( .A(b[288]), .B(n3965), .Z(n3966) );
  XOR U4706 ( .A(n3968), .B(n3969), .Z(n3965) );
  ANDN U4707 ( .B(n3970), .A(n798), .Z(n3968) );
  XNOR U4708 ( .A(a[287]), .B(n3971), .Z(n798) );
  IV U4709 ( .A(n3969), .Z(n3971) );
  XNOR U4710 ( .A(b[287]), .B(n3969), .Z(n3970) );
  XOR U4711 ( .A(n3972), .B(n3973), .Z(n3969) );
  ANDN U4712 ( .B(n3974), .A(n799), .Z(n3972) );
  XNOR U4713 ( .A(a[286]), .B(n3975), .Z(n799) );
  IV U4714 ( .A(n3973), .Z(n3975) );
  XNOR U4715 ( .A(b[286]), .B(n3973), .Z(n3974) );
  XOR U4716 ( .A(n3976), .B(n3977), .Z(n3973) );
  ANDN U4717 ( .B(n3978), .A(n800), .Z(n3976) );
  XNOR U4718 ( .A(a[285]), .B(n3979), .Z(n800) );
  IV U4719 ( .A(n3977), .Z(n3979) );
  XNOR U4720 ( .A(b[285]), .B(n3977), .Z(n3978) );
  XOR U4721 ( .A(n3980), .B(n3981), .Z(n3977) );
  ANDN U4722 ( .B(n3982), .A(n801), .Z(n3980) );
  XNOR U4723 ( .A(a[284]), .B(n3983), .Z(n801) );
  IV U4724 ( .A(n3981), .Z(n3983) );
  XNOR U4725 ( .A(b[284]), .B(n3981), .Z(n3982) );
  XOR U4726 ( .A(n3984), .B(n3985), .Z(n3981) );
  ANDN U4727 ( .B(n3986), .A(n802), .Z(n3984) );
  XNOR U4728 ( .A(a[283]), .B(n3987), .Z(n802) );
  IV U4729 ( .A(n3985), .Z(n3987) );
  XNOR U4730 ( .A(b[283]), .B(n3985), .Z(n3986) );
  XOR U4731 ( .A(n3988), .B(n3989), .Z(n3985) );
  ANDN U4732 ( .B(n3990), .A(n803), .Z(n3988) );
  XNOR U4733 ( .A(a[282]), .B(n3991), .Z(n803) );
  IV U4734 ( .A(n3989), .Z(n3991) );
  XNOR U4735 ( .A(b[282]), .B(n3989), .Z(n3990) );
  XOR U4736 ( .A(n3992), .B(n3993), .Z(n3989) );
  ANDN U4737 ( .B(n3994), .A(n804), .Z(n3992) );
  XNOR U4738 ( .A(a[281]), .B(n3995), .Z(n804) );
  IV U4739 ( .A(n3993), .Z(n3995) );
  XNOR U4740 ( .A(b[281]), .B(n3993), .Z(n3994) );
  XOR U4741 ( .A(n3996), .B(n3997), .Z(n3993) );
  ANDN U4742 ( .B(n3998), .A(n805), .Z(n3996) );
  XNOR U4743 ( .A(a[280]), .B(n3999), .Z(n805) );
  IV U4744 ( .A(n3997), .Z(n3999) );
  XNOR U4745 ( .A(b[280]), .B(n3997), .Z(n3998) );
  XOR U4746 ( .A(n4000), .B(n4001), .Z(n3997) );
  ANDN U4747 ( .B(n4002), .A(n807), .Z(n4000) );
  XNOR U4748 ( .A(a[279]), .B(n4003), .Z(n807) );
  IV U4749 ( .A(n4001), .Z(n4003) );
  XNOR U4750 ( .A(b[279]), .B(n4001), .Z(n4002) );
  XOR U4751 ( .A(n4004), .B(n4005), .Z(n4001) );
  ANDN U4752 ( .B(n4006), .A(n808), .Z(n4004) );
  XNOR U4753 ( .A(a[278]), .B(n4007), .Z(n808) );
  IV U4754 ( .A(n4005), .Z(n4007) );
  XNOR U4755 ( .A(b[278]), .B(n4005), .Z(n4006) );
  XOR U4756 ( .A(n4008), .B(n4009), .Z(n4005) );
  ANDN U4757 ( .B(n4010), .A(n809), .Z(n4008) );
  XNOR U4758 ( .A(a[277]), .B(n4011), .Z(n809) );
  IV U4759 ( .A(n4009), .Z(n4011) );
  XNOR U4760 ( .A(b[277]), .B(n4009), .Z(n4010) );
  XOR U4761 ( .A(n4012), .B(n4013), .Z(n4009) );
  ANDN U4762 ( .B(n4014), .A(n810), .Z(n4012) );
  XNOR U4763 ( .A(a[276]), .B(n4015), .Z(n810) );
  IV U4764 ( .A(n4013), .Z(n4015) );
  XNOR U4765 ( .A(b[276]), .B(n4013), .Z(n4014) );
  XOR U4766 ( .A(n4016), .B(n4017), .Z(n4013) );
  ANDN U4767 ( .B(n4018), .A(n811), .Z(n4016) );
  XNOR U4768 ( .A(a[275]), .B(n4019), .Z(n811) );
  IV U4769 ( .A(n4017), .Z(n4019) );
  XNOR U4770 ( .A(b[275]), .B(n4017), .Z(n4018) );
  XOR U4771 ( .A(n4020), .B(n4021), .Z(n4017) );
  ANDN U4772 ( .B(n4022), .A(n812), .Z(n4020) );
  XNOR U4773 ( .A(a[274]), .B(n4023), .Z(n812) );
  IV U4774 ( .A(n4021), .Z(n4023) );
  XNOR U4775 ( .A(b[274]), .B(n4021), .Z(n4022) );
  XOR U4776 ( .A(n4024), .B(n4025), .Z(n4021) );
  ANDN U4777 ( .B(n4026), .A(n813), .Z(n4024) );
  XNOR U4778 ( .A(a[273]), .B(n4027), .Z(n813) );
  IV U4779 ( .A(n4025), .Z(n4027) );
  XNOR U4780 ( .A(b[273]), .B(n4025), .Z(n4026) );
  XOR U4781 ( .A(n4028), .B(n4029), .Z(n4025) );
  ANDN U4782 ( .B(n4030), .A(n814), .Z(n4028) );
  XNOR U4783 ( .A(a[272]), .B(n4031), .Z(n814) );
  IV U4784 ( .A(n4029), .Z(n4031) );
  XNOR U4785 ( .A(b[272]), .B(n4029), .Z(n4030) );
  XOR U4786 ( .A(n4032), .B(n4033), .Z(n4029) );
  ANDN U4787 ( .B(n4034), .A(n815), .Z(n4032) );
  XNOR U4788 ( .A(a[271]), .B(n4035), .Z(n815) );
  IV U4789 ( .A(n4033), .Z(n4035) );
  XNOR U4790 ( .A(b[271]), .B(n4033), .Z(n4034) );
  XOR U4791 ( .A(n4036), .B(n4037), .Z(n4033) );
  ANDN U4792 ( .B(n4038), .A(n816), .Z(n4036) );
  XNOR U4793 ( .A(a[270]), .B(n4039), .Z(n816) );
  IV U4794 ( .A(n4037), .Z(n4039) );
  XNOR U4795 ( .A(b[270]), .B(n4037), .Z(n4038) );
  XOR U4796 ( .A(n4040), .B(n4041), .Z(n4037) );
  ANDN U4797 ( .B(n4042), .A(n818), .Z(n4040) );
  XNOR U4798 ( .A(a[269]), .B(n4043), .Z(n818) );
  IV U4799 ( .A(n4041), .Z(n4043) );
  XNOR U4800 ( .A(b[269]), .B(n4041), .Z(n4042) );
  XOR U4801 ( .A(n4044), .B(n4045), .Z(n4041) );
  ANDN U4802 ( .B(n4046), .A(n819), .Z(n4044) );
  XNOR U4803 ( .A(a[268]), .B(n4047), .Z(n819) );
  IV U4804 ( .A(n4045), .Z(n4047) );
  XNOR U4805 ( .A(b[268]), .B(n4045), .Z(n4046) );
  XOR U4806 ( .A(n4048), .B(n4049), .Z(n4045) );
  ANDN U4807 ( .B(n4050), .A(n820), .Z(n4048) );
  XNOR U4808 ( .A(a[267]), .B(n4051), .Z(n820) );
  IV U4809 ( .A(n4049), .Z(n4051) );
  XNOR U4810 ( .A(b[267]), .B(n4049), .Z(n4050) );
  XOR U4811 ( .A(n4052), .B(n4053), .Z(n4049) );
  ANDN U4812 ( .B(n4054), .A(n821), .Z(n4052) );
  XNOR U4813 ( .A(a[266]), .B(n4055), .Z(n821) );
  IV U4814 ( .A(n4053), .Z(n4055) );
  XNOR U4815 ( .A(b[266]), .B(n4053), .Z(n4054) );
  XOR U4816 ( .A(n4056), .B(n4057), .Z(n4053) );
  ANDN U4817 ( .B(n4058), .A(n822), .Z(n4056) );
  XNOR U4818 ( .A(a[265]), .B(n4059), .Z(n822) );
  IV U4819 ( .A(n4057), .Z(n4059) );
  XNOR U4820 ( .A(b[265]), .B(n4057), .Z(n4058) );
  XOR U4821 ( .A(n4060), .B(n4061), .Z(n4057) );
  ANDN U4822 ( .B(n4062), .A(n823), .Z(n4060) );
  XNOR U4823 ( .A(a[264]), .B(n4063), .Z(n823) );
  IV U4824 ( .A(n4061), .Z(n4063) );
  XNOR U4825 ( .A(b[264]), .B(n4061), .Z(n4062) );
  XOR U4826 ( .A(n4064), .B(n4065), .Z(n4061) );
  ANDN U4827 ( .B(n4066), .A(n824), .Z(n4064) );
  XNOR U4828 ( .A(a[263]), .B(n4067), .Z(n824) );
  IV U4829 ( .A(n4065), .Z(n4067) );
  XNOR U4830 ( .A(b[263]), .B(n4065), .Z(n4066) );
  XOR U4831 ( .A(n4068), .B(n4069), .Z(n4065) );
  ANDN U4832 ( .B(n4070), .A(n825), .Z(n4068) );
  XNOR U4833 ( .A(a[262]), .B(n4071), .Z(n825) );
  IV U4834 ( .A(n4069), .Z(n4071) );
  XNOR U4835 ( .A(b[262]), .B(n4069), .Z(n4070) );
  XOR U4836 ( .A(n4072), .B(n4073), .Z(n4069) );
  ANDN U4837 ( .B(n4074), .A(n826), .Z(n4072) );
  XNOR U4838 ( .A(a[261]), .B(n4075), .Z(n826) );
  IV U4839 ( .A(n4073), .Z(n4075) );
  XNOR U4840 ( .A(b[261]), .B(n4073), .Z(n4074) );
  XOR U4841 ( .A(n4076), .B(n4077), .Z(n4073) );
  ANDN U4842 ( .B(n4078), .A(n827), .Z(n4076) );
  XNOR U4843 ( .A(a[260]), .B(n4079), .Z(n827) );
  IV U4844 ( .A(n4077), .Z(n4079) );
  XNOR U4845 ( .A(b[260]), .B(n4077), .Z(n4078) );
  XOR U4846 ( .A(n4080), .B(n4081), .Z(n4077) );
  ANDN U4847 ( .B(n4082), .A(n829), .Z(n4080) );
  XNOR U4848 ( .A(a[259]), .B(n4083), .Z(n829) );
  IV U4849 ( .A(n4081), .Z(n4083) );
  XNOR U4850 ( .A(b[259]), .B(n4081), .Z(n4082) );
  XOR U4851 ( .A(n4084), .B(n4085), .Z(n4081) );
  ANDN U4852 ( .B(n4086), .A(n830), .Z(n4084) );
  XNOR U4853 ( .A(a[258]), .B(n4087), .Z(n830) );
  IV U4854 ( .A(n4085), .Z(n4087) );
  XNOR U4855 ( .A(b[258]), .B(n4085), .Z(n4086) );
  XOR U4856 ( .A(n4088), .B(n4089), .Z(n4085) );
  ANDN U4857 ( .B(n4090), .A(n831), .Z(n4088) );
  XNOR U4858 ( .A(a[257]), .B(n4091), .Z(n831) );
  IV U4859 ( .A(n4089), .Z(n4091) );
  XNOR U4860 ( .A(b[257]), .B(n4089), .Z(n4090) );
  XOR U4861 ( .A(n4092), .B(n4093), .Z(n4089) );
  ANDN U4862 ( .B(n4094), .A(n832), .Z(n4092) );
  XNOR U4863 ( .A(a[256]), .B(n4095), .Z(n832) );
  IV U4864 ( .A(n4093), .Z(n4095) );
  XNOR U4865 ( .A(b[256]), .B(n4093), .Z(n4094) );
  XOR U4866 ( .A(n4096), .B(n4097), .Z(n4093) );
  ANDN U4867 ( .B(n4098), .A(n833), .Z(n4096) );
  XNOR U4868 ( .A(a[255]), .B(n4099), .Z(n833) );
  IV U4869 ( .A(n4097), .Z(n4099) );
  XNOR U4870 ( .A(b[255]), .B(n4097), .Z(n4098) );
  XOR U4871 ( .A(n4100), .B(n4101), .Z(n4097) );
  ANDN U4872 ( .B(n4102), .A(n834), .Z(n4100) );
  XNOR U4873 ( .A(a[254]), .B(n4103), .Z(n834) );
  IV U4874 ( .A(n4101), .Z(n4103) );
  XNOR U4875 ( .A(b[254]), .B(n4101), .Z(n4102) );
  XOR U4876 ( .A(n4104), .B(n4105), .Z(n4101) );
  ANDN U4877 ( .B(n4106), .A(n835), .Z(n4104) );
  XNOR U4878 ( .A(a[253]), .B(n4107), .Z(n835) );
  IV U4879 ( .A(n4105), .Z(n4107) );
  XNOR U4880 ( .A(b[253]), .B(n4105), .Z(n4106) );
  XOR U4881 ( .A(n4108), .B(n4109), .Z(n4105) );
  ANDN U4882 ( .B(n4110), .A(n836), .Z(n4108) );
  XNOR U4883 ( .A(a[252]), .B(n4111), .Z(n836) );
  IV U4884 ( .A(n4109), .Z(n4111) );
  XNOR U4885 ( .A(b[252]), .B(n4109), .Z(n4110) );
  XOR U4886 ( .A(n4112), .B(n4113), .Z(n4109) );
  ANDN U4887 ( .B(n4114), .A(n837), .Z(n4112) );
  XNOR U4888 ( .A(a[251]), .B(n4115), .Z(n837) );
  IV U4889 ( .A(n4113), .Z(n4115) );
  XNOR U4890 ( .A(b[251]), .B(n4113), .Z(n4114) );
  XOR U4891 ( .A(n4116), .B(n4117), .Z(n4113) );
  ANDN U4892 ( .B(n4118), .A(n838), .Z(n4116) );
  XNOR U4893 ( .A(a[250]), .B(n4119), .Z(n838) );
  IV U4894 ( .A(n4117), .Z(n4119) );
  XNOR U4895 ( .A(b[250]), .B(n4117), .Z(n4118) );
  XOR U4896 ( .A(n4120), .B(n4121), .Z(n4117) );
  ANDN U4897 ( .B(n4122), .A(n840), .Z(n4120) );
  XNOR U4898 ( .A(a[249]), .B(n4123), .Z(n840) );
  IV U4899 ( .A(n4121), .Z(n4123) );
  XNOR U4900 ( .A(b[249]), .B(n4121), .Z(n4122) );
  XOR U4901 ( .A(n4124), .B(n4125), .Z(n4121) );
  ANDN U4902 ( .B(n4126), .A(n841), .Z(n4124) );
  XNOR U4903 ( .A(a[248]), .B(n4127), .Z(n841) );
  IV U4904 ( .A(n4125), .Z(n4127) );
  XNOR U4905 ( .A(b[248]), .B(n4125), .Z(n4126) );
  XOR U4906 ( .A(n4128), .B(n4129), .Z(n4125) );
  ANDN U4907 ( .B(n4130), .A(n842), .Z(n4128) );
  XNOR U4908 ( .A(a[247]), .B(n4131), .Z(n842) );
  IV U4909 ( .A(n4129), .Z(n4131) );
  XNOR U4910 ( .A(b[247]), .B(n4129), .Z(n4130) );
  XOR U4911 ( .A(n4132), .B(n4133), .Z(n4129) );
  ANDN U4912 ( .B(n4134), .A(n843), .Z(n4132) );
  XNOR U4913 ( .A(a[246]), .B(n4135), .Z(n843) );
  IV U4914 ( .A(n4133), .Z(n4135) );
  XNOR U4915 ( .A(b[246]), .B(n4133), .Z(n4134) );
  XOR U4916 ( .A(n4136), .B(n4137), .Z(n4133) );
  ANDN U4917 ( .B(n4138), .A(n844), .Z(n4136) );
  XNOR U4918 ( .A(a[245]), .B(n4139), .Z(n844) );
  IV U4919 ( .A(n4137), .Z(n4139) );
  XNOR U4920 ( .A(b[245]), .B(n4137), .Z(n4138) );
  XOR U4921 ( .A(n4140), .B(n4141), .Z(n4137) );
  ANDN U4922 ( .B(n4142), .A(n845), .Z(n4140) );
  XNOR U4923 ( .A(a[244]), .B(n4143), .Z(n845) );
  IV U4924 ( .A(n4141), .Z(n4143) );
  XNOR U4925 ( .A(b[244]), .B(n4141), .Z(n4142) );
  XOR U4926 ( .A(n4144), .B(n4145), .Z(n4141) );
  ANDN U4927 ( .B(n4146), .A(n846), .Z(n4144) );
  XNOR U4928 ( .A(a[243]), .B(n4147), .Z(n846) );
  IV U4929 ( .A(n4145), .Z(n4147) );
  XNOR U4930 ( .A(b[243]), .B(n4145), .Z(n4146) );
  XOR U4931 ( .A(n4148), .B(n4149), .Z(n4145) );
  ANDN U4932 ( .B(n4150), .A(n847), .Z(n4148) );
  XNOR U4933 ( .A(a[242]), .B(n4151), .Z(n847) );
  IV U4934 ( .A(n4149), .Z(n4151) );
  XNOR U4935 ( .A(b[242]), .B(n4149), .Z(n4150) );
  XOR U4936 ( .A(n4152), .B(n4153), .Z(n4149) );
  ANDN U4937 ( .B(n4154), .A(n848), .Z(n4152) );
  XNOR U4938 ( .A(a[241]), .B(n4155), .Z(n848) );
  IV U4939 ( .A(n4153), .Z(n4155) );
  XNOR U4940 ( .A(b[241]), .B(n4153), .Z(n4154) );
  XOR U4941 ( .A(n4156), .B(n4157), .Z(n4153) );
  ANDN U4942 ( .B(n4158), .A(n849), .Z(n4156) );
  XNOR U4943 ( .A(a[240]), .B(n4159), .Z(n849) );
  IV U4944 ( .A(n4157), .Z(n4159) );
  XNOR U4945 ( .A(b[240]), .B(n4157), .Z(n4158) );
  XOR U4946 ( .A(n4160), .B(n4161), .Z(n4157) );
  ANDN U4947 ( .B(n4162), .A(n851), .Z(n4160) );
  XNOR U4948 ( .A(a[239]), .B(n4163), .Z(n851) );
  IV U4949 ( .A(n4161), .Z(n4163) );
  XNOR U4950 ( .A(b[239]), .B(n4161), .Z(n4162) );
  XOR U4951 ( .A(n4164), .B(n4165), .Z(n4161) );
  ANDN U4952 ( .B(n4166), .A(n852), .Z(n4164) );
  XNOR U4953 ( .A(a[238]), .B(n4167), .Z(n852) );
  IV U4954 ( .A(n4165), .Z(n4167) );
  XNOR U4955 ( .A(b[238]), .B(n4165), .Z(n4166) );
  XOR U4956 ( .A(n4168), .B(n4169), .Z(n4165) );
  ANDN U4957 ( .B(n4170), .A(n853), .Z(n4168) );
  XNOR U4958 ( .A(a[237]), .B(n4171), .Z(n853) );
  IV U4959 ( .A(n4169), .Z(n4171) );
  XNOR U4960 ( .A(b[237]), .B(n4169), .Z(n4170) );
  XOR U4961 ( .A(n4172), .B(n4173), .Z(n4169) );
  ANDN U4962 ( .B(n4174), .A(n854), .Z(n4172) );
  XNOR U4963 ( .A(a[236]), .B(n4175), .Z(n854) );
  IV U4964 ( .A(n4173), .Z(n4175) );
  XNOR U4965 ( .A(b[236]), .B(n4173), .Z(n4174) );
  XOR U4966 ( .A(n4176), .B(n4177), .Z(n4173) );
  ANDN U4967 ( .B(n4178), .A(n855), .Z(n4176) );
  XNOR U4968 ( .A(a[235]), .B(n4179), .Z(n855) );
  IV U4969 ( .A(n4177), .Z(n4179) );
  XNOR U4970 ( .A(b[235]), .B(n4177), .Z(n4178) );
  XOR U4971 ( .A(n4180), .B(n4181), .Z(n4177) );
  ANDN U4972 ( .B(n4182), .A(n856), .Z(n4180) );
  XNOR U4973 ( .A(a[234]), .B(n4183), .Z(n856) );
  IV U4974 ( .A(n4181), .Z(n4183) );
  XNOR U4975 ( .A(b[234]), .B(n4181), .Z(n4182) );
  XOR U4976 ( .A(n4184), .B(n4185), .Z(n4181) );
  ANDN U4977 ( .B(n4186), .A(n857), .Z(n4184) );
  XNOR U4978 ( .A(a[233]), .B(n4187), .Z(n857) );
  IV U4979 ( .A(n4185), .Z(n4187) );
  XNOR U4980 ( .A(b[233]), .B(n4185), .Z(n4186) );
  XOR U4981 ( .A(n4188), .B(n4189), .Z(n4185) );
  ANDN U4982 ( .B(n4190), .A(n858), .Z(n4188) );
  XNOR U4983 ( .A(a[232]), .B(n4191), .Z(n858) );
  IV U4984 ( .A(n4189), .Z(n4191) );
  XNOR U4985 ( .A(b[232]), .B(n4189), .Z(n4190) );
  XOR U4986 ( .A(n4192), .B(n4193), .Z(n4189) );
  ANDN U4987 ( .B(n4194), .A(n859), .Z(n4192) );
  XNOR U4988 ( .A(a[231]), .B(n4195), .Z(n859) );
  IV U4989 ( .A(n4193), .Z(n4195) );
  XNOR U4990 ( .A(b[231]), .B(n4193), .Z(n4194) );
  XOR U4991 ( .A(n4196), .B(n4197), .Z(n4193) );
  ANDN U4992 ( .B(n4198), .A(n860), .Z(n4196) );
  XNOR U4993 ( .A(a[230]), .B(n4199), .Z(n860) );
  IV U4994 ( .A(n4197), .Z(n4199) );
  XNOR U4995 ( .A(b[230]), .B(n4197), .Z(n4198) );
  XOR U4996 ( .A(n4200), .B(n4201), .Z(n4197) );
  ANDN U4997 ( .B(n4202), .A(n862), .Z(n4200) );
  XNOR U4998 ( .A(a[229]), .B(n4203), .Z(n862) );
  IV U4999 ( .A(n4201), .Z(n4203) );
  XNOR U5000 ( .A(b[229]), .B(n4201), .Z(n4202) );
  XOR U5001 ( .A(n4204), .B(n4205), .Z(n4201) );
  ANDN U5002 ( .B(n4206), .A(n863), .Z(n4204) );
  XNOR U5003 ( .A(a[228]), .B(n4207), .Z(n863) );
  IV U5004 ( .A(n4205), .Z(n4207) );
  XNOR U5005 ( .A(b[228]), .B(n4205), .Z(n4206) );
  XOR U5006 ( .A(n4208), .B(n4209), .Z(n4205) );
  ANDN U5007 ( .B(n4210), .A(n864), .Z(n4208) );
  XNOR U5008 ( .A(a[227]), .B(n4211), .Z(n864) );
  IV U5009 ( .A(n4209), .Z(n4211) );
  XNOR U5010 ( .A(b[227]), .B(n4209), .Z(n4210) );
  XOR U5011 ( .A(n4212), .B(n4213), .Z(n4209) );
  ANDN U5012 ( .B(n4214), .A(n865), .Z(n4212) );
  XNOR U5013 ( .A(a[226]), .B(n4215), .Z(n865) );
  IV U5014 ( .A(n4213), .Z(n4215) );
  XNOR U5015 ( .A(b[226]), .B(n4213), .Z(n4214) );
  XOR U5016 ( .A(n4216), .B(n4217), .Z(n4213) );
  ANDN U5017 ( .B(n4218), .A(n866), .Z(n4216) );
  XNOR U5018 ( .A(a[225]), .B(n4219), .Z(n866) );
  IV U5019 ( .A(n4217), .Z(n4219) );
  XNOR U5020 ( .A(b[225]), .B(n4217), .Z(n4218) );
  XOR U5021 ( .A(n4220), .B(n4221), .Z(n4217) );
  ANDN U5022 ( .B(n4222), .A(n867), .Z(n4220) );
  XNOR U5023 ( .A(a[224]), .B(n4223), .Z(n867) );
  IV U5024 ( .A(n4221), .Z(n4223) );
  XNOR U5025 ( .A(b[224]), .B(n4221), .Z(n4222) );
  XOR U5026 ( .A(n4224), .B(n4225), .Z(n4221) );
  ANDN U5027 ( .B(n4226), .A(n868), .Z(n4224) );
  XNOR U5028 ( .A(a[223]), .B(n4227), .Z(n868) );
  IV U5029 ( .A(n4225), .Z(n4227) );
  XNOR U5030 ( .A(b[223]), .B(n4225), .Z(n4226) );
  XOR U5031 ( .A(n4228), .B(n4229), .Z(n4225) );
  ANDN U5032 ( .B(n4230), .A(n869), .Z(n4228) );
  XNOR U5033 ( .A(a[222]), .B(n4231), .Z(n869) );
  IV U5034 ( .A(n4229), .Z(n4231) );
  XNOR U5035 ( .A(b[222]), .B(n4229), .Z(n4230) );
  XOR U5036 ( .A(n4232), .B(n4233), .Z(n4229) );
  ANDN U5037 ( .B(n4234), .A(n870), .Z(n4232) );
  XNOR U5038 ( .A(a[221]), .B(n4235), .Z(n870) );
  IV U5039 ( .A(n4233), .Z(n4235) );
  XNOR U5040 ( .A(b[221]), .B(n4233), .Z(n4234) );
  XOR U5041 ( .A(n4236), .B(n4237), .Z(n4233) );
  ANDN U5042 ( .B(n4238), .A(n871), .Z(n4236) );
  XNOR U5043 ( .A(a[220]), .B(n4239), .Z(n871) );
  IV U5044 ( .A(n4237), .Z(n4239) );
  XNOR U5045 ( .A(b[220]), .B(n4237), .Z(n4238) );
  XOR U5046 ( .A(n4240), .B(n4241), .Z(n4237) );
  ANDN U5047 ( .B(n4242), .A(n873), .Z(n4240) );
  XNOR U5048 ( .A(a[219]), .B(n4243), .Z(n873) );
  IV U5049 ( .A(n4241), .Z(n4243) );
  XNOR U5050 ( .A(b[219]), .B(n4241), .Z(n4242) );
  XOR U5051 ( .A(n4244), .B(n4245), .Z(n4241) );
  ANDN U5052 ( .B(n4246), .A(n874), .Z(n4244) );
  XNOR U5053 ( .A(a[218]), .B(n4247), .Z(n874) );
  IV U5054 ( .A(n4245), .Z(n4247) );
  XNOR U5055 ( .A(b[218]), .B(n4245), .Z(n4246) );
  XOR U5056 ( .A(n4248), .B(n4249), .Z(n4245) );
  ANDN U5057 ( .B(n4250), .A(n875), .Z(n4248) );
  XNOR U5058 ( .A(a[217]), .B(n4251), .Z(n875) );
  IV U5059 ( .A(n4249), .Z(n4251) );
  XNOR U5060 ( .A(b[217]), .B(n4249), .Z(n4250) );
  XOR U5061 ( .A(n4252), .B(n4253), .Z(n4249) );
  ANDN U5062 ( .B(n4254), .A(n876), .Z(n4252) );
  XNOR U5063 ( .A(a[216]), .B(n4255), .Z(n876) );
  IV U5064 ( .A(n4253), .Z(n4255) );
  XNOR U5065 ( .A(b[216]), .B(n4253), .Z(n4254) );
  XOR U5066 ( .A(n4256), .B(n4257), .Z(n4253) );
  ANDN U5067 ( .B(n4258), .A(n877), .Z(n4256) );
  XNOR U5068 ( .A(a[215]), .B(n4259), .Z(n877) );
  IV U5069 ( .A(n4257), .Z(n4259) );
  XNOR U5070 ( .A(b[215]), .B(n4257), .Z(n4258) );
  XOR U5071 ( .A(n4260), .B(n4261), .Z(n4257) );
  ANDN U5072 ( .B(n4262), .A(n878), .Z(n4260) );
  XNOR U5073 ( .A(a[214]), .B(n4263), .Z(n878) );
  IV U5074 ( .A(n4261), .Z(n4263) );
  XNOR U5075 ( .A(b[214]), .B(n4261), .Z(n4262) );
  XOR U5076 ( .A(n4264), .B(n4265), .Z(n4261) );
  ANDN U5077 ( .B(n4266), .A(n879), .Z(n4264) );
  XNOR U5078 ( .A(a[213]), .B(n4267), .Z(n879) );
  IV U5079 ( .A(n4265), .Z(n4267) );
  XNOR U5080 ( .A(b[213]), .B(n4265), .Z(n4266) );
  XOR U5081 ( .A(n4268), .B(n4269), .Z(n4265) );
  ANDN U5082 ( .B(n4270), .A(n880), .Z(n4268) );
  XNOR U5083 ( .A(a[212]), .B(n4271), .Z(n880) );
  IV U5084 ( .A(n4269), .Z(n4271) );
  XNOR U5085 ( .A(b[212]), .B(n4269), .Z(n4270) );
  XOR U5086 ( .A(n4272), .B(n4273), .Z(n4269) );
  ANDN U5087 ( .B(n4274), .A(n881), .Z(n4272) );
  XNOR U5088 ( .A(a[211]), .B(n4275), .Z(n881) );
  IV U5089 ( .A(n4273), .Z(n4275) );
  XNOR U5090 ( .A(b[211]), .B(n4273), .Z(n4274) );
  XOR U5091 ( .A(n4276), .B(n4277), .Z(n4273) );
  ANDN U5092 ( .B(n4278), .A(n882), .Z(n4276) );
  XNOR U5093 ( .A(a[210]), .B(n4279), .Z(n882) );
  IV U5094 ( .A(n4277), .Z(n4279) );
  XNOR U5095 ( .A(b[210]), .B(n4277), .Z(n4278) );
  XOR U5096 ( .A(n4280), .B(n4281), .Z(n4277) );
  ANDN U5097 ( .B(n4282), .A(n884), .Z(n4280) );
  XNOR U5098 ( .A(a[209]), .B(n4283), .Z(n884) );
  IV U5099 ( .A(n4281), .Z(n4283) );
  XNOR U5100 ( .A(b[209]), .B(n4281), .Z(n4282) );
  XOR U5101 ( .A(n4284), .B(n4285), .Z(n4281) );
  ANDN U5102 ( .B(n4286), .A(n885), .Z(n4284) );
  XNOR U5103 ( .A(a[208]), .B(n4287), .Z(n885) );
  IV U5104 ( .A(n4285), .Z(n4287) );
  XNOR U5105 ( .A(b[208]), .B(n4285), .Z(n4286) );
  XOR U5106 ( .A(n4288), .B(n4289), .Z(n4285) );
  ANDN U5107 ( .B(n4290), .A(n886), .Z(n4288) );
  XNOR U5108 ( .A(a[207]), .B(n4291), .Z(n886) );
  IV U5109 ( .A(n4289), .Z(n4291) );
  XNOR U5110 ( .A(b[207]), .B(n4289), .Z(n4290) );
  XOR U5111 ( .A(n4292), .B(n4293), .Z(n4289) );
  ANDN U5112 ( .B(n4294), .A(n887), .Z(n4292) );
  XNOR U5113 ( .A(a[206]), .B(n4295), .Z(n887) );
  IV U5114 ( .A(n4293), .Z(n4295) );
  XNOR U5115 ( .A(b[206]), .B(n4293), .Z(n4294) );
  XOR U5116 ( .A(n4296), .B(n4297), .Z(n4293) );
  ANDN U5117 ( .B(n4298), .A(n888), .Z(n4296) );
  XNOR U5118 ( .A(a[205]), .B(n4299), .Z(n888) );
  IV U5119 ( .A(n4297), .Z(n4299) );
  XNOR U5120 ( .A(b[205]), .B(n4297), .Z(n4298) );
  XOR U5121 ( .A(n4300), .B(n4301), .Z(n4297) );
  ANDN U5122 ( .B(n4302), .A(n889), .Z(n4300) );
  XNOR U5123 ( .A(a[204]), .B(n4303), .Z(n889) );
  IV U5124 ( .A(n4301), .Z(n4303) );
  XNOR U5125 ( .A(b[204]), .B(n4301), .Z(n4302) );
  XOR U5126 ( .A(n4304), .B(n4305), .Z(n4301) );
  ANDN U5127 ( .B(n4306), .A(n890), .Z(n4304) );
  XNOR U5128 ( .A(a[203]), .B(n4307), .Z(n890) );
  IV U5129 ( .A(n4305), .Z(n4307) );
  XNOR U5130 ( .A(b[203]), .B(n4305), .Z(n4306) );
  XOR U5131 ( .A(n4308), .B(n4309), .Z(n4305) );
  ANDN U5132 ( .B(n4310), .A(n891), .Z(n4308) );
  XNOR U5133 ( .A(a[202]), .B(n4311), .Z(n891) );
  IV U5134 ( .A(n4309), .Z(n4311) );
  XNOR U5135 ( .A(b[202]), .B(n4309), .Z(n4310) );
  XOR U5136 ( .A(n4312), .B(n4313), .Z(n4309) );
  ANDN U5137 ( .B(n4314), .A(n892), .Z(n4312) );
  XNOR U5138 ( .A(a[201]), .B(n4315), .Z(n892) );
  IV U5139 ( .A(n4313), .Z(n4315) );
  XNOR U5140 ( .A(b[201]), .B(n4313), .Z(n4314) );
  XOR U5141 ( .A(n4316), .B(n4317), .Z(n4313) );
  ANDN U5142 ( .B(n4318), .A(n893), .Z(n4316) );
  XNOR U5143 ( .A(a[200]), .B(n4319), .Z(n893) );
  IV U5144 ( .A(n4317), .Z(n4319) );
  XNOR U5145 ( .A(b[200]), .B(n4317), .Z(n4318) );
  XOR U5146 ( .A(n4320), .B(n4321), .Z(n4317) );
  ANDN U5147 ( .B(n4322), .A(n896), .Z(n4320) );
  XNOR U5148 ( .A(a[199]), .B(n4323), .Z(n896) );
  IV U5149 ( .A(n4321), .Z(n4323) );
  XNOR U5150 ( .A(b[199]), .B(n4321), .Z(n4322) );
  XOR U5151 ( .A(n4324), .B(n4325), .Z(n4321) );
  ANDN U5152 ( .B(n4326), .A(n897), .Z(n4324) );
  XNOR U5153 ( .A(a[198]), .B(n4327), .Z(n897) );
  IV U5154 ( .A(n4325), .Z(n4327) );
  XNOR U5155 ( .A(b[198]), .B(n4325), .Z(n4326) );
  XOR U5156 ( .A(n4328), .B(n4329), .Z(n4325) );
  ANDN U5157 ( .B(n4330), .A(n898), .Z(n4328) );
  XNOR U5158 ( .A(a[197]), .B(n4331), .Z(n898) );
  IV U5159 ( .A(n4329), .Z(n4331) );
  XNOR U5160 ( .A(b[197]), .B(n4329), .Z(n4330) );
  XOR U5161 ( .A(n4332), .B(n4333), .Z(n4329) );
  ANDN U5162 ( .B(n4334), .A(n899), .Z(n4332) );
  XNOR U5163 ( .A(a[196]), .B(n4335), .Z(n899) );
  IV U5164 ( .A(n4333), .Z(n4335) );
  XNOR U5165 ( .A(b[196]), .B(n4333), .Z(n4334) );
  XOR U5166 ( .A(n4336), .B(n4337), .Z(n4333) );
  ANDN U5167 ( .B(n4338), .A(n900), .Z(n4336) );
  XNOR U5168 ( .A(a[195]), .B(n4339), .Z(n900) );
  IV U5169 ( .A(n4337), .Z(n4339) );
  XNOR U5170 ( .A(b[195]), .B(n4337), .Z(n4338) );
  XOR U5171 ( .A(n4340), .B(n4341), .Z(n4337) );
  ANDN U5172 ( .B(n4342), .A(n901), .Z(n4340) );
  XNOR U5173 ( .A(a[194]), .B(n4343), .Z(n901) );
  IV U5174 ( .A(n4341), .Z(n4343) );
  XNOR U5175 ( .A(b[194]), .B(n4341), .Z(n4342) );
  XOR U5176 ( .A(n4344), .B(n4345), .Z(n4341) );
  ANDN U5177 ( .B(n4346), .A(n902), .Z(n4344) );
  XNOR U5178 ( .A(a[193]), .B(n4347), .Z(n902) );
  IV U5179 ( .A(n4345), .Z(n4347) );
  XNOR U5180 ( .A(b[193]), .B(n4345), .Z(n4346) );
  XOR U5181 ( .A(n4348), .B(n4349), .Z(n4345) );
  ANDN U5182 ( .B(n4350), .A(n903), .Z(n4348) );
  XNOR U5183 ( .A(a[192]), .B(n4351), .Z(n903) );
  IV U5184 ( .A(n4349), .Z(n4351) );
  XNOR U5185 ( .A(b[192]), .B(n4349), .Z(n4350) );
  XOR U5186 ( .A(n4352), .B(n4353), .Z(n4349) );
  ANDN U5187 ( .B(n4354), .A(n904), .Z(n4352) );
  XNOR U5188 ( .A(a[191]), .B(n4355), .Z(n904) );
  IV U5189 ( .A(n4353), .Z(n4355) );
  XNOR U5190 ( .A(b[191]), .B(n4353), .Z(n4354) );
  XOR U5191 ( .A(n4356), .B(n4357), .Z(n4353) );
  ANDN U5192 ( .B(n4358), .A(n905), .Z(n4356) );
  XNOR U5193 ( .A(a[190]), .B(n4359), .Z(n905) );
  IV U5194 ( .A(n4357), .Z(n4359) );
  XNOR U5195 ( .A(b[190]), .B(n4357), .Z(n4358) );
  XOR U5196 ( .A(n4360), .B(n4361), .Z(n4357) );
  ANDN U5197 ( .B(n4362), .A(n907), .Z(n4360) );
  XNOR U5198 ( .A(a[189]), .B(n4363), .Z(n907) );
  IV U5199 ( .A(n4361), .Z(n4363) );
  XNOR U5200 ( .A(b[189]), .B(n4361), .Z(n4362) );
  XOR U5201 ( .A(n4364), .B(n4365), .Z(n4361) );
  ANDN U5202 ( .B(n4366), .A(n908), .Z(n4364) );
  XNOR U5203 ( .A(a[188]), .B(n4367), .Z(n908) );
  IV U5204 ( .A(n4365), .Z(n4367) );
  XNOR U5205 ( .A(b[188]), .B(n4365), .Z(n4366) );
  XOR U5206 ( .A(n4368), .B(n4369), .Z(n4365) );
  ANDN U5207 ( .B(n4370), .A(n909), .Z(n4368) );
  XNOR U5208 ( .A(a[187]), .B(n4371), .Z(n909) );
  IV U5209 ( .A(n4369), .Z(n4371) );
  XNOR U5210 ( .A(b[187]), .B(n4369), .Z(n4370) );
  XOR U5211 ( .A(n4372), .B(n4373), .Z(n4369) );
  ANDN U5212 ( .B(n4374), .A(n910), .Z(n4372) );
  XNOR U5213 ( .A(a[186]), .B(n4375), .Z(n910) );
  IV U5214 ( .A(n4373), .Z(n4375) );
  XNOR U5215 ( .A(b[186]), .B(n4373), .Z(n4374) );
  XOR U5216 ( .A(n4376), .B(n4377), .Z(n4373) );
  ANDN U5217 ( .B(n4378), .A(n911), .Z(n4376) );
  XNOR U5218 ( .A(a[185]), .B(n4379), .Z(n911) );
  IV U5219 ( .A(n4377), .Z(n4379) );
  XNOR U5220 ( .A(b[185]), .B(n4377), .Z(n4378) );
  XOR U5221 ( .A(n4380), .B(n4381), .Z(n4377) );
  ANDN U5222 ( .B(n4382), .A(n912), .Z(n4380) );
  XNOR U5223 ( .A(a[184]), .B(n4383), .Z(n912) );
  IV U5224 ( .A(n4381), .Z(n4383) );
  XNOR U5225 ( .A(b[184]), .B(n4381), .Z(n4382) );
  XOR U5226 ( .A(n4384), .B(n4385), .Z(n4381) );
  ANDN U5227 ( .B(n4386), .A(n913), .Z(n4384) );
  XNOR U5228 ( .A(a[183]), .B(n4387), .Z(n913) );
  IV U5229 ( .A(n4385), .Z(n4387) );
  XNOR U5230 ( .A(b[183]), .B(n4385), .Z(n4386) );
  XOR U5231 ( .A(n4388), .B(n4389), .Z(n4385) );
  ANDN U5232 ( .B(n4390), .A(n914), .Z(n4388) );
  XNOR U5233 ( .A(a[182]), .B(n4391), .Z(n914) );
  IV U5234 ( .A(n4389), .Z(n4391) );
  XNOR U5235 ( .A(b[182]), .B(n4389), .Z(n4390) );
  XOR U5236 ( .A(n4392), .B(n4393), .Z(n4389) );
  ANDN U5237 ( .B(n4394), .A(n915), .Z(n4392) );
  XNOR U5238 ( .A(a[181]), .B(n4395), .Z(n915) );
  IV U5239 ( .A(n4393), .Z(n4395) );
  XNOR U5240 ( .A(b[181]), .B(n4393), .Z(n4394) );
  XOR U5241 ( .A(n4396), .B(n4397), .Z(n4393) );
  ANDN U5242 ( .B(n4398), .A(n916), .Z(n4396) );
  XNOR U5243 ( .A(a[180]), .B(n4399), .Z(n916) );
  IV U5244 ( .A(n4397), .Z(n4399) );
  XNOR U5245 ( .A(b[180]), .B(n4397), .Z(n4398) );
  XOR U5246 ( .A(n4400), .B(n4401), .Z(n4397) );
  ANDN U5247 ( .B(n4402), .A(n918), .Z(n4400) );
  XNOR U5248 ( .A(a[179]), .B(n4403), .Z(n918) );
  IV U5249 ( .A(n4401), .Z(n4403) );
  XNOR U5250 ( .A(b[179]), .B(n4401), .Z(n4402) );
  XOR U5251 ( .A(n4404), .B(n4405), .Z(n4401) );
  ANDN U5252 ( .B(n4406), .A(n919), .Z(n4404) );
  XNOR U5253 ( .A(a[178]), .B(n4407), .Z(n919) );
  IV U5254 ( .A(n4405), .Z(n4407) );
  XNOR U5255 ( .A(b[178]), .B(n4405), .Z(n4406) );
  XOR U5256 ( .A(n4408), .B(n4409), .Z(n4405) );
  ANDN U5257 ( .B(n4410), .A(n920), .Z(n4408) );
  XNOR U5258 ( .A(a[177]), .B(n4411), .Z(n920) );
  IV U5259 ( .A(n4409), .Z(n4411) );
  XNOR U5260 ( .A(b[177]), .B(n4409), .Z(n4410) );
  XOR U5261 ( .A(n4412), .B(n4413), .Z(n4409) );
  ANDN U5262 ( .B(n4414), .A(n921), .Z(n4412) );
  XNOR U5263 ( .A(a[176]), .B(n4415), .Z(n921) );
  IV U5264 ( .A(n4413), .Z(n4415) );
  XNOR U5265 ( .A(b[176]), .B(n4413), .Z(n4414) );
  XOR U5266 ( .A(n4416), .B(n4417), .Z(n4413) );
  ANDN U5267 ( .B(n4418), .A(n922), .Z(n4416) );
  XNOR U5268 ( .A(a[175]), .B(n4419), .Z(n922) );
  IV U5269 ( .A(n4417), .Z(n4419) );
  XNOR U5270 ( .A(b[175]), .B(n4417), .Z(n4418) );
  XOR U5271 ( .A(n4420), .B(n4421), .Z(n4417) );
  ANDN U5272 ( .B(n4422), .A(n923), .Z(n4420) );
  XNOR U5273 ( .A(a[174]), .B(n4423), .Z(n923) );
  IV U5274 ( .A(n4421), .Z(n4423) );
  XNOR U5275 ( .A(b[174]), .B(n4421), .Z(n4422) );
  XOR U5276 ( .A(n4424), .B(n4425), .Z(n4421) );
  ANDN U5277 ( .B(n4426), .A(n924), .Z(n4424) );
  XNOR U5278 ( .A(a[173]), .B(n4427), .Z(n924) );
  IV U5279 ( .A(n4425), .Z(n4427) );
  XNOR U5280 ( .A(b[173]), .B(n4425), .Z(n4426) );
  XOR U5281 ( .A(n4428), .B(n4429), .Z(n4425) );
  ANDN U5282 ( .B(n4430), .A(n925), .Z(n4428) );
  XNOR U5283 ( .A(a[172]), .B(n4431), .Z(n925) );
  IV U5284 ( .A(n4429), .Z(n4431) );
  XNOR U5285 ( .A(b[172]), .B(n4429), .Z(n4430) );
  XOR U5286 ( .A(n4432), .B(n4433), .Z(n4429) );
  ANDN U5287 ( .B(n4434), .A(n926), .Z(n4432) );
  XNOR U5288 ( .A(a[171]), .B(n4435), .Z(n926) );
  IV U5289 ( .A(n4433), .Z(n4435) );
  XNOR U5290 ( .A(b[171]), .B(n4433), .Z(n4434) );
  XOR U5291 ( .A(n4436), .B(n4437), .Z(n4433) );
  ANDN U5292 ( .B(n4438), .A(n927), .Z(n4436) );
  XNOR U5293 ( .A(a[170]), .B(n4439), .Z(n927) );
  IV U5294 ( .A(n4437), .Z(n4439) );
  XNOR U5295 ( .A(b[170]), .B(n4437), .Z(n4438) );
  XOR U5296 ( .A(n4440), .B(n4441), .Z(n4437) );
  ANDN U5297 ( .B(n4442), .A(n929), .Z(n4440) );
  XNOR U5298 ( .A(a[169]), .B(n4443), .Z(n929) );
  IV U5299 ( .A(n4441), .Z(n4443) );
  XNOR U5300 ( .A(b[169]), .B(n4441), .Z(n4442) );
  XOR U5301 ( .A(n4444), .B(n4445), .Z(n4441) );
  ANDN U5302 ( .B(n4446), .A(n930), .Z(n4444) );
  XNOR U5303 ( .A(a[168]), .B(n4447), .Z(n930) );
  IV U5304 ( .A(n4445), .Z(n4447) );
  XNOR U5305 ( .A(b[168]), .B(n4445), .Z(n4446) );
  XOR U5306 ( .A(n4448), .B(n4449), .Z(n4445) );
  ANDN U5307 ( .B(n4450), .A(n931), .Z(n4448) );
  XNOR U5308 ( .A(a[167]), .B(n4451), .Z(n931) );
  IV U5309 ( .A(n4449), .Z(n4451) );
  XNOR U5310 ( .A(b[167]), .B(n4449), .Z(n4450) );
  XOR U5311 ( .A(n4452), .B(n4453), .Z(n4449) );
  ANDN U5312 ( .B(n4454), .A(n932), .Z(n4452) );
  XNOR U5313 ( .A(a[166]), .B(n4455), .Z(n932) );
  IV U5314 ( .A(n4453), .Z(n4455) );
  XNOR U5315 ( .A(b[166]), .B(n4453), .Z(n4454) );
  XOR U5316 ( .A(n4456), .B(n4457), .Z(n4453) );
  ANDN U5317 ( .B(n4458), .A(n933), .Z(n4456) );
  XNOR U5318 ( .A(a[165]), .B(n4459), .Z(n933) );
  IV U5319 ( .A(n4457), .Z(n4459) );
  XNOR U5320 ( .A(b[165]), .B(n4457), .Z(n4458) );
  XOR U5321 ( .A(n4460), .B(n4461), .Z(n4457) );
  ANDN U5322 ( .B(n4462), .A(n934), .Z(n4460) );
  XNOR U5323 ( .A(a[164]), .B(n4463), .Z(n934) );
  IV U5324 ( .A(n4461), .Z(n4463) );
  XNOR U5325 ( .A(b[164]), .B(n4461), .Z(n4462) );
  XOR U5326 ( .A(n4464), .B(n4465), .Z(n4461) );
  ANDN U5327 ( .B(n4466), .A(n935), .Z(n4464) );
  XNOR U5328 ( .A(a[163]), .B(n4467), .Z(n935) );
  IV U5329 ( .A(n4465), .Z(n4467) );
  XNOR U5330 ( .A(b[163]), .B(n4465), .Z(n4466) );
  XOR U5331 ( .A(n4468), .B(n4469), .Z(n4465) );
  ANDN U5332 ( .B(n4470), .A(n936), .Z(n4468) );
  XNOR U5333 ( .A(a[162]), .B(n4471), .Z(n936) );
  IV U5334 ( .A(n4469), .Z(n4471) );
  XNOR U5335 ( .A(b[162]), .B(n4469), .Z(n4470) );
  XOR U5336 ( .A(n4472), .B(n4473), .Z(n4469) );
  ANDN U5337 ( .B(n4474), .A(n937), .Z(n4472) );
  XNOR U5338 ( .A(a[161]), .B(n4475), .Z(n937) );
  IV U5339 ( .A(n4473), .Z(n4475) );
  XNOR U5340 ( .A(b[161]), .B(n4473), .Z(n4474) );
  XOR U5341 ( .A(n4476), .B(n4477), .Z(n4473) );
  ANDN U5342 ( .B(n4478), .A(n938), .Z(n4476) );
  XNOR U5343 ( .A(a[160]), .B(n4479), .Z(n938) );
  IV U5344 ( .A(n4477), .Z(n4479) );
  XNOR U5345 ( .A(b[160]), .B(n4477), .Z(n4478) );
  XOR U5346 ( .A(n4480), .B(n4481), .Z(n4477) );
  ANDN U5347 ( .B(n4482), .A(n940), .Z(n4480) );
  XNOR U5348 ( .A(a[159]), .B(n4483), .Z(n940) );
  IV U5349 ( .A(n4481), .Z(n4483) );
  XNOR U5350 ( .A(b[159]), .B(n4481), .Z(n4482) );
  XOR U5351 ( .A(n4484), .B(n4485), .Z(n4481) );
  ANDN U5352 ( .B(n4486), .A(n941), .Z(n4484) );
  XNOR U5353 ( .A(a[158]), .B(n4487), .Z(n941) );
  IV U5354 ( .A(n4485), .Z(n4487) );
  XNOR U5355 ( .A(b[158]), .B(n4485), .Z(n4486) );
  XOR U5356 ( .A(n4488), .B(n4489), .Z(n4485) );
  ANDN U5357 ( .B(n4490), .A(n942), .Z(n4488) );
  XNOR U5358 ( .A(a[157]), .B(n4491), .Z(n942) );
  IV U5359 ( .A(n4489), .Z(n4491) );
  XNOR U5360 ( .A(b[157]), .B(n4489), .Z(n4490) );
  XOR U5361 ( .A(n4492), .B(n4493), .Z(n4489) );
  ANDN U5362 ( .B(n4494), .A(n943), .Z(n4492) );
  XNOR U5363 ( .A(a[156]), .B(n4495), .Z(n943) );
  IV U5364 ( .A(n4493), .Z(n4495) );
  XNOR U5365 ( .A(b[156]), .B(n4493), .Z(n4494) );
  XOR U5366 ( .A(n4496), .B(n4497), .Z(n4493) );
  ANDN U5367 ( .B(n4498), .A(n944), .Z(n4496) );
  XNOR U5368 ( .A(a[155]), .B(n4499), .Z(n944) );
  IV U5369 ( .A(n4497), .Z(n4499) );
  XNOR U5370 ( .A(b[155]), .B(n4497), .Z(n4498) );
  XOR U5371 ( .A(n4500), .B(n4501), .Z(n4497) );
  ANDN U5372 ( .B(n4502), .A(n945), .Z(n4500) );
  XNOR U5373 ( .A(a[154]), .B(n4503), .Z(n945) );
  IV U5374 ( .A(n4501), .Z(n4503) );
  XNOR U5375 ( .A(b[154]), .B(n4501), .Z(n4502) );
  XOR U5376 ( .A(n4504), .B(n4505), .Z(n4501) );
  ANDN U5377 ( .B(n4506), .A(n946), .Z(n4504) );
  XNOR U5378 ( .A(a[153]), .B(n4507), .Z(n946) );
  IV U5379 ( .A(n4505), .Z(n4507) );
  XNOR U5380 ( .A(b[153]), .B(n4505), .Z(n4506) );
  XOR U5381 ( .A(n4508), .B(n4509), .Z(n4505) );
  ANDN U5382 ( .B(n4510), .A(n947), .Z(n4508) );
  XNOR U5383 ( .A(a[152]), .B(n4511), .Z(n947) );
  IV U5384 ( .A(n4509), .Z(n4511) );
  XNOR U5385 ( .A(b[152]), .B(n4509), .Z(n4510) );
  XOR U5386 ( .A(n4512), .B(n4513), .Z(n4509) );
  ANDN U5387 ( .B(n4514), .A(n948), .Z(n4512) );
  XNOR U5388 ( .A(a[151]), .B(n4515), .Z(n948) );
  IV U5389 ( .A(n4513), .Z(n4515) );
  XNOR U5390 ( .A(b[151]), .B(n4513), .Z(n4514) );
  XOR U5391 ( .A(n4516), .B(n4517), .Z(n4513) );
  ANDN U5392 ( .B(n4518), .A(n949), .Z(n4516) );
  XNOR U5393 ( .A(a[150]), .B(n4519), .Z(n949) );
  IV U5394 ( .A(n4517), .Z(n4519) );
  XNOR U5395 ( .A(b[150]), .B(n4517), .Z(n4518) );
  XOR U5396 ( .A(n4520), .B(n4521), .Z(n4517) );
  ANDN U5397 ( .B(n4522), .A(n951), .Z(n4520) );
  XNOR U5398 ( .A(a[149]), .B(n4523), .Z(n951) );
  IV U5399 ( .A(n4521), .Z(n4523) );
  XNOR U5400 ( .A(b[149]), .B(n4521), .Z(n4522) );
  XOR U5401 ( .A(n4524), .B(n4525), .Z(n4521) );
  ANDN U5402 ( .B(n4526), .A(n952), .Z(n4524) );
  XNOR U5403 ( .A(a[148]), .B(n4527), .Z(n952) );
  IV U5404 ( .A(n4525), .Z(n4527) );
  XNOR U5405 ( .A(b[148]), .B(n4525), .Z(n4526) );
  XOR U5406 ( .A(n4528), .B(n4529), .Z(n4525) );
  ANDN U5407 ( .B(n4530), .A(n953), .Z(n4528) );
  XNOR U5408 ( .A(a[147]), .B(n4531), .Z(n953) );
  IV U5409 ( .A(n4529), .Z(n4531) );
  XNOR U5410 ( .A(b[147]), .B(n4529), .Z(n4530) );
  XOR U5411 ( .A(n4532), .B(n4533), .Z(n4529) );
  ANDN U5412 ( .B(n4534), .A(n954), .Z(n4532) );
  XNOR U5413 ( .A(a[146]), .B(n4535), .Z(n954) );
  IV U5414 ( .A(n4533), .Z(n4535) );
  XNOR U5415 ( .A(b[146]), .B(n4533), .Z(n4534) );
  XOR U5416 ( .A(n4536), .B(n4537), .Z(n4533) );
  ANDN U5417 ( .B(n4538), .A(n955), .Z(n4536) );
  XNOR U5418 ( .A(a[145]), .B(n4539), .Z(n955) );
  IV U5419 ( .A(n4537), .Z(n4539) );
  XNOR U5420 ( .A(b[145]), .B(n4537), .Z(n4538) );
  XOR U5421 ( .A(n4540), .B(n4541), .Z(n4537) );
  ANDN U5422 ( .B(n4542), .A(n956), .Z(n4540) );
  XNOR U5423 ( .A(a[144]), .B(n4543), .Z(n956) );
  IV U5424 ( .A(n4541), .Z(n4543) );
  XNOR U5425 ( .A(b[144]), .B(n4541), .Z(n4542) );
  XOR U5426 ( .A(n4544), .B(n4545), .Z(n4541) );
  ANDN U5427 ( .B(n4546), .A(n957), .Z(n4544) );
  XNOR U5428 ( .A(a[143]), .B(n4547), .Z(n957) );
  IV U5429 ( .A(n4545), .Z(n4547) );
  XNOR U5430 ( .A(b[143]), .B(n4545), .Z(n4546) );
  XOR U5431 ( .A(n4548), .B(n4549), .Z(n4545) );
  ANDN U5432 ( .B(n4550), .A(n958), .Z(n4548) );
  XNOR U5433 ( .A(a[142]), .B(n4551), .Z(n958) );
  IV U5434 ( .A(n4549), .Z(n4551) );
  XNOR U5435 ( .A(b[142]), .B(n4549), .Z(n4550) );
  XOR U5436 ( .A(n4552), .B(n4553), .Z(n4549) );
  ANDN U5437 ( .B(n4554), .A(n959), .Z(n4552) );
  XNOR U5438 ( .A(a[141]), .B(n4555), .Z(n959) );
  IV U5439 ( .A(n4553), .Z(n4555) );
  XNOR U5440 ( .A(b[141]), .B(n4553), .Z(n4554) );
  XOR U5441 ( .A(n4556), .B(n4557), .Z(n4553) );
  ANDN U5442 ( .B(n4558), .A(n960), .Z(n4556) );
  XNOR U5443 ( .A(a[140]), .B(n4559), .Z(n960) );
  IV U5444 ( .A(n4557), .Z(n4559) );
  XNOR U5445 ( .A(b[140]), .B(n4557), .Z(n4558) );
  XOR U5446 ( .A(n4560), .B(n4561), .Z(n4557) );
  ANDN U5447 ( .B(n4562), .A(n962), .Z(n4560) );
  XNOR U5448 ( .A(a[139]), .B(n4563), .Z(n962) );
  IV U5449 ( .A(n4561), .Z(n4563) );
  XNOR U5450 ( .A(b[139]), .B(n4561), .Z(n4562) );
  XOR U5451 ( .A(n4564), .B(n4565), .Z(n4561) );
  ANDN U5452 ( .B(n4566), .A(n963), .Z(n4564) );
  XNOR U5453 ( .A(a[138]), .B(n4567), .Z(n963) );
  IV U5454 ( .A(n4565), .Z(n4567) );
  XNOR U5455 ( .A(b[138]), .B(n4565), .Z(n4566) );
  XOR U5456 ( .A(n4568), .B(n4569), .Z(n4565) );
  ANDN U5457 ( .B(n4570), .A(n964), .Z(n4568) );
  XNOR U5458 ( .A(a[137]), .B(n4571), .Z(n964) );
  IV U5459 ( .A(n4569), .Z(n4571) );
  XNOR U5460 ( .A(b[137]), .B(n4569), .Z(n4570) );
  XOR U5461 ( .A(n4572), .B(n4573), .Z(n4569) );
  ANDN U5462 ( .B(n4574), .A(n965), .Z(n4572) );
  XNOR U5463 ( .A(a[136]), .B(n4575), .Z(n965) );
  IV U5464 ( .A(n4573), .Z(n4575) );
  XNOR U5465 ( .A(b[136]), .B(n4573), .Z(n4574) );
  XOR U5466 ( .A(n4576), .B(n4577), .Z(n4573) );
  ANDN U5467 ( .B(n4578), .A(n966), .Z(n4576) );
  XNOR U5468 ( .A(a[135]), .B(n4579), .Z(n966) );
  IV U5469 ( .A(n4577), .Z(n4579) );
  XNOR U5470 ( .A(b[135]), .B(n4577), .Z(n4578) );
  XOR U5471 ( .A(n4580), .B(n4581), .Z(n4577) );
  ANDN U5472 ( .B(n4582), .A(n967), .Z(n4580) );
  XNOR U5473 ( .A(a[134]), .B(n4583), .Z(n967) );
  IV U5474 ( .A(n4581), .Z(n4583) );
  XNOR U5475 ( .A(b[134]), .B(n4581), .Z(n4582) );
  XOR U5476 ( .A(n4584), .B(n4585), .Z(n4581) );
  ANDN U5477 ( .B(n4586), .A(n968), .Z(n4584) );
  XNOR U5478 ( .A(a[133]), .B(n4587), .Z(n968) );
  IV U5479 ( .A(n4585), .Z(n4587) );
  XNOR U5480 ( .A(b[133]), .B(n4585), .Z(n4586) );
  XOR U5481 ( .A(n4588), .B(n4589), .Z(n4585) );
  ANDN U5482 ( .B(n4590), .A(n969), .Z(n4588) );
  XNOR U5483 ( .A(a[132]), .B(n4591), .Z(n969) );
  IV U5484 ( .A(n4589), .Z(n4591) );
  XNOR U5485 ( .A(b[132]), .B(n4589), .Z(n4590) );
  XOR U5486 ( .A(n4592), .B(n4593), .Z(n4589) );
  ANDN U5487 ( .B(n4594), .A(n970), .Z(n4592) );
  XNOR U5488 ( .A(a[131]), .B(n4595), .Z(n970) );
  IV U5489 ( .A(n4593), .Z(n4595) );
  XNOR U5490 ( .A(b[131]), .B(n4593), .Z(n4594) );
  XOR U5491 ( .A(n4596), .B(n4597), .Z(n4593) );
  ANDN U5492 ( .B(n4598), .A(n971), .Z(n4596) );
  XNOR U5493 ( .A(a[130]), .B(n4599), .Z(n971) );
  IV U5494 ( .A(n4597), .Z(n4599) );
  XNOR U5495 ( .A(b[130]), .B(n4597), .Z(n4598) );
  XOR U5496 ( .A(n4600), .B(n4601), .Z(n4597) );
  ANDN U5497 ( .B(n4602), .A(n973), .Z(n4600) );
  XNOR U5498 ( .A(a[129]), .B(n4603), .Z(n973) );
  IV U5499 ( .A(n4601), .Z(n4603) );
  XNOR U5500 ( .A(b[129]), .B(n4601), .Z(n4602) );
  XOR U5501 ( .A(n4604), .B(n4605), .Z(n4601) );
  ANDN U5502 ( .B(n4606), .A(n974), .Z(n4604) );
  XNOR U5503 ( .A(a[128]), .B(n4607), .Z(n974) );
  IV U5504 ( .A(n4605), .Z(n4607) );
  XNOR U5505 ( .A(b[128]), .B(n4605), .Z(n4606) );
  XOR U5506 ( .A(n4608), .B(n4609), .Z(n4605) );
  ANDN U5507 ( .B(n4610), .A(n975), .Z(n4608) );
  XNOR U5508 ( .A(a[127]), .B(n4611), .Z(n975) );
  IV U5509 ( .A(n4609), .Z(n4611) );
  XNOR U5510 ( .A(b[127]), .B(n4609), .Z(n4610) );
  XOR U5511 ( .A(n4612), .B(n4613), .Z(n4609) );
  ANDN U5512 ( .B(n4614), .A(n976), .Z(n4612) );
  XNOR U5513 ( .A(a[126]), .B(n4615), .Z(n976) );
  IV U5514 ( .A(n4613), .Z(n4615) );
  XNOR U5515 ( .A(b[126]), .B(n4613), .Z(n4614) );
  XOR U5516 ( .A(n4616), .B(n4617), .Z(n4613) );
  ANDN U5517 ( .B(n4618), .A(n977), .Z(n4616) );
  XNOR U5518 ( .A(a[125]), .B(n4619), .Z(n977) );
  IV U5519 ( .A(n4617), .Z(n4619) );
  XNOR U5520 ( .A(b[125]), .B(n4617), .Z(n4618) );
  XOR U5521 ( .A(n4620), .B(n4621), .Z(n4617) );
  ANDN U5522 ( .B(n4622), .A(n978), .Z(n4620) );
  XNOR U5523 ( .A(a[124]), .B(n4623), .Z(n978) );
  IV U5524 ( .A(n4621), .Z(n4623) );
  XNOR U5525 ( .A(b[124]), .B(n4621), .Z(n4622) );
  XOR U5526 ( .A(n4624), .B(n4625), .Z(n4621) );
  ANDN U5527 ( .B(n4626), .A(n979), .Z(n4624) );
  XNOR U5528 ( .A(a[123]), .B(n4627), .Z(n979) );
  IV U5529 ( .A(n4625), .Z(n4627) );
  XNOR U5530 ( .A(b[123]), .B(n4625), .Z(n4626) );
  XOR U5531 ( .A(n4628), .B(n4629), .Z(n4625) );
  ANDN U5532 ( .B(n4630), .A(n980), .Z(n4628) );
  XNOR U5533 ( .A(a[122]), .B(n4631), .Z(n980) );
  IV U5534 ( .A(n4629), .Z(n4631) );
  XNOR U5535 ( .A(b[122]), .B(n4629), .Z(n4630) );
  XOR U5536 ( .A(n4632), .B(n4633), .Z(n4629) );
  ANDN U5537 ( .B(n4634), .A(n981), .Z(n4632) );
  XNOR U5538 ( .A(a[121]), .B(n4635), .Z(n981) );
  IV U5539 ( .A(n4633), .Z(n4635) );
  XNOR U5540 ( .A(b[121]), .B(n4633), .Z(n4634) );
  XOR U5541 ( .A(n4636), .B(n4637), .Z(n4633) );
  ANDN U5542 ( .B(n4638), .A(n982), .Z(n4636) );
  XNOR U5543 ( .A(a[120]), .B(n4639), .Z(n982) );
  IV U5544 ( .A(n4637), .Z(n4639) );
  XNOR U5545 ( .A(b[120]), .B(n4637), .Z(n4638) );
  XOR U5546 ( .A(n4640), .B(n4641), .Z(n4637) );
  ANDN U5547 ( .B(n4642), .A(n984), .Z(n4640) );
  XNOR U5548 ( .A(a[119]), .B(n4643), .Z(n984) );
  IV U5549 ( .A(n4641), .Z(n4643) );
  XNOR U5550 ( .A(b[119]), .B(n4641), .Z(n4642) );
  XOR U5551 ( .A(n4644), .B(n4645), .Z(n4641) );
  ANDN U5552 ( .B(n4646), .A(n985), .Z(n4644) );
  XNOR U5553 ( .A(a[118]), .B(n4647), .Z(n985) );
  IV U5554 ( .A(n4645), .Z(n4647) );
  XNOR U5555 ( .A(b[118]), .B(n4645), .Z(n4646) );
  XOR U5556 ( .A(n4648), .B(n4649), .Z(n4645) );
  ANDN U5557 ( .B(n4650), .A(n986), .Z(n4648) );
  XNOR U5558 ( .A(a[117]), .B(n4651), .Z(n986) );
  IV U5559 ( .A(n4649), .Z(n4651) );
  XNOR U5560 ( .A(b[117]), .B(n4649), .Z(n4650) );
  XOR U5561 ( .A(n4652), .B(n4653), .Z(n4649) );
  ANDN U5562 ( .B(n4654), .A(n987), .Z(n4652) );
  XNOR U5563 ( .A(a[116]), .B(n4655), .Z(n987) );
  IV U5564 ( .A(n4653), .Z(n4655) );
  XNOR U5565 ( .A(b[116]), .B(n4653), .Z(n4654) );
  XOR U5566 ( .A(n4656), .B(n4657), .Z(n4653) );
  ANDN U5567 ( .B(n4658), .A(n988), .Z(n4656) );
  XNOR U5568 ( .A(a[115]), .B(n4659), .Z(n988) );
  IV U5569 ( .A(n4657), .Z(n4659) );
  XNOR U5570 ( .A(b[115]), .B(n4657), .Z(n4658) );
  XOR U5571 ( .A(n4660), .B(n4661), .Z(n4657) );
  ANDN U5572 ( .B(n4662), .A(n989), .Z(n4660) );
  XNOR U5573 ( .A(a[114]), .B(n4663), .Z(n989) );
  IV U5574 ( .A(n4661), .Z(n4663) );
  XNOR U5575 ( .A(b[114]), .B(n4661), .Z(n4662) );
  XOR U5576 ( .A(n4664), .B(n4665), .Z(n4661) );
  ANDN U5577 ( .B(n4666), .A(n990), .Z(n4664) );
  XNOR U5578 ( .A(a[113]), .B(n4667), .Z(n990) );
  IV U5579 ( .A(n4665), .Z(n4667) );
  XNOR U5580 ( .A(b[113]), .B(n4665), .Z(n4666) );
  XOR U5581 ( .A(n4668), .B(n4669), .Z(n4665) );
  ANDN U5582 ( .B(n4670), .A(n991), .Z(n4668) );
  XNOR U5583 ( .A(a[112]), .B(n4671), .Z(n991) );
  IV U5584 ( .A(n4669), .Z(n4671) );
  XNOR U5585 ( .A(b[112]), .B(n4669), .Z(n4670) );
  XOR U5586 ( .A(n4672), .B(n4673), .Z(n4669) );
  ANDN U5587 ( .B(n4674), .A(n992), .Z(n4672) );
  XNOR U5588 ( .A(a[111]), .B(n4675), .Z(n992) );
  IV U5589 ( .A(n4673), .Z(n4675) );
  XNOR U5590 ( .A(b[111]), .B(n4673), .Z(n4674) );
  XOR U5591 ( .A(n4676), .B(n4677), .Z(n4673) );
  ANDN U5592 ( .B(n4678), .A(n993), .Z(n4676) );
  XNOR U5593 ( .A(a[110]), .B(n4679), .Z(n993) );
  IV U5594 ( .A(n4677), .Z(n4679) );
  XNOR U5595 ( .A(b[110]), .B(n4677), .Z(n4678) );
  XOR U5596 ( .A(n4680), .B(n4681), .Z(n4677) );
  ANDN U5597 ( .B(n4682), .A(n995), .Z(n4680) );
  XNOR U5598 ( .A(a[109]), .B(n4683), .Z(n995) );
  IV U5599 ( .A(n4681), .Z(n4683) );
  XNOR U5600 ( .A(b[109]), .B(n4681), .Z(n4682) );
  XOR U5601 ( .A(n4684), .B(n4685), .Z(n4681) );
  ANDN U5602 ( .B(n4686), .A(n996), .Z(n4684) );
  XNOR U5603 ( .A(a[108]), .B(n4687), .Z(n996) );
  IV U5604 ( .A(n4685), .Z(n4687) );
  XNOR U5605 ( .A(b[108]), .B(n4685), .Z(n4686) );
  XOR U5606 ( .A(n4688), .B(n4689), .Z(n4685) );
  ANDN U5607 ( .B(n4690), .A(n997), .Z(n4688) );
  XNOR U5608 ( .A(a[107]), .B(n4691), .Z(n997) );
  IV U5609 ( .A(n4689), .Z(n4691) );
  XNOR U5610 ( .A(b[107]), .B(n4689), .Z(n4690) );
  XOR U5611 ( .A(n4692), .B(n4693), .Z(n4689) );
  ANDN U5612 ( .B(n4694), .A(n998), .Z(n4692) );
  XNOR U5613 ( .A(a[106]), .B(n4695), .Z(n998) );
  IV U5614 ( .A(n4693), .Z(n4695) );
  XNOR U5615 ( .A(b[106]), .B(n4693), .Z(n4694) );
  XOR U5616 ( .A(n4696), .B(n4697), .Z(n4693) );
  ANDN U5617 ( .B(n4698), .A(n999), .Z(n4696) );
  XNOR U5618 ( .A(a[105]), .B(n4699), .Z(n999) );
  IV U5619 ( .A(n4697), .Z(n4699) );
  XNOR U5620 ( .A(b[105]), .B(n4697), .Z(n4698) );
  XOR U5621 ( .A(n4700), .B(n4701), .Z(n4697) );
  ANDN U5622 ( .B(n4702), .A(n1000), .Z(n4700) );
  XNOR U5623 ( .A(a[104]), .B(n4703), .Z(n1000) );
  IV U5624 ( .A(n4701), .Z(n4703) );
  XNOR U5625 ( .A(b[104]), .B(n4701), .Z(n4702) );
  XOR U5626 ( .A(n4704), .B(n4705), .Z(n4701) );
  ANDN U5627 ( .B(n4706), .A(n1001), .Z(n4704) );
  XNOR U5628 ( .A(a[103]), .B(n4707), .Z(n1001) );
  IV U5629 ( .A(n4705), .Z(n4707) );
  XNOR U5630 ( .A(b[103]), .B(n4705), .Z(n4706) );
  XOR U5631 ( .A(n4708), .B(n4709), .Z(n4705) );
  ANDN U5632 ( .B(n4710), .A(n1002), .Z(n4708) );
  XNOR U5633 ( .A(a[102]), .B(n4711), .Z(n1002) );
  IV U5634 ( .A(n4709), .Z(n4711) );
  XNOR U5635 ( .A(b[102]), .B(n4709), .Z(n4710) );
  XOR U5636 ( .A(n4712), .B(n4713), .Z(n4709) );
  ANDN U5637 ( .B(n4714), .A(n1022), .Z(n4712) );
  XNOR U5638 ( .A(a[101]), .B(n4715), .Z(n1022) );
  IV U5639 ( .A(n4713), .Z(n4715) );
  XNOR U5640 ( .A(b[101]), .B(n4713), .Z(n4714) );
  XOR U5641 ( .A(n4716), .B(n4717), .Z(n4713) );
  ANDN U5642 ( .B(n4718), .A(n1073), .Z(n4716) );
  XNOR U5643 ( .A(a[100]), .B(n4719), .Z(n1073) );
  IV U5644 ( .A(n4717), .Z(n4719) );
  XNOR U5645 ( .A(b[100]), .B(n4717), .Z(n4718) );
  XOR U5646 ( .A(n4720), .B(n4721), .Z(n4717) );
  ANDN U5647 ( .B(n4722), .A(n7), .Z(n4720) );
  XNOR U5648 ( .A(a[99]), .B(n4723), .Z(n7) );
  IV U5649 ( .A(n4721), .Z(n4723) );
  XNOR U5650 ( .A(b[99]), .B(n4721), .Z(n4722) );
  XOR U5651 ( .A(n4724), .B(n4725), .Z(n4721) );
  ANDN U5652 ( .B(n4726), .A(n18), .Z(n4724) );
  XNOR U5653 ( .A(a[98]), .B(n4727), .Z(n18) );
  IV U5654 ( .A(n4725), .Z(n4727) );
  XNOR U5655 ( .A(b[98]), .B(n4725), .Z(n4726) );
  XOR U5656 ( .A(n4728), .B(n4729), .Z(n4725) );
  ANDN U5657 ( .B(n4730), .A(n29), .Z(n4728) );
  XNOR U5658 ( .A(a[97]), .B(n4731), .Z(n29) );
  IV U5659 ( .A(n4729), .Z(n4731) );
  XNOR U5660 ( .A(b[97]), .B(n4729), .Z(n4730) );
  XOR U5661 ( .A(n4732), .B(n4733), .Z(n4729) );
  ANDN U5662 ( .B(n4734), .A(n40), .Z(n4732) );
  XNOR U5663 ( .A(a[96]), .B(n4735), .Z(n40) );
  IV U5664 ( .A(n4733), .Z(n4735) );
  XNOR U5665 ( .A(b[96]), .B(n4733), .Z(n4734) );
  XOR U5666 ( .A(n4736), .B(n4737), .Z(n4733) );
  ANDN U5667 ( .B(n4738), .A(n51), .Z(n4736) );
  XNOR U5668 ( .A(a[95]), .B(n4739), .Z(n51) );
  IV U5669 ( .A(n4737), .Z(n4739) );
  XNOR U5670 ( .A(b[95]), .B(n4737), .Z(n4738) );
  XOR U5671 ( .A(n4740), .B(n4741), .Z(n4737) );
  ANDN U5672 ( .B(n4742), .A(n62), .Z(n4740) );
  XNOR U5673 ( .A(a[94]), .B(n4743), .Z(n62) );
  IV U5674 ( .A(n4741), .Z(n4743) );
  XNOR U5675 ( .A(b[94]), .B(n4741), .Z(n4742) );
  XOR U5676 ( .A(n4744), .B(n4745), .Z(n4741) );
  ANDN U5677 ( .B(n4746), .A(n73), .Z(n4744) );
  XNOR U5678 ( .A(a[93]), .B(n4747), .Z(n73) );
  IV U5679 ( .A(n4745), .Z(n4747) );
  XNOR U5680 ( .A(b[93]), .B(n4745), .Z(n4746) );
  XOR U5681 ( .A(n4748), .B(n4749), .Z(n4745) );
  ANDN U5682 ( .B(n4750), .A(n84), .Z(n4748) );
  XNOR U5683 ( .A(a[92]), .B(n4751), .Z(n84) );
  IV U5684 ( .A(n4749), .Z(n4751) );
  XNOR U5685 ( .A(b[92]), .B(n4749), .Z(n4750) );
  XOR U5686 ( .A(n4752), .B(n4753), .Z(n4749) );
  ANDN U5687 ( .B(n4754), .A(n95), .Z(n4752) );
  XNOR U5688 ( .A(a[91]), .B(n4755), .Z(n95) );
  IV U5689 ( .A(n4753), .Z(n4755) );
  XNOR U5690 ( .A(b[91]), .B(n4753), .Z(n4754) );
  XOR U5691 ( .A(n4756), .B(n4757), .Z(n4753) );
  ANDN U5692 ( .B(n4758), .A(n106), .Z(n4756) );
  XNOR U5693 ( .A(a[90]), .B(n4759), .Z(n106) );
  IV U5694 ( .A(n4757), .Z(n4759) );
  XNOR U5695 ( .A(b[90]), .B(n4757), .Z(n4758) );
  XOR U5696 ( .A(n4760), .B(n4761), .Z(n4757) );
  ANDN U5697 ( .B(n4762), .A(n118), .Z(n4760) );
  XNOR U5698 ( .A(a[89]), .B(n4763), .Z(n118) );
  IV U5699 ( .A(n4761), .Z(n4763) );
  XNOR U5700 ( .A(b[89]), .B(n4761), .Z(n4762) );
  XOR U5701 ( .A(n4764), .B(n4765), .Z(n4761) );
  ANDN U5702 ( .B(n4766), .A(n129), .Z(n4764) );
  XNOR U5703 ( .A(a[88]), .B(n4767), .Z(n129) );
  IV U5704 ( .A(n4765), .Z(n4767) );
  XNOR U5705 ( .A(b[88]), .B(n4765), .Z(n4766) );
  XOR U5706 ( .A(n4768), .B(n4769), .Z(n4765) );
  ANDN U5707 ( .B(n4770), .A(n140), .Z(n4768) );
  XNOR U5708 ( .A(a[87]), .B(n4771), .Z(n140) );
  IV U5709 ( .A(n4769), .Z(n4771) );
  XNOR U5710 ( .A(b[87]), .B(n4769), .Z(n4770) );
  XOR U5711 ( .A(n4772), .B(n4773), .Z(n4769) );
  ANDN U5712 ( .B(n4774), .A(n151), .Z(n4772) );
  XNOR U5713 ( .A(a[86]), .B(n4775), .Z(n151) );
  IV U5714 ( .A(n4773), .Z(n4775) );
  XNOR U5715 ( .A(b[86]), .B(n4773), .Z(n4774) );
  XOR U5716 ( .A(n4776), .B(n4777), .Z(n4773) );
  ANDN U5717 ( .B(n4778), .A(n162), .Z(n4776) );
  XNOR U5718 ( .A(a[85]), .B(n4779), .Z(n162) );
  IV U5719 ( .A(n4777), .Z(n4779) );
  XNOR U5720 ( .A(b[85]), .B(n4777), .Z(n4778) );
  XOR U5721 ( .A(n4780), .B(n4781), .Z(n4777) );
  ANDN U5722 ( .B(n4782), .A(n173), .Z(n4780) );
  XNOR U5723 ( .A(a[84]), .B(n4783), .Z(n173) );
  IV U5724 ( .A(n4781), .Z(n4783) );
  XNOR U5725 ( .A(b[84]), .B(n4781), .Z(n4782) );
  XOR U5726 ( .A(n4784), .B(n4785), .Z(n4781) );
  ANDN U5727 ( .B(n4786), .A(n184), .Z(n4784) );
  XNOR U5728 ( .A(a[83]), .B(n4787), .Z(n184) );
  IV U5729 ( .A(n4785), .Z(n4787) );
  XNOR U5730 ( .A(b[83]), .B(n4785), .Z(n4786) );
  XOR U5731 ( .A(n4788), .B(n4789), .Z(n4785) );
  ANDN U5732 ( .B(n4790), .A(n195), .Z(n4788) );
  XNOR U5733 ( .A(a[82]), .B(n4791), .Z(n195) );
  IV U5734 ( .A(n4789), .Z(n4791) );
  XNOR U5735 ( .A(b[82]), .B(n4789), .Z(n4790) );
  XOR U5736 ( .A(n4792), .B(n4793), .Z(n4789) );
  ANDN U5737 ( .B(n4794), .A(n206), .Z(n4792) );
  XNOR U5738 ( .A(a[81]), .B(n4795), .Z(n206) );
  IV U5739 ( .A(n4793), .Z(n4795) );
  XNOR U5740 ( .A(b[81]), .B(n4793), .Z(n4794) );
  XOR U5741 ( .A(n4796), .B(n4797), .Z(n4793) );
  ANDN U5742 ( .B(n4798), .A(n217), .Z(n4796) );
  XNOR U5743 ( .A(a[80]), .B(n4799), .Z(n217) );
  IV U5744 ( .A(n4797), .Z(n4799) );
  XNOR U5745 ( .A(b[80]), .B(n4797), .Z(n4798) );
  XOR U5746 ( .A(n4800), .B(n4801), .Z(n4797) );
  ANDN U5747 ( .B(n4802), .A(n229), .Z(n4800) );
  XNOR U5748 ( .A(a[79]), .B(n4803), .Z(n229) );
  IV U5749 ( .A(n4801), .Z(n4803) );
  XNOR U5750 ( .A(b[79]), .B(n4801), .Z(n4802) );
  XOR U5751 ( .A(n4804), .B(n4805), .Z(n4801) );
  ANDN U5752 ( .B(n4806), .A(n240), .Z(n4804) );
  XNOR U5753 ( .A(a[78]), .B(n4807), .Z(n240) );
  IV U5754 ( .A(n4805), .Z(n4807) );
  XNOR U5755 ( .A(b[78]), .B(n4805), .Z(n4806) );
  XOR U5756 ( .A(n4808), .B(n4809), .Z(n4805) );
  ANDN U5757 ( .B(n4810), .A(n251), .Z(n4808) );
  XNOR U5758 ( .A(a[77]), .B(n4811), .Z(n251) );
  IV U5759 ( .A(n4809), .Z(n4811) );
  XNOR U5760 ( .A(b[77]), .B(n4809), .Z(n4810) );
  XOR U5761 ( .A(n4812), .B(n4813), .Z(n4809) );
  ANDN U5762 ( .B(n4814), .A(n262), .Z(n4812) );
  XNOR U5763 ( .A(a[76]), .B(n4815), .Z(n262) );
  IV U5764 ( .A(n4813), .Z(n4815) );
  XNOR U5765 ( .A(b[76]), .B(n4813), .Z(n4814) );
  XOR U5766 ( .A(n4816), .B(n4817), .Z(n4813) );
  ANDN U5767 ( .B(n4818), .A(n273), .Z(n4816) );
  XNOR U5768 ( .A(a[75]), .B(n4819), .Z(n273) );
  IV U5769 ( .A(n4817), .Z(n4819) );
  XNOR U5770 ( .A(b[75]), .B(n4817), .Z(n4818) );
  XOR U5771 ( .A(n4820), .B(n4821), .Z(n4817) );
  ANDN U5772 ( .B(n4822), .A(n284), .Z(n4820) );
  XNOR U5773 ( .A(a[74]), .B(n4823), .Z(n284) );
  IV U5774 ( .A(n4821), .Z(n4823) );
  XNOR U5775 ( .A(b[74]), .B(n4821), .Z(n4822) );
  XOR U5776 ( .A(n4824), .B(n4825), .Z(n4821) );
  ANDN U5777 ( .B(n4826), .A(n295), .Z(n4824) );
  XNOR U5778 ( .A(a[73]), .B(n4827), .Z(n295) );
  IV U5779 ( .A(n4825), .Z(n4827) );
  XNOR U5780 ( .A(b[73]), .B(n4825), .Z(n4826) );
  XOR U5781 ( .A(n4828), .B(n4829), .Z(n4825) );
  ANDN U5782 ( .B(n4830), .A(n306), .Z(n4828) );
  XNOR U5783 ( .A(a[72]), .B(n4831), .Z(n306) );
  IV U5784 ( .A(n4829), .Z(n4831) );
  XNOR U5785 ( .A(b[72]), .B(n4829), .Z(n4830) );
  XOR U5786 ( .A(n4832), .B(n4833), .Z(n4829) );
  ANDN U5787 ( .B(n4834), .A(n317), .Z(n4832) );
  XNOR U5788 ( .A(a[71]), .B(n4835), .Z(n317) );
  IV U5789 ( .A(n4833), .Z(n4835) );
  XNOR U5790 ( .A(b[71]), .B(n4833), .Z(n4834) );
  XOR U5791 ( .A(n4836), .B(n4837), .Z(n4833) );
  ANDN U5792 ( .B(n4838), .A(n328), .Z(n4836) );
  XNOR U5793 ( .A(a[70]), .B(n4839), .Z(n328) );
  IV U5794 ( .A(n4837), .Z(n4839) );
  XNOR U5795 ( .A(b[70]), .B(n4837), .Z(n4838) );
  XOR U5796 ( .A(n4840), .B(n4841), .Z(n4837) );
  ANDN U5797 ( .B(n4842), .A(n340), .Z(n4840) );
  XNOR U5798 ( .A(a[69]), .B(n4843), .Z(n340) );
  IV U5799 ( .A(n4841), .Z(n4843) );
  XNOR U5800 ( .A(b[69]), .B(n4841), .Z(n4842) );
  XOR U5801 ( .A(n4844), .B(n4845), .Z(n4841) );
  ANDN U5802 ( .B(n4846), .A(n351), .Z(n4844) );
  XNOR U5803 ( .A(a[68]), .B(n4847), .Z(n351) );
  IV U5804 ( .A(n4845), .Z(n4847) );
  XNOR U5805 ( .A(b[68]), .B(n4845), .Z(n4846) );
  XOR U5806 ( .A(n4848), .B(n4849), .Z(n4845) );
  ANDN U5807 ( .B(n4850), .A(n362), .Z(n4848) );
  XNOR U5808 ( .A(a[67]), .B(n4851), .Z(n362) );
  IV U5809 ( .A(n4849), .Z(n4851) );
  XNOR U5810 ( .A(b[67]), .B(n4849), .Z(n4850) );
  XOR U5811 ( .A(n4852), .B(n4853), .Z(n4849) );
  ANDN U5812 ( .B(n4854), .A(n373), .Z(n4852) );
  XNOR U5813 ( .A(a[66]), .B(n4855), .Z(n373) );
  IV U5814 ( .A(n4853), .Z(n4855) );
  XNOR U5815 ( .A(b[66]), .B(n4853), .Z(n4854) );
  XOR U5816 ( .A(n4856), .B(n4857), .Z(n4853) );
  ANDN U5817 ( .B(n4858), .A(n384), .Z(n4856) );
  XNOR U5818 ( .A(a[65]), .B(n4859), .Z(n384) );
  IV U5819 ( .A(n4857), .Z(n4859) );
  XNOR U5820 ( .A(b[65]), .B(n4857), .Z(n4858) );
  XOR U5821 ( .A(n4860), .B(n4861), .Z(n4857) );
  ANDN U5822 ( .B(n4862), .A(n395), .Z(n4860) );
  XNOR U5823 ( .A(a[64]), .B(n4863), .Z(n395) );
  IV U5824 ( .A(n4861), .Z(n4863) );
  XNOR U5825 ( .A(b[64]), .B(n4861), .Z(n4862) );
  XOR U5826 ( .A(n4864), .B(n4865), .Z(n4861) );
  ANDN U5827 ( .B(n4866), .A(n406), .Z(n4864) );
  XNOR U5828 ( .A(a[63]), .B(n4867), .Z(n406) );
  IV U5829 ( .A(n4865), .Z(n4867) );
  XNOR U5830 ( .A(b[63]), .B(n4865), .Z(n4866) );
  XOR U5831 ( .A(n4868), .B(n4869), .Z(n4865) );
  ANDN U5832 ( .B(n4870), .A(n417), .Z(n4868) );
  XNOR U5833 ( .A(a[62]), .B(n4871), .Z(n417) );
  IV U5834 ( .A(n4869), .Z(n4871) );
  XNOR U5835 ( .A(b[62]), .B(n4869), .Z(n4870) );
  XOR U5836 ( .A(n4872), .B(n4873), .Z(n4869) );
  ANDN U5837 ( .B(n4874), .A(n428), .Z(n4872) );
  XNOR U5838 ( .A(a[61]), .B(n4875), .Z(n428) );
  IV U5839 ( .A(n4873), .Z(n4875) );
  XNOR U5840 ( .A(b[61]), .B(n4873), .Z(n4874) );
  XOR U5841 ( .A(n4876), .B(n4877), .Z(n4873) );
  ANDN U5842 ( .B(n4878), .A(n439), .Z(n4876) );
  XNOR U5843 ( .A(a[60]), .B(n4879), .Z(n439) );
  IV U5844 ( .A(n4877), .Z(n4879) );
  XNOR U5845 ( .A(b[60]), .B(n4877), .Z(n4878) );
  XOR U5846 ( .A(n4880), .B(n4881), .Z(n4877) );
  ANDN U5847 ( .B(n4882), .A(n451), .Z(n4880) );
  XNOR U5848 ( .A(a[59]), .B(n4883), .Z(n451) );
  IV U5849 ( .A(n4881), .Z(n4883) );
  XNOR U5850 ( .A(b[59]), .B(n4881), .Z(n4882) );
  XOR U5851 ( .A(n4884), .B(n4885), .Z(n4881) );
  ANDN U5852 ( .B(n4886), .A(n462), .Z(n4884) );
  XNOR U5853 ( .A(a[58]), .B(n4887), .Z(n462) );
  IV U5854 ( .A(n4885), .Z(n4887) );
  XNOR U5855 ( .A(b[58]), .B(n4885), .Z(n4886) );
  XOR U5856 ( .A(n4888), .B(n4889), .Z(n4885) );
  ANDN U5857 ( .B(n4890), .A(n473), .Z(n4888) );
  XNOR U5858 ( .A(a[57]), .B(n4891), .Z(n473) );
  IV U5859 ( .A(n4889), .Z(n4891) );
  XNOR U5860 ( .A(b[57]), .B(n4889), .Z(n4890) );
  XOR U5861 ( .A(n4892), .B(n4893), .Z(n4889) );
  ANDN U5862 ( .B(n4894), .A(n484), .Z(n4892) );
  XNOR U5863 ( .A(a[56]), .B(n4895), .Z(n484) );
  IV U5864 ( .A(n4893), .Z(n4895) );
  XNOR U5865 ( .A(b[56]), .B(n4893), .Z(n4894) );
  XOR U5866 ( .A(n4896), .B(n4897), .Z(n4893) );
  ANDN U5867 ( .B(n4898), .A(n495), .Z(n4896) );
  XNOR U5868 ( .A(a[55]), .B(n4899), .Z(n495) );
  IV U5869 ( .A(n4897), .Z(n4899) );
  XNOR U5870 ( .A(b[55]), .B(n4897), .Z(n4898) );
  XOR U5871 ( .A(n4900), .B(n4901), .Z(n4897) );
  ANDN U5872 ( .B(n4902), .A(n506), .Z(n4900) );
  XNOR U5873 ( .A(a[54]), .B(n4903), .Z(n506) );
  IV U5874 ( .A(n4901), .Z(n4903) );
  XNOR U5875 ( .A(b[54]), .B(n4901), .Z(n4902) );
  XOR U5876 ( .A(n4904), .B(n4905), .Z(n4901) );
  ANDN U5877 ( .B(n4906), .A(n517), .Z(n4904) );
  XNOR U5878 ( .A(a[53]), .B(n4907), .Z(n517) );
  IV U5879 ( .A(n4905), .Z(n4907) );
  XNOR U5880 ( .A(b[53]), .B(n4905), .Z(n4906) );
  XOR U5881 ( .A(n4908), .B(n4909), .Z(n4905) );
  ANDN U5882 ( .B(n4910), .A(n528), .Z(n4908) );
  XNOR U5883 ( .A(a[52]), .B(n4911), .Z(n528) );
  IV U5884 ( .A(n4909), .Z(n4911) );
  XNOR U5885 ( .A(b[52]), .B(n4909), .Z(n4910) );
  XOR U5886 ( .A(n4912), .B(n4913), .Z(n4909) );
  ANDN U5887 ( .B(n4914), .A(n539), .Z(n4912) );
  XNOR U5888 ( .A(a[51]), .B(n4915), .Z(n539) );
  IV U5889 ( .A(n4913), .Z(n4915) );
  XNOR U5890 ( .A(b[51]), .B(n4913), .Z(n4914) );
  XOR U5891 ( .A(n4916), .B(n4917), .Z(n4913) );
  ANDN U5892 ( .B(n4918), .A(n550), .Z(n4916) );
  XNOR U5893 ( .A(a[50]), .B(n4919), .Z(n550) );
  IV U5894 ( .A(n4917), .Z(n4919) );
  XNOR U5895 ( .A(b[50]), .B(n4917), .Z(n4918) );
  XOR U5896 ( .A(n4920), .B(n4921), .Z(n4917) );
  ANDN U5897 ( .B(n4922), .A(n562), .Z(n4920) );
  XNOR U5898 ( .A(a[49]), .B(n4923), .Z(n562) );
  IV U5899 ( .A(n4921), .Z(n4923) );
  XNOR U5900 ( .A(b[49]), .B(n4921), .Z(n4922) );
  XOR U5901 ( .A(n4924), .B(n4925), .Z(n4921) );
  ANDN U5902 ( .B(n4926), .A(n573), .Z(n4924) );
  XNOR U5903 ( .A(a[48]), .B(n4927), .Z(n573) );
  IV U5904 ( .A(n4925), .Z(n4927) );
  XNOR U5905 ( .A(b[48]), .B(n4925), .Z(n4926) );
  XOR U5906 ( .A(n4928), .B(n4929), .Z(n4925) );
  ANDN U5907 ( .B(n4930), .A(n584), .Z(n4928) );
  XNOR U5908 ( .A(a[47]), .B(n4931), .Z(n584) );
  IV U5909 ( .A(n4929), .Z(n4931) );
  XNOR U5910 ( .A(b[47]), .B(n4929), .Z(n4930) );
  XOR U5911 ( .A(n4932), .B(n4933), .Z(n4929) );
  ANDN U5912 ( .B(n4934), .A(n595), .Z(n4932) );
  XNOR U5913 ( .A(a[46]), .B(n4935), .Z(n595) );
  IV U5914 ( .A(n4933), .Z(n4935) );
  XNOR U5915 ( .A(b[46]), .B(n4933), .Z(n4934) );
  XOR U5916 ( .A(n4936), .B(n4937), .Z(n4933) );
  ANDN U5917 ( .B(n4938), .A(n606), .Z(n4936) );
  XNOR U5918 ( .A(a[45]), .B(n4939), .Z(n606) );
  IV U5919 ( .A(n4937), .Z(n4939) );
  XNOR U5920 ( .A(b[45]), .B(n4937), .Z(n4938) );
  XOR U5921 ( .A(n4940), .B(n4941), .Z(n4937) );
  ANDN U5922 ( .B(n4942), .A(n617), .Z(n4940) );
  XNOR U5923 ( .A(a[44]), .B(n4943), .Z(n617) );
  IV U5924 ( .A(n4941), .Z(n4943) );
  XNOR U5925 ( .A(b[44]), .B(n4941), .Z(n4942) );
  XOR U5926 ( .A(n4944), .B(n4945), .Z(n4941) );
  ANDN U5927 ( .B(n4946), .A(n628), .Z(n4944) );
  XNOR U5928 ( .A(a[43]), .B(n4947), .Z(n628) );
  IV U5929 ( .A(n4945), .Z(n4947) );
  XNOR U5930 ( .A(b[43]), .B(n4945), .Z(n4946) );
  XOR U5931 ( .A(n4948), .B(n4949), .Z(n4945) );
  ANDN U5932 ( .B(n4950), .A(n639), .Z(n4948) );
  XNOR U5933 ( .A(a[42]), .B(n4951), .Z(n639) );
  IV U5934 ( .A(n4949), .Z(n4951) );
  XNOR U5935 ( .A(b[42]), .B(n4949), .Z(n4950) );
  XOR U5936 ( .A(n4952), .B(n4953), .Z(n4949) );
  ANDN U5937 ( .B(n4954), .A(n650), .Z(n4952) );
  XNOR U5938 ( .A(a[41]), .B(n4955), .Z(n650) );
  IV U5939 ( .A(n4953), .Z(n4955) );
  XNOR U5940 ( .A(b[41]), .B(n4953), .Z(n4954) );
  XOR U5941 ( .A(n4956), .B(n4957), .Z(n4953) );
  ANDN U5942 ( .B(n4958), .A(n661), .Z(n4956) );
  XNOR U5943 ( .A(a[40]), .B(n4959), .Z(n661) );
  IV U5944 ( .A(n4957), .Z(n4959) );
  XNOR U5945 ( .A(b[40]), .B(n4957), .Z(n4958) );
  XOR U5946 ( .A(n4960), .B(n4961), .Z(n4957) );
  ANDN U5947 ( .B(n4962), .A(n673), .Z(n4960) );
  XNOR U5948 ( .A(a[39]), .B(n4963), .Z(n673) );
  IV U5949 ( .A(n4961), .Z(n4963) );
  XNOR U5950 ( .A(b[39]), .B(n4961), .Z(n4962) );
  XOR U5951 ( .A(n4964), .B(n4965), .Z(n4961) );
  ANDN U5952 ( .B(n4966), .A(n684), .Z(n4964) );
  XNOR U5953 ( .A(a[38]), .B(n4967), .Z(n684) );
  IV U5954 ( .A(n4965), .Z(n4967) );
  XNOR U5955 ( .A(b[38]), .B(n4965), .Z(n4966) );
  XOR U5956 ( .A(n4968), .B(n4969), .Z(n4965) );
  ANDN U5957 ( .B(n4970), .A(n695), .Z(n4968) );
  XNOR U5958 ( .A(a[37]), .B(n4971), .Z(n695) );
  IV U5959 ( .A(n4969), .Z(n4971) );
  XNOR U5960 ( .A(b[37]), .B(n4969), .Z(n4970) );
  XOR U5961 ( .A(n4972), .B(n4973), .Z(n4969) );
  ANDN U5962 ( .B(n4974), .A(n706), .Z(n4972) );
  XNOR U5963 ( .A(a[36]), .B(n4975), .Z(n706) );
  IV U5964 ( .A(n4973), .Z(n4975) );
  XNOR U5965 ( .A(b[36]), .B(n4973), .Z(n4974) );
  XOR U5966 ( .A(n4976), .B(n4977), .Z(n4973) );
  ANDN U5967 ( .B(n4978), .A(n717), .Z(n4976) );
  XNOR U5968 ( .A(a[35]), .B(n4979), .Z(n717) );
  IV U5969 ( .A(n4977), .Z(n4979) );
  XNOR U5970 ( .A(b[35]), .B(n4977), .Z(n4978) );
  XOR U5971 ( .A(n4980), .B(n4981), .Z(n4977) );
  ANDN U5972 ( .B(n4982), .A(n728), .Z(n4980) );
  XNOR U5973 ( .A(a[34]), .B(n4983), .Z(n728) );
  IV U5974 ( .A(n4981), .Z(n4983) );
  XNOR U5975 ( .A(b[34]), .B(n4981), .Z(n4982) );
  XOR U5976 ( .A(n4984), .B(n4985), .Z(n4981) );
  ANDN U5977 ( .B(n4986), .A(n739), .Z(n4984) );
  XNOR U5978 ( .A(a[33]), .B(n4987), .Z(n739) );
  IV U5979 ( .A(n4985), .Z(n4987) );
  XNOR U5980 ( .A(b[33]), .B(n4985), .Z(n4986) );
  XOR U5981 ( .A(n4988), .B(n4989), .Z(n4985) );
  ANDN U5982 ( .B(n4990), .A(n750), .Z(n4988) );
  XNOR U5983 ( .A(a[32]), .B(n4991), .Z(n750) );
  IV U5984 ( .A(n4989), .Z(n4991) );
  XNOR U5985 ( .A(b[32]), .B(n4989), .Z(n4990) );
  XOR U5986 ( .A(n4992), .B(n4993), .Z(n4989) );
  ANDN U5987 ( .B(n4994), .A(n761), .Z(n4992) );
  XNOR U5988 ( .A(a[31]), .B(n4995), .Z(n761) );
  IV U5989 ( .A(n4993), .Z(n4995) );
  XNOR U5990 ( .A(b[31]), .B(n4993), .Z(n4994) );
  XOR U5991 ( .A(n4996), .B(n4997), .Z(n4993) );
  ANDN U5992 ( .B(n4998), .A(n772), .Z(n4996) );
  XNOR U5993 ( .A(a[30]), .B(n4999), .Z(n772) );
  IV U5994 ( .A(n4997), .Z(n4999) );
  XNOR U5995 ( .A(b[30]), .B(n4997), .Z(n4998) );
  XOR U5996 ( .A(n5000), .B(n5001), .Z(n4997) );
  ANDN U5997 ( .B(n5002), .A(n784), .Z(n5000) );
  XNOR U5998 ( .A(a[29]), .B(n5003), .Z(n784) );
  IV U5999 ( .A(n5001), .Z(n5003) );
  XNOR U6000 ( .A(b[29]), .B(n5001), .Z(n5002) );
  XOR U6001 ( .A(n5004), .B(n5005), .Z(n5001) );
  ANDN U6002 ( .B(n5006), .A(n795), .Z(n5004) );
  XNOR U6003 ( .A(a[28]), .B(n5007), .Z(n795) );
  IV U6004 ( .A(n5005), .Z(n5007) );
  XNOR U6005 ( .A(b[28]), .B(n5005), .Z(n5006) );
  XOR U6006 ( .A(n5008), .B(n5009), .Z(n5005) );
  ANDN U6007 ( .B(n5010), .A(n806), .Z(n5008) );
  XNOR U6008 ( .A(a[27]), .B(n5011), .Z(n806) );
  IV U6009 ( .A(n5009), .Z(n5011) );
  XNOR U6010 ( .A(b[27]), .B(n5009), .Z(n5010) );
  XOR U6011 ( .A(n5012), .B(n5013), .Z(n5009) );
  ANDN U6012 ( .B(n5014), .A(n817), .Z(n5012) );
  XNOR U6013 ( .A(a[26]), .B(n5015), .Z(n817) );
  IV U6014 ( .A(n5013), .Z(n5015) );
  XNOR U6015 ( .A(b[26]), .B(n5013), .Z(n5014) );
  XOR U6016 ( .A(n5016), .B(n5017), .Z(n5013) );
  ANDN U6017 ( .B(n5018), .A(n828), .Z(n5016) );
  XNOR U6018 ( .A(a[25]), .B(n5019), .Z(n828) );
  IV U6019 ( .A(n5017), .Z(n5019) );
  XNOR U6020 ( .A(b[25]), .B(n5017), .Z(n5018) );
  XOR U6021 ( .A(n5020), .B(n5021), .Z(n5017) );
  ANDN U6022 ( .B(n5022), .A(n839), .Z(n5020) );
  XNOR U6023 ( .A(a[24]), .B(n5023), .Z(n839) );
  IV U6024 ( .A(n5021), .Z(n5023) );
  XNOR U6025 ( .A(b[24]), .B(n5021), .Z(n5022) );
  XOR U6026 ( .A(n5024), .B(n5025), .Z(n5021) );
  ANDN U6027 ( .B(n5026), .A(n850), .Z(n5024) );
  XNOR U6028 ( .A(a[23]), .B(n5027), .Z(n850) );
  IV U6029 ( .A(n5025), .Z(n5027) );
  XNOR U6030 ( .A(b[23]), .B(n5025), .Z(n5026) );
  XOR U6031 ( .A(n5028), .B(n5029), .Z(n5025) );
  ANDN U6032 ( .B(n5030), .A(n861), .Z(n5028) );
  XNOR U6033 ( .A(a[22]), .B(n5031), .Z(n861) );
  IV U6034 ( .A(n5029), .Z(n5031) );
  XNOR U6035 ( .A(b[22]), .B(n5029), .Z(n5030) );
  XOR U6036 ( .A(n5032), .B(n5033), .Z(n5029) );
  ANDN U6037 ( .B(n5034), .A(n872), .Z(n5032) );
  XNOR U6038 ( .A(a[21]), .B(n5035), .Z(n872) );
  IV U6039 ( .A(n5033), .Z(n5035) );
  XNOR U6040 ( .A(b[21]), .B(n5033), .Z(n5034) );
  XOR U6041 ( .A(n5036), .B(n5037), .Z(n5033) );
  ANDN U6042 ( .B(n5038), .A(n883), .Z(n5036) );
  XNOR U6043 ( .A(a[20]), .B(n5039), .Z(n883) );
  IV U6044 ( .A(n5037), .Z(n5039) );
  XNOR U6045 ( .A(b[20]), .B(n5037), .Z(n5038) );
  XOR U6046 ( .A(n5040), .B(n5041), .Z(n5037) );
  ANDN U6047 ( .B(n5042), .A(n895), .Z(n5040) );
  XNOR U6048 ( .A(a[19]), .B(n5043), .Z(n895) );
  IV U6049 ( .A(n5041), .Z(n5043) );
  XNOR U6050 ( .A(b[19]), .B(n5041), .Z(n5042) );
  XOR U6051 ( .A(n5044), .B(n5045), .Z(n5041) );
  ANDN U6052 ( .B(n5046), .A(n906), .Z(n5044) );
  XNOR U6053 ( .A(a[18]), .B(n5047), .Z(n906) );
  IV U6054 ( .A(n5045), .Z(n5047) );
  XNOR U6055 ( .A(b[18]), .B(n5045), .Z(n5046) );
  XOR U6056 ( .A(n5048), .B(n5049), .Z(n5045) );
  ANDN U6057 ( .B(n5050), .A(n917), .Z(n5048) );
  XNOR U6058 ( .A(a[17]), .B(n5051), .Z(n917) );
  IV U6059 ( .A(n5049), .Z(n5051) );
  XNOR U6060 ( .A(b[17]), .B(n5049), .Z(n5050) );
  XOR U6061 ( .A(n5052), .B(n5053), .Z(n5049) );
  ANDN U6062 ( .B(n5054), .A(n928), .Z(n5052) );
  XNOR U6063 ( .A(a[16]), .B(n5055), .Z(n928) );
  IV U6064 ( .A(n5053), .Z(n5055) );
  XNOR U6065 ( .A(b[16]), .B(n5053), .Z(n5054) );
  XOR U6066 ( .A(n5056), .B(n5057), .Z(n5053) );
  ANDN U6067 ( .B(n5058), .A(n939), .Z(n5056) );
  XNOR U6068 ( .A(a[15]), .B(n5059), .Z(n939) );
  IV U6069 ( .A(n5057), .Z(n5059) );
  XNOR U6070 ( .A(b[15]), .B(n5057), .Z(n5058) );
  XOR U6071 ( .A(n5060), .B(n5061), .Z(n5057) );
  ANDN U6072 ( .B(n5062), .A(n950), .Z(n5060) );
  XNOR U6073 ( .A(a[14]), .B(n5063), .Z(n950) );
  IV U6074 ( .A(n5061), .Z(n5063) );
  XNOR U6075 ( .A(b[14]), .B(n5061), .Z(n5062) );
  XOR U6076 ( .A(n5064), .B(n5065), .Z(n5061) );
  ANDN U6077 ( .B(n5066), .A(n961), .Z(n5064) );
  XNOR U6078 ( .A(a[13]), .B(n5067), .Z(n961) );
  IV U6079 ( .A(n5065), .Z(n5067) );
  XNOR U6080 ( .A(b[13]), .B(n5065), .Z(n5066) );
  XOR U6081 ( .A(n5068), .B(n5069), .Z(n5065) );
  ANDN U6082 ( .B(n5070), .A(n972), .Z(n5068) );
  XNOR U6083 ( .A(a[12]), .B(n5071), .Z(n972) );
  IV U6084 ( .A(n5069), .Z(n5071) );
  XNOR U6085 ( .A(b[12]), .B(n5069), .Z(n5070) );
  XOR U6086 ( .A(n5072), .B(n5073), .Z(n5069) );
  ANDN U6087 ( .B(n5074), .A(n983), .Z(n5072) );
  XNOR U6088 ( .A(a[11]), .B(n5075), .Z(n983) );
  IV U6089 ( .A(n5073), .Z(n5075) );
  XNOR U6090 ( .A(b[11]), .B(n5073), .Z(n5074) );
  XOR U6091 ( .A(n5076), .B(n5077), .Z(n5073) );
  ANDN U6092 ( .B(n5078), .A(n994), .Z(n5076) );
  XNOR U6093 ( .A(a[10]), .B(n5079), .Z(n994) );
  IV U6094 ( .A(n5077), .Z(n5079) );
  XNOR U6095 ( .A(b[10]), .B(n5077), .Z(n5078) );
  XOR U6096 ( .A(n5080), .B(n5081), .Z(n5077) );
  ANDN U6097 ( .B(n5082), .A(n6), .Z(n5080) );
  XNOR U6098 ( .A(a[9]), .B(n5083), .Z(n6) );
  IV U6099 ( .A(n5081), .Z(n5083) );
  XNOR U6100 ( .A(b[9]), .B(n5081), .Z(n5082) );
  XOR U6101 ( .A(n5084), .B(n5085), .Z(n5081) );
  ANDN U6102 ( .B(n5086), .A(n117), .Z(n5084) );
  XNOR U6103 ( .A(a[8]), .B(n5087), .Z(n117) );
  IV U6104 ( .A(n5085), .Z(n5087) );
  XNOR U6105 ( .A(b[8]), .B(n5085), .Z(n5086) );
  XOR U6106 ( .A(n5088), .B(n5089), .Z(n5085) );
  ANDN U6107 ( .B(n5090), .A(n228), .Z(n5088) );
  XNOR U6108 ( .A(a[7]), .B(n5091), .Z(n228) );
  IV U6109 ( .A(n5089), .Z(n5091) );
  XNOR U6110 ( .A(b[7]), .B(n5089), .Z(n5090) );
  XOR U6111 ( .A(n5092), .B(n5093), .Z(n5089) );
  ANDN U6112 ( .B(n5094), .A(n339), .Z(n5092) );
  XNOR U6113 ( .A(a[6]), .B(n5095), .Z(n339) );
  IV U6114 ( .A(n5093), .Z(n5095) );
  XNOR U6115 ( .A(b[6]), .B(n5093), .Z(n5094) );
  XOR U6116 ( .A(n5096), .B(n5097), .Z(n5093) );
  ANDN U6117 ( .B(n5098), .A(n450), .Z(n5096) );
  XNOR U6118 ( .A(a[5]), .B(n5099), .Z(n450) );
  IV U6119 ( .A(n5097), .Z(n5099) );
  XNOR U6120 ( .A(b[5]), .B(n5097), .Z(n5098) );
  XOR U6121 ( .A(n5100), .B(n5101), .Z(n5097) );
  ANDN U6122 ( .B(n5102), .A(n561), .Z(n5100) );
  XNOR U6123 ( .A(a[4]), .B(n5103), .Z(n561) );
  IV U6124 ( .A(n5101), .Z(n5103) );
  XNOR U6125 ( .A(b[4]), .B(n5101), .Z(n5102) );
  XOR U6126 ( .A(n5104), .B(n5105), .Z(n5101) );
  ANDN U6127 ( .B(n5106), .A(n672), .Z(n5104) );
  XNOR U6128 ( .A(a[3]), .B(n5107), .Z(n672) );
  IV U6129 ( .A(n5105), .Z(n5107) );
  XNOR U6130 ( .A(b[3]), .B(n5105), .Z(n5106) );
  XOR U6131 ( .A(n5108), .B(n5109), .Z(n5105) );
  ANDN U6132 ( .B(n5110), .A(n783), .Z(n5108) );
  XNOR U6133 ( .A(a[2]), .B(n5111), .Z(n783) );
  IV U6134 ( .A(n5109), .Z(n5111) );
  XNOR U6135 ( .A(b[2]), .B(n5109), .Z(n5110) );
  XOR U6136 ( .A(n5112), .B(n5113), .Z(n5109) );
  ANDN U6137 ( .B(n5114), .A(n894), .Z(n5112) );
  XNOR U6138 ( .A(a[1]), .B(n5115), .Z(n894) );
  IV U6139 ( .A(n5113), .Z(n5115) );
  XNOR U6140 ( .A(b[1]), .B(n5113), .Z(n5114) );
  XOR U6141 ( .A(carry_on), .B(n5116), .Z(n5113) );
  NANDN U6142 ( .A(n5117), .B(n5118), .Z(n5116) );
  XOR U6143 ( .A(carry_on), .B(b[0]), .Z(n5118) );
  XNOR U6144 ( .A(b[0]), .B(n5117), .Z(c[0]) );
  XNOR U6145 ( .A(a[0]), .B(carry_on), .Z(n5117) );
endmodule

