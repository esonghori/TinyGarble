
module SubBytes_2 ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986;

  XNOR U2962 ( .A(n328), .B(n339), .Z(n341) );
  XNOR U2963 ( .A(n170), .B(n162), .Z(n143) );
  XOR U2964 ( .A(n493), .B(n494), .Z(n646) );
  IV U2965 ( .A(x[1]), .Z(n1447) );
  XOR U2966 ( .A(x[0]), .B(x[6]), .Z(n2) );
  XOR U2967 ( .A(x[5]), .B(n2), .Z(n1446) );
  IV U2968 ( .A(n1446), .Z(n3) );
  AND U2969 ( .A(n1447), .B(n3), .Z(n10) );
  XNOR U2970 ( .A(x[3]), .B(n1447), .Z(n6) );
  XNOR U2971 ( .A(x[2]), .B(n6), .Z(n1) );
  XNOR U2972 ( .A(n2), .B(n1), .Z(n66) );
  IV U2973 ( .A(n66), .Z(n12) );
  XNOR U2974 ( .A(n12), .B(n1446), .Z(n65) );
  IV U2975 ( .A(x[7]), .Z(n4) );
  XNOR U2976 ( .A(x[1]), .B(n4), .Z(n1085) );
  NAND U2977 ( .A(n65), .B(n1085), .Z(n15) );
  XNOR U2978 ( .A(n4), .B(n3), .Z(n11) );
  IV U2979 ( .A(n11), .Z(n1083) );
  XOR U2980 ( .A(n66), .B(n1083), .Z(n31) );
  XNOR U2981 ( .A(n15), .B(n31), .Z(n8) );
  XOR U2982 ( .A(x[0]), .B(n12), .Z(n41) );
  XOR U2983 ( .A(x[4]), .B(n4), .Z(n5) );
  IV U2984 ( .A(n5), .Z(n790) );
  NANDN U2985 ( .A(n41), .B(n790), .Z(n14) );
  XNOR U2986 ( .A(n6), .B(n5), .Z(n59) );
  XNOR U2987 ( .A(n65), .B(n59), .Z(n57) );
  XOR U2988 ( .A(x[2]), .B(x[4]), .Z(n792) );
  NANDN U2989 ( .A(n57), .B(n792), .Z(n7) );
  XOR U2990 ( .A(n14), .B(n7), .Z(n33) );
  XNOR U2991 ( .A(n8), .B(n33), .Z(n9) );
  XOR U2992 ( .A(n10), .B(n9), .Z(n46) );
  IV U2993 ( .A(n46), .Z(n52) );
  AND U2994 ( .A(n12), .B(n11), .Z(n17) );
  XOR U2995 ( .A(x[0]), .B(n59), .Z(n60) );
  XNOR U2996 ( .A(n1446), .B(n60), .Z(n62) );
  XOR U2997 ( .A(x[2]), .B(x[7]), .Z(n807) );
  NANDN U2998 ( .A(n62), .B(n807), .Z(n13) );
  XNOR U2999 ( .A(n14), .B(n13), .Z(n22) );
  XNOR U3000 ( .A(n15), .B(n22), .Z(n16) );
  XOR U3001 ( .A(n17), .B(n16), .Z(n42) );
  XNOR U3002 ( .A(x[4]), .B(n1446), .Z(n800) );
  ANDN U3003 ( .B(x[0]), .A(n800), .Z(n24) );
  XOR U3004 ( .A(x[2]), .B(x[1]), .Z(n18) );
  XOR U3005 ( .A(n1083), .B(n18), .Z(n789) );
  XOR U3006 ( .A(n790), .B(n18), .Z(n795) );
  NAND U3007 ( .A(n59), .B(n795), .Z(n26) );
  XNOR U3008 ( .A(n789), .B(n26), .Z(n20) );
  XNOR U3009 ( .A(x[1]), .B(n60), .Z(n19) );
  XNOR U3010 ( .A(n20), .B(n19), .Z(n21) );
  XOR U3011 ( .A(n22), .B(n21), .Z(n23) );
  XOR U3012 ( .A(n24), .B(n23), .Z(n44) );
  NAND U3013 ( .A(n42), .B(n44), .Z(n25) );
  NAND U3014 ( .A(n52), .B(n25), .Z(n36) );
  IV U3015 ( .A(n42), .Z(n43) );
  IV U3016 ( .A(n44), .Z(n50) );
  XOR U3017 ( .A(n26), .B(n800), .Z(n29) );
  AND U3018 ( .A(n789), .B(n60), .Z(n27) );
  XNOR U3019 ( .A(x[0]), .B(n27), .Z(n28) );
  XNOR U3020 ( .A(n29), .B(n28), .Z(n30) );
  XNOR U3021 ( .A(n31), .B(n30), .Z(n32) );
  XNOR U3022 ( .A(n33), .B(n32), .Z(n54) );
  IV U3023 ( .A(n54), .Z(n49) );
  XOR U3024 ( .A(n50), .B(n49), .Z(n34) );
  NAND U3025 ( .A(n43), .B(n34), .Z(n35) );
  AND U3026 ( .A(n36), .B(n35), .Z(n1454) );
  NAND U3027 ( .A(n50), .B(n43), .Z(n37) );
  NAND U3028 ( .A(n49), .B(n37), .Z(n40) );
  XOR U3029 ( .A(n43), .B(n46), .Z(n38) );
  NAND U3030 ( .A(n44), .B(n38), .Z(n39) );
  AND U3031 ( .A(n40), .B(n39), .Z(n1084) );
  XNOR U3032 ( .A(n1454), .B(n1084), .Z(n791) );
  OR U3033 ( .A(n791), .B(n41), .Z(n64) );
  NAND U3034 ( .A(n52), .B(n42), .Z(n48) );
  AND U3035 ( .A(n44), .B(n43), .Z(n51) );
  XNOR U3036 ( .A(n49), .B(n51), .Z(n45) );
  NAND U3037 ( .A(n46), .B(n45), .Z(n47) );
  AND U3038 ( .A(n48), .B(n47), .Z(n788) );
  NAND U3039 ( .A(n50), .B(n49), .Z(n56) );
  XNOR U3040 ( .A(n52), .B(n51), .Z(n53) );
  NAND U3041 ( .A(n54), .B(n53), .Z(n55) );
  NAND U3042 ( .A(n56), .B(n55), .Z(n1448) );
  XNOR U3043 ( .A(n788), .B(n1448), .Z(n806) );
  XOR U3044 ( .A(n806), .B(n791), .Z(n793) );
  OR U3045 ( .A(n793), .B(n57), .Z(n58) );
  XNOR U3046 ( .A(n64), .B(n58), .Z(n810) );
  XOR U3047 ( .A(n788), .B(n1454), .Z(n796) );
  NANDN U3048 ( .A(n796), .B(n59), .Z(n1456) );
  NANDN U3049 ( .A(n788), .B(n60), .Z(n61) );
  XNOR U3050 ( .A(n1456), .B(n61), .Z(n953) );
  XOR U3051 ( .A(n810), .B(n953), .Z(n799) );
  NANDN U3052 ( .A(n62), .B(n806), .Z(n63) );
  XNOR U3053 ( .A(n64), .B(n63), .Z(n1730) );
  XNOR U3054 ( .A(n1448), .B(n1084), .Z(n1086) );
  NANDN U3055 ( .A(n1086), .B(n65), .Z(n802) );
  NAND U3056 ( .A(n66), .B(n1084), .Z(n67) );
  XNOR U3057 ( .A(n802), .B(n67), .Z(n1453) );
  XOR U3058 ( .A(n1730), .B(n1453), .Z(n1309) );
  XNOR U3059 ( .A(n799), .B(n1309), .Z(z[0]) );
  XOR U3060 ( .A(x[96]), .B(x[102]), .Z(n68) );
  XOR U3061 ( .A(x[101]), .B(n68), .Z(n135) );
  XOR U3062 ( .A(x[100]), .B(n135), .Z(n171) );
  AND U3063 ( .A(x[96]), .B(n171), .Z(n78) );
  XOR U3064 ( .A(x[97]), .B(x[99]), .Z(n71) );
  XNOR U3065 ( .A(n68), .B(x[98]), .Z(n69) );
  XOR U3066 ( .A(n71), .B(n69), .Z(n129) );
  XOR U3067 ( .A(x[96]), .B(n129), .Z(n128) );
  XNOR U3068 ( .A(x[103]), .B(x[100]), .Z(n70) );
  IV U3069 ( .A(n70), .Z(n142) );
  NANDN U3070 ( .A(n128), .B(n142), .Z(n80) );
  IV U3071 ( .A(n135), .Z(n91) );
  XNOR U3072 ( .A(n71), .B(n70), .Z(n123) );
  XOR U3073 ( .A(x[96]), .B(n123), .Z(n124) );
  XOR U3074 ( .A(n91), .B(n124), .Z(n126) );
  XOR U3075 ( .A(x[98]), .B(x[103]), .Z(n164) );
  NANDN U3076 ( .A(n126), .B(n164), .Z(n72) );
  XNOR U3077 ( .A(n80), .B(n72), .Z(n87) );
  XNOR U3078 ( .A(n135), .B(x[103]), .Z(n161) );
  XOR U3079 ( .A(x[97]), .B(x[98]), .Z(n73) );
  XNOR U3080 ( .A(n161), .B(n73), .Z(n151) );
  XOR U3081 ( .A(n142), .B(n73), .Z(n152) );
  NAND U3082 ( .A(n123), .B(n152), .Z(n81) );
  XNOR U3083 ( .A(n151), .B(n81), .Z(n75) );
  XNOR U3084 ( .A(x[97]), .B(n124), .Z(n74) );
  XNOR U3085 ( .A(n75), .B(n74), .Z(n76) );
  XOR U3086 ( .A(n87), .B(n76), .Z(n77) );
  XOR U3087 ( .A(n78), .B(n77), .Z(n115) );
  IV U3088 ( .A(n115), .Z(n108) );
  XNOR U3089 ( .A(n129), .B(n135), .Z(n105) );
  XNOR U3090 ( .A(n105), .B(n123), .Z(n158) );
  XNOR U3091 ( .A(x[98]), .B(x[100]), .Z(n144) );
  OR U3092 ( .A(n158), .B(n144), .Z(n79) );
  XOR U3093 ( .A(n80), .B(n79), .Z(n94) );
  XNOR U3094 ( .A(n129), .B(n161), .Z(n92) );
  XNOR U3095 ( .A(n81), .B(n171), .Z(n84) );
  AND U3096 ( .A(n151), .B(n124), .Z(n82) );
  XNOR U3097 ( .A(x[96]), .B(n82), .Z(n83) );
  XNOR U3098 ( .A(n84), .B(n83), .Z(n85) );
  XOR U3099 ( .A(n92), .B(n85), .Z(n86) );
  XOR U3100 ( .A(n94), .B(n86), .Z(n118) );
  AND U3101 ( .A(n129), .B(n161), .Z(n89) );
  IV U3102 ( .A(x[97]), .Z(n136) );
  XNOR U3103 ( .A(n136), .B(x[103]), .Z(n133) );
  NAND U3104 ( .A(n105), .B(n133), .Z(n93) );
  XNOR U3105 ( .A(n93), .B(n87), .Z(n88) );
  XOR U3106 ( .A(n89), .B(n88), .Z(n107) );
  NAND U3107 ( .A(n118), .B(n107), .Z(n90) );
  NAND U3108 ( .A(n108), .B(n90), .Z(n99) );
  IV U3109 ( .A(n118), .Z(n102) );
  NAND U3110 ( .A(n91), .B(n136), .Z(n97) );
  XOR U3111 ( .A(n93), .B(n92), .Z(n95) );
  XNOR U3112 ( .A(n95), .B(n94), .Z(n96) );
  XOR U3113 ( .A(n97), .B(n96), .Z(n114) );
  IV U3114 ( .A(n107), .Z(n116) );
  XOR U3115 ( .A(n114), .B(n116), .Z(n111) );
  NAND U3116 ( .A(n102), .B(n111), .Z(n98) );
  AND U3117 ( .A(n99), .B(n98), .Z(n127) );
  NAND U3118 ( .A(n118), .B(n108), .Z(n104) );
  AND U3119 ( .A(n115), .B(n116), .Z(n100) );
  XNOR U3120 ( .A(n114), .B(n100), .Z(n101) );
  NAND U3121 ( .A(n102), .B(n101), .Z(n103) );
  AND U3122 ( .A(n104), .B(n103), .Z(n138) );
  XNOR U3123 ( .A(n127), .B(n138), .Z(n134) );
  NANDN U3124 ( .A(n134), .B(n105), .Z(n131) );
  NANDN U3125 ( .A(n138), .B(n135), .Z(n106) );
  XNOR U3126 ( .A(n131), .B(n106), .Z(n173) );
  IV U3127 ( .A(n114), .Z(n120) );
  NAND U3128 ( .A(n120), .B(n107), .Z(n113) );
  AND U3129 ( .A(n120), .B(n118), .Z(n109) );
  XNOR U3130 ( .A(n109), .B(n108), .Z(n110) );
  NAND U3131 ( .A(n111), .B(n110), .Z(n112) );
  NAND U3132 ( .A(n113), .B(n112), .Z(n170) );
  NAND U3133 ( .A(n114), .B(n116), .Z(n122) );
  NAND U3134 ( .A(n116), .B(n115), .Z(n117) );
  XNOR U3135 ( .A(n118), .B(n117), .Z(n119) );
  NAND U3136 ( .A(n120), .B(n119), .Z(n121) );
  NAND U3137 ( .A(n122), .B(n121), .Z(n150) );
  XOR U3138 ( .A(n170), .B(n150), .Z(n153) );
  NANDN U3139 ( .A(n153), .B(n123), .Z(n147) );
  NANDN U3140 ( .A(n150), .B(n124), .Z(n125) );
  XNOR U3141 ( .A(n147), .B(n125), .Z(n160) );
  XNOR U3142 ( .A(n173), .B(n160), .Z(z[98]) );
  XOR U3143 ( .A(n150), .B(n138), .Z(n163) );
  ANDN U3144 ( .B(n163), .A(n126), .Z(n184) );
  IV U3145 ( .A(n127), .Z(n162) );
  OR U3146 ( .A(n143), .B(n128), .Z(n182) );
  NANDN U3147 ( .A(n129), .B(n162), .Z(n130) );
  XNOR U3148 ( .A(n131), .B(n130), .Z(n141) );
  XNOR U3149 ( .A(n182), .B(n141), .Z(n132) );
  XOR U3150 ( .A(n184), .B(n132), .Z(n1982) );
  XNOR U3151 ( .A(n1982), .B(z[98]), .Z(z[100]) );
  NANDN U3152 ( .A(n134), .B(n133), .Z(n167) );
  XNOR U3153 ( .A(n136), .B(n135), .Z(n137) );
  NANDN U3154 ( .A(n138), .B(n137), .Z(n139) );
  XOR U3155 ( .A(n167), .B(n139), .Z(n140) );
  XNOR U3156 ( .A(n141), .B(n140), .Z(n149) );
  NANDN U3157 ( .A(n143), .B(n142), .Z(n166) );
  XNOR U3158 ( .A(n143), .B(n163), .Z(n157) );
  NANDN U3159 ( .A(n144), .B(n157), .Z(n145) );
  XNOR U3160 ( .A(n166), .B(n145), .Z(n154) );
  NAND U3161 ( .A(n170), .B(x[96]), .Z(n146) );
  XNOR U3162 ( .A(n147), .B(n146), .Z(n181) );
  XNOR U3163 ( .A(n154), .B(n181), .Z(n148) );
  XOR U3164 ( .A(n149), .B(n148), .Z(z[101]) );
  ANDN U3165 ( .B(n151), .A(n150), .Z(n156) );
  NANDN U3166 ( .A(n153), .B(n152), .Z(n172) );
  XNOR U3167 ( .A(n172), .B(n154), .Z(n155) );
  XOR U3168 ( .A(n156), .B(n155), .Z(n1983) );
  NANDN U3169 ( .A(n158), .B(n157), .Z(n159) );
  XOR U3170 ( .A(n182), .B(n159), .Z(n176) );
  XOR U3171 ( .A(n176), .B(n160), .Z(n1981) );
  XNOR U3172 ( .A(n1983), .B(n1981), .Z(n180) );
  ANDN U3173 ( .B(n162), .A(n161), .Z(n169) );
  NAND U3174 ( .A(n164), .B(n163), .Z(n165) );
  XNOR U3175 ( .A(n166), .B(n165), .Z(n177) );
  XNOR U3176 ( .A(n177), .B(n167), .Z(n168) );
  XOR U3177 ( .A(n169), .B(n168), .Z(n1986) );
  XNOR U3178 ( .A(n180), .B(n1986), .Z(z[102]) );
  AND U3179 ( .A(n171), .B(n170), .Z(n175) );
  XNOR U3180 ( .A(n173), .B(n172), .Z(n174) );
  XNOR U3181 ( .A(n175), .B(n174), .Z(n179) );
  XOR U3182 ( .A(n177), .B(n176), .Z(n178) );
  XOR U3183 ( .A(n179), .B(n178), .Z(n1984) );
  XNOR U3184 ( .A(n1984), .B(n180), .Z(z[97]) );
  XNOR U3185 ( .A(n182), .B(n181), .Z(n183) );
  XNOR U3186 ( .A(n184), .B(n183), .Z(n185) );
  XOR U3187 ( .A(n185), .B(z[97]), .Z(z[103]) );
  IV U3188 ( .A(x[105]), .Z(n292) );
  XOR U3189 ( .A(x[104]), .B(x[110]), .Z(n187) );
  XOR U3190 ( .A(x[109]), .B(n187), .Z(n291) );
  IV U3191 ( .A(n291), .Z(n188) );
  AND U3192 ( .A(n292), .B(n188), .Z(n195) );
  XNOR U3193 ( .A(x[107]), .B(n292), .Z(n191) );
  XNOR U3194 ( .A(x[106]), .B(n191), .Z(n186) );
  XNOR U3195 ( .A(n187), .B(n186), .Z(n251) );
  IV U3196 ( .A(n251), .Z(n197) );
  XNOR U3197 ( .A(n197), .B(n291), .Z(n250) );
  IV U3198 ( .A(x[111]), .Z(n189) );
  XNOR U3199 ( .A(x[105]), .B(n189), .Z(n282) );
  NAND U3200 ( .A(n250), .B(n282), .Z(n200) );
  XNOR U3201 ( .A(n189), .B(n188), .Z(n196) );
  IV U3202 ( .A(n196), .Z(n280) );
  XOR U3203 ( .A(n251), .B(n280), .Z(n216) );
  XNOR U3204 ( .A(n200), .B(n216), .Z(n193) );
  XOR U3205 ( .A(x[104]), .B(n197), .Z(n226) );
  XOR U3206 ( .A(x[108]), .B(n189), .Z(n190) );
  IV U3207 ( .A(n190), .Z(n255) );
  NANDN U3208 ( .A(n226), .B(n255), .Z(n199) );
  XNOR U3209 ( .A(n191), .B(n190), .Z(n244) );
  XNOR U3210 ( .A(n250), .B(n244), .Z(n242) );
  XOR U3211 ( .A(x[106]), .B(x[108]), .Z(n257) );
  NANDN U3212 ( .A(n242), .B(n257), .Z(n192) );
  XOR U3213 ( .A(n199), .B(n192), .Z(n218) );
  XNOR U3214 ( .A(n193), .B(n218), .Z(n194) );
  XOR U3215 ( .A(n195), .B(n194), .Z(n231) );
  IV U3216 ( .A(n231), .Z(n237) );
  AND U3217 ( .A(n197), .B(n196), .Z(n202) );
  XOR U3218 ( .A(x[104]), .B(n244), .Z(n245) );
  XNOR U3219 ( .A(n291), .B(n245), .Z(n247) );
  XOR U3220 ( .A(x[106]), .B(x[111]), .Z(n272) );
  NANDN U3221 ( .A(n247), .B(n272), .Z(n198) );
  XNOR U3222 ( .A(n199), .B(n198), .Z(n207) );
  XNOR U3223 ( .A(n200), .B(n207), .Z(n201) );
  XOR U3224 ( .A(n202), .B(n201), .Z(n227) );
  XNOR U3225 ( .A(x[108]), .B(n291), .Z(n265) );
  ANDN U3226 ( .B(x[104]), .A(n265), .Z(n209) );
  XOR U3227 ( .A(x[106]), .B(x[105]), .Z(n203) );
  XOR U3228 ( .A(n280), .B(n203), .Z(n254) );
  XOR U3229 ( .A(n255), .B(n203), .Z(n260) );
  NAND U3230 ( .A(n244), .B(n260), .Z(n211) );
  XNOR U3231 ( .A(n254), .B(n211), .Z(n205) );
  XNOR U3232 ( .A(x[105]), .B(n245), .Z(n204) );
  XNOR U3233 ( .A(n205), .B(n204), .Z(n206) );
  XOR U3234 ( .A(n207), .B(n206), .Z(n208) );
  XOR U3235 ( .A(n209), .B(n208), .Z(n229) );
  NAND U3236 ( .A(n227), .B(n229), .Z(n210) );
  NAND U3237 ( .A(n237), .B(n210), .Z(n221) );
  IV U3238 ( .A(n227), .Z(n228) );
  IV U3239 ( .A(n229), .Z(n235) );
  XOR U3240 ( .A(n211), .B(n265), .Z(n214) );
  AND U3241 ( .A(n254), .B(n245), .Z(n212) );
  XNOR U3242 ( .A(x[104]), .B(n212), .Z(n213) );
  XNOR U3243 ( .A(n214), .B(n213), .Z(n215) );
  XNOR U3244 ( .A(n216), .B(n215), .Z(n217) );
  XNOR U3245 ( .A(n218), .B(n217), .Z(n239) );
  IV U3246 ( .A(n239), .Z(n234) );
  XOR U3247 ( .A(n235), .B(n234), .Z(n219) );
  NAND U3248 ( .A(n228), .B(n219), .Z(n220) );
  AND U3249 ( .A(n221), .B(n220), .Z(n299) );
  NAND U3250 ( .A(n235), .B(n228), .Z(n222) );
  NAND U3251 ( .A(n234), .B(n222), .Z(n225) );
  XOR U3252 ( .A(n228), .B(n231), .Z(n223) );
  NAND U3253 ( .A(n229), .B(n223), .Z(n224) );
  AND U3254 ( .A(n225), .B(n224), .Z(n281) );
  XNOR U3255 ( .A(n299), .B(n281), .Z(n256) );
  OR U3256 ( .A(n256), .B(n226), .Z(n249) );
  NAND U3257 ( .A(n237), .B(n227), .Z(n233) );
  AND U3258 ( .A(n229), .B(n228), .Z(n236) );
  XNOR U3259 ( .A(n234), .B(n236), .Z(n230) );
  NAND U3260 ( .A(n231), .B(n230), .Z(n232) );
  AND U3261 ( .A(n233), .B(n232), .Z(n253) );
  NAND U3262 ( .A(n235), .B(n234), .Z(n241) );
  XNOR U3263 ( .A(n237), .B(n236), .Z(n238) );
  NAND U3264 ( .A(n239), .B(n238), .Z(n240) );
  NAND U3265 ( .A(n241), .B(n240), .Z(n293) );
  XNOR U3266 ( .A(n253), .B(n293), .Z(n271) );
  XOR U3267 ( .A(n271), .B(n256), .Z(n258) );
  OR U3268 ( .A(n258), .B(n242), .Z(n243) );
  XNOR U3269 ( .A(n249), .B(n243), .Z(n275) );
  XOR U3270 ( .A(n253), .B(n299), .Z(n261) );
  NANDN U3271 ( .A(n261), .B(n244), .Z(n301) );
  NANDN U3272 ( .A(n253), .B(n245), .Z(n246) );
  XNOR U3273 ( .A(n301), .B(n246), .Z(n279) );
  XOR U3274 ( .A(n275), .B(n279), .Z(n264) );
  NANDN U3275 ( .A(n247), .B(n271), .Z(n248) );
  XNOR U3276 ( .A(n249), .B(n248), .Z(n366) );
  XNOR U3277 ( .A(n293), .B(n281), .Z(n283) );
  NANDN U3278 ( .A(n283), .B(n250), .Z(n267) );
  NAND U3279 ( .A(n251), .B(n281), .Z(n252) );
  XNOR U3280 ( .A(n267), .B(n252), .Z(n298) );
  XOR U3281 ( .A(n366), .B(n298), .Z(n290) );
  XNOR U3282 ( .A(n264), .B(n290), .Z(z[104]) );
  ANDN U3283 ( .B(n254), .A(n253), .Z(n263) );
  NANDN U3284 ( .A(n256), .B(n255), .Z(n274) );
  NANDN U3285 ( .A(n258), .B(n257), .Z(n259) );
  XNOR U3286 ( .A(n274), .B(n259), .Z(n302) );
  NANDN U3287 ( .A(n261), .B(n260), .Z(n268) );
  XNOR U3288 ( .A(n302), .B(n268), .Z(n262) );
  XOR U3289 ( .A(n263), .B(n262), .Z(n288) );
  XOR U3290 ( .A(n288), .B(n264), .Z(n365) );
  ANDN U3291 ( .B(n299), .A(n265), .Z(n270) );
  NAND U3292 ( .A(n291), .B(n293), .Z(n266) );
  XNOR U3293 ( .A(n267), .B(n266), .Z(n278) );
  XNOR U3294 ( .A(n268), .B(n278), .Z(n269) );
  XNOR U3295 ( .A(n270), .B(n269), .Z(n277) );
  NAND U3296 ( .A(n272), .B(n271), .Z(n273) );
  XNOR U3297 ( .A(n274), .B(n273), .Z(n284) );
  XNOR U3298 ( .A(n275), .B(n284), .Z(n276) );
  XOR U3299 ( .A(n277), .B(n276), .Z(n287) );
  XNOR U3300 ( .A(n365), .B(n287), .Z(z[105]) );
  XNOR U3301 ( .A(n279), .B(n278), .Z(z[106]) );
  AND U3302 ( .A(n281), .B(n280), .Z(n286) );
  NANDN U3303 ( .A(n283), .B(n282), .Z(n296) );
  XNOR U3304 ( .A(n284), .B(n296), .Z(n285) );
  XOR U3305 ( .A(n286), .B(n285), .Z(n364) );
  XOR U3306 ( .A(n288), .B(n287), .Z(n289) );
  XOR U3307 ( .A(n364), .B(n289), .Z(z[107]) );
  XOR U3308 ( .A(n290), .B(z[106]), .Z(z[108]) );
  XNOR U3309 ( .A(n292), .B(n291), .Z(n294) );
  NAND U3310 ( .A(n294), .B(n293), .Z(n295) );
  XOR U3311 ( .A(n296), .B(n295), .Z(n297) );
  XNOR U3312 ( .A(n298), .B(n297), .Z(n304) );
  NAND U3313 ( .A(n299), .B(x[104]), .Z(n300) );
  XNOR U3314 ( .A(n301), .B(n300), .Z(n367) );
  XNOR U3315 ( .A(n302), .B(n367), .Z(n303) );
  XOR U3316 ( .A(n304), .B(n303), .Z(z[109]) );
  IV U3317 ( .A(x[15]), .Z(n311) );
  IV U3318 ( .A(x[10]), .Z(n315) );
  XOR U3319 ( .A(x[11]), .B(x[9]), .Z(n307) );
  XOR U3320 ( .A(n315), .B(n307), .Z(n352) );
  IV U3321 ( .A(n352), .Z(n309) );
  XOR U3322 ( .A(x[13]), .B(n309), .Z(n305) );
  IV U3323 ( .A(x[9]), .Z(n655) );
  XNOR U3324 ( .A(n311), .B(n655), .Z(n515) );
  NAND U3325 ( .A(n305), .B(n515), .Z(n306) );
  XNOR U3326 ( .A(n311), .B(n306), .Z(n339) );
  XOR U3327 ( .A(x[12]), .B(n311), .Z(n314) );
  XNOR U3328 ( .A(x[14]), .B(n309), .Z(n497) );
  NOR U3329 ( .A(n314), .B(n497), .Z(n318) );
  IV U3330 ( .A(x[13]), .Z(n353) );
  XOR U3331 ( .A(x[8]), .B(x[14]), .Z(n310) );
  XOR U3332 ( .A(n353), .B(n310), .Z(n325) );
  IV U3333 ( .A(n325), .Z(n656) );
  XOR U3334 ( .A(n314), .B(n307), .Z(n316) );
  XNOR U3335 ( .A(x[8]), .B(n316), .Z(n350) );
  XNOR U3336 ( .A(n656), .B(n350), .Z(n648) );
  XNOR U3337 ( .A(x[15]), .B(n315), .Z(n673) );
  NANDN U3338 ( .A(n648), .B(n673), .Z(n308) );
  XOR U3339 ( .A(n318), .B(n308), .Z(n333) );
  XOR U3340 ( .A(n310), .B(n309), .Z(n313) );
  XNOR U3341 ( .A(n325), .B(n311), .Z(n516) );
  ANDN U3342 ( .B(n313), .A(n516), .Z(n312) );
  XOR U3343 ( .A(n333), .B(n312), .Z(n328) );
  IV U3344 ( .A(n313), .Z(n647) );
  IV U3345 ( .A(n314), .Z(n507) );
  XNOR U3346 ( .A(n655), .B(n315), .Z(n321) );
  XOR U3347 ( .A(n507), .B(n321), .Z(n501) );
  IV U3348 ( .A(n316), .Z(n344) );
  NANDN U3349 ( .A(n501), .B(n344), .Z(n329) );
  XNOR U3350 ( .A(x[12]), .B(x[10]), .Z(n508) );
  XNOR U3351 ( .A(n648), .B(n497), .Z(n498) );
  OR U3352 ( .A(n508), .B(n498), .Z(n317) );
  XOR U3353 ( .A(n318), .B(n317), .Z(n327) );
  XOR U3354 ( .A(n329), .B(n327), .Z(n320) );
  XNOR U3355 ( .A(x[8]), .B(n507), .Z(n319) );
  XNOR U3356 ( .A(n320), .B(n319), .Z(n323) );
  XOR U3357 ( .A(n321), .B(n516), .Z(n505) );
  NAND U3358 ( .A(n350), .B(n505), .Z(n322) );
  XNOR U3359 ( .A(n323), .B(n322), .Z(n324) );
  XOR U3360 ( .A(n647), .B(n324), .Z(n356) );
  IV U3361 ( .A(n356), .Z(n359) );
  NAND U3362 ( .A(n325), .B(n655), .Z(n326) );
  XOR U3363 ( .A(n327), .B(n326), .Z(n338) );
  XNOR U3364 ( .A(n328), .B(n338), .Z(n348) );
  NAND U3365 ( .A(n359), .B(n348), .Z(n337) );
  XOR U3366 ( .A(n656), .B(x[12]), .Z(n502) );
  AND U3367 ( .A(n502), .B(x[8]), .Z(n335) );
  XNOR U3368 ( .A(n505), .B(n329), .Z(n331) );
  XNOR U3369 ( .A(x[9]), .B(n350), .Z(n330) );
  XNOR U3370 ( .A(n331), .B(n330), .Z(n332) );
  XOR U3371 ( .A(n333), .B(n332), .Z(n334) );
  XNOR U3372 ( .A(n335), .B(n334), .Z(n358) );
  NANDN U3373 ( .A(n348), .B(n358), .Z(n336) );
  AND U3374 ( .A(n337), .B(n336), .Z(n342) );
  XNOR U3375 ( .A(n339), .B(n338), .Z(n345) );
  NANDN U3376 ( .A(n345), .B(n356), .Z(n340) );
  XNOR U3377 ( .A(n342), .B(n340), .Z(n354) );
  OR U3378 ( .A(n341), .B(n354), .Z(n495) );
  NANDN U3379 ( .A(n358), .B(n341), .Z(n347) );
  XOR U3380 ( .A(n345), .B(n342), .Z(n343) );
  XNOR U3381 ( .A(n347), .B(n343), .Z(n355) );
  NOR U3382 ( .A(n355), .B(n345), .Z(n349) );
  XOR U3383 ( .A(n495), .B(n349), .Z(n500) );
  NANDN U3384 ( .A(n500), .B(n344), .Z(n664) );
  ANDN U3385 ( .B(n359), .A(n345), .Z(n346) );
  XNOR U3386 ( .A(n347), .B(n346), .Z(n361) );
  OR U3387 ( .A(n361), .B(n348), .Z(n496) );
  XNOR U3388 ( .A(n496), .B(n349), .Z(n504) );
  AND U3389 ( .A(n504), .B(n350), .Z(n351) );
  XOR U3390 ( .A(n664), .B(n351), .Z(n670) );
  XOR U3391 ( .A(n353), .B(n352), .Z(n357) );
  ANDN U3392 ( .B(n358), .A(n354), .Z(n493) );
  NOR U3393 ( .A(n356), .B(n355), .Z(n362) );
  XOR U3394 ( .A(n493), .B(n362), .Z(n514) );
  NAND U3395 ( .A(n357), .B(n514), .Z(n651) );
  XOR U3396 ( .A(n359), .B(n358), .Z(n360) );
  NANDN U3397 ( .A(n361), .B(n360), .Z(n494) );
  XOR U3398 ( .A(n494), .B(n362), .Z(n658) );
  NANDN U3399 ( .A(n658), .B(n656), .Z(n363) );
  XNOR U3400 ( .A(n651), .B(n363), .Z(n519) );
  XOR U3401 ( .A(n670), .B(n519), .Z(n654) );
  IV U3402 ( .A(n654), .Z(z[10]) );
  XNOR U3403 ( .A(n365), .B(n364), .Z(z[110]) );
  XNOR U3404 ( .A(n367), .B(n366), .Z(n368) );
  XNOR U3405 ( .A(z[105]), .B(n368), .Z(z[111]) );
  IV U3406 ( .A(x[113]), .Z(n475) );
  XOR U3407 ( .A(x[112]), .B(x[118]), .Z(n370) );
  XOR U3408 ( .A(x[117]), .B(n370), .Z(n474) );
  IV U3409 ( .A(n474), .Z(n371) );
  AND U3410 ( .A(n475), .B(n371), .Z(n378) );
  XNOR U3411 ( .A(x[115]), .B(n475), .Z(n374) );
  XNOR U3412 ( .A(x[114]), .B(n374), .Z(n369) );
  XNOR U3413 ( .A(n370), .B(n369), .Z(n434) );
  IV U3414 ( .A(n434), .Z(n380) );
  XNOR U3415 ( .A(n380), .B(n474), .Z(n433) );
  IV U3416 ( .A(x[119]), .Z(n372) );
  XNOR U3417 ( .A(x[113]), .B(n372), .Z(n465) );
  NAND U3418 ( .A(n433), .B(n465), .Z(n383) );
  XNOR U3419 ( .A(n372), .B(n371), .Z(n379) );
  IV U3420 ( .A(n379), .Z(n463) );
  XOR U3421 ( .A(n434), .B(n463), .Z(n399) );
  XNOR U3422 ( .A(n383), .B(n399), .Z(n376) );
  XOR U3423 ( .A(x[112]), .B(n380), .Z(n409) );
  XOR U3424 ( .A(x[116]), .B(n372), .Z(n373) );
  IV U3425 ( .A(n373), .Z(n438) );
  NANDN U3426 ( .A(n409), .B(n438), .Z(n382) );
  XNOR U3427 ( .A(n374), .B(n373), .Z(n427) );
  XNOR U3428 ( .A(n433), .B(n427), .Z(n425) );
  XOR U3429 ( .A(x[114]), .B(x[116]), .Z(n440) );
  NANDN U3430 ( .A(n425), .B(n440), .Z(n375) );
  XOR U3431 ( .A(n382), .B(n375), .Z(n401) );
  XNOR U3432 ( .A(n376), .B(n401), .Z(n377) );
  XOR U3433 ( .A(n378), .B(n377), .Z(n414) );
  IV U3434 ( .A(n414), .Z(n420) );
  AND U3435 ( .A(n380), .B(n379), .Z(n385) );
  XOR U3436 ( .A(x[112]), .B(n427), .Z(n428) );
  XNOR U3437 ( .A(n474), .B(n428), .Z(n430) );
  XOR U3438 ( .A(x[114]), .B(x[119]), .Z(n455) );
  NANDN U3439 ( .A(n430), .B(n455), .Z(n381) );
  XNOR U3440 ( .A(n382), .B(n381), .Z(n390) );
  XNOR U3441 ( .A(n383), .B(n390), .Z(n384) );
  XOR U3442 ( .A(n385), .B(n384), .Z(n410) );
  XNOR U3443 ( .A(x[116]), .B(n474), .Z(n448) );
  ANDN U3444 ( .B(x[112]), .A(n448), .Z(n392) );
  XOR U3445 ( .A(x[114]), .B(x[113]), .Z(n386) );
  XOR U3446 ( .A(n463), .B(n386), .Z(n437) );
  XOR U3447 ( .A(n438), .B(n386), .Z(n443) );
  NAND U3448 ( .A(n427), .B(n443), .Z(n394) );
  XNOR U3449 ( .A(n437), .B(n394), .Z(n388) );
  XNOR U3450 ( .A(x[113]), .B(n428), .Z(n387) );
  XNOR U3451 ( .A(n388), .B(n387), .Z(n389) );
  XOR U3452 ( .A(n390), .B(n389), .Z(n391) );
  XOR U3453 ( .A(n392), .B(n391), .Z(n412) );
  NAND U3454 ( .A(n410), .B(n412), .Z(n393) );
  NAND U3455 ( .A(n420), .B(n393), .Z(n404) );
  IV U3456 ( .A(n410), .Z(n411) );
  IV U3457 ( .A(n412), .Z(n418) );
  XOR U3458 ( .A(n394), .B(n448), .Z(n397) );
  AND U3459 ( .A(n437), .B(n428), .Z(n395) );
  XNOR U3460 ( .A(x[112]), .B(n395), .Z(n396) );
  XNOR U3461 ( .A(n397), .B(n396), .Z(n398) );
  XNOR U3462 ( .A(n399), .B(n398), .Z(n400) );
  XNOR U3463 ( .A(n401), .B(n400), .Z(n422) );
  IV U3464 ( .A(n422), .Z(n417) );
  XOR U3465 ( .A(n418), .B(n417), .Z(n402) );
  NAND U3466 ( .A(n411), .B(n402), .Z(n403) );
  AND U3467 ( .A(n404), .B(n403), .Z(n482) );
  NAND U3468 ( .A(n418), .B(n411), .Z(n405) );
  NAND U3469 ( .A(n417), .B(n405), .Z(n408) );
  XOR U3470 ( .A(n411), .B(n414), .Z(n406) );
  NAND U3471 ( .A(n412), .B(n406), .Z(n407) );
  AND U3472 ( .A(n408), .B(n407), .Z(n464) );
  XNOR U3473 ( .A(n482), .B(n464), .Z(n439) );
  OR U3474 ( .A(n439), .B(n409), .Z(n432) );
  NAND U3475 ( .A(n420), .B(n410), .Z(n416) );
  AND U3476 ( .A(n412), .B(n411), .Z(n419) );
  XNOR U3477 ( .A(n417), .B(n419), .Z(n413) );
  NAND U3478 ( .A(n414), .B(n413), .Z(n415) );
  AND U3479 ( .A(n416), .B(n415), .Z(n436) );
  NAND U3480 ( .A(n418), .B(n417), .Z(n424) );
  XNOR U3481 ( .A(n420), .B(n419), .Z(n421) );
  NAND U3482 ( .A(n422), .B(n421), .Z(n423) );
  NAND U3483 ( .A(n424), .B(n423), .Z(n476) );
  XNOR U3484 ( .A(n436), .B(n476), .Z(n454) );
  XOR U3485 ( .A(n454), .B(n439), .Z(n441) );
  OR U3486 ( .A(n441), .B(n425), .Z(n426) );
  XNOR U3487 ( .A(n432), .B(n426), .Z(n458) );
  XOR U3488 ( .A(n436), .B(n482), .Z(n444) );
  NANDN U3489 ( .A(n444), .B(n427), .Z(n484) );
  NANDN U3490 ( .A(n436), .B(n428), .Z(n429) );
  XNOR U3491 ( .A(n484), .B(n429), .Z(n462) );
  XOR U3492 ( .A(n458), .B(n462), .Z(n447) );
  NANDN U3493 ( .A(n430), .B(n454), .Z(n431) );
  XNOR U3494 ( .A(n432), .B(n431), .Z(n490) );
  XNOR U3495 ( .A(n476), .B(n464), .Z(n466) );
  NANDN U3496 ( .A(n466), .B(n433), .Z(n450) );
  NAND U3497 ( .A(n434), .B(n464), .Z(n435) );
  XNOR U3498 ( .A(n450), .B(n435), .Z(n481) );
  XOR U3499 ( .A(n490), .B(n481), .Z(n473) );
  XNOR U3500 ( .A(n447), .B(n473), .Z(z[112]) );
  ANDN U3501 ( .B(n437), .A(n436), .Z(n446) );
  NANDN U3502 ( .A(n439), .B(n438), .Z(n457) );
  NANDN U3503 ( .A(n441), .B(n440), .Z(n442) );
  XNOR U3504 ( .A(n457), .B(n442), .Z(n485) );
  NANDN U3505 ( .A(n444), .B(n443), .Z(n451) );
  XNOR U3506 ( .A(n485), .B(n451), .Z(n445) );
  XOR U3507 ( .A(n446), .B(n445), .Z(n471) );
  XOR U3508 ( .A(n471), .B(n447), .Z(n489) );
  ANDN U3509 ( .B(n482), .A(n448), .Z(n453) );
  NAND U3510 ( .A(n474), .B(n476), .Z(n449) );
  XNOR U3511 ( .A(n450), .B(n449), .Z(n461) );
  XNOR U3512 ( .A(n451), .B(n461), .Z(n452) );
  XNOR U3513 ( .A(n453), .B(n452), .Z(n460) );
  NAND U3514 ( .A(n455), .B(n454), .Z(n456) );
  XNOR U3515 ( .A(n457), .B(n456), .Z(n467) );
  XNOR U3516 ( .A(n458), .B(n467), .Z(n459) );
  XOR U3517 ( .A(n460), .B(n459), .Z(n470) );
  XNOR U3518 ( .A(n489), .B(n470), .Z(z[113]) );
  XNOR U3519 ( .A(n462), .B(n461), .Z(z[114]) );
  AND U3520 ( .A(n464), .B(n463), .Z(n469) );
  NANDN U3521 ( .A(n466), .B(n465), .Z(n479) );
  XNOR U3522 ( .A(n467), .B(n479), .Z(n468) );
  XOR U3523 ( .A(n469), .B(n468), .Z(n488) );
  XOR U3524 ( .A(n471), .B(n470), .Z(n472) );
  XOR U3525 ( .A(n488), .B(n472), .Z(z[115]) );
  XOR U3526 ( .A(n473), .B(z[114]), .Z(z[116]) );
  XNOR U3527 ( .A(n475), .B(n474), .Z(n477) );
  NAND U3528 ( .A(n477), .B(n476), .Z(n478) );
  XOR U3529 ( .A(n479), .B(n478), .Z(n480) );
  XNOR U3530 ( .A(n481), .B(n480), .Z(n487) );
  NAND U3531 ( .A(n482), .B(x[112]), .Z(n483) );
  XNOR U3532 ( .A(n484), .B(n483), .Z(n491) );
  XNOR U3533 ( .A(n485), .B(n491), .Z(n486) );
  XOR U3534 ( .A(n487), .B(n486), .Z(z[117]) );
  XNOR U3535 ( .A(n489), .B(n488), .Z(z[118]) );
  XNOR U3536 ( .A(n491), .B(n490), .Z(n492) );
  XNOR U3537 ( .A(z[113]), .B(n492), .Z(z[119]) );
  XNOR U3538 ( .A(n496), .B(n495), .Z(n662) );
  XOR U3539 ( .A(n646), .B(n662), .Z(n506) );
  NANDN U3540 ( .A(n497), .B(n506), .Z(n650) );
  XNOR U3541 ( .A(n658), .B(n504), .Z(n672) );
  XNOR U3542 ( .A(n506), .B(n672), .Z(n509) );
  OR U3543 ( .A(n498), .B(n509), .Z(n499) );
  XNOR U3544 ( .A(n650), .B(n499), .Z(n671) );
  OR U3545 ( .A(n501), .B(n500), .Z(n511) );
  ANDN U3546 ( .B(n502), .A(n662), .Z(n503) );
  XNOR U3547 ( .A(n511), .B(n503), .Z(n678) );
  AND U3548 ( .A(n505), .B(n504), .Z(n513) );
  NAND U3549 ( .A(n507), .B(n506), .Z(n675) );
  OR U3550 ( .A(n509), .B(n508), .Z(n510) );
  XNOR U3551 ( .A(n675), .B(n510), .Z(n667) );
  XNOR U3552 ( .A(n667), .B(n511), .Z(n512) );
  XOR U3553 ( .A(n513), .B(n512), .Z(n682) );
  NANDN U3554 ( .A(n515), .B(n514), .Z(n660) );
  OR U3555 ( .A(n516), .B(n646), .Z(n517) );
  XOR U3556 ( .A(n660), .B(n517), .Z(n518) );
  XNOR U3557 ( .A(n682), .B(n518), .Z(n677) );
  XNOR U3558 ( .A(n519), .B(n677), .Z(n520) );
  XOR U3559 ( .A(n678), .B(n520), .Z(n521) );
  XOR U3560 ( .A(n671), .B(n521), .Z(z[11]) );
  IV U3561 ( .A(x[121]), .Z(n628) );
  XOR U3562 ( .A(x[120]), .B(x[126]), .Z(n523) );
  XOR U3563 ( .A(x[125]), .B(n523), .Z(n627) );
  IV U3564 ( .A(n627), .Z(n524) );
  AND U3565 ( .A(n628), .B(n524), .Z(n531) );
  XNOR U3566 ( .A(x[123]), .B(n628), .Z(n527) );
  XNOR U3567 ( .A(x[122]), .B(n527), .Z(n522) );
  XNOR U3568 ( .A(n523), .B(n522), .Z(n587) );
  IV U3569 ( .A(n587), .Z(n533) );
  XNOR U3570 ( .A(n533), .B(n627), .Z(n586) );
  IV U3571 ( .A(x[127]), .Z(n525) );
  XNOR U3572 ( .A(x[121]), .B(n525), .Z(n618) );
  NAND U3573 ( .A(n586), .B(n618), .Z(n536) );
  XNOR U3574 ( .A(n525), .B(n524), .Z(n532) );
  IV U3575 ( .A(n532), .Z(n616) );
  XOR U3576 ( .A(n587), .B(n616), .Z(n552) );
  XNOR U3577 ( .A(n536), .B(n552), .Z(n529) );
  XOR U3578 ( .A(x[120]), .B(n533), .Z(n562) );
  XOR U3579 ( .A(x[124]), .B(n525), .Z(n526) );
  IV U3580 ( .A(n526), .Z(n591) );
  NANDN U3581 ( .A(n562), .B(n591), .Z(n535) );
  XNOR U3582 ( .A(n527), .B(n526), .Z(n580) );
  XNOR U3583 ( .A(n586), .B(n580), .Z(n578) );
  XOR U3584 ( .A(x[122]), .B(x[124]), .Z(n593) );
  NANDN U3585 ( .A(n578), .B(n593), .Z(n528) );
  XOR U3586 ( .A(n535), .B(n528), .Z(n554) );
  XNOR U3587 ( .A(n529), .B(n554), .Z(n530) );
  XOR U3588 ( .A(n531), .B(n530), .Z(n567) );
  IV U3589 ( .A(n567), .Z(n573) );
  AND U3590 ( .A(n533), .B(n532), .Z(n538) );
  XOR U3591 ( .A(x[120]), .B(n580), .Z(n581) );
  XNOR U3592 ( .A(n627), .B(n581), .Z(n583) );
  XOR U3593 ( .A(x[122]), .B(x[127]), .Z(n608) );
  NANDN U3594 ( .A(n583), .B(n608), .Z(n534) );
  XNOR U3595 ( .A(n535), .B(n534), .Z(n543) );
  XNOR U3596 ( .A(n536), .B(n543), .Z(n537) );
  XOR U3597 ( .A(n538), .B(n537), .Z(n563) );
  XNOR U3598 ( .A(x[124]), .B(n627), .Z(n601) );
  ANDN U3599 ( .B(x[120]), .A(n601), .Z(n545) );
  XOR U3600 ( .A(x[122]), .B(x[121]), .Z(n539) );
  XOR U3601 ( .A(n616), .B(n539), .Z(n590) );
  XOR U3602 ( .A(n591), .B(n539), .Z(n596) );
  NAND U3603 ( .A(n580), .B(n596), .Z(n547) );
  XNOR U3604 ( .A(n590), .B(n547), .Z(n541) );
  XNOR U3605 ( .A(x[121]), .B(n581), .Z(n540) );
  XNOR U3606 ( .A(n541), .B(n540), .Z(n542) );
  XOR U3607 ( .A(n543), .B(n542), .Z(n544) );
  XOR U3608 ( .A(n545), .B(n544), .Z(n565) );
  NAND U3609 ( .A(n563), .B(n565), .Z(n546) );
  NAND U3610 ( .A(n573), .B(n546), .Z(n557) );
  IV U3611 ( .A(n563), .Z(n564) );
  IV U3612 ( .A(n565), .Z(n571) );
  XOR U3613 ( .A(n547), .B(n601), .Z(n550) );
  AND U3614 ( .A(n590), .B(n581), .Z(n548) );
  XNOR U3615 ( .A(x[120]), .B(n548), .Z(n549) );
  XNOR U3616 ( .A(n550), .B(n549), .Z(n551) );
  XNOR U3617 ( .A(n552), .B(n551), .Z(n553) );
  XNOR U3618 ( .A(n554), .B(n553), .Z(n575) );
  IV U3619 ( .A(n575), .Z(n570) );
  XOR U3620 ( .A(n571), .B(n570), .Z(n555) );
  NAND U3621 ( .A(n564), .B(n555), .Z(n556) );
  AND U3622 ( .A(n557), .B(n556), .Z(n635) );
  NAND U3623 ( .A(n571), .B(n564), .Z(n558) );
  NAND U3624 ( .A(n570), .B(n558), .Z(n561) );
  XOR U3625 ( .A(n564), .B(n567), .Z(n559) );
  NAND U3626 ( .A(n565), .B(n559), .Z(n560) );
  AND U3627 ( .A(n561), .B(n560), .Z(n617) );
  XNOR U3628 ( .A(n635), .B(n617), .Z(n592) );
  OR U3629 ( .A(n592), .B(n562), .Z(n585) );
  NAND U3630 ( .A(n573), .B(n563), .Z(n569) );
  AND U3631 ( .A(n565), .B(n564), .Z(n572) );
  XNOR U3632 ( .A(n570), .B(n572), .Z(n566) );
  NAND U3633 ( .A(n567), .B(n566), .Z(n568) );
  AND U3634 ( .A(n569), .B(n568), .Z(n589) );
  NAND U3635 ( .A(n571), .B(n570), .Z(n577) );
  XNOR U3636 ( .A(n573), .B(n572), .Z(n574) );
  NAND U3637 ( .A(n575), .B(n574), .Z(n576) );
  NAND U3638 ( .A(n577), .B(n576), .Z(n629) );
  XNOR U3639 ( .A(n589), .B(n629), .Z(n607) );
  XOR U3640 ( .A(n607), .B(n592), .Z(n594) );
  OR U3641 ( .A(n594), .B(n578), .Z(n579) );
  XNOR U3642 ( .A(n585), .B(n579), .Z(n611) );
  XOR U3643 ( .A(n589), .B(n635), .Z(n597) );
  NANDN U3644 ( .A(n597), .B(n580), .Z(n637) );
  NANDN U3645 ( .A(n589), .B(n581), .Z(n582) );
  XNOR U3646 ( .A(n637), .B(n582), .Z(n615) );
  XOR U3647 ( .A(n611), .B(n615), .Z(n600) );
  NANDN U3648 ( .A(n583), .B(n607), .Z(n584) );
  XNOR U3649 ( .A(n585), .B(n584), .Z(n643) );
  XNOR U3650 ( .A(n629), .B(n617), .Z(n619) );
  NANDN U3651 ( .A(n619), .B(n586), .Z(n603) );
  NAND U3652 ( .A(n587), .B(n617), .Z(n588) );
  XNOR U3653 ( .A(n603), .B(n588), .Z(n634) );
  XOR U3654 ( .A(n643), .B(n634), .Z(n626) );
  XNOR U3655 ( .A(n600), .B(n626), .Z(z[120]) );
  ANDN U3656 ( .B(n590), .A(n589), .Z(n599) );
  NANDN U3657 ( .A(n592), .B(n591), .Z(n610) );
  NANDN U3658 ( .A(n594), .B(n593), .Z(n595) );
  XNOR U3659 ( .A(n610), .B(n595), .Z(n638) );
  NANDN U3660 ( .A(n597), .B(n596), .Z(n604) );
  XNOR U3661 ( .A(n638), .B(n604), .Z(n598) );
  XOR U3662 ( .A(n599), .B(n598), .Z(n624) );
  XOR U3663 ( .A(n624), .B(n600), .Z(n642) );
  ANDN U3664 ( .B(n635), .A(n601), .Z(n606) );
  NAND U3665 ( .A(n627), .B(n629), .Z(n602) );
  XNOR U3666 ( .A(n603), .B(n602), .Z(n614) );
  XNOR U3667 ( .A(n604), .B(n614), .Z(n605) );
  XNOR U3668 ( .A(n606), .B(n605), .Z(n613) );
  NAND U3669 ( .A(n608), .B(n607), .Z(n609) );
  XNOR U3670 ( .A(n610), .B(n609), .Z(n620) );
  XNOR U3671 ( .A(n611), .B(n620), .Z(n612) );
  XOR U3672 ( .A(n613), .B(n612), .Z(n623) );
  XNOR U3673 ( .A(n642), .B(n623), .Z(z[121]) );
  XNOR U3674 ( .A(n615), .B(n614), .Z(z[122]) );
  AND U3675 ( .A(n617), .B(n616), .Z(n622) );
  NANDN U3676 ( .A(n619), .B(n618), .Z(n632) );
  XNOR U3677 ( .A(n620), .B(n632), .Z(n621) );
  XOR U3678 ( .A(n622), .B(n621), .Z(n641) );
  XOR U3679 ( .A(n624), .B(n623), .Z(n625) );
  XOR U3680 ( .A(n641), .B(n625), .Z(z[123]) );
  XOR U3681 ( .A(n626), .B(z[122]), .Z(z[124]) );
  XNOR U3682 ( .A(n628), .B(n627), .Z(n630) );
  NAND U3683 ( .A(n630), .B(n629), .Z(n631) );
  XOR U3684 ( .A(n632), .B(n631), .Z(n633) );
  XNOR U3685 ( .A(n634), .B(n633), .Z(n640) );
  NAND U3686 ( .A(n635), .B(x[120]), .Z(n636) );
  XNOR U3687 ( .A(n637), .B(n636), .Z(n644) );
  XNOR U3688 ( .A(n638), .B(n644), .Z(n639) );
  XOR U3689 ( .A(n640), .B(n639), .Z(z[125]) );
  XNOR U3690 ( .A(n642), .B(n641), .Z(z[126]) );
  XNOR U3691 ( .A(n644), .B(n643), .Z(n645) );
  XNOR U3692 ( .A(z[121]), .B(n645), .Z(z[127]) );
  NOR U3693 ( .A(n647), .B(n646), .Z(n653) );
  NANDN U3694 ( .A(n648), .B(n672), .Z(n649) );
  XNOR U3695 ( .A(n650), .B(n649), .Z(n663) );
  XNOR U3696 ( .A(n651), .B(n663), .Z(n652) );
  XOR U3697 ( .A(n653), .B(n652), .Z(n1947) );
  XOR U3698 ( .A(n1947), .B(n654), .Z(z[12]) );
  XNOR U3699 ( .A(n656), .B(n655), .Z(n657) );
  NANDN U3700 ( .A(n658), .B(n657), .Z(n659) );
  XOR U3701 ( .A(n660), .B(n659), .Z(n661) );
  XNOR U3702 ( .A(n1947), .B(n661), .Z(n669) );
  ANDN U3703 ( .B(x[8]), .A(n662), .Z(n666) );
  XNOR U3704 ( .A(n664), .B(n663), .Z(n665) );
  XOR U3705 ( .A(n666), .B(n665), .Z(n683) );
  XNOR U3706 ( .A(n667), .B(n683), .Z(n668) );
  XOR U3707 ( .A(n669), .B(n668), .Z(z[13]) );
  XNOR U3708 ( .A(n671), .B(n670), .Z(n1948) );
  NAND U3709 ( .A(n673), .B(n672), .Z(n674) );
  XNOR U3710 ( .A(n675), .B(n674), .Z(n679) );
  XNOR U3711 ( .A(n1948), .B(n679), .Z(n676) );
  XOR U3712 ( .A(n677), .B(n676), .Z(z[14]) );
  XNOR U3713 ( .A(n679), .B(n678), .Z(n680) );
  XNOR U3714 ( .A(z[10]), .B(n680), .Z(n681) );
  XOR U3715 ( .A(n682), .B(n681), .Z(z[9]) );
  XNOR U3716 ( .A(n683), .B(z[9]), .Z(z[15]) );
  IV U3717 ( .A(x[17]), .Z(n815) );
  XOR U3718 ( .A(x[16]), .B(x[22]), .Z(n685) );
  XOR U3719 ( .A(x[21]), .B(n685), .Z(n814) );
  IV U3720 ( .A(n814), .Z(n686) );
  AND U3721 ( .A(n815), .B(n686), .Z(n693) );
  XNOR U3722 ( .A(x[19]), .B(n815), .Z(n689) );
  XNOR U3723 ( .A(x[18]), .B(n689), .Z(n684) );
  XNOR U3724 ( .A(n685), .B(n684), .Z(n749) );
  IV U3725 ( .A(n749), .Z(n695) );
  XNOR U3726 ( .A(n695), .B(n814), .Z(n748) );
  IV U3727 ( .A(x[23]), .Z(n687) );
  XNOR U3728 ( .A(x[17]), .B(n687), .Z(n780) );
  NAND U3729 ( .A(n748), .B(n780), .Z(n698) );
  XNOR U3730 ( .A(n687), .B(n686), .Z(n694) );
  IV U3731 ( .A(n694), .Z(n778) );
  XOR U3732 ( .A(n749), .B(n778), .Z(n714) );
  XNOR U3733 ( .A(n698), .B(n714), .Z(n691) );
  XOR U3734 ( .A(x[16]), .B(n695), .Z(n724) );
  XOR U3735 ( .A(x[20]), .B(n687), .Z(n688) );
  IV U3736 ( .A(n688), .Z(n753) );
  NANDN U3737 ( .A(n724), .B(n753), .Z(n697) );
  XNOR U3738 ( .A(n689), .B(n688), .Z(n742) );
  XNOR U3739 ( .A(n748), .B(n742), .Z(n740) );
  XOR U3740 ( .A(x[18]), .B(x[20]), .Z(n755) );
  NANDN U3741 ( .A(n740), .B(n755), .Z(n690) );
  XOR U3742 ( .A(n697), .B(n690), .Z(n716) );
  XNOR U3743 ( .A(n691), .B(n716), .Z(n692) );
  XOR U3744 ( .A(n693), .B(n692), .Z(n729) );
  IV U3745 ( .A(n729), .Z(n735) );
  AND U3746 ( .A(n695), .B(n694), .Z(n700) );
  XOR U3747 ( .A(x[16]), .B(n742), .Z(n743) );
  XNOR U3748 ( .A(n814), .B(n743), .Z(n745) );
  XOR U3749 ( .A(x[18]), .B(x[23]), .Z(n770) );
  NANDN U3750 ( .A(n745), .B(n770), .Z(n696) );
  XNOR U3751 ( .A(n697), .B(n696), .Z(n705) );
  XNOR U3752 ( .A(n698), .B(n705), .Z(n699) );
  XOR U3753 ( .A(n700), .B(n699), .Z(n725) );
  XNOR U3754 ( .A(x[20]), .B(n814), .Z(n763) );
  ANDN U3755 ( .B(x[16]), .A(n763), .Z(n707) );
  XOR U3756 ( .A(x[18]), .B(x[17]), .Z(n701) );
  XOR U3757 ( .A(n778), .B(n701), .Z(n752) );
  XOR U3758 ( .A(n753), .B(n701), .Z(n758) );
  NAND U3759 ( .A(n742), .B(n758), .Z(n709) );
  XNOR U3760 ( .A(n752), .B(n709), .Z(n703) );
  XNOR U3761 ( .A(x[17]), .B(n743), .Z(n702) );
  XNOR U3762 ( .A(n703), .B(n702), .Z(n704) );
  XOR U3763 ( .A(n705), .B(n704), .Z(n706) );
  XOR U3764 ( .A(n707), .B(n706), .Z(n727) );
  NAND U3765 ( .A(n725), .B(n727), .Z(n708) );
  NAND U3766 ( .A(n735), .B(n708), .Z(n719) );
  IV U3767 ( .A(n725), .Z(n726) );
  IV U3768 ( .A(n727), .Z(n733) );
  XOR U3769 ( .A(n709), .B(n763), .Z(n712) );
  AND U3770 ( .A(n752), .B(n743), .Z(n710) );
  XNOR U3771 ( .A(x[16]), .B(n710), .Z(n711) );
  XNOR U3772 ( .A(n712), .B(n711), .Z(n713) );
  XNOR U3773 ( .A(n714), .B(n713), .Z(n715) );
  XNOR U3774 ( .A(n716), .B(n715), .Z(n737) );
  IV U3775 ( .A(n737), .Z(n732) );
  XOR U3776 ( .A(n733), .B(n732), .Z(n717) );
  NAND U3777 ( .A(n726), .B(n717), .Z(n718) );
  AND U3778 ( .A(n719), .B(n718), .Z(n822) );
  NAND U3779 ( .A(n733), .B(n726), .Z(n720) );
  NAND U3780 ( .A(n732), .B(n720), .Z(n723) );
  XOR U3781 ( .A(n726), .B(n729), .Z(n721) );
  NAND U3782 ( .A(n727), .B(n721), .Z(n722) );
  AND U3783 ( .A(n723), .B(n722), .Z(n779) );
  XNOR U3784 ( .A(n822), .B(n779), .Z(n754) );
  OR U3785 ( .A(n754), .B(n724), .Z(n747) );
  NAND U3786 ( .A(n735), .B(n725), .Z(n731) );
  AND U3787 ( .A(n727), .B(n726), .Z(n734) );
  XNOR U3788 ( .A(n732), .B(n734), .Z(n728) );
  NAND U3789 ( .A(n729), .B(n728), .Z(n730) );
  AND U3790 ( .A(n731), .B(n730), .Z(n751) );
  NAND U3791 ( .A(n733), .B(n732), .Z(n739) );
  XNOR U3792 ( .A(n735), .B(n734), .Z(n736) );
  NAND U3793 ( .A(n737), .B(n736), .Z(n738) );
  NAND U3794 ( .A(n739), .B(n738), .Z(n816) );
  XNOR U3795 ( .A(n751), .B(n816), .Z(n769) );
  XOR U3796 ( .A(n769), .B(n754), .Z(n756) );
  OR U3797 ( .A(n756), .B(n740), .Z(n741) );
  XNOR U3798 ( .A(n747), .B(n741), .Z(n773) );
  XOR U3799 ( .A(n751), .B(n822), .Z(n759) );
  NANDN U3800 ( .A(n759), .B(n742), .Z(n824) );
  NANDN U3801 ( .A(n751), .B(n743), .Z(n744) );
  XNOR U3802 ( .A(n824), .B(n744), .Z(n777) );
  XOR U3803 ( .A(n773), .B(n777), .Z(n762) );
  NANDN U3804 ( .A(n745), .B(n769), .Z(n746) );
  XNOR U3805 ( .A(n747), .B(n746), .Z(n830) );
  XNOR U3806 ( .A(n816), .B(n779), .Z(n781) );
  NANDN U3807 ( .A(n781), .B(n748), .Z(n765) );
  NAND U3808 ( .A(n749), .B(n779), .Z(n750) );
  XNOR U3809 ( .A(n765), .B(n750), .Z(n821) );
  XOR U3810 ( .A(n830), .B(n821), .Z(n813) );
  XNOR U3811 ( .A(n762), .B(n813), .Z(z[16]) );
  ANDN U3812 ( .B(n752), .A(n751), .Z(n761) );
  NANDN U3813 ( .A(n754), .B(n753), .Z(n772) );
  NANDN U3814 ( .A(n756), .B(n755), .Z(n757) );
  XNOR U3815 ( .A(n772), .B(n757), .Z(n825) );
  NANDN U3816 ( .A(n759), .B(n758), .Z(n766) );
  XNOR U3817 ( .A(n825), .B(n766), .Z(n760) );
  XOR U3818 ( .A(n761), .B(n760), .Z(n786) );
  XOR U3819 ( .A(n786), .B(n762), .Z(n829) );
  ANDN U3820 ( .B(n822), .A(n763), .Z(n768) );
  NAND U3821 ( .A(n814), .B(n816), .Z(n764) );
  XNOR U3822 ( .A(n765), .B(n764), .Z(n776) );
  XNOR U3823 ( .A(n766), .B(n776), .Z(n767) );
  XNOR U3824 ( .A(n768), .B(n767), .Z(n775) );
  NAND U3825 ( .A(n770), .B(n769), .Z(n771) );
  XNOR U3826 ( .A(n772), .B(n771), .Z(n782) );
  XNOR U3827 ( .A(n773), .B(n782), .Z(n774) );
  XOR U3828 ( .A(n775), .B(n774), .Z(n785) );
  XNOR U3829 ( .A(n829), .B(n785), .Z(z[17]) );
  XNOR U3830 ( .A(n777), .B(n776), .Z(z[18]) );
  AND U3831 ( .A(n779), .B(n778), .Z(n784) );
  NANDN U3832 ( .A(n781), .B(n780), .Z(n819) );
  XNOR U3833 ( .A(n782), .B(n819), .Z(n783) );
  XOR U3834 ( .A(n784), .B(n783), .Z(n828) );
  XOR U3835 ( .A(n786), .B(n785), .Z(n787) );
  XOR U3836 ( .A(n828), .B(n787), .Z(z[19]) );
  ANDN U3837 ( .B(n789), .A(n788), .Z(n798) );
  NANDN U3838 ( .A(n791), .B(n790), .Z(n809) );
  NANDN U3839 ( .A(n793), .B(n792), .Z(n794) );
  XNOR U3840 ( .A(n809), .B(n794), .Z(n1457) );
  NANDN U3841 ( .A(n796), .B(n795), .Z(n803) );
  XNOR U3842 ( .A(n1457), .B(n803), .Z(n797) );
  XOR U3843 ( .A(n798), .B(n797), .Z(n1091) );
  XOR U3844 ( .A(n1091), .B(n799), .Z(n1600) );
  ANDN U3845 ( .B(n1454), .A(n800), .Z(n805) );
  NAND U3846 ( .A(n1446), .B(n1448), .Z(n801) );
  XNOR U3847 ( .A(n802), .B(n801), .Z(n952) );
  XNOR U3848 ( .A(n803), .B(n952), .Z(n804) );
  XNOR U3849 ( .A(n805), .B(n804), .Z(n812) );
  NAND U3850 ( .A(n807), .B(n806), .Z(n808) );
  XNOR U3851 ( .A(n809), .B(n808), .Z(n1087) );
  XNOR U3852 ( .A(n810), .B(n1087), .Z(n811) );
  XOR U3853 ( .A(n812), .B(n811), .Z(n1090) );
  XNOR U3854 ( .A(n1600), .B(n1090), .Z(z[1]) );
  XOR U3855 ( .A(n813), .B(z[18]), .Z(z[20]) );
  XNOR U3856 ( .A(n815), .B(n814), .Z(n817) );
  NAND U3857 ( .A(n817), .B(n816), .Z(n818) );
  XOR U3858 ( .A(n819), .B(n818), .Z(n820) );
  XNOR U3859 ( .A(n821), .B(n820), .Z(n827) );
  NAND U3860 ( .A(n822), .B(x[16]), .Z(n823) );
  XNOR U3861 ( .A(n824), .B(n823), .Z(n831) );
  XNOR U3862 ( .A(n825), .B(n831), .Z(n826) );
  XOR U3863 ( .A(n827), .B(n826), .Z(z[21]) );
  XNOR U3864 ( .A(n829), .B(n828), .Z(z[22]) );
  XNOR U3865 ( .A(n831), .B(n830), .Z(n832) );
  XNOR U3866 ( .A(z[17]), .B(n832), .Z(z[23]) );
  IV U3867 ( .A(x[25]), .Z(n939) );
  XOR U3868 ( .A(x[24]), .B(x[30]), .Z(n834) );
  XOR U3869 ( .A(x[29]), .B(n834), .Z(n938) );
  IV U3870 ( .A(n938), .Z(n835) );
  AND U3871 ( .A(n939), .B(n835), .Z(n842) );
  XNOR U3872 ( .A(x[27]), .B(n939), .Z(n838) );
  XNOR U3873 ( .A(x[26]), .B(n838), .Z(n833) );
  XNOR U3874 ( .A(n834), .B(n833), .Z(n898) );
  IV U3875 ( .A(n898), .Z(n844) );
  XNOR U3876 ( .A(n844), .B(n938), .Z(n897) );
  IV U3877 ( .A(x[31]), .Z(n836) );
  XNOR U3878 ( .A(x[25]), .B(n836), .Z(n929) );
  NAND U3879 ( .A(n897), .B(n929), .Z(n847) );
  XNOR U3880 ( .A(n836), .B(n835), .Z(n843) );
  IV U3881 ( .A(n843), .Z(n927) );
  XOR U3882 ( .A(n898), .B(n927), .Z(n863) );
  XNOR U3883 ( .A(n847), .B(n863), .Z(n840) );
  XOR U3884 ( .A(x[24]), .B(n844), .Z(n873) );
  XOR U3885 ( .A(x[28]), .B(n836), .Z(n837) );
  IV U3886 ( .A(n837), .Z(n902) );
  NANDN U3887 ( .A(n873), .B(n902), .Z(n846) );
  XNOR U3888 ( .A(n838), .B(n837), .Z(n891) );
  XNOR U3889 ( .A(n897), .B(n891), .Z(n889) );
  XOR U3890 ( .A(x[26]), .B(x[28]), .Z(n904) );
  NANDN U3891 ( .A(n889), .B(n904), .Z(n839) );
  XOR U3892 ( .A(n846), .B(n839), .Z(n865) );
  XNOR U3893 ( .A(n840), .B(n865), .Z(n841) );
  XOR U3894 ( .A(n842), .B(n841), .Z(n878) );
  IV U3895 ( .A(n878), .Z(n884) );
  AND U3896 ( .A(n844), .B(n843), .Z(n849) );
  XOR U3897 ( .A(x[24]), .B(n891), .Z(n892) );
  XNOR U3898 ( .A(n938), .B(n892), .Z(n894) );
  XOR U3899 ( .A(x[26]), .B(x[31]), .Z(n919) );
  NANDN U3900 ( .A(n894), .B(n919), .Z(n845) );
  XNOR U3901 ( .A(n846), .B(n845), .Z(n854) );
  XNOR U3902 ( .A(n847), .B(n854), .Z(n848) );
  XOR U3903 ( .A(n849), .B(n848), .Z(n874) );
  XNOR U3904 ( .A(x[28]), .B(n938), .Z(n912) );
  ANDN U3905 ( .B(x[24]), .A(n912), .Z(n856) );
  XOR U3906 ( .A(x[26]), .B(x[25]), .Z(n850) );
  XOR U3907 ( .A(n927), .B(n850), .Z(n901) );
  XOR U3908 ( .A(n902), .B(n850), .Z(n907) );
  NAND U3909 ( .A(n891), .B(n907), .Z(n858) );
  XNOR U3910 ( .A(n901), .B(n858), .Z(n852) );
  XNOR U3911 ( .A(x[25]), .B(n892), .Z(n851) );
  XNOR U3912 ( .A(n852), .B(n851), .Z(n853) );
  XOR U3913 ( .A(n854), .B(n853), .Z(n855) );
  XOR U3914 ( .A(n856), .B(n855), .Z(n876) );
  NAND U3915 ( .A(n874), .B(n876), .Z(n857) );
  NAND U3916 ( .A(n884), .B(n857), .Z(n868) );
  IV U3917 ( .A(n874), .Z(n875) );
  IV U3918 ( .A(n876), .Z(n882) );
  XOR U3919 ( .A(n858), .B(n912), .Z(n861) );
  AND U3920 ( .A(n901), .B(n892), .Z(n859) );
  XNOR U3921 ( .A(x[24]), .B(n859), .Z(n860) );
  XNOR U3922 ( .A(n861), .B(n860), .Z(n862) );
  XNOR U3923 ( .A(n863), .B(n862), .Z(n864) );
  XNOR U3924 ( .A(n865), .B(n864), .Z(n886) );
  IV U3925 ( .A(n886), .Z(n881) );
  XOR U3926 ( .A(n882), .B(n881), .Z(n866) );
  NAND U3927 ( .A(n875), .B(n866), .Z(n867) );
  AND U3928 ( .A(n868), .B(n867), .Z(n946) );
  NAND U3929 ( .A(n882), .B(n875), .Z(n869) );
  NAND U3930 ( .A(n881), .B(n869), .Z(n872) );
  XOR U3931 ( .A(n875), .B(n878), .Z(n870) );
  NAND U3932 ( .A(n876), .B(n870), .Z(n871) );
  AND U3933 ( .A(n872), .B(n871), .Z(n928) );
  XNOR U3934 ( .A(n946), .B(n928), .Z(n903) );
  OR U3935 ( .A(n903), .B(n873), .Z(n896) );
  NAND U3936 ( .A(n884), .B(n874), .Z(n880) );
  AND U3937 ( .A(n876), .B(n875), .Z(n883) );
  XNOR U3938 ( .A(n881), .B(n883), .Z(n877) );
  NAND U3939 ( .A(n878), .B(n877), .Z(n879) );
  AND U3940 ( .A(n880), .B(n879), .Z(n900) );
  NAND U3941 ( .A(n882), .B(n881), .Z(n888) );
  XNOR U3942 ( .A(n884), .B(n883), .Z(n885) );
  NAND U3943 ( .A(n886), .B(n885), .Z(n887) );
  NAND U3944 ( .A(n888), .B(n887), .Z(n940) );
  XNOR U3945 ( .A(n900), .B(n940), .Z(n918) );
  XOR U3946 ( .A(n918), .B(n903), .Z(n905) );
  OR U3947 ( .A(n905), .B(n889), .Z(n890) );
  XNOR U3948 ( .A(n896), .B(n890), .Z(n922) );
  XOR U3949 ( .A(n900), .B(n946), .Z(n908) );
  NANDN U3950 ( .A(n908), .B(n891), .Z(n948) );
  NANDN U3951 ( .A(n900), .B(n892), .Z(n893) );
  XNOR U3952 ( .A(n948), .B(n893), .Z(n926) );
  XOR U3953 ( .A(n922), .B(n926), .Z(n911) );
  NANDN U3954 ( .A(n894), .B(n918), .Z(n895) );
  XNOR U3955 ( .A(n896), .B(n895), .Z(n956) );
  XNOR U3956 ( .A(n940), .B(n928), .Z(n930) );
  NANDN U3957 ( .A(n930), .B(n897), .Z(n914) );
  NAND U3958 ( .A(n898), .B(n928), .Z(n899) );
  XNOR U3959 ( .A(n914), .B(n899), .Z(n945) );
  XOR U3960 ( .A(n956), .B(n945), .Z(n937) );
  XNOR U3961 ( .A(n911), .B(n937), .Z(z[24]) );
  ANDN U3962 ( .B(n901), .A(n900), .Z(n910) );
  NANDN U3963 ( .A(n903), .B(n902), .Z(n921) );
  NANDN U3964 ( .A(n905), .B(n904), .Z(n906) );
  XNOR U3965 ( .A(n921), .B(n906), .Z(n949) );
  NANDN U3966 ( .A(n908), .B(n907), .Z(n915) );
  XNOR U3967 ( .A(n949), .B(n915), .Z(n909) );
  XOR U3968 ( .A(n910), .B(n909), .Z(n935) );
  XOR U3969 ( .A(n935), .B(n911), .Z(n955) );
  ANDN U3970 ( .B(n946), .A(n912), .Z(n917) );
  NAND U3971 ( .A(n938), .B(n940), .Z(n913) );
  XNOR U3972 ( .A(n914), .B(n913), .Z(n925) );
  XNOR U3973 ( .A(n915), .B(n925), .Z(n916) );
  XNOR U3974 ( .A(n917), .B(n916), .Z(n924) );
  NAND U3975 ( .A(n919), .B(n918), .Z(n920) );
  XNOR U3976 ( .A(n921), .B(n920), .Z(n931) );
  XNOR U3977 ( .A(n922), .B(n931), .Z(n923) );
  XOR U3978 ( .A(n924), .B(n923), .Z(n934) );
  XNOR U3979 ( .A(n955), .B(n934), .Z(z[25]) );
  XNOR U3980 ( .A(n926), .B(n925), .Z(z[26]) );
  AND U3981 ( .A(n928), .B(n927), .Z(n933) );
  NANDN U3982 ( .A(n930), .B(n929), .Z(n943) );
  XNOR U3983 ( .A(n931), .B(n943), .Z(n932) );
  XOR U3984 ( .A(n933), .B(n932), .Z(n954) );
  XOR U3985 ( .A(n935), .B(n934), .Z(n936) );
  XOR U3986 ( .A(n954), .B(n936), .Z(z[27]) );
  XOR U3987 ( .A(n937), .B(z[26]), .Z(z[28]) );
  XNOR U3988 ( .A(n939), .B(n938), .Z(n941) );
  NAND U3989 ( .A(n941), .B(n940), .Z(n942) );
  XOR U3990 ( .A(n943), .B(n942), .Z(n944) );
  XNOR U3991 ( .A(n945), .B(n944), .Z(n951) );
  NAND U3992 ( .A(n946), .B(x[24]), .Z(n947) );
  XNOR U3993 ( .A(n948), .B(n947), .Z(n957) );
  XNOR U3994 ( .A(n949), .B(n957), .Z(n950) );
  XOR U3995 ( .A(n951), .B(n950), .Z(z[29]) );
  XNOR U3996 ( .A(n953), .B(n952), .Z(z[2]) );
  XNOR U3997 ( .A(n955), .B(n954), .Z(z[30]) );
  XNOR U3998 ( .A(n957), .B(n956), .Z(n958) );
  XNOR U3999 ( .A(z[25]), .B(n958), .Z(z[31]) );
  IV U4000 ( .A(x[33]), .Z(n1065) );
  XOR U4001 ( .A(x[32]), .B(x[38]), .Z(n960) );
  XOR U4002 ( .A(x[37]), .B(n960), .Z(n1064) );
  IV U4003 ( .A(n1064), .Z(n961) );
  AND U4004 ( .A(n1065), .B(n961), .Z(n968) );
  XNOR U4005 ( .A(x[35]), .B(n1065), .Z(n964) );
  XNOR U4006 ( .A(x[34]), .B(n964), .Z(n959) );
  XNOR U4007 ( .A(n960), .B(n959), .Z(n1024) );
  IV U4008 ( .A(n1024), .Z(n970) );
  XNOR U4009 ( .A(n970), .B(n1064), .Z(n1023) );
  IV U4010 ( .A(x[39]), .Z(n962) );
  XNOR U4011 ( .A(x[33]), .B(n962), .Z(n1055) );
  NAND U4012 ( .A(n1023), .B(n1055), .Z(n973) );
  XNOR U4013 ( .A(n962), .B(n961), .Z(n969) );
  IV U4014 ( .A(n969), .Z(n1053) );
  XOR U4015 ( .A(n1024), .B(n1053), .Z(n989) );
  XNOR U4016 ( .A(n973), .B(n989), .Z(n966) );
  XOR U4017 ( .A(x[32]), .B(n970), .Z(n999) );
  XOR U4018 ( .A(x[36]), .B(n962), .Z(n963) );
  IV U4019 ( .A(n963), .Z(n1028) );
  NANDN U4020 ( .A(n999), .B(n1028), .Z(n972) );
  XNOR U4021 ( .A(n964), .B(n963), .Z(n1017) );
  XNOR U4022 ( .A(n1023), .B(n1017), .Z(n1015) );
  XOR U4023 ( .A(x[34]), .B(x[36]), .Z(n1030) );
  NANDN U4024 ( .A(n1015), .B(n1030), .Z(n965) );
  XOR U4025 ( .A(n972), .B(n965), .Z(n991) );
  XNOR U4026 ( .A(n966), .B(n991), .Z(n967) );
  XOR U4027 ( .A(n968), .B(n967), .Z(n1004) );
  IV U4028 ( .A(n1004), .Z(n1010) );
  AND U4029 ( .A(n970), .B(n969), .Z(n975) );
  XOR U4030 ( .A(x[32]), .B(n1017), .Z(n1018) );
  XNOR U4031 ( .A(n1064), .B(n1018), .Z(n1020) );
  XOR U4032 ( .A(x[34]), .B(x[39]), .Z(n1045) );
  NANDN U4033 ( .A(n1020), .B(n1045), .Z(n971) );
  XNOR U4034 ( .A(n972), .B(n971), .Z(n980) );
  XNOR U4035 ( .A(n973), .B(n980), .Z(n974) );
  XOR U4036 ( .A(n975), .B(n974), .Z(n1000) );
  XNOR U4037 ( .A(x[36]), .B(n1064), .Z(n1038) );
  ANDN U4038 ( .B(x[32]), .A(n1038), .Z(n982) );
  XOR U4039 ( .A(x[34]), .B(x[33]), .Z(n976) );
  XOR U4040 ( .A(n1053), .B(n976), .Z(n1027) );
  XOR U4041 ( .A(n1028), .B(n976), .Z(n1033) );
  NAND U4042 ( .A(n1017), .B(n1033), .Z(n984) );
  XNOR U4043 ( .A(n1027), .B(n984), .Z(n978) );
  XNOR U4044 ( .A(x[33]), .B(n1018), .Z(n977) );
  XNOR U4045 ( .A(n978), .B(n977), .Z(n979) );
  XOR U4046 ( .A(n980), .B(n979), .Z(n981) );
  XOR U4047 ( .A(n982), .B(n981), .Z(n1002) );
  NAND U4048 ( .A(n1000), .B(n1002), .Z(n983) );
  NAND U4049 ( .A(n1010), .B(n983), .Z(n994) );
  IV U4050 ( .A(n1000), .Z(n1001) );
  IV U4051 ( .A(n1002), .Z(n1008) );
  XOR U4052 ( .A(n984), .B(n1038), .Z(n987) );
  AND U4053 ( .A(n1027), .B(n1018), .Z(n985) );
  XNOR U4054 ( .A(x[32]), .B(n985), .Z(n986) );
  XNOR U4055 ( .A(n987), .B(n986), .Z(n988) );
  XNOR U4056 ( .A(n989), .B(n988), .Z(n990) );
  XNOR U4057 ( .A(n991), .B(n990), .Z(n1012) );
  IV U4058 ( .A(n1012), .Z(n1007) );
  XOR U4059 ( .A(n1008), .B(n1007), .Z(n992) );
  NAND U4060 ( .A(n1001), .B(n992), .Z(n993) );
  AND U4061 ( .A(n994), .B(n993), .Z(n1072) );
  NAND U4062 ( .A(n1008), .B(n1001), .Z(n995) );
  NAND U4063 ( .A(n1007), .B(n995), .Z(n998) );
  XOR U4064 ( .A(n1001), .B(n1004), .Z(n996) );
  NAND U4065 ( .A(n1002), .B(n996), .Z(n997) );
  AND U4066 ( .A(n998), .B(n997), .Z(n1054) );
  XNOR U4067 ( .A(n1072), .B(n1054), .Z(n1029) );
  OR U4068 ( .A(n1029), .B(n999), .Z(n1022) );
  NAND U4069 ( .A(n1010), .B(n1000), .Z(n1006) );
  AND U4070 ( .A(n1002), .B(n1001), .Z(n1009) );
  XNOR U4071 ( .A(n1007), .B(n1009), .Z(n1003) );
  NAND U4072 ( .A(n1004), .B(n1003), .Z(n1005) );
  AND U4073 ( .A(n1006), .B(n1005), .Z(n1026) );
  NAND U4074 ( .A(n1008), .B(n1007), .Z(n1014) );
  XNOR U4075 ( .A(n1010), .B(n1009), .Z(n1011) );
  NAND U4076 ( .A(n1012), .B(n1011), .Z(n1013) );
  NAND U4077 ( .A(n1014), .B(n1013), .Z(n1066) );
  XNOR U4078 ( .A(n1026), .B(n1066), .Z(n1044) );
  XOR U4079 ( .A(n1044), .B(n1029), .Z(n1031) );
  OR U4080 ( .A(n1031), .B(n1015), .Z(n1016) );
  XNOR U4081 ( .A(n1022), .B(n1016), .Z(n1048) );
  XOR U4082 ( .A(n1026), .B(n1072), .Z(n1034) );
  NANDN U4083 ( .A(n1034), .B(n1017), .Z(n1074) );
  NANDN U4084 ( .A(n1026), .B(n1018), .Z(n1019) );
  XNOR U4085 ( .A(n1074), .B(n1019), .Z(n1052) );
  XOR U4086 ( .A(n1048), .B(n1052), .Z(n1037) );
  NANDN U4087 ( .A(n1020), .B(n1044), .Z(n1021) );
  XNOR U4088 ( .A(n1022), .B(n1021), .Z(n1080) );
  XNOR U4089 ( .A(n1066), .B(n1054), .Z(n1056) );
  NANDN U4090 ( .A(n1056), .B(n1023), .Z(n1040) );
  NAND U4091 ( .A(n1024), .B(n1054), .Z(n1025) );
  XNOR U4092 ( .A(n1040), .B(n1025), .Z(n1071) );
  XOR U4093 ( .A(n1080), .B(n1071), .Z(n1063) );
  XNOR U4094 ( .A(n1037), .B(n1063), .Z(z[32]) );
  ANDN U4095 ( .B(n1027), .A(n1026), .Z(n1036) );
  NANDN U4096 ( .A(n1029), .B(n1028), .Z(n1047) );
  NANDN U4097 ( .A(n1031), .B(n1030), .Z(n1032) );
  XNOR U4098 ( .A(n1047), .B(n1032), .Z(n1075) );
  NANDN U4099 ( .A(n1034), .B(n1033), .Z(n1041) );
  XNOR U4100 ( .A(n1075), .B(n1041), .Z(n1035) );
  XOR U4101 ( .A(n1036), .B(n1035), .Z(n1061) );
  XOR U4102 ( .A(n1061), .B(n1037), .Z(n1079) );
  ANDN U4103 ( .B(n1072), .A(n1038), .Z(n1043) );
  NAND U4104 ( .A(n1064), .B(n1066), .Z(n1039) );
  XNOR U4105 ( .A(n1040), .B(n1039), .Z(n1051) );
  XNOR U4106 ( .A(n1041), .B(n1051), .Z(n1042) );
  XNOR U4107 ( .A(n1043), .B(n1042), .Z(n1050) );
  NAND U4108 ( .A(n1045), .B(n1044), .Z(n1046) );
  XNOR U4109 ( .A(n1047), .B(n1046), .Z(n1057) );
  XNOR U4110 ( .A(n1048), .B(n1057), .Z(n1049) );
  XOR U4111 ( .A(n1050), .B(n1049), .Z(n1060) );
  XNOR U4112 ( .A(n1079), .B(n1060), .Z(z[33]) );
  XNOR U4113 ( .A(n1052), .B(n1051), .Z(z[34]) );
  AND U4114 ( .A(n1054), .B(n1053), .Z(n1059) );
  NANDN U4115 ( .A(n1056), .B(n1055), .Z(n1069) );
  XNOR U4116 ( .A(n1057), .B(n1069), .Z(n1058) );
  XOR U4117 ( .A(n1059), .B(n1058), .Z(n1078) );
  XOR U4118 ( .A(n1061), .B(n1060), .Z(n1062) );
  XOR U4119 ( .A(n1078), .B(n1062), .Z(z[35]) );
  XOR U4120 ( .A(n1063), .B(z[34]), .Z(z[36]) );
  XNOR U4121 ( .A(n1065), .B(n1064), .Z(n1067) );
  NAND U4122 ( .A(n1067), .B(n1066), .Z(n1068) );
  XOR U4123 ( .A(n1069), .B(n1068), .Z(n1070) );
  XNOR U4124 ( .A(n1071), .B(n1070), .Z(n1077) );
  NAND U4125 ( .A(n1072), .B(x[32]), .Z(n1073) );
  XNOR U4126 ( .A(n1074), .B(n1073), .Z(n1081) );
  XNOR U4127 ( .A(n1075), .B(n1081), .Z(n1076) );
  XOR U4128 ( .A(n1077), .B(n1076), .Z(z[37]) );
  XNOR U4129 ( .A(n1079), .B(n1078), .Z(z[38]) );
  XNOR U4130 ( .A(n1081), .B(n1080), .Z(n1082) );
  XNOR U4131 ( .A(z[33]), .B(n1082), .Z(z[39]) );
  AND U4132 ( .A(n1084), .B(n1083), .Z(n1089) );
  NANDN U4133 ( .A(n1086), .B(n1085), .Z(n1451) );
  XNOR U4134 ( .A(n1087), .B(n1451), .Z(n1088) );
  XOR U4135 ( .A(n1089), .B(n1088), .Z(n1599) );
  XOR U4136 ( .A(n1091), .B(n1090), .Z(n1092) );
  XOR U4137 ( .A(n1599), .B(n1092), .Z(z[3]) );
  IV U4138 ( .A(x[41]), .Z(n1199) );
  XOR U4139 ( .A(x[40]), .B(x[46]), .Z(n1094) );
  XOR U4140 ( .A(x[45]), .B(n1094), .Z(n1198) );
  IV U4141 ( .A(n1198), .Z(n1095) );
  AND U4142 ( .A(n1199), .B(n1095), .Z(n1102) );
  XNOR U4143 ( .A(x[43]), .B(n1199), .Z(n1098) );
  XNOR U4144 ( .A(x[42]), .B(n1098), .Z(n1093) );
  XNOR U4145 ( .A(n1094), .B(n1093), .Z(n1158) );
  IV U4146 ( .A(n1158), .Z(n1104) );
  XNOR U4147 ( .A(n1104), .B(n1198), .Z(n1157) );
  IV U4148 ( .A(x[47]), .Z(n1096) );
  XNOR U4149 ( .A(x[41]), .B(n1096), .Z(n1189) );
  NAND U4150 ( .A(n1157), .B(n1189), .Z(n1107) );
  XNOR U4151 ( .A(n1096), .B(n1095), .Z(n1103) );
  IV U4152 ( .A(n1103), .Z(n1187) );
  XOR U4153 ( .A(n1158), .B(n1187), .Z(n1123) );
  XNOR U4154 ( .A(n1107), .B(n1123), .Z(n1100) );
  XOR U4155 ( .A(x[40]), .B(n1104), .Z(n1133) );
  XOR U4156 ( .A(x[44]), .B(n1096), .Z(n1097) );
  IV U4157 ( .A(n1097), .Z(n1162) );
  NANDN U4158 ( .A(n1133), .B(n1162), .Z(n1106) );
  XNOR U4159 ( .A(n1098), .B(n1097), .Z(n1151) );
  XNOR U4160 ( .A(n1157), .B(n1151), .Z(n1149) );
  XOR U4161 ( .A(x[42]), .B(x[44]), .Z(n1164) );
  NANDN U4162 ( .A(n1149), .B(n1164), .Z(n1099) );
  XOR U4163 ( .A(n1106), .B(n1099), .Z(n1125) );
  XNOR U4164 ( .A(n1100), .B(n1125), .Z(n1101) );
  XOR U4165 ( .A(n1102), .B(n1101), .Z(n1138) );
  IV U4166 ( .A(n1138), .Z(n1144) );
  AND U4167 ( .A(n1104), .B(n1103), .Z(n1109) );
  XOR U4168 ( .A(x[40]), .B(n1151), .Z(n1152) );
  XNOR U4169 ( .A(n1198), .B(n1152), .Z(n1154) );
  XOR U4170 ( .A(x[42]), .B(x[47]), .Z(n1179) );
  NANDN U4171 ( .A(n1154), .B(n1179), .Z(n1105) );
  XNOR U4172 ( .A(n1106), .B(n1105), .Z(n1114) );
  XNOR U4173 ( .A(n1107), .B(n1114), .Z(n1108) );
  XOR U4174 ( .A(n1109), .B(n1108), .Z(n1134) );
  XNOR U4175 ( .A(x[44]), .B(n1198), .Z(n1172) );
  ANDN U4176 ( .B(x[40]), .A(n1172), .Z(n1116) );
  XOR U4177 ( .A(x[42]), .B(x[41]), .Z(n1110) );
  XOR U4178 ( .A(n1187), .B(n1110), .Z(n1161) );
  XOR U4179 ( .A(n1162), .B(n1110), .Z(n1167) );
  NAND U4180 ( .A(n1151), .B(n1167), .Z(n1118) );
  XNOR U4181 ( .A(n1161), .B(n1118), .Z(n1112) );
  XNOR U4182 ( .A(x[41]), .B(n1152), .Z(n1111) );
  XNOR U4183 ( .A(n1112), .B(n1111), .Z(n1113) );
  XOR U4184 ( .A(n1114), .B(n1113), .Z(n1115) );
  XOR U4185 ( .A(n1116), .B(n1115), .Z(n1136) );
  NAND U4186 ( .A(n1134), .B(n1136), .Z(n1117) );
  NAND U4187 ( .A(n1144), .B(n1117), .Z(n1128) );
  IV U4188 ( .A(n1134), .Z(n1135) );
  IV U4189 ( .A(n1136), .Z(n1142) );
  XOR U4190 ( .A(n1118), .B(n1172), .Z(n1121) );
  AND U4191 ( .A(n1161), .B(n1152), .Z(n1119) );
  XNOR U4192 ( .A(x[40]), .B(n1119), .Z(n1120) );
  XNOR U4193 ( .A(n1121), .B(n1120), .Z(n1122) );
  XNOR U4194 ( .A(n1123), .B(n1122), .Z(n1124) );
  XNOR U4195 ( .A(n1125), .B(n1124), .Z(n1146) );
  IV U4196 ( .A(n1146), .Z(n1141) );
  XOR U4197 ( .A(n1142), .B(n1141), .Z(n1126) );
  NAND U4198 ( .A(n1135), .B(n1126), .Z(n1127) );
  AND U4199 ( .A(n1128), .B(n1127), .Z(n1206) );
  NAND U4200 ( .A(n1142), .B(n1135), .Z(n1129) );
  NAND U4201 ( .A(n1141), .B(n1129), .Z(n1132) );
  XOR U4202 ( .A(n1135), .B(n1138), .Z(n1130) );
  NAND U4203 ( .A(n1136), .B(n1130), .Z(n1131) );
  AND U4204 ( .A(n1132), .B(n1131), .Z(n1188) );
  XNOR U4205 ( .A(n1206), .B(n1188), .Z(n1163) );
  OR U4206 ( .A(n1163), .B(n1133), .Z(n1156) );
  NAND U4207 ( .A(n1144), .B(n1134), .Z(n1140) );
  AND U4208 ( .A(n1136), .B(n1135), .Z(n1143) );
  XNOR U4209 ( .A(n1141), .B(n1143), .Z(n1137) );
  NAND U4210 ( .A(n1138), .B(n1137), .Z(n1139) );
  AND U4211 ( .A(n1140), .B(n1139), .Z(n1160) );
  NAND U4212 ( .A(n1142), .B(n1141), .Z(n1148) );
  XNOR U4213 ( .A(n1144), .B(n1143), .Z(n1145) );
  NAND U4214 ( .A(n1146), .B(n1145), .Z(n1147) );
  NAND U4215 ( .A(n1148), .B(n1147), .Z(n1200) );
  XNOR U4216 ( .A(n1160), .B(n1200), .Z(n1178) );
  XOR U4217 ( .A(n1178), .B(n1163), .Z(n1165) );
  OR U4218 ( .A(n1165), .B(n1149), .Z(n1150) );
  XNOR U4219 ( .A(n1156), .B(n1150), .Z(n1182) );
  XOR U4220 ( .A(n1160), .B(n1206), .Z(n1168) );
  NANDN U4221 ( .A(n1168), .B(n1151), .Z(n1208) );
  NANDN U4222 ( .A(n1160), .B(n1152), .Z(n1153) );
  XNOR U4223 ( .A(n1208), .B(n1153), .Z(n1186) );
  XOR U4224 ( .A(n1182), .B(n1186), .Z(n1171) );
  NANDN U4225 ( .A(n1154), .B(n1178), .Z(n1155) );
  XNOR U4226 ( .A(n1156), .B(n1155), .Z(n1214) );
  XNOR U4227 ( .A(n1200), .B(n1188), .Z(n1190) );
  NANDN U4228 ( .A(n1190), .B(n1157), .Z(n1174) );
  NAND U4229 ( .A(n1158), .B(n1188), .Z(n1159) );
  XNOR U4230 ( .A(n1174), .B(n1159), .Z(n1205) );
  XOR U4231 ( .A(n1214), .B(n1205), .Z(n1197) );
  XNOR U4232 ( .A(n1171), .B(n1197), .Z(z[40]) );
  ANDN U4233 ( .B(n1161), .A(n1160), .Z(n1170) );
  NANDN U4234 ( .A(n1163), .B(n1162), .Z(n1181) );
  NANDN U4235 ( .A(n1165), .B(n1164), .Z(n1166) );
  XNOR U4236 ( .A(n1181), .B(n1166), .Z(n1209) );
  NANDN U4237 ( .A(n1168), .B(n1167), .Z(n1175) );
  XNOR U4238 ( .A(n1209), .B(n1175), .Z(n1169) );
  XOR U4239 ( .A(n1170), .B(n1169), .Z(n1195) );
  XOR U4240 ( .A(n1195), .B(n1171), .Z(n1213) );
  ANDN U4241 ( .B(n1206), .A(n1172), .Z(n1177) );
  NAND U4242 ( .A(n1198), .B(n1200), .Z(n1173) );
  XNOR U4243 ( .A(n1174), .B(n1173), .Z(n1185) );
  XNOR U4244 ( .A(n1175), .B(n1185), .Z(n1176) );
  XNOR U4245 ( .A(n1177), .B(n1176), .Z(n1184) );
  NAND U4246 ( .A(n1179), .B(n1178), .Z(n1180) );
  XNOR U4247 ( .A(n1181), .B(n1180), .Z(n1191) );
  XNOR U4248 ( .A(n1182), .B(n1191), .Z(n1183) );
  XOR U4249 ( .A(n1184), .B(n1183), .Z(n1194) );
  XNOR U4250 ( .A(n1213), .B(n1194), .Z(z[41]) );
  XNOR U4251 ( .A(n1186), .B(n1185), .Z(z[42]) );
  AND U4252 ( .A(n1188), .B(n1187), .Z(n1193) );
  NANDN U4253 ( .A(n1190), .B(n1189), .Z(n1203) );
  XNOR U4254 ( .A(n1191), .B(n1203), .Z(n1192) );
  XOR U4255 ( .A(n1193), .B(n1192), .Z(n1212) );
  XOR U4256 ( .A(n1195), .B(n1194), .Z(n1196) );
  XOR U4257 ( .A(n1212), .B(n1196), .Z(z[43]) );
  XOR U4258 ( .A(n1197), .B(z[42]), .Z(z[44]) );
  XNOR U4259 ( .A(n1199), .B(n1198), .Z(n1201) );
  NAND U4260 ( .A(n1201), .B(n1200), .Z(n1202) );
  XOR U4261 ( .A(n1203), .B(n1202), .Z(n1204) );
  XNOR U4262 ( .A(n1205), .B(n1204), .Z(n1211) );
  NAND U4263 ( .A(n1206), .B(x[40]), .Z(n1207) );
  XNOR U4264 ( .A(n1208), .B(n1207), .Z(n1215) );
  XNOR U4265 ( .A(n1209), .B(n1215), .Z(n1210) );
  XOR U4266 ( .A(n1211), .B(n1210), .Z(z[45]) );
  XNOR U4267 ( .A(n1213), .B(n1212), .Z(z[46]) );
  XNOR U4268 ( .A(n1215), .B(n1214), .Z(n1216) );
  XNOR U4269 ( .A(z[41]), .B(n1216), .Z(z[47]) );
  IV U4270 ( .A(x[49]), .Z(n1324) );
  XOR U4271 ( .A(x[48]), .B(x[54]), .Z(n1218) );
  XOR U4272 ( .A(x[53]), .B(n1218), .Z(n1323) );
  IV U4273 ( .A(n1323), .Z(n1219) );
  AND U4274 ( .A(n1324), .B(n1219), .Z(n1226) );
  XNOR U4275 ( .A(x[51]), .B(n1324), .Z(n1222) );
  XNOR U4276 ( .A(x[50]), .B(n1222), .Z(n1217) );
  XNOR U4277 ( .A(n1218), .B(n1217), .Z(n1282) );
  IV U4278 ( .A(n1282), .Z(n1228) );
  XNOR U4279 ( .A(n1228), .B(n1323), .Z(n1281) );
  IV U4280 ( .A(x[55]), .Z(n1220) );
  XNOR U4281 ( .A(x[49]), .B(n1220), .Z(n1314) );
  NAND U4282 ( .A(n1281), .B(n1314), .Z(n1231) );
  XNOR U4283 ( .A(n1220), .B(n1219), .Z(n1227) );
  IV U4284 ( .A(n1227), .Z(n1312) );
  XOR U4285 ( .A(n1282), .B(n1312), .Z(n1247) );
  XNOR U4286 ( .A(n1231), .B(n1247), .Z(n1224) );
  XOR U4287 ( .A(x[48]), .B(n1228), .Z(n1257) );
  XOR U4288 ( .A(x[52]), .B(n1220), .Z(n1221) );
  IV U4289 ( .A(n1221), .Z(n1286) );
  NANDN U4290 ( .A(n1257), .B(n1286), .Z(n1230) );
  XNOR U4291 ( .A(n1222), .B(n1221), .Z(n1275) );
  XNOR U4292 ( .A(n1281), .B(n1275), .Z(n1273) );
  XOR U4293 ( .A(x[50]), .B(x[52]), .Z(n1288) );
  NANDN U4294 ( .A(n1273), .B(n1288), .Z(n1223) );
  XOR U4295 ( .A(n1230), .B(n1223), .Z(n1249) );
  XNOR U4296 ( .A(n1224), .B(n1249), .Z(n1225) );
  XOR U4297 ( .A(n1226), .B(n1225), .Z(n1262) );
  IV U4298 ( .A(n1262), .Z(n1268) );
  AND U4299 ( .A(n1228), .B(n1227), .Z(n1233) );
  XOR U4300 ( .A(x[48]), .B(n1275), .Z(n1276) );
  XNOR U4301 ( .A(n1323), .B(n1276), .Z(n1278) );
  XOR U4302 ( .A(x[50]), .B(x[55]), .Z(n1303) );
  NANDN U4303 ( .A(n1278), .B(n1303), .Z(n1229) );
  XNOR U4304 ( .A(n1230), .B(n1229), .Z(n1238) );
  XNOR U4305 ( .A(n1231), .B(n1238), .Z(n1232) );
  XOR U4306 ( .A(n1233), .B(n1232), .Z(n1258) );
  XNOR U4307 ( .A(x[52]), .B(n1323), .Z(n1296) );
  ANDN U4308 ( .B(x[48]), .A(n1296), .Z(n1240) );
  XOR U4309 ( .A(x[50]), .B(x[49]), .Z(n1234) );
  XOR U4310 ( .A(n1312), .B(n1234), .Z(n1285) );
  XOR U4311 ( .A(n1286), .B(n1234), .Z(n1291) );
  NAND U4312 ( .A(n1275), .B(n1291), .Z(n1242) );
  XNOR U4313 ( .A(n1285), .B(n1242), .Z(n1236) );
  XNOR U4314 ( .A(x[49]), .B(n1276), .Z(n1235) );
  XNOR U4315 ( .A(n1236), .B(n1235), .Z(n1237) );
  XOR U4316 ( .A(n1238), .B(n1237), .Z(n1239) );
  XOR U4317 ( .A(n1240), .B(n1239), .Z(n1260) );
  NAND U4318 ( .A(n1258), .B(n1260), .Z(n1241) );
  NAND U4319 ( .A(n1268), .B(n1241), .Z(n1252) );
  IV U4320 ( .A(n1258), .Z(n1259) );
  IV U4321 ( .A(n1260), .Z(n1266) );
  XOR U4322 ( .A(n1242), .B(n1296), .Z(n1245) );
  AND U4323 ( .A(n1285), .B(n1276), .Z(n1243) );
  XNOR U4324 ( .A(x[48]), .B(n1243), .Z(n1244) );
  XNOR U4325 ( .A(n1245), .B(n1244), .Z(n1246) );
  XNOR U4326 ( .A(n1247), .B(n1246), .Z(n1248) );
  XNOR U4327 ( .A(n1249), .B(n1248), .Z(n1270) );
  IV U4328 ( .A(n1270), .Z(n1265) );
  XOR U4329 ( .A(n1266), .B(n1265), .Z(n1250) );
  NAND U4330 ( .A(n1259), .B(n1250), .Z(n1251) );
  AND U4331 ( .A(n1252), .B(n1251), .Z(n1331) );
  NAND U4332 ( .A(n1266), .B(n1259), .Z(n1253) );
  NAND U4333 ( .A(n1265), .B(n1253), .Z(n1256) );
  XOR U4334 ( .A(n1259), .B(n1262), .Z(n1254) );
  NAND U4335 ( .A(n1260), .B(n1254), .Z(n1255) );
  AND U4336 ( .A(n1256), .B(n1255), .Z(n1313) );
  XNOR U4337 ( .A(n1331), .B(n1313), .Z(n1287) );
  OR U4338 ( .A(n1287), .B(n1257), .Z(n1280) );
  NAND U4339 ( .A(n1268), .B(n1258), .Z(n1264) );
  AND U4340 ( .A(n1260), .B(n1259), .Z(n1267) );
  XNOR U4341 ( .A(n1265), .B(n1267), .Z(n1261) );
  NAND U4342 ( .A(n1262), .B(n1261), .Z(n1263) );
  AND U4343 ( .A(n1264), .B(n1263), .Z(n1284) );
  NAND U4344 ( .A(n1266), .B(n1265), .Z(n1272) );
  XNOR U4345 ( .A(n1268), .B(n1267), .Z(n1269) );
  NAND U4346 ( .A(n1270), .B(n1269), .Z(n1271) );
  NAND U4347 ( .A(n1272), .B(n1271), .Z(n1325) );
  XNOR U4348 ( .A(n1284), .B(n1325), .Z(n1302) );
  XOR U4349 ( .A(n1302), .B(n1287), .Z(n1289) );
  OR U4350 ( .A(n1289), .B(n1273), .Z(n1274) );
  XNOR U4351 ( .A(n1280), .B(n1274), .Z(n1306) );
  XOR U4352 ( .A(n1284), .B(n1331), .Z(n1292) );
  NANDN U4353 ( .A(n1292), .B(n1275), .Z(n1333) );
  NANDN U4354 ( .A(n1284), .B(n1276), .Z(n1277) );
  XNOR U4355 ( .A(n1333), .B(n1277), .Z(n1311) );
  XOR U4356 ( .A(n1306), .B(n1311), .Z(n1295) );
  NANDN U4357 ( .A(n1278), .B(n1302), .Z(n1279) );
  XNOR U4358 ( .A(n1280), .B(n1279), .Z(n1339) );
  XNOR U4359 ( .A(n1325), .B(n1313), .Z(n1315) );
  NANDN U4360 ( .A(n1315), .B(n1281), .Z(n1298) );
  NAND U4361 ( .A(n1282), .B(n1313), .Z(n1283) );
  XNOR U4362 ( .A(n1298), .B(n1283), .Z(n1330) );
  XOR U4363 ( .A(n1339), .B(n1330), .Z(n1322) );
  XNOR U4364 ( .A(n1295), .B(n1322), .Z(z[48]) );
  ANDN U4365 ( .B(n1285), .A(n1284), .Z(n1294) );
  NANDN U4366 ( .A(n1287), .B(n1286), .Z(n1305) );
  NANDN U4367 ( .A(n1289), .B(n1288), .Z(n1290) );
  XNOR U4368 ( .A(n1305), .B(n1290), .Z(n1334) );
  NANDN U4369 ( .A(n1292), .B(n1291), .Z(n1299) );
  XNOR U4370 ( .A(n1334), .B(n1299), .Z(n1293) );
  XOR U4371 ( .A(n1294), .B(n1293), .Z(n1320) );
  XOR U4372 ( .A(n1320), .B(n1295), .Z(n1338) );
  ANDN U4373 ( .B(n1331), .A(n1296), .Z(n1301) );
  NAND U4374 ( .A(n1323), .B(n1325), .Z(n1297) );
  XNOR U4375 ( .A(n1298), .B(n1297), .Z(n1310) );
  XNOR U4376 ( .A(n1299), .B(n1310), .Z(n1300) );
  XNOR U4377 ( .A(n1301), .B(n1300), .Z(n1308) );
  NAND U4378 ( .A(n1303), .B(n1302), .Z(n1304) );
  XNOR U4379 ( .A(n1305), .B(n1304), .Z(n1316) );
  XNOR U4380 ( .A(n1306), .B(n1316), .Z(n1307) );
  XOR U4381 ( .A(n1308), .B(n1307), .Z(n1319) );
  XNOR U4382 ( .A(n1338), .B(n1319), .Z(z[49]) );
  XOR U4383 ( .A(n1309), .B(z[2]), .Z(z[4]) );
  XNOR U4384 ( .A(n1311), .B(n1310), .Z(z[50]) );
  AND U4385 ( .A(n1313), .B(n1312), .Z(n1318) );
  NANDN U4386 ( .A(n1315), .B(n1314), .Z(n1328) );
  XNOR U4387 ( .A(n1316), .B(n1328), .Z(n1317) );
  XOR U4388 ( .A(n1318), .B(n1317), .Z(n1337) );
  XOR U4389 ( .A(n1320), .B(n1319), .Z(n1321) );
  XOR U4390 ( .A(n1337), .B(n1321), .Z(z[51]) );
  XOR U4391 ( .A(n1322), .B(z[50]), .Z(z[52]) );
  XNOR U4392 ( .A(n1324), .B(n1323), .Z(n1326) );
  NAND U4393 ( .A(n1326), .B(n1325), .Z(n1327) );
  XOR U4394 ( .A(n1328), .B(n1327), .Z(n1329) );
  XNOR U4395 ( .A(n1330), .B(n1329), .Z(n1336) );
  NAND U4396 ( .A(n1331), .B(x[48]), .Z(n1332) );
  XNOR U4397 ( .A(n1333), .B(n1332), .Z(n1340) );
  XNOR U4398 ( .A(n1334), .B(n1340), .Z(n1335) );
  XOR U4399 ( .A(n1336), .B(n1335), .Z(z[53]) );
  XNOR U4400 ( .A(n1338), .B(n1337), .Z(z[54]) );
  XNOR U4401 ( .A(n1340), .B(n1339), .Z(n1341) );
  XNOR U4402 ( .A(z[49]), .B(n1341), .Z(z[55]) );
  IV U4403 ( .A(x[57]), .Z(n1462) );
  XOR U4404 ( .A(x[56]), .B(x[62]), .Z(n1343) );
  XOR U4405 ( .A(x[61]), .B(n1343), .Z(n1461) );
  IV U4406 ( .A(n1461), .Z(n1344) );
  AND U4407 ( .A(n1462), .B(n1344), .Z(n1351) );
  XNOR U4408 ( .A(x[59]), .B(n1462), .Z(n1347) );
  XNOR U4409 ( .A(x[58]), .B(n1347), .Z(n1342) );
  XNOR U4410 ( .A(n1343), .B(n1342), .Z(n1407) );
  IV U4411 ( .A(n1407), .Z(n1353) );
  XNOR U4412 ( .A(n1353), .B(n1461), .Z(n1406) );
  IV U4413 ( .A(x[63]), .Z(n1345) );
  XNOR U4414 ( .A(x[57]), .B(n1345), .Z(n1438) );
  NAND U4415 ( .A(n1406), .B(n1438), .Z(n1356) );
  XNOR U4416 ( .A(n1345), .B(n1344), .Z(n1352) );
  IV U4417 ( .A(n1352), .Z(n1436) );
  XOR U4418 ( .A(n1407), .B(n1436), .Z(n1372) );
  XNOR U4419 ( .A(n1356), .B(n1372), .Z(n1349) );
  XOR U4420 ( .A(x[56]), .B(n1353), .Z(n1382) );
  XOR U4421 ( .A(x[60]), .B(n1345), .Z(n1346) );
  IV U4422 ( .A(n1346), .Z(n1411) );
  NANDN U4423 ( .A(n1382), .B(n1411), .Z(n1355) );
  XNOR U4424 ( .A(n1347), .B(n1346), .Z(n1400) );
  XNOR U4425 ( .A(n1406), .B(n1400), .Z(n1398) );
  XOR U4426 ( .A(x[58]), .B(x[60]), .Z(n1413) );
  NANDN U4427 ( .A(n1398), .B(n1413), .Z(n1348) );
  XOR U4428 ( .A(n1355), .B(n1348), .Z(n1374) );
  XNOR U4429 ( .A(n1349), .B(n1374), .Z(n1350) );
  XOR U4430 ( .A(n1351), .B(n1350), .Z(n1387) );
  IV U4431 ( .A(n1387), .Z(n1393) );
  AND U4432 ( .A(n1353), .B(n1352), .Z(n1358) );
  XOR U4433 ( .A(x[56]), .B(n1400), .Z(n1401) );
  XNOR U4434 ( .A(n1461), .B(n1401), .Z(n1403) );
  XOR U4435 ( .A(x[58]), .B(x[63]), .Z(n1428) );
  NANDN U4436 ( .A(n1403), .B(n1428), .Z(n1354) );
  XNOR U4437 ( .A(n1355), .B(n1354), .Z(n1363) );
  XNOR U4438 ( .A(n1356), .B(n1363), .Z(n1357) );
  XOR U4439 ( .A(n1358), .B(n1357), .Z(n1383) );
  XNOR U4440 ( .A(x[60]), .B(n1461), .Z(n1421) );
  ANDN U4441 ( .B(x[56]), .A(n1421), .Z(n1365) );
  XOR U4442 ( .A(x[58]), .B(x[57]), .Z(n1359) );
  XOR U4443 ( .A(n1436), .B(n1359), .Z(n1410) );
  XOR U4444 ( .A(n1411), .B(n1359), .Z(n1416) );
  NAND U4445 ( .A(n1400), .B(n1416), .Z(n1367) );
  XNOR U4446 ( .A(n1410), .B(n1367), .Z(n1361) );
  XNOR U4447 ( .A(x[57]), .B(n1401), .Z(n1360) );
  XNOR U4448 ( .A(n1361), .B(n1360), .Z(n1362) );
  XOR U4449 ( .A(n1363), .B(n1362), .Z(n1364) );
  XOR U4450 ( .A(n1365), .B(n1364), .Z(n1385) );
  NAND U4451 ( .A(n1383), .B(n1385), .Z(n1366) );
  NAND U4452 ( .A(n1393), .B(n1366), .Z(n1377) );
  IV U4453 ( .A(n1383), .Z(n1384) );
  IV U4454 ( .A(n1385), .Z(n1391) );
  XOR U4455 ( .A(n1367), .B(n1421), .Z(n1370) );
  AND U4456 ( .A(n1410), .B(n1401), .Z(n1368) );
  XNOR U4457 ( .A(x[56]), .B(n1368), .Z(n1369) );
  XNOR U4458 ( .A(n1370), .B(n1369), .Z(n1371) );
  XNOR U4459 ( .A(n1372), .B(n1371), .Z(n1373) );
  XNOR U4460 ( .A(n1374), .B(n1373), .Z(n1395) );
  IV U4461 ( .A(n1395), .Z(n1390) );
  XOR U4462 ( .A(n1391), .B(n1390), .Z(n1375) );
  NAND U4463 ( .A(n1384), .B(n1375), .Z(n1376) );
  AND U4464 ( .A(n1377), .B(n1376), .Z(n1469) );
  NAND U4465 ( .A(n1391), .B(n1384), .Z(n1378) );
  NAND U4466 ( .A(n1390), .B(n1378), .Z(n1381) );
  XOR U4467 ( .A(n1384), .B(n1387), .Z(n1379) );
  NAND U4468 ( .A(n1385), .B(n1379), .Z(n1380) );
  AND U4469 ( .A(n1381), .B(n1380), .Z(n1437) );
  XNOR U4470 ( .A(n1469), .B(n1437), .Z(n1412) );
  OR U4471 ( .A(n1412), .B(n1382), .Z(n1405) );
  NAND U4472 ( .A(n1393), .B(n1383), .Z(n1389) );
  AND U4473 ( .A(n1385), .B(n1384), .Z(n1392) );
  XNOR U4474 ( .A(n1390), .B(n1392), .Z(n1386) );
  NAND U4475 ( .A(n1387), .B(n1386), .Z(n1388) );
  AND U4476 ( .A(n1389), .B(n1388), .Z(n1409) );
  NAND U4477 ( .A(n1391), .B(n1390), .Z(n1397) );
  XNOR U4478 ( .A(n1393), .B(n1392), .Z(n1394) );
  NAND U4479 ( .A(n1395), .B(n1394), .Z(n1396) );
  NAND U4480 ( .A(n1397), .B(n1396), .Z(n1463) );
  XNOR U4481 ( .A(n1409), .B(n1463), .Z(n1427) );
  XOR U4482 ( .A(n1427), .B(n1412), .Z(n1414) );
  OR U4483 ( .A(n1414), .B(n1398), .Z(n1399) );
  XNOR U4484 ( .A(n1405), .B(n1399), .Z(n1431) );
  XOR U4485 ( .A(n1409), .B(n1469), .Z(n1417) );
  NANDN U4486 ( .A(n1417), .B(n1400), .Z(n1471) );
  NANDN U4487 ( .A(n1409), .B(n1401), .Z(n1402) );
  XNOR U4488 ( .A(n1471), .B(n1402), .Z(n1435) );
  XOR U4489 ( .A(n1431), .B(n1435), .Z(n1420) );
  NANDN U4490 ( .A(n1403), .B(n1427), .Z(n1404) );
  XNOR U4491 ( .A(n1405), .B(n1404), .Z(n1477) );
  XNOR U4492 ( .A(n1463), .B(n1437), .Z(n1439) );
  NANDN U4493 ( .A(n1439), .B(n1406), .Z(n1423) );
  NAND U4494 ( .A(n1407), .B(n1437), .Z(n1408) );
  XNOR U4495 ( .A(n1423), .B(n1408), .Z(n1468) );
  XOR U4496 ( .A(n1477), .B(n1468), .Z(n1460) );
  XNOR U4497 ( .A(n1420), .B(n1460), .Z(z[56]) );
  ANDN U4498 ( .B(n1410), .A(n1409), .Z(n1419) );
  NANDN U4499 ( .A(n1412), .B(n1411), .Z(n1430) );
  NANDN U4500 ( .A(n1414), .B(n1413), .Z(n1415) );
  XNOR U4501 ( .A(n1430), .B(n1415), .Z(n1472) );
  NANDN U4502 ( .A(n1417), .B(n1416), .Z(n1424) );
  XNOR U4503 ( .A(n1472), .B(n1424), .Z(n1418) );
  XOR U4504 ( .A(n1419), .B(n1418), .Z(n1444) );
  XOR U4505 ( .A(n1444), .B(n1420), .Z(n1476) );
  ANDN U4506 ( .B(n1469), .A(n1421), .Z(n1426) );
  NAND U4507 ( .A(n1461), .B(n1463), .Z(n1422) );
  XNOR U4508 ( .A(n1423), .B(n1422), .Z(n1434) );
  XNOR U4509 ( .A(n1424), .B(n1434), .Z(n1425) );
  XNOR U4510 ( .A(n1426), .B(n1425), .Z(n1433) );
  NAND U4511 ( .A(n1428), .B(n1427), .Z(n1429) );
  XNOR U4512 ( .A(n1430), .B(n1429), .Z(n1440) );
  XNOR U4513 ( .A(n1431), .B(n1440), .Z(n1432) );
  XOR U4514 ( .A(n1433), .B(n1432), .Z(n1443) );
  XNOR U4515 ( .A(n1476), .B(n1443), .Z(z[57]) );
  XNOR U4516 ( .A(n1435), .B(n1434), .Z(z[58]) );
  AND U4517 ( .A(n1437), .B(n1436), .Z(n1442) );
  NANDN U4518 ( .A(n1439), .B(n1438), .Z(n1466) );
  XNOR U4519 ( .A(n1440), .B(n1466), .Z(n1441) );
  XOR U4520 ( .A(n1442), .B(n1441), .Z(n1475) );
  XOR U4521 ( .A(n1444), .B(n1443), .Z(n1445) );
  XOR U4522 ( .A(n1475), .B(n1445), .Z(z[59]) );
  XNOR U4523 ( .A(n1447), .B(n1446), .Z(n1449) );
  NAND U4524 ( .A(n1449), .B(n1448), .Z(n1450) );
  XOR U4525 ( .A(n1451), .B(n1450), .Z(n1452) );
  XNOR U4526 ( .A(n1453), .B(n1452), .Z(n1459) );
  NAND U4527 ( .A(n1454), .B(x[0]), .Z(n1455) );
  XNOR U4528 ( .A(n1456), .B(n1455), .Z(n1731) );
  XNOR U4529 ( .A(n1457), .B(n1731), .Z(n1458) );
  XOR U4530 ( .A(n1459), .B(n1458), .Z(z[5]) );
  XOR U4531 ( .A(n1460), .B(z[58]), .Z(z[60]) );
  XNOR U4532 ( .A(n1462), .B(n1461), .Z(n1464) );
  NAND U4533 ( .A(n1464), .B(n1463), .Z(n1465) );
  XOR U4534 ( .A(n1466), .B(n1465), .Z(n1467) );
  XNOR U4535 ( .A(n1468), .B(n1467), .Z(n1474) );
  NAND U4536 ( .A(n1469), .B(x[56]), .Z(n1470) );
  XNOR U4537 ( .A(n1471), .B(n1470), .Z(n1478) );
  XNOR U4538 ( .A(n1472), .B(n1478), .Z(n1473) );
  XOR U4539 ( .A(n1474), .B(n1473), .Z(z[61]) );
  XNOR U4540 ( .A(n1476), .B(n1475), .Z(z[62]) );
  XNOR U4541 ( .A(n1478), .B(n1477), .Z(n1479) );
  XNOR U4542 ( .A(z[57]), .B(n1479), .Z(z[63]) );
  IV U4543 ( .A(x[65]), .Z(n1586) );
  XOR U4544 ( .A(x[64]), .B(x[70]), .Z(n1481) );
  XOR U4545 ( .A(x[69]), .B(n1481), .Z(n1585) );
  IV U4546 ( .A(n1585), .Z(n1482) );
  AND U4547 ( .A(n1586), .B(n1482), .Z(n1489) );
  XNOR U4548 ( .A(x[67]), .B(n1586), .Z(n1485) );
  XNOR U4549 ( .A(x[66]), .B(n1485), .Z(n1480) );
  XNOR U4550 ( .A(n1481), .B(n1480), .Z(n1545) );
  IV U4551 ( .A(n1545), .Z(n1491) );
  XNOR U4552 ( .A(n1491), .B(n1585), .Z(n1544) );
  IV U4553 ( .A(x[71]), .Z(n1483) );
  XNOR U4554 ( .A(x[65]), .B(n1483), .Z(n1576) );
  NAND U4555 ( .A(n1544), .B(n1576), .Z(n1494) );
  XNOR U4556 ( .A(n1483), .B(n1482), .Z(n1490) );
  IV U4557 ( .A(n1490), .Z(n1574) );
  XOR U4558 ( .A(n1545), .B(n1574), .Z(n1510) );
  XNOR U4559 ( .A(n1494), .B(n1510), .Z(n1487) );
  XOR U4560 ( .A(x[64]), .B(n1491), .Z(n1520) );
  XOR U4561 ( .A(x[68]), .B(n1483), .Z(n1484) );
  IV U4562 ( .A(n1484), .Z(n1549) );
  NANDN U4563 ( .A(n1520), .B(n1549), .Z(n1493) );
  XNOR U4564 ( .A(n1485), .B(n1484), .Z(n1538) );
  XNOR U4565 ( .A(n1544), .B(n1538), .Z(n1536) );
  XOR U4566 ( .A(x[66]), .B(x[68]), .Z(n1551) );
  NANDN U4567 ( .A(n1536), .B(n1551), .Z(n1486) );
  XOR U4568 ( .A(n1493), .B(n1486), .Z(n1512) );
  XNOR U4569 ( .A(n1487), .B(n1512), .Z(n1488) );
  XOR U4570 ( .A(n1489), .B(n1488), .Z(n1525) );
  IV U4571 ( .A(n1525), .Z(n1531) );
  AND U4572 ( .A(n1491), .B(n1490), .Z(n1496) );
  XOR U4573 ( .A(x[64]), .B(n1538), .Z(n1539) );
  XNOR U4574 ( .A(n1585), .B(n1539), .Z(n1541) );
  XOR U4575 ( .A(x[66]), .B(x[71]), .Z(n1566) );
  NANDN U4576 ( .A(n1541), .B(n1566), .Z(n1492) );
  XNOR U4577 ( .A(n1493), .B(n1492), .Z(n1501) );
  XNOR U4578 ( .A(n1494), .B(n1501), .Z(n1495) );
  XOR U4579 ( .A(n1496), .B(n1495), .Z(n1521) );
  XNOR U4580 ( .A(x[68]), .B(n1585), .Z(n1559) );
  ANDN U4581 ( .B(x[64]), .A(n1559), .Z(n1503) );
  XOR U4582 ( .A(x[66]), .B(x[65]), .Z(n1497) );
  XOR U4583 ( .A(n1574), .B(n1497), .Z(n1548) );
  XOR U4584 ( .A(n1549), .B(n1497), .Z(n1554) );
  NAND U4585 ( .A(n1538), .B(n1554), .Z(n1505) );
  XNOR U4586 ( .A(n1548), .B(n1505), .Z(n1499) );
  XNOR U4587 ( .A(x[65]), .B(n1539), .Z(n1498) );
  XNOR U4588 ( .A(n1499), .B(n1498), .Z(n1500) );
  XOR U4589 ( .A(n1501), .B(n1500), .Z(n1502) );
  XOR U4590 ( .A(n1503), .B(n1502), .Z(n1523) );
  NAND U4591 ( .A(n1521), .B(n1523), .Z(n1504) );
  NAND U4592 ( .A(n1531), .B(n1504), .Z(n1515) );
  IV U4593 ( .A(n1521), .Z(n1522) );
  IV U4594 ( .A(n1523), .Z(n1529) );
  XOR U4595 ( .A(n1505), .B(n1559), .Z(n1508) );
  AND U4596 ( .A(n1548), .B(n1539), .Z(n1506) );
  XNOR U4597 ( .A(x[64]), .B(n1506), .Z(n1507) );
  XNOR U4598 ( .A(n1508), .B(n1507), .Z(n1509) );
  XNOR U4599 ( .A(n1510), .B(n1509), .Z(n1511) );
  XNOR U4600 ( .A(n1512), .B(n1511), .Z(n1533) );
  IV U4601 ( .A(n1533), .Z(n1528) );
  XOR U4602 ( .A(n1529), .B(n1528), .Z(n1513) );
  NAND U4603 ( .A(n1522), .B(n1513), .Z(n1514) );
  AND U4604 ( .A(n1515), .B(n1514), .Z(n1593) );
  NAND U4605 ( .A(n1529), .B(n1522), .Z(n1516) );
  NAND U4606 ( .A(n1528), .B(n1516), .Z(n1519) );
  XOR U4607 ( .A(n1522), .B(n1525), .Z(n1517) );
  NAND U4608 ( .A(n1523), .B(n1517), .Z(n1518) );
  AND U4609 ( .A(n1519), .B(n1518), .Z(n1575) );
  XNOR U4610 ( .A(n1593), .B(n1575), .Z(n1550) );
  OR U4611 ( .A(n1550), .B(n1520), .Z(n1543) );
  NAND U4612 ( .A(n1531), .B(n1521), .Z(n1527) );
  AND U4613 ( .A(n1523), .B(n1522), .Z(n1530) );
  XNOR U4614 ( .A(n1528), .B(n1530), .Z(n1524) );
  NAND U4615 ( .A(n1525), .B(n1524), .Z(n1526) );
  AND U4616 ( .A(n1527), .B(n1526), .Z(n1547) );
  NAND U4617 ( .A(n1529), .B(n1528), .Z(n1535) );
  XNOR U4618 ( .A(n1531), .B(n1530), .Z(n1532) );
  NAND U4619 ( .A(n1533), .B(n1532), .Z(n1534) );
  NAND U4620 ( .A(n1535), .B(n1534), .Z(n1587) );
  XNOR U4621 ( .A(n1547), .B(n1587), .Z(n1565) );
  XOR U4622 ( .A(n1565), .B(n1550), .Z(n1552) );
  OR U4623 ( .A(n1552), .B(n1536), .Z(n1537) );
  XNOR U4624 ( .A(n1543), .B(n1537), .Z(n1569) );
  XOR U4625 ( .A(n1547), .B(n1593), .Z(n1555) );
  NANDN U4626 ( .A(n1555), .B(n1538), .Z(n1595) );
  NANDN U4627 ( .A(n1547), .B(n1539), .Z(n1540) );
  XNOR U4628 ( .A(n1595), .B(n1540), .Z(n1573) );
  XOR U4629 ( .A(n1569), .B(n1573), .Z(n1558) );
  NANDN U4630 ( .A(n1541), .B(n1565), .Z(n1542) );
  XNOR U4631 ( .A(n1543), .B(n1542), .Z(n1603) );
  XNOR U4632 ( .A(n1587), .B(n1575), .Z(n1577) );
  NANDN U4633 ( .A(n1577), .B(n1544), .Z(n1561) );
  NAND U4634 ( .A(n1545), .B(n1575), .Z(n1546) );
  XNOR U4635 ( .A(n1561), .B(n1546), .Z(n1592) );
  XOR U4636 ( .A(n1603), .B(n1592), .Z(n1584) );
  XNOR U4637 ( .A(n1558), .B(n1584), .Z(z[64]) );
  ANDN U4638 ( .B(n1548), .A(n1547), .Z(n1557) );
  NANDN U4639 ( .A(n1550), .B(n1549), .Z(n1568) );
  NANDN U4640 ( .A(n1552), .B(n1551), .Z(n1553) );
  XNOR U4641 ( .A(n1568), .B(n1553), .Z(n1596) );
  NANDN U4642 ( .A(n1555), .B(n1554), .Z(n1562) );
  XNOR U4643 ( .A(n1596), .B(n1562), .Z(n1556) );
  XOR U4644 ( .A(n1557), .B(n1556), .Z(n1582) );
  XOR U4645 ( .A(n1582), .B(n1558), .Z(n1602) );
  ANDN U4646 ( .B(n1593), .A(n1559), .Z(n1564) );
  NAND U4647 ( .A(n1585), .B(n1587), .Z(n1560) );
  XNOR U4648 ( .A(n1561), .B(n1560), .Z(n1572) );
  XNOR U4649 ( .A(n1562), .B(n1572), .Z(n1563) );
  XNOR U4650 ( .A(n1564), .B(n1563), .Z(n1571) );
  NAND U4651 ( .A(n1566), .B(n1565), .Z(n1567) );
  XNOR U4652 ( .A(n1568), .B(n1567), .Z(n1578) );
  XNOR U4653 ( .A(n1569), .B(n1578), .Z(n1570) );
  XOR U4654 ( .A(n1571), .B(n1570), .Z(n1581) );
  XNOR U4655 ( .A(n1602), .B(n1581), .Z(z[65]) );
  XNOR U4656 ( .A(n1573), .B(n1572), .Z(z[66]) );
  AND U4657 ( .A(n1575), .B(n1574), .Z(n1580) );
  NANDN U4658 ( .A(n1577), .B(n1576), .Z(n1590) );
  XNOR U4659 ( .A(n1578), .B(n1590), .Z(n1579) );
  XOR U4660 ( .A(n1580), .B(n1579), .Z(n1601) );
  XOR U4661 ( .A(n1582), .B(n1581), .Z(n1583) );
  XOR U4662 ( .A(n1601), .B(n1583), .Z(z[67]) );
  XOR U4663 ( .A(n1584), .B(z[66]), .Z(z[68]) );
  XNOR U4664 ( .A(n1586), .B(n1585), .Z(n1588) );
  NAND U4665 ( .A(n1588), .B(n1587), .Z(n1589) );
  XOR U4666 ( .A(n1590), .B(n1589), .Z(n1591) );
  XNOR U4667 ( .A(n1592), .B(n1591), .Z(n1598) );
  NAND U4668 ( .A(n1593), .B(x[64]), .Z(n1594) );
  XNOR U4669 ( .A(n1595), .B(n1594), .Z(n1604) );
  XNOR U4670 ( .A(n1596), .B(n1604), .Z(n1597) );
  XOR U4671 ( .A(n1598), .B(n1597), .Z(z[69]) );
  XNOR U4672 ( .A(n1600), .B(n1599), .Z(z[6]) );
  XNOR U4673 ( .A(n1602), .B(n1601), .Z(z[70]) );
  XNOR U4674 ( .A(n1604), .B(n1603), .Z(n1605) );
  XNOR U4675 ( .A(z[65]), .B(n1605), .Z(z[71]) );
  IV U4676 ( .A(x[73]), .Z(n1712) );
  XOR U4677 ( .A(x[72]), .B(x[78]), .Z(n1607) );
  XOR U4678 ( .A(x[77]), .B(n1607), .Z(n1711) );
  IV U4679 ( .A(n1711), .Z(n1608) );
  AND U4680 ( .A(n1712), .B(n1608), .Z(n1615) );
  XNOR U4681 ( .A(x[75]), .B(n1712), .Z(n1611) );
  XNOR U4682 ( .A(x[74]), .B(n1611), .Z(n1606) );
  XNOR U4683 ( .A(n1607), .B(n1606), .Z(n1671) );
  IV U4684 ( .A(n1671), .Z(n1617) );
  XNOR U4685 ( .A(n1617), .B(n1711), .Z(n1670) );
  IV U4686 ( .A(x[79]), .Z(n1609) );
  XNOR U4687 ( .A(x[73]), .B(n1609), .Z(n1702) );
  NAND U4688 ( .A(n1670), .B(n1702), .Z(n1620) );
  XNOR U4689 ( .A(n1609), .B(n1608), .Z(n1616) );
  IV U4690 ( .A(n1616), .Z(n1700) );
  XOR U4691 ( .A(n1671), .B(n1700), .Z(n1636) );
  XNOR U4692 ( .A(n1620), .B(n1636), .Z(n1613) );
  XOR U4693 ( .A(x[72]), .B(n1617), .Z(n1646) );
  XOR U4694 ( .A(x[76]), .B(n1609), .Z(n1610) );
  IV U4695 ( .A(n1610), .Z(n1675) );
  NANDN U4696 ( .A(n1646), .B(n1675), .Z(n1619) );
  XNOR U4697 ( .A(n1611), .B(n1610), .Z(n1664) );
  XNOR U4698 ( .A(n1670), .B(n1664), .Z(n1662) );
  XOR U4699 ( .A(x[74]), .B(x[76]), .Z(n1677) );
  NANDN U4700 ( .A(n1662), .B(n1677), .Z(n1612) );
  XOR U4701 ( .A(n1619), .B(n1612), .Z(n1638) );
  XNOR U4702 ( .A(n1613), .B(n1638), .Z(n1614) );
  XOR U4703 ( .A(n1615), .B(n1614), .Z(n1651) );
  IV U4704 ( .A(n1651), .Z(n1657) );
  AND U4705 ( .A(n1617), .B(n1616), .Z(n1622) );
  XOR U4706 ( .A(x[72]), .B(n1664), .Z(n1665) );
  XNOR U4707 ( .A(n1711), .B(n1665), .Z(n1667) );
  XOR U4708 ( .A(x[74]), .B(x[79]), .Z(n1692) );
  NANDN U4709 ( .A(n1667), .B(n1692), .Z(n1618) );
  XNOR U4710 ( .A(n1619), .B(n1618), .Z(n1627) );
  XNOR U4711 ( .A(n1620), .B(n1627), .Z(n1621) );
  XOR U4712 ( .A(n1622), .B(n1621), .Z(n1647) );
  XNOR U4713 ( .A(x[76]), .B(n1711), .Z(n1685) );
  ANDN U4714 ( .B(x[72]), .A(n1685), .Z(n1629) );
  XOR U4715 ( .A(x[74]), .B(x[73]), .Z(n1623) );
  XOR U4716 ( .A(n1700), .B(n1623), .Z(n1674) );
  XOR U4717 ( .A(n1675), .B(n1623), .Z(n1680) );
  NAND U4718 ( .A(n1664), .B(n1680), .Z(n1631) );
  XNOR U4719 ( .A(n1674), .B(n1631), .Z(n1625) );
  XNOR U4720 ( .A(x[73]), .B(n1665), .Z(n1624) );
  XNOR U4721 ( .A(n1625), .B(n1624), .Z(n1626) );
  XOR U4722 ( .A(n1627), .B(n1626), .Z(n1628) );
  XOR U4723 ( .A(n1629), .B(n1628), .Z(n1649) );
  NAND U4724 ( .A(n1647), .B(n1649), .Z(n1630) );
  NAND U4725 ( .A(n1657), .B(n1630), .Z(n1641) );
  IV U4726 ( .A(n1647), .Z(n1648) );
  IV U4727 ( .A(n1649), .Z(n1655) );
  XOR U4728 ( .A(n1631), .B(n1685), .Z(n1634) );
  AND U4729 ( .A(n1674), .B(n1665), .Z(n1632) );
  XNOR U4730 ( .A(x[72]), .B(n1632), .Z(n1633) );
  XNOR U4731 ( .A(n1634), .B(n1633), .Z(n1635) );
  XNOR U4732 ( .A(n1636), .B(n1635), .Z(n1637) );
  XNOR U4733 ( .A(n1638), .B(n1637), .Z(n1659) );
  IV U4734 ( .A(n1659), .Z(n1654) );
  XOR U4735 ( .A(n1655), .B(n1654), .Z(n1639) );
  NAND U4736 ( .A(n1648), .B(n1639), .Z(n1640) );
  AND U4737 ( .A(n1641), .B(n1640), .Z(n1719) );
  NAND U4738 ( .A(n1655), .B(n1648), .Z(n1642) );
  NAND U4739 ( .A(n1654), .B(n1642), .Z(n1645) );
  XOR U4740 ( .A(n1648), .B(n1651), .Z(n1643) );
  NAND U4741 ( .A(n1649), .B(n1643), .Z(n1644) );
  AND U4742 ( .A(n1645), .B(n1644), .Z(n1701) );
  XNOR U4743 ( .A(n1719), .B(n1701), .Z(n1676) );
  OR U4744 ( .A(n1676), .B(n1646), .Z(n1669) );
  NAND U4745 ( .A(n1657), .B(n1647), .Z(n1653) );
  AND U4746 ( .A(n1649), .B(n1648), .Z(n1656) );
  XNOR U4747 ( .A(n1654), .B(n1656), .Z(n1650) );
  NAND U4748 ( .A(n1651), .B(n1650), .Z(n1652) );
  AND U4749 ( .A(n1653), .B(n1652), .Z(n1673) );
  NAND U4750 ( .A(n1655), .B(n1654), .Z(n1661) );
  XNOR U4751 ( .A(n1657), .B(n1656), .Z(n1658) );
  NAND U4752 ( .A(n1659), .B(n1658), .Z(n1660) );
  NAND U4753 ( .A(n1661), .B(n1660), .Z(n1713) );
  XNOR U4754 ( .A(n1673), .B(n1713), .Z(n1691) );
  XOR U4755 ( .A(n1691), .B(n1676), .Z(n1678) );
  OR U4756 ( .A(n1678), .B(n1662), .Z(n1663) );
  XNOR U4757 ( .A(n1669), .B(n1663), .Z(n1695) );
  XOR U4758 ( .A(n1673), .B(n1719), .Z(n1681) );
  NANDN U4759 ( .A(n1681), .B(n1664), .Z(n1721) );
  NANDN U4760 ( .A(n1673), .B(n1665), .Z(n1666) );
  XNOR U4761 ( .A(n1721), .B(n1666), .Z(n1699) );
  XOR U4762 ( .A(n1695), .B(n1699), .Z(n1684) );
  NANDN U4763 ( .A(n1667), .B(n1691), .Z(n1668) );
  XNOR U4764 ( .A(n1669), .B(n1668), .Z(n1727) );
  XNOR U4765 ( .A(n1713), .B(n1701), .Z(n1703) );
  NANDN U4766 ( .A(n1703), .B(n1670), .Z(n1687) );
  NAND U4767 ( .A(n1671), .B(n1701), .Z(n1672) );
  XNOR U4768 ( .A(n1687), .B(n1672), .Z(n1718) );
  XOR U4769 ( .A(n1727), .B(n1718), .Z(n1710) );
  XNOR U4770 ( .A(n1684), .B(n1710), .Z(z[72]) );
  ANDN U4771 ( .B(n1674), .A(n1673), .Z(n1683) );
  NANDN U4772 ( .A(n1676), .B(n1675), .Z(n1694) );
  NANDN U4773 ( .A(n1678), .B(n1677), .Z(n1679) );
  XNOR U4774 ( .A(n1694), .B(n1679), .Z(n1722) );
  NANDN U4775 ( .A(n1681), .B(n1680), .Z(n1688) );
  XNOR U4776 ( .A(n1722), .B(n1688), .Z(n1682) );
  XOR U4777 ( .A(n1683), .B(n1682), .Z(n1708) );
  XOR U4778 ( .A(n1708), .B(n1684), .Z(n1726) );
  ANDN U4779 ( .B(n1719), .A(n1685), .Z(n1690) );
  NAND U4780 ( .A(n1711), .B(n1713), .Z(n1686) );
  XNOR U4781 ( .A(n1687), .B(n1686), .Z(n1698) );
  XNOR U4782 ( .A(n1688), .B(n1698), .Z(n1689) );
  XNOR U4783 ( .A(n1690), .B(n1689), .Z(n1697) );
  NAND U4784 ( .A(n1692), .B(n1691), .Z(n1693) );
  XNOR U4785 ( .A(n1694), .B(n1693), .Z(n1704) );
  XNOR U4786 ( .A(n1695), .B(n1704), .Z(n1696) );
  XOR U4787 ( .A(n1697), .B(n1696), .Z(n1707) );
  XNOR U4788 ( .A(n1726), .B(n1707), .Z(z[73]) );
  XNOR U4789 ( .A(n1699), .B(n1698), .Z(z[74]) );
  AND U4790 ( .A(n1701), .B(n1700), .Z(n1706) );
  NANDN U4791 ( .A(n1703), .B(n1702), .Z(n1716) );
  XNOR U4792 ( .A(n1704), .B(n1716), .Z(n1705) );
  XOR U4793 ( .A(n1706), .B(n1705), .Z(n1725) );
  XOR U4794 ( .A(n1708), .B(n1707), .Z(n1709) );
  XOR U4795 ( .A(n1725), .B(n1709), .Z(z[75]) );
  XOR U4796 ( .A(n1710), .B(z[74]), .Z(z[76]) );
  XNOR U4797 ( .A(n1712), .B(n1711), .Z(n1714) );
  NAND U4798 ( .A(n1714), .B(n1713), .Z(n1715) );
  XOR U4799 ( .A(n1716), .B(n1715), .Z(n1717) );
  XNOR U4800 ( .A(n1718), .B(n1717), .Z(n1724) );
  NAND U4801 ( .A(n1719), .B(x[72]), .Z(n1720) );
  XNOR U4802 ( .A(n1721), .B(n1720), .Z(n1728) );
  XNOR U4803 ( .A(n1722), .B(n1728), .Z(n1723) );
  XOR U4804 ( .A(n1724), .B(n1723), .Z(z[77]) );
  XNOR U4805 ( .A(n1726), .B(n1725), .Z(z[78]) );
  XNOR U4806 ( .A(n1728), .B(n1727), .Z(n1729) );
  XNOR U4807 ( .A(z[73]), .B(n1729), .Z(z[79]) );
  XNOR U4808 ( .A(n1731), .B(n1730), .Z(n1732) );
  XNOR U4809 ( .A(z[1]), .B(n1732), .Z(z[7]) );
  XOR U4810 ( .A(x[80]), .B(x[86]), .Z(n1733) );
  XOR U4811 ( .A(x[85]), .B(n1733), .Z(n1838) );
  IV U4812 ( .A(n1838), .Z(n1735) );
  IV U4813 ( .A(x[81]), .Z(n1837) );
  NAND U4814 ( .A(n1735), .B(n1837), .Z(n1742) );
  XOR U4815 ( .A(x[83]), .B(x[81]), .Z(n1738) );
  XNOR U4816 ( .A(x[82]), .B(n1733), .Z(n1734) );
  XNOR U4817 ( .A(n1738), .B(n1734), .Z(n1797) );
  XNOR U4818 ( .A(n1735), .B(n1797), .Z(n1796) );
  IV U4819 ( .A(x[87]), .Z(n1736) );
  XNOR U4820 ( .A(x[81]), .B(n1736), .Z(n1828) );
  NAND U4821 ( .A(n1796), .B(n1828), .Z(n1745) );
  XNOR U4822 ( .A(n1735), .B(n1736), .Z(n1826) );
  XOR U4823 ( .A(n1797), .B(n1826), .Z(n1753) );
  XOR U4824 ( .A(n1745), .B(n1753), .Z(n1740) );
  XNOR U4825 ( .A(x[80]), .B(n1797), .Z(n1772) );
  XOR U4826 ( .A(x[84]), .B(n1736), .Z(n1737) );
  IV U4827 ( .A(n1737), .Z(n1801) );
  NANDN U4828 ( .A(n1772), .B(n1801), .Z(n1744) );
  XOR U4829 ( .A(n1738), .B(n1737), .Z(n1790) );
  XOR U4830 ( .A(n1796), .B(n1790), .Z(n1788) );
  XOR U4831 ( .A(x[82]), .B(x[84]), .Z(n1803) );
  NANDN U4832 ( .A(n1788), .B(n1803), .Z(n1739) );
  XNOR U4833 ( .A(n1744), .B(n1739), .Z(n1749) );
  XOR U4834 ( .A(n1740), .B(n1749), .Z(n1741) );
  XOR U4835 ( .A(n1742), .B(n1741), .Z(n1783) );
  IV U4836 ( .A(n1783), .Z(n1777) );
  ANDN U4837 ( .B(n1826), .A(n1797), .Z(n1747) );
  XNOR U4838 ( .A(x[80]), .B(n1790), .Z(n1791) );
  XNOR U4839 ( .A(n1838), .B(n1791), .Z(n1793) );
  XOR U4840 ( .A(x[82]), .B(x[87]), .Z(n1818) );
  NANDN U4841 ( .A(n1793), .B(n1818), .Z(n1743) );
  XNOR U4842 ( .A(n1744), .B(n1743), .Z(n1760) );
  XNOR U4843 ( .A(n1745), .B(n1760), .Z(n1746) );
  XOR U4844 ( .A(n1747), .B(n1746), .Z(n1773) );
  NAND U4845 ( .A(n1777), .B(n1773), .Z(n1767) );
  IV U4846 ( .A(n1773), .Z(n1774) );
  XOR U4847 ( .A(n1783), .B(n1774), .Z(n1765) );
  XOR U4848 ( .A(x[82]), .B(x[81]), .Z(n1748) );
  XNOR U4849 ( .A(n1826), .B(n1748), .Z(n1800) );
  NAND U4850 ( .A(n1800), .B(n1791), .Z(n1755) );
  XNOR U4851 ( .A(x[84]), .B(n1838), .Z(n1811) );
  XOR U4852 ( .A(n1801), .B(n1748), .Z(n1806) );
  NANDN U4853 ( .A(n1790), .B(n1806), .Z(n1756) );
  XOR U4854 ( .A(n1811), .B(n1756), .Z(n1751) );
  XOR U4855 ( .A(x[80]), .B(n1749), .Z(n1750) );
  XNOR U4856 ( .A(n1751), .B(n1750), .Z(n1752) );
  XOR U4857 ( .A(n1753), .B(n1752), .Z(n1754) );
  XOR U4858 ( .A(n1755), .B(n1754), .Z(n1785) );
  IV U4859 ( .A(n1785), .Z(n1780) );
  AND U4860 ( .A(n1777), .B(n1780), .Z(n1763) );
  ANDN U4861 ( .B(x[80]), .A(n1811), .Z(n1762) );
  XNOR U4862 ( .A(n1800), .B(n1756), .Z(n1758) );
  XNOR U4863 ( .A(x[81]), .B(n1791), .Z(n1757) );
  XNOR U4864 ( .A(n1758), .B(n1757), .Z(n1759) );
  XOR U4865 ( .A(n1760), .B(n1759), .Z(n1761) );
  XOR U4866 ( .A(n1762), .B(n1761), .Z(n1775) );
  IV U4867 ( .A(n1775), .Z(n1781) );
  XNOR U4868 ( .A(n1763), .B(n1781), .Z(n1764) );
  NAND U4869 ( .A(n1765), .B(n1764), .Z(n1766) );
  NAND U4870 ( .A(n1767), .B(n1766), .Z(n1845) );
  NAND U4871 ( .A(n1781), .B(n1774), .Z(n1768) );
  NAND U4872 ( .A(n1780), .B(n1768), .Z(n1771) );
  XOR U4873 ( .A(n1774), .B(n1777), .Z(n1769) );
  NAND U4874 ( .A(n1775), .B(n1769), .Z(n1770) );
  AND U4875 ( .A(n1771), .B(n1770), .Z(n1827) );
  XNOR U4876 ( .A(n1845), .B(n1827), .Z(n1802) );
  OR U4877 ( .A(n1802), .B(n1772), .Z(n1795) );
  NAND U4878 ( .A(n1783), .B(n1773), .Z(n1779) );
  AND U4879 ( .A(n1775), .B(n1774), .Z(n1782) );
  XNOR U4880 ( .A(n1782), .B(n1780), .Z(n1776) );
  NAND U4881 ( .A(n1777), .B(n1776), .Z(n1778) );
  AND U4882 ( .A(n1779), .B(n1778), .Z(n1799) );
  NAND U4883 ( .A(n1781), .B(n1780), .Z(n1787) );
  XNOR U4884 ( .A(n1783), .B(n1782), .Z(n1784) );
  NAND U4885 ( .A(n1785), .B(n1784), .Z(n1786) );
  NAND U4886 ( .A(n1787), .B(n1786), .Z(n1839) );
  XNOR U4887 ( .A(n1799), .B(n1839), .Z(n1817) );
  XOR U4888 ( .A(n1817), .B(n1802), .Z(n1804) );
  OR U4889 ( .A(n1804), .B(n1788), .Z(n1789) );
  XNOR U4890 ( .A(n1795), .B(n1789), .Z(n1821) );
  XOR U4891 ( .A(n1799), .B(n1845), .Z(n1807) );
  OR U4892 ( .A(n1790), .B(n1807), .Z(n1847) );
  NANDN U4893 ( .A(n1799), .B(n1791), .Z(n1792) );
  XNOR U4894 ( .A(n1847), .B(n1792), .Z(n1825) );
  XOR U4895 ( .A(n1821), .B(n1825), .Z(n1810) );
  NANDN U4896 ( .A(n1793), .B(n1817), .Z(n1794) );
  XNOR U4897 ( .A(n1795), .B(n1794), .Z(n1853) );
  XNOR U4898 ( .A(n1839), .B(n1827), .Z(n1829) );
  NANDN U4899 ( .A(n1829), .B(n1796), .Z(n1813) );
  NAND U4900 ( .A(n1797), .B(n1827), .Z(n1798) );
  XNOR U4901 ( .A(n1813), .B(n1798), .Z(n1844) );
  XOR U4902 ( .A(n1853), .B(n1844), .Z(n1836) );
  XNOR U4903 ( .A(n1810), .B(n1836), .Z(z[80]) );
  ANDN U4904 ( .B(n1800), .A(n1799), .Z(n1809) );
  NANDN U4905 ( .A(n1802), .B(n1801), .Z(n1820) );
  NANDN U4906 ( .A(n1804), .B(n1803), .Z(n1805) );
  XNOR U4907 ( .A(n1820), .B(n1805), .Z(n1848) );
  NANDN U4908 ( .A(n1807), .B(n1806), .Z(n1814) );
  XNOR U4909 ( .A(n1848), .B(n1814), .Z(n1808) );
  XOR U4910 ( .A(n1809), .B(n1808), .Z(n1834) );
  XOR U4911 ( .A(n1834), .B(n1810), .Z(n1852) );
  ANDN U4912 ( .B(n1845), .A(n1811), .Z(n1816) );
  NAND U4913 ( .A(n1838), .B(n1839), .Z(n1812) );
  XNOR U4914 ( .A(n1813), .B(n1812), .Z(n1824) );
  XNOR U4915 ( .A(n1814), .B(n1824), .Z(n1815) );
  XNOR U4916 ( .A(n1816), .B(n1815), .Z(n1823) );
  NAND U4917 ( .A(n1818), .B(n1817), .Z(n1819) );
  XNOR U4918 ( .A(n1820), .B(n1819), .Z(n1830) );
  XNOR U4919 ( .A(n1821), .B(n1830), .Z(n1822) );
  XOR U4920 ( .A(n1823), .B(n1822), .Z(n1833) );
  XNOR U4921 ( .A(n1852), .B(n1833), .Z(z[81]) );
  XNOR U4922 ( .A(n1825), .B(n1824), .Z(z[82]) );
  ANDN U4923 ( .B(n1827), .A(n1826), .Z(n1832) );
  NANDN U4924 ( .A(n1829), .B(n1828), .Z(n1842) );
  XNOR U4925 ( .A(n1830), .B(n1842), .Z(n1831) );
  XOR U4926 ( .A(n1832), .B(n1831), .Z(n1851) );
  XOR U4927 ( .A(n1834), .B(n1833), .Z(n1835) );
  XOR U4928 ( .A(n1851), .B(n1835), .Z(z[83]) );
  XOR U4929 ( .A(n1836), .B(z[82]), .Z(z[84]) );
  XNOR U4930 ( .A(n1838), .B(n1837), .Z(n1840) );
  NAND U4931 ( .A(n1840), .B(n1839), .Z(n1841) );
  XOR U4932 ( .A(n1842), .B(n1841), .Z(n1843) );
  XNOR U4933 ( .A(n1844), .B(n1843), .Z(n1850) );
  NAND U4934 ( .A(x[80]), .B(n1845), .Z(n1846) );
  XNOR U4935 ( .A(n1847), .B(n1846), .Z(n1854) );
  XNOR U4936 ( .A(n1848), .B(n1854), .Z(n1849) );
  XOR U4937 ( .A(n1850), .B(n1849), .Z(z[85]) );
  XNOR U4938 ( .A(n1852), .B(n1851), .Z(z[86]) );
  XNOR U4939 ( .A(n1854), .B(n1853), .Z(n1855) );
  XNOR U4940 ( .A(z[81]), .B(n1855), .Z(z[87]) );
  XOR U4941 ( .A(x[88]), .B(x[94]), .Z(n1856) );
  XOR U4942 ( .A(x[93]), .B(n1856), .Z(n1963) );
  IV U4943 ( .A(n1963), .Z(n1858) );
  IV U4944 ( .A(x[89]), .Z(n1962) );
  NAND U4945 ( .A(n1858), .B(n1962), .Z(n1865) );
  XOR U4946 ( .A(x[91]), .B(x[89]), .Z(n1861) );
  XNOR U4947 ( .A(x[90]), .B(n1856), .Z(n1857) );
  XNOR U4948 ( .A(n1861), .B(n1857), .Z(n1920) );
  XNOR U4949 ( .A(n1858), .B(n1920), .Z(n1919) );
  IV U4950 ( .A(x[95]), .Z(n1859) );
  XNOR U4951 ( .A(x[89]), .B(n1859), .Z(n1953) );
  NAND U4952 ( .A(n1919), .B(n1953), .Z(n1868) );
  XNOR U4953 ( .A(n1858), .B(n1859), .Z(n1951) );
  XOR U4954 ( .A(n1920), .B(n1951), .Z(n1876) );
  XOR U4955 ( .A(n1868), .B(n1876), .Z(n1863) );
  XNOR U4956 ( .A(x[88]), .B(n1920), .Z(n1895) );
  XOR U4957 ( .A(x[92]), .B(n1859), .Z(n1860) );
  IV U4958 ( .A(n1860), .Z(n1924) );
  NANDN U4959 ( .A(n1895), .B(n1924), .Z(n1867) );
  XOR U4960 ( .A(n1861), .B(n1860), .Z(n1913) );
  XOR U4961 ( .A(n1919), .B(n1913), .Z(n1911) );
  XOR U4962 ( .A(x[90]), .B(x[92]), .Z(n1926) );
  NANDN U4963 ( .A(n1911), .B(n1926), .Z(n1862) );
  XNOR U4964 ( .A(n1867), .B(n1862), .Z(n1872) );
  XOR U4965 ( .A(n1863), .B(n1872), .Z(n1864) );
  XOR U4966 ( .A(n1865), .B(n1864), .Z(n1906) );
  IV U4967 ( .A(n1906), .Z(n1900) );
  ANDN U4968 ( .B(n1951), .A(n1920), .Z(n1870) );
  XNOR U4969 ( .A(x[88]), .B(n1913), .Z(n1914) );
  XNOR U4970 ( .A(n1963), .B(n1914), .Z(n1916) );
  XOR U4971 ( .A(x[90]), .B(x[95]), .Z(n1941) );
  NANDN U4972 ( .A(n1916), .B(n1941), .Z(n1866) );
  XNOR U4973 ( .A(n1867), .B(n1866), .Z(n1883) );
  XNOR U4974 ( .A(n1868), .B(n1883), .Z(n1869) );
  XOR U4975 ( .A(n1870), .B(n1869), .Z(n1896) );
  NAND U4976 ( .A(n1900), .B(n1896), .Z(n1890) );
  IV U4977 ( .A(n1896), .Z(n1897) );
  XOR U4978 ( .A(n1906), .B(n1897), .Z(n1888) );
  XOR U4979 ( .A(x[90]), .B(x[89]), .Z(n1871) );
  XNOR U4980 ( .A(n1951), .B(n1871), .Z(n1923) );
  NAND U4981 ( .A(n1923), .B(n1914), .Z(n1878) );
  XNOR U4982 ( .A(x[92]), .B(n1963), .Z(n1934) );
  XOR U4983 ( .A(n1924), .B(n1871), .Z(n1929) );
  NANDN U4984 ( .A(n1913), .B(n1929), .Z(n1879) );
  XOR U4985 ( .A(n1934), .B(n1879), .Z(n1874) );
  XOR U4986 ( .A(x[88]), .B(n1872), .Z(n1873) );
  XNOR U4987 ( .A(n1874), .B(n1873), .Z(n1875) );
  XOR U4988 ( .A(n1876), .B(n1875), .Z(n1877) );
  XOR U4989 ( .A(n1878), .B(n1877), .Z(n1908) );
  IV U4990 ( .A(n1908), .Z(n1903) );
  AND U4991 ( .A(n1900), .B(n1903), .Z(n1886) );
  ANDN U4992 ( .B(x[88]), .A(n1934), .Z(n1885) );
  XNOR U4993 ( .A(n1923), .B(n1879), .Z(n1881) );
  XNOR U4994 ( .A(x[89]), .B(n1914), .Z(n1880) );
  XNOR U4995 ( .A(n1881), .B(n1880), .Z(n1882) );
  XOR U4996 ( .A(n1883), .B(n1882), .Z(n1884) );
  XOR U4997 ( .A(n1885), .B(n1884), .Z(n1898) );
  IV U4998 ( .A(n1898), .Z(n1904) );
  XNOR U4999 ( .A(n1886), .B(n1904), .Z(n1887) );
  NAND U5000 ( .A(n1888), .B(n1887), .Z(n1889) );
  NAND U5001 ( .A(n1890), .B(n1889), .Z(n1970) );
  NAND U5002 ( .A(n1904), .B(n1897), .Z(n1891) );
  NAND U5003 ( .A(n1903), .B(n1891), .Z(n1894) );
  XOR U5004 ( .A(n1897), .B(n1900), .Z(n1892) );
  NAND U5005 ( .A(n1898), .B(n1892), .Z(n1893) );
  AND U5006 ( .A(n1894), .B(n1893), .Z(n1952) );
  XNOR U5007 ( .A(n1970), .B(n1952), .Z(n1925) );
  OR U5008 ( .A(n1925), .B(n1895), .Z(n1918) );
  NAND U5009 ( .A(n1906), .B(n1896), .Z(n1902) );
  AND U5010 ( .A(n1898), .B(n1897), .Z(n1905) );
  XNOR U5011 ( .A(n1905), .B(n1903), .Z(n1899) );
  NAND U5012 ( .A(n1900), .B(n1899), .Z(n1901) );
  AND U5013 ( .A(n1902), .B(n1901), .Z(n1922) );
  NAND U5014 ( .A(n1904), .B(n1903), .Z(n1910) );
  XNOR U5015 ( .A(n1906), .B(n1905), .Z(n1907) );
  NAND U5016 ( .A(n1908), .B(n1907), .Z(n1909) );
  NAND U5017 ( .A(n1910), .B(n1909), .Z(n1964) );
  XNOR U5018 ( .A(n1922), .B(n1964), .Z(n1940) );
  XOR U5019 ( .A(n1940), .B(n1925), .Z(n1927) );
  OR U5020 ( .A(n1927), .B(n1911), .Z(n1912) );
  XNOR U5021 ( .A(n1918), .B(n1912), .Z(n1944) );
  XOR U5022 ( .A(n1922), .B(n1970), .Z(n1930) );
  OR U5023 ( .A(n1913), .B(n1930), .Z(n1972) );
  NANDN U5024 ( .A(n1922), .B(n1914), .Z(n1915) );
  XNOR U5025 ( .A(n1972), .B(n1915), .Z(n1950) );
  XOR U5026 ( .A(n1944), .B(n1950), .Z(n1933) );
  NANDN U5027 ( .A(n1916), .B(n1940), .Z(n1917) );
  XNOR U5028 ( .A(n1918), .B(n1917), .Z(n1978) );
  XNOR U5029 ( .A(n1964), .B(n1952), .Z(n1954) );
  NANDN U5030 ( .A(n1954), .B(n1919), .Z(n1936) );
  NAND U5031 ( .A(n1920), .B(n1952), .Z(n1921) );
  XNOR U5032 ( .A(n1936), .B(n1921), .Z(n1969) );
  XOR U5033 ( .A(n1978), .B(n1969), .Z(n1961) );
  XNOR U5034 ( .A(n1933), .B(n1961), .Z(z[88]) );
  ANDN U5035 ( .B(n1923), .A(n1922), .Z(n1932) );
  NANDN U5036 ( .A(n1925), .B(n1924), .Z(n1943) );
  NANDN U5037 ( .A(n1927), .B(n1926), .Z(n1928) );
  XNOR U5038 ( .A(n1943), .B(n1928), .Z(n1973) );
  NANDN U5039 ( .A(n1930), .B(n1929), .Z(n1937) );
  XNOR U5040 ( .A(n1973), .B(n1937), .Z(n1931) );
  XOR U5041 ( .A(n1932), .B(n1931), .Z(n1959) );
  XOR U5042 ( .A(n1959), .B(n1933), .Z(n1977) );
  ANDN U5043 ( .B(n1970), .A(n1934), .Z(n1939) );
  NAND U5044 ( .A(n1963), .B(n1964), .Z(n1935) );
  XNOR U5045 ( .A(n1936), .B(n1935), .Z(n1949) );
  XNOR U5046 ( .A(n1937), .B(n1949), .Z(n1938) );
  XNOR U5047 ( .A(n1939), .B(n1938), .Z(n1946) );
  NAND U5048 ( .A(n1941), .B(n1940), .Z(n1942) );
  XNOR U5049 ( .A(n1943), .B(n1942), .Z(n1955) );
  XNOR U5050 ( .A(n1944), .B(n1955), .Z(n1945) );
  XOR U5051 ( .A(n1946), .B(n1945), .Z(n1958) );
  XNOR U5052 ( .A(n1977), .B(n1958), .Z(z[89]) );
  XNOR U5053 ( .A(n1948), .B(n1947), .Z(z[8]) );
  XNOR U5054 ( .A(n1950), .B(n1949), .Z(z[90]) );
  ANDN U5055 ( .B(n1952), .A(n1951), .Z(n1957) );
  NANDN U5056 ( .A(n1954), .B(n1953), .Z(n1967) );
  XNOR U5057 ( .A(n1955), .B(n1967), .Z(n1956) );
  XOR U5058 ( .A(n1957), .B(n1956), .Z(n1976) );
  XOR U5059 ( .A(n1959), .B(n1958), .Z(n1960) );
  XOR U5060 ( .A(n1976), .B(n1960), .Z(z[91]) );
  XOR U5061 ( .A(n1961), .B(z[90]), .Z(z[92]) );
  XNOR U5062 ( .A(n1963), .B(n1962), .Z(n1965) );
  NAND U5063 ( .A(n1965), .B(n1964), .Z(n1966) );
  XOR U5064 ( .A(n1967), .B(n1966), .Z(n1968) );
  XNOR U5065 ( .A(n1969), .B(n1968), .Z(n1975) );
  NAND U5066 ( .A(x[88]), .B(n1970), .Z(n1971) );
  XNOR U5067 ( .A(n1972), .B(n1971), .Z(n1979) );
  XNOR U5068 ( .A(n1973), .B(n1979), .Z(n1974) );
  XOR U5069 ( .A(n1975), .B(n1974), .Z(z[93]) );
  XNOR U5070 ( .A(n1977), .B(n1976), .Z(z[94]) );
  XNOR U5071 ( .A(n1979), .B(n1978), .Z(n1980) );
  XNOR U5072 ( .A(z[89]), .B(n1980), .Z(z[95]) );
  XNOR U5073 ( .A(n1982), .B(n1981), .Z(z[96]) );
  XOR U5074 ( .A(n1984), .B(n1983), .Z(n1985) );
  XOR U5075 ( .A(n1986), .B(n1985), .Z(z[99]) );
endmodule


module SubBytes_3 ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986;

  XNOR U2962 ( .A(n328), .B(n339), .Z(n341) );
  XNOR U2963 ( .A(n170), .B(n162), .Z(n143) );
  XOR U2964 ( .A(n493), .B(n494), .Z(n646) );
  IV U2965 ( .A(x[1]), .Z(n1447) );
  XOR U2966 ( .A(x[0]), .B(x[6]), .Z(n2) );
  XOR U2967 ( .A(x[5]), .B(n2), .Z(n1446) );
  IV U2968 ( .A(n1446), .Z(n3) );
  AND U2969 ( .A(n1447), .B(n3), .Z(n10) );
  XNOR U2970 ( .A(x[3]), .B(n1447), .Z(n6) );
  XNOR U2971 ( .A(x[2]), .B(n6), .Z(n1) );
  XNOR U2972 ( .A(n2), .B(n1), .Z(n66) );
  IV U2973 ( .A(n66), .Z(n12) );
  XNOR U2974 ( .A(n12), .B(n1446), .Z(n65) );
  IV U2975 ( .A(x[7]), .Z(n4) );
  XNOR U2976 ( .A(x[1]), .B(n4), .Z(n1085) );
  NAND U2977 ( .A(n65), .B(n1085), .Z(n15) );
  XNOR U2978 ( .A(n4), .B(n3), .Z(n11) );
  IV U2979 ( .A(n11), .Z(n1083) );
  XOR U2980 ( .A(n66), .B(n1083), .Z(n31) );
  XNOR U2981 ( .A(n15), .B(n31), .Z(n8) );
  XOR U2982 ( .A(x[0]), .B(n12), .Z(n41) );
  XOR U2983 ( .A(x[4]), .B(n4), .Z(n5) );
  IV U2984 ( .A(n5), .Z(n790) );
  NANDN U2985 ( .A(n41), .B(n790), .Z(n14) );
  XNOR U2986 ( .A(n6), .B(n5), .Z(n59) );
  XNOR U2987 ( .A(n65), .B(n59), .Z(n57) );
  XOR U2988 ( .A(x[2]), .B(x[4]), .Z(n792) );
  NANDN U2989 ( .A(n57), .B(n792), .Z(n7) );
  XOR U2990 ( .A(n14), .B(n7), .Z(n33) );
  XNOR U2991 ( .A(n8), .B(n33), .Z(n9) );
  XOR U2992 ( .A(n10), .B(n9), .Z(n46) );
  IV U2993 ( .A(n46), .Z(n52) );
  AND U2994 ( .A(n12), .B(n11), .Z(n17) );
  XOR U2995 ( .A(x[0]), .B(n59), .Z(n60) );
  XNOR U2996 ( .A(n1446), .B(n60), .Z(n62) );
  XOR U2997 ( .A(x[2]), .B(x[7]), .Z(n807) );
  NANDN U2998 ( .A(n62), .B(n807), .Z(n13) );
  XNOR U2999 ( .A(n14), .B(n13), .Z(n22) );
  XNOR U3000 ( .A(n15), .B(n22), .Z(n16) );
  XOR U3001 ( .A(n17), .B(n16), .Z(n42) );
  XNOR U3002 ( .A(x[4]), .B(n1446), .Z(n800) );
  ANDN U3003 ( .B(x[0]), .A(n800), .Z(n24) );
  XOR U3004 ( .A(x[2]), .B(x[1]), .Z(n18) );
  XOR U3005 ( .A(n1083), .B(n18), .Z(n789) );
  XOR U3006 ( .A(n790), .B(n18), .Z(n795) );
  NAND U3007 ( .A(n59), .B(n795), .Z(n26) );
  XNOR U3008 ( .A(n789), .B(n26), .Z(n20) );
  XNOR U3009 ( .A(x[1]), .B(n60), .Z(n19) );
  XNOR U3010 ( .A(n20), .B(n19), .Z(n21) );
  XOR U3011 ( .A(n22), .B(n21), .Z(n23) );
  XOR U3012 ( .A(n24), .B(n23), .Z(n44) );
  NAND U3013 ( .A(n42), .B(n44), .Z(n25) );
  NAND U3014 ( .A(n52), .B(n25), .Z(n36) );
  IV U3015 ( .A(n42), .Z(n43) );
  IV U3016 ( .A(n44), .Z(n50) );
  XOR U3017 ( .A(n26), .B(n800), .Z(n29) );
  AND U3018 ( .A(n789), .B(n60), .Z(n27) );
  XNOR U3019 ( .A(x[0]), .B(n27), .Z(n28) );
  XNOR U3020 ( .A(n29), .B(n28), .Z(n30) );
  XNOR U3021 ( .A(n31), .B(n30), .Z(n32) );
  XNOR U3022 ( .A(n33), .B(n32), .Z(n54) );
  IV U3023 ( .A(n54), .Z(n49) );
  XOR U3024 ( .A(n50), .B(n49), .Z(n34) );
  NAND U3025 ( .A(n43), .B(n34), .Z(n35) );
  AND U3026 ( .A(n36), .B(n35), .Z(n1454) );
  NAND U3027 ( .A(n50), .B(n43), .Z(n37) );
  NAND U3028 ( .A(n49), .B(n37), .Z(n40) );
  XOR U3029 ( .A(n43), .B(n46), .Z(n38) );
  NAND U3030 ( .A(n44), .B(n38), .Z(n39) );
  AND U3031 ( .A(n40), .B(n39), .Z(n1084) );
  XNOR U3032 ( .A(n1454), .B(n1084), .Z(n791) );
  OR U3033 ( .A(n791), .B(n41), .Z(n64) );
  NAND U3034 ( .A(n52), .B(n42), .Z(n48) );
  AND U3035 ( .A(n44), .B(n43), .Z(n51) );
  XNOR U3036 ( .A(n49), .B(n51), .Z(n45) );
  NAND U3037 ( .A(n46), .B(n45), .Z(n47) );
  AND U3038 ( .A(n48), .B(n47), .Z(n788) );
  NAND U3039 ( .A(n50), .B(n49), .Z(n56) );
  XNOR U3040 ( .A(n52), .B(n51), .Z(n53) );
  NAND U3041 ( .A(n54), .B(n53), .Z(n55) );
  NAND U3042 ( .A(n56), .B(n55), .Z(n1448) );
  XNOR U3043 ( .A(n788), .B(n1448), .Z(n806) );
  XOR U3044 ( .A(n806), .B(n791), .Z(n793) );
  OR U3045 ( .A(n793), .B(n57), .Z(n58) );
  XNOR U3046 ( .A(n64), .B(n58), .Z(n810) );
  XOR U3047 ( .A(n788), .B(n1454), .Z(n796) );
  NANDN U3048 ( .A(n796), .B(n59), .Z(n1456) );
  NANDN U3049 ( .A(n788), .B(n60), .Z(n61) );
  XNOR U3050 ( .A(n1456), .B(n61), .Z(n953) );
  XOR U3051 ( .A(n810), .B(n953), .Z(n799) );
  NANDN U3052 ( .A(n62), .B(n806), .Z(n63) );
  XNOR U3053 ( .A(n64), .B(n63), .Z(n1730) );
  XNOR U3054 ( .A(n1448), .B(n1084), .Z(n1086) );
  NANDN U3055 ( .A(n1086), .B(n65), .Z(n802) );
  NAND U3056 ( .A(n66), .B(n1084), .Z(n67) );
  XNOR U3057 ( .A(n802), .B(n67), .Z(n1453) );
  XOR U3058 ( .A(n1730), .B(n1453), .Z(n1309) );
  XNOR U3059 ( .A(n799), .B(n1309), .Z(z[0]) );
  XOR U3060 ( .A(x[96]), .B(x[102]), .Z(n68) );
  XOR U3061 ( .A(x[101]), .B(n68), .Z(n135) );
  XOR U3062 ( .A(x[100]), .B(n135), .Z(n171) );
  AND U3063 ( .A(x[96]), .B(n171), .Z(n78) );
  XOR U3064 ( .A(x[97]), .B(x[99]), .Z(n71) );
  XNOR U3065 ( .A(n68), .B(x[98]), .Z(n69) );
  XOR U3066 ( .A(n71), .B(n69), .Z(n129) );
  XOR U3067 ( .A(x[96]), .B(n129), .Z(n128) );
  XNOR U3068 ( .A(x[103]), .B(x[100]), .Z(n70) );
  IV U3069 ( .A(n70), .Z(n142) );
  NANDN U3070 ( .A(n128), .B(n142), .Z(n80) );
  IV U3071 ( .A(n135), .Z(n91) );
  XNOR U3072 ( .A(n71), .B(n70), .Z(n123) );
  XOR U3073 ( .A(x[96]), .B(n123), .Z(n124) );
  XOR U3074 ( .A(n91), .B(n124), .Z(n126) );
  XOR U3075 ( .A(x[98]), .B(x[103]), .Z(n164) );
  NANDN U3076 ( .A(n126), .B(n164), .Z(n72) );
  XNOR U3077 ( .A(n80), .B(n72), .Z(n87) );
  XNOR U3078 ( .A(n135), .B(x[103]), .Z(n161) );
  XOR U3079 ( .A(x[97]), .B(x[98]), .Z(n73) );
  XNOR U3080 ( .A(n161), .B(n73), .Z(n151) );
  XOR U3081 ( .A(n142), .B(n73), .Z(n152) );
  NAND U3082 ( .A(n123), .B(n152), .Z(n81) );
  XNOR U3083 ( .A(n151), .B(n81), .Z(n75) );
  XNOR U3084 ( .A(x[97]), .B(n124), .Z(n74) );
  XNOR U3085 ( .A(n75), .B(n74), .Z(n76) );
  XOR U3086 ( .A(n87), .B(n76), .Z(n77) );
  XOR U3087 ( .A(n78), .B(n77), .Z(n115) );
  IV U3088 ( .A(n115), .Z(n108) );
  XNOR U3089 ( .A(n129), .B(n135), .Z(n105) );
  XNOR U3090 ( .A(n105), .B(n123), .Z(n158) );
  XNOR U3091 ( .A(x[98]), .B(x[100]), .Z(n144) );
  OR U3092 ( .A(n158), .B(n144), .Z(n79) );
  XOR U3093 ( .A(n80), .B(n79), .Z(n94) );
  XNOR U3094 ( .A(n129), .B(n161), .Z(n92) );
  XNOR U3095 ( .A(n81), .B(n171), .Z(n84) );
  AND U3096 ( .A(n151), .B(n124), .Z(n82) );
  XNOR U3097 ( .A(x[96]), .B(n82), .Z(n83) );
  XNOR U3098 ( .A(n84), .B(n83), .Z(n85) );
  XOR U3099 ( .A(n92), .B(n85), .Z(n86) );
  XOR U3100 ( .A(n94), .B(n86), .Z(n118) );
  AND U3101 ( .A(n129), .B(n161), .Z(n89) );
  IV U3102 ( .A(x[97]), .Z(n136) );
  XNOR U3103 ( .A(n136), .B(x[103]), .Z(n133) );
  NAND U3104 ( .A(n105), .B(n133), .Z(n93) );
  XNOR U3105 ( .A(n93), .B(n87), .Z(n88) );
  XOR U3106 ( .A(n89), .B(n88), .Z(n107) );
  NAND U3107 ( .A(n118), .B(n107), .Z(n90) );
  NAND U3108 ( .A(n108), .B(n90), .Z(n99) );
  IV U3109 ( .A(n118), .Z(n102) );
  NAND U3110 ( .A(n91), .B(n136), .Z(n97) );
  XOR U3111 ( .A(n93), .B(n92), .Z(n95) );
  XNOR U3112 ( .A(n95), .B(n94), .Z(n96) );
  XOR U3113 ( .A(n97), .B(n96), .Z(n114) );
  IV U3114 ( .A(n107), .Z(n116) );
  XOR U3115 ( .A(n114), .B(n116), .Z(n111) );
  NAND U3116 ( .A(n102), .B(n111), .Z(n98) );
  AND U3117 ( .A(n99), .B(n98), .Z(n127) );
  NAND U3118 ( .A(n118), .B(n108), .Z(n104) );
  AND U3119 ( .A(n115), .B(n116), .Z(n100) );
  XNOR U3120 ( .A(n114), .B(n100), .Z(n101) );
  NAND U3121 ( .A(n102), .B(n101), .Z(n103) );
  AND U3122 ( .A(n104), .B(n103), .Z(n138) );
  XNOR U3123 ( .A(n127), .B(n138), .Z(n134) );
  NANDN U3124 ( .A(n134), .B(n105), .Z(n131) );
  NANDN U3125 ( .A(n138), .B(n135), .Z(n106) );
  XNOR U3126 ( .A(n131), .B(n106), .Z(n173) );
  IV U3127 ( .A(n114), .Z(n120) );
  NAND U3128 ( .A(n120), .B(n107), .Z(n113) );
  AND U3129 ( .A(n120), .B(n118), .Z(n109) );
  XNOR U3130 ( .A(n109), .B(n108), .Z(n110) );
  NAND U3131 ( .A(n111), .B(n110), .Z(n112) );
  NAND U3132 ( .A(n113), .B(n112), .Z(n170) );
  NAND U3133 ( .A(n114), .B(n116), .Z(n122) );
  NAND U3134 ( .A(n116), .B(n115), .Z(n117) );
  XNOR U3135 ( .A(n118), .B(n117), .Z(n119) );
  NAND U3136 ( .A(n120), .B(n119), .Z(n121) );
  NAND U3137 ( .A(n122), .B(n121), .Z(n150) );
  XOR U3138 ( .A(n170), .B(n150), .Z(n153) );
  NANDN U3139 ( .A(n153), .B(n123), .Z(n147) );
  NANDN U3140 ( .A(n150), .B(n124), .Z(n125) );
  XNOR U3141 ( .A(n147), .B(n125), .Z(n160) );
  XNOR U3142 ( .A(n173), .B(n160), .Z(z[98]) );
  XOR U3143 ( .A(n150), .B(n138), .Z(n163) );
  ANDN U3144 ( .B(n163), .A(n126), .Z(n184) );
  IV U3145 ( .A(n127), .Z(n162) );
  OR U3146 ( .A(n143), .B(n128), .Z(n182) );
  NANDN U3147 ( .A(n129), .B(n162), .Z(n130) );
  XNOR U3148 ( .A(n131), .B(n130), .Z(n141) );
  XNOR U3149 ( .A(n182), .B(n141), .Z(n132) );
  XOR U3150 ( .A(n184), .B(n132), .Z(n1982) );
  XNOR U3151 ( .A(n1982), .B(z[98]), .Z(z[100]) );
  NANDN U3152 ( .A(n134), .B(n133), .Z(n167) );
  XNOR U3153 ( .A(n136), .B(n135), .Z(n137) );
  NANDN U3154 ( .A(n138), .B(n137), .Z(n139) );
  XOR U3155 ( .A(n167), .B(n139), .Z(n140) );
  XNOR U3156 ( .A(n141), .B(n140), .Z(n149) );
  NANDN U3157 ( .A(n143), .B(n142), .Z(n166) );
  XNOR U3158 ( .A(n143), .B(n163), .Z(n157) );
  NANDN U3159 ( .A(n144), .B(n157), .Z(n145) );
  XNOR U3160 ( .A(n166), .B(n145), .Z(n154) );
  NAND U3161 ( .A(n170), .B(x[96]), .Z(n146) );
  XNOR U3162 ( .A(n147), .B(n146), .Z(n181) );
  XNOR U3163 ( .A(n154), .B(n181), .Z(n148) );
  XOR U3164 ( .A(n149), .B(n148), .Z(z[101]) );
  ANDN U3165 ( .B(n151), .A(n150), .Z(n156) );
  NANDN U3166 ( .A(n153), .B(n152), .Z(n172) );
  XNOR U3167 ( .A(n172), .B(n154), .Z(n155) );
  XOR U3168 ( .A(n156), .B(n155), .Z(n1983) );
  NANDN U3169 ( .A(n158), .B(n157), .Z(n159) );
  XOR U3170 ( .A(n182), .B(n159), .Z(n176) );
  XOR U3171 ( .A(n176), .B(n160), .Z(n1981) );
  XNOR U3172 ( .A(n1983), .B(n1981), .Z(n180) );
  ANDN U3173 ( .B(n162), .A(n161), .Z(n169) );
  NAND U3174 ( .A(n164), .B(n163), .Z(n165) );
  XNOR U3175 ( .A(n166), .B(n165), .Z(n177) );
  XNOR U3176 ( .A(n177), .B(n167), .Z(n168) );
  XOR U3177 ( .A(n169), .B(n168), .Z(n1986) );
  XNOR U3178 ( .A(n180), .B(n1986), .Z(z[102]) );
  AND U3179 ( .A(n171), .B(n170), .Z(n175) );
  XNOR U3180 ( .A(n173), .B(n172), .Z(n174) );
  XNOR U3181 ( .A(n175), .B(n174), .Z(n179) );
  XOR U3182 ( .A(n177), .B(n176), .Z(n178) );
  XOR U3183 ( .A(n179), .B(n178), .Z(n1984) );
  XNOR U3184 ( .A(n1984), .B(n180), .Z(z[97]) );
  XNOR U3185 ( .A(n182), .B(n181), .Z(n183) );
  XNOR U3186 ( .A(n184), .B(n183), .Z(n185) );
  XOR U3187 ( .A(n185), .B(z[97]), .Z(z[103]) );
  IV U3188 ( .A(x[105]), .Z(n292) );
  XOR U3189 ( .A(x[104]), .B(x[110]), .Z(n187) );
  XOR U3190 ( .A(x[109]), .B(n187), .Z(n291) );
  IV U3191 ( .A(n291), .Z(n188) );
  AND U3192 ( .A(n292), .B(n188), .Z(n195) );
  XNOR U3193 ( .A(x[107]), .B(n292), .Z(n191) );
  XNOR U3194 ( .A(x[106]), .B(n191), .Z(n186) );
  XNOR U3195 ( .A(n187), .B(n186), .Z(n251) );
  IV U3196 ( .A(n251), .Z(n197) );
  XNOR U3197 ( .A(n197), .B(n291), .Z(n250) );
  IV U3198 ( .A(x[111]), .Z(n189) );
  XNOR U3199 ( .A(x[105]), .B(n189), .Z(n282) );
  NAND U3200 ( .A(n250), .B(n282), .Z(n200) );
  XNOR U3201 ( .A(n189), .B(n188), .Z(n196) );
  IV U3202 ( .A(n196), .Z(n280) );
  XOR U3203 ( .A(n251), .B(n280), .Z(n216) );
  XNOR U3204 ( .A(n200), .B(n216), .Z(n193) );
  XOR U3205 ( .A(x[104]), .B(n197), .Z(n226) );
  XOR U3206 ( .A(x[108]), .B(n189), .Z(n190) );
  IV U3207 ( .A(n190), .Z(n255) );
  NANDN U3208 ( .A(n226), .B(n255), .Z(n199) );
  XNOR U3209 ( .A(n191), .B(n190), .Z(n244) );
  XNOR U3210 ( .A(n250), .B(n244), .Z(n242) );
  XOR U3211 ( .A(x[106]), .B(x[108]), .Z(n257) );
  NANDN U3212 ( .A(n242), .B(n257), .Z(n192) );
  XOR U3213 ( .A(n199), .B(n192), .Z(n218) );
  XNOR U3214 ( .A(n193), .B(n218), .Z(n194) );
  XOR U3215 ( .A(n195), .B(n194), .Z(n231) );
  IV U3216 ( .A(n231), .Z(n237) );
  AND U3217 ( .A(n197), .B(n196), .Z(n202) );
  XOR U3218 ( .A(x[104]), .B(n244), .Z(n245) );
  XNOR U3219 ( .A(n291), .B(n245), .Z(n247) );
  XOR U3220 ( .A(x[106]), .B(x[111]), .Z(n272) );
  NANDN U3221 ( .A(n247), .B(n272), .Z(n198) );
  XNOR U3222 ( .A(n199), .B(n198), .Z(n207) );
  XNOR U3223 ( .A(n200), .B(n207), .Z(n201) );
  XOR U3224 ( .A(n202), .B(n201), .Z(n227) );
  XNOR U3225 ( .A(x[108]), .B(n291), .Z(n265) );
  ANDN U3226 ( .B(x[104]), .A(n265), .Z(n209) );
  XOR U3227 ( .A(x[106]), .B(x[105]), .Z(n203) );
  XOR U3228 ( .A(n280), .B(n203), .Z(n254) );
  XOR U3229 ( .A(n255), .B(n203), .Z(n260) );
  NAND U3230 ( .A(n244), .B(n260), .Z(n211) );
  XNOR U3231 ( .A(n254), .B(n211), .Z(n205) );
  XNOR U3232 ( .A(x[105]), .B(n245), .Z(n204) );
  XNOR U3233 ( .A(n205), .B(n204), .Z(n206) );
  XOR U3234 ( .A(n207), .B(n206), .Z(n208) );
  XOR U3235 ( .A(n209), .B(n208), .Z(n229) );
  NAND U3236 ( .A(n227), .B(n229), .Z(n210) );
  NAND U3237 ( .A(n237), .B(n210), .Z(n221) );
  IV U3238 ( .A(n227), .Z(n228) );
  IV U3239 ( .A(n229), .Z(n235) );
  XOR U3240 ( .A(n211), .B(n265), .Z(n214) );
  AND U3241 ( .A(n254), .B(n245), .Z(n212) );
  XNOR U3242 ( .A(x[104]), .B(n212), .Z(n213) );
  XNOR U3243 ( .A(n214), .B(n213), .Z(n215) );
  XNOR U3244 ( .A(n216), .B(n215), .Z(n217) );
  XNOR U3245 ( .A(n218), .B(n217), .Z(n239) );
  IV U3246 ( .A(n239), .Z(n234) );
  XOR U3247 ( .A(n235), .B(n234), .Z(n219) );
  NAND U3248 ( .A(n228), .B(n219), .Z(n220) );
  AND U3249 ( .A(n221), .B(n220), .Z(n299) );
  NAND U3250 ( .A(n235), .B(n228), .Z(n222) );
  NAND U3251 ( .A(n234), .B(n222), .Z(n225) );
  XOR U3252 ( .A(n228), .B(n231), .Z(n223) );
  NAND U3253 ( .A(n229), .B(n223), .Z(n224) );
  AND U3254 ( .A(n225), .B(n224), .Z(n281) );
  XNOR U3255 ( .A(n299), .B(n281), .Z(n256) );
  OR U3256 ( .A(n256), .B(n226), .Z(n249) );
  NAND U3257 ( .A(n237), .B(n227), .Z(n233) );
  AND U3258 ( .A(n229), .B(n228), .Z(n236) );
  XNOR U3259 ( .A(n234), .B(n236), .Z(n230) );
  NAND U3260 ( .A(n231), .B(n230), .Z(n232) );
  AND U3261 ( .A(n233), .B(n232), .Z(n253) );
  NAND U3262 ( .A(n235), .B(n234), .Z(n241) );
  XNOR U3263 ( .A(n237), .B(n236), .Z(n238) );
  NAND U3264 ( .A(n239), .B(n238), .Z(n240) );
  NAND U3265 ( .A(n241), .B(n240), .Z(n293) );
  XNOR U3266 ( .A(n253), .B(n293), .Z(n271) );
  XOR U3267 ( .A(n271), .B(n256), .Z(n258) );
  OR U3268 ( .A(n258), .B(n242), .Z(n243) );
  XNOR U3269 ( .A(n249), .B(n243), .Z(n275) );
  XOR U3270 ( .A(n253), .B(n299), .Z(n261) );
  NANDN U3271 ( .A(n261), .B(n244), .Z(n301) );
  NANDN U3272 ( .A(n253), .B(n245), .Z(n246) );
  XNOR U3273 ( .A(n301), .B(n246), .Z(n279) );
  XOR U3274 ( .A(n275), .B(n279), .Z(n264) );
  NANDN U3275 ( .A(n247), .B(n271), .Z(n248) );
  XNOR U3276 ( .A(n249), .B(n248), .Z(n366) );
  XNOR U3277 ( .A(n293), .B(n281), .Z(n283) );
  NANDN U3278 ( .A(n283), .B(n250), .Z(n267) );
  NAND U3279 ( .A(n251), .B(n281), .Z(n252) );
  XNOR U3280 ( .A(n267), .B(n252), .Z(n298) );
  XOR U3281 ( .A(n366), .B(n298), .Z(n290) );
  XNOR U3282 ( .A(n264), .B(n290), .Z(z[104]) );
  ANDN U3283 ( .B(n254), .A(n253), .Z(n263) );
  NANDN U3284 ( .A(n256), .B(n255), .Z(n274) );
  NANDN U3285 ( .A(n258), .B(n257), .Z(n259) );
  XNOR U3286 ( .A(n274), .B(n259), .Z(n302) );
  NANDN U3287 ( .A(n261), .B(n260), .Z(n268) );
  XNOR U3288 ( .A(n302), .B(n268), .Z(n262) );
  XOR U3289 ( .A(n263), .B(n262), .Z(n288) );
  XOR U3290 ( .A(n288), .B(n264), .Z(n365) );
  ANDN U3291 ( .B(n299), .A(n265), .Z(n270) );
  NAND U3292 ( .A(n291), .B(n293), .Z(n266) );
  XNOR U3293 ( .A(n267), .B(n266), .Z(n278) );
  XNOR U3294 ( .A(n268), .B(n278), .Z(n269) );
  XNOR U3295 ( .A(n270), .B(n269), .Z(n277) );
  NAND U3296 ( .A(n272), .B(n271), .Z(n273) );
  XNOR U3297 ( .A(n274), .B(n273), .Z(n284) );
  XNOR U3298 ( .A(n275), .B(n284), .Z(n276) );
  XOR U3299 ( .A(n277), .B(n276), .Z(n287) );
  XNOR U3300 ( .A(n365), .B(n287), .Z(z[105]) );
  XNOR U3301 ( .A(n279), .B(n278), .Z(z[106]) );
  AND U3302 ( .A(n281), .B(n280), .Z(n286) );
  NANDN U3303 ( .A(n283), .B(n282), .Z(n296) );
  XNOR U3304 ( .A(n284), .B(n296), .Z(n285) );
  XOR U3305 ( .A(n286), .B(n285), .Z(n364) );
  XOR U3306 ( .A(n288), .B(n287), .Z(n289) );
  XOR U3307 ( .A(n364), .B(n289), .Z(z[107]) );
  XOR U3308 ( .A(n290), .B(z[106]), .Z(z[108]) );
  XNOR U3309 ( .A(n292), .B(n291), .Z(n294) );
  NAND U3310 ( .A(n294), .B(n293), .Z(n295) );
  XOR U3311 ( .A(n296), .B(n295), .Z(n297) );
  XNOR U3312 ( .A(n298), .B(n297), .Z(n304) );
  NAND U3313 ( .A(n299), .B(x[104]), .Z(n300) );
  XNOR U3314 ( .A(n301), .B(n300), .Z(n367) );
  XNOR U3315 ( .A(n302), .B(n367), .Z(n303) );
  XOR U3316 ( .A(n304), .B(n303), .Z(z[109]) );
  IV U3317 ( .A(x[15]), .Z(n311) );
  IV U3318 ( .A(x[10]), .Z(n315) );
  XOR U3319 ( .A(x[11]), .B(x[9]), .Z(n307) );
  XOR U3320 ( .A(n315), .B(n307), .Z(n352) );
  IV U3321 ( .A(n352), .Z(n309) );
  XOR U3322 ( .A(x[13]), .B(n309), .Z(n305) );
  IV U3323 ( .A(x[9]), .Z(n655) );
  XNOR U3324 ( .A(n311), .B(n655), .Z(n515) );
  NAND U3325 ( .A(n305), .B(n515), .Z(n306) );
  XNOR U3326 ( .A(n311), .B(n306), .Z(n339) );
  XOR U3327 ( .A(x[12]), .B(n311), .Z(n314) );
  XNOR U3328 ( .A(x[14]), .B(n309), .Z(n497) );
  NOR U3329 ( .A(n314), .B(n497), .Z(n318) );
  IV U3330 ( .A(x[13]), .Z(n353) );
  XOR U3331 ( .A(x[8]), .B(x[14]), .Z(n310) );
  XOR U3332 ( .A(n353), .B(n310), .Z(n325) );
  IV U3333 ( .A(n325), .Z(n656) );
  XOR U3334 ( .A(n314), .B(n307), .Z(n316) );
  XNOR U3335 ( .A(x[8]), .B(n316), .Z(n350) );
  XNOR U3336 ( .A(n656), .B(n350), .Z(n648) );
  XNOR U3337 ( .A(x[15]), .B(n315), .Z(n673) );
  NANDN U3338 ( .A(n648), .B(n673), .Z(n308) );
  XOR U3339 ( .A(n318), .B(n308), .Z(n333) );
  XOR U3340 ( .A(n310), .B(n309), .Z(n313) );
  XNOR U3341 ( .A(n325), .B(n311), .Z(n516) );
  ANDN U3342 ( .B(n313), .A(n516), .Z(n312) );
  XOR U3343 ( .A(n333), .B(n312), .Z(n328) );
  IV U3344 ( .A(n313), .Z(n647) );
  IV U3345 ( .A(n314), .Z(n507) );
  XNOR U3346 ( .A(n655), .B(n315), .Z(n321) );
  XOR U3347 ( .A(n507), .B(n321), .Z(n501) );
  IV U3348 ( .A(n316), .Z(n344) );
  NANDN U3349 ( .A(n501), .B(n344), .Z(n329) );
  XNOR U3350 ( .A(x[12]), .B(x[10]), .Z(n508) );
  XNOR U3351 ( .A(n648), .B(n497), .Z(n498) );
  OR U3352 ( .A(n508), .B(n498), .Z(n317) );
  XOR U3353 ( .A(n318), .B(n317), .Z(n327) );
  XOR U3354 ( .A(n329), .B(n327), .Z(n320) );
  XNOR U3355 ( .A(x[8]), .B(n507), .Z(n319) );
  XNOR U3356 ( .A(n320), .B(n319), .Z(n323) );
  XOR U3357 ( .A(n321), .B(n516), .Z(n505) );
  NAND U3358 ( .A(n350), .B(n505), .Z(n322) );
  XNOR U3359 ( .A(n323), .B(n322), .Z(n324) );
  XOR U3360 ( .A(n647), .B(n324), .Z(n356) );
  IV U3361 ( .A(n356), .Z(n359) );
  NAND U3362 ( .A(n325), .B(n655), .Z(n326) );
  XOR U3363 ( .A(n327), .B(n326), .Z(n338) );
  XNOR U3364 ( .A(n328), .B(n338), .Z(n348) );
  NAND U3365 ( .A(n359), .B(n348), .Z(n337) );
  XOR U3366 ( .A(n656), .B(x[12]), .Z(n502) );
  AND U3367 ( .A(n502), .B(x[8]), .Z(n335) );
  XNOR U3368 ( .A(n505), .B(n329), .Z(n331) );
  XNOR U3369 ( .A(x[9]), .B(n350), .Z(n330) );
  XNOR U3370 ( .A(n331), .B(n330), .Z(n332) );
  XOR U3371 ( .A(n333), .B(n332), .Z(n334) );
  XNOR U3372 ( .A(n335), .B(n334), .Z(n358) );
  NANDN U3373 ( .A(n348), .B(n358), .Z(n336) );
  AND U3374 ( .A(n337), .B(n336), .Z(n342) );
  XNOR U3375 ( .A(n339), .B(n338), .Z(n345) );
  NANDN U3376 ( .A(n345), .B(n356), .Z(n340) );
  XNOR U3377 ( .A(n342), .B(n340), .Z(n354) );
  OR U3378 ( .A(n341), .B(n354), .Z(n495) );
  NANDN U3379 ( .A(n358), .B(n341), .Z(n347) );
  XOR U3380 ( .A(n345), .B(n342), .Z(n343) );
  XNOR U3381 ( .A(n347), .B(n343), .Z(n355) );
  NOR U3382 ( .A(n355), .B(n345), .Z(n349) );
  XOR U3383 ( .A(n495), .B(n349), .Z(n500) );
  NANDN U3384 ( .A(n500), .B(n344), .Z(n664) );
  ANDN U3385 ( .B(n359), .A(n345), .Z(n346) );
  XNOR U3386 ( .A(n347), .B(n346), .Z(n361) );
  OR U3387 ( .A(n361), .B(n348), .Z(n496) );
  XNOR U3388 ( .A(n496), .B(n349), .Z(n504) );
  AND U3389 ( .A(n504), .B(n350), .Z(n351) );
  XOR U3390 ( .A(n664), .B(n351), .Z(n670) );
  XOR U3391 ( .A(n353), .B(n352), .Z(n357) );
  ANDN U3392 ( .B(n358), .A(n354), .Z(n493) );
  NOR U3393 ( .A(n356), .B(n355), .Z(n362) );
  XOR U3394 ( .A(n493), .B(n362), .Z(n514) );
  NAND U3395 ( .A(n357), .B(n514), .Z(n651) );
  XOR U3396 ( .A(n359), .B(n358), .Z(n360) );
  NANDN U3397 ( .A(n361), .B(n360), .Z(n494) );
  XOR U3398 ( .A(n494), .B(n362), .Z(n658) );
  NANDN U3399 ( .A(n658), .B(n656), .Z(n363) );
  XNOR U3400 ( .A(n651), .B(n363), .Z(n519) );
  XOR U3401 ( .A(n670), .B(n519), .Z(n654) );
  IV U3402 ( .A(n654), .Z(z[10]) );
  XNOR U3403 ( .A(n365), .B(n364), .Z(z[110]) );
  XNOR U3404 ( .A(n367), .B(n366), .Z(n368) );
  XNOR U3405 ( .A(z[105]), .B(n368), .Z(z[111]) );
  IV U3406 ( .A(x[113]), .Z(n475) );
  XOR U3407 ( .A(x[112]), .B(x[118]), .Z(n370) );
  XOR U3408 ( .A(x[117]), .B(n370), .Z(n474) );
  IV U3409 ( .A(n474), .Z(n371) );
  AND U3410 ( .A(n475), .B(n371), .Z(n378) );
  XNOR U3411 ( .A(x[115]), .B(n475), .Z(n374) );
  XNOR U3412 ( .A(x[114]), .B(n374), .Z(n369) );
  XNOR U3413 ( .A(n370), .B(n369), .Z(n434) );
  IV U3414 ( .A(n434), .Z(n380) );
  XNOR U3415 ( .A(n380), .B(n474), .Z(n433) );
  IV U3416 ( .A(x[119]), .Z(n372) );
  XNOR U3417 ( .A(x[113]), .B(n372), .Z(n465) );
  NAND U3418 ( .A(n433), .B(n465), .Z(n383) );
  XNOR U3419 ( .A(n372), .B(n371), .Z(n379) );
  IV U3420 ( .A(n379), .Z(n463) );
  XOR U3421 ( .A(n434), .B(n463), .Z(n399) );
  XNOR U3422 ( .A(n383), .B(n399), .Z(n376) );
  XOR U3423 ( .A(x[112]), .B(n380), .Z(n409) );
  XOR U3424 ( .A(x[116]), .B(n372), .Z(n373) );
  IV U3425 ( .A(n373), .Z(n438) );
  NANDN U3426 ( .A(n409), .B(n438), .Z(n382) );
  XNOR U3427 ( .A(n374), .B(n373), .Z(n427) );
  XNOR U3428 ( .A(n433), .B(n427), .Z(n425) );
  XOR U3429 ( .A(x[114]), .B(x[116]), .Z(n440) );
  NANDN U3430 ( .A(n425), .B(n440), .Z(n375) );
  XOR U3431 ( .A(n382), .B(n375), .Z(n401) );
  XNOR U3432 ( .A(n376), .B(n401), .Z(n377) );
  XOR U3433 ( .A(n378), .B(n377), .Z(n414) );
  IV U3434 ( .A(n414), .Z(n420) );
  AND U3435 ( .A(n380), .B(n379), .Z(n385) );
  XOR U3436 ( .A(x[112]), .B(n427), .Z(n428) );
  XNOR U3437 ( .A(n474), .B(n428), .Z(n430) );
  XOR U3438 ( .A(x[114]), .B(x[119]), .Z(n455) );
  NANDN U3439 ( .A(n430), .B(n455), .Z(n381) );
  XNOR U3440 ( .A(n382), .B(n381), .Z(n390) );
  XNOR U3441 ( .A(n383), .B(n390), .Z(n384) );
  XOR U3442 ( .A(n385), .B(n384), .Z(n410) );
  XNOR U3443 ( .A(x[116]), .B(n474), .Z(n448) );
  ANDN U3444 ( .B(x[112]), .A(n448), .Z(n392) );
  XOR U3445 ( .A(x[114]), .B(x[113]), .Z(n386) );
  XOR U3446 ( .A(n463), .B(n386), .Z(n437) );
  XOR U3447 ( .A(n438), .B(n386), .Z(n443) );
  NAND U3448 ( .A(n427), .B(n443), .Z(n394) );
  XNOR U3449 ( .A(n437), .B(n394), .Z(n388) );
  XNOR U3450 ( .A(x[113]), .B(n428), .Z(n387) );
  XNOR U3451 ( .A(n388), .B(n387), .Z(n389) );
  XOR U3452 ( .A(n390), .B(n389), .Z(n391) );
  XOR U3453 ( .A(n392), .B(n391), .Z(n412) );
  NAND U3454 ( .A(n410), .B(n412), .Z(n393) );
  NAND U3455 ( .A(n420), .B(n393), .Z(n404) );
  IV U3456 ( .A(n410), .Z(n411) );
  IV U3457 ( .A(n412), .Z(n418) );
  XOR U3458 ( .A(n394), .B(n448), .Z(n397) );
  AND U3459 ( .A(n437), .B(n428), .Z(n395) );
  XNOR U3460 ( .A(x[112]), .B(n395), .Z(n396) );
  XNOR U3461 ( .A(n397), .B(n396), .Z(n398) );
  XNOR U3462 ( .A(n399), .B(n398), .Z(n400) );
  XNOR U3463 ( .A(n401), .B(n400), .Z(n422) );
  IV U3464 ( .A(n422), .Z(n417) );
  XOR U3465 ( .A(n418), .B(n417), .Z(n402) );
  NAND U3466 ( .A(n411), .B(n402), .Z(n403) );
  AND U3467 ( .A(n404), .B(n403), .Z(n482) );
  NAND U3468 ( .A(n418), .B(n411), .Z(n405) );
  NAND U3469 ( .A(n417), .B(n405), .Z(n408) );
  XOR U3470 ( .A(n411), .B(n414), .Z(n406) );
  NAND U3471 ( .A(n412), .B(n406), .Z(n407) );
  AND U3472 ( .A(n408), .B(n407), .Z(n464) );
  XNOR U3473 ( .A(n482), .B(n464), .Z(n439) );
  OR U3474 ( .A(n439), .B(n409), .Z(n432) );
  NAND U3475 ( .A(n420), .B(n410), .Z(n416) );
  AND U3476 ( .A(n412), .B(n411), .Z(n419) );
  XNOR U3477 ( .A(n417), .B(n419), .Z(n413) );
  NAND U3478 ( .A(n414), .B(n413), .Z(n415) );
  AND U3479 ( .A(n416), .B(n415), .Z(n436) );
  NAND U3480 ( .A(n418), .B(n417), .Z(n424) );
  XNOR U3481 ( .A(n420), .B(n419), .Z(n421) );
  NAND U3482 ( .A(n422), .B(n421), .Z(n423) );
  NAND U3483 ( .A(n424), .B(n423), .Z(n476) );
  XNOR U3484 ( .A(n436), .B(n476), .Z(n454) );
  XOR U3485 ( .A(n454), .B(n439), .Z(n441) );
  OR U3486 ( .A(n441), .B(n425), .Z(n426) );
  XNOR U3487 ( .A(n432), .B(n426), .Z(n458) );
  XOR U3488 ( .A(n436), .B(n482), .Z(n444) );
  NANDN U3489 ( .A(n444), .B(n427), .Z(n484) );
  NANDN U3490 ( .A(n436), .B(n428), .Z(n429) );
  XNOR U3491 ( .A(n484), .B(n429), .Z(n462) );
  XOR U3492 ( .A(n458), .B(n462), .Z(n447) );
  NANDN U3493 ( .A(n430), .B(n454), .Z(n431) );
  XNOR U3494 ( .A(n432), .B(n431), .Z(n490) );
  XNOR U3495 ( .A(n476), .B(n464), .Z(n466) );
  NANDN U3496 ( .A(n466), .B(n433), .Z(n450) );
  NAND U3497 ( .A(n434), .B(n464), .Z(n435) );
  XNOR U3498 ( .A(n450), .B(n435), .Z(n481) );
  XOR U3499 ( .A(n490), .B(n481), .Z(n473) );
  XNOR U3500 ( .A(n447), .B(n473), .Z(z[112]) );
  ANDN U3501 ( .B(n437), .A(n436), .Z(n446) );
  NANDN U3502 ( .A(n439), .B(n438), .Z(n457) );
  NANDN U3503 ( .A(n441), .B(n440), .Z(n442) );
  XNOR U3504 ( .A(n457), .B(n442), .Z(n485) );
  NANDN U3505 ( .A(n444), .B(n443), .Z(n451) );
  XNOR U3506 ( .A(n485), .B(n451), .Z(n445) );
  XOR U3507 ( .A(n446), .B(n445), .Z(n471) );
  XOR U3508 ( .A(n471), .B(n447), .Z(n489) );
  ANDN U3509 ( .B(n482), .A(n448), .Z(n453) );
  NAND U3510 ( .A(n474), .B(n476), .Z(n449) );
  XNOR U3511 ( .A(n450), .B(n449), .Z(n461) );
  XNOR U3512 ( .A(n451), .B(n461), .Z(n452) );
  XNOR U3513 ( .A(n453), .B(n452), .Z(n460) );
  NAND U3514 ( .A(n455), .B(n454), .Z(n456) );
  XNOR U3515 ( .A(n457), .B(n456), .Z(n467) );
  XNOR U3516 ( .A(n458), .B(n467), .Z(n459) );
  XOR U3517 ( .A(n460), .B(n459), .Z(n470) );
  XNOR U3518 ( .A(n489), .B(n470), .Z(z[113]) );
  XNOR U3519 ( .A(n462), .B(n461), .Z(z[114]) );
  AND U3520 ( .A(n464), .B(n463), .Z(n469) );
  NANDN U3521 ( .A(n466), .B(n465), .Z(n479) );
  XNOR U3522 ( .A(n467), .B(n479), .Z(n468) );
  XOR U3523 ( .A(n469), .B(n468), .Z(n488) );
  XOR U3524 ( .A(n471), .B(n470), .Z(n472) );
  XOR U3525 ( .A(n488), .B(n472), .Z(z[115]) );
  XOR U3526 ( .A(n473), .B(z[114]), .Z(z[116]) );
  XNOR U3527 ( .A(n475), .B(n474), .Z(n477) );
  NAND U3528 ( .A(n477), .B(n476), .Z(n478) );
  XOR U3529 ( .A(n479), .B(n478), .Z(n480) );
  XNOR U3530 ( .A(n481), .B(n480), .Z(n487) );
  NAND U3531 ( .A(n482), .B(x[112]), .Z(n483) );
  XNOR U3532 ( .A(n484), .B(n483), .Z(n491) );
  XNOR U3533 ( .A(n485), .B(n491), .Z(n486) );
  XOR U3534 ( .A(n487), .B(n486), .Z(z[117]) );
  XNOR U3535 ( .A(n489), .B(n488), .Z(z[118]) );
  XNOR U3536 ( .A(n491), .B(n490), .Z(n492) );
  XNOR U3537 ( .A(z[113]), .B(n492), .Z(z[119]) );
  XNOR U3538 ( .A(n496), .B(n495), .Z(n662) );
  XOR U3539 ( .A(n646), .B(n662), .Z(n506) );
  NANDN U3540 ( .A(n497), .B(n506), .Z(n650) );
  XNOR U3541 ( .A(n658), .B(n504), .Z(n672) );
  XNOR U3542 ( .A(n506), .B(n672), .Z(n509) );
  OR U3543 ( .A(n498), .B(n509), .Z(n499) );
  XNOR U3544 ( .A(n650), .B(n499), .Z(n671) );
  OR U3545 ( .A(n501), .B(n500), .Z(n511) );
  ANDN U3546 ( .B(n502), .A(n662), .Z(n503) );
  XNOR U3547 ( .A(n511), .B(n503), .Z(n678) );
  AND U3548 ( .A(n505), .B(n504), .Z(n513) );
  NAND U3549 ( .A(n507), .B(n506), .Z(n675) );
  OR U3550 ( .A(n509), .B(n508), .Z(n510) );
  XNOR U3551 ( .A(n675), .B(n510), .Z(n667) );
  XNOR U3552 ( .A(n667), .B(n511), .Z(n512) );
  XOR U3553 ( .A(n513), .B(n512), .Z(n682) );
  NANDN U3554 ( .A(n515), .B(n514), .Z(n660) );
  OR U3555 ( .A(n516), .B(n646), .Z(n517) );
  XOR U3556 ( .A(n660), .B(n517), .Z(n518) );
  XNOR U3557 ( .A(n682), .B(n518), .Z(n677) );
  XNOR U3558 ( .A(n519), .B(n677), .Z(n520) );
  XOR U3559 ( .A(n678), .B(n520), .Z(n521) );
  XOR U3560 ( .A(n671), .B(n521), .Z(z[11]) );
  IV U3561 ( .A(x[121]), .Z(n628) );
  XOR U3562 ( .A(x[120]), .B(x[126]), .Z(n523) );
  XOR U3563 ( .A(x[125]), .B(n523), .Z(n627) );
  IV U3564 ( .A(n627), .Z(n524) );
  AND U3565 ( .A(n628), .B(n524), .Z(n531) );
  XNOR U3566 ( .A(x[123]), .B(n628), .Z(n527) );
  XNOR U3567 ( .A(x[122]), .B(n527), .Z(n522) );
  XNOR U3568 ( .A(n523), .B(n522), .Z(n587) );
  IV U3569 ( .A(n587), .Z(n533) );
  XNOR U3570 ( .A(n533), .B(n627), .Z(n586) );
  IV U3571 ( .A(x[127]), .Z(n525) );
  XNOR U3572 ( .A(x[121]), .B(n525), .Z(n618) );
  NAND U3573 ( .A(n586), .B(n618), .Z(n536) );
  XNOR U3574 ( .A(n525), .B(n524), .Z(n532) );
  IV U3575 ( .A(n532), .Z(n616) );
  XOR U3576 ( .A(n587), .B(n616), .Z(n552) );
  XNOR U3577 ( .A(n536), .B(n552), .Z(n529) );
  XOR U3578 ( .A(x[120]), .B(n533), .Z(n562) );
  XOR U3579 ( .A(x[124]), .B(n525), .Z(n526) );
  IV U3580 ( .A(n526), .Z(n591) );
  NANDN U3581 ( .A(n562), .B(n591), .Z(n535) );
  XNOR U3582 ( .A(n527), .B(n526), .Z(n580) );
  XNOR U3583 ( .A(n586), .B(n580), .Z(n578) );
  XOR U3584 ( .A(x[122]), .B(x[124]), .Z(n593) );
  NANDN U3585 ( .A(n578), .B(n593), .Z(n528) );
  XOR U3586 ( .A(n535), .B(n528), .Z(n554) );
  XNOR U3587 ( .A(n529), .B(n554), .Z(n530) );
  XOR U3588 ( .A(n531), .B(n530), .Z(n567) );
  IV U3589 ( .A(n567), .Z(n573) );
  AND U3590 ( .A(n533), .B(n532), .Z(n538) );
  XOR U3591 ( .A(x[120]), .B(n580), .Z(n581) );
  XNOR U3592 ( .A(n627), .B(n581), .Z(n583) );
  XOR U3593 ( .A(x[122]), .B(x[127]), .Z(n608) );
  NANDN U3594 ( .A(n583), .B(n608), .Z(n534) );
  XNOR U3595 ( .A(n535), .B(n534), .Z(n543) );
  XNOR U3596 ( .A(n536), .B(n543), .Z(n537) );
  XOR U3597 ( .A(n538), .B(n537), .Z(n563) );
  XNOR U3598 ( .A(x[124]), .B(n627), .Z(n601) );
  ANDN U3599 ( .B(x[120]), .A(n601), .Z(n545) );
  XOR U3600 ( .A(x[122]), .B(x[121]), .Z(n539) );
  XOR U3601 ( .A(n616), .B(n539), .Z(n590) );
  XOR U3602 ( .A(n591), .B(n539), .Z(n596) );
  NAND U3603 ( .A(n580), .B(n596), .Z(n547) );
  XNOR U3604 ( .A(n590), .B(n547), .Z(n541) );
  XNOR U3605 ( .A(x[121]), .B(n581), .Z(n540) );
  XNOR U3606 ( .A(n541), .B(n540), .Z(n542) );
  XOR U3607 ( .A(n543), .B(n542), .Z(n544) );
  XOR U3608 ( .A(n545), .B(n544), .Z(n565) );
  NAND U3609 ( .A(n563), .B(n565), .Z(n546) );
  NAND U3610 ( .A(n573), .B(n546), .Z(n557) );
  IV U3611 ( .A(n563), .Z(n564) );
  IV U3612 ( .A(n565), .Z(n571) );
  XOR U3613 ( .A(n547), .B(n601), .Z(n550) );
  AND U3614 ( .A(n590), .B(n581), .Z(n548) );
  XNOR U3615 ( .A(x[120]), .B(n548), .Z(n549) );
  XNOR U3616 ( .A(n550), .B(n549), .Z(n551) );
  XNOR U3617 ( .A(n552), .B(n551), .Z(n553) );
  XNOR U3618 ( .A(n554), .B(n553), .Z(n575) );
  IV U3619 ( .A(n575), .Z(n570) );
  XOR U3620 ( .A(n571), .B(n570), .Z(n555) );
  NAND U3621 ( .A(n564), .B(n555), .Z(n556) );
  AND U3622 ( .A(n557), .B(n556), .Z(n635) );
  NAND U3623 ( .A(n571), .B(n564), .Z(n558) );
  NAND U3624 ( .A(n570), .B(n558), .Z(n561) );
  XOR U3625 ( .A(n564), .B(n567), .Z(n559) );
  NAND U3626 ( .A(n565), .B(n559), .Z(n560) );
  AND U3627 ( .A(n561), .B(n560), .Z(n617) );
  XNOR U3628 ( .A(n635), .B(n617), .Z(n592) );
  OR U3629 ( .A(n592), .B(n562), .Z(n585) );
  NAND U3630 ( .A(n573), .B(n563), .Z(n569) );
  AND U3631 ( .A(n565), .B(n564), .Z(n572) );
  XNOR U3632 ( .A(n570), .B(n572), .Z(n566) );
  NAND U3633 ( .A(n567), .B(n566), .Z(n568) );
  AND U3634 ( .A(n569), .B(n568), .Z(n589) );
  NAND U3635 ( .A(n571), .B(n570), .Z(n577) );
  XNOR U3636 ( .A(n573), .B(n572), .Z(n574) );
  NAND U3637 ( .A(n575), .B(n574), .Z(n576) );
  NAND U3638 ( .A(n577), .B(n576), .Z(n629) );
  XNOR U3639 ( .A(n589), .B(n629), .Z(n607) );
  XOR U3640 ( .A(n607), .B(n592), .Z(n594) );
  OR U3641 ( .A(n594), .B(n578), .Z(n579) );
  XNOR U3642 ( .A(n585), .B(n579), .Z(n611) );
  XOR U3643 ( .A(n589), .B(n635), .Z(n597) );
  NANDN U3644 ( .A(n597), .B(n580), .Z(n637) );
  NANDN U3645 ( .A(n589), .B(n581), .Z(n582) );
  XNOR U3646 ( .A(n637), .B(n582), .Z(n615) );
  XOR U3647 ( .A(n611), .B(n615), .Z(n600) );
  NANDN U3648 ( .A(n583), .B(n607), .Z(n584) );
  XNOR U3649 ( .A(n585), .B(n584), .Z(n643) );
  XNOR U3650 ( .A(n629), .B(n617), .Z(n619) );
  NANDN U3651 ( .A(n619), .B(n586), .Z(n603) );
  NAND U3652 ( .A(n587), .B(n617), .Z(n588) );
  XNOR U3653 ( .A(n603), .B(n588), .Z(n634) );
  XOR U3654 ( .A(n643), .B(n634), .Z(n626) );
  XNOR U3655 ( .A(n600), .B(n626), .Z(z[120]) );
  ANDN U3656 ( .B(n590), .A(n589), .Z(n599) );
  NANDN U3657 ( .A(n592), .B(n591), .Z(n610) );
  NANDN U3658 ( .A(n594), .B(n593), .Z(n595) );
  XNOR U3659 ( .A(n610), .B(n595), .Z(n638) );
  NANDN U3660 ( .A(n597), .B(n596), .Z(n604) );
  XNOR U3661 ( .A(n638), .B(n604), .Z(n598) );
  XOR U3662 ( .A(n599), .B(n598), .Z(n624) );
  XOR U3663 ( .A(n624), .B(n600), .Z(n642) );
  ANDN U3664 ( .B(n635), .A(n601), .Z(n606) );
  NAND U3665 ( .A(n627), .B(n629), .Z(n602) );
  XNOR U3666 ( .A(n603), .B(n602), .Z(n614) );
  XNOR U3667 ( .A(n604), .B(n614), .Z(n605) );
  XNOR U3668 ( .A(n606), .B(n605), .Z(n613) );
  NAND U3669 ( .A(n608), .B(n607), .Z(n609) );
  XNOR U3670 ( .A(n610), .B(n609), .Z(n620) );
  XNOR U3671 ( .A(n611), .B(n620), .Z(n612) );
  XOR U3672 ( .A(n613), .B(n612), .Z(n623) );
  XNOR U3673 ( .A(n642), .B(n623), .Z(z[121]) );
  XNOR U3674 ( .A(n615), .B(n614), .Z(z[122]) );
  AND U3675 ( .A(n617), .B(n616), .Z(n622) );
  NANDN U3676 ( .A(n619), .B(n618), .Z(n632) );
  XNOR U3677 ( .A(n620), .B(n632), .Z(n621) );
  XOR U3678 ( .A(n622), .B(n621), .Z(n641) );
  XOR U3679 ( .A(n624), .B(n623), .Z(n625) );
  XOR U3680 ( .A(n641), .B(n625), .Z(z[123]) );
  XOR U3681 ( .A(n626), .B(z[122]), .Z(z[124]) );
  XNOR U3682 ( .A(n628), .B(n627), .Z(n630) );
  NAND U3683 ( .A(n630), .B(n629), .Z(n631) );
  XOR U3684 ( .A(n632), .B(n631), .Z(n633) );
  XNOR U3685 ( .A(n634), .B(n633), .Z(n640) );
  NAND U3686 ( .A(n635), .B(x[120]), .Z(n636) );
  XNOR U3687 ( .A(n637), .B(n636), .Z(n644) );
  XNOR U3688 ( .A(n638), .B(n644), .Z(n639) );
  XOR U3689 ( .A(n640), .B(n639), .Z(z[125]) );
  XNOR U3690 ( .A(n642), .B(n641), .Z(z[126]) );
  XNOR U3691 ( .A(n644), .B(n643), .Z(n645) );
  XNOR U3692 ( .A(z[121]), .B(n645), .Z(z[127]) );
  NOR U3693 ( .A(n647), .B(n646), .Z(n653) );
  NANDN U3694 ( .A(n648), .B(n672), .Z(n649) );
  XNOR U3695 ( .A(n650), .B(n649), .Z(n663) );
  XNOR U3696 ( .A(n651), .B(n663), .Z(n652) );
  XOR U3697 ( .A(n653), .B(n652), .Z(n1947) );
  XOR U3698 ( .A(n1947), .B(n654), .Z(z[12]) );
  XNOR U3699 ( .A(n656), .B(n655), .Z(n657) );
  NANDN U3700 ( .A(n658), .B(n657), .Z(n659) );
  XOR U3701 ( .A(n660), .B(n659), .Z(n661) );
  XNOR U3702 ( .A(n1947), .B(n661), .Z(n669) );
  ANDN U3703 ( .B(x[8]), .A(n662), .Z(n666) );
  XNOR U3704 ( .A(n664), .B(n663), .Z(n665) );
  XOR U3705 ( .A(n666), .B(n665), .Z(n683) );
  XNOR U3706 ( .A(n667), .B(n683), .Z(n668) );
  XOR U3707 ( .A(n669), .B(n668), .Z(z[13]) );
  XNOR U3708 ( .A(n671), .B(n670), .Z(n1948) );
  NAND U3709 ( .A(n673), .B(n672), .Z(n674) );
  XNOR U3710 ( .A(n675), .B(n674), .Z(n679) );
  XNOR U3711 ( .A(n1948), .B(n679), .Z(n676) );
  XOR U3712 ( .A(n677), .B(n676), .Z(z[14]) );
  XNOR U3713 ( .A(n679), .B(n678), .Z(n680) );
  XNOR U3714 ( .A(z[10]), .B(n680), .Z(n681) );
  XOR U3715 ( .A(n682), .B(n681), .Z(z[9]) );
  XNOR U3716 ( .A(n683), .B(z[9]), .Z(z[15]) );
  IV U3717 ( .A(x[17]), .Z(n815) );
  XOR U3718 ( .A(x[16]), .B(x[22]), .Z(n685) );
  XOR U3719 ( .A(x[21]), .B(n685), .Z(n814) );
  IV U3720 ( .A(n814), .Z(n686) );
  AND U3721 ( .A(n815), .B(n686), .Z(n693) );
  XNOR U3722 ( .A(x[19]), .B(n815), .Z(n689) );
  XNOR U3723 ( .A(x[18]), .B(n689), .Z(n684) );
  XNOR U3724 ( .A(n685), .B(n684), .Z(n749) );
  IV U3725 ( .A(n749), .Z(n695) );
  XNOR U3726 ( .A(n695), .B(n814), .Z(n748) );
  IV U3727 ( .A(x[23]), .Z(n687) );
  XNOR U3728 ( .A(x[17]), .B(n687), .Z(n780) );
  NAND U3729 ( .A(n748), .B(n780), .Z(n698) );
  XNOR U3730 ( .A(n687), .B(n686), .Z(n694) );
  IV U3731 ( .A(n694), .Z(n778) );
  XOR U3732 ( .A(n749), .B(n778), .Z(n714) );
  XNOR U3733 ( .A(n698), .B(n714), .Z(n691) );
  XOR U3734 ( .A(x[16]), .B(n695), .Z(n724) );
  XOR U3735 ( .A(x[20]), .B(n687), .Z(n688) );
  IV U3736 ( .A(n688), .Z(n753) );
  NANDN U3737 ( .A(n724), .B(n753), .Z(n697) );
  XNOR U3738 ( .A(n689), .B(n688), .Z(n742) );
  XNOR U3739 ( .A(n748), .B(n742), .Z(n740) );
  XOR U3740 ( .A(x[18]), .B(x[20]), .Z(n755) );
  NANDN U3741 ( .A(n740), .B(n755), .Z(n690) );
  XOR U3742 ( .A(n697), .B(n690), .Z(n716) );
  XNOR U3743 ( .A(n691), .B(n716), .Z(n692) );
  XOR U3744 ( .A(n693), .B(n692), .Z(n729) );
  IV U3745 ( .A(n729), .Z(n735) );
  AND U3746 ( .A(n695), .B(n694), .Z(n700) );
  XOR U3747 ( .A(x[16]), .B(n742), .Z(n743) );
  XNOR U3748 ( .A(n814), .B(n743), .Z(n745) );
  XOR U3749 ( .A(x[18]), .B(x[23]), .Z(n770) );
  NANDN U3750 ( .A(n745), .B(n770), .Z(n696) );
  XNOR U3751 ( .A(n697), .B(n696), .Z(n705) );
  XNOR U3752 ( .A(n698), .B(n705), .Z(n699) );
  XOR U3753 ( .A(n700), .B(n699), .Z(n725) );
  XNOR U3754 ( .A(x[20]), .B(n814), .Z(n763) );
  ANDN U3755 ( .B(x[16]), .A(n763), .Z(n707) );
  XOR U3756 ( .A(x[18]), .B(x[17]), .Z(n701) );
  XOR U3757 ( .A(n778), .B(n701), .Z(n752) );
  XOR U3758 ( .A(n753), .B(n701), .Z(n758) );
  NAND U3759 ( .A(n742), .B(n758), .Z(n709) );
  XNOR U3760 ( .A(n752), .B(n709), .Z(n703) );
  XNOR U3761 ( .A(x[17]), .B(n743), .Z(n702) );
  XNOR U3762 ( .A(n703), .B(n702), .Z(n704) );
  XOR U3763 ( .A(n705), .B(n704), .Z(n706) );
  XOR U3764 ( .A(n707), .B(n706), .Z(n727) );
  NAND U3765 ( .A(n725), .B(n727), .Z(n708) );
  NAND U3766 ( .A(n735), .B(n708), .Z(n719) );
  IV U3767 ( .A(n725), .Z(n726) );
  IV U3768 ( .A(n727), .Z(n733) );
  XOR U3769 ( .A(n709), .B(n763), .Z(n712) );
  AND U3770 ( .A(n752), .B(n743), .Z(n710) );
  XNOR U3771 ( .A(x[16]), .B(n710), .Z(n711) );
  XNOR U3772 ( .A(n712), .B(n711), .Z(n713) );
  XNOR U3773 ( .A(n714), .B(n713), .Z(n715) );
  XNOR U3774 ( .A(n716), .B(n715), .Z(n737) );
  IV U3775 ( .A(n737), .Z(n732) );
  XOR U3776 ( .A(n733), .B(n732), .Z(n717) );
  NAND U3777 ( .A(n726), .B(n717), .Z(n718) );
  AND U3778 ( .A(n719), .B(n718), .Z(n822) );
  NAND U3779 ( .A(n733), .B(n726), .Z(n720) );
  NAND U3780 ( .A(n732), .B(n720), .Z(n723) );
  XOR U3781 ( .A(n726), .B(n729), .Z(n721) );
  NAND U3782 ( .A(n727), .B(n721), .Z(n722) );
  AND U3783 ( .A(n723), .B(n722), .Z(n779) );
  XNOR U3784 ( .A(n822), .B(n779), .Z(n754) );
  OR U3785 ( .A(n754), .B(n724), .Z(n747) );
  NAND U3786 ( .A(n735), .B(n725), .Z(n731) );
  AND U3787 ( .A(n727), .B(n726), .Z(n734) );
  XNOR U3788 ( .A(n732), .B(n734), .Z(n728) );
  NAND U3789 ( .A(n729), .B(n728), .Z(n730) );
  AND U3790 ( .A(n731), .B(n730), .Z(n751) );
  NAND U3791 ( .A(n733), .B(n732), .Z(n739) );
  XNOR U3792 ( .A(n735), .B(n734), .Z(n736) );
  NAND U3793 ( .A(n737), .B(n736), .Z(n738) );
  NAND U3794 ( .A(n739), .B(n738), .Z(n816) );
  XNOR U3795 ( .A(n751), .B(n816), .Z(n769) );
  XOR U3796 ( .A(n769), .B(n754), .Z(n756) );
  OR U3797 ( .A(n756), .B(n740), .Z(n741) );
  XNOR U3798 ( .A(n747), .B(n741), .Z(n773) );
  XOR U3799 ( .A(n751), .B(n822), .Z(n759) );
  NANDN U3800 ( .A(n759), .B(n742), .Z(n824) );
  NANDN U3801 ( .A(n751), .B(n743), .Z(n744) );
  XNOR U3802 ( .A(n824), .B(n744), .Z(n777) );
  XOR U3803 ( .A(n773), .B(n777), .Z(n762) );
  NANDN U3804 ( .A(n745), .B(n769), .Z(n746) );
  XNOR U3805 ( .A(n747), .B(n746), .Z(n830) );
  XNOR U3806 ( .A(n816), .B(n779), .Z(n781) );
  NANDN U3807 ( .A(n781), .B(n748), .Z(n765) );
  NAND U3808 ( .A(n749), .B(n779), .Z(n750) );
  XNOR U3809 ( .A(n765), .B(n750), .Z(n821) );
  XOR U3810 ( .A(n830), .B(n821), .Z(n813) );
  XNOR U3811 ( .A(n762), .B(n813), .Z(z[16]) );
  ANDN U3812 ( .B(n752), .A(n751), .Z(n761) );
  NANDN U3813 ( .A(n754), .B(n753), .Z(n772) );
  NANDN U3814 ( .A(n756), .B(n755), .Z(n757) );
  XNOR U3815 ( .A(n772), .B(n757), .Z(n825) );
  NANDN U3816 ( .A(n759), .B(n758), .Z(n766) );
  XNOR U3817 ( .A(n825), .B(n766), .Z(n760) );
  XOR U3818 ( .A(n761), .B(n760), .Z(n786) );
  XOR U3819 ( .A(n786), .B(n762), .Z(n829) );
  ANDN U3820 ( .B(n822), .A(n763), .Z(n768) );
  NAND U3821 ( .A(n814), .B(n816), .Z(n764) );
  XNOR U3822 ( .A(n765), .B(n764), .Z(n776) );
  XNOR U3823 ( .A(n766), .B(n776), .Z(n767) );
  XNOR U3824 ( .A(n768), .B(n767), .Z(n775) );
  NAND U3825 ( .A(n770), .B(n769), .Z(n771) );
  XNOR U3826 ( .A(n772), .B(n771), .Z(n782) );
  XNOR U3827 ( .A(n773), .B(n782), .Z(n774) );
  XOR U3828 ( .A(n775), .B(n774), .Z(n785) );
  XNOR U3829 ( .A(n829), .B(n785), .Z(z[17]) );
  XNOR U3830 ( .A(n777), .B(n776), .Z(z[18]) );
  AND U3831 ( .A(n779), .B(n778), .Z(n784) );
  NANDN U3832 ( .A(n781), .B(n780), .Z(n819) );
  XNOR U3833 ( .A(n782), .B(n819), .Z(n783) );
  XOR U3834 ( .A(n784), .B(n783), .Z(n828) );
  XOR U3835 ( .A(n786), .B(n785), .Z(n787) );
  XOR U3836 ( .A(n828), .B(n787), .Z(z[19]) );
  ANDN U3837 ( .B(n789), .A(n788), .Z(n798) );
  NANDN U3838 ( .A(n791), .B(n790), .Z(n809) );
  NANDN U3839 ( .A(n793), .B(n792), .Z(n794) );
  XNOR U3840 ( .A(n809), .B(n794), .Z(n1457) );
  NANDN U3841 ( .A(n796), .B(n795), .Z(n803) );
  XNOR U3842 ( .A(n1457), .B(n803), .Z(n797) );
  XOR U3843 ( .A(n798), .B(n797), .Z(n1091) );
  XOR U3844 ( .A(n1091), .B(n799), .Z(n1600) );
  ANDN U3845 ( .B(n1454), .A(n800), .Z(n805) );
  NAND U3846 ( .A(n1446), .B(n1448), .Z(n801) );
  XNOR U3847 ( .A(n802), .B(n801), .Z(n952) );
  XNOR U3848 ( .A(n803), .B(n952), .Z(n804) );
  XNOR U3849 ( .A(n805), .B(n804), .Z(n812) );
  NAND U3850 ( .A(n807), .B(n806), .Z(n808) );
  XNOR U3851 ( .A(n809), .B(n808), .Z(n1087) );
  XNOR U3852 ( .A(n810), .B(n1087), .Z(n811) );
  XOR U3853 ( .A(n812), .B(n811), .Z(n1090) );
  XNOR U3854 ( .A(n1600), .B(n1090), .Z(z[1]) );
  XOR U3855 ( .A(n813), .B(z[18]), .Z(z[20]) );
  XNOR U3856 ( .A(n815), .B(n814), .Z(n817) );
  NAND U3857 ( .A(n817), .B(n816), .Z(n818) );
  XOR U3858 ( .A(n819), .B(n818), .Z(n820) );
  XNOR U3859 ( .A(n821), .B(n820), .Z(n827) );
  NAND U3860 ( .A(n822), .B(x[16]), .Z(n823) );
  XNOR U3861 ( .A(n824), .B(n823), .Z(n831) );
  XNOR U3862 ( .A(n825), .B(n831), .Z(n826) );
  XOR U3863 ( .A(n827), .B(n826), .Z(z[21]) );
  XNOR U3864 ( .A(n829), .B(n828), .Z(z[22]) );
  XNOR U3865 ( .A(n831), .B(n830), .Z(n832) );
  XNOR U3866 ( .A(z[17]), .B(n832), .Z(z[23]) );
  IV U3867 ( .A(x[25]), .Z(n939) );
  XOR U3868 ( .A(x[24]), .B(x[30]), .Z(n834) );
  XOR U3869 ( .A(x[29]), .B(n834), .Z(n938) );
  IV U3870 ( .A(n938), .Z(n835) );
  AND U3871 ( .A(n939), .B(n835), .Z(n842) );
  XNOR U3872 ( .A(x[27]), .B(n939), .Z(n838) );
  XNOR U3873 ( .A(x[26]), .B(n838), .Z(n833) );
  XNOR U3874 ( .A(n834), .B(n833), .Z(n898) );
  IV U3875 ( .A(n898), .Z(n844) );
  XNOR U3876 ( .A(n844), .B(n938), .Z(n897) );
  IV U3877 ( .A(x[31]), .Z(n836) );
  XNOR U3878 ( .A(x[25]), .B(n836), .Z(n929) );
  NAND U3879 ( .A(n897), .B(n929), .Z(n847) );
  XNOR U3880 ( .A(n836), .B(n835), .Z(n843) );
  IV U3881 ( .A(n843), .Z(n927) );
  XOR U3882 ( .A(n898), .B(n927), .Z(n863) );
  XNOR U3883 ( .A(n847), .B(n863), .Z(n840) );
  XOR U3884 ( .A(x[24]), .B(n844), .Z(n873) );
  XOR U3885 ( .A(x[28]), .B(n836), .Z(n837) );
  IV U3886 ( .A(n837), .Z(n902) );
  NANDN U3887 ( .A(n873), .B(n902), .Z(n846) );
  XNOR U3888 ( .A(n838), .B(n837), .Z(n891) );
  XNOR U3889 ( .A(n897), .B(n891), .Z(n889) );
  XOR U3890 ( .A(x[26]), .B(x[28]), .Z(n904) );
  NANDN U3891 ( .A(n889), .B(n904), .Z(n839) );
  XOR U3892 ( .A(n846), .B(n839), .Z(n865) );
  XNOR U3893 ( .A(n840), .B(n865), .Z(n841) );
  XOR U3894 ( .A(n842), .B(n841), .Z(n878) );
  IV U3895 ( .A(n878), .Z(n884) );
  AND U3896 ( .A(n844), .B(n843), .Z(n849) );
  XOR U3897 ( .A(x[24]), .B(n891), .Z(n892) );
  XNOR U3898 ( .A(n938), .B(n892), .Z(n894) );
  XOR U3899 ( .A(x[26]), .B(x[31]), .Z(n919) );
  NANDN U3900 ( .A(n894), .B(n919), .Z(n845) );
  XNOR U3901 ( .A(n846), .B(n845), .Z(n854) );
  XNOR U3902 ( .A(n847), .B(n854), .Z(n848) );
  XOR U3903 ( .A(n849), .B(n848), .Z(n874) );
  XNOR U3904 ( .A(x[28]), .B(n938), .Z(n912) );
  ANDN U3905 ( .B(x[24]), .A(n912), .Z(n856) );
  XOR U3906 ( .A(x[26]), .B(x[25]), .Z(n850) );
  XOR U3907 ( .A(n927), .B(n850), .Z(n901) );
  XOR U3908 ( .A(n902), .B(n850), .Z(n907) );
  NAND U3909 ( .A(n891), .B(n907), .Z(n858) );
  XNOR U3910 ( .A(n901), .B(n858), .Z(n852) );
  XNOR U3911 ( .A(x[25]), .B(n892), .Z(n851) );
  XNOR U3912 ( .A(n852), .B(n851), .Z(n853) );
  XOR U3913 ( .A(n854), .B(n853), .Z(n855) );
  XOR U3914 ( .A(n856), .B(n855), .Z(n876) );
  NAND U3915 ( .A(n874), .B(n876), .Z(n857) );
  NAND U3916 ( .A(n884), .B(n857), .Z(n868) );
  IV U3917 ( .A(n874), .Z(n875) );
  IV U3918 ( .A(n876), .Z(n882) );
  XOR U3919 ( .A(n858), .B(n912), .Z(n861) );
  AND U3920 ( .A(n901), .B(n892), .Z(n859) );
  XNOR U3921 ( .A(x[24]), .B(n859), .Z(n860) );
  XNOR U3922 ( .A(n861), .B(n860), .Z(n862) );
  XNOR U3923 ( .A(n863), .B(n862), .Z(n864) );
  XNOR U3924 ( .A(n865), .B(n864), .Z(n886) );
  IV U3925 ( .A(n886), .Z(n881) );
  XOR U3926 ( .A(n882), .B(n881), .Z(n866) );
  NAND U3927 ( .A(n875), .B(n866), .Z(n867) );
  AND U3928 ( .A(n868), .B(n867), .Z(n946) );
  NAND U3929 ( .A(n882), .B(n875), .Z(n869) );
  NAND U3930 ( .A(n881), .B(n869), .Z(n872) );
  XOR U3931 ( .A(n875), .B(n878), .Z(n870) );
  NAND U3932 ( .A(n876), .B(n870), .Z(n871) );
  AND U3933 ( .A(n872), .B(n871), .Z(n928) );
  XNOR U3934 ( .A(n946), .B(n928), .Z(n903) );
  OR U3935 ( .A(n903), .B(n873), .Z(n896) );
  NAND U3936 ( .A(n884), .B(n874), .Z(n880) );
  AND U3937 ( .A(n876), .B(n875), .Z(n883) );
  XNOR U3938 ( .A(n881), .B(n883), .Z(n877) );
  NAND U3939 ( .A(n878), .B(n877), .Z(n879) );
  AND U3940 ( .A(n880), .B(n879), .Z(n900) );
  NAND U3941 ( .A(n882), .B(n881), .Z(n888) );
  XNOR U3942 ( .A(n884), .B(n883), .Z(n885) );
  NAND U3943 ( .A(n886), .B(n885), .Z(n887) );
  NAND U3944 ( .A(n888), .B(n887), .Z(n940) );
  XNOR U3945 ( .A(n900), .B(n940), .Z(n918) );
  XOR U3946 ( .A(n918), .B(n903), .Z(n905) );
  OR U3947 ( .A(n905), .B(n889), .Z(n890) );
  XNOR U3948 ( .A(n896), .B(n890), .Z(n922) );
  XOR U3949 ( .A(n900), .B(n946), .Z(n908) );
  NANDN U3950 ( .A(n908), .B(n891), .Z(n948) );
  NANDN U3951 ( .A(n900), .B(n892), .Z(n893) );
  XNOR U3952 ( .A(n948), .B(n893), .Z(n926) );
  XOR U3953 ( .A(n922), .B(n926), .Z(n911) );
  NANDN U3954 ( .A(n894), .B(n918), .Z(n895) );
  XNOR U3955 ( .A(n896), .B(n895), .Z(n956) );
  XNOR U3956 ( .A(n940), .B(n928), .Z(n930) );
  NANDN U3957 ( .A(n930), .B(n897), .Z(n914) );
  NAND U3958 ( .A(n898), .B(n928), .Z(n899) );
  XNOR U3959 ( .A(n914), .B(n899), .Z(n945) );
  XOR U3960 ( .A(n956), .B(n945), .Z(n937) );
  XNOR U3961 ( .A(n911), .B(n937), .Z(z[24]) );
  ANDN U3962 ( .B(n901), .A(n900), .Z(n910) );
  NANDN U3963 ( .A(n903), .B(n902), .Z(n921) );
  NANDN U3964 ( .A(n905), .B(n904), .Z(n906) );
  XNOR U3965 ( .A(n921), .B(n906), .Z(n949) );
  NANDN U3966 ( .A(n908), .B(n907), .Z(n915) );
  XNOR U3967 ( .A(n949), .B(n915), .Z(n909) );
  XOR U3968 ( .A(n910), .B(n909), .Z(n935) );
  XOR U3969 ( .A(n935), .B(n911), .Z(n955) );
  ANDN U3970 ( .B(n946), .A(n912), .Z(n917) );
  NAND U3971 ( .A(n938), .B(n940), .Z(n913) );
  XNOR U3972 ( .A(n914), .B(n913), .Z(n925) );
  XNOR U3973 ( .A(n915), .B(n925), .Z(n916) );
  XNOR U3974 ( .A(n917), .B(n916), .Z(n924) );
  NAND U3975 ( .A(n919), .B(n918), .Z(n920) );
  XNOR U3976 ( .A(n921), .B(n920), .Z(n931) );
  XNOR U3977 ( .A(n922), .B(n931), .Z(n923) );
  XOR U3978 ( .A(n924), .B(n923), .Z(n934) );
  XNOR U3979 ( .A(n955), .B(n934), .Z(z[25]) );
  XNOR U3980 ( .A(n926), .B(n925), .Z(z[26]) );
  AND U3981 ( .A(n928), .B(n927), .Z(n933) );
  NANDN U3982 ( .A(n930), .B(n929), .Z(n943) );
  XNOR U3983 ( .A(n931), .B(n943), .Z(n932) );
  XOR U3984 ( .A(n933), .B(n932), .Z(n954) );
  XOR U3985 ( .A(n935), .B(n934), .Z(n936) );
  XOR U3986 ( .A(n954), .B(n936), .Z(z[27]) );
  XOR U3987 ( .A(n937), .B(z[26]), .Z(z[28]) );
  XNOR U3988 ( .A(n939), .B(n938), .Z(n941) );
  NAND U3989 ( .A(n941), .B(n940), .Z(n942) );
  XOR U3990 ( .A(n943), .B(n942), .Z(n944) );
  XNOR U3991 ( .A(n945), .B(n944), .Z(n951) );
  NAND U3992 ( .A(n946), .B(x[24]), .Z(n947) );
  XNOR U3993 ( .A(n948), .B(n947), .Z(n957) );
  XNOR U3994 ( .A(n949), .B(n957), .Z(n950) );
  XOR U3995 ( .A(n951), .B(n950), .Z(z[29]) );
  XNOR U3996 ( .A(n953), .B(n952), .Z(z[2]) );
  XNOR U3997 ( .A(n955), .B(n954), .Z(z[30]) );
  XNOR U3998 ( .A(n957), .B(n956), .Z(n958) );
  XNOR U3999 ( .A(z[25]), .B(n958), .Z(z[31]) );
  IV U4000 ( .A(x[33]), .Z(n1065) );
  XOR U4001 ( .A(x[32]), .B(x[38]), .Z(n960) );
  XOR U4002 ( .A(x[37]), .B(n960), .Z(n1064) );
  IV U4003 ( .A(n1064), .Z(n961) );
  AND U4004 ( .A(n1065), .B(n961), .Z(n968) );
  XNOR U4005 ( .A(x[35]), .B(n1065), .Z(n964) );
  XNOR U4006 ( .A(x[34]), .B(n964), .Z(n959) );
  XNOR U4007 ( .A(n960), .B(n959), .Z(n1024) );
  IV U4008 ( .A(n1024), .Z(n970) );
  XNOR U4009 ( .A(n970), .B(n1064), .Z(n1023) );
  IV U4010 ( .A(x[39]), .Z(n962) );
  XNOR U4011 ( .A(x[33]), .B(n962), .Z(n1055) );
  NAND U4012 ( .A(n1023), .B(n1055), .Z(n973) );
  XNOR U4013 ( .A(n962), .B(n961), .Z(n969) );
  IV U4014 ( .A(n969), .Z(n1053) );
  XOR U4015 ( .A(n1024), .B(n1053), .Z(n989) );
  XNOR U4016 ( .A(n973), .B(n989), .Z(n966) );
  XOR U4017 ( .A(x[32]), .B(n970), .Z(n999) );
  XOR U4018 ( .A(x[36]), .B(n962), .Z(n963) );
  IV U4019 ( .A(n963), .Z(n1028) );
  NANDN U4020 ( .A(n999), .B(n1028), .Z(n972) );
  XNOR U4021 ( .A(n964), .B(n963), .Z(n1017) );
  XNOR U4022 ( .A(n1023), .B(n1017), .Z(n1015) );
  XOR U4023 ( .A(x[34]), .B(x[36]), .Z(n1030) );
  NANDN U4024 ( .A(n1015), .B(n1030), .Z(n965) );
  XOR U4025 ( .A(n972), .B(n965), .Z(n991) );
  XNOR U4026 ( .A(n966), .B(n991), .Z(n967) );
  XOR U4027 ( .A(n968), .B(n967), .Z(n1004) );
  IV U4028 ( .A(n1004), .Z(n1010) );
  AND U4029 ( .A(n970), .B(n969), .Z(n975) );
  XOR U4030 ( .A(x[32]), .B(n1017), .Z(n1018) );
  XNOR U4031 ( .A(n1064), .B(n1018), .Z(n1020) );
  XOR U4032 ( .A(x[34]), .B(x[39]), .Z(n1045) );
  NANDN U4033 ( .A(n1020), .B(n1045), .Z(n971) );
  XNOR U4034 ( .A(n972), .B(n971), .Z(n980) );
  XNOR U4035 ( .A(n973), .B(n980), .Z(n974) );
  XOR U4036 ( .A(n975), .B(n974), .Z(n1000) );
  XNOR U4037 ( .A(x[36]), .B(n1064), .Z(n1038) );
  ANDN U4038 ( .B(x[32]), .A(n1038), .Z(n982) );
  XOR U4039 ( .A(x[34]), .B(x[33]), .Z(n976) );
  XOR U4040 ( .A(n1053), .B(n976), .Z(n1027) );
  XOR U4041 ( .A(n1028), .B(n976), .Z(n1033) );
  NAND U4042 ( .A(n1017), .B(n1033), .Z(n984) );
  XNOR U4043 ( .A(n1027), .B(n984), .Z(n978) );
  XNOR U4044 ( .A(x[33]), .B(n1018), .Z(n977) );
  XNOR U4045 ( .A(n978), .B(n977), .Z(n979) );
  XOR U4046 ( .A(n980), .B(n979), .Z(n981) );
  XOR U4047 ( .A(n982), .B(n981), .Z(n1002) );
  NAND U4048 ( .A(n1000), .B(n1002), .Z(n983) );
  NAND U4049 ( .A(n1010), .B(n983), .Z(n994) );
  IV U4050 ( .A(n1000), .Z(n1001) );
  IV U4051 ( .A(n1002), .Z(n1008) );
  XOR U4052 ( .A(n984), .B(n1038), .Z(n987) );
  AND U4053 ( .A(n1027), .B(n1018), .Z(n985) );
  XNOR U4054 ( .A(x[32]), .B(n985), .Z(n986) );
  XNOR U4055 ( .A(n987), .B(n986), .Z(n988) );
  XNOR U4056 ( .A(n989), .B(n988), .Z(n990) );
  XNOR U4057 ( .A(n991), .B(n990), .Z(n1012) );
  IV U4058 ( .A(n1012), .Z(n1007) );
  XOR U4059 ( .A(n1008), .B(n1007), .Z(n992) );
  NAND U4060 ( .A(n1001), .B(n992), .Z(n993) );
  AND U4061 ( .A(n994), .B(n993), .Z(n1072) );
  NAND U4062 ( .A(n1008), .B(n1001), .Z(n995) );
  NAND U4063 ( .A(n1007), .B(n995), .Z(n998) );
  XOR U4064 ( .A(n1001), .B(n1004), .Z(n996) );
  NAND U4065 ( .A(n1002), .B(n996), .Z(n997) );
  AND U4066 ( .A(n998), .B(n997), .Z(n1054) );
  XNOR U4067 ( .A(n1072), .B(n1054), .Z(n1029) );
  OR U4068 ( .A(n1029), .B(n999), .Z(n1022) );
  NAND U4069 ( .A(n1010), .B(n1000), .Z(n1006) );
  AND U4070 ( .A(n1002), .B(n1001), .Z(n1009) );
  XNOR U4071 ( .A(n1007), .B(n1009), .Z(n1003) );
  NAND U4072 ( .A(n1004), .B(n1003), .Z(n1005) );
  AND U4073 ( .A(n1006), .B(n1005), .Z(n1026) );
  NAND U4074 ( .A(n1008), .B(n1007), .Z(n1014) );
  XNOR U4075 ( .A(n1010), .B(n1009), .Z(n1011) );
  NAND U4076 ( .A(n1012), .B(n1011), .Z(n1013) );
  NAND U4077 ( .A(n1014), .B(n1013), .Z(n1066) );
  XNOR U4078 ( .A(n1026), .B(n1066), .Z(n1044) );
  XOR U4079 ( .A(n1044), .B(n1029), .Z(n1031) );
  OR U4080 ( .A(n1031), .B(n1015), .Z(n1016) );
  XNOR U4081 ( .A(n1022), .B(n1016), .Z(n1048) );
  XOR U4082 ( .A(n1026), .B(n1072), .Z(n1034) );
  NANDN U4083 ( .A(n1034), .B(n1017), .Z(n1074) );
  NANDN U4084 ( .A(n1026), .B(n1018), .Z(n1019) );
  XNOR U4085 ( .A(n1074), .B(n1019), .Z(n1052) );
  XOR U4086 ( .A(n1048), .B(n1052), .Z(n1037) );
  NANDN U4087 ( .A(n1020), .B(n1044), .Z(n1021) );
  XNOR U4088 ( .A(n1022), .B(n1021), .Z(n1080) );
  XNOR U4089 ( .A(n1066), .B(n1054), .Z(n1056) );
  NANDN U4090 ( .A(n1056), .B(n1023), .Z(n1040) );
  NAND U4091 ( .A(n1024), .B(n1054), .Z(n1025) );
  XNOR U4092 ( .A(n1040), .B(n1025), .Z(n1071) );
  XOR U4093 ( .A(n1080), .B(n1071), .Z(n1063) );
  XNOR U4094 ( .A(n1037), .B(n1063), .Z(z[32]) );
  ANDN U4095 ( .B(n1027), .A(n1026), .Z(n1036) );
  NANDN U4096 ( .A(n1029), .B(n1028), .Z(n1047) );
  NANDN U4097 ( .A(n1031), .B(n1030), .Z(n1032) );
  XNOR U4098 ( .A(n1047), .B(n1032), .Z(n1075) );
  NANDN U4099 ( .A(n1034), .B(n1033), .Z(n1041) );
  XNOR U4100 ( .A(n1075), .B(n1041), .Z(n1035) );
  XOR U4101 ( .A(n1036), .B(n1035), .Z(n1061) );
  XOR U4102 ( .A(n1061), .B(n1037), .Z(n1079) );
  ANDN U4103 ( .B(n1072), .A(n1038), .Z(n1043) );
  NAND U4104 ( .A(n1064), .B(n1066), .Z(n1039) );
  XNOR U4105 ( .A(n1040), .B(n1039), .Z(n1051) );
  XNOR U4106 ( .A(n1041), .B(n1051), .Z(n1042) );
  XNOR U4107 ( .A(n1043), .B(n1042), .Z(n1050) );
  NAND U4108 ( .A(n1045), .B(n1044), .Z(n1046) );
  XNOR U4109 ( .A(n1047), .B(n1046), .Z(n1057) );
  XNOR U4110 ( .A(n1048), .B(n1057), .Z(n1049) );
  XOR U4111 ( .A(n1050), .B(n1049), .Z(n1060) );
  XNOR U4112 ( .A(n1079), .B(n1060), .Z(z[33]) );
  XNOR U4113 ( .A(n1052), .B(n1051), .Z(z[34]) );
  AND U4114 ( .A(n1054), .B(n1053), .Z(n1059) );
  NANDN U4115 ( .A(n1056), .B(n1055), .Z(n1069) );
  XNOR U4116 ( .A(n1057), .B(n1069), .Z(n1058) );
  XOR U4117 ( .A(n1059), .B(n1058), .Z(n1078) );
  XOR U4118 ( .A(n1061), .B(n1060), .Z(n1062) );
  XOR U4119 ( .A(n1078), .B(n1062), .Z(z[35]) );
  XOR U4120 ( .A(n1063), .B(z[34]), .Z(z[36]) );
  XNOR U4121 ( .A(n1065), .B(n1064), .Z(n1067) );
  NAND U4122 ( .A(n1067), .B(n1066), .Z(n1068) );
  XOR U4123 ( .A(n1069), .B(n1068), .Z(n1070) );
  XNOR U4124 ( .A(n1071), .B(n1070), .Z(n1077) );
  NAND U4125 ( .A(n1072), .B(x[32]), .Z(n1073) );
  XNOR U4126 ( .A(n1074), .B(n1073), .Z(n1081) );
  XNOR U4127 ( .A(n1075), .B(n1081), .Z(n1076) );
  XOR U4128 ( .A(n1077), .B(n1076), .Z(z[37]) );
  XNOR U4129 ( .A(n1079), .B(n1078), .Z(z[38]) );
  XNOR U4130 ( .A(n1081), .B(n1080), .Z(n1082) );
  XNOR U4131 ( .A(z[33]), .B(n1082), .Z(z[39]) );
  AND U4132 ( .A(n1084), .B(n1083), .Z(n1089) );
  NANDN U4133 ( .A(n1086), .B(n1085), .Z(n1451) );
  XNOR U4134 ( .A(n1087), .B(n1451), .Z(n1088) );
  XOR U4135 ( .A(n1089), .B(n1088), .Z(n1599) );
  XOR U4136 ( .A(n1091), .B(n1090), .Z(n1092) );
  XOR U4137 ( .A(n1599), .B(n1092), .Z(z[3]) );
  IV U4138 ( .A(x[41]), .Z(n1199) );
  XOR U4139 ( .A(x[40]), .B(x[46]), .Z(n1094) );
  XOR U4140 ( .A(x[45]), .B(n1094), .Z(n1198) );
  IV U4141 ( .A(n1198), .Z(n1095) );
  AND U4142 ( .A(n1199), .B(n1095), .Z(n1102) );
  XNOR U4143 ( .A(x[43]), .B(n1199), .Z(n1098) );
  XNOR U4144 ( .A(x[42]), .B(n1098), .Z(n1093) );
  XNOR U4145 ( .A(n1094), .B(n1093), .Z(n1158) );
  IV U4146 ( .A(n1158), .Z(n1104) );
  XNOR U4147 ( .A(n1104), .B(n1198), .Z(n1157) );
  IV U4148 ( .A(x[47]), .Z(n1096) );
  XNOR U4149 ( .A(x[41]), .B(n1096), .Z(n1189) );
  NAND U4150 ( .A(n1157), .B(n1189), .Z(n1107) );
  XNOR U4151 ( .A(n1096), .B(n1095), .Z(n1103) );
  IV U4152 ( .A(n1103), .Z(n1187) );
  XOR U4153 ( .A(n1158), .B(n1187), .Z(n1123) );
  XNOR U4154 ( .A(n1107), .B(n1123), .Z(n1100) );
  XOR U4155 ( .A(x[40]), .B(n1104), .Z(n1133) );
  XOR U4156 ( .A(x[44]), .B(n1096), .Z(n1097) );
  IV U4157 ( .A(n1097), .Z(n1162) );
  NANDN U4158 ( .A(n1133), .B(n1162), .Z(n1106) );
  XNOR U4159 ( .A(n1098), .B(n1097), .Z(n1151) );
  XNOR U4160 ( .A(n1157), .B(n1151), .Z(n1149) );
  XOR U4161 ( .A(x[42]), .B(x[44]), .Z(n1164) );
  NANDN U4162 ( .A(n1149), .B(n1164), .Z(n1099) );
  XOR U4163 ( .A(n1106), .B(n1099), .Z(n1125) );
  XNOR U4164 ( .A(n1100), .B(n1125), .Z(n1101) );
  XOR U4165 ( .A(n1102), .B(n1101), .Z(n1138) );
  IV U4166 ( .A(n1138), .Z(n1144) );
  AND U4167 ( .A(n1104), .B(n1103), .Z(n1109) );
  XOR U4168 ( .A(x[40]), .B(n1151), .Z(n1152) );
  XNOR U4169 ( .A(n1198), .B(n1152), .Z(n1154) );
  XOR U4170 ( .A(x[42]), .B(x[47]), .Z(n1179) );
  NANDN U4171 ( .A(n1154), .B(n1179), .Z(n1105) );
  XNOR U4172 ( .A(n1106), .B(n1105), .Z(n1114) );
  XNOR U4173 ( .A(n1107), .B(n1114), .Z(n1108) );
  XOR U4174 ( .A(n1109), .B(n1108), .Z(n1134) );
  XNOR U4175 ( .A(x[44]), .B(n1198), .Z(n1172) );
  ANDN U4176 ( .B(x[40]), .A(n1172), .Z(n1116) );
  XOR U4177 ( .A(x[42]), .B(x[41]), .Z(n1110) );
  XOR U4178 ( .A(n1187), .B(n1110), .Z(n1161) );
  XOR U4179 ( .A(n1162), .B(n1110), .Z(n1167) );
  NAND U4180 ( .A(n1151), .B(n1167), .Z(n1118) );
  XNOR U4181 ( .A(n1161), .B(n1118), .Z(n1112) );
  XNOR U4182 ( .A(x[41]), .B(n1152), .Z(n1111) );
  XNOR U4183 ( .A(n1112), .B(n1111), .Z(n1113) );
  XOR U4184 ( .A(n1114), .B(n1113), .Z(n1115) );
  XOR U4185 ( .A(n1116), .B(n1115), .Z(n1136) );
  NAND U4186 ( .A(n1134), .B(n1136), .Z(n1117) );
  NAND U4187 ( .A(n1144), .B(n1117), .Z(n1128) );
  IV U4188 ( .A(n1134), .Z(n1135) );
  IV U4189 ( .A(n1136), .Z(n1142) );
  XOR U4190 ( .A(n1118), .B(n1172), .Z(n1121) );
  AND U4191 ( .A(n1161), .B(n1152), .Z(n1119) );
  XNOR U4192 ( .A(x[40]), .B(n1119), .Z(n1120) );
  XNOR U4193 ( .A(n1121), .B(n1120), .Z(n1122) );
  XNOR U4194 ( .A(n1123), .B(n1122), .Z(n1124) );
  XNOR U4195 ( .A(n1125), .B(n1124), .Z(n1146) );
  IV U4196 ( .A(n1146), .Z(n1141) );
  XOR U4197 ( .A(n1142), .B(n1141), .Z(n1126) );
  NAND U4198 ( .A(n1135), .B(n1126), .Z(n1127) );
  AND U4199 ( .A(n1128), .B(n1127), .Z(n1206) );
  NAND U4200 ( .A(n1142), .B(n1135), .Z(n1129) );
  NAND U4201 ( .A(n1141), .B(n1129), .Z(n1132) );
  XOR U4202 ( .A(n1135), .B(n1138), .Z(n1130) );
  NAND U4203 ( .A(n1136), .B(n1130), .Z(n1131) );
  AND U4204 ( .A(n1132), .B(n1131), .Z(n1188) );
  XNOR U4205 ( .A(n1206), .B(n1188), .Z(n1163) );
  OR U4206 ( .A(n1163), .B(n1133), .Z(n1156) );
  NAND U4207 ( .A(n1144), .B(n1134), .Z(n1140) );
  AND U4208 ( .A(n1136), .B(n1135), .Z(n1143) );
  XNOR U4209 ( .A(n1141), .B(n1143), .Z(n1137) );
  NAND U4210 ( .A(n1138), .B(n1137), .Z(n1139) );
  AND U4211 ( .A(n1140), .B(n1139), .Z(n1160) );
  NAND U4212 ( .A(n1142), .B(n1141), .Z(n1148) );
  XNOR U4213 ( .A(n1144), .B(n1143), .Z(n1145) );
  NAND U4214 ( .A(n1146), .B(n1145), .Z(n1147) );
  NAND U4215 ( .A(n1148), .B(n1147), .Z(n1200) );
  XNOR U4216 ( .A(n1160), .B(n1200), .Z(n1178) );
  XOR U4217 ( .A(n1178), .B(n1163), .Z(n1165) );
  OR U4218 ( .A(n1165), .B(n1149), .Z(n1150) );
  XNOR U4219 ( .A(n1156), .B(n1150), .Z(n1182) );
  XOR U4220 ( .A(n1160), .B(n1206), .Z(n1168) );
  NANDN U4221 ( .A(n1168), .B(n1151), .Z(n1208) );
  NANDN U4222 ( .A(n1160), .B(n1152), .Z(n1153) );
  XNOR U4223 ( .A(n1208), .B(n1153), .Z(n1186) );
  XOR U4224 ( .A(n1182), .B(n1186), .Z(n1171) );
  NANDN U4225 ( .A(n1154), .B(n1178), .Z(n1155) );
  XNOR U4226 ( .A(n1156), .B(n1155), .Z(n1214) );
  XNOR U4227 ( .A(n1200), .B(n1188), .Z(n1190) );
  NANDN U4228 ( .A(n1190), .B(n1157), .Z(n1174) );
  NAND U4229 ( .A(n1158), .B(n1188), .Z(n1159) );
  XNOR U4230 ( .A(n1174), .B(n1159), .Z(n1205) );
  XOR U4231 ( .A(n1214), .B(n1205), .Z(n1197) );
  XNOR U4232 ( .A(n1171), .B(n1197), .Z(z[40]) );
  ANDN U4233 ( .B(n1161), .A(n1160), .Z(n1170) );
  NANDN U4234 ( .A(n1163), .B(n1162), .Z(n1181) );
  NANDN U4235 ( .A(n1165), .B(n1164), .Z(n1166) );
  XNOR U4236 ( .A(n1181), .B(n1166), .Z(n1209) );
  NANDN U4237 ( .A(n1168), .B(n1167), .Z(n1175) );
  XNOR U4238 ( .A(n1209), .B(n1175), .Z(n1169) );
  XOR U4239 ( .A(n1170), .B(n1169), .Z(n1195) );
  XOR U4240 ( .A(n1195), .B(n1171), .Z(n1213) );
  ANDN U4241 ( .B(n1206), .A(n1172), .Z(n1177) );
  NAND U4242 ( .A(n1198), .B(n1200), .Z(n1173) );
  XNOR U4243 ( .A(n1174), .B(n1173), .Z(n1185) );
  XNOR U4244 ( .A(n1175), .B(n1185), .Z(n1176) );
  XNOR U4245 ( .A(n1177), .B(n1176), .Z(n1184) );
  NAND U4246 ( .A(n1179), .B(n1178), .Z(n1180) );
  XNOR U4247 ( .A(n1181), .B(n1180), .Z(n1191) );
  XNOR U4248 ( .A(n1182), .B(n1191), .Z(n1183) );
  XOR U4249 ( .A(n1184), .B(n1183), .Z(n1194) );
  XNOR U4250 ( .A(n1213), .B(n1194), .Z(z[41]) );
  XNOR U4251 ( .A(n1186), .B(n1185), .Z(z[42]) );
  AND U4252 ( .A(n1188), .B(n1187), .Z(n1193) );
  NANDN U4253 ( .A(n1190), .B(n1189), .Z(n1203) );
  XNOR U4254 ( .A(n1191), .B(n1203), .Z(n1192) );
  XOR U4255 ( .A(n1193), .B(n1192), .Z(n1212) );
  XOR U4256 ( .A(n1195), .B(n1194), .Z(n1196) );
  XOR U4257 ( .A(n1212), .B(n1196), .Z(z[43]) );
  XOR U4258 ( .A(n1197), .B(z[42]), .Z(z[44]) );
  XNOR U4259 ( .A(n1199), .B(n1198), .Z(n1201) );
  NAND U4260 ( .A(n1201), .B(n1200), .Z(n1202) );
  XOR U4261 ( .A(n1203), .B(n1202), .Z(n1204) );
  XNOR U4262 ( .A(n1205), .B(n1204), .Z(n1211) );
  NAND U4263 ( .A(n1206), .B(x[40]), .Z(n1207) );
  XNOR U4264 ( .A(n1208), .B(n1207), .Z(n1215) );
  XNOR U4265 ( .A(n1209), .B(n1215), .Z(n1210) );
  XOR U4266 ( .A(n1211), .B(n1210), .Z(z[45]) );
  XNOR U4267 ( .A(n1213), .B(n1212), .Z(z[46]) );
  XNOR U4268 ( .A(n1215), .B(n1214), .Z(n1216) );
  XNOR U4269 ( .A(z[41]), .B(n1216), .Z(z[47]) );
  IV U4270 ( .A(x[49]), .Z(n1324) );
  XOR U4271 ( .A(x[48]), .B(x[54]), .Z(n1218) );
  XOR U4272 ( .A(x[53]), .B(n1218), .Z(n1323) );
  IV U4273 ( .A(n1323), .Z(n1219) );
  AND U4274 ( .A(n1324), .B(n1219), .Z(n1226) );
  XNOR U4275 ( .A(x[51]), .B(n1324), .Z(n1222) );
  XNOR U4276 ( .A(x[50]), .B(n1222), .Z(n1217) );
  XNOR U4277 ( .A(n1218), .B(n1217), .Z(n1282) );
  IV U4278 ( .A(n1282), .Z(n1228) );
  XNOR U4279 ( .A(n1228), .B(n1323), .Z(n1281) );
  IV U4280 ( .A(x[55]), .Z(n1220) );
  XNOR U4281 ( .A(x[49]), .B(n1220), .Z(n1314) );
  NAND U4282 ( .A(n1281), .B(n1314), .Z(n1231) );
  XNOR U4283 ( .A(n1220), .B(n1219), .Z(n1227) );
  IV U4284 ( .A(n1227), .Z(n1312) );
  XOR U4285 ( .A(n1282), .B(n1312), .Z(n1247) );
  XNOR U4286 ( .A(n1231), .B(n1247), .Z(n1224) );
  XOR U4287 ( .A(x[48]), .B(n1228), .Z(n1257) );
  XOR U4288 ( .A(x[52]), .B(n1220), .Z(n1221) );
  IV U4289 ( .A(n1221), .Z(n1286) );
  NANDN U4290 ( .A(n1257), .B(n1286), .Z(n1230) );
  XNOR U4291 ( .A(n1222), .B(n1221), .Z(n1275) );
  XNOR U4292 ( .A(n1281), .B(n1275), .Z(n1273) );
  XOR U4293 ( .A(x[50]), .B(x[52]), .Z(n1288) );
  NANDN U4294 ( .A(n1273), .B(n1288), .Z(n1223) );
  XOR U4295 ( .A(n1230), .B(n1223), .Z(n1249) );
  XNOR U4296 ( .A(n1224), .B(n1249), .Z(n1225) );
  XOR U4297 ( .A(n1226), .B(n1225), .Z(n1262) );
  IV U4298 ( .A(n1262), .Z(n1268) );
  AND U4299 ( .A(n1228), .B(n1227), .Z(n1233) );
  XOR U4300 ( .A(x[48]), .B(n1275), .Z(n1276) );
  XNOR U4301 ( .A(n1323), .B(n1276), .Z(n1278) );
  XOR U4302 ( .A(x[50]), .B(x[55]), .Z(n1303) );
  NANDN U4303 ( .A(n1278), .B(n1303), .Z(n1229) );
  XNOR U4304 ( .A(n1230), .B(n1229), .Z(n1238) );
  XNOR U4305 ( .A(n1231), .B(n1238), .Z(n1232) );
  XOR U4306 ( .A(n1233), .B(n1232), .Z(n1258) );
  XNOR U4307 ( .A(x[52]), .B(n1323), .Z(n1296) );
  ANDN U4308 ( .B(x[48]), .A(n1296), .Z(n1240) );
  XOR U4309 ( .A(x[50]), .B(x[49]), .Z(n1234) );
  XOR U4310 ( .A(n1312), .B(n1234), .Z(n1285) );
  XOR U4311 ( .A(n1286), .B(n1234), .Z(n1291) );
  NAND U4312 ( .A(n1275), .B(n1291), .Z(n1242) );
  XNOR U4313 ( .A(n1285), .B(n1242), .Z(n1236) );
  XNOR U4314 ( .A(x[49]), .B(n1276), .Z(n1235) );
  XNOR U4315 ( .A(n1236), .B(n1235), .Z(n1237) );
  XOR U4316 ( .A(n1238), .B(n1237), .Z(n1239) );
  XOR U4317 ( .A(n1240), .B(n1239), .Z(n1260) );
  NAND U4318 ( .A(n1258), .B(n1260), .Z(n1241) );
  NAND U4319 ( .A(n1268), .B(n1241), .Z(n1252) );
  IV U4320 ( .A(n1258), .Z(n1259) );
  IV U4321 ( .A(n1260), .Z(n1266) );
  XOR U4322 ( .A(n1242), .B(n1296), .Z(n1245) );
  AND U4323 ( .A(n1285), .B(n1276), .Z(n1243) );
  XNOR U4324 ( .A(x[48]), .B(n1243), .Z(n1244) );
  XNOR U4325 ( .A(n1245), .B(n1244), .Z(n1246) );
  XNOR U4326 ( .A(n1247), .B(n1246), .Z(n1248) );
  XNOR U4327 ( .A(n1249), .B(n1248), .Z(n1270) );
  IV U4328 ( .A(n1270), .Z(n1265) );
  XOR U4329 ( .A(n1266), .B(n1265), .Z(n1250) );
  NAND U4330 ( .A(n1259), .B(n1250), .Z(n1251) );
  AND U4331 ( .A(n1252), .B(n1251), .Z(n1331) );
  NAND U4332 ( .A(n1266), .B(n1259), .Z(n1253) );
  NAND U4333 ( .A(n1265), .B(n1253), .Z(n1256) );
  XOR U4334 ( .A(n1259), .B(n1262), .Z(n1254) );
  NAND U4335 ( .A(n1260), .B(n1254), .Z(n1255) );
  AND U4336 ( .A(n1256), .B(n1255), .Z(n1313) );
  XNOR U4337 ( .A(n1331), .B(n1313), .Z(n1287) );
  OR U4338 ( .A(n1287), .B(n1257), .Z(n1280) );
  NAND U4339 ( .A(n1268), .B(n1258), .Z(n1264) );
  AND U4340 ( .A(n1260), .B(n1259), .Z(n1267) );
  XNOR U4341 ( .A(n1265), .B(n1267), .Z(n1261) );
  NAND U4342 ( .A(n1262), .B(n1261), .Z(n1263) );
  AND U4343 ( .A(n1264), .B(n1263), .Z(n1284) );
  NAND U4344 ( .A(n1266), .B(n1265), .Z(n1272) );
  XNOR U4345 ( .A(n1268), .B(n1267), .Z(n1269) );
  NAND U4346 ( .A(n1270), .B(n1269), .Z(n1271) );
  NAND U4347 ( .A(n1272), .B(n1271), .Z(n1325) );
  XNOR U4348 ( .A(n1284), .B(n1325), .Z(n1302) );
  XOR U4349 ( .A(n1302), .B(n1287), .Z(n1289) );
  OR U4350 ( .A(n1289), .B(n1273), .Z(n1274) );
  XNOR U4351 ( .A(n1280), .B(n1274), .Z(n1306) );
  XOR U4352 ( .A(n1284), .B(n1331), .Z(n1292) );
  NANDN U4353 ( .A(n1292), .B(n1275), .Z(n1333) );
  NANDN U4354 ( .A(n1284), .B(n1276), .Z(n1277) );
  XNOR U4355 ( .A(n1333), .B(n1277), .Z(n1311) );
  XOR U4356 ( .A(n1306), .B(n1311), .Z(n1295) );
  NANDN U4357 ( .A(n1278), .B(n1302), .Z(n1279) );
  XNOR U4358 ( .A(n1280), .B(n1279), .Z(n1339) );
  XNOR U4359 ( .A(n1325), .B(n1313), .Z(n1315) );
  NANDN U4360 ( .A(n1315), .B(n1281), .Z(n1298) );
  NAND U4361 ( .A(n1282), .B(n1313), .Z(n1283) );
  XNOR U4362 ( .A(n1298), .B(n1283), .Z(n1330) );
  XOR U4363 ( .A(n1339), .B(n1330), .Z(n1322) );
  XNOR U4364 ( .A(n1295), .B(n1322), .Z(z[48]) );
  ANDN U4365 ( .B(n1285), .A(n1284), .Z(n1294) );
  NANDN U4366 ( .A(n1287), .B(n1286), .Z(n1305) );
  NANDN U4367 ( .A(n1289), .B(n1288), .Z(n1290) );
  XNOR U4368 ( .A(n1305), .B(n1290), .Z(n1334) );
  NANDN U4369 ( .A(n1292), .B(n1291), .Z(n1299) );
  XNOR U4370 ( .A(n1334), .B(n1299), .Z(n1293) );
  XOR U4371 ( .A(n1294), .B(n1293), .Z(n1320) );
  XOR U4372 ( .A(n1320), .B(n1295), .Z(n1338) );
  ANDN U4373 ( .B(n1331), .A(n1296), .Z(n1301) );
  NAND U4374 ( .A(n1323), .B(n1325), .Z(n1297) );
  XNOR U4375 ( .A(n1298), .B(n1297), .Z(n1310) );
  XNOR U4376 ( .A(n1299), .B(n1310), .Z(n1300) );
  XNOR U4377 ( .A(n1301), .B(n1300), .Z(n1308) );
  NAND U4378 ( .A(n1303), .B(n1302), .Z(n1304) );
  XNOR U4379 ( .A(n1305), .B(n1304), .Z(n1316) );
  XNOR U4380 ( .A(n1306), .B(n1316), .Z(n1307) );
  XOR U4381 ( .A(n1308), .B(n1307), .Z(n1319) );
  XNOR U4382 ( .A(n1338), .B(n1319), .Z(z[49]) );
  XOR U4383 ( .A(n1309), .B(z[2]), .Z(z[4]) );
  XNOR U4384 ( .A(n1311), .B(n1310), .Z(z[50]) );
  AND U4385 ( .A(n1313), .B(n1312), .Z(n1318) );
  NANDN U4386 ( .A(n1315), .B(n1314), .Z(n1328) );
  XNOR U4387 ( .A(n1316), .B(n1328), .Z(n1317) );
  XOR U4388 ( .A(n1318), .B(n1317), .Z(n1337) );
  XOR U4389 ( .A(n1320), .B(n1319), .Z(n1321) );
  XOR U4390 ( .A(n1337), .B(n1321), .Z(z[51]) );
  XOR U4391 ( .A(n1322), .B(z[50]), .Z(z[52]) );
  XNOR U4392 ( .A(n1324), .B(n1323), .Z(n1326) );
  NAND U4393 ( .A(n1326), .B(n1325), .Z(n1327) );
  XOR U4394 ( .A(n1328), .B(n1327), .Z(n1329) );
  XNOR U4395 ( .A(n1330), .B(n1329), .Z(n1336) );
  NAND U4396 ( .A(n1331), .B(x[48]), .Z(n1332) );
  XNOR U4397 ( .A(n1333), .B(n1332), .Z(n1340) );
  XNOR U4398 ( .A(n1334), .B(n1340), .Z(n1335) );
  XOR U4399 ( .A(n1336), .B(n1335), .Z(z[53]) );
  XNOR U4400 ( .A(n1338), .B(n1337), .Z(z[54]) );
  XNOR U4401 ( .A(n1340), .B(n1339), .Z(n1341) );
  XNOR U4402 ( .A(z[49]), .B(n1341), .Z(z[55]) );
  IV U4403 ( .A(x[57]), .Z(n1462) );
  XOR U4404 ( .A(x[56]), .B(x[62]), .Z(n1343) );
  XOR U4405 ( .A(x[61]), .B(n1343), .Z(n1461) );
  IV U4406 ( .A(n1461), .Z(n1344) );
  AND U4407 ( .A(n1462), .B(n1344), .Z(n1351) );
  XNOR U4408 ( .A(x[59]), .B(n1462), .Z(n1347) );
  XNOR U4409 ( .A(x[58]), .B(n1347), .Z(n1342) );
  XNOR U4410 ( .A(n1343), .B(n1342), .Z(n1407) );
  IV U4411 ( .A(n1407), .Z(n1353) );
  XNOR U4412 ( .A(n1353), .B(n1461), .Z(n1406) );
  IV U4413 ( .A(x[63]), .Z(n1345) );
  XNOR U4414 ( .A(x[57]), .B(n1345), .Z(n1438) );
  NAND U4415 ( .A(n1406), .B(n1438), .Z(n1356) );
  XNOR U4416 ( .A(n1345), .B(n1344), .Z(n1352) );
  IV U4417 ( .A(n1352), .Z(n1436) );
  XOR U4418 ( .A(n1407), .B(n1436), .Z(n1372) );
  XNOR U4419 ( .A(n1356), .B(n1372), .Z(n1349) );
  XOR U4420 ( .A(x[56]), .B(n1353), .Z(n1382) );
  XOR U4421 ( .A(x[60]), .B(n1345), .Z(n1346) );
  IV U4422 ( .A(n1346), .Z(n1411) );
  NANDN U4423 ( .A(n1382), .B(n1411), .Z(n1355) );
  XNOR U4424 ( .A(n1347), .B(n1346), .Z(n1400) );
  XNOR U4425 ( .A(n1406), .B(n1400), .Z(n1398) );
  XOR U4426 ( .A(x[58]), .B(x[60]), .Z(n1413) );
  NANDN U4427 ( .A(n1398), .B(n1413), .Z(n1348) );
  XOR U4428 ( .A(n1355), .B(n1348), .Z(n1374) );
  XNOR U4429 ( .A(n1349), .B(n1374), .Z(n1350) );
  XOR U4430 ( .A(n1351), .B(n1350), .Z(n1387) );
  IV U4431 ( .A(n1387), .Z(n1393) );
  AND U4432 ( .A(n1353), .B(n1352), .Z(n1358) );
  XOR U4433 ( .A(x[56]), .B(n1400), .Z(n1401) );
  XNOR U4434 ( .A(n1461), .B(n1401), .Z(n1403) );
  XOR U4435 ( .A(x[58]), .B(x[63]), .Z(n1428) );
  NANDN U4436 ( .A(n1403), .B(n1428), .Z(n1354) );
  XNOR U4437 ( .A(n1355), .B(n1354), .Z(n1363) );
  XNOR U4438 ( .A(n1356), .B(n1363), .Z(n1357) );
  XOR U4439 ( .A(n1358), .B(n1357), .Z(n1383) );
  XNOR U4440 ( .A(x[60]), .B(n1461), .Z(n1421) );
  ANDN U4441 ( .B(x[56]), .A(n1421), .Z(n1365) );
  XOR U4442 ( .A(x[58]), .B(x[57]), .Z(n1359) );
  XOR U4443 ( .A(n1436), .B(n1359), .Z(n1410) );
  XOR U4444 ( .A(n1411), .B(n1359), .Z(n1416) );
  NAND U4445 ( .A(n1400), .B(n1416), .Z(n1367) );
  XNOR U4446 ( .A(n1410), .B(n1367), .Z(n1361) );
  XNOR U4447 ( .A(x[57]), .B(n1401), .Z(n1360) );
  XNOR U4448 ( .A(n1361), .B(n1360), .Z(n1362) );
  XOR U4449 ( .A(n1363), .B(n1362), .Z(n1364) );
  XOR U4450 ( .A(n1365), .B(n1364), .Z(n1385) );
  NAND U4451 ( .A(n1383), .B(n1385), .Z(n1366) );
  NAND U4452 ( .A(n1393), .B(n1366), .Z(n1377) );
  IV U4453 ( .A(n1383), .Z(n1384) );
  IV U4454 ( .A(n1385), .Z(n1391) );
  XOR U4455 ( .A(n1367), .B(n1421), .Z(n1370) );
  AND U4456 ( .A(n1410), .B(n1401), .Z(n1368) );
  XNOR U4457 ( .A(x[56]), .B(n1368), .Z(n1369) );
  XNOR U4458 ( .A(n1370), .B(n1369), .Z(n1371) );
  XNOR U4459 ( .A(n1372), .B(n1371), .Z(n1373) );
  XNOR U4460 ( .A(n1374), .B(n1373), .Z(n1395) );
  IV U4461 ( .A(n1395), .Z(n1390) );
  XOR U4462 ( .A(n1391), .B(n1390), .Z(n1375) );
  NAND U4463 ( .A(n1384), .B(n1375), .Z(n1376) );
  AND U4464 ( .A(n1377), .B(n1376), .Z(n1469) );
  NAND U4465 ( .A(n1391), .B(n1384), .Z(n1378) );
  NAND U4466 ( .A(n1390), .B(n1378), .Z(n1381) );
  XOR U4467 ( .A(n1384), .B(n1387), .Z(n1379) );
  NAND U4468 ( .A(n1385), .B(n1379), .Z(n1380) );
  AND U4469 ( .A(n1381), .B(n1380), .Z(n1437) );
  XNOR U4470 ( .A(n1469), .B(n1437), .Z(n1412) );
  OR U4471 ( .A(n1412), .B(n1382), .Z(n1405) );
  NAND U4472 ( .A(n1393), .B(n1383), .Z(n1389) );
  AND U4473 ( .A(n1385), .B(n1384), .Z(n1392) );
  XNOR U4474 ( .A(n1390), .B(n1392), .Z(n1386) );
  NAND U4475 ( .A(n1387), .B(n1386), .Z(n1388) );
  AND U4476 ( .A(n1389), .B(n1388), .Z(n1409) );
  NAND U4477 ( .A(n1391), .B(n1390), .Z(n1397) );
  XNOR U4478 ( .A(n1393), .B(n1392), .Z(n1394) );
  NAND U4479 ( .A(n1395), .B(n1394), .Z(n1396) );
  NAND U4480 ( .A(n1397), .B(n1396), .Z(n1463) );
  XNOR U4481 ( .A(n1409), .B(n1463), .Z(n1427) );
  XOR U4482 ( .A(n1427), .B(n1412), .Z(n1414) );
  OR U4483 ( .A(n1414), .B(n1398), .Z(n1399) );
  XNOR U4484 ( .A(n1405), .B(n1399), .Z(n1431) );
  XOR U4485 ( .A(n1409), .B(n1469), .Z(n1417) );
  NANDN U4486 ( .A(n1417), .B(n1400), .Z(n1471) );
  NANDN U4487 ( .A(n1409), .B(n1401), .Z(n1402) );
  XNOR U4488 ( .A(n1471), .B(n1402), .Z(n1435) );
  XOR U4489 ( .A(n1431), .B(n1435), .Z(n1420) );
  NANDN U4490 ( .A(n1403), .B(n1427), .Z(n1404) );
  XNOR U4491 ( .A(n1405), .B(n1404), .Z(n1477) );
  XNOR U4492 ( .A(n1463), .B(n1437), .Z(n1439) );
  NANDN U4493 ( .A(n1439), .B(n1406), .Z(n1423) );
  NAND U4494 ( .A(n1407), .B(n1437), .Z(n1408) );
  XNOR U4495 ( .A(n1423), .B(n1408), .Z(n1468) );
  XOR U4496 ( .A(n1477), .B(n1468), .Z(n1460) );
  XNOR U4497 ( .A(n1420), .B(n1460), .Z(z[56]) );
  ANDN U4498 ( .B(n1410), .A(n1409), .Z(n1419) );
  NANDN U4499 ( .A(n1412), .B(n1411), .Z(n1430) );
  NANDN U4500 ( .A(n1414), .B(n1413), .Z(n1415) );
  XNOR U4501 ( .A(n1430), .B(n1415), .Z(n1472) );
  NANDN U4502 ( .A(n1417), .B(n1416), .Z(n1424) );
  XNOR U4503 ( .A(n1472), .B(n1424), .Z(n1418) );
  XOR U4504 ( .A(n1419), .B(n1418), .Z(n1444) );
  XOR U4505 ( .A(n1444), .B(n1420), .Z(n1476) );
  ANDN U4506 ( .B(n1469), .A(n1421), .Z(n1426) );
  NAND U4507 ( .A(n1461), .B(n1463), .Z(n1422) );
  XNOR U4508 ( .A(n1423), .B(n1422), .Z(n1434) );
  XNOR U4509 ( .A(n1424), .B(n1434), .Z(n1425) );
  XNOR U4510 ( .A(n1426), .B(n1425), .Z(n1433) );
  NAND U4511 ( .A(n1428), .B(n1427), .Z(n1429) );
  XNOR U4512 ( .A(n1430), .B(n1429), .Z(n1440) );
  XNOR U4513 ( .A(n1431), .B(n1440), .Z(n1432) );
  XOR U4514 ( .A(n1433), .B(n1432), .Z(n1443) );
  XNOR U4515 ( .A(n1476), .B(n1443), .Z(z[57]) );
  XNOR U4516 ( .A(n1435), .B(n1434), .Z(z[58]) );
  AND U4517 ( .A(n1437), .B(n1436), .Z(n1442) );
  NANDN U4518 ( .A(n1439), .B(n1438), .Z(n1466) );
  XNOR U4519 ( .A(n1440), .B(n1466), .Z(n1441) );
  XOR U4520 ( .A(n1442), .B(n1441), .Z(n1475) );
  XOR U4521 ( .A(n1444), .B(n1443), .Z(n1445) );
  XOR U4522 ( .A(n1475), .B(n1445), .Z(z[59]) );
  XNOR U4523 ( .A(n1447), .B(n1446), .Z(n1449) );
  NAND U4524 ( .A(n1449), .B(n1448), .Z(n1450) );
  XOR U4525 ( .A(n1451), .B(n1450), .Z(n1452) );
  XNOR U4526 ( .A(n1453), .B(n1452), .Z(n1459) );
  NAND U4527 ( .A(n1454), .B(x[0]), .Z(n1455) );
  XNOR U4528 ( .A(n1456), .B(n1455), .Z(n1731) );
  XNOR U4529 ( .A(n1457), .B(n1731), .Z(n1458) );
  XOR U4530 ( .A(n1459), .B(n1458), .Z(z[5]) );
  XOR U4531 ( .A(n1460), .B(z[58]), .Z(z[60]) );
  XNOR U4532 ( .A(n1462), .B(n1461), .Z(n1464) );
  NAND U4533 ( .A(n1464), .B(n1463), .Z(n1465) );
  XOR U4534 ( .A(n1466), .B(n1465), .Z(n1467) );
  XNOR U4535 ( .A(n1468), .B(n1467), .Z(n1474) );
  NAND U4536 ( .A(n1469), .B(x[56]), .Z(n1470) );
  XNOR U4537 ( .A(n1471), .B(n1470), .Z(n1478) );
  XNOR U4538 ( .A(n1472), .B(n1478), .Z(n1473) );
  XOR U4539 ( .A(n1474), .B(n1473), .Z(z[61]) );
  XNOR U4540 ( .A(n1476), .B(n1475), .Z(z[62]) );
  XNOR U4541 ( .A(n1478), .B(n1477), .Z(n1479) );
  XNOR U4542 ( .A(z[57]), .B(n1479), .Z(z[63]) );
  IV U4543 ( .A(x[65]), .Z(n1586) );
  XOR U4544 ( .A(x[64]), .B(x[70]), .Z(n1481) );
  XOR U4545 ( .A(x[69]), .B(n1481), .Z(n1585) );
  IV U4546 ( .A(n1585), .Z(n1482) );
  AND U4547 ( .A(n1586), .B(n1482), .Z(n1489) );
  XNOR U4548 ( .A(x[67]), .B(n1586), .Z(n1485) );
  XNOR U4549 ( .A(x[66]), .B(n1485), .Z(n1480) );
  XNOR U4550 ( .A(n1481), .B(n1480), .Z(n1545) );
  IV U4551 ( .A(n1545), .Z(n1491) );
  XNOR U4552 ( .A(n1491), .B(n1585), .Z(n1544) );
  IV U4553 ( .A(x[71]), .Z(n1483) );
  XNOR U4554 ( .A(x[65]), .B(n1483), .Z(n1576) );
  NAND U4555 ( .A(n1544), .B(n1576), .Z(n1494) );
  XNOR U4556 ( .A(n1483), .B(n1482), .Z(n1490) );
  IV U4557 ( .A(n1490), .Z(n1574) );
  XOR U4558 ( .A(n1545), .B(n1574), .Z(n1510) );
  XNOR U4559 ( .A(n1494), .B(n1510), .Z(n1487) );
  XOR U4560 ( .A(x[64]), .B(n1491), .Z(n1520) );
  XOR U4561 ( .A(x[68]), .B(n1483), .Z(n1484) );
  IV U4562 ( .A(n1484), .Z(n1549) );
  NANDN U4563 ( .A(n1520), .B(n1549), .Z(n1493) );
  XNOR U4564 ( .A(n1485), .B(n1484), .Z(n1538) );
  XNOR U4565 ( .A(n1544), .B(n1538), .Z(n1536) );
  XOR U4566 ( .A(x[66]), .B(x[68]), .Z(n1551) );
  NANDN U4567 ( .A(n1536), .B(n1551), .Z(n1486) );
  XOR U4568 ( .A(n1493), .B(n1486), .Z(n1512) );
  XNOR U4569 ( .A(n1487), .B(n1512), .Z(n1488) );
  XOR U4570 ( .A(n1489), .B(n1488), .Z(n1525) );
  IV U4571 ( .A(n1525), .Z(n1531) );
  AND U4572 ( .A(n1491), .B(n1490), .Z(n1496) );
  XOR U4573 ( .A(x[64]), .B(n1538), .Z(n1539) );
  XNOR U4574 ( .A(n1585), .B(n1539), .Z(n1541) );
  XOR U4575 ( .A(x[66]), .B(x[71]), .Z(n1566) );
  NANDN U4576 ( .A(n1541), .B(n1566), .Z(n1492) );
  XNOR U4577 ( .A(n1493), .B(n1492), .Z(n1501) );
  XNOR U4578 ( .A(n1494), .B(n1501), .Z(n1495) );
  XOR U4579 ( .A(n1496), .B(n1495), .Z(n1521) );
  XNOR U4580 ( .A(x[68]), .B(n1585), .Z(n1559) );
  ANDN U4581 ( .B(x[64]), .A(n1559), .Z(n1503) );
  XOR U4582 ( .A(x[66]), .B(x[65]), .Z(n1497) );
  XOR U4583 ( .A(n1574), .B(n1497), .Z(n1548) );
  XOR U4584 ( .A(n1549), .B(n1497), .Z(n1554) );
  NAND U4585 ( .A(n1538), .B(n1554), .Z(n1505) );
  XNOR U4586 ( .A(n1548), .B(n1505), .Z(n1499) );
  XNOR U4587 ( .A(x[65]), .B(n1539), .Z(n1498) );
  XNOR U4588 ( .A(n1499), .B(n1498), .Z(n1500) );
  XOR U4589 ( .A(n1501), .B(n1500), .Z(n1502) );
  XOR U4590 ( .A(n1503), .B(n1502), .Z(n1523) );
  NAND U4591 ( .A(n1521), .B(n1523), .Z(n1504) );
  NAND U4592 ( .A(n1531), .B(n1504), .Z(n1515) );
  IV U4593 ( .A(n1521), .Z(n1522) );
  IV U4594 ( .A(n1523), .Z(n1529) );
  XOR U4595 ( .A(n1505), .B(n1559), .Z(n1508) );
  AND U4596 ( .A(n1548), .B(n1539), .Z(n1506) );
  XNOR U4597 ( .A(x[64]), .B(n1506), .Z(n1507) );
  XNOR U4598 ( .A(n1508), .B(n1507), .Z(n1509) );
  XNOR U4599 ( .A(n1510), .B(n1509), .Z(n1511) );
  XNOR U4600 ( .A(n1512), .B(n1511), .Z(n1533) );
  IV U4601 ( .A(n1533), .Z(n1528) );
  XOR U4602 ( .A(n1529), .B(n1528), .Z(n1513) );
  NAND U4603 ( .A(n1522), .B(n1513), .Z(n1514) );
  AND U4604 ( .A(n1515), .B(n1514), .Z(n1593) );
  NAND U4605 ( .A(n1529), .B(n1522), .Z(n1516) );
  NAND U4606 ( .A(n1528), .B(n1516), .Z(n1519) );
  XOR U4607 ( .A(n1522), .B(n1525), .Z(n1517) );
  NAND U4608 ( .A(n1523), .B(n1517), .Z(n1518) );
  AND U4609 ( .A(n1519), .B(n1518), .Z(n1575) );
  XNOR U4610 ( .A(n1593), .B(n1575), .Z(n1550) );
  OR U4611 ( .A(n1550), .B(n1520), .Z(n1543) );
  NAND U4612 ( .A(n1531), .B(n1521), .Z(n1527) );
  AND U4613 ( .A(n1523), .B(n1522), .Z(n1530) );
  XNOR U4614 ( .A(n1528), .B(n1530), .Z(n1524) );
  NAND U4615 ( .A(n1525), .B(n1524), .Z(n1526) );
  AND U4616 ( .A(n1527), .B(n1526), .Z(n1547) );
  NAND U4617 ( .A(n1529), .B(n1528), .Z(n1535) );
  XNOR U4618 ( .A(n1531), .B(n1530), .Z(n1532) );
  NAND U4619 ( .A(n1533), .B(n1532), .Z(n1534) );
  NAND U4620 ( .A(n1535), .B(n1534), .Z(n1587) );
  XNOR U4621 ( .A(n1547), .B(n1587), .Z(n1565) );
  XOR U4622 ( .A(n1565), .B(n1550), .Z(n1552) );
  OR U4623 ( .A(n1552), .B(n1536), .Z(n1537) );
  XNOR U4624 ( .A(n1543), .B(n1537), .Z(n1569) );
  XOR U4625 ( .A(n1547), .B(n1593), .Z(n1555) );
  NANDN U4626 ( .A(n1555), .B(n1538), .Z(n1595) );
  NANDN U4627 ( .A(n1547), .B(n1539), .Z(n1540) );
  XNOR U4628 ( .A(n1595), .B(n1540), .Z(n1573) );
  XOR U4629 ( .A(n1569), .B(n1573), .Z(n1558) );
  NANDN U4630 ( .A(n1541), .B(n1565), .Z(n1542) );
  XNOR U4631 ( .A(n1543), .B(n1542), .Z(n1603) );
  XNOR U4632 ( .A(n1587), .B(n1575), .Z(n1577) );
  NANDN U4633 ( .A(n1577), .B(n1544), .Z(n1561) );
  NAND U4634 ( .A(n1545), .B(n1575), .Z(n1546) );
  XNOR U4635 ( .A(n1561), .B(n1546), .Z(n1592) );
  XOR U4636 ( .A(n1603), .B(n1592), .Z(n1584) );
  XNOR U4637 ( .A(n1558), .B(n1584), .Z(z[64]) );
  ANDN U4638 ( .B(n1548), .A(n1547), .Z(n1557) );
  NANDN U4639 ( .A(n1550), .B(n1549), .Z(n1568) );
  NANDN U4640 ( .A(n1552), .B(n1551), .Z(n1553) );
  XNOR U4641 ( .A(n1568), .B(n1553), .Z(n1596) );
  NANDN U4642 ( .A(n1555), .B(n1554), .Z(n1562) );
  XNOR U4643 ( .A(n1596), .B(n1562), .Z(n1556) );
  XOR U4644 ( .A(n1557), .B(n1556), .Z(n1582) );
  XOR U4645 ( .A(n1582), .B(n1558), .Z(n1602) );
  ANDN U4646 ( .B(n1593), .A(n1559), .Z(n1564) );
  NAND U4647 ( .A(n1585), .B(n1587), .Z(n1560) );
  XNOR U4648 ( .A(n1561), .B(n1560), .Z(n1572) );
  XNOR U4649 ( .A(n1562), .B(n1572), .Z(n1563) );
  XNOR U4650 ( .A(n1564), .B(n1563), .Z(n1571) );
  NAND U4651 ( .A(n1566), .B(n1565), .Z(n1567) );
  XNOR U4652 ( .A(n1568), .B(n1567), .Z(n1578) );
  XNOR U4653 ( .A(n1569), .B(n1578), .Z(n1570) );
  XOR U4654 ( .A(n1571), .B(n1570), .Z(n1581) );
  XNOR U4655 ( .A(n1602), .B(n1581), .Z(z[65]) );
  XNOR U4656 ( .A(n1573), .B(n1572), .Z(z[66]) );
  AND U4657 ( .A(n1575), .B(n1574), .Z(n1580) );
  NANDN U4658 ( .A(n1577), .B(n1576), .Z(n1590) );
  XNOR U4659 ( .A(n1578), .B(n1590), .Z(n1579) );
  XOR U4660 ( .A(n1580), .B(n1579), .Z(n1601) );
  XOR U4661 ( .A(n1582), .B(n1581), .Z(n1583) );
  XOR U4662 ( .A(n1601), .B(n1583), .Z(z[67]) );
  XOR U4663 ( .A(n1584), .B(z[66]), .Z(z[68]) );
  XNOR U4664 ( .A(n1586), .B(n1585), .Z(n1588) );
  NAND U4665 ( .A(n1588), .B(n1587), .Z(n1589) );
  XOR U4666 ( .A(n1590), .B(n1589), .Z(n1591) );
  XNOR U4667 ( .A(n1592), .B(n1591), .Z(n1598) );
  NAND U4668 ( .A(n1593), .B(x[64]), .Z(n1594) );
  XNOR U4669 ( .A(n1595), .B(n1594), .Z(n1604) );
  XNOR U4670 ( .A(n1596), .B(n1604), .Z(n1597) );
  XOR U4671 ( .A(n1598), .B(n1597), .Z(z[69]) );
  XNOR U4672 ( .A(n1600), .B(n1599), .Z(z[6]) );
  XNOR U4673 ( .A(n1602), .B(n1601), .Z(z[70]) );
  XNOR U4674 ( .A(n1604), .B(n1603), .Z(n1605) );
  XNOR U4675 ( .A(z[65]), .B(n1605), .Z(z[71]) );
  IV U4676 ( .A(x[73]), .Z(n1712) );
  XOR U4677 ( .A(x[72]), .B(x[78]), .Z(n1607) );
  XOR U4678 ( .A(x[77]), .B(n1607), .Z(n1711) );
  IV U4679 ( .A(n1711), .Z(n1608) );
  AND U4680 ( .A(n1712), .B(n1608), .Z(n1615) );
  XNOR U4681 ( .A(x[75]), .B(n1712), .Z(n1611) );
  XNOR U4682 ( .A(x[74]), .B(n1611), .Z(n1606) );
  XNOR U4683 ( .A(n1607), .B(n1606), .Z(n1671) );
  IV U4684 ( .A(n1671), .Z(n1617) );
  XNOR U4685 ( .A(n1617), .B(n1711), .Z(n1670) );
  IV U4686 ( .A(x[79]), .Z(n1609) );
  XNOR U4687 ( .A(x[73]), .B(n1609), .Z(n1702) );
  NAND U4688 ( .A(n1670), .B(n1702), .Z(n1620) );
  XNOR U4689 ( .A(n1609), .B(n1608), .Z(n1616) );
  IV U4690 ( .A(n1616), .Z(n1700) );
  XOR U4691 ( .A(n1671), .B(n1700), .Z(n1636) );
  XNOR U4692 ( .A(n1620), .B(n1636), .Z(n1613) );
  XOR U4693 ( .A(x[72]), .B(n1617), .Z(n1646) );
  XOR U4694 ( .A(x[76]), .B(n1609), .Z(n1610) );
  IV U4695 ( .A(n1610), .Z(n1675) );
  NANDN U4696 ( .A(n1646), .B(n1675), .Z(n1619) );
  XNOR U4697 ( .A(n1611), .B(n1610), .Z(n1664) );
  XNOR U4698 ( .A(n1670), .B(n1664), .Z(n1662) );
  XOR U4699 ( .A(x[74]), .B(x[76]), .Z(n1677) );
  NANDN U4700 ( .A(n1662), .B(n1677), .Z(n1612) );
  XOR U4701 ( .A(n1619), .B(n1612), .Z(n1638) );
  XNOR U4702 ( .A(n1613), .B(n1638), .Z(n1614) );
  XOR U4703 ( .A(n1615), .B(n1614), .Z(n1651) );
  IV U4704 ( .A(n1651), .Z(n1657) );
  AND U4705 ( .A(n1617), .B(n1616), .Z(n1622) );
  XOR U4706 ( .A(x[72]), .B(n1664), .Z(n1665) );
  XNOR U4707 ( .A(n1711), .B(n1665), .Z(n1667) );
  XOR U4708 ( .A(x[74]), .B(x[79]), .Z(n1692) );
  NANDN U4709 ( .A(n1667), .B(n1692), .Z(n1618) );
  XNOR U4710 ( .A(n1619), .B(n1618), .Z(n1627) );
  XNOR U4711 ( .A(n1620), .B(n1627), .Z(n1621) );
  XOR U4712 ( .A(n1622), .B(n1621), .Z(n1647) );
  XNOR U4713 ( .A(x[76]), .B(n1711), .Z(n1685) );
  ANDN U4714 ( .B(x[72]), .A(n1685), .Z(n1629) );
  XOR U4715 ( .A(x[74]), .B(x[73]), .Z(n1623) );
  XOR U4716 ( .A(n1700), .B(n1623), .Z(n1674) );
  XOR U4717 ( .A(n1675), .B(n1623), .Z(n1680) );
  NAND U4718 ( .A(n1664), .B(n1680), .Z(n1631) );
  XNOR U4719 ( .A(n1674), .B(n1631), .Z(n1625) );
  XNOR U4720 ( .A(x[73]), .B(n1665), .Z(n1624) );
  XNOR U4721 ( .A(n1625), .B(n1624), .Z(n1626) );
  XOR U4722 ( .A(n1627), .B(n1626), .Z(n1628) );
  XOR U4723 ( .A(n1629), .B(n1628), .Z(n1649) );
  NAND U4724 ( .A(n1647), .B(n1649), .Z(n1630) );
  NAND U4725 ( .A(n1657), .B(n1630), .Z(n1641) );
  IV U4726 ( .A(n1647), .Z(n1648) );
  IV U4727 ( .A(n1649), .Z(n1655) );
  XOR U4728 ( .A(n1631), .B(n1685), .Z(n1634) );
  AND U4729 ( .A(n1674), .B(n1665), .Z(n1632) );
  XNOR U4730 ( .A(x[72]), .B(n1632), .Z(n1633) );
  XNOR U4731 ( .A(n1634), .B(n1633), .Z(n1635) );
  XNOR U4732 ( .A(n1636), .B(n1635), .Z(n1637) );
  XNOR U4733 ( .A(n1638), .B(n1637), .Z(n1659) );
  IV U4734 ( .A(n1659), .Z(n1654) );
  XOR U4735 ( .A(n1655), .B(n1654), .Z(n1639) );
  NAND U4736 ( .A(n1648), .B(n1639), .Z(n1640) );
  AND U4737 ( .A(n1641), .B(n1640), .Z(n1719) );
  NAND U4738 ( .A(n1655), .B(n1648), .Z(n1642) );
  NAND U4739 ( .A(n1654), .B(n1642), .Z(n1645) );
  XOR U4740 ( .A(n1648), .B(n1651), .Z(n1643) );
  NAND U4741 ( .A(n1649), .B(n1643), .Z(n1644) );
  AND U4742 ( .A(n1645), .B(n1644), .Z(n1701) );
  XNOR U4743 ( .A(n1719), .B(n1701), .Z(n1676) );
  OR U4744 ( .A(n1676), .B(n1646), .Z(n1669) );
  NAND U4745 ( .A(n1657), .B(n1647), .Z(n1653) );
  AND U4746 ( .A(n1649), .B(n1648), .Z(n1656) );
  XNOR U4747 ( .A(n1654), .B(n1656), .Z(n1650) );
  NAND U4748 ( .A(n1651), .B(n1650), .Z(n1652) );
  AND U4749 ( .A(n1653), .B(n1652), .Z(n1673) );
  NAND U4750 ( .A(n1655), .B(n1654), .Z(n1661) );
  XNOR U4751 ( .A(n1657), .B(n1656), .Z(n1658) );
  NAND U4752 ( .A(n1659), .B(n1658), .Z(n1660) );
  NAND U4753 ( .A(n1661), .B(n1660), .Z(n1713) );
  XNOR U4754 ( .A(n1673), .B(n1713), .Z(n1691) );
  XOR U4755 ( .A(n1691), .B(n1676), .Z(n1678) );
  OR U4756 ( .A(n1678), .B(n1662), .Z(n1663) );
  XNOR U4757 ( .A(n1669), .B(n1663), .Z(n1695) );
  XOR U4758 ( .A(n1673), .B(n1719), .Z(n1681) );
  NANDN U4759 ( .A(n1681), .B(n1664), .Z(n1721) );
  NANDN U4760 ( .A(n1673), .B(n1665), .Z(n1666) );
  XNOR U4761 ( .A(n1721), .B(n1666), .Z(n1699) );
  XOR U4762 ( .A(n1695), .B(n1699), .Z(n1684) );
  NANDN U4763 ( .A(n1667), .B(n1691), .Z(n1668) );
  XNOR U4764 ( .A(n1669), .B(n1668), .Z(n1727) );
  XNOR U4765 ( .A(n1713), .B(n1701), .Z(n1703) );
  NANDN U4766 ( .A(n1703), .B(n1670), .Z(n1687) );
  NAND U4767 ( .A(n1671), .B(n1701), .Z(n1672) );
  XNOR U4768 ( .A(n1687), .B(n1672), .Z(n1718) );
  XOR U4769 ( .A(n1727), .B(n1718), .Z(n1710) );
  XNOR U4770 ( .A(n1684), .B(n1710), .Z(z[72]) );
  ANDN U4771 ( .B(n1674), .A(n1673), .Z(n1683) );
  NANDN U4772 ( .A(n1676), .B(n1675), .Z(n1694) );
  NANDN U4773 ( .A(n1678), .B(n1677), .Z(n1679) );
  XNOR U4774 ( .A(n1694), .B(n1679), .Z(n1722) );
  NANDN U4775 ( .A(n1681), .B(n1680), .Z(n1688) );
  XNOR U4776 ( .A(n1722), .B(n1688), .Z(n1682) );
  XOR U4777 ( .A(n1683), .B(n1682), .Z(n1708) );
  XOR U4778 ( .A(n1708), .B(n1684), .Z(n1726) );
  ANDN U4779 ( .B(n1719), .A(n1685), .Z(n1690) );
  NAND U4780 ( .A(n1711), .B(n1713), .Z(n1686) );
  XNOR U4781 ( .A(n1687), .B(n1686), .Z(n1698) );
  XNOR U4782 ( .A(n1688), .B(n1698), .Z(n1689) );
  XNOR U4783 ( .A(n1690), .B(n1689), .Z(n1697) );
  NAND U4784 ( .A(n1692), .B(n1691), .Z(n1693) );
  XNOR U4785 ( .A(n1694), .B(n1693), .Z(n1704) );
  XNOR U4786 ( .A(n1695), .B(n1704), .Z(n1696) );
  XOR U4787 ( .A(n1697), .B(n1696), .Z(n1707) );
  XNOR U4788 ( .A(n1726), .B(n1707), .Z(z[73]) );
  XNOR U4789 ( .A(n1699), .B(n1698), .Z(z[74]) );
  AND U4790 ( .A(n1701), .B(n1700), .Z(n1706) );
  NANDN U4791 ( .A(n1703), .B(n1702), .Z(n1716) );
  XNOR U4792 ( .A(n1704), .B(n1716), .Z(n1705) );
  XOR U4793 ( .A(n1706), .B(n1705), .Z(n1725) );
  XOR U4794 ( .A(n1708), .B(n1707), .Z(n1709) );
  XOR U4795 ( .A(n1725), .B(n1709), .Z(z[75]) );
  XOR U4796 ( .A(n1710), .B(z[74]), .Z(z[76]) );
  XNOR U4797 ( .A(n1712), .B(n1711), .Z(n1714) );
  NAND U4798 ( .A(n1714), .B(n1713), .Z(n1715) );
  XOR U4799 ( .A(n1716), .B(n1715), .Z(n1717) );
  XNOR U4800 ( .A(n1718), .B(n1717), .Z(n1724) );
  NAND U4801 ( .A(n1719), .B(x[72]), .Z(n1720) );
  XNOR U4802 ( .A(n1721), .B(n1720), .Z(n1728) );
  XNOR U4803 ( .A(n1722), .B(n1728), .Z(n1723) );
  XOR U4804 ( .A(n1724), .B(n1723), .Z(z[77]) );
  XNOR U4805 ( .A(n1726), .B(n1725), .Z(z[78]) );
  XNOR U4806 ( .A(n1728), .B(n1727), .Z(n1729) );
  XNOR U4807 ( .A(z[73]), .B(n1729), .Z(z[79]) );
  XNOR U4808 ( .A(n1731), .B(n1730), .Z(n1732) );
  XNOR U4809 ( .A(z[1]), .B(n1732), .Z(z[7]) );
  XOR U4810 ( .A(x[80]), .B(x[86]), .Z(n1733) );
  XOR U4811 ( .A(x[85]), .B(n1733), .Z(n1838) );
  IV U4812 ( .A(n1838), .Z(n1735) );
  IV U4813 ( .A(x[81]), .Z(n1837) );
  NAND U4814 ( .A(n1735), .B(n1837), .Z(n1742) );
  XOR U4815 ( .A(x[83]), .B(x[81]), .Z(n1738) );
  XNOR U4816 ( .A(x[82]), .B(n1733), .Z(n1734) );
  XNOR U4817 ( .A(n1738), .B(n1734), .Z(n1797) );
  XNOR U4818 ( .A(n1735), .B(n1797), .Z(n1796) );
  IV U4819 ( .A(x[87]), .Z(n1736) );
  XNOR U4820 ( .A(x[81]), .B(n1736), .Z(n1828) );
  NAND U4821 ( .A(n1796), .B(n1828), .Z(n1745) );
  XNOR U4822 ( .A(n1735), .B(n1736), .Z(n1826) );
  XOR U4823 ( .A(n1797), .B(n1826), .Z(n1753) );
  XOR U4824 ( .A(n1745), .B(n1753), .Z(n1740) );
  XNOR U4825 ( .A(x[80]), .B(n1797), .Z(n1772) );
  XOR U4826 ( .A(x[84]), .B(n1736), .Z(n1737) );
  IV U4827 ( .A(n1737), .Z(n1801) );
  NANDN U4828 ( .A(n1772), .B(n1801), .Z(n1744) );
  XOR U4829 ( .A(n1738), .B(n1737), .Z(n1790) );
  XOR U4830 ( .A(n1796), .B(n1790), .Z(n1788) );
  XOR U4831 ( .A(x[82]), .B(x[84]), .Z(n1803) );
  NANDN U4832 ( .A(n1788), .B(n1803), .Z(n1739) );
  XNOR U4833 ( .A(n1744), .B(n1739), .Z(n1749) );
  XOR U4834 ( .A(n1740), .B(n1749), .Z(n1741) );
  XOR U4835 ( .A(n1742), .B(n1741), .Z(n1783) );
  IV U4836 ( .A(n1783), .Z(n1777) );
  ANDN U4837 ( .B(n1826), .A(n1797), .Z(n1747) );
  XNOR U4838 ( .A(x[80]), .B(n1790), .Z(n1791) );
  XNOR U4839 ( .A(n1838), .B(n1791), .Z(n1793) );
  XOR U4840 ( .A(x[82]), .B(x[87]), .Z(n1818) );
  NANDN U4841 ( .A(n1793), .B(n1818), .Z(n1743) );
  XNOR U4842 ( .A(n1744), .B(n1743), .Z(n1760) );
  XNOR U4843 ( .A(n1745), .B(n1760), .Z(n1746) );
  XOR U4844 ( .A(n1747), .B(n1746), .Z(n1773) );
  NAND U4845 ( .A(n1777), .B(n1773), .Z(n1767) );
  IV U4846 ( .A(n1773), .Z(n1774) );
  XOR U4847 ( .A(n1783), .B(n1774), .Z(n1765) );
  XOR U4848 ( .A(x[82]), .B(x[81]), .Z(n1748) );
  XNOR U4849 ( .A(n1826), .B(n1748), .Z(n1800) );
  NAND U4850 ( .A(n1800), .B(n1791), .Z(n1755) );
  XNOR U4851 ( .A(x[84]), .B(n1838), .Z(n1811) );
  XOR U4852 ( .A(n1801), .B(n1748), .Z(n1806) );
  NANDN U4853 ( .A(n1790), .B(n1806), .Z(n1756) );
  XOR U4854 ( .A(n1811), .B(n1756), .Z(n1751) );
  XOR U4855 ( .A(x[80]), .B(n1749), .Z(n1750) );
  XNOR U4856 ( .A(n1751), .B(n1750), .Z(n1752) );
  XOR U4857 ( .A(n1753), .B(n1752), .Z(n1754) );
  XOR U4858 ( .A(n1755), .B(n1754), .Z(n1785) );
  IV U4859 ( .A(n1785), .Z(n1780) );
  AND U4860 ( .A(n1777), .B(n1780), .Z(n1763) );
  ANDN U4861 ( .B(x[80]), .A(n1811), .Z(n1762) );
  XNOR U4862 ( .A(n1800), .B(n1756), .Z(n1758) );
  XNOR U4863 ( .A(x[81]), .B(n1791), .Z(n1757) );
  XNOR U4864 ( .A(n1758), .B(n1757), .Z(n1759) );
  XOR U4865 ( .A(n1760), .B(n1759), .Z(n1761) );
  XOR U4866 ( .A(n1762), .B(n1761), .Z(n1775) );
  IV U4867 ( .A(n1775), .Z(n1781) );
  XNOR U4868 ( .A(n1763), .B(n1781), .Z(n1764) );
  NAND U4869 ( .A(n1765), .B(n1764), .Z(n1766) );
  NAND U4870 ( .A(n1767), .B(n1766), .Z(n1845) );
  NAND U4871 ( .A(n1781), .B(n1774), .Z(n1768) );
  NAND U4872 ( .A(n1780), .B(n1768), .Z(n1771) );
  XOR U4873 ( .A(n1774), .B(n1777), .Z(n1769) );
  NAND U4874 ( .A(n1775), .B(n1769), .Z(n1770) );
  AND U4875 ( .A(n1771), .B(n1770), .Z(n1827) );
  XNOR U4876 ( .A(n1845), .B(n1827), .Z(n1802) );
  OR U4877 ( .A(n1802), .B(n1772), .Z(n1795) );
  NAND U4878 ( .A(n1783), .B(n1773), .Z(n1779) );
  AND U4879 ( .A(n1775), .B(n1774), .Z(n1782) );
  XNOR U4880 ( .A(n1782), .B(n1780), .Z(n1776) );
  NAND U4881 ( .A(n1777), .B(n1776), .Z(n1778) );
  AND U4882 ( .A(n1779), .B(n1778), .Z(n1799) );
  NAND U4883 ( .A(n1781), .B(n1780), .Z(n1787) );
  XNOR U4884 ( .A(n1783), .B(n1782), .Z(n1784) );
  NAND U4885 ( .A(n1785), .B(n1784), .Z(n1786) );
  NAND U4886 ( .A(n1787), .B(n1786), .Z(n1839) );
  XNOR U4887 ( .A(n1799), .B(n1839), .Z(n1817) );
  XOR U4888 ( .A(n1817), .B(n1802), .Z(n1804) );
  OR U4889 ( .A(n1804), .B(n1788), .Z(n1789) );
  XNOR U4890 ( .A(n1795), .B(n1789), .Z(n1821) );
  XOR U4891 ( .A(n1799), .B(n1845), .Z(n1807) );
  OR U4892 ( .A(n1790), .B(n1807), .Z(n1847) );
  NANDN U4893 ( .A(n1799), .B(n1791), .Z(n1792) );
  XNOR U4894 ( .A(n1847), .B(n1792), .Z(n1825) );
  XOR U4895 ( .A(n1821), .B(n1825), .Z(n1810) );
  NANDN U4896 ( .A(n1793), .B(n1817), .Z(n1794) );
  XNOR U4897 ( .A(n1795), .B(n1794), .Z(n1853) );
  XNOR U4898 ( .A(n1839), .B(n1827), .Z(n1829) );
  NANDN U4899 ( .A(n1829), .B(n1796), .Z(n1813) );
  NAND U4900 ( .A(n1797), .B(n1827), .Z(n1798) );
  XNOR U4901 ( .A(n1813), .B(n1798), .Z(n1844) );
  XOR U4902 ( .A(n1853), .B(n1844), .Z(n1836) );
  XNOR U4903 ( .A(n1810), .B(n1836), .Z(z[80]) );
  ANDN U4904 ( .B(n1800), .A(n1799), .Z(n1809) );
  NANDN U4905 ( .A(n1802), .B(n1801), .Z(n1820) );
  NANDN U4906 ( .A(n1804), .B(n1803), .Z(n1805) );
  XNOR U4907 ( .A(n1820), .B(n1805), .Z(n1848) );
  NANDN U4908 ( .A(n1807), .B(n1806), .Z(n1814) );
  XNOR U4909 ( .A(n1848), .B(n1814), .Z(n1808) );
  XOR U4910 ( .A(n1809), .B(n1808), .Z(n1834) );
  XOR U4911 ( .A(n1834), .B(n1810), .Z(n1852) );
  ANDN U4912 ( .B(n1845), .A(n1811), .Z(n1816) );
  NAND U4913 ( .A(n1838), .B(n1839), .Z(n1812) );
  XNOR U4914 ( .A(n1813), .B(n1812), .Z(n1824) );
  XNOR U4915 ( .A(n1814), .B(n1824), .Z(n1815) );
  XNOR U4916 ( .A(n1816), .B(n1815), .Z(n1823) );
  NAND U4917 ( .A(n1818), .B(n1817), .Z(n1819) );
  XNOR U4918 ( .A(n1820), .B(n1819), .Z(n1830) );
  XNOR U4919 ( .A(n1821), .B(n1830), .Z(n1822) );
  XOR U4920 ( .A(n1823), .B(n1822), .Z(n1833) );
  XNOR U4921 ( .A(n1852), .B(n1833), .Z(z[81]) );
  XNOR U4922 ( .A(n1825), .B(n1824), .Z(z[82]) );
  ANDN U4923 ( .B(n1827), .A(n1826), .Z(n1832) );
  NANDN U4924 ( .A(n1829), .B(n1828), .Z(n1842) );
  XNOR U4925 ( .A(n1830), .B(n1842), .Z(n1831) );
  XOR U4926 ( .A(n1832), .B(n1831), .Z(n1851) );
  XOR U4927 ( .A(n1834), .B(n1833), .Z(n1835) );
  XOR U4928 ( .A(n1851), .B(n1835), .Z(z[83]) );
  XOR U4929 ( .A(n1836), .B(z[82]), .Z(z[84]) );
  XNOR U4930 ( .A(n1838), .B(n1837), .Z(n1840) );
  NAND U4931 ( .A(n1840), .B(n1839), .Z(n1841) );
  XOR U4932 ( .A(n1842), .B(n1841), .Z(n1843) );
  XNOR U4933 ( .A(n1844), .B(n1843), .Z(n1850) );
  NAND U4934 ( .A(x[80]), .B(n1845), .Z(n1846) );
  XNOR U4935 ( .A(n1847), .B(n1846), .Z(n1854) );
  XNOR U4936 ( .A(n1848), .B(n1854), .Z(n1849) );
  XOR U4937 ( .A(n1850), .B(n1849), .Z(z[85]) );
  XNOR U4938 ( .A(n1852), .B(n1851), .Z(z[86]) );
  XNOR U4939 ( .A(n1854), .B(n1853), .Z(n1855) );
  XNOR U4940 ( .A(z[81]), .B(n1855), .Z(z[87]) );
  XOR U4941 ( .A(x[88]), .B(x[94]), .Z(n1856) );
  XOR U4942 ( .A(x[93]), .B(n1856), .Z(n1963) );
  IV U4943 ( .A(n1963), .Z(n1858) );
  IV U4944 ( .A(x[89]), .Z(n1962) );
  NAND U4945 ( .A(n1858), .B(n1962), .Z(n1865) );
  XOR U4946 ( .A(x[91]), .B(x[89]), .Z(n1861) );
  XNOR U4947 ( .A(x[90]), .B(n1856), .Z(n1857) );
  XNOR U4948 ( .A(n1861), .B(n1857), .Z(n1920) );
  XNOR U4949 ( .A(n1858), .B(n1920), .Z(n1919) );
  IV U4950 ( .A(x[95]), .Z(n1859) );
  XNOR U4951 ( .A(x[89]), .B(n1859), .Z(n1953) );
  NAND U4952 ( .A(n1919), .B(n1953), .Z(n1868) );
  XNOR U4953 ( .A(n1858), .B(n1859), .Z(n1951) );
  XOR U4954 ( .A(n1920), .B(n1951), .Z(n1876) );
  XOR U4955 ( .A(n1868), .B(n1876), .Z(n1863) );
  XNOR U4956 ( .A(x[88]), .B(n1920), .Z(n1895) );
  XOR U4957 ( .A(x[92]), .B(n1859), .Z(n1860) );
  IV U4958 ( .A(n1860), .Z(n1924) );
  NANDN U4959 ( .A(n1895), .B(n1924), .Z(n1867) );
  XOR U4960 ( .A(n1861), .B(n1860), .Z(n1913) );
  XOR U4961 ( .A(n1919), .B(n1913), .Z(n1911) );
  XOR U4962 ( .A(x[90]), .B(x[92]), .Z(n1926) );
  NANDN U4963 ( .A(n1911), .B(n1926), .Z(n1862) );
  XNOR U4964 ( .A(n1867), .B(n1862), .Z(n1872) );
  XOR U4965 ( .A(n1863), .B(n1872), .Z(n1864) );
  XOR U4966 ( .A(n1865), .B(n1864), .Z(n1906) );
  IV U4967 ( .A(n1906), .Z(n1900) );
  ANDN U4968 ( .B(n1951), .A(n1920), .Z(n1870) );
  XNOR U4969 ( .A(x[88]), .B(n1913), .Z(n1914) );
  XNOR U4970 ( .A(n1963), .B(n1914), .Z(n1916) );
  XOR U4971 ( .A(x[90]), .B(x[95]), .Z(n1941) );
  NANDN U4972 ( .A(n1916), .B(n1941), .Z(n1866) );
  XNOR U4973 ( .A(n1867), .B(n1866), .Z(n1883) );
  XNOR U4974 ( .A(n1868), .B(n1883), .Z(n1869) );
  XOR U4975 ( .A(n1870), .B(n1869), .Z(n1896) );
  NAND U4976 ( .A(n1900), .B(n1896), .Z(n1890) );
  IV U4977 ( .A(n1896), .Z(n1897) );
  XOR U4978 ( .A(n1906), .B(n1897), .Z(n1888) );
  XOR U4979 ( .A(x[90]), .B(x[89]), .Z(n1871) );
  XNOR U4980 ( .A(n1951), .B(n1871), .Z(n1923) );
  NAND U4981 ( .A(n1923), .B(n1914), .Z(n1878) );
  XNOR U4982 ( .A(x[92]), .B(n1963), .Z(n1934) );
  XOR U4983 ( .A(n1924), .B(n1871), .Z(n1929) );
  NANDN U4984 ( .A(n1913), .B(n1929), .Z(n1879) );
  XOR U4985 ( .A(n1934), .B(n1879), .Z(n1874) );
  XOR U4986 ( .A(x[88]), .B(n1872), .Z(n1873) );
  XNOR U4987 ( .A(n1874), .B(n1873), .Z(n1875) );
  XOR U4988 ( .A(n1876), .B(n1875), .Z(n1877) );
  XOR U4989 ( .A(n1878), .B(n1877), .Z(n1908) );
  IV U4990 ( .A(n1908), .Z(n1903) );
  AND U4991 ( .A(n1900), .B(n1903), .Z(n1886) );
  ANDN U4992 ( .B(x[88]), .A(n1934), .Z(n1885) );
  XNOR U4993 ( .A(n1923), .B(n1879), .Z(n1881) );
  XNOR U4994 ( .A(x[89]), .B(n1914), .Z(n1880) );
  XNOR U4995 ( .A(n1881), .B(n1880), .Z(n1882) );
  XOR U4996 ( .A(n1883), .B(n1882), .Z(n1884) );
  XOR U4997 ( .A(n1885), .B(n1884), .Z(n1898) );
  IV U4998 ( .A(n1898), .Z(n1904) );
  XNOR U4999 ( .A(n1886), .B(n1904), .Z(n1887) );
  NAND U5000 ( .A(n1888), .B(n1887), .Z(n1889) );
  NAND U5001 ( .A(n1890), .B(n1889), .Z(n1970) );
  NAND U5002 ( .A(n1904), .B(n1897), .Z(n1891) );
  NAND U5003 ( .A(n1903), .B(n1891), .Z(n1894) );
  XOR U5004 ( .A(n1897), .B(n1900), .Z(n1892) );
  NAND U5005 ( .A(n1898), .B(n1892), .Z(n1893) );
  AND U5006 ( .A(n1894), .B(n1893), .Z(n1952) );
  XNOR U5007 ( .A(n1970), .B(n1952), .Z(n1925) );
  OR U5008 ( .A(n1925), .B(n1895), .Z(n1918) );
  NAND U5009 ( .A(n1906), .B(n1896), .Z(n1902) );
  AND U5010 ( .A(n1898), .B(n1897), .Z(n1905) );
  XNOR U5011 ( .A(n1905), .B(n1903), .Z(n1899) );
  NAND U5012 ( .A(n1900), .B(n1899), .Z(n1901) );
  AND U5013 ( .A(n1902), .B(n1901), .Z(n1922) );
  NAND U5014 ( .A(n1904), .B(n1903), .Z(n1910) );
  XNOR U5015 ( .A(n1906), .B(n1905), .Z(n1907) );
  NAND U5016 ( .A(n1908), .B(n1907), .Z(n1909) );
  NAND U5017 ( .A(n1910), .B(n1909), .Z(n1964) );
  XNOR U5018 ( .A(n1922), .B(n1964), .Z(n1940) );
  XOR U5019 ( .A(n1940), .B(n1925), .Z(n1927) );
  OR U5020 ( .A(n1927), .B(n1911), .Z(n1912) );
  XNOR U5021 ( .A(n1918), .B(n1912), .Z(n1944) );
  XOR U5022 ( .A(n1922), .B(n1970), .Z(n1930) );
  OR U5023 ( .A(n1913), .B(n1930), .Z(n1972) );
  NANDN U5024 ( .A(n1922), .B(n1914), .Z(n1915) );
  XNOR U5025 ( .A(n1972), .B(n1915), .Z(n1950) );
  XOR U5026 ( .A(n1944), .B(n1950), .Z(n1933) );
  NANDN U5027 ( .A(n1916), .B(n1940), .Z(n1917) );
  XNOR U5028 ( .A(n1918), .B(n1917), .Z(n1978) );
  XNOR U5029 ( .A(n1964), .B(n1952), .Z(n1954) );
  NANDN U5030 ( .A(n1954), .B(n1919), .Z(n1936) );
  NAND U5031 ( .A(n1920), .B(n1952), .Z(n1921) );
  XNOR U5032 ( .A(n1936), .B(n1921), .Z(n1969) );
  XOR U5033 ( .A(n1978), .B(n1969), .Z(n1961) );
  XNOR U5034 ( .A(n1933), .B(n1961), .Z(z[88]) );
  ANDN U5035 ( .B(n1923), .A(n1922), .Z(n1932) );
  NANDN U5036 ( .A(n1925), .B(n1924), .Z(n1943) );
  NANDN U5037 ( .A(n1927), .B(n1926), .Z(n1928) );
  XNOR U5038 ( .A(n1943), .B(n1928), .Z(n1973) );
  NANDN U5039 ( .A(n1930), .B(n1929), .Z(n1937) );
  XNOR U5040 ( .A(n1973), .B(n1937), .Z(n1931) );
  XOR U5041 ( .A(n1932), .B(n1931), .Z(n1959) );
  XOR U5042 ( .A(n1959), .B(n1933), .Z(n1977) );
  ANDN U5043 ( .B(n1970), .A(n1934), .Z(n1939) );
  NAND U5044 ( .A(n1963), .B(n1964), .Z(n1935) );
  XNOR U5045 ( .A(n1936), .B(n1935), .Z(n1949) );
  XNOR U5046 ( .A(n1937), .B(n1949), .Z(n1938) );
  XNOR U5047 ( .A(n1939), .B(n1938), .Z(n1946) );
  NAND U5048 ( .A(n1941), .B(n1940), .Z(n1942) );
  XNOR U5049 ( .A(n1943), .B(n1942), .Z(n1955) );
  XNOR U5050 ( .A(n1944), .B(n1955), .Z(n1945) );
  XOR U5051 ( .A(n1946), .B(n1945), .Z(n1958) );
  XNOR U5052 ( .A(n1977), .B(n1958), .Z(z[89]) );
  XNOR U5053 ( .A(n1948), .B(n1947), .Z(z[8]) );
  XNOR U5054 ( .A(n1950), .B(n1949), .Z(z[90]) );
  ANDN U5055 ( .B(n1952), .A(n1951), .Z(n1957) );
  NANDN U5056 ( .A(n1954), .B(n1953), .Z(n1967) );
  XNOR U5057 ( .A(n1955), .B(n1967), .Z(n1956) );
  XOR U5058 ( .A(n1957), .B(n1956), .Z(n1976) );
  XOR U5059 ( .A(n1959), .B(n1958), .Z(n1960) );
  XOR U5060 ( .A(n1976), .B(n1960), .Z(z[91]) );
  XOR U5061 ( .A(n1961), .B(z[90]), .Z(z[92]) );
  XNOR U5062 ( .A(n1963), .B(n1962), .Z(n1965) );
  NAND U5063 ( .A(n1965), .B(n1964), .Z(n1966) );
  XOR U5064 ( .A(n1967), .B(n1966), .Z(n1968) );
  XNOR U5065 ( .A(n1969), .B(n1968), .Z(n1975) );
  NAND U5066 ( .A(x[88]), .B(n1970), .Z(n1971) );
  XNOR U5067 ( .A(n1972), .B(n1971), .Z(n1979) );
  XNOR U5068 ( .A(n1973), .B(n1979), .Z(n1974) );
  XOR U5069 ( .A(n1975), .B(n1974), .Z(z[93]) );
  XNOR U5070 ( .A(n1977), .B(n1976), .Z(z[94]) );
  XNOR U5071 ( .A(n1979), .B(n1978), .Z(n1980) );
  XNOR U5072 ( .A(z[89]), .B(n1980), .Z(z[95]) );
  XNOR U5073 ( .A(n1982), .B(n1981), .Z(z[96]) );
  XOR U5074 ( .A(n1984), .B(n1983), .Z(n1985) );
  XOR U5075 ( .A(n1986), .B(n1985), .Z(z[99]) );
endmodule


module SubBytes_4 ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986;

  XOR U2962 ( .A(x[16]), .B(x[22]), .Z(n685) );
  XNOR U2963 ( .A(n328), .B(n339), .Z(n341) );
  XOR U2964 ( .A(x[81]), .B(x[83]), .Z(n1738) );
  XNOR U2965 ( .A(n1324), .B(x[51]), .Z(n1222) );
  XNOR U2966 ( .A(n170), .B(n162), .Z(n143) );
  XOR U2967 ( .A(n493), .B(n494), .Z(n646) );
  XOR U2968 ( .A(x[85]), .B(n1733), .Z(n1838) );
  XOR U2969 ( .A(x[21]), .B(n685), .Z(n814) );
  XOR U2970 ( .A(x[53]), .B(n1218), .Z(n1323) );
  IV U2971 ( .A(x[1]), .Z(n1447) );
  XOR U2972 ( .A(x[0]), .B(x[6]), .Z(n2) );
  XOR U2973 ( .A(x[5]), .B(n2), .Z(n1446) );
  IV U2974 ( .A(n1446), .Z(n3) );
  AND U2975 ( .A(n1447), .B(n3), .Z(n10) );
  XNOR U2976 ( .A(x[3]), .B(n1447), .Z(n6) );
  XNOR U2977 ( .A(x[2]), .B(n6), .Z(n1) );
  XNOR U2978 ( .A(n2), .B(n1), .Z(n66) );
  IV U2979 ( .A(n66), .Z(n12) );
  XNOR U2980 ( .A(n12), .B(n1446), .Z(n65) );
  IV U2981 ( .A(x[7]), .Z(n4) );
  XNOR U2982 ( .A(x[1]), .B(n4), .Z(n1085) );
  NAND U2983 ( .A(n65), .B(n1085), .Z(n15) );
  XNOR U2984 ( .A(n4), .B(n3), .Z(n11) );
  IV U2985 ( .A(n11), .Z(n1083) );
  XOR U2986 ( .A(n66), .B(n1083), .Z(n31) );
  XNOR U2987 ( .A(n15), .B(n31), .Z(n8) );
  XOR U2988 ( .A(x[0]), .B(n12), .Z(n41) );
  XOR U2989 ( .A(x[4]), .B(n4), .Z(n5) );
  IV U2990 ( .A(n5), .Z(n790) );
  NANDN U2991 ( .A(n41), .B(n790), .Z(n14) );
  XNOR U2992 ( .A(n6), .B(n5), .Z(n59) );
  XNOR U2993 ( .A(n65), .B(n59), .Z(n57) );
  XOR U2994 ( .A(x[2]), .B(x[4]), .Z(n792) );
  NANDN U2995 ( .A(n57), .B(n792), .Z(n7) );
  XOR U2996 ( .A(n14), .B(n7), .Z(n33) );
  XNOR U2997 ( .A(n8), .B(n33), .Z(n9) );
  XOR U2998 ( .A(n10), .B(n9), .Z(n46) );
  IV U2999 ( .A(n46), .Z(n52) );
  AND U3000 ( .A(n12), .B(n11), .Z(n17) );
  XOR U3001 ( .A(x[0]), .B(n59), .Z(n60) );
  XNOR U3002 ( .A(n1446), .B(n60), .Z(n62) );
  XOR U3003 ( .A(x[2]), .B(x[7]), .Z(n807) );
  NANDN U3004 ( .A(n62), .B(n807), .Z(n13) );
  XNOR U3005 ( .A(n14), .B(n13), .Z(n22) );
  XNOR U3006 ( .A(n15), .B(n22), .Z(n16) );
  XOR U3007 ( .A(n17), .B(n16), .Z(n42) );
  XNOR U3008 ( .A(x[4]), .B(n1446), .Z(n800) );
  ANDN U3009 ( .B(x[0]), .A(n800), .Z(n24) );
  XOR U3010 ( .A(x[2]), .B(x[1]), .Z(n18) );
  XOR U3011 ( .A(n1083), .B(n18), .Z(n789) );
  XOR U3012 ( .A(n790), .B(n18), .Z(n795) );
  NAND U3013 ( .A(n59), .B(n795), .Z(n26) );
  XNOR U3014 ( .A(n789), .B(n26), .Z(n20) );
  XNOR U3015 ( .A(x[1]), .B(n60), .Z(n19) );
  XNOR U3016 ( .A(n20), .B(n19), .Z(n21) );
  XOR U3017 ( .A(n22), .B(n21), .Z(n23) );
  XOR U3018 ( .A(n24), .B(n23), .Z(n44) );
  NAND U3019 ( .A(n42), .B(n44), .Z(n25) );
  NAND U3020 ( .A(n52), .B(n25), .Z(n36) );
  IV U3021 ( .A(n42), .Z(n43) );
  IV U3022 ( .A(n44), .Z(n50) );
  XOR U3023 ( .A(n26), .B(n800), .Z(n29) );
  AND U3024 ( .A(n789), .B(n60), .Z(n27) );
  XNOR U3025 ( .A(x[0]), .B(n27), .Z(n28) );
  XNOR U3026 ( .A(n29), .B(n28), .Z(n30) );
  XNOR U3027 ( .A(n31), .B(n30), .Z(n32) );
  XNOR U3028 ( .A(n33), .B(n32), .Z(n54) );
  IV U3029 ( .A(n54), .Z(n49) );
  XOR U3030 ( .A(n50), .B(n49), .Z(n34) );
  NAND U3031 ( .A(n43), .B(n34), .Z(n35) );
  AND U3032 ( .A(n36), .B(n35), .Z(n1454) );
  NAND U3033 ( .A(n50), .B(n43), .Z(n37) );
  NAND U3034 ( .A(n49), .B(n37), .Z(n40) );
  XOR U3035 ( .A(n43), .B(n46), .Z(n38) );
  NAND U3036 ( .A(n44), .B(n38), .Z(n39) );
  AND U3037 ( .A(n40), .B(n39), .Z(n1084) );
  XNOR U3038 ( .A(n1454), .B(n1084), .Z(n791) );
  OR U3039 ( .A(n791), .B(n41), .Z(n64) );
  NAND U3040 ( .A(n52), .B(n42), .Z(n48) );
  AND U3041 ( .A(n44), .B(n43), .Z(n51) );
  XNOR U3042 ( .A(n49), .B(n51), .Z(n45) );
  NAND U3043 ( .A(n46), .B(n45), .Z(n47) );
  AND U3044 ( .A(n48), .B(n47), .Z(n788) );
  NAND U3045 ( .A(n50), .B(n49), .Z(n56) );
  XNOR U3046 ( .A(n52), .B(n51), .Z(n53) );
  NAND U3047 ( .A(n54), .B(n53), .Z(n55) );
  NAND U3048 ( .A(n56), .B(n55), .Z(n1448) );
  XNOR U3049 ( .A(n788), .B(n1448), .Z(n806) );
  XOR U3050 ( .A(n806), .B(n791), .Z(n793) );
  OR U3051 ( .A(n793), .B(n57), .Z(n58) );
  XNOR U3052 ( .A(n64), .B(n58), .Z(n810) );
  XOR U3053 ( .A(n788), .B(n1454), .Z(n796) );
  NANDN U3054 ( .A(n796), .B(n59), .Z(n1456) );
  NANDN U3055 ( .A(n788), .B(n60), .Z(n61) );
  XNOR U3056 ( .A(n1456), .B(n61), .Z(n953) );
  XOR U3057 ( .A(n810), .B(n953), .Z(n799) );
  NANDN U3058 ( .A(n62), .B(n806), .Z(n63) );
  XNOR U3059 ( .A(n64), .B(n63), .Z(n1730) );
  XNOR U3060 ( .A(n1448), .B(n1084), .Z(n1086) );
  NANDN U3061 ( .A(n1086), .B(n65), .Z(n802) );
  NAND U3062 ( .A(n66), .B(n1084), .Z(n67) );
  XNOR U3063 ( .A(n802), .B(n67), .Z(n1453) );
  XOR U3064 ( .A(n1730), .B(n1453), .Z(n1309) );
  XNOR U3065 ( .A(n799), .B(n1309), .Z(z[0]) );
  XOR U3066 ( .A(x[96]), .B(x[102]), .Z(n68) );
  XOR U3067 ( .A(x[101]), .B(n68), .Z(n135) );
  XOR U3068 ( .A(x[100]), .B(n135), .Z(n171) );
  AND U3069 ( .A(x[96]), .B(n171), .Z(n78) );
  XOR U3070 ( .A(x[97]), .B(x[99]), .Z(n71) );
  XNOR U3071 ( .A(n68), .B(x[98]), .Z(n69) );
  XOR U3072 ( .A(n71), .B(n69), .Z(n129) );
  XOR U3073 ( .A(x[96]), .B(n129), .Z(n128) );
  XNOR U3074 ( .A(x[103]), .B(x[100]), .Z(n70) );
  IV U3075 ( .A(n70), .Z(n142) );
  NANDN U3076 ( .A(n128), .B(n142), .Z(n80) );
  IV U3077 ( .A(n135), .Z(n91) );
  XNOR U3078 ( .A(n71), .B(n70), .Z(n123) );
  XOR U3079 ( .A(x[96]), .B(n123), .Z(n124) );
  XOR U3080 ( .A(n91), .B(n124), .Z(n126) );
  XOR U3081 ( .A(x[98]), .B(x[103]), .Z(n164) );
  NANDN U3082 ( .A(n126), .B(n164), .Z(n72) );
  XNOR U3083 ( .A(n80), .B(n72), .Z(n87) );
  XNOR U3084 ( .A(n135), .B(x[103]), .Z(n161) );
  XOR U3085 ( .A(x[97]), .B(x[98]), .Z(n73) );
  XNOR U3086 ( .A(n161), .B(n73), .Z(n151) );
  XOR U3087 ( .A(n142), .B(n73), .Z(n152) );
  NAND U3088 ( .A(n123), .B(n152), .Z(n81) );
  XNOR U3089 ( .A(n151), .B(n81), .Z(n75) );
  XNOR U3090 ( .A(x[97]), .B(n124), .Z(n74) );
  XNOR U3091 ( .A(n75), .B(n74), .Z(n76) );
  XOR U3092 ( .A(n87), .B(n76), .Z(n77) );
  XOR U3093 ( .A(n78), .B(n77), .Z(n115) );
  IV U3094 ( .A(n115), .Z(n108) );
  XNOR U3095 ( .A(n129), .B(n135), .Z(n105) );
  XNOR U3096 ( .A(n105), .B(n123), .Z(n158) );
  XNOR U3097 ( .A(x[98]), .B(x[100]), .Z(n144) );
  OR U3098 ( .A(n158), .B(n144), .Z(n79) );
  XOR U3099 ( .A(n80), .B(n79), .Z(n94) );
  XNOR U3100 ( .A(n129), .B(n161), .Z(n92) );
  XNOR U3101 ( .A(n81), .B(n171), .Z(n84) );
  AND U3102 ( .A(n151), .B(n124), .Z(n82) );
  XNOR U3103 ( .A(x[96]), .B(n82), .Z(n83) );
  XNOR U3104 ( .A(n84), .B(n83), .Z(n85) );
  XOR U3105 ( .A(n92), .B(n85), .Z(n86) );
  XOR U3106 ( .A(n94), .B(n86), .Z(n118) );
  AND U3107 ( .A(n129), .B(n161), .Z(n89) );
  IV U3108 ( .A(x[97]), .Z(n136) );
  XNOR U3109 ( .A(n136), .B(x[103]), .Z(n133) );
  NAND U3110 ( .A(n105), .B(n133), .Z(n93) );
  XNOR U3111 ( .A(n93), .B(n87), .Z(n88) );
  XOR U3112 ( .A(n89), .B(n88), .Z(n107) );
  NAND U3113 ( .A(n118), .B(n107), .Z(n90) );
  NAND U3114 ( .A(n108), .B(n90), .Z(n99) );
  IV U3115 ( .A(n118), .Z(n102) );
  NAND U3116 ( .A(n91), .B(n136), .Z(n97) );
  XOR U3117 ( .A(n93), .B(n92), .Z(n95) );
  XNOR U3118 ( .A(n95), .B(n94), .Z(n96) );
  XOR U3119 ( .A(n97), .B(n96), .Z(n114) );
  IV U3120 ( .A(n107), .Z(n116) );
  XOR U3121 ( .A(n114), .B(n116), .Z(n111) );
  NAND U3122 ( .A(n102), .B(n111), .Z(n98) );
  AND U3123 ( .A(n99), .B(n98), .Z(n127) );
  NAND U3124 ( .A(n118), .B(n108), .Z(n104) );
  AND U3125 ( .A(n115), .B(n116), .Z(n100) );
  XNOR U3126 ( .A(n114), .B(n100), .Z(n101) );
  NAND U3127 ( .A(n102), .B(n101), .Z(n103) );
  AND U3128 ( .A(n104), .B(n103), .Z(n138) );
  XNOR U3129 ( .A(n127), .B(n138), .Z(n134) );
  NANDN U3130 ( .A(n134), .B(n105), .Z(n131) );
  NANDN U3131 ( .A(n138), .B(n135), .Z(n106) );
  XNOR U3132 ( .A(n131), .B(n106), .Z(n173) );
  IV U3133 ( .A(n114), .Z(n120) );
  NAND U3134 ( .A(n120), .B(n107), .Z(n113) );
  AND U3135 ( .A(n120), .B(n118), .Z(n109) );
  XNOR U3136 ( .A(n109), .B(n108), .Z(n110) );
  NAND U3137 ( .A(n111), .B(n110), .Z(n112) );
  NAND U3138 ( .A(n113), .B(n112), .Z(n170) );
  NAND U3139 ( .A(n114), .B(n116), .Z(n122) );
  NAND U3140 ( .A(n116), .B(n115), .Z(n117) );
  XNOR U3141 ( .A(n118), .B(n117), .Z(n119) );
  NAND U3142 ( .A(n120), .B(n119), .Z(n121) );
  NAND U3143 ( .A(n122), .B(n121), .Z(n150) );
  XOR U3144 ( .A(n170), .B(n150), .Z(n153) );
  NANDN U3145 ( .A(n153), .B(n123), .Z(n147) );
  NANDN U3146 ( .A(n150), .B(n124), .Z(n125) );
  XNOR U3147 ( .A(n147), .B(n125), .Z(n160) );
  XNOR U3148 ( .A(n173), .B(n160), .Z(z[98]) );
  XOR U3149 ( .A(n150), .B(n138), .Z(n163) );
  ANDN U3150 ( .B(n163), .A(n126), .Z(n184) );
  IV U3151 ( .A(n127), .Z(n162) );
  OR U3152 ( .A(n143), .B(n128), .Z(n182) );
  NANDN U3153 ( .A(n129), .B(n162), .Z(n130) );
  XNOR U3154 ( .A(n131), .B(n130), .Z(n141) );
  XNOR U3155 ( .A(n182), .B(n141), .Z(n132) );
  XOR U3156 ( .A(n184), .B(n132), .Z(n1982) );
  XNOR U3157 ( .A(n1982), .B(z[98]), .Z(z[100]) );
  NANDN U3158 ( .A(n134), .B(n133), .Z(n167) );
  XNOR U3159 ( .A(n136), .B(n135), .Z(n137) );
  NANDN U3160 ( .A(n138), .B(n137), .Z(n139) );
  XOR U3161 ( .A(n167), .B(n139), .Z(n140) );
  XNOR U3162 ( .A(n141), .B(n140), .Z(n149) );
  NANDN U3163 ( .A(n143), .B(n142), .Z(n166) );
  XNOR U3164 ( .A(n143), .B(n163), .Z(n157) );
  NANDN U3165 ( .A(n144), .B(n157), .Z(n145) );
  XNOR U3166 ( .A(n166), .B(n145), .Z(n154) );
  NAND U3167 ( .A(n170), .B(x[96]), .Z(n146) );
  XNOR U3168 ( .A(n147), .B(n146), .Z(n181) );
  XNOR U3169 ( .A(n154), .B(n181), .Z(n148) );
  XOR U3170 ( .A(n149), .B(n148), .Z(z[101]) );
  ANDN U3171 ( .B(n151), .A(n150), .Z(n156) );
  NANDN U3172 ( .A(n153), .B(n152), .Z(n172) );
  XNOR U3173 ( .A(n172), .B(n154), .Z(n155) );
  XOR U3174 ( .A(n156), .B(n155), .Z(n1983) );
  NANDN U3175 ( .A(n158), .B(n157), .Z(n159) );
  XOR U3176 ( .A(n182), .B(n159), .Z(n176) );
  XOR U3177 ( .A(n176), .B(n160), .Z(n1981) );
  XNOR U3178 ( .A(n1983), .B(n1981), .Z(n180) );
  ANDN U3179 ( .B(n162), .A(n161), .Z(n169) );
  NAND U3180 ( .A(n164), .B(n163), .Z(n165) );
  XNOR U3181 ( .A(n166), .B(n165), .Z(n177) );
  XNOR U3182 ( .A(n177), .B(n167), .Z(n168) );
  XOR U3183 ( .A(n169), .B(n168), .Z(n1986) );
  XNOR U3184 ( .A(n180), .B(n1986), .Z(z[102]) );
  AND U3185 ( .A(n171), .B(n170), .Z(n175) );
  XNOR U3186 ( .A(n173), .B(n172), .Z(n174) );
  XNOR U3187 ( .A(n175), .B(n174), .Z(n179) );
  XOR U3188 ( .A(n177), .B(n176), .Z(n178) );
  XOR U3189 ( .A(n179), .B(n178), .Z(n1984) );
  XNOR U3190 ( .A(n1984), .B(n180), .Z(z[97]) );
  XNOR U3191 ( .A(n182), .B(n181), .Z(n183) );
  XNOR U3192 ( .A(n184), .B(n183), .Z(n185) );
  XOR U3193 ( .A(n185), .B(z[97]), .Z(z[103]) );
  IV U3194 ( .A(x[105]), .Z(n292) );
  XOR U3195 ( .A(x[104]), .B(x[110]), .Z(n187) );
  XOR U3196 ( .A(x[109]), .B(n187), .Z(n291) );
  IV U3197 ( .A(n291), .Z(n188) );
  AND U3198 ( .A(n292), .B(n188), .Z(n195) );
  XNOR U3199 ( .A(x[107]), .B(n292), .Z(n191) );
  XNOR U3200 ( .A(x[106]), .B(n191), .Z(n186) );
  XNOR U3201 ( .A(n187), .B(n186), .Z(n251) );
  IV U3202 ( .A(n251), .Z(n197) );
  XNOR U3203 ( .A(n197), .B(n291), .Z(n250) );
  IV U3204 ( .A(x[111]), .Z(n189) );
  XNOR U3205 ( .A(x[105]), .B(n189), .Z(n282) );
  NAND U3206 ( .A(n250), .B(n282), .Z(n200) );
  XNOR U3207 ( .A(n189), .B(n188), .Z(n196) );
  IV U3208 ( .A(n196), .Z(n280) );
  XOR U3209 ( .A(n251), .B(n280), .Z(n216) );
  XNOR U3210 ( .A(n200), .B(n216), .Z(n193) );
  XOR U3211 ( .A(x[104]), .B(n197), .Z(n226) );
  XOR U3212 ( .A(x[108]), .B(n189), .Z(n190) );
  IV U3213 ( .A(n190), .Z(n255) );
  NANDN U3214 ( .A(n226), .B(n255), .Z(n199) );
  XNOR U3215 ( .A(n191), .B(n190), .Z(n244) );
  XNOR U3216 ( .A(n250), .B(n244), .Z(n242) );
  XOR U3217 ( .A(x[106]), .B(x[108]), .Z(n257) );
  NANDN U3218 ( .A(n242), .B(n257), .Z(n192) );
  XOR U3219 ( .A(n199), .B(n192), .Z(n218) );
  XNOR U3220 ( .A(n193), .B(n218), .Z(n194) );
  XOR U3221 ( .A(n195), .B(n194), .Z(n231) );
  IV U3222 ( .A(n231), .Z(n237) );
  AND U3223 ( .A(n197), .B(n196), .Z(n202) );
  XOR U3224 ( .A(x[104]), .B(n244), .Z(n245) );
  XNOR U3225 ( .A(n291), .B(n245), .Z(n247) );
  XOR U3226 ( .A(x[106]), .B(x[111]), .Z(n272) );
  NANDN U3227 ( .A(n247), .B(n272), .Z(n198) );
  XNOR U3228 ( .A(n199), .B(n198), .Z(n207) );
  XNOR U3229 ( .A(n200), .B(n207), .Z(n201) );
  XOR U3230 ( .A(n202), .B(n201), .Z(n227) );
  XNOR U3231 ( .A(x[108]), .B(n291), .Z(n265) );
  ANDN U3232 ( .B(x[104]), .A(n265), .Z(n209) );
  XOR U3233 ( .A(x[106]), .B(x[105]), .Z(n203) );
  XOR U3234 ( .A(n280), .B(n203), .Z(n254) );
  XOR U3235 ( .A(n255), .B(n203), .Z(n260) );
  NAND U3236 ( .A(n244), .B(n260), .Z(n211) );
  XNOR U3237 ( .A(n254), .B(n211), .Z(n205) );
  XNOR U3238 ( .A(x[105]), .B(n245), .Z(n204) );
  XNOR U3239 ( .A(n205), .B(n204), .Z(n206) );
  XOR U3240 ( .A(n207), .B(n206), .Z(n208) );
  XOR U3241 ( .A(n209), .B(n208), .Z(n229) );
  NAND U3242 ( .A(n227), .B(n229), .Z(n210) );
  NAND U3243 ( .A(n237), .B(n210), .Z(n221) );
  IV U3244 ( .A(n227), .Z(n228) );
  IV U3245 ( .A(n229), .Z(n235) );
  XOR U3246 ( .A(n211), .B(n265), .Z(n214) );
  AND U3247 ( .A(n254), .B(n245), .Z(n212) );
  XNOR U3248 ( .A(x[104]), .B(n212), .Z(n213) );
  XNOR U3249 ( .A(n214), .B(n213), .Z(n215) );
  XNOR U3250 ( .A(n216), .B(n215), .Z(n217) );
  XNOR U3251 ( .A(n218), .B(n217), .Z(n239) );
  IV U3252 ( .A(n239), .Z(n234) );
  XOR U3253 ( .A(n235), .B(n234), .Z(n219) );
  NAND U3254 ( .A(n228), .B(n219), .Z(n220) );
  AND U3255 ( .A(n221), .B(n220), .Z(n299) );
  NAND U3256 ( .A(n235), .B(n228), .Z(n222) );
  NAND U3257 ( .A(n234), .B(n222), .Z(n225) );
  XOR U3258 ( .A(n228), .B(n231), .Z(n223) );
  NAND U3259 ( .A(n229), .B(n223), .Z(n224) );
  AND U3260 ( .A(n225), .B(n224), .Z(n281) );
  XNOR U3261 ( .A(n299), .B(n281), .Z(n256) );
  OR U3262 ( .A(n256), .B(n226), .Z(n249) );
  NAND U3263 ( .A(n237), .B(n227), .Z(n233) );
  AND U3264 ( .A(n229), .B(n228), .Z(n236) );
  XNOR U3265 ( .A(n234), .B(n236), .Z(n230) );
  NAND U3266 ( .A(n231), .B(n230), .Z(n232) );
  AND U3267 ( .A(n233), .B(n232), .Z(n253) );
  NAND U3268 ( .A(n235), .B(n234), .Z(n241) );
  XNOR U3269 ( .A(n237), .B(n236), .Z(n238) );
  NAND U3270 ( .A(n239), .B(n238), .Z(n240) );
  NAND U3271 ( .A(n241), .B(n240), .Z(n293) );
  XNOR U3272 ( .A(n253), .B(n293), .Z(n271) );
  XOR U3273 ( .A(n271), .B(n256), .Z(n258) );
  OR U3274 ( .A(n258), .B(n242), .Z(n243) );
  XNOR U3275 ( .A(n249), .B(n243), .Z(n275) );
  XOR U3276 ( .A(n253), .B(n299), .Z(n261) );
  NANDN U3277 ( .A(n261), .B(n244), .Z(n301) );
  NANDN U3278 ( .A(n253), .B(n245), .Z(n246) );
  XNOR U3279 ( .A(n301), .B(n246), .Z(n279) );
  XOR U3280 ( .A(n275), .B(n279), .Z(n264) );
  NANDN U3281 ( .A(n247), .B(n271), .Z(n248) );
  XNOR U3282 ( .A(n249), .B(n248), .Z(n366) );
  XNOR U3283 ( .A(n293), .B(n281), .Z(n283) );
  NANDN U3284 ( .A(n283), .B(n250), .Z(n267) );
  NAND U3285 ( .A(n251), .B(n281), .Z(n252) );
  XNOR U3286 ( .A(n267), .B(n252), .Z(n298) );
  XOR U3287 ( .A(n366), .B(n298), .Z(n290) );
  XNOR U3288 ( .A(n264), .B(n290), .Z(z[104]) );
  ANDN U3289 ( .B(n254), .A(n253), .Z(n263) );
  NANDN U3290 ( .A(n256), .B(n255), .Z(n274) );
  NANDN U3291 ( .A(n258), .B(n257), .Z(n259) );
  XNOR U3292 ( .A(n274), .B(n259), .Z(n302) );
  NANDN U3293 ( .A(n261), .B(n260), .Z(n268) );
  XNOR U3294 ( .A(n302), .B(n268), .Z(n262) );
  XOR U3295 ( .A(n263), .B(n262), .Z(n288) );
  XOR U3296 ( .A(n288), .B(n264), .Z(n365) );
  ANDN U3297 ( .B(n299), .A(n265), .Z(n270) );
  NAND U3298 ( .A(n291), .B(n293), .Z(n266) );
  XNOR U3299 ( .A(n267), .B(n266), .Z(n278) );
  XNOR U3300 ( .A(n268), .B(n278), .Z(n269) );
  XNOR U3301 ( .A(n270), .B(n269), .Z(n277) );
  NAND U3302 ( .A(n272), .B(n271), .Z(n273) );
  XNOR U3303 ( .A(n274), .B(n273), .Z(n284) );
  XNOR U3304 ( .A(n275), .B(n284), .Z(n276) );
  XOR U3305 ( .A(n277), .B(n276), .Z(n287) );
  XNOR U3306 ( .A(n365), .B(n287), .Z(z[105]) );
  XNOR U3307 ( .A(n279), .B(n278), .Z(z[106]) );
  AND U3308 ( .A(n281), .B(n280), .Z(n286) );
  NANDN U3309 ( .A(n283), .B(n282), .Z(n296) );
  XNOR U3310 ( .A(n284), .B(n296), .Z(n285) );
  XOR U3311 ( .A(n286), .B(n285), .Z(n364) );
  XOR U3312 ( .A(n288), .B(n287), .Z(n289) );
  XOR U3313 ( .A(n364), .B(n289), .Z(z[107]) );
  XOR U3314 ( .A(n290), .B(z[106]), .Z(z[108]) );
  XNOR U3315 ( .A(n292), .B(n291), .Z(n294) );
  NAND U3316 ( .A(n294), .B(n293), .Z(n295) );
  XOR U3317 ( .A(n296), .B(n295), .Z(n297) );
  XNOR U3318 ( .A(n298), .B(n297), .Z(n304) );
  NAND U3319 ( .A(n299), .B(x[104]), .Z(n300) );
  XNOR U3320 ( .A(n301), .B(n300), .Z(n367) );
  XNOR U3321 ( .A(n302), .B(n367), .Z(n303) );
  XOR U3322 ( .A(n304), .B(n303), .Z(z[109]) );
  IV U3323 ( .A(x[15]), .Z(n311) );
  IV U3324 ( .A(x[10]), .Z(n315) );
  XOR U3325 ( .A(x[11]), .B(x[9]), .Z(n307) );
  XOR U3326 ( .A(n315), .B(n307), .Z(n352) );
  IV U3327 ( .A(n352), .Z(n309) );
  XOR U3328 ( .A(x[13]), .B(n309), .Z(n305) );
  IV U3329 ( .A(x[9]), .Z(n655) );
  XNOR U3330 ( .A(n311), .B(n655), .Z(n515) );
  NAND U3331 ( .A(n305), .B(n515), .Z(n306) );
  XNOR U3332 ( .A(n311), .B(n306), .Z(n339) );
  XOR U3333 ( .A(x[12]), .B(n311), .Z(n314) );
  XNOR U3334 ( .A(x[14]), .B(n309), .Z(n497) );
  NOR U3335 ( .A(n314), .B(n497), .Z(n318) );
  IV U3336 ( .A(x[13]), .Z(n353) );
  XOR U3337 ( .A(x[8]), .B(x[14]), .Z(n310) );
  XOR U3338 ( .A(n353), .B(n310), .Z(n325) );
  IV U3339 ( .A(n325), .Z(n656) );
  XOR U3340 ( .A(n314), .B(n307), .Z(n316) );
  XNOR U3341 ( .A(x[8]), .B(n316), .Z(n350) );
  XNOR U3342 ( .A(n656), .B(n350), .Z(n648) );
  XNOR U3343 ( .A(x[15]), .B(n315), .Z(n673) );
  NANDN U3344 ( .A(n648), .B(n673), .Z(n308) );
  XOR U3345 ( .A(n318), .B(n308), .Z(n333) );
  XOR U3346 ( .A(n310), .B(n309), .Z(n313) );
  XNOR U3347 ( .A(n325), .B(n311), .Z(n516) );
  ANDN U3348 ( .B(n313), .A(n516), .Z(n312) );
  XOR U3349 ( .A(n333), .B(n312), .Z(n328) );
  IV U3350 ( .A(n313), .Z(n647) );
  IV U3351 ( .A(n314), .Z(n507) );
  XNOR U3352 ( .A(n655), .B(n315), .Z(n321) );
  XOR U3353 ( .A(n507), .B(n321), .Z(n501) );
  IV U3354 ( .A(n316), .Z(n344) );
  NANDN U3355 ( .A(n501), .B(n344), .Z(n329) );
  XNOR U3356 ( .A(x[12]), .B(x[10]), .Z(n508) );
  XNOR U3357 ( .A(n648), .B(n497), .Z(n498) );
  OR U3358 ( .A(n508), .B(n498), .Z(n317) );
  XOR U3359 ( .A(n318), .B(n317), .Z(n327) );
  XOR U3360 ( .A(n329), .B(n327), .Z(n320) );
  XNOR U3361 ( .A(x[8]), .B(n507), .Z(n319) );
  XNOR U3362 ( .A(n320), .B(n319), .Z(n323) );
  XOR U3363 ( .A(n321), .B(n516), .Z(n505) );
  NAND U3364 ( .A(n350), .B(n505), .Z(n322) );
  XNOR U3365 ( .A(n323), .B(n322), .Z(n324) );
  XOR U3366 ( .A(n647), .B(n324), .Z(n356) );
  IV U3367 ( .A(n356), .Z(n359) );
  NAND U3368 ( .A(n325), .B(n655), .Z(n326) );
  XOR U3369 ( .A(n327), .B(n326), .Z(n338) );
  XNOR U3370 ( .A(n328), .B(n338), .Z(n348) );
  NAND U3371 ( .A(n359), .B(n348), .Z(n337) );
  XOR U3372 ( .A(n656), .B(x[12]), .Z(n502) );
  AND U3373 ( .A(n502), .B(x[8]), .Z(n335) );
  XNOR U3374 ( .A(n505), .B(n329), .Z(n331) );
  XNOR U3375 ( .A(x[9]), .B(n350), .Z(n330) );
  XNOR U3376 ( .A(n331), .B(n330), .Z(n332) );
  XOR U3377 ( .A(n333), .B(n332), .Z(n334) );
  XNOR U3378 ( .A(n335), .B(n334), .Z(n358) );
  NANDN U3379 ( .A(n348), .B(n358), .Z(n336) );
  AND U3380 ( .A(n337), .B(n336), .Z(n342) );
  XNOR U3381 ( .A(n339), .B(n338), .Z(n345) );
  NANDN U3382 ( .A(n345), .B(n356), .Z(n340) );
  XNOR U3383 ( .A(n342), .B(n340), .Z(n354) );
  OR U3384 ( .A(n341), .B(n354), .Z(n495) );
  NANDN U3385 ( .A(n358), .B(n341), .Z(n347) );
  XOR U3386 ( .A(n345), .B(n342), .Z(n343) );
  XNOR U3387 ( .A(n347), .B(n343), .Z(n355) );
  NOR U3388 ( .A(n355), .B(n345), .Z(n349) );
  XOR U3389 ( .A(n495), .B(n349), .Z(n500) );
  NANDN U3390 ( .A(n500), .B(n344), .Z(n664) );
  ANDN U3391 ( .B(n359), .A(n345), .Z(n346) );
  XNOR U3392 ( .A(n347), .B(n346), .Z(n361) );
  OR U3393 ( .A(n361), .B(n348), .Z(n496) );
  XNOR U3394 ( .A(n496), .B(n349), .Z(n504) );
  AND U3395 ( .A(n504), .B(n350), .Z(n351) );
  XOR U3396 ( .A(n664), .B(n351), .Z(n670) );
  XOR U3397 ( .A(n353), .B(n352), .Z(n357) );
  ANDN U3398 ( .B(n358), .A(n354), .Z(n493) );
  NOR U3399 ( .A(n356), .B(n355), .Z(n362) );
  XOR U3400 ( .A(n493), .B(n362), .Z(n514) );
  NAND U3401 ( .A(n357), .B(n514), .Z(n651) );
  XOR U3402 ( .A(n359), .B(n358), .Z(n360) );
  NANDN U3403 ( .A(n361), .B(n360), .Z(n494) );
  XOR U3404 ( .A(n494), .B(n362), .Z(n658) );
  NANDN U3405 ( .A(n658), .B(n656), .Z(n363) );
  XNOR U3406 ( .A(n651), .B(n363), .Z(n519) );
  XOR U3407 ( .A(n670), .B(n519), .Z(n654) );
  IV U3408 ( .A(n654), .Z(z[10]) );
  XNOR U3409 ( .A(n365), .B(n364), .Z(z[110]) );
  XNOR U3410 ( .A(n367), .B(n366), .Z(n368) );
  XNOR U3411 ( .A(z[105]), .B(n368), .Z(z[111]) );
  IV U3412 ( .A(x[113]), .Z(n475) );
  XOR U3413 ( .A(x[112]), .B(x[118]), .Z(n370) );
  XOR U3414 ( .A(x[117]), .B(n370), .Z(n474) );
  IV U3415 ( .A(n474), .Z(n371) );
  AND U3416 ( .A(n475), .B(n371), .Z(n378) );
  XNOR U3417 ( .A(x[115]), .B(n475), .Z(n374) );
  XNOR U3418 ( .A(x[114]), .B(n374), .Z(n369) );
  XNOR U3419 ( .A(n370), .B(n369), .Z(n434) );
  IV U3420 ( .A(n434), .Z(n380) );
  XNOR U3421 ( .A(n380), .B(n474), .Z(n433) );
  IV U3422 ( .A(x[119]), .Z(n372) );
  XNOR U3423 ( .A(x[113]), .B(n372), .Z(n465) );
  NAND U3424 ( .A(n433), .B(n465), .Z(n383) );
  XNOR U3425 ( .A(n372), .B(n371), .Z(n379) );
  IV U3426 ( .A(n379), .Z(n463) );
  XOR U3427 ( .A(n434), .B(n463), .Z(n399) );
  XNOR U3428 ( .A(n383), .B(n399), .Z(n376) );
  XOR U3429 ( .A(x[112]), .B(n380), .Z(n409) );
  XOR U3430 ( .A(x[116]), .B(n372), .Z(n373) );
  IV U3431 ( .A(n373), .Z(n438) );
  NANDN U3432 ( .A(n409), .B(n438), .Z(n382) );
  XNOR U3433 ( .A(n374), .B(n373), .Z(n427) );
  XNOR U3434 ( .A(n433), .B(n427), .Z(n425) );
  XOR U3435 ( .A(x[114]), .B(x[116]), .Z(n440) );
  NANDN U3436 ( .A(n425), .B(n440), .Z(n375) );
  XOR U3437 ( .A(n382), .B(n375), .Z(n401) );
  XNOR U3438 ( .A(n376), .B(n401), .Z(n377) );
  XOR U3439 ( .A(n378), .B(n377), .Z(n414) );
  IV U3440 ( .A(n414), .Z(n420) );
  AND U3441 ( .A(n380), .B(n379), .Z(n385) );
  XOR U3442 ( .A(x[112]), .B(n427), .Z(n428) );
  XNOR U3443 ( .A(n474), .B(n428), .Z(n430) );
  XOR U3444 ( .A(x[114]), .B(x[119]), .Z(n455) );
  NANDN U3445 ( .A(n430), .B(n455), .Z(n381) );
  XNOR U3446 ( .A(n382), .B(n381), .Z(n390) );
  XNOR U3447 ( .A(n383), .B(n390), .Z(n384) );
  XOR U3448 ( .A(n385), .B(n384), .Z(n410) );
  XNOR U3449 ( .A(x[116]), .B(n474), .Z(n448) );
  ANDN U3450 ( .B(x[112]), .A(n448), .Z(n392) );
  XOR U3451 ( .A(x[114]), .B(x[113]), .Z(n386) );
  XOR U3452 ( .A(n463), .B(n386), .Z(n437) );
  XOR U3453 ( .A(n438), .B(n386), .Z(n443) );
  NAND U3454 ( .A(n427), .B(n443), .Z(n394) );
  XNOR U3455 ( .A(n437), .B(n394), .Z(n388) );
  XNOR U3456 ( .A(x[113]), .B(n428), .Z(n387) );
  XNOR U3457 ( .A(n388), .B(n387), .Z(n389) );
  XOR U3458 ( .A(n390), .B(n389), .Z(n391) );
  XOR U3459 ( .A(n392), .B(n391), .Z(n412) );
  NAND U3460 ( .A(n410), .B(n412), .Z(n393) );
  NAND U3461 ( .A(n420), .B(n393), .Z(n404) );
  IV U3462 ( .A(n410), .Z(n411) );
  IV U3463 ( .A(n412), .Z(n418) );
  XOR U3464 ( .A(n394), .B(n448), .Z(n397) );
  AND U3465 ( .A(n437), .B(n428), .Z(n395) );
  XNOR U3466 ( .A(x[112]), .B(n395), .Z(n396) );
  XNOR U3467 ( .A(n397), .B(n396), .Z(n398) );
  XNOR U3468 ( .A(n399), .B(n398), .Z(n400) );
  XNOR U3469 ( .A(n401), .B(n400), .Z(n422) );
  IV U3470 ( .A(n422), .Z(n417) );
  XOR U3471 ( .A(n418), .B(n417), .Z(n402) );
  NAND U3472 ( .A(n411), .B(n402), .Z(n403) );
  AND U3473 ( .A(n404), .B(n403), .Z(n482) );
  NAND U3474 ( .A(n418), .B(n411), .Z(n405) );
  NAND U3475 ( .A(n417), .B(n405), .Z(n408) );
  XOR U3476 ( .A(n411), .B(n414), .Z(n406) );
  NAND U3477 ( .A(n412), .B(n406), .Z(n407) );
  AND U3478 ( .A(n408), .B(n407), .Z(n464) );
  XNOR U3479 ( .A(n482), .B(n464), .Z(n439) );
  OR U3480 ( .A(n439), .B(n409), .Z(n432) );
  NAND U3481 ( .A(n420), .B(n410), .Z(n416) );
  AND U3482 ( .A(n412), .B(n411), .Z(n419) );
  XNOR U3483 ( .A(n417), .B(n419), .Z(n413) );
  NAND U3484 ( .A(n414), .B(n413), .Z(n415) );
  AND U3485 ( .A(n416), .B(n415), .Z(n436) );
  NAND U3486 ( .A(n418), .B(n417), .Z(n424) );
  XNOR U3487 ( .A(n420), .B(n419), .Z(n421) );
  NAND U3488 ( .A(n422), .B(n421), .Z(n423) );
  NAND U3489 ( .A(n424), .B(n423), .Z(n476) );
  XNOR U3490 ( .A(n436), .B(n476), .Z(n454) );
  XOR U3491 ( .A(n454), .B(n439), .Z(n441) );
  OR U3492 ( .A(n441), .B(n425), .Z(n426) );
  XNOR U3493 ( .A(n432), .B(n426), .Z(n458) );
  XOR U3494 ( .A(n436), .B(n482), .Z(n444) );
  NANDN U3495 ( .A(n444), .B(n427), .Z(n484) );
  NANDN U3496 ( .A(n436), .B(n428), .Z(n429) );
  XNOR U3497 ( .A(n484), .B(n429), .Z(n462) );
  XOR U3498 ( .A(n458), .B(n462), .Z(n447) );
  NANDN U3499 ( .A(n430), .B(n454), .Z(n431) );
  XNOR U3500 ( .A(n432), .B(n431), .Z(n490) );
  XNOR U3501 ( .A(n476), .B(n464), .Z(n466) );
  NANDN U3502 ( .A(n466), .B(n433), .Z(n450) );
  NAND U3503 ( .A(n434), .B(n464), .Z(n435) );
  XNOR U3504 ( .A(n450), .B(n435), .Z(n481) );
  XOR U3505 ( .A(n490), .B(n481), .Z(n473) );
  XNOR U3506 ( .A(n447), .B(n473), .Z(z[112]) );
  ANDN U3507 ( .B(n437), .A(n436), .Z(n446) );
  NANDN U3508 ( .A(n439), .B(n438), .Z(n457) );
  NANDN U3509 ( .A(n441), .B(n440), .Z(n442) );
  XNOR U3510 ( .A(n457), .B(n442), .Z(n485) );
  NANDN U3511 ( .A(n444), .B(n443), .Z(n451) );
  XNOR U3512 ( .A(n485), .B(n451), .Z(n445) );
  XOR U3513 ( .A(n446), .B(n445), .Z(n471) );
  XOR U3514 ( .A(n471), .B(n447), .Z(n489) );
  ANDN U3515 ( .B(n482), .A(n448), .Z(n453) );
  NAND U3516 ( .A(n474), .B(n476), .Z(n449) );
  XNOR U3517 ( .A(n450), .B(n449), .Z(n461) );
  XNOR U3518 ( .A(n451), .B(n461), .Z(n452) );
  XNOR U3519 ( .A(n453), .B(n452), .Z(n460) );
  NAND U3520 ( .A(n455), .B(n454), .Z(n456) );
  XNOR U3521 ( .A(n457), .B(n456), .Z(n467) );
  XNOR U3522 ( .A(n458), .B(n467), .Z(n459) );
  XOR U3523 ( .A(n460), .B(n459), .Z(n470) );
  XNOR U3524 ( .A(n489), .B(n470), .Z(z[113]) );
  XNOR U3525 ( .A(n462), .B(n461), .Z(z[114]) );
  AND U3526 ( .A(n464), .B(n463), .Z(n469) );
  NANDN U3527 ( .A(n466), .B(n465), .Z(n479) );
  XNOR U3528 ( .A(n467), .B(n479), .Z(n468) );
  XOR U3529 ( .A(n469), .B(n468), .Z(n488) );
  XOR U3530 ( .A(n471), .B(n470), .Z(n472) );
  XOR U3531 ( .A(n488), .B(n472), .Z(z[115]) );
  XOR U3532 ( .A(n473), .B(z[114]), .Z(z[116]) );
  XNOR U3533 ( .A(n475), .B(n474), .Z(n477) );
  NAND U3534 ( .A(n477), .B(n476), .Z(n478) );
  XOR U3535 ( .A(n479), .B(n478), .Z(n480) );
  XNOR U3536 ( .A(n481), .B(n480), .Z(n487) );
  NAND U3537 ( .A(n482), .B(x[112]), .Z(n483) );
  XNOR U3538 ( .A(n484), .B(n483), .Z(n491) );
  XNOR U3539 ( .A(n485), .B(n491), .Z(n486) );
  XOR U3540 ( .A(n487), .B(n486), .Z(z[117]) );
  XNOR U3541 ( .A(n489), .B(n488), .Z(z[118]) );
  XNOR U3542 ( .A(n491), .B(n490), .Z(n492) );
  XNOR U3543 ( .A(z[113]), .B(n492), .Z(z[119]) );
  XNOR U3544 ( .A(n496), .B(n495), .Z(n662) );
  XOR U3545 ( .A(n646), .B(n662), .Z(n506) );
  NANDN U3546 ( .A(n497), .B(n506), .Z(n650) );
  XNOR U3547 ( .A(n658), .B(n504), .Z(n672) );
  XNOR U3548 ( .A(n506), .B(n672), .Z(n509) );
  OR U3549 ( .A(n498), .B(n509), .Z(n499) );
  XNOR U3550 ( .A(n650), .B(n499), .Z(n671) );
  OR U3551 ( .A(n501), .B(n500), .Z(n511) );
  ANDN U3552 ( .B(n502), .A(n662), .Z(n503) );
  XNOR U3553 ( .A(n511), .B(n503), .Z(n678) );
  AND U3554 ( .A(n505), .B(n504), .Z(n513) );
  NAND U3555 ( .A(n507), .B(n506), .Z(n675) );
  OR U3556 ( .A(n509), .B(n508), .Z(n510) );
  XNOR U3557 ( .A(n675), .B(n510), .Z(n667) );
  XNOR U3558 ( .A(n667), .B(n511), .Z(n512) );
  XOR U3559 ( .A(n513), .B(n512), .Z(n682) );
  NANDN U3560 ( .A(n515), .B(n514), .Z(n660) );
  OR U3561 ( .A(n516), .B(n646), .Z(n517) );
  XOR U3562 ( .A(n660), .B(n517), .Z(n518) );
  XNOR U3563 ( .A(n682), .B(n518), .Z(n677) );
  XNOR U3564 ( .A(n519), .B(n677), .Z(n520) );
  XOR U3565 ( .A(n678), .B(n520), .Z(n521) );
  XOR U3566 ( .A(n671), .B(n521), .Z(z[11]) );
  IV U3567 ( .A(x[121]), .Z(n628) );
  XOR U3568 ( .A(x[120]), .B(x[126]), .Z(n523) );
  XOR U3569 ( .A(x[125]), .B(n523), .Z(n627) );
  IV U3570 ( .A(n627), .Z(n524) );
  AND U3571 ( .A(n628), .B(n524), .Z(n531) );
  XNOR U3572 ( .A(x[123]), .B(n628), .Z(n527) );
  XNOR U3573 ( .A(x[122]), .B(n527), .Z(n522) );
  XNOR U3574 ( .A(n523), .B(n522), .Z(n587) );
  IV U3575 ( .A(n587), .Z(n533) );
  XNOR U3576 ( .A(n533), .B(n627), .Z(n586) );
  IV U3577 ( .A(x[127]), .Z(n525) );
  XNOR U3578 ( .A(x[121]), .B(n525), .Z(n618) );
  NAND U3579 ( .A(n586), .B(n618), .Z(n536) );
  XNOR U3580 ( .A(n525), .B(n524), .Z(n532) );
  IV U3581 ( .A(n532), .Z(n616) );
  XOR U3582 ( .A(n587), .B(n616), .Z(n552) );
  XNOR U3583 ( .A(n536), .B(n552), .Z(n529) );
  XOR U3584 ( .A(x[120]), .B(n533), .Z(n562) );
  XOR U3585 ( .A(x[124]), .B(n525), .Z(n526) );
  IV U3586 ( .A(n526), .Z(n591) );
  NANDN U3587 ( .A(n562), .B(n591), .Z(n535) );
  XNOR U3588 ( .A(n527), .B(n526), .Z(n580) );
  XNOR U3589 ( .A(n586), .B(n580), .Z(n578) );
  XOR U3590 ( .A(x[122]), .B(x[124]), .Z(n593) );
  NANDN U3591 ( .A(n578), .B(n593), .Z(n528) );
  XOR U3592 ( .A(n535), .B(n528), .Z(n554) );
  XNOR U3593 ( .A(n529), .B(n554), .Z(n530) );
  XOR U3594 ( .A(n531), .B(n530), .Z(n567) );
  IV U3595 ( .A(n567), .Z(n573) );
  AND U3596 ( .A(n533), .B(n532), .Z(n538) );
  XOR U3597 ( .A(x[120]), .B(n580), .Z(n581) );
  XNOR U3598 ( .A(n627), .B(n581), .Z(n583) );
  XOR U3599 ( .A(x[122]), .B(x[127]), .Z(n608) );
  NANDN U3600 ( .A(n583), .B(n608), .Z(n534) );
  XNOR U3601 ( .A(n535), .B(n534), .Z(n543) );
  XNOR U3602 ( .A(n536), .B(n543), .Z(n537) );
  XOR U3603 ( .A(n538), .B(n537), .Z(n563) );
  XNOR U3604 ( .A(x[124]), .B(n627), .Z(n601) );
  ANDN U3605 ( .B(x[120]), .A(n601), .Z(n545) );
  XOR U3606 ( .A(x[122]), .B(x[121]), .Z(n539) );
  XOR U3607 ( .A(n616), .B(n539), .Z(n590) );
  XOR U3608 ( .A(n591), .B(n539), .Z(n596) );
  NAND U3609 ( .A(n580), .B(n596), .Z(n547) );
  XNOR U3610 ( .A(n590), .B(n547), .Z(n541) );
  XNOR U3611 ( .A(x[121]), .B(n581), .Z(n540) );
  XNOR U3612 ( .A(n541), .B(n540), .Z(n542) );
  XOR U3613 ( .A(n543), .B(n542), .Z(n544) );
  XOR U3614 ( .A(n545), .B(n544), .Z(n565) );
  NAND U3615 ( .A(n563), .B(n565), .Z(n546) );
  NAND U3616 ( .A(n573), .B(n546), .Z(n557) );
  IV U3617 ( .A(n563), .Z(n564) );
  IV U3618 ( .A(n565), .Z(n571) );
  XOR U3619 ( .A(n547), .B(n601), .Z(n550) );
  AND U3620 ( .A(n590), .B(n581), .Z(n548) );
  XNOR U3621 ( .A(x[120]), .B(n548), .Z(n549) );
  XNOR U3622 ( .A(n550), .B(n549), .Z(n551) );
  XNOR U3623 ( .A(n552), .B(n551), .Z(n553) );
  XNOR U3624 ( .A(n554), .B(n553), .Z(n575) );
  IV U3625 ( .A(n575), .Z(n570) );
  XOR U3626 ( .A(n571), .B(n570), .Z(n555) );
  NAND U3627 ( .A(n564), .B(n555), .Z(n556) );
  AND U3628 ( .A(n557), .B(n556), .Z(n635) );
  NAND U3629 ( .A(n571), .B(n564), .Z(n558) );
  NAND U3630 ( .A(n570), .B(n558), .Z(n561) );
  XOR U3631 ( .A(n564), .B(n567), .Z(n559) );
  NAND U3632 ( .A(n565), .B(n559), .Z(n560) );
  AND U3633 ( .A(n561), .B(n560), .Z(n617) );
  XNOR U3634 ( .A(n635), .B(n617), .Z(n592) );
  OR U3635 ( .A(n592), .B(n562), .Z(n585) );
  NAND U3636 ( .A(n573), .B(n563), .Z(n569) );
  AND U3637 ( .A(n565), .B(n564), .Z(n572) );
  XNOR U3638 ( .A(n570), .B(n572), .Z(n566) );
  NAND U3639 ( .A(n567), .B(n566), .Z(n568) );
  AND U3640 ( .A(n569), .B(n568), .Z(n589) );
  NAND U3641 ( .A(n571), .B(n570), .Z(n577) );
  XNOR U3642 ( .A(n573), .B(n572), .Z(n574) );
  NAND U3643 ( .A(n575), .B(n574), .Z(n576) );
  NAND U3644 ( .A(n577), .B(n576), .Z(n629) );
  XNOR U3645 ( .A(n589), .B(n629), .Z(n607) );
  XOR U3646 ( .A(n607), .B(n592), .Z(n594) );
  OR U3647 ( .A(n594), .B(n578), .Z(n579) );
  XNOR U3648 ( .A(n585), .B(n579), .Z(n611) );
  XOR U3649 ( .A(n589), .B(n635), .Z(n597) );
  NANDN U3650 ( .A(n597), .B(n580), .Z(n637) );
  NANDN U3651 ( .A(n589), .B(n581), .Z(n582) );
  XNOR U3652 ( .A(n637), .B(n582), .Z(n615) );
  XOR U3653 ( .A(n611), .B(n615), .Z(n600) );
  NANDN U3654 ( .A(n583), .B(n607), .Z(n584) );
  XNOR U3655 ( .A(n585), .B(n584), .Z(n643) );
  XNOR U3656 ( .A(n629), .B(n617), .Z(n619) );
  NANDN U3657 ( .A(n619), .B(n586), .Z(n603) );
  NAND U3658 ( .A(n587), .B(n617), .Z(n588) );
  XNOR U3659 ( .A(n603), .B(n588), .Z(n634) );
  XOR U3660 ( .A(n643), .B(n634), .Z(n626) );
  XNOR U3661 ( .A(n600), .B(n626), .Z(z[120]) );
  ANDN U3662 ( .B(n590), .A(n589), .Z(n599) );
  NANDN U3663 ( .A(n592), .B(n591), .Z(n610) );
  NANDN U3664 ( .A(n594), .B(n593), .Z(n595) );
  XNOR U3665 ( .A(n610), .B(n595), .Z(n638) );
  NANDN U3666 ( .A(n597), .B(n596), .Z(n604) );
  XNOR U3667 ( .A(n638), .B(n604), .Z(n598) );
  XOR U3668 ( .A(n599), .B(n598), .Z(n624) );
  XOR U3669 ( .A(n624), .B(n600), .Z(n642) );
  ANDN U3670 ( .B(n635), .A(n601), .Z(n606) );
  NAND U3671 ( .A(n627), .B(n629), .Z(n602) );
  XNOR U3672 ( .A(n603), .B(n602), .Z(n614) );
  XNOR U3673 ( .A(n604), .B(n614), .Z(n605) );
  XNOR U3674 ( .A(n606), .B(n605), .Z(n613) );
  NAND U3675 ( .A(n608), .B(n607), .Z(n609) );
  XNOR U3676 ( .A(n610), .B(n609), .Z(n620) );
  XNOR U3677 ( .A(n611), .B(n620), .Z(n612) );
  XOR U3678 ( .A(n613), .B(n612), .Z(n623) );
  XNOR U3679 ( .A(n642), .B(n623), .Z(z[121]) );
  XNOR U3680 ( .A(n615), .B(n614), .Z(z[122]) );
  AND U3681 ( .A(n617), .B(n616), .Z(n622) );
  NANDN U3682 ( .A(n619), .B(n618), .Z(n632) );
  XNOR U3683 ( .A(n620), .B(n632), .Z(n621) );
  XOR U3684 ( .A(n622), .B(n621), .Z(n641) );
  XOR U3685 ( .A(n624), .B(n623), .Z(n625) );
  XOR U3686 ( .A(n641), .B(n625), .Z(z[123]) );
  XOR U3687 ( .A(n626), .B(z[122]), .Z(z[124]) );
  XNOR U3688 ( .A(n628), .B(n627), .Z(n630) );
  NAND U3689 ( .A(n630), .B(n629), .Z(n631) );
  XOR U3690 ( .A(n632), .B(n631), .Z(n633) );
  XNOR U3691 ( .A(n634), .B(n633), .Z(n640) );
  NAND U3692 ( .A(n635), .B(x[120]), .Z(n636) );
  XNOR U3693 ( .A(n637), .B(n636), .Z(n644) );
  XNOR U3694 ( .A(n638), .B(n644), .Z(n639) );
  XOR U3695 ( .A(n640), .B(n639), .Z(z[125]) );
  XNOR U3696 ( .A(n642), .B(n641), .Z(z[126]) );
  XNOR U3697 ( .A(n644), .B(n643), .Z(n645) );
  XNOR U3698 ( .A(z[121]), .B(n645), .Z(z[127]) );
  NOR U3699 ( .A(n647), .B(n646), .Z(n653) );
  NANDN U3700 ( .A(n648), .B(n672), .Z(n649) );
  XNOR U3701 ( .A(n650), .B(n649), .Z(n663) );
  XNOR U3702 ( .A(n651), .B(n663), .Z(n652) );
  XOR U3703 ( .A(n653), .B(n652), .Z(n1947) );
  XOR U3704 ( .A(n1947), .B(n654), .Z(z[12]) );
  XNOR U3705 ( .A(n656), .B(n655), .Z(n657) );
  NANDN U3706 ( .A(n658), .B(n657), .Z(n659) );
  XOR U3707 ( .A(n660), .B(n659), .Z(n661) );
  XNOR U3708 ( .A(n1947), .B(n661), .Z(n669) );
  ANDN U3709 ( .B(x[8]), .A(n662), .Z(n666) );
  XNOR U3710 ( .A(n664), .B(n663), .Z(n665) );
  XOR U3711 ( .A(n666), .B(n665), .Z(n683) );
  XNOR U3712 ( .A(n667), .B(n683), .Z(n668) );
  XOR U3713 ( .A(n669), .B(n668), .Z(z[13]) );
  XNOR U3714 ( .A(n671), .B(n670), .Z(n1948) );
  NAND U3715 ( .A(n673), .B(n672), .Z(n674) );
  XNOR U3716 ( .A(n675), .B(n674), .Z(n679) );
  XNOR U3717 ( .A(n1948), .B(n679), .Z(n676) );
  XOR U3718 ( .A(n677), .B(n676), .Z(z[14]) );
  XNOR U3719 ( .A(n679), .B(n678), .Z(n680) );
  XNOR U3720 ( .A(z[10]), .B(n680), .Z(n681) );
  XOR U3721 ( .A(n682), .B(n681), .Z(z[9]) );
  XNOR U3722 ( .A(n683), .B(z[9]), .Z(z[15]) );
  IV U3723 ( .A(x[17]), .Z(n815) );
  IV U3724 ( .A(n814), .Z(n686) );
  AND U3725 ( .A(n815), .B(n686), .Z(n693) );
  XNOR U3726 ( .A(x[19]), .B(n815), .Z(n689) );
  XNOR U3727 ( .A(x[18]), .B(n689), .Z(n684) );
  XNOR U3728 ( .A(n685), .B(n684), .Z(n749) );
  IV U3729 ( .A(n749), .Z(n695) );
  XNOR U3730 ( .A(n695), .B(n814), .Z(n748) );
  IV U3731 ( .A(x[23]), .Z(n687) );
  XNOR U3732 ( .A(x[17]), .B(n687), .Z(n780) );
  NAND U3733 ( .A(n748), .B(n780), .Z(n698) );
  XNOR U3734 ( .A(n687), .B(n686), .Z(n694) );
  IV U3735 ( .A(n694), .Z(n778) );
  XOR U3736 ( .A(n749), .B(n778), .Z(n714) );
  XNOR U3737 ( .A(n698), .B(n714), .Z(n691) );
  XOR U3738 ( .A(x[16]), .B(n695), .Z(n724) );
  XOR U3739 ( .A(x[20]), .B(n687), .Z(n688) );
  IV U3740 ( .A(n688), .Z(n753) );
  NANDN U3741 ( .A(n724), .B(n753), .Z(n697) );
  XNOR U3742 ( .A(n689), .B(n688), .Z(n742) );
  XNOR U3743 ( .A(n748), .B(n742), .Z(n740) );
  XOR U3744 ( .A(x[18]), .B(x[20]), .Z(n755) );
  NANDN U3745 ( .A(n740), .B(n755), .Z(n690) );
  XOR U3746 ( .A(n697), .B(n690), .Z(n716) );
  XNOR U3747 ( .A(n691), .B(n716), .Z(n692) );
  XOR U3748 ( .A(n693), .B(n692), .Z(n729) );
  IV U3749 ( .A(n729), .Z(n735) );
  AND U3750 ( .A(n695), .B(n694), .Z(n700) );
  XOR U3751 ( .A(x[16]), .B(n742), .Z(n743) );
  XNOR U3752 ( .A(n814), .B(n743), .Z(n745) );
  XOR U3753 ( .A(x[18]), .B(x[23]), .Z(n770) );
  NANDN U3754 ( .A(n745), .B(n770), .Z(n696) );
  XNOR U3755 ( .A(n697), .B(n696), .Z(n705) );
  XNOR U3756 ( .A(n698), .B(n705), .Z(n699) );
  XOR U3757 ( .A(n700), .B(n699), .Z(n725) );
  XNOR U3758 ( .A(x[20]), .B(n814), .Z(n763) );
  ANDN U3759 ( .B(x[16]), .A(n763), .Z(n707) );
  XOR U3760 ( .A(x[18]), .B(x[17]), .Z(n701) );
  XOR U3761 ( .A(n778), .B(n701), .Z(n752) );
  XOR U3762 ( .A(n753), .B(n701), .Z(n758) );
  NAND U3763 ( .A(n742), .B(n758), .Z(n709) );
  XNOR U3764 ( .A(n752), .B(n709), .Z(n703) );
  XNOR U3765 ( .A(x[17]), .B(n743), .Z(n702) );
  XNOR U3766 ( .A(n703), .B(n702), .Z(n704) );
  XOR U3767 ( .A(n705), .B(n704), .Z(n706) );
  XOR U3768 ( .A(n707), .B(n706), .Z(n727) );
  NAND U3769 ( .A(n725), .B(n727), .Z(n708) );
  NAND U3770 ( .A(n735), .B(n708), .Z(n719) );
  IV U3771 ( .A(n725), .Z(n726) );
  IV U3772 ( .A(n727), .Z(n733) );
  XOR U3773 ( .A(n709), .B(n763), .Z(n712) );
  AND U3774 ( .A(n752), .B(n743), .Z(n710) );
  XNOR U3775 ( .A(x[16]), .B(n710), .Z(n711) );
  XNOR U3776 ( .A(n712), .B(n711), .Z(n713) );
  XNOR U3777 ( .A(n714), .B(n713), .Z(n715) );
  XNOR U3778 ( .A(n716), .B(n715), .Z(n737) );
  IV U3779 ( .A(n737), .Z(n732) );
  XOR U3780 ( .A(n733), .B(n732), .Z(n717) );
  NAND U3781 ( .A(n726), .B(n717), .Z(n718) );
  AND U3782 ( .A(n719), .B(n718), .Z(n822) );
  NAND U3783 ( .A(n733), .B(n726), .Z(n720) );
  NAND U3784 ( .A(n732), .B(n720), .Z(n723) );
  XOR U3785 ( .A(n726), .B(n729), .Z(n721) );
  NAND U3786 ( .A(n727), .B(n721), .Z(n722) );
  AND U3787 ( .A(n723), .B(n722), .Z(n779) );
  XNOR U3788 ( .A(n822), .B(n779), .Z(n754) );
  OR U3789 ( .A(n754), .B(n724), .Z(n747) );
  NAND U3790 ( .A(n735), .B(n725), .Z(n731) );
  AND U3791 ( .A(n727), .B(n726), .Z(n734) );
  XNOR U3792 ( .A(n732), .B(n734), .Z(n728) );
  NAND U3793 ( .A(n729), .B(n728), .Z(n730) );
  AND U3794 ( .A(n731), .B(n730), .Z(n751) );
  NAND U3795 ( .A(n733), .B(n732), .Z(n739) );
  XNOR U3796 ( .A(n735), .B(n734), .Z(n736) );
  NAND U3797 ( .A(n737), .B(n736), .Z(n738) );
  NAND U3798 ( .A(n739), .B(n738), .Z(n816) );
  XNOR U3799 ( .A(n751), .B(n816), .Z(n769) );
  XOR U3800 ( .A(n769), .B(n754), .Z(n756) );
  OR U3801 ( .A(n756), .B(n740), .Z(n741) );
  XNOR U3802 ( .A(n747), .B(n741), .Z(n773) );
  XOR U3803 ( .A(n751), .B(n822), .Z(n759) );
  NANDN U3804 ( .A(n759), .B(n742), .Z(n824) );
  NANDN U3805 ( .A(n751), .B(n743), .Z(n744) );
  XNOR U3806 ( .A(n824), .B(n744), .Z(n777) );
  XOR U3807 ( .A(n773), .B(n777), .Z(n762) );
  NANDN U3808 ( .A(n745), .B(n769), .Z(n746) );
  XNOR U3809 ( .A(n747), .B(n746), .Z(n830) );
  XNOR U3810 ( .A(n816), .B(n779), .Z(n781) );
  NANDN U3811 ( .A(n781), .B(n748), .Z(n765) );
  NAND U3812 ( .A(n749), .B(n779), .Z(n750) );
  XNOR U3813 ( .A(n765), .B(n750), .Z(n821) );
  XOR U3814 ( .A(n830), .B(n821), .Z(n813) );
  XNOR U3815 ( .A(n762), .B(n813), .Z(z[16]) );
  ANDN U3816 ( .B(n752), .A(n751), .Z(n761) );
  NANDN U3817 ( .A(n754), .B(n753), .Z(n772) );
  NANDN U3818 ( .A(n756), .B(n755), .Z(n757) );
  XNOR U3819 ( .A(n772), .B(n757), .Z(n825) );
  NANDN U3820 ( .A(n759), .B(n758), .Z(n766) );
  XNOR U3821 ( .A(n825), .B(n766), .Z(n760) );
  XOR U3822 ( .A(n761), .B(n760), .Z(n786) );
  XOR U3823 ( .A(n786), .B(n762), .Z(n829) );
  ANDN U3824 ( .B(n822), .A(n763), .Z(n768) );
  NAND U3825 ( .A(n814), .B(n816), .Z(n764) );
  XNOR U3826 ( .A(n765), .B(n764), .Z(n776) );
  XNOR U3827 ( .A(n766), .B(n776), .Z(n767) );
  XNOR U3828 ( .A(n768), .B(n767), .Z(n775) );
  NAND U3829 ( .A(n770), .B(n769), .Z(n771) );
  XNOR U3830 ( .A(n772), .B(n771), .Z(n782) );
  XNOR U3831 ( .A(n773), .B(n782), .Z(n774) );
  XOR U3832 ( .A(n775), .B(n774), .Z(n785) );
  XNOR U3833 ( .A(n829), .B(n785), .Z(z[17]) );
  XNOR U3834 ( .A(n777), .B(n776), .Z(z[18]) );
  AND U3835 ( .A(n779), .B(n778), .Z(n784) );
  NANDN U3836 ( .A(n781), .B(n780), .Z(n819) );
  XNOR U3837 ( .A(n782), .B(n819), .Z(n783) );
  XOR U3838 ( .A(n784), .B(n783), .Z(n828) );
  XOR U3839 ( .A(n786), .B(n785), .Z(n787) );
  XOR U3840 ( .A(n828), .B(n787), .Z(z[19]) );
  ANDN U3841 ( .B(n789), .A(n788), .Z(n798) );
  NANDN U3842 ( .A(n791), .B(n790), .Z(n809) );
  NANDN U3843 ( .A(n793), .B(n792), .Z(n794) );
  XNOR U3844 ( .A(n809), .B(n794), .Z(n1457) );
  NANDN U3845 ( .A(n796), .B(n795), .Z(n803) );
  XNOR U3846 ( .A(n1457), .B(n803), .Z(n797) );
  XOR U3847 ( .A(n798), .B(n797), .Z(n1091) );
  XOR U3848 ( .A(n1091), .B(n799), .Z(n1600) );
  ANDN U3849 ( .B(n1454), .A(n800), .Z(n805) );
  NAND U3850 ( .A(n1446), .B(n1448), .Z(n801) );
  XNOR U3851 ( .A(n802), .B(n801), .Z(n952) );
  XNOR U3852 ( .A(n803), .B(n952), .Z(n804) );
  XNOR U3853 ( .A(n805), .B(n804), .Z(n812) );
  NAND U3854 ( .A(n807), .B(n806), .Z(n808) );
  XNOR U3855 ( .A(n809), .B(n808), .Z(n1087) );
  XNOR U3856 ( .A(n810), .B(n1087), .Z(n811) );
  XOR U3857 ( .A(n812), .B(n811), .Z(n1090) );
  XNOR U3858 ( .A(n1600), .B(n1090), .Z(z[1]) );
  XOR U3859 ( .A(n813), .B(z[18]), .Z(z[20]) );
  XNOR U3860 ( .A(n815), .B(n814), .Z(n817) );
  NAND U3861 ( .A(n817), .B(n816), .Z(n818) );
  XOR U3862 ( .A(n819), .B(n818), .Z(n820) );
  XNOR U3863 ( .A(n821), .B(n820), .Z(n827) );
  NAND U3864 ( .A(n822), .B(x[16]), .Z(n823) );
  XNOR U3865 ( .A(n824), .B(n823), .Z(n831) );
  XNOR U3866 ( .A(n825), .B(n831), .Z(n826) );
  XOR U3867 ( .A(n827), .B(n826), .Z(z[21]) );
  XNOR U3868 ( .A(n829), .B(n828), .Z(z[22]) );
  XNOR U3869 ( .A(n831), .B(n830), .Z(n832) );
  XNOR U3870 ( .A(z[17]), .B(n832), .Z(z[23]) );
  IV U3871 ( .A(x[25]), .Z(n939) );
  XOR U3872 ( .A(x[24]), .B(x[30]), .Z(n834) );
  XOR U3873 ( .A(x[29]), .B(n834), .Z(n938) );
  IV U3874 ( .A(n938), .Z(n835) );
  AND U3875 ( .A(n939), .B(n835), .Z(n842) );
  XNOR U3876 ( .A(x[27]), .B(n939), .Z(n838) );
  XNOR U3877 ( .A(x[26]), .B(n838), .Z(n833) );
  XNOR U3878 ( .A(n834), .B(n833), .Z(n898) );
  IV U3879 ( .A(n898), .Z(n844) );
  XNOR U3880 ( .A(n844), .B(n938), .Z(n897) );
  IV U3881 ( .A(x[31]), .Z(n836) );
  XNOR U3882 ( .A(x[25]), .B(n836), .Z(n929) );
  NAND U3883 ( .A(n897), .B(n929), .Z(n847) );
  XNOR U3884 ( .A(n836), .B(n835), .Z(n843) );
  IV U3885 ( .A(n843), .Z(n927) );
  XOR U3886 ( .A(n898), .B(n927), .Z(n863) );
  XNOR U3887 ( .A(n847), .B(n863), .Z(n840) );
  XOR U3888 ( .A(x[24]), .B(n844), .Z(n873) );
  XOR U3889 ( .A(x[28]), .B(n836), .Z(n837) );
  IV U3890 ( .A(n837), .Z(n902) );
  NANDN U3891 ( .A(n873), .B(n902), .Z(n846) );
  XNOR U3892 ( .A(n838), .B(n837), .Z(n891) );
  XNOR U3893 ( .A(n897), .B(n891), .Z(n889) );
  XOR U3894 ( .A(x[26]), .B(x[28]), .Z(n904) );
  NANDN U3895 ( .A(n889), .B(n904), .Z(n839) );
  XOR U3896 ( .A(n846), .B(n839), .Z(n865) );
  XNOR U3897 ( .A(n840), .B(n865), .Z(n841) );
  XOR U3898 ( .A(n842), .B(n841), .Z(n878) );
  IV U3899 ( .A(n878), .Z(n884) );
  AND U3900 ( .A(n844), .B(n843), .Z(n849) );
  XOR U3901 ( .A(x[24]), .B(n891), .Z(n892) );
  XNOR U3902 ( .A(n938), .B(n892), .Z(n894) );
  XOR U3903 ( .A(x[26]), .B(x[31]), .Z(n919) );
  NANDN U3904 ( .A(n894), .B(n919), .Z(n845) );
  XNOR U3905 ( .A(n846), .B(n845), .Z(n854) );
  XNOR U3906 ( .A(n847), .B(n854), .Z(n848) );
  XOR U3907 ( .A(n849), .B(n848), .Z(n874) );
  XNOR U3908 ( .A(x[28]), .B(n938), .Z(n912) );
  ANDN U3909 ( .B(x[24]), .A(n912), .Z(n856) );
  XOR U3910 ( .A(x[26]), .B(x[25]), .Z(n850) );
  XOR U3911 ( .A(n927), .B(n850), .Z(n901) );
  XOR U3912 ( .A(n902), .B(n850), .Z(n907) );
  NAND U3913 ( .A(n891), .B(n907), .Z(n858) );
  XNOR U3914 ( .A(n901), .B(n858), .Z(n852) );
  XNOR U3915 ( .A(x[25]), .B(n892), .Z(n851) );
  XNOR U3916 ( .A(n852), .B(n851), .Z(n853) );
  XOR U3917 ( .A(n854), .B(n853), .Z(n855) );
  XOR U3918 ( .A(n856), .B(n855), .Z(n876) );
  NAND U3919 ( .A(n874), .B(n876), .Z(n857) );
  NAND U3920 ( .A(n884), .B(n857), .Z(n868) );
  IV U3921 ( .A(n874), .Z(n875) );
  IV U3922 ( .A(n876), .Z(n882) );
  XOR U3923 ( .A(n858), .B(n912), .Z(n861) );
  AND U3924 ( .A(n901), .B(n892), .Z(n859) );
  XNOR U3925 ( .A(x[24]), .B(n859), .Z(n860) );
  XNOR U3926 ( .A(n861), .B(n860), .Z(n862) );
  XNOR U3927 ( .A(n863), .B(n862), .Z(n864) );
  XNOR U3928 ( .A(n865), .B(n864), .Z(n886) );
  IV U3929 ( .A(n886), .Z(n881) );
  XOR U3930 ( .A(n882), .B(n881), .Z(n866) );
  NAND U3931 ( .A(n875), .B(n866), .Z(n867) );
  AND U3932 ( .A(n868), .B(n867), .Z(n946) );
  NAND U3933 ( .A(n882), .B(n875), .Z(n869) );
  NAND U3934 ( .A(n881), .B(n869), .Z(n872) );
  XOR U3935 ( .A(n875), .B(n878), .Z(n870) );
  NAND U3936 ( .A(n876), .B(n870), .Z(n871) );
  AND U3937 ( .A(n872), .B(n871), .Z(n928) );
  XNOR U3938 ( .A(n946), .B(n928), .Z(n903) );
  OR U3939 ( .A(n903), .B(n873), .Z(n896) );
  NAND U3940 ( .A(n884), .B(n874), .Z(n880) );
  AND U3941 ( .A(n876), .B(n875), .Z(n883) );
  XNOR U3942 ( .A(n881), .B(n883), .Z(n877) );
  NAND U3943 ( .A(n878), .B(n877), .Z(n879) );
  AND U3944 ( .A(n880), .B(n879), .Z(n900) );
  NAND U3945 ( .A(n882), .B(n881), .Z(n888) );
  XNOR U3946 ( .A(n884), .B(n883), .Z(n885) );
  NAND U3947 ( .A(n886), .B(n885), .Z(n887) );
  NAND U3948 ( .A(n888), .B(n887), .Z(n940) );
  XNOR U3949 ( .A(n900), .B(n940), .Z(n918) );
  XOR U3950 ( .A(n918), .B(n903), .Z(n905) );
  OR U3951 ( .A(n905), .B(n889), .Z(n890) );
  XNOR U3952 ( .A(n896), .B(n890), .Z(n922) );
  XOR U3953 ( .A(n900), .B(n946), .Z(n908) );
  NANDN U3954 ( .A(n908), .B(n891), .Z(n948) );
  NANDN U3955 ( .A(n900), .B(n892), .Z(n893) );
  XNOR U3956 ( .A(n948), .B(n893), .Z(n926) );
  XOR U3957 ( .A(n922), .B(n926), .Z(n911) );
  NANDN U3958 ( .A(n894), .B(n918), .Z(n895) );
  XNOR U3959 ( .A(n896), .B(n895), .Z(n956) );
  XNOR U3960 ( .A(n940), .B(n928), .Z(n930) );
  NANDN U3961 ( .A(n930), .B(n897), .Z(n914) );
  NAND U3962 ( .A(n898), .B(n928), .Z(n899) );
  XNOR U3963 ( .A(n914), .B(n899), .Z(n945) );
  XOR U3964 ( .A(n956), .B(n945), .Z(n937) );
  XNOR U3965 ( .A(n911), .B(n937), .Z(z[24]) );
  ANDN U3966 ( .B(n901), .A(n900), .Z(n910) );
  NANDN U3967 ( .A(n903), .B(n902), .Z(n921) );
  NANDN U3968 ( .A(n905), .B(n904), .Z(n906) );
  XNOR U3969 ( .A(n921), .B(n906), .Z(n949) );
  NANDN U3970 ( .A(n908), .B(n907), .Z(n915) );
  XNOR U3971 ( .A(n949), .B(n915), .Z(n909) );
  XOR U3972 ( .A(n910), .B(n909), .Z(n935) );
  XOR U3973 ( .A(n935), .B(n911), .Z(n955) );
  ANDN U3974 ( .B(n946), .A(n912), .Z(n917) );
  NAND U3975 ( .A(n938), .B(n940), .Z(n913) );
  XNOR U3976 ( .A(n914), .B(n913), .Z(n925) );
  XNOR U3977 ( .A(n915), .B(n925), .Z(n916) );
  XNOR U3978 ( .A(n917), .B(n916), .Z(n924) );
  NAND U3979 ( .A(n919), .B(n918), .Z(n920) );
  XNOR U3980 ( .A(n921), .B(n920), .Z(n931) );
  XNOR U3981 ( .A(n922), .B(n931), .Z(n923) );
  XOR U3982 ( .A(n924), .B(n923), .Z(n934) );
  XNOR U3983 ( .A(n955), .B(n934), .Z(z[25]) );
  XNOR U3984 ( .A(n926), .B(n925), .Z(z[26]) );
  AND U3985 ( .A(n928), .B(n927), .Z(n933) );
  NANDN U3986 ( .A(n930), .B(n929), .Z(n943) );
  XNOR U3987 ( .A(n931), .B(n943), .Z(n932) );
  XOR U3988 ( .A(n933), .B(n932), .Z(n954) );
  XOR U3989 ( .A(n935), .B(n934), .Z(n936) );
  XOR U3990 ( .A(n954), .B(n936), .Z(z[27]) );
  XOR U3991 ( .A(n937), .B(z[26]), .Z(z[28]) );
  XNOR U3992 ( .A(n939), .B(n938), .Z(n941) );
  NAND U3993 ( .A(n941), .B(n940), .Z(n942) );
  XOR U3994 ( .A(n943), .B(n942), .Z(n944) );
  XNOR U3995 ( .A(n945), .B(n944), .Z(n951) );
  NAND U3996 ( .A(n946), .B(x[24]), .Z(n947) );
  XNOR U3997 ( .A(n948), .B(n947), .Z(n957) );
  XNOR U3998 ( .A(n949), .B(n957), .Z(n950) );
  XOR U3999 ( .A(n951), .B(n950), .Z(z[29]) );
  XNOR U4000 ( .A(n953), .B(n952), .Z(z[2]) );
  XNOR U4001 ( .A(n955), .B(n954), .Z(z[30]) );
  XNOR U4002 ( .A(n957), .B(n956), .Z(n958) );
  XNOR U4003 ( .A(z[25]), .B(n958), .Z(z[31]) );
  IV U4004 ( .A(x[33]), .Z(n1065) );
  XOR U4005 ( .A(x[32]), .B(x[38]), .Z(n960) );
  XOR U4006 ( .A(x[37]), .B(n960), .Z(n1064) );
  IV U4007 ( .A(n1064), .Z(n961) );
  AND U4008 ( .A(n1065), .B(n961), .Z(n968) );
  XNOR U4009 ( .A(x[35]), .B(n1065), .Z(n964) );
  XNOR U4010 ( .A(x[34]), .B(n964), .Z(n959) );
  XNOR U4011 ( .A(n960), .B(n959), .Z(n1024) );
  IV U4012 ( .A(n1024), .Z(n970) );
  XNOR U4013 ( .A(n970), .B(n1064), .Z(n1023) );
  IV U4014 ( .A(x[39]), .Z(n962) );
  XNOR U4015 ( .A(x[33]), .B(n962), .Z(n1055) );
  NAND U4016 ( .A(n1023), .B(n1055), .Z(n973) );
  XNOR U4017 ( .A(n962), .B(n961), .Z(n969) );
  IV U4018 ( .A(n969), .Z(n1053) );
  XOR U4019 ( .A(n1024), .B(n1053), .Z(n989) );
  XNOR U4020 ( .A(n973), .B(n989), .Z(n966) );
  XOR U4021 ( .A(x[32]), .B(n970), .Z(n999) );
  XOR U4022 ( .A(x[36]), .B(n962), .Z(n963) );
  IV U4023 ( .A(n963), .Z(n1028) );
  NANDN U4024 ( .A(n999), .B(n1028), .Z(n972) );
  XNOR U4025 ( .A(n964), .B(n963), .Z(n1017) );
  XNOR U4026 ( .A(n1023), .B(n1017), .Z(n1015) );
  XOR U4027 ( .A(x[34]), .B(x[36]), .Z(n1030) );
  NANDN U4028 ( .A(n1015), .B(n1030), .Z(n965) );
  XOR U4029 ( .A(n972), .B(n965), .Z(n991) );
  XNOR U4030 ( .A(n966), .B(n991), .Z(n967) );
  XOR U4031 ( .A(n968), .B(n967), .Z(n1004) );
  IV U4032 ( .A(n1004), .Z(n1010) );
  AND U4033 ( .A(n970), .B(n969), .Z(n975) );
  XOR U4034 ( .A(x[32]), .B(n1017), .Z(n1018) );
  XNOR U4035 ( .A(n1064), .B(n1018), .Z(n1020) );
  XOR U4036 ( .A(x[34]), .B(x[39]), .Z(n1045) );
  NANDN U4037 ( .A(n1020), .B(n1045), .Z(n971) );
  XNOR U4038 ( .A(n972), .B(n971), .Z(n980) );
  XNOR U4039 ( .A(n973), .B(n980), .Z(n974) );
  XOR U4040 ( .A(n975), .B(n974), .Z(n1000) );
  XNOR U4041 ( .A(x[36]), .B(n1064), .Z(n1038) );
  ANDN U4042 ( .B(x[32]), .A(n1038), .Z(n982) );
  XOR U4043 ( .A(x[34]), .B(x[33]), .Z(n976) );
  XOR U4044 ( .A(n1053), .B(n976), .Z(n1027) );
  XOR U4045 ( .A(n1028), .B(n976), .Z(n1033) );
  NAND U4046 ( .A(n1017), .B(n1033), .Z(n984) );
  XNOR U4047 ( .A(n1027), .B(n984), .Z(n978) );
  XNOR U4048 ( .A(x[33]), .B(n1018), .Z(n977) );
  XNOR U4049 ( .A(n978), .B(n977), .Z(n979) );
  XOR U4050 ( .A(n980), .B(n979), .Z(n981) );
  XOR U4051 ( .A(n982), .B(n981), .Z(n1002) );
  NAND U4052 ( .A(n1000), .B(n1002), .Z(n983) );
  NAND U4053 ( .A(n1010), .B(n983), .Z(n994) );
  IV U4054 ( .A(n1000), .Z(n1001) );
  IV U4055 ( .A(n1002), .Z(n1008) );
  XOR U4056 ( .A(n984), .B(n1038), .Z(n987) );
  AND U4057 ( .A(n1027), .B(n1018), .Z(n985) );
  XNOR U4058 ( .A(x[32]), .B(n985), .Z(n986) );
  XNOR U4059 ( .A(n987), .B(n986), .Z(n988) );
  XNOR U4060 ( .A(n989), .B(n988), .Z(n990) );
  XNOR U4061 ( .A(n991), .B(n990), .Z(n1012) );
  IV U4062 ( .A(n1012), .Z(n1007) );
  XOR U4063 ( .A(n1008), .B(n1007), .Z(n992) );
  NAND U4064 ( .A(n1001), .B(n992), .Z(n993) );
  AND U4065 ( .A(n994), .B(n993), .Z(n1072) );
  NAND U4066 ( .A(n1008), .B(n1001), .Z(n995) );
  NAND U4067 ( .A(n1007), .B(n995), .Z(n998) );
  XOR U4068 ( .A(n1001), .B(n1004), .Z(n996) );
  NAND U4069 ( .A(n1002), .B(n996), .Z(n997) );
  AND U4070 ( .A(n998), .B(n997), .Z(n1054) );
  XNOR U4071 ( .A(n1072), .B(n1054), .Z(n1029) );
  OR U4072 ( .A(n1029), .B(n999), .Z(n1022) );
  NAND U4073 ( .A(n1010), .B(n1000), .Z(n1006) );
  AND U4074 ( .A(n1002), .B(n1001), .Z(n1009) );
  XNOR U4075 ( .A(n1007), .B(n1009), .Z(n1003) );
  NAND U4076 ( .A(n1004), .B(n1003), .Z(n1005) );
  AND U4077 ( .A(n1006), .B(n1005), .Z(n1026) );
  NAND U4078 ( .A(n1008), .B(n1007), .Z(n1014) );
  XNOR U4079 ( .A(n1010), .B(n1009), .Z(n1011) );
  NAND U4080 ( .A(n1012), .B(n1011), .Z(n1013) );
  NAND U4081 ( .A(n1014), .B(n1013), .Z(n1066) );
  XNOR U4082 ( .A(n1026), .B(n1066), .Z(n1044) );
  XOR U4083 ( .A(n1044), .B(n1029), .Z(n1031) );
  OR U4084 ( .A(n1031), .B(n1015), .Z(n1016) );
  XNOR U4085 ( .A(n1022), .B(n1016), .Z(n1048) );
  XOR U4086 ( .A(n1026), .B(n1072), .Z(n1034) );
  NANDN U4087 ( .A(n1034), .B(n1017), .Z(n1074) );
  NANDN U4088 ( .A(n1026), .B(n1018), .Z(n1019) );
  XNOR U4089 ( .A(n1074), .B(n1019), .Z(n1052) );
  XOR U4090 ( .A(n1048), .B(n1052), .Z(n1037) );
  NANDN U4091 ( .A(n1020), .B(n1044), .Z(n1021) );
  XNOR U4092 ( .A(n1022), .B(n1021), .Z(n1080) );
  XNOR U4093 ( .A(n1066), .B(n1054), .Z(n1056) );
  NANDN U4094 ( .A(n1056), .B(n1023), .Z(n1040) );
  NAND U4095 ( .A(n1024), .B(n1054), .Z(n1025) );
  XNOR U4096 ( .A(n1040), .B(n1025), .Z(n1071) );
  XOR U4097 ( .A(n1080), .B(n1071), .Z(n1063) );
  XNOR U4098 ( .A(n1037), .B(n1063), .Z(z[32]) );
  ANDN U4099 ( .B(n1027), .A(n1026), .Z(n1036) );
  NANDN U4100 ( .A(n1029), .B(n1028), .Z(n1047) );
  NANDN U4101 ( .A(n1031), .B(n1030), .Z(n1032) );
  XNOR U4102 ( .A(n1047), .B(n1032), .Z(n1075) );
  NANDN U4103 ( .A(n1034), .B(n1033), .Z(n1041) );
  XNOR U4104 ( .A(n1075), .B(n1041), .Z(n1035) );
  XOR U4105 ( .A(n1036), .B(n1035), .Z(n1061) );
  XOR U4106 ( .A(n1061), .B(n1037), .Z(n1079) );
  ANDN U4107 ( .B(n1072), .A(n1038), .Z(n1043) );
  NAND U4108 ( .A(n1064), .B(n1066), .Z(n1039) );
  XNOR U4109 ( .A(n1040), .B(n1039), .Z(n1051) );
  XNOR U4110 ( .A(n1041), .B(n1051), .Z(n1042) );
  XNOR U4111 ( .A(n1043), .B(n1042), .Z(n1050) );
  NAND U4112 ( .A(n1045), .B(n1044), .Z(n1046) );
  XNOR U4113 ( .A(n1047), .B(n1046), .Z(n1057) );
  XNOR U4114 ( .A(n1048), .B(n1057), .Z(n1049) );
  XOR U4115 ( .A(n1050), .B(n1049), .Z(n1060) );
  XNOR U4116 ( .A(n1079), .B(n1060), .Z(z[33]) );
  XNOR U4117 ( .A(n1052), .B(n1051), .Z(z[34]) );
  AND U4118 ( .A(n1054), .B(n1053), .Z(n1059) );
  NANDN U4119 ( .A(n1056), .B(n1055), .Z(n1069) );
  XNOR U4120 ( .A(n1057), .B(n1069), .Z(n1058) );
  XOR U4121 ( .A(n1059), .B(n1058), .Z(n1078) );
  XOR U4122 ( .A(n1061), .B(n1060), .Z(n1062) );
  XOR U4123 ( .A(n1078), .B(n1062), .Z(z[35]) );
  XOR U4124 ( .A(n1063), .B(z[34]), .Z(z[36]) );
  XNOR U4125 ( .A(n1065), .B(n1064), .Z(n1067) );
  NAND U4126 ( .A(n1067), .B(n1066), .Z(n1068) );
  XOR U4127 ( .A(n1069), .B(n1068), .Z(n1070) );
  XNOR U4128 ( .A(n1071), .B(n1070), .Z(n1077) );
  NAND U4129 ( .A(n1072), .B(x[32]), .Z(n1073) );
  XNOR U4130 ( .A(n1074), .B(n1073), .Z(n1081) );
  XNOR U4131 ( .A(n1075), .B(n1081), .Z(n1076) );
  XOR U4132 ( .A(n1077), .B(n1076), .Z(z[37]) );
  XNOR U4133 ( .A(n1079), .B(n1078), .Z(z[38]) );
  XNOR U4134 ( .A(n1081), .B(n1080), .Z(n1082) );
  XNOR U4135 ( .A(z[33]), .B(n1082), .Z(z[39]) );
  AND U4136 ( .A(n1084), .B(n1083), .Z(n1089) );
  NANDN U4137 ( .A(n1086), .B(n1085), .Z(n1451) );
  XNOR U4138 ( .A(n1087), .B(n1451), .Z(n1088) );
  XOR U4139 ( .A(n1089), .B(n1088), .Z(n1599) );
  XOR U4140 ( .A(n1091), .B(n1090), .Z(n1092) );
  XOR U4141 ( .A(n1599), .B(n1092), .Z(z[3]) );
  IV U4142 ( .A(x[41]), .Z(n1199) );
  XOR U4143 ( .A(x[40]), .B(x[46]), .Z(n1094) );
  XOR U4144 ( .A(x[45]), .B(n1094), .Z(n1198) );
  IV U4145 ( .A(n1198), .Z(n1095) );
  AND U4146 ( .A(n1199), .B(n1095), .Z(n1102) );
  XNOR U4147 ( .A(x[43]), .B(n1199), .Z(n1098) );
  XNOR U4148 ( .A(x[42]), .B(n1098), .Z(n1093) );
  XNOR U4149 ( .A(n1094), .B(n1093), .Z(n1158) );
  IV U4150 ( .A(n1158), .Z(n1104) );
  XNOR U4151 ( .A(n1104), .B(n1198), .Z(n1157) );
  IV U4152 ( .A(x[47]), .Z(n1096) );
  XNOR U4153 ( .A(x[41]), .B(n1096), .Z(n1189) );
  NAND U4154 ( .A(n1157), .B(n1189), .Z(n1107) );
  XNOR U4155 ( .A(n1096), .B(n1095), .Z(n1103) );
  IV U4156 ( .A(n1103), .Z(n1187) );
  XOR U4157 ( .A(n1158), .B(n1187), .Z(n1123) );
  XNOR U4158 ( .A(n1107), .B(n1123), .Z(n1100) );
  XOR U4159 ( .A(x[40]), .B(n1104), .Z(n1133) );
  XOR U4160 ( .A(x[44]), .B(n1096), .Z(n1097) );
  IV U4161 ( .A(n1097), .Z(n1162) );
  NANDN U4162 ( .A(n1133), .B(n1162), .Z(n1106) );
  XNOR U4163 ( .A(n1098), .B(n1097), .Z(n1151) );
  XNOR U4164 ( .A(n1157), .B(n1151), .Z(n1149) );
  XOR U4165 ( .A(x[42]), .B(x[44]), .Z(n1164) );
  NANDN U4166 ( .A(n1149), .B(n1164), .Z(n1099) );
  XOR U4167 ( .A(n1106), .B(n1099), .Z(n1125) );
  XNOR U4168 ( .A(n1100), .B(n1125), .Z(n1101) );
  XOR U4169 ( .A(n1102), .B(n1101), .Z(n1138) );
  IV U4170 ( .A(n1138), .Z(n1144) );
  AND U4171 ( .A(n1104), .B(n1103), .Z(n1109) );
  XOR U4172 ( .A(x[40]), .B(n1151), .Z(n1152) );
  XNOR U4173 ( .A(n1198), .B(n1152), .Z(n1154) );
  XOR U4174 ( .A(x[42]), .B(x[47]), .Z(n1179) );
  NANDN U4175 ( .A(n1154), .B(n1179), .Z(n1105) );
  XNOR U4176 ( .A(n1106), .B(n1105), .Z(n1114) );
  XNOR U4177 ( .A(n1107), .B(n1114), .Z(n1108) );
  XOR U4178 ( .A(n1109), .B(n1108), .Z(n1134) );
  XNOR U4179 ( .A(x[44]), .B(n1198), .Z(n1172) );
  ANDN U4180 ( .B(x[40]), .A(n1172), .Z(n1116) );
  XOR U4181 ( .A(x[42]), .B(x[41]), .Z(n1110) );
  XOR U4182 ( .A(n1187), .B(n1110), .Z(n1161) );
  XOR U4183 ( .A(n1162), .B(n1110), .Z(n1167) );
  NAND U4184 ( .A(n1151), .B(n1167), .Z(n1118) );
  XNOR U4185 ( .A(n1161), .B(n1118), .Z(n1112) );
  XNOR U4186 ( .A(x[41]), .B(n1152), .Z(n1111) );
  XNOR U4187 ( .A(n1112), .B(n1111), .Z(n1113) );
  XOR U4188 ( .A(n1114), .B(n1113), .Z(n1115) );
  XOR U4189 ( .A(n1116), .B(n1115), .Z(n1136) );
  NAND U4190 ( .A(n1134), .B(n1136), .Z(n1117) );
  NAND U4191 ( .A(n1144), .B(n1117), .Z(n1128) );
  IV U4192 ( .A(n1134), .Z(n1135) );
  IV U4193 ( .A(n1136), .Z(n1142) );
  XOR U4194 ( .A(n1118), .B(n1172), .Z(n1121) );
  AND U4195 ( .A(n1161), .B(n1152), .Z(n1119) );
  XNOR U4196 ( .A(x[40]), .B(n1119), .Z(n1120) );
  XNOR U4197 ( .A(n1121), .B(n1120), .Z(n1122) );
  XNOR U4198 ( .A(n1123), .B(n1122), .Z(n1124) );
  XNOR U4199 ( .A(n1125), .B(n1124), .Z(n1146) );
  IV U4200 ( .A(n1146), .Z(n1141) );
  XOR U4201 ( .A(n1142), .B(n1141), .Z(n1126) );
  NAND U4202 ( .A(n1135), .B(n1126), .Z(n1127) );
  AND U4203 ( .A(n1128), .B(n1127), .Z(n1206) );
  NAND U4204 ( .A(n1142), .B(n1135), .Z(n1129) );
  NAND U4205 ( .A(n1141), .B(n1129), .Z(n1132) );
  XOR U4206 ( .A(n1135), .B(n1138), .Z(n1130) );
  NAND U4207 ( .A(n1136), .B(n1130), .Z(n1131) );
  AND U4208 ( .A(n1132), .B(n1131), .Z(n1188) );
  XNOR U4209 ( .A(n1206), .B(n1188), .Z(n1163) );
  OR U4210 ( .A(n1163), .B(n1133), .Z(n1156) );
  NAND U4211 ( .A(n1144), .B(n1134), .Z(n1140) );
  AND U4212 ( .A(n1136), .B(n1135), .Z(n1143) );
  XNOR U4213 ( .A(n1141), .B(n1143), .Z(n1137) );
  NAND U4214 ( .A(n1138), .B(n1137), .Z(n1139) );
  AND U4215 ( .A(n1140), .B(n1139), .Z(n1160) );
  NAND U4216 ( .A(n1142), .B(n1141), .Z(n1148) );
  XNOR U4217 ( .A(n1144), .B(n1143), .Z(n1145) );
  NAND U4218 ( .A(n1146), .B(n1145), .Z(n1147) );
  NAND U4219 ( .A(n1148), .B(n1147), .Z(n1200) );
  XNOR U4220 ( .A(n1160), .B(n1200), .Z(n1178) );
  XOR U4221 ( .A(n1178), .B(n1163), .Z(n1165) );
  OR U4222 ( .A(n1165), .B(n1149), .Z(n1150) );
  XNOR U4223 ( .A(n1156), .B(n1150), .Z(n1182) );
  XOR U4224 ( .A(n1160), .B(n1206), .Z(n1168) );
  NANDN U4225 ( .A(n1168), .B(n1151), .Z(n1208) );
  NANDN U4226 ( .A(n1160), .B(n1152), .Z(n1153) );
  XNOR U4227 ( .A(n1208), .B(n1153), .Z(n1186) );
  XOR U4228 ( .A(n1182), .B(n1186), .Z(n1171) );
  NANDN U4229 ( .A(n1154), .B(n1178), .Z(n1155) );
  XNOR U4230 ( .A(n1156), .B(n1155), .Z(n1214) );
  XNOR U4231 ( .A(n1200), .B(n1188), .Z(n1190) );
  NANDN U4232 ( .A(n1190), .B(n1157), .Z(n1174) );
  NAND U4233 ( .A(n1158), .B(n1188), .Z(n1159) );
  XNOR U4234 ( .A(n1174), .B(n1159), .Z(n1205) );
  XOR U4235 ( .A(n1214), .B(n1205), .Z(n1197) );
  XNOR U4236 ( .A(n1171), .B(n1197), .Z(z[40]) );
  ANDN U4237 ( .B(n1161), .A(n1160), .Z(n1170) );
  NANDN U4238 ( .A(n1163), .B(n1162), .Z(n1181) );
  NANDN U4239 ( .A(n1165), .B(n1164), .Z(n1166) );
  XNOR U4240 ( .A(n1181), .B(n1166), .Z(n1209) );
  NANDN U4241 ( .A(n1168), .B(n1167), .Z(n1175) );
  XNOR U4242 ( .A(n1209), .B(n1175), .Z(n1169) );
  XOR U4243 ( .A(n1170), .B(n1169), .Z(n1195) );
  XOR U4244 ( .A(n1195), .B(n1171), .Z(n1213) );
  ANDN U4245 ( .B(n1206), .A(n1172), .Z(n1177) );
  NAND U4246 ( .A(n1198), .B(n1200), .Z(n1173) );
  XNOR U4247 ( .A(n1174), .B(n1173), .Z(n1185) );
  XNOR U4248 ( .A(n1175), .B(n1185), .Z(n1176) );
  XNOR U4249 ( .A(n1177), .B(n1176), .Z(n1184) );
  NAND U4250 ( .A(n1179), .B(n1178), .Z(n1180) );
  XNOR U4251 ( .A(n1181), .B(n1180), .Z(n1191) );
  XNOR U4252 ( .A(n1182), .B(n1191), .Z(n1183) );
  XOR U4253 ( .A(n1184), .B(n1183), .Z(n1194) );
  XNOR U4254 ( .A(n1213), .B(n1194), .Z(z[41]) );
  XNOR U4255 ( .A(n1186), .B(n1185), .Z(z[42]) );
  AND U4256 ( .A(n1188), .B(n1187), .Z(n1193) );
  NANDN U4257 ( .A(n1190), .B(n1189), .Z(n1203) );
  XNOR U4258 ( .A(n1191), .B(n1203), .Z(n1192) );
  XOR U4259 ( .A(n1193), .B(n1192), .Z(n1212) );
  XOR U4260 ( .A(n1195), .B(n1194), .Z(n1196) );
  XOR U4261 ( .A(n1212), .B(n1196), .Z(z[43]) );
  XOR U4262 ( .A(n1197), .B(z[42]), .Z(z[44]) );
  XNOR U4263 ( .A(n1199), .B(n1198), .Z(n1201) );
  NAND U4264 ( .A(n1201), .B(n1200), .Z(n1202) );
  XOR U4265 ( .A(n1203), .B(n1202), .Z(n1204) );
  XNOR U4266 ( .A(n1205), .B(n1204), .Z(n1211) );
  NAND U4267 ( .A(n1206), .B(x[40]), .Z(n1207) );
  XNOR U4268 ( .A(n1208), .B(n1207), .Z(n1215) );
  XNOR U4269 ( .A(n1209), .B(n1215), .Z(n1210) );
  XOR U4270 ( .A(n1211), .B(n1210), .Z(z[45]) );
  XNOR U4271 ( .A(n1213), .B(n1212), .Z(z[46]) );
  XNOR U4272 ( .A(n1215), .B(n1214), .Z(n1216) );
  XNOR U4273 ( .A(z[41]), .B(n1216), .Z(z[47]) );
  IV U4274 ( .A(x[49]), .Z(n1324) );
  XOR U4275 ( .A(x[48]), .B(x[54]), .Z(n1218) );
  IV U4276 ( .A(n1323), .Z(n1219) );
  AND U4277 ( .A(n1324), .B(n1219), .Z(n1226) );
  XNOR U4278 ( .A(x[50]), .B(n1222), .Z(n1217) );
  XNOR U4279 ( .A(n1218), .B(n1217), .Z(n1282) );
  IV U4280 ( .A(n1282), .Z(n1228) );
  XNOR U4281 ( .A(n1228), .B(n1323), .Z(n1281) );
  IV U4282 ( .A(x[55]), .Z(n1220) );
  XNOR U4283 ( .A(x[49]), .B(n1220), .Z(n1314) );
  NAND U4284 ( .A(n1281), .B(n1314), .Z(n1231) );
  XNOR U4285 ( .A(n1220), .B(n1219), .Z(n1227) );
  IV U4286 ( .A(n1227), .Z(n1312) );
  XOR U4287 ( .A(n1282), .B(n1312), .Z(n1247) );
  XNOR U4288 ( .A(n1231), .B(n1247), .Z(n1224) );
  XOR U4289 ( .A(x[48]), .B(n1228), .Z(n1257) );
  XOR U4290 ( .A(x[52]), .B(n1220), .Z(n1221) );
  IV U4291 ( .A(n1221), .Z(n1286) );
  NANDN U4292 ( .A(n1257), .B(n1286), .Z(n1230) );
  XNOR U4293 ( .A(n1222), .B(n1221), .Z(n1275) );
  XNOR U4294 ( .A(n1281), .B(n1275), .Z(n1273) );
  XOR U4295 ( .A(x[50]), .B(x[52]), .Z(n1288) );
  NANDN U4296 ( .A(n1273), .B(n1288), .Z(n1223) );
  XOR U4297 ( .A(n1230), .B(n1223), .Z(n1249) );
  XNOR U4298 ( .A(n1224), .B(n1249), .Z(n1225) );
  XOR U4299 ( .A(n1226), .B(n1225), .Z(n1262) );
  IV U4300 ( .A(n1262), .Z(n1268) );
  AND U4301 ( .A(n1228), .B(n1227), .Z(n1233) );
  XOR U4302 ( .A(x[48]), .B(n1275), .Z(n1276) );
  XNOR U4303 ( .A(n1323), .B(n1276), .Z(n1278) );
  XOR U4304 ( .A(x[50]), .B(x[55]), .Z(n1303) );
  NANDN U4305 ( .A(n1278), .B(n1303), .Z(n1229) );
  XNOR U4306 ( .A(n1230), .B(n1229), .Z(n1238) );
  XNOR U4307 ( .A(n1231), .B(n1238), .Z(n1232) );
  XOR U4308 ( .A(n1233), .B(n1232), .Z(n1258) );
  XNOR U4309 ( .A(x[52]), .B(n1323), .Z(n1296) );
  ANDN U4310 ( .B(x[48]), .A(n1296), .Z(n1240) );
  XOR U4311 ( .A(x[50]), .B(x[49]), .Z(n1234) );
  XOR U4312 ( .A(n1312), .B(n1234), .Z(n1285) );
  XOR U4313 ( .A(n1286), .B(n1234), .Z(n1291) );
  NAND U4314 ( .A(n1275), .B(n1291), .Z(n1242) );
  XNOR U4315 ( .A(n1285), .B(n1242), .Z(n1236) );
  XNOR U4316 ( .A(x[49]), .B(n1276), .Z(n1235) );
  XNOR U4317 ( .A(n1236), .B(n1235), .Z(n1237) );
  XOR U4318 ( .A(n1238), .B(n1237), .Z(n1239) );
  XOR U4319 ( .A(n1240), .B(n1239), .Z(n1260) );
  NAND U4320 ( .A(n1258), .B(n1260), .Z(n1241) );
  NAND U4321 ( .A(n1268), .B(n1241), .Z(n1252) );
  IV U4322 ( .A(n1258), .Z(n1259) );
  IV U4323 ( .A(n1260), .Z(n1266) );
  XOR U4324 ( .A(n1242), .B(n1296), .Z(n1245) );
  AND U4325 ( .A(n1285), .B(n1276), .Z(n1243) );
  XNOR U4326 ( .A(x[48]), .B(n1243), .Z(n1244) );
  XNOR U4327 ( .A(n1245), .B(n1244), .Z(n1246) );
  XNOR U4328 ( .A(n1247), .B(n1246), .Z(n1248) );
  XNOR U4329 ( .A(n1249), .B(n1248), .Z(n1270) );
  IV U4330 ( .A(n1270), .Z(n1265) );
  XOR U4331 ( .A(n1266), .B(n1265), .Z(n1250) );
  NAND U4332 ( .A(n1259), .B(n1250), .Z(n1251) );
  AND U4333 ( .A(n1252), .B(n1251), .Z(n1331) );
  NAND U4334 ( .A(n1266), .B(n1259), .Z(n1253) );
  NAND U4335 ( .A(n1265), .B(n1253), .Z(n1256) );
  XOR U4336 ( .A(n1259), .B(n1262), .Z(n1254) );
  NAND U4337 ( .A(n1260), .B(n1254), .Z(n1255) );
  AND U4338 ( .A(n1256), .B(n1255), .Z(n1313) );
  XNOR U4339 ( .A(n1331), .B(n1313), .Z(n1287) );
  OR U4340 ( .A(n1287), .B(n1257), .Z(n1280) );
  NAND U4341 ( .A(n1268), .B(n1258), .Z(n1264) );
  AND U4342 ( .A(n1260), .B(n1259), .Z(n1267) );
  XNOR U4343 ( .A(n1265), .B(n1267), .Z(n1261) );
  NAND U4344 ( .A(n1262), .B(n1261), .Z(n1263) );
  AND U4345 ( .A(n1264), .B(n1263), .Z(n1284) );
  NAND U4346 ( .A(n1266), .B(n1265), .Z(n1272) );
  XNOR U4347 ( .A(n1268), .B(n1267), .Z(n1269) );
  NAND U4348 ( .A(n1270), .B(n1269), .Z(n1271) );
  NAND U4349 ( .A(n1272), .B(n1271), .Z(n1325) );
  XNOR U4350 ( .A(n1284), .B(n1325), .Z(n1302) );
  XOR U4351 ( .A(n1302), .B(n1287), .Z(n1289) );
  OR U4352 ( .A(n1289), .B(n1273), .Z(n1274) );
  XNOR U4353 ( .A(n1280), .B(n1274), .Z(n1306) );
  XOR U4354 ( .A(n1284), .B(n1331), .Z(n1292) );
  NANDN U4355 ( .A(n1292), .B(n1275), .Z(n1333) );
  NANDN U4356 ( .A(n1284), .B(n1276), .Z(n1277) );
  XNOR U4357 ( .A(n1333), .B(n1277), .Z(n1311) );
  XOR U4358 ( .A(n1306), .B(n1311), .Z(n1295) );
  NANDN U4359 ( .A(n1278), .B(n1302), .Z(n1279) );
  XNOR U4360 ( .A(n1280), .B(n1279), .Z(n1339) );
  XNOR U4361 ( .A(n1325), .B(n1313), .Z(n1315) );
  NANDN U4362 ( .A(n1315), .B(n1281), .Z(n1298) );
  NAND U4363 ( .A(n1282), .B(n1313), .Z(n1283) );
  XNOR U4364 ( .A(n1298), .B(n1283), .Z(n1330) );
  XOR U4365 ( .A(n1339), .B(n1330), .Z(n1322) );
  XNOR U4366 ( .A(n1295), .B(n1322), .Z(z[48]) );
  ANDN U4367 ( .B(n1285), .A(n1284), .Z(n1294) );
  NANDN U4368 ( .A(n1287), .B(n1286), .Z(n1305) );
  NANDN U4369 ( .A(n1289), .B(n1288), .Z(n1290) );
  XNOR U4370 ( .A(n1305), .B(n1290), .Z(n1334) );
  NANDN U4371 ( .A(n1292), .B(n1291), .Z(n1299) );
  XNOR U4372 ( .A(n1334), .B(n1299), .Z(n1293) );
  XOR U4373 ( .A(n1294), .B(n1293), .Z(n1320) );
  XOR U4374 ( .A(n1320), .B(n1295), .Z(n1338) );
  ANDN U4375 ( .B(n1331), .A(n1296), .Z(n1301) );
  NAND U4376 ( .A(n1323), .B(n1325), .Z(n1297) );
  XNOR U4377 ( .A(n1298), .B(n1297), .Z(n1310) );
  XNOR U4378 ( .A(n1299), .B(n1310), .Z(n1300) );
  XNOR U4379 ( .A(n1301), .B(n1300), .Z(n1308) );
  NAND U4380 ( .A(n1303), .B(n1302), .Z(n1304) );
  XNOR U4381 ( .A(n1305), .B(n1304), .Z(n1316) );
  XNOR U4382 ( .A(n1306), .B(n1316), .Z(n1307) );
  XOR U4383 ( .A(n1308), .B(n1307), .Z(n1319) );
  XNOR U4384 ( .A(n1338), .B(n1319), .Z(z[49]) );
  XOR U4385 ( .A(n1309), .B(z[2]), .Z(z[4]) );
  XNOR U4386 ( .A(n1311), .B(n1310), .Z(z[50]) );
  AND U4387 ( .A(n1313), .B(n1312), .Z(n1318) );
  NANDN U4388 ( .A(n1315), .B(n1314), .Z(n1328) );
  XNOR U4389 ( .A(n1316), .B(n1328), .Z(n1317) );
  XOR U4390 ( .A(n1318), .B(n1317), .Z(n1337) );
  XOR U4391 ( .A(n1320), .B(n1319), .Z(n1321) );
  XOR U4392 ( .A(n1337), .B(n1321), .Z(z[51]) );
  XOR U4393 ( .A(n1322), .B(z[50]), .Z(z[52]) );
  XNOR U4394 ( .A(n1324), .B(n1323), .Z(n1326) );
  NAND U4395 ( .A(n1326), .B(n1325), .Z(n1327) );
  XOR U4396 ( .A(n1328), .B(n1327), .Z(n1329) );
  XNOR U4397 ( .A(n1330), .B(n1329), .Z(n1336) );
  NAND U4398 ( .A(n1331), .B(x[48]), .Z(n1332) );
  XNOR U4399 ( .A(n1333), .B(n1332), .Z(n1340) );
  XNOR U4400 ( .A(n1334), .B(n1340), .Z(n1335) );
  XOR U4401 ( .A(n1336), .B(n1335), .Z(z[53]) );
  XNOR U4402 ( .A(n1338), .B(n1337), .Z(z[54]) );
  XNOR U4403 ( .A(n1340), .B(n1339), .Z(n1341) );
  XNOR U4404 ( .A(z[49]), .B(n1341), .Z(z[55]) );
  IV U4405 ( .A(x[57]), .Z(n1462) );
  XOR U4406 ( .A(x[56]), .B(x[62]), .Z(n1343) );
  XOR U4407 ( .A(x[61]), .B(n1343), .Z(n1461) );
  IV U4408 ( .A(n1461), .Z(n1344) );
  AND U4409 ( .A(n1462), .B(n1344), .Z(n1351) );
  XNOR U4410 ( .A(x[59]), .B(n1462), .Z(n1347) );
  XNOR U4411 ( .A(x[58]), .B(n1347), .Z(n1342) );
  XNOR U4412 ( .A(n1343), .B(n1342), .Z(n1407) );
  IV U4413 ( .A(n1407), .Z(n1353) );
  XNOR U4414 ( .A(n1353), .B(n1461), .Z(n1406) );
  IV U4415 ( .A(x[63]), .Z(n1345) );
  XNOR U4416 ( .A(x[57]), .B(n1345), .Z(n1438) );
  NAND U4417 ( .A(n1406), .B(n1438), .Z(n1356) );
  XNOR U4418 ( .A(n1345), .B(n1344), .Z(n1352) );
  IV U4419 ( .A(n1352), .Z(n1436) );
  XOR U4420 ( .A(n1407), .B(n1436), .Z(n1372) );
  XNOR U4421 ( .A(n1356), .B(n1372), .Z(n1349) );
  XOR U4422 ( .A(x[56]), .B(n1353), .Z(n1382) );
  XOR U4423 ( .A(x[60]), .B(n1345), .Z(n1346) );
  IV U4424 ( .A(n1346), .Z(n1411) );
  NANDN U4425 ( .A(n1382), .B(n1411), .Z(n1355) );
  XNOR U4426 ( .A(n1347), .B(n1346), .Z(n1400) );
  XNOR U4427 ( .A(n1406), .B(n1400), .Z(n1398) );
  XOR U4428 ( .A(x[58]), .B(x[60]), .Z(n1413) );
  NANDN U4429 ( .A(n1398), .B(n1413), .Z(n1348) );
  XOR U4430 ( .A(n1355), .B(n1348), .Z(n1374) );
  XNOR U4431 ( .A(n1349), .B(n1374), .Z(n1350) );
  XOR U4432 ( .A(n1351), .B(n1350), .Z(n1387) );
  IV U4433 ( .A(n1387), .Z(n1393) );
  AND U4434 ( .A(n1353), .B(n1352), .Z(n1358) );
  XOR U4435 ( .A(x[56]), .B(n1400), .Z(n1401) );
  XNOR U4436 ( .A(n1461), .B(n1401), .Z(n1403) );
  XOR U4437 ( .A(x[58]), .B(x[63]), .Z(n1428) );
  NANDN U4438 ( .A(n1403), .B(n1428), .Z(n1354) );
  XNOR U4439 ( .A(n1355), .B(n1354), .Z(n1363) );
  XNOR U4440 ( .A(n1356), .B(n1363), .Z(n1357) );
  XOR U4441 ( .A(n1358), .B(n1357), .Z(n1383) );
  XNOR U4442 ( .A(x[60]), .B(n1461), .Z(n1421) );
  ANDN U4443 ( .B(x[56]), .A(n1421), .Z(n1365) );
  XOR U4444 ( .A(x[58]), .B(x[57]), .Z(n1359) );
  XOR U4445 ( .A(n1436), .B(n1359), .Z(n1410) );
  XOR U4446 ( .A(n1411), .B(n1359), .Z(n1416) );
  NAND U4447 ( .A(n1400), .B(n1416), .Z(n1367) );
  XNOR U4448 ( .A(n1410), .B(n1367), .Z(n1361) );
  XNOR U4449 ( .A(x[57]), .B(n1401), .Z(n1360) );
  XNOR U4450 ( .A(n1361), .B(n1360), .Z(n1362) );
  XOR U4451 ( .A(n1363), .B(n1362), .Z(n1364) );
  XOR U4452 ( .A(n1365), .B(n1364), .Z(n1385) );
  NAND U4453 ( .A(n1383), .B(n1385), .Z(n1366) );
  NAND U4454 ( .A(n1393), .B(n1366), .Z(n1377) );
  IV U4455 ( .A(n1383), .Z(n1384) );
  IV U4456 ( .A(n1385), .Z(n1391) );
  XOR U4457 ( .A(n1367), .B(n1421), .Z(n1370) );
  AND U4458 ( .A(n1410), .B(n1401), .Z(n1368) );
  XNOR U4459 ( .A(x[56]), .B(n1368), .Z(n1369) );
  XNOR U4460 ( .A(n1370), .B(n1369), .Z(n1371) );
  XNOR U4461 ( .A(n1372), .B(n1371), .Z(n1373) );
  XNOR U4462 ( .A(n1374), .B(n1373), .Z(n1395) );
  IV U4463 ( .A(n1395), .Z(n1390) );
  XOR U4464 ( .A(n1391), .B(n1390), .Z(n1375) );
  NAND U4465 ( .A(n1384), .B(n1375), .Z(n1376) );
  AND U4466 ( .A(n1377), .B(n1376), .Z(n1469) );
  NAND U4467 ( .A(n1391), .B(n1384), .Z(n1378) );
  NAND U4468 ( .A(n1390), .B(n1378), .Z(n1381) );
  XOR U4469 ( .A(n1384), .B(n1387), .Z(n1379) );
  NAND U4470 ( .A(n1385), .B(n1379), .Z(n1380) );
  AND U4471 ( .A(n1381), .B(n1380), .Z(n1437) );
  XNOR U4472 ( .A(n1469), .B(n1437), .Z(n1412) );
  OR U4473 ( .A(n1412), .B(n1382), .Z(n1405) );
  NAND U4474 ( .A(n1393), .B(n1383), .Z(n1389) );
  AND U4475 ( .A(n1385), .B(n1384), .Z(n1392) );
  XNOR U4476 ( .A(n1390), .B(n1392), .Z(n1386) );
  NAND U4477 ( .A(n1387), .B(n1386), .Z(n1388) );
  AND U4478 ( .A(n1389), .B(n1388), .Z(n1409) );
  NAND U4479 ( .A(n1391), .B(n1390), .Z(n1397) );
  XNOR U4480 ( .A(n1393), .B(n1392), .Z(n1394) );
  NAND U4481 ( .A(n1395), .B(n1394), .Z(n1396) );
  NAND U4482 ( .A(n1397), .B(n1396), .Z(n1463) );
  XNOR U4483 ( .A(n1409), .B(n1463), .Z(n1427) );
  XOR U4484 ( .A(n1427), .B(n1412), .Z(n1414) );
  OR U4485 ( .A(n1414), .B(n1398), .Z(n1399) );
  XNOR U4486 ( .A(n1405), .B(n1399), .Z(n1431) );
  XOR U4487 ( .A(n1409), .B(n1469), .Z(n1417) );
  NANDN U4488 ( .A(n1417), .B(n1400), .Z(n1471) );
  NANDN U4489 ( .A(n1409), .B(n1401), .Z(n1402) );
  XNOR U4490 ( .A(n1471), .B(n1402), .Z(n1435) );
  XOR U4491 ( .A(n1431), .B(n1435), .Z(n1420) );
  NANDN U4492 ( .A(n1403), .B(n1427), .Z(n1404) );
  XNOR U4493 ( .A(n1405), .B(n1404), .Z(n1477) );
  XNOR U4494 ( .A(n1463), .B(n1437), .Z(n1439) );
  NANDN U4495 ( .A(n1439), .B(n1406), .Z(n1423) );
  NAND U4496 ( .A(n1407), .B(n1437), .Z(n1408) );
  XNOR U4497 ( .A(n1423), .B(n1408), .Z(n1468) );
  XOR U4498 ( .A(n1477), .B(n1468), .Z(n1460) );
  XNOR U4499 ( .A(n1420), .B(n1460), .Z(z[56]) );
  ANDN U4500 ( .B(n1410), .A(n1409), .Z(n1419) );
  NANDN U4501 ( .A(n1412), .B(n1411), .Z(n1430) );
  NANDN U4502 ( .A(n1414), .B(n1413), .Z(n1415) );
  XNOR U4503 ( .A(n1430), .B(n1415), .Z(n1472) );
  NANDN U4504 ( .A(n1417), .B(n1416), .Z(n1424) );
  XNOR U4505 ( .A(n1472), .B(n1424), .Z(n1418) );
  XOR U4506 ( .A(n1419), .B(n1418), .Z(n1444) );
  XOR U4507 ( .A(n1444), .B(n1420), .Z(n1476) );
  ANDN U4508 ( .B(n1469), .A(n1421), .Z(n1426) );
  NAND U4509 ( .A(n1461), .B(n1463), .Z(n1422) );
  XNOR U4510 ( .A(n1423), .B(n1422), .Z(n1434) );
  XNOR U4511 ( .A(n1424), .B(n1434), .Z(n1425) );
  XNOR U4512 ( .A(n1426), .B(n1425), .Z(n1433) );
  NAND U4513 ( .A(n1428), .B(n1427), .Z(n1429) );
  XNOR U4514 ( .A(n1430), .B(n1429), .Z(n1440) );
  XNOR U4515 ( .A(n1431), .B(n1440), .Z(n1432) );
  XOR U4516 ( .A(n1433), .B(n1432), .Z(n1443) );
  XNOR U4517 ( .A(n1476), .B(n1443), .Z(z[57]) );
  XNOR U4518 ( .A(n1435), .B(n1434), .Z(z[58]) );
  AND U4519 ( .A(n1437), .B(n1436), .Z(n1442) );
  NANDN U4520 ( .A(n1439), .B(n1438), .Z(n1466) );
  XNOR U4521 ( .A(n1440), .B(n1466), .Z(n1441) );
  XOR U4522 ( .A(n1442), .B(n1441), .Z(n1475) );
  XOR U4523 ( .A(n1444), .B(n1443), .Z(n1445) );
  XOR U4524 ( .A(n1475), .B(n1445), .Z(z[59]) );
  XNOR U4525 ( .A(n1447), .B(n1446), .Z(n1449) );
  NAND U4526 ( .A(n1449), .B(n1448), .Z(n1450) );
  XOR U4527 ( .A(n1451), .B(n1450), .Z(n1452) );
  XNOR U4528 ( .A(n1453), .B(n1452), .Z(n1459) );
  NAND U4529 ( .A(n1454), .B(x[0]), .Z(n1455) );
  XNOR U4530 ( .A(n1456), .B(n1455), .Z(n1731) );
  XNOR U4531 ( .A(n1457), .B(n1731), .Z(n1458) );
  XOR U4532 ( .A(n1459), .B(n1458), .Z(z[5]) );
  XOR U4533 ( .A(n1460), .B(z[58]), .Z(z[60]) );
  XNOR U4534 ( .A(n1462), .B(n1461), .Z(n1464) );
  NAND U4535 ( .A(n1464), .B(n1463), .Z(n1465) );
  XOR U4536 ( .A(n1466), .B(n1465), .Z(n1467) );
  XNOR U4537 ( .A(n1468), .B(n1467), .Z(n1474) );
  NAND U4538 ( .A(n1469), .B(x[56]), .Z(n1470) );
  XNOR U4539 ( .A(n1471), .B(n1470), .Z(n1478) );
  XNOR U4540 ( .A(n1472), .B(n1478), .Z(n1473) );
  XOR U4541 ( .A(n1474), .B(n1473), .Z(z[61]) );
  XNOR U4542 ( .A(n1476), .B(n1475), .Z(z[62]) );
  XNOR U4543 ( .A(n1478), .B(n1477), .Z(n1479) );
  XNOR U4544 ( .A(z[57]), .B(n1479), .Z(z[63]) );
  IV U4545 ( .A(x[65]), .Z(n1586) );
  XOR U4546 ( .A(x[64]), .B(x[70]), .Z(n1481) );
  XOR U4547 ( .A(x[69]), .B(n1481), .Z(n1585) );
  IV U4548 ( .A(n1585), .Z(n1482) );
  AND U4549 ( .A(n1586), .B(n1482), .Z(n1489) );
  XNOR U4550 ( .A(x[67]), .B(n1586), .Z(n1485) );
  XNOR U4551 ( .A(x[66]), .B(n1485), .Z(n1480) );
  XNOR U4552 ( .A(n1481), .B(n1480), .Z(n1545) );
  IV U4553 ( .A(n1545), .Z(n1491) );
  XNOR U4554 ( .A(n1491), .B(n1585), .Z(n1544) );
  IV U4555 ( .A(x[71]), .Z(n1483) );
  XNOR U4556 ( .A(x[65]), .B(n1483), .Z(n1576) );
  NAND U4557 ( .A(n1544), .B(n1576), .Z(n1494) );
  XNOR U4558 ( .A(n1483), .B(n1482), .Z(n1490) );
  IV U4559 ( .A(n1490), .Z(n1574) );
  XOR U4560 ( .A(n1545), .B(n1574), .Z(n1510) );
  XNOR U4561 ( .A(n1494), .B(n1510), .Z(n1487) );
  XOR U4562 ( .A(x[64]), .B(n1491), .Z(n1520) );
  XOR U4563 ( .A(x[68]), .B(n1483), .Z(n1484) );
  IV U4564 ( .A(n1484), .Z(n1549) );
  NANDN U4565 ( .A(n1520), .B(n1549), .Z(n1493) );
  XNOR U4566 ( .A(n1485), .B(n1484), .Z(n1538) );
  XNOR U4567 ( .A(n1544), .B(n1538), .Z(n1536) );
  XOR U4568 ( .A(x[66]), .B(x[68]), .Z(n1551) );
  NANDN U4569 ( .A(n1536), .B(n1551), .Z(n1486) );
  XOR U4570 ( .A(n1493), .B(n1486), .Z(n1512) );
  XNOR U4571 ( .A(n1487), .B(n1512), .Z(n1488) );
  XOR U4572 ( .A(n1489), .B(n1488), .Z(n1525) );
  IV U4573 ( .A(n1525), .Z(n1531) );
  AND U4574 ( .A(n1491), .B(n1490), .Z(n1496) );
  XOR U4575 ( .A(x[64]), .B(n1538), .Z(n1539) );
  XNOR U4576 ( .A(n1585), .B(n1539), .Z(n1541) );
  XOR U4577 ( .A(x[66]), .B(x[71]), .Z(n1566) );
  NANDN U4578 ( .A(n1541), .B(n1566), .Z(n1492) );
  XNOR U4579 ( .A(n1493), .B(n1492), .Z(n1501) );
  XNOR U4580 ( .A(n1494), .B(n1501), .Z(n1495) );
  XOR U4581 ( .A(n1496), .B(n1495), .Z(n1521) );
  XNOR U4582 ( .A(x[68]), .B(n1585), .Z(n1559) );
  ANDN U4583 ( .B(x[64]), .A(n1559), .Z(n1503) );
  XOR U4584 ( .A(x[66]), .B(x[65]), .Z(n1497) );
  XOR U4585 ( .A(n1574), .B(n1497), .Z(n1548) );
  XOR U4586 ( .A(n1549), .B(n1497), .Z(n1554) );
  NAND U4587 ( .A(n1538), .B(n1554), .Z(n1505) );
  XNOR U4588 ( .A(n1548), .B(n1505), .Z(n1499) );
  XNOR U4589 ( .A(x[65]), .B(n1539), .Z(n1498) );
  XNOR U4590 ( .A(n1499), .B(n1498), .Z(n1500) );
  XOR U4591 ( .A(n1501), .B(n1500), .Z(n1502) );
  XOR U4592 ( .A(n1503), .B(n1502), .Z(n1523) );
  NAND U4593 ( .A(n1521), .B(n1523), .Z(n1504) );
  NAND U4594 ( .A(n1531), .B(n1504), .Z(n1515) );
  IV U4595 ( .A(n1521), .Z(n1522) );
  IV U4596 ( .A(n1523), .Z(n1529) );
  XOR U4597 ( .A(n1505), .B(n1559), .Z(n1508) );
  AND U4598 ( .A(n1548), .B(n1539), .Z(n1506) );
  XNOR U4599 ( .A(x[64]), .B(n1506), .Z(n1507) );
  XNOR U4600 ( .A(n1508), .B(n1507), .Z(n1509) );
  XNOR U4601 ( .A(n1510), .B(n1509), .Z(n1511) );
  XNOR U4602 ( .A(n1512), .B(n1511), .Z(n1533) );
  IV U4603 ( .A(n1533), .Z(n1528) );
  XOR U4604 ( .A(n1529), .B(n1528), .Z(n1513) );
  NAND U4605 ( .A(n1522), .B(n1513), .Z(n1514) );
  AND U4606 ( .A(n1515), .B(n1514), .Z(n1593) );
  NAND U4607 ( .A(n1529), .B(n1522), .Z(n1516) );
  NAND U4608 ( .A(n1528), .B(n1516), .Z(n1519) );
  XOR U4609 ( .A(n1522), .B(n1525), .Z(n1517) );
  NAND U4610 ( .A(n1523), .B(n1517), .Z(n1518) );
  AND U4611 ( .A(n1519), .B(n1518), .Z(n1575) );
  XNOR U4612 ( .A(n1593), .B(n1575), .Z(n1550) );
  OR U4613 ( .A(n1550), .B(n1520), .Z(n1543) );
  NAND U4614 ( .A(n1531), .B(n1521), .Z(n1527) );
  AND U4615 ( .A(n1523), .B(n1522), .Z(n1530) );
  XNOR U4616 ( .A(n1528), .B(n1530), .Z(n1524) );
  NAND U4617 ( .A(n1525), .B(n1524), .Z(n1526) );
  AND U4618 ( .A(n1527), .B(n1526), .Z(n1547) );
  NAND U4619 ( .A(n1529), .B(n1528), .Z(n1535) );
  XNOR U4620 ( .A(n1531), .B(n1530), .Z(n1532) );
  NAND U4621 ( .A(n1533), .B(n1532), .Z(n1534) );
  NAND U4622 ( .A(n1535), .B(n1534), .Z(n1587) );
  XNOR U4623 ( .A(n1547), .B(n1587), .Z(n1565) );
  XOR U4624 ( .A(n1565), .B(n1550), .Z(n1552) );
  OR U4625 ( .A(n1552), .B(n1536), .Z(n1537) );
  XNOR U4626 ( .A(n1543), .B(n1537), .Z(n1569) );
  XOR U4627 ( .A(n1547), .B(n1593), .Z(n1555) );
  NANDN U4628 ( .A(n1555), .B(n1538), .Z(n1595) );
  NANDN U4629 ( .A(n1547), .B(n1539), .Z(n1540) );
  XNOR U4630 ( .A(n1595), .B(n1540), .Z(n1573) );
  XOR U4631 ( .A(n1569), .B(n1573), .Z(n1558) );
  NANDN U4632 ( .A(n1541), .B(n1565), .Z(n1542) );
  XNOR U4633 ( .A(n1543), .B(n1542), .Z(n1603) );
  XNOR U4634 ( .A(n1587), .B(n1575), .Z(n1577) );
  NANDN U4635 ( .A(n1577), .B(n1544), .Z(n1561) );
  NAND U4636 ( .A(n1545), .B(n1575), .Z(n1546) );
  XNOR U4637 ( .A(n1561), .B(n1546), .Z(n1592) );
  XOR U4638 ( .A(n1603), .B(n1592), .Z(n1584) );
  XNOR U4639 ( .A(n1558), .B(n1584), .Z(z[64]) );
  ANDN U4640 ( .B(n1548), .A(n1547), .Z(n1557) );
  NANDN U4641 ( .A(n1550), .B(n1549), .Z(n1568) );
  NANDN U4642 ( .A(n1552), .B(n1551), .Z(n1553) );
  XNOR U4643 ( .A(n1568), .B(n1553), .Z(n1596) );
  NANDN U4644 ( .A(n1555), .B(n1554), .Z(n1562) );
  XNOR U4645 ( .A(n1596), .B(n1562), .Z(n1556) );
  XOR U4646 ( .A(n1557), .B(n1556), .Z(n1582) );
  XOR U4647 ( .A(n1582), .B(n1558), .Z(n1602) );
  ANDN U4648 ( .B(n1593), .A(n1559), .Z(n1564) );
  NAND U4649 ( .A(n1585), .B(n1587), .Z(n1560) );
  XNOR U4650 ( .A(n1561), .B(n1560), .Z(n1572) );
  XNOR U4651 ( .A(n1562), .B(n1572), .Z(n1563) );
  XNOR U4652 ( .A(n1564), .B(n1563), .Z(n1571) );
  NAND U4653 ( .A(n1566), .B(n1565), .Z(n1567) );
  XNOR U4654 ( .A(n1568), .B(n1567), .Z(n1578) );
  XNOR U4655 ( .A(n1569), .B(n1578), .Z(n1570) );
  XOR U4656 ( .A(n1571), .B(n1570), .Z(n1581) );
  XNOR U4657 ( .A(n1602), .B(n1581), .Z(z[65]) );
  XNOR U4658 ( .A(n1573), .B(n1572), .Z(z[66]) );
  AND U4659 ( .A(n1575), .B(n1574), .Z(n1580) );
  NANDN U4660 ( .A(n1577), .B(n1576), .Z(n1590) );
  XNOR U4661 ( .A(n1578), .B(n1590), .Z(n1579) );
  XOR U4662 ( .A(n1580), .B(n1579), .Z(n1601) );
  XOR U4663 ( .A(n1582), .B(n1581), .Z(n1583) );
  XOR U4664 ( .A(n1601), .B(n1583), .Z(z[67]) );
  XOR U4665 ( .A(n1584), .B(z[66]), .Z(z[68]) );
  XNOR U4666 ( .A(n1586), .B(n1585), .Z(n1588) );
  NAND U4667 ( .A(n1588), .B(n1587), .Z(n1589) );
  XOR U4668 ( .A(n1590), .B(n1589), .Z(n1591) );
  XNOR U4669 ( .A(n1592), .B(n1591), .Z(n1598) );
  NAND U4670 ( .A(n1593), .B(x[64]), .Z(n1594) );
  XNOR U4671 ( .A(n1595), .B(n1594), .Z(n1604) );
  XNOR U4672 ( .A(n1596), .B(n1604), .Z(n1597) );
  XOR U4673 ( .A(n1598), .B(n1597), .Z(z[69]) );
  XNOR U4674 ( .A(n1600), .B(n1599), .Z(z[6]) );
  XNOR U4675 ( .A(n1602), .B(n1601), .Z(z[70]) );
  XNOR U4676 ( .A(n1604), .B(n1603), .Z(n1605) );
  XNOR U4677 ( .A(z[65]), .B(n1605), .Z(z[71]) );
  IV U4678 ( .A(x[73]), .Z(n1712) );
  XOR U4679 ( .A(x[72]), .B(x[78]), .Z(n1607) );
  XOR U4680 ( .A(x[77]), .B(n1607), .Z(n1711) );
  IV U4681 ( .A(n1711), .Z(n1608) );
  AND U4682 ( .A(n1712), .B(n1608), .Z(n1615) );
  XNOR U4683 ( .A(x[75]), .B(n1712), .Z(n1611) );
  XNOR U4684 ( .A(x[74]), .B(n1611), .Z(n1606) );
  XNOR U4685 ( .A(n1607), .B(n1606), .Z(n1671) );
  IV U4686 ( .A(n1671), .Z(n1617) );
  XNOR U4687 ( .A(n1617), .B(n1711), .Z(n1670) );
  IV U4688 ( .A(x[79]), .Z(n1609) );
  XNOR U4689 ( .A(x[73]), .B(n1609), .Z(n1702) );
  NAND U4690 ( .A(n1670), .B(n1702), .Z(n1620) );
  XNOR U4691 ( .A(n1609), .B(n1608), .Z(n1616) );
  IV U4692 ( .A(n1616), .Z(n1700) );
  XOR U4693 ( .A(n1671), .B(n1700), .Z(n1636) );
  XNOR U4694 ( .A(n1620), .B(n1636), .Z(n1613) );
  XOR U4695 ( .A(x[72]), .B(n1617), .Z(n1646) );
  XOR U4696 ( .A(x[76]), .B(n1609), .Z(n1610) );
  IV U4697 ( .A(n1610), .Z(n1675) );
  NANDN U4698 ( .A(n1646), .B(n1675), .Z(n1619) );
  XNOR U4699 ( .A(n1611), .B(n1610), .Z(n1664) );
  XNOR U4700 ( .A(n1670), .B(n1664), .Z(n1662) );
  XOR U4701 ( .A(x[74]), .B(x[76]), .Z(n1677) );
  NANDN U4702 ( .A(n1662), .B(n1677), .Z(n1612) );
  XOR U4703 ( .A(n1619), .B(n1612), .Z(n1638) );
  XNOR U4704 ( .A(n1613), .B(n1638), .Z(n1614) );
  XOR U4705 ( .A(n1615), .B(n1614), .Z(n1651) );
  IV U4706 ( .A(n1651), .Z(n1657) );
  AND U4707 ( .A(n1617), .B(n1616), .Z(n1622) );
  XOR U4708 ( .A(x[72]), .B(n1664), .Z(n1665) );
  XNOR U4709 ( .A(n1711), .B(n1665), .Z(n1667) );
  XOR U4710 ( .A(x[74]), .B(x[79]), .Z(n1692) );
  NANDN U4711 ( .A(n1667), .B(n1692), .Z(n1618) );
  XNOR U4712 ( .A(n1619), .B(n1618), .Z(n1627) );
  XNOR U4713 ( .A(n1620), .B(n1627), .Z(n1621) );
  XOR U4714 ( .A(n1622), .B(n1621), .Z(n1647) );
  XNOR U4715 ( .A(x[76]), .B(n1711), .Z(n1685) );
  ANDN U4716 ( .B(x[72]), .A(n1685), .Z(n1629) );
  XOR U4717 ( .A(x[74]), .B(x[73]), .Z(n1623) );
  XOR U4718 ( .A(n1700), .B(n1623), .Z(n1674) );
  XOR U4719 ( .A(n1675), .B(n1623), .Z(n1680) );
  NAND U4720 ( .A(n1664), .B(n1680), .Z(n1631) );
  XNOR U4721 ( .A(n1674), .B(n1631), .Z(n1625) );
  XNOR U4722 ( .A(x[73]), .B(n1665), .Z(n1624) );
  XNOR U4723 ( .A(n1625), .B(n1624), .Z(n1626) );
  XOR U4724 ( .A(n1627), .B(n1626), .Z(n1628) );
  XOR U4725 ( .A(n1629), .B(n1628), .Z(n1649) );
  NAND U4726 ( .A(n1647), .B(n1649), .Z(n1630) );
  NAND U4727 ( .A(n1657), .B(n1630), .Z(n1641) );
  IV U4728 ( .A(n1647), .Z(n1648) );
  IV U4729 ( .A(n1649), .Z(n1655) );
  XOR U4730 ( .A(n1631), .B(n1685), .Z(n1634) );
  AND U4731 ( .A(n1674), .B(n1665), .Z(n1632) );
  XNOR U4732 ( .A(x[72]), .B(n1632), .Z(n1633) );
  XNOR U4733 ( .A(n1634), .B(n1633), .Z(n1635) );
  XNOR U4734 ( .A(n1636), .B(n1635), .Z(n1637) );
  XNOR U4735 ( .A(n1638), .B(n1637), .Z(n1659) );
  IV U4736 ( .A(n1659), .Z(n1654) );
  XOR U4737 ( .A(n1655), .B(n1654), .Z(n1639) );
  NAND U4738 ( .A(n1648), .B(n1639), .Z(n1640) );
  AND U4739 ( .A(n1641), .B(n1640), .Z(n1719) );
  NAND U4740 ( .A(n1655), .B(n1648), .Z(n1642) );
  NAND U4741 ( .A(n1654), .B(n1642), .Z(n1645) );
  XOR U4742 ( .A(n1648), .B(n1651), .Z(n1643) );
  NAND U4743 ( .A(n1649), .B(n1643), .Z(n1644) );
  AND U4744 ( .A(n1645), .B(n1644), .Z(n1701) );
  XNOR U4745 ( .A(n1719), .B(n1701), .Z(n1676) );
  OR U4746 ( .A(n1676), .B(n1646), .Z(n1669) );
  NAND U4747 ( .A(n1657), .B(n1647), .Z(n1653) );
  AND U4748 ( .A(n1649), .B(n1648), .Z(n1656) );
  XNOR U4749 ( .A(n1654), .B(n1656), .Z(n1650) );
  NAND U4750 ( .A(n1651), .B(n1650), .Z(n1652) );
  AND U4751 ( .A(n1653), .B(n1652), .Z(n1673) );
  NAND U4752 ( .A(n1655), .B(n1654), .Z(n1661) );
  XNOR U4753 ( .A(n1657), .B(n1656), .Z(n1658) );
  NAND U4754 ( .A(n1659), .B(n1658), .Z(n1660) );
  NAND U4755 ( .A(n1661), .B(n1660), .Z(n1713) );
  XNOR U4756 ( .A(n1673), .B(n1713), .Z(n1691) );
  XOR U4757 ( .A(n1691), .B(n1676), .Z(n1678) );
  OR U4758 ( .A(n1678), .B(n1662), .Z(n1663) );
  XNOR U4759 ( .A(n1669), .B(n1663), .Z(n1695) );
  XOR U4760 ( .A(n1673), .B(n1719), .Z(n1681) );
  NANDN U4761 ( .A(n1681), .B(n1664), .Z(n1721) );
  NANDN U4762 ( .A(n1673), .B(n1665), .Z(n1666) );
  XNOR U4763 ( .A(n1721), .B(n1666), .Z(n1699) );
  XOR U4764 ( .A(n1695), .B(n1699), .Z(n1684) );
  NANDN U4765 ( .A(n1667), .B(n1691), .Z(n1668) );
  XNOR U4766 ( .A(n1669), .B(n1668), .Z(n1727) );
  XNOR U4767 ( .A(n1713), .B(n1701), .Z(n1703) );
  NANDN U4768 ( .A(n1703), .B(n1670), .Z(n1687) );
  NAND U4769 ( .A(n1671), .B(n1701), .Z(n1672) );
  XNOR U4770 ( .A(n1687), .B(n1672), .Z(n1718) );
  XOR U4771 ( .A(n1727), .B(n1718), .Z(n1710) );
  XNOR U4772 ( .A(n1684), .B(n1710), .Z(z[72]) );
  ANDN U4773 ( .B(n1674), .A(n1673), .Z(n1683) );
  NANDN U4774 ( .A(n1676), .B(n1675), .Z(n1694) );
  NANDN U4775 ( .A(n1678), .B(n1677), .Z(n1679) );
  XNOR U4776 ( .A(n1694), .B(n1679), .Z(n1722) );
  NANDN U4777 ( .A(n1681), .B(n1680), .Z(n1688) );
  XNOR U4778 ( .A(n1722), .B(n1688), .Z(n1682) );
  XOR U4779 ( .A(n1683), .B(n1682), .Z(n1708) );
  XOR U4780 ( .A(n1708), .B(n1684), .Z(n1726) );
  ANDN U4781 ( .B(n1719), .A(n1685), .Z(n1690) );
  NAND U4782 ( .A(n1711), .B(n1713), .Z(n1686) );
  XNOR U4783 ( .A(n1687), .B(n1686), .Z(n1698) );
  XNOR U4784 ( .A(n1688), .B(n1698), .Z(n1689) );
  XNOR U4785 ( .A(n1690), .B(n1689), .Z(n1697) );
  NAND U4786 ( .A(n1692), .B(n1691), .Z(n1693) );
  XNOR U4787 ( .A(n1694), .B(n1693), .Z(n1704) );
  XNOR U4788 ( .A(n1695), .B(n1704), .Z(n1696) );
  XOR U4789 ( .A(n1697), .B(n1696), .Z(n1707) );
  XNOR U4790 ( .A(n1726), .B(n1707), .Z(z[73]) );
  XNOR U4791 ( .A(n1699), .B(n1698), .Z(z[74]) );
  AND U4792 ( .A(n1701), .B(n1700), .Z(n1706) );
  NANDN U4793 ( .A(n1703), .B(n1702), .Z(n1716) );
  XNOR U4794 ( .A(n1704), .B(n1716), .Z(n1705) );
  XOR U4795 ( .A(n1706), .B(n1705), .Z(n1725) );
  XOR U4796 ( .A(n1708), .B(n1707), .Z(n1709) );
  XOR U4797 ( .A(n1725), .B(n1709), .Z(z[75]) );
  XOR U4798 ( .A(n1710), .B(z[74]), .Z(z[76]) );
  XNOR U4799 ( .A(n1712), .B(n1711), .Z(n1714) );
  NAND U4800 ( .A(n1714), .B(n1713), .Z(n1715) );
  XOR U4801 ( .A(n1716), .B(n1715), .Z(n1717) );
  XNOR U4802 ( .A(n1718), .B(n1717), .Z(n1724) );
  NAND U4803 ( .A(n1719), .B(x[72]), .Z(n1720) );
  XNOR U4804 ( .A(n1721), .B(n1720), .Z(n1728) );
  XNOR U4805 ( .A(n1722), .B(n1728), .Z(n1723) );
  XOR U4806 ( .A(n1724), .B(n1723), .Z(z[77]) );
  XNOR U4807 ( .A(n1726), .B(n1725), .Z(z[78]) );
  XNOR U4808 ( .A(n1728), .B(n1727), .Z(n1729) );
  XNOR U4809 ( .A(z[73]), .B(n1729), .Z(z[79]) );
  XNOR U4810 ( .A(n1731), .B(n1730), .Z(n1732) );
  XNOR U4811 ( .A(z[1]), .B(n1732), .Z(z[7]) );
  XOR U4812 ( .A(x[80]), .B(x[86]), .Z(n1733) );
  IV U4813 ( .A(n1838), .Z(n1735) );
  IV U4814 ( .A(x[81]), .Z(n1837) );
  NAND U4815 ( .A(n1735), .B(n1837), .Z(n1742) );
  XNOR U4816 ( .A(x[82]), .B(n1733), .Z(n1734) );
  XNOR U4817 ( .A(n1738), .B(n1734), .Z(n1797) );
  XNOR U4818 ( .A(n1735), .B(n1797), .Z(n1796) );
  IV U4819 ( .A(x[87]), .Z(n1736) );
  XNOR U4820 ( .A(x[81]), .B(n1736), .Z(n1828) );
  NAND U4821 ( .A(n1796), .B(n1828), .Z(n1745) );
  XNOR U4822 ( .A(n1735), .B(n1736), .Z(n1826) );
  XOR U4823 ( .A(n1797), .B(n1826), .Z(n1753) );
  XOR U4824 ( .A(n1745), .B(n1753), .Z(n1740) );
  XNOR U4825 ( .A(x[80]), .B(n1797), .Z(n1772) );
  XOR U4826 ( .A(x[84]), .B(n1736), .Z(n1737) );
  IV U4827 ( .A(n1737), .Z(n1801) );
  NANDN U4828 ( .A(n1772), .B(n1801), .Z(n1744) );
  XOR U4829 ( .A(n1738), .B(n1737), .Z(n1790) );
  XOR U4830 ( .A(n1796), .B(n1790), .Z(n1788) );
  XOR U4831 ( .A(x[82]), .B(x[84]), .Z(n1803) );
  NANDN U4832 ( .A(n1788), .B(n1803), .Z(n1739) );
  XNOR U4833 ( .A(n1744), .B(n1739), .Z(n1749) );
  XOR U4834 ( .A(n1740), .B(n1749), .Z(n1741) );
  XOR U4835 ( .A(n1742), .B(n1741), .Z(n1783) );
  IV U4836 ( .A(n1783), .Z(n1777) );
  ANDN U4837 ( .B(n1826), .A(n1797), .Z(n1747) );
  XNOR U4838 ( .A(x[80]), .B(n1790), .Z(n1791) );
  XNOR U4839 ( .A(n1838), .B(n1791), .Z(n1793) );
  XOR U4840 ( .A(x[82]), .B(x[87]), .Z(n1818) );
  NANDN U4841 ( .A(n1793), .B(n1818), .Z(n1743) );
  XNOR U4842 ( .A(n1744), .B(n1743), .Z(n1760) );
  XNOR U4843 ( .A(n1745), .B(n1760), .Z(n1746) );
  XOR U4844 ( .A(n1747), .B(n1746), .Z(n1773) );
  NAND U4845 ( .A(n1777), .B(n1773), .Z(n1767) );
  IV U4846 ( .A(n1773), .Z(n1774) );
  XOR U4847 ( .A(n1783), .B(n1774), .Z(n1765) );
  XOR U4848 ( .A(x[82]), .B(x[81]), .Z(n1748) );
  XNOR U4849 ( .A(n1826), .B(n1748), .Z(n1800) );
  NAND U4850 ( .A(n1800), .B(n1791), .Z(n1755) );
  XNOR U4851 ( .A(x[84]), .B(n1838), .Z(n1811) );
  XOR U4852 ( .A(n1801), .B(n1748), .Z(n1806) );
  NANDN U4853 ( .A(n1790), .B(n1806), .Z(n1756) );
  XOR U4854 ( .A(n1811), .B(n1756), .Z(n1751) );
  XOR U4855 ( .A(x[80]), .B(n1749), .Z(n1750) );
  XNOR U4856 ( .A(n1751), .B(n1750), .Z(n1752) );
  XOR U4857 ( .A(n1753), .B(n1752), .Z(n1754) );
  XOR U4858 ( .A(n1755), .B(n1754), .Z(n1785) );
  IV U4859 ( .A(n1785), .Z(n1780) );
  AND U4860 ( .A(n1777), .B(n1780), .Z(n1763) );
  ANDN U4861 ( .B(x[80]), .A(n1811), .Z(n1762) );
  XNOR U4862 ( .A(n1800), .B(n1756), .Z(n1758) );
  XNOR U4863 ( .A(x[81]), .B(n1791), .Z(n1757) );
  XNOR U4864 ( .A(n1758), .B(n1757), .Z(n1759) );
  XOR U4865 ( .A(n1760), .B(n1759), .Z(n1761) );
  XOR U4866 ( .A(n1762), .B(n1761), .Z(n1775) );
  IV U4867 ( .A(n1775), .Z(n1781) );
  XNOR U4868 ( .A(n1763), .B(n1781), .Z(n1764) );
  NAND U4869 ( .A(n1765), .B(n1764), .Z(n1766) );
  NAND U4870 ( .A(n1767), .B(n1766), .Z(n1845) );
  NAND U4871 ( .A(n1781), .B(n1774), .Z(n1768) );
  NAND U4872 ( .A(n1780), .B(n1768), .Z(n1771) );
  XOR U4873 ( .A(n1774), .B(n1777), .Z(n1769) );
  NAND U4874 ( .A(n1775), .B(n1769), .Z(n1770) );
  AND U4875 ( .A(n1771), .B(n1770), .Z(n1827) );
  XNOR U4876 ( .A(n1845), .B(n1827), .Z(n1802) );
  OR U4877 ( .A(n1802), .B(n1772), .Z(n1795) );
  NAND U4878 ( .A(n1783), .B(n1773), .Z(n1779) );
  AND U4879 ( .A(n1775), .B(n1774), .Z(n1782) );
  XNOR U4880 ( .A(n1782), .B(n1780), .Z(n1776) );
  NAND U4881 ( .A(n1777), .B(n1776), .Z(n1778) );
  AND U4882 ( .A(n1779), .B(n1778), .Z(n1799) );
  NAND U4883 ( .A(n1781), .B(n1780), .Z(n1787) );
  XNOR U4884 ( .A(n1783), .B(n1782), .Z(n1784) );
  NAND U4885 ( .A(n1785), .B(n1784), .Z(n1786) );
  NAND U4886 ( .A(n1787), .B(n1786), .Z(n1839) );
  XNOR U4887 ( .A(n1799), .B(n1839), .Z(n1817) );
  XOR U4888 ( .A(n1817), .B(n1802), .Z(n1804) );
  OR U4889 ( .A(n1804), .B(n1788), .Z(n1789) );
  XNOR U4890 ( .A(n1795), .B(n1789), .Z(n1821) );
  XOR U4891 ( .A(n1799), .B(n1845), .Z(n1807) );
  OR U4892 ( .A(n1790), .B(n1807), .Z(n1847) );
  NANDN U4893 ( .A(n1799), .B(n1791), .Z(n1792) );
  XNOR U4894 ( .A(n1847), .B(n1792), .Z(n1825) );
  XOR U4895 ( .A(n1821), .B(n1825), .Z(n1810) );
  NANDN U4896 ( .A(n1793), .B(n1817), .Z(n1794) );
  XNOR U4897 ( .A(n1795), .B(n1794), .Z(n1853) );
  XNOR U4898 ( .A(n1839), .B(n1827), .Z(n1829) );
  NANDN U4899 ( .A(n1829), .B(n1796), .Z(n1813) );
  NAND U4900 ( .A(n1797), .B(n1827), .Z(n1798) );
  XNOR U4901 ( .A(n1813), .B(n1798), .Z(n1844) );
  XOR U4902 ( .A(n1853), .B(n1844), .Z(n1836) );
  XNOR U4903 ( .A(n1810), .B(n1836), .Z(z[80]) );
  ANDN U4904 ( .B(n1800), .A(n1799), .Z(n1809) );
  NANDN U4905 ( .A(n1802), .B(n1801), .Z(n1820) );
  NANDN U4906 ( .A(n1804), .B(n1803), .Z(n1805) );
  XNOR U4907 ( .A(n1820), .B(n1805), .Z(n1848) );
  NANDN U4908 ( .A(n1807), .B(n1806), .Z(n1814) );
  XNOR U4909 ( .A(n1848), .B(n1814), .Z(n1808) );
  XOR U4910 ( .A(n1809), .B(n1808), .Z(n1834) );
  XOR U4911 ( .A(n1834), .B(n1810), .Z(n1852) );
  ANDN U4912 ( .B(n1845), .A(n1811), .Z(n1816) );
  NAND U4913 ( .A(n1838), .B(n1839), .Z(n1812) );
  XNOR U4914 ( .A(n1813), .B(n1812), .Z(n1824) );
  XNOR U4915 ( .A(n1814), .B(n1824), .Z(n1815) );
  XNOR U4916 ( .A(n1816), .B(n1815), .Z(n1823) );
  NAND U4917 ( .A(n1818), .B(n1817), .Z(n1819) );
  XNOR U4918 ( .A(n1820), .B(n1819), .Z(n1830) );
  XNOR U4919 ( .A(n1821), .B(n1830), .Z(n1822) );
  XOR U4920 ( .A(n1823), .B(n1822), .Z(n1833) );
  XNOR U4921 ( .A(n1852), .B(n1833), .Z(z[81]) );
  XNOR U4922 ( .A(n1825), .B(n1824), .Z(z[82]) );
  ANDN U4923 ( .B(n1827), .A(n1826), .Z(n1832) );
  NANDN U4924 ( .A(n1829), .B(n1828), .Z(n1842) );
  XNOR U4925 ( .A(n1830), .B(n1842), .Z(n1831) );
  XOR U4926 ( .A(n1832), .B(n1831), .Z(n1851) );
  XOR U4927 ( .A(n1834), .B(n1833), .Z(n1835) );
  XOR U4928 ( .A(n1851), .B(n1835), .Z(z[83]) );
  XOR U4929 ( .A(n1836), .B(z[82]), .Z(z[84]) );
  XNOR U4930 ( .A(n1838), .B(n1837), .Z(n1840) );
  NAND U4931 ( .A(n1840), .B(n1839), .Z(n1841) );
  XOR U4932 ( .A(n1842), .B(n1841), .Z(n1843) );
  XNOR U4933 ( .A(n1844), .B(n1843), .Z(n1850) );
  NAND U4934 ( .A(x[80]), .B(n1845), .Z(n1846) );
  XNOR U4935 ( .A(n1847), .B(n1846), .Z(n1854) );
  XNOR U4936 ( .A(n1848), .B(n1854), .Z(n1849) );
  XOR U4937 ( .A(n1850), .B(n1849), .Z(z[85]) );
  XNOR U4938 ( .A(n1852), .B(n1851), .Z(z[86]) );
  XNOR U4939 ( .A(n1854), .B(n1853), .Z(n1855) );
  XNOR U4940 ( .A(z[81]), .B(n1855), .Z(z[87]) );
  XOR U4941 ( .A(x[88]), .B(x[94]), .Z(n1856) );
  XOR U4942 ( .A(x[93]), .B(n1856), .Z(n1963) );
  IV U4943 ( .A(n1963), .Z(n1858) );
  IV U4944 ( .A(x[89]), .Z(n1962) );
  NAND U4945 ( .A(n1858), .B(n1962), .Z(n1865) );
  XOR U4946 ( .A(x[91]), .B(x[89]), .Z(n1861) );
  XNOR U4947 ( .A(x[90]), .B(n1856), .Z(n1857) );
  XNOR U4948 ( .A(n1861), .B(n1857), .Z(n1920) );
  XNOR U4949 ( .A(n1858), .B(n1920), .Z(n1919) );
  IV U4950 ( .A(x[95]), .Z(n1859) );
  XNOR U4951 ( .A(x[89]), .B(n1859), .Z(n1953) );
  NAND U4952 ( .A(n1919), .B(n1953), .Z(n1868) );
  XNOR U4953 ( .A(n1858), .B(n1859), .Z(n1951) );
  XOR U4954 ( .A(n1920), .B(n1951), .Z(n1876) );
  XOR U4955 ( .A(n1868), .B(n1876), .Z(n1863) );
  XNOR U4956 ( .A(x[88]), .B(n1920), .Z(n1895) );
  XOR U4957 ( .A(x[92]), .B(n1859), .Z(n1860) );
  IV U4958 ( .A(n1860), .Z(n1924) );
  NANDN U4959 ( .A(n1895), .B(n1924), .Z(n1867) );
  XOR U4960 ( .A(n1861), .B(n1860), .Z(n1913) );
  XOR U4961 ( .A(n1919), .B(n1913), .Z(n1911) );
  XOR U4962 ( .A(x[90]), .B(x[92]), .Z(n1926) );
  NANDN U4963 ( .A(n1911), .B(n1926), .Z(n1862) );
  XNOR U4964 ( .A(n1867), .B(n1862), .Z(n1872) );
  XOR U4965 ( .A(n1863), .B(n1872), .Z(n1864) );
  XOR U4966 ( .A(n1865), .B(n1864), .Z(n1906) );
  IV U4967 ( .A(n1906), .Z(n1900) );
  ANDN U4968 ( .B(n1951), .A(n1920), .Z(n1870) );
  XNOR U4969 ( .A(x[88]), .B(n1913), .Z(n1914) );
  XNOR U4970 ( .A(n1963), .B(n1914), .Z(n1916) );
  XOR U4971 ( .A(x[90]), .B(x[95]), .Z(n1941) );
  NANDN U4972 ( .A(n1916), .B(n1941), .Z(n1866) );
  XNOR U4973 ( .A(n1867), .B(n1866), .Z(n1883) );
  XNOR U4974 ( .A(n1868), .B(n1883), .Z(n1869) );
  XOR U4975 ( .A(n1870), .B(n1869), .Z(n1896) );
  NAND U4976 ( .A(n1900), .B(n1896), .Z(n1890) );
  IV U4977 ( .A(n1896), .Z(n1897) );
  XOR U4978 ( .A(n1906), .B(n1897), .Z(n1888) );
  XOR U4979 ( .A(x[90]), .B(x[89]), .Z(n1871) );
  XNOR U4980 ( .A(n1951), .B(n1871), .Z(n1923) );
  NAND U4981 ( .A(n1923), .B(n1914), .Z(n1878) );
  XNOR U4982 ( .A(x[92]), .B(n1963), .Z(n1934) );
  XOR U4983 ( .A(n1924), .B(n1871), .Z(n1929) );
  NANDN U4984 ( .A(n1913), .B(n1929), .Z(n1879) );
  XOR U4985 ( .A(n1934), .B(n1879), .Z(n1874) );
  XOR U4986 ( .A(x[88]), .B(n1872), .Z(n1873) );
  XNOR U4987 ( .A(n1874), .B(n1873), .Z(n1875) );
  XOR U4988 ( .A(n1876), .B(n1875), .Z(n1877) );
  XOR U4989 ( .A(n1878), .B(n1877), .Z(n1908) );
  IV U4990 ( .A(n1908), .Z(n1903) );
  AND U4991 ( .A(n1900), .B(n1903), .Z(n1886) );
  ANDN U4992 ( .B(x[88]), .A(n1934), .Z(n1885) );
  XNOR U4993 ( .A(n1923), .B(n1879), .Z(n1881) );
  XNOR U4994 ( .A(x[89]), .B(n1914), .Z(n1880) );
  XNOR U4995 ( .A(n1881), .B(n1880), .Z(n1882) );
  XOR U4996 ( .A(n1883), .B(n1882), .Z(n1884) );
  XOR U4997 ( .A(n1885), .B(n1884), .Z(n1898) );
  IV U4998 ( .A(n1898), .Z(n1904) );
  XNOR U4999 ( .A(n1886), .B(n1904), .Z(n1887) );
  NAND U5000 ( .A(n1888), .B(n1887), .Z(n1889) );
  NAND U5001 ( .A(n1890), .B(n1889), .Z(n1970) );
  NAND U5002 ( .A(n1904), .B(n1897), .Z(n1891) );
  NAND U5003 ( .A(n1903), .B(n1891), .Z(n1894) );
  XOR U5004 ( .A(n1897), .B(n1900), .Z(n1892) );
  NAND U5005 ( .A(n1898), .B(n1892), .Z(n1893) );
  AND U5006 ( .A(n1894), .B(n1893), .Z(n1952) );
  XNOR U5007 ( .A(n1970), .B(n1952), .Z(n1925) );
  OR U5008 ( .A(n1925), .B(n1895), .Z(n1918) );
  NAND U5009 ( .A(n1906), .B(n1896), .Z(n1902) );
  AND U5010 ( .A(n1898), .B(n1897), .Z(n1905) );
  XNOR U5011 ( .A(n1905), .B(n1903), .Z(n1899) );
  NAND U5012 ( .A(n1900), .B(n1899), .Z(n1901) );
  AND U5013 ( .A(n1902), .B(n1901), .Z(n1922) );
  NAND U5014 ( .A(n1904), .B(n1903), .Z(n1910) );
  XNOR U5015 ( .A(n1906), .B(n1905), .Z(n1907) );
  NAND U5016 ( .A(n1908), .B(n1907), .Z(n1909) );
  NAND U5017 ( .A(n1910), .B(n1909), .Z(n1964) );
  XNOR U5018 ( .A(n1922), .B(n1964), .Z(n1940) );
  XOR U5019 ( .A(n1940), .B(n1925), .Z(n1927) );
  OR U5020 ( .A(n1927), .B(n1911), .Z(n1912) );
  XNOR U5021 ( .A(n1918), .B(n1912), .Z(n1944) );
  XOR U5022 ( .A(n1922), .B(n1970), .Z(n1930) );
  OR U5023 ( .A(n1913), .B(n1930), .Z(n1972) );
  NANDN U5024 ( .A(n1922), .B(n1914), .Z(n1915) );
  XNOR U5025 ( .A(n1972), .B(n1915), .Z(n1950) );
  XOR U5026 ( .A(n1944), .B(n1950), .Z(n1933) );
  NANDN U5027 ( .A(n1916), .B(n1940), .Z(n1917) );
  XNOR U5028 ( .A(n1918), .B(n1917), .Z(n1978) );
  XNOR U5029 ( .A(n1964), .B(n1952), .Z(n1954) );
  NANDN U5030 ( .A(n1954), .B(n1919), .Z(n1936) );
  NAND U5031 ( .A(n1920), .B(n1952), .Z(n1921) );
  XNOR U5032 ( .A(n1936), .B(n1921), .Z(n1969) );
  XOR U5033 ( .A(n1978), .B(n1969), .Z(n1961) );
  XNOR U5034 ( .A(n1933), .B(n1961), .Z(z[88]) );
  ANDN U5035 ( .B(n1923), .A(n1922), .Z(n1932) );
  NANDN U5036 ( .A(n1925), .B(n1924), .Z(n1943) );
  NANDN U5037 ( .A(n1927), .B(n1926), .Z(n1928) );
  XNOR U5038 ( .A(n1943), .B(n1928), .Z(n1973) );
  NANDN U5039 ( .A(n1930), .B(n1929), .Z(n1937) );
  XNOR U5040 ( .A(n1973), .B(n1937), .Z(n1931) );
  XOR U5041 ( .A(n1932), .B(n1931), .Z(n1959) );
  XOR U5042 ( .A(n1959), .B(n1933), .Z(n1977) );
  ANDN U5043 ( .B(n1970), .A(n1934), .Z(n1939) );
  NAND U5044 ( .A(n1963), .B(n1964), .Z(n1935) );
  XNOR U5045 ( .A(n1936), .B(n1935), .Z(n1949) );
  XNOR U5046 ( .A(n1937), .B(n1949), .Z(n1938) );
  XNOR U5047 ( .A(n1939), .B(n1938), .Z(n1946) );
  NAND U5048 ( .A(n1941), .B(n1940), .Z(n1942) );
  XNOR U5049 ( .A(n1943), .B(n1942), .Z(n1955) );
  XNOR U5050 ( .A(n1944), .B(n1955), .Z(n1945) );
  XOR U5051 ( .A(n1946), .B(n1945), .Z(n1958) );
  XNOR U5052 ( .A(n1977), .B(n1958), .Z(z[89]) );
  XNOR U5053 ( .A(n1948), .B(n1947), .Z(z[8]) );
  XNOR U5054 ( .A(n1950), .B(n1949), .Z(z[90]) );
  ANDN U5055 ( .B(n1952), .A(n1951), .Z(n1957) );
  NANDN U5056 ( .A(n1954), .B(n1953), .Z(n1967) );
  XNOR U5057 ( .A(n1955), .B(n1967), .Z(n1956) );
  XOR U5058 ( .A(n1957), .B(n1956), .Z(n1976) );
  XOR U5059 ( .A(n1959), .B(n1958), .Z(n1960) );
  XOR U5060 ( .A(n1976), .B(n1960), .Z(z[91]) );
  XOR U5061 ( .A(n1961), .B(z[90]), .Z(z[92]) );
  XNOR U5062 ( .A(n1963), .B(n1962), .Z(n1965) );
  NAND U5063 ( .A(n1965), .B(n1964), .Z(n1966) );
  XOR U5064 ( .A(n1967), .B(n1966), .Z(n1968) );
  XNOR U5065 ( .A(n1969), .B(n1968), .Z(n1975) );
  NAND U5066 ( .A(x[88]), .B(n1970), .Z(n1971) );
  XNOR U5067 ( .A(n1972), .B(n1971), .Z(n1979) );
  XNOR U5068 ( .A(n1973), .B(n1979), .Z(n1974) );
  XOR U5069 ( .A(n1975), .B(n1974), .Z(z[93]) );
  XNOR U5070 ( .A(n1977), .B(n1976), .Z(z[94]) );
  XNOR U5071 ( .A(n1979), .B(n1978), .Z(n1980) );
  XNOR U5072 ( .A(z[89]), .B(n1980), .Z(z[95]) );
  XNOR U5073 ( .A(n1982), .B(n1981), .Z(z[96]) );
  XOR U5074 ( .A(n1984), .B(n1983), .Z(n1985) );
  XOR U5075 ( .A(n1986), .B(n1985), .Z(z[99]) );
endmodule


module SubBytes_5 ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986;

  XOR U2962 ( .A(x[21]), .B(n685), .Z(n814) );
  XOR U2963 ( .A(x[53]), .B(n1218), .Z(n1323) );
  XNOR U2964 ( .A(n328), .B(n339), .Z(n341) );
  XNOR U2965 ( .A(n1324), .B(x[51]), .Z(n1222) );
  XOR U2966 ( .A(x[81]), .B(x[83]), .Z(n1738) );
  XNOR U2967 ( .A(n170), .B(n162), .Z(n143) );
  XOR U2968 ( .A(x[16]), .B(x[22]), .Z(n685) );
  XOR U2969 ( .A(n493), .B(n494), .Z(n646) );
  XOR U2970 ( .A(x[85]), .B(n1733), .Z(n1838) );
  IV U2971 ( .A(x[1]), .Z(n1447) );
  XOR U2972 ( .A(x[0]), .B(x[6]), .Z(n2) );
  XOR U2973 ( .A(x[5]), .B(n2), .Z(n1446) );
  IV U2974 ( .A(n1446), .Z(n3) );
  AND U2975 ( .A(n1447), .B(n3), .Z(n10) );
  XNOR U2976 ( .A(x[3]), .B(n1447), .Z(n6) );
  XNOR U2977 ( .A(x[2]), .B(n6), .Z(n1) );
  XNOR U2978 ( .A(n2), .B(n1), .Z(n66) );
  IV U2979 ( .A(n66), .Z(n12) );
  XNOR U2980 ( .A(n12), .B(n1446), .Z(n65) );
  IV U2981 ( .A(x[7]), .Z(n4) );
  XNOR U2982 ( .A(x[1]), .B(n4), .Z(n1085) );
  NAND U2983 ( .A(n65), .B(n1085), .Z(n15) );
  XNOR U2984 ( .A(n4), .B(n3), .Z(n11) );
  IV U2985 ( .A(n11), .Z(n1083) );
  XOR U2986 ( .A(n66), .B(n1083), .Z(n31) );
  XNOR U2987 ( .A(n15), .B(n31), .Z(n8) );
  XOR U2988 ( .A(x[0]), .B(n12), .Z(n41) );
  XOR U2989 ( .A(x[4]), .B(n4), .Z(n5) );
  IV U2990 ( .A(n5), .Z(n790) );
  NANDN U2991 ( .A(n41), .B(n790), .Z(n14) );
  XNOR U2992 ( .A(n6), .B(n5), .Z(n59) );
  XNOR U2993 ( .A(n65), .B(n59), .Z(n57) );
  XOR U2994 ( .A(x[2]), .B(x[4]), .Z(n792) );
  NANDN U2995 ( .A(n57), .B(n792), .Z(n7) );
  XOR U2996 ( .A(n14), .B(n7), .Z(n33) );
  XNOR U2997 ( .A(n8), .B(n33), .Z(n9) );
  XOR U2998 ( .A(n10), .B(n9), .Z(n46) );
  IV U2999 ( .A(n46), .Z(n52) );
  AND U3000 ( .A(n12), .B(n11), .Z(n17) );
  XOR U3001 ( .A(x[0]), .B(n59), .Z(n60) );
  XNOR U3002 ( .A(n1446), .B(n60), .Z(n62) );
  XOR U3003 ( .A(x[2]), .B(x[7]), .Z(n807) );
  NANDN U3004 ( .A(n62), .B(n807), .Z(n13) );
  XNOR U3005 ( .A(n14), .B(n13), .Z(n22) );
  XNOR U3006 ( .A(n15), .B(n22), .Z(n16) );
  XOR U3007 ( .A(n17), .B(n16), .Z(n42) );
  XNOR U3008 ( .A(x[4]), .B(n1446), .Z(n800) );
  ANDN U3009 ( .B(x[0]), .A(n800), .Z(n24) );
  XOR U3010 ( .A(x[2]), .B(x[1]), .Z(n18) );
  XOR U3011 ( .A(n1083), .B(n18), .Z(n789) );
  XOR U3012 ( .A(n790), .B(n18), .Z(n795) );
  NAND U3013 ( .A(n59), .B(n795), .Z(n26) );
  XNOR U3014 ( .A(n789), .B(n26), .Z(n20) );
  XNOR U3015 ( .A(x[1]), .B(n60), .Z(n19) );
  XNOR U3016 ( .A(n20), .B(n19), .Z(n21) );
  XOR U3017 ( .A(n22), .B(n21), .Z(n23) );
  XOR U3018 ( .A(n24), .B(n23), .Z(n44) );
  NAND U3019 ( .A(n42), .B(n44), .Z(n25) );
  NAND U3020 ( .A(n52), .B(n25), .Z(n36) );
  IV U3021 ( .A(n42), .Z(n43) );
  IV U3022 ( .A(n44), .Z(n50) );
  XOR U3023 ( .A(n26), .B(n800), .Z(n29) );
  AND U3024 ( .A(n789), .B(n60), .Z(n27) );
  XNOR U3025 ( .A(x[0]), .B(n27), .Z(n28) );
  XNOR U3026 ( .A(n29), .B(n28), .Z(n30) );
  XNOR U3027 ( .A(n31), .B(n30), .Z(n32) );
  XNOR U3028 ( .A(n33), .B(n32), .Z(n54) );
  IV U3029 ( .A(n54), .Z(n49) );
  XOR U3030 ( .A(n50), .B(n49), .Z(n34) );
  NAND U3031 ( .A(n43), .B(n34), .Z(n35) );
  AND U3032 ( .A(n36), .B(n35), .Z(n1454) );
  NAND U3033 ( .A(n50), .B(n43), .Z(n37) );
  NAND U3034 ( .A(n49), .B(n37), .Z(n40) );
  XOR U3035 ( .A(n43), .B(n46), .Z(n38) );
  NAND U3036 ( .A(n44), .B(n38), .Z(n39) );
  AND U3037 ( .A(n40), .B(n39), .Z(n1084) );
  XNOR U3038 ( .A(n1454), .B(n1084), .Z(n791) );
  OR U3039 ( .A(n791), .B(n41), .Z(n64) );
  NAND U3040 ( .A(n52), .B(n42), .Z(n48) );
  AND U3041 ( .A(n44), .B(n43), .Z(n51) );
  XNOR U3042 ( .A(n49), .B(n51), .Z(n45) );
  NAND U3043 ( .A(n46), .B(n45), .Z(n47) );
  AND U3044 ( .A(n48), .B(n47), .Z(n788) );
  NAND U3045 ( .A(n50), .B(n49), .Z(n56) );
  XNOR U3046 ( .A(n52), .B(n51), .Z(n53) );
  NAND U3047 ( .A(n54), .B(n53), .Z(n55) );
  NAND U3048 ( .A(n56), .B(n55), .Z(n1448) );
  XNOR U3049 ( .A(n788), .B(n1448), .Z(n806) );
  XOR U3050 ( .A(n806), .B(n791), .Z(n793) );
  OR U3051 ( .A(n793), .B(n57), .Z(n58) );
  XNOR U3052 ( .A(n64), .B(n58), .Z(n810) );
  XOR U3053 ( .A(n788), .B(n1454), .Z(n796) );
  NANDN U3054 ( .A(n796), .B(n59), .Z(n1456) );
  NANDN U3055 ( .A(n788), .B(n60), .Z(n61) );
  XNOR U3056 ( .A(n1456), .B(n61), .Z(n953) );
  XOR U3057 ( .A(n810), .B(n953), .Z(n799) );
  NANDN U3058 ( .A(n62), .B(n806), .Z(n63) );
  XNOR U3059 ( .A(n64), .B(n63), .Z(n1730) );
  XNOR U3060 ( .A(n1448), .B(n1084), .Z(n1086) );
  NANDN U3061 ( .A(n1086), .B(n65), .Z(n802) );
  NAND U3062 ( .A(n66), .B(n1084), .Z(n67) );
  XNOR U3063 ( .A(n802), .B(n67), .Z(n1453) );
  XOR U3064 ( .A(n1730), .B(n1453), .Z(n1309) );
  XNOR U3065 ( .A(n799), .B(n1309), .Z(z[0]) );
  XOR U3066 ( .A(x[96]), .B(x[102]), .Z(n68) );
  XOR U3067 ( .A(x[101]), .B(n68), .Z(n135) );
  XOR U3068 ( .A(x[100]), .B(n135), .Z(n171) );
  AND U3069 ( .A(x[96]), .B(n171), .Z(n78) );
  XOR U3070 ( .A(x[97]), .B(x[99]), .Z(n71) );
  XNOR U3071 ( .A(n68), .B(x[98]), .Z(n69) );
  XOR U3072 ( .A(n71), .B(n69), .Z(n129) );
  XOR U3073 ( .A(x[96]), .B(n129), .Z(n128) );
  XNOR U3074 ( .A(x[103]), .B(x[100]), .Z(n70) );
  IV U3075 ( .A(n70), .Z(n142) );
  NANDN U3076 ( .A(n128), .B(n142), .Z(n80) );
  IV U3077 ( .A(n135), .Z(n91) );
  XNOR U3078 ( .A(n71), .B(n70), .Z(n123) );
  XOR U3079 ( .A(x[96]), .B(n123), .Z(n124) );
  XOR U3080 ( .A(n91), .B(n124), .Z(n126) );
  XOR U3081 ( .A(x[98]), .B(x[103]), .Z(n164) );
  NANDN U3082 ( .A(n126), .B(n164), .Z(n72) );
  XNOR U3083 ( .A(n80), .B(n72), .Z(n87) );
  XNOR U3084 ( .A(n135), .B(x[103]), .Z(n161) );
  XOR U3085 ( .A(x[97]), .B(x[98]), .Z(n73) );
  XNOR U3086 ( .A(n161), .B(n73), .Z(n151) );
  XOR U3087 ( .A(n142), .B(n73), .Z(n152) );
  NAND U3088 ( .A(n123), .B(n152), .Z(n81) );
  XNOR U3089 ( .A(n151), .B(n81), .Z(n75) );
  XNOR U3090 ( .A(x[97]), .B(n124), .Z(n74) );
  XNOR U3091 ( .A(n75), .B(n74), .Z(n76) );
  XOR U3092 ( .A(n87), .B(n76), .Z(n77) );
  XOR U3093 ( .A(n78), .B(n77), .Z(n115) );
  IV U3094 ( .A(n115), .Z(n108) );
  XNOR U3095 ( .A(n129), .B(n135), .Z(n105) );
  XNOR U3096 ( .A(n105), .B(n123), .Z(n158) );
  XNOR U3097 ( .A(x[98]), .B(x[100]), .Z(n144) );
  OR U3098 ( .A(n158), .B(n144), .Z(n79) );
  XOR U3099 ( .A(n80), .B(n79), .Z(n94) );
  XNOR U3100 ( .A(n129), .B(n161), .Z(n92) );
  XNOR U3101 ( .A(n81), .B(n171), .Z(n84) );
  AND U3102 ( .A(n151), .B(n124), .Z(n82) );
  XNOR U3103 ( .A(x[96]), .B(n82), .Z(n83) );
  XNOR U3104 ( .A(n84), .B(n83), .Z(n85) );
  XOR U3105 ( .A(n92), .B(n85), .Z(n86) );
  XOR U3106 ( .A(n94), .B(n86), .Z(n118) );
  AND U3107 ( .A(n129), .B(n161), .Z(n89) );
  IV U3108 ( .A(x[97]), .Z(n136) );
  XNOR U3109 ( .A(n136), .B(x[103]), .Z(n133) );
  NAND U3110 ( .A(n105), .B(n133), .Z(n93) );
  XNOR U3111 ( .A(n93), .B(n87), .Z(n88) );
  XOR U3112 ( .A(n89), .B(n88), .Z(n107) );
  NAND U3113 ( .A(n118), .B(n107), .Z(n90) );
  NAND U3114 ( .A(n108), .B(n90), .Z(n99) );
  IV U3115 ( .A(n118), .Z(n102) );
  NAND U3116 ( .A(n91), .B(n136), .Z(n97) );
  XOR U3117 ( .A(n93), .B(n92), .Z(n95) );
  XNOR U3118 ( .A(n95), .B(n94), .Z(n96) );
  XOR U3119 ( .A(n97), .B(n96), .Z(n114) );
  IV U3120 ( .A(n107), .Z(n116) );
  XOR U3121 ( .A(n114), .B(n116), .Z(n111) );
  NAND U3122 ( .A(n102), .B(n111), .Z(n98) );
  AND U3123 ( .A(n99), .B(n98), .Z(n127) );
  NAND U3124 ( .A(n118), .B(n108), .Z(n104) );
  AND U3125 ( .A(n115), .B(n116), .Z(n100) );
  XNOR U3126 ( .A(n114), .B(n100), .Z(n101) );
  NAND U3127 ( .A(n102), .B(n101), .Z(n103) );
  AND U3128 ( .A(n104), .B(n103), .Z(n138) );
  XNOR U3129 ( .A(n127), .B(n138), .Z(n134) );
  NANDN U3130 ( .A(n134), .B(n105), .Z(n131) );
  NANDN U3131 ( .A(n138), .B(n135), .Z(n106) );
  XNOR U3132 ( .A(n131), .B(n106), .Z(n173) );
  IV U3133 ( .A(n114), .Z(n120) );
  NAND U3134 ( .A(n120), .B(n107), .Z(n113) );
  AND U3135 ( .A(n120), .B(n118), .Z(n109) );
  XNOR U3136 ( .A(n109), .B(n108), .Z(n110) );
  NAND U3137 ( .A(n111), .B(n110), .Z(n112) );
  NAND U3138 ( .A(n113), .B(n112), .Z(n170) );
  NAND U3139 ( .A(n114), .B(n116), .Z(n122) );
  NAND U3140 ( .A(n116), .B(n115), .Z(n117) );
  XNOR U3141 ( .A(n118), .B(n117), .Z(n119) );
  NAND U3142 ( .A(n120), .B(n119), .Z(n121) );
  NAND U3143 ( .A(n122), .B(n121), .Z(n150) );
  XOR U3144 ( .A(n170), .B(n150), .Z(n153) );
  NANDN U3145 ( .A(n153), .B(n123), .Z(n147) );
  NANDN U3146 ( .A(n150), .B(n124), .Z(n125) );
  XNOR U3147 ( .A(n147), .B(n125), .Z(n160) );
  XNOR U3148 ( .A(n173), .B(n160), .Z(z[98]) );
  XOR U3149 ( .A(n150), .B(n138), .Z(n163) );
  ANDN U3150 ( .B(n163), .A(n126), .Z(n184) );
  IV U3151 ( .A(n127), .Z(n162) );
  OR U3152 ( .A(n143), .B(n128), .Z(n182) );
  NANDN U3153 ( .A(n129), .B(n162), .Z(n130) );
  XNOR U3154 ( .A(n131), .B(n130), .Z(n141) );
  XNOR U3155 ( .A(n182), .B(n141), .Z(n132) );
  XOR U3156 ( .A(n184), .B(n132), .Z(n1982) );
  XNOR U3157 ( .A(n1982), .B(z[98]), .Z(z[100]) );
  NANDN U3158 ( .A(n134), .B(n133), .Z(n167) );
  XNOR U3159 ( .A(n136), .B(n135), .Z(n137) );
  NANDN U3160 ( .A(n138), .B(n137), .Z(n139) );
  XOR U3161 ( .A(n167), .B(n139), .Z(n140) );
  XNOR U3162 ( .A(n141), .B(n140), .Z(n149) );
  NANDN U3163 ( .A(n143), .B(n142), .Z(n166) );
  XNOR U3164 ( .A(n143), .B(n163), .Z(n157) );
  NANDN U3165 ( .A(n144), .B(n157), .Z(n145) );
  XNOR U3166 ( .A(n166), .B(n145), .Z(n154) );
  NAND U3167 ( .A(n170), .B(x[96]), .Z(n146) );
  XNOR U3168 ( .A(n147), .B(n146), .Z(n181) );
  XNOR U3169 ( .A(n154), .B(n181), .Z(n148) );
  XOR U3170 ( .A(n149), .B(n148), .Z(z[101]) );
  ANDN U3171 ( .B(n151), .A(n150), .Z(n156) );
  NANDN U3172 ( .A(n153), .B(n152), .Z(n172) );
  XNOR U3173 ( .A(n172), .B(n154), .Z(n155) );
  XOR U3174 ( .A(n156), .B(n155), .Z(n1983) );
  NANDN U3175 ( .A(n158), .B(n157), .Z(n159) );
  XOR U3176 ( .A(n182), .B(n159), .Z(n176) );
  XOR U3177 ( .A(n176), .B(n160), .Z(n1981) );
  XNOR U3178 ( .A(n1983), .B(n1981), .Z(n180) );
  ANDN U3179 ( .B(n162), .A(n161), .Z(n169) );
  NAND U3180 ( .A(n164), .B(n163), .Z(n165) );
  XNOR U3181 ( .A(n166), .B(n165), .Z(n177) );
  XNOR U3182 ( .A(n177), .B(n167), .Z(n168) );
  XOR U3183 ( .A(n169), .B(n168), .Z(n1986) );
  XNOR U3184 ( .A(n180), .B(n1986), .Z(z[102]) );
  AND U3185 ( .A(n171), .B(n170), .Z(n175) );
  XNOR U3186 ( .A(n173), .B(n172), .Z(n174) );
  XNOR U3187 ( .A(n175), .B(n174), .Z(n179) );
  XOR U3188 ( .A(n177), .B(n176), .Z(n178) );
  XOR U3189 ( .A(n179), .B(n178), .Z(n1984) );
  XNOR U3190 ( .A(n1984), .B(n180), .Z(z[97]) );
  XNOR U3191 ( .A(n182), .B(n181), .Z(n183) );
  XNOR U3192 ( .A(n184), .B(n183), .Z(n185) );
  XOR U3193 ( .A(n185), .B(z[97]), .Z(z[103]) );
  IV U3194 ( .A(x[105]), .Z(n292) );
  XOR U3195 ( .A(x[104]), .B(x[110]), .Z(n187) );
  XOR U3196 ( .A(x[109]), .B(n187), .Z(n291) );
  IV U3197 ( .A(n291), .Z(n188) );
  AND U3198 ( .A(n292), .B(n188), .Z(n195) );
  XNOR U3199 ( .A(x[107]), .B(n292), .Z(n191) );
  XNOR U3200 ( .A(x[106]), .B(n191), .Z(n186) );
  XNOR U3201 ( .A(n187), .B(n186), .Z(n251) );
  IV U3202 ( .A(n251), .Z(n197) );
  XNOR U3203 ( .A(n197), .B(n291), .Z(n250) );
  IV U3204 ( .A(x[111]), .Z(n189) );
  XNOR U3205 ( .A(x[105]), .B(n189), .Z(n282) );
  NAND U3206 ( .A(n250), .B(n282), .Z(n200) );
  XNOR U3207 ( .A(n189), .B(n188), .Z(n196) );
  IV U3208 ( .A(n196), .Z(n280) );
  XOR U3209 ( .A(n251), .B(n280), .Z(n216) );
  XNOR U3210 ( .A(n200), .B(n216), .Z(n193) );
  XOR U3211 ( .A(x[104]), .B(n197), .Z(n226) );
  XOR U3212 ( .A(x[108]), .B(n189), .Z(n190) );
  IV U3213 ( .A(n190), .Z(n255) );
  NANDN U3214 ( .A(n226), .B(n255), .Z(n199) );
  XNOR U3215 ( .A(n191), .B(n190), .Z(n244) );
  XNOR U3216 ( .A(n250), .B(n244), .Z(n242) );
  XOR U3217 ( .A(x[106]), .B(x[108]), .Z(n257) );
  NANDN U3218 ( .A(n242), .B(n257), .Z(n192) );
  XOR U3219 ( .A(n199), .B(n192), .Z(n218) );
  XNOR U3220 ( .A(n193), .B(n218), .Z(n194) );
  XOR U3221 ( .A(n195), .B(n194), .Z(n231) );
  IV U3222 ( .A(n231), .Z(n237) );
  AND U3223 ( .A(n197), .B(n196), .Z(n202) );
  XOR U3224 ( .A(x[104]), .B(n244), .Z(n245) );
  XNOR U3225 ( .A(n291), .B(n245), .Z(n247) );
  XOR U3226 ( .A(x[106]), .B(x[111]), .Z(n272) );
  NANDN U3227 ( .A(n247), .B(n272), .Z(n198) );
  XNOR U3228 ( .A(n199), .B(n198), .Z(n207) );
  XNOR U3229 ( .A(n200), .B(n207), .Z(n201) );
  XOR U3230 ( .A(n202), .B(n201), .Z(n227) );
  XNOR U3231 ( .A(x[108]), .B(n291), .Z(n265) );
  ANDN U3232 ( .B(x[104]), .A(n265), .Z(n209) );
  XOR U3233 ( .A(x[106]), .B(x[105]), .Z(n203) );
  XOR U3234 ( .A(n280), .B(n203), .Z(n254) );
  XOR U3235 ( .A(n255), .B(n203), .Z(n260) );
  NAND U3236 ( .A(n244), .B(n260), .Z(n211) );
  XNOR U3237 ( .A(n254), .B(n211), .Z(n205) );
  XNOR U3238 ( .A(x[105]), .B(n245), .Z(n204) );
  XNOR U3239 ( .A(n205), .B(n204), .Z(n206) );
  XOR U3240 ( .A(n207), .B(n206), .Z(n208) );
  XOR U3241 ( .A(n209), .B(n208), .Z(n229) );
  NAND U3242 ( .A(n227), .B(n229), .Z(n210) );
  NAND U3243 ( .A(n237), .B(n210), .Z(n221) );
  IV U3244 ( .A(n227), .Z(n228) );
  IV U3245 ( .A(n229), .Z(n235) );
  XOR U3246 ( .A(n211), .B(n265), .Z(n214) );
  AND U3247 ( .A(n254), .B(n245), .Z(n212) );
  XNOR U3248 ( .A(x[104]), .B(n212), .Z(n213) );
  XNOR U3249 ( .A(n214), .B(n213), .Z(n215) );
  XNOR U3250 ( .A(n216), .B(n215), .Z(n217) );
  XNOR U3251 ( .A(n218), .B(n217), .Z(n239) );
  IV U3252 ( .A(n239), .Z(n234) );
  XOR U3253 ( .A(n235), .B(n234), .Z(n219) );
  NAND U3254 ( .A(n228), .B(n219), .Z(n220) );
  AND U3255 ( .A(n221), .B(n220), .Z(n299) );
  NAND U3256 ( .A(n235), .B(n228), .Z(n222) );
  NAND U3257 ( .A(n234), .B(n222), .Z(n225) );
  XOR U3258 ( .A(n228), .B(n231), .Z(n223) );
  NAND U3259 ( .A(n229), .B(n223), .Z(n224) );
  AND U3260 ( .A(n225), .B(n224), .Z(n281) );
  XNOR U3261 ( .A(n299), .B(n281), .Z(n256) );
  OR U3262 ( .A(n256), .B(n226), .Z(n249) );
  NAND U3263 ( .A(n237), .B(n227), .Z(n233) );
  AND U3264 ( .A(n229), .B(n228), .Z(n236) );
  XNOR U3265 ( .A(n234), .B(n236), .Z(n230) );
  NAND U3266 ( .A(n231), .B(n230), .Z(n232) );
  AND U3267 ( .A(n233), .B(n232), .Z(n253) );
  NAND U3268 ( .A(n235), .B(n234), .Z(n241) );
  XNOR U3269 ( .A(n237), .B(n236), .Z(n238) );
  NAND U3270 ( .A(n239), .B(n238), .Z(n240) );
  NAND U3271 ( .A(n241), .B(n240), .Z(n293) );
  XNOR U3272 ( .A(n253), .B(n293), .Z(n271) );
  XOR U3273 ( .A(n271), .B(n256), .Z(n258) );
  OR U3274 ( .A(n258), .B(n242), .Z(n243) );
  XNOR U3275 ( .A(n249), .B(n243), .Z(n275) );
  XOR U3276 ( .A(n253), .B(n299), .Z(n261) );
  NANDN U3277 ( .A(n261), .B(n244), .Z(n301) );
  NANDN U3278 ( .A(n253), .B(n245), .Z(n246) );
  XNOR U3279 ( .A(n301), .B(n246), .Z(n279) );
  XOR U3280 ( .A(n275), .B(n279), .Z(n264) );
  NANDN U3281 ( .A(n247), .B(n271), .Z(n248) );
  XNOR U3282 ( .A(n249), .B(n248), .Z(n366) );
  XNOR U3283 ( .A(n293), .B(n281), .Z(n283) );
  NANDN U3284 ( .A(n283), .B(n250), .Z(n267) );
  NAND U3285 ( .A(n251), .B(n281), .Z(n252) );
  XNOR U3286 ( .A(n267), .B(n252), .Z(n298) );
  XOR U3287 ( .A(n366), .B(n298), .Z(n290) );
  XNOR U3288 ( .A(n264), .B(n290), .Z(z[104]) );
  ANDN U3289 ( .B(n254), .A(n253), .Z(n263) );
  NANDN U3290 ( .A(n256), .B(n255), .Z(n274) );
  NANDN U3291 ( .A(n258), .B(n257), .Z(n259) );
  XNOR U3292 ( .A(n274), .B(n259), .Z(n302) );
  NANDN U3293 ( .A(n261), .B(n260), .Z(n268) );
  XNOR U3294 ( .A(n302), .B(n268), .Z(n262) );
  XOR U3295 ( .A(n263), .B(n262), .Z(n288) );
  XOR U3296 ( .A(n288), .B(n264), .Z(n365) );
  ANDN U3297 ( .B(n299), .A(n265), .Z(n270) );
  NAND U3298 ( .A(n291), .B(n293), .Z(n266) );
  XNOR U3299 ( .A(n267), .B(n266), .Z(n278) );
  XNOR U3300 ( .A(n268), .B(n278), .Z(n269) );
  XNOR U3301 ( .A(n270), .B(n269), .Z(n277) );
  NAND U3302 ( .A(n272), .B(n271), .Z(n273) );
  XNOR U3303 ( .A(n274), .B(n273), .Z(n284) );
  XNOR U3304 ( .A(n275), .B(n284), .Z(n276) );
  XOR U3305 ( .A(n277), .B(n276), .Z(n287) );
  XNOR U3306 ( .A(n365), .B(n287), .Z(z[105]) );
  XNOR U3307 ( .A(n279), .B(n278), .Z(z[106]) );
  AND U3308 ( .A(n281), .B(n280), .Z(n286) );
  NANDN U3309 ( .A(n283), .B(n282), .Z(n296) );
  XNOR U3310 ( .A(n284), .B(n296), .Z(n285) );
  XOR U3311 ( .A(n286), .B(n285), .Z(n364) );
  XOR U3312 ( .A(n288), .B(n287), .Z(n289) );
  XOR U3313 ( .A(n364), .B(n289), .Z(z[107]) );
  XOR U3314 ( .A(n290), .B(z[106]), .Z(z[108]) );
  XNOR U3315 ( .A(n292), .B(n291), .Z(n294) );
  NAND U3316 ( .A(n294), .B(n293), .Z(n295) );
  XOR U3317 ( .A(n296), .B(n295), .Z(n297) );
  XNOR U3318 ( .A(n298), .B(n297), .Z(n304) );
  NAND U3319 ( .A(n299), .B(x[104]), .Z(n300) );
  XNOR U3320 ( .A(n301), .B(n300), .Z(n367) );
  XNOR U3321 ( .A(n302), .B(n367), .Z(n303) );
  XOR U3322 ( .A(n304), .B(n303), .Z(z[109]) );
  IV U3323 ( .A(x[15]), .Z(n311) );
  IV U3324 ( .A(x[10]), .Z(n315) );
  XOR U3325 ( .A(x[11]), .B(x[9]), .Z(n307) );
  XOR U3326 ( .A(n315), .B(n307), .Z(n352) );
  IV U3327 ( .A(n352), .Z(n309) );
  XOR U3328 ( .A(x[13]), .B(n309), .Z(n305) );
  IV U3329 ( .A(x[9]), .Z(n655) );
  XNOR U3330 ( .A(n311), .B(n655), .Z(n515) );
  NAND U3331 ( .A(n305), .B(n515), .Z(n306) );
  XNOR U3332 ( .A(n311), .B(n306), .Z(n339) );
  XOR U3333 ( .A(x[12]), .B(n311), .Z(n314) );
  XNOR U3334 ( .A(x[14]), .B(n309), .Z(n497) );
  NOR U3335 ( .A(n314), .B(n497), .Z(n318) );
  IV U3336 ( .A(x[13]), .Z(n353) );
  XOR U3337 ( .A(x[8]), .B(x[14]), .Z(n310) );
  XOR U3338 ( .A(n353), .B(n310), .Z(n325) );
  IV U3339 ( .A(n325), .Z(n656) );
  XOR U3340 ( .A(n314), .B(n307), .Z(n316) );
  XNOR U3341 ( .A(x[8]), .B(n316), .Z(n350) );
  XNOR U3342 ( .A(n656), .B(n350), .Z(n648) );
  XNOR U3343 ( .A(x[15]), .B(n315), .Z(n673) );
  NANDN U3344 ( .A(n648), .B(n673), .Z(n308) );
  XOR U3345 ( .A(n318), .B(n308), .Z(n333) );
  XOR U3346 ( .A(n310), .B(n309), .Z(n313) );
  XNOR U3347 ( .A(n325), .B(n311), .Z(n516) );
  ANDN U3348 ( .B(n313), .A(n516), .Z(n312) );
  XOR U3349 ( .A(n333), .B(n312), .Z(n328) );
  IV U3350 ( .A(n313), .Z(n647) );
  IV U3351 ( .A(n314), .Z(n507) );
  XNOR U3352 ( .A(n655), .B(n315), .Z(n321) );
  XOR U3353 ( .A(n507), .B(n321), .Z(n501) );
  IV U3354 ( .A(n316), .Z(n344) );
  NANDN U3355 ( .A(n501), .B(n344), .Z(n329) );
  XNOR U3356 ( .A(x[12]), .B(x[10]), .Z(n508) );
  XNOR U3357 ( .A(n648), .B(n497), .Z(n498) );
  OR U3358 ( .A(n508), .B(n498), .Z(n317) );
  XOR U3359 ( .A(n318), .B(n317), .Z(n327) );
  XOR U3360 ( .A(n329), .B(n327), .Z(n320) );
  XNOR U3361 ( .A(x[8]), .B(n507), .Z(n319) );
  XNOR U3362 ( .A(n320), .B(n319), .Z(n323) );
  XOR U3363 ( .A(n321), .B(n516), .Z(n505) );
  NAND U3364 ( .A(n350), .B(n505), .Z(n322) );
  XNOR U3365 ( .A(n323), .B(n322), .Z(n324) );
  XOR U3366 ( .A(n647), .B(n324), .Z(n356) );
  IV U3367 ( .A(n356), .Z(n359) );
  NAND U3368 ( .A(n325), .B(n655), .Z(n326) );
  XOR U3369 ( .A(n327), .B(n326), .Z(n338) );
  XNOR U3370 ( .A(n328), .B(n338), .Z(n348) );
  NAND U3371 ( .A(n359), .B(n348), .Z(n337) );
  XOR U3372 ( .A(n656), .B(x[12]), .Z(n502) );
  AND U3373 ( .A(n502), .B(x[8]), .Z(n335) );
  XNOR U3374 ( .A(n505), .B(n329), .Z(n331) );
  XNOR U3375 ( .A(x[9]), .B(n350), .Z(n330) );
  XNOR U3376 ( .A(n331), .B(n330), .Z(n332) );
  XOR U3377 ( .A(n333), .B(n332), .Z(n334) );
  XNOR U3378 ( .A(n335), .B(n334), .Z(n358) );
  NANDN U3379 ( .A(n348), .B(n358), .Z(n336) );
  AND U3380 ( .A(n337), .B(n336), .Z(n342) );
  XNOR U3381 ( .A(n339), .B(n338), .Z(n345) );
  NANDN U3382 ( .A(n345), .B(n356), .Z(n340) );
  XNOR U3383 ( .A(n342), .B(n340), .Z(n354) );
  OR U3384 ( .A(n341), .B(n354), .Z(n495) );
  NANDN U3385 ( .A(n358), .B(n341), .Z(n347) );
  XOR U3386 ( .A(n345), .B(n342), .Z(n343) );
  XNOR U3387 ( .A(n347), .B(n343), .Z(n355) );
  NOR U3388 ( .A(n355), .B(n345), .Z(n349) );
  XOR U3389 ( .A(n495), .B(n349), .Z(n500) );
  NANDN U3390 ( .A(n500), .B(n344), .Z(n664) );
  ANDN U3391 ( .B(n359), .A(n345), .Z(n346) );
  XNOR U3392 ( .A(n347), .B(n346), .Z(n361) );
  OR U3393 ( .A(n361), .B(n348), .Z(n496) );
  XNOR U3394 ( .A(n496), .B(n349), .Z(n504) );
  AND U3395 ( .A(n504), .B(n350), .Z(n351) );
  XOR U3396 ( .A(n664), .B(n351), .Z(n670) );
  XOR U3397 ( .A(n353), .B(n352), .Z(n357) );
  ANDN U3398 ( .B(n358), .A(n354), .Z(n493) );
  NOR U3399 ( .A(n356), .B(n355), .Z(n362) );
  XOR U3400 ( .A(n493), .B(n362), .Z(n514) );
  NAND U3401 ( .A(n357), .B(n514), .Z(n651) );
  XOR U3402 ( .A(n359), .B(n358), .Z(n360) );
  NANDN U3403 ( .A(n361), .B(n360), .Z(n494) );
  XOR U3404 ( .A(n494), .B(n362), .Z(n658) );
  NANDN U3405 ( .A(n658), .B(n656), .Z(n363) );
  XNOR U3406 ( .A(n651), .B(n363), .Z(n519) );
  XOR U3407 ( .A(n670), .B(n519), .Z(n654) );
  IV U3408 ( .A(n654), .Z(z[10]) );
  XNOR U3409 ( .A(n365), .B(n364), .Z(z[110]) );
  XNOR U3410 ( .A(n367), .B(n366), .Z(n368) );
  XNOR U3411 ( .A(z[105]), .B(n368), .Z(z[111]) );
  IV U3412 ( .A(x[113]), .Z(n475) );
  XOR U3413 ( .A(x[112]), .B(x[118]), .Z(n370) );
  XOR U3414 ( .A(x[117]), .B(n370), .Z(n474) );
  IV U3415 ( .A(n474), .Z(n371) );
  AND U3416 ( .A(n475), .B(n371), .Z(n378) );
  XNOR U3417 ( .A(x[115]), .B(n475), .Z(n374) );
  XNOR U3418 ( .A(x[114]), .B(n374), .Z(n369) );
  XNOR U3419 ( .A(n370), .B(n369), .Z(n434) );
  IV U3420 ( .A(n434), .Z(n380) );
  XNOR U3421 ( .A(n380), .B(n474), .Z(n433) );
  IV U3422 ( .A(x[119]), .Z(n372) );
  XNOR U3423 ( .A(x[113]), .B(n372), .Z(n465) );
  NAND U3424 ( .A(n433), .B(n465), .Z(n383) );
  XNOR U3425 ( .A(n372), .B(n371), .Z(n379) );
  IV U3426 ( .A(n379), .Z(n463) );
  XOR U3427 ( .A(n434), .B(n463), .Z(n399) );
  XNOR U3428 ( .A(n383), .B(n399), .Z(n376) );
  XOR U3429 ( .A(x[112]), .B(n380), .Z(n409) );
  XOR U3430 ( .A(x[116]), .B(n372), .Z(n373) );
  IV U3431 ( .A(n373), .Z(n438) );
  NANDN U3432 ( .A(n409), .B(n438), .Z(n382) );
  XNOR U3433 ( .A(n374), .B(n373), .Z(n427) );
  XNOR U3434 ( .A(n433), .B(n427), .Z(n425) );
  XOR U3435 ( .A(x[114]), .B(x[116]), .Z(n440) );
  NANDN U3436 ( .A(n425), .B(n440), .Z(n375) );
  XOR U3437 ( .A(n382), .B(n375), .Z(n401) );
  XNOR U3438 ( .A(n376), .B(n401), .Z(n377) );
  XOR U3439 ( .A(n378), .B(n377), .Z(n414) );
  IV U3440 ( .A(n414), .Z(n420) );
  AND U3441 ( .A(n380), .B(n379), .Z(n385) );
  XOR U3442 ( .A(x[112]), .B(n427), .Z(n428) );
  XNOR U3443 ( .A(n474), .B(n428), .Z(n430) );
  XOR U3444 ( .A(x[114]), .B(x[119]), .Z(n455) );
  NANDN U3445 ( .A(n430), .B(n455), .Z(n381) );
  XNOR U3446 ( .A(n382), .B(n381), .Z(n390) );
  XNOR U3447 ( .A(n383), .B(n390), .Z(n384) );
  XOR U3448 ( .A(n385), .B(n384), .Z(n410) );
  XNOR U3449 ( .A(x[116]), .B(n474), .Z(n448) );
  ANDN U3450 ( .B(x[112]), .A(n448), .Z(n392) );
  XOR U3451 ( .A(x[114]), .B(x[113]), .Z(n386) );
  XOR U3452 ( .A(n463), .B(n386), .Z(n437) );
  XOR U3453 ( .A(n438), .B(n386), .Z(n443) );
  NAND U3454 ( .A(n427), .B(n443), .Z(n394) );
  XNOR U3455 ( .A(n437), .B(n394), .Z(n388) );
  XNOR U3456 ( .A(x[113]), .B(n428), .Z(n387) );
  XNOR U3457 ( .A(n388), .B(n387), .Z(n389) );
  XOR U3458 ( .A(n390), .B(n389), .Z(n391) );
  XOR U3459 ( .A(n392), .B(n391), .Z(n412) );
  NAND U3460 ( .A(n410), .B(n412), .Z(n393) );
  NAND U3461 ( .A(n420), .B(n393), .Z(n404) );
  IV U3462 ( .A(n410), .Z(n411) );
  IV U3463 ( .A(n412), .Z(n418) );
  XOR U3464 ( .A(n394), .B(n448), .Z(n397) );
  AND U3465 ( .A(n437), .B(n428), .Z(n395) );
  XNOR U3466 ( .A(x[112]), .B(n395), .Z(n396) );
  XNOR U3467 ( .A(n397), .B(n396), .Z(n398) );
  XNOR U3468 ( .A(n399), .B(n398), .Z(n400) );
  XNOR U3469 ( .A(n401), .B(n400), .Z(n422) );
  IV U3470 ( .A(n422), .Z(n417) );
  XOR U3471 ( .A(n418), .B(n417), .Z(n402) );
  NAND U3472 ( .A(n411), .B(n402), .Z(n403) );
  AND U3473 ( .A(n404), .B(n403), .Z(n482) );
  NAND U3474 ( .A(n418), .B(n411), .Z(n405) );
  NAND U3475 ( .A(n417), .B(n405), .Z(n408) );
  XOR U3476 ( .A(n411), .B(n414), .Z(n406) );
  NAND U3477 ( .A(n412), .B(n406), .Z(n407) );
  AND U3478 ( .A(n408), .B(n407), .Z(n464) );
  XNOR U3479 ( .A(n482), .B(n464), .Z(n439) );
  OR U3480 ( .A(n439), .B(n409), .Z(n432) );
  NAND U3481 ( .A(n420), .B(n410), .Z(n416) );
  AND U3482 ( .A(n412), .B(n411), .Z(n419) );
  XNOR U3483 ( .A(n417), .B(n419), .Z(n413) );
  NAND U3484 ( .A(n414), .B(n413), .Z(n415) );
  AND U3485 ( .A(n416), .B(n415), .Z(n436) );
  NAND U3486 ( .A(n418), .B(n417), .Z(n424) );
  XNOR U3487 ( .A(n420), .B(n419), .Z(n421) );
  NAND U3488 ( .A(n422), .B(n421), .Z(n423) );
  NAND U3489 ( .A(n424), .B(n423), .Z(n476) );
  XNOR U3490 ( .A(n436), .B(n476), .Z(n454) );
  XOR U3491 ( .A(n454), .B(n439), .Z(n441) );
  OR U3492 ( .A(n441), .B(n425), .Z(n426) );
  XNOR U3493 ( .A(n432), .B(n426), .Z(n458) );
  XOR U3494 ( .A(n436), .B(n482), .Z(n444) );
  NANDN U3495 ( .A(n444), .B(n427), .Z(n484) );
  NANDN U3496 ( .A(n436), .B(n428), .Z(n429) );
  XNOR U3497 ( .A(n484), .B(n429), .Z(n462) );
  XOR U3498 ( .A(n458), .B(n462), .Z(n447) );
  NANDN U3499 ( .A(n430), .B(n454), .Z(n431) );
  XNOR U3500 ( .A(n432), .B(n431), .Z(n490) );
  XNOR U3501 ( .A(n476), .B(n464), .Z(n466) );
  NANDN U3502 ( .A(n466), .B(n433), .Z(n450) );
  NAND U3503 ( .A(n434), .B(n464), .Z(n435) );
  XNOR U3504 ( .A(n450), .B(n435), .Z(n481) );
  XOR U3505 ( .A(n490), .B(n481), .Z(n473) );
  XNOR U3506 ( .A(n447), .B(n473), .Z(z[112]) );
  ANDN U3507 ( .B(n437), .A(n436), .Z(n446) );
  NANDN U3508 ( .A(n439), .B(n438), .Z(n457) );
  NANDN U3509 ( .A(n441), .B(n440), .Z(n442) );
  XNOR U3510 ( .A(n457), .B(n442), .Z(n485) );
  NANDN U3511 ( .A(n444), .B(n443), .Z(n451) );
  XNOR U3512 ( .A(n485), .B(n451), .Z(n445) );
  XOR U3513 ( .A(n446), .B(n445), .Z(n471) );
  XOR U3514 ( .A(n471), .B(n447), .Z(n489) );
  ANDN U3515 ( .B(n482), .A(n448), .Z(n453) );
  NAND U3516 ( .A(n474), .B(n476), .Z(n449) );
  XNOR U3517 ( .A(n450), .B(n449), .Z(n461) );
  XNOR U3518 ( .A(n451), .B(n461), .Z(n452) );
  XNOR U3519 ( .A(n453), .B(n452), .Z(n460) );
  NAND U3520 ( .A(n455), .B(n454), .Z(n456) );
  XNOR U3521 ( .A(n457), .B(n456), .Z(n467) );
  XNOR U3522 ( .A(n458), .B(n467), .Z(n459) );
  XOR U3523 ( .A(n460), .B(n459), .Z(n470) );
  XNOR U3524 ( .A(n489), .B(n470), .Z(z[113]) );
  XNOR U3525 ( .A(n462), .B(n461), .Z(z[114]) );
  AND U3526 ( .A(n464), .B(n463), .Z(n469) );
  NANDN U3527 ( .A(n466), .B(n465), .Z(n479) );
  XNOR U3528 ( .A(n467), .B(n479), .Z(n468) );
  XOR U3529 ( .A(n469), .B(n468), .Z(n488) );
  XOR U3530 ( .A(n471), .B(n470), .Z(n472) );
  XOR U3531 ( .A(n488), .B(n472), .Z(z[115]) );
  XOR U3532 ( .A(n473), .B(z[114]), .Z(z[116]) );
  XNOR U3533 ( .A(n475), .B(n474), .Z(n477) );
  NAND U3534 ( .A(n477), .B(n476), .Z(n478) );
  XOR U3535 ( .A(n479), .B(n478), .Z(n480) );
  XNOR U3536 ( .A(n481), .B(n480), .Z(n487) );
  NAND U3537 ( .A(n482), .B(x[112]), .Z(n483) );
  XNOR U3538 ( .A(n484), .B(n483), .Z(n491) );
  XNOR U3539 ( .A(n485), .B(n491), .Z(n486) );
  XOR U3540 ( .A(n487), .B(n486), .Z(z[117]) );
  XNOR U3541 ( .A(n489), .B(n488), .Z(z[118]) );
  XNOR U3542 ( .A(n491), .B(n490), .Z(n492) );
  XNOR U3543 ( .A(z[113]), .B(n492), .Z(z[119]) );
  XNOR U3544 ( .A(n496), .B(n495), .Z(n662) );
  XOR U3545 ( .A(n646), .B(n662), .Z(n506) );
  NANDN U3546 ( .A(n497), .B(n506), .Z(n650) );
  XNOR U3547 ( .A(n658), .B(n504), .Z(n672) );
  XNOR U3548 ( .A(n506), .B(n672), .Z(n509) );
  OR U3549 ( .A(n498), .B(n509), .Z(n499) );
  XNOR U3550 ( .A(n650), .B(n499), .Z(n671) );
  OR U3551 ( .A(n501), .B(n500), .Z(n511) );
  ANDN U3552 ( .B(n502), .A(n662), .Z(n503) );
  XNOR U3553 ( .A(n511), .B(n503), .Z(n678) );
  AND U3554 ( .A(n505), .B(n504), .Z(n513) );
  NAND U3555 ( .A(n507), .B(n506), .Z(n675) );
  OR U3556 ( .A(n509), .B(n508), .Z(n510) );
  XNOR U3557 ( .A(n675), .B(n510), .Z(n667) );
  XNOR U3558 ( .A(n667), .B(n511), .Z(n512) );
  XOR U3559 ( .A(n513), .B(n512), .Z(n682) );
  NANDN U3560 ( .A(n515), .B(n514), .Z(n660) );
  OR U3561 ( .A(n516), .B(n646), .Z(n517) );
  XOR U3562 ( .A(n660), .B(n517), .Z(n518) );
  XNOR U3563 ( .A(n682), .B(n518), .Z(n677) );
  XNOR U3564 ( .A(n519), .B(n677), .Z(n520) );
  XOR U3565 ( .A(n678), .B(n520), .Z(n521) );
  XOR U3566 ( .A(n671), .B(n521), .Z(z[11]) );
  IV U3567 ( .A(x[121]), .Z(n628) );
  XOR U3568 ( .A(x[120]), .B(x[126]), .Z(n523) );
  XOR U3569 ( .A(x[125]), .B(n523), .Z(n627) );
  IV U3570 ( .A(n627), .Z(n524) );
  AND U3571 ( .A(n628), .B(n524), .Z(n531) );
  XNOR U3572 ( .A(x[123]), .B(n628), .Z(n527) );
  XNOR U3573 ( .A(x[122]), .B(n527), .Z(n522) );
  XNOR U3574 ( .A(n523), .B(n522), .Z(n587) );
  IV U3575 ( .A(n587), .Z(n533) );
  XNOR U3576 ( .A(n533), .B(n627), .Z(n586) );
  IV U3577 ( .A(x[127]), .Z(n525) );
  XNOR U3578 ( .A(x[121]), .B(n525), .Z(n618) );
  NAND U3579 ( .A(n586), .B(n618), .Z(n536) );
  XNOR U3580 ( .A(n525), .B(n524), .Z(n532) );
  IV U3581 ( .A(n532), .Z(n616) );
  XOR U3582 ( .A(n587), .B(n616), .Z(n552) );
  XNOR U3583 ( .A(n536), .B(n552), .Z(n529) );
  XOR U3584 ( .A(x[120]), .B(n533), .Z(n562) );
  XOR U3585 ( .A(x[124]), .B(n525), .Z(n526) );
  IV U3586 ( .A(n526), .Z(n591) );
  NANDN U3587 ( .A(n562), .B(n591), .Z(n535) );
  XNOR U3588 ( .A(n527), .B(n526), .Z(n580) );
  XNOR U3589 ( .A(n586), .B(n580), .Z(n578) );
  XOR U3590 ( .A(x[122]), .B(x[124]), .Z(n593) );
  NANDN U3591 ( .A(n578), .B(n593), .Z(n528) );
  XOR U3592 ( .A(n535), .B(n528), .Z(n554) );
  XNOR U3593 ( .A(n529), .B(n554), .Z(n530) );
  XOR U3594 ( .A(n531), .B(n530), .Z(n567) );
  IV U3595 ( .A(n567), .Z(n573) );
  AND U3596 ( .A(n533), .B(n532), .Z(n538) );
  XOR U3597 ( .A(x[120]), .B(n580), .Z(n581) );
  XNOR U3598 ( .A(n627), .B(n581), .Z(n583) );
  XOR U3599 ( .A(x[122]), .B(x[127]), .Z(n608) );
  NANDN U3600 ( .A(n583), .B(n608), .Z(n534) );
  XNOR U3601 ( .A(n535), .B(n534), .Z(n543) );
  XNOR U3602 ( .A(n536), .B(n543), .Z(n537) );
  XOR U3603 ( .A(n538), .B(n537), .Z(n563) );
  XNOR U3604 ( .A(x[124]), .B(n627), .Z(n601) );
  ANDN U3605 ( .B(x[120]), .A(n601), .Z(n545) );
  XOR U3606 ( .A(x[122]), .B(x[121]), .Z(n539) );
  XOR U3607 ( .A(n616), .B(n539), .Z(n590) );
  XOR U3608 ( .A(n591), .B(n539), .Z(n596) );
  NAND U3609 ( .A(n580), .B(n596), .Z(n547) );
  XNOR U3610 ( .A(n590), .B(n547), .Z(n541) );
  XNOR U3611 ( .A(x[121]), .B(n581), .Z(n540) );
  XNOR U3612 ( .A(n541), .B(n540), .Z(n542) );
  XOR U3613 ( .A(n543), .B(n542), .Z(n544) );
  XOR U3614 ( .A(n545), .B(n544), .Z(n565) );
  NAND U3615 ( .A(n563), .B(n565), .Z(n546) );
  NAND U3616 ( .A(n573), .B(n546), .Z(n557) );
  IV U3617 ( .A(n563), .Z(n564) );
  IV U3618 ( .A(n565), .Z(n571) );
  XOR U3619 ( .A(n547), .B(n601), .Z(n550) );
  AND U3620 ( .A(n590), .B(n581), .Z(n548) );
  XNOR U3621 ( .A(x[120]), .B(n548), .Z(n549) );
  XNOR U3622 ( .A(n550), .B(n549), .Z(n551) );
  XNOR U3623 ( .A(n552), .B(n551), .Z(n553) );
  XNOR U3624 ( .A(n554), .B(n553), .Z(n575) );
  IV U3625 ( .A(n575), .Z(n570) );
  XOR U3626 ( .A(n571), .B(n570), .Z(n555) );
  NAND U3627 ( .A(n564), .B(n555), .Z(n556) );
  AND U3628 ( .A(n557), .B(n556), .Z(n635) );
  NAND U3629 ( .A(n571), .B(n564), .Z(n558) );
  NAND U3630 ( .A(n570), .B(n558), .Z(n561) );
  XOR U3631 ( .A(n564), .B(n567), .Z(n559) );
  NAND U3632 ( .A(n565), .B(n559), .Z(n560) );
  AND U3633 ( .A(n561), .B(n560), .Z(n617) );
  XNOR U3634 ( .A(n635), .B(n617), .Z(n592) );
  OR U3635 ( .A(n592), .B(n562), .Z(n585) );
  NAND U3636 ( .A(n573), .B(n563), .Z(n569) );
  AND U3637 ( .A(n565), .B(n564), .Z(n572) );
  XNOR U3638 ( .A(n570), .B(n572), .Z(n566) );
  NAND U3639 ( .A(n567), .B(n566), .Z(n568) );
  AND U3640 ( .A(n569), .B(n568), .Z(n589) );
  NAND U3641 ( .A(n571), .B(n570), .Z(n577) );
  XNOR U3642 ( .A(n573), .B(n572), .Z(n574) );
  NAND U3643 ( .A(n575), .B(n574), .Z(n576) );
  NAND U3644 ( .A(n577), .B(n576), .Z(n629) );
  XNOR U3645 ( .A(n589), .B(n629), .Z(n607) );
  XOR U3646 ( .A(n607), .B(n592), .Z(n594) );
  OR U3647 ( .A(n594), .B(n578), .Z(n579) );
  XNOR U3648 ( .A(n585), .B(n579), .Z(n611) );
  XOR U3649 ( .A(n589), .B(n635), .Z(n597) );
  NANDN U3650 ( .A(n597), .B(n580), .Z(n637) );
  NANDN U3651 ( .A(n589), .B(n581), .Z(n582) );
  XNOR U3652 ( .A(n637), .B(n582), .Z(n615) );
  XOR U3653 ( .A(n611), .B(n615), .Z(n600) );
  NANDN U3654 ( .A(n583), .B(n607), .Z(n584) );
  XNOR U3655 ( .A(n585), .B(n584), .Z(n643) );
  XNOR U3656 ( .A(n629), .B(n617), .Z(n619) );
  NANDN U3657 ( .A(n619), .B(n586), .Z(n603) );
  NAND U3658 ( .A(n587), .B(n617), .Z(n588) );
  XNOR U3659 ( .A(n603), .B(n588), .Z(n634) );
  XOR U3660 ( .A(n643), .B(n634), .Z(n626) );
  XNOR U3661 ( .A(n600), .B(n626), .Z(z[120]) );
  ANDN U3662 ( .B(n590), .A(n589), .Z(n599) );
  NANDN U3663 ( .A(n592), .B(n591), .Z(n610) );
  NANDN U3664 ( .A(n594), .B(n593), .Z(n595) );
  XNOR U3665 ( .A(n610), .B(n595), .Z(n638) );
  NANDN U3666 ( .A(n597), .B(n596), .Z(n604) );
  XNOR U3667 ( .A(n638), .B(n604), .Z(n598) );
  XOR U3668 ( .A(n599), .B(n598), .Z(n624) );
  XOR U3669 ( .A(n624), .B(n600), .Z(n642) );
  ANDN U3670 ( .B(n635), .A(n601), .Z(n606) );
  NAND U3671 ( .A(n627), .B(n629), .Z(n602) );
  XNOR U3672 ( .A(n603), .B(n602), .Z(n614) );
  XNOR U3673 ( .A(n604), .B(n614), .Z(n605) );
  XNOR U3674 ( .A(n606), .B(n605), .Z(n613) );
  NAND U3675 ( .A(n608), .B(n607), .Z(n609) );
  XNOR U3676 ( .A(n610), .B(n609), .Z(n620) );
  XNOR U3677 ( .A(n611), .B(n620), .Z(n612) );
  XOR U3678 ( .A(n613), .B(n612), .Z(n623) );
  XNOR U3679 ( .A(n642), .B(n623), .Z(z[121]) );
  XNOR U3680 ( .A(n615), .B(n614), .Z(z[122]) );
  AND U3681 ( .A(n617), .B(n616), .Z(n622) );
  NANDN U3682 ( .A(n619), .B(n618), .Z(n632) );
  XNOR U3683 ( .A(n620), .B(n632), .Z(n621) );
  XOR U3684 ( .A(n622), .B(n621), .Z(n641) );
  XOR U3685 ( .A(n624), .B(n623), .Z(n625) );
  XOR U3686 ( .A(n641), .B(n625), .Z(z[123]) );
  XOR U3687 ( .A(n626), .B(z[122]), .Z(z[124]) );
  XNOR U3688 ( .A(n628), .B(n627), .Z(n630) );
  NAND U3689 ( .A(n630), .B(n629), .Z(n631) );
  XOR U3690 ( .A(n632), .B(n631), .Z(n633) );
  XNOR U3691 ( .A(n634), .B(n633), .Z(n640) );
  NAND U3692 ( .A(n635), .B(x[120]), .Z(n636) );
  XNOR U3693 ( .A(n637), .B(n636), .Z(n644) );
  XNOR U3694 ( .A(n638), .B(n644), .Z(n639) );
  XOR U3695 ( .A(n640), .B(n639), .Z(z[125]) );
  XNOR U3696 ( .A(n642), .B(n641), .Z(z[126]) );
  XNOR U3697 ( .A(n644), .B(n643), .Z(n645) );
  XNOR U3698 ( .A(z[121]), .B(n645), .Z(z[127]) );
  NOR U3699 ( .A(n647), .B(n646), .Z(n653) );
  NANDN U3700 ( .A(n648), .B(n672), .Z(n649) );
  XNOR U3701 ( .A(n650), .B(n649), .Z(n663) );
  XNOR U3702 ( .A(n651), .B(n663), .Z(n652) );
  XOR U3703 ( .A(n653), .B(n652), .Z(n1947) );
  XOR U3704 ( .A(n1947), .B(n654), .Z(z[12]) );
  XNOR U3705 ( .A(n656), .B(n655), .Z(n657) );
  NANDN U3706 ( .A(n658), .B(n657), .Z(n659) );
  XOR U3707 ( .A(n660), .B(n659), .Z(n661) );
  XNOR U3708 ( .A(n1947), .B(n661), .Z(n669) );
  ANDN U3709 ( .B(x[8]), .A(n662), .Z(n666) );
  XNOR U3710 ( .A(n664), .B(n663), .Z(n665) );
  XOR U3711 ( .A(n666), .B(n665), .Z(n683) );
  XNOR U3712 ( .A(n667), .B(n683), .Z(n668) );
  XOR U3713 ( .A(n669), .B(n668), .Z(z[13]) );
  XNOR U3714 ( .A(n671), .B(n670), .Z(n1948) );
  NAND U3715 ( .A(n673), .B(n672), .Z(n674) );
  XNOR U3716 ( .A(n675), .B(n674), .Z(n679) );
  XNOR U3717 ( .A(n1948), .B(n679), .Z(n676) );
  XOR U3718 ( .A(n677), .B(n676), .Z(z[14]) );
  XNOR U3719 ( .A(n679), .B(n678), .Z(n680) );
  XNOR U3720 ( .A(z[10]), .B(n680), .Z(n681) );
  XOR U3721 ( .A(n682), .B(n681), .Z(z[9]) );
  XNOR U3722 ( .A(n683), .B(z[9]), .Z(z[15]) );
  IV U3723 ( .A(x[17]), .Z(n815) );
  IV U3724 ( .A(n814), .Z(n686) );
  AND U3725 ( .A(n815), .B(n686), .Z(n693) );
  XNOR U3726 ( .A(x[19]), .B(n815), .Z(n689) );
  XNOR U3727 ( .A(x[18]), .B(n689), .Z(n684) );
  XNOR U3728 ( .A(n685), .B(n684), .Z(n749) );
  IV U3729 ( .A(n749), .Z(n695) );
  XNOR U3730 ( .A(n695), .B(n814), .Z(n748) );
  IV U3731 ( .A(x[23]), .Z(n687) );
  XNOR U3732 ( .A(x[17]), .B(n687), .Z(n780) );
  NAND U3733 ( .A(n748), .B(n780), .Z(n698) );
  XNOR U3734 ( .A(n687), .B(n686), .Z(n694) );
  IV U3735 ( .A(n694), .Z(n778) );
  XOR U3736 ( .A(n749), .B(n778), .Z(n714) );
  XNOR U3737 ( .A(n698), .B(n714), .Z(n691) );
  XOR U3738 ( .A(x[16]), .B(n695), .Z(n724) );
  XOR U3739 ( .A(x[20]), .B(n687), .Z(n688) );
  IV U3740 ( .A(n688), .Z(n753) );
  NANDN U3741 ( .A(n724), .B(n753), .Z(n697) );
  XNOR U3742 ( .A(n689), .B(n688), .Z(n742) );
  XNOR U3743 ( .A(n748), .B(n742), .Z(n740) );
  XOR U3744 ( .A(x[18]), .B(x[20]), .Z(n755) );
  NANDN U3745 ( .A(n740), .B(n755), .Z(n690) );
  XOR U3746 ( .A(n697), .B(n690), .Z(n716) );
  XNOR U3747 ( .A(n691), .B(n716), .Z(n692) );
  XOR U3748 ( .A(n693), .B(n692), .Z(n729) );
  IV U3749 ( .A(n729), .Z(n735) );
  AND U3750 ( .A(n695), .B(n694), .Z(n700) );
  XOR U3751 ( .A(x[16]), .B(n742), .Z(n743) );
  XNOR U3752 ( .A(n814), .B(n743), .Z(n745) );
  XOR U3753 ( .A(x[18]), .B(x[23]), .Z(n770) );
  NANDN U3754 ( .A(n745), .B(n770), .Z(n696) );
  XNOR U3755 ( .A(n697), .B(n696), .Z(n705) );
  XNOR U3756 ( .A(n698), .B(n705), .Z(n699) );
  XOR U3757 ( .A(n700), .B(n699), .Z(n725) );
  XNOR U3758 ( .A(x[20]), .B(n814), .Z(n763) );
  ANDN U3759 ( .B(x[16]), .A(n763), .Z(n707) );
  XOR U3760 ( .A(x[18]), .B(x[17]), .Z(n701) );
  XOR U3761 ( .A(n778), .B(n701), .Z(n752) );
  XOR U3762 ( .A(n753), .B(n701), .Z(n758) );
  NAND U3763 ( .A(n742), .B(n758), .Z(n709) );
  XNOR U3764 ( .A(n752), .B(n709), .Z(n703) );
  XNOR U3765 ( .A(x[17]), .B(n743), .Z(n702) );
  XNOR U3766 ( .A(n703), .B(n702), .Z(n704) );
  XOR U3767 ( .A(n705), .B(n704), .Z(n706) );
  XOR U3768 ( .A(n707), .B(n706), .Z(n727) );
  NAND U3769 ( .A(n725), .B(n727), .Z(n708) );
  NAND U3770 ( .A(n735), .B(n708), .Z(n719) );
  IV U3771 ( .A(n725), .Z(n726) );
  IV U3772 ( .A(n727), .Z(n733) );
  XOR U3773 ( .A(n709), .B(n763), .Z(n712) );
  AND U3774 ( .A(n752), .B(n743), .Z(n710) );
  XNOR U3775 ( .A(x[16]), .B(n710), .Z(n711) );
  XNOR U3776 ( .A(n712), .B(n711), .Z(n713) );
  XNOR U3777 ( .A(n714), .B(n713), .Z(n715) );
  XNOR U3778 ( .A(n716), .B(n715), .Z(n737) );
  IV U3779 ( .A(n737), .Z(n732) );
  XOR U3780 ( .A(n733), .B(n732), .Z(n717) );
  NAND U3781 ( .A(n726), .B(n717), .Z(n718) );
  AND U3782 ( .A(n719), .B(n718), .Z(n822) );
  NAND U3783 ( .A(n733), .B(n726), .Z(n720) );
  NAND U3784 ( .A(n732), .B(n720), .Z(n723) );
  XOR U3785 ( .A(n726), .B(n729), .Z(n721) );
  NAND U3786 ( .A(n727), .B(n721), .Z(n722) );
  AND U3787 ( .A(n723), .B(n722), .Z(n779) );
  XNOR U3788 ( .A(n822), .B(n779), .Z(n754) );
  OR U3789 ( .A(n754), .B(n724), .Z(n747) );
  NAND U3790 ( .A(n735), .B(n725), .Z(n731) );
  AND U3791 ( .A(n727), .B(n726), .Z(n734) );
  XNOR U3792 ( .A(n732), .B(n734), .Z(n728) );
  NAND U3793 ( .A(n729), .B(n728), .Z(n730) );
  AND U3794 ( .A(n731), .B(n730), .Z(n751) );
  NAND U3795 ( .A(n733), .B(n732), .Z(n739) );
  XNOR U3796 ( .A(n735), .B(n734), .Z(n736) );
  NAND U3797 ( .A(n737), .B(n736), .Z(n738) );
  NAND U3798 ( .A(n739), .B(n738), .Z(n816) );
  XNOR U3799 ( .A(n751), .B(n816), .Z(n769) );
  XOR U3800 ( .A(n769), .B(n754), .Z(n756) );
  OR U3801 ( .A(n756), .B(n740), .Z(n741) );
  XNOR U3802 ( .A(n747), .B(n741), .Z(n773) );
  XOR U3803 ( .A(n751), .B(n822), .Z(n759) );
  NANDN U3804 ( .A(n759), .B(n742), .Z(n824) );
  NANDN U3805 ( .A(n751), .B(n743), .Z(n744) );
  XNOR U3806 ( .A(n824), .B(n744), .Z(n777) );
  XOR U3807 ( .A(n773), .B(n777), .Z(n762) );
  NANDN U3808 ( .A(n745), .B(n769), .Z(n746) );
  XNOR U3809 ( .A(n747), .B(n746), .Z(n830) );
  XNOR U3810 ( .A(n816), .B(n779), .Z(n781) );
  NANDN U3811 ( .A(n781), .B(n748), .Z(n765) );
  NAND U3812 ( .A(n749), .B(n779), .Z(n750) );
  XNOR U3813 ( .A(n765), .B(n750), .Z(n821) );
  XOR U3814 ( .A(n830), .B(n821), .Z(n813) );
  XNOR U3815 ( .A(n762), .B(n813), .Z(z[16]) );
  ANDN U3816 ( .B(n752), .A(n751), .Z(n761) );
  NANDN U3817 ( .A(n754), .B(n753), .Z(n772) );
  NANDN U3818 ( .A(n756), .B(n755), .Z(n757) );
  XNOR U3819 ( .A(n772), .B(n757), .Z(n825) );
  NANDN U3820 ( .A(n759), .B(n758), .Z(n766) );
  XNOR U3821 ( .A(n825), .B(n766), .Z(n760) );
  XOR U3822 ( .A(n761), .B(n760), .Z(n786) );
  XOR U3823 ( .A(n786), .B(n762), .Z(n829) );
  ANDN U3824 ( .B(n822), .A(n763), .Z(n768) );
  NAND U3825 ( .A(n814), .B(n816), .Z(n764) );
  XNOR U3826 ( .A(n765), .B(n764), .Z(n776) );
  XNOR U3827 ( .A(n766), .B(n776), .Z(n767) );
  XNOR U3828 ( .A(n768), .B(n767), .Z(n775) );
  NAND U3829 ( .A(n770), .B(n769), .Z(n771) );
  XNOR U3830 ( .A(n772), .B(n771), .Z(n782) );
  XNOR U3831 ( .A(n773), .B(n782), .Z(n774) );
  XOR U3832 ( .A(n775), .B(n774), .Z(n785) );
  XNOR U3833 ( .A(n829), .B(n785), .Z(z[17]) );
  XNOR U3834 ( .A(n777), .B(n776), .Z(z[18]) );
  AND U3835 ( .A(n779), .B(n778), .Z(n784) );
  NANDN U3836 ( .A(n781), .B(n780), .Z(n819) );
  XNOR U3837 ( .A(n782), .B(n819), .Z(n783) );
  XOR U3838 ( .A(n784), .B(n783), .Z(n828) );
  XOR U3839 ( .A(n786), .B(n785), .Z(n787) );
  XOR U3840 ( .A(n828), .B(n787), .Z(z[19]) );
  ANDN U3841 ( .B(n789), .A(n788), .Z(n798) );
  NANDN U3842 ( .A(n791), .B(n790), .Z(n809) );
  NANDN U3843 ( .A(n793), .B(n792), .Z(n794) );
  XNOR U3844 ( .A(n809), .B(n794), .Z(n1457) );
  NANDN U3845 ( .A(n796), .B(n795), .Z(n803) );
  XNOR U3846 ( .A(n1457), .B(n803), .Z(n797) );
  XOR U3847 ( .A(n798), .B(n797), .Z(n1091) );
  XOR U3848 ( .A(n1091), .B(n799), .Z(n1600) );
  ANDN U3849 ( .B(n1454), .A(n800), .Z(n805) );
  NAND U3850 ( .A(n1446), .B(n1448), .Z(n801) );
  XNOR U3851 ( .A(n802), .B(n801), .Z(n952) );
  XNOR U3852 ( .A(n803), .B(n952), .Z(n804) );
  XNOR U3853 ( .A(n805), .B(n804), .Z(n812) );
  NAND U3854 ( .A(n807), .B(n806), .Z(n808) );
  XNOR U3855 ( .A(n809), .B(n808), .Z(n1087) );
  XNOR U3856 ( .A(n810), .B(n1087), .Z(n811) );
  XOR U3857 ( .A(n812), .B(n811), .Z(n1090) );
  XNOR U3858 ( .A(n1600), .B(n1090), .Z(z[1]) );
  XOR U3859 ( .A(n813), .B(z[18]), .Z(z[20]) );
  XNOR U3860 ( .A(n815), .B(n814), .Z(n817) );
  NAND U3861 ( .A(n817), .B(n816), .Z(n818) );
  XOR U3862 ( .A(n819), .B(n818), .Z(n820) );
  XNOR U3863 ( .A(n821), .B(n820), .Z(n827) );
  NAND U3864 ( .A(n822), .B(x[16]), .Z(n823) );
  XNOR U3865 ( .A(n824), .B(n823), .Z(n831) );
  XNOR U3866 ( .A(n825), .B(n831), .Z(n826) );
  XOR U3867 ( .A(n827), .B(n826), .Z(z[21]) );
  XNOR U3868 ( .A(n829), .B(n828), .Z(z[22]) );
  XNOR U3869 ( .A(n831), .B(n830), .Z(n832) );
  XNOR U3870 ( .A(z[17]), .B(n832), .Z(z[23]) );
  IV U3871 ( .A(x[25]), .Z(n939) );
  XOR U3872 ( .A(x[24]), .B(x[30]), .Z(n834) );
  XOR U3873 ( .A(x[29]), .B(n834), .Z(n938) );
  IV U3874 ( .A(n938), .Z(n835) );
  AND U3875 ( .A(n939), .B(n835), .Z(n842) );
  XNOR U3876 ( .A(x[27]), .B(n939), .Z(n838) );
  XNOR U3877 ( .A(x[26]), .B(n838), .Z(n833) );
  XNOR U3878 ( .A(n834), .B(n833), .Z(n898) );
  IV U3879 ( .A(n898), .Z(n844) );
  XNOR U3880 ( .A(n844), .B(n938), .Z(n897) );
  IV U3881 ( .A(x[31]), .Z(n836) );
  XNOR U3882 ( .A(x[25]), .B(n836), .Z(n929) );
  NAND U3883 ( .A(n897), .B(n929), .Z(n847) );
  XNOR U3884 ( .A(n836), .B(n835), .Z(n843) );
  IV U3885 ( .A(n843), .Z(n927) );
  XOR U3886 ( .A(n898), .B(n927), .Z(n863) );
  XNOR U3887 ( .A(n847), .B(n863), .Z(n840) );
  XOR U3888 ( .A(x[24]), .B(n844), .Z(n873) );
  XOR U3889 ( .A(x[28]), .B(n836), .Z(n837) );
  IV U3890 ( .A(n837), .Z(n902) );
  NANDN U3891 ( .A(n873), .B(n902), .Z(n846) );
  XNOR U3892 ( .A(n838), .B(n837), .Z(n891) );
  XNOR U3893 ( .A(n897), .B(n891), .Z(n889) );
  XOR U3894 ( .A(x[26]), .B(x[28]), .Z(n904) );
  NANDN U3895 ( .A(n889), .B(n904), .Z(n839) );
  XOR U3896 ( .A(n846), .B(n839), .Z(n865) );
  XNOR U3897 ( .A(n840), .B(n865), .Z(n841) );
  XOR U3898 ( .A(n842), .B(n841), .Z(n878) );
  IV U3899 ( .A(n878), .Z(n884) );
  AND U3900 ( .A(n844), .B(n843), .Z(n849) );
  XOR U3901 ( .A(x[24]), .B(n891), .Z(n892) );
  XNOR U3902 ( .A(n938), .B(n892), .Z(n894) );
  XOR U3903 ( .A(x[26]), .B(x[31]), .Z(n919) );
  NANDN U3904 ( .A(n894), .B(n919), .Z(n845) );
  XNOR U3905 ( .A(n846), .B(n845), .Z(n854) );
  XNOR U3906 ( .A(n847), .B(n854), .Z(n848) );
  XOR U3907 ( .A(n849), .B(n848), .Z(n874) );
  XNOR U3908 ( .A(x[28]), .B(n938), .Z(n912) );
  ANDN U3909 ( .B(x[24]), .A(n912), .Z(n856) );
  XOR U3910 ( .A(x[26]), .B(x[25]), .Z(n850) );
  XOR U3911 ( .A(n927), .B(n850), .Z(n901) );
  XOR U3912 ( .A(n902), .B(n850), .Z(n907) );
  NAND U3913 ( .A(n891), .B(n907), .Z(n858) );
  XNOR U3914 ( .A(n901), .B(n858), .Z(n852) );
  XNOR U3915 ( .A(x[25]), .B(n892), .Z(n851) );
  XNOR U3916 ( .A(n852), .B(n851), .Z(n853) );
  XOR U3917 ( .A(n854), .B(n853), .Z(n855) );
  XOR U3918 ( .A(n856), .B(n855), .Z(n876) );
  NAND U3919 ( .A(n874), .B(n876), .Z(n857) );
  NAND U3920 ( .A(n884), .B(n857), .Z(n868) );
  IV U3921 ( .A(n874), .Z(n875) );
  IV U3922 ( .A(n876), .Z(n882) );
  XOR U3923 ( .A(n858), .B(n912), .Z(n861) );
  AND U3924 ( .A(n901), .B(n892), .Z(n859) );
  XNOR U3925 ( .A(x[24]), .B(n859), .Z(n860) );
  XNOR U3926 ( .A(n861), .B(n860), .Z(n862) );
  XNOR U3927 ( .A(n863), .B(n862), .Z(n864) );
  XNOR U3928 ( .A(n865), .B(n864), .Z(n886) );
  IV U3929 ( .A(n886), .Z(n881) );
  XOR U3930 ( .A(n882), .B(n881), .Z(n866) );
  NAND U3931 ( .A(n875), .B(n866), .Z(n867) );
  AND U3932 ( .A(n868), .B(n867), .Z(n946) );
  NAND U3933 ( .A(n882), .B(n875), .Z(n869) );
  NAND U3934 ( .A(n881), .B(n869), .Z(n872) );
  XOR U3935 ( .A(n875), .B(n878), .Z(n870) );
  NAND U3936 ( .A(n876), .B(n870), .Z(n871) );
  AND U3937 ( .A(n872), .B(n871), .Z(n928) );
  XNOR U3938 ( .A(n946), .B(n928), .Z(n903) );
  OR U3939 ( .A(n903), .B(n873), .Z(n896) );
  NAND U3940 ( .A(n884), .B(n874), .Z(n880) );
  AND U3941 ( .A(n876), .B(n875), .Z(n883) );
  XNOR U3942 ( .A(n881), .B(n883), .Z(n877) );
  NAND U3943 ( .A(n878), .B(n877), .Z(n879) );
  AND U3944 ( .A(n880), .B(n879), .Z(n900) );
  NAND U3945 ( .A(n882), .B(n881), .Z(n888) );
  XNOR U3946 ( .A(n884), .B(n883), .Z(n885) );
  NAND U3947 ( .A(n886), .B(n885), .Z(n887) );
  NAND U3948 ( .A(n888), .B(n887), .Z(n940) );
  XNOR U3949 ( .A(n900), .B(n940), .Z(n918) );
  XOR U3950 ( .A(n918), .B(n903), .Z(n905) );
  OR U3951 ( .A(n905), .B(n889), .Z(n890) );
  XNOR U3952 ( .A(n896), .B(n890), .Z(n922) );
  XOR U3953 ( .A(n900), .B(n946), .Z(n908) );
  NANDN U3954 ( .A(n908), .B(n891), .Z(n948) );
  NANDN U3955 ( .A(n900), .B(n892), .Z(n893) );
  XNOR U3956 ( .A(n948), .B(n893), .Z(n926) );
  XOR U3957 ( .A(n922), .B(n926), .Z(n911) );
  NANDN U3958 ( .A(n894), .B(n918), .Z(n895) );
  XNOR U3959 ( .A(n896), .B(n895), .Z(n956) );
  XNOR U3960 ( .A(n940), .B(n928), .Z(n930) );
  NANDN U3961 ( .A(n930), .B(n897), .Z(n914) );
  NAND U3962 ( .A(n898), .B(n928), .Z(n899) );
  XNOR U3963 ( .A(n914), .B(n899), .Z(n945) );
  XOR U3964 ( .A(n956), .B(n945), .Z(n937) );
  XNOR U3965 ( .A(n911), .B(n937), .Z(z[24]) );
  ANDN U3966 ( .B(n901), .A(n900), .Z(n910) );
  NANDN U3967 ( .A(n903), .B(n902), .Z(n921) );
  NANDN U3968 ( .A(n905), .B(n904), .Z(n906) );
  XNOR U3969 ( .A(n921), .B(n906), .Z(n949) );
  NANDN U3970 ( .A(n908), .B(n907), .Z(n915) );
  XNOR U3971 ( .A(n949), .B(n915), .Z(n909) );
  XOR U3972 ( .A(n910), .B(n909), .Z(n935) );
  XOR U3973 ( .A(n935), .B(n911), .Z(n955) );
  ANDN U3974 ( .B(n946), .A(n912), .Z(n917) );
  NAND U3975 ( .A(n938), .B(n940), .Z(n913) );
  XNOR U3976 ( .A(n914), .B(n913), .Z(n925) );
  XNOR U3977 ( .A(n915), .B(n925), .Z(n916) );
  XNOR U3978 ( .A(n917), .B(n916), .Z(n924) );
  NAND U3979 ( .A(n919), .B(n918), .Z(n920) );
  XNOR U3980 ( .A(n921), .B(n920), .Z(n931) );
  XNOR U3981 ( .A(n922), .B(n931), .Z(n923) );
  XOR U3982 ( .A(n924), .B(n923), .Z(n934) );
  XNOR U3983 ( .A(n955), .B(n934), .Z(z[25]) );
  XNOR U3984 ( .A(n926), .B(n925), .Z(z[26]) );
  AND U3985 ( .A(n928), .B(n927), .Z(n933) );
  NANDN U3986 ( .A(n930), .B(n929), .Z(n943) );
  XNOR U3987 ( .A(n931), .B(n943), .Z(n932) );
  XOR U3988 ( .A(n933), .B(n932), .Z(n954) );
  XOR U3989 ( .A(n935), .B(n934), .Z(n936) );
  XOR U3990 ( .A(n954), .B(n936), .Z(z[27]) );
  XOR U3991 ( .A(n937), .B(z[26]), .Z(z[28]) );
  XNOR U3992 ( .A(n939), .B(n938), .Z(n941) );
  NAND U3993 ( .A(n941), .B(n940), .Z(n942) );
  XOR U3994 ( .A(n943), .B(n942), .Z(n944) );
  XNOR U3995 ( .A(n945), .B(n944), .Z(n951) );
  NAND U3996 ( .A(n946), .B(x[24]), .Z(n947) );
  XNOR U3997 ( .A(n948), .B(n947), .Z(n957) );
  XNOR U3998 ( .A(n949), .B(n957), .Z(n950) );
  XOR U3999 ( .A(n951), .B(n950), .Z(z[29]) );
  XNOR U4000 ( .A(n953), .B(n952), .Z(z[2]) );
  XNOR U4001 ( .A(n955), .B(n954), .Z(z[30]) );
  XNOR U4002 ( .A(n957), .B(n956), .Z(n958) );
  XNOR U4003 ( .A(z[25]), .B(n958), .Z(z[31]) );
  IV U4004 ( .A(x[33]), .Z(n1065) );
  XOR U4005 ( .A(x[32]), .B(x[38]), .Z(n960) );
  XOR U4006 ( .A(x[37]), .B(n960), .Z(n1064) );
  IV U4007 ( .A(n1064), .Z(n961) );
  AND U4008 ( .A(n1065), .B(n961), .Z(n968) );
  XNOR U4009 ( .A(x[35]), .B(n1065), .Z(n964) );
  XNOR U4010 ( .A(x[34]), .B(n964), .Z(n959) );
  XNOR U4011 ( .A(n960), .B(n959), .Z(n1024) );
  IV U4012 ( .A(n1024), .Z(n970) );
  XNOR U4013 ( .A(n970), .B(n1064), .Z(n1023) );
  IV U4014 ( .A(x[39]), .Z(n962) );
  XNOR U4015 ( .A(x[33]), .B(n962), .Z(n1055) );
  NAND U4016 ( .A(n1023), .B(n1055), .Z(n973) );
  XNOR U4017 ( .A(n962), .B(n961), .Z(n969) );
  IV U4018 ( .A(n969), .Z(n1053) );
  XOR U4019 ( .A(n1024), .B(n1053), .Z(n989) );
  XNOR U4020 ( .A(n973), .B(n989), .Z(n966) );
  XOR U4021 ( .A(x[32]), .B(n970), .Z(n999) );
  XOR U4022 ( .A(x[36]), .B(n962), .Z(n963) );
  IV U4023 ( .A(n963), .Z(n1028) );
  NANDN U4024 ( .A(n999), .B(n1028), .Z(n972) );
  XNOR U4025 ( .A(n964), .B(n963), .Z(n1017) );
  XNOR U4026 ( .A(n1023), .B(n1017), .Z(n1015) );
  XOR U4027 ( .A(x[34]), .B(x[36]), .Z(n1030) );
  NANDN U4028 ( .A(n1015), .B(n1030), .Z(n965) );
  XOR U4029 ( .A(n972), .B(n965), .Z(n991) );
  XNOR U4030 ( .A(n966), .B(n991), .Z(n967) );
  XOR U4031 ( .A(n968), .B(n967), .Z(n1004) );
  IV U4032 ( .A(n1004), .Z(n1010) );
  AND U4033 ( .A(n970), .B(n969), .Z(n975) );
  XOR U4034 ( .A(x[32]), .B(n1017), .Z(n1018) );
  XNOR U4035 ( .A(n1064), .B(n1018), .Z(n1020) );
  XOR U4036 ( .A(x[34]), .B(x[39]), .Z(n1045) );
  NANDN U4037 ( .A(n1020), .B(n1045), .Z(n971) );
  XNOR U4038 ( .A(n972), .B(n971), .Z(n980) );
  XNOR U4039 ( .A(n973), .B(n980), .Z(n974) );
  XOR U4040 ( .A(n975), .B(n974), .Z(n1000) );
  XNOR U4041 ( .A(x[36]), .B(n1064), .Z(n1038) );
  ANDN U4042 ( .B(x[32]), .A(n1038), .Z(n982) );
  XOR U4043 ( .A(x[34]), .B(x[33]), .Z(n976) );
  XOR U4044 ( .A(n1053), .B(n976), .Z(n1027) );
  XOR U4045 ( .A(n1028), .B(n976), .Z(n1033) );
  NAND U4046 ( .A(n1017), .B(n1033), .Z(n984) );
  XNOR U4047 ( .A(n1027), .B(n984), .Z(n978) );
  XNOR U4048 ( .A(x[33]), .B(n1018), .Z(n977) );
  XNOR U4049 ( .A(n978), .B(n977), .Z(n979) );
  XOR U4050 ( .A(n980), .B(n979), .Z(n981) );
  XOR U4051 ( .A(n982), .B(n981), .Z(n1002) );
  NAND U4052 ( .A(n1000), .B(n1002), .Z(n983) );
  NAND U4053 ( .A(n1010), .B(n983), .Z(n994) );
  IV U4054 ( .A(n1000), .Z(n1001) );
  IV U4055 ( .A(n1002), .Z(n1008) );
  XOR U4056 ( .A(n984), .B(n1038), .Z(n987) );
  AND U4057 ( .A(n1027), .B(n1018), .Z(n985) );
  XNOR U4058 ( .A(x[32]), .B(n985), .Z(n986) );
  XNOR U4059 ( .A(n987), .B(n986), .Z(n988) );
  XNOR U4060 ( .A(n989), .B(n988), .Z(n990) );
  XNOR U4061 ( .A(n991), .B(n990), .Z(n1012) );
  IV U4062 ( .A(n1012), .Z(n1007) );
  XOR U4063 ( .A(n1008), .B(n1007), .Z(n992) );
  NAND U4064 ( .A(n1001), .B(n992), .Z(n993) );
  AND U4065 ( .A(n994), .B(n993), .Z(n1072) );
  NAND U4066 ( .A(n1008), .B(n1001), .Z(n995) );
  NAND U4067 ( .A(n1007), .B(n995), .Z(n998) );
  XOR U4068 ( .A(n1001), .B(n1004), .Z(n996) );
  NAND U4069 ( .A(n1002), .B(n996), .Z(n997) );
  AND U4070 ( .A(n998), .B(n997), .Z(n1054) );
  XNOR U4071 ( .A(n1072), .B(n1054), .Z(n1029) );
  OR U4072 ( .A(n1029), .B(n999), .Z(n1022) );
  NAND U4073 ( .A(n1010), .B(n1000), .Z(n1006) );
  AND U4074 ( .A(n1002), .B(n1001), .Z(n1009) );
  XNOR U4075 ( .A(n1007), .B(n1009), .Z(n1003) );
  NAND U4076 ( .A(n1004), .B(n1003), .Z(n1005) );
  AND U4077 ( .A(n1006), .B(n1005), .Z(n1026) );
  NAND U4078 ( .A(n1008), .B(n1007), .Z(n1014) );
  XNOR U4079 ( .A(n1010), .B(n1009), .Z(n1011) );
  NAND U4080 ( .A(n1012), .B(n1011), .Z(n1013) );
  NAND U4081 ( .A(n1014), .B(n1013), .Z(n1066) );
  XNOR U4082 ( .A(n1026), .B(n1066), .Z(n1044) );
  XOR U4083 ( .A(n1044), .B(n1029), .Z(n1031) );
  OR U4084 ( .A(n1031), .B(n1015), .Z(n1016) );
  XNOR U4085 ( .A(n1022), .B(n1016), .Z(n1048) );
  XOR U4086 ( .A(n1026), .B(n1072), .Z(n1034) );
  NANDN U4087 ( .A(n1034), .B(n1017), .Z(n1074) );
  NANDN U4088 ( .A(n1026), .B(n1018), .Z(n1019) );
  XNOR U4089 ( .A(n1074), .B(n1019), .Z(n1052) );
  XOR U4090 ( .A(n1048), .B(n1052), .Z(n1037) );
  NANDN U4091 ( .A(n1020), .B(n1044), .Z(n1021) );
  XNOR U4092 ( .A(n1022), .B(n1021), .Z(n1080) );
  XNOR U4093 ( .A(n1066), .B(n1054), .Z(n1056) );
  NANDN U4094 ( .A(n1056), .B(n1023), .Z(n1040) );
  NAND U4095 ( .A(n1024), .B(n1054), .Z(n1025) );
  XNOR U4096 ( .A(n1040), .B(n1025), .Z(n1071) );
  XOR U4097 ( .A(n1080), .B(n1071), .Z(n1063) );
  XNOR U4098 ( .A(n1037), .B(n1063), .Z(z[32]) );
  ANDN U4099 ( .B(n1027), .A(n1026), .Z(n1036) );
  NANDN U4100 ( .A(n1029), .B(n1028), .Z(n1047) );
  NANDN U4101 ( .A(n1031), .B(n1030), .Z(n1032) );
  XNOR U4102 ( .A(n1047), .B(n1032), .Z(n1075) );
  NANDN U4103 ( .A(n1034), .B(n1033), .Z(n1041) );
  XNOR U4104 ( .A(n1075), .B(n1041), .Z(n1035) );
  XOR U4105 ( .A(n1036), .B(n1035), .Z(n1061) );
  XOR U4106 ( .A(n1061), .B(n1037), .Z(n1079) );
  ANDN U4107 ( .B(n1072), .A(n1038), .Z(n1043) );
  NAND U4108 ( .A(n1064), .B(n1066), .Z(n1039) );
  XNOR U4109 ( .A(n1040), .B(n1039), .Z(n1051) );
  XNOR U4110 ( .A(n1041), .B(n1051), .Z(n1042) );
  XNOR U4111 ( .A(n1043), .B(n1042), .Z(n1050) );
  NAND U4112 ( .A(n1045), .B(n1044), .Z(n1046) );
  XNOR U4113 ( .A(n1047), .B(n1046), .Z(n1057) );
  XNOR U4114 ( .A(n1048), .B(n1057), .Z(n1049) );
  XOR U4115 ( .A(n1050), .B(n1049), .Z(n1060) );
  XNOR U4116 ( .A(n1079), .B(n1060), .Z(z[33]) );
  XNOR U4117 ( .A(n1052), .B(n1051), .Z(z[34]) );
  AND U4118 ( .A(n1054), .B(n1053), .Z(n1059) );
  NANDN U4119 ( .A(n1056), .B(n1055), .Z(n1069) );
  XNOR U4120 ( .A(n1057), .B(n1069), .Z(n1058) );
  XOR U4121 ( .A(n1059), .B(n1058), .Z(n1078) );
  XOR U4122 ( .A(n1061), .B(n1060), .Z(n1062) );
  XOR U4123 ( .A(n1078), .B(n1062), .Z(z[35]) );
  XOR U4124 ( .A(n1063), .B(z[34]), .Z(z[36]) );
  XNOR U4125 ( .A(n1065), .B(n1064), .Z(n1067) );
  NAND U4126 ( .A(n1067), .B(n1066), .Z(n1068) );
  XOR U4127 ( .A(n1069), .B(n1068), .Z(n1070) );
  XNOR U4128 ( .A(n1071), .B(n1070), .Z(n1077) );
  NAND U4129 ( .A(n1072), .B(x[32]), .Z(n1073) );
  XNOR U4130 ( .A(n1074), .B(n1073), .Z(n1081) );
  XNOR U4131 ( .A(n1075), .B(n1081), .Z(n1076) );
  XOR U4132 ( .A(n1077), .B(n1076), .Z(z[37]) );
  XNOR U4133 ( .A(n1079), .B(n1078), .Z(z[38]) );
  XNOR U4134 ( .A(n1081), .B(n1080), .Z(n1082) );
  XNOR U4135 ( .A(z[33]), .B(n1082), .Z(z[39]) );
  AND U4136 ( .A(n1084), .B(n1083), .Z(n1089) );
  NANDN U4137 ( .A(n1086), .B(n1085), .Z(n1451) );
  XNOR U4138 ( .A(n1087), .B(n1451), .Z(n1088) );
  XOR U4139 ( .A(n1089), .B(n1088), .Z(n1599) );
  XOR U4140 ( .A(n1091), .B(n1090), .Z(n1092) );
  XOR U4141 ( .A(n1599), .B(n1092), .Z(z[3]) );
  IV U4142 ( .A(x[41]), .Z(n1199) );
  XOR U4143 ( .A(x[40]), .B(x[46]), .Z(n1094) );
  XOR U4144 ( .A(x[45]), .B(n1094), .Z(n1198) );
  IV U4145 ( .A(n1198), .Z(n1095) );
  AND U4146 ( .A(n1199), .B(n1095), .Z(n1102) );
  XNOR U4147 ( .A(x[43]), .B(n1199), .Z(n1098) );
  XNOR U4148 ( .A(x[42]), .B(n1098), .Z(n1093) );
  XNOR U4149 ( .A(n1094), .B(n1093), .Z(n1158) );
  IV U4150 ( .A(n1158), .Z(n1104) );
  XNOR U4151 ( .A(n1104), .B(n1198), .Z(n1157) );
  IV U4152 ( .A(x[47]), .Z(n1096) );
  XNOR U4153 ( .A(x[41]), .B(n1096), .Z(n1189) );
  NAND U4154 ( .A(n1157), .B(n1189), .Z(n1107) );
  XNOR U4155 ( .A(n1096), .B(n1095), .Z(n1103) );
  IV U4156 ( .A(n1103), .Z(n1187) );
  XOR U4157 ( .A(n1158), .B(n1187), .Z(n1123) );
  XNOR U4158 ( .A(n1107), .B(n1123), .Z(n1100) );
  XOR U4159 ( .A(x[40]), .B(n1104), .Z(n1133) );
  XOR U4160 ( .A(x[44]), .B(n1096), .Z(n1097) );
  IV U4161 ( .A(n1097), .Z(n1162) );
  NANDN U4162 ( .A(n1133), .B(n1162), .Z(n1106) );
  XNOR U4163 ( .A(n1098), .B(n1097), .Z(n1151) );
  XNOR U4164 ( .A(n1157), .B(n1151), .Z(n1149) );
  XOR U4165 ( .A(x[42]), .B(x[44]), .Z(n1164) );
  NANDN U4166 ( .A(n1149), .B(n1164), .Z(n1099) );
  XOR U4167 ( .A(n1106), .B(n1099), .Z(n1125) );
  XNOR U4168 ( .A(n1100), .B(n1125), .Z(n1101) );
  XOR U4169 ( .A(n1102), .B(n1101), .Z(n1138) );
  IV U4170 ( .A(n1138), .Z(n1144) );
  AND U4171 ( .A(n1104), .B(n1103), .Z(n1109) );
  XOR U4172 ( .A(x[40]), .B(n1151), .Z(n1152) );
  XNOR U4173 ( .A(n1198), .B(n1152), .Z(n1154) );
  XOR U4174 ( .A(x[42]), .B(x[47]), .Z(n1179) );
  NANDN U4175 ( .A(n1154), .B(n1179), .Z(n1105) );
  XNOR U4176 ( .A(n1106), .B(n1105), .Z(n1114) );
  XNOR U4177 ( .A(n1107), .B(n1114), .Z(n1108) );
  XOR U4178 ( .A(n1109), .B(n1108), .Z(n1134) );
  XNOR U4179 ( .A(x[44]), .B(n1198), .Z(n1172) );
  ANDN U4180 ( .B(x[40]), .A(n1172), .Z(n1116) );
  XOR U4181 ( .A(x[42]), .B(x[41]), .Z(n1110) );
  XOR U4182 ( .A(n1187), .B(n1110), .Z(n1161) );
  XOR U4183 ( .A(n1162), .B(n1110), .Z(n1167) );
  NAND U4184 ( .A(n1151), .B(n1167), .Z(n1118) );
  XNOR U4185 ( .A(n1161), .B(n1118), .Z(n1112) );
  XNOR U4186 ( .A(x[41]), .B(n1152), .Z(n1111) );
  XNOR U4187 ( .A(n1112), .B(n1111), .Z(n1113) );
  XOR U4188 ( .A(n1114), .B(n1113), .Z(n1115) );
  XOR U4189 ( .A(n1116), .B(n1115), .Z(n1136) );
  NAND U4190 ( .A(n1134), .B(n1136), .Z(n1117) );
  NAND U4191 ( .A(n1144), .B(n1117), .Z(n1128) );
  IV U4192 ( .A(n1134), .Z(n1135) );
  IV U4193 ( .A(n1136), .Z(n1142) );
  XOR U4194 ( .A(n1118), .B(n1172), .Z(n1121) );
  AND U4195 ( .A(n1161), .B(n1152), .Z(n1119) );
  XNOR U4196 ( .A(x[40]), .B(n1119), .Z(n1120) );
  XNOR U4197 ( .A(n1121), .B(n1120), .Z(n1122) );
  XNOR U4198 ( .A(n1123), .B(n1122), .Z(n1124) );
  XNOR U4199 ( .A(n1125), .B(n1124), .Z(n1146) );
  IV U4200 ( .A(n1146), .Z(n1141) );
  XOR U4201 ( .A(n1142), .B(n1141), .Z(n1126) );
  NAND U4202 ( .A(n1135), .B(n1126), .Z(n1127) );
  AND U4203 ( .A(n1128), .B(n1127), .Z(n1206) );
  NAND U4204 ( .A(n1142), .B(n1135), .Z(n1129) );
  NAND U4205 ( .A(n1141), .B(n1129), .Z(n1132) );
  XOR U4206 ( .A(n1135), .B(n1138), .Z(n1130) );
  NAND U4207 ( .A(n1136), .B(n1130), .Z(n1131) );
  AND U4208 ( .A(n1132), .B(n1131), .Z(n1188) );
  XNOR U4209 ( .A(n1206), .B(n1188), .Z(n1163) );
  OR U4210 ( .A(n1163), .B(n1133), .Z(n1156) );
  NAND U4211 ( .A(n1144), .B(n1134), .Z(n1140) );
  AND U4212 ( .A(n1136), .B(n1135), .Z(n1143) );
  XNOR U4213 ( .A(n1141), .B(n1143), .Z(n1137) );
  NAND U4214 ( .A(n1138), .B(n1137), .Z(n1139) );
  AND U4215 ( .A(n1140), .B(n1139), .Z(n1160) );
  NAND U4216 ( .A(n1142), .B(n1141), .Z(n1148) );
  XNOR U4217 ( .A(n1144), .B(n1143), .Z(n1145) );
  NAND U4218 ( .A(n1146), .B(n1145), .Z(n1147) );
  NAND U4219 ( .A(n1148), .B(n1147), .Z(n1200) );
  XNOR U4220 ( .A(n1160), .B(n1200), .Z(n1178) );
  XOR U4221 ( .A(n1178), .B(n1163), .Z(n1165) );
  OR U4222 ( .A(n1165), .B(n1149), .Z(n1150) );
  XNOR U4223 ( .A(n1156), .B(n1150), .Z(n1182) );
  XOR U4224 ( .A(n1160), .B(n1206), .Z(n1168) );
  NANDN U4225 ( .A(n1168), .B(n1151), .Z(n1208) );
  NANDN U4226 ( .A(n1160), .B(n1152), .Z(n1153) );
  XNOR U4227 ( .A(n1208), .B(n1153), .Z(n1186) );
  XOR U4228 ( .A(n1182), .B(n1186), .Z(n1171) );
  NANDN U4229 ( .A(n1154), .B(n1178), .Z(n1155) );
  XNOR U4230 ( .A(n1156), .B(n1155), .Z(n1214) );
  XNOR U4231 ( .A(n1200), .B(n1188), .Z(n1190) );
  NANDN U4232 ( .A(n1190), .B(n1157), .Z(n1174) );
  NAND U4233 ( .A(n1158), .B(n1188), .Z(n1159) );
  XNOR U4234 ( .A(n1174), .B(n1159), .Z(n1205) );
  XOR U4235 ( .A(n1214), .B(n1205), .Z(n1197) );
  XNOR U4236 ( .A(n1171), .B(n1197), .Z(z[40]) );
  ANDN U4237 ( .B(n1161), .A(n1160), .Z(n1170) );
  NANDN U4238 ( .A(n1163), .B(n1162), .Z(n1181) );
  NANDN U4239 ( .A(n1165), .B(n1164), .Z(n1166) );
  XNOR U4240 ( .A(n1181), .B(n1166), .Z(n1209) );
  NANDN U4241 ( .A(n1168), .B(n1167), .Z(n1175) );
  XNOR U4242 ( .A(n1209), .B(n1175), .Z(n1169) );
  XOR U4243 ( .A(n1170), .B(n1169), .Z(n1195) );
  XOR U4244 ( .A(n1195), .B(n1171), .Z(n1213) );
  ANDN U4245 ( .B(n1206), .A(n1172), .Z(n1177) );
  NAND U4246 ( .A(n1198), .B(n1200), .Z(n1173) );
  XNOR U4247 ( .A(n1174), .B(n1173), .Z(n1185) );
  XNOR U4248 ( .A(n1175), .B(n1185), .Z(n1176) );
  XNOR U4249 ( .A(n1177), .B(n1176), .Z(n1184) );
  NAND U4250 ( .A(n1179), .B(n1178), .Z(n1180) );
  XNOR U4251 ( .A(n1181), .B(n1180), .Z(n1191) );
  XNOR U4252 ( .A(n1182), .B(n1191), .Z(n1183) );
  XOR U4253 ( .A(n1184), .B(n1183), .Z(n1194) );
  XNOR U4254 ( .A(n1213), .B(n1194), .Z(z[41]) );
  XNOR U4255 ( .A(n1186), .B(n1185), .Z(z[42]) );
  AND U4256 ( .A(n1188), .B(n1187), .Z(n1193) );
  NANDN U4257 ( .A(n1190), .B(n1189), .Z(n1203) );
  XNOR U4258 ( .A(n1191), .B(n1203), .Z(n1192) );
  XOR U4259 ( .A(n1193), .B(n1192), .Z(n1212) );
  XOR U4260 ( .A(n1195), .B(n1194), .Z(n1196) );
  XOR U4261 ( .A(n1212), .B(n1196), .Z(z[43]) );
  XOR U4262 ( .A(n1197), .B(z[42]), .Z(z[44]) );
  XNOR U4263 ( .A(n1199), .B(n1198), .Z(n1201) );
  NAND U4264 ( .A(n1201), .B(n1200), .Z(n1202) );
  XOR U4265 ( .A(n1203), .B(n1202), .Z(n1204) );
  XNOR U4266 ( .A(n1205), .B(n1204), .Z(n1211) );
  NAND U4267 ( .A(n1206), .B(x[40]), .Z(n1207) );
  XNOR U4268 ( .A(n1208), .B(n1207), .Z(n1215) );
  XNOR U4269 ( .A(n1209), .B(n1215), .Z(n1210) );
  XOR U4270 ( .A(n1211), .B(n1210), .Z(z[45]) );
  XNOR U4271 ( .A(n1213), .B(n1212), .Z(z[46]) );
  XNOR U4272 ( .A(n1215), .B(n1214), .Z(n1216) );
  XNOR U4273 ( .A(z[41]), .B(n1216), .Z(z[47]) );
  IV U4274 ( .A(x[49]), .Z(n1324) );
  XOR U4275 ( .A(x[48]), .B(x[54]), .Z(n1218) );
  IV U4276 ( .A(n1323), .Z(n1219) );
  AND U4277 ( .A(n1324), .B(n1219), .Z(n1226) );
  XNOR U4278 ( .A(x[50]), .B(n1222), .Z(n1217) );
  XNOR U4279 ( .A(n1218), .B(n1217), .Z(n1282) );
  IV U4280 ( .A(n1282), .Z(n1228) );
  XNOR U4281 ( .A(n1228), .B(n1323), .Z(n1281) );
  IV U4282 ( .A(x[55]), .Z(n1220) );
  XNOR U4283 ( .A(x[49]), .B(n1220), .Z(n1314) );
  NAND U4284 ( .A(n1281), .B(n1314), .Z(n1231) );
  XNOR U4285 ( .A(n1220), .B(n1219), .Z(n1227) );
  IV U4286 ( .A(n1227), .Z(n1312) );
  XOR U4287 ( .A(n1282), .B(n1312), .Z(n1247) );
  XNOR U4288 ( .A(n1231), .B(n1247), .Z(n1224) );
  XOR U4289 ( .A(x[48]), .B(n1228), .Z(n1257) );
  XOR U4290 ( .A(x[52]), .B(n1220), .Z(n1221) );
  IV U4291 ( .A(n1221), .Z(n1286) );
  NANDN U4292 ( .A(n1257), .B(n1286), .Z(n1230) );
  XNOR U4293 ( .A(n1222), .B(n1221), .Z(n1275) );
  XNOR U4294 ( .A(n1281), .B(n1275), .Z(n1273) );
  XOR U4295 ( .A(x[50]), .B(x[52]), .Z(n1288) );
  NANDN U4296 ( .A(n1273), .B(n1288), .Z(n1223) );
  XOR U4297 ( .A(n1230), .B(n1223), .Z(n1249) );
  XNOR U4298 ( .A(n1224), .B(n1249), .Z(n1225) );
  XOR U4299 ( .A(n1226), .B(n1225), .Z(n1262) );
  IV U4300 ( .A(n1262), .Z(n1268) );
  AND U4301 ( .A(n1228), .B(n1227), .Z(n1233) );
  XOR U4302 ( .A(x[48]), .B(n1275), .Z(n1276) );
  XNOR U4303 ( .A(n1323), .B(n1276), .Z(n1278) );
  XOR U4304 ( .A(x[50]), .B(x[55]), .Z(n1303) );
  NANDN U4305 ( .A(n1278), .B(n1303), .Z(n1229) );
  XNOR U4306 ( .A(n1230), .B(n1229), .Z(n1238) );
  XNOR U4307 ( .A(n1231), .B(n1238), .Z(n1232) );
  XOR U4308 ( .A(n1233), .B(n1232), .Z(n1258) );
  XNOR U4309 ( .A(x[52]), .B(n1323), .Z(n1296) );
  ANDN U4310 ( .B(x[48]), .A(n1296), .Z(n1240) );
  XOR U4311 ( .A(x[50]), .B(x[49]), .Z(n1234) );
  XOR U4312 ( .A(n1312), .B(n1234), .Z(n1285) );
  XOR U4313 ( .A(n1286), .B(n1234), .Z(n1291) );
  NAND U4314 ( .A(n1275), .B(n1291), .Z(n1242) );
  XNOR U4315 ( .A(n1285), .B(n1242), .Z(n1236) );
  XNOR U4316 ( .A(x[49]), .B(n1276), .Z(n1235) );
  XNOR U4317 ( .A(n1236), .B(n1235), .Z(n1237) );
  XOR U4318 ( .A(n1238), .B(n1237), .Z(n1239) );
  XOR U4319 ( .A(n1240), .B(n1239), .Z(n1260) );
  NAND U4320 ( .A(n1258), .B(n1260), .Z(n1241) );
  NAND U4321 ( .A(n1268), .B(n1241), .Z(n1252) );
  IV U4322 ( .A(n1258), .Z(n1259) );
  IV U4323 ( .A(n1260), .Z(n1266) );
  XOR U4324 ( .A(n1242), .B(n1296), .Z(n1245) );
  AND U4325 ( .A(n1285), .B(n1276), .Z(n1243) );
  XNOR U4326 ( .A(x[48]), .B(n1243), .Z(n1244) );
  XNOR U4327 ( .A(n1245), .B(n1244), .Z(n1246) );
  XNOR U4328 ( .A(n1247), .B(n1246), .Z(n1248) );
  XNOR U4329 ( .A(n1249), .B(n1248), .Z(n1270) );
  IV U4330 ( .A(n1270), .Z(n1265) );
  XOR U4331 ( .A(n1266), .B(n1265), .Z(n1250) );
  NAND U4332 ( .A(n1259), .B(n1250), .Z(n1251) );
  AND U4333 ( .A(n1252), .B(n1251), .Z(n1331) );
  NAND U4334 ( .A(n1266), .B(n1259), .Z(n1253) );
  NAND U4335 ( .A(n1265), .B(n1253), .Z(n1256) );
  XOR U4336 ( .A(n1259), .B(n1262), .Z(n1254) );
  NAND U4337 ( .A(n1260), .B(n1254), .Z(n1255) );
  AND U4338 ( .A(n1256), .B(n1255), .Z(n1313) );
  XNOR U4339 ( .A(n1331), .B(n1313), .Z(n1287) );
  OR U4340 ( .A(n1287), .B(n1257), .Z(n1280) );
  NAND U4341 ( .A(n1268), .B(n1258), .Z(n1264) );
  AND U4342 ( .A(n1260), .B(n1259), .Z(n1267) );
  XNOR U4343 ( .A(n1265), .B(n1267), .Z(n1261) );
  NAND U4344 ( .A(n1262), .B(n1261), .Z(n1263) );
  AND U4345 ( .A(n1264), .B(n1263), .Z(n1284) );
  NAND U4346 ( .A(n1266), .B(n1265), .Z(n1272) );
  XNOR U4347 ( .A(n1268), .B(n1267), .Z(n1269) );
  NAND U4348 ( .A(n1270), .B(n1269), .Z(n1271) );
  NAND U4349 ( .A(n1272), .B(n1271), .Z(n1325) );
  XNOR U4350 ( .A(n1284), .B(n1325), .Z(n1302) );
  XOR U4351 ( .A(n1302), .B(n1287), .Z(n1289) );
  OR U4352 ( .A(n1289), .B(n1273), .Z(n1274) );
  XNOR U4353 ( .A(n1280), .B(n1274), .Z(n1306) );
  XOR U4354 ( .A(n1284), .B(n1331), .Z(n1292) );
  NANDN U4355 ( .A(n1292), .B(n1275), .Z(n1333) );
  NANDN U4356 ( .A(n1284), .B(n1276), .Z(n1277) );
  XNOR U4357 ( .A(n1333), .B(n1277), .Z(n1311) );
  XOR U4358 ( .A(n1306), .B(n1311), .Z(n1295) );
  NANDN U4359 ( .A(n1278), .B(n1302), .Z(n1279) );
  XNOR U4360 ( .A(n1280), .B(n1279), .Z(n1339) );
  XNOR U4361 ( .A(n1325), .B(n1313), .Z(n1315) );
  NANDN U4362 ( .A(n1315), .B(n1281), .Z(n1298) );
  NAND U4363 ( .A(n1282), .B(n1313), .Z(n1283) );
  XNOR U4364 ( .A(n1298), .B(n1283), .Z(n1330) );
  XOR U4365 ( .A(n1339), .B(n1330), .Z(n1322) );
  XNOR U4366 ( .A(n1295), .B(n1322), .Z(z[48]) );
  ANDN U4367 ( .B(n1285), .A(n1284), .Z(n1294) );
  NANDN U4368 ( .A(n1287), .B(n1286), .Z(n1305) );
  NANDN U4369 ( .A(n1289), .B(n1288), .Z(n1290) );
  XNOR U4370 ( .A(n1305), .B(n1290), .Z(n1334) );
  NANDN U4371 ( .A(n1292), .B(n1291), .Z(n1299) );
  XNOR U4372 ( .A(n1334), .B(n1299), .Z(n1293) );
  XOR U4373 ( .A(n1294), .B(n1293), .Z(n1320) );
  XOR U4374 ( .A(n1320), .B(n1295), .Z(n1338) );
  ANDN U4375 ( .B(n1331), .A(n1296), .Z(n1301) );
  NAND U4376 ( .A(n1323), .B(n1325), .Z(n1297) );
  XNOR U4377 ( .A(n1298), .B(n1297), .Z(n1310) );
  XNOR U4378 ( .A(n1299), .B(n1310), .Z(n1300) );
  XNOR U4379 ( .A(n1301), .B(n1300), .Z(n1308) );
  NAND U4380 ( .A(n1303), .B(n1302), .Z(n1304) );
  XNOR U4381 ( .A(n1305), .B(n1304), .Z(n1316) );
  XNOR U4382 ( .A(n1306), .B(n1316), .Z(n1307) );
  XOR U4383 ( .A(n1308), .B(n1307), .Z(n1319) );
  XNOR U4384 ( .A(n1338), .B(n1319), .Z(z[49]) );
  XOR U4385 ( .A(n1309), .B(z[2]), .Z(z[4]) );
  XNOR U4386 ( .A(n1311), .B(n1310), .Z(z[50]) );
  AND U4387 ( .A(n1313), .B(n1312), .Z(n1318) );
  NANDN U4388 ( .A(n1315), .B(n1314), .Z(n1328) );
  XNOR U4389 ( .A(n1316), .B(n1328), .Z(n1317) );
  XOR U4390 ( .A(n1318), .B(n1317), .Z(n1337) );
  XOR U4391 ( .A(n1320), .B(n1319), .Z(n1321) );
  XOR U4392 ( .A(n1337), .B(n1321), .Z(z[51]) );
  XOR U4393 ( .A(n1322), .B(z[50]), .Z(z[52]) );
  XNOR U4394 ( .A(n1324), .B(n1323), .Z(n1326) );
  NAND U4395 ( .A(n1326), .B(n1325), .Z(n1327) );
  XOR U4396 ( .A(n1328), .B(n1327), .Z(n1329) );
  XNOR U4397 ( .A(n1330), .B(n1329), .Z(n1336) );
  NAND U4398 ( .A(n1331), .B(x[48]), .Z(n1332) );
  XNOR U4399 ( .A(n1333), .B(n1332), .Z(n1340) );
  XNOR U4400 ( .A(n1334), .B(n1340), .Z(n1335) );
  XOR U4401 ( .A(n1336), .B(n1335), .Z(z[53]) );
  XNOR U4402 ( .A(n1338), .B(n1337), .Z(z[54]) );
  XNOR U4403 ( .A(n1340), .B(n1339), .Z(n1341) );
  XNOR U4404 ( .A(z[49]), .B(n1341), .Z(z[55]) );
  IV U4405 ( .A(x[57]), .Z(n1462) );
  XOR U4406 ( .A(x[56]), .B(x[62]), .Z(n1343) );
  XOR U4407 ( .A(x[61]), .B(n1343), .Z(n1461) );
  IV U4408 ( .A(n1461), .Z(n1344) );
  AND U4409 ( .A(n1462), .B(n1344), .Z(n1351) );
  XNOR U4410 ( .A(x[59]), .B(n1462), .Z(n1347) );
  XNOR U4411 ( .A(x[58]), .B(n1347), .Z(n1342) );
  XNOR U4412 ( .A(n1343), .B(n1342), .Z(n1407) );
  IV U4413 ( .A(n1407), .Z(n1353) );
  XNOR U4414 ( .A(n1353), .B(n1461), .Z(n1406) );
  IV U4415 ( .A(x[63]), .Z(n1345) );
  XNOR U4416 ( .A(x[57]), .B(n1345), .Z(n1438) );
  NAND U4417 ( .A(n1406), .B(n1438), .Z(n1356) );
  XNOR U4418 ( .A(n1345), .B(n1344), .Z(n1352) );
  IV U4419 ( .A(n1352), .Z(n1436) );
  XOR U4420 ( .A(n1407), .B(n1436), .Z(n1372) );
  XNOR U4421 ( .A(n1356), .B(n1372), .Z(n1349) );
  XOR U4422 ( .A(x[56]), .B(n1353), .Z(n1382) );
  XOR U4423 ( .A(x[60]), .B(n1345), .Z(n1346) );
  IV U4424 ( .A(n1346), .Z(n1411) );
  NANDN U4425 ( .A(n1382), .B(n1411), .Z(n1355) );
  XNOR U4426 ( .A(n1347), .B(n1346), .Z(n1400) );
  XNOR U4427 ( .A(n1406), .B(n1400), .Z(n1398) );
  XOR U4428 ( .A(x[58]), .B(x[60]), .Z(n1413) );
  NANDN U4429 ( .A(n1398), .B(n1413), .Z(n1348) );
  XOR U4430 ( .A(n1355), .B(n1348), .Z(n1374) );
  XNOR U4431 ( .A(n1349), .B(n1374), .Z(n1350) );
  XOR U4432 ( .A(n1351), .B(n1350), .Z(n1387) );
  IV U4433 ( .A(n1387), .Z(n1393) );
  AND U4434 ( .A(n1353), .B(n1352), .Z(n1358) );
  XOR U4435 ( .A(x[56]), .B(n1400), .Z(n1401) );
  XNOR U4436 ( .A(n1461), .B(n1401), .Z(n1403) );
  XOR U4437 ( .A(x[58]), .B(x[63]), .Z(n1428) );
  NANDN U4438 ( .A(n1403), .B(n1428), .Z(n1354) );
  XNOR U4439 ( .A(n1355), .B(n1354), .Z(n1363) );
  XNOR U4440 ( .A(n1356), .B(n1363), .Z(n1357) );
  XOR U4441 ( .A(n1358), .B(n1357), .Z(n1383) );
  XNOR U4442 ( .A(x[60]), .B(n1461), .Z(n1421) );
  ANDN U4443 ( .B(x[56]), .A(n1421), .Z(n1365) );
  XOR U4444 ( .A(x[58]), .B(x[57]), .Z(n1359) );
  XOR U4445 ( .A(n1436), .B(n1359), .Z(n1410) );
  XOR U4446 ( .A(n1411), .B(n1359), .Z(n1416) );
  NAND U4447 ( .A(n1400), .B(n1416), .Z(n1367) );
  XNOR U4448 ( .A(n1410), .B(n1367), .Z(n1361) );
  XNOR U4449 ( .A(x[57]), .B(n1401), .Z(n1360) );
  XNOR U4450 ( .A(n1361), .B(n1360), .Z(n1362) );
  XOR U4451 ( .A(n1363), .B(n1362), .Z(n1364) );
  XOR U4452 ( .A(n1365), .B(n1364), .Z(n1385) );
  NAND U4453 ( .A(n1383), .B(n1385), .Z(n1366) );
  NAND U4454 ( .A(n1393), .B(n1366), .Z(n1377) );
  IV U4455 ( .A(n1383), .Z(n1384) );
  IV U4456 ( .A(n1385), .Z(n1391) );
  XOR U4457 ( .A(n1367), .B(n1421), .Z(n1370) );
  AND U4458 ( .A(n1410), .B(n1401), .Z(n1368) );
  XNOR U4459 ( .A(x[56]), .B(n1368), .Z(n1369) );
  XNOR U4460 ( .A(n1370), .B(n1369), .Z(n1371) );
  XNOR U4461 ( .A(n1372), .B(n1371), .Z(n1373) );
  XNOR U4462 ( .A(n1374), .B(n1373), .Z(n1395) );
  IV U4463 ( .A(n1395), .Z(n1390) );
  XOR U4464 ( .A(n1391), .B(n1390), .Z(n1375) );
  NAND U4465 ( .A(n1384), .B(n1375), .Z(n1376) );
  AND U4466 ( .A(n1377), .B(n1376), .Z(n1469) );
  NAND U4467 ( .A(n1391), .B(n1384), .Z(n1378) );
  NAND U4468 ( .A(n1390), .B(n1378), .Z(n1381) );
  XOR U4469 ( .A(n1384), .B(n1387), .Z(n1379) );
  NAND U4470 ( .A(n1385), .B(n1379), .Z(n1380) );
  AND U4471 ( .A(n1381), .B(n1380), .Z(n1437) );
  XNOR U4472 ( .A(n1469), .B(n1437), .Z(n1412) );
  OR U4473 ( .A(n1412), .B(n1382), .Z(n1405) );
  NAND U4474 ( .A(n1393), .B(n1383), .Z(n1389) );
  AND U4475 ( .A(n1385), .B(n1384), .Z(n1392) );
  XNOR U4476 ( .A(n1390), .B(n1392), .Z(n1386) );
  NAND U4477 ( .A(n1387), .B(n1386), .Z(n1388) );
  AND U4478 ( .A(n1389), .B(n1388), .Z(n1409) );
  NAND U4479 ( .A(n1391), .B(n1390), .Z(n1397) );
  XNOR U4480 ( .A(n1393), .B(n1392), .Z(n1394) );
  NAND U4481 ( .A(n1395), .B(n1394), .Z(n1396) );
  NAND U4482 ( .A(n1397), .B(n1396), .Z(n1463) );
  XNOR U4483 ( .A(n1409), .B(n1463), .Z(n1427) );
  XOR U4484 ( .A(n1427), .B(n1412), .Z(n1414) );
  OR U4485 ( .A(n1414), .B(n1398), .Z(n1399) );
  XNOR U4486 ( .A(n1405), .B(n1399), .Z(n1431) );
  XOR U4487 ( .A(n1409), .B(n1469), .Z(n1417) );
  NANDN U4488 ( .A(n1417), .B(n1400), .Z(n1471) );
  NANDN U4489 ( .A(n1409), .B(n1401), .Z(n1402) );
  XNOR U4490 ( .A(n1471), .B(n1402), .Z(n1435) );
  XOR U4491 ( .A(n1431), .B(n1435), .Z(n1420) );
  NANDN U4492 ( .A(n1403), .B(n1427), .Z(n1404) );
  XNOR U4493 ( .A(n1405), .B(n1404), .Z(n1477) );
  XNOR U4494 ( .A(n1463), .B(n1437), .Z(n1439) );
  NANDN U4495 ( .A(n1439), .B(n1406), .Z(n1423) );
  NAND U4496 ( .A(n1407), .B(n1437), .Z(n1408) );
  XNOR U4497 ( .A(n1423), .B(n1408), .Z(n1468) );
  XOR U4498 ( .A(n1477), .B(n1468), .Z(n1460) );
  XNOR U4499 ( .A(n1420), .B(n1460), .Z(z[56]) );
  ANDN U4500 ( .B(n1410), .A(n1409), .Z(n1419) );
  NANDN U4501 ( .A(n1412), .B(n1411), .Z(n1430) );
  NANDN U4502 ( .A(n1414), .B(n1413), .Z(n1415) );
  XNOR U4503 ( .A(n1430), .B(n1415), .Z(n1472) );
  NANDN U4504 ( .A(n1417), .B(n1416), .Z(n1424) );
  XNOR U4505 ( .A(n1472), .B(n1424), .Z(n1418) );
  XOR U4506 ( .A(n1419), .B(n1418), .Z(n1444) );
  XOR U4507 ( .A(n1444), .B(n1420), .Z(n1476) );
  ANDN U4508 ( .B(n1469), .A(n1421), .Z(n1426) );
  NAND U4509 ( .A(n1461), .B(n1463), .Z(n1422) );
  XNOR U4510 ( .A(n1423), .B(n1422), .Z(n1434) );
  XNOR U4511 ( .A(n1424), .B(n1434), .Z(n1425) );
  XNOR U4512 ( .A(n1426), .B(n1425), .Z(n1433) );
  NAND U4513 ( .A(n1428), .B(n1427), .Z(n1429) );
  XNOR U4514 ( .A(n1430), .B(n1429), .Z(n1440) );
  XNOR U4515 ( .A(n1431), .B(n1440), .Z(n1432) );
  XOR U4516 ( .A(n1433), .B(n1432), .Z(n1443) );
  XNOR U4517 ( .A(n1476), .B(n1443), .Z(z[57]) );
  XNOR U4518 ( .A(n1435), .B(n1434), .Z(z[58]) );
  AND U4519 ( .A(n1437), .B(n1436), .Z(n1442) );
  NANDN U4520 ( .A(n1439), .B(n1438), .Z(n1466) );
  XNOR U4521 ( .A(n1440), .B(n1466), .Z(n1441) );
  XOR U4522 ( .A(n1442), .B(n1441), .Z(n1475) );
  XOR U4523 ( .A(n1444), .B(n1443), .Z(n1445) );
  XOR U4524 ( .A(n1475), .B(n1445), .Z(z[59]) );
  XNOR U4525 ( .A(n1447), .B(n1446), .Z(n1449) );
  NAND U4526 ( .A(n1449), .B(n1448), .Z(n1450) );
  XOR U4527 ( .A(n1451), .B(n1450), .Z(n1452) );
  XNOR U4528 ( .A(n1453), .B(n1452), .Z(n1459) );
  NAND U4529 ( .A(n1454), .B(x[0]), .Z(n1455) );
  XNOR U4530 ( .A(n1456), .B(n1455), .Z(n1731) );
  XNOR U4531 ( .A(n1457), .B(n1731), .Z(n1458) );
  XOR U4532 ( .A(n1459), .B(n1458), .Z(z[5]) );
  XOR U4533 ( .A(n1460), .B(z[58]), .Z(z[60]) );
  XNOR U4534 ( .A(n1462), .B(n1461), .Z(n1464) );
  NAND U4535 ( .A(n1464), .B(n1463), .Z(n1465) );
  XOR U4536 ( .A(n1466), .B(n1465), .Z(n1467) );
  XNOR U4537 ( .A(n1468), .B(n1467), .Z(n1474) );
  NAND U4538 ( .A(n1469), .B(x[56]), .Z(n1470) );
  XNOR U4539 ( .A(n1471), .B(n1470), .Z(n1478) );
  XNOR U4540 ( .A(n1472), .B(n1478), .Z(n1473) );
  XOR U4541 ( .A(n1474), .B(n1473), .Z(z[61]) );
  XNOR U4542 ( .A(n1476), .B(n1475), .Z(z[62]) );
  XNOR U4543 ( .A(n1478), .B(n1477), .Z(n1479) );
  XNOR U4544 ( .A(z[57]), .B(n1479), .Z(z[63]) );
  IV U4545 ( .A(x[65]), .Z(n1586) );
  XOR U4546 ( .A(x[64]), .B(x[70]), .Z(n1481) );
  XOR U4547 ( .A(x[69]), .B(n1481), .Z(n1585) );
  IV U4548 ( .A(n1585), .Z(n1482) );
  AND U4549 ( .A(n1586), .B(n1482), .Z(n1489) );
  XNOR U4550 ( .A(x[67]), .B(n1586), .Z(n1485) );
  XNOR U4551 ( .A(x[66]), .B(n1485), .Z(n1480) );
  XNOR U4552 ( .A(n1481), .B(n1480), .Z(n1545) );
  IV U4553 ( .A(n1545), .Z(n1491) );
  XNOR U4554 ( .A(n1491), .B(n1585), .Z(n1544) );
  IV U4555 ( .A(x[71]), .Z(n1483) );
  XNOR U4556 ( .A(x[65]), .B(n1483), .Z(n1576) );
  NAND U4557 ( .A(n1544), .B(n1576), .Z(n1494) );
  XNOR U4558 ( .A(n1483), .B(n1482), .Z(n1490) );
  IV U4559 ( .A(n1490), .Z(n1574) );
  XOR U4560 ( .A(n1545), .B(n1574), .Z(n1510) );
  XNOR U4561 ( .A(n1494), .B(n1510), .Z(n1487) );
  XOR U4562 ( .A(x[64]), .B(n1491), .Z(n1520) );
  XOR U4563 ( .A(x[68]), .B(n1483), .Z(n1484) );
  IV U4564 ( .A(n1484), .Z(n1549) );
  NANDN U4565 ( .A(n1520), .B(n1549), .Z(n1493) );
  XNOR U4566 ( .A(n1485), .B(n1484), .Z(n1538) );
  XNOR U4567 ( .A(n1544), .B(n1538), .Z(n1536) );
  XOR U4568 ( .A(x[66]), .B(x[68]), .Z(n1551) );
  NANDN U4569 ( .A(n1536), .B(n1551), .Z(n1486) );
  XOR U4570 ( .A(n1493), .B(n1486), .Z(n1512) );
  XNOR U4571 ( .A(n1487), .B(n1512), .Z(n1488) );
  XOR U4572 ( .A(n1489), .B(n1488), .Z(n1525) );
  IV U4573 ( .A(n1525), .Z(n1531) );
  AND U4574 ( .A(n1491), .B(n1490), .Z(n1496) );
  XOR U4575 ( .A(x[64]), .B(n1538), .Z(n1539) );
  XNOR U4576 ( .A(n1585), .B(n1539), .Z(n1541) );
  XOR U4577 ( .A(x[66]), .B(x[71]), .Z(n1566) );
  NANDN U4578 ( .A(n1541), .B(n1566), .Z(n1492) );
  XNOR U4579 ( .A(n1493), .B(n1492), .Z(n1501) );
  XNOR U4580 ( .A(n1494), .B(n1501), .Z(n1495) );
  XOR U4581 ( .A(n1496), .B(n1495), .Z(n1521) );
  XNOR U4582 ( .A(x[68]), .B(n1585), .Z(n1559) );
  ANDN U4583 ( .B(x[64]), .A(n1559), .Z(n1503) );
  XOR U4584 ( .A(x[66]), .B(x[65]), .Z(n1497) );
  XOR U4585 ( .A(n1574), .B(n1497), .Z(n1548) );
  XOR U4586 ( .A(n1549), .B(n1497), .Z(n1554) );
  NAND U4587 ( .A(n1538), .B(n1554), .Z(n1505) );
  XNOR U4588 ( .A(n1548), .B(n1505), .Z(n1499) );
  XNOR U4589 ( .A(x[65]), .B(n1539), .Z(n1498) );
  XNOR U4590 ( .A(n1499), .B(n1498), .Z(n1500) );
  XOR U4591 ( .A(n1501), .B(n1500), .Z(n1502) );
  XOR U4592 ( .A(n1503), .B(n1502), .Z(n1523) );
  NAND U4593 ( .A(n1521), .B(n1523), .Z(n1504) );
  NAND U4594 ( .A(n1531), .B(n1504), .Z(n1515) );
  IV U4595 ( .A(n1521), .Z(n1522) );
  IV U4596 ( .A(n1523), .Z(n1529) );
  XOR U4597 ( .A(n1505), .B(n1559), .Z(n1508) );
  AND U4598 ( .A(n1548), .B(n1539), .Z(n1506) );
  XNOR U4599 ( .A(x[64]), .B(n1506), .Z(n1507) );
  XNOR U4600 ( .A(n1508), .B(n1507), .Z(n1509) );
  XNOR U4601 ( .A(n1510), .B(n1509), .Z(n1511) );
  XNOR U4602 ( .A(n1512), .B(n1511), .Z(n1533) );
  IV U4603 ( .A(n1533), .Z(n1528) );
  XOR U4604 ( .A(n1529), .B(n1528), .Z(n1513) );
  NAND U4605 ( .A(n1522), .B(n1513), .Z(n1514) );
  AND U4606 ( .A(n1515), .B(n1514), .Z(n1593) );
  NAND U4607 ( .A(n1529), .B(n1522), .Z(n1516) );
  NAND U4608 ( .A(n1528), .B(n1516), .Z(n1519) );
  XOR U4609 ( .A(n1522), .B(n1525), .Z(n1517) );
  NAND U4610 ( .A(n1523), .B(n1517), .Z(n1518) );
  AND U4611 ( .A(n1519), .B(n1518), .Z(n1575) );
  XNOR U4612 ( .A(n1593), .B(n1575), .Z(n1550) );
  OR U4613 ( .A(n1550), .B(n1520), .Z(n1543) );
  NAND U4614 ( .A(n1531), .B(n1521), .Z(n1527) );
  AND U4615 ( .A(n1523), .B(n1522), .Z(n1530) );
  XNOR U4616 ( .A(n1528), .B(n1530), .Z(n1524) );
  NAND U4617 ( .A(n1525), .B(n1524), .Z(n1526) );
  AND U4618 ( .A(n1527), .B(n1526), .Z(n1547) );
  NAND U4619 ( .A(n1529), .B(n1528), .Z(n1535) );
  XNOR U4620 ( .A(n1531), .B(n1530), .Z(n1532) );
  NAND U4621 ( .A(n1533), .B(n1532), .Z(n1534) );
  NAND U4622 ( .A(n1535), .B(n1534), .Z(n1587) );
  XNOR U4623 ( .A(n1547), .B(n1587), .Z(n1565) );
  XOR U4624 ( .A(n1565), .B(n1550), .Z(n1552) );
  OR U4625 ( .A(n1552), .B(n1536), .Z(n1537) );
  XNOR U4626 ( .A(n1543), .B(n1537), .Z(n1569) );
  XOR U4627 ( .A(n1547), .B(n1593), .Z(n1555) );
  NANDN U4628 ( .A(n1555), .B(n1538), .Z(n1595) );
  NANDN U4629 ( .A(n1547), .B(n1539), .Z(n1540) );
  XNOR U4630 ( .A(n1595), .B(n1540), .Z(n1573) );
  XOR U4631 ( .A(n1569), .B(n1573), .Z(n1558) );
  NANDN U4632 ( .A(n1541), .B(n1565), .Z(n1542) );
  XNOR U4633 ( .A(n1543), .B(n1542), .Z(n1603) );
  XNOR U4634 ( .A(n1587), .B(n1575), .Z(n1577) );
  NANDN U4635 ( .A(n1577), .B(n1544), .Z(n1561) );
  NAND U4636 ( .A(n1545), .B(n1575), .Z(n1546) );
  XNOR U4637 ( .A(n1561), .B(n1546), .Z(n1592) );
  XOR U4638 ( .A(n1603), .B(n1592), .Z(n1584) );
  XNOR U4639 ( .A(n1558), .B(n1584), .Z(z[64]) );
  ANDN U4640 ( .B(n1548), .A(n1547), .Z(n1557) );
  NANDN U4641 ( .A(n1550), .B(n1549), .Z(n1568) );
  NANDN U4642 ( .A(n1552), .B(n1551), .Z(n1553) );
  XNOR U4643 ( .A(n1568), .B(n1553), .Z(n1596) );
  NANDN U4644 ( .A(n1555), .B(n1554), .Z(n1562) );
  XNOR U4645 ( .A(n1596), .B(n1562), .Z(n1556) );
  XOR U4646 ( .A(n1557), .B(n1556), .Z(n1582) );
  XOR U4647 ( .A(n1582), .B(n1558), .Z(n1602) );
  ANDN U4648 ( .B(n1593), .A(n1559), .Z(n1564) );
  NAND U4649 ( .A(n1585), .B(n1587), .Z(n1560) );
  XNOR U4650 ( .A(n1561), .B(n1560), .Z(n1572) );
  XNOR U4651 ( .A(n1562), .B(n1572), .Z(n1563) );
  XNOR U4652 ( .A(n1564), .B(n1563), .Z(n1571) );
  NAND U4653 ( .A(n1566), .B(n1565), .Z(n1567) );
  XNOR U4654 ( .A(n1568), .B(n1567), .Z(n1578) );
  XNOR U4655 ( .A(n1569), .B(n1578), .Z(n1570) );
  XOR U4656 ( .A(n1571), .B(n1570), .Z(n1581) );
  XNOR U4657 ( .A(n1602), .B(n1581), .Z(z[65]) );
  XNOR U4658 ( .A(n1573), .B(n1572), .Z(z[66]) );
  AND U4659 ( .A(n1575), .B(n1574), .Z(n1580) );
  NANDN U4660 ( .A(n1577), .B(n1576), .Z(n1590) );
  XNOR U4661 ( .A(n1578), .B(n1590), .Z(n1579) );
  XOR U4662 ( .A(n1580), .B(n1579), .Z(n1601) );
  XOR U4663 ( .A(n1582), .B(n1581), .Z(n1583) );
  XOR U4664 ( .A(n1601), .B(n1583), .Z(z[67]) );
  XOR U4665 ( .A(n1584), .B(z[66]), .Z(z[68]) );
  XNOR U4666 ( .A(n1586), .B(n1585), .Z(n1588) );
  NAND U4667 ( .A(n1588), .B(n1587), .Z(n1589) );
  XOR U4668 ( .A(n1590), .B(n1589), .Z(n1591) );
  XNOR U4669 ( .A(n1592), .B(n1591), .Z(n1598) );
  NAND U4670 ( .A(n1593), .B(x[64]), .Z(n1594) );
  XNOR U4671 ( .A(n1595), .B(n1594), .Z(n1604) );
  XNOR U4672 ( .A(n1596), .B(n1604), .Z(n1597) );
  XOR U4673 ( .A(n1598), .B(n1597), .Z(z[69]) );
  XNOR U4674 ( .A(n1600), .B(n1599), .Z(z[6]) );
  XNOR U4675 ( .A(n1602), .B(n1601), .Z(z[70]) );
  XNOR U4676 ( .A(n1604), .B(n1603), .Z(n1605) );
  XNOR U4677 ( .A(z[65]), .B(n1605), .Z(z[71]) );
  IV U4678 ( .A(x[73]), .Z(n1712) );
  XOR U4679 ( .A(x[72]), .B(x[78]), .Z(n1607) );
  XOR U4680 ( .A(x[77]), .B(n1607), .Z(n1711) );
  IV U4681 ( .A(n1711), .Z(n1608) );
  AND U4682 ( .A(n1712), .B(n1608), .Z(n1615) );
  XNOR U4683 ( .A(x[75]), .B(n1712), .Z(n1611) );
  XNOR U4684 ( .A(x[74]), .B(n1611), .Z(n1606) );
  XNOR U4685 ( .A(n1607), .B(n1606), .Z(n1671) );
  IV U4686 ( .A(n1671), .Z(n1617) );
  XNOR U4687 ( .A(n1617), .B(n1711), .Z(n1670) );
  IV U4688 ( .A(x[79]), .Z(n1609) );
  XNOR U4689 ( .A(x[73]), .B(n1609), .Z(n1702) );
  NAND U4690 ( .A(n1670), .B(n1702), .Z(n1620) );
  XNOR U4691 ( .A(n1609), .B(n1608), .Z(n1616) );
  IV U4692 ( .A(n1616), .Z(n1700) );
  XOR U4693 ( .A(n1671), .B(n1700), .Z(n1636) );
  XNOR U4694 ( .A(n1620), .B(n1636), .Z(n1613) );
  XOR U4695 ( .A(x[72]), .B(n1617), .Z(n1646) );
  XOR U4696 ( .A(x[76]), .B(n1609), .Z(n1610) );
  IV U4697 ( .A(n1610), .Z(n1675) );
  NANDN U4698 ( .A(n1646), .B(n1675), .Z(n1619) );
  XNOR U4699 ( .A(n1611), .B(n1610), .Z(n1664) );
  XNOR U4700 ( .A(n1670), .B(n1664), .Z(n1662) );
  XOR U4701 ( .A(x[74]), .B(x[76]), .Z(n1677) );
  NANDN U4702 ( .A(n1662), .B(n1677), .Z(n1612) );
  XOR U4703 ( .A(n1619), .B(n1612), .Z(n1638) );
  XNOR U4704 ( .A(n1613), .B(n1638), .Z(n1614) );
  XOR U4705 ( .A(n1615), .B(n1614), .Z(n1651) );
  IV U4706 ( .A(n1651), .Z(n1657) );
  AND U4707 ( .A(n1617), .B(n1616), .Z(n1622) );
  XOR U4708 ( .A(x[72]), .B(n1664), .Z(n1665) );
  XNOR U4709 ( .A(n1711), .B(n1665), .Z(n1667) );
  XOR U4710 ( .A(x[74]), .B(x[79]), .Z(n1692) );
  NANDN U4711 ( .A(n1667), .B(n1692), .Z(n1618) );
  XNOR U4712 ( .A(n1619), .B(n1618), .Z(n1627) );
  XNOR U4713 ( .A(n1620), .B(n1627), .Z(n1621) );
  XOR U4714 ( .A(n1622), .B(n1621), .Z(n1647) );
  XNOR U4715 ( .A(x[76]), .B(n1711), .Z(n1685) );
  ANDN U4716 ( .B(x[72]), .A(n1685), .Z(n1629) );
  XOR U4717 ( .A(x[74]), .B(x[73]), .Z(n1623) );
  XOR U4718 ( .A(n1700), .B(n1623), .Z(n1674) );
  XOR U4719 ( .A(n1675), .B(n1623), .Z(n1680) );
  NAND U4720 ( .A(n1664), .B(n1680), .Z(n1631) );
  XNOR U4721 ( .A(n1674), .B(n1631), .Z(n1625) );
  XNOR U4722 ( .A(x[73]), .B(n1665), .Z(n1624) );
  XNOR U4723 ( .A(n1625), .B(n1624), .Z(n1626) );
  XOR U4724 ( .A(n1627), .B(n1626), .Z(n1628) );
  XOR U4725 ( .A(n1629), .B(n1628), .Z(n1649) );
  NAND U4726 ( .A(n1647), .B(n1649), .Z(n1630) );
  NAND U4727 ( .A(n1657), .B(n1630), .Z(n1641) );
  IV U4728 ( .A(n1647), .Z(n1648) );
  IV U4729 ( .A(n1649), .Z(n1655) );
  XOR U4730 ( .A(n1631), .B(n1685), .Z(n1634) );
  AND U4731 ( .A(n1674), .B(n1665), .Z(n1632) );
  XNOR U4732 ( .A(x[72]), .B(n1632), .Z(n1633) );
  XNOR U4733 ( .A(n1634), .B(n1633), .Z(n1635) );
  XNOR U4734 ( .A(n1636), .B(n1635), .Z(n1637) );
  XNOR U4735 ( .A(n1638), .B(n1637), .Z(n1659) );
  IV U4736 ( .A(n1659), .Z(n1654) );
  XOR U4737 ( .A(n1655), .B(n1654), .Z(n1639) );
  NAND U4738 ( .A(n1648), .B(n1639), .Z(n1640) );
  AND U4739 ( .A(n1641), .B(n1640), .Z(n1719) );
  NAND U4740 ( .A(n1655), .B(n1648), .Z(n1642) );
  NAND U4741 ( .A(n1654), .B(n1642), .Z(n1645) );
  XOR U4742 ( .A(n1648), .B(n1651), .Z(n1643) );
  NAND U4743 ( .A(n1649), .B(n1643), .Z(n1644) );
  AND U4744 ( .A(n1645), .B(n1644), .Z(n1701) );
  XNOR U4745 ( .A(n1719), .B(n1701), .Z(n1676) );
  OR U4746 ( .A(n1676), .B(n1646), .Z(n1669) );
  NAND U4747 ( .A(n1657), .B(n1647), .Z(n1653) );
  AND U4748 ( .A(n1649), .B(n1648), .Z(n1656) );
  XNOR U4749 ( .A(n1654), .B(n1656), .Z(n1650) );
  NAND U4750 ( .A(n1651), .B(n1650), .Z(n1652) );
  AND U4751 ( .A(n1653), .B(n1652), .Z(n1673) );
  NAND U4752 ( .A(n1655), .B(n1654), .Z(n1661) );
  XNOR U4753 ( .A(n1657), .B(n1656), .Z(n1658) );
  NAND U4754 ( .A(n1659), .B(n1658), .Z(n1660) );
  NAND U4755 ( .A(n1661), .B(n1660), .Z(n1713) );
  XNOR U4756 ( .A(n1673), .B(n1713), .Z(n1691) );
  XOR U4757 ( .A(n1691), .B(n1676), .Z(n1678) );
  OR U4758 ( .A(n1678), .B(n1662), .Z(n1663) );
  XNOR U4759 ( .A(n1669), .B(n1663), .Z(n1695) );
  XOR U4760 ( .A(n1673), .B(n1719), .Z(n1681) );
  NANDN U4761 ( .A(n1681), .B(n1664), .Z(n1721) );
  NANDN U4762 ( .A(n1673), .B(n1665), .Z(n1666) );
  XNOR U4763 ( .A(n1721), .B(n1666), .Z(n1699) );
  XOR U4764 ( .A(n1695), .B(n1699), .Z(n1684) );
  NANDN U4765 ( .A(n1667), .B(n1691), .Z(n1668) );
  XNOR U4766 ( .A(n1669), .B(n1668), .Z(n1727) );
  XNOR U4767 ( .A(n1713), .B(n1701), .Z(n1703) );
  NANDN U4768 ( .A(n1703), .B(n1670), .Z(n1687) );
  NAND U4769 ( .A(n1671), .B(n1701), .Z(n1672) );
  XNOR U4770 ( .A(n1687), .B(n1672), .Z(n1718) );
  XOR U4771 ( .A(n1727), .B(n1718), .Z(n1710) );
  XNOR U4772 ( .A(n1684), .B(n1710), .Z(z[72]) );
  ANDN U4773 ( .B(n1674), .A(n1673), .Z(n1683) );
  NANDN U4774 ( .A(n1676), .B(n1675), .Z(n1694) );
  NANDN U4775 ( .A(n1678), .B(n1677), .Z(n1679) );
  XNOR U4776 ( .A(n1694), .B(n1679), .Z(n1722) );
  NANDN U4777 ( .A(n1681), .B(n1680), .Z(n1688) );
  XNOR U4778 ( .A(n1722), .B(n1688), .Z(n1682) );
  XOR U4779 ( .A(n1683), .B(n1682), .Z(n1708) );
  XOR U4780 ( .A(n1708), .B(n1684), .Z(n1726) );
  ANDN U4781 ( .B(n1719), .A(n1685), .Z(n1690) );
  NAND U4782 ( .A(n1711), .B(n1713), .Z(n1686) );
  XNOR U4783 ( .A(n1687), .B(n1686), .Z(n1698) );
  XNOR U4784 ( .A(n1688), .B(n1698), .Z(n1689) );
  XNOR U4785 ( .A(n1690), .B(n1689), .Z(n1697) );
  NAND U4786 ( .A(n1692), .B(n1691), .Z(n1693) );
  XNOR U4787 ( .A(n1694), .B(n1693), .Z(n1704) );
  XNOR U4788 ( .A(n1695), .B(n1704), .Z(n1696) );
  XOR U4789 ( .A(n1697), .B(n1696), .Z(n1707) );
  XNOR U4790 ( .A(n1726), .B(n1707), .Z(z[73]) );
  XNOR U4791 ( .A(n1699), .B(n1698), .Z(z[74]) );
  AND U4792 ( .A(n1701), .B(n1700), .Z(n1706) );
  NANDN U4793 ( .A(n1703), .B(n1702), .Z(n1716) );
  XNOR U4794 ( .A(n1704), .B(n1716), .Z(n1705) );
  XOR U4795 ( .A(n1706), .B(n1705), .Z(n1725) );
  XOR U4796 ( .A(n1708), .B(n1707), .Z(n1709) );
  XOR U4797 ( .A(n1725), .B(n1709), .Z(z[75]) );
  XOR U4798 ( .A(n1710), .B(z[74]), .Z(z[76]) );
  XNOR U4799 ( .A(n1712), .B(n1711), .Z(n1714) );
  NAND U4800 ( .A(n1714), .B(n1713), .Z(n1715) );
  XOR U4801 ( .A(n1716), .B(n1715), .Z(n1717) );
  XNOR U4802 ( .A(n1718), .B(n1717), .Z(n1724) );
  NAND U4803 ( .A(n1719), .B(x[72]), .Z(n1720) );
  XNOR U4804 ( .A(n1721), .B(n1720), .Z(n1728) );
  XNOR U4805 ( .A(n1722), .B(n1728), .Z(n1723) );
  XOR U4806 ( .A(n1724), .B(n1723), .Z(z[77]) );
  XNOR U4807 ( .A(n1726), .B(n1725), .Z(z[78]) );
  XNOR U4808 ( .A(n1728), .B(n1727), .Z(n1729) );
  XNOR U4809 ( .A(z[73]), .B(n1729), .Z(z[79]) );
  XNOR U4810 ( .A(n1731), .B(n1730), .Z(n1732) );
  XNOR U4811 ( .A(z[1]), .B(n1732), .Z(z[7]) );
  XOR U4812 ( .A(x[80]), .B(x[86]), .Z(n1733) );
  IV U4813 ( .A(n1838), .Z(n1735) );
  IV U4814 ( .A(x[81]), .Z(n1837) );
  NAND U4815 ( .A(n1735), .B(n1837), .Z(n1742) );
  XNOR U4816 ( .A(x[82]), .B(n1733), .Z(n1734) );
  XNOR U4817 ( .A(n1738), .B(n1734), .Z(n1797) );
  XNOR U4818 ( .A(n1735), .B(n1797), .Z(n1796) );
  IV U4819 ( .A(x[87]), .Z(n1736) );
  XNOR U4820 ( .A(x[81]), .B(n1736), .Z(n1828) );
  NAND U4821 ( .A(n1796), .B(n1828), .Z(n1745) );
  XNOR U4822 ( .A(n1735), .B(n1736), .Z(n1826) );
  XOR U4823 ( .A(n1797), .B(n1826), .Z(n1753) );
  XOR U4824 ( .A(n1745), .B(n1753), .Z(n1740) );
  XNOR U4825 ( .A(x[80]), .B(n1797), .Z(n1772) );
  XOR U4826 ( .A(x[84]), .B(n1736), .Z(n1737) );
  IV U4827 ( .A(n1737), .Z(n1801) );
  NANDN U4828 ( .A(n1772), .B(n1801), .Z(n1744) );
  XOR U4829 ( .A(n1738), .B(n1737), .Z(n1790) );
  XOR U4830 ( .A(n1796), .B(n1790), .Z(n1788) );
  XOR U4831 ( .A(x[82]), .B(x[84]), .Z(n1803) );
  NANDN U4832 ( .A(n1788), .B(n1803), .Z(n1739) );
  XNOR U4833 ( .A(n1744), .B(n1739), .Z(n1749) );
  XOR U4834 ( .A(n1740), .B(n1749), .Z(n1741) );
  XOR U4835 ( .A(n1742), .B(n1741), .Z(n1783) );
  IV U4836 ( .A(n1783), .Z(n1777) );
  ANDN U4837 ( .B(n1826), .A(n1797), .Z(n1747) );
  XNOR U4838 ( .A(x[80]), .B(n1790), .Z(n1791) );
  XNOR U4839 ( .A(n1838), .B(n1791), .Z(n1793) );
  XOR U4840 ( .A(x[82]), .B(x[87]), .Z(n1818) );
  NANDN U4841 ( .A(n1793), .B(n1818), .Z(n1743) );
  XNOR U4842 ( .A(n1744), .B(n1743), .Z(n1760) );
  XNOR U4843 ( .A(n1745), .B(n1760), .Z(n1746) );
  XOR U4844 ( .A(n1747), .B(n1746), .Z(n1773) );
  NAND U4845 ( .A(n1777), .B(n1773), .Z(n1767) );
  IV U4846 ( .A(n1773), .Z(n1774) );
  XOR U4847 ( .A(n1783), .B(n1774), .Z(n1765) );
  XOR U4848 ( .A(x[82]), .B(x[81]), .Z(n1748) );
  XNOR U4849 ( .A(n1826), .B(n1748), .Z(n1800) );
  NAND U4850 ( .A(n1800), .B(n1791), .Z(n1755) );
  XNOR U4851 ( .A(x[84]), .B(n1838), .Z(n1811) );
  XOR U4852 ( .A(n1801), .B(n1748), .Z(n1806) );
  NANDN U4853 ( .A(n1790), .B(n1806), .Z(n1756) );
  XOR U4854 ( .A(n1811), .B(n1756), .Z(n1751) );
  XOR U4855 ( .A(x[80]), .B(n1749), .Z(n1750) );
  XNOR U4856 ( .A(n1751), .B(n1750), .Z(n1752) );
  XOR U4857 ( .A(n1753), .B(n1752), .Z(n1754) );
  XOR U4858 ( .A(n1755), .B(n1754), .Z(n1785) );
  IV U4859 ( .A(n1785), .Z(n1780) );
  AND U4860 ( .A(n1777), .B(n1780), .Z(n1763) );
  ANDN U4861 ( .B(x[80]), .A(n1811), .Z(n1762) );
  XNOR U4862 ( .A(n1800), .B(n1756), .Z(n1758) );
  XNOR U4863 ( .A(x[81]), .B(n1791), .Z(n1757) );
  XNOR U4864 ( .A(n1758), .B(n1757), .Z(n1759) );
  XOR U4865 ( .A(n1760), .B(n1759), .Z(n1761) );
  XOR U4866 ( .A(n1762), .B(n1761), .Z(n1775) );
  IV U4867 ( .A(n1775), .Z(n1781) );
  XNOR U4868 ( .A(n1763), .B(n1781), .Z(n1764) );
  NAND U4869 ( .A(n1765), .B(n1764), .Z(n1766) );
  NAND U4870 ( .A(n1767), .B(n1766), .Z(n1845) );
  NAND U4871 ( .A(n1781), .B(n1774), .Z(n1768) );
  NAND U4872 ( .A(n1780), .B(n1768), .Z(n1771) );
  XOR U4873 ( .A(n1774), .B(n1777), .Z(n1769) );
  NAND U4874 ( .A(n1775), .B(n1769), .Z(n1770) );
  AND U4875 ( .A(n1771), .B(n1770), .Z(n1827) );
  XNOR U4876 ( .A(n1845), .B(n1827), .Z(n1802) );
  OR U4877 ( .A(n1802), .B(n1772), .Z(n1795) );
  NAND U4878 ( .A(n1783), .B(n1773), .Z(n1779) );
  AND U4879 ( .A(n1775), .B(n1774), .Z(n1782) );
  XNOR U4880 ( .A(n1782), .B(n1780), .Z(n1776) );
  NAND U4881 ( .A(n1777), .B(n1776), .Z(n1778) );
  AND U4882 ( .A(n1779), .B(n1778), .Z(n1799) );
  NAND U4883 ( .A(n1781), .B(n1780), .Z(n1787) );
  XNOR U4884 ( .A(n1783), .B(n1782), .Z(n1784) );
  NAND U4885 ( .A(n1785), .B(n1784), .Z(n1786) );
  NAND U4886 ( .A(n1787), .B(n1786), .Z(n1839) );
  XNOR U4887 ( .A(n1799), .B(n1839), .Z(n1817) );
  XOR U4888 ( .A(n1817), .B(n1802), .Z(n1804) );
  OR U4889 ( .A(n1804), .B(n1788), .Z(n1789) );
  XNOR U4890 ( .A(n1795), .B(n1789), .Z(n1821) );
  XOR U4891 ( .A(n1799), .B(n1845), .Z(n1807) );
  OR U4892 ( .A(n1790), .B(n1807), .Z(n1847) );
  NANDN U4893 ( .A(n1799), .B(n1791), .Z(n1792) );
  XNOR U4894 ( .A(n1847), .B(n1792), .Z(n1825) );
  XOR U4895 ( .A(n1821), .B(n1825), .Z(n1810) );
  NANDN U4896 ( .A(n1793), .B(n1817), .Z(n1794) );
  XNOR U4897 ( .A(n1795), .B(n1794), .Z(n1853) );
  XNOR U4898 ( .A(n1839), .B(n1827), .Z(n1829) );
  NANDN U4899 ( .A(n1829), .B(n1796), .Z(n1813) );
  NAND U4900 ( .A(n1797), .B(n1827), .Z(n1798) );
  XNOR U4901 ( .A(n1813), .B(n1798), .Z(n1844) );
  XOR U4902 ( .A(n1853), .B(n1844), .Z(n1836) );
  XNOR U4903 ( .A(n1810), .B(n1836), .Z(z[80]) );
  ANDN U4904 ( .B(n1800), .A(n1799), .Z(n1809) );
  NANDN U4905 ( .A(n1802), .B(n1801), .Z(n1820) );
  NANDN U4906 ( .A(n1804), .B(n1803), .Z(n1805) );
  XNOR U4907 ( .A(n1820), .B(n1805), .Z(n1848) );
  NANDN U4908 ( .A(n1807), .B(n1806), .Z(n1814) );
  XNOR U4909 ( .A(n1848), .B(n1814), .Z(n1808) );
  XOR U4910 ( .A(n1809), .B(n1808), .Z(n1834) );
  XOR U4911 ( .A(n1834), .B(n1810), .Z(n1852) );
  ANDN U4912 ( .B(n1845), .A(n1811), .Z(n1816) );
  NAND U4913 ( .A(n1838), .B(n1839), .Z(n1812) );
  XNOR U4914 ( .A(n1813), .B(n1812), .Z(n1824) );
  XNOR U4915 ( .A(n1814), .B(n1824), .Z(n1815) );
  XNOR U4916 ( .A(n1816), .B(n1815), .Z(n1823) );
  NAND U4917 ( .A(n1818), .B(n1817), .Z(n1819) );
  XNOR U4918 ( .A(n1820), .B(n1819), .Z(n1830) );
  XNOR U4919 ( .A(n1821), .B(n1830), .Z(n1822) );
  XOR U4920 ( .A(n1823), .B(n1822), .Z(n1833) );
  XNOR U4921 ( .A(n1852), .B(n1833), .Z(z[81]) );
  XNOR U4922 ( .A(n1825), .B(n1824), .Z(z[82]) );
  ANDN U4923 ( .B(n1827), .A(n1826), .Z(n1832) );
  NANDN U4924 ( .A(n1829), .B(n1828), .Z(n1842) );
  XNOR U4925 ( .A(n1830), .B(n1842), .Z(n1831) );
  XOR U4926 ( .A(n1832), .B(n1831), .Z(n1851) );
  XOR U4927 ( .A(n1834), .B(n1833), .Z(n1835) );
  XOR U4928 ( .A(n1851), .B(n1835), .Z(z[83]) );
  XOR U4929 ( .A(n1836), .B(z[82]), .Z(z[84]) );
  XNOR U4930 ( .A(n1838), .B(n1837), .Z(n1840) );
  NAND U4931 ( .A(n1840), .B(n1839), .Z(n1841) );
  XOR U4932 ( .A(n1842), .B(n1841), .Z(n1843) );
  XNOR U4933 ( .A(n1844), .B(n1843), .Z(n1850) );
  NAND U4934 ( .A(x[80]), .B(n1845), .Z(n1846) );
  XNOR U4935 ( .A(n1847), .B(n1846), .Z(n1854) );
  XNOR U4936 ( .A(n1848), .B(n1854), .Z(n1849) );
  XOR U4937 ( .A(n1850), .B(n1849), .Z(z[85]) );
  XNOR U4938 ( .A(n1852), .B(n1851), .Z(z[86]) );
  XNOR U4939 ( .A(n1854), .B(n1853), .Z(n1855) );
  XNOR U4940 ( .A(z[81]), .B(n1855), .Z(z[87]) );
  XOR U4941 ( .A(x[88]), .B(x[94]), .Z(n1856) );
  XOR U4942 ( .A(x[93]), .B(n1856), .Z(n1963) );
  IV U4943 ( .A(n1963), .Z(n1858) );
  IV U4944 ( .A(x[89]), .Z(n1962) );
  NAND U4945 ( .A(n1858), .B(n1962), .Z(n1865) );
  XOR U4946 ( .A(x[91]), .B(x[89]), .Z(n1861) );
  XNOR U4947 ( .A(x[90]), .B(n1856), .Z(n1857) );
  XNOR U4948 ( .A(n1861), .B(n1857), .Z(n1920) );
  XNOR U4949 ( .A(n1858), .B(n1920), .Z(n1919) );
  IV U4950 ( .A(x[95]), .Z(n1859) );
  XNOR U4951 ( .A(x[89]), .B(n1859), .Z(n1953) );
  NAND U4952 ( .A(n1919), .B(n1953), .Z(n1868) );
  XNOR U4953 ( .A(n1858), .B(n1859), .Z(n1951) );
  XOR U4954 ( .A(n1920), .B(n1951), .Z(n1876) );
  XOR U4955 ( .A(n1868), .B(n1876), .Z(n1863) );
  XNOR U4956 ( .A(x[88]), .B(n1920), .Z(n1895) );
  XOR U4957 ( .A(x[92]), .B(n1859), .Z(n1860) );
  IV U4958 ( .A(n1860), .Z(n1924) );
  NANDN U4959 ( .A(n1895), .B(n1924), .Z(n1867) );
  XOR U4960 ( .A(n1861), .B(n1860), .Z(n1913) );
  XOR U4961 ( .A(n1919), .B(n1913), .Z(n1911) );
  XOR U4962 ( .A(x[90]), .B(x[92]), .Z(n1926) );
  NANDN U4963 ( .A(n1911), .B(n1926), .Z(n1862) );
  XNOR U4964 ( .A(n1867), .B(n1862), .Z(n1872) );
  XOR U4965 ( .A(n1863), .B(n1872), .Z(n1864) );
  XOR U4966 ( .A(n1865), .B(n1864), .Z(n1906) );
  IV U4967 ( .A(n1906), .Z(n1900) );
  ANDN U4968 ( .B(n1951), .A(n1920), .Z(n1870) );
  XNOR U4969 ( .A(x[88]), .B(n1913), .Z(n1914) );
  XNOR U4970 ( .A(n1963), .B(n1914), .Z(n1916) );
  XOR U4971 ( .A(x[90]), .B(x[95]), .Z(n1941) );
  NANDN U4972 ( .A(n1916), .B(n1941), .Z(n1866) );
  XNOR U4973 ( .A(n1867), .B(n1866), .Z(n1883) );
  XNOR U4974 ( .A(n1868), .B(n1883), .Z(n1869) );
  XOR U4975 ( .A(n1870), .B(n1869), .Z(n1896) );
  NAND U4976 ( .A(n1900), .B(n1896), .Z(n1890) );
  IV U4977 ( .A(n1896), .Z(n1897) );
  XOR U4978 ( .A(n1906), .B(n1897), .Z(n1888) );
  XOR U4979 ( .A(x[90]), .B(x[89]), .Z(n1871) );
  XNOR U4980 ( .A(n1951), .B(n1871), .Z(n1923) );
  NAND U4981 ( .A(n1923), .B(n1914), .Z(n1878) );
  XNOR U4982 ( .A(x[92]), .B(n1963), .Z(n1934) );
  XOR U4983 ( .A(n1924), .B(n1871), .Z(n1929) );
  NANDN U4984 ( .A(n1913), .B(n1929), .Z(n1879) );
  XOR U4985 ( .A(n1934), .B(n1879), .Z(n1874) );
  XOR U4986 ( .A(x[88]), .B(n1872), .Z(n1873) );
  XNOR U4987 ( .A(n1874), .B(n1873), .Z(n1875) );
  XOR U4988 ( .A(n1876), .B(n1875), .Z(n1877) );
  XOR U4989 ( .A(n1878), .B(n1877), .Z(n1908) );
  IV U4990 ( .A(n1908), .Z(n1903) );
  AND U4991 ( .A(n1900), .B(n1903), .Z(n1886) );
  ANDN U4992 ( .B(x[88]), .A(n1934), .Z(n1885) );
  XNOR U4993 ( .A(n1923), .B(n1879), .Z(n1881) );
  XNOR U4994 ( .A(x[89]), .B(n1914), .Z(n1880) );
  XNOR U4995 ( .A(n1881), .B(n1880), .Z(n1882) );
  XOR U4996 ( .A(n1883), .B(n1882), .Z(n1884) );
  XOR U4997 ( .A(n1885), .B(n1884), .Z(n1898) );
  IV U4998 ( .A(n1898), .Z(n1904) );
  XNOR U4999 ( .A(n1886), .B(n1904), .Z(n1887) );
  NAND U5000 ( .A(n1888), .B(n1887), .Z(n1889) );
  NAND U5001 ( .A(n1890), .B(n1889), .Z(n1970) );
  NAND U5002 ( .A(n1904), .B(n1897), .Z(n1891) );
  NAND U5003 ( .A(n1903), .B(n1891), .Z(n1894) );
  XOR U5004 ( .A(n1897), .B(n1900), .Z(n1892) );
  NAND U5005 ( .A(n1898), .B(n1892), .Z(n1893) );
  AND U5006 ( .A(n1894), .B(n1893), .Z(n1952) );
  XNOR U5007 ( .A(n1970), .B(n1952), .Z(n1925) );
  OR U5008 ( .A(n1925), .B(n1895), .Z(n1918) );
  NAND U5009 ( .A(n1906), .B(n1896), .Z(n1902) );
  AND U5010 ( .A(n1898), .B(n1897), .Z(n1905) );
  XNOR U5011 ( .A(n1905), .B(n1903), .Z(n1899) );
  NAND U5012 ( .A(n1900), .B(n1899), .Z(n1901) );
  AND U5013 ( .A(n1902), .B(n1901), .Z(n1922) );
  NAND U5014 ( .A(n1904), .B(n1903), .Z(n1910) );
  XNOR U5015 ( .A(n1906), .B(n1905), .Z(n1907) );
  NAND U5016 ( .A(n1908), .B(n1907), .Z(n1909) );
  NAND U5017 ( .A(n1910), .B(n1909), .Z(n1964) );
  XNOR U5018 ( .A(n1922), .B(n1964), .Z(n1940) );
  XOR U5019 ( .A(n1940), .B(n1925), .Z(n1927) );
  OR U5020 ( .A(n1927), .B(n1911), .Z(n1912) );
  XNOR U5021 ( .A(n1918), .B(n1912), .Z(n1944) );
  XOR U5022 ( .A(n1922), .B(n1970), .Z(n1930) );
  OR U5023 ( .A(n1913), .B(n1930), .Z(n1972) );
  NANDN U5024 ( .A(n1922), .B(n1914), .Z(n1915) );
  XNOR U5025 ( .A(n1972), .B(n1915), .Z(n1950) );
  XOR U5026 ( .A(n1944), .B(n1950), .Z(n1933) );
  NANDN U5027 ( .A(n1916), .B(n1940), .Z(n1917) );
  XNOR U5028 ( .A(n1918), .B(n1917), .Z(n1978) );
  XNOR U5029 ( .A(n1964), .B(n1952), .Z(n1954) );
  NANDN U5030 ( .A(n1954), .B(n1919), .Z(n1936) );
  NAND U5031 ( .A(n1920), .B(n1952), .Z(n1921) );
  XNOR U5032 ( .A(n1936), .B(n1921), .Z(n1969) );
  XOR U5033 ( .A(n1978), .B(n1969), .Z(n1961) );
  XNOR U5034 ( .A(n1933), .B(n1961), .Z(z[88]) );
  ANDN U5035 ( .B(n1923), .A(n1922), .Z(n1932) );
  NANDN U5036 ( .A(n1925), .B(n1924), .Z(n1943) );
  NANDN U5037 ( .A(n1927), .B(n1926), .Z(n1928) );
  XNOR U5038 ( .A(n1943), .B(n1928), .Z(n1973) );
  NANDN U5039 ( .A(n1930), .B(n1929), .Z(n1937) );
  XNOR U5040 ( .A(n1973), .B(n1937), .Z(n1931) );
  XOR U5041 ( .A(n1932), .B(n1931), .Z(n1959) );
  XOR U5042 ( .A(n1959), .B(n1933), .Z(n1977) );
  ANDN U5043 ( .B(n1970), .A(n1934), .Z(n1939) );
  NAND U5044 ( .A(n1963), .B(n1964), .Z(n1935) );
  XNOR U5045 ( .A(n1936), .B(n1935), .Z(n1949) );
  XNOR U5046 ( .A(n1937), .B(n1949), .Z(n1938) );
  XNOR U5047 ( .A(n1939), .B(n1938), .Z(n1946) );
  NAND U5048 ( .A(n1941), .B(n1940), .Z(n1942) );
  XNOR U5049 ( .A(n1943), .B(n1942), .Z(n1955) );
  XNOR U5050 ( .A(n1944), .B(n1955), .Z(n1945) );
  XOR U5051 ( .A(n1946), .B(n1945), .Z(n1958) );
  XNOR U5052 ( .A(n1977), .B(n1958), .Z(z[89]) );
  XNOR U5053 ( .A(n1948), .B(n1947), .Z(z[8]) );
  XNOR U5054 ( .A(n1950), .B(n1949), .Z(z[90]) );
  ANDN U5055 ( .B(n1952), .A(n1951), .Z(n1957) );
  NANDN U5056 ( .A(n1954), .B(n1953), .Z(n1967) );
  XNOR U5057 ( .A(n1955), .B(n1967), .Z(n1956) );
  XOR U5058 ( .A(n1957), .B(n1956), .Z(n1976) );
  XOR U5059 ( .A(n1959), .B(n1958), .Z(n1960) );
  XOR U5060 ( .A(n1976), .B(n1960), .Z(z[91]) );
  XOR U5061 ( .A(n1961), .B(z[90]), .Z(z[92]) );
  XNOR U5062 ( .A(n1963), .B(n1962), .Z(n1965) );
  NAND U5063 ( .A(n1965), .B(n1964), .Z(n1966) );
  XOR U5064 ( .A(n1967), .B(n1966), .Z(n1968) );
  XNOR U5065 ( .A(n1969), .B(n1968), .Z(n1975) );
  NAND U5066 ( .A(x[88]), .B(n1970), .Z(n1971) );
  XNOR U5067 ( .A(n1972), .B(n1971), .Z(n1979) );
  XNOR U5068 ( .A(n1973), .B(n1979), .Z(n1974) );
  XOR U5069 ( .A(n1975), .B(n1974), .Z(z[93]) );
  XNOR U5070 ( .A(n1977), .B(n1976), .Z(z[94]) );
  XNOR U5071 ( .A(n1979), .B(n1978), .Z(n1980) );
  XNOR U5072 ( .A(z[89]), .B(n1980), .Z(z[95]) );
  XNOR U5073 ( .A(n1982), .B(n1981), .Z(z[96]) );
  XOR U5074 ( .A(n1984), .B(n1983), .Z(n1985) );
  XOR U5075 ( .A(n1986), .B(n1985), .Z(z[99]) );
endmodule


module SubBytes_6 ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986;

  XOR U2962 ( .A(x[24]), .B(x[30]), .Z(n834) );
  XOR U2963 ( .A(x[16]), .B(x[22]), .Z(n685) );
  XOR U2964 ( .A(x[53]), .B(n1218), .Z(n1323) );
  XNOR U2965 ( .A(n328), .B(n339), .Z(n341) );
  XNOR U2966 ( .A(n815), .B(x[19]), .Z(n689) );
  XNOR U2967 ( .A(n1324), .B(x[51]), .Z(n1222) );
  XNOR U2968 ( .A(n170), .B(n162), .Z(n143) );
  XOR U2969 ( .A(x[81]), .B(x[83]), .Z(n1738) );
  XOR U2970 ( .A(n493), .B(n494), .Z(n646) );
  XOR U2971 ( .A(x[21]), .B(n685), .Z(n814) );
  XOR U2972 ( .A(x[85]), .B(n1733), .Z(n1838) );
  IV U2973 ( .A(x[1]), .Z(n1447) );
  XOR U2974 ( .A(x[0]), .B(x[6]), .Z(n2) );
  XOR U2975 ( .A(x[5]), .B(n2), .Z(n1446) );
  IV U2976 ( .A(n1446), .Z(n3) );
  AND U2977 ( .A(n1447), .B(n3), .Z(n10) );
  XNOR U2978 ( .A(x[3]), .B(n1447), .Z(n6) );
  XNOR U2979 ( .A(x[2]), .B(n6), .Z(n1) );
  XNOR U2980 ( .A(n2), .B(n1), .Z(n66) );
  IV U2981 ( .A(n66), .Z(n12) );
  XNOR U2982 ( .A(n12), .B(n1446), .Z(n65) );
  IV U2983 ( .A(x[7]), .Z(n4) );
  XNOR U2984 ( .A(x[1]), .B(n4), .Z(n1085) );
  NAND U2985 ( .A(n65), .B(n1085), .Z(n15) );
  XNOR U2986 ( .A(n4), .B(n3), .Z(n11) );
  IV U2987 ( .A(n11), .Z(n1083) );
  XOR U2988 ( .A(n66), .B(n1083), .Z(n31) );
  XNOR U2989 ( .A(n15), .B(n31), .Z(n8) );
  XOR U2990 ( .A(x[0]), .B(n12), .Z(n41) );
  XOR U2991 ( .A(x[4]), .B(n4), .Z(n5) );
  IV U2992 ( .A(n5), .Z(n790) );
  NANDN U2993 ( .A(n41), .B(n790), .Z(n14) );
  XNOR U2994 ( .A(n6), .B(n5), .Z(n59) );
  XNOR U2995 ( .A(n65), .B(n59), .Z(n57) );
  XOR U2996 ( .A(x[2]), .B(x[4]), .Z(n792) );
  NANDN U2997 ( .A(n57), .B(n792), .Z(n7) );
  XOR U2998 ( .A(n14), .B(n7), .Z(n33) );
  XNOR U2999 ( .A(n8), .B(n33), .Z(n9) );
  XOR U3000 ( .A(n10), .B(n9), .Z(n46) );
  IV U3001 ( .A(n46), .Z(n52) );
  AND U3002 ( .A(n12), .B(n11), .Z(n17) );
  XOR U3003 ( .A(x[0]), .B(n59), .Z(n60) );
  XNOR U3004 ( .A(n1446), .B(n60), .Z(n62) );
  XOR U3005 ( .A(x[2]), .B(x[7]), .Z(n807) );
  NANDN U3006 ( .A(n62), .B(n807), .Z(n13) );
  XNOR U3007 ( .A(n14), .B(n13), .Z(n22) );
  XNOR U3008 ( .A(n15), .B(n22), .Z(n16) );
  XOR U3009 ( .A(n17), .B(n16), .Z(n42) );
  XNOR U3010 ( .A(x[4]), .B(n1446), .Z(n800) );
  ANDN U3011 ( .B(x[0]), .A(n800), .Z(n24) );
  XOR U3012 ( .A(x[2]), .B(x[1]), .Z(n18) );
  XOR U3013 ( .A(n1083), .B(n18), .Z(n789) );
  XOR U3014 ( .A(n790), .B(n18), .Z(n795) );
  NAND U3015 ( .A(n59), .B(n795), .Z(n26) );
  XNOR U3016 ( .A(n789), .B(n26), .Z(n20) );
  XNOR U3017 ( .A(x[1]), .B(n60), .Z(n19) );
  XNOR U3018 ( .A(n20), .B(n19), .Z(n21) );
  XOR U3019 ( .A(n22), .B(n21), .Z(n23) );
  XOR U3020 ( .A(n24), .B(n23), .Z(n44) );
  NAND U3021 ( .A(n42), .B(n44), .Z(n25) );
  NAND U3022 ( .A(n52), .B(n25), .Z(n36) );
  IV U3023 ( .A(n42), .Z(n43) );
  IV U3024 ( .A(n44), .Z(n50) );
  XOR U3025 ( .A(n26), .B(n800), .Z(n29) );
  AND U3026 ( .A(n789), .B(n60), .Z(n27) );
  XNOR U3027 ( .A(x[0]), .B(n27), .Z(n28) );
  XNOR U3028 ( .A(n29), .B(n28), .Z(n30) );
  XNOR U3029 ( .A(n31), .B(n30), .Z(n32) );
  XNOR U3030 ( .A(n33), .B(n32), .Z(n54) );
  IV U3031 ( .A(n54), .Z(n49) );
  XOR U3032 ( .A(n50), .B(n49), .Z(n34) );
  NAND U3033 ( .A(n43), .B(n34), .Z(n35) );
  AND U3034 ( .A(n36), .B(n35), .Z(n1454) );
  NAND U3035 ( .A(n50), .B(n43), .Z(n37) );
  NAND U3036 ( .A(n49), .B(n37), .Z(n40) );
  XOR U3037 ( .A(n43), .B(n46), .Z(n38) );
  NAND U3038 ( .A(n44), .B(n38), .Z(n39) );
  AND U3039 ( .A(n40), .B(n39), .Z(n1084) );
  XNOR U3040 ( .A(n1454), .B(n1084), .Z(n791) );
  OR U3041 ( .A(n791), .B(n41), .Z(n64) );
  NAND U3042 ( .A(n52), .B(n42), .Z(n48) );
  AND U3043 ( .A(n44), .B(n43), .Z(n51) );
  XNOR U3044 ( .A(n49), .B(n51), .Z(n45) );
  NAND U3045 ( .A(n46), .B(n45), .Z(n47) );
  AND U3046 ( .A(n48), .B(n47), .Z(n788) );
  NAND U3047 ( .A(n50), .B(n49), .Z(n56) );
  XNOR U3048 ( .A(n52), .B(n51), .Z(n53) );
  NAND U3049 ( .A(n54), .B(n53), .Z(n55) );
  NAND U3050 ( .A(n56), .B(n55), .Z(n1448) );
  XNOR U3051 ( .A(n788), .B(n1448), .Z(n806) );
  XOR U3052 ( .A(n806), .B(n791), .Z(n793) );
  OR U3053 ( .A(n793), .B(n57), .Z(n58) );
  XNOR U3054 ( .A(n64), .B(n58), .Z(n810) );
  XOR U3055 ( .A(n788), .B(n1454), .Z(n796) );
  NANDN U3056 ( .A(n796), .B(n59), .Z(n1456) );
  NANDN U3057 ( .A(n788), .B(n60), .Z(n61) );
  XNOR U3058 ( .A(n1456), .B(n61), .Z(n953) );
  XOR U3059 ( .A(n810), .B(n953), .Z(n799) );
  NANDN U3060 ( .A(n62), .B(n806), .Z(n63) );
  XNOR U3061 ( .A(n64), .B(n63), .Z(n1730) );
  XNOR U3062 ( .A(n1448), .B(n1084), .Z(n1086) );
  NANDN U3063 ( .A(n1086), .B(n65), .Z(n802) );
  NAND U3064 ( .A(n66), .B(n1084), .Z(n67) );
  XNOR U3065 ( .A(n802), .B(n67), .Z(n1453) );
  XOR U3066 ( .A(n1730), .B(n1453), .Z(n1309) );
  XNOR U3067 ( .A(n799), .B(n1309), .Z(z[0]) );
  XOR U3068 ( .A(x[96]), .B(x[102]), .Z(n68) );
  XOR U3069 ( .A(x[101]), .B(n68), .Z(n135) );
  XOR U3070 ( .A(x[100]), .B(n135), .Z(n171) );
  AND U3071 ( .A(x[96]), .B(n171), .Z(n78) );
  XOR U3072 ( .A(x[97]), .B(x[99]), .Z(n71) );
  XNOR U3073 ( .A(n68), .B(x[98]), .Z(n69) );
  XOR U3074 ( .A(n71), .B(n69), .Z(n129) );
  XOR U3075 ( .A(x[96]), .B(n129), .Z(n128) );
  XNOR U3076 ( .A(x[103]), .B(x[100]), .Z(n70) );
  IV U3077 ( .A(n70), .Z(n142) );
  NANDN U3078 ( .A(n128), .B(n142), .Z(n80) );
  IV U3079 ( .A(n135), .Z(n91) );
  XNOR U3080 ( .A(n71), .B(n70), .Z(n123) );
  XOR U3081 ( .A(x[96]), .B(n123), .Z(n124) );
  XOR U3082 ( .A(n91), .B(n124), .Z(n126) );
  XOR U3083 ( .A(x[98]), .B(x[103]), .Z(n164) );
  NANDN U3084 ( .A(n126), .B(n164), .Z(n72) );
  XNOR U3085 ( .A(n80), .B(n72), .Z(n87) );
  XNOR U3086 ( .A(n135), .B(x[103]), .Z(n161) );
  XOR U3087 ( .A(x[97]), .B(x[98]), .Z(n73) );
  XNOR U3088 ( .A(n161), .B(n73), .Z(n151) );
  XOR U3089 ( .A(n142), .B(n73), .Z(n152) );
  NAND U3090 ( .A(n123), .B(n152), .Z(n81) );
  XNOR U3091 ( .A(n151), .B(n81), .Z(n75) );
  XNOR U3092 ( .A(x[97]), .B(n124), .Z(n74) );
  XNOR U3093 ( .A(n75), .B(n74), .Z(n76) );
  XOR U3094 ( .A(n87), .B(n76), .Z(n77) );
  XOR U3095 ( .A(n78), .B(n77), .Z(n115) );
  IV U3096 ( .A(n115), .Z(n108) );
  XNOR U3097 ( .A(n129), .B(n135), .Z(n105) );
  XNOR U3098 ( .A(n105), .B(n123), .Z(n158) );
  XNOR U3099 ( .A(x[98]), .B(x[100]), .Z(n144) );
  OR U3100 ( .A(n158), .B(n144), .Z(n79) );
  XOR U3101 ( .A(n80), .B(n79), .Z(n94) );
  XNOR U3102 ( .A(n129), .B(n161), .Z(n92) );
  XNOR U3103 ( .A(n81), .B(n171), .Z(n84) );
  AND U3104 ( .A(n151), .B(n124), .Z(n82) );
  XNOR U3105 ( .A(x[96]), .B(n82), .Z(n83) );
  XNOR U3106 ( .A(n84), .B(n83), .Z(n85) );
  XOR U3107 ( .A(n92), .B(n85), .Z(n86) );
  XOR U3108 ( .A(n94), .B(n86), .Z(n118) );
  AND U3109 ( .A(n129), .B(n161), .Z(n89) );
  IV U3110 ( .A(x[97]), .Z(n136) );
  XNOR U3111 ( .A(n136), .B(x[103]), .Z(n133) );
  NAND U3112 ( .A(n105), .B(n133), .Z(n93) );
  XNOR U3113 ( .A(n93), .B(n87), .Z(n88) );
  XOR U3114 ( .A(n89), .B(n88), .Z(n107) );
  NAND U3115 ( .A(n118), .B(n107), .Z(n90) );
  NAND U3116 ( .A(n108), .B(n90), .Z(n99) );
  IV U3117 ( .A(n118), .Z(n102) );
  NAND U3118 ( .A(n91), .B(n136), .Z(n97) );
  XOR U3119 ( .A(n93), .B(n92), .Z(n95) );
  XNOR U3120 ( .A(n95), .B(n94), .Z(n96) );
  XOR U3121 ( .A(n97), .B(n96), .Z(n114) );
  IV U3122 ( .A(n107), .Z(n116) );
  XOR U3123 ( .A(n114), .B(n116), .Z(n111) );
  NAND U3124 ( .A(n102), .B(n111), .Z(n98) );
  AND U3125 ( .A(n99), .B(n98), .Z(n127) );
  NAND U3126 ( .A(n118), .B(n108), .Z(n104) );
  AND U3127 ( .A(n115), .B(n116), .Z(n100) );
  XNOR U3128 ( .A(n114), .B(n100), .Z(n101) );
  NAND U3129 ( .A(n102), .B(n101), .Z(n103) );
  AND U3130 ( .A(n104), .B(n103), .Z(n138) );
  XNOR U3131 ( .A(n127), .B(n138), .Z(n134) );
  NANDN U3132 ( .A(n134), .B(n105), .Z(n131) );
  NANDN U3133 ( .A(n138), .B(n135), .Z(n106) );
  XNOR U3134 ( .A(n131), .B(n106), .Z(n173) );
  IV U3135 ( .A(n114), .Z(n120) );
  NAND U3136 ( .A(n120), .B(n107), .Z(n113) );
  AND U3137 ( .A(n120), .B(n118), .Z(n109) );
  XNOR U3138 ( .A(n109), .B(n108), .Z(n110) );
  NAND U3139 ( .A(n111), .B(n110), .Z(n112) );
  NAND U3140 ( .A(n113), .B(n112), .Z(n170) );
  NAND U3141 ( .A(n114), .B(n116), .Z(n122) );
  NAND U3142 ( .A(n116), .B(n115), .Z(n117) );
  XNOR U3143 ( .A(n118), .B(n117), .Z(n119) );
  NAND U3144 ( .A(n120), .B(n119), .Z(n121) );
  NAND U3145 ( .A(n122), .B(n121), .Z(n150) );
  XOR U3146 ( .A(n170), .B(n150), .Z(n153) );
  NANDN U3147 ( .A(n153), .B(n123), .Z(n147) );
  NANDN U3148 ( .A(n150), .B(n124), .Z(n125) );
  XNOR U3149 ( .A(n147), .B(n125), .Z(n160) );
  XNOR U3150 ( .A(n173), .B(n160), .Z(z[98]) );
  XOR U3151 ( .A(n150), .B(n138), .Z(n163) );
  ANDN U3152 ( .B(n163), .A(n126), .Z(n184) );
  IV U3153 ( .A(n127), .Z(n162) );
  OR U3154 ( .A(n143), .B(n128), .Z(n182) );
  NANDN U3155 ( .A(n129), .B(n162), .Z(n130) );
  XNOR U3156 ( .A(n131), .B(n130), .Z(n141) );
  XNOR U3157 ( .A(n182), .B(n141), .Z(n132) );
  XOR U3158 ( .A(n184), .B(n132), .Z(n1982) );
  XNOR U3159 ( .A(n1982), .B(z[98]), .Z(z[100]) );
  NANDN U3160 ( .A(n134), .B(n133), .Z(n167) );
  XNOR U3161 ( .A(n136), .B(n135), .Z(n137) );
  NANDN U3162 ( .A(n138), .B(n137), .Z(n139) );
  XOR U3163 ( .A(n167), .B(n139), .Z(n140) );
  XNOR U3164 ( .A(n141), .B(n140), .Z(n149) );
  NANDN U3165 ( .A(n143), .B(n142), .Z(n166) );
  XNOR U3166 ( .A(n143), .B(n163), .Z(n157) );
  NANDN U3167 ( .A(n144), .B(n157), .Z(n145) );
  XNOR U3168 ( .A(n166), .B(n145), .Z(n154) );
  NAND U3169 ( .A(n170), .B(x[96]), .Z(n146) );
  XNOR U3170 ( .A(n147), .B(n146), .Z(n181) );
  XNOR U3171 ( .A(n154), .B(n181), .Z(n148) );
  XOR U3172 ( .A(n149), .B(n148), .Z(z[101]) );
  ANDN U3173 ( .B(n151), .A(n150), .Z(n156) );
  NANDN U3174 ( .A(n153), .B(n152), .Z(n172) );
  XNOR U3175 ( .A(n172), .B(n154), .Z(n155) );
  XOR U3176 ( .A(n156), .B(n155), .Z(n1983) );
  NANDN U3177 ( .A(n158), .B(n157), .Z(n159) );
  XOR U3178 ( .A(n182), .B(n159), .Z(n176) );
  XOR U3179 ( .A(n176), .B(n160), .Z(n1981) );
  XNOR U3180 ( .A(n1983), .B(n1981), .Z(n180) );
  ANDN U3181 ( .B(n162), .A(n161), .Z(n169) );
  NAND U3182 ( .A(n164), .B(n163), .Z(n165) );
  XNOR U3183 ( .A(n166), .B(n165), .Z(n177) );
  XNOR U3184 ( .A(n177), .B(n167), .Z(n168) );
  XOR U3185 ( .A(n169), .B(n168), .Z(n1986) );
  XNOR U3186 ( .A(n180), .B(n1986), .Z(z[102]) );
  AND U3187 ( .A(n171), .B(n170), .Z(n175) );
  XNOR U3188 ( .A(n173), .B(n172), .Z(n174) );
  XNOR U3189 ( .A(n175), .B(n174), .Z(n179) );
  XOR U3190 ( .A(n177), .B(n176), .Z(n178) );
  XOR U3191 ( .A(n179), .B(n178), .Z(n1984) );
  XNOR U3192 ( .A(n1984), .B(n180), .Z(z[97]) );
  XNOR U3193 ( .A(n182), .B(n181), .Z(n183) );
  XNOR U3194 ( .A(n184), .B(n183), .Z(n185) );
  XOR U3195 ( .A(n185), .B(z[97]), .Z(z[103]) );
  IV U3196 ( .A(x[105]), .Z(n292) );
  XOR U3197 ( .A(x[104]), .B(x[110]), .Z(n187) );
  XOR U3198 ( .A(x[109]), .B(n187), .Z(n291) );
  IV U3199 ( .A(n291), .Z(n188) );
  AND U3200 ( .A(n292), .B(n188), .Z(n195) );
  XNOR U3201 ( .A(x[107]), .B(n292), .Z(n191) );
  XNOR U3202 ( .A(x[106]), .B(n191), .Z(n186) );
  XNOR U3203 ( .A(n187), .B(n186), .Z(n251) );
  IV U3204 ( .A(n251), .Z(n197) );
  XNOR U3205 ( .A(n197), .B(n291), .Z(n250) );
  IV U3206 ( .A(x[111]), .Z(n189) );
  XNOR U3207 ( .A(x[105]), .B(n189), .Z(n282) );
  NAND U3208 ( .A(n250), .B(n282), .Z(n200) );
  XNOR U3209 ( .A(n189), .B(n188), .Z(n196) );
  IV U3210 ( .A(n196), .Z(n280) );
  XOR U3211 ( .A(n251), .B(n280), .Z(n216) );
  XNOR U3212 ( .A(n200), .B(n216), .Z(n193) );
  XOR U3213 ( .A(x[104]), .B(n197), .Z(n226) );
  XOR U3214 ( .A(x[108]), .B(n189), .Z(n190) );
  IV U3215 ( .A(n190), .Z(n255) );
  NANDN U3216 ( .A(n226), .B(n255), .Z(n199) );
  XNOR U3217 ( .A(n191), .B(n190), .Z(n244) );
  XNOR U3218 ( .A(n250), .B(n244), .Z(n242) );
  XOR U3219 ( .A(x[106]), .B(x[108]), .Z(n257) );
  NANDN U3220 ( .A(n242), .B(n257), .Z(n192) );
  XOR U3221 ( .A(n199), .B(n192), .Z(n218) );
  XNOR U3222 ( .A(n193), .B(n218), .Z(n194) );
  XOR U3223 ( .A(n195), .B(n194), .Z(n231) );
  IV U3224 ( .A(n231), .Z(n237) );
  AND U3225 ( .A(n197), .B(n196), .Z(n202) );
  XOR U3226 ( .A(x[104]), .B(n244), .Z(n245) );
  XNOR U3227 ( .A(n291), .B(n245), .Z(n247) );
  XOR U3228 ( .A(x[106]), .B(x[111]), .Z(n272) );
  NANDN U3229 ( .A(n247), .B(n272), .Z(n198) );
  XNOR U3230 ( .A(n199), .B(n198), .Z(n207) );
  XNOR U3231 ( .A(n200), .B(n207), .Z(n201) );
  XOR U3232 ( .A(n202), .B(n201), .Z(n227) );
  XNOR U3233 ( .A(x[108]), .B(n291), .Z(n265) );
  ANDN U3234 ( .B(x[104]), .A(n265), .Z(n209) );
  XOR U3235 ( .A(x[106]), .B(x[105]), .Z(n203) );
  XOR U3236 ( .A(n280), .B(n203), .Z(n254) );
  XOR U3237 ( .A(n255), .B(n203), .Z(n260) );
  NAND U3238 ( .A(n244), .B(n260), .Z(n211) );
  XNOR U3239 ( .A(n254), .B(n211), .Z(n205) );
  XNOR U3240 ( .A(x[105]), .B(n245), .Z(n204) );
  XNOR U3241 ( .A(n205), .B(n204), .Z(n206) );
  XOR U3242 ( .A(n207), .B(n206), .Z(n208) );
  XOR U3243 ( .A(n209), .B(n208), .Z(n229) );
  NAND U3244 ( .A(n227), .B(n229), .Z(n210) );
  NAND U3245 ( .A(n237), .B(n210), .Z(n221) );
  IV U3246 ( .A(n227), .Z(n228) );
  IV U3247 ( .A(n229), .Z(n235) );
  XOR U3248 ( .A(n211), .B(n265), .Z(n214) );
  AND U3249 ( .A(n254), .B(n245), .Z(n212) );
  XNOR U3250 ( .A(x[104]), .B(n212), .Z(n213) );
  XNOR U3251 ( .A(n214), .B(n213), .Z(n215) );
  XNOR U3252 ( .A(n216), .B(n215), .Z(n217) );
  XNOR U3253 ( .A(n218), .B(n217), .Z(n239) );
  IV U3254 ( .A(n239), .Z(n234) );
  XOR U3255 ( .A(n235), .B(n234), .Z(n219) );
  NAND U3256 ( .A(n228), .B(n219), .Z(n220) );
  AND U3257 ( .A(n221), .B(n220), .Z(n299) );
  NAND U3258 ( .A(n235), .B(n228), .Z(n222) );
  NAND U3259 ( .A(n234), .B(n222), .Z(n225) );
  XOR U3260 ( .A(n228), .B(n231), .Z(n223) );
  NAND U3261 ( .A(n229), .B(n223), .Z(n224) );
  AND U3262 ( .A(n225), .B(n224), .Z(n281) );
  XNOR U3263 ( .A(n299), .B(n281), .Z(n256) );
  OR U3264 ( .A(n256), .B(n226), .Z(n249) );
  NAND U3265 ( .A(n237), .B(n227), .Z(n233) );
  AND U3266 ( .A(n229), .B(n228), .Z(n236) );
  XNOR U3267 ( .A(n234), .B(n236), .Z(n230) );
  NAND U3268 ( .A(n231), .B(n230), .Z(n232) );
  AND U3269 ( .A(n233), .B(n232), .Z(n253) );
  NAND U3270 ( .A(n235), .B(n234), .Z(n241) );
  XNOR U3271 ( .A(n237), .B(n236), .Z(n238) );
  NAND U3272 ( .A(n239), .B(n238), .Z(n240) );
  NAND U3273 ( .A(n241), .B(n240), .Z(n293) );
  XNOR U3274 ( .A(n253), .B(n293), .Z(n271) );
  XOR U3275 ( .A(n271), .B(n256), .Z(n258) );
  OR U3276 ( .A(n258), .B(n242), .Z(n243) );
  XNOR U3277 ( .A(n249), .B(n243), .Z(n275) );
  XOR U3278 ( .A(n253), .B(n299), .Z(n261) );
  NANDN U3279 ( .A(n261), .B(n244), .Z(n301) );
  NANDN U3280 ( .A(n253), .B(n245), .Z(n246) );
  XNOR U3281 ( .A(n301), .B(n246), .Z(n279) );
  XOR U3282 ( .A(n275), .B(n279), .Z(n264) );
  NANDN U3283 ( .A(n247), .B(n271), .Z(n248) );
  XNOR U3284 ( .A(n249), .B(n248), .Z(n366) );
  XNOR U3285 ( .A(n293), .B(n281), .Z(n283) );
  NANDN U3286 ( .A(n283), .B(n250), .Z(n267) );
  NAND U3287 ( .A(n251), .B(n281), .Z(n252) );
  XNOR U3288 ( .A(n267), .B(n252), .Z(n298) );
  XOR U3289 ( .A(n366), .B(n298), .Z(n290) );
  XNOR U3290 ( .A(n264), .B(n290), .Z(z[104]) );
  ANDN U3291 ( .B(n254), .A(n253), .Z(n263) );
  NANDN U3292 ( .A(n256), .B(n255), .Z(n274) );
  NANDN U3293 ( .A(n258), .B(n257), .Z(n259) );
  XNOR U3294 ( .A(n274), .B(n259), .Z(n302) );
  NANDN U3295 ( .A(n261), .B(n260), .Z(n268) );
  XNOR U3296 ( .A(n302), .B(n268), .Z(n262) );
  XOR U3297 ( .A(n263), .B(n262), .Z(n288) );
  XOR U3298 ( .A(n288), .B(n264), .Z(n365) );
  ANDN U3299 ( .B(n299), .A(n265), .Z(n270) );
  NAND U3300 ( .A(n291), .B(n293), .Z(n266) );
  XNOR U3301 ( .A(n267), .B(n266), .Z(n278) );
  XNOR U3302 ( .A(n268), .B(n278), .Z(n269) );
  XNOR U3303 ( .A(n270), .B(n269), .Z(n277) );
  NAND U3304 ( .A(n272), .B(n271), .Z(n273) );
  XNOR U3305 ( .A(n274), .B(n273), .Z(n284) );
  XNOR U3306 ( .A(n275), .B(n284), .Z(n276) );
  XOR U3307 ( .A(n277), .B(n276), .Z(n287) );
  XNOR U3308 ( .A(n365), .B(n287), .Z(z[105]) );
  XNOR U3309 ( .A(n279), .B(n278), .Z(z[106]) );
  AND U3310 ( .A(n281), .B(n280), .Z(n286) );
  NANDN U3311 ( .A(n283), .B(n282), .Z(n296) );
  XNOR U3312 ( .A(n284), .B(n296), .Z(n285) );
  XOR U3313 ( .A(n286), .B(n285), .Z(n364) );
  XOR U3314 ( .A(n288), .B(n287), .Z(n289) );
  XOR U3315 ( .A(n364), .B(n289), .Z(z[107]) );
  XOR U3316 ( .A(n290), .B(z[106]), .Z(z[108]) );
  XNOR U3317 ( .A(n292), .B(n291), .Z(n294) );
  NAND U3318 ( .A(n294), .B(n293), .Z(n295) );
  XOR U3319 ( .A(n296), .B(n295), .Z(n297) );
  XNOR U3320 ( .A(n298), .B(n297), .Z(n304) );
  NAND U3321 ( .A(n299), .B(x[104]), .Z(n300) );
  XNOR U3322 ( .A(n301), .B(n300), .Z(n367) );
  XNOR U3323 ( .A(n302), .B(n367), .Z(n303) );
  XOR U3324 ( .A(n304), .B(n303), .Z(z[109]) );
  IV U3325 ( .A(x[15]), .Z(n311) );
  IV U3326 ( .A(x[10]), .Z(n315) );
  XOR U3327 ( .A(x[11]), .B(x[9]), .Z(n307) );
  XOR U3328 ( .A(n315), .B(n307), .Z(n352) );
  IV U3329 ( .A(n352), .Z(n309) );
  XOR U3330 ( .A(x[13]), .B(n309), .Z(n305) );
  IV U3331 ( .A(x[9]), .Z(n655) );
  XNOR U3332 ( .A(n311), .B(n655), .Z(n515) );
  NAND U3333 ( .A(n305), .B(n515), .Z(n306) );
  XNOR U3334 ( .A(n311), .B(n306), .Z(n339) );
  XOR U3335 ( .A(x[12]), .B(n311), .Z(n314) );
  XNOR U3336 ( .A(x[14]), .B(n309), .Z(n497) );
  NOR U3337 ( .A(n314), .B(n497), .Z(n318) );
  IV U3338 ( .A(x[13]), .Z(n353) );
  XOR U3339 ( .A(x[8]), .B(x[14]), .Z(n310) );
  XOR U3340 ( .A(n353), .B(n310), .Z(n325) );
  IV U3341 ( .A(n325), .Z(n656) );
  XOR U3342 ( .A(n314), .B(n307), .Z(n316) );
  XNOR U3343 ( .A(x[8]), .B(n316), .Z(n350) );
  XNOR U3344 ( .A(n656), .B(n350), .Z(n648) );
  XNOR U3345 ( .A(x[15]), .B(n315), .Z(n673) );
  NANDN U3346 ( .A(n648), .B(n673), .Z(n308) );
  XOR U3347 ( .A(n318), .B(n308), .Z(n333) );
  XOR U3348 ( .A(n310), .B(n309), .Z(n313) );
  XNOR U3349 ( .A(n325), .B(n311), .Z(n516) );
  ANDN U3350 ( .B(n313), .A(n516), .Z(n312) );
  XOR U3351 ( .A(n333), .B(n312), .Z(n328) );
  IV U3352 ( .A(n313), .Z(n647) );
  IV U3353 ( .A(n314), .Z(n507) );
  XNOR U3354 ( .A(n655), .B(n315), .Z(n321) );
  XOR U3355 ( .A(n507), .B(n321), .Z(n501) );
  IV U3356 ( .A(n316), .Z(n344) );
  NANDN U3357 ( .A(n501), .B(n344), .Z(n329) );
  XNOR U3358 ( .A(x[12]), .B(x[10]), .Z(n508) );
  XNOR U3359 ( .A(n648), .B(n497), .Z(n498) );
  OR U3360 ( .A(n508), .B(n498), .Z(n317) );
  XOR U3361 ( .A(n318), .B(n317), .Z(n327) );
  XOR U3362 ( .A(n329), .B(n327), .Z(n320) );
  XNOR U3363 ( .A(x[8]), .B(n507), .Z(n319) );
  XNOR U3364 ( .A(n320), .B(n319), .Z(n323) );
  XOR U3365 ( .A(n321), .B(n516), .Z(n505) );
  NAND U3366 ( .A(n350), .B(n505), .Z(n322) );
  XNOR U3367 ( .A(n323), .B(n322), .Z(n324) );
  XOR U3368 ( .A(n647), .B(n324), .Z(n356) );
  IV U3369 ( .A(n356), .Z(n359) );
  NAND U3370 ( .A(n325), .B(n655), .Z(n326) );
  XOR U3371 ( .A(n327), .B(n326), .Z(n338) );
  XNOR U3372 ( .A(n328), .B(n338), .Z(n348) );
  NAND U3373 ( .A(n359), .B(n348), .Z(n337) );
  XOR U3374 ( .A(n656), .B(x[12]), .Z(n502) );
  AND U3375 ( .A(n502), .B(x[8]), .Z(n335) );
  XNOR U3376 ( .A(n505), .B(n329), .Z(n331) );
  XNOR U3377 ( .A(x[9]), .B(n350), .Z(n330) );
  XNOR U3378 ( .A(n331), .B(n330), .Z(n332) );
  XOR U3379 ( .A(n333), .B(n332), .Z(n334) );
  XNOR U3380 ( .A(n335), .B(n334), .Z(n358) );
  NANDN U3381 ( .A(n348), .B(n358), .Z(n336) );
  AND U3382 ( .A(n337), .B(n336), .Z(n342) );
  XNOR U3383 ( .A(n339), .B(n338), .Z(n345) );
  NANDN U3384 ( .A(n345), .B(n356), .Z(n340) );
  XNOR U3385 ( .A(n342), .B(n340), .Z(n354) );
  OR U3386 ( .A(n341), .B(n354), .Z(n495) );
  NANDN U3387 ( .A(n358), .B(n341), .Z(n347) );
  XOR U3388 ( .A(n345), .B(n342), .Z(n343) );
  XNOR U3389 ( .A(n347), .B(n343), .Z(n355) );
  NOR U3390 ( .A(n355), .B(n345), .Z(n349) );
  XOR U3391 ( .A(n495), .B(n349), .Z(n500) );
  NANDN U3392 ( .A(n500), .B(n344), .Z(n664) );
  ANDN U3393 ( .B(n359), .A(n345), .Z(n346) );
  XNOR U3394 ( .A(n347), .B(n346), .Z(n361) );
  OR U3395 ( .A(n361), .B(n348), .Z(n496) );
  XNOR U3396 ( .A(n496), .B(n349), .Z(n504) );
  AND U3397 ( .A(n504), .B(n350), .Z(n351) );
  XOR U3398 ( .A(n664), .B(n351), .Z(n670) );
  XOR U3399 ( .A(n353), .B(n352), .Z(n357) );
  ANDN U3400 ( .B(n358), .A(n354), .Z(n493) );
  NOR U3401 ( .A(n356), .B(n355), .Z(n362) );
  XOR U3402 ( .A(n493), .B(n362), .Z(n514) );
  NAND U3403 ( .A(n357), .B(n514), .Z(n651) );
  XOR U3404 ( .A(n359), .B(n358), .Z(n360) );
  NANDN U3405 ( .A(n361), .B(n360), .Z(n494) );
  XOR U3406 ( .A(n494), .B(n362), .Z(n658) );
  NANDN U3407 ( .A(n658), .B(n656), .Z(n363) );
  XNOR U3408 ( .A(n651), .B(n363), .Z(n519) );
  XOR U3409 ( .A(n670), .B(n519), .Z(n654) );
  IV U3410 ( .A(n654), .Z(z[10]) );
  XNOR U3411 ( .A(n365), .B(n364), .Z(z[110]) );
  XNOR U3412 ( .A(n367), .B(n366), .Z(n368) );
  XNOR U3413 ( .A(z[105]), .B(n368), .Z(z[111]) );
  IV U3414 ( .A(x[113]), .Z(n475) );
  XOR U3415 ( .A(x[112]), .B(x[118]), .Z(n370) );
  XOR U3416 ( .A(x[117]), .B(n370), .Z(n474) );
  IV U3417 ( .A(n474), .Z(n371) );
  AND U3418 ( .A(n475), .B(n371), .Z(n378) );
  XNOR U3419 ( .A(x[115]), .B(n475), .Z(n374) );
  XNOR U3420 ( .A(x[114]), .B(n374), .Z(n369) );
  XNOR U3421 ( .A(n370), .B(n369), .Z(n434) );
  IV U3422 ( .A(n434), .Z(n380) );
  XNOR U3423 ( .A(n380), .B(n474), .Z(n433) );
  IV U3424 ( .A(x[119]), .Z(n372) );
  XNOR U3425 ( .A(x[113]), .B(n372), .Z(n465) );
  NAND U3426 ( .A(n433), .B(n465), .Z(n383) );
  XNOR U3427 ( .A(n372), .B(n371), .Z(n379) );
  IV U3428 ( .A(n379), .Z(n463) );
  XOR U3429 ( .A(n434), .B(n463), .Z(n399) );
  XNOR U3430 ( .A(n383), .B(n399), .Z(n376) );
  XOR U3431 ( .A(x[112]), .B(n380), .Z(n409) );
  XOR U3432 ( .A(x[116]), .B(n372), .Z(n373) );
  IV U3433 ( .A(n373), .Z(n438) );
  NANDN U3434 ( .A(n409), .B(n438), .Z(n382) );
  XNOR U3435 ( .A(n374), .B(n373), .Z(n427) );
  XNOR U3436 ( .A(n433), .B(n427), .Z(n425) );
  XOR U3437 ( .A(x[114]), .B(x[116]), .Z(n440) );
  NANDN U3438 ( .A(n425), .B(n440), .Z(n375) );
  XOR U3439 ( .A(n382), .B(n375), .Z(n401) );
  XNOR U3440 ( .A(n376), .B(n401), .Z(n377) );
  XOR U3441 ( .A(n378), .B(n377), .Z(n414) );
  IV U3442 ( .A(n414), .Z(n420) );
  AND U3443 ( .A(n380), .B(n379), .Z(n385) );
  XOR U3444 ( .A(x[112]), .B(n427), .Z(n428) );
  XNOR U3445 ( .A(n474), .B(n428), .Z(n430) );
  XOR U3446 ( .A(x[114]), .B(x[119]), .Z(n455) );
  NANDN U3447 ( .A(n430), .B(n455), .Z(n381) );
  XNOR U3448 ( .A(n382), .B(n381), .Z(n390) );
  XNOR U3449 ( .A(n383), .B(n390), .Z(n384) );
  XOR U3450 ( .A(n385), .B(n384), .Z(n410) );
  XNOR U3451 ( .A(x[116]), .B(n474), .Z(n448) );
  ANDN U3452 ( .B(x[112]), .A(n448), .Z(n392) );
  XOR U3453 ( .A(x[114]), .B(x[113]), .Z(n386) );
  XOR U3454 ( .A(n463), .B(n386), .Z(n437) );
  XOR U3455 ( .A(n438), .B(n386), .Z(n443) );
  NAND U3456 ( .A(n427), .B(n443), .Z(n394) );
  XNOR U3457 ( .A(n437), .B(n394), .Z(n388) );
  XNOR U3458 ( .A(x[113]), .B(n428), .Z(n387) );
  XNOR U3459 ( .A(n388), .B(n387), .Z(n389) );
  XOR U3460 ( .A(n390), .B(n389), .Z(n391) );
  XOR U3461 ( .A(n392), .B(n391), .Z(n412) );
  NAND U3462 ( .A(n410), .B(n412), .Z(n393) );
  NAND U3463 ( .A(n420), .B(n393), .Z(n404) );
  IV U3464 ( .A(n410), .Z(n411) );
  IV U3465 ( .A(n412), .Z(n418) );
  XOR U3466 ( .A(n394), .B(n448), .Z(n397) );
  AND U3467 ( .A(n437), .B(n428), .Z(n395) );
  XNOR U3468 ( .A(x[112]), .B(n395), .Z(n396) );
  XNOR U3469 ( .A(n397), .B(n396), .Z(n398) );
  XNOR U3470 ( .A(n399), .B(n398), .Z(n400) );
  XNOR U3471 ( .A(n401), .B(n400), .Z(n422) );
  IV U3472 ( .A(n422), .Z(n417) );
  XOR U3473 ( .A(n418), .B(n417), .Z(n402) );
  NAND U3474 ( .A(n411), .B(n402), .Z(n403) );
  AND U3475 ( .A(n404), .B(n403), .Z(n482) );
  NAND U3476 ( .A(n418), .B(n411), .Z(n405) );
  NAND U3477 ( .A(n417), .B(n405), .Z(n408) );
  XOR U3478 ( .A(n411), .B(n414), .Z(n406) );
  NAND U3479 ( .A(n412), .B(n406), .Z(n407) );
  AND U3480 ( .A(n408), .B(n407), .Z(n464) );
  XNOR U3481 ( .A(n482), .B(n464), .Z(n439) );
  OR U3482 ( .A(n439), .B(n409), .Z(n432) );
  NAND U3483 ( .A(n420), .B(n410), .Z(n416) );
  AND U3484 ( .A(n412), .B(n411), .Z(n419) );
  XNOR U3485 ( .A(n417), .B(n419), .Z(n413) );
  NAND U3486 ( .A(n414), .B(n413), .Z(n415) );
  AND U3487 ( .A(n416), .B(n415), .Z(n436) );
  NAND U3488 ( .A(n418), .B(n417), .Z(n424) );
  XNOR U3489 ( .A(n420), .B(n419), .Z(n421) );
  NAND U3490 ( .A(n422), .B(n421), .Z(n423) );
  NAND U3491 ( .A(n424), .B(n423), .Z(n476) );
  XNOR U3492 ( .A(n436), .B(n476), .Z(n454) );
  XOR U3493 ( .A(n454), .B(n439), .Z(n441) );
  OR U3494 ( .A(n441), .B(n425), .Z(n426) );
  XNOR U3495 ( .A(n432), .B(n426), .Z(n458) );
  XOR U3496 ( .A(n436), .B(n482), .Z(n444) );
  NANDN U3497 ( .A(n444), .B(n427), .Z(n484) );
  NANDN U3498 ( .A(n436), .B(n428), .Z(n429) );
  XNOR U3499 ( .A(n484), .B(n429), .Z(n462) );
  XOR U3500 ( .A(n458), .B(n462), .Z(n447) );
  NANDN U3501 ( .A(n430), .B(n454), .Z(n431) );
  XNOR U3502 ( .A(n432), .B(n431), .Z(n490) );
  XNOR U3503 ( .A(n476), .B(n464), .Z(n466) );
  NANDN U3504 ( .A(n466), .B(n433), .Z(n450) );
  NAND U3505 ( .A(n434), .B(n464), .Z(n435) );
  XNOR U3506 ( .A(n450), .B(n435), .Z(n481) );
  XOR U3507 ( .A(n490), .B(n481), .Z(n473) );
  XNOR U3508 ( .A(n447), .B(n473), .Z(z[112]) );
  ANDN U3509 ( .B(n437), .A(n436), .Z(n446) );
  NANDN U3510 ( .A(n439), .B(n438), .Z(n457) );
  NANDN U3511 ( .A(n441), .B(n440), .Z(n442) );
  XNOR U3512 ( .A(n457), .B(n442), .Z(n485) );
  NANDN U3513 ( .A(n444), .B(n443), .Z(n451) );
  XNOR U3514 ( .A(n485), .B(n451), .Z(n445) );
  XOR U3515 ( .A(n446), .B(n445), .Z(n471) );
  XOR U3516 ( .A(n471), .B(n447), .Z(n489) );
  ANDN U3517 ( .B(n482), .A(n448), .Z(n453) );
  NAND U3518 ( .A(n474), .B(n476), .Z(n449) );
  XNOR U3519 ( .A(n450), .B(n449), .Z(n461) );
  XNOR U3520 ( .A(n451), .B(n461), .Z(n452) );
  XNOR U3521 ( .A(n453), .B(n452), .Z(n460) );
  NAND U3522 ( .A(n455), .B(n454), .Z(n456) );
  XNOR U3523 ( .A(n457), .B(n456), .Z(n467) );
  XNOR U3524 ( .A(n458), .B(n467), .Z(n459) );
  XOR U3525 ( .A(n460), .B(n459), .Z(n470) );
  XNOR U3526 ( .A(n489), .B(n470), .Z(z[113]) );
  XNOR U3527 ( .A(n462), .B(n461), .Z(z[114]) );
  AND U3528 ( .A(n464), .B(n463), .Z(n469) );
  NANDN U3529 ( .A(n466), .B(n465), .Z(n479) );
  XNOR U3530 ( .A(n467), .B(n479), .Z(n468) );
  XOR U3531 ( .A(n469), .B(n468), .Z(n488) );
  XOR U3532 ( .A(n471), .B(n470), .Z(n472) );
  XOR U3533 ( .A(n488), .B(n472), .Z(z[115]) );
  XOR U3534 ( .A(n473), .B(z[114]), .Z(z[116]) );
  XNOR U3535 ( .A(n475), .B(n474), .Z(n477) );
  NAND U3536 ( .A(n477), .B(n476), .Z(n478) );
  XOR U3537 ( .A(n479), .B(n478), .Z(n480) );
  XNOR U3538 ( .A(n481), .B(n480), .Z(n487) );
  NAND U3539 ( .A(n482), .B(x[112]), .Z(n483) );
  XNOR U3540 ( .A(n484), .B(n483), .Z(n491) );
  XNOR U3541 ( .A(n485), .B(n491), .Z(n486) );
  XOR U3542 ( .A(n487), .B(n486), .Z(z[117]) );
  XNOR U3543 ( .A(n489), .B(n488), .Z(z[118]) );
  XNOR U3544 ( .A(n491), .B(n490), .Z(n492) );
  XNOR U3545 ( .A(z[113]), .B(n492), .Z(z[119]) );
  XNOR U3546 ( .A(n496), .B(n495), .Z(n662) );
  XOR U3547 ( .A(n646), .B(n662), .Z(n506) );
  NANDN U3548 ( .A(n497), .B(n506), .Z(n650) );
  XNOR U3549 ( .A(n658), .B(n504), .Z(n672) );
  XNOR U3550 ( .A(n506), .B(n672), .Z(n509) );
  OR U3551 ( .A(n498), .B(n509), .Z(n499) );
  XNOR U3552 ( .A(n650), .B(n499), .Z(n671) );
  OR U3553 ( .A(n501), .B(n500), .Z(n511) );
  ANDN U3554 ( .B(n502), .A(n662), .Z(n503) );
  XNOR U3555 ( .A(n511), .B(n503), .Z(n678) );
  AND U3556 ( .A(n505), .B(n504), .Z(n513) );
  NAND U3557 ( .A(n507), .B(n506), .Z(n675) );
  OR U3558 ( .A(n509), .B(n508), .Z(n510) );
  XNOR U3559 ( .A(n675), .B(n510), .Z(n667) );
  XNOR U3560 ( .A(n667), .B(n511), .Z(n512) );
  XOR U3561 ( .A(n513), .B(n512), .Z(n682) );
  NANDN U3562 ( .A(n515), .B(n514), .Z(n660) );
  OR U3563 ( .A(n516), .B(n646), .Z(n517) );
  XOR U3564 ( .A(n660), .B(n517), .Z(n518) );
  XNOR U3565 ( .A(n682), .B(n518), .Z(n677) );
  XNOR U3566 ( .A(n519), .B(n677), .Z(n520) );
  XOR U3567 ( .A(n678), .B(n520), .Z(n521) );
  XOR U3568 ( .A(n671), .B(n521), .Z(z[11]) );
  IV U3569 ( .A(x[121]), .Z(n628) );
  XOR U3570 ( .A(x[120]), .B(x[126]), .Z(n523) );
  XOR U3571 ( .A(x[125]), .B(n523), .Z(n627) );
  IV U3572 ( .A(n627), .Z(n524) );
  AND U3573 ( .A(n628), .B(n524), .Z(n531) );
  XNOR U3574 ( .A(x[123]), .B(n628), .Z(n527) );
  XNOR U3575 ( .A(x[122]), .B(n527), .Z(n522) );
  XNOR U3576 ( .A(n523), .B(n522), .Z(n587) );
  IV U3577 ( .A(n587), .Z(n533) );
  XNOR U3578 ( .A(n533), .B(n627), .Z(n586) );
  IV U3579 ( .A(x[127]), .Z(n525) );
  XNOR U3580 ( .A(x[121]), .B(n525), .Z(n618) );
  NAND U3581 ( .A(n586), .B(n618), .Z(n536) );
  XNOR U3582 ( .A(n525), .B(n524), .Z(n532) );
  IV U3583 ( .A(n532), .Z(n616) );
  XOR U3584 ( .A(n587), .B(n616), .Z(n552) );
  XNOR U3585 ( .A(n536), .B(n552), .Z(n529) );
  XOR U3586 ( .A(x[120]), .B(n533), .Z(n562) );
  XOR U3587 ( .A(x[124]), .B(n525), .Z(n526) );
  IV U3588 ( .A(n526), .Z(n591) );
  NANDN U3589 ( .A(n562), .B(n591), .Z(n535) );
  XNOR U3590 ( .A(n527), .B(n526), .Z(n580) );
  XNOR U3591 ( .A(n586), .B(n580), .Z(n578) );
  XOR U3592 ( .A(x[122]), .B(x[124]), .Z(n593) );
  NANDN U3593 ( .A(n578), .B(n593), .Z(n528) );
  XOR U3594 ( .A(n535), .B(n528), .Z(n554) );
  XNOR U3595 ( .A(n529), .B(n554), .Z(n530) );
  XOR U3596 ( .A(n531), .B(n530), .Z(n567) );
  IV U3597 ( .A(n567), .Z(n573) );
  AND U3598 ( .A(n533), .B(n532), .Z(n538) );
  XOR U3599 ( .A(x[120]), .B(n580), .Z(n581) );
  XNOR U3600 ( .A(n627), .B(n581), .Z(n583) );
  XOR U3601 ( .A(x[122]), .B(x[127]), .Z(n608) );
  NANDN U3602 ( .A(n583), .B(n608), .Z(n534) );
  XNOR U3603 ( .A(n535), .B(n534), .Z(n543) );
  XNOR U3604 ( .A(n536), .B(n543), .Z(n537) );
  XOR U3605 ( .A(n538), .B(n537), .Z(n563) );
  XNOR U3606 ( .A(x[124]), .B(n627), .Z(n601) );
  ANDN U3607 ( .B(x[120]), .A(n601), .Z(n545) );
  XOR U3608 ( .A(x[122]), .B(x[121]), .Z(n539) );
  XOR U3609 ( .A(n616), .B(n539), .Z(n590) );
  XOR U3610 ( .A(n591), .B(n539), .Z(n596) );
  NAND U3611 ( .A(n580), .B(n596), .Z(n547) );
  XNOR U3612 ( .A(n590), .B(n547), .Z(n541) );
  XNOR U3613 ( .A(x[121]), .B(n581), .Z(n540) );
  XNOR U3614 ( .A(n541), .B(n540), .Z(n542) );
  XOR U3615 ( .A(n543), .B(n542), .Z(n544) );
  XOR U3616 ( .A(n545), .B(n544), .Z(n565) );
  NAND U3617 ( .A(n563), .B(n565), .Z(n546) );
  NAND U3618 ( .A(n573), .B(n546), .Z(n557) );
  IV U3619 ( .A(n563), .Z(n564) );
  IV U3620 ( .A(n565), .Z(n571) );
  XOR U3621 ( .A(n547), .B(n601), .Z(n550) );
  AND U3622 ( .A(n590), .B(n581), .Z(n548) );
  XNOR U3623 ( .A(x[120]), .B(n548), .Z(n549) );
  XNOR U3624 ( .A(n550), .B(n549), .Z(n551) );
  XNOR U3625 ( .A(n552), .B(n551), .Z(n553) );
  XNOR U3626 ( .A(n554), .B(n553), .Z(n575) );
  IV U3627 ( .A(n575), .Z(n570) );
  XOR U3628 ( .A(n571), .B(n570), .Z(n555) );
  NAND U3629 ( .A(n564), .B(n555), .Z(n556) );
  AND U3630 ( .A(n557), .B(n556), .Z(n635) );
  NAND U3631 ( .A(n571), .B(n564), .Z(n558) );
  NAND U3632 ( .A(n570), .B(n558), .Z(n561) );
  XOR U3633 ( .A(n564), .B(n567), .Z(n559) );
  NAND U3634 ( .A(n565), .B(n559), .Z(n560) );
  AND U3635 ( .A(n561), .B(n560), .Z(n617) );
  XNOR U3636 ( .A(n635), .B(n617), .Z(n592) );
  OR U3637 ( .A(n592), .B(n562), .Z(n585) );
  NAND U3638 ( .A(n573), .B(n563), .Z(n569) );
  AND U3639 ( .A(n565), .B(n564), .Z(n572) );
  XNOR U3640 ( .A(n570), .B(n572), .Z(n566) );
  NAND U3641 ( .A(n567), .B(n566), .Z(n568) );
  AND U3642 ( .A(n569), .B(n568), .Z(n589) );
  NAND U3643 ( .A(n571), .B(n570), .Z(n577) );
  XNOR U3644 ( .A(n573), .B(n572), .Z(n574) );
  NAND U3645 ( .A(n575), .B(n574), .Z(n576) );
  NAND U3646 ( .A(n577), .B(n576), .Z(n629) );
  XNOR U3647 ( .A(n589), .B(n629), .Z(n607) );
  XOR U3648 ( .A(n607), .B(n592), .Z(n594) );
  OR U3649 ( .A(n594), .B(n578), .Z(n579) );
  XNOR U3650 ( .A(n585), .B(n579), .Z(n611) );
  XOR U3651 ( .A(n589), .B(n635), .Z(n597) );
  NANDN U3652 ( .A(n597), .B(n580), .Z(n637) );
  NANDN U3653 ( .A(n589), .B(n581), .Z(n582) );
  XNOR U3654 ( .A(n637), .B(n582), .Z(n615) );
  XOR U3655 ( .A(n611), .B(n615), .Z(n600) );
  NANDN U3656 ( .A(n583), .B(n607), .Z(n584) );
  XNOR U3657 ( .A(n585), .B(n584), .Z(n643) );
  XNOR U3658 ( .A(n629), .B(n617), .Z(n619) );
  NANDN U3659 ( .A(n619), .B(n586), .Z(n603) );
  NAND U3660 ( .A(n587), .B(n617), .Z(n588) );
  XNOR U3661 ( .A(n603), .B(n588), .Z(n634) );
  XOR U3662 ( .A(n643), .B(n634), .Z(n626) );
  XNOR U3663 ( .A(n600), .B(n626), .Z(z[120]) );
  ANDN U3664 ( .B(n590), .A(n589), .Z(n599) );
  NANDN U3665 ( .A(n592), .B(n591), .Z(n610) );
  NANDN U3666 ( .A(n594), .B(n593), .Z(n595) );
  XNOR U3667 ( .A(n610), .B(n595), .Z(n638) );
  NANDN U3668 ( .A(n597), .B(n596), .Z(n604) );
  XNOR U3669 ( .A(n638), .B(n604), .Z(n598) );
  XOR U3670 ( .A(n599), .B(n598), .Z(n624) );
  XOR U3671 ( .A(n624), .B(n600), .Z(n642) );
  ANDN U3672 ( .B(n635), .A(n601), .Z(n606) );
  NAND U3673 ( .A(n627), .B(n629), .Z(n602) );
  XNOR U3674 ( .A(n603), .B(n602), .Z(n614) );
  XNOR U3675 ( .A(n604), .B(n614), .Z(n605) );
  XNOR U3676 ( .A(n606), .B(n605), .Z(n613) );
  NAND U3677 ( .A(n608), .B(n607), .Z(n609) );
  XNOR U3678 ( .A(n610), .B(n609), .Z(n620) );
  XNOR U3679 ( .A(n611), .B(n620), .Z(n612) );
  XOR U3680 ( .A(n613), .B(n612), .Z(n623) );
  XNOR U3681 ( .A(n642), .B(n623), .Z(z[121]) );
  XNOR U3682 ( .A(n615), .B(n614), .Z(z[122]) );
  AND U3683 ( .A(n617), .B(n616), .Z(n622) );
  NANDN U3684 ( .A(n619), .B(n618), .Z(n632) );
  XNOR U3685 ( .A(n620), .B(n632), .Z(n621) );
  XOR U3686 ( .A(n622), .B(n621), .Z(n641) );
  XOR U3687 ( .A(n624), .B(n623), .Z(n625) );
  XOR U3688 ( .A(n641), .B(n625), .Z(z[123]) );
  XOR U3689 ( .A(n626), .B(z[122]), .Z(z[124]) );
  XNOR U3690 ( .A(n628), .B(n627), .Z(n630) );
  NAND U3691 ( .A(n630), .B(n629), .Z(n631) );
  XOR U3692 ( .A(n632), .B(n631), .Z(n633) );
  XNOR U3693 ( .A(n634), .B(n633), .Z(n640) );
  NAND U3694 ( .A(n635), .B(x[120]), .Z(n636) );
  XNOR U3695 ( .A(n637), .B(n636), .Z(n644) );
  XNOR U3696 ( .A(n638), .B(n644), .Z(n639) );
  XOR U3697 ( .A(n640), .B(n639), .Z(z[125]) );
  XNOR U3698 ( .A(n642), .B(n641), .Z(z[126]) );
  XNOR U3699 ( .A(n644), .B(n643), .Z(n645) );
  XNOR U3700 ( .A(z[121]), .B(n645), .Z(z[127]) );
  NOR U3701 ( .A(n647), .B(n646), .Z(n653) );
  NANDN U3702 ( .A(n648), .B(n672), .Z(n649) );
  XNOR U3703 ( .A(n650), .B(n649), .Z(n663) );
  XNOR U3704 ( .A(n651), .B(n663), .Z(n652) );
  XOR U3705 ( .A(n653), .B(n652), .Z(n1947) );
  XOR U3706 ( .A(n1947), .B(n654), .Z(z[12]) );
  XNOR U3707 ( .A(n656), .B(n655), .Z(n657) );
  NANDN U3708 ( .A(n658), .B(n657), .Z(n659) );
  XOR U3709 ( .A(n660), .B(n659), .Z(n661) );
  XNOR U3710 ( .A(n1947), .B(n661), .Z(n669) );
  ANDN U3711 ( .B(x[8]), .A(n662), .Z(n666) );
  XNOR U3712 ( .A(n664), .B(n663), .Z(n665) );
  XOR U3713 ( .A(n666), .B(n665), .Z(n683) );
  XNOR U3714 ( .A(n667), .B(n683), .Z(n668) );
  XOR U3715 ( .A(n669), .B(n668), .Z(z[13]) );
  XNOR U3716 ( .A(n671), .B(n670), .Z(n1948) );
  NAND U3717 ( .A(n673), .B(n672), .Z(n674) );
  XNOR U3718 ( .A(n675), .B(n674), .Z(n679) );
  XNOR U3719 ( .A(n1948), .B(n679), .Z(n676) );
  XOR U3720 ( .A(n677), .B(n676), .Z(z[14]) );
  XNOR U3721 ( .A(n679), .B(n678), .Z(n680) );
  XNOR U3722 ( .A(z[10]), .B(n680), .Z(n681) );
  XOR U3723 ( .A(n682), .B(n681), .Z(z[9]) );
  XNOR U3724 ( .A(n683), .B(z[9]), .Z(z[15]) );
  IV U3725 ( .A(x[17]), .Z(n815) );
  IV U3726 ( .A(n814), .Z(n686) );
  AND U3727 ( .A(n815), .B(n686), .Z(n693) );
  XNOR U3728 ( .A(x[18]), .B(n689), .Z(n684) );
  XNOR U3729 ( .A(n685), .B(n684), .Z(n749) );
  IV U3730 ( .A(n749), .Z(n695) );
  XNOR U3731 ( .A(n695), .B(n814), .Z(n748) );
  IV U3732 ( .A(x[23]), .Z(n687) );
  XNOR U3733 ( .A(x[17]), .B(n687), .Z(n780) );
  NAND U3734 ( .A(n748), .B(n780), .Z(n698) );
  XNOR U3735 ( .A(n687), .B(n686), .Z(n694) );
  IV U3736 ( .A(n694), .Z(n778) );
  XOR U3737 ( .A(n749), .B(n778), .Z(n714) );
  XNOR U3738 ( .A(n698), .B(n714), .Z(n691) );
  XOR U3739 ( .A(x[16]), .B(n695), .Z(n724) );
  XOR U3740 ( .A(x[20]), .B(n687), .Z(n688) );
  IV U3741 ( .A(n688), .Z(n753) );
  NANDN U3742 ( .A(n724), .B(n753), .Z(n697) );
  XNOR U3743 ( .A(n689), .B(n688), .Z(n742) );
  XNOR U3744 ( .A(n748), .B(n742), .Z(n740) );
  XOR U3745 ( .A(x[18]), .B(x[20]), .Z(n755) );
  NANDN U3746 ( .A(n740), .B(n755), .Z(n690) );
  XOR U3747 ( .A(n697), .B(n690), .Z(n716) );
  XNOR U3748 ( .A(n691), .B(n716), .Z(n692) );
  XOR U3749 ( .A(n693), .B(n692), .Z(n729) );
  IV U3750 ( .A(n729), .Z(n735) );
  AND U3751 ( .A(n695), .B(n694), .Z(n700) );
  XOR U3752 ( .A(x[16]), .B(n742), .Z(n743) );
  XNOR U3753 ( .A(n814), .B(n743), .Z(n745) );
  XOR U3754 ( .A(x[18]), .B(x[23]), .Z(n770) );
  NANDN U3755 ( .A(n745), .B(n770), .Z(n696) );
  XNOR U3756 ( .A(n697), .B(n696), .Z(n705) );
  XNOR U3757 ( .A(n698), .B(n705), .Z(n699) );
  XOR U3758 ( .A(n700), .B(n699), .Z(n725) );
  XNOR U3759 ( .A(x[20]), .B(n814), .Z(n763) );
  ANDN U3760 ( .B(x[16]), .A(n763), .Z(n707) );
  XOR U3761 ( .A(x[18]), .B(x[17]), .Z(n701) );
  XOR U3762 ( .A(n778), .B(n701), .Z(n752) );
  XOR U3763 ( .A(n753), .B(n701), .Z(n758) );
  NAND U3764 ( .A(n742), .B(n758), .Z(n709) );
  XNOR U3765 ( .A(n752), .B(n709), .Z(n703) );
  XNOR U3766 ( .A(x[17]), .B(n743), .Z(n702) );
  XNOR U3767 ( .A(n703), .B(n702), .Z(n704) );
  XOR U3768 ( .A(n705), .B(n704), .Z(n706) );
  XOR U3769 ( .A(n707), .B(n706), .Z(n727) );
  NAND U3770 ( .A(n725), .B(n727), .Z(n708) );
  NAND U3771 ( .A(n735), .B(n708), .Z(n719) );
  IV U3772 ( .A(n725), .Z(n726) );
  IV U3773 ( .A(n727), .Z(n733) );
  XOR U3774 ( .A(n709), .B(n763), .Z(n712) );
  AND U3775 ( .A(n752), .B(n743), .Z(n710) );
  XNOR U3776 ( .A(x[16]), .B(n710), .Z(n711) );
  XNOR U3777 ( .A(n712), .B(n711), .Z(n713) );
  XNOR U3778 ( .A(n714), .B(n713), .Z(n715) );
  XNOR U3779 ( .A(n716), .B(n715), .Z(n737) );
  IV U3780 ( .A(n737), .Z(n732) );
  XOR U3781 ( .A(n733), .B(n732), .Z(n717) );
  NAND U3782 ( .A(n726), .B(n717), .Z(n718) );
  AND U3783 ( .A(n719), .B(n718), .Z(n822) );
  NAND U3784 ( .A(n733), .B(n726), .Z(n720) );
  NAND U3785 ( .A(n732), .B(n720), .Z(n723) );
  XOR U3786 ( .A(n726), .B(n729), .Z(n721) );
  NAND U3787 ( .A(n727), .B(n721), .Z(n722) );
  AND U3788 ( .A(n723), .B(n722), .Z(n779) );
  XNOR U3789 ( .A(n822), .B(n779), .Z(n754) );
  OR U3790 ( .A(n754), .B(n724), .Z(n747) );
  NAND U3791 ( .A(n735), .B(n725), .Z(n731) );
  AND U3792 ( .A(n727), .B(n726), .Z(n734) );
  XNOR U3793 ( .A(n732), .B(n734), .Z(n728) );
  NAND U3794 ( .A(n729), .B(n728), .Z(n730) );
  AND U3795 ( .A(n731), .B(n730), .Z(n751) );
  NAND U3796 ( .A(n733), .B(n732), .Z(n739) );
  XNOR U3797 ( .A(n735), .B(n734), .Z(n736) );
  NAND U3798 ( .A(n737), .B(n736), .Z(n738) );
  NAND U3799 ( .A(n739), .B(n738), .Z(n816) );
  XNOR U3800 ( .A(n751), .B(n816), .Z(n769) );
  XOR U3801 ( .A(n769), .B(n754), .Z(n756) );
  OR U3802 ( .A(n756), .B(n740), .Z(n741) );
  XNOR U3803 ( .A(n747), .B(n741), .Z(n773) );
  XOR U3804 ( .A(n751), .B(n822), .Z(n759) );
  NANDN U3805 ( .A(n759), .B(n742), .Z(n824) );
  NANDN U3806 ( .A(n751), .B(n743), .Z(n744) );
  XNOR U3807 ( .A(n824), .B(n744), .Z(n777) );
  XOR U3808 ( .A(n773), .B(n777), .Z(n762) );
  NANDN U3809 ( .A(n745), .B(n769), .Z(n746) );
  XNOR U3810 ( .A(n747), .B(n746), .Z(n830) );
  XNOR U3811 ( .A(n816), .B(n779), .Z(n781) );
  NANDN U3812 ( .A(n781), .B(n748), .Z(n765) );
  NAND U3813 ( .A(n749), .B(n779), .Z(n750) );
  XNOR U3814 ( .A(n765), .B(n750), .Z(n821) );
  XOR U3815 ( .A(n830), .B(n821), .Z(n813) );
  XNOR U3816 ( .A(n762), .B(n813), .Z(z[16]) );
  ANDN U3817 ( .B(n752), .A(n751), .Z(n761) );
  NANDN U3818 ( .A(n754), .B(n753), .Z(n772) );
  NANDN U3819 ( .A(n756), .B(n755), .Z(n757) );
  XNOR U3820 ( .A(n772), .B(n757), .Z(n825) );
  NANDN U3821 ( .A(n759), .B(n758), .Z(n766) );
  XNOR U3822 ( .A(n825), .B(n766), .Z(n760) );
  XOR U3823 ( .A(n761), .B(n760), .Z(n786) );
  XOR U3824 ( .A(n786), .B(n762), .Z(n829) );
  ANDN U3825 ( .B(n822), .A(n763), .Z(n768) );
  NAND U3826 ( .A(n814), .B(n816), .Z(n764) );
  XNOR U3827 ( .A(n765), .B(n764), .Z(n776) );
  XNOR U3828 ( .A(n766), .B(n776), .Z(n767) );
  XNOR U3829 ( .A(n768), .B(n767), .Z(n775) );
  NAND U3830 ( .A(n770), .B(n769), .Z(n771) );
  XNOR U3831 ( .A(n772), .B(n771), .Z(n782) );
  XNOR U3832 ( .A(n773), .B(n782), .Z(n774) );
  XOR U3833 ( .A(n775), .B(n774), .Z(n785) );
  XNOR U3834 ( .A(n829), .B(n785), .Z(z[17]) );
  XNOR U3835 ( .A(n777), .B(n776), .Z(z[18]) );
  AND U3836 ( .A(n779), .B(n778), .Z(n784) );
  NANDN U3837 ( .A(n781), .B(n780), .Z(n819) );
  XNOR U3838 ( .A(n782), .B(n819), .Z(n783) );
  XOR U3839 ( .A(n784), .B(n783), .Z(n828) );
  XOR U3840 ( .A(n786), .B(n785), .Z(n787) );
  XOR U3841 ( .A(n828), .B(n787), .Z(z[19]) );
  ANDN U3842 ( .B(n789), .A(n788), .Z(n798) );
  NANDN U3843 ( .A(n791), .B(n790), .Z(n809) );
  NANDN U3844 ( .A(n793), .B(n792), .Z(n794) );
  XNOR U3845 ( .A(n809), .B(n794), .Z(n1457) );
  NANDN U3846 ( .A(n796), .B(n795), .Z(n803) );
  XNOR U3847 ( .A(n1457), .B(n803), .Z(n797) );
  XOR U3848 ( .A(n798), .B(n797), .Z(n1091) );
  XOR U3849 ( .A(n1091), .B(n799), .Z(n1600) );
  ANDN U3850 ( .B(n1454), .A(n800), .Z(n805) );
  NAND U3851 ( .A(n1446), .B(n1448), .Z(n801) );
  XNOR U3852 ( .A(n802), .B(n801), .Z(n952) );
  XNOR U3853 ( .A(n803), .B(n952), .Z(n804) );
  XNOR U3854 ( .A(n805), .B(n804), .Z(n812) );
  NAND U3855 ( .A(n807), .B(n806), .Z(n808) );
  XNOR U3856 ( .A(n809), .B(n808), .Z(n1087) );
  XNOR U3857 ( .A(n810), .B(n1087), .Z(n811) );
  XOR U3858 ( .A(n812), .B(n811), .Z(n1090) );
  XNOR U3859 ( .A(n1600), .B(n1090), .Z(z[1]) );
  XOR U3860 ( .A(n813), .B(z[18]), .Z(z[20]) );
  XNOR U3861 ( .A(n815), .B(n814), .Z(n817) );
  NAND U3862 ( .A(n817), .B(n816), .Z(n818) );
  XOR U3863 ( .A(n819), .B(n818), .Z(n820) );
  XNOR U3864 ( .A(n821), .B(n820), .Z(n827) );
  NAND U3865 ( .A(n822), .B(x[16]), .Z(n823) );
  XNOR U3866 ( .A(n824), .B(n823), .Z(n831) );
  XNOR U3867 ( .A(n825), .B(n831), .Z(n826) );
  XOR U3868 ( .A(n827), .B(n826), .Z(z[21]) );
  XNOR U3869 ( .A(n829), .B(n828), .Z(z[22]) );
  XNOR U3870 ( .A(n831), .B(n830), .Z(n832) );
  XNOR U3871 ( .A(z[17]), .B(n832), .Z(z[23]) );
  IV U3872 ( .A(x[25]), .Z(n939) );
  XOR U3873 ( .A(x[29]), .B(n834), .Z(n938) );
  IV U3874 ( .A(n938), .Z(n835) );
  AND U3875 ( .A(n939), .B(n835), .Z(n842) );
  XNOR U3876 ( .A(x[27]), .B(n939), .Z(n838) );
  XNOR U3877 ( .A(x[26]), .B(n838), .Z(n833) );
  XNOR U3878 ( .A(n834), .B(n833), .Z(n898) );
  IV U3879 ( .A(n898), .Z(n844) );
  XNOR U3880 ( .A(n844), .B(n938), .Z(n897) );
  IV U3881 ( .A(x[31]), .Z(n836) );
  XNOR U3882 ( .A(x[25]), .B(n836), .Z(n929) );
  NAND U3883 ( .A(n897), .B(n929), .Z(n847) );
  XNOR U3884 ( .A(n836), .B(n835), .Z(n843) );
  IV U3885 ( .A(n843), .Z(n927) );
  XOR U3886 ( .A(n898), .B(n927), .Z(n863) );
  XNOR U3887 ( .A(n847), .B(n863), .Z(n840) );
  XOR U3888 ( .A(x[24]), .B(n844), .Z(n873) );
  XOR U3889 ( .A(x[28]), .B(n836), .Z(n837) );
  IV U3890 ( .A(n837), .Z(n902) );
  NANDN U3891 ( .A(n873), .B(n902), .Z(n846) );
  XNOR U3892 ( .A(n838), .B(n837), .Z(n891) );
  XNOR U3893 ( .A(n897), .B(n891), .Z(n889) );
  XOR U3894 ( .A(x[26]), .B(x[28]), .Z(n904) );
  NANDN U3895 ( .A(n889), .B(n904), .Z(n839) );
  XOR U3896 ( .A(n846), .B(n839), .Z(n865) );
  XNOR U3897 ( .A(n840), .B(n865), .Z(n841) );
  XOR U3898 ( .A(n842), .B(n841), .Z(n878) );
  IV U3899 ( .A(n878), .Z(n884) );
  AND U3900 ( .A(n844), .B(n843), .Z(n849) );
  XOR U3901 ( .A(x[24]), .B(n891), .Z(n892) );
  XNOR U3902 ( .A(n938), .B(n892), .Z(n894) );
  XOR U3903 ( .A(x[26]), .B(x[31]), .Z(n919) );
  NANDN U3904 ( .A(n894), .B(n919), .Z(n845) );
  XNOR U3905 ( .A(n846), .B(n845), .Z(n854) );
  XNOR U3906 ( .A(n847), .B(n854), .Z(n848) );
  XOR U3907 ( .A(n849), .B(n848), .Z(n874) );
  XNOR U3908 ( .A(x[28]), .B(n938), .Z(n912) );
  ANDN U3909 ( .B(x[24]), .A(n912), .Z(n856) );
  XOR U3910 ( .A(x[26]), .B(x[25]), .Z(n850) );
  XOR U3911 ( .A(n927), .B(n850), .Z(n901) );
  XOR U3912 ( .A(n902), .B(n850), .Z(n907) );
  NAND U3913 ( .A(n891), .B(n907), .Z(n858) );
  XNOR U3914 ( .A(n901), .B(n858), .Z(n852) );
  XNOR U3915 ( .A(x[25]), .B(n892), .Z(n851) );
  XNOR U3916 ( .A(n852), .B(n851), .Z(n853) );
  XOR U3917 ( .A(n854), .B(n853), .Z(n855) );
  XOR U3918 ( .A(n856), .B(n855), .Z(n876) );
  NAND U3919 ( .A(n874), .B(n876), .Z(n857) );
  NAND U3920 ( .A(n884), .B(n857), .Z(n868) );
  IV U3921 ( .A(n874), .Z(n875) );
  IV U3922 ( .A(n876), .Z(n882) );
  XOR U3923 ( .A(n858), .B(n912), .Z(n861) );
  AND U3924 ( .A(n901), .B(n892), .Z(n859) );
  XNOR U3925 ( .A(x[24]), .B(n859), .Z(n860) );
  XNOR U3926 ( .A(n861), .B(n860), .Z(n862) );
  XNOR U3927 ( .A(n863), .B(n862), .Z(n864) );
  XNOR U3928 ( .A(n865), .B(n864), .Z(n886) );
  IV U3929 ( .A(n886), .Z(n881) );
  XOR U3930 ( .A(n882), .B(n881), .Z(n866) );
  NAND U3931 ( .A(n875), .B(n866), .Z(n867) );
  AND U3932 ( .A(n868), .B(n867), .Z(n946) );
  NAND U3933 ( .A(n882), .B(n875), .Z(n869) );
  NAND U3934 ( .A(n881), .B(n869), .Z(n872) );
  XOR U3935 ( .A(n875), .B(n878), .Z(n870) );
  NAND U3936 ( .A(n876), .B(n870), .Z(n871) );
  AND U3937 ( .A(n872), .B(n871), .Z(n928) );
  XNOR U3938 ( .A(n946), .B(n928), .Z(n903) );
  OR U3939 ( .A(n903), .B(n873), .Z(n896) );
  NAND U3940 ( .A(n884), .B(n874), .Z(n880) );
  AND U3941 ( .A(n876), .B(n875), .Z(n883) );
  XNOR U3942 ( .A(n881), .B(n883), .Z(n877) );
  NAND U3943 ( .A(n878), .B(n877), .Z(n879) );
  AND U3944 ( .A(n880), .B(n879), .Z(n900) );
  NAND U3945 ( .A(n882), .B(n881), .Z(n888) );
  XNOR U3946 ( .A(n884), .B(n883), .Z(n885) );
  NAND U3947 ( .A(n886), .B(n885), .Z(n887) );
  NAND U3948 ( .A(n888), .B(n887), .Z(n940) );
  XNOR U3949 ( .A(n900), .B(n940), .Z(n918) );
  XOR U3950 ( .A(n918), .B(n903), .Z(n905) );
  OR U3951 ( .A(n905), .B(n889), .Z(n890) );
  XNOR U3952 ( .A(n896), .B(n890), .Z(n922) );
  XOR U3953 ( .A(n900), .B(n946), .Z(n908) );
  NANDN U3954 ( .A(n908), .B(n891), .Z(n948) );
  NANDN U3955 ( .A(n900), .B(n892), .Z(n893) );
  XNOR U3956 ( .A(n948), .B(n893), .Z(n926) );
  XOR U3957 ( .A(n922), .B(n926), .Z(n911) );
  NANDN U3958 ( .A(n894), .B(n918), .Z(n895) );
  XNOR U3959 ( .A(n896), .B(n895), .Z(n956) );
  XNOR U3960 ( .A(n940), .B(n928), .Z(n930) );
  NANDN U3961 ( .A(n930), .B(n897), .Z(n914) );
  NAND U3962 ( .A(n898), .B(n928), .Z(n899) );
  XNOR U3963 ( .A(n914), .B(n899), .Z(n945) );
  XOR U3964 ( .A(n956), .B(n945), .Z(n937) );
  XNOR U3965 ( .A(n911), .B(n937), .Z(z[24]) );
  ANDN U3966 ( .B(n901), .A(n900), .Z(n910) );
  NANDN U3967 ( .A(n903), .B(n902), .Z(n921) );
  NANDN U3968 ( .A(n905), .B(n904), .Z(n906) );
  XNOR U3969 ( .A(n921), .B(n906), .Z(n949) );
  NANDN U3970 ( .A(n908), .B(n907), .Z(n915) );
  XNOR U3971 ( .A(n949), .B(n915), .Z(n909) );
  XOR U3972 ( .A(n910), .B(n909), .Z(n935) );
  XOR U3973 ( .A(n935), .B(n911), .Z(n955) );
  ANDN U3974 ( .B(n946), .A(n912), .Z(n917) );
  NAND U3975 ( .A(n938), .B(n940), .Z(n913) );
  XNOR U3976 ( .A(n914), .B(n913), .Z(n925) );
  XNOR U3977 ( .A(n915), .B(n925), .Z(n916) );
  XNOR U3978 ( .A(n917), .B(n916), .Z(n924) );
  NAND U3979 ( .A(n919), .B(n918), .Z(n920) );
  XNOR U3980 ( .A(n921), .B(n920), .Z(n931) );
  XNOR U3981 ( .A(n922), .B(n931), .Z(n923) );
  XOR U3982 ( .A(n924), .B(n923), .Z(n934) );
  XNOR U3983 ( .A(n955), .B(n934), .Z(z[25]) );
  XNOR U3984 ( .A(n926), .B(n925), .Z(z[26]) );
  AND U3985 ( .A(n928), .B(n927), .Z(n933) );
  NANDN U3986 ( .A(n930), .B(n929), .Z(n943) );
  XNOR U3987 ( .A(n931), .B(n943), .Z(n932) );
  XOR U3988 ( .A(n933), .B(n932), .Z(n954) );
  XOR U3989 ( .A(n935), .B(n934), .Z(n936) );
  XOR U3990 ( .A(n954), .B(n936), .Z(z[27]) );
  XOR U3991 ( .A(n937), .B(z[26]), .Z(z[28]) );
  XNOR U3992 ( .A(n939), .B(n938), .Z(n941) );
  NAND U3993 ( .A(n941), .B(n940), .Z(n942) );
  XOR U3994 ( .A(n943), .B(n942), .Z(n944) );
  XNOR U3995 ( .A(n945), .B(n944), .Z(n951) );
  NAND U3996 ( .A(n946), .B(x[24]), .Z(n947) );
  XNOR U3997 ( .A(n948), .B(n947), .Z(n957) );
  XNOR U3998 ( .A(n949), .B(n957), .Z(n950) );
  XOR U3999 ( .A(n951), .B(n950), .Z(z[29]) );
  XNOR U4000 ( .A(n953), .B(n952), .Z(z[2]) );
  XNOR U4001 ( .A(n955), .B(n954), .Z(z[30]) );
  XNOR U4002 ( .A(n957), .B(n956), .Z(n958) );
  XNOR U4003 ( .A(z[25]), .B(n958), .Z(z[31]) );
  IV U4004 ( .A(x[33]), .Z(n1065) );
  XOR U4005 ( .A(x[32]), .B(x[38]), .Z(n960) );
  XOR U4006 ( .A(x[37]), .B(n960), .Z(n1064) );
  IV U4007 ( .A(n1064), .Z(n961) );
  AND U4008 ( .A(n1065), .B(n961), .Z(n968) );
  XNOR U4009 ( .A(x[35]), .B(n1065), .Z(n964) );
  XNOR U4010 ( .A(x[34]), .B(n964), .Z(n959) );
  XNOR U4011 ( .A(n960), .B(n959), .Z(n1024) );
  IV U4012 ( .A(n1024), .Z(n970) );
  XNOR U4013 ( .A(n970), .B(n1064), .Z(n1023) );
  IV U4014 ( .A(x[39]), .Z(n962) );
  XNOR U4015 ( .A(x[33]), .B(n962), .Z(n1055) );
  NAND U4016 ( .A(n1023), .B(n1055), .Z(n973) );
  XNOR U4017 ( .A(n962), .B(n961), .Z(n969) );
  IV U4018 ( .A(n969), .Z(n1053) );
  XOR U4019 ( .A(n1024), .B(n1053), .Z(n989) );
  XNOR U4020 ( .A(n973), .B(n989), .Z(n966) );
  XOR U4021 ( .A(x[32]), .B(n970), .Z(n999) );
  XOR U4022 ( .A(x[36]), .B(n962), .Z(n963) );
  IV U4023 ( .A(n963), .Z(n1028) );
  NANDN U4024 ( .A(n999), .B(n1028), .Z(n972) );
  XNOR U4025 ( .A(n964), .B(n963), .Z(n1017) );
  XNOR U4026 ( .A(n1023), .B(n1017), .Z(n1015) );
  XOR U4027 ( .A(x[34]), .B(x[36]), .Z(n1030) );
  NANDN U4028 ( .A(n1015), .B(n1030), .Z(n965) );
  XOR U4029 ( .A(n972), .B(n965), .Z(n991) );
  XNOR U4030 ( .A(n966), .B(n991), .Z(n967) );
  XOR U4031 ( .A(n968), .B(n967), .Z(n1004) );
  IV U4032 ( .A(n1004), .Z(n1010) );
  AND U4033 ( .A(n970), .B(n969), .Z(n975) );
  XOR U4034 ( .A(x[32]), .B(n1017), .Z(n1018) );
  XNOR U4035 ( .A(n1064), .B(n1018), .Z(n1020) );
  XOR U4036 ( .A(x[34]), .B(x[39]), .Z(n1045) );
  NANDN U4037 ( .A(n1020), .B(n1045), .Z(n971) );
  XNOR U4038 ( .A(n972), .B(n971), .Z(n980) );
  XNOR U4039 ( .A(n973), .B(n980), .Z(n974) );
  XOR U4040 ( .A(n975), .B(n974), .Z(n1000) );
  XNOR U4041 ( .A(x[36]), .B(n1064), .Z(n1038) );
  ANDN U4042 ( .B(x[32]), .A(n1038), .Z(n982) );
  XOR U4043 ( .A(x[34]), .B(x[33]), .Z(n976) );
  XOR U4044 ( .A(n1053), .B(n976), .Z(n1027) );
  XOR U4045 ( .A(n1028), .B(n976), .Z(n1033) );
  NAND U4046 ( .A(n1017), .B(n1033), .Z(n984) );
  XNOR U4047 ( .A(n1027), .B(n984), .Z(n978) );
  XNOR U4048 ( .A(x[33]), .B(n1018), .Z(n977) );
  XNOR U4049 ( .A(n978), .B(n977), .Z(n979) );
  XOR U4050 ( .A(n980), .B(n979), .Z(n981) );
  XOR U4051 ( .A(n982), .B(n981), .Z(n1002) );
  NAND U4052 ( .A(n1000), .B(n1002), .Z(n983) );
  NAND U4053 ( .A(n1010), .B(n983), .Z(n994) );
  IV U4054 ( .A(n1000), .Z(n1001) );
  IV U4055 ( .A(n1002), .Z(n1008) );
  XOR U4056 ( .A(n984), .B(n1038), .Z(n987) );
  AND U4057 ( .A(n1027), .B(n1018), .Z(n985) );
  XNOR U4058 ( .A(x[32]), .B(n985), .Z(n986) );
  XNOR U4059 ( .A(n987), .B(n986), .Z(n988) );
  XNOR U4060 ( .A(n989), .B(n988), .Z(n990) );
  XNOR U4061 ( .A(n991), .B(n990), .Z(n1012) );
  IV U4062 ( .A(n1012), .Z(n1007) );
  XOR U4063 ( .A(n1008), .B(n1007), .Z(n992) );
  NAND U4064 ( .A(n1001), .B(n992), .Z(n993) );
  AND U4065 ( .A(n994), .B(n993), .Z(n1072) );
  NAND U4066 ( .A(n1008), .B(n1001), .Z(n995) );
  NAND U4067 ( .A(n1007), .B(n995), .Z(n998) );
  XOR U4068 ( .A(n1001), .B(n1004), .Z(n996) );
  NAND U4069 ( .A(n1002), .B(n996), .Z(n997) );
  AND U4070 ( .A(n998), .B(n997), .Z(n1054) );
  XNOR U4071 ( .A(n1072), .B(n1054), .Z(n1029) );
  OR U4072 ( .A(n1029), .B(n999), .Z(n1022) );
  NAND U4073 ( .A(n1010), .B(n1000), .Z(n1006) );
  AND U4074 ( .A(n1002), .B(n1001), .Z(n1009) );
  XNOR U4075 ( .A(n1007), .B(n1009), .Z(n1003) );
  NAND U4076 ( .A(n1004), .B(n1003), .Z(n1005) );
  AND U4077 ( .A(n1006), .B(n1005), .Z(n1026) );
  NAND U4078 ( .A(n1008), .B(n1007), .Z(n1014) );
  XNOR U4079 ( .A(n1010), .B(n1009), .Z(n1011) );
  NAND U4080 ( .A(n1012), .B(n1011), .Z(n1013) );
  NAND U4081 ( .A(n1014), .B(n1013), .Z(n1066) );
  XNOR U4082 ( .A(n1026), .B(n1066), .Z(n1044) );
  XOR U4083 ( .A(n1044), .B(n1029), .Z(n1031) );
  OR U4084 ( .A(n1031), .B(n1015), .Z(n1016) );
  XNOR U4085 ( .A(n1022), .B(n1016), .Z(n1048) );
  XOR U4086 ( .A(n1026), .B(n1072), .Z(n1034) );
  NANDN U4087 ( .A(n1034), .B(n1017), .Z(n1074) );
  NANDN U4088 ( .A(n1026), .B(n1018), .Z(n1019) );
  XNOR U4089 ( .A(n1074), .B(n1019), .Z(n1052) );
  XOR U4090 ( .A(n1048), .B(n1052), .Z(n1037) );
  NANDN U4091 ( .A(n1020), .B(n1044), .Z(n1021) );
  XNOR U4092 ( .A(n1022), .B(n1021), .Z(n1080) );
  XNOR U4093 ( .A(n1066), .B(n1054), .Z(n1056) );
  NANDN U4094 ( .A(n1056), .B(n1023), .Z(n1040) );
  NAND U4095 ( .A(n1024), .B(n1054), .Z(n1025) );
  XNOR U4096 ( .A(n1040), .B(n1025), .Z(n1071) );
  XOR U4097 ( .A(n1080), .B(n1071), .Z(n1063) );
  XNOR U4098 ( .A(n1037), .B(n1063), .Z(z[32]) );
  ANDN U4099 ( .B(n1027), .A(n1026), .Z(n1036) );
  NANDN U4100 ( .A(n1029), .B(n1028), .Z(n1047) );
  NANDN U4101 ( .A(n1031), .B(n1030), .Z(n1032) );
  XNOR U4102 ( .A(n1047), .B(n1032), .Z(n1075) );
  NANDN U4103 ( .A(n1034), .B(n1033), .Z(n1041) );
  XNOR U4104 ( .A(n1075), .B(n1041), .Z(n1035) );
  XOR U4105 ( .A(n1036), .B(n1035), .Z(n1061) );
  XOR U4106 ( .A(n1061), .B(n1037), .Z(n1079) );
  ANDN U4107 ( .B(n1072), .A(n1038), .Z(n1043) );
  NAND U4108 ( .A(n1064), .B(n1066), .Z(n1039) );
  XNOR U4109 ( .A(n1040), .B(n1039), .Z(n1051) );
  XNOR U4110 ( .A(n1041), .B(n1051), .Z(n1042) );
  XNOR U4111 ( .A(n1043), .B(n1042), .Z(n1050) );
  NAND U4112 ( .A(n1045), .B(n1044), .Z(n1046) );
  XNOR U4113 ( .A(n1047), .B(n1046), .Z(n1057) );
  XNOR U4114 ( .A(n1048), .B(n1057), .Z(n1049) );
  XOR U4115 ( .A(n1050), .B(n1049), .Z(n1060) );
  XNOR U4116 ( .A(n1079), .B(n1060), .Z(z[33]) );
  XNOR U4117 ( .A(n1052), .B(n1051), .Z(z[34]) );
  AND U4118 ( .A(n1054), .B(n1053), .Z(n1059) );
  NANDN U4119 ( .A(n1056), .B(n1055), .Z(n1069) );
  XNOR U4120 ( .A(n1057), .B(n1069), .Z(n1058) );
  XOR U4121 ( .A(n1059), .B(n1058), .Z(n1078) );
  XOR U4122 ( .A(n1061), .B(n1060), .Z(n1062) );
  XOR U4123 ( .A(n1078), .B(n1062), .Z(z[35]) );
  XOR U4124 ( .A(n1063), .B(z[34]), .Z(z[36]) );
  XNOR U4125 ( .A(n1065), .B(n1064), .Z(n1067) );
  NAND U4126 ( .A(n1067), .B(n1066), .Z(n1068) );
  XOR U4127 ( .A(n1069), .B(n1068), .Z(n1070) );
  XNOR U4128 ( .A(n1071), .B(n1070), .Z(n1077) );
  NAND U4129 ( .A(n1072), .B(x[32]), .Z(n1073) );
  XNOR U4130 ( .A(n1074), .B(n1073), .Z(n1081) );
  XNOR U4131 ( .A(n1075), .B(n1081), .Z(n1076) );
  XOR U4132 ( .A(n1077), .B(n1076), .Z(z[37]) );
  XNOR U4133 ( .A(n1079), .B(n1078), .Z(z[38]) );
  XNOR U4134 ( .A(n1081), .B(n1080), .Z(n1082) );
  XNOR U4135 ( .A(z[33]), .B(n1082), .Z(z[39]) );
  AND U4136 ( .A(n1084), .B(n1083), .Z(n1089) );
  NANDN U4137 ( .A(n1086), .B(n1085), .Z(n1451) );
  XNOR U4138 ( .A(n1087), .B(n1451), .Z(n1088) );
  XOR U4139 ( .A(n1089), .B(n1088), .Z(n1599) );
  XOR U4140 ( .A(n1091), .B(n1090), .Z(n1092) );
  XOR U4141 ( .A(n1599), .B(n1092), .Z(z[3]) );
  IV U4142 ( .A(x[41]), .Z(n1199) );
  XOR U4143 ( .A(x[40]), .B(x[46]), .Z(n1094) );
  XOR U4144 ( .A(x[45]), .B(n1094), .Z(n1198) );
  IV U4145 ( .A(n1198), .Z(n1095) );
  AND U4146 ( .A(n1199), .B(n1095), .Z(n1102) );
  XNOR U4147 ( .A(x[43]), .B(n1199), .Z(n1098) );
  XNOR U4148 ( .A(x[42]), .B(n1098), .Z(n1093) );
  XNOR U4149 ( .A(n1094), .B(n1093), .Z(n1158) );
  IV U4150 ( .A(n1158), .Z(n1104) );
  XNOR U4151 ( .A(n1104), .B(n1198), .Z(n1157) );
  IV U4152 ( .A(x[47]), .Z(n1096) );
  XNOR U4153 ( .A(x[41]), .B(n1096), .Z(n1189) );
  NAND U4154 ( .A(n1157), .B(n1189), .Z(n1107) );
  XNOR U4155 ( .A(n1096), .B(n1095), .Z(n1103) );
  IV U4156 ( .A(n1103), .Z(n1187) );
  XOR U4157 ( .A(n1158), .B(n1187), .Z(n1123) );
  XNOR U4158 ( .A(n1107), .B(n1123), .Z(n1100) );
  XOR U4159 ( .A(x[40]), .B(n1104), .Z(n1133) );
  XOR U4160 ( .A(x[44]), .B(n1096), .Z(n1097) );
  IV U4161 ( .A(n1097), .Z(n1162) );
  NANDN U4162 ( .A(n1133), .B(n1162), .Z(n1106) );
  XNOR U4163 ( .A(n1098), .B(n1097), .Z(n1151) );
  XNOR U4164 ( .A(n1157), .B(n1151), .Z(n1149) );
  XOR U4165 ( .A(x[42]), .B(x[44]), .Z(n1164) );
  NANDN U4166 ( .A(n1149), .B(n1164), .Z(n1099) );
  XOR U4167 ( .A(n1106), .B(n1099), .Z(n1125) );
  XNOR U4168 ( .A(n1100), .B(n1125), .Z(n1101) );
  XOR U4169 ( .A(n1102), .B(n1101), .Z(n1138) );
  IV U4170 ( .A(n1138), .Z(n1144) );
  AND U4171 ( .A(n1104), .B(n1103), .Z(n1109) );
  XOR U4172 ( .A(x[40]), .B(n1151), .Z(n1152) );
  XNOR U4173 ( .A(n1198), .B(n1152), .Z(n1154) );
  XOR U4174 ( .A(x[42]), .B(x[47]), .Z(n1179) );
  NANDN U4175 ( .A(n1154), .B(n1179), .Z(n1105) );
  XNOR U4176 ( .A(n1106), .B(n1105), .Z(n1114) );
  XNOR U4177 ( .A(n1107), .B(n1114), .Z(n1108) );
  XOR U4178 ( .A(n1109), .B(n1108), .Z(n1134) );
  XNOR U4179 ( .A(x[44]), .B(n1198), .Z(n1172) );
  ANDN U4180 ( .B(x[40]), .A(n1172), .Z(n1116) );
  XOR U4181 ( .A(x[42]), .B(x[41]), .Z(n1110) );
  XOR U4182 ( .A(n1187), .B(n1110), .Z(n1161) );
  XOR U4183 ( .A(n1162), .B(n1110), .Z(n1167) );
  NAND U4184 ( .A(n1151), .B(n1167), .Z(n1118) );
  XNOR U4185 ( .A(n1161), .B(n1118), .Z(n1112) );
  XNOR U4186 ( .A(x[41]), .B(n1152), .Z(n1111) );
  XNOR U4187 ( .A(n1112), .B(n1111), .Z(n1113) );
  XOR U4188 ( .A(n1114), .B(n1113), .Z(n1115) );
  XOR U4189 ( .A(n1116), .B(n1115), .Z(n1136) );
  NAND U4190 ( .A(n1134), .B(n1136), .Z(n1117) );
  NAND U4191 ( .A(n1144), .B(n1117), .Z(n1128) );
  IV U4192 ( .A(n1134), .Z(n1135) );
  IV U4193 ( .A(n1136), .Z(n1142) );
  XOR U4194 ( .A(n1118), .B(n1172), .Z(n1121) );
  AND U4195 ( .A(n1161), .B(n1152), .Z(n1119) );
  XNOR U4196 ( .A(x[40]), .B(n1119), .Z(n1120) );
  XNOR U4197 ( .A(n1121), .B(n1120), .Z(n1122) );
  XNOR U4198 ( .A(n1123), .B(n1122), .Z(n1124) );
  XNOR U4199 ( .A(n1125), .B(n1124), .Z(n1146) );
  IV U4200 ( .A(n1146), .Z(n1141) );
  XOR U4201 ( .A(n1142), .B(n1141), .Z(n1126) );
  NAND U4202 ( .A(n1135), .B(n1126), .Z(n1127) );
  AND U4203 ( .A(n1128), .B(n1127), .Z(n1206) );
  NAND U4204 ( .A(n1142), .B(n1135), .Z(n1129) );
  NAND U4205 ( .A(n1141), .B(n1129), .Z(n1132) );
  XOR U4206 ( .A(n1135), .B(n1138), .Z(n1130) );
  NAND U4207 ( .A(n1136), .B(n1130), .Z(n1131) );
  AND U4208 ( .A(n1132), .B(n1131), .Z(n1188) );
  XNOR U4209 ( .A(n1206), .B(n1188), .Z(n1163) );
  OR U4210 ( .A(n1163), .B(n1133), .Z(n1156) );
  NAND U4211 ( .A(n1144), .B(n1134), .Z(n1140) );
  AND U4212 ( .A(n1136), .B(n1135), .Z(n1143) );
  XNOR U4213 ( .A(n1141), .B(n1143), .Z(n1137) );
  NAND U4214 ( .A(n1138), .B(n1137), .Z(n1139) );
  AND U4215 ( .A(n1140), .B(n1139), .Z(n1160) );
  NAND U4216 ( .A(n1142), .B(n1141), .Z(n1148) );
  XNOR U4217 ( .A(n1144), .B(n1143), .Z(n1145) );
  NAND U4218 ( .A(n1146), .B(n1145), .Z(n1147) );
  NAND U4219 ( .A(n1148), .B(n1147), .Z(n1200) );
  XNOR U4220 ( .A(n1160), .B(n1200), .Z(n1178) );
  XOR U4221 ( .A(n1178), .B(n1163), .Z(n1165) );
  OR U4222 ( .A(n1165), .B(n1149), .Z(n1150) );
  XNOR U4223 ( .A(n1156), .B(n1150), .Z(n1182) );
  XOR U4224 ( .A(n1160), .B(n1206), .Z(n1168) );
  NANDN U4225 ( .A(n1168), .B(n1151), .Z(n1208) );
  NANDN U4226 ( .A(n1160), .B(n1152), .Z(n1153) );
  XNOR U4227 ( .A(n1208), .B(n1153), .Z(n1186) );
  XOR U4228 ( .A(n1182), .B(n1186), .Z(n1171) );
  NANDN U4229 ( .A(n1154), .B(n1178), .Z(n1155) );
  XNOR U4230 ( .A(n1156), .B(n1155), .Z(n1214) );
  XNOR U4231 ( .A(n1200), .B(n1188), .Z(n1190) );
  NANDN U4232 ( .A(n1190), .B(n1157), .Z(n1174) );
  NAND U4233 ( .A(n1158), .B(n1188), .Z(n1159) );
  XNOR U4234 ( .A(n1174), .B(n1159), .Z(n1205) );
  XOR U4235 ( .A(n1214), .B(n1205), .Z(n1197) );
  XNOR U4236 ( .A(n1171), .B(n1197), .Z(z[40]) );
  ANDN U4237 ( .B(n1161), .A(n1160), .Z(n1170) );
  NANDN U4238 ( .A(n1163), .B(n1162), .Z(n1181) );
  NANDN U4239 ( .A(n1165), .B(n1164), .Z(n1166) );
  XNOR U4240 ( .A(n1181), .B(n1166), .Z(n1209) );
  NANDN U4241 ( .A(n1168), .B(n1167), .Z(n1175) );
  XNOR U4242 ( .A(n1209), .B(n1175), .Z(n1169) );
  XOR U4243 ( .A(n1170), .B(n1169), .Z(n1195) );
  XOR U4244 ( .A(n1195), .B(n1171), .Z(n1213) );
  ANDN U4245 ( .B(n1206), .A(n1172), .Z(n1177) );
  NAND U4246 ( .A(n1198), .B(n1200), .Z(n1173) );
  XNOR U4247 ( .A(n1174), .B(n1173), .Z(n1185) );
  XNOR U4248 ( .A(n1175), .B(n1185), .Z(n1176) );
  XNOR U4249 ( .A(n1177), .B(n1176), .Z(n1184) );
  NAND U4250 ( .A(n1179), .B(n1178), .Z(n1180) );
  XNOR U4251 ( .A(n1181), .B(n1180), .Z(n1191) );
  XNOR U4252 ( .A(n1182), .B(n1191), .Z(n1183) );
  XOR U4253 ( .A(n1184), .B(n1183), .Z(n1194) );
  XNOR U4254 ( .A(n1213), .B(n1194), .Z(z[41]) );
  XNOR U4255 ( .A(n1186), .B(n1185), .Z(z[42]) );
  AND U4256 ( .A(n1188), .B(n1187), .Z(n1193) );
  NANDN U4257 ( .A(n1190), .B(n1189), .Z(n1203) );
  XNOR U4258 ( .A(n1191), .B(n1203), .Z(n1192) );
  XOR U4259 ( .A(n1193), .B(n1192), .Z(n1212) );
  XOR U4260 ( .A(n1195), .B(n1194), .Z(n1196) );
  XOR U4261 ( .A(n1212), .B(n1196), .Z(z[43]) );
  XOR U4262 ( .A(n1197), .B(z[42]), .Z(z[44]) );
  XNOR U4263 ( .A(n1199), .B(n1198), .Z(n1201) );
  NAND U4264 ( .A(n1201), .B(n1200), .Z(n1202) );
  XOR U4265 ( .A(n1203), .B(n1202), .Z(n1204) );
  XNOR U4266 ( .A(n1205), .B(n1204), .Z(n1211) );
  NAND U4267 ( .A(n1206), .B(x[40]), .Z(n1207) );
  XNOR U4268 ( .A(n1208), .B(n1207), .Z(n1215) );
  XNOR U4269 ( .A(n1209), .B(n1215), .Z(n1210) );
  XOR U4270 ( .A(n1211), .B(n1210), .Z(z[45]) );
  XNOR U4271 ( .A(n1213), .B(n1212), .Z(z[46]) );
  XNOR U4272 ( .A(n1215), .B(n1214), .Z(n1216) );
  XNOR U4273 ( .A(z[41]), .B(n1216), .Z(z[47]) );
  IV U4274 ( .A(x[49]), .Z(n1324) );
  XOR U4275 ( .A(x[48]), .B(x[54]), .Z(n1218) );
  IV U4276 ( .A(n1323), .Z(n1219) );
  AND U4277 ( .A(n1324), .B(n1219), .Z(n1226) );
  XNOR U4278 ( .A(x[50]), .B(n1222), .Z(n1217) );
  XNOR U4279 ( .A(n1218), .B(n1217), .Z(n1282) );
  IV U4280 ( .A(n1282), .Z(n1228) );
  XNOR U4281 ( .A(n1228), .B(n1323), .Z(n1281) );
  IV U4282 ( .A(x[55]), .Z(n1220) );
  XNOR U4283 ( .A(x[49]), .B(n1220), .Z(n1314) );
  NAND U4284 ( .A(n1281), .B(n1314), .Z(n1231) );
  XNOR U4285 ( .A(n1220), .B(n1219), .Z(n1227) );
  IV U4286 ( .A(n1227), .Z(n1312) );
  XOR U4287 ( .A(n1282), .B(n1312), .Z(n1247) );
  XNOR U4288 ( .A(n1231), .B(n1247), .Z(n1224) );
  XOR U4289 ( .A(x[48]), .B(n1228), .Z(n1257) );
  XOR U4290 ( .A(x[52]), .B(n1220), .Z(n1221) );
  IV U4291 ( .A(n1221), .Z(n1286) );
  NANDN U4292 ( .A(n1257), .B(n1286), .Z(n1230) );
  XNOR U4293 ( .A(n1222), .B(n1221), .Z(n1275) );
  XNOR U4294 ( .A(n1281), .B(n1275), .Z(n1273) );
  XOR U4295 ( .A(x[50]), .B(x[52]), .Z(n1288) );
  NANDN U4296 ( .A(n1273), .B(n1288), .Z(n1223) );
  XOR U4297 ( .A(n1230), .B(n1223), .Z(n1249) );
  XNOR U4298 ( .A(n1224), .B(n1249), .Z(n1225) );
  XOR U4299 ( .A(n1226), .B(n1225), .Z(n1262) );
  IV U4300 ( .A(n1262), .Z(n1268) );
  AND U4301 ( .A(n1228), .B(n1227), .Z(n1233) );
  XOR U4302 ( .A(x[48]), .B(n1275), .Z(n1276) );
  XNOR U4303 ( .A(n1323), .B(n1276), .Z(n1278) );
  XOR U4304 ( .A(x[50]), .B(x[55]), .Z(n1303) );
  NANDN U4305 ( .A(n1278), .B(n1303), .Z(n1229) );
  XNOR U4306 ( .A(n1230), .B(n1229), .Z(n1238) );
  XNOR U4307 ( .A(n1231), .B(n1238), .Z(n1232) );
  XOR U4308 ( .A(n1233), .B(n1232), .Z(n1258) );
  XNOR U4309 ( .A(x[52]), .B(n1323), .Z(n1296) );
  ANDN U4310 ( .B(x[48]), .A(n1296), .Z(n1240) );
  XOR U4311 ( .A(x[50]), .B(x[49]), .Z(n1234) );
  XOR U4312 ( .A(n1312), .B(n1234), .Z(n1285) );
  XOR U4313 ( .A(n1286), .B(n1234), .Z(n1291) );
  NAND U4314 ( .A(n1275), .B(n1291), .Z(n1242) );
  XNOR U4315 ( .A(n1285), .B(n1242), .Z(n1236) );
  XNOR U4316 ( .A(x[49]), .B(n1276), .Z(n1235) );
  XNOR U4317 ( .A(n1236), .B(n1235), .Z(n1237) );
  XOR U4318 ( .A(n1238), .B(n1237), .Z(n1239) );
  XOR U4319 ( .A(n1240), .B(n1239), .Z(n1260) );
  NAND U4320 ( .A(n1258), .B(n1260), .Z(n1241) );
  NAND U4321 ( .A(n1268), .B(n1241), .Z(n1252) );
  IV U4322 ( .A(n1258), .Z(n1259) );
  IV U4323 ( .A(n1260), .Z(n1266) );
  XOR U4324 ( .A(n1242), .B(n1296), .Z(n1245) );
  AND U4325 ( .A(n1285), .B(n1276), .Z(n1243) );
  XNOR U4326 ( .A(x[48]), .B(n1243), .Z(n1244) );
  XNOR U4327 ( .A(n1245), .B(n1244), .Z(n1246) );
  XNOR U4328 ( .A(n1247), .B(n1246), .Z(n1248) );
  XNOR U4329 ( .A(n1249), .B(n1248), .Z(n1270) );
  IV U4330 ( .A(n1270), .Z(n1265) );
  XOR U4331 ( .A(n1266), .B(n1265), .Z(n1250) );
  NAND U4332 ( .A(n1259), .B(n1250), .Z(n1251) );
  AND U4333 ( .A(n1252), .B(n1251), .Z(n1331) );
  NAND U4334 ( .A(n1266), .B(n1259), .Z(n1253) );
  NAND U4335 ( .A(n1265), .B(n1253), .Z(n1256) );
  XOR U4336 ( .A(n1259), .B(n1262), .Z(n1254) );
  NAND U4337 ( .A(n1260), .B(n1254), .Z(n1255) );
  AND U4338 ( .A(n1256), .B(n1255), .Z(n1313) );
  XNOR U4339 ( .A(n1331), .B(n1313), .Z(n1287) );
  OR U4340 ( .A(n1287), .B(n1257), .Z(n1280) );
  NAND U4341 ( .A(n1268), .B(n1258), .Z(n1264) );
  AND U4342 ( .A(n1260), .B(n1259), .Z(n1267) );
  XNOR U4343 ( .A(n1265), .B(n1267), .Z(n1261) );
  NAND U4344 ( .A(n1262), .B(n1261), .Z(n1263) );
  AND U4345 ( .A(n1264), .B(n1263), .Z(n1284) );
  NAND U4346 ( .A(n1266), .B(n1265), .Z(n1272) );
  XNOR U4347 ( .A(n1268), .B(n1267), .Z(n1269) );
  NAND U4348 ( .A(n1270), .B(n1269), .Z(n1271) );
  NAND U4349 ( .A(n1272), .B(n1271), .Z(n1325) );
  XNOR U4350 ( .A(n1284), .B(n1325), .Z(n1302) );
  XOR U4351 ( .A(n1302), .B(n1287), .Z(n1289) );
  OR U4352 ( .A(n1289), .B(n1273), .Z(n1274) );
  XNOR U4353 ( .A(n1280), .B(n1274), .Z(n1306) );
  XOR U4354 ( .A(n1284), .B(n1331), .Z(n1292) );
  NANDN U4355 ( .A(n1292), .B(n1275), .Z(n1333) );
  NANDN U4356 ( .A(n1284), .B(n1276), .Z(n1277) );
  XNOR U4357 ( .A(n1333), .B(n1277), .Z(n1311) );
  XOR U4358 ( .A(n1306), .B(n1311), .Z(n1295) );
  NANDN U4359 ( .A(n1278), .B(n1302), .Z(n1279) );
  XNOR U4360 ( .A(n1280), .B(n1279), .Z(n1339) );
  XNOR U4361 ( .A(n1325), .B(n1313), .Z(n1315) );
  NANDN U4362 ( .A(n1315), .B(n1281), .Z(n1298) );
  NAND U4363 ( .A(n1282), .B(n1313), .Z(n1283) );
  XNOR U4364 ( .A(n1298), .B(n1283), .Z(n1330) );
  XOR U4365 ( .A(n1339), .B(n1330), .Z(n1322) );
  XNOR U4366 ( .A(n1295), .B(n1322), .Z(z[48]) );
  ANDN U4367 ( .B(n1285), .A(n1284), .Z(n1294) );
  NANDN U4368 ( .A(n1287), .B(n1286), .Z(n1305) );
  NANDN U4369 ( .A(n1289), .B(n1288), .Z(n1290) );
  XNOR U4370 ( .A(n1305), .B(n1290), .Z(n1334) );
  NANDN U4371 ( .A(n1292), .B(n1291), .Z(n1299) );
  XNOR U4372 ( .A(n1334), .B(n1299), .Z(n1293) );
  XOR U4373 ( .A(n1294), .B(n1293), .Z(n1320) );
  XOR U4374 ( .A(n1320), .B(n1295), .Z(n1338) );
  ANDN U4375 ( .B(n1331), .A(n1296), .Z(n1301) );
  NAND U4376 ( .A(n1323), .B(n1325), .Z(n1297) );
  XNOR U4377 ( .A(n1298), .B(n1297), .Z(n1310) );
  XNOR U4378 ( .A(n1299), .B(n1310), .Z(n1300) );
  XNOR U4379 ( .A(n1301), .B(n1300), .Z(n1308) );
  NAND U4380 ( .A(n1303), .B(n1302), .Z(n1304) );
  XNOR U4381 ( .A(n1305), .B(n1304), .Z(n1316) );
  XNOR U4382 ( .A(n1306), .B(n1316), .Z(n1307) );
  XOR U4383 ( .A(n1308), .B(n1307), .Z(n1319) );
  XNOR U4384 ( .A(n1338), .B(n1319), .Z(z[49]) );
  XOR U4385 ( .A(n1309), .B(z[2]), .Z(z[4]) );
  XNOR U4386 ( .A(n1311), .B(n1310), .Z(z[50]) );
  AND U4387 ( .A(n1313), .B(n1312), .Z(n1318) );
  NANDN U4388 ( .A(n1315), .B(n1314), .Z(n1328) );
  XNOR U4389 ( .A(n1316), .B(n1328), .Z(n1317) );
  XOR U4390 ( .A(n1318), .B(n1317), .Z(n1337) );
  XOR U4391 ( .A(n1320), .B(n1319), .Z(n1321) );
  XOR U4392 ( .A(n1337), .B(n1321), .Z(z[51]) );
  XOR U4393 ( .A(n1322), .B(z[50]), .Z(z[52]) );
  XNOR U4394 ( .A(n1324), .B(n1323), .Z(n1326) );
  NAND U4395 ( .A(n1326), .B(n1325), .Z(n1327) );
  XOR U4396 ( .A(n1328), .B(n1327), .Z(n1329) );
  XNOR U4397 ( .A(n1330), .B(n1329), .Z(n1336) );
  NAND U4398 ( .A(n1331), .B(x[48]), .Z(n1332) );
  XNOR U4399 ( .A(n1333), .B(n1332), .Z(n1340) );
  XNOR U4400 ( .A(n1334), .B(n1340), .Z(n1335) );
  XOR U4401 ( .A(n1336), .B(n1335), .Z(z[53]) );
  XNOR U4402 ( .A(n1338), .B(n1337), .Z(z[54]) );
  XNOR U4403 ( .A(n1340), .B(n1339), .Z(n1341) );
  XNOR U4404 ( .A(z[49]), .B(n1341), .Z(z[55]) );
  IV U4405 ( .A(x[57]), .Z(n1462) );
  XOR U4406 ( .A(x[56]), .B(x[62]), .Z(n1343) );
  XOR U4407 ( .A(x[61]), .B(n1343), .Z(n1461) );
  IV U4408 ( .A(n1461), .Z(n1344) );
  AND U4409 ( .A(n1462), .B(n1344), .Z(n1351) );
  XNOR U4410 ( .A(x[59]), .B(n1462), .Z(n1347) );
  XNOR U4411 ( .A(x[58]), .B(n1347), .Z(n1342) );
  XNOR U4412 ( .A(n1343), .B(n1342), .Z(n1407) );
  IV U4413 ( .A(n1407), .Z(n1353) );
  XNOR U4414 ( .A(n1353), .B(n1461), .Z(n1406) );
  IV U4415 ( .A(x[63]), .Z(n1345) );
  XNOR U4416 ( .A(x[57]), .B(n1345), .Z(n1438) );
  NAND U4417 ( .A(n1406), .B(n1438), .Z(n1356) );
  XNOR U4418 ( .A(n1345), .B(n1344), .Z(n1352) );
  IV U4419 ( .A(n1352), .Z(n1436) );
  XOR U4420 ( .A(n1407), .B(n1436), .Z(n1372) );
  XNOR U4421 ( .A(n1356), .B(n1372), .Z(n1349) );
  XOR U4422 ( .A(x[56]), .B(n1353), .Z(n1382) );
  XOR U4423 ( .A(x[60]), .B(n1345), .Z(n1346) );
  IV U4424 ( .A(n1346), .Z(n1411) );
  NANDN U4425 ( .A(n1382), .B(n1411), .Z(n1355) );
  XNOR U4426 ( .A(n1347), .B(n1346), .Z(n1400) );
  XNOR U4427 ( .A(n1406), .B(n1400), .Z(n1398) );
  XOR U4428 ( .A(x[58]), .B(x[60]), .Z(n1413) );
  NANDN U4429 ( .A(n1398), .B(n1413), .Z(n1348) );
  XOR U4430 ( .A(n1355), .B(n1348), .Z(n1374) );
  XNOR U4431 ( .A(n1349), .B(n1374), .Z(n1350) );
  XOR U4432 ( .A(n1351), .B(n1350), .Z(n1387) );
  IV U4433 ( .A(n1387), .Z(n1393) );
  AND U4434 ( .A(n1353), .B(n1352), .Z(n1358) );
  XOR U4435 ( .A(x[56]), .B(n1400), .Z(n1401) );
  XNOR U4436 ( .A(n1461), .B(n1401), .Z(n1403) );
  XOR U4437 ( .A(x[58]), .B(x[63]), .Z(n1428) );
  NANDN U4438 ( .A(n1403), .B(n1428), .Z(n1354) );
  XNOR U4439 ( .A(n1355), .B(n1354), .Z(n1363) );
  XNOR U4440 ( .A(n1356), .B(n1363), .Z(n1357) );
  XOR U4441 ( .A(n1358), .B(n1357), .Z(n1383) );
  XNOR U4442 ( .A(x[60]), .B(n1461), .Z(n1421) );
  ANDN U4443 ( .B(x[56]), .A(n1421), .Z(n1365) );
  XOR U4444 ( .A(x[58]), .B(x[57]), .Z(n1359) );
  XOR U4445 ( .A(n1436), .B(n1359), .Z(n1410) );
  XOR U4446 ( .A(n1411), .B(n1359), .Z(n1416) );
  NAND U4447 ( .A(n1400), .B(n1416), .Z(n1367) );
  XNOR U4448 ( .A(n1410), .B(n1367), .Z(n1361) );
  XNOR U4449 ( .A(x[57]), .B(n1401), .Z(n1360) );
  XNOR U4450 ( .A(n1361), .B(n1360), .Z(n1362) );
  XOR U4451 ( .A(n1363), .B(n1362), .Z(n1364) );
  XOR U4452 ( .A(n1365), .B(n1364), .Z(n1385) );
  NAND U4453 ( .A(n1383), .B(n1385), .Z(n1366) );
  NAND U4454 ( .A(n1393), .B(n1366), .Z(n1377) );
  IV U4455 ( .A(n1383), .Z(n1384) );
  IV U4456 ( .A(n1385), .Z(n1391) );
  XOR U4457 ( .A(n1367), .B(n1421), .Z(n1370) );
  AND U4458 ( .A(n1410), .B(n1401), .Z(n1368) );
  XNOR U4459 ( .A(x[56]), .B(n1368), .Z(n1369) );
  XNOR U4460 ( .A(n1370), .B(n1369), .Z(n1371) );
  XNOR U4461 ( .A(n1372), .B(n1371), .Z(n1373) );
  XNOR U4462 ( .A(n1374), .B(n1373), .Z(n1395) );
  IV U4463 ( .A(n1395), .Z(n1390) );
  XOR U4464 ( .A(n1391), .B(n1390), .Z(n1375) );
  NAND U4465 ( .A(n1384), .B(n1375), .Z(n1376) );
  AND U4466 ( .A(n1377), .B(n1376), .Z(n1469) );
  NAND U4467 ( .A(n1391), .B(n1384), .Z(n1378) );
  NAND U4468 ( .A(n1390), .B(n1378), .Z(n1381) );
  XOR U4469 ( .A(n1384), .B(n1387), .Z(n1379) );
  NAND U4470 ( .A(n1385), .B(n1379), .Z(n1380) );
  AND U4471 ( .A(n1381), .B(n1380), .Z(n1437) );
  XNOR U4472 ( .A(n1469), .B(n1437), .Z(n1412) );
  OR U4473 ( .A(n1412), .B(n1382), .Z(n1405) );
  NAND U4474 ( .A(n1393), .B(n1383), .Z(n1389) );
  AND U4475 ( .A(n1385), .B(n1384), .Z(n1392) );
  XNOR U4476 ( .A(n1390), .B(n1392), .Z(n1386) );
  NAND U4477 ( .A(n1387), .B(n1386), .Z(n1388) );
  AND U4478 ( .A(n1389), .B(n1388), .Z(n1409) );
  NAND U4479 ( .A(n1391), .B(n1390), .Z(n1397) );
  XNOR U4480 ( .A(n1393), .B(n1392), .Z(n1394) );
  NAND U4481 ( .A(n1395), .B(n1394), .Z(n1396) );
  NAND U4482 ( .A(n1397), .B(n1396), .Z(n1463) );
  XNOR U4483 ( .A(n1409), .B(n1463), .Z(n1427) );
  XOR U4484 ( .A(n1427), .B(n1412), .Z(n1414) );
  OR U4485 ( .A(n1414), .B(n1398), .Z(n1399) );
  XNOR U4486 ( .A(n1405), .B(n1399), .Z(n1431) );
  XOR U4487 ( .A(n1409), .B(n1469), .Z(n1417) );
  NANDN U4488 ( .A(n1417), .B(n1400), .Z(n1471) );
  NANDN U4489 ( .A(n1409), .B(n1401), .Z(n1402) );
  XNOR U4490 ( .A(n1471), .B(n1402), .Z(n1435) );
  XOR U4491 ( .A(n1431), .B(n1435), .Z(n1420) );
  NANDN U4492 ( .A(n1403), .B(n1427), .Z(n1404) );
  XNOR U4493 ( .A(n1405), .B(n1404), .Z(n1477) );
  XNOR U4494 ( .A(n1463), .B(n1437), .Z(n1439) );
  NANDN U4495 ( .A(n1439), .B(n1406), .Z(n1423) );
  NAND U4496 ( .A(n1407), .B(n1437), .Z(n1408) );
  XNOR U4497 ( .A(n1423), .B(n1408), .Z(n1468) );
  XOR U4498 ( .A(n1477), .B(n1468), .Z(n1460) );
  XNOR U4499 ( .A(n1420), .B(n1460), .Z(z[56]) );
  ANDN U4500 ( .B(n1410), .A(n1409), .Z(n1419) );
  NANDN U4501 ( .A(n1412), .B(n1411), .Z(n1430) );
  NANDN U4502 ( .A(n1414), .B(n1413), .Z(n1415) );
  XNOR U4503 ( .A(n1430), .B(n1415), .Z(n1472) );
  NANDN U4504 ( .A(n1417), .B(n1416), .Z(n1424) );
  XNOR U4505 ( .A(n1472), .B(n1424), .Z(n1418) );
  XOR U4506 ( .A(n1419), .B(n1418), .Z(n1444) );
  XOR U4507 ( .A(n1444), .B(n1420), .Z(n1476) );
  ANDN U4508 ( .B(n1469), .A(n1421), .Z(n1426) );
  NAND U4509 ( .A(n1461), .B(n1463), .Z(n1422) );
  XNOR U4510 ( .A(n1423), .B(n1422), .Z(n1434) );
  XNOR U4511 ( .A(n1424), .B(n1434), .Z(n1425) );
  XNOR U4512 ( .A(n1426), .B(n1425), .Z(n1433) );
  NAND U4513 ( .A(n1428), .B(n1427), .Z(n1429) );
  XNOR U4514 ( .A(n1430), .B(n1429), .Z(n1440) );
  XNOR U4515 ( .A(n1431), .B(n1440), .Z(n1432) );
  XOR U4516 ( .A(n1433), .B(n1432), .Z(n1443) );
  XNOR U4517 ( .A(n1476), .B(n1443), .Z(z[57]) );
  XNOR U4518 ( .A(n1435), .B(n1434), .Z(z[58]) );
  AND U4519 ( .A(n1437), .B(n1436), .Z(n1442) );
  NANDN U4520 ( .A(n1439), .B(n1438), .Z(n1466) );
  XNOR U4521 ( .A(n1440), .B(n1466), .Z(n1441) );
  XOR U4522 ( .A(n1442), .B(n1441), .Z(n1475) );
  XOR U4523 ( .A(n1444), .B(n1443), .Z(n1445) );
  XOR U4524 ( .A(n1475), .B(n1445), .Z(z[59]) );
  XNOR U4525 ( .A(n1447), .B(n1446), .Z(n1449) );
  NAND U4526 ( .A(n1449), .B(n1448), .Z(n1450) );
  XOR U4527 ( .A(n1451), .B(n1450), .Z(n1452) );
  XNOR U4528 ( .A(n1453), .B(n1452), .Z(n1459) );
  NAND U4529 ( .A(n1454), .B(x[0]), .Z(n1455) );
  XNOR U4530 ( .A(n1456), .B(n1455), .Z(n1731) );
  XNOR U4531 ( .A(n1457), .B(n1731), .Z(n1458) );
  XOR U4532 ( .A(n1459), .B(n1458), .Z(z[5]) );
  XOR U4533 ( .A(n1460), .B(z[58]), .Z(z[60]) );
  XNOR U4534 ( .A(n1462), .B(n1461), .Z(n1464) );
  NAND U4535 ( .A(n1464), .B(n1463), .Z(n1465) );
  XOR U4536 ( .A(n1466), .B(n1465), .Z(n1467) );
  XNOR U4537 ( .A(n1468), .B(n1467), .Z(n1474) );
  NAND U4538 ( .A(n1469), .B(x[56]), .Z(n1470) );
  XNOR U4539 ( .A(n1471), .B(n1470), .Z(n1478) );
  XNOR U4540 ( .A(n1472), .B(n1478), .Z(n1473) );
  XOR U4541 ( .A(n1474), .B(n1473), .Z(z[61]) );
  XNOR U4542 ( .A(n1476), .B(n1475), .Z(z[62]) );
  XNOR U4543 ( .A(n1478), .B(n1477), .Z(n1479) );
  XNOR U4544 ( .A(z[57]), .B(n1479), .Z(z[63]) );
  IV U4545 ( .A(x[65]), .Z(n1586) );
  XOR U4546 ( .A(x[64]), .B(x[70]), .Z(n1481) );
  XOR U4547 ( .A(x[69]), .B(n1481), .Z(n1585) );
  IV U4548 ( .A(n1585), .Z(n1482) );
  AND U4549 ( .A(n1586), .B(n1482), .Z(n1489) );
  XNOR U4550 ( .A(x[67]), .B(n1586), .Z(n1485) );
  XNOR U4551 ( .A(x[66]), .B(n1485), .Z(n1480) );
  XNOR U4552 ( .A(n1481), .B(n1480), .Z(n1545) );
  IV U4553 ( .A(n1545), .Z(n1491) );
  XNOR U4554 ( .A(n1491), .B(n1585), .Z(n1544) );
  IV U4555 ( .A(x[71]), .Z(n1483) );
  XNOR U4556 ( .A(x[65]), .B(n1483), .Z(n1576) );
  NAND U4557 ( .A(n1544), .B(n1576), .Z(n1494) );
  XNOR U4558 ( .A(n1483), .B(n1482), .Z(n1490) );
  IV U4559 ( .A(n1490), .Z(n1574) );
  XOR U4560 ( .A(n1545), .B(n1574), .Z(n1510) );
  XNOR U4561 ( .A(n1494), .B(n1510), .Z(n1487) );
  XOR U4562 ( .A(x[64]), .B(n1491), .Z(n1520) );
  XOR U4563 ( .A(x[68]), .B(n1483), .Z(n1484) );
  IV U4564 ( .A(n1484), .Z(n1549) );
  NANDN U4565 ( .A(n1520), .B(n1549), .Z(n1493) );
  XNOR U4566 ( .A(n1485), .B(n1484), .Z(n1538) );
  XNOR U4567 ( .A(n1544), .B(n1538), .Z(n1536) );
  XOR U4568 ( .A(x[66]), .B(x[68]), .Z(n1551) );
  NANDN U4569 ( .A(n1536), .B(n1551), .Z(n1486) );
  XOR U4570 ( .A(n1493), .B(n1486), .Z(n1512) );
  XNOR U4571 ( .A(n1487), .B(n1512), .Z(n1488) );
  XOR U4572 ( .A(n1489), .B(n1488), .Z(n1525) );
  IV U4573 ( .A(n1525), .Z(n1531) );
  AND U4574 ( .A(n1491), .B(n1490), .Z(n1496) );
  XOR U4575 ( .A(x[64]), .B(n1538), .Z(n1539) );
  XNOR U4576 ( .A(n1585), .B(n1539), .Z(n1541) );
  XOR U4577 ( .A(x[66]), .B(x[71]), .Z(n1566) );
  NANDN U4578 ( .A(n1541), .B(n1566), .Z(n1492) );
  XNOR U4579 ( .A(n1493), .B(n1492), .Z(n1501) );
  XNOR U4580 ( .A(n1494), .B(n1501), .Z(n1495) );
  XOR U4581 ( .A(n1496), .B(n1495), .Z(n1521) );
  XNOR U4582 ( .A(x[68]), .B(n1585), .Z(n1559) );
  ANDN U4583 ( .B(x[64]), .A(n1559), .Z(n1503) );
  XOR U4584 ( .A(x[66]), .B(x[65]), .Z(n1497) );
  XOR U4585 ( .A(n1574), .B(n1497), .Z(n1548) );
  XOR U4586 ( .A(n1549), .B(n1497), .Z(n1554) );
  NAND U4587 ( .A(n1538), .B(n1554), .Z(n1505) );
  XNOR U4588 ( .A(n1548), .B(n1505), .Z(n1499) );
  XNOR U4589 ( .A(x[65]), .B(n1539), .Z(n1498) );
  XNOR U4590 ( .A(n1499), .B(n1498), .Z(n1500) );
  XOR U4591 ( .A(n1501), .B(n1500), .Z(n1502) );
  XOR U4592 ( .A(n1503), .B(n1502), .Z(n1523) );
  NAND U4593 ( .A(n1521), .B(n1523), .Z(n1504) );
  NAND U4594 ( .A(n1531), .B(n1504), .Z(n1515) );
  IV U4595 ( .A(n1521), .Z(n1522) );
  IV U4596 ( .A(n1523), .Z(n1529) );
  XOR U4597 ( .A(n1505), .B(n1559), .Z(n1508) );
  AND U4598 ( .A(n1548), .B(n1539), .Z(n1506) );
  XNOR U4599 ( .A(x[64]), .B(n1506), .Z(n1507) );
  XNOR U4600 ( .A(n1508), .B(n1507), .Z(n1509) );
  XNOR U4601 ( .A(n1510), .B(n1509), .Z(n1511) );
  XNOR U4602 ( .A(n1512), .B(n1511), .Z(n1533) );
  IV U4603 ( .A(n1533), .Z(n1528) );
  XOR U4604 ( .A(n1529), .B(n1528), .Z(n1513) );
  NAND U4605 ( .A(n1522), .B(n1513), .Z(n1514) );
  AND U4606 ( .A(n1515), .B(n1514), .Z(n1593) );
  NAND U4607 ( .A(n1529), .B(n1522), .Z(n1516) );
  NAND U4608 ( .A(n1528), .B(n1516), .Z(n1519) );
  XOR U4609 ( .A(n1522), .B(n1525), .Z(n1517) );
  NAND U4610 ( .A(n1523), .B(n1517), .Z(n1518) );
  AND U4611 ( .A(n1519), .B(n1518), .Z(n1575) );
  XNOR U4612 ( .A(n1593), .B(n1575), .Z(n1550) );
  OR U4613 ( .A(n1550), .B(n1520), .Z(n1543) );
  NAND U4614 ( .A(n1531), .B(n1521), .Z(n1527) );
  AND U4615 ( .A(n1523), .B(n1522), .Z(n1530) );
  XNOR U4616 ( .A(n1528), .B(n1530), .Z(n1524) );
  NAND U4617 ( .A(n1525), .B(n1524), .Z(n1526) );
  AND U4618 ( .A(n1527), .B(n1526), .Z(n1547) );
  NAND U4619 ( .A(n1529), .B(n1528), .Z(n1535) );
  XNOR U4620 ( .A(n1531), .B(n1530), .Z(n1532) );
  NAND U4621 ( .A(n1533), .B(n1532), .Z(n1534) );
  NAND U4622 ( .A(n1535), .B(n1534), .Z(n1587) );
  XNOR U4623 ( .A(n1547), .B(n1587), .Z(n1565) );
  XOR U4624 ( .A(n1565), .B(n1550), .Z(n1552) );
  OR U4625 ( .A(n1552), .B(n1536), .Z(n1537) );
  XNOR U4626 ( .A(n1543), .B(n1537), .Z(n1569) );
  XOR U4627 ( .A(n1547), .B(n1593), .Z(n1555) );
  NANDN U4628 ( .A(n1555), .B(n1538), .Z(n1595) );
  NANDN U4629 ( .A(n1547), .B(n1539), .Z(n1540) );
  XNOR U4630 ( .A(n1595), .B(n1540), .Z(n1573) );
  XOR U4631 ( .A(n1569), .B(n1573), .Z(n1558) );
  NANDN U4632 ( .A(n1541), .B(n1565), .Z(n1542) );
  XNOR U4633 ( .A(n1543), .B(n1542), .Z(n1603) );
  XNOR U4634 ( .A(n1587), .B(n1575), .Z(n1577) );
  NANDN U4635 ( .A(n1577), .B(n1544), .Z(n1561) );
  NAND U4636 ( .A(n1545), .B(n1575), .Z(n1546) );
  XNOR U4637 ( .A(n1561), .B(n1546), .Z(n1592) );
  XOR U4638 ( .A(n1603), .B(n1592), .Z(n1584) );
  XNOR U4639 ( .A(n1558), .B(n1584), .Z(z[64]) );
  ANDN U4640 ( .B(n1548), .A(n1547), .Z(n1557) );
  NANDN U4641 ( .A(n1550), .B(n1549), .Z(n1568) );
  NANDN U4642 ( .A(n1552), .B(n1551), .Z(n1553) );
  XNOR U4643 ( .A(n1568), .B(n1553), .Z(n1596) );
  NANDN U4644 ( .A(n1555), .B(n1554), .Z(n1562) );
  XNOR U4645 ( .A(n1596), .B(n1562), .Z(n1556) );
  XOR U4646 ( .A(n1557), .B(n1556), .Z(n1582) );
  XOR U4647 ( .A(n1582), .B(n1558), .Z(n1602) );
  ANDN U4648 ( .B(n1593), .A(n1559), .Z(n1564) );
  NAND U4649 ( .A(n1585), .B(n1587), .Z(n1560) );
  XNOR U4650 ( .A(n1561), .B(n1560), .Z(n1572) );
  XNOR U4651 ( .A(n1562), .B(n1572), .Z(n1563) );
  XNOR U4652 ( .A(n1564), .B(n1563), .Z(n1571) );
  NAND U4653 ( .A(n1566), .B(n1565), .Z(n1567) );
  XNOR U4654 ( .A(n1568), .B(n1567), .Z(n1578) );
  XNOR U4655 ( .A(n1569), .B(n1578), .Z(n1570) );
  XOR U4656 ( .A(n1571), .B(n1570), .Z(n1581) );
  XNOR U4657 ( .A(n1602), .B(n1581), .Z(z[65]) );
  XNOR U4658 ( .A(n1573), .B(n1572), .Z(z[66]) );
  AND U4659 ( .A(n1575), .B(n1574), .Z(n1580) );
  NANDN U4660 ( .A(n1577), .B(n1576), .Z(n1590) );
  XNOR U4661 ( .A(n1578), .B(n1590), .Z(n1579) );
  XOR U4662 ( .A(n1580), .B(n1579), .Z(n1601) );
  XOR U4663 ( .A(n1582), .B(n1581), .Z(n1583) );
  XOR U4664 ( .A(n1601), .B(n1583), .Z(z[67]) );
  XOR U4665 ( .A(n1584), .B(z[66]), .Z(z[68]) );
  XNOR U4666 ( .A(n1586), .B(n1585), .Z(n1588) );
  NAND U4667 ( .A(n1588), .B(n1587), .Z(n1589) );
  XOR U4668 ( .A(n1590), .B(n1589), .Z(n1591) );
  XNOR U4669 ( .A(n1592), .B(n1591), .Z(n1598) );
  NAND U4670 ( .A(n1593), .B(x[64]), .Z(n1594) );
  XNOR U4671 ( .A(n1595), .B(n1594), .Z(n1604) );
  XNOR U4672 ( .A(n1596), .B(n1604), .Z(n1597) );
  XOR U4673 ( .A(n1598), .B(n1597), .Z(z[69]) );
  XNOR U4674 ( .A(n1600), .B(n1599), .Z(z[6]) );
  XNOR U4675 ( .A(n1602), .B(n1601), .Z(z[70]) );
  XNOR U4676 ( .A(n1604), .B(n1603), .Z(n1605) );
  XNOR U4677 ( .A(z[65]), .B(n1605), .Z(z[71]) );
  IV U4678 ( .A(x[73]), .Z(n1712) );
  XOR U4679 ( .A(x[72]), .B(x[78]), .Z(n1607) );
  XOR U4680 ( .A(x[77]), .B(n1607), .Z(n1711) );
  IV U4681 ( .A(n1711), .Z(n1608) );
  AND U4682 ( .A(n1712), .B(n1608), .Z(n1615) );
  XNOR U4683 ( .A(x[75]), .B(n1712), .Z(n1611) );
  XNOR U4684 ( .A(x[74]), .B(n1611), .Z(n1606) );
  XNOR U4685 ( .A(n1607), .B(n1606), .Z(n1671) );
  IV U4686 ( .A(n1671), .Z(n1617) );
  XNOR U4687 ( .A(n1617), .B(n1711), .Z(n1670) );
  IV U4688 ( .A(x[79]), .Z(n1609) );
  XNOR U4689 ( .A(x[73]), .B(n1609), .Z(n1702) );
  NAND U4690 ( .A(n1670), .B(n1702), .Z(n1620) );
  XNOR U4691 ( .A(n1609), .B(n1608), .Z(n1616) );
  IV U4692 ( .A(n1616), .Z(n1700) );
  XOR U4693 ( .A(n1671), .B(n1700), .Z(n1636) );
  XNOR U4694 ( .A(n1620), .B(n1636), .Z(n1613) );
  XOR U4695 ( .A(x[72]), .B(n1617), .Z(n1646) );
  XOR U4696 ( .A(x[76]), .B(n1609), .Z(n1610) );
  IV U4697 ( .A(n1610), .Z(n1675) );
  NANDN U4698 ( .A(n1646), .B(n1675), .Z(n1619) );
  XNOR U4699 ( .A(n1611), .B(n1610), .Z(n1664) );
  XNOR U4700 ( .A(n1670), .B(n1664), .Z(n1662) );
  XOR U4701 ( .A(x[74]), .B(x[76]), .Z(n1677) );
  NANDN U4702 ( .A(n1662), .B(n1677), .Z(n1612) );
  XOR U4703 ( .A(n1619), .B(n1612), .Z(n1638) );
  XNOR U4704 ( .A(n1613), .B(n1638), .Z(n1614) );
  XOR U4705 ( .A(n1615), .B(n1614), .Z(n1651) );
  IV U4706 ( .A(n1651), .Z(n1657) );
  AND U4707 ( .A(n1617), .B(n1616), .Z(n1622) );
  XOR U4708 ( .A(x[72]), .B(n1664), .Z(n1665) );
  XNOR U4709 ( .A(n1711), .B(n1665), .Z(n1667) );
  XOR U4710 ( .A(x[74]), .B(x[79]), .Z(n1692) );
  NANDN U4711 ( .A(n1667), .B(n1692), .Z(n1618) );
  XNOR U4712 ( .A(n1619), .B(n1618), .Z(n1627) );
  XNOR U4713 ( .A(n1620), .B(n1627), .Z(n1621) );
  XOR U4714 ( .A(n1622), .B(n1621), .Z(n1647) );
  XNOR U4715 ( .A(x[76]), .B(n1711), .Z(n1685) );
  ANDN U4716 ( .B(x[72]), .A(n1685), .Z(n1629) );
  XOR U4717 ( .A(x[74]), .B(x[73]), .Z(n1623) );
  XOR U4718 ( .A(n1700), .B(n1623), .Z(n1674) );
  XOR U4719 ( .A(n1675), .B(n1623), .Z(n1680) );
  NAND U4720 ( .A(n1664), .B(n1680), .Z(n1631) );
  XNOR U4721 ( .A(n1674), .B(n1631), .Z(n1625) );
  XNOR U4722 ( .A(x[73]), .B(n1665), .Z(n1624) );
  XNOR U4723 ( .A(n1625), .B(n1624), .Z(n1626) );
  XOR U4724 ( .A(n1627), .B(n1626), .Z(n1628) );
  XOR U4725 ( .A(n1629), .B(n1628), .Z(n1649) );
  NAND U4726 ( .A(n1647), .B(n1649), .Z(n1630) );
  NAND U4727 ( .A(n1657), .B(n1630), .Z(n1641) );
  IV U4728 ( .A(n1647), .Z(n1648) );
  IV U4729 ( .A(n1649), .Z(n1655) );
  XOR U4730 ( .A(n1631), .B(n1685), .Z(n1634) );
  AND U4731 ( .A(n1674), .B(n1665), .Z(n1632) );
  XNOR U4732 ( .A(x[72]), .B(n1632), .Z(n1633) );
  XNOR U4733 ( .A(n1634), .B(n1633), .Z(n1635) );
  XNOR U4734 ( .A(n1636), .B(n1635), .Z(n1637) );
  XNOR U4735 ( .A(n1638), .B(n1637), .Z(n1659) );
  IV U4736 ( .A(n1659), .Z(n1654) );
  XOR U4737 ( .A(n1655), .B(n1654), .Z(n1639) );
  NAND U4738 ( .A(n1648), .B(n1639), .Z(n1640) );
  AND U4739 ( .A(n1641), .B(n1640), .Z(n1719) );
  NAND U4740 ( .A(n1655), .B(n1648), .Z(n1642) );
  NAND U4741 ( .A(n1654), .B(n1642), .Z(n1645) );
  XOR U4742 ( .A(n1648), .B(n1651), .Z(n1643) );
  NAND U4743 ( .A(n1649), .B(n1643), .Z(n1644) );
  AND U4744 ( .A(n1645), .B(n1644), .Z(n1701) );
  XNOR U4745 ( .A(n1719), .B(n1701), .Z(n1676) );
  OR U4746 ( .A(n1676), .B(n1646), .Z(n1669) );
  NAND U4747 ( .A(n1657), .B(n1647), .Z(n1653) );
  AND U4748 ( .A(n1649), .B(n1648), .Z(n1656) );
  XNOR U4749 ( .A(n1654), .B(n1656), .Z(n1650) );
  NAND U4750 ( .A(n1651), .B(n1650), .Z(n1652) );
  AND U4751 ( .A(n1653), .B(n1652), .Z(n1673) );
  NAND U4752 ( .A(n1655), .B(n1654), .Z(n1661) );
  XNOR U4753 ( .A(n1657), .B(n1656), .Z(n1658) );
  NAND U4754 ( .A(n1659), .B(n1658), .Z(n1660) );
  NAND U4755 ( .A(n1661), .B(n1660), .Z(n1713) );
  XNOR U4756 ( .A(n1673), .B(n1713), .Z(n1691) );
  XOR U4757 ( .A(n1691), .B(n1676), .Z(n1678) );
  OR U4758 ( .A(n1678), .B(n1662), .Z(n1663) );
  XNOR U4759 ( .A(n1669), .B(n1663), .Z(n1695) );
  XOR U4760 ( .A(n1673), .B(n1719), .Z(n1681) );
  NANDN U4761 ( .A(n1681), .B(n1664), .Z(n1721) );
  NANDN U4762 ( .A(n1673), .B(n1665), .Z(n1666) );
  XNOR U4763 ( .A(n1721), .B(n1666), .Z(n1699) );
  XOR U4764 ( .A(n1695), .B(n1699), .Z(n1684) );
  NANDN U4765 ( .A(n1667), .B(n1691), .Z(n1668) );
  XNOR U4766 ( .A(n1669), .B(n1668), .Z(n1727) );
  XNOR U4767 ( .A(n1713), .B(n1701), .Z(n1703) );
  NANDN U4768 ( .A(n1703), .B(n1670), .Z(n1687) );
  NAND U4769 ( .A(n1671), .B(n1701), .Z(n1672) );
  XNOR U4770 ( .A(n1687), .B(n1672), .Z(n1718) );
  XOR U4771 ( .A(n1727), .B(n1718), .Z(n1710) );
  XNOR U4772 ( .A(n1684), .B(n1710), .Z(z[72]) );
  ANDN U4773 ( .B(n1674), .A(n1673), .Z(n1683) );
  NANDN U4774 ( .A(n1676), .B(n1675), .Z(n1694) );
  NANDN U4775 ( .A(n1678), .B(n1677), .Z(n1679) );
  XNOR U4776 ( .A(n1694), .B(n1679), .Z(n1722) );
  NANDN U4777 ( .A(n1681), .B(n1680), .Z(n1688) );
  XNOR U4778 ( .A(n1722), .B(n1688), .Z(n1682) );
  XOR U4779 ( .A(n1683), .B(n1682), .Z(n1708) );
  XOR U4780 ( .A(n1708), .B(n1684), .Z(n1726) );
  ANDN U4781 ( .B(n1719), .A(n1685), .Z(n1690) );
  NAND U4782 ( .A(n1711), .B(n1713), .Z(n1686) );
  XNOR U4783 ( .A(n1687), .B(n1686), .Z(n1698) );
  XNOR U4784 ( .A(n1688), .B(n1698), .Z(n1689) );
  XNOR U4785 ( .A(n1690), .B(n1689), .Z(n1697) );
  NAND U4786 ( .A(n1692), .B(n1691), .Z(n1693) );
  XNOR U4787 ( .A(n1694), .B(n1693), .Z(n1704) );
  XNOR U4788 ( .A(n1695), .B(n1704), .Z(n1696) );
  XOR U4789 ( .A(n1697), .B(n1696), .Z(n1707) );
  XNOR U4790 ( .A(n1726), .B(n1707), .Z(z[73]) );
  XNOR U4791 ( .A(n1699), .B(n1698), .Z(z[74]) );
  AND U4792 ( .A(n1701), .B(n1700), .Z(n1706) );
  NANDN U4793 ( .A(n1703), .B(n1702), .Z(n1716) );
  XNOR U4794 ( .A(n1704), .B(n1716), .Z(n1705) );
  XOR U4795 ( .A(n1706), .B(n1705), .Z(n1725) );
  XOR U4796 ( .A(n1708), .B(n1707), .Z(n1709) );
  XOR U4797 ( .A(n1725), .B(n1709), .Z(z[75]) );
  XOR U4798 ( .A(n1710), .B(z[74]), .Z(z[76]) );
  XNOR U4799 ( .A(n1712), .B(n1711), .Z(n1714) );
  NAND U4800 ( .A(n1714), .B(n1713), .Z(n1715) );
  XOR U4801 ( .A(n1716), .B(n1715), .Z(n1717) );
  XNOR U4802 ( .A(n1718), .B(n1717), .Z(n1724) );
  NAND U4803 ( .A(n1719), .B(x[72]), .Z(n1720) );
  XNOR U4804 ( .A(n1721), .B(n1720), .Z(n1728) );
  XNOR U4805 ( .A(n1722), .B(n1728), .Z(n1723) );
  XOR U4806 ( .A(n1724), .B(n1723), .Z(z[77]) );
  XNOR U4807 ( .A(n1726), .B(n1725), .Z(z[78]) );
  XNOR U4808 ( .A(n1728), .B(n1727), .Z(n1729) );
  XNOR U4809 ( .A(z[73]), .B(n1729), .Z(z[79]) );
  XNOR U4810 ( .A(n1731), .B(n1730), .Z(n1732) );
  XNOR U4811 ( .A(z[1]), .B(n1732), .Z(z[7]) );
  XOR U4812 ( .A(x[80]), .B(x[86]), .Z(n1733) );
  IV U4813 ( .A(n1838), .Z(n1735) );
  IV U4814 ( .A(x[81]), .Z(n1837) );
  NAND U4815 ( .A(n1735), .B(n1837), .Z(n1742) );
  XNOR U4816 ( .A(x[82]), .B(n1733), .Z(n1734) );
  XNOR U4817 ( .A(n1738), .B(n1734), .Z(n1797) );
  XNOR U4818 ( .A(n1735), .B(n1797), .Z(n1796) );
  IV U4819 ( .A(x[87]), .Z(n1736) );
  XNOR U4820 ( .A(x[81]), .B(n1736), .Z(n1828) );
  NAND U4821 ( .A(n1796), .B(n1828), .Z(n1745) );
  XNOR U4822 ( .A(n1735), .B(n1736), .Z(n1826) );
  XOR U4823 ( .A(n1797), .B(n1826), .Z(n1753) );
  XOR U4824 ( .A(n1745), .B(n1753), .Z(n1740) );
  XNOR U4825 ( .A(x[80]), .B(n1797), .Z(n1772) );
  XOR U4826 ( .A(x[84]), .B(n1736), .Z(n1737) );
  IV U4827 ( .A(n1737), .Z(n1801) );
  NANDN U4828 ( .A(n1772), .B(n1801), .Z(n1744) );
  XOR U4829 ( .A(n1738), .B(n1737), .Z(n1790) );
  XOR U4830 ( .A(n1796), .B(n1790), .Z(n1788) );
  XOR U4831 ( .A(x[82]), .B(x[84]), .Z(n1803) );
  NANDN U4832 ( .A(n1788), .B(n1803), .Z(n1739) );
  XNOR U4833 ( .A(n1744), .B(n1739), .Z(n1749) );
  XOR U4834 ( .A(n1740), .B(n1749), .Z(n1741) );
  XOR U4835 ( .A(n1742), .B(n1741), .Z(n1783) );
  IV U4836 ( .A(n1783), .Z(n1777) );
  ANDN U4837 ( .B(n1826), .A(n1797), .Z(n1747) );
  XNOR U4838 ( .A(x[80]), .B(n1790), .Z(n1791) );
  XNOR U4839 ( .A(n1838), .B(n1791), .Z(n1793) );
  XOR U4840 ( .A(x[82]), .B(x[87]), .Z(n1818) );
  NANDN U4841 ( .A(n1793), .B(n1818), .Z(n1743) );
  XNOR U4842 ( .A(n1744), .B(n1743), .Z(n1760) );
  XNOR U4843 ( .A(n1745), .B(n1760), .Z(n1746) );
  XOR U4844 ( .A(n1747), .B(n1746), .Z(n1773) );
  NAND U4845 ( .A(n1777), .B(n1773), .Z(n1767) );
  IV U4846 ( .A(n1773), .Z(n1774) );
  XOR U4847 ( .A(n1783), .B(n1774), .Z(n1765) );
  XOR U4848 ( .A(x[82]), .B(x[81]), .Z(n1748) );
  XNOR U4849 ( .A(n1826), .B(n1748), .Z(n1800) );
  NAND U4850 ( .A(n1800), .B(n1791), .Z(n1755) );
  XNOR U4851 ( .A(x[84]), .B(n1838), .Z(n1811) );
  XOR U4852 ( .A(n1801), .B(n1748), .Z(n1806) );
  NANDN U4853 ( .A(n1790), .B(n1806), .Z(n1756) );
  XOR U4854 ( .A(n1811), .B(n1756), .Z(n1751) );
  XOR U4855 ( .A(x[80]), .B(n1749), .Z(n1750) );
  XNOR U4856 ( .A(n1751), .B(n1750), .Z(n1752) );
  XOR U4857 ( .A(n1753), .B(n1752), .Z(n1754) );
  XOR U4858 ( .A(n1755), .B(n1754), .Z(n1785) );
  IV U4859 ( .A(n1785), .Z(n1780) );
  AND U4860 ( .A(n1777), .B(n1780), .Z(n1763) );
  ANDN U4861 ( .B(x[80]), .A(n1811), .Z(n1762) );
  XNOR U4862 ( .A(n1800), .B(n1756), .Z(n1758) );
  XNOR U4863 ( .A(x[81]), .B(n1791), .Z(n1757) );
  XNOR U4864 ( .A(n1758), .B(n1757), .Z(n1759) );
  XOR U4865 ( .A(n1760), .B(n1759), .Z(n1761) );
  XOR U4866 ( .A(n1762), .B(n1761), .Z(n1775) );
  IV U4867 ( .A(n1775), .Z(n1781) );
  XNOR U4868 ( .A(n1763), .B(n1781), .Z(n1764) );
  NAND U4869 ( .A(n1765), .B(n1764), .Z(n1766) );
  NAND U4870 ( .A(n1767), .B(n1766), .Z(n1845) );
  NAND U4871 ( .A(n1781), .B(n1774), .Z(n1768) );
  NAND U4872 ( .A(n1780), .B(n1768), .Z(n1771) );
  XOR U4873 ( .A(n1774), .B(n1777), .Z(n1769) );
  NAND U4874 ( .A(n1775), .B(n1769), .Z(n1770) );
  AND U4875 ( .A(n1771), .B(n1770), .Z(n1827) );
  XNOR U4876 ( .A(n1845), .B(n1827), .Z(n1802) );
  OR U4877 ( .A(n1802), .B(n1772), .Z(n1795) );
  NAND U4878 ( .A(n1783), .B(n1773), .Z(n1779) );
  AND U4879 ( .A(n1775), .B(n1774), .Z(n1782) );
  XNOR U4880 ( .A(n1782), .B(n1780), .Z(n1776) );
  NAND U4881 ( .A(n1777), .B(n1776), .Z(n1778) );
  AND U4882 ( .A(n1779), .B(n1778), .Z(n1799) );
  NAND U4883 ( .A(n1781), .B(n1780), .Z(n1787) );
  XNOR U4884 ( .A(n1783), .B(n1782), .Z(n1784) );
  NAND U4885 ( .A(n1785), .B(n1784), .Z(n1786) );
  NAND U4886 ( .A(n1787), .B(n1786), .Z(n1839) );
  XNOR U4887 ( .A(n1799), .B(n1839), .Z(n1817) );
  XOR U4888 ( .A(n1817), .B(n1802), .Z(n1804) );
  OR U4889 ( .A(n1804), .B(n1788), .Z(n1789) );
  XNOR U4890 ( .A(n1795), .B(n1789), .Z(n1821) );
  XOR U4891 ( .A(n1799), .B(n1845), .Z(n1807) );
  OR U4892 ( .A(n1790), .B(n1807), .Z(n1847) );
  NANDN U4893 ( .A(n1799), .B(n1791), .Z(n1792) );
  XNOR U4894 ( .A(n1847), .B(n1792), .Z(n1825) );
  XOR U4895 ( .A(n1821), .B(n1825), .Z(n1810) );
  NANDN U4896 ( .A(n1793), .B(n1817), .Z(n1794) );
  XNOR U4897 ( .A(n1795), .B(n1794), .Z(n1853) );
  XNOR U4898 ( .A(n1839), .B(n1827), .Z(n1829) );
  NANDN U4899 ( .A(n1829), .B(n1796), .Z(n1813) );
  NAND U4900 ( .A(n1797), .B(n1827), .Z(n1798) );
  XNOR U4901 ( .A(n1813), .B(n1798), .Z(n1844) );
  XOR U4902 ( .A(n1853), .B(n1844), .Z(n1836) );
  XNOR U4903 ( .A(n1810), .B(n1836), .Z(z[80]) );
  ANDN U4904 ( .B(n1800), .A(n1799), .Z(n1809) );
  NANDN U4905 ( .A(n1802), .B(n1801), .Z(n1820) );
  NANDN U4906 ( .A(n1804), .B(n1803), .Z(n1805) );
  XNOR U4907 ( .A(n1820), .B(n1805), .Z(n1848) );
  NANDN U4908 ( .A(n1807), .B(n1806), .Z(n1814) );
  XNOR U4909 ( .A(n1848), .B(n1814), .Z(n1808) );
  XOR U4910 ( .A(n1809), .B(n1808), .Z(n1834) );
  XOR U4911 ( .A(n1834), .B(n1810), .Z(n1852) );
  ANDN U4912 ( .B(n1845), .A(n1811), .Z(n1816) );
  NAND U4913 ( .A(n1838), .B(n1839), .Z(n1812) );
  XNOR U4914 ( .A(n1813), .B(n1812), .Z(n1824) );
  XNOR U4915 ( .A(n1814), .B(n1824), .Z(n1815) );
  XNOR U4916 ( .A(n1816), .B(n1815), .Z(n1823) );
  NAND U4917 ( .A(n1818), .B(n1817), .Z(n1819) );
  XNOR U4918 ( .A(n1820), .B(n1819), .Z(n1830) );
  XNOR U4919 ( .A(n1821), .B(n1830), .Z(n1822) );
  XOR U4920 ( .A(n1823), .B(n1822), .Z(n1833) );
  XNOR U4921 ( .A(n1852), .B(n1833), .Z(z[81]) );
  XNOR U4922 ( .A(n1825), .B(n1824), .Z(z[82]) );
  ANDN U4923 ( .B(n1827), .A(n1826), .Z(n1832) );
  NANDN U4924 ( .A(n1829), .B(n1828), .Z(n1842) );
  XNOR U4925 ( .A(n1830), .B(n1842), .Z(n1831) );
  XOR U4926 ( .A(n1832), .B(n1831), .Z(n1851) );
  XOR U4927 ( .A(n1834), .B(n1833), .Z(n1835) );
  XOR U4928 ( .A(n1851), .B(n1835), .Z(z[83]) );
  XOR U4929 ( .A(n1836), .B(z[82]), .Z(z[84]) );
  XNOR U4930 ( .A(n1838), .B(n1837), .Z(n1840) );
  NAND U4931 ( .A(n1840), .B(n1839), .Z(n1841) );
  XOR U4932 ( .A(n1842), .B(n1841), .Z(n1843) );
  XNOR U4933 ( .A(n1844), .B(n1843), .Z(n1850) );
  NAND U4934 ( .A(x[80]), .B(n1845), .Z(n1846) );
  XNOR U4935 ( .A(n1847), .B(n1846), .Z(n1854) );
  XNOR U4936 ( .A(n1848), .B(n1854), .Z(n1849) );
  XOR U4937 ( .A(n1850), .B(n1849), .Z(z[85]) );
  XNOR U4938 ( .A(n1852), .B(n1851), .Z(z[86]) );
  XNOR U4939 ( .A(n1854), .B(n1853), .Z(n1855) );
  XNOR U4940 ( .A(z[81]), .B(n1855), .Z(z[87]) );
  XOR U4941 ( .A(x[88]), .B(x[94]), .Z(n1856) );
  XOR U4942 ( .A(x[93]), .B(n1856), .Z(n1963) );
  IV U4943 ( .A(n1963), .Z(n1858) );
  IV U4944 ( .A(x[89]), .Z(n1962) );
  NAND U4945 ( .A(n1858), .B(n1962), .Z(n1865) );
  XOR U4946 ( .A(x[91]), .B(x[89]), .Z(n1861) );
  XNOR U4947 ( .A(x[90]), .B(n1856), .Z(n1857) );
  XNOR U4948 ( .A(n1861), .B(n1857), .Z(n1920) );
  XNOR U4949 ( .A(n1858), .B(n1920), .Z(n1919) );
  IV U4950 ( .A(x[95]), .Z(n1859) );
  XNOR U4951 ( .A(x[89]), .B(n1859), .Z(n1953) );
  NAND U4952 ( .A(n1919), .B(n1953), .Z(n1868) );
  XNOR U4953 ( .A(n1858), .B(n1859), .Z(n1951) );
  XOR U4954 ( .A(n1920), .B(n1951), .Z(n1876) );
  XOR U4955 ( .A(n1868), .B(n1876), .Z(n1863) );
  XNOR U4956 ( .A(x[88]), .B(n1920), .Z(n1895) );
  XOR U4957 ( .A(x[92]), .B(n1859), .Z(n1860) );
  IV U4958 ( .A(n1860), .Z(n1924) );
  NANDN U4959 ( .A(n1895), .B(n1924), .Z(n1867) );
  XOR U4960 ( .A(n1861), .B(n1860), .Z(n1913) );
  XOR U4961 ( .A(n1919), .B(n1913), .Z(n1911) );
  XOR U4962 ( .A(x[90]), .B(x[92]), .Z(n1926) );
  NANDN U4963 ( .A(n1911), .B(n1926), .Z(n1862) );
  XNOR U4964 ( .A(n1867), .B(n1862), .Z(n1872) );
  XOR U4965 ( .A(n1863), .B(n1872), .Z(n1864) );
  XOR U4966 ( .A(n1865), .B(n1864), .Z(n1906) );
  IV U4967 ( .A(n1906), .Z(n1900) );
  ANDN U4968 ( .B(n1951), .A(n1920), .Z(n1870) );
  XNOR U4969 ( .A(x[88]), .B(n1913), .Z(n1914) );
  XNOR U4970 ( .A(n1963), .B(n1914), .Z(n1916) );
  XOR U4971 ( .A(x[90]), .B(x[95]), .Z(n1941) );
  NANDN U4972 ( .A(n1916), .B(n1941), .Z(n1866) );
  XNOR U4973 ( .A(n1867), .B(n1866), .Z(n1883) );
  XNOR U4974 ( .A(n1868), .B(n1883), .Z(n1869) );
  XOR U4975 ( .A(n1870), .B(n1869), .Z(n1896) );
  NAND U4976 ( .A(n1900), .B(n1896), .Z(n1890) );
  IV U4977 ( .A(n1896), .Z(n1897) );
  XOR U4978 ( .A(n1906), .B(n1897), .Z(n1888) );
  XOR U4979 ( .A(x[90]), .B(x[89]), .Z(n1871) );
  XNOR U4980 ( .A(n1951), .B(n1871), .Z(n1923) );
  NAND U4981 ( .A(n1923), .B(n1914), .Z(n1878) );
  XNOR U4982 ( .A(x[92]), .B(n1963), .Z(n1934) );
  XOR U4983 ( .A(n1924), .B(n1871), .Z(n1929) );
  NANDN U4984 ( .A(n1913), .B(n1929), .Z(n1879) );
  XOR U4985 ( .A(n1934), .B(n1879), .Z(n1874) );
  XOR U4986 ( .A(x[88]), .B(n1872), .Z(n1873) );
  XNOR U4987 ( .A(n1874), .B(n1873), .Z(n1875) );
  XOR U4988 ( .A(n1876), .B(n1875), .Z(n1877) );
  XOR U4989 ( .A(n1878), .B(n1877), .Z(n1908) );
  IV U4990 ( .A(n1908), .Z(n1903) );
  AND U4991 ( .A(n1900), .B(n1903), .Z(n1886) );
  ANDN U4992 ( .B(x[88]), .A(n1934), .Z(n1885) );
  XNOR U4993 ( .A(n1923), .B(n1879), .Z(n1881) );
  XNOR U4994 ( .A(x[89]), .B(n1914), .Z(n1880) );
  XNOR U4995 ( .A(n1881), .B(n1880), .Z(n1882) );
  XOR U4996 ( .A(n1883), .B(n1882), .Z(n1884) );
  XOR U4997 ( .A(n1885), .B(n1884), .Z(n1898) );
  IV U4998 ( .A(n1898), .Z(n1904) );
  XNOR U4999 ( .A(n1886), .B(n1904), .Z(n1887) );
  NAND U5000 ( .A(n1888), .B(n1887), .Z(n1889) );
  NAND U5001 ( .A(n1890), .B(n1889), .Z(n1970) );
  NAND U5002 ( .A(n1904), .B(n1897), .Z(n1891) );
  NAND U5003 ( .A(n1903), .B(n1891), .Z(n1894) );
  XOR U5004 ( .A(n1897), .B(n1900), .Z(n1892) );
  NAND U5005 ( .A(n1898), .B(n1892), .Z(n1893) );
  AND U5006 ( .A(n1894), .B(n1893), .Z(n1952) );
  XNOR U5007 ( .A(n1970), .B(n1952), .Z(n1925) );
  OR U5008 ( .A(n1925), .B(n1895), .Z(n1918) );
  NAND U5009 ( .A(n1906), .B(n1896), .Z(n1902) );
  AND U5010 ( .A(n1898), .B(n1897), .Z(n1905) );
  XNOR U5011 ( .A(n1905), .B(n1903), .Z(n1899) );
  NAND U5012 ( .A(n1900), .B(n1899), .Z(n1901) );
  AND U5013 ( .A(n1902), .B(n1901), .Z(n1922) );
  NAND U5014 ( .A(n1904), .B(n1903), .Z(n1910) );
  XNOR U5015 ( .A(n1906), .B(n1905), .Z(n1907) );
  NAND U5016 ( .A(n1908), .B(n1907), .Z(n1909) );
  NAND U5017 ( .A(n1910), .B(n1909), .Z(n1964) );
  XNOR U5018 ( .A(n1922), .B(n1964), .Z(n1940) );
  XOR U5019 ( .A(n1940), .B(n1925), .Z(n1927) );
  OR U5020 ( .A(n1927), .B(n1911), .Z(n1912) );
  XNOR U5021 ( .A(n1918), .B(n1912), .Z(n1944) );
  XOR U5022 ( .A(n1922), .B(n1970), .Z(n1930) );
  OR U5023 ( .A(n1913), .B(n1930), .Z(n1972) );
  NANDN U5024 ( .A(n1922), .B(n1914), .Z(n1915) );
  XNOR U5025 ( .A(n1972), .B(n1915), .Z(n1950) );
  XOR U5026 ( .A(n1944), .B(n1950), .Z(n1933) );
  NANDN U5027 ( .A(n1916), .B(n1940), .Z(n1917) );
  XNOR U5028 ( .A(n1918), .B(n1917), .Z(n1978) );
  XNOR U5029 ( .A(n1964), .B(n1952), .Z(n1954) );
  NANDN U5030 ( .A(n1954), .B(n1919), .Z(n1936) );
  NAND U5031 ( .A(n1920), .B(n1952), .Z(n1921) );
  XNOR U5032 ( .A(n1936), .B(n1921), .Z(n1969) );
  XOR U5033 ( .A(n1978), .B(n1969), .Z(n1961) );
  XNOR U5034 ( .A(n1933), .B(n1961), .Z(z[88]) );
  ANDN U5035 ( .B(n1923), .A(n1922), .Z(n1932) );
  NANDN U5036 ( .A(n1925), .B(n1924), .Z(n1943) );
  NANDN U5037 ( .A(n1927), .B(n1926), .Z(n1928) );
  XNOR U5038 ( .A(n1943), .B(n1928), .Z(n1973) );
  NANDN U5039 ( .A(n1930), .B(n1929), .Z(n1937) );
  XNOR U5040 ( .A(n1973), .B(n1937), .Z(n1931) );
  XOR U5041 ( .A(n1932), .B(n1931), .Z(n1959) );
  XOR U5042 ( .A(n1959), .B(n1933), .Z(n1977) );
  ANDN U5043 ( .B(n1970), .A(n1934), .Z(n1939) );
  NAND U5044 ( .A(n1963), .B(n1964), .Z(n1935) );
  XNOR U5045 ( .A(n1936), .B(n1935), .Z(n1949) );
  XNOR U5046 ( .A(n1937), .B(n1949), .Z(n1938) );
  XNOR U5047 ( .A(n1939), .B(n1938), .Z(n1946) );
  NAND U5048 ( .A(n1941), .B(n1940), .Z(n1942) );
  XNOR U5049 ( .A(n1943), .B(n1942), .Z(n1955) );
  XNOR U5050 ( .A(n1944), .B(n1955), .Z(n1945) );
  XOR U5051 ( .A(n1946), .B(n1945), .Z(n1958) );
  XNOR U5052 ( .A(n1977), .B(n1958), .Z(z[89]) );
  XNOR U5053 ( .A(n1948), .B(n1947), .Z(z[8]) );
  XNOR U5054 ( .A(n1950), .B(n1949), .Z(z[90]) );
  ANDN U5055 ( .B(n1952), .A(n1951), .Z(n1957) );
  NANDN U5056 ( .A(n1954), .B(n1953), .Z(n1967) );
  XNOR U5057 ( .A(n1955), .B(n1967), .Z(n1956) );
  XOR U5058 ( .A(n1957), .B(n1956), .Z(n1976) );
  XOR U5059 ( .A(n1959), .B(n1958), .Z(n1960) );
  XOR U5060 ( .A(n1976), .B(n1960), .Z(z[91]) );
  XOR U5061 ( .A(n1961), .B(z[90]), .Z(z[92]) );
  XNOR U5062 ( .A(n1963), .B(n1962), .Z(n1965) );
  NAND U5063 ( .A(n1965), .B(n1964), .Z(n1966) );
  XOR U5064 ( .A(n1967), .B(n1966), .Z(n1968) );
  XNOR U5065 ( .A(n1969), .B(n1968), .Z(n1975) );
  NAND U5066 ( .A(x[88]), .B(n1970), .Z(n1971) );
  XNOR U5067 ( .A(n1972), .B(n1971), .Z(n1979) );
  XNOR U5068 ( .A(n1973), .B(n1979), .Z(n1974) );
  XOR U5069 ( .A(n1975), .B(n1974), .Z(z[93]) );
  XNOR U5070 ( .A(n1977), .B(n1976), .Z(z[94]) );
  XNOR U5071 ( .A(n1979), .B(n1978), .Z(n1980) );
  XNOR U5072 ( .A(z[89]), .B(n1980), .Z(z[95]) );
  XNOR U5073 ( .A(n1982), .B(n1981), .Z(z[96]) );
  XOR U5074 ( .A(n1984), .B(n1983), .Z(n1985) );
  XOR U5075 ( .A(n1986), .B(n1985), .Z(z[99]) );
endmodule


module aes_seq_CC2 ( clk, rst, msg, key, out );
  input [127:0] msg;
  input [639:0] key;
  output [127:0] out;
  input clk, rst;
  wire   init, \w0[4][127] , \w0[4][126] , \w0[4][125] , \w0[4][124] ,
         \w0[4][123] , \w0[4][122] , \w0[4][121] , \w0[4][120] , \w0[4][119] ,
         \w0[4][118] , \w0[4][117] , \w0[4][116] , \w0[4][115] , \w0[4][114] ,
         \w0[4][113] , \w0[4][112] , \w0[4][111] , \w0[4][110] , \w0[4][109] ,
         \w0[4][108] , \w0[4][107] , \w0[4][106] , \w0[4][105] , \w0[4][104] ,
         \w0[4][103] , \w0[4][102] , \w0[4][101] , \w0[4][100] , \w0[4][99] ,
         \w0[4][98] , \w0[4][97] , \w0[4][96] , \w0[4][95] , \w0[4][94] ,
         \w0[4][93] , \w0[4][92] , \w0[4][91] , \w0[4][90] , \w0[4][89] ,
         \w0[4][88] , \w0[4][87] , \w0[4][86] , \w0[4][85] , \w0[4][84] ,
         \w0[4][83] , \w0[4][82] , \w0[4][81] , \w0[4][80] , \w0[4][79] ,
         \w0[4][78] , \w0[4][77] , \w0[4][76] , \w0[4][75] , \w0[4][74] ,
         \w0[4][73] , \w0[4][72] , \w0[4][71] , \w0[4][70] , \w0[4][69] ,
         \w0[4][68] , \w0[4][67] , \w0[4][66] , \w0[4][65] , \w0[4][64] ,
         \w0[4][63] , \w0[4][62] , \w0[4][61] , \w0[4][60] , \w0[4][59] ,
         \w0[4][58] , \w0[4][57] , \w0[4][56] , \w0[4][55] , \w0[4][54] ,
         \w0[4][53] , \w0[4][52] , \w0[4][51] , \w0[4][50] , \w0[4][49] ,
         \w0[4][48] , \w0[4][47] , \w0[4][46] , \w0[4][45] , \w0[4][44] ,
         \w0[4][43] , \w0[4][42] , \w0[4][41] , \w0[4][40] , \w0[4][39] ,
         \w0[4][38] , \w0[4][37] , \w0[4][36] , \w0[4][35] , \w0[4][34] ,
         \w0[4][33] , \w0[4][32] , \w0[4][31] , \w0[4][30] , \w0[4][29] ,
         \w0[4][28] , \w0[4][27] , \w0[4][26] , \w0[4][25] , \w0[4][24] ,
         \w0[4][23] , \w0[4][22] , \w0[4][21] , \w0[4][20] , \w0[4][19] ,
         \w0[4][18] , \w0[4][17] , \w0[4][16] , \w0[4][15] , \w0[4][14] ,
         \w0[4][13] , \w0[4][12] , \w0[4][11] , \w0[4][10] , \w0[4][9] ,
         \w0[4][8] , \w0[4][7] , \w0[4][6] , \w0[4][5] , \w0[4][4] ,
         \w0[4][3] , \w0[4][2] , \w0[4][1] , \w0[4][0] , \w1[4][127] ,
         \w1[4][126] , \w1[4][125] , \w1[4][124] , \w1[4][123] , \w1[4][122] ,
         \w1[4][121] , \w1[4][120] , \w1[4][119] , \w1[4][118] , \w1[4][117] ,
         \w1[4][116] , \w1[4][115] , \w1[4][114] , \w1[4][113] , \w1[4][112] ,
         \w1[4][111] , \w1[4][110] , \w1[4][109] , \w1[4][108] , \w1[4][107] ,
         \w1[4][106] , \w1[4][105] , \w1[4][104] , \w1[4][103] , \w1[4][102] ,
         \w1[4][101] , \w1[4][100] , \w1[4][99] , \w1[4][98] , \w1[4][97] ,
         \w1[4][96] , \w1[4][95] , \w1[4][94] , \w1[4][93] , \w1[4][92] ,
         \w1[4][91] , \w1[4][90] , \w1[4][89] , \w1[4][88] , \w1[4][87] ,
         \w1[4][86] , \w1[4][85] , \w1[4][84] , \w1[4][83] , \w1[4][82] ,
         \w1[4][81] , \w1[4][80] , \w1[4][79] , \w1[4][78] , \w1[4][77] ,
         \w1[4][76] , \w1[4][75] , \w1[4][74] , \w1[4][73] , \w1[4][72] ,
         \w1[4][71] , \w1[4][70] , \w1[4][69] , \w1[4][68] , \w1[4][67] ,
         \w1[4][66] , \w1[4][65] , \w1[4][64] , \w1[4][63] , \w1[4][62] ,
         \w1[4][61] , \w1[4][60] , \w1[4][59] , \w1[4][58] , \w1[4][57] ,
         \w1[4][56] , \w1[4][55] , \w1[4][54] , \w1[4][53] , \w1[4][52] ,
         \w1[4][51] , \w1[4][50] , \w1[4][49] , \w1[4][48] , \w1[4][47] ,
         \w1[4][46] , \w1[4][45] , \w1[4][44] , \w1[4][43] , \w1[4][42] ,
         \w1[4][41] , \w1[4][40] , \w1[4][39] , \w1[4][38] , \w1[4][37] ,
         \w1[4][36] , \w1[4][35] , \w1[4][34] , \w1[4][33] , \w1[4][32] ,
         \w1[4][31] , \w1[4][30] , \w1[4][29] , \w1[4][28] , \w1[4][27] ,
         \w1[4][26] , \w1[4][25] , \w1[4][24] , \w1[4][23] , \w1[4][22] ,
         \w1[4][21] , \w1[4][20] , \w1[4][19] , \w1[4][18] , \w1[4][17] ,
         \w1[4][16] , \w1[4][15] , \w1[4][14] , \w1[4][13] , \w1[4][12] ,
         \w1[4][11] , \w1[4][10] , \w1[4][9] , \w1[4][8] , \w1[4][7] ,
         \w1[4][6] , \w1[4][5] , \w1[4][4] , \w1[4][3] , \w1[4][2] ,
         \w1[4][1] , \w1[4][0] , \w1[3][127] , \w1[3][126] , \w1[3][125] ,
         \w1[3][124] , \w1[3][123] , \w1[3][122] , \w1[3][121] , \w1[3][120] ,
         \w1[3][119] , \w1[3][118] , \w1[3][117] , \w1[3][116] , \w1[3][115] ,
         \w1[3][114] , \w1[3][113] , \w1[3][112] , \w1[3][111] , \w1[3][110] ,
         \w1[3][109] , \w1[3][108] , \w1[3][107] , \w1[3][106] , \w1[3][105] ,
         \w1[3][104] , \w1[3][103] , \w1[3][102] , \w1[3][101] , \w1[3][100] ,
         \w1[3][99] , \w1[3][98] , \w1[3][97] , \w1[3][96] , \w1[3][95] ,
         \w1[3][94] , \w1[3][93] , \w1[3][92] , \w1[3][91] , \w1[3][90] ,
         \w1[3][89] , \w1[3][88] , \w1[3][87] , \w1[3][86] , \w1[3][85] ,
         \w1[3][84] , \w1[3][83] , \w1[3][82] , \w1[3][81] , \w1[3][80] ,
         \w1[3][79] , \w1[3][78] , \w1[3][77] , \w1[3][76] , \w1[3][75] ,
         \w1[3][74] , \w1[3][73] , \w1[3][72] , \w1[3][71] , \w1[3][70] ,
         \w1[3][69] , \w1[3][68] , \w1[3][67] , \w1[3][66] , \w1[3][65] ,
         \w1[3][64] , \w1[3][63] , \w1[3][62] , \w1[3][61] , \w1[3][60] ,
         \w1[3][59] , \w1[3][58] , \w1[3][57] , \w1[3][56] , \w1[3][55] ,
         \w1[3][54] , \w1[3][53] , \w1[3][52] , \w1[3][51] , \w1[3][50] ,
         \w1[3][49] , \w1[3][48] , \w1[3][47] , \w1[3][46] , \w1[3][45] ,
         \w1[3][44] , \w1[3][43] , \w1[3][42] , \w1[3][41] , \w1[3][40] ,
         \w1[3][39] , \w1[3][38] , \w1[3][37] , \w1[3][36] , \w1[3][35] ,
         \w1[3][34] , \w1[3][33] , \w1[3][32] , \w1[3][31] , \w1[3][30] ,
         \w1[3][29] , \w1[3][28] , \w1[3][27] , \w1[3][26] , \w1[3][25] ,
         \w1[3][24] , \w1[3][23] , \w1[3][22] , \w1[3][21] , \w1[3][20] ,
         \w1[3][19] , \w1[3][18] , \w1[3][17] , \w1[3][16] , \w1[3][15] ,
         \w1[3][14] , \w1[3][13] , \w1[3][12] , \w1[3][11] , \w1[3][10] ,
         \w1[3][9] , \w1[3][8] , \w1[3][7] , \w1[3][6] , \w1[3][5] ,
         \w1[3][4] , \w1[3][3] , \w1[3][2] , \w1[3][1] , \w1[3][0] ,
         \w1[2][127] , \w1[2][126] , \w1[2][125] , \w1[2][124] , \w1[2][123] ,
         \w1[2][122] , \w1[2][121] , \w1[2][120] , \w1[2][119] , \w1[2][118] ,
         \w1[2][117] , \w1[2][116] , \w1[2][115] , \w1[2][114] , \w1[2][113] ,
         \w1[2][112] , \w1[2][111] , \w1[2][110] , \w1[2][109] , \w1[2][108] ,
         \w1[2][107] , \w1[2][106] , \w1[2][105] , \w1[2][104] , \w1[2][103] ,
         \w1[2][102] , \w1[2][101] , \w1[2][100] , \w1[2][99] , \w1[2][98] ,
         \w1[2][97] , \w1[2][96] , \w1[2][95] , \w1[2][94] , \w1[2][93] ,
         \w1[2][92] , \w1[2][91] , \w1[2][90] , \w1[2][89] , \w1[2][88] ,
         \w1[2][87] , \w1[2][86] , \w1[2][85] , \w1[2][84] , \w1[2][83] ,
         \w1[2][82] , \w1[2][81] , \w1[2][80] , \w1[2][79] , \w1[2][78] ,
         \w1[2][77] , \w1[2][76] , \w1[2][75] , \w1[2][74] , \w1[2][73] ,
         \w1[2][72] , \w1[2][71] , \w1[2][70] , \w1[2][69] , \w1[2][68] ,
         \w1[2][67] , \w1[2][66] , \w1[2][65] , \w1[2][64] , \w1[2][63] ,
         \w1[2][62] , \w1[2][61] , \w1[2][60] , \w1[2][59] , \w1[2][58] ,
         \w1[2][57] , \w1[2][56] , \w1[2][55] , \w1[2][54] , \w1[2][53] ,
         \w1[2][52] , \w1[2][51] , \w1[2][50] , \w1[2][49] , \w1[2][48] ,
         \w1[2][47] , \w1[2][46] , \w1[2][45] , \w1[2][44] , \w1[2][43] ,
         \w1[2][42] , \w1[2][41] , \w1[2][40] , \w1[2][39] , \w1[2][38] ,
         \w1[2][37] , \w1[2][36] , \w1[2][35] , \w1[2][34] , \w1[2][33] ,
         \w1[2][32] , \w1[2][31] , \w1[2][30] , \w1[2][29] , \w1[2][28] ,
         \w1[2][27] , \w1[2][26] , \w1[2][25] , \w1[2][24] , \w1[2][23] ,
         \w1[2][22] , \w1[2][21] , \w1[2][20] , \w1[2][19] , \w1[2][18] ,
         \w1[2][17] , \w1[2][16] , \w1[2][15] , \w1[2][14] , \w1[2][13] ,
         \w1[2][12] , \w1[2][11] , \w1[2][10] , \w1[2][9] , \w1[2][8] ,
         \w1[2][7] , \w1[2][6] , \w1[2][5] , \w1[2][4] , \w1[2][3] ,
         \w1[2][2] , \w1[2][1] , \w1[2][0] , \w1[1][127] , \w1[1][126] ,
         \w1[1][125] , \w1[1][124] , \w1[1][123] , \w1[1][122] , \w1[1][121] ,
         \w1[1][120] , \w1[1][119] , \w1[1][118] , \w1[1][117] , \w1[1][116] ,
         \w1[1][115] , \w1[1][114] , \w1[1][113] , \w1[1][112] , \w1[1][111] ,
         \w1[1][110] , \w1[1][109] , \w1[1][108] , \w1[1][107] , \w1[1][106] ,
         \w1[1][105] , \w1[1][104] , \w1[1][103] , \w1[1][102] , \w1[1][101] ,
         \w1[1][100] , \w1[1][99] , \w1[1][98] , \w1[1][97] , \w1[1][96] ,
         \w1[1][95] , \w1[1][94] , \w1[1][93] , \w1[1][92] , \w1[1][91] ,
         \w1[1][90] , \w1[1][89] , \w1[1][88] , \w1[1][87] , \w1[1][86] ,
         \w1[1][85] , \w1[1][84] , \w1[1][83] , \w1[1][82] , \w1[1][81] ,
         \w1[1][80] , \w1[1][79] , \w1[1][78] , \w1[1][77] , \w1[1][76] ,
         \w1[1][75] , \w1[1][74] , \w1[1][73] , \w1[1][72] , \w1[1][71] ,
         \w1[1][70] , \w1[1][69] , \w1[1][68] , \w1[1][67] , \w1[1][66] ,
         \w1[1][65] , \w1[1][64] , \w1[1][63] , \w1[1][62] , \w1[1][61] ,
         \w1[1][60] , \w1[1][59] , \w1[1][58] , \w1[1][57] , \w1[1][56] ,
         \w1[1][55] , \w1[1][54] , \w1[1][53] , \w1[1][52] , \w1[1][51] ,
         \w1[1][50] , \w1[1][49] , \w1[1][48] , \w1[1][47] , \w1[1][46] ,
         \w1[1][45] , \w1[1][44] , \w1[1][43] , \w1[1][42] , \w1[1][41] ,
         \w1[1][40] , \w1[1][39] , \w1[1][38] , \w1[1][37] , \w1[1][36] ,
         \w1[1][35] , \w1[1][34] , \w1[1][33] , \w1[1][32] , \w1[1][31] ,
         \w1[1][30] , \w1[1][29] , \w1[1][28] , \w1[1][27] , \w1[1][26] ,
         \w1[1][25] , \w1[1][24] , \w1[1][23] , \w1[1][22] , \w1[1][21] ,
         \w1[1][20] , \w1[1][19] , \w1[1][18] , \w1[1][17] , \w1[1][16] ,
         \w1[1][15] , \w1[1][14] , \w1[1][13] , \w1[1][12] , \w1[1][11] ,
         \w1[1][10] , \w1[1][9] , \w1[1][8] , \w1[1][7] , \w1[1][6] ,
         \w1[1][5] , \w1[1][4] , \w1[1][3] , \w1[1][2] , \w1[1][1] ,
         \w1[1][0] , \w1[0][127] , \w1[0][126] , \w1[0][125] , \w1[0][124] ,
         \w1[0][123] , \w1[0][122] , \w1[0][121] , \w1[0][120] , \w1[0][119] ,
         \w1[0][118] , \w1[0][117] , \w1[0][116] , \w1[0][115] , \w1[0][114] ,
         \w1[0][113] , \w1[0][112] , \w1[0][111] , \w1[0][110] , \w1[0][109] ,
         \w1[0][108] , \w1[0][107] , \w1[0][106] , \w1[0][105] , \w1[0][104] ,
         \w1[0][103] , \w1[0][102] , \w1[0][101] , \w1[0][100] , \w1[0][99] ,
         \w1[0][98] , \w1[0][97] , \w1[0][96] , \w1[0][95] , \w1[0][94] ,
         \w1[0][93] , \w1[0][92] , \w1[0][91] , \w1[0][90] , \w1[0][89] ,
         \w1[0][88] , \w1[0][87] , \w1[0][86] , \w1[0][85] , \w1[0][84] ,
         \w1[0][83] , \w1[0][82] , \w1[0][81] , \w1[0][80] , \w1[0][79] ,
         \w1[0][78] , \w1[0][77] , \w1[0][76] , \w1[0][75] , \w1[0][74] ,
         \w1[0][73] , \w1[0][72] , \w1[0][71] , \w1[0][70] , \w1[0][69] ,
         \w1[0][68] , \w1[0][67] , \w1[0][66] , \w1[0][65] , \w1[0][64] ,
         \w1[0][63] , \w1[0][62] , \w1[0][61] , \w1[0][60] , \w1[0][59] ,
         \w1[0][58] , \w1[0][57] , \w1[0][56] , \w1[0][55] , \w1[0][54] ,
         \w1[0][53] , \w1[0][52] , \w1[0][51] , \w1[0][50] , \w1[0][49] ,
         \w1[0][48] , \w1[0][47] , \w1[0][46] , \w1[0][45] , \w1[0][44] ,
         \w1[0][43] , \w1[0][42] , \w1[0][41] , \w1[0][40] , \w1[0][39] ,
         \w1[0][38] , \w1[0][37] , \w1[0][36] , \w1[0][35] , \w1[0][34] ,
         \w1[0][33] , \w1[0][32] , \w1[0][31] , \w1[0][30] , \w1[0][29] ,
         \w1[0][28] , \w1[0][27] , \w1[0][26] , \w1[0][25] , \w1[0][24] ,
         \w1[0][23] , \w1[0][22] , \w1[0][21] , \w1[0][20] , \w1[0][19] ,
         \w1[0][18] , \w1[0][17] , \w1[0][16] , \w1[0][15] , \w1[0][14] ,
         \w1[0][13] , \w1[0][12] , \w1[0][11] , \w1[0][10] , \w1[0][9] ,
         \w1[0][8] , \w1[0][7] , \w1[0][6] , \w1[0][5] , \w1[0][4] ,
         \w1[0][3] , \w1[0][2] , \w1[0][1] , \w1[0][0] , \w3[4][127] ,
         \w3[4][126] , \w3[4][125] , \w3[4][124] , \w3[4][123] , \w3[4][122] ,
         \w3[4][121] , \w3[4][120] , \w3[4][119] , \w3[4][118] , \w3[4][117] ,
         \w3[4][116] , \w3[4][115] , \w3[4][114] , \w3[4][113] , \w3[4][112] ,
         \w3[4][111] , \w3[4][110] , \w3[4][109] , \w3[4][108] , \w3[4][107] ,
         \w3[4][106] , \w3[4][105] , \w3[4][104] , \w3[4][103] , \w3[4][102] ,
         \w3[4][101] , \w3[4][100] , \w3[4][99] , \w3[4][98] , \w3[4][97] ,
         \w3[4][96] , \w3[4][95] , \w3[4][94] , \w3[4][93] , \w3[4][92] ,
         \w3[4][91] , \w3[4][90] , \w3[4][89] , \w3[4][88] , \w3[4][87] ,
         \w3[4][86] , \w3[4][85] , \w3[4][84] , \w3[4][83] , \w3[4][82] ,
         \w3[4][81] , \w3[4][80] , \w3[4][79] , \w3[4][78] , \w3[4][77] ,
         \w3[4][76] , \w3[4][75] , \w3[4][74] , \w3[4][73] , \w3[4][72] ,
         \w3[4][71] , \w3[4][70] , \w3[4][69] , \w3[4][68] , \w3[4][67] ,
         \w3[4][66] , \w3[4][65] , \w3[4][64] , \w3[4][63] , \w3[4][62] ,
         \w3[4][61] , \w3[4][60] , \w3[4][59] , \w3[4][58] , \w3[4][57] ,
         \w3[4][56] , \w3[4][55] , \w3[4][54] , \w3[4][53] , \w3[4][52] ,
         \w3[4][51] , \w3[4][50] , \w3[4][49] , \w3[4][48] , \w3[4][47] ,
         \w3[4][46] , \w3[4][45] , \w3[4][44] , \w3[4][43] , \w3[4][42] ,
         \w3[4][41] , \w3[4][40] , \w3[4][39] , \w3[4][38] , \w3[4][37] ,
         \w3[4][36] , \w3[4][35] , \w3[4][34] , \w3[4][33] , \w3[4][32] ,
         \w3[4][31] , \w3[4][30] , \w3[4][29] , \w3[4][28] , \w3[4][27] ,
         \w3[4][26] , \w3[4][25] , \w3[4][24] , \w3[4][23] , \w3[4][22] ,
         \w3[4][21] , \w3[4][20] , \w3[4][19] , \w3[4][18] , \w3[4][17] ,
         \w3[4][16] , \w3[4][15] , \w3[4][14] , \w3[4][13] , \w3[4][12] ,
         \w3[4][11] , \w3[4][10] , \w3[4][9] , \w3[4][8] , \w3[4][7] ,
         \w3[4][6] , \w3[4][5] , \w3[4][4] , \w3[4][3] , \w3[4][2] ,
         \w3[4][1] , \w3[4][0] , \w3[3][127] , \w3[3][126] , \w3[3][125] ,
         \w3[3][124] , \w3[3][123] , \w3[3][122] , \w3[3][121] , \w3[3][120] ,
         \w3[3][119] , \w3[3][118] , \w3[3][117] , \w3[3][116] , \w3[3][115] ,
         \w3[3][114] , \w3[3][113] , \w3[3][112] , \w3[3][111] , \w3[3][110] ,
         \w3[3][109] , \w3[3][108] , \w3[3][107] , \w3[3][106] , \w3[3][105] ,
         \w3[3][104] , \w3[3][103] , \w3[3][102] , \w3[3][101] , \w3[3][100] ,
         \w3[3][99] , \w3[3][98] , \w3[3][97] , \w3[3][96] , \w3[3][95] ,
         \w3[3][94] , \w3[3][93] , \w3[3][92] , \w3[3][91] , \w3[3][90] ,
         \w3[3][89] , \w3[3][88] , \w3[3][87] , \w3[3][86] , \w3[3][85] ,
         \w3[3][84] , \w3[3][83] , \w3[3][82] , \w3[3][81] , \w3[3][80] ,
         \w3[3][79] , \w3[3][78] , \w3[3][77] , \w3[3][76] , \w3[3][75] ,
         \w3[3][74] , \w3[3][73] , \w3[3][72] , \w3[3][71] , \w3[3][70] ,
         \w3[3][69] , \w3[3][68] , \w3[3][67] , \w3[3][66] , \w3[3][65] ,
         \w3[3][64] , \w3[3][63] , \w3[3][62] , \w3[3][61] , \w3[3][60] ,
         \w3[3][59] , \w3[3][58] , \w3[3][57] , \w3[3][56] , \w3[3][55] ,
         \w3[3][54] , \w3[3][53] , \w3[3][52] , \w3[3][51] , \w3[3][50] ,
         \w3[3][49] , \w3[3][48] , \w3[3][47] , \w3[3][46] , \w3[3][45] ,
         \w3[3][44] , \w3[3][43] , \w3[3][42] , \w3[3][41] , \w3[3][40] ,
         \w3[3][39] , \w3[3][38] , \w3[3][37] , \w3[3][36] , \w3[3][35] ,
         \w3[3][34] , \w3[3][33] , \w3[3][32] , \w3[3][31] , \w3[3][30] ,
         \w3[3][29] , \w3[3][28] , \w3[3][27] , \w3[3][26] , \w3[3][25] ,
         \w3[3][24] , \w3[3][23] , \w3[3][22] , \w3[3][21] , \w3[3][20] ,
         \w3[3][19] , \w3[3][18] , \w3[3][17] , \w3[3][16] , \w3[3][15] ,
         \w3[3][14] , \w3[3][13] , \w3[3][12] , \w3[3][11] , \w3[3][10] ,
         \w3[3][9] , \w3[3][8] , \w3[3][7] , \w3[3][6] , \w3[3][5] ,
         \w3[3][4] , \w3[3][3] , \w3[3][2] , \w3[3][1] , \w3[3][0] ,
         \w3[2][127] , \w3[2][126] , \w3[2][125] , \w3[2][124] , \w3[2][123] ,
         \w3[2][122] , \w3[2][121] , \w3[2][120] , \w3[2][119] , \w3[2][118] ,
         \w3[2][117] , \w3[2][116] , \w3[2][115] , \w3[2][114] , \w3[2][113] ,
         \w3[2][112] , \w3[2][111] , \w3[2][110] , \w3[2][109] , \w3[2][108] ,
         \w3[2][107] , \w3[2][106] , \w3[2][105] , \w3[2][104] , \w3[2][103] ,
         \w3[2][102] , \w3[2][101] , \w3[2][100] , \w3[2][99] , \w3[2][98] ,
         \w3[2][97] , \w3[2][96] , \w3[2][95] , \w3[2][94] , \w3[2][93] ,
         \w3[2][92] , \w3[2][91] , \w3[2][90] , \w3[2][89] , \w3[2][88] ,
         \w3[2][87] , \w3[2][86] , \w3[2][85] , \w3[2][84] , \w3[2][83] ,
         \w3[2][82] , \w3[2][81] , \w3[2][80] , \w3[2][79] , \w3[2][78] ,
         \w3[2][77] , \w3[2][76] , \w3[2][75] , \w3[2][74] , \w3[2][73] ,
         \w3[2][72] , \w3[2][71] , \w3[2][70] , \w3[2][69] , \w3[2][68] ,
         \w3[2][67] , \w3[2][66] , \w3[2][65] , \w3[2][64] , \w3[2][63] ,
         \w3[2][62] , \w3[2][61] , \w3[2][60] , \w3[2][59] , \w3[2][58] ,
         \w3[2][57] , \w3[2][56] , \w3[2][55] , \w3[2][54] , \w3[2][53] ,
         \w3[2][52] , \w3[2][51] , \w3[2][50] , \w3[2][49] , \w3[2][48] ,
         \w3[2][47] , \w3[2][46] , \w3[2][45] , \w3[2][44] , \w3[2][43] ,
         \w3[2][42] , \w3[2][41] , \w3[2][40] , \w3[2][39] , \w3[2][38] ,
         \w3[2][37] , \w3[2][36] , \w3[2][35] , \w3[2][34] , \w3[2][33] ,
         \w3[2][32] , \w3[2][31] , \w3[2][30] , \w3[2][29] , \w3[2][28] ,
         \w3[2][27] , \w3[2][26] , \w3[2][25] , \w3[2][24] , \w3[2][23] ,
         \w3[2][22] , \w3[2][21] , \w3[2][20] , \w3[2][19] , \w3[2][18] ,
         \w3[2][17] , \w3[2][16] , \w3[2][15] , \w3[2][14] , \w3[2][13] ,
         \w3[2][12] , \w3[2][11] , \w3[2][10] , \w3[2][9] , \w3[2][8] ,
         \w3[2][7] , \w3[2][6] , \w3[2][5] , \w3[2][4] , \w3[2][3] ,
         \w3[2][2] , \w3[2][1] , \w3[2][0] , \w3[1][127] , \w3[1][126] ,
         \w3[1][125] , \w3[1][124] , \w3[1][123] , \w3[1][122] , \w3[1][121] ,
         \w3[1][120] , \w3[1][119] , \w3[1][118] , \w3[1][117] , \w3[1][116] ,
         \w3[1][115] , \w3[1][114] , \w3[1][113] , \w3[1][112] , \w3[1][111] ,
         \w3[1][110] , \w3[1][109] , \w3[1][108] , \w3[1][107] , \w3[1][106] ,
         \w3[1][105] , \w3[1][104] , \w3[1][103] , \w3[1][102] , \w3[1][101] ,
         \w3[1][100] , \w3[1][99] , \w3[1][98] , \w3[1][97] , \w3[1][96] ,
         \w3[1][95] , \w3[1][94] , \w3[1][93] , \w3[1][92] , \w3[1][91] ,
         \w3[1][90] , \w3[1][89] , \w3[1][88] , \w3[1][87] , \w3[1][86] ,
         \w3[1][85] , \w3[1][84] , \w3[1][83] , \w3[1][82] , \w3[1][81] ,
         \w3[1][80] , \w3[1][79] , \w3[1][78] , \w3[1][77] , \w3[1][76] ,
         \w3[1][75] , \w3[1][74] , \w3[1][73] , \w3[1][72] , \w3[1][71] ,
         \w3[1][70] , \w3[1][69] , \w3[1][68] , \w3[1][67] , \w3[1][66] ,
         \w3[1][65] , \w3[1][64] , \w3[1][63] , \w3[1][62] , \w3[1][61] ,
         \w3[1][60] , \w3[1][59] , \w3[1][58] , \w3[1][57] , \w3[1][56] ,
         \w3[1][55] , \w3[1][54] , \w3[1][53] , \w3[1][52] , \w3[1][51] ,
         \w3[1][50] , \w3[1][49] , \w3[1][48] , \w3[1][47] , \w3[1][46] ,
         \w3[1][45] , \w3[1][44] , \w3[1][43] , \w3[1][42] , \w3[1][41] ,
         \w3[1][40] , \w3[1][39] , \w3[1][38] , \w3[1][37] , \w3[1][36] ,
         \w3[1][35] , \w3[1][34] , \w3[1][33] , \w3[1][32] , \w3[1][31] ,
         \w3[1][30] , \w3[1][29] , \w3[1][28] , \w3[1][27] , \w3[1][26] ,
         \w3[1][25] , \w3[1][24] , \w3[1][23] , \w3[1][22] , \w3[1][21] ,
         \w3[1][20] , \w3[1][19] , \w3[1][18] , \w3[1][17] , \w3[1][16] ,
         \w3[1][15] , \w3[1][14] , \w3[1][13] , \w3[1][12] , \w3[1][11] ,
         \w3[1][10] , \w3[1][9] , \w3[1][8] , \w3[1][7] , \w3[1][6] ,
         \w3[1][5] , \w3[1][4] , \w3[1][3] , \w3[1][2] , \w3[1][1] ,
         \w3[1][0] , \w3[0][127] , \w3[0][126] , \w3[0][125] , \w3[0][124] ,
         \w3[0][123] , \w3[0][122] , \w3[0][121] , \w3[0][120] , \w3[0][119] ,
         \w3[0][118] , \w3[0][117] , \w3[0][116] , \w3[0][115] , \w3[0][114] ,
         \w3[0][113] , \w3[0][112] , \w3[0][111] , \w3[0][110] , \w3[0][109] ,
         \w3[0][108] , \w3[0][107] , \w3[0][106] , \w3[0][105] , \w3[0][104] ,
         \w3[0][103] , \w3[0][102] , \w3[0][101] , \w3[0][100] , \w3[0][99] ,
         \w3[0][98] , \w3[0][97] , \w3[0][96] , \w3[0][95] , \w3[0][94] ,
         \w3[0][93] , \w3[0][92] , \w3[0][91] , \w3[0][90] , \w3[0][89] ,
         \w3[0][88] , \w3[0][87] , \w3[0][86] , \w3[0][85] , \w3[0][84] ,
         \w3[0][83] , \w3[0][82] , \w3[0][81] , \w3[0][80] , \w3[0][79] ,
         \w3[0][78] , \w3[0][77] , \w3[0][76] , \w3[0][75] , \w3[0][74] ,
         \w3[0][73] , \w3[0][72] , \w3[0][71] , \w3[0][70] , \w3[0][69] ,
         \w3[0][68] , \w3[0][67] , \w3[0][66] , \w3[0][65] , \w3[0][64] ,
         \w3[0][63] , \w3[0][62] , \w3[0][61] , \w3[0][60] , \w3[0][59] ,
         \w3[0][58] , \w3[0][57] , \w3[0][56] , \w3[0][55] , \w3[0][54] ,
         \w3[0][53] , \w3[0][52] , \w3[0][51] , \w3[0][50] , \w3[0][49] ,
         \w3[0][48] , \w3[0][47] , \w3[0][46] , \w3[0][45] , \w3[0][44] ,
         \w3[0][43] , \w3[0][42] , \w3[0][41] , \w3[0][40] , \w3[0][39] ,
         \w3[0][38] , \w3[0][37] , \w3[0][36] , \w3[0][35] , \w3[0][34] ,
         \w3[0][33] , \w3[0][32] , \w3[0][31] , \w3[0][30] , \w3[0][29] ,
         \w3[0][28] , \w3[0][27] , \w3[0][26] , \w3[0][25] , \w3[0][24] ,
         \w3[0][23] , \w3[0][22] , \w3[0][21] , \w3[0][20] , \w3[0][19] ,
         \w3[0][18] , \w3[0][17] , \w3[0][16] , \w3[0][15] , \w3[0][14] ,
         \w3[0][13] , \w3[0][12] , \w3[0][11] , \w3[0][10] , \w3[0][9] ,
         \w3[0][8] , \w3[0][7] , \w3[0][6] , \w3[0][5] , \w3[0][4] ,
         \w3[0][3] , \w3[0][2] , \w3[0][1] , \w3[0][0] , n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136;
  wire   [127:0] state;

  SubBytes_2 \SUBBYTES[0].a  ( .x({\w1[0][127] , \w1[0][126] , \w1[0][125] , 
        \w1[0][124] , \w1[0][123] , \w1[0][122] , \w1[0][121] , \w1[0][120] , 
        \w1[0][119] , \w1[0][118] , \w1[0][117] , \w1[0][116] , \w1[0][115] , 
        \w1[0][114] , \w1[0][113] , \w1[0][112] , \w1[0][111] , \w1[0][110] , 
        \w1[0][109] , \w1[0][108] , \w1[0][107] , \w1[0][106] , \w1[0][105] , 
        \w1[0][104] , \w1[0][103] , \w1[0][102] , \w1[0][101] , \w1[0][100] , 
        \w1[0][99] , \w1[0][98] , \w1[0][97] , \w1[0][96] , \w1[0][95] , 
        \w1[0][94] , \w1[0][93] , \w1[0][92] , \w1[0][91] , \w1[0][90] , 
        \w1[0][89] , \w1[0][88] , \w1[0][87] , \w1[0][86] , \w1[0][85] , 
        \w1[0][84] , \w1[0][83] , \w1[0][82] , \w1[0][81] , \w1[0][80] , 
        \w1[0][79] , \w1[0][78] , \w1[0][77] , \w1[0][76] , \w1[0][75] , 
        \w1[0][74] , \w1[0][73] , \w1[0][72] , \w1[0][71] , \w1[0][70] , 
        \w1[0][69] , \w1[0][68] , \w1[0][67] , \w1[0][66] , \w1[0][65] , 
        \w1[0][64] , \w1[0][63] , \w1[0][62] , \w1[0][61] , \w1[0][60] , 
        \w1[0][59] , \w1[0][58] , \w1[0][57] , \w1[0][56] , \w1[0][55] , 
        \w1[0][54] , \w1[0][53] , \w1[0][52] , \w1[0][51] , \w1[0][50] , 
        \w1[0][49] , \w1[0][48] , \w1[0][47] , \w1[0][46] , \w1[0][45] , 
        \w1[0][44] , \w1[0][43] , \w1[0][42] , \w1[0][41] , \w1[0][40] , 
        \w1[0][39] , \w1[0][38] , \w1[0][37] , \w1[0][36] , \w1[0][35] , 
        \w1[0][34] , \w1[0][33] , \w1[0][32] , \w1[0][31] , \w1[0][30] , 
        \w1[0][29] , \w1[0][28] , \w1[0][27] , \w1[0][26] , \w1[0][25] , 
        \w1[0][24] , \w1[0][23] , \w1[0][22] , \w1[0][21] , \w1[0][20] , 
        \w1[0][19] , \w1[0][18] , \w1[0][17] , \w1[0][16] , \w1[0][15] , 
        \w1[0][14] , \w1[0][13] , \w1[0][12] , \w1[0][11] , \w1[0][10] , 
        \w1[0][9] , \w1[0][8] , \w1[0][7] , \w1[0][6] , \w1[0][5] , \w1[0][4] , 
        \w1[0][3] , \w1[0][2] , \w1[0][1] , \w1[0][0] }), .z({\w3[0][127] , 
        \w3[0][126] , \w3[0][125] , \w3[0][124] , \w3[0][123] , \w3[0][122] , 
        \w3[0][121] , \w3[0][120] , \w3[0][23] , \w3[0][22] , \w3[0][21] , 
        \w3[0][20] , \w3[0][19] , \w3[0][18] , \w3[0][17] , \w3[0][16] , 
        \w3[0][47] , \w3[0][46] , \w3[0][45] , \w3[0][44] , \w3[0][43] , 
        \w3[0][42] , \w3[0][41] , \w3[0][40] , \w3[0][71] , \w3[0][70] , 
        \w3[0][69] , \w3[0][68] , \w3[0][67] , \w3[0][66] , \w3[0][65] , 
        \w3[0][64] , \w3[0][95] , \w3[0][94] , \w3[0][93] , \w3[0][92] , 
        \w3[0][91] , \w3[0][90] , \w3[0][89] , \w3[0][88] , \w3[0][119] , 
        \w3[0][118] , \w3[0][117] , \w3[0][116] , \w3[0][115] , \w3[0][114] , 
        \w3[0][113] , \w3[0][112] , \w3[0][15] , \w3[0][14] , \w3[0][13] , 
        \w3[0][12] , \w3[0][11] , \w3[0][10] , \w3[0][9] , \w3[0][8] , 
        \w3[0][39] , \w3[0][38] , \w3[0][37] , \w3[0][36] , \w3[0][35] , 
        \w3[0][34] , \w3[0][33] , \w3[0][32] , \w3[0][63] , \w3[0][62] , 
        \w3[0][61] , \w3[0][60] , \w3[0][59] , \w3[0][58] , \w3[0][57] , 
        \w3[0][56] , \w3[0][87] , \w3[0][86] , \w3[0][85] , \w3[0][84] , 
        \w3[0][83] , \w3[0][82] , \w3[0][81] , \w3[0][80] , \w3[0][111] , 
        \w3[0][110] , \w3[0][109] , \w3[0][108] , \w3[0][107] , \w3[0][106] , 
        \w3[0][105] , \w3[0][104] , \w3[0][7] , \w3[0][6] , \w3[0][5] , 
        \w3[0][4] , \w3[0][3] , \w3[0][2] , \w3[0][1] , \w3[0][0] , 
        \w3[0][31] , \w3[0][30] , \w3[0][29] , \w3[0][28] , \w3[0][27] , 
        \w3[0][26] , \w3[0][25] , \w3[0][24] , \w3[0][55] , \w3[0][54] , 
        \w3[0][53] , \w3[0][52] , \w3[0][51] , \w3[0][50] , \w3[0][49] , 
        \w3[0][48] , \w3[0][79] , \w3[0][78] , \w3[0][77] , \w3[0][76] , 
        \w3[0][75] , \w3[0][74] , \w3[0][73] , \w3[0][72] , \w3[0][103] , 
        \w3[0][102] , \w3[0][101] , \w3[0][100] , \w3[0][99] , \w3[0][98] , 
        \w3[0][97] , \w3[0][96] }) );
  SubBytes_6 \SUBBYTES[1].a  ( .x({\w1[1][127] , \w1[1][126] , \w1[1][125] , 
        \w1[1][124] , \w1[1][123] , \w1[1][122] , \w1[1][121] , \w1[1][120] , 
        \w1[1][119] , \w1[1][118] , \w1[1][117] , \w1[1][116] , \w1[1][115] , 
        \w1[1][114] , \w1[1][113] , \w1[1][112] , \w1[1][111] , \w1[1][110] , 
        \w1[1][109] , \w1[1][108] , \w1[1][107] , \w1[1][106] , \w1[1][105] , 
        \w1[1][104] , \w1[1][103] , \w1[1][102] , \w1[1][101] , \w1[1][100] , 
        \w1[1][99] , \w1[1][98] , \w1[1][97] , \w1[1][96] , \w1[1][95] , 
        \w1[1][94] , \w1[1][93] , \w1[1][92] , \w1[1][91] , \w1[1][90] , 
        \w1[1][89] , \w1[1][88] , \w1[1][87] , \w1[1][86] , \w1[1][85] , 
        \w1[1][84] , \w1[1][83] , \w1[1][82] , \w1[1][81] , \w1[1][80] , 
        \w1[1][79] , \w1[1][78] , \w1[1][77] , \w1[1][76] , \w1[1][75] , 
        \w1[1][74] , \w1[1][73] , \w1[1][72] , \w1[1][71] , \w1[1][70] , 
        \w1[1][69] , \w1[1][68] , \w1[1][67] , \w1[1][66] , \w1[1][65] , 
        \w1[1][64] , \w1[1][63] , \w1[1][62] , \w1[1][61] , \w1[1][60] , 
        \w1[1][59] , \w1[1][58] , \w1[1][57] , \w1[1][56] , \w1[1][55] , 
        \w1[1][54] , \w1[1][53] , \w1[1][52] , \w1[1][51] , \w1[1][50] , 
        \w1[1][49] , \w1[1][48] , \w1[1][47] , \w1[1][46] , \w1[1][45] , 
        \w1[1][44] , \w1[1][43] , \w1[1][42] , \w1[1][41] , \w1[1][40] , 
        \w1[1][39] , \w1[1][38] , \w1[1][37] , \w1[1][36] , \w1[1][35] , 
        \w1[1][34] , \w1[1][33] , \w1[1][32] , \w1[1][31] , \w1[1][30] , 
        \w1[1][29] , \w1[1][28] , \w1[1][27] , \w1[1][26] , \w1[1][25] , 
        \w1[1][24] , \w1[1][23] , \w1[1][22] , \w1[1][21] , \w1[1][20] , 
        \w1[1][19] , \w1[1][18] , \w1[1][17] , \w1[1][16] , \w1[1][15] , 
        \w1[1][14] , \w1[1][13] , \w1[1][12] , \w1[1][11] , \w1[1][10] , 
        \w1[1][9] , \w1[1][8] , \w1[1][7] , \w1[1][6] , \w1[1][5] , \w1[1][4] , 
        \w1[1][3] , \w1[1][2] , \w1[1][1] , \w1[1][0] }), .z({\w3[1][127] , 
        \w3[1][126] , \w3[1][125] , \w3[1][124] , \w3[1][123] , \w3[1][122] , 
        \w3[1][121] , \w3[1][120] , \w3[1][23] , \w3[1][22] , \w3[1][21] , 
        \w3[1][20] , \w3[1][19] , \w3[1][18] , \w3[1][17] , \w3[1][16] , 
        \w3[1][47] , \w3[1][46] , \w3[1][45] , \w3[1][44] , \w3[1][43] , 
        \w3[1][42] , \w3[1][41] , \w3[1][40] , \w3[1][71] , \w3[1][70] , 
        \w3[1][69] , \w3[1][68] , \w3[1][67] , \w3[1][66] , \w3[1][65] , 
        \w3[1][64] , \w3[1][95] , \w3[1][94] , \w3[1][93] , \w3[1][92] , 
        \w3[1][91] , \w3[1][90] , \w3[1][89] , \w3[1][88] , \w3[1][119] , 
        \w3[1][118] , \w3[1][117] , \w3[1][116] , \w3[1][115] , \w3[1][114] , 
        \w3[1][113] , \w3[1][112] , \w3[1][15] , \w3[1][14] , \w3[1][13] , 
        \w3[1][12] , \w3[1][11] , \w3[1][10] , \w3[1][9] , \w3[1][8] , 
        \w3[1][39] , \w3[1][38] , \w3[1][37] , \w3[1][36] , \w3[1][35] , 
        \w3[1][34] , \w3[1][33] , \w3[1][32] , \w3[1][63] , \w3[1][62] , 
        \w3[1][61] , \w3[1][60] , \w3[1][59] , \w3[1][58] , \w3[1][57] , 
        \w3[1][56] , \w3[1][87] , \w3[1][86] , \w3[1][85] , \w3[1][84] , 
        \w3[1][83] , \w3[1][82] , \w3[1][81] , \w3[1][80] , \w3[1][111] , 
        \w3[1][110] , \w3[1][109] , \w3[1][108] , \w3[1][107] , \w3[1][106] , 
        \w3[1][105] , \w3[1][104] , \w3[1][7] , \w3[1][6] , \w3[1][5] , 
        \w3[1][4] , \w3[1][3] , \w3[1][2] , \w3[1][1] , \w3[1][0] , 
        \w3[1][31] , \w3[1][30] , \w3[1][29] , \w3[1][28] , \w3[1][27] , 
        \w3[1][26] , \w3[1][25] , \w3[1][24] , \w3[1][55] , \w3[1][54] , 
        \w3[1][53] , \w3[1][52] , \w3[1][51] , \w3[1][50] , \w3[1][49] , 
        \w3[1][48] , \w3[1][79] , \w3[1][78] , \w3[1][77] , \w3[1][76] , 
        \w3[1][75] , \w3[1][74] , \w3[1][73] , \w3[1][72] , \w3[1][103] , 
        \w3[1][102] , \w3[1][101] , \w3[1][100] , \w3[1][99] , \w3[1][98] , 
        \w3[1][97] , \w3[1][96] }) );
  SubBytes_5 \SUBBYTES[2].a  ( .x({\w1[2][127] , \w1[2][126] , \w1[2][125] , 
        \w1[2][124] , \w1[2][123] , \w1[2][122] , \w1[2][121] , \w1[2][120] , 
        \w1[2][119] , \w1[2][118] , \w1[2][117] , \w1[2][116] , \w1[2][115] , 
        \w1[2][114] , \w1[2][113] , \w1[2][112] , \w1[2][111] , \w1[2][110] , 
        \w1[2][109] , \w1[2][108] , \w1[2][107] , \w1[2][106] , \w1[2][105] , 
        \w1[2][104] , \w1[2][103] , \w1[2][102] , \w1[2][101] , \w1[2][100] , 
        \w1[2][99] , \w1[2][98] , \w1[2][97] , \w1[2][96] , \w1[2][95] , 
        \w1[2][94] , \w1[2][93] , \w1[2][92] , \w1[2][91] , \w1[2][90] , 
        \w1[2][89] , \w1[2][88] , \w1[2][87] , \w1[2][86] , \w1[2][85] , 
        \w1[2][84] , \w1[2][83] , \w1[2][82] , \w1[2][81] , \w1[2][80] , 
        \w1[2][79] , \w1[2][78] , \w1[2][77] , \w1[2][76] , \w1[2][75] , 
        \w1[2][74] , \w1[2][73] , \w1[2][72] , \w1[2][71] , \w1[2][70] , 
        \w1[2][69] , \w1[2][68] , \w1[2][67] , \w1[2][66] , \w1[2][65] , 
        \w1[2][64] , \w1[2][63] , \w1[2][62] , \w1[2][61] , \w1[2][60] , 
        \w1[2][59] , \w1[2][58] , \w1[2][57] , \w1[2][56] , \w1[2][55] , 
        \w1[2][54] , \w1[2][53] , \w1[2][52] , \w1[2][51] , \w1[2][50] , 
        \w1[2][49] , \w1[2][48] , \w1[2][47] , \w1[2][46] , \w1[2][45] , 
        \w1[2][44] , \w1[2][43] , \w1[2][42] , \w1[2][41] , \w1[2][40] , 
        \w1[2][39] , \w1[2][38] , \w1[2][37] , \w1[2][36] , \w1[2][35] , 
        \w1[2][34] , \w1[2][33] , \w1[2][32] , \w1[2][31] , \w1[2][30] , 
        \w1[2][29] , \w1[2][28] , \w1[2][27] , \w1[2][26] , \w1[2][25] , 
        \w1[2][24] , \w1[2][23] , \w1[2][22] , \w1[2][21] , \w1[2][20] , 
        \w1[2][19] , \w1[2][18] , \w1[2][17] , \w1[2][16] , \w1[2][15] , 
        \w1[2][14] , \w1[2][13] , \w1[2][12] , \w1[2][11] , \w1[2][10] , 
        \w1[2][9] , \w1[2][8] , \w1[2][7] , \w1[2][6] , \w1[2][5] , \w1[2][4] , 
        \w1[2][3] , \w1[2][2] , \w1[2][1] , \w1[2][0] }), .z({\w3[2][127] , 
        \w3[2][126] , \w3[2][125] , \w3[2][124] , \w3[2][123] , \w3[2][122] , 
        \w3[2][121] , \w3[2][120] , \w3[2][23] , \w3[2][22] , \w3[2][21] , 
        \w3[2][20] , \w3[2][19] , \w3[2][18] , \w3[2][17] , \w3[2][16] , 
        \w3[2][47] , \w3[2][46] , \w3[2][45] , \w3[2][44] , \w3[2][43] , 
        \w3[2][42] , \w3[2][41] , \w3[2][40] , \w3[2][71] , \w3[2][70] , 
        \w3[2][69] , \w3[2][68] , \w3[2][67] , \w3[2][66] , \w3[2][65] , 
        \w3[2][64] , \w3[2][95] , \w3[2][94] , \w3[2][93] , \w3[2][92] , 
        \w3[2][91] , \w3[2][90] , \w3[2][89] , \w3[2][88] , \w3[2][119] , 
        \w3[2][118] , \w3[2][117] , \w3[2][116] , \w3[2][115] , \w3[2][114] , 
        \w3[2][113] , \w3[2][112] , \w3[2][15] , \w3[2][14] , \w3[2][13] , 
        \w3[2][12] , \w3[2][11] , \w3[2][10] , \w3[2][9] , \w3[2][8] , 
        \w3[2][39] , \w3[2][38] , \w3[2][37] , \w3[2][36] , \w3[2][35] , 
        \w3[2][34] , \w3[2][33] , \w3[2][32] , \w3[2][63] , \w3[2][62] , 
        \w3[2][61] , \w3[2][60] , \w3[2][59] , \w3[2][58] , \w3[2][57] , 
        \w3[2][56] , \w3[2][87] , \w3[2][86] , \w3[2][85] , \w3[2][84] , 
        \w3[2][83] , \w3[2][82] , \w3[2][81] , \w3[2][80] , \w3[2][111] , 
        \w3[2][110] , \w3[2][109] , \w3[2][108] , \w3[2][107] , \w3[2][106] , 
        \w3[2][105] , \w3[2][104] , \w3[2][7] , \w3[2][6] , \w3[2][5] , 
        \w3[2][4] , \w3[2][3] , \w3[2][2] , \w3[2][1] , \w3[2][0] , 
        \w3[2][31] , \w3[2][30] , \w3[2][29] , \w3[2][28] , \w3[2][27] , 
        \w3[2][26] , \w3[2][25] , \w3[2][24] , \w3[2][55] , \w3[2][54] , 
        \w3[2][53] , \w3[2][52] , \w3[2][51] , \w3[2][50] , \w3[2][49] , 
        \w3[2][48] , \w3[2][79] , \w3[2][78] , \w3[2][77] , \w3[2][76] , 
        \w3[2][75] , \w3[2][74] , \w3[2][73] , \w3[2][72] , \w3[2][103] , 
        \w3[2][102] , \w3[2][101] , \w3[2][100] , \w3[2][99] , \w3[2][98] , 
        \w3[2][97] , \w3[2][96] }) );
  SubBytes_4 \SUBBYTES[3].a  ( .x({\w1[3][127] , \w1[3][126] , \w1[3][125] , 
        \w1[3][124] , \w1[3][123] , \w1[3][122] , \w1[3][121] , \w1[3][120] , 
        \w1[3][119] , \w1[3][118] , \w1[3][117] , \w1[3][116] , \w1[3][115] , 
        \w1[3][114] , \w1[3][113] , \w1[3][112] , \w1[3][111] , \w1[3][110] , 
        \w1[3][109] , \w1[3][108] , \w1[3][107] , \w1[3][106] , \w1[3][105] , 
        \w1[3][104] , \w1[3][103] , \w1[3][102] , \w1[3][101] , \w1[3][100] , 
        \w1[3][99] , \w1[3][98] , \w1[3][97] , \w1[3][96] , \w1[3][95] , 
        \w1[3][94] , \w1[3][93] , \w1[3][92] , \w1[3][91] , \w1[3][90] , 
        \w1[3][89] , \w1[3][88] , \w1[3][87] , \w1[3][86] , \w1[3][85] , 
        \w1[3][84] , \w1[3][83] , \w1[3][82] , \w1[3][81] , \w1[3][80] , 
        \w1[3][79] , \w1[3][78] , \w1[3][77] , \w1[3][76] , \w1[3][75] , 
        \w1[3][74] , \w1[3][73] , \w1[3][72] , \w1[3][71] , \w1[3][70] , 
        \w1[3][69] , \w1[3][68] , \w1[3][67] , \w1[3][66] , \w1[3][65] , 
        \w1[3][64] , \w1[3][63] , \w1[3][62] , \w1[3][61] , \w1[3][60] , 
        \w1[3][59] , \w1[3][58] , \w1[3][57] , \w1[3][56] , \w1[3][55] , 
        \w1[3][54] , \w1[3][53] , \w1[3][52] , \w1[3][51] , \w1[3][50] , 
        \w1[3][49] , \w1[3][48] , \w1[3][47] , \w1[3][46] , \w1[3][45] , 
        \w1[3][44] , \w1[3][43] , \w1[3][42] , \w1[3][41] , \w1[3][40] , 
        \w1[3][39] , \w1[3][38] , \w1[3][37] , \w1[3][36] , \w1[3][35] , 
        \w1[3][34] , \w1[3][33] , \w1[3][32] , \w1[3][31] , \w1[3][30] , 
        \w1[3][29] , \w1[3][28] , \w1[3][27] , \w1[3][26] , \w1[3][25] , 
        \w1[3][24] , \w1[3][23] , \w1[3][22] , \w1[3][21] , \w1[3][20] , 
        \w1[3][19] , \w1[3][18] , \w1[3][17] , \w1[3][16] , \w1[3][15] , 
        \w1[3][14] , \w1[3][13] , \w1[3][12] , \w1[3][11] , \w1[3][10] , 
        \w1[3][9] , \w1[3][8] , \w1[3][7] , \w1[3][6] , \w1[3][5] , \w1[3][4] , 
        \w1[3][3] , \w1[3][2] , \w1[3][1] , \w1[3][0] }), .z({\w3[3][127] , 
        \w3[3][126] , \w3[3][125] , \w3[3][124] , \w3[3][123] , \w3[3][122] , 
        \w3[3][121] , \w3[3][120] , \w3[3][23] , \w3[3][22] , \w3[3][21] , 
        \w3[3][20] , \w3[3][19] , \w3[3][18] , \w3[3][17] , \w3[3][16] , 
        \w3[3][47] , \w3[3][46] , \w3[3][45] , \w3[3][44] , \w3[3][43] , 
        \w3[3][42] , \w3[3][41] , \w3[3][40] , \w3[3][71] , \w3[3][70] , 
        \w3[3][69] , \w3[3][68] , \w3[3][67] , \w3[3][66] , \w3[3][65] , 
        \w3[3][64] , \w3[3][95] , \w3[3][94] , \w3[3][93] , \w3[3][92] , 
        \w3[3][91] , \w3[3][90] , \w3[3][89] , \w3[3][88] , \w3[3][119] , 
        \w3[3][118] , \w3[3][117] , \w3[3][116] , \w3[3][115] , \w3[3][114] , 
        \w3[3][113] , \w3[3][112] , \w3[3][15] , \w3[3][14] , \w3[3][13] , 
        \w3[3][12] , \w3[3][11] , \w3[3][10] , \w3[3][9] , \w3[3][8] , 
        \w3[3][39] , \w3[3][38] , \w3[3][37] , \w3[3][36] , \w3[3][35] , 
        \w3[3][34] , \w3[3][33] , \w3[3][32] , \w3[3][63] , \w3[3][62] , 
        \w3[3][61] , \w3[3][60] , \w3[3][59] , \w3[3][58] , \w3[3][57] , 
        \w3[3][56] , \w3[3][87] , \w3[3][86] , \w3[3][85] , \w3[3][84] , 
        \w3[3][83] , \w3[3][82] , \w3[3][81] , \w3[3][80] , \w3[3][111] , 
        \w3[3][110] , \w3[3][109] , \w3[3][108] , \w3[3][107] , \w3[3][106] , 
        \w3[3][105] , \w3[3][104] , \w3[3][7] , \w3[3][6] , \w3[3][5] , 
        \w3[3][4] , \w3[3][3] , \w3[3][2] , \w3[3][1] , \w3[3][0] , 
        \w3[3][31] , \w3[3][30] , \w3[3][29] , \w3[3][28] , \w3[3][27] , 
        \w3[3][26] , \w3[3][25] , \w3[3][24] , \w3[3][55] , \w3[3][54] , 
        \w3[3][53] , \w3[3][52] , \w3[3][51] , \w3[3][50] , \w3[3][49] , 
        \w3[3][48] , \w3[3][79] , \w3[3][78] , \w3[3][77] , \w3[3][76] , 
        \w3[3][75] , \w3[3][74] , \w3[3][73] , \w3[3][72] , \w3[3][103] , 
        \w3[3][102] , \w3[3][101] , \w3[3][100] , \w3[3][99] , \w3[3][98] , 
        \w3[3][97] , \w3[3][96] }) );
  SubBytes_3 \SUBBYTES[4].a  ( .x({\w1[4][127] , \w1[4][126] , \w1[4][125] , 
        \w1[4][124] , \w1[4][123] , \w1[4][122] , \w1[4][121] , \w1[4][120] , 
        \w1[4][119] , \w1[4][118] , \w1[4][117] , \w1[4][116] , \w1[4][115] , 
        \w1[4][114] , \w1[4][113] , \w1[4][112] , \w1[4][111] , \w1[4][110] , 
        \w1[4][109] , \w1[4][108] , \w1[4][107] , \w1[4][106] , \w1[4][105] , 
        \w1[4][104] , \w1[4][103] , \w1[4][102] , \w1[4][101] , \w1[4][100] , 
        \w1[4][99] , \w1[4][98] , \w1[4][97] , \w1[4][96] , \w1[4][95] , 
        \w1[4][94] , \w1[4][93] , \w1[4][92] , \w1[4][91] , \w1[4][90] , 
        \w1[4][89] , \w1[4][88] , \w1[4][87] , \w1[4][86] , \w1[4][85] , 
        \w1[4][84] , \w1[4][83] , \w1[4][82] , \w1[4][81] , \w1[4][80] , 
        \w1[4][79] , \w1[4][78] , \w1[4][77] , \w1[4][76] , \w1[4][75] , 
        \w1[4][74] , \w1[4][73] , \w1[4][72] , \w1[4][71] , \w1[4][70] , 
        \w1[4][69] , \w1[4][68] , \w1[4][67] , \w1[4][66] , \w1[4][65] , 
        \w1[4][64] , \w1[4][63] , \w1[4][62] , \w1[4][61] , \w1[4][60] , 
        \w1[4][59] , \w1[4][58] , \w1[4][57] , \w1[4][56] , \w1[4][55] , 
        \w1[4][54] , \w1[4][53] , \w1[4][52] , \w1[4][51] , \w1[4][50] , 
        \w1[4][49] , \w1[4][48] , \w1[4][47] , \w1[4][46] , \w1[4][45] , 
        \w1[4][44] , \w1[4][43] , \w1[4][42] , \w1[4][41] , \w1[4][40] , 
        \w1[4][39] , \w1[4][38] , \w1[4][37] , \w1[4][36] , \w1[4][35] , 
        \w1[4][34] , \w1[4][33] , \w1[4][32] , \w1[4][31] , \w1[4][30] , 
        \w1[4][29] , \w1[4][28] , \w1[4][27] , \w1[4][26] , \w1[4][25] , 
        \w1[4][24] , \w1[4][23] , \w1[4][22] , \w1[4][21] , \w1[4][20] , 
        \w1[4][19] , \w1[4][18] , \w1[4][17] , \w1[4][16] , \w1[4][15] , 
        \w1[4][14] , \w1[4][13] , \w1[4][12] , \w1[4][11] , \w1[4][10] , 
        \w1[4][9] , \w1[4][8] , \w1[4][7] , \w1[4][6] , \w1[4][5] , \w1[4][4] , 
        \w1[4][3] , \w1[4][2] , \w1[4][1] , \w1[4][0] }), .z({\w3[4][127] , 
        \w3[4][126] , \w3[4][125] , \w3[4][124] , \w3[4][123] , \w3[4][122] , 
        \w3[4][121] , \w3[4][120] , \w3[4][23] , \w3[4][22] , \w3[4][21] , 
        \w3[4][20] , \w3[4][19] , \w3[4][18] , \w3[4][17] , \w3[4][16] , 
        \w3[4][47] , \w3[4][46] , \w3[4][45] , \w3[4][44] , \w3[4][43] , 
        \w3[4][42] , \w3[4][41] , \w3[4][40] , \w3[4][71] , \w3[4][70] , 
        \w3[4][69] , \w3[4][68] , \w3[4][67] , \w3[4][66] , \w3[4][65] , 
        \w3[4][64] , \w3[4][95] , \w3[4][94] , \w3[4][93] , \w3[4][92] , 
        \w3[4][91] , \w3[4][90] , \w3[4][89] , \w3[4][88] , \w3[4][119] , 
        \w3[4][118] , \w3[4][117] , \w3[4][116] , \w3[4][115] , \w3[4][114] , 
        \w3[4][113] , \w3[4][112] , \w3[4][15] , \w3[4][14] , \w3[4][13] , 
        \w3[4][12] , \w3[4][11] , \w3[4][10] , \w3[4][9] , \w3[4][8] , 
        \w3[4][39] , \w3[4][38] , \w3[4][37] , \w3[4][36] , \w3[4][35] , 
        \w3[4][34] , \w3[4][33] , \w3[4][32] , \w3[4][63] , \w3[4][62] , 
        \w3[4][61] , \w3[4][60] , \w3[4][59] , \w3[4][58] , \w3[4][57] , 
        \w3[4][56] , \w3[4][87] , \w3[4][86] , \w3[4][85] , \w3[4][84] , 
        \w3[4][83] , \w3[4][82] , \w3[4][81] , \w3[4][80] , \w3[4][111] , 
        \w3[4][110] , \w3[4][109] , \w3[4][108] , \w3[4][107] , \w3[4][106] , 
        \w3[4][105] , \w3[4][104] , \w3[4][7] , \w3[4][6] , \w3[4][5] , 
        \w3[4][4] , \w3[4][3] , \w3[4][2] , \w3[4][1] , \w3[4][0] , 
        \w3[4][31] , \w3[4][30] , \w3[4][29] , \w3[4][28] , \w3[4][27] , 
        \w3[4][26] , \w3[4][25] , \w3[4][24] , \w3[4][55] , \w3[4][54] , 
        \w3[4][53] , \w3[4][52] , \w3[4][51] , \w3[4][50] , \w3[4][49] , 
        \w3[4][48] , \w3[4][79] , \w3[4][78] , \w3[4][77] , \w3[4][76] , 
        \w3[4][75] , \w3[4][74] , \w3[4][73] , \w3[4][72] , \w3[4][103] , 
        \w3[4][102] , \w3[4][101] , \w3[4][100] , \w3[4][99] , \w3[4][98] , 
        \w3[4][97] , \w3[4][96] }) );
  DFF init_reg ( .D(1'b1), .CLK(clk), .RST(rst), .Q(init) );
  DFF \state_reg[0]  ( .D(\w0[4][0] ), .CLK(clk), .RST(rst), .Q(state[0]) );
  DFF \state_reg[71]  ( .D(\w0[4][71] ), .CLK(clk), .RST(rst), .Q(state[71])
         );
  DFF \state_reg[88]  ( .D(\w0[4][88] ), .CLK(clk), .RST(rst), .Q(state[88])
         );
  DFF \state_reg[80]  ( .D(\w0[4][80] ), .CLK(clk), .RST(rst), .Q(state[80])
         );
  DFF \state_reg[81]  ( .D(\w0[4][81] ), .CLK(clk), .RST(rst), .Q(state[81])
         );
  DFF \state_reg[64]  ( .D(\w0[4][64] ), .CLK(clk), .RST(rst), .Q(state[64])
         );
  DFF \state_reg[72]  ( .D(\w0[4][72] ), .CLK(clk), .RST(rst), .Q(state[72])
         );
  DFF \state_reg[89]  ( .D(\w0[4][89] ), .CLK(clk), .RST(rst), .Q(state[89])
         );
  DFF \state_reg[82]  ( .D(\w0[4][82] ), .CLK(clk), .RST(rst), .Q(state[82])
         );
  DFF \state_reg[65]  ( .D(\w0[4][65] ), .CLK(clk), .RST(rst), .Q(state[65])
         );
  DFF \state_reg[73]  ( .D(\w0[4][73] ), .CLK(clk), .RST(rst), .Q(state[73])
         );
  DFF \state_reg[90]  ( .D(\w0[4][90] ), .CLK(clk), .RST(rst), .Q(state[90])
         );
  DFF \state_reg[83]  ( .D(\w0[4][83] ), .CLK(clk), .RST(rst), .Q(state[83])
         );
  DFF \state_reg[66]  ( .D(\w0[4][66] ), .CLK(clk), .RST(rst), .Q(state[66])
         );
  DFF \state_reg[74]  ( .D(\w0[4][74] ), .CLK(clk), .RST(rst), .Q(state[74])
         );
  DFF \state_reg[91]  ( .D(\w0[4][91] ), .CLK(clk), .RST(rst), .Q(state[91])
         );
  DFF \state_reg[75]  ( .D(\w0[4][75] ), .CLK(clk), .RST(rst), .Q(state[75])
         );
  DFF \state_reg[67]  ( .D(\w0[4][67] ), .CLK(clk), .RST(rst), .Q(state[67])
         );
  DFF \state_reg[84]  ( .D(\w0[4][84] ), .CLK(clk), .RST(rst), .Q(state[84])
         );
  DFF \state_reg[92]  ( .D(\w0[4][92] ), .CLK(clk), .RST(rst), .Q(state[92])
         );
  DFF \state_reg[76]  ( .D(\w0[4][76] ), .CLK(clk), .RST(rst), .Q(state[76])
         );
  DFF \state_reg[68]  ( .D(\w0[4][68] ), .CLK(clk), .RST(rst), .Q(state[68])
         );
  DFF \state_reg[85]  ( .D(\w0[4][85] ), .CLK(clk), .RST(rst), .Q(state[85])
         );
  DFF \state_reg[93]  ( .D(\w0[4][93] ), .CLK(clk), .RST(rst), .Q(state[93])
         );
  DFF \state_reg[86]  ( .D(\w0[4][86] ), .CLK(clk), .RST(rst), .Q(state[86])
         );
  DFF \state_reg[69]  ( .D(\w0[4][69] ), .CLK(clk), .RST(rst), .Q(state[69])
         );
  DFF \state_reg[77]  ( .D(\w0[4][77] ), .CLK(clk), .RST(rst), .Q(state[77])
         );
  DFF \state_reg[94]  ( .D(\w0[4][94] ), .CLK(clk), .RST(rst), .Q(state[94])
         );
  DFF \state_reg[78]  ( .D(\w0[4][78] ), .CLK(clk), .RST(rst), .Q(state[78])
         );
  DFF \state_reg[70]  ( .D(\w0[4][70] ), .CLK(clk), .RST(rst), .Q(state[70])
         );
  DFF \state_reg[87]  ( .D(\w0[4][87] ), .CLK(clk), .RST(rst), .Q(state[87])
         );
  DFF \state_reg[79]  ( .D(\w0[4][79] ), .CLK(clk), .RST(rst), .Q(state[79])
         );
  DFF \state_reg[95]  ( .D(\w0[4][95] ), .CLK(clk), .RST(rst), .Q(state[95])
         );
  DFF \state_reg[32]  ( .D(\w0[4][32] ), .CLK(clk), .RST(rst), .Q(state[32])
         );
  DFF \state_reg[56]  ( .D(\w0[4][56] ), .CLK(clk), .RST(rst), .Q(state[56])
         );
  DFF \state_reg[47]  ( .D(\w0[4][47] ), .CLK(clk), .RST(rst), .Q(state[47])
         );
  DFF \state_reg[57]  ( .D(\w0[4][57] ), .CLK(clk), .RST(rst), .Q(state[57])
         );
  DFF \state_reg[48]  ( .D(\w0[4][48] ), .CLK(clk), .RST(rst), .Q(state[48])
         );
  DFF \state_reg[33]  ( .D(\w0[4][33] ), .CLK(clk), .RST(rst), .Q(state[33])
         );
  DFF \state_reg[40]  ( .D(\w0[4][40] ), .CLK(clk), .RST(rst), .Q(state[40])
         );
  DFF \state_reg[58]  ( .D(\w0[4][58] ), .CLK(clk), .RST(rst), .Q(state[58])
         );
  DFF \state_reg[49]  ( .D(\w0[4][49] ), .CLK(clk), .RST(rst), .Q(state[49])
         );
  DFF \state_reg[34]  ( .D(\w0[4][34] ), .CLK(clk), .RST(rst), .Q(state[34])
         );
  DFF \state_reg[41]  ( .D(\w0[4][41] ), .CLK(clk), .RST(rst), .Q(state[41])
         );
  DFF \state_reg[50]  ( .D(\w0[4][50] ), .CLK(clk), .RST(rst), .Q(state[50])
         );
  DFF \state_reg[59]  ( .D(\w0[4][59] ), .CLK(clk), .RST(rst), .Q(state[59])
         );
  DFF \state_reg[35]  ( .D(\w0[4][35] ), .CLK(clk), .RST(rst), .Q(state[35])
         );
  DFF \state_reg[42]  ( .D(\w0[4][42] ), .CLK(clk), .RST(rst), .Q(state[42])
         );
  DFF \state_reg[60]  ( .D(\w0[4][60] ), .CLK(clk), .RST(rst), .Q(state[60])
         );
  DFF \state_reg[36]  ( .D(\w0[4][36] ), .CLK(clk), .RST(rst), .Q(state[36])
         );
  DFF \state_reg[51]  ( .D(\w0[4][51] ), .CLK(clk), .RST(rst), .Q(state[51])
         );
  DFF \state_reg[43]  ( .D(\w0[4][43] ), .CLK(clk), .RST(rst), .Q(state[43])
         );
  DFF \state_reg[61]  ( .D(\w0[4][61] ), .CLK(clk), .RST(rst), .Q(state[61])
         );
  DFF \state_reg[37]  ( .D(\w0[4][37] ), .CLK(clk), .RST(rst), .Q(state[37])
         );
  DFF \state_reg[52]  ( .D(\w0[4][52] ), .CLK(clk), .RST(rst), .Q(state[52])
         );
  DFF \state_reg[44]  ( .D(\w0[4][44] ), .CLK(clk), .RST(rst), .Q(state[44])
         );
  DFF \state_reg[53]  ( .D(\w0[4][53] ), .CLK(clk), .RST(rst), .Q(state[53])
         );
  DFF \state_reg[62]  ( .D(\w0[4][62] ), .CLK(clk), .RST(rst), .Q(state[62])
         );
  DFF \state_reg[38]  ( .D(\w0[4][38] ), .CLK(clk), .RST(rst), .Q(state[38])
         );
  DFF \state_reg[45]  ( .D(\w0[4][45] ), .CLK(clk), .RST(rst), .Q(state[45])
         );
  DFF \state_reg[63]  ( .D(\w0[4][63] ), .CLK(clk), .RST(rst), .Q(state[63])
         );
  DFF \state_reg[39]  ( .D(\w0[4][39] ), .CLK(clk), .RST(rst), .Q(state[39])
         );
  DFF \state_reg[55]  ( .D(\w0[4][55] ), .CLK(clk), .RST(rst), .Q(state[55])
         );
  DFF \state_reg[54]  ( .D(\w0[4][54] ), .CLK(clk), .RST(rst), .Q(state[54])
         );
  DFF \state_reg[46]  ( .D(\w0[4][46] ), .CLK(clk), .RST(rst), .Q(state[46])
         );
  DFF \state_reg[8]  ( .D(\w0[4][8] ), .CLK(clk), .RST(rst), .Q(state[8]) );
  DFF \state_reg[23]  ( .D(\w0[4][23] ), .CLK(clk), .RST(rst), .Q(state[23])
         );
  DFF \state_reg[1]  ( .D(\w0[4][1] ), .CLK(clk), .RST(rst), .Q(state[1]) );
  DFF \state_reg[16]  ( .D(\w0[4][16] ), .CLK(clk), .RST(rst), .Q(state[16])
         );
  DFF \state_reg[24]  ( .D(\w0[4][24] ), .CLK(clk), .RST(rst), .Q(state[24])
         );
  DFF \state_reg[9]  ( .D(\w0[4][9] ), .CLK(clk), .RST(rst), .Q(state[9]) );
  DFF \state_reg[10]  ( .D(\w0[4][10] ), .CLK(clk), .RST(rst), .Q(state[10])
         );
  DFF \state_reg[2]  ( .D(\w0[4][2] ), .CLK(clk), .RST(rst), .Q(state[2]) );
  DFF \state_reg[17]  ( .D(\w0[4][17] ), .CLK(clk), .RST(rst), .Q(state[17])
         );
  DFF \state_reg[25]  ( .D(\w0[4][25] ), .CLK(clk), .RST(rst), .Q(state[25])
         );
  DFF \state_reg[11]  ( .D(\w0[4][11] ), .CLK(clk), .RST(rst), .Q(state[11])
         );
  DFF \state_reg[3]  ( .D(\w0[4][3] ), .CLK(clk), .RST(rst), .Q(state[3]) );
  DFF \state_reg[18]  ( .D(\w0[4][18] ), .CLK(clk), .RST(rst), .Q(state[18])
         );
  DFF \state_reg[26]  ( .D(\w0[4][26] ), .CLK(clk), .RST(rst), .Q(state[26])
         );
  DFF \state_reg[12]  ( .D(\w0[4][12] ), .CLK(clk), .RST(rst), .Q(state[12])
         );
  DFF \state_reg[27]  ( .D(\w0[4][27] ), .CLK(clk), .RST(rst), .Q(state[27])
         );
  DFF \state_reg[19]  ( .D(\w0[4][19] ), .CLK(clk), .RST(rst), .Q(state[19])
         );
  DFF \state_reg[4]  ( .D(\w0[4][4] ), .CLK(clk), .RST(rst), .Q(state[4]) );
  DFF \state_reg[13]  ( .D(\w0[4][13] ), .CLK(clk), .RST(rst), .Q(state[13])
         );
  DFF \state_reg[28]  ( .D(\w0[4][28] ), .CLK(clk), .RST(rst), .Q(state[28])
         );
  DFF \state_reg[20]  ( .D(\w0[4][20] ), .CLK(clk), .RST(rst), .Q(state[20])
         );
  DFF \state_reg[5]  ( .D(\w0[4][5] ), .CLK(clk), .RST(rst), .Q(state[5]) );
  DFF \state_reg[14]  ( .D(\w0[4][14] ), .CLK(clk), .RST(rst), .Q(state[14])
         );
  DFF \state_reg[6]  ( .D(\w0[4][6] ), .CLK(clk), .RST(rst), .Q(state[6]) );
  DFF \state_reg[21]  ( .D(\w0[4][21] ), .CLK(clk), .RST(rst), .Q(state[21])
         );
  DFF \state_reg[29]  ( .D(\w0[4][29] ), .CLK(clk), .RST(rst), .Q(state[29])
         );
  DFF \state_reg[15]  ( .D(\w0[4][15] ), .CLK(clk), .RST(rst), .Q(state[15])
         );
  DFF \state_reg[30]  ( .D(\w0[4][30] ), .CLK(clk), .RST(rst), .Q(state[30])
         );
  DFF \state_reg[22]  ( .D(\w0[4][22] ), .CLK(clk), .RST(rst), .Q(state[22])
         );
  DFF \state_reg[7]  ( .D(\w0[4][7] ), .CLK(clk), .RST(rst), .Q(state[7]) );
  DFF \state_reg[31]  ( .D(\w0[4][31] ), .CLK(clk), .RST(rst), .Q(state[31])
         );
  DFF \state_reg[127]  ( .D(\w0[4][127] ), .CLK(clk), .RST(rst), .Q(state[127]) );
  DFF \state_reg[104]  ( .D(\w0[4][104] ), .CLK(clk), .RST(rst), .Q(state[104]) );
  DFF \state_reg[112]  ( .D(\w0[4][112] ), .CLK(clk), .RST(rst), .Q(state[112]) );
  DFF \state_reg[96]  ( .D(\w0[4][96] ), .CLK(clk), .RST(rst), .Q(state[96])
         );
  DFF \state_reg[113]  ( .D(\w0[4][113] ), .CLK(clk), .RST(rst), .Q(state[113]) );
  DFF \state_reg[105]  ( .D(\w0[4][105] ), .CLK(clk), .RST(rst), .Q(state[105]) );
  DFF \state_reg[120]  ( .D(\w0[4][120] ), .CLK(clk), .RST(rst), .Q(state[120]) );
  DFF \state_reg[97]  ( .D(\w0[4][97] ), .CLK(clk), .RST(rst), .Q(state[97])
         );
  DFF \state_reg[114]  ( .D(\w0[4][114] ), .CLK(clk), .RST(rst), .Q(state[114]) );
  DFF \state_reg[106]  ( .D(\w0[4][106] ), .CLK(clk), .RST(rst), .Q(state[106]) );
  DFF \state_reg[121]  ( .D(\w0[4][121] ), .CLK(clk), .RST(rst), .Q(state[121]) );
  DFF \state_reg[98]  ( .D(\w0[4][98] ), .CLK(clk), .RST(rst), .Q(state[98])
         );
  DFF \state_reg[115]  ( .D(\w0[4][115] ), .CLK(clk), .RST(rst), .Q(state[115]) );
  DFF \state_reg[107]  ( .D(\w0[4][107] ), .CLK(clk), .RST(rst), .Q(state[107]) );
  DFF \state_reg[122]  ( .D(\w0[4][122] ), .CLK(clk), .RST(rst), .Q(state[122]) );
  DFF \state_reg[116]  ( .D(\w0[4][116] ), .CLK(clk), .RST(rst), .Q(state[116]) );
  DFF \state_reg[108]  ( .D(\w0[4][108] ), .CLK(clk), .RST(rst), .Q(state[108]) );
  DFF \state_reg[99]  ( .D(\w0[4][99] ), .CLK(clk), .RST(rst), .Q(state[99])
         );
  DFF \state_reg[123]  ( .D(\w0[4][123] ), .CLK(clk), .RST(rst), .Q(state[123]) );
  DFF \state_reg[124]  ( .D(\w0[4][124] ), .CLK(clk), .RST(rst), .Q(state[124]) );
  DFF \state_reg[100]  ( .D(\w0[4][100] ), .CLK(clk), .RST(rst), .Q(state[100]) );
  DFF \state_reg[117]  ( .D(\w0[4][117] ), .CLK(clk), .RST(rst), .Q(state[117]) );
  DFF \state_reg[109]  ( .D(\w0[4][109] ), .CLK(clk), .RST(rst), .Q(state[109]) );
  DFF \state_reg[118]  ( .D(\w0[4][118] ), .CLK(clk), .RST(rst), .Q(state[118]) );
  DFF \state_reg[110]  ( .D(\w0[4][110] ), .CLK(clk), .RST(rst), .Q(state[110]) );
  DFF \state_reg[101]  ( .D(\w0[4][101] ), .CLK(clk), .RST(rst), .Q(state[101]) );
  DFF \state_reg[125]  ( .D(\w0[4][125] ), .CLK(clk), .RST(rst), .Q(state[125]) );
  DFF \state_reg[103]  ( .D(\w0[4][103] ), .CLK(clk), .RST(rst), .Q(state[103]) );
  DFF \state_reg[126]  ( .D(\w0[4][126] ), .CLK(clk), .RST(rst), .Q(state[126]) );
  DFF \state_reg[102]  ( .D(\w0[4][102] ), .CLK(clk), .RST(rst), .Q(state[102]) );
  DFF \state_reg[119]  ( .D(\w0[4][119] ), .CLK(clk), .RST(rst), .Q(state[119]) );
  DFF \state_reg[111]  ( .D(\w0[4][111] ), .CLK(clk), .RST(rst), .Q(state[111]) );
  XOR U2988 ( .A(key[158]), .B(n3053), .Z(n2090) );
  XNOR U2989 ( .A(\w3[0][6] ), .B(n3186), .Z(n2091) );
  XNOR U2990 ( .A(n2090), .B(n2091), .Z(\w1[1][30] ) );
  XNOR U2991 ( .A(\w3[0][59] ), .B(\w3[0][35] ), .Z(n3086) );
  XNOR U2992 ( .A(\w3[0][91] ), .B(\w3[0][67] ), .Z(n3202) );
  XNOR U2993 ( .A(\w3[0][8] ), .B(\w3[0][12] ), .Z(n2092) );
  XNOR U2994 ( .A(n3048), .B(n2092), .Z(n3005) );
  XOR U2995 ( .A(n3139), .B(\w3[0][41] ), .Z(n2093) );
  XNOR U2996 ( .A(\w3[0][32] ), .B(key[168]), .Z(n2094) );
  XNOR U2997 ( .A(n2093), .B(n2094), .Z(n2095) );
  XOR U2998 ( .A(n3168), .B(n2095), .Z(\w1[1][40] ) );
  XOR U2999 ( .A(n3255), .B(\w3[0][73] ), .Z(n2096) );
  XNOR U3000 ( .A(\w3[0][64] ), .B(key[200]), .Z(n2097) );
  XNOR U3001 ( .A(n2096), .B(n2097), .Z(n2098) );
  XOR U3002 ( .A(n3282), .B(n2098), .Z(\w1[1][72] ) );
  XNOR U3003 ( .A(\w3[1][59] ), .B(\w3[1][35] ), .Z(n3502) );
  XOR U3004 ( .A(key[150]), .B(n3013), .Z(n2099) );
  XNOR U3005 ( .A(\w3[0][14] ), .B(n3053), .Z(n2100) );
  XOR U3006 ( .A(n2099), .B(n2100), .Z(\w1[1][22] ) );
  XOR U3007 ( .A(key[136]), .B(\w3[0][1] ), .Z(n2101) );
  XNOR U3008 ( .A(\w3[0][0] ), .B(n3256), .Z(n2102) );
  XNOR U3009 ( .A(n2101), .B(n2102), .Z(n2103) );
  XOR U3010 ( .A(n2103), .B(n3257), .Z(\w1[1][8] ) );
  XNOR U3011 ( .A(\w3[1][91] ), .B(\w3[1][67] ), .Z(n3618) );
  XOR U3012 ( .A(key[181]), .B(n3125), .Z(n2104) );
  XNOR U3013 ( .A(\w3[0][45] ), .B(n3124), .Z(n2105) );
  XOR U3014 ( .A(n2104), .B(n2105), .Z(\w1[1][53] ) );
  XOR U3015 ( .A(key[264]), .B(\w3[1][1] ), .Z(n2106) );
  XNOR U3016 ( .A(\w3[1][0] ), .B(n3672), .Z(n2107) );
  XNOR U3017 ( .A(n2106), .B(n2107), .Z(n2108) );
  XOR U3018 ( .A(n2108), .B(n3673), .Z(\w1[2][8] ) );
  XOR U3019 ( .A(n3554), .B(\w3[1][58] ), .Z(n2109) );
  XNOR U3020 ( .A(\w3[1][50] ), .B(key[313]), .Z(n2110) );
  XNOR U3021 ( .A(n2109), .B(n2110), .Z(n2111) );
  XOR U3022 ( .A(n3555), .B(n2111), .Z(\w1[2][57] ) );
  XNOR U3023 ( .A(\w3[2][59] ), .B(\w3[2][35] ), .Z(n3918) );
  XOR U3024 ( .A(n3671), .B(\w3[1][73] ), .Z(n2112) );
  XNOR U3025 ( .A(\w3[1][64] ), .B(key[328]), .Z(n2113) );
  XNOR U3026 ( .A(n2112), .B(n2113), .Z(n2114) );
  XOR U3027 ( .A(n3698), .B(n2114), .Z(\w1[2][72] ) );
  XNOR U3028 ( .A(\w3[2][91] ), .B(\w3[2][67] ), .Z(n4034) );
  XOR U3029 ( .A(key[277]), .B(n3430), .Z(n2115) );
  XNOR U3030 ( .A(\w3[1][13] ), .B(n3465), .Z(n2116) );
  XNOR U3031 ( .A(n2115), .B(n2116), .Z(\w1[2][21] ) );
  XOR U3032 ( .A(key[309]), .B(n3541), .Z(n2117) );
  XNOR U3033 ( .A(\w3[1][45] ), .B(n3540), .Z(n2118) );
  XOR U3034 ( .A(n2117), .B(n2118), .Z(\w1[2][53] ) );
  XOR U3035 ( .A(n3971), .B(\w3[2][41] ), .Z(n2119) );
  XNOR U3036 ( .A(\w3[2][32] ), .B(key[424]), .Z(n2120) );
  XNOR U3037 ( .A(n2119), .B(n2120), .Z(n2121) );
  XOR U3038 ( .A(n4000), .B(n2121), .Z(\w1[3][40] ) );
  XOR U3039 ( .A(n4087), .B(\w3[2][73] ), .Z(n2122) );
  XNOR U3040 ( .A(\w3[2][64] ), .B(key[456]), .Z(n2123) );
  XNOR U3041 ( .A(n2122), .B(n2123), .Z(n2124) );
  XOR U3042 ( .A(n4114), .B(n2124), .Z(\w1[3][72] ) );
  XOR U3043 ( .A(key[406]), .B(n3847), .Z(n2125) );
  XNOR U3044 ( .A(\w3[2][14] ), .B(n3882), .Z(n2126) );
  XOR U3045 ( .A(n2125), .B(n2126), .Z(\w1[3][22] ) );
  XOR U3046 ( .A(key[392]), .B(\w3[2][1] ), .Z(n2127) );
  XNOR U3047 ( .A(\w3[2][0] ), .B(n4088), .Z(n2128) );
  XNOR U3048 ( .A(n2127), .B(n2128), .Z(n2129) );
  XOR U3049 ( .A(n2129), .B(n4089), .Z(\w1[3][8] ) );
  XNOR U3050 ( .A(\w3[3][97] ), .B(\w3[3][105] ), .Z(n2250) );
  XNOR U3051 ( .A(\w3[3][107] ), .B(n2259), .Z(n2130) );
  XNOR U3052 ( .A(n2235), .B(n2130), .Z(\w0[4][115] ) );
  XOR U3053 ( .A(n2469), .B(\w3[3][7] ), .Z(n2131) );
  XNOR U3054 ( .A(n2443), .B(n2131), .Z(\w0[4][31] ) );
  XNOR U3055 ( .A(\w3[3][74] ), .B(n2449), .Z(n2132) );
  XNOR U3056 ( .A(n2448), .B(n2132), .Z(\w0[4][82] ) );
  XOR U3057 ( .A(key[147]), .B(n3005), .Z(n2133) );
  XNOR U3058 ( .A(\w3[0][11] ), .B(n3034), .Z(n2134) );
  XNOR U3059 ( .A(n2133), .B(n2134), .Z(\w1[1][19] ) );
  XOR U3060 ( .A(key[179]), .B(n3119), .Z(n2135) );
  XNOR U3061 ( .A(\w3[0][43] ), .B(n3146), .Z(n2136) );
  XNOR U3062 ( .A(n2135), .B(n2136), .Z(\w1[1][51] ) );
  XOR U3063 ( .A(key[211]), .B(n3235), .Z(n2137) );
  XNOR U3064 ( .A(\w3[0][75] ), .B(n3264), .Z(n2138) );
  XNOR U3065 ( .A(n2137), .B(n2138), .Z(\w1[1][83] ) );
  XNOR U3066 ( .A(\w3[1][8] ), .B(\w3[1][12] ), .Z(n2139) );
  XNOR U3067 ( .A(n3461), .B(n2139), .Z(n3421) );
  XOR U3068 ( .A(\w3[0][96] ), .B(n2962), .Z(n2140) );
  XNOR U3069 ( .A(key[232]), .B(\w3[0][105] ), .Z(n2141) );
  XNOR U3070 ( .A(n2140), .B(n2141), .Z(n2142) );
  XOR U3071 ( .A(n2142), .B(n3286), .Z(\w1[1][104] ) );
  XOR U3072 ( .A(n3138), .B(\w3[0][58] ), .Z(n2143) );
  XNOR U3073 ( .A(\w3[0][50] ), .B(key[185]), .Z(n2144) );
  XNOR U3074 ( .A(n2143), .B(n2144), .Z(n2145) );
  XOR U3075 ( .A(n3139), .B(n2145), .Z(\w1[1][57] ) );
  XOR U3076 ( .A(n3254), .B(\w3[0][90] ), .Z(n2146) );
  XNOR U3077 ( .A(\w3[0][82] ), .B(key[217]), .Z(n2147) );
  XNOR U3078 ( .A(n2146), .B(n2147), .Z(n2148) );
  XOR U3079 ( .A(n3255), .B(n2148), .Z(\w1[1][89] ) );
  XOR U3080 ( .A(key[307]), .B(n3535), .Z(n2149) );
  XNOR U3081 ( .A(\w3[1][43] ), .B(n3562), .Z(n2150) );
  XNOR U3082 ( .A(n2149), .B(n2150), .Z(\w1[2][51] ) );
  XOR U3083 ( .A(key[149]), .B(n3012), .Z(n2151) );
  XNOR U3084 ( .A(\w3[0][13] ), .B(n3052), .Z(n2152) );
  XNOR U3085 ( .A(n2151), .B(n2152), .Z(\w1[1][21] ) );
  XOR U3086 ( .A(key[339]), .B(n3651), .Z(n2153) );
  XNOR U3087 ( .A(\w3[1][75] ), .B(n3680), .Z(n2154) );
  XNOR U3088 ( .A(n2153), .B(n2154), .Z(\w1[2][83] ) );
  XOR U3089 ( .A(key[213]), .B(n3241), .Z(n2155) );
  XNOR U3090 ( .A(\w3[0][77] ), .B(n3240), .Z(n2156) );
  XNOR U3091 ( .A(n2155), .B(n2156), .Z(\w1[1][85] ) );
  XOR U3092 ( .A(\w3[1][1] ), .B(\w3[1][26] ), .Z(n2157) );
  XNOR U3093 ( .A(n3441), .B(key[281]), .Z(n2158) );
  XNOR U3094 ( .A(n2157), .B(n2158), .Z(n2159) );
  XNOR U3095 ( .A(n2159), .B(\w3[1][18] ), .Z(\w1[2][25] ) );
  XOR U3096 ( .A(key[278]), .B(n3431), .Z(n2160) );
  XNOR U3097 ( .A(\w3[1][14] ), .B(n3466), .Z(n2161) );
  XOR U3098 ( .A(n2160), .B(n2161), .Z(\w1[2][22] ) );
  XOR U3099 ( .A(n3555), .B(\w3[1][41] ), .Z(n2162) );
  XNOR U3100 ( .A(\w3[1][32] ), .B(key[296]), .Z(n2163) );
  XNOR U3101 ( .A(n2162), .B(n2163), .Z(n2164) );
  XOR U3102 ( .A(n3584), .B(n2164), .Z(\w1[2][40] ) );
  XNOR U3103 ( .A(\w3[2][8] ), .B(\w3[2][12] ), .Z(n2165) );
  XNOR U3104 ( .A(n3877), .B(n2165), .Z(n3837) );
  XOR U3105 ( .A(n3670), .B(\w3[1][90] ), .Z(n2166) );
  XNOR U3106 ( .A(\w3[1][82] ), .B(key[345]), .Z(n2167) );
  XNOR U3107 ( .A(n2166), .B(n2167), .Z(n2168) );
  XOR U3108 ( .A(n3671), .B(n2168), .Z(\w1[2][89] ) );
  XOR U3109 ( .A(\w3[1][96] ), .B(n3377), .Z(n2169) );
  XNOR U3110 ( .A(key[360]), .B(\w3[1][105] ), .Z(n2170) );
  XNOR U3111 ( .A(n2169), .B(n2170), .Z(n2171) );
  XOR U3112 ( .A(n2171), .B(n3702), .Z(\w1[2][104] ) );
  XOR U3113 ( .A(key[467]), .B(n4067), .Z(n2172) );
  XNOR U3114 ( .A(\w3[2][75] ), .B(n4096), .Z(n2173) );
  XNOR U3115 ( .A(n2172), .B(n2173), .Z(\w1[3][83] ) );
  XOR U3116 ( .A(key[341]), .B(n3657), .Z(n2174) );
  XNOR U3117 ( .A(\w3[1][77] ), .B(n3656), .Z(n2175) );
  XOR U3118 ( .A(n2174), .B(n2175), .Z(\w1[2][85] ) );
  XOR U3119 ( .A(key[435]), .B(n3951), .Z(n2176) );
  XNOR U3120 ( .A(\w3[2][43] ), .B(n3978), .Z(n2177) );
  XNOR U3121 ( .A(n2176), .B(n2177), .Z(\w1[3][51] ) );
  XOR U3122 ( .A(\w3[2][1] ), .B(\w3[2][26] ), .Z(n2178) );
  XNOR U3123 ( .A(n3857), .B(key[409]), .Z(n2179) );
  XNOR U3124 ( .A(n2178), .B(n2179), .Z(n2180) );
  XNOR U3125 ( .A(n2180), .B(\w3[2][18] ), .Z(\w1[3][25] ) );
  XOR U3126 ( .A(\w3[2][96] ), .B(n3794), .Z(n2181) );
  XNOR U3127 ( .A(key[488]), .B(\w3[2][105] ), .Z(n2182) );
  XNOR U3128 ( .A(n2181), .B(n2182), .Z(n2183) );
  XOR U3129 ( .A(n2183), .B(n4118), .Z(\w1[3][104] ) );
  XOR U3130 ( .A(n3970), .B(\w3[2][58] ), .Z(n2184) );
  XNOR U3131 ( .A(\w3[2][50] ), .B(key[441]), .Z(n2185) );
  XNOR U3132 ( .A(n2184), .B(n2185), .Z(n2186) );
  XOR U3133 ( .A(n3971), .B(n2186), .Z(\w1[3][57] ) );
  XOR U3134 ( .A(n4086), .B(\w3[2][90] ), .Z(n2187) );
  XNOR U3135 ( .A(\w3[2][82] ), .B(key[473]), .Z(n2188) );
  XNOR U3136 ( .A(n2187), .B(n2188), .Z(n2189) );
  XOR U3137 ( .A(n4087), .B(n2189), .Z(\w1[3][89] ) );
  XOR U3138 ( .A(key[469]), .B(n4073), .Z(n2190) );
  XNOR U3139 ( .A(\w3[2][77] ), .B(n4072), .Z(n2191) );
  XOR U3140 ( .A(n2190), .B(n2191), .Z(\w1[3][85] ) );
  XOR U3141 ( .A(key[405]), .B(n3846), .Z(n2192) );
  XNOR U3142 ( .A(\w3[2][13] ), .B(n3881), .Z(n2193) );
  XNOR U3143 ( .A(n2192), .B(n2193), .Z(\w1[3][21] ) );
  XOR U3144 ( .A(key[437]), .B(n3957), .Z(n2194) );
  XNOR U3145 ( .A(\w3[2][45] ), .B(n3956), .Z(n2195) );
  XOR U3146 ( .A(n2194), .B(n2195), .Z(\w1[3][53] ) );
  XNOR U3147 ( .A(\w3[3][96] ), .B(n2250), .Z(n2196) );
  XNOR U3148 ( .A(n2489), .B(n2196), .Z(\w0[4][104] ) );
  XNOR U3149 ( .A(\w3[3][13] ), .B(n2319), .Z(n2197) );
  XNOR U3150 ( .A(n2290), .B(n2197), .Z(\w0[4][21] ) );
  XOR U3151 ( .A(n2469), .B(n2468), .Z(n2198) );
  XNOR U3152 ( .A(\w3[3][0] ), .B(\w3[3][1] ), .Z(n2199) );
  XOR U3153 ( .A(n2198), .B(n2199), .Z(\w0[4][8] ) );
  XOR U3154 ( .A(\w3[3][45] ), .B(n2371), .Z(n2200) );
  XNOR U3155 ( .A(n2372), .B(n2200), .Z(\w0[4][53] ) );
  XOR U3156 ( .A(\w3[3][41] ), .B(n2386), .Z(n2201) );
  XNOR U3157 ( .A(n2359), .B(n2201), .Z(\w0[4][49] ) );
  XOR U3158 ( .A(\w3[3][73] ), .B(n2470), .Z(n2202) );
  XNOR U3159 ( .A(n2447), .B(n2202), .Z(\w0[4][81] ) );
  IV U3160 ( .A(init), .Z(n2203) );
  XOR U3161 ( .A(key[512]), .B(\w3[4][0] ), .Z(out[0]) );
  XOR U3162 ( .A(key[612]), .B(\w3[4][100] ), .Z(out[100]) );
  XOR U3163 ( .A(key[613]), .B(\w3[4][101] ), .Z(out[101]) );
  XOR U3164 ( .A(key[614]), .B(\w3[4][102] ), .Z(out[102]) );
  XOR U3165 ( .A(key[615]), .B(\w3[4][103] ), .Z(out[103]) );
  XOR U3166 ( .A(key[616]), .B(\w3[4][104] ), .Z(out[104]) );
  XOR U3167 ( .A(key[617]), .B(\w3[4][105] ), .Z(out[105]) );
  XOR U3168 ( .A(key[618]), .B(\w3[4][106] ), .Z(out[106]) );
  XOR U3169 ( .A(key[619]), .B(\w3[4][107] ), .Z(out[107]) );
  XOR U3170 ( .A(key[620]), .B(\w3[4][108] ), .Z(out[108]) );
  XOR U3171 ( .A(key[621]), .B(\w3[4][109] ), .Z(out[109]) );
  XOR U3172 ( .A(key[522]), .B(\w3[4][10] ), .Z(out[10]) );
  XOR U3173 ( .A(key[622]), .B(\w3[4][110] ), .Z(out[110]) );
  XOR U3174 ( .A(key[623]), .B(\w3[4][111] ), .Z(out[111]) );
  XOR U3175 ( .A(key[624]), .B(\w3[4][112] ), .Z(out[112]) );
  XOR U3176 ( .A(key[625]), .B(\w3[4][113] ), .Z(out[113]) );
  XOR U3177 ( .A(key[626]), .B(\w3[4][114] ), .Z(out[114]) );
  XOR U3178 ( .A(key[627]), .B(\w3[4][115] ), .Z(out[115]) );
  XOR U3179 ( .A(key[628]), .B(\w3[4][116] ), .Z(out[116]) );
  XOR U3180 ( .A(key[629]), .B(\w3[4][117] ), .Z(out[117]) );
  XOR U3181 ( .A(key[630]), .B(\w3[4][118] ), .Z(out[118]) );
  XOR U3182 ( .A(key[631]), .B(\w3[4][119] ), .Z(out[119]) );
  XOR U3183 ( .A(key[523]), .B(\w3[4][11] ), .Z(out[11]) );
  XOR U3184 ( .A(key[632]), .B(\w3[4][120] ), .Z(out[120]) );
  XOR U3185 ( .A(key[633]), .B(\w3[4][121] ), .Z(out[121]) );
  XOR U3186 ( .A(key[634]), .B(\w3[4][122] ), .Z(out[122]) );
  XOR U3187 ( .A(key[635]), .B(\w3[4][123] ), .Z(out[123]) );
  XOR U3188 ( .A(key[636]), .B(\w3[4][124] ), .Z(out[124]) );
  XOR U3189 ( .A(key[637]), .B(\w3[4][125] ), .Z(out[125]) );
  XOR U3190 ( .A(key[638]), .B(\w3[4][126] ), .Z(out[126]) );
  XOR U3191 ( .A(key[639]), .B(\w3[4][127] ), .Z(out[127]) );
  XOR U3192 ( .A(key[524]), .B(\w3[4][12] ), .Z(out[12]) );
  XOR U3193 ( .A(key[525]), .B(\w3[4][13] ), .Z(out[13]) );
  XOR U3194 ( .A(key[526]), .B(\w3[4][14] ), .Z(out[14]) );
  XOR U3195 ( .A(key[527]), .B(\w3[4][15] ), .Z(out[15]) );
  XOR U3196 ( .A(key[528]), .B(\w3[4][16] ), .Z(out[16]) );
  XOR U3197 ( .A(key[529]), .B(\w3[4][17] ), .Z(out[17]) );
  XOR U3198 ( .A(key[530]), .B(\w3[4][18] ), .Z(out[18]) );
  XOR U3199 ( .A(key[531]), .B(\w3[4][19] ), .Z(out[19]) );
  XOR U3200 ( .A(key[513]), .B(\w3[4][1] ), .Z(out[1]) );
  XOR U3201 ( .A(key[532]), .B(\w3[4][20] ), .Z(out[20]) );
  XOR U3202 ( .A(key[533]), .B(\w3[4][21] ), .Z(out[21]) );
  XOR U3203 ( .A(key[534]), .B(\w3[4][22] ), .Z(out[22]) );
  XOR U3204 ( .A(key[535]), .B(\w3[4][23] ), .Z(out[23]) );
  XOR U3205 ( .A(key[536]), .B(\w3[4][24] ), .Z(out[24]) );
  XOR U3206 ( .A(key[537]), .B(\w3[4][25] ), .Z(out[25]) );
  XOR U3207 ( .A(key[538]), .B(\w3[4][26] ), .Z(out[26]) );
  XOR U3208 ( .A(key[539]), .B(\w3[4][27] ), .Z(out[27]) );
  XOR U3209 ( .A(key[540]), .B(\w3[4][28] ), .Z(out[28]) );
  XOR U3210 ( .A(key[541]), .B(\w3[4][29] ), .Z(out[29]) );
  XOR U3211 ( .A(key[514]), .B(\w3[4][2] ), .Z(out[2]) );
  XOR U3212 ( .A(key[542]), .B(\w3[4][30] ), .Z(out[30]) );
  XOR U3213 ( .A(key[543]), .B(\w3[4][31] ), .Z(out[31]) );
  XOR U3214 ( .A(key[544]), .B(\w3[4][32] ), .Z(out[32]) );
  XOR U3215 ( .A(key[545]), .B(\w3[4][33] ), .Z(out[33]) );
  XOR U3216 ( .A(key[546]), .B(\w3[4][34] ), .Z(out[34]) );
  XOR U3217 ( .A(key[547]), .B(\w3[4][35] ), .Z(out[35]) );
  XOR U3218 ( .A(key[548]), .B(\w3[4][36] ), .Z(out[36]) );
  XOR U3219 ( .A(key[549]), .B(\w3[4][37] ), .Z(out[37]) );
  XOR U3220 ( .A(key[550]), .B(\w3[4][38] ), .Z(out[38]) );
  XOR U3221 ( .A(key[551]), .B(\w3[4][39] ), .Z(out[39]) );
  XOR U3222 ( .A(key[515]), .B(\w3[4][3] ), .Z(out[3]) );
  XOR U3223 ( .A(key[552]), .B(\w3[4][40] ), .Z(out[40]) );
  XOR U3224 ( .A(key[553]), .B(\w3[4][41] ), .Z(out[41]) );
  XOR U3225 ( .A(key[554]), .B(\w3[4][42] ), .Z(out[42]) );
  XOR U3226 ( .A(key[555]), .B(\w3[4][43] ), .Z(out[43]) );
  XOR U3227 ( .A(key[556]), .B(\w3[4][44] ), .Z(out[44]) );
  XOR U3228 ( .A(key[557]), .B(\w3[4][45] ), .Z(out[45]) );
  XOR U3229 ( .A(key[558]), .B(\w3[4][46] ), .Z(out[46]) );
  XOR U3230 ( .A(key[559]), .B(\w3[4][47] ), .Z(out[47]) );
  XOR U3231 ( .A(key[560]), .B(\w3[4][48] ), .Z(out[48]) );
  XOR U3232 ( .A(key[561]), .B(\w3[4][49] ), .Z(out[49]) );
  XOR U3233 ( .A(key[516]), .B(\w3[4][4] ), .Z(out[4]) );
  XOR U3234 ( .A(key[562]), .B(\w3[4][50] ), .Z(out[50]) );
  XOR U3235 ( .A(key[563]), .B(\w3[4][51] ), .Z(out[51]) );
  XOR U3236 ( .A(key[564]), .B(\w3[4][52] ), .Z(out[52]) );
  XOR U3237 ( .A(key[565]), .B(\w3[4][53] ), .Z(out[53]) );
  XOR U3238 ( .A(key[566]), .B(\w3[4][54] ), .Z(out[54]) );
  XOR U3239 ( .A(key[567]), .B(\w3[4][55] ), .Z(out[55]) );
  XOR U3240 ( .A(key[568]), .B(\w3[4][56] ), .Z(out[56]) );
  XOR U3241 ( .A(key[569]), .B(\w3[4][57] ), .Z(out[57]) );
  XOR U3242 ( .A(key[570]), .B(\w3[4][58] ), .Z(out[58]) );
  XOR U3243 ( .A(key[571]), .B(\w3[4][59] ), .Z(out[59]) );
  XOR U3244 ( .A(key[517]), .B(\w3[4][5] ), .Z(out[5]) );
  XOR U3245 ( .A(key[572]), .B(\w3[4][60] ), .Z(out[60]) );
  XOR U3246 ( .A(key[573]), .B(\w3[4][61] ), .Z(out[61]) );
  XOR U3247 ( .A(key[574]), .B(\w3[4][62] ), .Z(out[62]) );
  XOR U3248 ( .A(key[575]), .B(\w3[4][63] ), .Z(out[63]) );
  XOR U3249 ( .A(key[576]), .B(\w3[4][64] ), .Z(out[64]) );
  XOR U3250 ( .A(key[577]), .B(\w3[4][65] ), .Z(out[65]) );
  XOR U3251 ( .A(key[578]), .B(\w3[4][66] ), .Z(out[66]) );
  XOR U3252 ( .A(key[579]), .B(\w3[4][67] ), .Z(out[67]) );
  XOR U3253 ( .A(key[580]), .B(\w3[4][68] ), .Z(out[68]) );
  XOR U3254 ( .A(key[581]), .B(\w3[4][69] ), .Z(out[69]) );
  XOR U3255 ( .A(key[518]), .B(\w3[4][6] ), .Z(out[6]) );
  XOR U3256 ( .A(key[582]), .B(\w3[4][70] ), .Z(out[70]) );
  XOR U3257 ( .A(key[583]), .B(\w3[4][71] ), .Z(out[71]) );
  XOR U3258 ( .A(key[584]), .B(\w3[4][72] ), .Z(out[72]) );
  XOR U3259 ( .A(key[585]), .B(\w3[4][73] ), .Z(out[73]) );
  XOR U3260 ( .A(key[586]), .B(\w3[4][74] ), .Z(out[74]) );
  XOR U3261 ( .A(key[587]), .B(\w3[4][75] ), .Z(out[75]) );
  XOR U3262 ( .A(key[588]), .B(\w3[4][76] ), .Z(out[76]) );
  XOR U3263 ( .A(key[589]), .B(\w3[4][77] ), .Z(out[77]) );
  XOR U3264 ( .A(key[590]), .B(\w3[4][78] ), .Z(out[78]) );
  XOR U3265 ( .A(key[591]), .B(\w3[4][79] ), .Z(out[79]) );
  XOR U3266 ( .A(key[519]), .B(\w3[4][7] ), .Z(out[7]) );
  XOR U3267 ( .A(key[592]), .B(\w3[4][80] ), .Z(out[80]) );
  XOR U3268 ( .A(key[593]), .B(\w3[4][81] ), .Z(out[81]) );
  XOR U3269 ( .A(key[594]), .B(\w3[4][82] ), .Z(out[82]) );
  XOR U3270 ( .A(key[595]), .B(\w3[4][83] ), .Z(out[83]) );
  XOR U3271 ( .A(key[596]), .B(\w3[4][84] ), .Z(out[84]) );
  XOR U3272 ( .A(key[597]), .B(\w3[4][85] ), .Z(out[85]) );
  XOR U3273 ( .A(key[598]), .B(\w3[4][86] ), .Z(out[86]) );
  XOR U3274 ( .A(key[599]), .B(\w3[4][87] ), .Z(out[87]) );
  XOR U3275 ( .A(key[600]), .B(\w3[4][88] ), .Z(out[88]) );
  XOR U3276 ( .A(key[601]), .B(\w3[4][89] ), .Z(out[89]) );
  XOR U3277 ( .A(key[520]), .B(\w3[4][8] ), .Z(out[8]) );
  XOR U3278 ( .A(key[602]), .B(\w3[4][90] ), .Z(out[90]) );
  XOR U3279 ( .A(key[603]), .B(\w3[4][91] ), .Z(out[91]) );
  XOR U3280 ( .A(key[604]), .B(\w3[4][92] ), .Z(out[92]) );
  XOR U3281 ( .A(key[605]), .B(\w3[4][93] ), .Z(out[93]) );
  XOR U3282 ( .A(key[606]), .B(\w3[4][94] ), .Z(out[94]) );
  XOR U3283 ( .A(key[607]), .B(\w3[4][95] ), .Z(out[95]) );
  XOR U3284 ( .A(key[608]), .B(\w3[4][96] ), .Z(out[96]) );
  XOR U3285 ( .A(key[609]), .B(\w3[4][97] ), .Z(out[97]) );
  XOR U3286 ( .A(key[610]), .B(\w3[4][98] ), .Z(out[98]) );
  XOR U3287 ( .A(key[611]), .B(\w3[4][99] ), .Z(out[99]) );
  XOR U3288 ( .A(key[521]), .B(\w3[4][9] ), .Z(out[9]) );
  XNOR U3289 ( .A(\w3[3][1] ), .B(\w3[3][25] ), .Z(n2503) );
  XOR U3290 ( .A(\w3[3][16] ), .B(\w3[3][24] ), .Z(n2469) );
  XOR U3291 ( .A(n2503), .B(n2469), .Z(n2204) );
  XNOR U3292 ( .A(\w3[3][8] ), .B(n2204), .Z(\w0[4][0] ) );
  XOR U3293 ( .A(\w3[3][96] ), .B(\w3[3][101] ), .Z(n2219) );
  XOR U3294 ( .A(\w3[3][108] ), .B(\w3[3][116] ), .Z(n2206) );
  IV U3295 ( .A(\w3[3][120] ), .Z(n2256) );
  XOR U3296 ( .A(n2256), .B(\w3[3][125] ), .Z(n2205) );
  XOR U3297 ( .A(n2206), .B(n2205), .Z(n2263) );
  XOR U3298 ( .A(\w3[3][124] ), .B(n2263), .Z(n2207) );
  XNOR U3299 ( .A(n2219), .B(n2207), .Z(\w0[4][100] ) );
  XNOR U3300 ( .A(\w3[3][102] ), .B(\w3[3][126] ), .Z(n2225) );
  XNOR U3301 ( .A(\w3[3][109] ), .B(\w3[3][117] ), .Z(n2266) );
  XOR U3302 ( .A(\w3[3][125] ), .B(n2266), .Z(n2208) );
  XOR U3303 ( .A(n2225), .B(n2208), .Z(\w0[4][101] ) );
  XOR U3304 ( .A(\w3[3][96] ), .B(\w3[3][103] ), .Z(n2226) );
  XOR U3305 ( .A(n2256), .B(\w3[3][127] ), .Z(n2210) );
  XOR U3306 ( .A(\w3[3][110] ), .B(\w3[3][118] ), .Z(n2240) );
  XOR U3307 ( .A(n2210), .B(n2240), .Z(n2269) );
  XOR U3308 ( .A(\w3[3][126] ), .B(n2269), .Z(n2209) );
  XNOR U3309 ( .A(n2226), .B(n2209), .Z(\w0[4][102] ) );
  XNOR U3310 ( .A(\w3[3][111] ), .B(\w3[3][119] ), .Z(n2272) );
  XOR U3311 ( .A(\w3[3][96] ), .B(n2210), .Z(n2211) );
  XOR U3312 ( .A(n2272), .B(n2211), .Z(\w0[4][103] ) );
  XNOR U3313 ( .A(\w3[3][120] ), .B(\w3[3][112] ), .Z(n2489) );
  XOR U3314 ( .A(\w3[3][106] ), .B(\w3[3][98] ), .Z(n2253) );
  XNOR U3315 ( .A(\w3[3][113] ), .B(\w3[3][121] ), .Z(n2492) );
  XOR U3316 ( .A(\w3[3][97] ), .B(n2492), .Z(n2212) );
  XNOR U3317 ( .A(n2253), .B(n2212), .Z(\w0[4][105] ) );
  XOR U3318 ( .A(\w3[3][98] ), .B(\w3[3][122] ), .Z(n2494) );
  XOR U3319 ( .A(\w3[3][114] ), .B(n2494), .Z(n2214) );
  IV U3320 ( .A(\w3[3][99] ), .Z(n2260) );
  XOR U3321 ( .A(\w3[3][107] ), .B(n2260), .Z(n2213) );
  XNOR U3322 ( .A(n2214), .B(n2213), .Z(\w0[4][106] ) );
  IV U3323 ( .A(\w3[3][123] ), .Z(n2499) );
  XOR U3324 ( .A(\w3[3][99] ), .B(n2499), .Z(n2495) );
  XOR U3325 ( .A(\w3[3][108] ), .B(n2495), .Z(n2215) );
  XOR U3326 ( .A(\w3[3][104] ), .B(n2215), .Z(n2235) );
  IV U3327 ( .A(\w3[3][100] ), .Z(n2262) );
  XOR U3328 ( .A(\w3[3][96] ), .B(n2262), .Z(n2500) );
  XOR U3329 ( .A(\w3[3][115] ), .B(n2500), .Z(n2216) );
  XOR U3330 ( .A(n2235), .B(n2216), .Z(\w0[4][107] ) );
  XOR U3331 ( .A(\w3[3][100] ), .B(\w3[3][104] ), .Z(n2218) );
  XNOR U3332 ( .A(\w3[3][124] ), .B(\w3[3][109] ), .Z(n2217) );
  XOR U3333 ( .A(n2218), .B(n2217), .Z(n2236) );
  XNOR U3334 ( .A(\w3[3][116] ), .B(n2219), .Z(n2220) );
  XOR U3335 ( .A(n2236), .B(n2220), .Z(\w0[4][108] ) );
  XNOR U3336 ( .A(\w3[3][125] ), .B(\w3[3][101] ), .Z(n2238) );
  XNOR U3337 ( .A(\w3[3][110] ), .B(n2238), .Z(n2222) );
  XNOR U3338 ( .A(\w3[3][117] ), .B(\w3[3][102] ), .Z(n2221) );
  XNOR U3339 ( .A(n2222), .B(n2221), .Z(\w0[4][109] ) );
  XNOR U3340 ( .A(\w3[3][2] ), .B(\w3[3][26] ), .Z(n2286) );
  XNOR U3341 ( .A(\w3[3][3] ), .B(n2286), .Z(n2224) );
  XNOR U3342 ( .A(\w3[3][11] ), .B(\w3[3][18] ), .Z(n2223) );
  XNOR U3343 ( .A(n2224), .B(n2223), .Z(\w0[4][10] ) );
  XOR U3344 ( .A(\w3[3][111] ), .B(\w3[3][104] ), .Z(n2245) );
  XOR U3345 ( .A(n2225), .B(n2245), .Z(n2241) );
  XNOR U3346 ( .A(\w3[3][118] ), .B(n2226), .Z(n2227) );
  XOR U3347 ( .A(n2241), .B(n2227), .Z(\w0[4][110] ) );
  XOR U3348 ( .A(\w3[3][127] ), .B(\w3[3][103] ), .Z(n2243) );
  XNOR U3349 ( .A(\w3[3][96] ), .B(\w3[3][104] ), .Z(n2249) );
  XOR U3350 ( .A(\w3[3][119] ), .B(n2249), .Z(n2228) );
  XNOR U3351 ( .A(n2243), .B(n2228), .Z(\w0[4][111] ) );
  XNOR U3352 ( .A(\w3[3][113] ), .B(n2249), .Z(n2230) );
  IV U3353 ( .A(\w3[3][105] ), .Z(n2231) );
  XOR U3354 ( .A(\w3[3][120] ), .B(n2231), .Z(n2229) );
  XNOR U3355 ( .A(n2230), .B(n2229), .Z(\w0[4][112] ) );
  XOR U3356 ( .A(\w3[3][97] ), .B(\w3[3][121] ), .Z(n2491) );
  XOR U3357 ( .A(\w3[3][114] ), .B(n2491), .Z(n2233) );
  IV U3358 ( .A(\w3[3][106] ), .Z(n2496) );
  XNOR U3359 ( .A(n2231), .B(n2496), .Z(n2232) );
  XNOR U3360 ( .A(n2233), .B(n2232), .Z(\w0[4][113] ) );
  IV U3361 ( .A(\w3[3][115] ), .Z(n2252) );
  XOR U3362 ( .A(\w3[3][107] ), .B(n2252), .Z(n2258) );
  XOR U3363 ( .A(n2496), .B(n2494), .Z(n2234) );
  XOR U3364 ( .A(n2258), .B(n2234), .Z(\w0[4][114] ) );
  XNOR U3365 ( .A(\w3[3][116] ), .B(\w3[3][112] ), .Z(n2259) );
  XNOR U3366 ( .A(\w3[3][117] ), .B(\w3[3][112] ), .Z(n2265) );
  XOR U3367 ( .A(\w3[3][108] ), .B(n2236), .Z(n2237) );
  XOR U3368 ( .A(n2265), .B(n2237), .Z(\w0[4][116] ) );
  XNOR U3369 ( .A(\w3[3][109] ), .B(n2238), .Z(n2239) );
  XOR U3370 ( .A(n2240), .B(n2239), .Z(\w0[4][117] ) );
  XNOR U3371 ( .A(\w3[3][119] ), .B(\w3[3][112] ), .Z(n2271) );
  XOR U3372 ( .A(\w3[3][110] ), .B(n2241), .Z(n2242) );
  XOR U3373 ( .A(n2271), .B(n2242), .Z(\w0[4][118] ) );
  XOR U3374 ( .A(\w3[3][112] ), .B(n2243), .Z(n2244) );
  XOR U3375 ( .A(n2245), .B(n2244), .Z(\w0[4][119] ) );
  XNOR U3376 ( .A(\w3[3][3] ), .B(\w3[3][27] ), .Z(n2315) );
  XNOR U3377 ( .A(\w3[3][8] ), .B(\w3[3][12] ), .Z(n2246) );
  XNOR U3378 ( .A(n2315), .B(n2246), .Z(n2284) );
  XNOR U3379 ( .A(\w3[3][0] ), .B(\w3[3][4] ), .Z(n2334) );
  XOR U3380 ( .A(\w3[3][19] ), .B(n2334), .Z(n2247) );
  XOR U3381 ( .A(n2284), .B(n2247), .Z(\w0[4][11] ) );
  XOR U3382 ( .A(\w3[3][112] ), .B(n2492), .Z(n2248) );
  XOR U3383 ( .A(n2249), .B(n2248), .Z(\w0[4][120] ) );
  XNOR U3384 ( .A(\w3[3][114] ), .B(\w3[3][122] ), .Z(n2498) );
  XOR U3385 ( .A(n2250), .B(\w3[3][113] ), .Z(n2251) );
  XOR U3386 ( .A(n2498), .B(n2251), .Z(\w0[4][121] ) );
  XOR U3387 ( .A(n2252), .B(n2499), .Z(n2255) );
  XNOR U3388 ( .A(n2253), .B(\w3[3][114] ), .Z(n2254) );
  XNOR U3389 ( .A(n2255), .B(n2254), .Z(\w0[4][122] ) );
  XOR U3390 ( .A(\w3[3][124] ), .B(n2256), .Z(n2257) );
  XOR U3391 ( .A(n2258), .B(n2257), .Z(n2502) );
  XNOR U3392 ( .A(n2260), .B(n2259), .Z(n2261) );
  XNOR U3393 ( .A(n2502), .B(n2261), .Z(\w0[4][123] ) );
  XNOR U3394 ( .A(n2263), .B(n2262), .Z(n2264) );
  XOR U3395 ( .A(n2265), .B(n2264), .Z(\w0[4][124] ) );
  XOR U3396 ( .A(\w3[3][126] ), .B(\w3[3][118] ), .Z(n2268) );
  XOR U3397 ( .A(\w3[3][101] ), .B(n2266), .Z(n2267) );
  XNOR U3398 ( .A(n2268), .B(n2267), .Z(\w0[4][125] ) );
  XOR U3399 ( .A(\w3[3][102] ), .B(n2269), .Z(n2270) );
  XOR U3400 ( .A(n2271), .B(n2270), .Z(\w0[4][126] ) );
  XOR U3401 ( .A(\w3[3][103] ), .B(n2272), .Z(n2273) );
  XOR U3402 ( .A(n2489), .B(n2273), .Z(\w0[4][127] ) );
  XOR U3403 ( .A(\w3[3][13] ), .B(\w3[3][28] ), .Z(n2275) );
  XNOR U3404 ( .A(\w3[3][8] ), .B(\w3[3][4] ), .Z(n2274) );
  XOR U3405 ( .A(n2275), .B(n2274), .Z(n2288) );
  XNOR U3406 ( .A(\w3[3][0] ), .B(\w3[3][5] ), .Z(n2360) );
  XOR U3407 ( .A(\w3[3][20] ), .B(n2360), .Z(n2276) );
  XOR U3408 ( .A(n2288), .B(n2276), .Z(\w0[4][12] ) );
  XNOR U3409 ( .A(\w3[3][5] ), .B(\w3[3][29] ), .Z(n2290) );
  XNOR U3410 ( .A(\w3[3][21] ), .B(n2290), .Z(n2278) );
  XNOR U3411 ( .A(\w3[3][14] ), .B(\w3[3][6] ), .Z(n2277) );
  XNOR U3412 ( .A(n2278), .B(n2277), .Z(\w0[4][13] ) );
  XNOR U3413 ( .A(\w3[3][6] ), .B(\w3[3][30] ), .Z(n2392) );
  XOR U3414 ( .A(\w3[3][8] ), .B(\w3[3][15] ), .Z(n2295) );
  XOR U3415 ( .A(n2392), .B(n2295), .Z(n2291) );
  XNOR U3416 ( .A(\w3[3][0] ), .B(\w3[3][7] ), .Z(n2416) );
  XOR U3417 ( .A(\w3[3][22] ), .B(n2416), .Z(n2279) );
  XOR U3418 ( .A(n2291), .B(n2279), .Z(\w0[4][14] ) );
  XNOR U3419 ( .A(\w3[3][7] ), .B(\w3[3][31] ), .Z(n2293) );
  XOR U3420 ( .A(\w3[3][8] ), .B(\w3[3][0] ), .Z(n2296) );
  XNOR U3421 ( .A(\w3[3][23] ), .B(n2296), .Z(n2280) );
  XOR U3422 ( .A(n2293), .B(n2280), .Z(\w0[4][15] ) );
  XOR U3423 ( .A(\w3[3][17] ), .B(\w3[3][9] ), .Z(n2299) );
  XNOR U3424 ( .A(\w3[3][24] ), .B(n2296), .Z(n2281) );
  XNOR U3425 ( .A(n2299), .B(n2281), .Z(\w0[4][16] ) );
  XOR U3426 ( .A(\w3[3][18] ), .B(\w3[3][10] ), .Z(n2317) );
  IV U3427 ( .A(\w3[3][9] ), .Z(n2468) );
  XNOR U3428 ( .A(n2503), .B(n2468), .Z(n2282) );
  XNOR U3429 ( .A(n2317), .B(n2282), .Z(\w0[4][17] ) );
  XNOR U3430 ( .A(\w3[3][11] ), .B(\w3[3][19] ), .Z(n2305) );
  XOR U3431 ( .A(n2286), .B(\w3[3][10] ), .Z(n2283) );
  XOR U3432 ( .A(n2305), .B(n2283), .Z(\w0[4][18] ) );
  XNOR U3433 ( .A(\w3[3][16] ), .B(\w3[3][20] ), .Z(n2306) );
  XOR U3434 ( .A(\w3[3][11] ), .B(n2284), .Z(n2285) );
  XOR U3435 ( .A(n2306), .B(n2285), .Z(\w0[4][19] ) );
  XOR U3436 ( .A(\w3[3][25] ), .B(n2286), .Z(n2287) );
  XNOR U3437 ( .A(n2299), .B(n2287), .Z(\w0[4][1] ) );
  IV U3438 ( .A(\w3[3][21] ), .Z(n2312) );
  XOR U3439 ( .A(\w3[3][16] ), .B(n2312), .Z(n2310) );
  XOR U3440 ( .A(\w3[3][12] ), .B(n2288), .Z(n2289) );
  XOR U3441 ( .A(n2310), .B(n2289), .Z(\w0[4][20] ) );
  XNOR U3442 ( .A(\w3[3][14] ), .B(\w3[3][22] ), .Z(n2319) );
  XNOR U3443 ( .A(\w3[3][16] ), .B(\w3[3][23] ), .Z(n2320) );
  XOR U3444 ( .A(\w3[3][14] ), .B(n2291), .Z(n2292) );
  XOR U3445 ( .A(n2320), .B(n2292), .Z(\w0[4][22] ) );
  XNOR U3446 ( .A(\w3[3][16] ), .B(n2293), .Z(n2294) );
  XOR U3447 ( .A(n2295), .B(n2294), .Z(\w0[4][23] ) );
  XOR U3448 ( .A(n2296), .B(\w3[3][17] ), .Z(n2298) );
  XNOR U3449 ( .A(\w3[3][25] ), .B(\w3[3][16] ), .Z(n2297) );
  XNOR U3450 ( .A(n2298), .B(n2297), .Z(\w0[4][24] ) );
  XOR U3451 ( .A(\w3[3][26] ), .B(n2299), .Z(n2301) );
  XNOR U3452 ( .A(\w3[3][1] ), .B(\w3[3][18] ), .Z(n2300) );
  XNOR U3453 ( .A(n2301), .B(n2300), .Z(\w0[4][25] ) );
  XOR U3454 ( .A(\w3[3][27] ), .B(n2317), .Z(n2303) );
  XNOR U3455 ( .A(\w3[3][2] ), .B(\w3[3][19] ), .Z(n2302) );
  XNOR U3456 ( .A(n2303), .B(n2302), .Z(\w0[4][26] ) );
  IV U3457 ( .A(\w3[3][24] ), .Z(n2318) );
  XOR U3458 ( .A(n2318), .B(\w3[3][28] ), .Z(n2304) );
  XOR U3459 ( .A(n2305), .B(n2304), .Z(n2336) );
  XOR U3460 ( .A(\w3[3][3] ), .B(n2306), .Z(n2307) );
  XNOR U3461 ( .A(n2336), .B(n2307), .Z(\w0[4][27] ) );
  XOR U3462 ( .A(\w3[3][20] ), .B(\w3[3][29] ), .Z(n2309) );
  XOR U3463 ( .A(n2318), .B(\w3[3][12] ), .Z(n2308) );
  XOR U3464 ( .A(n2309), .B(n2308), .Z(n2362) );
  XOR U3465 ( .A(\w3[3][4] ), .B(n2310), .Z(n2311) );
  XOR U3466 ( .A(n2362), .B(n2311), .Z(\w0[4][28] ) );
  XOR U3467 ( .A(\w3[3][13] ), .B(n2312), .Z(n2394) );
  XNOR U3468 ( .A(\w3[3][30] ), .B(n2394), .Z(n2314) );
  XNOR U3469 ( .A(\w3[3][5] ), .B(\w3[3][22] ), .Z(n2313) );
  XNOR U3470 ( .A(n2314), .B(n2313), .Z(\w0[4][29] ) );
  XOR U3471 ( .A(\w3[3][26] ), .B(n2315), .Z(n2316) );
  XNOR U3472 ( .A(n2317), .B(n2316), .Z(\w0[4][2] ) );
  XNOR U3473 ( .A(n2318), .B(\w3[3][31] ), .Z(n2445) );
  XOR U3474 ( .A(n2319), .B(n2445), .Z(n2418) );
  XOR U3475 ( .A(\w3[3][6] ), .B(n2320), .Z(n2321) );
  XOR U3476 ( .A(n2418), .B(n2321), .Z(\w0[4][30] ) );
  XNOR U3477 ( .A(\w3[3][15] ), .B(\w3[3][23] ), .Z(n2443) );
  XOR U3478 ( .A(\w3[3][33] ), .B(\w3[3][57] ), .Z(n2359) );
  XNOR U3479 ( .A(\w3[3][48] ), .B(\w3[3][56] ), .Z(n2404) );
  XOR U3480 ( .A(n2404), .B(\w3[3][40] ), .Z(n2322) );
  XNOR U3481 ( .A(n2359), .B(n2322), .Z(\w0[4][32] ) );
  XOR U3482 ( .A(\w3[3][34] ), .B(\w3[3][58] ), .Z(n2363) );
  XOR U3483 ( .A(\w3[3][41] ), .B(\w3[3][49] ), .Z(n2382) );
  XNOR U3484 ( .A(\w3[3][57] ), .B(n2382), .Z(n2323) );
  XNOR U3485 ( .A(n2363), .B(n2323), .Z(\w0[4][33] ) );
  XNOR U3486 ( .A(\w3[3][35] ), .B(\w3[3][59] ), .Z(n2343) );
  XNOR U3487 ( .A(\w3[3][42] ), .B(\w3[3][50] ), .Z(n2386) );
  XOR U3488 ( .A(\w3[3][58] ), .B(n2386), .Z(n2324) );
  XOR U3489 ( .A(n2343), .B(n2324), .Z(\w0[4][34] ) );
  XOR U3490 ( .A(\w3[3][36] ), .B(\w3[3][32] ), .Z(n2345) );
  XNOR U3491 ( .A(\w3[3][43] ), .B(\w3[3][51] ), .Z(n2365) );
  XOR U3492 ( .A(\w3[3][56] ), .B(n2365), .Z(n2325) );
  XNOR U3493 ( .A(\w3[3][60] ), .B(n2325), .Z(n2389) );
  XNOR U3494 ( .A(\w3[3][59] ), .B(n2389), .Z(n2326) );
  XNOR U3495 ( .A(n2345), .B(n2326), .Z(\w0[4][35] ) );
  XOR U3496 ( .A(\w3[3][32] ), .B(\w3[3][37] ), .Z(n2350) );
  XOR U3497 ( .A(\w3[3][44] ), .B(\w3[3][52] ), .Z(n2328) );
  XNOR U3498 ( .A(\w3[3][56] ), .B(\w3[3][61] ), .Z(n2327) );
  XOR U3499 ( .A(n2328), .B(n2327), .Z(n2395) );
  XOR U3500 ( .A(\w3[3][60] ), .B(n2395), .Z(n2329) );
  XNOR U3501 ( .A(n2350), .B(n2329), .Z(\w0[4][36] ) );
  XNOR U3502 ( .A(\w3[3][38] ), .B(\w3[3][62] ), .Z(n2354) );
  IV U3503 ( .A(\w3[3][53] ), .Z(n2368) );
  XOR U3504 ( .A(\w3[3][45] ), .B(n2368), .Z(n2398) );
  XOR U3505 ( .A(\w3[3][61] ), .B(n2398), .Z(n2330) );
  XOR U3506 ( .A(n2354), .B(n2330), .Z(\w0[4][37] ) );
  XOR U3507 ( .A(\w3[3][32] ), .B(\w3[3][39] ), .Z(n2355) );
  XNOR U3508 ( .A(\w3[3][56] ), .B(\w3[3][63] ), .Z(n2332) );
  XOR U3509 ( .A(\w3[3][46] ), .B(\w3[3][54] ), .Z(n2372) );
  XOR U3510 ( .A(n2332), .B(n2372), .Z(n2401) );
  XOR U3511 ( .A(\w3[3][62] ), .B(n2401), .Z(n2331) );
  XNOR U3512 ( .A(n2355), .B(n2331), .Z(\w0[4][38] ) );
  XNOR U3513 ( .A(\w3[3][47] ), .B(\w3[3][55] ), .Z(n2406) );
  XOR U3514 ( .A(\w3[3][32] ), .B(n2332), .Z(n2333) );
  XOR U3515 ( .A(n2406), .B(n2333), .Z(\w0[4][39] ) );
  XOR U3516 ( .A(n2334), .B(\w3[3][27] ), .Z(n2335) );
  XNOR U3517 ( .A(n2336), .B(n2335), .Z(\w0[4][3] ) );
  XOR U3518 ( .A(\w3[3][41] ), .B(\w3[3][32] ), .Z(n2338) );
  IV U3519 ( .A(\w3[3][33] ), .Z(n2383) );
  XNOR U3520 ( .A(n2404), .B(n2383), .Z(n2337) );
  XNOR U3521 ( .A(n2338), .B(n2337), .Z(\w0[4][40] ) );
  XOR U3522 ( .A(\w3[3][34] ), .B(\w3[3][42] ), .Z(n2340) );
  XNOR U3523 ( .A(n2359), .B(\w3[3][49] ), .Z(n2339) );
  XNOR U3524 ( .A(n2340), .B(n2339), .Z(\w0[4][41] ) );
  XOR U3525 ( .A(\w3[3][35] ), .B(\w3[3][43] ), .Z(n2342) );
  XNOR U3526 ( .A(n2363), .B(\w3[3][50] ), .Z(n2341) );
  XNOR U3527 ( .A(n2342), .B(n2341), .Z(\w0[4][42] ) );
  IV U3528 ( .A(\w3[3][40] ), .Z(n2347) );
  XNOR U3529 ( .A(n2347), .B(n2343), .Z(n2344) );
  XOR U3530 ( .A(\w3[3][44] ), .B(n2344), .Z(n2366) );
  XNOR U3531 ( .A(\w3[3][51] ), .B(n2345), .Z(n2346) );
  XOR U3532 ( .A(n2366), .B(n2346), .Z(\w0[4][43] ) );
  XOR U3533 ( .A(\w3[3][36] ), .B(\w3[3][45] ), .Z(n2349) );
  XOR U3534 ( .A(n2347), .B(\w3[3][60] ), .Z(n2348) );
  XOR U3535 ( .A(n2349), .B(n2348), .Z(n2369) );
  XNOR U3536 ( .A(\w3[3][52] ), .B(n2350), .Z(n2351) );
  XOR U3537 ( .A(n2369), .B(n2351), .Z(\w0[4][44] ) );
  XNOR U3538 ( .A(\w3[3][61] ), .B(\w3[3][37] ), .Z(n2371) );
  XNOR U3539 ( .A(\w3[3][46] ), .B(n2371), .Z(n2353) );
  XOR U3540 ( .A(n2368), .B(\w3[3][38] ), .Z(n2352) );
  XNOR U3541 ( .A(n2353), .B(n2352), .Z(\w0[4][45] ) );
  XOR U3542 ( .A(\w3[3][40] ), .B(\w3[3][47] ), .Z(n2377) );
  XOR U3543 ( .A(n2354), .B(n2377), .Z(n2373) );
  XNOR U3544 ( .A(\w3[3][54] ), .B(n2355), .Z(n2356) );
  XOR U3545 ( .A(n2373), .B(n2356), .Z(\w0[4][46] ) );
  XOR U3546 ( .A(\w3[3][63] ), .B(\w3[3][39] ), .Z(n2375) );
  XNOR U3547 ( .A(\w3[3][40] ), .B(\w3[3][32] ), .Z(n2378) );
  XOR U3548 ( .A(\w3[3][55] ), .B(n2378), .Z(n2357) );
  XNOR U3549 ( .A(n2375), .B(n2357), .Z(\w0[4][47] ) );
  XNOR U3550 ( .A(\w3[3][56] ), .B(n2382), .Z(n2358) );
  XOR U3551 ( .A(n2378), .B(n2358), .Z(\w0[4][48] ) );
  XOR U3552 ( .A(n2360), .B(\w3[3][28] ), .Z(n2361) );
  XOR U3553 ( .A(n2362), .B(n2361), .Z(\w0[4][4] ) );
  XNOR U3554 ( .A(n2363), .B(\w3[3][42] ), .Z(n2364) );
  XOR U3555 ( .A(n2365), .B(n2364), .Z(\w0[4][50] ) );
  IV U3556 ( .A(\w3[3][48] ), .Z(n2379) );
  XOR U3557 ( .A(n2379), .B(\w3[3][52] ), .Z(n2391) );
  XOR U3558 ( .A(\w3[3][43] ), .B(n2366), .Z(n2367) );
  XOR U3559 ( .A(n2391), .B(n2367), .Z(\w0[4][51] ) );
  XOR U3560 ( .A(\w3[3][48] ), .B(n2368), .Z(n2397) );
  XOR U3561 ( .A(\w3[3][44] ), .B(n2369), .Z(n2370) );
  XOR U3562 ( .A(n2397), .B(n2370), .Z(\w0[4][52] ) );
  XOR U3563 ( .A(n2379), .B(\w3[3][55] ), .Z(n2403) );
  XOR U3564 ( .A(\w3[3][46] ), .B(n2373), .Z(n2374) );
  XOR U3565 ( .A(n2403), .B(n2374), .Z(\w0[4][54] ) );
  XOR U3566 ( .A(\w3[3][48] ), .B(n2375), .Z(n2376) );
  XOR U3567 ( .A(n2377), .B(n2376), .Z(\w0[4][55] ) );
  XNOR U3568 ( .A(\w3[3][49] ), .B(n2378), .Z(n2381) );
  XOR U3569 ( .A(n2379), .B(\w3[3][57] ), .Z(n2380) );
  XNOR U3570 ( .A(n2381), .B(n2380), .Z(\w0[4][56] ) );
  XOR U3571 ( .A(\w3[3][58] ), .B(\w3[3][50] ), .Z(n2385) );
  XOR U3572 ( .A(n2383), .B(n2382), .Z(n2384) );
  XNOR U3573 ( .A(n2385), .B(n2384), .Z(\w0[4][57] ) );
  XOR U3574 ( .A(\w3[3][59] ), .B(\w3[3][51] ), .Z(n2388) );
  XOR U3575 ( .A(\w3[3][34] ), .B(n2386), .Z(n2387) );
  XNOR U3576 ( .A(n2388), .B(n2387), .Z(\w0[4][58] ) );
  XNOR U3577 ( .A(\w3[3][35] ), .B(n2389), .Z(n2390) );
  XOR U3578 ( .A(n2391), .B(n2390), .Z(\w0[4][59] ) );
  XOR U3579 ( .A(\w3[3][29] ), .B(n2392), .Z(n2393) );
  XOR U3580 ( .A(n2394), .B(n2393), .Z(\w0[4][5] ) );
  XOR U3581 ( .A(\w3[3][36] ), .B(n2395), .Z(n2396) );
  XOR U3582 ( .A(n2397), .B(n2396), .Z(\w0[4][60] ) );
  XOR U3583 ( .A(\w3[3][62] ), .B(\w3[3][54] ), .Z(n2400) );
  XOR U3584 ( .A(\w3[3][37] ), .B(n2398), .Z(n2399) );
  XNOR U3585 ( .A(n2400), .B(n2399), .Z(\w0[4][61] ) );
  XOR U3586 ( .A(\w3[3][38] ), .B(n2401), .Z(n2402) );
  XOR U3587 ( .A(n2403), .B(n2402), .Z(\w0[4][62] ) );
  XOR U3588 ( .A(n2404), .B(\w3[3][39] ), .Z(n2405) );
  XOR U3589 ( .A(n2406), .B(n2405), .Z(\w0[4][63] ) );
  XOR U3590 ( .A(\w3[3][80] ), .B(\w3[3][88] ), .Z(n2488) );
  XOR U3591 ( .A(\w3[3][65] ), .B(n2488), .Z(n2422) );
  XNOR U3592 ( .A(\w3[3][89] ), .B(\w3[3][72] ), .Z(n2407) );
  XNOR U3593 ( .A(n2422), .B(n2407), .Z(\w0[4][64] ) );
  IV U3594 ( .A(\w3[3][66] ), .Z(n2471) );
  XOR U3595 ( .A(n2471), .B(\w3[3][90] ), .Z(n2448) );
  XNOR U3596 ( .A(\w3[3][73] ), .B(\w3[3][81] ), .Z(n2465) );
  XOR U3597 ( .A(\w3[3][89] ), .B(n2465), .Z(n2408) );
  XOR U3598 ( .A(n2448), .B(n2408), .Z(\w0[4][65] ) );
  XNOR U3599 ( .A(\w3[3][67] ), .B(\w3[3][91] ), .Z(n2428) );
  XOR U3600 ( .A(\w3[3][74] ), .B(\w3[3][82] ), .Z(n2470) );
  XNOR U3601 ( .A(\w3[3][90] ), .B(n2470), .Z(n2409) );
  XOR U3602 ( .A(n2428), .B(n2409), .Z(\w0[4][66] ) );
  XOR U3603 ( .A(\w3[3][68] ), .B(\w3[3][64] ), .Z(n2430) );
  XNOR U3604 ( .A(\w3[3][75] ), .B(\w3[3][83] ), .Z(n2449) );
  XOR U3605 ( .A(\w3[3][88] ), .B(n2449), .Z(n2410) );
  XNOR U3606 ( .A(\w3[3][92] ), .B(n2410), .Z(n2474) );
  XNOR U3607 ( .A(\w3[3][91] ), .B(n2474), .Z(n2411) );
  XNOR U3608 ( .A(n2430), .B(n2411), .Z(\w0[4][67] ) );
  XOR U3609 ( .A(\w3[3][64] ), .B(\w3[3][69] ), .Z(n2434) );
  XOR U3610 ( .A(\w3[3][76] ), .B(\w3[3][84] ), .Z(n2413) );
  XNOR U3611 ( .A(\w3[3][88] ), .B(\w3[3][93] ), .Z(n2412) );
  XOR U3612 ( .A(n2413), .B(n2412), .Z(n2477) );
  XOR U3613 ( .A(\w3[3][92] ), .B(n2477), .Z(n2414) );
  XNOR U3614 ( .A(n2434), .B(n2414), .Z(\w0[4][68] ) );
  XNOR U3615 ( .A(\w3[3][70] ), .B(\w3[3][94] ), .Z(n2438) );
  XNOR U3616 ( .A(\w3[3][77] ), .B(\w3[3][85] ), .Z(n2480) );
  XOR U3617 ( .A(\w3[3][93] ), .B(n2480), .Z(n2415) );
  XOR U3618 ( .A(n2438), .B(n2415), .Z(\w0[4][69] ) );
  XOR U3619 ( .A(n2416), .B(\w3[3][30] ), .Z(n2417) );
  XOR U3620 ( .A(n2418), .B(n2417), .Z(\w0[4][6] ) );
  XOR U3621 ( .A(\w3[3][64] ), .B(\w3[3][71] ), .Z(n2439) );
  XNOR U3622 ( .A(\w3[3][88] ), .B(\w3[3][95] ), .Z(n2420) );
  XOR U3623 ( .A(\w3[3][78] ), .B(\w3[3][86] ), .Z(n2456) );
  XOR U3624 ( .A(n2420), .B(n2456), .Z(n2483) );
  XOR U3625 ( .A(\w3[3][94] ), .B(n2483), .Z(n2419) );
  XNOR U3626 ( .A(n2439), .B(n2419), .Z(\w0[4][70] ) );
  XNOR U3627 ( .A(\w3[3][79] ), .B(\w3[3][87] ), .Z(n2486) );
  XOR U3628 ( .A(\w3[3][64] ), .B(n2420), .Z(n2421) );
  XOR U3629 ( .A(n2486), .B(n2421), .Z(\w0[4][71] ) );
  IV U3630 ( .A(\w3[3][64] ), .Z(n2441) );
  XNOR U3631 ( .A(n2422), .B(\w3[3][73] ), .Z(n2423) );
  XOR U3632 ( .A(n2441), .B(n2423), .Z(\w0[4][72] ) );
  XNOR U3633 ( .A(\w3[3][89] ), .B(\w3[3][65] ), .Z(n2447) );
  XNOR U3634 ( .A(\w3[3][74] ), .B(n2447), .Z(n2425) );
  XOR U3635 ( .A(\w3[3][81] ), .B(n2471), .Z(n2424) );
  XNOR U3636 ( .A(n2425), .B(n2424), .Z(\w0[4][73] ) );
  XOR U3637 ( .A(\w3[3][90] ), .B(\w3[3][82] ), .Z(n2467) );
  XOR U3638 ( .A(\w3[3][75] ), .B(n2467), .Z(n2427) );
  XNOR U3639 ( .A(\w3[3][66] ), .B(\w3[3][67] ), .Z(n2426) );
  XNOR U3640 ( .A(n2427), .B(n2426), .Z(\w0[4][74] ) );
  XOR U3641 ( .A(\w3[3][72] ), .B(n2428), .Z(n2429) );
  XOR U3642 ( .A(\w3[3][76] ), .B(n2429), .Z(n2450) );
  XNOR U3643 ( .A(\w3[3][83] ), .B(n2430), .Z(n2431) );
  XOR U3644 ( .A(n2450), .B(n2431), .Z(\w0[4][75] ) );
  XOR U3645 ( .A(\w3[3][68] ), .B(\w3[3][77] ), .Z(n2433) );
  XNOR U3646 ( .A(\w3[3][72] ), .B(\w3[3][92] ), .Z(n2432) );
  XOR U3647 ( .A(n2433), .B(n2432), .Z(n2452) );
  XNOR U3648 ( .A(\w3[3][84] ), .B(n2434), .Z(n2435) );
  XOR U3649 ( .A(n2452), .B(n2435), .Z(\w0[4][76] ) );
  XNOR U3650 ( .A(\w3[3][93] ), .B(\w3[3][69] ), .Z(n2454) );
  XNOR U3651 ( .A(\w3[3][78] ), .B(n2454), .Z(n2437) );
  XNOR U3652 ( .A(\w3[3][85] ), .B(\w3[3][70] ), .Z(n2436) );
  XNOR U3653 ( .A(n2437), .B(n2436), .Z(\w0[4][77] ) );
  XOR U3654 ( .A(\w3[3][72] ), .B(\w3[3][79] ), .Z(n2461) );
  XOR U3655 ( .A(n2438), .B(n2461), .Z(n2457) );
  XNOR U3656 ( .A(\w3[3][86] ), .B(n2439), .Z(n2440) );
  XOR U3657 ( .A(n2457), .B(n2440), .Z(\w0[4][78] ) );
  XOR U3658 ( .A(\w3[3][95] ), .B(\w3[3][71] ), .Z(n2459) );
  XOR U3659 ( .A(\w3[3][72] ), .B(n2441), .Z(n2462) );
  XOR U3660 ( .A(\w3[3][87] ), .B(n2462), .Z(n2442) );
  XNOR U3661 ( .A(n2459), .B(n2442), .Z(\w0[4][79] ) );
  XNOR U3662 ( .A(\w3[3][0] ), .B(n2443), .Z(n2444) );
  XOR U3663 ( .A(n2445), .B(n2444), .Z(\w0[4][7] ) );
  XOR U3664 ( .A(\w3[3][88] ), .B(n2465), .Z(n2446) );
  XOR U3665 ( .A(n2462), .B(n2446), .Z(\w0[4][80] ) );
  XNOR U3666 ( .A(\w3[3][80] ), .B(\w3[3][84] ), .Z(n2476) );
  XOR U3667 ( .A(\w3[3][75] ), .B(n2450), .Z(n2451) );
  XOR U3668 ( .A(n2476), .B(n2451), .Z(\w0[4][83] ) );
  XNOR U3669 ( .A(\w3[3][80] ), .B(\w3[3][85] ), .Z(n2479) );
  XOR U3670 ( .A(\w3[3][76] ), .B(n2452), .Z(n2453) );
  XOR U3671 ( .A(n2479), .B(n2453), .Z(\w0[4][84] ) );
  XNOR U3672 ( .A(\w3[3][77] ), .B(n2454), .Z(n2455) );
  XOR U3673 ( .A(n2456), .B(n2455), .Z(\w0[4][85] ) );
  XNOR U3674 ( .A(\w3[3][80] ), .B(\w3[3][87] ), .Z(n2485) );
  XOR U3675 ( .A(\w3[3][78] ), .B(n2457), .Z(n2458) );
  XOR U3676 ( .A(n2485), .B(n2458), .Z(\w0[4][86] ) );
  XOR U3677 ( .A(\w3[3][80] ), .B(n2459), .Z(n2460) );
  XOR U3678 ( .A(n2461), .B(n2460), .Z(\w0[4][87] ) );
  XNOR U3679 ( .A(\w3[3][81] ), .B(n2462), .Z(n2464) );
  XNOR U3680 ( .A(\w3[3][89] ), .B(\w3[3][80] ), .Z(n2463) );
  XNOR U3681 ( .A(n2464), .B(n2463), .Z(\w0[4][88] ) );
  XOR U3682 ( .A(\w3[3][65] ), .B(n2465), .Z(n2466) );
  XNOR U3683 ( .A(n2467), .B(n2466), .Z(\w0[4][89] ) );
  XOR U3684 ( .A(\w3[3][91] ), .B(\w3[3][83] ), .Z(n2473) );
  XOR U3685 ( .A(n2471), .B(n2470), .Z(n2472) );
  XNOR U3686 ( .A(n2473), .B(n2472), .Z(\w0[4][90] ) );
  XNOR U3687 ( .A(\w3[3][67] ), .B(n2474), .Z(n2475) );
  XOR U3688 ( .A(n2476), .B(n2475), .Z(\w0[4][91] ) );
  XOR U3689 ( .A(\w3[3][68] ), .B(n2477), .Z(n2478) );
  XOR U3690 ( .A(n2479), .B(n2478), .Z(\w0[4][92] ) );
  XOR U3691 ( .A(\w3[3][94] ), .B(\w3[3][86] ), .Z(n2482) );
  XOR U3692 ( .A(\w3[3][69] ), .B(n2480), .Z(n2481) );
  XNOR U3693 ( .A(n2482), .B(n2481), .Z(\w0[4][93] ) );
  XOR U3694 ( .A(\w3[3][70] ), .B(n2483), .Z(n2484) );
  XOR U3695 ( .A(n2485), .B(n2484), .Z(\w0[4][94] ) );
  XNOR U3696 ( .A(\w3[3][71] ), .B(n2486), .Z(n2487) );
  XOR U3697 ( .A(n2488), .B(n2487), .Z(\w0[4][95] ) );
  XOR U3698 ( .A(n2489), .B(\w3[3][104] ), .Z(n2490) );
  XNOR U3699 ( .A(n2491), .B(n2490), .Z(\w0[4][96] ) );
  XOR U3700 ( .A(\w3[3][105] ), .B(n2492), .Z(n2493) );
  XNOR U3701 ( .A(n2494), .B(n2493), .Z(\w0[4][97] ) );
  XNOR U3702 ( .A(n2496), .B(n2495), .Z(n2497) );
  XOR U3703 ( .A(n2498), .B(n2497), .Z(\w0[4][98] ) );
  XNOR U3704 ( .A(n2500), .B(n2499), .Z(n2501) );
  XNOR U3705 ( .A(n2502), .B(n2501), .Z(\w0[4][99] ) );
  XOR U3706 ( .A(\w3[3][17] ), .B(\w3[3][10] ), .Z(n2505) );
  XOR U3707 ( .A(n2503), .B(\w3[3][2] ), .Z(n2504) );
  XNOR U3708 ( .A(n2505), .B(n2504), .Z(\w0[4][9] ) );
  NANDN U3709 ( .A(n2203), .B(state[0]), .Z(n2507) );
  NANDN U3710 ( .A(init), .B(msg[0]), .Z(n2506) );
  NAND U3711 ( .A(n2507), .B(n2506), .Z(n2508) );
  XOR U3712 ( .A(key[0]), .B(n2508), .Z(\w1[0][0] ) );
  NANDN U3713 ( .A(n2203), .B(state[100]), .Z(n2510) );
  NANDN U3714 ( .A(init), .B(msg[100]), .Z(n2509) );
  NAND U3715 ( .A(n2510), .B(n2509), .Z(n2511) );
  XOR U3716 ( .A(key[100]), .B(n2511), .Z(\w1[0][100] ) );
  NANDN U3717 ( .A(n2203), .B(state[101]), .Z(n2513) );
  NANDN U3718 ( .A(init), .B(msg[101]), .Z(n2512) );
  NAND U3719 ( .A(n2513), .B(n2512), .Z(n2514) );
  XOR U3720 ( .A(key[101]), .B(n2514), .Z(\w1[0][101] ) );
  NANDN U3721 ( .A(n2203), .B(state[102]), .Z(n2516) );
  NANDN U3722 ( .A(init), .B(msg[102]), .Z(n2515) );
  NAND U3723 ( .A(n2516), .B(n2515), .Z(n2517) );
  XOR U3724 ( .A(key[102]), .B(n2517), .Z(\w1[0][102] ) );
  NANDN U3725 ( .A(n2203), .B(state[103]), .Z(n2519) );
  NANDN U3726 ( .A(init), .B(msg[103]), .Z(n2518) );
  NAND U3727 ( .A(n2519), .B(n2518), .Z(n2520) );
  XOR U3728 ( .A(key[103]), .B(n2520), .Z(\w1[0][103] ) );
  NANDN U3729 ( .A(n2203), .B(state[104]), .Z(n2522) );
  NANDN U3730 ( .A(init), .B(msg[104]), .Z(n2521) );
  NAND U3731 ( .A(n2522), .B(n2521), .Z(n2523) );
  XOR U3732 ( .A(key[104]), .B(n2523), .Z(\w1[0][104] ) );
  NANDN U3733 ( .A(n2203), .B(state[105]), .Z(n2525) );
  NANDN U3734 ( .A(init), .B(msg[105]), .Z(n2524) );
  NAND U3735 ( .A(n2525), .B(n2524), .Z(n2526) );
  XOR U3736 ( .A(key[105]), .B(n2526), .Z(\w1[0][105] ) );
  NANDN U3737 ( .A(n2203), .B(state[106]), .Z(n2528) );
  NANDN U3738 ( .A(init), .B(msg[106]), .Z(n2527) );
  NAND U3739 ( .A(n2528), .B(n2527), .Z(n2529) );
  XOR U3740 ( .A(key[106]), .B(n2529), .Z(\w1[0][106] ) );
  NANDN U3741 ( .A(n2203), .B(state[107]), .Z(n2531) );
  NANDN U3742 ( .A(init), .B(msg[107]), .Z(n2530) );
  NAND U3743 ( .A(n2531), .B(n2530), .Z(n2532) );
  XOR U3744 ( .A(key[107]), .B(n2532), .Z(\w1[0][107] ) );
  NANDN U3745 ( .A(n2203), .B(state[108]), .Z(n2534) );
  NANDN U3746 ( .A(init), .B(msg[108]), .Z(n2533) );
  NAND U3747 ( .A(n2534), .B(n2533), .Z(n2535) );
  XOR U3748 ( .A(key[108]), .B(n2535), .Z(\w1[0][108] ) );
  NANDN U3749 ( .A(n2203), .B(state[109]), .Z(n2537) );
  NANDN U3750 ( .A(init), .B(msg[109]), .Z(n2536) );
  NAND U3751 ( .A(n2537), .B(n2536), .Z(n2538) );
  XOR U3752 ( .A(key[109]), .B(n2538), .Z(\w1[0][109] ) );
  NANDN U3753 ( .A(n2203), .B(state[10]), .Z(n2540) );
  NANDN U3754 ( .A(init), .B(msg[10]), .Z(n2539) );
  NAND U3755 ( .A(n2540), .B(n2539), .Z(n2541) );
  XOR U3756 ( .A(key[10]), .B(n2541), .Z(\w1[0][10] ) );
  NANDN U3757 ( .A(n2203), .B(state[110]), .Z(n2543) );
  NANDN U3758 ( .A(init), .B(msg[110]), .Z(n2542) );
  NAND U3759 ( .A(n2543), .B(n2542), .Z(n2544) );
  XOR U3760 ( .A(key[110]), .B(n2544), .Z(\w1[0][110] ) );
  NANDN U3761 ( .A(n2203), .B(state[111]), .Z(n2546) );
  NANDN U3762 ( .A(init), .B(msg[111]), .Z(n2545) );
  NAND U3763 ( .A(n2546), .B(n2545), .Z(n2547) );
  XOR U3764 ( .A(key[111]), .B(n2547), .Z(\w1[0][111] ) );
  NANDN U3765 ( .A(n2203), .B(state[112]), .Z(n2549) );
  NANDN U3766 ( .A(init), .B(msg[112]), .Z(n2548) );
  NAND U3767 ( .A(n2549), .B(n2548), .Z(n2550) );
  XOR U3768 ( .A(key[112]), .B(n2550), .Z(\w1[0][112] ) );
  NANDN U3769 ( .A(n2203), .B(state[113]), .Z(n2552) );
  NANDN U3770 ( .A(init), .B(msg[113]), .Z(n2551) );
  NAND U3771 ( .A(n2552), .B(n2551), .Z(n2553) );
  XOR U3772 ( .A(key[113]), .B(n2553), .Z(\w1[0][113] ) );
  NANDN U3773 ( .A(n2203), .B(state[114]), .Z(n2555) );
  NANDN U3774 ( .A(init), .B(msg[114]), .Z(n2554) );
  NAND U3775 ( .A(n2555), .B(n2554), .Z(n2556) );
  XOR U3776 ( .A(key[114]), .B(n2556), .Z(\w1[0][114] ) );
  NANDN U3777 ( .A(n2203), .B(state[115]), .Z(n2558) );
  NANDN U3778 ( .A(init), .B(msg[115]), .Z(n2557) );
  NAND U3779 ( .A(n2558), .B(n2557), .Z(n2559) );
  XOR U3780 ( .A(key[115]), .B(n2559), .Z(\w1[0][115] ) );
  NANDN U3781 ( .A(n2203), .B(state[116]), .Z(n2561) );
  NANDN U3782 ( .A(init), .B(msg[116]), .Z(n2560) );
  NAND U3783 ( .A(n2561), .B(n2560), .Z(n2562) );
  XOR U3784 ( .A(key[116]), .B(n2562), .Z(\w1[0][116] ) );
  NANDN U3785 ( .A(n2203), .B(state[117]), .Z(n2564) );
  NANDN U3786 ( .A(init), .B(msg[117]), .Z(n2563) );
  NAND U3787 ( .A(n2564), .B(n2563), .Z(n2565) );
  XOR U3788 ( .A(key[117]), .B(n2565), .Z(\w1[0][117] ) );
  NANDN U3789 ( .A(n2203), .B(state[118]), .Z(n2567) );
  NANDN U3790 ( .A(init), .B(msg[118]), .Z(n2566) );
  NAND U3791 ( .A(n2567), .B(n2566), .Z(n2568) );
  XOR U3792 ( .A(key[118]), .B(n2568), .Z(\w1[0][118] ) );
  NANDN U3793 ( .A(n2203), .B(state[119]), .Z(n2570) );
  NANDN U3794 ( .A(init), .B(msg[119]), .Z(n2569) );
  NAND U3795 ( .A(n2570), .B(n2569), .Z(n2571) );
  XOR U3796 ( .A(key[119]), .B(n2571), .Z(\w1[0][119] ) );
  NANDN U3797 ( .A(n2203), .B(state[11]), .Z(n2573) );
  NANDN U3798 ( .A(init), .B(msg[11]), .Z(n2572) );
  NAND U3799 ( .A(n2573), .B(n2572), .Z(n2574) );
  XOR U3800 ( .A(key[11]), .B(n2574), .Z(\w1[0][11] ) );
  NANDN U3801 ( .A(n2203), .B(state[120]), .Z(n2576) );
  NANDN U3802 ( .A(init), .B(msg[120]), .Z(n2575) );
  NAND U3803 ( .A(n2576), .B(n2575), .Z(n2577) );
  XOR U3804 ( .A(key[120]), .B(n2577), .Z(\w1[0][120] ) );
  NANDN U3805 ( .A(n2203), .B(state[121]), .Z(n2579) );
  NANDN U3806 ( .A(init), .B(msg[121]), .Z(n2578) );
  NAND U3807 ( .A(n2579), .B(n2578), .Z(n2580) );
  XOR U3808 ( .A(key[121]), .B(n2580), .Z(\w1[0][121] ) );
  NANDN U3809 ( .A(n2203), .B(state[122]), .Z(n2582) );
  NANDN U3810 ( .A(init), .B(msg[122]), .Z(n2581) );
  NAND U3811 ( .A(n2582), .B(n2581), .Z(n2583) );
  XOR U3812 ( .A(key[122]), .B(n2583), .Z(\w1[0][122] ) );
  NANDN U3813 ( .A(n2203), .B(state[123]), .Z(n2585) );
  NANDN U3814 ( .A(init), .B(msg[123]), .Z(n2584) );
  NAND U3815 ( .A(n2585), .B(n2584), .Z(n2586) );
  XOR U3816 ( .A(key[123]), .B(n2586), .Z(\w1[0][123] ) );
  NANDN U3817 ( .A(n2203), .B(state[124]), .Z(n2588) );
  NANDN U3818 ( .A(init), .B(msg[124]), .Z(n2587) );
  NAND U3819 ( .A(n2588), .B(n2587), .Z(n2589) );
  XOR U3820 ( .A(key[124]), .B(n2589), .Z(\w1[0][124] ) );
  NANDN U3821 ( .A(n2203), .B(state[125]), .Z(n2591) );
  NANDN U3822 ( .A(init), .B(msg[125]), .Z(n2590) );
  NAND U3823 ( .A(n2591), .B(n2590), .Z(n2592) );
  XOR U3824 ( .A(key[125]), .B(n2592), .Z(\w1[0][125] ) );
  NANDN U3825 ( .A(n2203), .B(state[126]), .Z(n2594) );
  NANDN U3826 ( .A(init), .B(msg[126]), .Z(n2593) );
  NAND U3827 ( .A(n2594), .B(n2593), .Z(n2595) );
  XOR U3828 ( .A(key[126]), .B(n2595), .Z(\w1[0][126] ) );
  NANDN U3829 ( .A(n2203), .B(state[127]), .Z(n2597) );
  NANDN U3830 ( .A(init), .B(msg[127]), .Z(n2596) );
  NAND U3831 ( .A(n2597), .B(n2596), .Z(n2598) );
  XOR U3832 ( .A(key[127]), .B(n2598), .Z(\w1[0][127] ) );
  NANDN U3833 ( .A(n2203), .B(state[12]), .Z(n2600) );
  NANDN U3834 ( .A(init), .B(msg[12]), .Z(n2599) );
  NAND U3835 ( .A(n2600), .B(n2599), .Z(n2601) );
  XOR U3836 ( .A(key[12]), .B(n2601), .Z(\w1[0][12] ) );
  NANDN U3837 ( .A(n2203), .B(state[13]), .Z(n2603) );
  NANDN U3838 ( .A(init), .B(msg[13]), .Z(n2602) );
  NAND U3839 ( .A(n2603), .B(n2602), .Z(n2604) );
  XOR U3840 ( .A(key[13]), .B(n2604), .Z(\w1[0][13] ) );
  NANDN U3841 ( .A(n2203), .B(state[14]), .Z(n2606) );
  NANDN U3842 ( .A(init), .B(msg[14]), .Z(n2605) );
  NAND U3843 ( .A(n2606), .B(n2605), .Z(n2607) );
  XOR U3844 ( .A(key[14]), .B(n2607), .Z(\w1[0][14] ) );
  NANDN U3845 ( .A(n2203), .B(state[15]), .Z(n2609) );
  NANDN U3846 ( .A(init), .B(msg[15]), .Z(n2608) );
  NAND U3847 ( .A(n2609), .B(n2608), .Z(n2610) );
  XOR U3848 ( .A(key[15]), .B(n2610), .Z(\w1[0][15] ) );
  NANDN U3849 ( .A(n2203), .B(state[16]), .Z(n2612) );
  NANDN U3850 ( .A(init), .B(msg[16]), .Z(n2611) );
  NAND U3851 ( .A(n2612), .B(n2611), .Z(n2613) );
  XOR U3852 ( .A(key[16]), .B(n2613), .Z(\w1[0][16] ) );
  NANDN U3853 ( .A(n2203), .B(state[17]), .Z(n2615) );
  NANDN U3854 ( .A(init), .B(msg[17]), .Z(n2614) );
  NAND U3855 ( .A(n2615), .B(n2614), .Z(n2616) );
  XOR U3856 ( .A(key[17]), .B(n2616), .Z(\w1[0][17] ) );
  NANDN U3857 ( .A(n2203), .B(state[18]), .Z(n2618) );
  NANDN U3858 ( .A(init), .B(msg[18]), .Z(n2617) );
  NAND U3859 ( .A(n2618), .B(n2617), .Z(n2619) );
  XOR U3860 ( .A(key[18]), .B(n2619), .Z(\w1[0][18] ) );
  NANDN U3861 ( .A(n2203), .B(state[19]), .Z(n2621) );
  NANDN U3862 ( .A(init), .B(msg[19]), .Z(n2620) );
  NAND U3863 ( .A(n2621), .B(n2620), .Z(n2622) );
  XOR U3864 ( .A(key[19]), .B(n2622), .Z(\w1[0][19] ) );
  NANDN U3865 ( .A(n2203), .B(state[1]), .Z(n2624) );
  NANDN U3866 ( .A(init), .B(msg[1]), .Z(n2623) );
  NAND U3867 ( .A(n2624), .B(n2623), .Z(n2625) );
  XOR U3868 ( .A(key[1]), .B(n2625), .Z(\w1[0][1] ) );
  NANDN U3869 ( .A(n2203), .B(state[20]), .Z(n2627) );
  NANDN U3870 ( .A(init), .B(msg[20]), .Z(n2626) );
  NAND U3871 ( .A(n2627), .B(n2626), .Z(n2628) );
  XOR U3872 ( .A(key[20]), .B(n2628), .Z(\w1[0][20] ) );
  NANDN U3873 ( .A(n2203), .B(state[21]), .Z(n2630) );
  NANDN U3874 ( .A(init), .B(msg[21]), .Z(n2629) );
  NAND U3875 ( .A(n2630), .B(n2629), .Z(n2631) );
  XOR U3876 ( .A(key[21]), .B(n2631), .Z(\w1[0][21] ) );
  NANDN U3877 ( .A(n2203), .B(state[22]), .Z(n2633) );
  NANDN U3878 ( .A(init), .B(msg[22]), .Z(n2632) );
  NAND U3879 ( .A(n2633), .B(n2632), .Z(n2634) );
  XOR U3880 ( .A(key[22]), .B(n2634), .Z(\w1[0][22] ) );
  NANDN U3881 ( .A(n2203), .B(state[23]), .Z(n2636) );
  NANDN U3882 ( .A(init), .B(msg[23]), .Z(n2635) );
  NAND U3883 ( .A(n2636), .B(n2635), .Z(n2637) );
  XOR U3884 ( .A(key[23]), .B(n2637), .Z(\w1[0][23] ) );
  NANDN U3885 ( .A(n2203), .B(state[24]), .Z(n2639) );
  NANDN U3886 ( .A(init), .B(msg[24]), .Z(n2638) );
  NAND U3887 ( .A(n2639), .B(n2638), .Z(n2640) );
  XOR U3888 ( .A(key[24]), .B(n2640), .Z(\w1[0][24] ) );
  NANDN U3889 ( .A(n2203), .B(state[25]), .Z(n2642) );
  NANDN U3890 ( .A(init), .B(msg[25]), .Z(n2641) );
  NAND U3891 ( .A(n2642), .B(n2641), .Z(n2643) );
  XOR U3892 ( .A(key[25]), .B(n2643), .Z(\w1[0][25] ) );
  NANDN U3893 ( .A(n2203), .B(state[26]), .Z(n2645) );
  NANDN U3894 ( .A(init), .B(msg[26]), .Z(n2644) );
  NAND U3895 ( .A(n2645), .B(n2644), .Z(n2646) );
  XOR U3896 ( .A(key[26]), .B(n2646), .Z(\w1[0][26] ) );
  NANDN U3897 ( .A(n2203), .B(state[27]), .Z(n2648) );
  NANDN U3898 ( .A(init), .B(msg[27]), .Z(n2647) );
  NAND U3899 ( .A(n2648), .B(n2647), .Z(n2649) );
  XOR U3900 ( .A(key[27]), .B(n2649), .Z(\w1[0][27] ) );
  NANDN U3901 ( .A(n2203), .B(state[28]), .Z(n2651) );
  NANDN U3902 ( .A(init), .B(msg[28]), .Z(n2650) );
  NAND U3903 ( .A(n2651), .B(n2650), .Z(n2652) );
  XOR U3904 ( .A(key[28]), .B(n2652), .Z(\w1[0][28] ) );
  NANDN U3905 ( .A(n2203), .B(state[29]), .Z(n2654) );
  NANDN U3906 ( .A(init), .B(msg[29]), .Z(n2653) );
  NAND U3907 ( .A(n2654), .B(n2653), .Z(n2655) );
  XOR U3908 ( .A(key[29]), .B(n2655), .Z(\w1[0][29] ) );
  NANDN U3909 ( .A(n2203), .B(state[2]), .Z(n2657) );
  NANDN U3910 ( .A(init), .B(msg[2]), .Z(n2656) );
  NAND U3911 ( .A(n2657), .B(n2656), .Z(n2658) );
  XOR U3912 ( .A(key[2]), .B(n2658), .Z(\w1[0][2] ) );
  NANDN U3913 ( .A(n2203), .B(state[30]), .Z(n2660) );
  NANDN U3914 ( .A(init), .B(msg[30]), .Z(n2659) );
  NAND U3915 ( .A(n2660), .B(n2659), .Z(n2661) );
  XOR U3916 ( .A(key[30]), .B(n2661), .Z(\w1[0][30] ) );
  NANDN U3917 ( .A(n2203), .B(state[31]), .Z(n2663) );
  NANDN U3918 ( .A(init), .B(msg[31]), .Z(n2662) );
  NAND U3919 ( .A(n2663), .B(n2662), .Z(n2664) );
  XOR U3920 ( .A(key[31]), .B(n2664), .Z(\w1[0][31] ) );
  NANDN U3921 ( .A(n2203), .B(state[32]), .Z(n2666) );
  NANDN U3922 ( .A(init), .B(msg[32]), .Z(n2665) );
  NAND U3923 ( .A(n2666), .B(n2665), .Z(n2667) );
  XOR U3924 ( .A(key[32]), .B(n2667), .Z(\w1[0][32] ) );
  NANDN U3925 ( .A(n2203), .B(state[33]), .Z(n2669) );
  NANDN U3926 ( .A(init), .B(msg[33]), .Z(n2668) );
  NAND U3927 ( .A(n2669), .B(n2668), .Z(n2670) );
  XOR U3928 ( .A(key[33]), .B(n2670), .Z(\w1[0][33] ) );
  NANDN U3929 ( .A(n2203), .B(state[34]), .Z(n2672) );
  NANDN U3930 ( .A(init), .B(msg[34]), .Z(n2671) );
  NAND U3931 ( .A(n2672), .B(n2671), .Z(n2673) );
  XOR U3932 ( .A(key[34]), .B(n2673), .Z(\w1[0][34] ) );
  NANDN U3933 ( .A(n2203), .B(state[35]), .Z(n2675) );
  NANDN U3934 ( .A(init), .B(msg[35]), .Z(n2674) );
  NAND U3935 ( .A(n2675), .B(n2674), .Z(n2676) );
  XOR U3936 ( .A(key[35]), .B(n2676), .Z(\w1[0][35] ) );
  NANDN U3937 ( .A(n2203), .B(state[36]), .Z(n2678) );
  NANDN U3938 ( .A(init), .B(msg[36]), .Z(n2677) );
  NAND U3939 ( .A(n2678), .B(n2677), .Z(n2679) );
  XOR U3940 ( .A(key[36]), .B(n2679), .Z(\w1[0][36] ) );
  NANDN U3941 ( .A(n2203), .B(state[37]), .Z(n2681) );
  NANDN U3942 ( .A(init), .B(msg[37]), .Z(n2680) );
  NAND U3943 ( .A(n2681), .B(n2680), .Z(n2682) );
  XOR U3944 ( .A(key[37]), .B(n2682), .Z(\w1[0][37] ) );
  NANDN U3945 ( .A(n2203), .B(state[38]), .Z(n2684) );
  NANDN U3946 ( .A(init), .B(msg[38]), .Z(n2683) );
  NAND U3947 ( .A(n2684), .B(n2683), .Z(n2685) );
  XOR U3948 ( .A(key[38]), .B(n2685), .Z(\w1[0][38] ) );
  NANDN U3949 ( .A(n2203), .B(state[39]), .Z(n2687) );
  NANDN U3950 ( .A(init), .B(msg[39]), .Z(n2686) );
  NAND U3951 ( .A(n2687), .B(n2686), .Z(n2688) );
  XOR U3952 ( .A(key[39]), .B(n2688), .Z(\w1[0][39] ) );
  NANDN U3953 ( .A(n2203), .B(state[3]), .Z(n2690) );
  NANDN U3954 ( .A(init), .B(msg[3]), .Z(n2689) );
  NAND U3955 ( .A(n2690), .B(n2689), .Z(n2691) );
  XOR U3956 ( .A(key[3]), .B(n2691), .Z(\w1[0][3] ) );
  NANDN U3957 ( .A(n2203), .B(state[40]), .Z(n2693) );
  NANDN U3958 ( .A(init), .B(msg[40]), .Z(n2692) );
  NAND U3959 ( .A(n2693), .B(n2692), .Z(n2694) );
  XOR U3960 ( .A(key[40]), .B(n2694), .Z(\w1[0][40] ) );
  NANDN U3961 ( .A(n2203), .B(state[41]), .Z(n2696) );
  NANDN U3962 ( .A(init), .B(msg[41]), .Z(n2695) );
  NAND U3963 ( .A(n2696), .B(n2695), .Z(n2697) );
  XOR U3964 ( .A(key[41]), .B(n2697), .Z(\w1[0][41] ) );
  NANDN U3965 ( .A(n2203), .B(state[42]), .Z(n2699) );
  NANDN U3966 ( .A(init), .B(msg[42]), .Z(n2698) );
  NAND U3967 ( .A(n2699), .B(n2698), .Z(n2700) );
  XOR U3968 ( .A(key[42]), .B(n2700), .Z(\w1[0][42] ) );
  NANDN U3969 ( .A(n2203), .B(state[43]), .Z(n2702) );
  NANDN U3970 ( .A(init), .B(msg[43]), .Z(n2701) );
  NAND U3971 ( .A(n2702), .B(n2701), .Z(n2703) );
  XOR U3972 ( .A(key[43]), .B(n2703), .Z(\w1[0][43] ) );
  NANDN U3973 ( .A(n2203), .B(state[44]), .Z(n2705) );
  NANDN U3974 ( .A(init), .B(msg[44]), .Z(n2704) );
  NAND U3975 ( .A(n2705), .B(n2704), .Z(n2706) );
  XOR U3976 ( .A(key[44]), .B(n2706), .Z(\w1[0][44] ) );
  NANDN U3977 ( .A(n2203), .B(state[45]), .Z(n2708) );
  NANDN U3978 ( .A(init), .B(msg[45]), .Z(n2707) );
  NAND U3979 ( .A(n2708), .B(n2707), .Z(n2709) );
  XOR U3980 ( .A(key[45]), .B(n2709), .Z(\w1[0][45] ) );
  NANDN U3981 ( .A(n2203), .B(state[46]), .Z(n2711) );
  NANDN U3982 ( .A(init), .B(msg[46]), .Z(n2710) );
  NAND U3983 ( .A(n2711), .B(n2710), .Z(n2712) );
  XOR U3984 ( .A(key[46]), .B(n2712), .Z(\w1[0][46] ) );
  NANDN U3985 ( .A(n2203), .B(state[47]), .Z(n2714) );
  NANDN U3986 ( .A(init), .B(msg[47]), .Z(n2713) );
  NAND U3987 ( .A(n2714), .B(n2713), .Z(n2715) );
  XOR U3988 ( .A(key[47]), .B(n2715), .Z(\w1[0][47] ) );
  NANDN U3989 ( .A(n2203), .B(state[48]), .Z(n2717) );
  NANDN U3990 ( .A(init), .B(msg[48]), .Z(n2716) );
  NAND U3991 ( .A(n2717), .B(n2716), .Z(n2718) );
  XOR U3992 ( .A(key[48]), .B(n2718), .Z(\w1[0][48] ) );
  NANDN U3993 ( .A(n2203), .B(state[49]), .Z(n2720) );
  NANDN U3994 ( .A(init), .B(msg[49]), .Z(n2719) );
  NAND U3995 ( .A(n2720), .B(n2719), .Z(n2721) );
  XOR U3996 ( .A(key[49]), .B(n2721), .Z(\w1[0][49] ) );
  NANDN U3997 ( .A(n2203), .B(state[4]), .Z(n2723) );
  NANDN U3998 ( .A(init), .B(msg[4]), .Z(n2722) );
  NAND U3999 ( .A(n2723), .B(n2722), .Z(n2724) );
  XOR U4000 ( .A(key[4]), .B(n2724), .Z(\w1[0][4] ) );
  NANDN U4001 ( .A(n2203), .B(state[50]), .Z(n2726) );
  NANDN U4002 ( .A(init), .B(msg[50]), .Z(n2725) );
  NAND U4003 ( .A(n2726), .B(n2725), .Z(n2727) );
  XOR U4004 ( .A(key[50]), .B(n2727), .Z(\w1[0][50] ) );
  NANDN U4005 ( .A(n2203), .B(state[51]), .Z(n2729) );
  NANDN U4006 ( .A(init), .B(msg[51]), .Z(n2728) );
  NAND U4007 ( .A(n2729), .B(n2728), .Z(n2730) );
  XOR U4008 ( .A(key[51]), .B(n2730), .Z(\w1[0][51] ) );
  NANDN U4009 ( .A(n2203), .B(state[52]), .Z(n2732) );
  NANDN U4010 ( .A(init), .B(msg[52]), .Z(n2731) );
  NAND U4011 ( .A(n2732), .B(n2731), .Z(n2733) );
  XOR U4012 ( .A(key[52]), .B(n2733), .Z(\w1[0][52] ) );
  NANDN U4013 ( .A(n2203), .B(state[53]), .Z(n2735) );
  NANDN U4014 ( .A(init), .B(msg[53]), .Z(n2734) );
  NAND U4015 ( .A(n2735), .B(n2734), .Z(n2736) );
  XOR U4016 ( .A(key[53]), .B(n2736), .Z(\w1[0][53] ) );
  NANDN U4017 ( .A(n2203), .B(state[54]), .Z(n2738) );
  NANDN U4018 ( .A(init), .B(msg[54]), .Z(n2737) );
  NAND U4019 ( .A(n2738), .B(n2737), .Z(n2739) );
  XOR U4020 ( .A(key[54]), .B(n2739), .Z(\w1[0][54] ) );
  NANDN U4021 ( .A(n2203), .B(state[55]), .Z(n2741) );
  NANDN U4022 ( .A(init), .B(msg[55]), .Z(n2740) );
  NAND U4023 ( .A(n2741), .B(n2740), .Z(n2742) );
  XOR U4024 ( .A(key[55]), .B(n2742), .Z(\w1[0][55] ) );
  NANDN U4025 ( .A(n2203), .B(state[56]), .Z(n2744) );
  NANDN U4026 ( .A(init), .B(msg[56]), .Z(n2743) );
  NAND U4027 ( .A(n2744), .B(n2743), .Z(n2745) );
  XOR U4028 ( .A(key[56]), .B(n2745), .Z(\w1[0][56] ) );
  NANDN U4029 ( .A(n2203), .B(state[57]), .Z(n2747) );
  NANDN U4030 ( .A(init), .B(msg[57]), .Z(n2746) );
  NAND U4031 ( .A(n2747), .B(n2746), .Z(n2748) );
  XOR U4032 ( .A(key[57]), .B(n2748), .Z(\w1[0][57] ) );
  NANDN U4033 ( .A(n2203), .B(state[58]), .Z(n2750) );
  NANDN U4034 ( .A(init), .B(msg[58]), .Z(n2749) );
  NAND U4035 ( .A(n2750), .B(n2749), .Z(n2751) );
  XOR U4036 ( .A(key[58]), .B(n2751), .Z(\w1[0][58] ) );
  NANDN U4037 ( .A(n2203), .B(state[59]), .Z(n2753) );
  NANDN U4038 ( .A(init), .B(msg[59]), .Z(n2752) );
  NAND U4039 ( .A(n2753), .B(n2752), .Z(n2754) );
  XOR U4040 ( .A(key[59]), .B(n2754), .Z(\w1[0][59] ) );
  NANDN U4041 ( .A(n2203), .B(state[5]), .Z(n2756) );
  NANDN U4042 ( .A(init), .B(msg[5]), .Z(n2755) );
  NAND U4043 ( .A(n2756), .B(n2755), .Z(n2757) );
  XOR U4044 ( .A(key[5]), .B(n2757), .Z(\w1[0][5] ) );
  NANDN U4045 ( .A(n2203), .B(state[60]), .Z(n2759) );
  NANDN U4046 ( .A(init), .B(msg[60]), .Z(n2758) );
  NAND U4047 ( .A(n2759), .B(n2758), .Z(n2760) );
  XOR U4048 ( .A(key[60]), .B(n2760), .Z(\w1[0][60] ) );
  NANDN U4049 ( .A(n2203), .B(state[61]), .Z(n2762) );
  NANDN U4050 ( .A(init), .B(msg[61]), .Z(n2761) );
  NAND U4051 ( .A(n2762), .B(n2761), .Z(n2763) );
  XOR U4052 ( .A(key[61]), .B(n2763), .Z(\w1[0][61] ) );
  NANDN U4053 ( .A(n2203), .B(state[62]), .Z(n2765) );
  NANDN U4054 ( .A(init), .B(msg[62]), .Z(n2764) );
  NAND U4055 ( .A(n2765), .B(n2764), .Z(n2766) );
  XOR U4056 ( .A(key[62]), .B(n2766), .Z(\w1[0][62] ) );
  NANDN U4057 ( .A(n2203), .B(state[63]), .Z(n2768) );
  NANDN U4058 ( .A(init), .B(msg[63]), .Z(n2767) );
  NAND U4059 ( .A(n2768), .B(n2767), .Z(n2769) );
  XOR U4060 ( .A(key[63]), .B(n2769), .Z(\w1[0][63] ) );
  NANDN U4061 ( .A(n2203), .B(state[64]), .Z(n2771) );
  NANDN U4062 ( .A(init), .B(msg[64]), .Z(n2770) );
  NAND U4063 ( .A(n2771), .B(n2770), .Z(n2772) );
  XOR U4064 ( .A(key[64]), .B(n2772), .Z(\w1[0][64] ) );
  NANDN U4065 ( .A(n2203), .B(state[65]), .Z(n2774) );
  NANDN U4066 ( .A(init), .B(msg[65]), .Z(n2773) );
  NAND U4067 ( .A(n2774), .B(n2773), .Z(n2775) );
  XOR U4068 ( .A(key[65]), .B(n2775), .Z(\w1[0][65] ) );
  NANDN U4069 ( .A(n2203), .B(state[66]), .Z(n2777) );
  NANDN U4070 ( .A(init), .B(msg[66]), .Z(n2776) );
  NAND U4071 ( .A(n2777), .B(n2776), .Z(n2778) );
  XOR U4072 ( .A(key[66]), .B(n2778), .Z(\w1[0][66] ) );
  NANDN U4073 ( .A(n2203), .B(state[67]), .Z(n2780) );
  NANDN U4074 ( .A(init), .B(msg[67]), .Z(n2779) );
  NAND U4075 ( .A(n2780), .B(n2779), .Z(n2781) );
  XOR U4076 ( .A(key[67]), .B(n2781), .Z(\w1[0][67] ) );
  NANDN U4077 ( .A(n2203), .B(state[68]), .Z(n2783) );
  NANDN U4078 ( .A(init), .B(msg[68]), .Z(n2782) );
  NAND U4079 ( .A(n2783), .B(n2782), .Z(n2784) );
  XOR U4080 ( .A(key[68]), .B(n2784), .Z(\w1[0][68] ) );
  NANDN U4081 ( .A(n2203), .B(state[69]), .Z(n2786) );
  NANDN U4082 ( .A(init), .B(msg[69]), .Z(n2785) );
  NAND U4083 ( .A(n2786), .B(n2785), .Z(n2787) );
  XOR U4084 ( .A(key[69]), .B(n2787), .Z(\w1[0][69] ) );
  NANDN U4085 ( .A(n2203), .B(state[6]), .Z(n2789) );
  NANDN U4086 ( .A(init), .B(msg[6]), .Z(n2788) );
  NAND U4087 ( .A(n2789), .B(n2788), .Z(n2790) );
  XOR U4088 ( .A(key[6]), .B(n2790), .Z(\w1[0][6] ) );
  NANDN U4089 ( .A(n2203), .B(state[70]), .Z(n2792) );
  NANDN U4090 ( .A(init), .B(msg[70]), .Z(n2791) );
  NAND U4091 ( .A(n2792), .B(n2791), .Z(n2793) );
  XOR U4092 ( .A(key[70]), .B(n2793), .Z(\w1[0][70] ) );
  NANDN U4093 ( .A(n2203), .B(state[71]), .Z(n2795) );
  NANDN U4094 ( .A(init), .B(msg[71]), .Z(n2794) );
  NAND U4095 ( .A(n2795), .B(n2794), .Z(n2796) );
  XOR U4096 ( .A(key[71]), .B(n2796), .Z(\w1[0][71] ) );
  NANDN U4097 ( .A(n2203), .B(state[72]), .Z(n2798) );
  NANDN U4098 ( .A(init), .B(msg[72]), .Z(n2797) );
  NAND U4099 ( .A(n2798), .B(n2797), .Z(n2799) );
  XOR U4100 ( .A(key[72]), .B(n2799), .Z(\w1[0][72] ) );
  NANDN U4101 ( .A(n2203), .B(state[73]), .Z(n2801) );
  NANDN U4102 ( .A(init), .B(msg[73]), .Z(n2800) );
  NAND U4103 ( .A(n2801), .B(n2800), .Z(n2802) );
  XOR U4104 ( .A(key[73]), .B(n2802), .Z(\w1[0][73] ) );
  NANDN U4105 ( .A(n2203), .B(state[74]), .Z(n2804) );
  NANDN U4106 ( .A(init), .B(msg[74]), .Z(n2803) );
  NAND U4107 ( .A(n2804), .B(n2803), .Z(n2805) );
  XOR U4108 ( .A(key[74]), .B(n2805), .Z(\w1[0][74] ) );
  NANDN U4109 ( .A(n2203), .B(state[75]), .Z(n2807) );
  NANDN U4110 ( .A(init), .B(msg[75]), .Z(n2806) );
  NAND U4111 ( .A(n2807), .B(n2806), .Z(n2808) );
  XOR U4112 ( .A(key[75]), .B(n2808), .Z(\w1[0][75] ) );
  NANDN U4113 ( .A(n2203), .B(state[76]), .Z(n2810) );
  NANDN U4114 ( .A(init), .B(msg[76]), .Z(n2809) );
  NAND U4115 ( .A(n2810), .B(n2809), .Z(n2811) );
  XOR U4116 ( .A(key[76]), .B(n2811), .Z(\w1[0][76] ) );
  NANDN U4117 ( .A(n2203), .B(state[77]), .Z(n2813) );
  NANDN U4118 ( .A(init), .B(msg[77]), .Z(n2812) );
  NAND U4119 ( .A(n2813), .B(n2812), .Z(n2814) );
  XOR U4120 ( .A(key[77]), .B(n2814), .Z(\w1[0][77] ) );
  NANDN U4121 ( .A(n2203), .B(state[78]), .Z(n2816) );
  NANDN U4122 ( .A(init), .B(msg[78]), .Z(n2815) );
  NAND U4123 ( .A(n2816), .B(n2815), .Z(n2817) );
  XOR U4124 ( .A(key[78]), .B(n2817), .Z(\w1[0][78] ) );
  NANDN U4125 ( .A(n2203), .B(state[79]), .Z(n2819) );
  NANDN U4126 ( .A(init), .B(msg[79]), .Z(n2818) );
  NAND U4127 ( .A(n2819), .B(n2818), .Z(n2820) );
  XOR U4128 ( .A(key[79]), .B(n2820), .Z(\w1[0][79] ) );
  NANDN U4129 ( .A(n2203), .B(state[7]), .Z(n2822) );
  NANDN U4130 ( .A(init), .B(msg[7]), .Z(n2821) );
  NAND U4131 ( .A(n2822), .B(n2821), .Z(n2823) );
  XOR U4132 ( .A(key[7]), .B(n2823), .Z(\w1[0][7] ) );
  NANDN U4133 ( .A(n2203), .B(state[80]), .Z(n2825) );
  NANDN U4134 ( .A(init), .B(msg[80]), .Z(n2824) );
  NAND U4135 ( .A(n2825), .B(n2824), .Z(n2826) );
  XOR U4136 ( .A(key[80]), .B(n2826), .Z(\w1[0][80] ) );
  NANDN U4137 ( .A(n2203), .B(state[81]), .Z(n2828) );
  NANDN U4138 ( .A(init), .B(msg[81]), .Z(n2827) );
  NAND U4139 ( .A(n2828), .B(n2827), .Z(n2829) );
  XOR U4140 ( .A(key[81]), .B(n2829), .Z(\w1[0][81] ) );
  NANDN U4141 ( .A(n2203), .B(state[82]), .Z(n2831) );
  NANDN U4142 ( .A(init), .B(msg[82]), .Z(n2830) );
  NAND U4143 ( .A(n2831), .B(n2830), .Z(n2832) );
  XOR U4144 ( .A(key[82]), .B(n2832), .Z(\w1[0][82] ) );
  NANDN U4145 ( .A(n2203), .B(state[83]), .Z(n2834) );
  NANDN U4146 ( .A(init), .B(msg[83]), .Z(n2833) );
  NAND U4147 ( .A(n2834), .B(n2833), .Z(n2835) );
  XOR U4148 ( .A(key[83]), .B(n2835), .Z(\w1[0][83] ) );
  NANDN U4149 ( .A(n2203), .B(state[84]), .Z(n2837) );
  NANDN U4150 ( .A(init), .B(msg[84]), .Z(n2836) );
  NAND U4151 ( .A(n2837), .B(n2836), .Z(n2838) );
  XOR U4152 ( .A(key[84]), .B(n2838), .Z(\w1[0][84] ) );
  NANDN U4153 ( .A(n2203), .B(state[85]), .Z(n2840) );
  NANDN U4154 ( .A(init), .B(msg[85]), .Z(n2839) );
  NAND U4155 ( .A(n2840), .B(n2839), .Z(n2841) );
  XOR U4156 ( .A(key[85]), .B(n2841), .Z(\w1[0][85] ) );
  NANDN U4157 ( .A(n2203), .B(state[86]), .Z(n2843) );
  NANDN U4158 ( .A(init), .B(msg[86]), .Z(n2842) );
  NAND U4159 ( .A(n2843), .B(n2842), .Z(n2844) );
  XOR U4160 ( .A(key[86]), .B(n2844), .Z(\w1[0][86] ) );
  NANDN U4161 ( .A(n2203), .B(state[87]), .Z(n2846) );
  NANDN U4162 ( .A(init), .B(msg[87]), .Z(n2845) );
  NAND U4163 ( .A(n2846), .B(n2845), .Z(n2847) );
  XOR U4164 ( .A(key[87]), .B(n2847), .Z(\w1[0][87] ) );
  NANDN U4165 ( .A(n2203), .B(state[88]), .Z(n2849) );
  NANDN U4166 ( .A(init), .B(msg[88]), .Z(n2848) );
  NAND U4167 ( .A(n2849), .B(n2848), .Z(n2850) );
  XOR U4168 ( .A(key[88]), .B(n2850), .Z(\w1[0][88] ) );
  NANDN U4169 ( .A(n2203), .B(state[89]), .Z(n2852) );
  NANDN U4170 ( .A(init), .B(msg[89]), .Z(n2851) );
  NAND U4171 ( .A(n2852), .B(n2851), .Z(n2853) );
  XOR U4172 ( .A(key[89]), .B(n2853), .Z(\w1[0][89] ) );
  NANDN U4173 ( .A(n2203), .B(state[8]), .Z(n2855) );
  NANDN U4174 ( .A(init), .B(msg[8]), .Z(n2854) );
  NAND U4175 ( .A(n2855), .B(n2854), .Z(n2856) );
  XOR U4176 ( .A(key[8]), .B(n2856), .Z(\w1[0][8] ) );
  NANDN U4177 ( .A(n2203), .B(state[90]), .Z(n2858) );
  NANDN U4178 ( .A(init), .B(msg[90]), .Z(n2857) );
  NAND U4179 ( .A(n2858), .B(n2857), .Z(n2859) );
  XOR U4180 ( .A(key[90]), .B(n2859), .Z(\w1[0][90] ) );
  NANDN U4181 ( .A(n2203), .B(state[91]), .Z(n2861) );
  NANDN U4182 ( .A(init), .B(msg[91]), .Z(n2860) );
  NAND U4183 ( .A(n2861), .B(n2860), .Z(n2862) );
  XOR U4184 ( .A(key[91]), .B(n2862), .Z(\w1[0][91] ) );
  NANDN U4185 ( .A(n2203), .B(state[92]), .Z(n2864) );
  NANDN U4186 ( .A(init), .B(msg[92]), .Z(n2863) );
  NAND U4187 ( .A(n2864), .B(n2863), .Z(n2865) );
  XOR U4188 ( .A(key[92]), .B(n2865), .Z(\w1[0][92] ) );
  NANDN U4189 ( .A(n2203), .B(state[93]), .Z(n2867) );
  NANDN U4190 ( .A(init), .B(msg[93]), .Z(n2866) );
  NAND U4191 ( .A(n2867), .B(n2866), .Z(n2868) );
  XOR U4192 ( .A(key[93]), .B(n2868), .Z(\w1[0][93] ) );
  NANDN U4193 ( .A(n2203), .B(state[94]), .Z(n2870) );
  NANDN U4194 ( .A(init), .B(msg[94]), .Z(n2869) );
  NAND U4195 ( .A(n2870), .B(n2869), .Z(n2871) );
  XOR U4196 ( .A(key[94]), .B(n2871), .Z(\w1[0][94] ) );
  NANDN U4197 ( .A(n2203), .B(state[95]), .Z(n2873) );
  NANDN U4198 ( .A(init), .B(msg[95]), .Z(n2872) );
  NAND U4199 ( .A(n2873), .B(n2872), .Z(n2874) );
  XOR U4200 ( .A(key[95]), .B(n2874), .Z(\w1[0][95] ) );
  NANDN U4201 ( .A(n2203), .B(state[96]), .Z(n2876) );
  NANDN U4202 ( .A(init), .B(msg[96]), .Z(n2875) );
  NAND U4203 ( .A(n2876), .B(n2875), .Z(n2877) );
  XOR U4204 ( .A(key[96]), .B(n2877), .Z(\w1[0][96] ) );
  NANDN U4205 ( .A(n2203), .B(state[97]), .Z(n2879) );
  NANDN U4206 ( .A(init), .B(msg[97]), .Z(n2878) );
  NAND U4207 ( .A(n2879), .B(n2878), .Z(n2880) );
  XOR U4208 ( .A(key[97]), .B(n2880), .Z(\w1[0][97] ) );
  NANDN U4209 ( .A(n2203), .B(state[98]), .Z(n2882) );
  NANDN U4210 ( .A(init), .B(msg[98]), .Z(n2881) );
  NAND U4211 ( .A(n2882), .B(n2881), .Z(n2883) );
  XOR U4212 ( .A(key[98]), .B(n2883), .Z(\w1[0][98] ) );
  NANDN U4213 ( .A(n2203), .B(state[99]), .Z(n2885) );
  NANDN U4214 ( .A(init), .B(msg[99]), .Z(n2884) );
  NAND U4215 ( .A(n2885), .B(n2884), .Z(n2886) );
  XOR U4216 ( .A(key[99]), .B(n2886), .Z(\w1[0][99] ) );
  NANDN U4217 ( .A(n2203), .B(state[9]), .Z(n2888) );
  NANDN U4218 ( .A(init), .B(msg[9]), .Z(n2887) );
  NAND U4219 ( .A(n2888), .B(n2887), .Z(n2889) );
  XOR U4220 ( .A(key[9]), .B(n2889), .Z(\w1[0][9] ) );
  XNOR U4221 ( .A(\w3[0][1] ), .B(\w3[0][25] ), .Z(n3305) );
  IV U4222 ( .A(\w3[0][24] ), .Z(n3051) );
  XOR U4223 ( .A(\w3[0][16] ), .B(n3051), .Z(n3257) );
  XNOR U4224 ( .A(\w3[0][8] ), .B(key[128]), .Z(n2890) );
  XNOR U4225 ( .A(n3257), .B(n2890), .Z(n2891) );
  XOR U4226 ( .A(n3305), .B(n2891), .Z(\w1[1][0] ) );
  XOR U4227 ( .A(\w3[0][96] ), .B(\w3[0][101] ), .Z(n2914) );
  XOR U4228 ( .A(\w3[0][116] ), .B(\w3[0][125] ), .Z(n2893) );
  IV U4229 ( .A(\w3[0][120] ), .Z(n2966) );
  XOR U4230 ( .A(n2966), .B(\w3[0][108] ), .Z(n2892) );
  XOR U4231 ( .A(n2893), .B(n2892), .Z(n2974) );
  XOR U4232 ( .A(n2974), .B(key[228]), .Z(n2894) );
  XOR U4233 ( .A(n2914), .B(n2894), .Z(n2895) );
  XNOR U4234 ( .A(\w3[0][124] ), .B(n2895), .Z(\w1[1][100] ) );
  XNOR U4235 ( .A(\w3[0][102] ), .B(\w3[0][126] ), .Z(n2923) );
  XNOR U4236 ( .A(n2923), .B(key[229]), .Z(n2897) );
  XNOR U4237 ( .A(\w3[0][109] ), .B(\w3[0][117] ), .Z(n2977) );
  XOR U4238 ( .A(\w3[0][125] ), .B(n2977), .Z(n2896) );
  XNOR U4239 ( .A(n2897), .B(n2896), .Z(\w1[1][101] ) );
  XOR U4240 ( .A(\w3[0][96] ), .B(\w3[0][103] ), .Z(n2924) );
  XOR U4241 ( .A(n2924), .B(key[230]), .Z(n2899) );
  XNOR U4242 ( .A(\w3[0][110] ), .B(\w3[0][118] ), .Z(n2942) );
  XNOR U4243 ( .A(n2966), .B(\w3[0][127] ), .Z(n2900) );
  XOR U4244 ( .A(n2942), .B(n2900), .Z(n2982) );
  XOR U4245 ( .A(\w3[0][126] ), .B(n2982), .Z(n2898) );
  XNOR U4246 ( .A(n2899), .B(n2898), .Z(\w1[1][102] ) );
  XNOR U4247 ( .A(\w3[0][111] ), .B(\w3[0][119] ), .Z(n2985) );
  XNOR U4248 ( .A(n2985), .B(key[231]), .Z(n2902) );
  XNOR U4249 ( .A(\w3[0][96] ), .B(n2900), .Z(n2901) );
  XNOR U4250 ( .A(n2902), .B(n2901), .Z(\w1[1][103] ) );
  IV U4251 ( .A(\w3[0][97] ), .Z(n2962) );
  IV U4252 ( .A(\w3[0][112] ), .Z(n2958) );
  XOR U4253 ( .A(\w3[0][120] ), .B(n2958), .Z(n3286) );
  XOR U4254 ( .A(\w3[0][106] ), .B(\w3[0][113] ), .Z(n2904) );
  XNOR U4255 ( .A(\w3[0][97] ), .B(\w3[0][121] ), .Z(n3285) );
  XOR U4256 ( .A(n3285), .B(key[233]), .Z(n2903) );
  XNOR U4257 ( .A(n2904), .B(n2903), .Z(n2905) );
  XOR U4258 ( .A(\w3[0][98] ), .B(n2905), .Z(\w1[1][105] ) );
  XOR U4259 ( .A(\w3[0][107] ), .B(\w3[0][114] ), .Z(n2907) );
  XOR U4260 ( .A(\w3[0][98] ), .B(\w3[0][122] ), .Z(n3290) );
  XNOR U4261 ( .A(n3290), .B(key[234]), .Z(n2906) );
  XNOR U4262 ( .A(n2907), .B(n2906), .Z(n2908) );
  XOR U4263 ( .A(\w3[0][99] ), .B(n2908), .Z(\w1[1][106] ) );
  XNOR U4264 ( .A(\w3[0][99] ), .B(\w3[0][123] ), .Z(n3294) );
  XOR U4265 ( .A(\w3[0][108] ), .B(n3294), .Z(n2909) );
  XOR U4266 ( .A(\w3[0][104] ), .B(n2909), .Z(n2935) );
  XNOR U4267 ( .A(n2935), .B(key[235]), .Z(n2911) );
  IV U4268 ( .A(\w3[0][100] ), .Z(n2973) );
  XOR U4269 ( .A(\w3[0][96] ), .B(n2973), .Z(n3298) );
  XOR U4270 ( .A(\w3[0][115] ), .B(n3298), .Z(n2910) );
  XNOR U4271 ( .A(n2911), .B(n2910), .Z(\w1[1][107] ) );
  XOR U4272 ( .A(\w3[0][100] ), .B(\w3[0][104] ), .Z(n2913) );
  XNOR U4273 ( .A(\w3[0][124] ), .B(\w3[0][109] ), .Z(n2912) );
  XOR U4274 ( .A(n2913), .B(n2912), .Z(n2938) );
  XNOR U4275 ( .A(n2938), .B(key[236]), .Z(n2916) );
  XNOR U4276 ( .A(\w3[0][116] ), .B(n2914), .Z(n2915) );
  XNOR U4277 ( .A(n2916), .B(n2915), .Z(\w1[1][108] ) );
  XNOR U4278 ( .A(\w3[0][125] ), .B(\w3[0][101] ), .Z(n2941) );
  XNOR U4279 ( .A(n2941), .B(key[237]), .Z(n2918) );
  XNOR U4280 ( .A(\w3[0][102] ), .B(\w3[0][110] ), .Z(n2917) );
  XNOR U4281 ( .A(n2918), .B(n2917), .Z(n2919) );
  XOR U4282 ( .A(\w3[0][117] ), .B(n2919), .Z(\w1[1][109] ) );
  IV U4283 ( .A(\w3[0][18] ), .Z(n3027) );
  XNOR U4284 ( .A(\w3[0][11] ), .B(n3027), .Z(n2921) );
  XNOR U4285 ( .A(\w3[0][2] ), .B(\w3[0][26] ), .Z(n3006) );
  XOR U4286 ( .A(n3006), .B(key[138]), .Z(n2920) );
  XNOR U4287 ( .A(n2921), .B(n2920), .Z(n2922) );
  XOR U4288 ( .A(\w3[0][3] ), .B(n2922), .Z(\w1[1][10] ) );
  XOR U4289 ( .A(\w3[0][111] ), .B(\w3[0][104] ), .Z(n2949) );
  XOR U4290 ( .A(n2923), .B(n2949), .Z(n2945) );
  XNOR U4291 ( .A(n2945), .B(key[238]), .Z(n2926) );
  XNOR U4292 ( .A(\w3[0][118] ), .B(n2924), .Z(n2925) );
  XNOR U4293 ( .A(n2926), .B(n2925), .Z(\w1[1][110] ) );
  XOR U4294 ( .A(\w3[0][127] ), .B(\w3[0][103] ), .Z(n2948) );
  XOR U4295 ( .A(n2948), .B(key[239]), .Z(n2928) );
  XNOR U4296 ( .A(\w3[0][96] ), .B(\w3[0][104] ), .Z(n2954) );
  XOR U4297 ( .A(\w3[0][119] ), .B(n2954), .Z(n2927) );
  XNOR U4298 ( .A(n2928), .B(n2927), .Z(\w1[1][111] ) );
  XNOR U4299 ( .A(\w3[0][105] ), .B(\w3[0][113] ), .Z(n3289) );
  XNOR U4300 ( .A(n3289), .B(key[240]), .Z(n2930) );
  XNOR U4301 ( .A(n2966), .B(n2954), .Z(n2929) );
  XNOR U4302 ( .A(n2930), .B(n2929), .Z(\w1[1][112] ) );
  XNOR U4303 ( .A(\w3[0][106] ), .B(\w3[0][114] ), .Z(n3293) );
  XNOR U4304 ( .A(n3293), .B(key[241]), .Z(n2932) );
  XOR U4305 ( .A(\w3[0][105] ), .B(n3285), .Z(n2931) );
  XNOR U4306 ( .A(n2932), .B(n2931), .Z(\w1[1][113] ) );
  XNOR U4307 ( .A(\w3[0][107] ), .B(\w3[0][115] ), .Z(n2968) );
  XNOR U4308 ( .A(n2968), .B(key[242]), .Z(n2934) );
  XNOR U4309 ( .A(\w3[0][106] ), .B(n3290), .Z(n2933) );
  XNOR U4310 ( .A(n2934), .B(n2933), .Z(\w1[1][114] ) );
  XOR U4311 ( .A(\w3[0][116] ), .B(n2958), .Z(n2969) );
  XNOR U4312 ( .A(n2969), .B(key[243]), .Z(n2937) );
  XOR U4313 ( .A(\w3[0][107] ), .B(n2935), .Z(n2936) );
  XNOR U4314 ( .A(n2937), .B(n2936), .Z(\w1[1][115] ) );
  XOR U4315 ( .A(\w3[0][117] ), .B(n2958), .Z(n2972) );
  XNOR U4316 ( .A(n2972), .B(key[244]), .Z(n2940) );
  XOR U4317 ( .A(\w3[0][108] ), .B(n2938), .Z(n2939) );
  XNOR U4318 ( .A(n2940), .B(n2939), .Z(\w1[1][116] ) );
  XNOR U4319 ( .A(n2941), .B(key[245]), .Z(n2944) );
  XOR U4320 ( .A(\w3[0][109] ), .B(n2942), .Z(n2943) );
  XNOR U4321 ( .A(n2944), .B(n2943), .Z(\w1[1][117] ) );
  XOR U4322 ( .A(\w3[0][119] ), .B(n2958), .Z(n2981) );
  XNOR U4323 ( .A(n2981), .B(key[246]), .Z(n2947) );
  XOR U4324 ( .A(\w3[0][110] ), .B(n2945), .Z(n2946) );
  XNOR U4325 ( .A(n2947), .B(n2946), .Z(\w1[1][118] ) );
  XOR U4326 ( .A(n2948), .B(key[247]), .Z(n2951) );
  XNOR U4327 ( .A(\w3[0][112] ), .B(n2949), .Z(n2950) );
  XNOR U4328 ( .A(n2951), .B(n2950), .Z(\w1[1][119] ) );
  XNOR U4329 ( .A(\w3[0][3] ), .B(\w3[0][27] ), .Z(n3048) );
  XNOR U4330 ( .A(n3005), .B(key[139]), .Z(n2953) );
  XNOR U4331 ( .A(\w3[0][0] ), .B(\w3[0][4] ), .Z(n3077) );
  XOR U4332 ( .A(\w3[0][19] ), .B(n3077), .Z(n2952) );
  XNOR U4333 ( .A(n2953), .B(n2952), .Z(\w1[1][11] ) );
  XNOR U4334 ( .A(n2954), .B(key[248]), .Z(n2956) );
  XNOR U4335 ( .A(\w3[0][121] ), .B(\w3[0][113] ), .Z(n2955) );
  XNOR U4336 ( .A(n2956), .B(n2955), .Z(n2957) );
  XNOR U4337 ( .A(n2958), .B(n2957), .Z(\w1[1][120] ) );
  XNOR U4338 ( .A(n3289), .B(key[249]), .Z(n2960) );
  XNOR U4339 ( .A(\w3[0][122] ), .B(\w3[0][114] ), .Z(n2959) );
  XNOR U4340 ( .A(n2960), .B(n2959), .Z(n2961) );
  XNOR U4341 ( .A(n2962), .B(n2961), .Z(\w1[1][121] ) );
  XNOR U4342 ( .A(n3293), .B(key[250]), .Z(n2964) );
  XNOR U4343 ( .A(\w3[0][115] ), .B(\w3[0][123] ), .Z(n2963) );
  XNOR U4344 ( .A(n2964), .B(n2963), .Z(n2965) );
  XOR U4345 ( .A(\w3[0][98] ), .B(n2965), .Z(\w1[1][122] ) );
  XOR U4346 ( .A(\w3[0][124] ), .B(n2966), .Z(n2967) );
  XOR U4347 ( .A(n2968), .B(n2967), .Z(n3297) );
  XOR U4348 ( .A(n3297), .B(key[251]), .Z(n2971) );
  XOR U4349 ( .A(\w3[0][99] ), .B(n2969), .Z(n2970) );
  XNOR U4350 ( .A(n2971), .B(n2970), .Z(\w1[1][123] ) );
  XNOR U4351 ( .A(n2972), .B(key[252]), .Z(n2976) );
  XNOR U4352 ( .A(n2974), .B(n2973), .Z(n2975) );
  XNOR U4353 ( .A(n2976), .B(n2975), .Z(\w1[1][124] ) );
  XOR U4354 ( .A(\w3[0][118] ), .B(key[253]), .Z(n2979) );
  XOR U4355 ( .A(n2977), .B(\w3[0][126] ), .Z(n2978) );
  XNOR U4356 ( .A(n2979), .B(n2978), .Z(n2980) );
  XOR U4357 ( .A(\w3[0][101] ), .B(n2980), .Z(\w1[1][125] ) );
  XNOR U4358 ( .A(n2981), .B(key[254]), .Z(n2984) );
  XOR U4359 ( .A(\w3[0][102] ), .B(n2982), .Z(n2983) );
  XNOR U4360 ( .A(n2984), .B(n2983), .Z(\w1[1][126] ) );
  XNOR U4361 ( .A(n3286), .B(key[255]), .Z(n2987) );
  XOR U4362 ( .A(\w3[0][103] ), .B(n2985), .Z(n2986) );
  XNOR U4363 ( .A(n2987), .B(n2986), .Z(\w1[1][127] ) );
  XOR U4364 ( .A(\w3[0][13] ), .B(\w3[0][28] ), .Z(n2989) );
  XNOR U4365 ( .A(\w3[0][8] ), .B(\w3[0][4] ), .Z(n2988) );
  XOR U4366 ( .A(n2989), .B(n2988), .Z(n3009) );
  XNOR U4367 ( .A(n3009), .B(key[140]), .Z(n2991) );
  XNOR U4368 ( .A(\w3[0][0] ), .B(\w3[0][5] ), .Z(n3112) );
  XOR U4369 ( .A(\w3[0][20] ), .B(n3112), .Z(n2990) );
  XNOR U4370 ( .A(n2991), .B(n2990), .Z(\w1[1][12] ) );
  IV U4371 ( .A(\w3[0][21] ), .Z(n3042) );
  XNOR U4372 ( .A(\w3[0][14] ), .B(n3042), .Z(n2993) );
  XNOR U4373 ( .A(\w3[0][5] ), .B(\w3[0][29] ), .Z(n3012) );
  XOR U4374 ( .A(n3012), .B(key[141]), .Z(n2992) );
  XNOR U4375 ( .A(n2993), .B(n2992), .Z(n2994) );
  XOR U4376 ( .A(\w3[0][6] ), .B(n2994), .Z(\w1[1][13] ) );
  IV U4377 ( .A(\w3[0][30] ), .Z(n3187) );
  XOR U4378 ( .A(\w3[0][6] ), .B(n3187), .Z(n3152) );
  XOR U4379 ( .A(\w3[0][8] ), .B(\w3[0][15] ), .Z(n3015) );
  XNOR U4380 ( .A(n3152), .B(n3015), .Z(n3013) );
  XOR U4381 ( .A(n3013), .B(key[142]), .Z(n2996) );
  XNOR U4382 ( .A(\w3[0][0] ), .B(\w3[0][7] ), .Z(n3188) );
  XOR U4383 ( .A(\w3[0][22] ), .B(n3188), .Z(n2995) );
  XNOR U4384 ( .A(n2996), .B(n2995), .Z(\w1[1][14] ) );
  XNOR U4385 ( .A(\w3[0][7] ), .B(\w3[0][31] ), .Z(n3014) );
  XNOR U4386 ( .A(n3014), .B(key[143]), .Z(n2998) );
  XOR U4387 ( .A(\w3[0][8] ), .B(\w3[0][0] ), .Z(n3019) );
  XNOR U4388 ( .A(\w3[0][23] ), .B(n3019), .Z(n2997) );
  XNOR U4389 ( .A(n2998), .B(n2997), .Z(\w1[1][15] ) );
  IV U4390 ( .A(\w3[0][9] ), .Z(n3256) );
  XOR U4391 ( .A(\w3[0][17] ), .B(n3256), .Z(n3023) );
  XNOR U4392 ( .A(n3023), .B(key[144]), .Z(n3000) );
  XNOR U4393 ( .A(\w3[0][24] ), .B(n3019), .Z(n2999) );
  XNOR U4394 ( .A(n3000), .B(n2999), .Z(\w1[1][16] ) );
  XNOR U4395 ( .A(\w3[0][18] ), .B(\w3[0][10] ), .Z(n3047) );
  XNOR U4396 ( .A(n3047), .B(key[145]), .Z(n3002) );
  XNOR U4397 ( .A(n3305), .B(n3256), .Z(n3001) );
  XNOR U4398 ( .A(n3002), .B(n3001), .Z(\w1[1][17] ) );
  IV U4399 ( .A(\w3[0][19] ), .Z(n3028) );
  XOR U4400 ( .A(\w3[0][11] ), .B(n3028), .Z(n3033) );
  XNOR U4401 ( .A(n3033), .B(key[146]), .Z(n3004) );
  XOR U4402 ( .A(n3006), .B(\w3[0][10] ), .Z(n3003) );
  XNOR U4403 ( .A(n3004), .B(n3003), .Z(\w1[1][18] ) );
  IV U4404 ( .A(\w3[0][16] ), .Z(n3020) );
  XOR U4405 ( .A(n3020), .B(\w3[0][20] ), .Z(n3034) );
  IV U4406 ( .A(\w3[0][17] ), .Z(n3301) );
  XOR U4407 ( .A(\w3[0][25] ), .B(n3301), .Z(n3018) );
  XNOR U4408 ( .A(n3018), .B(key[129]), .Z(n3008) );
  XNOR U4409 ( .A(n3006), .B(n3256), .Z(n3007) );
  XNOR U4410 ( .A(n3008), .B(n3007), .Z(\w1[1][1] ) );
  XOR U4411 ( .A(\w3[0][16] ), .B(n3042), .Z(n3039) );
  XNOR U4412 ( .A(n3039), .B(key[148]), .Z(n3011) );
  XOR U4413 ( .A(\w3[0][12] ), .B(n3009), .Z(n3010) );
  XNOR U4414 ( .A(n3011), .B(n3010), .Z(\w1[1][20] ) );
  IV U4415 ( .A(\w3[0][22] ), .Z(n3043) );
  XOR U4416 ( .A(\w3[0][14] ), .B(n3043), .Z(n3052) );
  XOR U4417 ( .A(n3020), .B(\w3[0][23] ), .Z(n3053) );
  XNOR U4418 ( .A(n3014), .B(key[151]), .Z(n3017) );
  XNOR U4419 ( .A(\w3[0][16] ), .B(n3015), .Z(n3016) );
  XNOR U4420 ( .A(n3017), .B(n3016), .Z(\w1[1][23] ) );
  XNOR U4421 ( .A(n3018), .B(key[152]), .Z(n3022) );
  XOR U4422 ( .A(n3020), .B(n3019), .Z(n3021) );
  XNOR U4423 ( .A(n3022), .B(n3021), .Z(\w1[1][24] ) );
  XNOR U4424 ( .A(n3023), .B(key[153]), .Z(n3025) );
  XNOR U4425 ( .A(\w3[0][1] ), .B(\w3[0][26] ), .Z(n3024) );
  XNOR U4426 ( .A(n3025), .B(n3024), .Z(n3026) );
  XNOR U4427 ( .A(n3027), .B(n3026), .Z(\w1[1][25] ) );
  XNOR U4428 ( .A(n3047), .B(key[154]), .Z(n3030) );
  XOR U4429 ( .A(\w3[0][2] ), .B(n3028), .Z(n3029) );
  XNOR U4430 ( .A(n3030), .B(n3029), .Z(n3031) );
  XOR U4431 ( .A(\w3[0][27] ), .B(n3031), .Z(\w1[1][26] ) );
  XOR U4432 ( .A(n3051), .B(\w3[0][28] ), .Z(n3032) );
  XOR U4433 ( .A(n3033), .B(n3032), .Z(n3076) );
  XOR U4434 ( .A(n3076), .B(key[155]), .Z(n3036) );
  XOR U4435 ( .A(\w3[0][3] ), .B(n3034), .Z(n3035) );
  XNOR U4436 ( .A(n3036), .B(n3035), .Z(\w1[1][27] ) );
  XOR U4437 ( .A(\w3[0][20] ), .B(\w3[0][29] ), .Z(n3038) );
  XOR U4438 ( .A(n3051), .B(\w3[0][12] ), .Z(n3037) );
  XOR U4439 ( .A(n3038), .B(n3037), .Z(n3111) );
  XNOR U4440 ( .A(n3111), .B(key[156]), .Z(n3041) );
  XOR U4441 ( .A(\w3[0][4] ), .B(n3039), .Z(n3040) );
  XNOR U4442 ( .A(n3041), .B(n3040), .Z(\w1[1][28] ) );
  XOR U4443 ( .A(\w3[0][13] ), .B(n3042), .Z(n3151) );
  XNOR U4444 ( .A(n3151), .B(key[157]), .Z(n3045) );
  XNOR U4445 ( .A(n3043), .B(n3187), .Z(n3044) );
  XNOR U4446 ( .A(n3045), .B(n3044), .Z(n3046) );
  XOR U4447 ( .A(\w3[0][5] ), .B(n3046), .Z(\w1[1][29] ) );
  XNOR U4448 ( .A(n3047), .B(key[130]), .Z(n3050) );
  XOR U4449 ( .A(\w3[0][26] ), .B(n3048), .Z(n3049) );
  XNOR U4450 ( .A(n3050), .B(n3049), .Z(\w1[1][2] ) );
  XOR U4451 ( .A(n3051), .B(\w3[0][31] ), .Z(n3223) );
  XNOR U4452 ( .A(n3052), .B(n3223), .Z(n3186) );
  XNOR U4453 ( .A(\w3[0][15] ), .B(\w3[0][23] ), .Z(n3222) );
  XNOR U4454 ( .A(n3222), .B(key[159]), .Z(n3055) );
  XOR U4455 ( .A(n3257), .B(\w3[0][7] ), .Z(n3054) );
  XNOR U4456 ( .A(n3055), .B(n3054), .Z(\w1[1][31] ) );
  XNOR U4457 ( .A(\w3[0][48] ), .B(\w3[0][56] ), .Z(n3168) );
  XNOR U4458 ( .A(\w3[0][33] ), .B(\w3[0][57] ), .Z(n3108) );
  XNOR U4459 ( .A(\w3[0][40] ), .B(key[160]), .Z(n3056) );
  XNOR U4460 ( .A(n3108), .B(n3056), .Z(n3057) );
  XOR U4461 ( .A(n3168), .B(n3057), .Z(\w1[1][32] ) );
  XNOR U4462 ( .A(\w3[0][34] ), .B(\w3[0][58] ), .Z(n3116) );
  XNOR U4463 ( .A(\w3[0][41] ), .B(\w3[0][49] ), .Z(n3138) );
  XOR U4464 ( .A(n3138), .B(key[161]), .Z(n3058) );
  XNOR U4465 ( .A(n3116), .B(n3058), .Z(n3059) );
  XNOR U4466 ( .A(\w3[0][57] ), .B(n3059), .Z(\w1[1][33] ) );
  XNOR U4467 ( .A(n3086), .B(key[162]), .Z(n3061) );
  XNOR U4468 ( .A(\w3[0][42] ), .B(\w3[0][50] ), .Z(n3141) );
  XOR U4469 ( .A(\w3[0][58] ), .B(n3141), .Z(n3060) );
  XNOR U4470 ( .A(n3061), .B(n3060), .Z(\w1[1][34] ) );
  XOR U4471 ( .A(\w3[0][36] ), .B(\w3[0][32] ), .Z(n3088) );
  XOR U4472 ( .A(n3088), .B(key[163]), .Z(n3064) );
  IV U4473 ( .A(\w3[0][51] ), .Z(n3140) );
  XOR U4474 ( .A(\w3[0][43] ), .B(n3140), .Z(n3115) );
  XOR U4475 ( .A(\w3[0][56] ), .B(n3115), .Z(n3062) );
  XNOR U4476 ( .A(\w3[0][60] ), .B(n3062), .Z(n3147) );
  XNOR U4477 ( .A(\w3[0][59] ), .B(n3147), .Z(n3063) );
  XNOR U4478 ( .A(n3064), .B(n3063), .Z(\w1[1][35] ) );
  XOR U4479 ( .A(\w3[0][32] ), .B(\w3[0][37] ), .Z(n3094) );
  XOR U4480 ( .A(\w3[0][52] ), .B(\w3[0][61] ), .Z(n3066) );
  XNOR U4481 ( .A(\w3[0][56] ), .B(\w3[0][44] ), .Z(n3065) );
  XOR U4482 ( .A(n3066), .B(n3065), .Z(n3156) );
  XOR U4483 ( .A(n3156), .B(key[164]), .Z(n3067) );
  XOR U4484 ( .A(n3094), .B(n3067), .Z(n3068) );
  XNOR U4485 ( .A(\w3[0][60] ), .B(n3068), .Z(\w1[1][36] ) );
  XNOR U4486 ( .A(\w3[0][38] ), .B(\w3[0][62] ), .Z(n3100) );
  XNOR U4487 ( .A(n3100), .B(key[165]), .Z(n3070) );
  IV U4488 ( .A(\w3[0][53] ), .Z(n3120) );
  XOR U4489 ( .A(\w3[0][45] ), .B(n3120), .Z(n3159) );
  XOR U4490 ( .A(\w3[0][61] ), .B(n3159), .Z(n3069) );
  XNOR U4491 ( .A(n3070), .B(n3069), .Z(\w1[1][37] ) );
  XOR U4492 ( .A(\w3[0][32] ), .B(\w3[0][39] ), .Z(n3101) );
  XOR U4493 ( .A(n3101), .B(key[166]), .Z(n3072) );
  XNOR U4494 ( .A(\w3[0][56] ), .B(\w3[0][63] ), .Z(n3073) );
  XOR U4495 ( .A(\w3[0][46] ), .B(\w3[0][54] ), .Z(n3125) );
  XOR U4496 ( .A(n3073), .B(n3125), .Z(n3164) );
  XOR U4497 ( .A(\w3[0][62] ), .B(n3164), .Z(n3071) );
  XNOR U4498 ( .A(n3072), .B(n3071), .Z(\w1[1][38] ) );
  XNOR U4499 ( .A(\w3[0][47] ), .B(\w3[0][55] ), .Z(n3167) );
  XNOR U4500 ( .A(n3167), .B(key[167]), .Z(n3075) );
  XOR U4501 ( .A(\w3[0][32] ), .B(n3073), .Z(n3074) );
  XNOR U4502 ( .A(n3075), .B(n3074), .Z(\w1[1][39] ) );
  XOR U4503 ( .A(n3076), .B(key[131]), .Z(n3079) );
  XOR U4504 ( .A(n3077), .B(\w3[0][27] ), .Z(n3078) );
  XNOR U4505 ( .A(n3079), .B(n3078), .Z(\w1[1][3] ) );
  IV U4506 ( .A(\w3[0][33] ), .Z(n3139) );
  XOR U4507 ( .A(\w3[0][42] ), .B(key[169]), .Z(n3081) );
  IV U4508 ( .A(\w3[0][34] ), .Z(n3145) );
  XOR U4509 ( .A(\w3[0][49] ), .B(n3145), .Z(n3080) );
  XNOR U4510 ( .A(n3081), .B(n3080), .Z(n3082) );
  XNOR U4511 ( .A(n3082), .B(n3108), .Z(\w1[1][41] ) );
  XOR U4512 ( .A(\w3[0][43] ), .B(key[170]), .Z(n3084) );
  IV U4513 ( .A(\w3[0][35] ), .Z(n3148) );
  XOR U4514 ( .A(\w3[0][50] ), .B(n3148), .Z(n3083) );
  XNOR U4515 ( .A(n3084), .B(n3083), .Z(n3085) );
  XNOR U4516 ( .A(n3085), .B(n3116), .Z(\w1[1][42] ) );
  IV U4517 ( .A(\w3[0][40] ), .Z(n3091) );
  XNOR U4518 ( .A(n3091), .B(n3086), .Z(n3087) );
  XOR U4519 ( .A(\w3[0][44] ), .B(n3087), .Z(n3119) );
  XNOR U4520 ( .A(n3119), .B(key[171]), .Z(n3090) );
  XNOR U4521 ( .A(\w3[0][51] ), .B(n3088), .Z(n3089) );
  XNOR U4522 ( .A(n3090), .B(n3089), .Z(\w1[1][43] ) );
  XOR U4523 ( .A(\w3[0][36] ), .B(\w3[0][45] ), .Z(n3093) );
  XOR U4524 ( .A(n3091), .B(\w3[0][60] ), .Z(n3092) );
  XOR U4525 ( .A(n3093), .B(n3092), .Z(n3121) );
  XNOR U4526 ( .A(n3121), .B(key[172]), .Z(n3096) );
  XNOR U4527 ( .A(\w3[0][52] ), .B(n3094), .Z(n3095) );
  XNOR U4528 ( .A(n3096), .B(n3095), .Z(\w1[1][44] ) );
  XNOR U4529 ( .A(\w3[0][61] ), .B(\w3[0][37] ), .Z(n3124) );
  XNOR U4530 ( .A(n3124), .B(key[173]), .Z(n3098) );
  XNOR U4531 ( .A(\w3[0][38] ), .B(\w3[0][46] ), .Z(n3097) );
  XNOR U4532 ( .A(n3098), .B(n3097), .Z(n3099) );
  XOR U4533 ( .A(\w3[0][53] ), .B(n3099), .Z(\w1[1][45] ) );
  XOR U4534 ( .A(\w3[0][40] ), .B(\w3[0][47] ), .Z(n3130) );
  XOR U4535 ( .A(n3100), .B(n3130), .Z(n3126) );
  XNOR U4536 ( .A(n3126), .B(key[174]), .Z(n3103) );
  XNOR U4537 ( .A(\w3[0][54] ), .B(n3101), .Z(n3102) );
  XNOR U4538 ( .A(n3103), .B(n3102), .Z(\w1[1][46] ) );
  XOR U4539 ( .A(\w3[0][63] ), .B(\w3[0][39] ), .Z(n3129) );
  XOR U4540 ( .A(n3129), .B(key[175]), .Z(n3105) );
  XNOR U4541 ( .A(\w3[0][40] ), .B(\w3[0][32] ), .Z(n3133) );
  XOR U4542 ( .A(\w3[0][55] ), .B(n3133), .Z(n3104) );
  XNOR U4543 ( .A(n3105), .B(n3104), .Z(\w1[1][47] ) );
  XNOR U4544 ( .A(n3133), .B(key[176]), .Z(n3107) );
  XOR U4545 ( .A(\w3[0][56] ), .B(n3138), .Z(n3106) );
  XNOR U4546 ( .A(n3107), .B(n3106), .Z(\w1[1][48] ) );
  XNOR U4547 ( .A(n3141), .B(key[177]), .Z(n3110) );
  XOR U4548 ( .A(n3108), .B(\w3[0][41] ), .Z(n3109) );
  XNOR U4549 ( .A(n3110), .B(n3109), .Z(\w1[1][49] ) );
  XNOR U4550 ( .A(n3111), .B(key[132]), .Z(n3114) );
  XOR U4551 ( .A(n3112), .B(\w3[0][28] ), .Z(n3113) );
  XNOR U4552 ( .A(n3114), .B(n3113), .Z(\w1[1][4] ) );
  XNOR U4553 ( .A(n3115), .B(key[178]), .Z(n3118) );
  XOR U4554 ( .A(n3116), .B(\w3[0][42] ), .Z(n3117) );
  XNOR U4555 ( .A(n3118), .B(n3117), .Z(\w1[1][50] ) );
  IV U4556 ( .A(\w3[0][48] ), .Z(n3134) );
  XOR U4557 ( .A(n3134), .B(\w3[0][52] ), .Z(n3146) );
  XOR U4558 ( .A(\w3[0][48] ), .B(n3120), .Z(n3155) );
  XNOR U4559 ( .A(n3155), .B(key[180]), .Z(n3123) );
  XOR U4560 ( .A(\w3[0][44] ), .B(n3121), .Z(n3122) );
  XNOR U4561 ( .A(n3123), .B(n3122), .Z(\w1[1][52] ) );
  XOR U4562 ( .A(n3134), .B(\w3[0][55] ), .Z(n3163) );
  XNOR U4563 ( .A(n3163), .B(key[182]), .Z(n3128) );
  XOR U4564 ( .A(\w3[0][46] ), .B(n3126), .Z(n3127) );
  XNOR U4565 ( .A(n3128), .B(n3127), .Z(\w1[1][54] ) );
  XOR U4566 ( .A(n3129), .B(key[183]), .Z(n3132) );
  XNOR U4567 ( .A(\w3[0][48] ), .B(n3130), .Z(n3131) );
  XNOR U4568 ( .A(n3132), .B(n3131), .Z(\w1[1][55] ) );
  XNOR U4569 ( .A(n3133), .B(key[184]), .Z(n3136) );
  XOR U4570 ( .A(n3134), .B(\w3[0][49] ), .Z(n3135) );
  XNOR U4571 ( .A(n3136), .B(n3135), .Z(n3137) );
  XOR U4572 ( .A(\w3[0][57] ), .B(n3137), .Z(\w1[1][56] ) );
  XNOR U4573 ( .A(n3140), .B(key[186]), .Z(n3143) );
  XOR U4574 ( .A(n3141), .B(\w3[0][59] ), .Z(n3142) );
  XNOR U4575 ( .A(n3143), .B(n3142), .Z(n3144) );
  XNOR U4576 ( .A(n3145), .B(n3144), .Z(\w1[1][58] ) );
  XNOR U4577 ( .A(n3146), .B(key[187]), .Z(n3150) );
  XOR U4578 ( .A(n3148), .B(n3147), .Z(n3149) );
  XNOR U4579 ( .A(n3150), .B(n3149), .Z(\w1[1][59] ) );
  XNOR U4580 ( .A(n3151), .B(key[133]), .Z(n3154) );
  XOR U4581 ( .A(\w3[0][29] ), .B(n3152), .Z(n3153) );
  XNOR U4582 ( .A(n3154), .B(n3153), .Z(\w1[1][5] ) );
  XNOR U4583 ( .A(n3155), .B(key[188]), .Z(n3158) );
  XOR U4584 ( .A(\w3[0][36] ), .B(n3156), .Z(n3157) );
  XNOR U4585 ( .A(n3158), .B(n3157), .Z(\w1[1][60] ) );
  XOR U4586 ( .A(\w3[0][54] ), .B(key[189]), .Z(n3161) );
  XOR U4587 ( .A(n3159), .B(\w3[0][62] ), .Z(n3160) );
  XNOR U4588 ( .A(n3161), .B(n3160), .Z(n3162) );
  XOR U4589 ( .A(\w3[0][37] ), .B(n3162), .Z(\w1[1][61] ) );
  XNOR U4590 ( .A(n3163), .B(key[190]), .Z(n3166) );
  XOR U4591 ( .A(\w3[0][38] ), .B(n3164), .Z(n3165) );
  XNOR U4592 ( .A(n3166), .B(n3165), .Z(\w1[1][62] ) );
  XNOR U4593 ( .A(n3167), .B(key[191]), .Z(n3170) );
  XOR U4594 ( .A(n3168), .B(\w3[0][39] ), .Z(n3169) );
  XNOR U4595 ( .A(n3170), .B(n3169), .Z(\w1[1][63] ) );
  XNOR U4596 ( .A(\w3[0][80] ), .B(\w3[0][88] ), .Z(n3282) );
  XNOR U4597 ( .A(\w3[0][65] ), .B(\w3[0][89] ), .Z(n3228) );
  XNOR U4598 ( .A(\w3[0][72] ), .B(key[192]), .Z(n3171) );
  XNOR U4599 ( .A(n3228), .B(n3171), .Z(n3172) );
  XOR U4600 ( .A(n3282), .B(n3172), .Z(\w1[1][64] ) );
  XNOR U4601 ( .A(\w3[0][66] ), .B(\w3[0][90] ), .Z(n3232) );
  XNOR U4602 ( .A(\w3[0][73] ), .B(\w3[0][81] ), .Z(n3254) );
  XOR U4603 ( .A(n3254), .B(key[193]), .Z(n3173) );
  XNOR U4604 ( .A(n3232), .B(n3173), .Z(n3174) );
  XNOR U4605 ( .A(\w3[0][89] ), .B(n3174), .Z(\w1[1][65] ) );
  XNOR U4606 ( .A(n3202), .B(key[194]), .Z(n3176) );
  XNOR U4607 ( .A(\w3[0][74] ), .B(\w3[0][82] ), .Z(n3259) );
  XOR U4608 ( .A(\w3[0][90] ), .B(n3259), .Z(n3175) );
  XNOR U4609 ( .A(n3176), .B(n3175), .Z(\w1[1][66] ) );
  XOR U4610 ( .A(\w3[0][68] ), .B(\w3[0][64] ), .Z(n3204) );
  XOR U4611 ( .A(n3204), .B(key[195]), .Z(n3179) );
  IV U4612 ( .A(\w3[0][83] ), .Z(n3258) );
  XOR U4613 ( .A(\w3[0][75] ), .B(n3258), .Z(n3231) );
  XOR U4614 ( .A(\w3[0][88] ), .B(n3231), .Z(n3177) );
  XNOR U4615 ( .A(\w3[0][92] ), .B(n3177), .Z(n3265) );
  XNOR U4616 ( .A(\w3[0][91] ), .B(n3265), .Z(n3178) );
  XNOR U4617 ( .A(n3179), .B(n3178), .Z(\w1[1][67] ) );
  XOR U4618 ( .A(\w3[0][64] ), .B(\w3[0][69] ), .Z(n3210) );
  XOR U4619 ( .A(\w3[0][84] ), .B(\w3[0][93] ), .Z(n3181) );
  XNOR U4620 ( .A(\w3[0][88] ), .B(\w3[0][76] ), .Z(n3180) );
  XOR U4621 ( .A(n3181), .B(n3180), .Z(n3270) );
  XOR U4622 ( .A(n3270), .B(key[196]), .Z(n3182) );
  XOR U4623 ( .A(n3210), .B(n3182), .Z(n3183) );
  XNOR U4624 ( .A(\w3[0][92] ), .B(n3183), .Z(\w1[1][68] ) );
  XNOR U4625 ( .A(\w3[0][70] ), .B(\w3[0][94] ), .Z(n3216) );
  XNOR U4626 ( .A(n3216), .B(key[197]), .Z(n3185) );
  IV U4627 ( .A(\w3[0][85] ), .Z(n3236) );
  XOR U4628 ( .A(\w3[0][77] ), .B(n3236), .Z(n3273) );
  XOR U4629 ( .A(\w3[0][93] ), .B(n3273), .Z(n3184) );
  XNOR U4630 ( .A(n3185), .B(n3184), .Z(\w1[1][69] ) );
  XNOR U4631 ( .A(n3186), .B(key[134]), .Z(n3190) );
  XNOR U4632 ( .A(n3188), .B(n3187), .Z(n3189) );
  XNOR U4633 ( .A(n3190), .B(n3189), .Z(\w1[1][6] ) );
  XOR U4634 ( .A(\w3[0][64] ), .B(\w3[0][71] ), .Z(n3217) );
  XOR U4635 ( .A(n3217), .B(key[198]), .Z(n3192) );
  XNOR U4636 ( .A(\w3[0][78] ), .B(\w3[0][86] ), .Z(n3241) );
  XOR U4637 ( .A(\w3[0][88] ), .B(\w3[0][95] ), .Z(n3193) );
  XOR U4638 ( .A(n3241), .B(n3193), .Z(n3278) );
  XOR U4639 ( .A(\w3[0][94] ), .B(n3278), .Z(n3191) );
  XNOR U4640 ( .A(n3192), .B(n3191), .Z(\w1[1][70] ) );
  XNOR U4641 ( .A(\w3[0][79] ), .B(\w3[0][87] ), .Z(n3281) );
  XNOR U4642 ( .A(n3281), .B(key[199]), .Z(n3195) );
  XNOR U4643 ( .A(\w3[0][64] ), .B(n3193), .Z(n3194) );
  XNOR U4644 ( .A(n3195), .B(n3194), .Z(\w1[1][71] ) );
  IV U4645 ( .A(\w3[0][65] ), .Z(n3255) );
  XOR U4646 ( .A(\w3[0][74] ), .B(key[201]), .Z(n3197) );
  IV U4647 ( .A(\w3[0][66] ), .Z(n3263) );
  XOR U4648 ( .A(\w3[0][81] ), .B(n3263), .Z(n3196) );
  XNOR U4649 ( .A(n3197), .B(n3196), .Z(n3198) );
  XNOR U4650 ( .A(n3198), .B(n3228), .Z(\w1[1][73] ) );
  XOR U4651 ( .A(\w3[0][75] ), .B(key[202]), .Z(n3200) );
  IV U4652 ( .A(\w3[0][67] ), .Z(n3266) );
  XOR U4653 ( .A(\w3[0][82] ), .B(n3266), .Z(n3199) );
  XNOR U4654 ( .A(n3200), .B(n3199), .Z(n3201) );
  XNOR U4655 ( .A(n3201), .B(n3232), .Z(\w1[1][74] ) );
  IV U4656 ( .A(\w3[0][72] ), .Z(n3207) );
  XNOR U4657 ( .A(n3207), .B(n3202), .Z(n3203) );
  XOR U4658 ( .A(\w3[0][76] ), .B(n3203), .Z(n3235) );
  XNOR U4659 ( .A(n3235), .B(key[203]), .Z(n3206) );
  XNOR U4660 ( .A(\w3[0][83] ), .B(n3204), .Z(n3205) );
  XNOR U4661 ( .A(n3206), .B(n3205), .Z(\w1[1][75] ) );
  XOR U4662 ( .A(\w3[0][68] ), .B(\w3[0][77] ), .Z(n3209) );
  XOR U4663 ( .A(n3207), .B(\w3[0][92] ), .Z(n3208) );
  XOR U4664 ( .A(n3209), .B(n3208), .Z(n3237) );
  XNOR U4665 ( .A(n3237), .B(key[204]), .Z(n3212) );
  XNOR U4666 ( .A(\w3[0][84] ), .B(n3210), .Z(n3211) );
  XNOR U4667 ( .A(n3212), .B(n3211), .Z(\w1[1][76] ) );
  XNOR U4668 ( .A(\w3[0][93] ), .B(\w3[0][69] ), .Z(n3240) );
  XNOR U4669 ( .A(n3240), .B(key[205]), .Z(n3214) );
  XNOR U4670 ( .A(\w3[0][70] ), .B(\w3[0][78] ), .Z(n3213) );
  XNOR U4671 ( .A(n3214), .B(n3213), .Z(n3215) );
  XOR U4672 ( .A(\w3[0][85] ), .B(n3215), .Z(\w1[1][77] ) );
  XOR U4673 ( .A(\w3[0][72] ), .B(\w3[0][79] ), .Z(n3246) );
  XOR U4674 ( .A(n3216), .B(n3246), .Z(n3242) );
  XNOR U4675 ( .A(n3242), .B(key[206]), .Z(n3219) );
  XNOR U4676 ( .A(\w3[0][86] ), .B(n3217), .Z(n3218) );
  XNOR U4677 ( .A(n3219), .B(n3218), .Z(\w1[1][78] ) );
  XOR U4678 ( .A(\w3[0][95] ), .B(\w3[0][71] ), .Z(n3245) );
  XOR U4679 ( .A(n3245), .B(key[207]), .Z(n3221) );
  XNOR U4680 ( .A(\w3[0][72] ), .B(\w3[0][64] ), .Z(n3249) );
  XOR U4681 ( .A(\w3[0][87] ), .B(n3249), .Z(n3220) );
  XNOR U4682 ( .A(n3221), .B(n3220), .Z(\w1[1][79] ) );
  XNOR U4683 ( .A(n3222), .B(key[135]), .Z(n3225) );
  XOR U4684 ( .A(\w3[0][0] ), .B(n3223), .Z(n3224) );
  XNOR U4685 ( .A(n3225), .B(n3224), .Z(\w1[1][7] ) );
  XNOR U4686 ( .A(n3249), .B(key[208]), .Z(n3227) );
  XOR U4687 ( .A(\w3[0][88] ), .B(n3254), .Z(n3226) );
  XNOR U4688 ( .A(n3227), .B(n3226), .Z(\w1[1][80] ) );
  XNOR U4689 ( .A(n3259), .B(key[209]), .Z(n3230) );
  XOR U4690 ( .A(n3228), .B(\w3[0][73] ), .Z(n3229) );
  XNOR U4691 ( .A(n3230), .B(n3229), .Z(\w1[1][81] ) );
  XNOR U4692 ( .A(n3231), .B(key[210]), .Z(n3234) );
  XOR U4693 ( .A(n3232), .B(\w3[0][74] ), .Z(n3233) );
  XNOR U4694 ( .A(n3234), .B(n3233), .Z(\w1[1][82] ) );
  IV U4695 ( .A(\w3[0][80] ), .Z(n3250) );
  XOR U4696 ( .A(n3250), .B(\w3[0][84] ), .Z(n3264) );
  XOR U4697 ( .A(\w3[0][80] ), .B(n3236), .Z(n3269) );
  XNOR U4698 ( .A(n3269), .B(key[212]), .Z(n3239) );
  XOR U4699 ( .A(\w3[0][76] ), .B(n3237), .Z(n3238) );
  XNOR U4700 ( .A(n3239), .B(n3238), .Z(\w1[1][84] ) );
  XOR U4701 ( .A(n3250), .B(\w3[0][87] ), .Z(n3277) );
  XNOR U4702 ( .A(n3277), .B(key[214]), .Z(n3244) );
  XOR U4703 ( .A(\w3[0][78] ), .B(n3242), .Z(n3243) );
  XNOR U4704 ( .A(n3244), .B(n3243), .Z(\w1[1][86] ) );
  XOR U4705 ( .A(n3245), .B(key[215]), .Z(n3248) );
  XNOR U4706 ( .A(\w3[0][80] ), .B(n3246), .Z(n3247) );
  XNOR U4707 ( .A(n3248), .B(n3247), .Z(\w1[1][87] ) );
  XNOR U4708 ( .A(n3249), .B(key[216]), .Z(n3252) );
  XOR U4709 ( .A(n3250), .B(\w3[0][81] ), .Z(n3251) );
  XNOR U4710 ( .A(n3252), .B(n3251), .Z(n3253) );
  XOR U4711 ( .A(\w3[0][89] ), .B(n3253), .Z(\w1[1][88] ) );
  XNOR U4712 ( .A(n3258), .B(key[218]), .Z(n3261) );
  XOR U4713 ( .A(n3259), .B(\w3[0][91] ), .Z(n3260) );
  XNOR U4714 ( .A(n3261), .B(n3260), .Z(n3262) );
  XNOR U4715 ( .A(n3263), .B(n3262), .Z(\w1[1][90] ) );
  XNOR U4716 ( .A(n3264), .B(key[219]), .Z(n3268) );
  XOR U4717 ( .A(n3266), .B(n3265), .Z(n3267) );
  XNOR U4718 ( .A(n3268), .B(n3267), .Z(\w1[1][91] ) );
  XNOR U4719 ( .A(n3269), .B(key[220]), .Z(n3272) );
  XOR U4720 ( .A(\w3[0][68] ), .B(n3270), .Z(n3271) );
  XNOR U4721 ( .A(n3272), .B(n3271), .Z(\w1[1][92] ) );
  XOR U4722 ( .A(\w3[0][86] ), .B(key[221]), .Z(n3275) );
  XOR U4723 ( .A(n3273), .B(\w3[0][94] ), .Z(n3274) );
  XNOR U4724 ( .A(n3275), .B(n3274), .Z(n3276) );
  XOR U4725 ( .A(\w3[0][69] ), .B(n3276), .Z(\w1[1][93] ) );
  XNOR U4726 ( .A(n3277), .B(key[222]), .Z(n3280) );
  XOR U4727 ( .A(\w3[0][70] ), .B(n3278), .Z(n3279) );
  XNOR U4728 ( .A(n3280), .B(n3279), .Z(\w1[1][94] ) );
  XNOR U4729 ( .A(n3281), .B(key[223]), .Z(n3284) );
  XOR U4730 ( .A(n3282), .B(\w3[0][71] ), .Z(n3283) );
  XNOR U4731 ( .A(n3284), .B(n3283), .Z(\w1[1][95] ) );
  XOR U4732 ( .A(\w3[0][104] ), .B(key[224]), .Z(n3288) );
  XNOR U4733 ( .A(n3286), .B(n3285), .Z(n3287) );
  XNOR U4734 ( .A(n3288), .B(n3287), .Z(\w1[1][96] ) );
  XNOR U4735 ( .A(n3289), .B(key[225]), .Z(n3292) );
  XNOR U4736 ( .A(\w3[0][121] ), .B(n3290), .Z(n3291) );
  XNOR U4737 ( .A(n3292), .B(n3291), .Z(\w1[1][97] ) );
  XNOR U4738 ( .A(n3293), .B(key[226]), .Z(n3296) );
  XOR U4739 ( .A(\w3[0][122] ), .B(n3294), .Z(n3295) );
  XNOR U4740 ( .A(n3296), .B(n3295), .Z(\w1[1][98] ) );
  XOR U4741 ( .A(n3297), .B(key[227]), .Z(n3300) );
  XOR U4742 ( .A(n3298), .B(\w3[0][123] ), .Z(n3299) );
  XNOR U4743 ( .A(n3300), .B(n3299), .Z(\w1[1][99] ) );
  XOR U4744 ( .A(\w3[0][10] ), .B(key[137]), .Z(n3303) );
  XOR U4745 ( .A(\w3[0][2] ), .B(n3301), .Z(n3302) );
  XNOR U4746 ( .A(n3303), .B(n3302), .Z(n3304) );
  XNOR U4747 ( .A(n3305), .B(n3304), .Z(\w1[1][9] ) );
  XNOR U4748 ( .A(\w3[1][1] ), .B(\w3[1][25] ), .Z(n3721) );
  IV U4749 ( .A(\w3[1][24] ), .Z(n3464) );
  XOR U4750 ( .A(\w3[1][16] ), .B(n3464), .Z(n3673) );
  XNOR U4751 ( .A(\w3[1][8] ), .B(key[256]), .Z(n3306) );
  XNOR U4752 ( .A(n3673), .B(n3306), .Z(n3307) );
  XOR U4753 ( .A(n3721), .B(n3307), .Z(\w1[2][0] ) );
  XOR U4754 ( .A(\w3[1][96] ), .B(\w3[1][101] ), .Z(n3329) );
  XOR U4755 ( .A(\w3[1][116] ), .B(\w3[1][125] ), .Z(n3309) );
  IV U4756 ( .A(\w3[1][120] ), .Z(n3382) );
  XOR U4757 ( .A(n3382), .B(\w3[1][108] ), .Z(n3308) );
  XOR U4758 ( .A(n3309), .B(n3308), .Z(n3390) );
  XOR U4759 ( .A(n3390), .B(key[356]), .Z(n3310) );
  XOR U4760 ( .A(n3329), .B(n3310), .Z(n3311) );
  XNOR U4761 ( .A(\w3[1][124] ), .B(n3311), .Z(\w1[2][100] ) );
  XNOR U4762 ( .A(\w3[1][102] ), .B(\w3[1][126] ), .Z(n3338) );
  XNOR U4763 ( .A(n3338), .B(key[357]), .Z(n3313) );
  XNOR U4764 ( .A(\w3[1][109] ), .B(\w3[1][117] ), .Z(n3393) );
  XOR U4765 ( .A(\w3[1][125] ), .B(n3393), .Z(n3312) );
  XNOR U4766 ( .A(n3313), .B(n3312), .Z(\w1[2][101] ) );
  XOR U4767 ( .A(\w3[1][96] ), .B(\w3[1][103] ), .Z(n3339) );
  XOR U4768 ( .A(n3339), .B(key[358]), .Z(n3315) );
  XOR U4769 ( .A(n3382), .B(\w3[1][127] ), .Z(n3316) );
  XOR U4770 ( .A(\w3[1][110] ), .B(\w3[1][118] ), .Z(n3357) );
  XOR U4771 ( .A(n3316), .B(n3357), .Z(n3398) );
  XOR U4772 ( .A(\w3[1][126] ), .B(n3398), .Z(n3314) );
  XNOR U4773 ( .A(n3315), .B(n3314), .Z(\w1[2][102] ) );
  XNOR U4774 ( .A(\w3[1][111] ), .B(\w3[1][119] ), .Z(n3401) );
  XNOR U4775 ( .A(n3401), .B(key[359]), .Z(n3318) );
  XOR U4776 ( .A(\w3[1][96] ), .B(n3316), .Z(n3317) );
  XNOR U4777 ( .A(n3318), .B(n3317), .Z(\w1[2][103] ) );
  IV U4778 ( .A(\w3[1][97] ), .Z(n3377) );
  IV U4779 ( .A(\w3[1][112] ), .Z(n3373) );
  XOR U4780 ( .A(\w3[1][120] ), .B(n3373), .Z(n3702) );
  XOR U4781 ( .A(\w3[1][106] ), .B(\w3[1][98] ), .Z(n3380) );
  XNOR U4782 ( .A(\w3[1][97] ), .B(\w3[1][121] ), .Z(n3701) );
  XOR U4783 ( .A(n3701), .B(key[361]), .Z(n3319) );
  XOR U4784 ( .A(n3380), .B(n3319), .Z(n3320) );
  XNOR U4785 ( .A(\w3[1][113] ), .B(n3320), .Z(\w1[2][105] ) );
  XOR U4786 ( .A(\w3[1][107] ), .B(\w3[1][99] ), .Z(n3322) );
  XNOR U4787 ( .A(\w3[1][98] ), .B(\w3[1][122] ), .Z(n3706) );
  XOR U4788 ( .A(n3706), .B(key[362]), .Z(n3321) );
  XNOR U4789 ( .A(n3322), .B(n3321), .Z(n3323) );
  XOR U4790 ( .A(\w3[1][114] ), .B(n3323), .Z(\w1[2][106] ) );
  XNOR U4791 ( .A(\w3[1][99] ), .B(\w3[1][123] ), .Z(n3710) );
  XOR U4792 ( .A(\w3[1][108] ), .B(n3710), .Z(n3324) );
  XOR U4793 ( .A(\w3[1][104] ), .B(n3324), .Z(n3350) );
  XNOR U4794 ( .A(n3350), .B(key[363]), .Z(n3326) );
  IV U4795 ( .A(\w3[1][100] ), .Z(n3389) );
  XOR U4796 ( .A(\w3[1][96] ), .B(n3389), .Z(n3714) );
  XOR U4797 ( .A(\w3[1][115] ), .B(n3714), .Z(n3325) );
  XNOR U4798 ( .A(n3326), .B(n3325), .Z(\w1[2][107] ) );
  XOR U4799 ( .A(\w3[1][100] ), .B(\w3[1][104] ), .Z(n3328) );
  XNOR U4800 ( .A(\w3[1][124] ), .B(\w3[1][109] ), .Z(n3327) );
  XOR U4801 ( .A(n3328), .B(n3327), .Z(n3353) );
  XNOR U4802 ( .A(n3353), .B(key[364]), .Z(n3331) );
  XNOR U4803 ( .A(\w3[1][116] ), .B(n3329), .Z(n3330) );
  XNOR U4804 ( .A(n3331), .B(n3330), .Z(\w1[2][108] ) );
  XNOR U4805 ( .A(\w3[1][125] ), .B(\w3[1][101] ), .Z(n3356) );
  XNOR U4806 ( .A(n3356), .B(key[365]), .Z(n3333) );
  XNOR U4807 ( .A(\w3[1][102] ), .B(\w3[1][110] ), .Z(n3332) );
  XNOR U4808 ( .A(n3333), .B(n3332), .Z(n3334) );
  XOR U4809 ( .A(\w3[1][117] ), .B(n3334), .Z(\w1[2][109] ) );
  XOR U4810 ( .A(\w3[1][11] ), .B(\w3[1][3] ), .Z(n3336) );
  XNOR U4811 ( .A(\w3[1][2] ), .B(\w3[1][26] ), .Z(n3424) );
  XOR U4812 ( .A(n3424), .B(key[266]), .Z(n3335) );
  XNOR U4813 ( .A(n3336), .B(n3335), .Z(n3337) );
  XOR U4814 ( .A(\w3[1][18] ), .B(n3337), .Z(\w1[2][10] ) );
  XOR U4815 ( .A(\w3[1][111] ), .B(\w3[1][104] ), .Z(n3364) );
  XOR U4816 ( .A(n3338), .B(n3364), .Z(n3360) );
  XNOR U4817 ( .A(n3360), .B(key[366]), .Z(n3341) );
  XNOR U4818 ( .A(\w3[1][118] ), .B(n3339), .Z(n3340) );
  XNOR U4819 ( .A(n3341), .B(n3340), .Z(\w1[2][110] ) );
  XOR U4820 ( .A(\w3[1][127] ), .B(\w3[1][103] ), .Z(n3363) );
  XOR U4821 ( .A(n3363), .B(key[367]), .Z(n3343) );
  XNOR U4822 ( .A(\w3[1][96] ), .B(\w3[1][104] ), .Z(n3369) );
  XOR U4823 ( .A(\w3[1][119] ), .B(n3369), .Z(n3342) );
  XNOR U4824 ( .A(n3343), .B(n3342), .Z(\w1[2][111] ) );
  XNOR U4825 ( .A(\w3[1][105] ), .B(\w3[1][113] ), .Z(n3705) );
  XNOR U4826 ( .A(n3705), .B(key[368]), .Z(n3345) );
  XNOR U4827 ( .A(n3382), .B(n3369), .Z(n3344) );
  XNOR U4828 ( .A(n3345), .B(n3344), .Z(\w1[2][112] ) );
  XNOR U4829 ( .A(\w3[1][106] ), .B(\w3[1][114] ), .Z(n3709) );
  XNOR U4830 ( .A(n3709), .B(key[369]), .Z(n3347) );
  XOR U4831 ( .A(\w3[1][105] ), .B(n3701), .Z(n3346) );
  XNOR U4832 ( .A(n3347), .B(n3346), .Z(\w1[2][113] ) );
  XNOR U4833 ( .A(\w3[1][107] ), .B(\w3[1][115] ), .Z(n3384) );
  XNOR U4834 ( .A(n3384), .B(key[370]), .Z(n3349) );
  XNOR U4835 ( .A(n3380), .B(\w3[1][122] ), .Z(n3348) );
  XNOR U4836 ( .A(n3349), .B(n3348), .Z(\w1[2][114] ) );
  XOR U4837 ( .A(\w3[1][116] ), .B(n3373), .Z(n3385) );
  XNOR U4838 ( .A(n3385), .B(key[371]), .Z(n3352) );
  XOR U4839 ( .A(\w3[1][107] ), .B(n3350), .Z(n3351) );
  XNOR U4840 ( .A(n3352), .B(n3351), .Z(\w1[2][115] ) );
  XOR U4841 ( .A(\w3[1][117] ), .B(n3373), .Z(n3388) );
  XNOR U4842 ( .A(n3388), .B(key[372]), .Z(n3355) );
  XOR U4843 ( .A(\w3[1][108] ), .B(n3353), .Z(n3354) );
  XNOR U4844 ( .A(n3355), .B(n3354), .Z(\w1[2][116] ) );
  XNOR U4845 ( .A(n3356), .B(key[373]), .Z(n3359) );
  XNOR U4846 ( .A(\w3[1][109] ), .B(n3357), .Z(n3358) );
  XNOR U4847 ( .A(n3359), .B(n3358), .Z(\w1[2][117] ) );
  XOR U4848 ( .A(\w3[1][119] ), .B(n3373), .Z(n3397) );
  XNOR U4849 ( .A(n3397), .B(key[374]), .Z(n3362) );
  XOR U4850 ( .A(\w3[1][110] ), .B(n3360), .Z(n3361) );
  XNOR U4851 ( .A(n3362), .B(n3361), .Z(\w1[2][118] ) );
  XOR U4852 ( .A(n3363), .B(key[375]), .Z(n3366) );
  XNOR U4853 ( .A(\w3[1][112] ), .B(n3364), .Z(n3365) );
  XNOR U4854 ( .A(n3366), .B(n3365), .Z(\w1[2][119] ) );
  XNOR U4855 ( .A(\w3[1][3] ), .B(\w3[1][27] ), .Z(n3461) );
  XNOR U4856 ( .A(n3421), .B(key[267]), .Z(n3368) );
  XNOR U4857 ( .A(\w3[1][0] ), .B(\w3[1][4] ), .Z(n3493) );
  XOR U4858 ( .A(\w3[1][19] ), .B(n3493), .Z(n3367) );
  XNOR U4859 ( .A(n3368), .B(n3367), .Z(\w1[2][11] ) );
  XNOR U4860 ( .A(n3369), .B(key[376]), .Z(n3371) );
  XNOR U4861 ( .A(\w3[1][113] ), .B(\w3[1][121] ), .Z(n3370) );
  XNOR U4862 ( .A(n3371), .B(n3370), .Z(n3372) );
  XNOR U4863 ( .A(n3373), .B(n3372), .Z(\w1[2][120] ) );
  XNOR U4864 ( .A(n3705), .B(key[377]), .Z(n3375) );
  XNOR U4865 ( .A(\w3[1][114] ), .B(\w3[1][122] ), .Z(n3374) );
  XNOR U4866 ( .A(n3375), .B(n3374), .Z(n3376) );
  XNOR U4867 ( .A(n3377), .B(n3376), .Z(\w1[2][121] ) );
  XOR U4868 ( .A(\w3[1][123] ), .B(key[378]), .Z(n3379) );
  XNOR U4869 ( .A(\w3[1][114] ), .B(\w3[1][115] ), .Z(n3378) );
  XNOR U4870 ( .A(n3379), .B(n3378), .Z(n3381) );
  XOR U4871 ( .A(n3381), .B(n3380), .Z(\w1[2][122] ) );
  XOR U4872 ( .A(\w3[1][124] ), .B(n3382), .Z(n3383) );
  XOR U4873 ( .A(n3384), .B(n3383), .Z(n3713) );
  XOR U4874 ( .A(n3713), .B(key[379]), .Z(n3387) );
  XOR U4875 ( .A(\w3[1][99] ), .B(n3385), .Z(n3386) );
  XNOR U4876 ( .A(n3387), .B(n3386), .Z(\w1[2][123] ) );
  XNOR U4877 ( .A(n3388), .B(key[380]), .Z(n3392) );
  XNOR U4878 ( .A(n3390), .B(n3389), .Z(n3391) );
  XNOR U4879 ( .A(n3392), .B(n3391), .Z(\w1[2][124] ) );
  XOR U4880 ( .A(\w3[1][118] ), .B(key[381]), .Z(n3395) );
  XOR U4881 ( .A(n3393), .B(\w3[1][126] ), .Z(n3394) );
  XNOR U4882 ( .A(n3395), .B(n3394), .Z(n3396) );
  XOR U4883 ( .A(\w3[1][101] ), .B(n3396), .Z(\w1[2][125] ) );
  XNOR U4884 ( .A(n3397), .B(key[382]), .Z(n3400) );
  XOR U4885 ( .A(\w3[1][102] ), .B(n3398), .Z(n3399) );
  XNOR U4886 ( .A(n3400), .B(n3399), .Z(\w1[2][126] ) );
  XNOR U4887 ( .A(n3702), .B(key[383]), .Z(n3403) );
  XOR U4888 ( .A(\w3[1][103] ), .B(n3401), .Z(n3402) );
  XNOR U4889 ( .A(n3403), .B(n3402), .Z(\w1[2][127] ) );
  XOR U4890 ( .A(\w3[1][13] ), .B(\w3[1][28] ), .Z(n3405) );
  XNOR U4891 ( .A(\w3[1][8] ), .B(\w3[1][4] ), .Z(n3404) );
  XOR U4892 ( .A(n3405), .B(n3404), .Z(n3427) );
  XNOR U4893 ( .A(n3427), .B(key[268]), .Z(n3407) );
  XNOR U4894 ( .A(\w3[1][0] ), .B(\w3[1][5] ), .Z(n3528) );
  XOR U4895 ( .A(\w3[1][20] ), .B(n3528), .Z(n3406) );
  XNOR U4896 ( .A(n3407), .B(n3406), .Z(\w1[2][12] ) );
  IV U4897 ( .A(\w3[1][6] ), .Z(n3467) );
  XNOR U4898 ( .A(\w3[1][14] ), .B(n3467), .Z(n3409) );
  XNOR U4899 ( .A(\w3[1][5] ), .B(\w3[1][29] ), .Z(n3430) );
  XOR U4900 ( .A(n3430), .B(key[269]), .Z(n3408) );
  XNOR U4901 ( .A(n3409), .B(n3408), .Z(n3410) );
  XOR U4902 ( .A(\w3[1][21] ), .B(n3410), .Z(\w1[2][13] ) );
  IV U4903 ( .A(\w3[1][30] ), .Z(n3603) );
  XOR U4904 ( .A(\w3[1][6] ), .B(n3603), .Z(n3568) );
  XOR U4905 ( .A(\w3[1][8] ), .B(\w3[1][15] ), .Z(n3433) );
  XNOR U4906 ( .A(n3568), .B(n3433), .Z(n3431) );
  XOR U4907 ( .A(n3431), .B(key[270]), .Z(n3412) );
  XNOR U4908 ( .A(\w3[1][0] ), .B(\w3[1][7] ), .Z(n3604) );
  XOR U4909 ( .A(\w3[1][22] ), .B(n3604), .Z(n3411) );
  XNOR U4910 ( .A(n3412), .B(n3411), .Z(\w1[2][14] ) );
  XNOR U4911 ( .A(\w3[1][7] ), .B(\w3[1][31] ), .Z(n3432) );
  XNOR U4912 ( .A(n3432), .B(key[271]), .Z(n3414) );
  XOR U4913 ( .A(\w3[1][8] ), .B(\w3[1][0] ), .Z(n3437) );
  XNOR U4914 ( .A(\w3[1][23] ), .B(n3437), .Z(n3413) );
  XNOR U4915 ( .A(n3414), .B(n3413), .Z(\w1[2][15] ) );
  IV U4916 ( .A(\w3[1][9] ), .Z(n3672) );
  XOR U4917 ( .A(\w3[1][17] ), .B(n3672), .Z(n3441) );
  XNOR U4918 ( .A(n3441), .B(key[272]), .Z(n3416) );
  XNOR U4919 ( .A(\w3[1][24] ), .B(n3437), .Z(n3415) );
  XNOR U4920 ( .A(n3416), .B(n3415), .Z(\w1[2][16] ) );
  XNOR U4921 ( .A(\w3[1][18] ), .B(\w3[1][10] ), .Z(n3460) );
  XNOR U4922 ( .A(n3460), .B(key[273]), .Z(n3418) );
  XNOR U4923 ( .A(n3721), .B(n3672), .Z(n3417) );
  XNOR U4924 ( .A(n3418), .B(n3417), .Z(\w1[2][17] ) );
  XNOR U4925 ( .A(\w3[1][11] ), .B(\w3[1][19] ), .Z(n3446) );
  XNOR U4926 ( .A(n3446), .B(key[274]), .Z(n3420) );
  XOR U4927 ( .A(n3424), .B(\w3[1][10] ), .Z(n3419) );
  XNOR U4928 ( .A(n3420), .B(n3419), .Z(\w1[2][18] ) );
  IV U4929 ( .A(\w3[1][16] ), .Z(n3438) );
  XOR U4930 ( .A(n3438), .B(\w3[1][20] ), .Z(n3447) );
  XNOR U4931 ( .A(n3447), .B(key[275]), .Z(n3423) );
  XOR U4932 ( .A(\w3[1][11] ), .B(n3421), .Z(n3422) );
  XNOR U4933 ( .A(n3423), .B(n3422), .Z(\w1[2][19] ) );
  IV U4934 ( .A(\w3[1][17] ), .Z(n3717) );
  XOR U4935 ( .A(\w3[1][25] ), .B(n3717), .Z(n3436) );
  XNOR U4936 ( .A(n3436), .B(key[257]), .Z(n3426) );
  XNOR U4937 ( .A(n3424), .B(n3672), .Z(n3425) );
  XNOR U4938 ( .A(n3426), .B(n3425), .Z(\w1[2][1] ) );
  IV U4939 ( .A(\w3[1][21] ), .Z(n3455) );
  XOR U4940 ( .A(\w3[1][16] ), .B(n3455), .Z(n3452) );
  XNOR U4941 ( .A(n3452), .B(key[276]), .Z(n3429) );
  XOR U4942 ( .A(\w3[1][12] ), .B(n3427), .Z(n3428) );
  XNOR U4943 ( .A(n3429), .B(n3428), .Z(\w1[2][20] ) );
  IV U4944 ( .A(\w3[1][22] ), .Z(n3456) );
  XOR U4945 ( .A(\w3[1][14] ), .B(n3456), .Z(n3465) );
  XOR U4946 ( .A(n3438), .B(\w3[1][23] ), .Z(n3466) );
  XNOR U4947 ( .A(n3432), .B(key[279]), .Z(n3435) );
  XNOR U4948 ( .A(\w3[1][16] ), .B(n3433), .Z(n3434) );
  XNOR U4949 ( .A(n3435), .B(n3434), .Z(\w1[2][23] ) );
  XNOR U4950 ( .A(n3436), .B(key[280]), .Z(n3440) );
  XOR U4951 ( .A(n3438), .B(n3437), .Z(n3439) );
  XNOR U4952 ( .A(n3440), .B(n3439), .Z(\w1[2][24] ) );
  XNOR U4953 ( .A(n3460), .B(key[282]), .Z(n3443) );
  XNOR U4954 ( .A(\w3[1][2] ), .B(\w3[1][19] ), .Z(n3442) );
  XNOR U4955 ( .A(n3443), .B(n3442), .Z(n3444) );
  XOR U4956 ( .A(\w3[1][27] ), .B(n3444), .Z(\w1[2][26] ) );
  XOR U4957 ( .A(n3464), .B(\w3[1][28] ), .Z(n3445) );
  XOR U4958 ( .A(n3446), .B(n3445), .Z(n3492) );
  XOR U4959 ( .A(n3492), .B(key[283]), .Z(n3449) );
  XOR U4960 ( .A(\w3[1][3] ), .B(n3447), .Z(n3448) );
  XNOR U4961 ( .A(n3449), .B(n3448), .Z(\w1[2][27] ) );
  XOR U4962 ( .A(\w3[1][20] ), .B(\w3[1][29] ), .Z(n3451) );
  XOR U4963 ( .A(n3464), .B(\w3[1][12] ), .Z(n3450) );
  XOR U4964 ( .A(n3451), .B(n3450), .Z(n3527) );
  XNOR U4965 ( .A(n3527), .B(key[284]), .Z(n3454) );
  XOR U4966 ( .A(\w3[1][4] ), .B(n3452), .Z(n3453) );
  XNOR U4967 ( .A(n3454), .B(n3453), .Z(\w1[2][28] ) );
  XOR U4968 ( .A(\w3[1][13] ), .B(n3455), .Z(n3567) );
  XNOR U4969 ( .A(n3567), .B(key[285]), .Z(n3458) );
  XNOR U4970 ( .A(n3456), .B(n3603), .Z(n3457) );
  XNOR U4971 ( .A(n3458), .B(n3457), .Z(n3459) );
  XOR U4972 ( .A(\w3[1][5] ), .B(n3459), .Z(\w1[2][29] ) );
  XNOR U4973 ( .A(n3460), .B(key[258]), .Z(n3463) );
  XOR U4974 ( .A(\w3[1][26] ), .B(n3461), .Z(n3462) );
  XNOR U4975 ( .A(n3463), .B(n3462), .Z(\w1[2][2] ) );
  XOR U4976 ( .A(n3464), .B(\w3[1][31] ), .Z(n3639) );
  XNOR U4977 ( .A(n3465), .B(n3639), .Z(n3602) );
  XNOR U4978 ( .A(n3602), .B(key[286]), .Z(n3469) );
  XNOR U4979 ( .A(n3467), .B(n3466), .Z(n3468) );
  XNOR U4980 ( .A(n3469), .B(n3468), .Z(\w1[2][30] ) );
  XNOR U4981 ( .A(\w3[1][15] ), .B(\w3[1][23] ), .Z(n3638) );
  XNOR U4982 ( .A(n3638), .B(key[287]), .Z(n3471) );
  XOR U4983 ( .A(n3673), .B(\w3[1][7] ), .Z(n3470) );
  XNOR U4984 ( .A(n3471), .B(n3470), .Z(\w1[2][31] ) );
  XNOR U4985 ( .A(\w3[1][48] ), .B(\w3[1][56] ), .Z(n3584) );
  XNOR U4986 ( .A(\w3[1][33] ), .B(\w3[1][57] ), .Z(n3524) );
  XNOR U4987 ( .A(\w3[1][40] ), .B(key[288]), .Z(n3472) );
  XNOR U4988 ( .A(n3524), .B(n3472), .Z(n3473) );
  XOR U4989 ( .A(n3584), .B(n3473), .Z(\w1[2][32] ) );
  XNOR U4990 ( .A(\w3[1][34] ), .B(\w3[1][58] ), .Z(n3532) );
  XNOR U4991 ( .A(\w3[1][41] ), .B(\w3[1][49] ), .Z(n3554) );
  XOR U4992 ( .A(n3554), .B(key[289]), .Z(n3474) );
  XNOR U4993 ( .A(n3532), .B(n3474), .Z(n3475) );
  XNOR U4994 ( .A(\w3[1][57] ), .B(n3475), .Z(\w1[2][33] ) );
  XNOR U4995 ( .A(n3502), .B(key[290]), .Z(n3477) );
  XNOR U4996 ( .A(\w3[1][42] ), .B(\w3[1][50] ), .Z(n3557) );
  XOR U4997 ( .A(\w3[1][58] ), .B(n3557), .Z(n3476) );
  XNOR U4998 ( .A(n3477), .B(n3476), .Z(\w1[2][34] ) );
  XOR U4999 ( .A(\w3[1][36] ), .B(\w3[1][32] ), .Z(n3504) );
  XOR U5000 ( .A(n3504), .B(key[291]), .Z(n3480) );
  IV U5001 ( .A(\w3[1][51] ), .Z(n3556) );
  XOR U5002 ( .A(\w3[1][43] ), .B(n3556), .Z(n3531) );
  XOR U5003 ( .A(\w3[1][56] ), .B(n3531), .Z(n3478) );
  XNOR U5004 ( .A(\w3[1][60] ), .B(n3478), .Z(n3563) );
  XNOR U5005 ( .A(\w3[1][59] ), .B(n3563), .Z(n3479) );
  XNOR U5006 ( .A(n3480), .B(n3479), .Z(\w1[2][35] ) );
  XOR U5007 ( .A(\w3[1][32] ), .B(\w3[1][37] ), .Z(n3510) );
  XOR U5008 ( .A(\w3[1][52] ), .B(\w3[1][61] ), .Z(n3482) );
  XNOR U5009 ( .A(\w3[1][56] ), .B(\w3[1][44] ), .Z(n3481) );
  XOR U5010 ( .A(n3482), .B(n3481), .Z(n3572) );
  XOR U5011 ( .A(n3572), .B(key[292]), .Z(n3483) );
  XOR U5012 ( .A(n3510), .B(n3483), .Z(n3484) );
  XNOR U5013 ( .A(\w3[1][60] ), .B(n3484), .Z(\w1[2][36] ) );
  XNOR U5014 ( .A(\w3[1][38] ), .B(\w3[1][62] ), .Z(n3516) );
  XNOR U5015 ( .A(n3516), .B(key[293]), .Z(n3486) );
  IV U5016 ( .A(\w3[1][53] ), .Z(n3536) );
  XOR U5017 ( .A(\w3[1][45] ), .B(n3536), .Z(n3575) );
  XOR U5018 ( .A(\w3[1][61] ), .B(n3575), .Z(n3485) );
  XNOR U5019 ( .A(n3486), .B(n3485), .Z(\w1[2][37] ) );
  XOR U5020 ( .A(\w3[1][32] ), .B(\w3[1][39] ), .Z(n3517) );
  XOR U5021 ( .A(n3517), .B(key[294]), .Z(n3488) );
  XNOR U5022 ( .A(\w3[1][56] ), .B(\w3[1][63] ), .Z(n3489) );
  XOR U5023 ( .A(\w3[1][46] ), .B(\w3[1][54] ), .Z(n3541) );
  XOR U5024 ( .A(n3489), .B(n3541), .Z(n3580) );
  XOR U5025 ( .A(\w3[1][62] ), .B(n3580), .Z(n3487) );
  XNOR U5026 ( .A(n3488), .B(n3487), .Z(\w1[2][38] ) );
  XNOR U5027 ( .A(\w3[1][47] ), .B(\w3[1][55] ), .Z(n3583) );
  XNOR U5028 ( .A(n3583), .B(key[295]), .Z(n3491) );
  XOR U5029 ( .A(\w3[1][32] ), .B(n3489), .Z(n3490) );
  XNOR U5030 ( .A(n3491), .B(n3490), .Z(\w1[2][39] ) );
  XOR U5031 ( .A(n3492), .B(key[259]), .Z(n3495) );
  XOR U5032 ( .A(n3493), .B(\w3[1][27] ), .Z(n3494) );
  XNOR U5033 ( .A(n3495), .B(n3494), .Z(\w1[2][3] ) );
  IV U5034 ( .A(\w3[1][33] ), .Z(n3555) );
  XOR U5035 ( .A(\w3[1][42] ), .B(key[297]), .Z(n3497) );
  IV U5036 ( .A(\w3[1][34] ), .Z(n3561) );
  XOR U5037 ( .A(\w3[1][49] ), .B(n3561), .Z(n3496) );
  XNOR U5038 ( .A(n3497), .B(n3496), .Z(n3498) );
  XNOR U5039 ( .A(n3498), .B(n3524), .Z(\w1[2][41] ) );
  XOR U5040 ( .A(\w3[1][43] ), .B(key[298]), .Z(n3500) );
  IV U5041 ( .A(\w3[1][35] ), .Z(n3564) );
  XOR U5042 ( .A(\w3[1][50] ), .B(n3564), .Z(n3499) );
  XNOR U5043 ( .A(n3500), .B(n3499), .Z(n3501) );
  XNOR U5044 ( .A(n3501), .B(n3532), .Z(\w1[2][42] ) );
  IV U5045 ( .A(\w3[1][40] ), .Z(n3507) );
  XNOR U5046 ( .A(n3507), .B(n3502), .Z(n3503) );
  XOR U5047 ( .A(\w3[1][44] ), .B(n3503), .Z(n3535) );
  XNOR U5048 ( .A(n3535), .B(key[299]), .Z(n3506) );
  XNOR U5049 ( .A(\w3[1][51] ), .B(n3504), .Z(n3505) );
  XNOR U5050 ( .A(n3506), .B(n3505), .Z(\w1[2][43] ) );
  XOR U5051 ( .A(\w3[1][36] ), .B(\w3[1][45] ), .Z(n3509) );
  XOR U5052 ( .A(n3507), .B(\w3[1][60] ), .Z(n3508) );
  XOR U5053 ( .A(n3509), .B(n3508), .Z(n3537) );
  XNOR U5054 ( .A(n3537), .B(key[300]), .Z(n3512) );
  XNOR U5055 ( .A(\w3[1][52] ), .B(n3510), .Z(n3511) );
  XNOR U5056 ( .A(n3512), .B(n3511), .Z(\w1[2][44] ) );
  XNOR U5057 ( .A(\w3[1][61] ), .B(\w3[1][37] ), .Z(n3540) );
  XNOR U5058 ( .A(n3540), .B(key[301]), .Z(n3514) );
  XNOR U5059 ( .A(\w3[1][38] ), .B(\w3[1][46] ), .Z(n3513) );
  XNOR U5060 ( .A(n3514), .B(n3513), .Z(n3515) );
  XOR U5061 ( .A(\w3[1][53] ), .B(n3515), .Z(\w1[2][45] ) );
  XOR U5062 ( .A(\w3[1][40] ), .B(\w3[1][47] ), .Z(n3546) );
  XOR U5063 ( .A(n3516), .B(n3546), .Z(n3542) );
  XNOR U5064 ( .A(n3542), .B(key[302]), .Z(n3519) );
  XNOR U5065 ( .A(\w3[1][54] ), .B(n3517), .Z(n3518) );
  XNOR U5066 ( .A(n3519), .B(n3518), .Z(\w1[2][46] ) );
  XOR U5067 ( .A(\w3[1][63] ), .B(\w3[1][39] ), .Z(n3545) );
  XOR U5068 ( .A(n3545), .B(key[303]), .Z(n3521) );
  XNOR U5069 ( .A(\w3[1][40] ), .B(\w3[1][32] ), .Z(n3549) );
  XOR U5070 ( .A(\w3[1][55] ), .B(n3549), .Z(n3520) );
  XNOR U5071 ( .A(n3521), .B(n3520), .Z(\w1[2][47] ) );
  XNOR U5072 ( .A(n3549), .B(key[304]), .Z(n3523) );
  XOR U5073 ( .A(\w3[1][56] ), .B(n3554), .Z(n3522) );
  XNOR U5074 ( .A(n3523), .B(n3522), .Z(\w1[2][48] ) );
  XNOR U5075 ( .A(n3557), .B(key[305]), .Z(n3526) );
  XOR U5076 ( .A(n3524), .B(\w3[1][41] ), .Z(n3525) );
  XNOR U5077 ( .A(n3526), .B(n3525), .Z(\w1[2][49] ) );
  XNOR U5078 ( .A(n3527), .B(key[260]), .Z(n3530) );
  XOR U5079 ( .A(n3528), .B(\w3[1][28] ), .Z(n3529) );
  XNOR U5080 ( .A(n3530), .B(n3529), .Z(\w1[2][4] ) );
  XNOR U5081 ( .A(n3531), .B(key[306]), .Z(n3534) );
  XOR U5082 ( .A(n3532), .B(\w3[1][42] ), .Z(n3533) );
  XNOR U5083 ( .A(n3534), .B(n3533), .Z(\w1[2][50] ) );
  IV U5084 ( .A(\w3[1][48] ), .Z(n3550) );
  XOR U5085 ( .A(n3550), .B(\w3[1][52] ), .Z(n3562) );
  XOR U5086 ( .A(\w3[1][48] ), .B(n3536), .Z(n3571) );
  XNOR U5087 ( .A(n3571), .B(key[308]), .Z(n3539) );
  XOR U5088 ( .A(\w3[1][44] ), .B(n3537), .Z(n3538) );
  XNOR U5089 ( .A(n3539), .B(n3538), .Z(\w1[2][52] ) );
  XOR U5090 ( .A(n3550), .B(\w3[1][55] ), .Z(n3579) );
  XNOR U5091 ( .A(n3579), .B(key[310]), .Z(n3544) );
  XOR U5092 ( .A(\w3[1][46] ), .B(n3542), .Z(n3543) );
  XNOR U5093 ( .A(n3544), .B(n3543), .Z(\w1[2][54] ) );
  XOR U5094 ( .A(n3545), .B(key[311]), .Z(n3548) );
  XNOR U5095 ( .A(\w3[1][48] ), .B(n3546), .Z(n3547) );
  XNOR U5096 ( .A(n3548), .B(n3547), .Z(\w1[2][55] ) );
  XNOR U5097 ( .A(n3549), .B(key[312]), .Z(n3552) );
  XOR U5098 ( .A(n3550), .B(\w3[1][49] ), .Z(n3551) );
  XNOR U5099 ( .A(n3552), .B(n3551), .Z(n3553) );
  XOR U5100 ( .A(\w3[1][57] ), .B(n3553), .Z(\w1[2][56] ) );
  XNOR U5101 ( .A(n3556), .B(key[314]), .Z(n3559) );
  XOR U5102 ( .A(n3557), .B(\w3[1][59] ), .Z(n3558) );
  XNOR U5103 ( .A(n3559), .B(n3558), .Z(n3560) );
  XNOR U5104 ( .A(n3561), .B(n3560), .Z(\w1[2][58] ) );
  XNOR U5105 ( .A(n3562), .B(key[315]), .Z(n3566) );
  XOR U5106 ( .A(n3564), .B(n3563), .Z(n3565) );
  XNOR U5107 ( .A(n3566), .B(n3565), .Z(\w1[2][59] ) );
  XNOR U5108 ( .A(n3567), .B(key[261]), .Z(n3570) );
  XOR U5109 ( .A(\w3[1][29] ), .B(n3568), .Z(n3569) );
  XNOR U5110 ( .A(n3570), .B(n3569), .Z(\w1[2][5] ) );
  XNOR U5111 ( .A(n3571), .B(key[316]), .Z(n3574) );
  XOR U5112 ( .A(\w3[1][36] ), .B(n3572), .Z(n3573) );
  XNOR U5113 ( .A(n3574), .B(n3573), .Z(\w1[2][60] ) );
  XOR U5114 ( .A(\w3[1][54] ), .B(key[317]), .Z(n3577) );
  XOR U5115 ( .A(n3575), .B(\w3[1][62] ), .Z(n3576) );
  XNOR U5116 ( .A(n3577), .B(n3576), .Z(n3578) );
  XOR U5117 ( .A(\w3[1][37] ), .B(n3578), .Z(\w1[2][61] ) );
  XNOR U5118 ( .A(n3579), .B(key[318]), .Z(n3582) );
  XOR U5119 ( .A(\w3[1][38] ), .B(n3580), .Z(n3581) );
  XNOR U5120 ( .A(n3582), .B(n3581), .Z(\w1[2][62] ) );
  XNOR U5121 ( .A(n3583), .B(key[319]), .Z(n3586) );
  XOR U5122 ( .A(n3584), .B(\w3[1][39] ), .Z(n3585) );
  XNOR U5123 ( .A(n3586), .B(n3585), .Z(\w1[2][63] ) );
  XNOR U5124 ( .A(\w3[1][80] ), .B(\w3[1][88] ), .Z(n3698) );
  XNOR U5125 ( .A(\w3[1][65] ), .B(\w3[1][89] ), .Z(n3644) );
  XNOR U5126 ( .A(\w3[1][72] ), .B(key[320]), .Z(n3587) );
  XNOR U5127 ( .A(n3644), .B(n3587), .Z(n3588) );
  XOR U5128 ( .A(n3698), .B(n3588), .Z(\w1[2][64] ) );
  XNOR U5129 ( .A(\w3[1][66] ), .B(\w3[1][90] ), .Z(n3648) );
  XNOR U5130 ( .A(\w3[1][73] ), .B(\w3[1][81] ), .Z(n3670) );
  XOR U5131 ( .A(n3670), .B(key[321]), .Z(n3589) );
  XNOR U5132 ( .A(n3648), .B(n3589), .Z(n3590) );
  XNOR U5133 ( .A(\w3[1][89] ), .B(n3590), .Z(\w1[2][65] ) );
  XNOR U5134 ( .A(n3618), .B(key[322]), .Z(n3592) );
  XNOR U5135 ( .A(\w3[1][74] ), .B(\w3[1][82] ), .Z(n3675) );
  XOR U5136 ( .A(\w3[1][90] ), .B(n3675), .Z(n3591) );
  XNOR U5137 ( .A(n3592), .B(n3591), .Z(\w1[2][66] ) );
  XOR U5138 ( .A(\w3[1][68] ), .B(\w3[1][64] ), .Z(n3620) );
  XOR U5139 ( .A(n3620), .B(key[323]), .Z(n3595) );
  IV U5140 ( .A(\w3[1][83] ), .Z(n3674) );
  XOR U5141 ( .A(\w3[1][75] ), .B(n3674), .Z(n3647) );
  XOR U5142 ( .A(\w3[1][88] ), .B(n3647), .Z(n3593) );
  XNOR U5143 ( .A(\w3[1][92] ), .B(n3593), .Z(n3681) );
  XNOR U5144 ( .A(\w3[1][91] ), .B(n3681), .Z(n3594) );
  XNOR U5145 ( .A(n3595), .B(n3594), .Z(\w1[2][67] ) );
  XOR U5146 ( .A(\w3[1][64] ), .B(\w3[1][69] ), .Z(n3626) );
  XOR U5147 ( .A(\w3[1][84] ), .B(\w3[1][93] ), .Z(n3597) );
  XNOR U5148 ( .A(\w3[1][88] ), .B(\w3[1][76] ), .Z(n3596) );
  XOR U5149 ( .A(n3597), .B(n3596), .Z(n3686) );
  XOR U5150 ( .A(n3686), .B(key[324]), .Z(n3598) );
  XOR U5151 ( .A(n3626), .B(n3598), .Z(n3599) );
  XNOR U5152 ( .A(\w3[1][92] ), .B(n3599), .Z(\w1[2][68] ) );
  XNOR U5153 ( .A(\w3[1][70] ), .B(\w3[1][94] ), .Z(n3632) );
  XNOR U5154 ( .A(n3632), .B(key[325]), .Z(n3601) );
  IV U5155 ( .A(\w3[1][85] ), .Z(n3652) );
  XOR U5156 ( .A(\w3[1][77] ), .B(n3652), .Z(n3689) );
  XOR U5157 ( .A(\w3[1][93] ), .B(n3689), .Z(n3600) );
  XNOR U5158 ( .A(n3601), .B(n3600), .Z(\w1[2][69] ) );
  XNOR U5159 ( .A(n3602), .B(key[262]), .Z(n3606) );
  XNOR U5160 ( .A(n3604), .B(n3603), .Z(n3605) );
  XNOR U5161 ( .A(n3606), .B(n3605), .Z(\w1[2][6] ) );
  XOR U5162 ( .A(\w3[1][64] ), .B(\w3[1][71] ), .Z(n3633) );
  XOR U5163 ( .A(n3633), .B(key[326]), .Z(n3608) );
  XNOR U5164 ( .A(\w3[1][88] ), .B(\w3[1][95] ), .Z(n3609) );
  XOR U5165 ( .A(\w3[1][78] ), .B(\w3[1][86] ), .Z(n3657) );
  XOR U5166 ( .A(n3609), .B(n3657), .Z(n3694) );
  XOR U5167 ( .A(\w3[1][94] ), .B(n3694), .Z(n3607) );
  XNOR U5168 ( .A(n3608), .B(n3607), .Z(\w1[2][70] ) );
  XNOR U5169 ( .A(\w3[1][79] ), .B(\w3[1][87] ), .Z(n3697) );
  XNOR U5170 ( .A(n3697), .B(key[327]), .Z(n3611) );
  XOR U5171 ( .A(\w3[1][64] ), .B(n3609), .Z(n3610) );
  XNOR U5172 ( .A(n3611), .B(n3610), .Z(\w1[2][71] ) );
  IV U5173 ( .A(\w3[1][65] ), .Z(n3671) );
  XOR U5174 ( .A(\w3[1][74] ), .B(key[329]), .Z(n3613) );
  IV U5175 ( .A(\w3[1][66] ), .Z(n3679) );
  XOR U5176 ( .A(\w3[1][81] ), .B(n3679), .Z(n3612) );
  XNOR U5177 ( .A(n3613), .B(n3612), .Z(n3614) );
  XNOR U5178 ( .A(n3614), .B(n3644), .Z(\w1[2][73] ) );
  XOR U5179 ( .A(\w3[1][75] ), .B(key[330]), .Z(n3616) );
  IV U5180 ( .A(\w3[1][67] ), .Z(n3682) );
  XOR U5181 ( .A(\w3[1][82] ), .B(n3682), .Z(n3615) );
  XNOR U5182 ( .A(n3616), .B(n3615), .Z(n3617) );
  XNOR U5183 ( .A(n3617), .B(n3648), .Z(\w1[2][74] ) );
  IV U5184 ( .A(\w3[1][72] ), .Z(n3623) );
  XNOR U5185 ( .A(n3623), .B(n3618), .Z(n3619) );
  XOR U5186 ( .A(\w3[1][76] ), .B(n3619), .Z(n3651) );
  XNOR U5187 ( .A(n3651), .B(key[331]), .Z(n3622) );
  XNOR U5188 ( .A(\w3[1][83] ), .B(n3620), .Z(n3621) );
  XNOR U5189 ( .A(n3622), .B(n3621), .Z(\w1[2][75] ) );
  XOR U5190 ( .A(\w3[1][68] ), .B(\w3[1][77] ), .Z(n3625) );
  XOR U5191 ( .A(n3623), .B(\w3[1][92] ), .Z(n3624) );
  XOR U5192 ( .A(n3625), .B(n3624), .Z(n3653) );
  XNOR U5193 ( .A(n3653), .B(key[332]), .Z(n3628) );
  XNOR U5194 ( .A(\w3[1][84] ), .B(n3626), .Z(n3627) );
  XNOR U5195 ( .A(n3628), .B(n3627), .Z(\w1[2][76] ) );
  XNOR U5196 ( .A(\w3[1][93] ), .B(\w3[1][69] ), .Z(n3656) );
  XNOR U5197 ( .A(n3656), .B(key[333]), .Z(n3630) );
  XNOR U5198 ( .A(\w3[1][70] ), .B(\w3[1][78] ), .Z(n3629) );
  XNOR U5199 ( .A(n3630), .B(n3629), .Z(n3631) );
  XOR U5200 ( .A(\w3[1][85] ), .B(n3631), .Z(\w1[2][77] ) );
  XOR U5201 ( .A(\w3[1][72] ), .B(\w3[1][79] ), .Z(n3662) );
  XOR U5202 ( .A(n3632), .B(n3662), .Z(n3658) );
  XNOR U5203 ( .A(n3658), .B(key[334]), .Z(n3635) );
  XNOR U5204 ( .A(\w3[1][86] ), .B(n3633), .Z(n3634) );
  XNOR U5205 ( .A(n3635), .B(n3634), .Z(\w1[2][78] ) );
  XOR U5206 ( .A(\w3[1][95] ), .B(\w3[1][71] ), .Z(n3661) );
  XOR U5207 ( .A(n3661), .B(key[335]), .Z(n3637) );
  XNOR U5208 ( .A(\w3[1][72] ), .B(\w3[1][64] ), .Z(n3665) );
  XOR U5209 ( .A(\w3[1][87] ), .B(n3665), .Z(n3636) );
  XNOR U5210 ( .A(n3637), .B(n3636), .Z(\w1[2][79] ) );
  XNOR U5211 ( .A(n3638), .B(key[263]), .Z(n3641) );
  XOR U5212 ( .A(\w3[1][0] ), .B(n3639), .Z(n3640) );
  XNOR U5213 ( .A(n3641), .B(n3640), .Z(\w1[2][7] ) );
  XNOR U5214 ( .A(n3665), .B(key[336]), .Z(n3643) );
  XOR U5215 ( .A(\w3[1][88] ), .B(n3670), .Z(n3642) );
  XNOR U5216 ( .A(n3643), .B(n3642), .Z(\w1[2][80] ) );
  XNOR U5217 ( .A(n3675), .B(key[337]), .Z(n3646) );
  XOR U5218 ( .A(n3644), .B(\w3[1][73] ), .Z(n3645) );
  XNOR U5219 ( .A(n3646), .B(n3645), .Z(\w1[2][81] ) );
  XNOR U5220 ( .A(n3647), .B(key[338]), .Z(n3650) );
  XOR U5221 ( .A(n3648), .B(\w3[1][74] ), .Z(n3649) );
  XNOR U5222 ( .A(n3650), .B(n3649), .Z(\w1[2][82] ) );
  IV U5223 ( .A(\w3[1][80] ), .Z(n3666) );
  XOR U5224 ( .A(n3666), .B(\w3[1][84] ), .Z(n3680) );
  XOR U5225 ( .A(\w3[1][80] ), .B(n3652), .Z(n3685) );
  XNOR U5226 ( .A(n3685), .B(key[340]), .Z(n3655) );
  XOR U5227 ( .A(\w3[1][76] ), .B(n3653), .Z(n3654) );
  XNOR U5228 ( .A(n3655), .B(n3654), .Z(\w1[2][84] ) );
  XOR U5229 ( .A(n3666), .B(\w3[1][87] ), .Z(n3693) );
  XNOR U5230 ( .A(n3693), .B(key[342]), .Z(n3660) );
  XOR U5231 ( .A(\w3[1][78] ), .B(n3658), .Z(n3659) );
  XNOR U5232 ( .A(n3660), .B(n3659), .Z(\w1[2][86] ) );
  XOR U5233 ( .A(n3661), .B(key[343]), .Z(n3664) );
  XNOR U5234 ( .A(\w3[1][80] ), .B(n3662), .Z(n3663) );
  XNOR U5235 ( .A(n3664), .B(n3663), .Z(\w1[2][87] ) );
  XNOR U5236 ( .A(n3665), .B(key[344]), .Z(n3668) );
  XOR U5237 ( .A(n3666), .B(\w3[1][81] ), .Z(n3667) );
  XNOR U5238 ( .A(n3668), .B(n3667), .Z(n3669) );
  XOR U5239 ( .A(\w3[1][89] ), .B(n3669), .Z(\w1[2][88] ) );
  XNOR U5240 ( .A(n3674), .B(key[346]), .Z(n3677) );
  XOR U5241 ( .A(n3675), .B(\w3[1][91] ), .Z(n3676) );
  XNOR U5242 ( .A(n3677), .B(n3676), .Z(n3678) );
  XNOR U5243 ( .A(n3679), .B(n3678), .Z(\w1[2][90] ) );
  XNOR U5244 ( .A(n3680), .B(key[347]), .Z(n3684) );
  XOR U5245 ( .A(n3682), .B(n3681), .Z(n3683) );
  XNOR U5246 ( .A(n3684), .B(n3683), .Z(\w1[2][91] ) );
  XNOR U5247 ( .A(n3685), .B(key[348]), .Z(n3688) );
  XOR U5248 ( .A(\w3[1][68] ), .B(n3686), .Z(n3687) );
  XNOR U5249 ( .A(n3688), .B(n3687), .Z(\w1[2][92] ) );
  XOR U5250 ( .A(\w3[1][86] ), .B(key[349]), .Z(n3691) );
  XOR U5251 ( .A(n3689), .B(\w3[1][94] ), .Z(n3690) );
  XNOR U5252 ( .A(n3691), .B(n3690), .Z(n3692) );
  XOR U5253 ( .A(\w3[1][69] ), .B(n3692), .Z(\w1[2][93] ) );
  XNOR U5254 ( .A(n3693), .B(key[350]), .Z(n3696) );
  XOR U5255 ( .A(\w3[1][70] ), .B(n3694), .Z(n3695) );
  XNOR U5256 ( .A(n3696), .B(n3695), .Z(\w1[2][94] ) );
  XNOR U5257 ( .A(n3697), .B(key[351]), .Z(n3700) );
  XOR U5258 ( .A(n3698), .B(\w3[1][71] ), .Z(n3699) );
  XNOR U5259 ( .A(n3700), .B(n3699), .Z(\w1[2][95] ) );
  XOR U5260 ( .A(\w3[1][104] ), .B(key[352]), .Z(n3704) );
  XNOR U5261 ( .A(n3702), .B(n3701), .Z(n3703) );
  XNOR U5262 ( .A(n3704), .B(n3703), .Z(\w1[2][96] ) );
  XNOR U5263 ( .A(n3705), .B(key[353]), .Z(n3708) );
  XOR U5264 ( .A(\w3[1][121] ), .B(n3706), .Z(n3707) );
  XNOR U5265 ( .A(n3708), .B(n3707), .Z(\w1[2][97] ) );
  XNOR U5266 ( .A(n3709), .B(key[354]), .Z(n3712) );
  XOR U5267 ( .A(\w3[1][122] ), .B(n3710), .Z(n3711) );
  XNOR U5268 ( .A(n3712), .B(n3711), .Z(\w1[2][98] ) );
  XOR U5269 ( .A(n3713), .B(key[355]), .Z(n3716) );
  XOR U5270 ( .A(n3714), .B(\w3[1][123] ), .Z(n3715) );
  XNOR U5271 ( .A(n3716), .B(n3715), .Z(\w1[2][99] ) );
  XOR U5272 ( .A(\w3[1][10] ), .B(key[265]), .Z(n3719) );
  XOR U5273 ( .A(\w3[1][2] ), .B(n3717), .Z(n3718) );
  XNOR U5274 ( .A(n3719), .B(n3718), .Z(n3720) );
  XNOR U5275 ( .A(n3721), .B(n3720), .Z(\w1[2][9] ) );
  XNOR U5276 ( .A(\w3[2][1] ), .B(\w3[2][25] ), .Z(n4136) );
  IV U5277 ( .A(\w3[2][24] ), .Z(n3880) );
  XOR U5278 ( .A(\w3[2][16] ), .B(n3880), .Z(n4089) );
  XNOR U5279 ( .A(\w3[2][8] ), .B(key[384]), .Z(n3722) );
  XNOR U5280 ( .A(n4089), .B(n3722), .Z(n3723) );
  XOR U5281 ( .A(n4136), .B(n3723), .Z(\w1[3][0] ) );
  XOR U5282 ( .A(\w3[2][96] ), .B(\w3[2][101] ), .Z(n3746) );
  XOR U5283 ( .A(\w3[2][116] ), .B(\w3[2][125] ), .Z(n3725) );
  IV U5284 ( .A(\w3[2][120] ), .Z(n3798) );
  XOR U5285 ( .A(n3798), .B(\w3[2][108] ), .Z(n3724) );
  XOR U5286 ( .A(n3725), .B(n3724), .Z(n3806) );
  XOR U5287 ( .A(n3806), .B(key[484]), .Z(n3726) );
  XOR U5288 ( .A(n3746), .B(n3726), .Z(n3727) );
  XNOR U5289 ( .A(\w3[2][124] ), .B(n3727), .Z(\w1[3][100] ) );
  XNOR U5290 ( .A(\w3[2][102] ), .B(\w3[2][126] ), .Z(n3755) );
  XNOR U5291 ( .A(n3755), .B(key[485]), .Z(n3729) );
  XNOR U5292 ( .A(\w3[2][109] ), .B(\w3[2][117] ), .Z(n3809) );
  XOR U5293 ( .A(\w3[2][125] ), .B(n3809), .Z(n3728) );
  XNOR U5294 ( .A(n3729), .B(n3728), .Z(\w1[3][101] ) );
  XOR U5295 ( .A(\w3[2][96] ), .B(\w3[2][103] ), .Z(n3756) );
  XOR U5296 ( .A(n3756), .B(key[486]), .Z(n3731) );
  XOR U5297 ( .A(n3798), .B(\w3[2][127] ), .Z(n3732) );
  XOR U5298 ( .A(\w3[2][110] ), .B(\w3[2][118] ), .Z(n3774) );
  XOR U5299 ( .A(n3732), .B(n3774), .Z(n3814) );
  XOR U5300 ( .A(\w3[2][126] ), .B(n3814), .Z(n3730) );
  XNOR U5301 ( .A(n3731), .B(n3730), .Z(\w1[3][102] ) );
  XNOR U5302 ( .A(\w3[2][111] ), .B(\w3[2][119] ), .Z(n3817) );
  XNOR U5303 ( .A(n3817), .B(key[487]), .Z(n3734) );
  XOR U5304 ( .A(\w3[2][96] ), .B(n3732), .Z(n3733) );
  XNOR U5305 ( .A(n3734), .B(n3733), .Z(\w1[3][103] ) );
  IV U5306 ( .A(\w3[2][97] ), .Z(n3794) );
  IV U5307 ( .A(\w3[2][112] ), .Z(n3790) );
  XOR U5308 ( .A(\w3[2][120] ), .B(n3790), .Z(n4118) );
  XOR U5309 ( .A(\w3[2][106] ), .B(\w3[2][113] ), .Z(n3736) );
  XNOR U5310 ( .A(\w3[2][97] ), .B(\w3[2][121] ), .Z(n4117) );
  XOR U5311 ( .A(n4117), .B(key[489]), .Z(n3735) );
  XNOR U5312 ( .A(n3736), .B(n3735), .Z(n3737) );
  XOR U5313 ( .A(\w3[2][98] ), .B(n3737), .Z(\w1[3][105] ) );
  XOR U5314 ( .A(\w3[2][107] ), .B(\w3[2][114] ), .Z(n3739) );
  XOR U5315 ( .A(\w3[2][98] ), .B(\w3[2][122] ), .Z(n4122) );
  XNOR U5316 ( .A(n4122), .B(key[490]), .Z(n3738) );
  XNOR U5317 ( .A(n3739), .B(n3738), .Z(n3740) );
  XOR U5318 ( .A(\w3[2][99] ), .B(n3740), .Z(\w1[3][106] ) );
  XNOR U5319 ( .A(\w3[2][99] ), .B(\w3[2][123] ), .Z(n4126) );
  XOR U5320 ( .A(\w3[2][108] ), .B(n4126), .Z(n3741) );
  XOR U5321 ( .A(\w3[2][104] ), .B(n3741), .Z(n3767) );
  XNOR U5322 ( .A(n3767), .B(key[491]), .Z(n3743) );
  IV U5323 ( .A(\w3[2][100] ), .Z(n3805) );
  XOR U5324 ( .A(\w3[2][96] ), .B(n3805), .Z(n4130) );
  XOR U5325 ( .A(\w3[2][115] ), .B(n4130), .Z(n3742) );
  XNOR U5326 ( .A(n3743), .B(n3742), .Z(\w1[3][107] ) );
  XOR U5327 ( .A(\w3[2][100] ), .B(\w3[2][104] ), .Z(n3745) );
  XNOR U5328 ( .A(\w3[2][124] ), .B(\w3[2][109] ), .Z(n3744) );
  XOR U5329 ( .A(n3745), .B(n3744), .Z(n3770) );
  XNOR U5330 ( .A(n3770), .B(key[492]), .Z(n3748) );
  XNOR U5331 ( .A(\w3[2][116] ), .B(n3746), .Z(n3747) );
  XNOR U5332 ( .A(n3748), .B(n3747), .Z(\w1[3][108] ) );
  XNOR U5333 ( .A(\w3[2][125] ), .B(\w3[2][101] ), .Z(n3773) );
  XNOR U5334 ( .A(n3773), .B(key[493]), .Z(n3750) );
  XNOR U5335 ( .A(\w3[2][102] ), .B(\w3[2][110] ), .Z(n3749) );
  XNOR U5336 ( .A(n3750), .B(n3749), .Z(n3751) );
  XOR U5337 ( .A(\w3[2][117] ), .B(n3751), .Z(\w1[3][109] ) );
  XOR U5338 ( .A(\w3[2][11] ), .B(\w3[2][3] ), .Z(n3753) );
  XNOR U5339 ( .A(\w3[2][2] ), .B(\w3[2][26] ), .Z(n3840) );
  XOR U5340 ( .A(n3840), .B(key[394]), .Z(n3752) );
  XNOR U5341 ( .A(n3753), .B(n3752), .Z(n3754) );
  XOR U5342 ( .A(\w3[2][18] ), .B(n3754), .Z(\w1[3][10] ) );
  XOR U5343 ( .A(\w3[2][111] ), .B(\w3[2][104] ), .Z(n3781) );
  XOR U5344 ( .A(n3755), .B(n3781), .Z(n3777) );
  XNOR U5345 ( .A(n3777), .B(key[494]), .Z(n3758) );
  XNOR U5346 ( .A(\w3[2][118] ), .B(n3756), .Z(n3757) );
  XNOR U5347 ( .A(n3758), .B(n3757), .Z(\w1[3][110] ) );
  XOR U5348 ( .A(\w3[2][127] ), .B(\w3[2][103] ), .Z(n3780) );
  XOR U5349 ( .A(n3780), .B(key[495]), .Z(n3760) );
  XNOR U5350 ( .A(\w3[2][96] ), .B(\w3[2][104] ), .Z(n3786) );
  XOR U5351 ( .A(\w3[2][119] ), .B(n3786), .Z(n3759) );
  XNOR U5352 ( .A(n3760), .B(n3759), .Z(\w1[3][111] ) );
  XNOR U5353 ( .A(\w3[2][105] ), .B(\w3[2][113] ), .Z(n4121) );
  XNOR U5354 ( .A(n4121), .B(key[496]), .Z(n3762) );
  XNOR U5355 ( .A(n3798), .B(n3786), .Z(n3761) );
  XNOR U5356 ( .A(n3762), .B(n3761), .Z(\w1[3][112] ) );
  XNOR U5357 ( .A(\w3[2][106] ), .B(\w3[2][114] ), .Z(n4125) );
  XNOR U5358 ( .A(n4125), .B(key[497]), .Z(n3764) );
  XOR U5359 ( .A(\w3[2][105] ), .B(n4117), .Z(n3763) );
  XNOR U5360 ( .A(n3764), .B(n3763), .Z(\w1[3][113] ) );
  XNOR U5361 ( .A(\w3[2][107] ), .B(\w3[2][115] ), .Z(n3800) );
  XNOR U5362 ( .A(n3800), .B(key[498]), .Z(n3766) );
  XNOR U5363 ( .A(\w3[2][106] ), .B(n4122), .Z(n3765) );
  XNOR U5364 ( .A(n3766), .B(n3765), .Z(\w1[3][114] ) );
  XOR U5365 ( .A(\w3[2][116] ), .B(n3790), .Z(n3801) );
  XNOR U5366 ( .A(n3801), .B(key[499]), .Z(n3769) );
  XOR U5367 ( .A(\w3[2][107] ), .B(n3767), .Z(n3768) );
  XNOR U5368 ( .A(n3769), .B(n3768), .Z(\w1[3][115] ) );
  XOR U5369 ( .A(\w3[2][117] ), .B(n3790), .Z(n3804) );
  XNOR U5370 ( .A(n3804), .B(key[500]), .Z(n3772) );
  XOR U5371 ( .A(\w3[2][108] ), .B(n3770), .Z(n3771) );
  XNOR U5372 ( .A(n3772), .B(n3771), .Z(\w1[3][116] ) );
  XNOR U5373 ( .A(n3773), .B(key[501]), .Z(n3776) );
  XNOR U5374 ( .A(\w3[2][109] ), .B(n3774), .Z(n3775) );
  XNOR U5375 ( .A(n3776), .B(n3775), .Z(\w1[3][117] ) );
  XOR U5376 ( .A(\w3[2][119] ), .B(n3790), .Z(n3813) );
  XNOR U5377 ( .A(n3813), .B(key[502]), .Z(n3779) );
  XOR U5378 ( .A(\w3[2][110] ), .B(n3777), .Z(n3778) );
  XNOR U5379 ( .A(n3779), .B(n3778), .Z(\w1[3][118] ) );
  XOR U5380 ( .A(n3780), .B(key[503]), .Z(n3783) );
  XNOR U5381 ( .A(\w3[2][112] ), .B(n3781), .Z(n3782) );
  XNOR U5382 ( .A(n3783), .B(n3782), .Z(\w1[3][119] ) );
  XNOR U5383 ( .A(\w3[2][3] ), .B(\w3[2][27] ), .Z(n3877) );
  XNOR U5384 ( .A(n3837), .B(key[395]), .Z(n3785) );
  XNOR U5385 ( .A(\w3[2][0] ), .B(\w3[2][4] ), .Z(n3909) );
  XOR U5386 ( .A(\w3[2][19] ), .B(n3909), .Z(n3784) );
  XNOR U5387 ( .A(n3785), .B(n3784), .Z(\w1[3][11] ) );
  XNOR U5388 ( .A(n3786), .B(key[504]), .Z(n3788) );
  XNOR U5389 ( .A(\w3[2][121] ), .B(\w3[2][113] ), .Z(n3787) );
  XNOR U5390 ( .A(n3788), .B(n3787), .Z(n3789) );
  XNOR U5391 ( .A(n3790), .B(n3789), .Z(\w1[3][120] ) );
  XNOR U5392 ( .A(n4121), .B(key[505]), .Z(n3792) );
  XNOR U5393 ( .A(\w3[2][122] ), .B(\w3[2][114] ), .Z(n3791) );
  XNOR U5394 ( .A(n3792), .B(n3791), .Z(n3793) );
  XNOR U5395 ( .A(n3794), .B(n3793), .Z(\w1[3][121] ) );
  XNOR U5396 ( .A(n4125), .B(key[506]), .Z(n3796) );
  XNOR U5397 ( .A(\w3[2][115] ), .B(\w3[2][123] ), .Z(n3795) );
  XNOR U5398 ( .A(n3796), .B(n3795), .Z(n3797) );
  XOR U5399 ( .A(\w3[2][98] ), .B(n3797), .Z(\w1[3][122] ) );
  XOR U5400 ( .A(\w3[2][124] ), .B(n3798), .Z(n3799) );
  XOR U5401 ( .A(n3800), .B(n3799), .Z(n4129) );
  XOR U5402 ( .A(n4129), .B(key[507]), .Z(n3803) );
  XOR U5403 ( .A(\w3[2][99] ), .B(n3801), .Z(n3802) );
  XNOR U5404 ( .A(n3803), .B(n3802), .Z(\w1[3][123] ) );
  XNOR U5405 ( .A(n3804), .B(key[508]), .Z(n3808) );
  XNOR U5406 ( .A(n3806), .B(n3805), .Z(n3807) );
  XNOR U5407 ( .A(n3808), .B(n3807), .Z(\w1[3][124] ) );
  XOR U5408 ( .A(\w3[2][118] ), .B(key[509]), .Z(n3811) );
  XOR U5409 ( .A(n3809), .B(\w3[2][126] ), .Z(n3810) );
  XNOR U5410 ( .A(n3811), .B(n3810), .Z(n3812) );
  XOR U5411 ( .A(\w3[2][101] ), .B(n3812), .Z(\w1[3][125] ) );
  XNOR U5412 ( .A(n3813), .B(key[510]), .Z(n3816) );
  XOR U5413 ( .A(\w3[2][102] ), .B(n3814), .Z(n3815) );
  XNOR U5414 ( .A(n3816), .B(n3815), .Z(\w1[3][126] ) );
  XNOR U5415 ( .A(n4118), .B(key[511]), .Z(n3819) );
  XOR U5416 ( .A(\w3[2][103] ), .B(n3817), .Z(n3818) );
  XNOR U5417 ( .A(n3819), .B(n3818), .Z(\w1[3][127] ) );
  XOR U5418 ( .A(\w3[2][13] ), .B(\w3[2][28] ), .Z(n3821) );
  XNOR U5419 ( .A(\w3[2][8] ), .B(\w3[2][4] ), .Z(n3820) );
  XOR U5420 ( .A(n3821), .B(n3820), .Z(n3843) );
  XNOR U5421 ( .A(n3843), .B(key[396]), .Z(n3823) );
  XNOR U5422 ( .A(\w3[2][0] ), .B(\w3[2][5] ), .Z(n3944) );
  XOR U5423 ( .A(\w3[2][20] ), .B(n3944), .Z(n3822) );
  XNOR U5424 ( .A(n3823), .B(n3822), .Z(\w1[3][12] ) );
  IV U5425 ( .A(\w3[2][6] ), .Z(n3883) );
  XNOR U5426 ( .A(\w3[2][14] ), .B(n3883), .Z(n3825) );
  XNOR U5427 ( .A(\w3[2][5] ), .B(\w3[2][29] ), .Z(n3846) );
  XOR U5428 ( .A(n3846), .B(key[397]), .Z(n3824) );
  XNOR U5429 ( .A(n3825), .B(n3824), .Z(n3826) );
  XOR U5430 ( .A(\w3[2][21] ), .B(n3826), .Z(\w1[3][13] ) );
  IV U5431 ( .A(\w3[2][30] ), .Z(n4019) );
  XOR U5432 ( .A(\w3[2][6] ), .B(n4019), .Z(n3984) );
  XOR U5433 ( .A(\w3[2][8] ), .B(\w3[2][15] ), .Z(n3849) );
  XNOR U5434 ( .A(n3984), .B(n3849), .Z(n3847) );
  XOR U5435 ( .A(n3847), .B(key[398]), .Z(n3828) );
  XNOR U5436 ( .A(\w3[2][0] ), .B(\w3[2][7] ), .Z(n4020) );
  XOR U5437 ( .A(\w3[2][22] ), .B(n4020), .Z(n3827) );
  XNOR U5438 ( .A(n3828), .B(n3827), .Z(\w1[3][14] ) );
  XNOR U5439 ( .A(\w3[2][7] ), .B(\w3[2][31] ), .Z(n3848) );
  XNOR U5440 ( .A(n3848), .B(key[399]), .Z(n3830) );
  XOR U5441 ( .A(\w3[2][8] ), .B(\w3[2][0] ), .Z(n3852) );
  XNOR U5442 ( .A(\w3[2][23] ), .B(n3852), .Z(n3829) );
  XNOR U5443 ( .A(n3830), .B(n3829), .Z(\w1[3][15] ) );
  XNOR U5444 ( .A(\w3[2][17] ), .B(\w3[2][9] ), .Z(n3857) );
  XNOR U5445 ( .A(n3857), .B(key[400]), .Z(n3832) );
  XNOR U5446 ( .A(\w3[2][24] ), .B(n3852), .Z(n3831) );
  XNOR U5447 ( .A(n3832), .B(n3831), .Z(\w1[3][16] ) );
  XNOR U5448 ( .A(\w3[2][18] ), .B(\w3[2][10] ), .Z(n3876) );
  XNOR U5449 ( .A(n3876), .B(key[401]), .Z(n3834) );
  IV U5450 ( .A(\w3[2][9] ), .Z(n4088) );
  XNOR U5451 ( .A(n4136), .B(n4088), .Z(n3833) );
  XNOR U5452 ( .A(n3834), .B(n3833), .Z(\w1[3][17] ) );
  XNOR U5453 ( .A(\w3[2][11] ), .B(\w3[2][19] ), .Z(n3862) );
  XNOR U5454 ( .A(n3862), .B(key[402]), .Z(n3836) );
  XOR U5455 ( .A(n3840), .B(\w3[2][10] ), .Z(n3835) );
  XNOR U5456 ( .A(n3836), .B(n3835), .Z(\w1[3][18] ) );
  IV U5457 ( .A(\w3[2][16] ), .Z(n3856) );
  XOR U5458 ( .A(n3856), .B(\w3[2][20] ), .Z(n3863) );
  XNOR U5459 ( .A(n3863), .B(key[403]), .Z(n3839) );
  XOR U5460 ( .A(\w3[2][11] ), .B(n3837), .Z(n3838) );
  XNOR U5461 ( .A(n3839), .B(n3838), .Z(\w1[3][19] ) );
  XNOR U5462 ( .A(n3857), .B(key[385]), .Z(n3842) );
  XOR U5463 ( .A(\w3[2][25] ), .B(n3840), .Z(n3841) );
  XNOR U5464 ( .A(n3842), .B(n3841), .Z(\w1[3][1] ) );
  IV U5465 ( .A(\w3[2][21] ), .Z(n3871) );
  XOR U5466 ( .A(\w3[2][16] ), .B(n3871), .Z(n3868) );
  XNOR U5467 ( .A(n3868), .B(key[404]), .Z(n3845) );
  XOR U5468 ( .A(\w3[2][12] ), .B(n3843), .Z(n3844) );
  XNOR U5469 ( .A(n3845), .B(n3844), .Z(\w1[3][20] ) );
  IV U5470 ( .A(\w3[2][22] ), .Z(n3872) );
  XOR U5471 ( .A(\w3[2][14] ), .B(n3872), .Z(n3881) );
  XOR U5472 ( .A(n3856), .B(\w3[2][23] ), .Z(n3882) );
  XNOR U5473 ( .A(n3848), .B(key[407]), .Z(n3851) );
  XNOR U5474 ( .A(\w3[2][16] ), .B(n3849), .Z(n3850) );
  XNOR U5475 ( .A(n3851), .B(n3850), .Z(\w1[3][23] ) );
  XOR U5476 ( .A(\w3[2][17] ), .B(key[408]), .Z(n3854) );
  XNOR U5477 ( .A(\w3[2][25] ), .B(n3852), .Z(n3853) );
  XNOR U5478 ( .A(n3854), .B(n3853), .Z(n3855) );
  XNOR U5479 ( .A(n3856), .B(n3855), .Z(\w1[3][24] ) );
  XNOR U5480 ( .A(n3876), .B(key[410]), .Z(n3859) );
  XNOR U5481 ( .A(\w3[2][2] ), .B(\w3[2][19] ), .Z(n3858) );
  XNOR U5482 ( .A(n3859), .B(n3858), .Z(n3860) );
  XOR U5483 ( .A(\w3[2][27] ), .B(n3860), .Z(\w1[3][26] ) );
  XOR U5484 ( .A(n3880), .B(\w3[2][28] ), .Z(n3861) );
  XOR U5485 ( .A(n3862), .B(n3861), .Z(n3908) );
  XOR U5486 ( .A(n3908), .B(key[411]), .Z(n3865) );
  XOR U5487 ( .A(\w3[2][3] ), .B(n3863), .Z(n3864) );
  XNOR U5488 ( .A(n3865), .B(n3864), .Z(\w1[3][27] ) );
  XOR U5489 ( .A(\w3[2][20] ), .B(\w3[2][29] ), .Z(n3867) );
  XOR U5490 ( .A(n3880), .B(\w3[2][12] ), .Z(n3866) );
  XOR U5491 ( .A(n3867), .B(n3866), .Z(n3943) );
  XNOR U5492 ( .A(n3943), .B(key[412]), .Z(n3870) );
  XOR U5493 ( .A(\w3[2][4] ), .B(n3868), .Z(n3869) );
  XNOR U5494 ( .A(n3870), .B(n3869), .Z(\w1[3][28] ) );
  XOR U5495 ( .A(\w3[2][13] ), .B(n3871), .Z(n3983) );
  XNOR U5496 ( .A(n3983), .B(key[413]), .Z(n3874) );
  XNOR U5497 ( .A(n3872), .B(n4019), .Z(n3873) );
  XNOR U5498 ( .A(n3874), .B(n3873), .Z(n3875) );
  XOR U5499 ( .A(\w3[2][5] ), .B(n3875), .Z(\w1[3][29] ) );
  XNOR U5500 ( .A(n3876), .B(key[386]), .Z(n3879) );
  XOR U5501 ( .A(\w3[2][26] ), .B(n3877), .Z(n3878) );
  XNOR U5502 ( .A(n3879), .B(n3878), .Z(\w1[3][2] ) );
  XOR U5503 ( .A(n3880), .B(\w3[2][31] ), .Z(n4055) );
  XNOR U5504 ( .A(n3881), .B(n4055), .Z(n4018) );
  XNOR U5505 ( .A(n4018), .B(key[414]), .Z(n3885) );
  XNOR U5506 ( .A(n3883), .B(n3882), .Z(n3884) );
  XNOR U5507 ( .A(n3885), .B(n3884), .Z(\w1[3][30] ) );
  XNOR U5508 ( .A(\w3[2][15] ), .B(\w3[2][23] ), .Z(n4054) );
  XNOR U5509 ( .A(n4054), .B(key[415]), .Z(n3887) );
  XOR U5510 ( .A(n4089), .B(\w3[2][7] ), .Z(n3886) );
  XNOR U5511 ( .A(n3887), .B(n3886), .Z(\w1[3][31] ) );
  XNOR U5512 ( .A(\w3[2][48] ), .B(\w3[2][56] ), .Z(n4000) );
  XNOR U5513 ( .A(\w3[2][33] ), .B(\w3[2][57] ), .Z(n3940) );
  XNOR U5514 ( .A(\w3[2][40] ), .B(key[416]), .Z(n3888) );
  XNOR U5515 ( .A(n3940), .B(n3888), .Z(n3889) );
  XOR U5516 ( .A(n4000), .B(n3889), .Z(\w1[3][32] ) );
  XNOR U5517 ( .A(\w3[2][34] ), .B(\w3[2][58] ), .Z(n3948) );
  XNOR U5518 ( .A(\w3[2][41] ), .B(\w3[2][49] ), .Z(n3970) );
  XOR U5519 ( .A(n3970), .B(key[417]), .Z(n3890) );
  XNOR U5520 ( .A(n3948), .B(n3890), .Z(n3891) );
  XNOR U5521 ( .A(\w3[2][57] ), .B(n3891), .Z(\w1[3][33] ) );
  XNOR U5522 ( .A(n3918), .B(key[418]), .Z(n3893) );
  XNOR U5523 ( .A(\w3[2][42] ), .B(\w3[2][50] ), .Z(n3973) );
  XOR U5524 ( .A(\w3[2][58] ), .B(n3973), .Z(n3892) );
  XNOR U5525 ( .A(n3893), .B(n3892), .Z(\w1[3][34] ) );
  XOR U5526 ( .A(\w3[2][36] ), .B(\w3[2][32] ), .Z(n3920) );
  XOR U5527 ( .A(n3920), .B(key[419]), .Z(n3896) );
  IV U5528 ( .A(\w3[2][51] ), .Z(n3972) );
  XOR U5529 ( .A(\w3[2][43] ), .B(n3972), .Z(n3947) );
  XOR U5530 ( .A(\w3[2][56] ), .B(n3947), .Z(n3894) );
  XNOR U5531 ( .A(\w3[2][60] ), .B(n3894), .Z(n3979) );
  XNOR U5532 ( .A(\w3[2][59] ), .B(n3979), .Z(n3895) );
  XNOR U5533 ( .A(n3896), .B(n3895), .Z(\w1[3][35] ) );
  XOR U5534 ( .A(\w3[2][32] ), .B(\w3[2][37] ), .Z(n3926) );
  XOR U5535 ( .A(\w3[2][52] ), .B(\w3[2][61] ), .Z(n3898) );
  XNOR U5536 ( .A(\w3[2][56] ), .B(\w3[2][44] ), .Z(n3897) );
  XOR U5537 ( .A(n3898), .B(n3897), .Z(n3988) );
  XOR U5538 ( .A(n3988), .B(key[420]), .Z(n3899) );
  XOR U5539 ( .A(n3926), .B(n3899), .Z(n3900) );
  XNOR U5540 ( .A(\w3[2][60] ), .B(n3900), .Z(\w1[3][36] ) );
  XNOR U5541 ( .A(\w3[2][38] ), .B(\w3[2][62] ), .Z(n3932) );
  XNOR U5542 ( .A(n3932), .B(key[421]), .Z(n3902) );
  IV U5543 ( .A(\w3[2][53] ), .Z(n3952) );
  XOR U5544 ( .A(\w3[2][45] ), .B(n3952), .Z(n3991) );
  XOR U5545 ( .A(\w3[2][61] ), .B(n3991), .Z(n3901) );
  XNOR U5546 ( .A(n3902), .B(n3901), .Z(\w1[3][37] ) );
  XOR U5547 ( .A(\w3[2][32] ), .B(\w3[2][39] ), .Z(n3933) );
  XOR U5548 ( .A(n3933), .B(key[422]), .Z(n3904) );
  XNOR U5549 ( .A(\w3[2][56] ), .B(\w3[2][63] ), .Z(n3905) );
  XOR U5550 ( .A(\w3[2][46] ), .B(\w3[2][54] ), .Z(n3957) );
  XOR U5551 ( .A(n3905), .B(n3957), .Z(n3996) );
  XOR U5552 ( .A(\w3[2][62] ), .B(n3996), .Z(n3903) );
  XNOR U5553 ( .A(n3904), .B(n3903), .Z(\w1[3][38] ) );
  XNOR U5554 ( .A(\w3[2][47] ), .B(\w3[2][55] ), .Z(n3999) );
  XNOR U5555 ( .A(n3999), .B(key[423]), .Z(n3907) );
  XOR U5556 ( .A(\w3[2][32] ), .B(n3905), .Z(n3906) );
  XNOR U5557 ( .A(n3907), .B(n3906), .Z(\w1[3][39] ) );
  XOR U5558 ( .A(n3908), .B(key[387]), .Z(n3911) );
  XOR U5559 ( .A(n3909), .B(\w3[2][27] ), .Z(n3910) );
  XNOR U5560 ( .A(n3911), .B(n3910), .Z(\w1[3][3] ) );
  IV U5561 ( .A(\w3[2][33] ), .Z(n3971) );
  XOR U5562 ( .A(\w3[2][42] ), .B(key[425]), .Z(n3913) );
  IV U5563 ( .A(\w3[2][34] ), .Z(n3977) );
  XOR U5564 ( .A(\w3[2][49] ), .B(n3977), .Z(n3912) );
  XNOR U5565 ( .A(n3913), .B(n3912), .Z(n3914) );
  XNOR U5566 ( .A(n3914), .B(n3940), .Z(\w1[3][41] ) );
  XOR U5567 ( .A(\w3[2][43] ), .B(key[426]), .Z(n3916) );
  IV U5568 ( .A(\w3[2][35] ), .Z(n3980) );
  XOR U5569 ( .A(\w3[2][50] ), .B(n3980), .Z(n3915) );
  XNOR U5570 ( .A(n3916), .B(n3915), .Z(n3917) );
  XNOR U5571 ( .A(n3917), .B(n3948), .Z(\w1[3][42] ) );
  IV U5572 ( .A(\w3[2][40] ), .Z(n3923) );
  XNOR U5573 ( .A(n3923), .B(n3918), .Z(n3919) );
  XOR U5574 ( .A(\w3[2][44] ), .B(n3919), .Z(n3951) );
  XNOR U5575 ( .A(n3951), .B(key[427]), .Z(n3922) );
  XNOR U5576 ( .A(\w3[2][51] ), .B(n3920), .Z(n3921) );
  XNOR U5577 ( .A(n3922), .B(n3921), .Z(\w1[3][43] ) );
  XOR U5578 ( .A(\w3[2][36] ), .B(\w3[2][45] ), .Z(n3925) );
  XOR U5579 ( .A(n3923), .B(\w3[2][60] ), .Z(n3924) );
  XOR U5580 ( .A(n3925), .B(n3924), .Z(n3953) );
  XNOR U5581 ( .A(n3953), .B(key[428]), .Z(n3928) );
  XNOR U5582 ( .A(\w3[2][52] ), .B(n3926), .Z(n3927) );
  XNOR U5583 ( .A(n3928), .B(n3927), .Z(\w1[3][44] ) );
  XNOR U5584 ( .A(\w3[2][61] ), .B(\w3[2][37] ), .Z(n3956) );
  XNOR U5585 ( .A(n3956), .B(key[429]), .Z(n3930) );
  XNOR U5586 ( .A(\w3[2][38] ), .B(\w3[2][46] ), .Z(n3929) );
  XNOR U5587 ( .A(n3930), .B(n3929), .Z(n3931) );
  XOR U5588 ( .A(\w3[2][53] ), .B(n3931), .Z(\w1[3][45] ) );
  XOR U5589 ( .A(\w3[2][40] ), .B(\w3[2][47] ), .Z(n3962) );
  XOR U5590 ( .A(n3932), .B(n3962), .Z(n3958) );
  XNOR U5591 ( .A(n3958), .B(key[430]), .Z(n3935) );
  XNOR U5592 ( .A(\w3[2][54] ), .B(n3933), .Z(n3934) );
  XNOR U5593 ( .A(n3935), .B(n3934), .Z(\w1[3][46] ) );
  XOR U5594 ( .A(\w3[2][63] ), .B(\w3[2][39] ), .Z(n3961) );
  XOR U5595 ( .A(n3961), .B(key[431]), .Z(n3937) );
  XNOR U5596 ( .A(\w3[2][40] ), .B(\w3[2][32] ), .Z(n3965) );
  XOR U5597 ( .A(\w3[2][55] ), .B(n3965), .Z(n3936) );
  XNOR U5598 ( .A(n3937), .B(n3936), .Z(\w1[3][47] ) );
  XNOR U5599 ( .A(n3965), .B(key[432]), .Z(n3939) );
  XOR U5600 ( .A(\w3[2][56] ), .B(n3970), .Z(n3938) );
  XNOR U5601 ( .A(n3939), .B(n3938), .Z(\w1[3][48] ) );
  XNOR U5602 ( .A(n3973), .B(key[433]), .Z(n3942) );
  XOR U5603 ( .A(n3940), .B(\w3[2][41] ), .Z(n3941) );
  XNOR U5604 ( .A(n3942), .B(n3941), .Z(\w1[3][49] ) );
  XNOR U5605 ( .A(n3943), .B(key[388]), .Z(n3946) );
  XOR U5606 ( .A(n3944), .B(\w3[2][28] ), .Z(n3945) );
  XNOR U5607 ( .A(n3946), .B(n3945), .Z(\w1[3][4] ) );
  XNOR U5608 ( .A(n3947), .B(key[434]), .Z(n3950) );
  XOR U5609 ( .A(n3948), .B(\w3[2][42] ), .Z(n3949) );
  XNOR U5610 ( .A(n3950), .B(n3949), .Z(\w1[3][50] ) );
  IV U5611 ( .A(\w3[2][48] ), .Z(n3966) );
  XOR U5612 ( .A(n3966), .B(\w3[2][52] ), .Z(n3978) );
  XOR U5613 ( .A(\w3[2][48] ), .B(n3952), .Z(n3987) );
  XNOR U5614 ( .A(n3987), .B(key[436]), .Z(n3955) );
  XOR U5615 ( .A(\w3[2][44] ), .B(n3953), .Z(n3954) );
  XNOR U5616 ( .A(n3955), .B(n3954), .Z(\w1[3][52] ) );
  XOR U5617 ( .A(n3966), .B(\w3[2][55] ), .Z(n3995) );
  XNOR U5618 ( .A(n3995), .B(key[438]), .Z(n3960) );
  XOR U5619 ( .A(\w3[2][46] ), .B(n3958), .Z(n3959) );
  XNOR U5620 ( .A(n3960), .B(n3959), .Z(\w1[3][54] ) );
  XOR U5621 ( .A(n3961), .B(key[439]), .Z(n3964) );
  XNOR U5622 ( .A(\w3[2][48] ), .B(n3962), .Z(n3963) );
  XNOR U5623 ( .A(n3964), .B(n3963), .Z(\w1[3][55] ) );
  XNOR U5624 ( .A(n3965), .B(key[440]), .Z(n3968) );
  XOR U5625 ( .A(n3966), .B(\w3[2][49] ), .Z(n3967) );
  XNOR U5626 ( .A(n3968), .B(n3967), .Z(n3969) );
  XOR U5627 ( .A(\w3[2][57] ), .B(n3969), .Z(\w1[3][56] ) );
  XNOR U5628 ( .A(n3972), .B(key[442]), .Z(n3975) );
  XOR U5629 ( .A(n3973), .B(\w3[2][59] ), .Z(n3974) );
  XNOR U5630 ( .A(n3975), .B(n3974), .Z(n3976) );
  XNOR U5631 ( .A(n3977), .B(n3976), .Z(\w1[3][58] ) );
  XNOR U5632 ( .A(n3978), .B(key[443]), .Z(n3982) );
  XOR U5633 ( .A(n3980), .B(n3979), .Z(n3981) );
  XNOR U5634 ( .A(n3982), .B(n3981), .Z(\w1[3][59] ) );
  XNOR U5635 ( .A(n3983), .B(key[389]), .Z(n3986) );
  XOR U5636 ( .A(\w3[2][29] ), .B(n3984), .Z(n3985) );
  XNOR U5637 ( .A(n3986), .B(n3985), .Z(\w1[3][5] ) );
  XNOR U5638 ( .A(n3987), .B(key[444]), .Z(n3990) );
  XOR U5639 ( .A(\w3[2][36] ), .B(n3988), .Z(n3989) );
  XNOR U5640 ( .A(n3990), .B(n3989), .Z(\w1[3][60] ) );
  XOR U5641 ( .A(\w3[2][54] ), .B(key[445]), .Z(n3993) );
  XOR U5642 ( .A(n3991), .B(\w3[2][62] ), .Z(n3992) );
  XNOR U5643 ( .A(n3993), .B(n3992), .Z(n3994) );
  XOR U5644 ( .A(\w3[2][37] ), .B(n3994), .Z(\w1[3][61] ) );
  XNOR U5645 ( .A(n3995), .B(key[446]), .Z(n3998) );
  XOR U5646 ( .A(\w3[2][38] ), .B(n3996), .Z(n3997) );
  XNOR U5647 ( .A(n3998), .B(n3997), .Z(\w1[3][62] ) );
  XNOR U5648 ( .A(n3999), .B(key[447]), .Z(n4002) );
  XOR U5649 ( .A(n4000), .B(\w3[2][39] ), .Z(n4001) );
  XNOR U5650 ( .A(n4002), .B(n4001), .Z(\w1[3][63] ) );
  XNOR U5651 ( .A(\w3[2][80] ), .B(\w3[2][88] ), .Z(n4114) );
  XNOR U5652 ( .A(\w3[2][65] ), .B(\w3[2][89] ), .Z(n4060) );
  XNOR U5653 ( .A(\w3[2][72] ), .B(key[448]), .Z(n4003) );
  XNOR U5654 ( .A(n4060), .B(n4003), .Z(n4004) );
  XOR U5655 ( .A(n4114), .B(n4004), .Z(\w1[3][64] ) );
  XNOR U5656 ( .A(\w3[2][66] ), .B(\w3[2][90] ), .Z(n4064) );
  XNOR U5657 ( .A(\w3[2][73] ), .B(\w3[2][81] ), .Z(n4086) );
  XOR U5658 ( .A(n4086), .B(key[449]), .Z(n4005) );
  XNOR U5659 ( .A(n4064), .B(n4005), .Z(n4006) );
  XNOR U5660 ( .A(\w3[2][89] ), .B(n4006), .Z(\w1[3][65] ) );
  XNOR U5661 ( .A(n4034), .B(key[450]), .Z(n4008) );
  XNOR U5662 ( .A(\w3[2][74] ), .B(\w3[2][82] ), .Z(n4091) );
  XOR U5663 ( .A(\w3[2][90] ), .B(n4091), .Z(n4007) );
  XNOR U5664 ( .A(n4008), .B(n4007), .Z(\w1[3][66] ) );
  XOR U5665 ( .A(\w3[2][68] ), .B(\w3[2][64] ), .Z(n4036) );
  XOR U5666 ( .A(n4036), .B(key[451]), .Z(n4011) );
  IV U5667 ( .A(\w3[2][83] ), .Z(n4090) );
  XOR U5668 ( .A(\w3[2][75] ), .B(n4090), .Z(n4063) );
  XOR U5669 ( .A(\w3[2][88] ), .B(n4063), .Z(n4009) );
  XNOR U5670 ( .A(\w3[2][92] ), .B(n4009), .Z(n4097) );
  XNOR U5671 ( .A(\w3[2][91] ), .B(n4097), .Z(n4010) );
  XNOR U5672 ( .A(n4011), .B(n4010), .Z(\w1[3][67] ) );
  XOR U5673 ( .A(\w3[2][64] ), .B(\w3[2][69] ), .Z(n4042) );
  XOR U5674 ( .A(\w3[2][84] ), .B(\w3[2][93] ), .Z(n4013) );
  XNOR U5675 ( .A(\w3[2][88] ), .B(\w3[2][76] ), .Z(n4012) );
  XOR U5676 ( .A(n4013), .B(n4012), .Z(n4102) );
  XOR U5677 ( .A(n4102), .B(key[452]), .Z(n4014) );
  XOR U5678 ( .A(n4042), .B(n4014), .Z(n4015) );
  XNOR U5679 ( .A(\w3[2][92] ), .B(n4015), .Z(\w1[3][68] ) );
  XNOR U5680 ( .A(\w3[2][70] ), .B(\w3[2][94] ), .Z(n4048) );
  XNOR U5681 ( .A(n4048), .B(key[453]), .Z(n4017) );
  IV U5682 ( .A(\w3[2][85] ), .Z(n4068) );
  XOR U5683 ( .A(\w3[2][77] ), .B(n4068), .Z(n4105) );
  XOR U5684 ( .A(\w3[2][93] ), .B(n4105), .Z(n4016) );
  XNOR U5685 ( .A(n4017), .B(n4016), .Z(\w1[3][69] ) );
  XNOR U5686 ( .A(n4018), .B(key[390]), .Z(n4022) );
  XNOR U5687 ( .A(n4020), .B(n4019), .Z(n4021) );
  XNOR U5688 ( .A(n4022), .B(n4021), .Z(\w1[3][6] ) );
  XOR U5689 ( .A(\w3[2][64] ), .B(\w3[2][71] ), .Z(n4049) );
  XOR U5690 ( .A(n4049), .B(key[454]), .Z(n4024) );
  XNOR U5691 ( .A(\w3[2][88] ), .B(\w3[2][95] ), .Z(n4025) );
  XOR U5692 ( .A(\w3[2][78] ), .B(\w3[2][86] ), .Z(n4073) );
  XOR U5693 ( .A(n4025), .B(n4073), .Z(n4110) );
  XOR U5694 ( .A(\w3[2][94] ), .B(n4110), .Z(n4023) );
  XNOR U5695 ( .A(n4024), .B(n4023), .Z(\w1[3][70] ) );
  XNOR U5696 ( .A(\w3[2][79] ), .B(\w3[2][87] ), .Z(n4113) );
  XNOR U5697 ( .A(n4113), .B(key[455]), .Z(n4027) );
  XOR U5698 ( .A(\w3[2][64] ), .B(n4025), .Z(n4026) );
  XNOR U5699 ( .A(n4027), .B(n4026), .Z(\w1[3][71] ) );
  IV U5700 ( .A(\w3[2][65] ), .Z(n4087) );
  XOR U5701 ( .A(\w3[2][74] ), .B(key[457]), .Z(n4029) );
  IV U5702 ( .A(\w3[2][66] ), .Z(n4095) );
  XOR U5703 ( .A(\w3[2][81] ), .B(n4095), .Z(n4028) );
  XNOR U5704 ( .A(n4029), .B(n4028), .Z(n4030) );
  XNOR U5705 ( .A(n4030), .B(n4060), .Z(\w1[3][73] ) );
  XOR U5706 ( .A(\w3[2][75] ), .B(key[458]), .Z(n4032) );
  IV U5707 ( .A(\w3[2][67] ), .Z(n4098) );
  XOR U5708 ( .A(\w3[2][82] ), .B(n4098), .Z(n4031) );
  XNOR U5709 ( .A(n4032), .B(n4031), .Z(n4033) );
  XNOR U5710 ( .A(n4033), .B(n4064), .Z(\w1[3][74] ) );
  IV U5711 ( .A(\w3[2][72] ), .Z(n4039) );
  XNOR U5712 ( .A(n4039), .B(n4034), .Z(n4035) );
  XOR U5713 ( .A(\w3[2][76] ), .B(n4035), .Z(n4067) );
  XNOR U5714 ( .A(n4067), .B(key[459]), .Z(n4038) );
  XNOR U5715 ( .A(\w3[2][83] ), .B(n4036), .Z(n4037) );
  XNOR U5716 ( .A(n4038), .B(n4037), .Z(\w1[3][75] ) );
  XOR U5717 ( .A(\w3[2][68] ), .B(\w3[2][77] ), .Z(n4041) );
  XOR U5718 ( .A(n4039), .B(\w3[2][92] ), .Z(n4040) );
  XOR U5719 ( .A(n4041), .B(n4040), .Z(n4069) );
  XNOR U5720 ( .A(n4069), .B(key[460]), .Z(n4044) );
  XNOR U5721 ( .A(\w3[2][84] ), .B(n4042), .Z(n4043) );
  XNOR U5722 ( .A(n4044), .B(n4043), .Z(\w1[3][76] ) );
  XNOR U5723 ( .A(\w3[2][93] ), .B(\w3[2][69] ), .Z(n4072) );
  XNOR U5724 ( .A(n4072), .B(key[461]), .Z(n4046) );
  XNOR U5725 ( .A(\w3[2][70] ), .B(\w3[2][78] ), .Z(n4045) );
  XNOR U5726 ( .A(n4046), .B(n4045), .Z(n4047) );
  XOR U5727 ( .A(\w3[2][85] ), .B(n4047), .Z(\w1[3][77] ) );
  XOR U5728 ( .A(\w3[2][72] ), .B(\w3[2][79] ), .Z(n4078) );
  XOR U5729 ( .A(n4048), .B(n4078), .Z(n4074) );
  XNOR U5730 ( .A(n4074), .B(key[462]), .Z(n4051) );
  XNOR U5731 ( .A(\w3[2][86] ), .B(n4049), .Z(n4050) );
  XNOR U5732 ( .A(n4051), .B(n4050), .Z(\w1[3][78] ) );
  XOR U5733 ( .A(\w3[2][95] ), .B(\w3[2][71] ), .Z(n4077) );
  XOR U5734 ( .A(n4077), .B(key[463]), .Z(n4053) );
  XNOR U5735 ( .A(\w3[2][72] ), .B(\w3[2][64] ), .Z(n4081) );
  XOR U5736 ( .A(\w3[2][87] ), .B(n4081), .Z(n4052) );
  XNOR U5737 ( .A(n4053), .B(n4052), .Z(\w1[3][79] ) );
  XNOR U5738 ( .A(n4054), .B(key[391]), .Z(n4057) );
  XOR U5739 ( .A(\w3[2][0] ), .B(n4055), .Z(n4056) );
  XNOR U5740 ( .A(n4057), .B(n4056), .Z(\w1[3][7] ) );
  XNOR U5741 ( .A(n4081), .B(key[464]), .Z(n4059) );
  XOR U5742 ( .A(\w3[2][88] ), .B(n4086), .Z(n4058) );
  XNOR U5743 ( .A(n4059), .B(n4058), .Z(\w1[3][80] ) );
  XNOR U5744 ( .A(n4091), .B(key[465]), .Z(n4062) );
  XOR U5745 ( .A(n4060), .B(\w3[2][73] ), .Z(n4061) );
  XNOR U5746 ( .A(n4062), .B(n4061), .Z(\w1[3][81] ) );
  XNOR U5747 ( .A(n4063), .B(key[466]), .Z(n4066) );
  XOR U5748 ( .A(n4064), .B(\w3[2][74] ), .Z(n4065) );
  XNOR U5749 ( .A(n4066), .B(n4065), .Z(\w1[3][82] ) );
  IV U5750 ( .A(\w3[2][80] ), .Z(n4082) );
  XOR U5751 ( .A(n4082), .B(\w3[2][84] ), .Z(n4096) );
  XOR U5752 ( .A(\w3[2][80] ), .B(n4068), .Z(n4101) );
  XNOR U5753 ( .A(n4101), .B(key[468]), .Z(n4071) );
  XOR U5754 ( .A(\w3[2][76] ), .B(n4069), .Z(n4070) );
  XNOR U5755 ( .A(n4071), .B(n4070), .Z(\w1[3][84] ) );
  XOR U5756 ( .A(n4082), .B(\w3[2][87] ), .Z(n4109) );
  XNOR U5757 ( .A(n4109), .B(key[470]), .Z(n4076) );
  XOR U5758 ( .A(\w3[2][78] ), .B(n4074), .Z(n4075) );
  XNOR U5759 ( .A(n4076), .B(n4075), .Z(\w1[3][86] ) );
  XOR U5760 ( .A(n4077), .B(key[471]), .Z(n4080) );
  XNOR U5761 ( .A(\w3[2][80] ), .B(n4078), .Z(n4079) );
  XNOR U5762 ( .A(n4080), .B(n4079), .Z(\w1[3][87] ) );
  XNOR U5763 ( .A(n4081), .B(key[472]), .Z(n4084) );
  XOR U5764 ( .A(n4082), .B(\w3[2][81] ), .Z(n4083) );
  XNOR U5765 ( .A(n4084), .B(n4083), .Z(n4085) );
  XOR U5766 ( .A(\w3[2][89] ), .B(n4085), .Z(\w1[3][88] ) );
  XNOR U5767 ( .A(n4090), .B(key[474]), .Z(n4093) );
  XOR U5768 ( .A(n4091), .B(\w3[2][91] ), .Z(n4092) );
  XNOR U5769 ( .A(n4093), .B(n4092), .Z(n4094) );
  XNOR U5770 ( .A(n4095), .B(n4094), .Z(\w1[3][90] ) );
  XNOR U5771 ( .A(n4096), .B(key[475]), .Z(n4100) );
  XOR U5772 ( .A(n4098), .B(n4097), .Z(n4099) );
  XNOR U5773 ( .A(n4100), .B(n4099), .Z(\w1[3][91] ) );
  XNOR U5774 ( .A(n4101), .B(key[476]), .Z(n4104) );
  XOR U5775 ( .A(\w3[2][68] ), .B(n4102), .Z(n4103) );
  XNOR U5776 ( .A(n4104), .B(n4103), .Z(\w1[3][92] ) );
  XOR U5777 ( .A(\w3[2][86] ), .B(key[477]), .Z(n4107) );
  XOR U5778 ( .A(n4105), .B(\w3[2][94] ), .Z(n4106) );
  XNOR U5779 ( .A(n4107), .B(n4106), .Z(n4108) );
  XOR U5780 ( .A(\w3[2][69] ), .B(n4108), .Z(\w1[3][93] ) );
  XNOR U5781 ( .A(n4109), .B(key[478]), .Z(n4112) );
  XOR U5782 ( .A(\w3[2][70] ), .B(n4110), .Z(n4111) );
  XNOR U5783 ( .A(n4112), .B(n4111), .Z(\w1[3][94] ) );
  XNOR U5784 ( .A(n4113), .B(key[479]), .Z(n4116) );
  XOR U5785 ( .A(n4114), .B(\w3[2][71] ), .Z(n4115) );
  XNOR U5786 ( .A(n4116), .B(n4115), .Z(\w1[3][95] ) );
  XOR U5787 ( .A(\w3[2][104] ), .B(key[480]), .Z(n4120) );
  XNOR U5788 ( .A(n4118), .B(n4117), .Z(n4119) );
  XNOR U5789 ( .A(n4120), .B(n4119), .Z(\w1[3][96] ) );
  XNOR U5790 ( .A(n4121), .B(key[481]), .Z(n4124) );
  XNOR U5791 ( .A(\w3[2][121] ), .B(n4122), .Z(n4123) );
  XNOR U5792 ( .A(n4124), .B(n4123), .Z(\w1[3][97] ) );
  XNOR U5793 ( .A(n4125), .B(key[482]), .Z(n4128) );
  XOR U5794 ( .A(\w3[2][122] ), .B(n4126), .Z(n4127) );
  XNOR U5795 ( .A(n4128), .B(n4127), .Z(\w1[3][98] ) );
  XOR U5796 ( .A(n4129), .B(key[483]), .Z(n4132) );
  XOR U5797 ( .A(n4130), .B(\w3[2][123] ), .Z(n4131) );
  XNOR U5798 ( .A(n4132), .B(n4131), .Z(\w1[3][99] ) );
  XOR U5799 ( .A(\w3[2][10] ), .B(key[393]), .Z(n4134) );
  XNOR U5800 ( .A(\w3[2][2] ), .B(\w3[2][17] ), .Z(n4133) );
  XNOR U5801 ( .A(n4134), .B(n4133), .Z(n4135) );
  XNOR U5802 ( .A(n4136), .B(n4135), .Z(\w1[3][9] ) );
  XOR U5803 ( .A(key[512]), .B(\w0[4][0] ), .Z(\w1[4][0] ) );
  XOR U5804 ( .A(key[612]), .B(\w0[4][100] ), .Z(\w1[4][100] ) );
  XOR U5805 ( .A(key[613]), .B(\w0[4][101] ), .Z(\w1[4][101] ) );
  XOR U5806 ( .A(key[614]), .B(\w0[4][102] ), .Z(\w1[4][102] ) );
  XOR U5807 ( .A(key[615]), .B(\w0[4][103] ), .Z(\w1[4][103] ) );
  XOR U5808 ( .A(key[616]), .B(\w0[4][104] ), .Z(\w1[4][104] ) );
  XOR U5809 ( .A(key[617]), .B(\w0[4][105] ), .Z(\w1[4][105] ) );
  XOR U5810 ( .A(key[618]), .B(\w0[4][106] ), .Z(\w1[4][106] ) );
  XOR U5811 ( .A(key[619]), .B(\w0[4][107] ), .Z(\w1[4][107] ) );
  XOR U5812 ( .A(key[620]), .B(\w0[4][108] ), .Z(\w1[4][108] ) );
  XOR U5813 ( .A(key[621]), .B(\w0[4][109] ), .Z(\w1[4][109] ) );
  XOR U5814 ( .A(key[522]), .B(\w0[4][10] ), .Z(\w1[4][10] ) );
  XOR U5815 ( .A(key[622]), .B(\w0[4][110] ), .Z(\w1[4][110] ) );
  XOR U5816 ( .A(key[623]), .B(\w0[4][111] ), .Z(\w1[4][111] ) );
  XOR U5817 ( .A(key[624]), .B(\w0[4][112] ), .Z(\w1[4][112] ) );
  XOR U5818 ( .A(key[625]), .B(\w0[4][113] ), .Z(\w1[4][113] ) );
  XOR U5819 ( .A(key[626]), .B(\w0[4][114] ), .Z(\w1[4][114] ) );
  XOR U5820 ( .A(key[627]), .B(\w0[4][115] ), .Z(\w1[4][115] ) );
  XOR U5821 ( .A(key[628]), .B(\w0[4][116] ), .Z(\w1[4][116] ) );
  XOR U5822 ( .A(key[629]), .B(\w0[4][117] ), .Z(\w1[4][117] ) );
  XOR U5823 ( .A(key[630]), .B(\w0[4][118] ), .Z(\w1[4][118] ) );
  XOR U5824 ( .A(key[631]), .B(\w0[4][119] ), .Z(\w1[4][119] ) );
  XOR U5825 ( .A(key[523]), .B(\w0[4][11] ), .Z(\w1[4][11] ) );
  XOR U5826 ( .A(key[632]), .B(\w0[4][120] ), .Z(\w1[4][120] ) );
  XOR U5827 ( .A(key[633]), .B(\w0[4][121] ), .Z(\w1[4][121] ) );
  XOR U5828 ( .A(key[634]), .B(\w0[4][122] ), .Z(\w1[4][122] ) );
  XOR U5829 ( .A(key[635]), .B(\w0[4][123] ), .Z(\w1[4][123] ) );
  XOR U5830 ( .A(key[636]), .B(\w0[4][124] ), .Z(\w1[4][124] ) );
  XOR U5831 ( .A(key[637]), .B(\w0[4][125] ), .Z(\w1[4][125] ) );
  XOR U5832 ( .A(key[638]), .B(\w0[4][126] ), .Z(\w1[4][126] ) );
  XOR U5833 ( .A(key[639]), .B(\w0[4][127] ), .Z(\w1[4][127] ) );
  XOR U5834 ( .A(key[524]), .B(\w0[4][12] ), .Z(\w1[4][12] ) );
  XOR U5835 ( .A(key[525]), .B(\w0[4][13] ), .Z(\w1[4][13] ) );
  XOR U5836 ( .A(key[526]), .B(\w0[4][14] ), .Z(\w1[4][14] ) );
  XOR U5837 ( .A(key[527]), .B(\w0[4][15] ), .Z(\w1[4][15] ) );
  XOR U5838 ( .A(key[528]), .B(\w0[4][16] ), .Z(\w1[4][16] ) );
  XOR U5839 ( .A(key[529]), .B(\w0[4][17] ), .Z(\w1[4][17] ) );
  XOR U5840 ( .A(key[530]), .B(\w0[4][18] ), .Z(\w1[4][18] ) );
  XOR U5841 ( .A(key[531]), .B(\w0[4][19] ), .Z(\w1[4][19] ) );
  XOR U5842 ( .A(key[513]), .B(\w0[4][1] ), .Z(\w1[4][1] ) );
  XOR U5843 ( .A(key[532]), .B(\w0[4][20] ), .Z(\w1[4][20] ) );
  XOR U5844 ( .A(key[533]), .B(\w0[4][21] ), .Z(\w1[4][21] ) );
  XOR U5845 ( .A(key[534]), .B(\w0[4][22] ), .Z(\w1[4][22] ) );
  XOR U5846 ( .A(key[535]), .B(\w0[4][23] ), .Z(\w1[4][23] ) );
  XOR U5847 ( .A(key[536]), .B(\w0[4][24] ), .Z(\w1[4][24] ) );
  XOR U5848 ( .A(key[537]), .B(\w0[4][25] ), .Z(\w1[4][25] ) );
  XOR U5849 ( .A(key[538]), .B(\w0[4][26] ), .Z(\w1[4][26] ) );
  XOR U5850 ( .A(key[539]), .B(\w0[4][27] ), .Z(\w1[4][27] ) );
  XOR U5851 ( .A(key[540]), .B(\w0[4][28] ), .Z(\w1[4][28] ) );
  XOR U5852 ( .A(key[541]), .B(\w0[4][29] ), .Z(\w1[4][29] ) );
  XOR U5853 ( .A(key[514]), .B(\w0[4][2] ), .Z(\w1[4][2] ) );
  XOR U5854 ( .A(key[542]), .B(\w0[4][30] ), .Z(\w1[4][30] ) );
  XOR U5855 ( .A(key[543]), .B(\w0[4][31] ), .Z(\w1[4][31] ) );
  XOR U5856 ( .A(key[544]), .B(\w0[4][32] ), .Z(\w1[4][32] ) );
  XOR U5857 ( .A(key[545]), .B(\w0[4][33] ), .Z(\w1[4][33] ) );
  XOR U5858 ( .A(key[546]), .B(\w0[4][34] ), .Z(\w1[4][34] ) );
  XOR U5859 ( .A(key[547]), .B(\w0[4][35] ), .Z(\w1[4][35] ) );
  XOR U5860 ( .A(key[548]), .B(\w0[4][36] ), .Z(\w1[4][36] ) );
  XOR U5861 ( .A(key[549]), .B(\w0[4][37] ), .Z(\w1[4][37] ) );
  XOR U5862 ( .A(key[550]), .B(\w0[4][38] ), .Z(\w1[4][38] ) );
  XOR U5863 ( .A(key[551]), .B(\w0[4][39] ), .Z(\w1[4][39] ) );
  XOR U5864 ( .A(key[515]), .B(\w0[4][3] ), .Z(\w1[4][3] ) );
  XOR U5865 ( .A(key[552]), .B(\w0[4][40] ), .Z(\w1[4][40] ) );
  XOR U5866 ( .A(key[553]), .B(\w0[4][41] ), .Z(\w1[4][41] ) );
  XOR U5867 ( .A(key[554]), .B(\w0[4][42] ), .Z(\w1[4][42] ) );
  XOR U5868 ( .A(key[555]), .B(\w0[4][43] ), .Z(\w1[4][43] ) );
  XOR U5869 ( .A(key[556]), .B(\w0[4][44] ), .Z(\w1[4][44] ) );
  XOR U5870 ( .A(key[557]), .B(\w0[4][45] ), .Z(\w1[4][45] ) );
  XOR U5871 ( .A(key[558]), .B(\w0[4][46] ), .Z(\w1[4][46] ) );
  XOR U5872 ( .A(key[559]), .B(\w0[4][47] ), .Z(\w1[4][47] ) );
  XOR U5873 ( .A(key[560]), .B(\w0[4][48] ), .Z(\w1[4][48] ) );
  XOR U5874 ( .A(key[561]), .B(\w0[4][49] ), .Z(\w1[4][49] ) );
  XOR U5875 ( .A(key[516]), .B(\w0[4][4] ), .Z(\w1[4][4] ) );
  XOR U5876 ( .A(key[562]), .B(\w0[4][50] ), .Z(\w1[4][50] ) );
  XOR U5877 ( .A(key[563]), .B(\w0[4][51] ), .Z(\w1[4][51] ) );
  XOR U5878 ( .A(key[564]), .B(\w0[4][52] ), .Z(\w1[4][52] ) );
  XOR U5879 ( .A(key[565]), .B(\w0[4][53] ), .Z(\w1[4][53] ) );
  XOR U5880 ( .A(key[566]), .B(\w0[4][54] ), .Z(\w1[4][54] ) );
  XOR U5881 ( .A(key[567]), .B(\w0[4][55] ), .Z(\w1[4][55] ) );
  XOR U5882 ( .A(key[568]), .B(\w0[4][56] ), .Z(\w1[4][56] ) );
  XOR U5883 ( .A(key[569]), .B(\w0[4][57] ), .Z(\w1[4][57] ) );
  XOR U5884 ( .A(key[570]), .B(\w0[4][58] ), .Z(\w1[4][58] ) );
  XOR U5885 ( .A(key[571]), .B(\w0[4][59] ), .Z(\w1[4][59] ) );
  XOR U5886 ( .A(key[517]), .B(\w0[4][5] ), .Z(\w1[4][5] ) );
  XOR U5887 ( .A(key[572]), .B(\w0[4][60] ), .Z(\w1[4][60] ) );
  XOR U5888 ( .A(key[573]), .B(\w0[4][61] ), .Z(\w1[4][61] ) );
  XOR U5889 ( .A(key[574]), .B(\w0[4][62] ), .Z(\w1[4][62] ) );
  XOR U5890 ( .A(key[575]), .B(\w0[4][63] ), .Z(\w1[4][63] ) );
  XOR U5891 ( .A(key[576]), .B(\w0[4][64] ), .Z(\w1[4][64] ) );
  XOR U5892 ( .A(key[577]), .B(\w0[4][65] ), .Z(\w1[4][65] ) );
  XOR U5893 ( .A(key[578]), .B(\w0[4][66] ), .Z(\w1[4][66] ) );
  XOR U5894 ( .A(key[579]), .B(\w0[4][67] ), .Z(\w1[4][67] ) );
  XOR U5895 ( .A(key[580]), .B(\w0[4][68] ), .Z(\w1[4][68] ) );
  XOR U5896 ( .A(key[581]), .B(\w0[4][69] ), .Z(\w1[4][69] ) );
  XOR U5897 ( .A(key[518]), .B(\w0[4][6] ), .Z(\w1[4][6] ) );
  XOR U5898 ( .A(key[582]), .B(\w0[4][70] ), .Z(\w1[4][70] ) );
  XOR U5899 ( .A(key[583]), .B(\w0[4][71] ), .Z(\w1[4][71] ) );
  XOR U5900 ( .A(key[584]), .B(\w0[4][72] ), .Z(\w1[4][72] ) );
  XOR U5901 ( .A(key[585]), .B(\w0[4][73] ), .Z(\w1[4][73] ) );
  XOR U5902 ( .A(key[586]), .B(\w0[4][74] ), .Z(\w1[4][74] ) );
  XOR U5903 ( .A(key[587]), .B(\w0[4][75] ), .Z(\w1[4][75] ) );
  XOR U5904 ( .A(key[588]), .B(\w0[4][76] ), .Z(\w1[4][76] ) );
  XOR U5905 ( .A(key[589]), .B(\w0[4][77] ), .Z(\w1[4][77] ) );
  XOR U5906 ( .A(key[590]), .B(\w0[4][78] ), .Z(\w1[4][78] ) );
  XOR U5907 ( .A(key[591]), .B(\w0[4][79] ), .Z(\w1[4][79] ) );
  XOR U5908 ( .A(key[519]), .B(\w0[4][7] ), .Z(\w1[4][7] ) );
  XOR U5909 ( .A(key[592]), .B(\w0[4][80] ), .Z(\w1[4][80] ) );
  XOR U5910 ( .A(key[593]), .B(\w0[4][81] ), .Z(\w1[4][81] ) );
  XOR U5911 ( .A(key[594]), .B(\w0[4][82] ), .Z(\w1[4][82] ) );
  XOR U5912 ( .A(key[595]), .B(\w0[4][83] ), .Z(\w1[4][83] ) );
  XOR U5913 ( .A(key[596]), .B(\w0[4][84] ), .Z(\w1[4][84] ) );
  XOR U5914 ( .A(key[597]), .B(\w0[4][85] ), .Z(\w1[4][85] ) );
  XOR U5915 ( .A(key[598]), .B(\w0[4][86] ), .Z(\w1[4][86] ) );
  XOR U5916 ( .A(key[599]), .B(\w0[4][87] ), .Z(\w1[4][87] ) );
  XOR U5917 ( .A(key[600]), .B(\w0[4][88] ), .Z(\w1[4][88] ) );
  XOR U5918 ( .A(key[601]), .B(\w0[4][89] ), .Z(\w1[4][89] ) );
  XOR U5919 ( .A(key[520]), .B(\w0[4][8] ), .Z(\w1[4][8] ) );
  XOR U5920 ( .A(key[602]), .B(\w0[4][90] ), .Z(\w1[4][90] ) );
  XOR U5921 ( .A(key[603]), .B(\w0[4][91] ), .Z(\w1[4][91] ) );
  XOR U5922 ( .A(key[604]), .B(\w0[4][92] ), .Z(\w1[4][92] ) );
  XOR U5923 ( .A(key[605]), .B(\w0[4][93] ), .Z(\w1[4][93] ) );
  XOR U5924 ( .A(key[606]), .B(\w0[4][94] ), .Z(\w1[4][94] ) );
  XOR U5925 ( .A(key[607]), .B(\w0[4][95] ), .Z(\w1[4][95] ) );
  XOR U5926 ( .A(key[608]), .B(\w0[4][96] ), .Z(\w1[4][96] ) );
  XOR U5927 ( .A(key[609]), .B(\w0[4][97] ), .Z(\w1[4][97] ) );
  XOR U5928 ( .A(key[610]), .B(\w0[4][98] ), .Z(\w1[4][98] ) );
  XOR U5929 ( .A(key[611]), .B(\w0[4][99] ), .Z(\w1[4][99] ) );
  XOR U5930 ( .A(key[521]), .B(\w0[4][9] ), .Z(\w1[4][9] ) );
endmodule

