
module mult_N128_CC16 ( clk, rst, a, b, c );
  input [127:0] a;
  input [7:0] b;
  output [255:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345;
  wire   [255:0] sreg;

  DFF \sreg_reg[247]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(sreg[247]) );
  DFF \sreg_reg[246]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(sreg[246]) );
  DFF \sreg_reg[245]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(sreg[245]) );
  DFF \sreg_reg[244]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(sreg[244]) );
  DFF \sreg_reg[243]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(sreg[243]) );
  DFF \sreg_reg[242]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(sreg[242]) );
  DFF \sreg_reg[241]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(sreg[241]) );
  DFF \sreg_reg[240]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(sreg[240]) );
  DFF \sreg_reg[239]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(sreg[239]) );
  DFF \sreg_reg[238]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(sreg[238]) );
  DFF \sreg_reg[237]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(sreg[237]) );
  DFF \sreg_reg[236]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(sreg[236]) );
  DFF \sreg_reg[235]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(sreg[235]) );
  DFF \sreg_reg[234]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(sreg[234]) );
  DFF \sreg_reg[233]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(sreg[233]) );
  DFF \sreg_reg[232]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(sreg[232]) );
  DFF \sreg_reg[231]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(sreg[231]) );
  DFF \sreg_reg[230]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(sreg[230]) );
  DFF \sreg_reg[229]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(sreg[229]) );
  DFF \sreg_reg[228]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(sreg[228]) );
  DFF \sreg_reg[227]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(sreg[227]) );
  DFF \sreg_reg[226]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(sreg[226]) );
  DFF \sreg_reg[225]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(sreg[225]) );
  DFF \sreg_reg[224]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(sreg[224]) );
  DFF \sreg_reg[223]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(sreg[223]) );
  DFF \sreg_reg[222]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(sreg[222]) );
  DFF \sreg_reg[221]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(sreg[221]) );
  DFF \sreg_reg[220]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(sreg[220]) );
  DFF \sreg_reg[219]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(sreg[219]) );
  DFF \sreg_reg[218]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(sreg[218]) );
  DFF \sreg_reg[217]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(sreg[217]) );
  DFF \sreg_reg[216]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(sreg[216]) );
  DFF \sreg_reg[215]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(sreg[215]) );
  DFF \sreg_reg[214]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(sreg[214]) );
  DFF \sreg_reg[213]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(sreg[213]) );
  DFF \sreg_reg[212]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(sreg[212]) );
  DFF \sreg_reg[211]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(sreg[211]) );
  DFF \sreg_reg[210]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(sreg[210]) );
  DFF \sreg_reg[209]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(sreg[209]) );
  DFF \sreg_reg[208]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(sreg[208]) );
  DFF \sreg_reg[207]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(sreg[207]) );
  DFF \sreg_reg[206]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(sreg[206]) );
  DFF \sreg_reg[205]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(sreg[205]) );
  DFF \sreg_reg[204]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(sreg[204]) );
  DFF \sreg_reg[203]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(sreg[203]) );
  DFF \sreg_reg[202]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(sreg[202]) );
  DFF \sreg_reg[201]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(sreg[201]) );
  DFF \sreg_reg[200]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(sreg[200]) );
  DFF \sreg_reg[199]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(sreg[199]) );
  DFF \sreg_reg[198]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(sreg[198]) );
  DFF \sreg_reg[197]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(sreg[197]) );
  DFF \sreg_reg[196]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(sreg[196]) );
  DFF \sreg_reg[195]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(sreg[195]) );
  DFF \sreg_reg[194]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(sreg[194]) );
  DFF \sreg_reg[193]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(sreg[193]) );
  DFF \sreg_reg[192]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(sreg[192]) );
  DFF \sreg_reg[191]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(sreg[191]) );
  DFF \sreg_reg[190]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(sreg[190]) );
  DFF \sreg_reg[189]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(sreg[189]) );
  DFF \sreg_reg[188]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(sreg[188]) );
  DFF \sreg_reg[187]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(sreg[187]) );
  DFF \sreg_reg[186]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(sreg[186]) );
  DFF \sreg_reg[185]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(sreg[185]) );
  DFF \sreg_reg[184]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(sreg[184]) );
  DFF \sreg_reg[183]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(sreg[183]) );
  DFF \sreg_reg[182]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(sreg[182]) );
  DFF \sreg_reg[181]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(sreg[181]) );
  DFF \sreg_reg[180]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(sreg[180]) );
  DFF \sreg_reg[179]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(sreg[179]) );
  DFF \sreg_reg[178]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(sreg[178]) );
  DFF \sreg_reg[177]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(sreg[177]) );
  DFF \sreg_reg[176]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(sreg[176]) );
  DFF \sreg_reg[175]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(sreg[175]) );
  DFF \sreg_reg[174]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(sreg[174]) );
  DFF \sreg_reg[173]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(sreg[173]) );
  DFF \sreg_reg[172]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(sreg[172]) );
  DFF \sreg_reg[171]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(sreg[171]) );
  DFF \sreg_reg[170]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(sreg[170]) );
  DFF \sreg_reg[169]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(sreg[169]) );
  DFF \sreg_reg[168]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(sreg[168]) );
  DFF \sreg_reg[167]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(sreg[167]) );
  DFF \sreg_reg[166]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(sreg[166]) );
  DFF \sreg_reg[165]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(sreg[165]) );
  DFF \sreg_reg[164]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(sreg[164]) );
  DFF \sreg_reg[163]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(sreg[163]) );
  DFF \sreg_reg[162]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(sreg[162]) );
  DFF \sreg_reg[161]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(sreg[161]) );
  DFF \sreg_reg[160]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(sreg[160]) );
  DFF \sreg_reg[159]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(sreg[159]) );
  DFF \sreg_reg[158]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(sreg[158]) );
  DFF \sreg_reg[157]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(sreg[157]) );
  DFF \sreg_reg[156]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(sreg[156]) );
  DFF \sreg_reg[155]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(sreg[155]) );
  DFF \sreg_reg[154]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(sreg[154]) );
  DFF \sreg_reg[153]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(sreg[153]) );
  DFF \sreg_reg[152]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(sreg[152]) );
  DFF \sreg_reg[151]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(sreg[151]) );
  DFF \sreg_reg[150]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(sreg[150]) );
  DFF \sreg_reg[149]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(sreg[149]) );
  DFF \sreg_reg[148]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(sreg[148]) );
  DFF \sreg_reg[147]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(sreg[147]) );
  DFF \sreg_reg[146]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(sreg[146]) );
  DFF \sreg_reg[145]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(sreg[145]) );
  DFF \sreg_reg[144]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(sreg[144]) );
  DFF \sreg_reg[143]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(sreg[143]) );
  DFF \sreg_reg[142]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(sreg[142]) );
  DFF \sreg_reg[141]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(sreg[141]) );
  DFF \sreg_reg[140]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(sreg[140]) );
  DFF \sreg_reg[139]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(sreg[139]) );
  DFF \sreg_reg[138]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(sreg[138]) );
  DFF \sreg_reg[137]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(sreg[137]) );
  DFF \sreg_reg[136]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(sreg[136]) );
  DFF \sreg_reg[135]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(sreg[135]) );
  DFF \sreg_reg[134]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(sreg[134]) );
  DFF \sreg_reg[133]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(sreg[133]) );
  DFF \sreg_reg[132]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(sreg[132]) );
  DFF \sreg_reg[131]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(sreg[131]) );
  DFF \sreg_reg[130]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(sreg[130]) );
  DFF \sreg_reg[129]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(sreg[129]) );
  DFF \sreg_reg[128]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(sreg[128]) );
  DFF \sreg_reg[127]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(sreg[127]) );
  DFF \sreg_reg[126]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(sreg[126]) );
  DFF \sreg_reg[125]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(sreg[125]) );
  DFF \sreg_reg[124]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(sreg[124]) );
  DFF \sreg_reg[123]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(sreg[123]) );
  DFF \sreg_reg[122]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(sreg[122]) );
  DFF \sreg_reg[121]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(sreg[121]) );
  DFF \sreg_reg[120]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(sreg[120]) );
  DFF \sreg_reg[119]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[118]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[117]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[116]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[115]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[114]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[113]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[112]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[111]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[110]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[109]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[108]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[107]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[106]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[105]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[104]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[103]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[102]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[101]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[100]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[99]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[98]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[97]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[96]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[95]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[94]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[93]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[92]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[91]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[90]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[89]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[88]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[87]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[86]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[85]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[84]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[83]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[82]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[81]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[80]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[79]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[78]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[77]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[76]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[75]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[74]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[73]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[72]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[71]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[70]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[69]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[68]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[67]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[66]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[65]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[64]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[63]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[62]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[0]) );
  NAND U11 ( .A(n1832), .B(n1831), .Z(n1) );
  NAND U12 ( .A(n1829), .B(n1830), .Z(n2) );
  NAND U13 ( .A(n1), .B(n2), .Z(n1839) );
  NAND U14 ( .A(n2454), .B(n2453), .Z(n3) );
  NAND U15 ( .A(n2451), .B(n2452), .Z(n4) );
  NAND U16 ( .A(n3), .B(n4), .Z(n2461) );
  NAND U17 ( .A(n2647), .B(n2648), .Z(n5) );
  NANDN U18 ( .A(n2646), .B(n2645), .Z(n6) );
  NAND U19 ( .A(n5), .B(n6), .Z(n2655) );
  NAND U20 ( .A(n3231), .B(n3230), .Z(n7) );
  NAND U21 ( .A(n3228), .B(n3229), .Z(n8) );
  NAND U22 ( .A(n7), .B(n8), .Z(n3238) );
  NAND U23 ( .A(n4204), .B(n4205), .Z(n9) );
  NANDN U24 ( .A(n4203), .B(n4202), .Z(n10) );
  NAND U25 ( .A(n9), .B(n10), .Z(n4212) );
  NAND U26 ( .A(n4476), .B(n4475), .Z(n11) );
  NAND U27 ( .A(n4473), .B(n4474), .Z(n12) );
  NAND U28 ( .A(n11), .B(n12), .Z(n4483) );
  NAND U29 ( .A(n2026), .B(n2027), .Z(n13) );
  NANDN U30 ( .A(n2025), .B(n2024), .Z(n14) );
  NAND U31 ( .A(n13), .B(n14), .Z(n2034) );
  XOR U32 ( .A(n345), .B(n344), .Z(n15) );
  NANDN U33 ( .A(n343), .B(n15), .Z(n16) );
  NAND U34 ( .A(n345), .B(n344), .Z(n17) );
  AND U35 ( .A(n16), .B(n17), .Z(n372) );
  NAND U36 ( .A(n594), .B(n595), .Z(n18) );
  NANDN U37 ( .A(n593), .B(n592), .Z(n19) );
  NAND U38 ( .A(n18), .B(n19), .Z(n634) );
  NAND U39 ( .A(n711), .B(n712), .Z(n20) );
  NANDN U40 ( .A(n710), .B(n709), .Z(n21) );
  NAND U41 ( .A(n20), .B(n21), .Z(n751) );
  NAND U42 ( .A(n828), .B(n829), .Z(n22) );
  NANDN U43 ( .A(n827), .B(n826), .Z(n23) );
  NAND U44 ( .A(n22), .B(n23), .Z(n868) );
  NAND U45 ( .A(n945), .B(n946), .Z(n24) );
  NANDN U46 ( .A(n944), .B(n943), .Z(n25) );
  NAND U47 ( .A(n24), .B(n25), .Z(n985) );
  NAND U48 ( .A(n1062), .B(n1063), .Z(n26) );
  NANDN U49 ( .A(n1061), .B(n1060), .Z(n27) );
  NAND U50 ( .A(n26), .B(n27), .Z(n1102) );
  NAND U51 ( .A(n1179), .B(n1180), .Z(n28) );
  NANDN U52 ( .A(n1178), .B(n1177), .Z(n29) );
  NAND U53 ( .A(n28), .B(n29), .Z(n1219) );
  NAND U54 ( .A(n1296), .B(n1297), .Z(n30) );
  NANDN U55 ( .A(n1295), .B(n1294), .Z(n31) );
  NAND U56 ( .A(n30), .B(n31), .Z(n1336) );
  NAND U57 ( .A(n1413), .B(n1414), .Z(n32) );
  NANDN U58 ( .A(n1412), .B(n1411), .Z(n33) );
  NAND U59 ( .A(n32), .B(n33), .Z(n1453) );
  NAND U60 ( .A(n1530), .B(n1531), .Z(n34) );
  NANDN U61 ( .A(n1529), .B(n1528), .Z(n35) );
  NAND U62 ( .A(n34), .B(n35), .Z(n1570) );
  NAND U63 ( .A(n1647), .B(n1648), .Z(n36) );
  NANDN U64 ( .A(n1646), .B(n1645), .Z(n37) );
  NAND U65 ( .A(n36), .B(n37), .Z(n1687) );
  NAND U66 ( .A(n1764), .B(n1765), .Z(n38) );
  NANDN U67 ( .A(n1763), .B(n1762), .Z(n39) );
  NAND U68 ( .A(n38), .B(n39), .Z(n1804) );
  NAND U69 ( .A(n1879), .B(n1880), .Z(n40) );
  NANDN U70 ( .A(n1878), .B(n1877), .Z(n41) );
  NAND U71 ( .A(n40), .B(n41), .Z(n1919) );
  NAND U72 ( .A(n2113), .B(n2114), .Z(n42) );
  NANDN U73 ( .A(n2112), .B(n2111), .Z(n43) );
  NAND U74 ( .A(n42), .B(n43), .Z(n2153) );
  NAND U75 ( .A(n2230), .B(n2231), .Z(n44) );
  NANDN U76 ( .A(n2229), .B(n2228), .Z(n45) );
  NAND U77 ( .A(n44), .B(n45), .Z(n2270) );
  NAND U78 ( .A(n2347), .B(n2348), .Z(n46) );
  NANDN U79 ( .A(n2346), .B(n2345), .Z(n47) );
  NAND U80 ( .A(n46), .B(n47), .Z(n2387) );
  NAND U81 ( .A(n2462), .B(n2463), .Z(n48) );
  NANDN U82 ( .A(n2461), .B(n2460), .Z(n49) );
  NAND U83 ( .A(n48), .B(n49), .Z(n2502) );
  NAND U84 ( .A(n2580), .B(n2581), .Z(n50) );
  NANDN U85 ( .A(n2579), .B(n2578), .Z(n51) );
  NAND U86 ( .A(n50), .B(n51), .Z(n2620) );
  NAND U87 ( .A(n2695), .B(n2696), .Z(n52) );
  NANDN U88 ( .A(n2694), .B(n2693), .Z(n53) );
  NAND U89 ( .A(n52), .B(n53), .Z(n2735) );
  NAND U90 ( .A(n2812), .B(n2813), .Z(n54) );
  NANDN U91 ( .A(n2811), .B(n2810), .Z(n55) );
  NAND U92 ( .A(n54), .B(n55), .Z(n2852) );
  NAND U93 ( .A(n2929), .B(n2930), .Z(n56) );
  NANDN U94 ( .A(n2928), .B(n2927), .Z(n57) );
  NAND U95 ( .A(n56), .B(n57), .Z(n2969) );
  NAND U96 ( .A(n3046), .B(n3047), .Z(n58) );
  NANDN U97 ( .A(n3045), .B(n3044), .Z(n59) );
  NAND U98 ( .A(n58), .B(n59), .Z(n3086) );
  NAND U99 ( .A(n3163), .B(n3164), .Z(n60) );
  NANDN U100 ( .A(n3162), .B(n3161), .Z(n61) );
  NAND U101 ( .A(n60), .B(n61), .Z(n3203) );
  NAND U102 ( .A(n3278), .B(n3279), .Z(n62) );
  NANDN U103 ( .A(n3277), .B(n3276), .Z(n63) );
  NAND U104 ( .A(n62), .B(n63), .Z(n3318) );
  NAND U105 ( .A(n3395), .B(n3396), .Z(n64) );
  NANDN U106 ( .A(n3394), .B(n3393), .Z(n65) );
  NAND U107 ( .A(n64), .B(n65), .Z(n3435) );
  NAND U108 ( .A(n3512), .B(n3513), .Z(n66) );
  NANDN U109 ( .A(n3511), .B(n3510), .Z(n67) );
  NAND U110 ( .A(n66), .B(n67), .Z(n3552) );
  NAND U111 ( .A(n3629), .B(n3630), .Z(n68) );
  NANDN U112 ( .A(n3628), .B(n3627), .Z(n69) );
  NAND U113 ( .A(n68), .B(n69), .Z(n3669) );
  NAND U114 ( .A(n3746), .B(n3747), .Z(n70) );
  NANDN U115 ( .A(n3745), .B(n3744), .Z(n71) );
  NAND U116 ( .A(n70), .B(n71), .Z(n3786) );
  NAND U117 ( .A(n3863), .B(n3864), .Z(n72) );
  NANDN U118 ( .A(n3862), .B(n3861), .Z(n73) );
  NAND U119 ( .A(n72), .B(n73), .Z(n3903) );
  NAND U120 ( .A(n3980), .B(n3981), .Z(n74) );
  NANDN U121 ( .A(n3979), .B(n3978), .Z(n75) );
  NAND U122 ( .A(n74), .B(n75), .Z(n4020) );
  NAND U123 ( .A(n4097), .B(n4098), .Z(n76) );
  NANDN U124 ( .A(n4096), .B(n4095), .Z(n77) );
  NAND U125 ( .A(n76), .B(n77), .Z(n4138) );
  NAND U126 ( .A(n4213), .B(n4214), .Z(n78) );
  NANDN U127 ( .A(n4212), .B(n4211), .Z(n79) );
  NAND U128 ( .A(n78), .B(n79), .Z(n4253) );
  NAND U129 ( .A(n4330), .B(n4331), .Z(n80) );
  NANDN U130 ( .A(n4329), .B(n4328), .Z(n81) );
  NAND U131 ( .A(n80), .B(n81), .Z(n4370) );
  NAND U132 ( .A(n4447), .B(n4448), .Z(n82) );
  NANDN U133 ( .A(n4446), .B(n4445), .Z(n83) );
  NAND U134 ( .A(n82), .B(n83), .Z(n4485) );
  NAND U135 ( .A(n4562), .B(n4563), .Z(n84) );
  NANDN U136 ( .A(n4561), .B(n4560), .Z(n85) );
  NAND U137 ( .A(n84), .B(n85), .Z(n4602) );
  NAND U138 ( .A(n4679), .B(n4680), .Z(n86) );
  NANDN U139 ( .A(n4678), .B(n4677), .Z(n87) );
  NAND U140 ( .A(n86), .B(n87), .Z(n4719) );
  NAND U141 ( .A(n4796), .B(n4797), .Z(n88) );
  NANDN U142 ( .A(n4795), .B(n4794), .Z(n89) );
  NAND U143 ( .A(n88), .B(n89), .Z(n4836) );
  NAND U144 ( .A(n4913), .B(n4914), .Z(n90) );
  NANDN U145 ( .A(n4912), .B(n4911), .Z(n91) );
  NAND U146 ( .A(n90), .B(n91), .Z(n4953) );
  NAND U147 ( .A(n5030), .B(n5031), .Z(n92) );
  NANDN U148 ( .A(n5029), .B(n5028), .Z(n93) );
  NAND U149 ( .A(n92), .B(n93), .Z(n5070) );
  NAND U150 ( .A(n5225), .B(n5224), .Z(n94) );
  XOR U151 ( .A(n5224), .B(n5225), .Z(n95) );
  NAND U152 ( .A(n95), .B(n5223), .Z(n96) );
  NAND U153 ( .A(n94), .B(n96), .Z(n5255) );
  XOR U154 ( .A(n5319), .B(n5320), .Z(n5330) );
  NANDN U155 ( .A(a[0]), .B(n294), .Z(n97) );
  XNOR U156 ( .A(n294), .B(a[0]), .Z(n98) );
  NAND U157 ( .A(n98), .B(n5336), .Z(n99) );
  NAND U158 ( .A(n97), .B(n99), .Z(n100) );
  AND U159 ( .A(b[7]), .B(n100), .Z(n448) );
  NOR U160 ( .A(n376), .B(n377), .Z(n423) );
  NAND U161 ( .A(n633), .B(n634), .Z(n101) );
  NANDN U162 ( .A(n632), .B(n631), .Z(n102) );
  NAND U163 ( .A(n101), .B(n102), .Z(n673) );
  NAND U164 ( .A(n750), .B(n751), .Z(n103) );
  NANDN U165 ( .A(n749), .B(n748), .Z(n104) );
  NAND U166 ( .A(n103), .B(n104), .Z(n790) );
  NAND U167 ( .A(n867), .B(n868), .Z(n105) );
  NANDN U168 ( .A(n866), .B(n865), .Z(n106) );
  NAND U169 ( .A(n105), .B(n106), .Z(n907) );
  NAND U170 ( .A(n984), .B(n985), .Z(n107) );
  NANDN U171 ( .A(n983), .B(n982), .Z(n108) );
  NAND U172 ( .A(n107), .B(n108), .Z(n1024) );
  NAND U173 ( .A(n1101), .B(n1102), .Z(n109) );
  NANDN U174 ( .A(n1100), .B(n1099), .Z(n110) );
  NAND U175 ( .A(n109), .B(n110), .Z(n1141) );
  NAND U176 ( .A(n1218), .B(n1219), .Z(n111) );
  NANDN U177 ( .A(n1217), .B(n1216), .Z(n112) );
  NAND U178 ( .A(n111), .B(n112), .Z(n1258) );
  NAND U179 ( .A(n1335), .B(n1336), .Z(n113) );
  NANDN U180 ( .A(n1334), .B(n1333), .Z(n114) );
  NAND U181 ( .A(n113), .B(n114), .Z(n1375) );
  NAND U182 ( .A(n1452), .B(n1453), .Z(n115) );
  NANDN U183 ( .A(n1451), .B(n1450), .Z(n116) );
  NAND U184 ( .A(n115), .B(n116), .Z(n1492) );
  NAND U185 ( .A(n1569), .B(n1570), .Z(n117) );
  NANDN U186 ( .A(n1568), .B(n1567), .Z(n118) );
  NAND U187 ( .A(n117), .B(n118), .Z(n1609) );
  NAND U188 ( .A(n1686), .B(n1687), .Z(n119) );
  NANDN U189 ( .A(n1685), .B(n1684), .Z(n120) );
  NAND U190 ( .A(n119), .B(n120), .Z(n1726) );
  NAND U191 ( .A(n1803), .B(n1804), .Z(n121) );
  NANDN U192 ( .A(n1802), .B(n1801), .Z(n122) );
  NAND U193 ( .A(n121), .B(n122), .Z(n1841) );
  NAND U194 ( .A(n1918), .B(n1919), .Z(n123) );
  NANDN U195 ( .A(n1917), .B(n1916), .Z(n124) );
  NAND U196 ( .A(n123), .B(n124), .Z(n1958) );
  NAND U197 ( .A(n2035), .B(n2036), .Z(n125) );
  NANDN U198 ( .A(n2034), .B(n2033), .Z(n126) );
  NAND U199 ( .A(n125), .B(n126), .Z(n2075) );
  NAND U200 ( .A(n2152), .B(n2153), .Z(n127) );
  NANDN U201 ( .A(n2151), .B(n2150), .Z(n128) );
  NAND U202 ( .A(n127), .B(n128), .Z(n2192) );
  NAND U203 ( .A(n2269), .B(n2270), .Z(n129) );
  NANDN U204 ( .A(n2268), .B(n2267), .Z(n130) );
  NAND U205 ( .A(n129), .B(n130), .Z(n2309) );
  NAND U206 ( .A(n2386), .B(n2387), .Z(n131) );
  NANDN U207 ( .A(n2385), .B(n2384), .Z(n132) );
  NAND U208 ( .A(n131), .B(n132), .Z(n2426) );
  NAND U209 ( .A(n2501), .B(n2502), .Z(n133) );
  NANDN U210 ( .A(n2500), .B(n2499), .Z(n134) );
  NAND U211 ( .A(n133), .B(n134), .Z(n2541) );
  NAND U212 ( .A(n2619), .B(n2620), .Z(n135) );
  NANDN U213 ( .A(n2618), .B(n2617), .Z(n136) );
  NAND U214 ( .A(n135), .B(n136), .Z(n2657) );
  NAND U215 ( .A(n2734), .B(n2735), .Z(n137) );
  NANDN U216 ( .A(n2733), .B(n2732), .Z(n138) );
  NAND U217 ( .A(n137), .B(n138), .Z(n2774) );
  NAND U218 ( .A(n2851), .B(n2852), .Z(n139) );
  NANDN U219 ( .A(n2850), .B(n2849), .Z(n140) );
  NAND U220 ( .A(n139), .B(n140), .Z(n2891) );
  NAND U221 ( .A(n2968), .B(n2969), .Z(n141) );
  NANDN U222 ( .A(n2967), .B(n2966), .Z(n142) );
  NAND U223 ( .A(n141), .B(n142), .Z(n3008) );
  NAND U224 ( .A(n3085), .B(n3086), .Z(n143) );
  NANDN U225 ( .A(n3084), .B(n3083), .Z(n144) );
  NAND U226 ( .A(n143), .B(n144), .Z(n3125) );
  NAND U227 ( .A(n3202), .B(n3203), .Z(n145) );
  NANDN U228 ( .A(n3201), .B(n3200), .Z(n146) );
  NAND U229 ( .A(n145), .B(n146), .Z(n3240) );
  NAND U230 ( .A(n3317), .B(n3318), .Z(n147) );
  NANDN U231 ( .A(n3316), .B(n3315), .Z(n148) );
  NAND U232 ( .A(n147), .B(n148), .Z(n3357) );
  NAND U233 ( .A(n3434), .B(n3435), .Z(n149) );
  NANDN U234 ( .A(n3433), .B(n3432), .Z(n150) );
  NAND U235 ( .A(n149), .B(n150), .Z(n3474) );
  NAND U236 ( .A(n3551), .B(n3552), .Z(n151) );
  NANDN U237 ( .A(n3550), .B(n3549), .Z(n152) );
  NAND U238 ( .A(n151), .B(n152), .Z(n3591) );
  NAND U239 ( .A(n3668), .B(n3669), .Z(n153) );
  NANDN U240 ( .A(n3667), .B(n3666), .Z(n154) );
  NAND U241 ( .A(n153), .B(n154), .Z(n3708) );
  NAND U242 ( .A(n3785), .B(n3786), .Z(n155) );
  NANDN U243 ( .A(n3784), .B(n3783), .Z(n156) );
  NAND U244 ( .A(n155), .B(n156), .Z(n3825) );
  NAND U245 ( .A(n3902), .B(n3903), .Z(n157) );
  NANDN U246 ( .A(n3901), .B(n3900), .Z(n158) );
  NAND U247 ( .A(n157), .B(n158), .Z(n3942) );
  NAND U248 ( .A(n4019), .B(n4020), .Z(n159) );
  NANDN U249 ( .A(n4018), .B(n4017), .Z(n160) );
  NAND U250 ( .A(n159), .B(n160), .Z(n4059) );
  NAND U251 ( .A(n4137), .B(n4138), .Z(n161) );
  NANDN U252 ( .A(n4136), .B(n4135), .Z(n162) );
  NAND U253 ( .A(n161), .B(n162), .Z(n4177) );
  NAND U254 ( .A(n4252), .B(n4253), .Z(n163) );
  NANDN U255 ( .A(n4251), .B(n4250), .Z(n164) );
  NAND U256 ( .A(n163), .B(n164), .Z(n4292) );
  NAND U257 ( .A(n4369), .B(n4370), .Z(n165) );
  NANDN U258 ( .A(n4368), .B(n4367), .Z(n166) );
  NAND U259 ( .A(n165), .B(n166), .Z(n4409) );
  NAND U260 ( .A(n4484), .B(n4485), .Z(n167) );
  NANDN U261 ( .A(n4483), .B(n4482), .Z(n168) );
  NAND U262 ( .A(n167), .B(n168), .Z(n4524) );
  NAND U263 ( .A(n4601), .B(n4602), .Z(n169) );
  NANDN U264 ( .A(n4600), .B(n4599), .Z(n170) );
  NAND U265 ( .A(n169), .B(n170), .Z(n4641) );
  NAND U266 ( .A(n4718), .B(n4719), .Z(n171) );
  NANDN U267 ( .A(n4717), .B(n4716), .Z(n172) );
  NAND U268 ( .A(n171), .B(n172), .Z(n4758) );
  NAND U269 ( .A(n4835), .B(n4836), .Z(n173) );
  NANDN U270 ( .A(n4834), .B(n4833), .Z(n174) );
  NAND U271 ( .A(n173), .B(n174), .Z(n4875) );
  NAND U272 ( .A(n4952), .B(n4953), .Z(n175) );
  NANDN U273 ( .A(n4951), .B(n4950), .Z(n176) );
  NAND U274 ( .A(n175), .B(n176), .Z(n4992) );
  NAND U275 ( .A(n5069), .B(n5070), .Z(n177) );
  NANDN U276 ( .A(n5068), .B(n5067), .Z(n178) );
  NAND U277 ( .A(n177), .B(n178), .Z(n5116) );
  XOR U278 ( .A(n341), .B(n340), .Z(n179) );
  NAND U279 ( .A(n179), .B(n339), .Z(n180) );
  NAND U280 ( .A(n341), .B(n340), .Z(n181) );
  AND U281 ( .A(n180), .B(n181), .Z(n345) );
  NAND U282 ( .A(n5227), .B(n5226), .Z(n182) );
  NANDN U283 ( .A(n5229), .B(n5228), .Z(n183) );
  AND U284 ( .A(n182), .B(n183), .Z(n5254) );
  NAND U285 ( .A(n5326), .B(n5325), .Z(n184) );
  XOR U286 ( .A(n5325), .B(n5326), .Z(n185) );
  NANDN U287 ( .A(n5324), .B(n185), .Z(n186) );
  NAND U288 ( .A(n184), .B(n186), .Z(n5338) );
  NAND U289 ( .A(n404), .B(n405), .Z(n187) );
  NANDN U290 ( .A(n403), .B(n402), .Z(n188) );
  NAND U291 ( .A(n187), .B(n188), .Z(n445) );
  XNOR U292 ( .A(n5173), .B(n5174), .Z(n5166) );
  NANDN U293 ( .A(a[0]), .B(n5160), .Z(n189) );
  NANDN U294 ( .A(b[2]), .B(n5199), .Z(n190) );
  NAND U295 ( .A(n190), .B(n189), .Z(n191) );
  NANDN U296 ( .A(n293), .B(n191), .Z(n339) );
  XOR U297 ( .A(n401), .B(n400), .Z(n192) );
  NANDN U298 ( .A(n399), .B(n192), .Z(n193) );
  NAND U299 ( .A(n401), .B(n400), .Z(n194) );
  AND U300 ( .A(n193), .B(n194), .Z(n438) );
  NAND U301 ( .A(n672), .B(n673), .Z(n195) );
  NANDN U302 ( .A(n671), .B(n670), .Z(n196) );
  NAND U303 ( .A(n195), .B(n196), .Z(n712) );
  NAND U304 ( .A(n789), .B(n790), .Z(n197) );
  NANDN U305 ( .A(n788), .B(n787), .Z(n198) );
  NAND U306 ( .A(n197), .B(n198), .Z(n829) );
  NAND U307 ( .A(n906), .B(n907), .Z(n199) );
  NANDN U308 ( .A(n905), .B(n904), .Z(n200) );
  NAND U309 ( .A(n199), .B(n200), .Z(n946) );
  NAND U310 ( .A(n1023), .B(n1024), .Z(n201) );
  NANDN U311 ( .A(n1022), .B(n1021), .Z(n202) );
  NAND U312 ( .A(n201), .B(n202), .Z(n1063) );
  NAND U313 ( .A(n1140), .B(n1141), .Z(n203) );
  NANDN U314 ( .A(n1139), .B(n1138), .Z(n204) );
  NAND U315 ( .A(n203), .B(n204), .Z(n1180) );
  NAND U316 ( .A(n1257), .B(n1258), .Z(n205) );
  NANDN U317 ( .A(n1256), .B(n1255), .Z(n206) );
  NAND U318 ( .A(n205), .B(n206), .Z(n1297) );
  NAND U319 ( .A(n1374), .B(n1375), .Z(n207) );
  NANDN U320 ( .A(n1373), .B(n1372), .Z(n208) );
  NAND U321 ( .A(n207), .B(n208), .Z(n1414) );
  NAND U322 ( .A(n1491), .B(n1492), .Z(n209) );
  NANDN U323 ( .A(n1490), .B(n1489), .Z(n210) );
  NAND U324 ( .A(n209), .B(n210), .Z(n1531) );
  NAND U325 ( .A(n1608), .B(n1609), .Z(n211) );
  NANDN U326 ( .A(n1607), .B(n1606), .Z(n212) );
  NAND U327 ( .A(n211), .B(n212), .Z(n1648) );
  NAND U328 ( .A(n1725), .B(n1726), .Z(n213) );
  NANDN U329 ( .A(n1724), .B(n1723), .Z(n214) );
  NAND U330 ( .A(n213), .B(n214), .Z(n1765) );
  NAND U331 ( .A(n1840), .B(n1841), .Z(n215) );
  NANDN U332 ( .A(n1839), .B(n1838), .Z(n216) );
  NAND U333 ( .A(n215), .B(n216), .Z(n1880) );
  NAND U334 ( .A(n1957), .B(n1958), .Z(n217) );
  NANDN U335 ( .A(n1956), .B(n1955), .Z(n218) );
  NAND U336 ( .A(n217), .B(n218), .Z(n1997) );
  NAND U337 ( .A(n2074), .B(n2075), .Z(n219) );
  NANDN U338 ( .A(n2073), .B(n2072), .Z(n220) );
  NAND U339 ( .A(n219), .B(n220), .Z(n2114) );
  NAND U340 ( .A(n2191), .B(n2192), .Z(n221) );
  NANDN U341 ( .A(n2190), .B(n2189), .Z(n222) );
  NAND U342 ( .A(n221), .B(n222), .Z(n2231) );
  NAND U343 ( .A(n2308), .B(n2309), .Z(n223) );
  NANDN U344 ( .A(n2307), .B(n2306), .Z(n224) );
  NAND U345 ( .A(n223), .B(n224), .Z(n2348) );
  NAND U346 ( .A(n2425), .B(n2426), .Z(n225) );
  NANDN U347 ( .A(n2424), .B(n2423), .Z(n226) );
  NAND U348 ( .A(n225), .B(n226), .Z(n2463) );
  NAND U349 ( .A(n2540), .B(n2541), .Z(n227) );
  NANDN U350 ( .A(n2539), .B(n2538), .Z(n228) );
  NAND U351 ( .A(n227), .B(n228), .Z(n2581) );
  NAND U352 ( .A(n2656), .B(n2657), .Z(n229) );
  NANDN U353 ( .A(n2655), .B(n2654), .Z(n230) );
  NAND U354 ( .A(n229), .B(n230), .Z(n2696) );
  NAND U355 ( .A(n2773), .B(n2774), .Z(n231) );
  NANDN U356 ( .A(n2772), .B(n2771), .Z(n232) );
  NAND U357 ( .A(n231), .B(n232), .Z(n2813) );
  NAND U358 ( .A(n2890), .B(n2891), .Z(n233) );
  NANDN U359 ( .A(n2889), .B(n2888), .Z(n234) );
  NAND U360 ( .A(n233), .B(n234), .Z(n2930) );
  NAND U361 ( .A(n3007), .B(n3008), .Z(n235) );
  NANDN U362 ( .A(n3006), .B(n3005), .Z(n236) );
  NAND U363 ( .A(n235), .B(n236), .Z(n3047) );
  NAND U364 ( .A(n3124), .B(n3125), .Z(n237) );
  NANDN U365 ( .A(n3123), .B(n3122), .Z(n238) );
  NAND U366 ( .A(n237), .B(n238), .Z(n3164) );
  NAND U367 ( .A(n3239), .B(n3240), .Z(n239) );
  NANDN U368 ( .A(n3238), .B(n3237), .Z(n240) );
  NAND U369 ( .A(n239), .B(n240), .Z(n3279) );
  NAND U370 ( .A(n3356), .B(n3357), .Z(n241) );
  NANDN U371 ( .A(n3355), .B(n3354), .Z(n242) );
  NAND U372 ( .A(n241), .B(n242), .Z(n3396) );
  NAND U373 ( .A(n3473), .B(n3474), .Z(n243) );
  NANDN U374 ( .A(n3472), .B(n3471), .Z(n244) );
  NAND U375 ( .A(n243), .B(n244), .Z(n3513) );
  NAND U376 ( .A(n3590), .B(n3591), .Z(n245) );
  NANDN U377 ( .A(n3589), .B(n3588), .Z(n246) );
  NAND U378 ( .A(n245), .B(n246), .Z(n3630) );
  NAND U379 ( .A(n3707), .B(n3708), .Z(n247) );
  NANDN U380 ( .A(n3706), .B(n3705), .Z(n248) );
  NAND U381 ( .A(n247), .B(n248), .Z(n3747) );
  NAND U382 ( .A(n3824), .B(n3825), .Z(n249) );
  NANDN U383 ( .A(n3823), .B(n3822), .Z(n250) );
  NAND U384 ( .A(n249), .B(n250), .Z(n3864) );
  NAND U385 ( .A(n3941), .B(n3942), .Z(n251) );
  NANDN U386 ( .A(n3940), .B(n3939), .Z(n252) );
  NAND U387 ( .A(n251), .B(n252), .Z(n3981) );
  NAND U388 ( .A(n4058), .B(n4059), .Z(n253) );
  NANDN U389 ( .A(n4057), .B(n4056), .Z(n254) );
  NAND U390 ( .A(n253), .B(n254), .Z(n4098) );
  NAND U391 ( .A(n4176), .B(n4177), .Z(n255) );
  NANDN U392 ( .A(n4175), .B(n4174), .Z(n256) );
  NAND U393 ( .A(n255), .B(n256), .Z(n4214) );
  NAND U394 ( .A(n4291), .B(n4292), .Z(n257) );
  NANDN U395 ( .A(n4290), .B(n4289), .Z(n258) );
  NAND U396 ( .A(n257), .B(n258), .Z(n4331) );
  NAND U397 ( .A(n4408), .B(n4409), .Z(n259) );
  NANDN U398 ( .A(n4407), .B(n4406), .Z(n260) );
  NAND U399 ( .A(n259), .B(n260), .Z(n4448) );
  NAND U400 ( .A(n4523), .B(n4524), .Z(n261) );
  NANDN U401 ( .A(n4522), .B(n4521), .Z(n262) );
  NAND U402 ( .A(n261), .B(n262), .Z(n4563) );
  NAND U403 ( .A(n4640), .B(n4641), .Z(n263) );
  NANDN U404 ( .A(n4639), .B(n4638), .Z(n264) );
  NAND U405 ( .A(n263), .B(n264), .Z(n4680) );
  NAND U406 ( .A(n4757), .B(n4758), .Z(n265) );
  NANDN U407 ( .A(n4756), .B(n4755), .Z(n266) );
  NAND U408 ( .A(n265), .B(n266), .Z(n4797) );
  NAND U409 ( .A(n4874), .B(n4875), .Z(n267) );
  NANDN U410 ( .A(n4873), .B(n4872), .Z(n268) );
  NAND U411 ( .A(n267), .B(n268), .Z(n4914) );
  NAND U412 ( .A(n4991), .B(n4992), .Z(n269) );
  NANDN U413 ( .A(n4990), .B(n4989), .Z(n270) );
  NAND U414 ( .A(n269), .B(n270), .Z(n5031) );
  ANDN U415 ( .B(n338), .A(n337), .Z(n344) );
  NAND U416 ( .A(n5115), .B(n5116), .Z(n271) );
  NANDN U417 ( .A(n5114), .B(n5113), .Z(n272) );
  NAND U418 ( .A(n271), .B(n272), .Z(n5151) );
  XOR U419 ( .A(n5255), .B(n5254), .Z(n273) );
  NANDN U420 ( .A(n5253), .B(n273), .Z(n274) );
  NAND U421 ( .A(n5255), .B(n5254), .Z(n275) );
  AND U422 ( .A(n274), .B(n275), .Z(n5302) );
  XNOR U423 ( .A(n294), .B(b[7]), .Z(n276) );
  ANDN U424 ( .B(n276), .A(n5336), .Z(n277) );
  NANDN U425 ( .A(n295), .B(b[5]), .Z(n278) );
  NANDN U426 ( .A(n277), .B(n278), .Z(n279) );
  AND U427 ( .A(a[127]), .B(n279), .Z(n280) );
  NANDN U428 ( .A(n5339), .B(n5338), .Z(n281) );
  XNOR U429 ( .A(n5339), .B(n5338), .Z(n282) );
  NAND U430 ( .A(n282), .B(n5337), .Z(n283) );
  NAND U431 ( .A(n281), .B(n283), .Z(n284) );
  XNOR U432 ( .A(n280), .B(n284), .Z(n285) );
  OR U433 ( .A(n5340), .B(n5341), .Z(n286) );
  XNOR U434 ( .A(n5341), .B(n5342), .Z(n287) );
  NANDN U435 ( .A(n5343), .B(n287), .Z(n288) );
  NAND U436 ( .A(n286), .B(n288), .Z(n289) );
  XNOR U437 ( .A(n285), .B(n289), .Z(n290) );
  NANDN U438 ( .A(n5345), .B(n5344), .Z(n291) );
  XNOR U439 ( .A(n290), .B(n291), .Z(c[255]) );
  IV U440 ( .A(b[0]), .Z(n292) );
  IV U441 ( .A(b[3]), .Z(n293) );
  IV U442 ( .A(b[5]), .Z(n294) );
  IV U443 ( .A(b[7]), .Z(n295) );
  NANDN U444 ( .A(n292), .B(a[0]), .Z(n297) );
  XNOR U445 ( .A(n297), .B(sreg[120]), .Z(c[120]) );
  IV U446 ( .A(b[1]), .Z(n5199) );
  ANDN U447 ( .B(a[0]), .A(n5199), .Z(n296) );
  NANDN U448 ( .A(n292), .B(a[1]), .Z(n302) );
  XNOR U449 ( .A(n296), .B(n302), .Z(n305) );
  XNOR U450 ( .A(sreg[121]), .B(n305), .Z(n307) );
  NANDN U451 ( .A(n297), .B(sreg[120]), .Z(n306) );
  XOR U452 ( .A(n307), .B(n306), .Z(c[121]) );
  NANDN U453 ( .A(n292), .B(a[2]), .Z(n298) );
  XOR U454 ( .A(n5199), .B(n298), .Z(n300) );
  NANDN U455 ( .A(b[0]), .B(a[1]), .Z(n299) );
  AND U456 ( .A(n300), .B(n299), .Z(n310) );
  IV U457 ( .A(a[0]), .Z(n465) );
  NANDN U458 ( .A(n465), .B(b[2]), .Z(n301) );
  XOR U459 ( .A(n5199), .B(n301), .Z(n304) );
  OR U460 ( .A(n302), .B(a[0]), .Z(n303) );
  AND U461 ( .A(n304), .B(n303), .Z(n311) );
  XOR U462 ( .A(n310), .B(n311), .Z(n322) );
  NAND U463 ( .A(sreg[121]), .B(n305), .Z(n309) );
  OR U464 ( .A(n307), .B(n306), .Z(n308) );
  NAND U465 ( .A(n309), .B(n308), .Z(n321) );
  XNOR U466 ( .A(n321), .B(sreg[122]), .Z(n323) );
  XNOR U467 ( .A(n322), .B(n323), .Z(c[122]) );
  NAND U468 ( .A(n311), .B(n310), .Z(n341) );
  XNOR U469 ( .A(n5199), .B(b[2]), .Z(n5160) );
  XNOR U470 ( .A(n293), .B(a[0]), .Z(n314) );
  XNOR U471 ( .A(n293), .B(b[1]), .Z(n313) );
  XNOR U472 ( .A(n293), .B(b[2]), .Z(n312) );
  AND U473 ( .A(n313), .B(n312), .Z(n5161) );
  NAND U474 ( .A(n314), .B(n5161), .Z(n316) );
  XNOR U475 ( .A(n293), .B(a[1]), .Z(n334) );
  NAND U476 ( .A(n334), .B(n5160), .Z(n315) );
  AND U477 ( .A(n316), .B(n315), .Z(n337) );
  NANDN U478 ( .A(n292), .B(a[3]), .Z(n317) );
  XOR U479 ( .A(n5199), .B(n317), .Z(n319) );
  NANDN U480 ( .A(b[0]), .B(a[2]), .Z(n318) );
  AND U481 ( .A(n319), .B(n318), .Z(n338) );
  XOR U482 ( .A(n337), .B(n338), .Z(n340) );
  XOR U483 ( .A(n339), .B(n340), .Z(n320) );
  XNOR U484 ( .A(n341), .B(n320), .Z(n326) );
  XNOR U485 ( .A(sreg[123]), .B(n326), .Z(n328) );
  NAND U486 ( .A(n321), .B(sreg[122]), .Z(n325) );
  NANDN U487 ( .A(n323), .B(n322), .Z(n324) );
  AND U488 ( .A(n325), .B(n324), .Z(n327) );
  XOR U489 ( .A(n328), .B(n327), .Z(c[123]) );
  NAND U490 ( .A(sreg[123]), .B(n326), .Z(n330) );
  OR U491 ( .A(n328), .B(n327), .Z(n329) );
  NAND U492 ( .A(n330), .B(n329), .Z(n365) );
  XNOR U493 ( .A(n365), .B(sreg[124]), .Z(n367) );
  NANDN U494 ( .A(n292), .B(a[4]), .Z(n331) );
  XOR U495 ( .A(n5199), .B(n331), .Z(n333) );
  NANDN U496 ( .A(b[0]), .B(a[3]), .Z(n332) );
  AND U497 ( .A(n333), .B(n332), .Z(n359) );
  XNOR U498 ( .A(b[3]), .B(a[2]), .Z(n346) );
  NANDN U499 ( .A(n346), .B(n5160), .Z(n336) );
  NAND U500 ( .A(n334), .B(n5161), .Z(n335) );
  AND U501 ( .A(n336), .B(n335), .Z(n360) );
  XOR U502 ( .A(n359), .B(n360), .Z(n362) );
  IV U503 ( .A(b[4]), .Z(n5269) );
  XOR U504 ( .A(n293), .B(n5269), .Z(n5240) );
  NANDN U505 ( .A(n465), .B(n5240), .Z(n361) );
  XNOR U506 ( .A(n362), .B(n361), .Z(n343) );
  XOR U507 ( .A(n344), .B(n345), .Z(n342) );
  XNOR U508 ( .A(n343), .B(n342), .Z(n366) );
  XNOR U509 ( .A(n367), .B(n366), .Z(c[124]) );
  XNOR U510 ( .A(b[3]), .B(a[3]), .Z(n378) );
  NANDN U511 ( .A(n378), .B(n5160), .Z(n348) );
  NANDN U512 ( .A(n346), .B(n5161), .Z(n347) );
  NAND U513 ( .A(n348), .B(n347), .Z(n387) );
  NANDN U514 ( .A(n293), .B(b[4]), .Z(n5268) );
  ANDN U515 ( .B(n5268), .A(n294), .Z(n5317) );
  XNOR U516 ( .A(n5269), .B(b[3]), .Z(n349) );
  NANDN U517 ( .A(n465), .B(n349), .Z(n350) );
  NAND U518 ( .A(n5317), .B(n350), .Z(n388) );
  XNOR U519 ( .A(n387), .B(n388), .Z(n389) );
  NANDN U520 ( .A(n292), .B(a[5]), .Z(n351) );
  XOR U521 ( .A(n5199), .B(n351), .Z(n353) );
  NANDN U522 ( .A(b[0]), .B(a[4]), .Z(n352) );
  NAND U523 ( .A(n353), .B(n352), .Z(n376) );
  XNOR U524 ( .A(n294), .B(a[0]), .Z(n356) );
  XNOR U525 ( .A(n294), .B(b[3]), .Z(n355) );
  XNOR U526 ( .A(n294), .B(b[4]), .Z(n354) );
  AND U527 ( .A(n355), .B(n354), .Z(n5241) );
  NAND U528 ( .A(n356), .B(n5241), .Z(n358) );
  XNOR U529 ( .A(n294), .B(a[1]), .Z(n384) );
  AND U530 ( .A(n5240), .B(n384), .Z(n357) );
  ANDN U531 ( .B(n358), .A(n357), .Z(n377) );
  XNOR U532 ( .A(n376), .B(n377), .Z(n390) );
  XOR U533 ( .A(n389), .B(n390), .Z(n370) );
  NANDN U534 ( .A(n360), .B(n359), .Z(n364) );
  OR U535 ( .A(n362), .B(n361), .Z(n363) );
  NAND U536 ( .A(n364), .B(n363), .Z(n371) );
  XNOR U537 ( .A(n370), .B(n371), .Z(n373) );
  XOR U538 ( .A(n372), .B(n373), .Z(n394) );
  XOR U539 ( .A(n394), .B(sreg[125]), .Z(n396) );
  NAND U540 ( .A(n365), .B(sreg[124]), .Z(n369) );
  NANDN U541 ( .A(n367), .B(n366), .Z(n368) );
  AND U542 ( .A(n369), .B(n368), .Z(n395) );
  XOR U543 ( .A(n396), .B(n395), .Z(c[125]) );
  NANDN U544 ( .A(n371), .B(n370), .Z(n375) );
  NAND U545 ( .A(n373), .B(n372), .Z(n374) );
  NAND U546 ( .A(n375), .B(n374), .Z(n401) );
  XNOR U547 ( .A(n293), .B(a[4]), .Z(n417) );
  NAND U548 ( .A(n417), .B(n5160), .Z(n380) );
  NANDN U549 ( .A(n378), .B(n5161), .Z(n379) );
  NAND U550 ( .A(n380), .B(n379), .Z(n405) );
  IV U551 ( .A(b[6]), .Z(n5336) );
  XOR U552 ( .A(n294), .B(n5336), .Z(n5293) );
  NANDN U553 ( .A(n465), .B(n5293), .Z(n403) );
  NANDN U554 ( .A(n292), .B(a[6]), .Z(n381) );
  XOR U555 ( .A(n5199), .B(n381), .Z(n383) );
  NANDN U556 ( .A(b[0]), .B(a[5]), .Z(n382) );
  AND U557 ( .A(n383), .B(n382), .Z(n402) );
  XNOR U558 ( .A(n403), .B(n402), .Z(n404) );
  XNOR U559 ( .A(n405), .B(n404), .Z(n420) );
  XNOR U560 ( .A(b[5]), .B(a[2]), .Z(n406) );
  NANDN U561 ( .A(n406), .B(n5240), .Z(n386) );
  NAND U562 ( .A(n5241), .B(n384), .Z(n385) );
  NAND U563 ( .A(n386), .B(n385), .Z(n421) );
  XNOR U564 ( .A(n420), .B(n421), .Z(n422) );
  XOR U565 ( .A(n423), .B(n422), .Z(n399) );
  NANDN U566 ( .A(n388), .B(n387), .Z(n392) );
  NANDN U567 ( .A(n390), .B(n389), .Z(n391) );
  AND U568 ( .A(n392), .B(n391), .Z(n400) );
  XOR U569 ( .A(n399), .B(n400), .Z(n393) );
  XNOR U570 ( .A(n401), .B(n393), .Z(n428) );
  NANDN U571 ( .A(n394), .B(sreg[125]), .Z(n398) );
  OR U572 ( .A(n396), .B(n395), .Z(n397) );
  NAND U573 ( .A(n398), .B(n397), .Z(n426) );
  XNOR U574 ( .A(n426), .B(sreg[126]), .Z(n427) );
  XOR U575 ( .A(n428), .B(n427), .Z(c[126]) );
  XNOR U576 ( .A(n294), .B(a[3]), .Z(n466) );
  NAND U577 ( .A(n466), .B(n5240), .Z(n408) );
  NANDN U578 ( .A(n406), .B(n5241), .Z(n407) );
  NAND U579 ( .A(n408), .B(n407), .Z(n455) );
  XNOR U580 ( .A(n295), .B(a[1]), .Z(n459) );
  AND U581 ( .A(n5293), .B(n459), .Z(n413) );
  XNOR U582 ( .A(n295), .B(a[0]), .Z(n411) );
  XNOR U583 ( .A(n295), .B(b[5]), .Z(n410) );
  XNOR U584 ( .A(n295), .B(b[6]), .Z(n409) );
  AND U585 ( .A(n410), .B(n409), .Z(n5294) );
  NAND U586 ( .A(n411), .B(n5294), .Z(n412) );
  NANDN U587 ( .A(n413), .B(n412), .Z(n454) );
  XNOR U588 ( .A(n455), .B(n454), .Z(n451) );
  NANDN U589 ( .A(n292), .B(a[7]), .Z(n414) );
  XOR U590 ( .A(n5199), .B(n414), .Z(n416) );
  NANDN U591 ( .A(b[0]), .B(a[6]), .Z(n415) );
  AND U592 ( .A(n416), .B(n415), .Z(n449) );
  XOR U593 ( .A(n448), .B(n449), .Z(n450) );
  XOR U594 ( .A(n451), .B(n450), .Z(n442) );
  XOR U595 ( .A(n293), .B(a[5]), .Z(n456) );
  NANDN U596 ( .A(n456), .B(n5160), .Z(n419) );
  NAND U597 ( .A(n5161), .B(n417), .Z(n418) );
  AND U598 ( .A(n419), .B(n418), .Z(n443) );
  XNOR U599 ( .A(n442), .B(n443), .Z(n444) );
  XNOR U600 ( .A(n445), .B(n444), .Z(n436) );
  NANDN U601 ( .A(n421), .B(n420), .Z(n425) );
  NANDN U602 ( .A(n423), .B(n422), .Z(n424) );
  NAND U603 ( .A(n425), .B(n424), .Z(n437) );
  XNOR U604 ( .A(n436), .B(n437), .Z(n439) );
  XOR U605 ( .A(n438), .B(n439), .Z(n431) );
  XNOR U606 ( .A(sreg[127]), .B(n431), .Z(n433) );
  NAND U607 ( .A(n426), .B(sreg[126]), .Z(n430) );
  OR U608 ( .A(n428), .B(n427), .Z(n429) );
  AND U609 ( .A(n430), .B(n429), .Z(n432) );
  XOR U610 ( .A(n433), .B(n432), .Z(c[127]) );
  NAND U611 ( .A(sreg[127]), .B(n431), .Z(n435) );
  OR U612 ( .A(n433), .B(n432), .Z(n434) );
  NAND U613 ( .A(n435), .B(n434), .Z(n505) );
  XNOR U614 ( .A(n505), .B(sreg[128]), .Z(n507) );
  NANDN U615 ( .A(n437), .B(n436), .Z(n441) );
  NAND U616 ( .A(n439), .B(n438), .Z(n440) );
  NAND U617 ( .A(n441), .B(n440), .Z(n502) );
  NAND U618 ( .A(n443), .B(n442), .Z(n447) );
  OR U619 ( .A(n445), .B(n444), .Z(n446) );
  NAND U620 ( .A(n447), .B(n446), .Z(n500) );
  OR U621 ( .A(n449), .B(n448), .Z(n453) );
  NAND U622 ( .A(n451), .B(n450), .Z(n452) );
  NAND U623 ( .A(n453), .B(n452), .Z(n493) );
  NAND U624 ( .A(n455), .B(n454), .Z(n490) );
  XNOR U625 ( .A(b[3]), .B(a[6]), .Z(n472) );
  NANDN U626 ( .A(n472), .B(n5160), .Z(n458) );
  NANDN U627 ( .A(n456), .B(n5161), .Z(n457) );
  NAND U628 ( .A(n458), .B(n457), .Z(n488) );
  XNOR U629 ( .A(b[7]), .B(a[2]), .Z(n469) );
  NANDN U630 ( .A(n469), .B(n5293), .Z(n461) );
  NAND U631 ( .A(n5294), .B(n459), .Z(n460) );
  AND U632 ( .A(n461), .B(n460), .Z(n487) );
  XNOR U633 ( .A(n488), .B(n487), .Z(n489) );
  XNOR U634 ( .A(n490), .B(n489), .Z(n494) );
  XNOR U635 ( .A(n493), .B(n494), .Z(n495) );
  NANDN U636 ( .A(n292), .B(a[8]), .Z(n462) );
  XOR U637 ( .A(n5199), .B(n462), .Z(n464) );
  NANDN U638 ( .A(b[0]), .B(a[7]), .Z(n463) );
  AND U639 ( .A(n464), .B(n463), .Z(n484) );
  ANDN U640 ( .B(b[7]), .A(n465), .Z(n481) );
  XNOR U641 ( .A(b[5]), .B(a[4]), .Z(n478) );
  NANDN U642 ( .A(n478), .B(n5240), .Z(n468) );
  NAND U643 ( .A(n5241), .B(n466), .Z(n467) );
  NAND U644 ( .A(n468), .B(n467), .Z(n482) );
  XOR U645 ( .A(n481), .B(n482), .Z(n483) );
  XOR U646 ( .A(n484), .B(n483), .Z(n496) );
  XNOR U647 ( .A(n495), .B(n496), .Z(n499) );
  XNOR U648 ( .A(n500), .B(n499), .Z(n501) );
  XOR U649 ( .A(n502), .B(n501), .Z(n506) );
  XOR U650 ( .A(n507), .B(n506), .Z(c[128]) );
  XNOR U651 ( .A(b[7]), .B(a[3]), .Z(n528) );
  NANDN U652 ( .A(n528), .B(n5293), .Z(n471) );
  NANDN U653 ( .A(n469), .B(n5294), .Z(n470) );
  NAND U654 ( .A(n471), .B(n470), .Z(n516) );
  XNOR U655 ( .A(b[3]), .B(a[7]), .Z(n531) );
  NANDN U656 ( .A(n531), .B(n5160), .Z(n474) );
  NANDN U657 ( .A(n472), .B(n5161), .Z(n473) );
  AND U658 ( .A(n474), .B(n473), .Z(n517) );
  XNOR U659 ( .A(n516), .B(n517), .Z(n518) );
  NANDN U660 ( .A(n292), .B(a[9]), .Z(n475) );
  XOR U661 ( .A(n5199), .B(n475), .Z(n477) );
  NANDN U662 ( .A(b[0]), .B(a[8]), .Z(n476) );
  AND U663 ( .A(n477), .B(n476), .Z(n524) );
  XNOR U664 ( .A(b[5]), .B(a[5]), .Z(n537) );
  NANDN U665 ( .A(n537), .B(n5240), .Z(n480) );
  NANDN U666 ( .A(n478), .B(n5241), .Z(n479) );
  NAND U667 ( .A(n480), .B(n479), .Z(n522) );
  NANDN U668 ( .A(n295), .B(a[1]), .Z(n523) );
  XNOR U669 ( .A(n522), .B(n523), .Z(n525) );
  XOR U670 ( .A(n524), .B(n525), .Z(n519) );
  XOR U671 ( .A(n518), .B(n519), .Z(n540) );
  OR U672 ( .A(n482), .B(n481), .Z(n486) );
  NANDN U673 ( .A(n484), .B(n483), .Z(n485) );
  AND U674 ( .A(n486), .B(n485), .Z(n541) );
  XNOR U675 ( .A(n540), .B(n541), .Z(n543) );
  NANDN U676 ( .A(n488), .B(n487), .Z(n492) );
  NAND U677 ( .A(n490), .B(n489), .Z(n491) );
  AND U678 ( .A(n492), .B(n491), .Z(n542) );
  XNOR U679 ( .A(n543), .B(n542), .Z(n510) );
  NANDN U680 ( .A(n494), .B(n493), .Z(n498) );
  NANDN U681 ( .A(n496), .B(n495), .Z(n497) );
  AND U682 ( .A(n498), .B(n497), .Z(n511) );
  XNOR U683 ( .A(n510), .B(n511), .Z(n513) );
  NAND U684 ( .A(n500), .B(n499), .Z(n504) );
  OR U685 ( .A(n502), .B(n501), .Z(n503) );
  AND U686 ( .A(n504), .B(n503), .Z(n512) );
  XNOR U687 ( .A(n513), .B(n512), .Z(n546) );
  XNOR U688 ( .A(sreg[129]), .B(n546), .Z(n548) );
  NAND U689 ( .A(n505), .B(sreg[128]), .Z(n509) );
  OR U690 ( .A(n507), .B(n506), .Z(n508) );
  AND U691 ( .A(n509), .B(n508), .Z(n547) );
  XOR U692 ( .A(n548), .B(n547), .Z(c[129]) );
  NAND U693 ( .A(n511), .B(n510), .Z(n515) );
  NANDN U694 ( .A(n513), .B(n512), .Z(n514) );
  NAND U695 ( .A(n515), .B(n514), .Z(n553) );
  NANDN U696 ( .A(n517), .B(n516), .Z(n521) );
  NAND U697 ( .A(n519), .B(n518), .Z(n520) );
  NAND U698 ( .A(n521), .B(n520), .Z(n584) );
  NANDN U699 ( .A(n523), .B(n522), .Z(n527) );
  NAND U700 ( .A(n525), .B(n524), .Z(n526) );
  NAND U701 ( .A(n527), .B(n526), .Z(n582) );
  XNOR U702 ( .A(b[7]), .B(a[4]), .Z(n569) );
  NANDN U703 ( .A(n569), .B(n5293), .Z(n530) );
  NANDN U704 ( .A(n528), .B(n5294), .Z(n529) );
  NAND U705 ( .A(n530), .B(n529), .Z(n557) );
  XNOR U706 ( .A(b[3]), .B(a[8]), .Z(n572) );
  NANDN U707 ( .A(n572), .B(n5160), .Z(n533) );
  NANDN U708 ( .A(n531), .B(n5161), .Z(n532) );
  AND U709 ( .A(n533), .B(n532), .Z(n558) );
  XNOR U710 ( .A(n557), .B(n558), .Z(n559) );
  NANDN U711 ( .A(n292), .B(a[10]), .Z(n534) );
  XOR U712 ( .A(n5199), .B(n534), .Z(n536) );
  NANDN U713 ( .A(b[0]), .B(a[9]), .Z(n535) );
  AND U714 ( .A(n536), .B(n535), .Z(n565) );
  XNOR U715 ( .A(b[5]), .B(a[6]), .Z(n578) );
  NANDN U716 ( .A(n578), .B(n5240), .Z(n539) );
  NANDN U717 ( .A(n537), .B(n5241), .Z(n538) );
  NAND U718 ( .A(n539), .B(n538), .Z(n563) );
  NANDN U719 ( .A(n295), .B(a[2]), .Z(n564) );
  XNOR U720 ( .A(n563), .B(n564), .Z(n566) );
  XOR U721 ( .A(n565), .B(n566), .Z(n560) );
  XOR U722 ( .A(n559), .B(n560), .Z(n581) );
  XOR U723 ( .A(n582), .B(n581), .Z(n583) );
  XNOR U724 ( .A(n584), .B(n583), .Z(n551) );
  NAND U725 ( .A(n541), .B(n540), .Z(n545) );
  NANDN U726 ( .A(n543), .B(n542), .Z(n544) );
  NAND U727 ( .A(n545), .B(n544), .Z(n552) );
  XOR U728 ( .A(n551), .B(n552), .Z(n554) );
  XNOR U729 ( .A(n553), .B(n554), .Z(n587) );
  XNOR U730 ( .A(n587), .B(sreg[130]), .Z(n589) );
  NAND U731 ( .A(sreg[129]), .B(n546), .Z(n550) );
  OR U732 ( .A(n548), .B(n547), .Z(n549) );
  AND U733 ( .A(n550), .B(n549), .Z(n588) );
  XOR U734 ( .A(n589), .B(n588), .Z(c[130]) );
  NANDN U735 ( .A(n552), .B(n551), .Z(n556) );
  OR U736 ( .A(n554), .B(n553), .Z(n555) );
  NAND U737 ( .A(n556), .B(n555), .Z(n595) );
  NANDN U738 ( .A(n558), .B(n557), .Z(n562) );
  NAND U739 ( .A(n560), .B(n559), .Z(n561) );
  NAND U740 ( .A(n562), .B(n561), .Z(n623) );
  NANDN U741 ( .A(n564), .B(n563), .Z(n568) );
  NAND U742 ( .A(n566), .B(n565), .Z(n567) );
  NAND U743 ( .A(n568), .B(n567), .Z(n621) );
  XNOR U744 ( .A(b[7]), .B(a[5]), .Z(n608) );
  NANDN U745 ( .A(n608), .B(n5293), .Z(n571) );
  NANDN U746 ( .A(n569), .B(n5294), .Z(n570) );
  NAND U747 ( .A(n571), .B(n570), .Z(n596) );
  XNOR U748 ( .A(b[3]), .B(a[9]), .Z(n611) );
  NANDN U749 ( .A(n611), .B(n5160), .Z(n574) );
  NANDN U750 ( .A(n572), .B(n5161), .Z(n573) );
  AND U751 ( .A(n574), .B(n573), .Z(n597) );
  XNOR U752 ( .A(n596), .B(n597), .Z(n598) );
  NANDN U753 ( .A(n292), .B(a[11]), .Z(n575) );
  XOR U754 ( .A(n5199), .B(n575), .Z(n577) );
  NANDN U755 ( .A(b[0]), .B(a[10]), .Z(n576) );
  AND U756 ( .A(n577), .B(n576), .Z(n604) );
  XNOR U757 ( .A(b[5]), .B(a[7]), .Z(n617) );
  NANDN U758 ( .A(n617), .B(n5240), .Z(n580) );
  NANDN U759 ( .A(n578), .B(n5241), .Z(n579) );
  NAND U760 ( .A(n580), .B(n579), .Z(n602) );
  NANDN U761 ( .A(n295), .B(a[3]), .Z(n603) );
  XNOR U762 ( .A(n602), .B(n603), .Z(n605) );
  XOR U763 ( .A(n604), .B(n605), .Z(n599) );
  XOR U764 ( .A(n598), .B(n599), .Z(n620) );
  XOR U765 ( .A(n621), .B(n620), .Z(n622) );
  XNOR U766 ( .A(n623), .B(n622), .Z(n592) );
  NAND U767 ( .A(n582), .B(n581), .Z(n586) );
  NAND U768 ( .A(n584), .B(n583), .Z(n585) );
  NAND U769 ( .A(n586), .B(n585), .Z(n593) );
  XNOR U770 ( .A(n592), .B(n593), .Z(n594) );
  XNOR U771 ( .A(n595), .B(n594), .Z(n626) );
  XNOR U772 ( .A(n626), .B(sreg[131]), .Z(n628) );
  NAND U773 ( .A(n587), .B(sreg[130]), .Z(n591) );
  OR U774 ( .A(n589), .B(n588), .Z(n590) );
  AND U775 ( .A(n591), .B(n590), .Z(n627) );
  XOR U776 ( .A(n628), .B(n627), .Z(c[131]) );
  NANDN U777 ( .A(n597), .B(n596), .Z(n601) );
  NAND U778 ( .A(n599), .B(n598), .Z(n600) );
  NAND U779 ( .A(n601), .B(n600), .Z(n662) );
  NANDN U780 ( .A(n603), .B(n602), .Z(n607) );
  NAND U781 ( .A(n605), .B(n604), .Z(n606) );
  NAND U782 ( .A(n607), .B(n606), .Z(n660) );
  XNOR U783 ( .A(b[7]), .B(a[6]), .Z(n647) );
  NANDN U784 ( .A(n647), .B(n5293), .Z(n610) );
  NANDN U785 ( .A(n608), .B(n5294), .Z(n609) );
  NAND U786 ( .A(n610), .B(n609), .Z(n635) );
  XNOR U787 ( .A(b[3]), .B(a[10]), .Z(n650) );
  NANDN U788 ( .A(n650), .B(n5160), .Z(n613) );
  NANDN U789 ( .A(n611), .B(n5161), .Z(n612) );
  AND U790 ( .A(n613), .B(n612), .Z(n636) );
  XNOR U791 ( .A(n635), .B(n636), .Z(n637) );
  NANDN U792 ( .A(n292), .B(a[12]), .Z(n614) );
  XOR U793 ( .A(n5199), .B(n614), .Z(n616) );
  NANDN U794 ( .A(b[0]), .B(a[11]), .Z(n615) );
  AND U795 ( .A(n616), .B(n615), .Z(n643) );
  XNOR U796 ( .A(b[5]), .B(a[8]), .Z(n656) );
  NANDN U797 ( .A(n656), .B(n5240), .Z(n619) );
  NANDN U798 ( .A(n617), .B(n5241), .Z(n618) );
  NAND U799 ( .A(n619), .B(n618), .Z(n641) );
  NANDN U800 ( .A(n295), .B(a[4]), .Z(n642) );
  XNOR U801 ( .A(n641), .B(n642), .Z(n644) );
  XOR U802 ( .A(n643), .B(n644), .Z(n638) );
  XOR U803 ( .A(n637), .B(n638), .Z(n659) );
  XOR U804 ( .A(n660), .B(n659), .Z(n661) );
  XNOR U805 ( .A(n662), .B(n661), .Z(n631) );
  NAND U806 ( .A(n621), .B(n620), .Z(n625) );
  NAND U807 ( .A(n623), .B(n622), .Z(n624) );
  NAND U808 ( .A(n625), .B(n624), .Z(n632) );
  XNOR U809 ( .A(n631), .B(n632), .Z(n633) );
  XNOR U810 ( .A(n634), .B(n633), .Z(n665) );
  XNOR U811 ( .A(n665), .B(sreg[132]), .Z(n667) );
  NAND U812 ( .A(n626), .B(sreg[131]), .Z(n630) );
  OR U813 ( .A(n628), .B(n627), .Z(n629) );
  AND U814 ( .A(n630), .B(n629), .Z(n666) );
  XOR U815 ( .A(n667), .B(n666), .Z(c[132]) );
  NANDN U816 ( .A(n636), .B(n635), .Z(n640) );
  NAND U817 ( .A(n638), .B(n637), .Z(n639) );
  NAND U818 ( .A(n640), .B(n639), .Z(n701) );
  NANDN U819 ( .A(n642), .B(n641), .Z(n646) );
  NAND U820 ( .A(n644), .B(n643), .Z(n645) );
  NAND U821 ( .A(n646), .B(n645), .Z(n699) );
  XNOR U822 ( .A(b[7]), .B(a[7]), .Z(n686) );
  NANDN U823 ( .A(n686), .B(n5293), .Z(n649) );
  NANDN U824 ( .A(n647), .B(n5294), .Z(n648) );
  NAND U825 ( .A(n649), .B(n648), .Z(n674) );
  XNOR U826 ( .A(b[3]), .B(a[11]), .Z(n689) );
  NANDN U827 ( .A(n689), .B(n5160), .Z(n652) );
  NANDN U828 ( .A(n650), .B(n5161), .Z(n651) );
  AND U829 ( .A(n652), .B(n651), .Z(n675) );
  XNOR U830 ( .A(n674), .B(n675), .Z(n676) );
  NANDN U831 ( .A(n292), .B(a[13]), .Z(n653) );
  XOR U832 ( .A(n5199), .B(n653), .Z(n655) );
  NANDN U833 ( .A(b[0]), .B(a[12]), .Z(n654) );
  AND U834 ( .A(n655), .B(n654), .Z(n682) );
  XNOR U835 ( .A(b[5]), .B(a[9]), .Z(n695) );
  NANDN U836 ( .A(n695), .B(n5240), .Z(n658) );
  NANDN U837 ( .A(n656), .B(n5241), .Z(n657) );
  NAND U838 ( .A(n658), .B(n657), .Z(n680) );
  NANDN U839 ( .A(n295), .B(a[5]), .Z(n681) );
  XNOR U840 ( .A(n680), .B(n681), .Z(n683) );
  XOR U841 ( .A(n682), .B(n683), .Z(n677) );
  XOR U842 ( .A(n676), .B(n677), .Z(n698) );
  XOR U843 ( .A(n699), .B(n698), .Z(n700) );
  XNOR U844 ( .A(n701), .B(n700), .Z(n670) );
  NAND U845 ( .A(n660), .B(n659), .Z(n664) );
  NAND U846 ( .A(n662), .B(n661), .Z(n663) );
  NAND U847 ( .A(n664), .B(n663), .Z(n671) );
  XNOR U848 ( .A(n670), .B(n671), .Z(n672) );
  XNOR U849 ( .A(n673), .B(n672), .Z(n704) );
  XNOR U850 ( .A(n704), .B(sreg[133]), .Z(n706) );
  NAND U851 ( .A(n665), .B(sreg[132]), .Z(n669) );
  OR U852 ( .A(n667), .B(n666), .Z(n668) );
  AND U853 ( .A(n669), .B(n668), .Z(n705) );
  XOR U854 ( .A(n706), .B(n705), .Z(c[133]) );
  NANDN U855 ( .A(n675), .B(n674), .Z(n679) );
  NAND U856 ( .A(n677), .B(n676), .Z(n678) );
  NAND U857 ( .A(n679), .B(n678), .Z(n740) );
  NANDN U858 ( .A(n681), .B(n680), .Z(n685) );
  NAND U859 ( .A(n683), .B(n682), .Z(n684) );
  NAND U860 ( .A(n685), .B(n684), .Z(n738) );
  XNOR U861 ( .A(b[7]), .B(a[8]), .Z(n725) );
  NANDN U862 ( .A(n725), .B(n5293), .Z(n688) );
  NANDN U863 ( .A(n686), .B(n5294), .Z(n687) );
  NAND U864 ( .A(n688), .B(n687), .Z(n713) );
  XNOR U865 ( .A(b[3]), .B(a[12]), .Z(n728) );
  NANDN U866 ( .A(n728), .B(n5160), .Z(n691) );
  NANDN U867 ( .A(n689), .B(n5161), .Z(n690) );
  AND U868 ( .A(n691), .B(n690), .Z(n714) );
  XNOR U869 ( .A(n713), .B(n714), .Z(n715) );
  NANDN U870 ( .A(n292), .B(a[14]), .Z(n692) );
  XOR U871 ( .A(n5199), .B(n692), .Z(n694) );
  NANDN U872 ( .A(b[0]), .B(a[13]), .Z(n693) );
  AND U873 ( .A(n694), .B(n693), .Z(n721) );
  XNOR U874 ( .A(b[5]), .B(a[10]), .Z(n734) );
  NANDN U875 ( .A(n734), .B(n5240), .Z(n697) );
  NANDN U876 ( .A(n695), .B(n5241), .Z(n696) );
  NAND U877 ( .A(n697), .B(n696), .Z(n719) );
  NANDN U878 ( .A(n295), .B(a[6]), .Z(n720) );
  XNOR U879 ( .A(n719), .B(n720), .Z(n722) );
  XOR U880 ( .A(n721), .B(n722), .Z(n716) );
  XOR U881 ( .A(n715), .B(n716), .Z(n737) );
  XOR U882 ( .A(n738), .B(n737), .Z(n739) );
  XNOR U883 ( .A(n740), .B(n739), .Z(n709) );
  NAND U884 ( .A(n699), .B(n698), .Z(n703) );
  NAND U885 ( .A(n701), .B(n700), .Z(n702) );
  NAND U886 ( .A(n703), .B(n702), .Z(n710) );
  XNOR U887 ( .A(n709), .B(n710), .Z(n711) );
  XNOR U888 ( .A(n712), .B(n711), .Z(n743) );
  XNOR U889 ( .A(n743), .B(sreg[134]), .Z(n745) );
  NAND U890 ( .A(n704), .B(sreg[133]), .Z(n708) );
  OR U891 ( .A(n706), .B(n705), .Z(n707) );
  AND U892 ( .A(n708), .B(n707), .Z(n744) );
  XOR U893 ( .A(n745), .B(n744), .Z(c[134]) );
  NANDN U894 ( .A(n714), .B(n713), .Z(n718) );
  NAND U895 ( .A(n716), .B(n715), .Z(n717) );
  NAND U896 ( .A(n718), .B(n717), .Z(n779) );
  NANDN U897 ( .A(n720), .B(n719), .Z(n724) );
  NAND U898 ( .A(n722), .B(n721), .Z(n723) );
  NAND U899 ( .A(n724), .B(n723), .Z(n777) );
  XNOR U900 ( .A(b[7]), .B(a[9]), .Z(n764) );
  NANDN U901 ( .A(n764), .B(n5293), .Z(n727) );
  NANDN U902 ( .A(n725), .B(n5294), .Z(n726) );
  NAND U903 ( .A(n727), .B(n726), .Z(n752) );
  XNOR U904 ( .A(b[3]), .B(a[13]), .Z(n767) );
  NANDN U905 ( .A(n767), .B(n5160), .Z(n730) );
  NANDN U906 ( .A(n728), .B(n5161), .Z(n729) );
  AND U907 ( .A(n730), .B(n729), .Z(n753) );
  XNOR U908 ( .A(n752), .B(n753), .Z(n754) );
  NANDN U909 ( .A(n292), .B(a[15]), .Z(n731) );
  XOR U910 ( .A(n5199), .B(n731), .Z(n733) );
  NANDN U911 ( .A(b[0]), .B(a[14]), .Z(n732) );
  AND U912 ( .A(n733), .B(n732), .Z(n760) );
  XNOR U913 ( .A(b[5]), .B(a[11]), .Z(n773) );
  NANDN U914 ( .A(n773), .B(n5240), .Z(n736) );
  NANDN U915 ( .A(n734), .B(n5241), .Z(n735) );
  NAND U916 ( .A(n736), .B(n735), .Z(n758) );
  NANDN U917 ( .A(n295), .B(a[7]), .Z(n759) );
  XNOR U918 ( .A(n758), .B(n759), .Z(n761) );
  XOR U919 ( .A(n760), .B(n761), .Z(n755) );
  XOR U920 ( .A(n754), .B(n755), .Z(n776) );
  XOR U921 ( .A(n777), .B(n776), .Z(n778) );
  XNOR U922 ( .A(n779), .B(n778), .Z(n748) );
  NAND U923 ( .A(n738), .B(n737), .Z(n742) );
  NAND U924 ( .A(n740), .B(n739), .Z(n741) );
  NAND U925 ( .A(n742), .B(n741), .Z(n749) );
  XNOR U926 ( .A(n748), .B(n749), .Z(n750) );
  XNOR U927 ( .A(n751), .B(n750), .Z(n782) );
  XNOR U928 ( .A(n782), .B(sreg[135]), .Z(n784) );
  NAND U929 ( .A(n743), .B(sreg[134]), .Z(n747) );
  OR U930 ( .A(n745), .B(n744), .Z(n746) );
  AND U931 ( .A(n747), .B(n746), .Z(n783) );
  XOR U932 ( .A(n784), .B(n783), .Z(c[135]) );
  NANDN U933 ( .A(n753), .B(n752), .Z(n757) );
  NAND U934 ( .A(n755), .B(n754), .Z(n756) );
  NAND U935 ( .A(n757), .B(n756), .Z(n818) );
  NANDN U936 ( .A(n759), .B(n758), .Z(n763) );
  NAND U937 ( .A(n761), .B(n760), .Z(n762) );
  NAND U938 ( .A(n763), .B(n762), .Z(n816) );
  XNOR U939 ( .A(b[7]), .B(a[10]), .Z(n803) );
  NANDN U940 ( .A(n803), .B(n5293), .Z(n766) );
  NANDN U941 ( .A(n764), .B(n5294), .Z(n765) );
  NAND U942 ( .A(n766), .B(n765), .Z(n791) );
  XNOR U943 ( .A(b[3]), .B(a[14]), .Z(n806) );
  NANDN U944 ( .A(n806), .B(n5160), .Z(n769) );
  NANDN U945 ( .A(n767), .B(n5161), .Z(n768) );
  AND U946 ( .A(n769), .B(n768), .Z(n792) );
  XNOR U947 ( .A(n791), .B(n792), .Z(n793) );
  NANDN U948 ( .A(n292), .B(a[16]), .Z(n770) );
  XOR U949 ( .A(n5199), .B(n770), .Z(n772) );
  NANDN U950 ( .A(b[0]), .B(a[15]), .Z(n771) );
  AND U951 ( .A(n772), .B(n771), .Z(n799) );
  XNOR U952 ( .A(b[5]), .B(a[12]), .Z(n812) );
  NANDN U953 ( .A(n812), .B(n5240), .Z(n775) );
  NANDN U954 ( .A(n773), .B(n5241), .Z(n774) );
  NAND U955 ( .A(n775), .B(n774), .Z(n797) );
  NANDN U956 ( .A(n295), .B(a[8]), .Z(n798) );
  XNOR U957 ( .A(n797), .B(n798), .Z(n800) );
  XOR U958 ( .A(n799), .B(n800), .Z(n794) );
  XOR U959 ( .A(n793), .B(n794), .Z(n815) );
  XOR U960 ( .A(n816), .B(n815), .Z(n817) );
  XNOR U961 ( .A(n818), .B(n817), .Z(n787) );
  NAND U962 ( .A(n777), .B(n776), .Z(n781) );
  NAND U963 ( .A(n779), .B(n778), .Z(n780) );
  NAND U964 ( .A(n781), .B(n780), .Z(n788) );
  XNOR U965 ( .A(n787), .B(n788), .Z(n789) );
  XNOR U966 ( .A(n790), .B(n789), .Z(n821) );
  XNOR U967 ( .A(n821), .B(sreg[136]), .Z(n823) );
  NAND U968 ( .A(n782), .B(sreg[135]), .Z(n786) );
  OR U969 ( .A(n784), .B(n783), .Z(n785) );
  AND U970 ( .A(n786), .B(n785), .Z(n822) );
  XOR U971 ( .A(n823), .B(n822), .Z(c[136]) );
  NANDN U972 ( .A(n792), .B(n791), .Z(n796) );
  NAND U973 ( .A(n794), .B(n793), .Z(n795) );
  NAND U974 ( .A(n796), .B(n795), .Z(n857) );
  NANDN U975 ( .A(n798), .B(n797), .Z(n802) );
  NAND U976 ( .A(n800), .B(n799), .Z(n801) );
  NAND U977 ( .A(n802), .B(n801), .Z(n855) );
  XNOR U978 ( .A(b[7]), .B(a[11]), .Z(n842) );
  NANDN U979 ( .A(n842), .B(n5293), .Z(n805) );
  NANDN U980 ( .A(n803), .B(n5294), .Z(n804) );
  NAND U981 ( .A(n805), .B(n804), .Z(n830) );
  XNOR U982 ( .A(b[3]), .B(a[15]), .Z(n845) );
  NANDN U983 ( .A(n845), .B(n5160), .Z(n808) );
  NANDN U984 ( .A(n806), .B(n5161), .Z(n807) );
  AND U985 ( .A(n808), .B(n807), .Z(n831) );
  XNOR U986 ( .A(n830), .B(n831), .Z(n832) );
  NANDN U987 ( .A(n292), .B(a[17]), .Z(n809) );
  XOR U988 ( .A(n5199), .B(n809), .Z(n811) );
  NANDN U989 ( .A(b[0]), .B(a[16]), .Z(n810) );
  AND U990 ( .A(n811), .B(n810), .Z(n838) );
  XNOR U991 ( .A(b[5]), .B(a[13]), .Z(n851) );
  NANDN U992 ( .A(n851), .B(n5240), .Z(n814) );
  NANDN U993 ( .A(n812), .B(n5241), .Z(n813) );
  NAND U994 ( .A(n814), .B(n813), .Z(n836) );
  NANDN U995 ( .A(n295), .B(a[9]), .Z(n837) );
  XNOR U996 ( .A(n836), .B(n837), .Z(n839) );
  XOR U997 ( .A(n838), .B(n839), .Z(n833) );
  XOR U998 ( .A(n832), .B(n833), .Z(n854) );
  XOR U999 ( .A(n855), .B(n854), .Z(n856) );
  XNOR U1000 ( .A(n857), .B(n856), .Z(n826) );
  NAND U1001 ( .A(n816), .B(n815), .Z(n820) );
  NAND U1002 ( .A(n818), .B(n817), .Z(n819) );
  NAND U1003 ( .A(n820), .B(n819), .Z(n827) );
  XNOR U1004 ( .A(n826), .B(n827), .Z(n828) );
  XNOR U1005 ( .A(n829), .B(n828), .Z(n860) );
  XNOR U1006 ( .A(n860), .B(sreg[137]), .Z(n862) );
  NAND U1007 ( .A(n821), .B(sreg[136]), .Z(n825) );
  OR U1008 ( .A(n823), .B(n822), .Z(n824) );
  AND U1009 ( .A(n825), .B(n824), .Z(n861) );
  XOR U1010 ( .A(n862), .B(n861), .Z(c[137]) );
  NANDN U1011 ( .A(n831), .B(n830), .Z(n835) );
  NAND U1012 ( .A(n833), .B(n832), .Z(n834) );
  NAND U1013 ( .A(n835), .B(n834), .Z(n896) );
  NANDN U1014 ( .A(n837), .B(n836), .Z(n841) );
  NAND U1015 ( .A(n839), .B(n838), .Z(n840) );
  NAND U1016 ( .A(n841), .B(n840), .Z(n894) );
  XNOR U1017 ( .A(b[7]), .B(a[12]), .Z(n881) );
  NANDN U1018 ( .A(n881), .B(n5293), .Z(n844) );
  NANDN U1019 ( .A(n842), .B(n5294), .Z(n843) );
  NAND U1020 ( .A(n844), .B(n843), .Z(n869) );
  XNOR U1021 ( .A(b[3]), .B(a[16]), .Z(n884) );
  NANDN U1022 ( .A(n884), .B(n5160), .Z(n847) );
  NANDN U1023 ( .A(n845), .B(n5161), .Z(n846) );
  AND U1024 ( .A(n847), .B(n846), .Z(n870) );
  XNOR U1025 ( .A(n869), .B(n870), .Z(n871) );
  NANDN U1026 ( .A(n292), .B(a[18]), .Z(n848) );
  XOR U1027 ( .A(n5199), .B(n848), .Z(n850) );
  NANDN U1028 ( .A(b[0]), .B(a[17]), .Z(n849) );
  AND U1029 ( .A(n850), .B(n849), .Z(n877) );
  XNOR U1030 ( .A(b[5]), .B(a[14]), .Z(n890) );
  NANDN U1031 ( .A(n890), .B(n5240), .Z(n853) );
  NANDN U1032 ( .A(n851), .B(n5241), .Z(n852) );
  NAND U1033 ( .A(n853), .B(n852), .Z(n875) );
  NANDN U1034 ( .A(n295), .B(a[10]), .Z(n876) );
  XNOR U1035 ( .A(n875), .B(n876), .Z(n878) );
  XOR U1036 ( .A(n877), .B(n878), .Z(n872) );
  XOR U1037 ( .A(n871), .B(n872), .Z(n893) );
  XOR U1038 ( .A(n894), .B(n893), .Z(n895) );
  XNOR U1039 ( .A(n896), .B(n895), .Z(n865) );
  NAND U1040 ( .A(n855), .B(n854), .Z(n859) );
  NAND U1041 ( .A(n857), .B(n856), .Z(n858) );
  NAND U1042 ( .A(n859), .B(n858), .Z(n866) );
  XNOR U1043 ( .A(n865), .B(n866), .Z(n867) );
  XNOR U1044 ( .A(n868), .B(n867), .Z(n899) );
  XNOR U1045 ( .A(n899), .B(sreg[138]), .Z(n901) );
  NAND U1046 ( .A(n860), .B(sreg[137]), .Z(n864) );
  OR U1047 ( .A(n862), .B(n861), .Z(n863) );
  AND U1048 ( .A(n864), .B(n863), .Z(n900) );
  XOR U1049 ( .A(n901), .B(n900), .Z(c[138]) );
  NANDN U1050 ( .A(n870), .B(n869), .Z(n874) );
  NAND U1051 ( .A(n872), .B(n871), .Z(n873) );
  NAND U1052 ( .A(n874), .B(n873), .Z(n935) );
  NANDN U1053 ( .A(n876), .B(n875), .Z(n880) );
  NAND U1054 ( .A(n878), .B(n877), .Z(n879) );
  NAND U1055 ( .A(n880), .B(n879), .Z(n933) );
  XNOR U1056 ( .A(b[7]), .B(a[13]), .Z(n920) );
  NANDN U1057 ( .A(n920), .B(n5293), .Z(n883) );
  NANDN U1058 ( .A(n881), .B(n5294), .Z(n882) );
  NAND U1059 ( .A(n883), .B(n882), .Z(n908) );
  XNOR U1060 ( .A(b[3]), .B(a[17]), .Z(n923) );
  NANDN U1061 ( .A(n923), .B(n5160), .Z(n886) );
  NANDN U1062 ( .A(n884), .B(n5161), .Z(n885) );
  AND U1063 ( .A(n886), .B(n885), .Z(n909) );
  XNOR U1064 ( .A(n908), .B(n909), .Z(n910) );
  NANDN U1065 ( .A(n292), .B(a[19]), .Z(n887) );
  XOR U1066 ( .A(n5199), .B(n887), .Z(n889) );
  NANDN U1067 ( .A(b[0]), .B(a[18]), .Z(n888) );
  AND U1068 ( .A(n889), .B(n888), .Z(n916) );
  XNOR U1069 ( .A(b[5]), .B(a[15]), .Z(n929) );
  NANDN U1070 ( .A(n929), .B(n5240), .Z(n892) );
  NANDN U1071 ( .A(n890), .B(n5241), .Z(n891) );
  NAND U1072 ( .A(n892), .B(n891), .Z(n914) );
  NANDN U1073 ( .A(n295), .B(a[11]), .Z(n915) );
  XNOR U1074 ( .A(n914), .B(n915), .Z(n917) );
  XOR U1075 ( .A(n916), .B(n917), .Z(n911) );
  XOR U1076 ( .A(n910), .B(n911), .Z(n932) );
  XOR U1077 ( .A(n933), .B(n932), .Z(n934) );
  XNOR U1078 ( .A(n935), .B(n934), .Z(n904) );
  NAND U1079 ( .A(n894), .B(n893), .Z(n898) );
  NAND U1080 ( .A(n896), .B(n895), .Z(n897) );
  NAND U1081 ( .A(n898), .B(n897), .Z(n905) );
  XNOR U1082 ( .A(n904), .B(n905), .Z(n906) );
  XNOR U1083 ( .A(n907), .B(n906), .Z(n938) );
  XNOR U1084 ( .A(n938), .B(sreg[139]), .Z(n940) );
  NAND U1085 ( .A(n899), .B(sreg[138]), .Z(n903) );
  OR U1086 ( .A(n901), .B(n900), .Z(n902) );
  AND U1087 ( .A(n903), .B(n902), .Z(n939) );
  XOR U1088 ( .A(n940), .B(n939), .Z(c[139]) );
  NANDN U1089 ( .A(n909), .B(n908), .Z(n913) );
  NAND U1090 ( .A(n911), .B(n910), .Z(n912) );
  NAND U1091 ( .A(n913), .B(n912), .Z(n974) );
  NANDN U1092 ( .A(n915), .B(n914), .Z(n919) );
  NAND U1093 ( .A(n917), .B(n916), .Z(n918) );
  NAND U1094 ( .A(n919), .B(n918), .Z(n972) );
  XNOR U1095 ( .A(b[7]), .B(a[14]), .Z(n959) );
  NANDN U1096 ( .A(n959), .B(n5293), .Z(n922) );
  NANDN U1097 ( .A(n920), .B(n5294), .Z(n921) );
  NAND U1098 ( .A(n922), .B(n921), .Z(n947) );
  XNOR U1099 ( .A(b[3]), .B(a[18]), .Z(n962) );
  NANDN U1100 ( .A(n962), .B(n5160), .Z(n925) );
  NANDN U1101 ( .A(n923), .B(n5161), .Z(n924) );
  AND U1102 ( .A(n925), .B(n924), .Z(n948) );
  XNOR U1103 ( .A(n947), .B(n948), .Z(n949) );
  NANDN U1104 ( .A(n292), .B(a[20]), .Z(n926) );
  XOR U1105 ( .A(n5199), .B(n926), .Z(n928) );
  NANDN U1106 ( .A(b[0]), .B(a[19]), .Z(n927) );
  AND U1107 ( .A(n928), .B(n927), .Z(n955) );
  XNOR U1108 ( .A(b[5]), .B(a[16]), .Z(n968) );
  NANDN U1109 ( .A(n968), .B(n5240), .Z(n931) );
  NANDN U1110 ( .A(n929), .B(n5241), .Z(n930) );
  NAND U1111 ( .A(n931), .B(n930), .Z(n953) );
  NANDN U1112 ( .A(n295), .B(a[12]), .Z(n954) );
  XNOR U1113 ( .A(n953), .B(n954), .Z(n956) );
  XOR U1114 ( .A(n955), .B(n956), .Z(n950) );
  XOR U1115 ( .A(n949), .B(n950), .Z(n971) );
  XOR U1116 ( .A(n972), .B(n971), .Z(n973) );
  XNOR U1117 ( .A(n974), .B(n973), .Z(n943) );
  NAND U1118 ( .A(n933), .B(n932), .Z(n937) );
  NAND U1119 ( .A(n935), .B(n934), .Z(n936) );
  NAND U1120 ( .A(n937), .B(n936), .Z(n944) );
  XNOR U1121 ( .A(n943), .B(n944), .Z(n945) );
  XNOR U1122 ( .A(n946), .B(n945), .Z(n977) );
  XNOR U1123 ( .A(n977), .B(sreg[140]), .Z(n979) );
  NAND U1124 ( .A(n938), .B(sreg[139]), .Z(n942) );
  OR U1125 ( .A(n940), .B(n939), .Z(n941) );
  AND U1126 ( .A(n942), .B(n941), .Z(n978) );
  XOR U1127 ( .A(n979), .B(n978), .Z(c[140]) );
  NANDN U1128 ( .A(n948), .B(n947), .Z(n952) );
  NAND U1129 ( .A(n950), .B(n949), .Z(n951) );
  NAND U1130 ( .A(n952), .B(n951), .Z(n1013) );
  NANDN U1131 ( .A(n954), .B(n953), .Z(n958) );
  NAND U1132 ( .A(n956), .B(n955), .Z(n957) );
  NAND U1133 ( .A(n958), .B(n957), .Z(n1011) );
  XNOR U1134 ( .A(b[7]), .B(a[15]), .Z(n998) );
  NANDN U1135 ( .A(n998), .B(n5293), .Z(n961) );
  NANDN U1136 ( .A(n959), .B(n5294), .Z(n960) );
  NAND U1137 ( .A(n961), .B(n960), .Z(n986) );
  XNOR U1138 ( .A(b[3]), .B(a[19]), .Z(n1001) );
  NANDN U1139 ( .A(n1001), .B(n5160), .Z(n964) );
  NANDN U1140 ( .A(n962), .B(n5161), .Z(n963) );
  AND U1141 ( .A(n964), .B(n963), .Z(n987) );
  XNOR U1142 ( .A(n986), .B(n987), .Z(n988) );
  NANDN U1143 ( .A(n292), .B(a[21]), .Z(n965) );
  XOR U1144 ( .A(n5199), .B(n965), .Z(n967) );
  NANDN U1145 ( .A(b[0]), .B(a[20]), .Z(n966) );
  AND U1146 ( .A(n967), .B(n966), .Z(n994) );
  XNOR U1147 ( .A(b[5]), .B(a[17]), .Z(n1007) );
  NANDN U1148 ( .A(n1007), .B(n5240), .Z(n970) );
  NANDN U1149 ( .A(n968), .B(n5241), .Z(n969) );
  NAND U1150 ( .A(n970), .B(n969), .Z(n992) );
  NANDN U1151 ( .A(n295), .B(a[13]), .Z(n993) );
  XNOR U1152 ( .A(n992), .B(n993), .Z(n995) );
  XOR U1153 ( .A(n994), .B(n995), .Z(n989) );
  XOR U1154 ( .A(n988), .B(n989), .Z(n1010) );
  XOR U1155 ( .A(n1011), .B(n1010), .Z(n1012) );
  XNOR U1156 ( .A(n1013), .B(n1012), .Z(n982) );
  NAND U1157 ( .A(n972), .B(n971), .Z(n976) );
  NAND U1158 ( .A(n974), .B(n973), .Z(n975) );
  NAND U1159 ( .A(n976), .B(n975), .Z(n983) );
  XNOR U1160 ( .A(n982), .B(n983), .Z(n984) );
  XNOR U1161 ( .A(n985), .B(n984), .Z(n1016) );
  XNOR U1162 ( .A(n1016), .B(sreg[141]), .Z(n1018) );
  NAND U1163 ( .A(n977), .B(sreg[140]), .Z(n981) );
  OR U1164 ( .A(n979), .B(n978), .Z(n980) );
  AND U1165 ( .A(n981), .B(n980), .Z(n1017) );
  XOR U1166 ( .A(n1018), .B(n1017), .Z(c[141]) );
  NANDN U1167 ( .A(n987), .B(n986), .Z(n991) );
  NAND U1168 ( .A(n989), .B(n988), .Z(n990) );
  NAND U1169 ( .A(n991), .B(n990), .Z(n1052) );
  NANDN U1170 ( .A(n993), .B(n992), .Z(n997) );
  NAND U1171 ( .A(n995), .B(n994), .Z(n996) );
  NAND U1172 ( .A(n997), .B(n996), .Z(n1050) );
  XNOR U1173 ( .A(b[7]), .B(a[16]), .Z(n1025) );
  NANDN U1174 ( .A(n1025), .B(n5293), .Z(n1000) );
  NANDN U1175 ( .A(n998), .B(n5294), .Z(n999) );
  NAND U1176 ( .A(n1000), .B(n999), .Z(n1043) );
  XNOR U1177 ( .A(b[3]), .B(a[20]), .Z(n1028) );
  NANDN U1178 ( .A(n1028), .B(n5160), .Z(n1003) );
  NANDN U1179 ( .A(n1001), .B(n5161), .Z(n1002) );
  AND U1180 ( .A(n1003), .B(n1002), .Z(n1044) );
  XNOR U1181 ( .A(n1043), .B(n1044), .Z(n1045) );
  NANDN U1182 ( .A(n292), .B(a[22]), .Z(n1004) );
  XOR U1183 ( .A(n5199), .B(n1004), .Z(n1006) );
  NANDN U1184 ( .A(b[0]), .B(a[21]), .Z(n1005) );
  AND U1185 ( .A(n1006), .B(n1005), .Z(n1039) );
  XNOR U1186 ( .A(b[5]), .B(a[18]), .Z(n1034) );
  NANDN U1187 ( .A(n1034), .B(n5240), .Z(n1009) );
  NANDN U1188 ( .A(n1007), .B(n5241), .Z(n1008) );
  NAND U1189 ( .A(n1009), .B(n1008), .Z(n1037) );
  NANDN U1190 ( .A(n295), .B(a[14]), .Z(n1038) );
  XNOR U1191 ( .A(n1037), .B(n1038), .Z(n1040) );
  XOR U1192 ( .A(n1039), .B(n1040), .Z(n1046) );
  XOR U1193 ( .A(n1045), .B(n1046), .Z(n1049) );
  XOR U1194 ( .A(n1050), .B(n1049), .Z(n1051) );
  XNOR U1195 ( .A(n1052), .B(n1051), .Z(n1021) );
  NAND U1196 ( .A(n1011), .B(n1010), .Z(n1015) );
  NAND U1197 ( .A(n1013), .B(n1012), .Z(n1014) );
  NAND U1198 ( .A(n1015), .B(n1014), .Z(n1022) );
  XNOR U1199 ( .A(n1021), .B(n1022), .Z(n1023) );
  XNOR U1200 ( .A(n1024), .B(n1023), .Z(n1055) );
  XNOR U1201 ( .A(n1055), .B(sreg[142]), .Z(n1057) );
  NAND U1202 ( .A(n1016), .B(sreg[141]), .Z(n1020) );
  OR U1203 ( .A(n1018), .B(n1017), .Z(n1019) );
  AND U1204 ( .A(n1020), .B(n1019), .Z(n1056) );
  XOR U1205 ( .A(n1057), .B(n1056), .Z(c[142]) );
  XNOR U1206 ( .A(b[7]), .B(a[17]), .Z(n1076) );
  NANDN U1207 ( .A(n1076), .B(n5293), .Z(n1027) );
  NANDN U1208 ( .A(n1025), .B(n5294), .Z(n1026) );
  NAND U1209 ( .A(n1027), .B(n1026), .Z(n1064) );
  XNOR U1210 ( .A(b[3]), .B(a[21]), .Z(n1079) );
  NANDN U1211 ( .A(n1079), .B(n5160), .Z(n1030) );
  NANDN U1212 ( .A(n1028), .B(n5161), .Z(n1029) );
  AND U1213 ( .A(n1030), .B(n1029), .Z(n1065) );
  XNOR U1214 ( .A(n1064), .B(n1065), .Z(n1066) );
  NANDN U1215 ( .A(n292), .B(a[23]), .Z(n1031) );
  XOR U1216 ( .A(n5199), .B(n1031), .Z(n1033) );
  NANDN U1217 ( .A(b[0]), .B(a[22]), .Z(n1032) );
  AND U1218 ( .A(n1033), .B(n1032), .Z(n1072) );
  XNOR U1219 ( .A(b[5]), .B(a[19]), .Z(n1085) );
  NANDN U1220 ( .A(n1085), .B(n5240), .Z(n1036) );
  NANDN U1221 ( .A(n1034), .B(n5241), .Z(n1035) );
  NAND U1222 ( .A(n1036), .B(n1035), .Z(n1070) );
  NANDN U1223 ( .A(n295), .B(a[15]), .Z(n1071) );
  XNOR U1224 ( .A(n1070), .B(n1071), .Z(n1073) );
  XOR U1225 ( .A(n1072), .B(n1073), .Z(n1067) );
  XOR U1226 ( .A(n1066), .B(n1067), .Z(n1090) );
  NANDN U1227 ( .A(n1038), .B(n1037), .Z(n1042) );
  NAND U1228 ( .A(n1040), .B(n1039), .Z(n1041) );
  NAND U1229 ( .A(n1042), .B(n1041), .Z(n1088) );
  NANDN U1230 ( .A(n1044), .B(n1043), .Z(n1048) );
  NAND U1231 ( .A(n1046), .B(n1045), .Z(n1047) );
  AND U1232 ( .A(n1048), .B(n1047), .Z(n1089) );
  XNOR U1233 ( .A(n1088), .B(n1089), .Z(n1091) );
  XNOR U1234 ( .A(n1090), .B(n1091), .Z(n1060) );
  NAND U1235 ( .A(n1050), .B(n1049), .Z(n1054) );
  NAND U1236 ( .A(n1052), .B(n1051), .Z(n1053) );
  NAND U1237 ( .A(n1054), .B(n1053), .Z(n1061) );
  XNOR U1238 ( .A(n1060), .B(n1061), .Z(n1062) );
  XNOR U1239 ( .A(n1063), .B(n1062), .Z(n1094) );
  XNOR U1240 ( .A(n1094), .B(sreg[143]), .Z(n1096) );
  NAND U1241 ( .A(n1055), .B(sreg[142]), .Z(n1059) );
  OR U1242 ( .A(n1057), .B(n1056), .Z(n1058) );
  AND U1243 ( .A(n1059), .B(n1058), .Z(n1095) );
  XOR U1244 ( .A(n1096), .B(n1095), .Z(c[143]) );
  NANDN U1245 ( .A(n1065), .B(n1064), .Z(n1069) );
  NAND U1246 ( .A(n1067), .B(n1066), .Z(n1068) );
  NAND U1247 ( .A(n1069), .B(n1068), .Z(n1130) );
  NANDN U1248 ( .A(n1071), .B(n1070), .Z(n1075) );
  NAND U1249 ( .A(n1073), .B(n1072), .Z(n1074) );
  NAND U1250 ( .A(n1075), .B(n1074), .Z(n1128) );
  XNOR U1251 ( .A(b[7]), .B(a[18]), .Z(n1115) );
  NANDN U1252 ( .A(n1115), .B(n5293), .Z(n1078) );
  NANDN U1253 ( .A(n1076), .B(n5294), .Z(n1077) );
  NAND U1254 ( .A(n1078), .B(n1077), .Z(n1103) );
  XNOR U1255 ( .A(b[3]), .B(a[22]), .Z(n1118) );
  NANDN U1256 ( .A(n1118), .B(n5160), .Z(n1081) );
  NANDN U1257 ( .A(n1079), .B(n5161), .Z(n1080) );
  AND U1258 ( .A(n1081), .B(n1080), .Z(n1104) );
  XNOR U1259 ( .A(n1103), .B(n1104), .Z(n1105) );
  NANDN U1260 ( .A(n292), .B(a[24]), .Z(n1082) );
  XOR U1261 ( .A(n5199), .B(n1082), .Z(n1084) );
  NANDN U1262 ( .A(b[0]), .B(a[23]), .Z(n1083) );
  AND U1263 ( .A(n1084), .B(n1083), .Z(n1111) );
  XNOR U1264 ( .A(b[5]), .B(a[20]), .Z(n1124) );
  NANDN U1265 ( .A(n1124), .B(n5240), .Z(n1087) );
  NANDN U1266 ( .A(n1085), .B(n5241), .Z(n1086) );
  NAND U1267 ( .A(n1087), .B(n1086), .Z(n1109) );
  NANDN U1268 ( .A(n295), .B(a[16]), .Z(n1110) );
  XNOR U1269 ( .A(n1109), .B(n1110), .Z(n1112) );
  XOR U1270 ( .A(n1111), .B(n1112), .Z(n1106) );
  XOR U1271 ( .A(n1105), .B(n1106), .Z(n1127) );
  XOR U1272 ( .A(n1128), .B(n1127), .Z(n1129) );
  XNOR U1273 ( .A(n1130), .B(n1129), .Z(n1099) );
  NANDN U1274 ( .A(n1089), .B(n1088), .Z(n1093) );
  NAND U1275 ( .A(n1091), .B(n1090), .Z(n1092) );
  NAND U1276 ( .A(n1093), .B(n1092), .Z(n1100) );
  XNOR U1277 ( .A(n1099), .B(n1100), .Z(n1101) );
  XNOR U1278 ( .A(n1102), .B(n1101), .Z(n1133) );
  XNOR U1279 ( .A(n1133), .B(sreg[144]), .Z(n1135) );
  NAND U1280 ( .A(n1094), .B(sreg[143]), .Z(n1098) );
  OR U1281 ( .A(n1096), .B(n1095), .Z(n1097) );
  AND U1282 ( .A(n1098), .B(n1097), .Z(n1134) );
  XOR U1283 ( .A(n1135), .B(n1134), .Z(c[144]) );
  NANDN U1284 ( .A(n1104), .B(n1103), .Z(n1108) );
  NAND U1285 ( .A(n1106), .B(n1105), .Z(n1107) );
  NAND U1286 ( .A(n1108), .B(n1107), .Z(n1169) );
  NANDN U1287 ( .A(n1110), .B(n1109), .Z(n1114) );
  NAND U1288 ( .A(n1112), .B(n1111), .Z(n1113) );
  NAND U1289 ( .A(n1114), .B(n1113), .Z(n1167) );
  XNOR U1290 ( .A(b[7]), .B(a[19]), .Z(n1154) );
  NANDN U1291 ( .A(n1154), .B(n5293), .Z(n1117) );
  NANDN U1292 ( .A(n1115), .B(n5294), .Z(n1116) );
  NAND U1293 ( .A(n1117), .B(n1116), .Z(n1142) );
  XNOR U1294 ( .A(b[3]), .B(a[23]), .Z(n1157) );
  NANDN U1295 ( .A(n1157), .B(n5160), .Z(n1120) );
  NANDN U1296 ( .A(n1118), .B(n5161), .Z(n1119) );
  AND U1297 ( .A(n1120), .B(n1119), .Z(n1143) );
  XNOR U1298 ( .A(n1142), .B(n1143), .Z(n1144) );
  NANDN U1299 ( .A(n292), .B(a[25]), .Z(n1121) );
  XOR U1300 ( .A(n5199), .B(n1121), .Z(n1123) );
  NANDN U1301 ( .A(b[0]), .B(a[24]), .Z(n1122) );
  AND U1302 ( .A(n1123), .B(n1122), .Z(n1150) );
  XNOR U1303 ( .A(b[5]), .B(a[21]), .Z(n1163) );
  NANDN U1304 ( .A(n1163), .B(n5240), .Z(n1126) );
  NANDN U1305 ( .A(n1124), .B(n5241), .Z(n1125) );
  NAND U1306 ( .A(n1126), .B(n1125), .Z(n1148) );
  NANDN U1307 ( .A(n295), .B(a[17]), .Z(n1149) );
  XNOR U1308 ( .A(n1148), .B(n1149), .Z(n1151) );
  XOR U1309 ( .A(n1150), .B(n1151), .Z(n1145) );
  XOR U1310 ( .A(n1144), .B(n1145), .Z(n1166) );
  XOR U1311 ( .A(n1167), .B(n1166), .Z(n1168) );
  XNOR U1312 ( .A(n1169), .B(n1168), .Z(n1138) );
  NAND U1313 ( .A(n1128), .B(n1127), .Z(n1132) );
  NAND U1314 ( .A(n1130), .B(n1129), .Z(n1131) );
  NAND U1315 ( .A(n1132), .B(n1131), .Z(n1139) );
  XNOR U1316 ( .A(n1138), .B(n1139), .Z(n1140) );
  XNOR U1317 ( .A(n1141), .B(n1140), .Z(n1172) );
  XNOR U1318 ( .A(n1172), .B(sreg[145]), .Z(n1174) );
  NAND U1319 ( .A(n1133), .B(sreg[144]), .Z(n1137) );
  OR U1320 ( .A(n1135), .B(n1134), .Z(n1136) );
  AND U1321 ( .A(n1137), .B(n1136), .Z(n1173) );
  XOR U1322 ( .A(n1174), .B(n1173), .Z(c[145]) );
  NANDN U1323 ( .A(n1143), .B(n1142), .Z(n1147) );
  NAND U1324 ( .A(n1145), .B(n1144), .Z(n1146) );
  NAND U1325 ( .A(n1147), .B(n1146), .Z(n1208) );
  NANDN U1326 ( .A(n1149), .B(n1148), .Z(n1153) );
  NAND U1327 ( .A(n1151), .B(n1150), .Z(n1152) );
  NAND U1328 ( .A(n1153), .B(n1152), .Z(n1206) );
  XNOR U1329 ( .A(b[7]), .B(a[20]), .Z(n1193) );
  NANDN U1330 ( .A(n1193), .B(n5293), .Z(n1156) );
  NANDN U1331 ( .A(n1154), .B(n5294), .Z(n1155) );
  NAND U1332 ( .A(n1156), .B(n1155), .Z(n1181) );
  XNOR U1333 ( .A(b[3]), .B(a[24]), .Z(n1196) );
  NANDN U1334 ( .A(n1196), .B(n5160), .Z(n1159) );
  NANDN U1335 ( .A(n1157), .B(n5161), .Z(n1158) );
  AND U1336 ( .A(n1159), .B(n1158), .Z(n1182) );
  XNOR U1337 ( .A(n1181), .B(n1182), .Z(n1183) );
  NANDN U1338 ( .A(n292), .B(a[26]), .Z(n1160) );
  XOR U1339 ( .A(n5199), .B(n1160), .Z(n1162) );
  NANDN U1340 ( .A(b[0]), .B(a[25]), .Z(n1161) );
  AND U1341 ( .A(n1162), .B(n1161), .Z(n1189) );
  XNOR U1342 ( .A(b[5]), .B(a[22]), .Z(n1202) );
  NANDN U1343 ( .A(n1202), .B(n5240), .Z(n1165) );
  NANDN U1344 ( .A(n1163), .B(n5241), .Z(n1164) );
  NAND U1345 ( .A(n1165), .B(n1164), .Z(n1187) );
  NANDN U1346 ( .A(n295), .B(a[18]), .Z(n1188) );
  XNOR U1347 ( .A(n1187), .B(n1188), .Z(n1190) );
  XOR U1348 ( .A(n1189), .B(n1190), .Z(n1184) );
  XOR U1349 ( .A(n1183), .B(n1184), .Z(n1205) );
  XOR U1350 ( .A(n1206), .B(n1205), .Z(n1207) );
  XNOR U1351 ( .A(n1208), .B(n1207), .Z(n1177) );
  NAND U1352 ( .A(n1167), .B(n1166), .Z(n1171) );
  NAND U1353 ( .A(n1169), .B(n1168), .Z(n1170) );
  NAND U1354 ( .A(n1171), .B(n1170), .Z(n1178) );
  XNOR U1355 ( .A(n1177), .B(n1178), .Z(n1179) );
  XNOR U1356 ( .A(n1180), .B(n1179), .Z(n1211) );
  XNOR U1357 ( .A(n1211), .B(sreg[146]), .Z(n1213) );
  NAND U1358 ( .A(n1172), .B(sreg[145]), .Z(n1176) );
  OR U1359 ( .A(n1174), .B(n1173), .Z(n1175) );
  AND U1360 ( .A(n1176), .B(n1175), .Z(n1212) );
  XOR U1361 ( .A(n1213), .B(n1212), .Z(c[146]) );
  NANDN U1362 ( .A(n1182), .B(n1181), .Z(n1186) );
  NAND U1363 ( .A(n1184), .B(n1183), .Z(n1185) );
  NAND U1364 ( .A(n1186), .B(n1185), .Z(n1247) );
  NANDN U1365 ( .A(n1188), .B(n1187), .Z(n1192) );
  NAND U1366 ( .A(n1190), .B(n1189), .Z(n1191) );
  NAND U1367 ( .A(n1192), .B(n1191), .Z(n1245) );
  XNOR U1368 ( .A(b[7]), .B(a[21]), .Z(n1238) );
  NANDN U1369 ( .A(n1238), .B(n5293), .Z(n1195) );
  NANDN U1370 ( .A(n1193), .B(n5294), .Z(n1194) );
  NAND U1371 ( .A(n1195), .B(n1194), .Z(n1220) );
  XNOR U1372 ( .A(b[3]), .B(a[25]), .Z(n1241) );
  NANDN U1373 ( .A(n1241), .B(n5160), .Z(n1198) );
  NANDN U1374 ( .A(n1196), .B(n5161), .Z(n1197) );
  AND U1375 ( .A(n1198), .B(n1197), .Z(n1221) );
  XNOR U1376 ( .A(n1220), .B(n1221), .Z(n1222) );
  NANDN U1377 ( .A(n292), .B(a[27]), .Z(n1199) );
  XOR U1378 ( .A(n5199), .B(n1199), .Z(n1201) );
  NANDN U1379 ( .A(b[0]), .B(a[26]), .Z(n1200) );
  AND U1380 ( .A(n1201), .B(n1200), .Z(n1228) );
  XNOR U1381 ( .A(b[5]), .B(a[23]), .Z(n1235) );
  NANDN U1382 ( .A(n1235), .B(n5240), .Z(n1204) );
  NANDN U1383 ( .A(n1202), .B(n5241), .Z(n1203) );
  NAND U1384 ( .A(n1204), .B(n1203), .Z(n1226) );
  NANDN U1385 ( .A(n295), .B(a[19]), .Z(n1227) );
  XNOR U1386 ( .A(n1226), .B(n1227), .Z(n1229) );
  XOR U1387 ( .A(n1228), .B(n1229), .Z(n1223) );
  XOR U1388 ( .A(n1222), .B(n1223), .Z(n1244) );
  XOR U1389 ( .A(n1245), .B(n1244), .Z(n1246) );
  XNOR U1390 ( .A(n1247), .B(n1246), .Z(n1216) );
  NAND U1391 ( .A(n1206), .B(n1205), .Z(n1210) );
  NAND U1392 ( .A(n1208), .B(n1207), .Z(n1209) );
  NAND U1393 ( .A(n1210), .B(n1209), .Z(n1217) );
  XNOR U1394 ( .A(n1216), .B(n1217), .Z(n1218) );
  XNOR U1395 ( .A(n1219), .B(n1218), .Z(n1250) );
  XNOR U1396 ( .A(n1250), .B(sreg[147]), .Z(n1252) );
  NAND U1397 ( .A(n1211), .B(sreg[146]), .Z(n1215) );
  OR U1398 ( .A(n1213), .B(n1212), .Z(n1214) );
  AND U1399 ( .A(n1215), .B(n1214), .Z(n1251) );
  XOR U1400 ( .A(n1252), .B(n1251), .Z(c[147]) );
  NANDN U1401 ( .A(n1221), .B(n1220), .Z(n1225) );
  NAND U1402 ( .A(n1223), .B(n1222), .Z(n1224) );
  NAND U1403 ( .A(n1225), .B(n1224), .Z(n1286) );
  NANDN U1404 ( .A(n1227), .B(n1226), .Z(n1231) );
  NAND U1405 ( .A(n1229), .B(n1228), .Z(n1230) );
  NAND U1406 ( .A(n1231), .B(n1230), .Z(n1284) );
  NANDN U1407 ( .A(n292), .B(a[28]), .Z(n1232) );
  XOR U1408 ( .A(n5199), .B(n1232), .Z(n1234) );
  NANDN U1409 ( .A(b[0]), .B(a[27]), .Z(n1233) );
  AND U1410 ( .A(n1234), .B(n1233), .Z(n1267) );
  XNOR U1411 ( .A(b[5]), .B(a[24]), .Z(n1280) );
  NANDN U1412 ( .A(n1280), .B(n5240), .Z(n1237) );
  NANDN U1413 ( .A(n1235), .B(n5241), .Z(n1236) );
  NAND U1414 ( .A(n1237), .B(n1236), .Z(n1265) );
  NANDN U1415 ( .A(n295), .B(a[20]), .Z(n1266) );
  XNOR U1416 ( .A(n1265), .B(n1266), .Z(n1268) );
  XOR U1417 ( .A(n1267), .B(n1268), .Z(n1261) );
  XNOR U1418 ( .A(b[7]), .B(a[22]), .Z(n1271) );
  NANDN U1419 ( .A(n1271), .B(n5293), .Z(n1240) );
  NANDN U1420 ( .A(n1238), .B(n5294), .Z(n1239) );
  NAND U1421 ( .A(n1240), .B(n1239), .Z(n1259) );
  XNOR U1422 ( .A(b[3]), .B(a[26]), .Z(n1274) );
  NANDN U1423 ( .A(n1274), .B(n5160), .Z(n1243) );
  NANDN U1424 ( .A(n1241), .B(n5161), .Z(n1242) );
  AND U1425 ( .A(n1243), .B(n1242), .Z(n1260) );
  XNOR U1426 ( .A(n1259), .B(n1260), .Z(n1262) );
  XOR U1427 ( .A(n1261), .B(n1262), .Z(n1283) );
  XOR U1428 ( .A(n1284), .B(n1283), .Z(n1285) );
  XNOR U1429 ( .A(n1286), .B(n1285), .Z(n1255) );
  NAND U1430 ( .A(n1245), .B(n1244), .Z(n1249) );
  NAND U1431 ( .A(n1247), .B(n1246), .Z(n1248) );
  NAND U1432 ( .A(n1249), .B(n1248), .Z(n1256) );
  XNOR U1433 ( .A(n1255), .B(n1256), .Z(n1257) );
  XNOR U1434 ( .A(n1258), .B(n1257), .Z(n1289) );
  XNOR U1435 ( .A(n1289), .B(sreg[148]), .Z(n1291) );
  NAND U1436 ( .A(n1250), .B(sreg[147]), .Z(n1254) );
  OR U1437 ( .A(n1252), .B(n1251), .Z(n1253) );
  AND U1438 ( .A(n1254), .B(n1253), .Z(n1290) );
  XOR U1439 ( .A(n1291), .B(n1290), .Z(c[148]) );
  NANDN U1440 ( .A(n1260), .B(n1259), .Z(n1264) );
  NAND U1441 ( .A(n1262), .B(n1261), .Z(n1263) );
  NAND U1442 ( .A(n1264), .B(n1263), .Z(n1325) );
  NANDN U1443 ( .A(n1266), .B(n1265), .Z(n1270) );
  NAND U1444 ( .A(n1268), .B(n1267), .Z(n1269) );
  NAND U1445 ( .A(n1270), .B(n1269), .Z(n1323) );
  XNOR U1446 ( .A(b[7]), .B(a[23]), .Z(n1310) );
  NANDN U1447 ( .A(n1310), .B(n5293), .Z(n1273) );
  NANDN U1448 ( .A(n1271), .B(n5294), .Z(n1272) );
  NAND U1449 ( .A(n1273), .B(n1272), .Z(n1298) );
  XNOR U1450 ( .A(b[3]), .B(a[27]), .Z(n1313) );
  NANDN U1451 ( .A(n1313), .B(n5160), .Z(n1276) );
  NANDN U1452 ( .A(n1274), .B(n5161), .Z(n1275) );
  AND U1453 ( .A(n1276), .B(n1275), .Z(n1299) );
  XNOR U1454 ( .A(n1298), .B(n1299), .Z(n1300) );
  NANDN U1455 ( .A(n292), .B(a[29]), .Z(n1277) );
  XOR U1456 ( .A(n5199), .B(n1277), .Z(n1279) );
  NANDN U1457 ( .A(b[0]), .B(a[28]), .Z(n1278) );
  AND U1458 ( .A(n1279), .B(n1278), .Z(n1306) );
  XNOR U1459 ( .A(b[5]), .B(a[25]), .Z(n1319) );
  NANDN U1460 ( .A(n1319), .B(n5240), .Z(n1282) );
  NANDN U1461 ( .A(n1280), .B(n5241), .Z(n1281) );
  NAND U1462 ( .A(n1282), .B(n1281), .Z(n1304) );
  NANDN U1463 ( .A(n295), .B(a[21]), .Z(n1305) );
  XNOR U1464 ( .A(n1304), .B(n1305), .Z(n1307) );
  XOR U1465 ( .A(n1306), .B(n1307), .Z(n1301) );
  XOR U1466 ( .A(n1300), .B(n1301), .Z(n1322) );
  XOR U1467 ( .A(n1323), .B(n1322), .Z(n1324) );
  XNOR U1468 ( .A(n1325), .B(n1324), .Z(n1294) );
  NAND U1469 ( .A(n1284), .B(n1283), .Z(n1288) );
  NAND U1470 ( .A(n1286), .B(n1285), .Z(n1287) );
  NAND U1471 ( .A(n1288), .B(n1287), .Z(n1295) );
  XNOR U1472 ( .A(n1294), .B(n1295), .Z(n1296) );
  XNOR U1473 ( .A(n1297), .B(n1296), .Z(n1328) );
  XNOR U1474 ( .A(n1328), .B(sreg[149]), .Z(n1330) );
  NAND U1475 ( .A(n1289), .B(sreg[148]), .Z(n1293) );
  OR U1476 ( .A(n1291), .B(n1290), .Z(n1292) );
  AND U1477 ( .A(n1293), .B(n1292), .Z(n1329) );
  XOR U1478 ( .A(n1330), .B(n1329), .Z(c[149]) );
  NANDN U1479 ( .A(n1299), .B(n1298), .Z(n1303) );
  NAND U1480 ( .A(n1301), .B(n1300), .Z(n1302) );
  NAND U1481 ( .A(n1303), .B(n1302), .Z(n1364) );
  NANDN U1482 ( .A(n1305), .B(n1304), .Z(n1309) );
  NAND U1483 ( .A(n1307), .B(n1306), .Z(n1308) );
  NAND U1484 ( .A(n1309), .B(n1308), .Z(n1362) );
  XNOR U1485 ( .A(b[7]), .B(a[24]), .Z(n1355) );
  NANDN U1486 ( .A(n1355), .B(n5293), .Z(n1312) );
  NANDN U1487 ( .A(n1310), .B(n5294), .Z(n1311) );
  NAND U1488 ( .A(n1312), .B(n1311), .Z(n1337) );
  XNOR U1489 ( .A(b[3]), .B(a[28]), .Z(n1358) );
  NANDN U1490 ( .A(n1358), .B(n5160), .Z(n1315) );
  NANDN U1491 ( .A(n1313), .B(n5161), .Z(n1314) );
  AND U1492 ( .A(n1315), .B(n1314), .Z(n1338) );
  XNOR U1493 ( .A(n1337), .B(n1338), .Z(n1339) );
  NANDN U1494 ( .A(n292), .B(a[30]), .Z(n1316) );
  XOR U1495 ( .A(n5199), .B(n1316), .Z(n1318) );
  NANDN U1496 ( .A(b[0]), .B(a[29]), .Z(n1317) );
  AND U1497 ( .A(n1318), .B(n1317), .Z(n1345) );
  XNOR U1498 ( .A(b[5]), .B(a[26]), .Z(n1352) );
  NANDN U1499 ( .A(n1352), .B(n5240), .Z(n1321) );
  NANDN U1500 ( .A(n1319), .B(n5241), .Z(n1320) );
  NAND U1501 ( .A(n1321), .B(n1320), .Z(n1343) );
  NANDN U1502 ( .A(n295), .B(a[22]), .Z(n1344) );
  XNOR U1503 ( .A(n1343), .B(n1344), .Z(n1346) );
  XOR U1504 ( .A(n1345), .B(n1346), .Z(n1340) );
  XOR U1505 ( .A(n1339), .B(n1340), .Z(n1361) );
  XOR U1506 ( .A(n1362), .B(n1361), .Z(n1363) );
  XNOR U1507 ( .A(n1364), .B(n1363), .Z(n1333) );
  NAND U1508 ( .A(n1323), .B(n1322), .Z(n1327) );
  NAND U1509 ( .A(n1325), .B(n1324), .Z(n1326) );
  NAND U1510 ( .A(n1327), .B(n1326), .Z(n1334) );
  XNOR U1511 ( .A(n1333), .B(n1334), .Z(n1335) );
  XNOR U1512 ( .A(n1336), .B(n1335), .Z(n1367) );
  XNOR U1513 ( .A(n1367), .B(sreg[150]), .Z(n1369) );
  NAND U1514 ( .A(n1328), .B(sreg[149]), .Z(n1332) );
  OR U1515 ( .A(n1330), .B(n1329), .Z(n1331) );
  AND U1516 ( .A(n1332), .B(n1331), .Z(n1368) );
  XOR U1517 ( .A(n1369), .B(n1368), .Z(c[150]) );
  NANDN U1518 ( .A(n1338), .B(n1337), .Z(n1342) );
  NAND U1519 ( .A(n1340), .B(n1339), .Z(n1341) );
  NAND U1520 ( .A(n1342), .B(n1341), .Z(n1403) );
  NANDN U1521 ( .A(n1344), .B(n1343), .Z(n1348) );
  NAND U1522 ( .A(n1346), .B(n1345), .Z(n1347) );
  NAND U1523 ( .A(n1348), .B(n1347), .Z(n1401) );
  NANDN U1524 ( .A(n292), .B(a[31]), .Z(n1349) );
  XOR U1525 ( .A(n5199), .B(n1349), .Z(n1351) );
  NANDN U1526 ( .A(b[0]), .B(a[30]), .Z(n1350) );
  AND U1527 ( .A(n1351), .B(n1350), .Z(n1384) );
  XNOR U1528 ( .A(b[5]), .B(a[27]), .Z(n1397) );
  NANDN U1529 ( .A(n1397), .B(n5240), .Z(n1354) );
  NANDN U1530 ( .A(n1352), .B(n5241), .Z(n1353) );
  NAND U1531 ( .A(n1354), .B(n1353), .Z(n1382) );
  NANDN U1532 ( .A(n295), .B(a[23]), .Z(n1383) );
  XNOR U1533 ( .A(n1382), .B(n1383), .Z(n1385) );
  XOR U1534 ( .A(n1384), .B(n1385), .Z(n1378) );
  XNOR U1535 ( .A(b[7]), .B(a[25]), .Z(n1388) );
  NANDN U1536 ( .A(n1388), .B(n5293), .Z(n1357) );
  NANDN U1537 ( .A(n1355), .B(n5294), .Z(n1356) );
  NAND U1538 ( .A(n1357), .B(n1356), .Z(n1376) );
  XNOR U1539 ( .A(b[3]), .B(a[29]), .Z(n1391) );
  NANDN U1540 ( .A(n1391), .B(n5160), .Z(n1360) );
  NANDN U1541 ( .A(n1358), .B(n5161), .Z(n1359) );
  AND U1542 ( .A(n1360), .B(n1359), .Z(n1377) );
  XNOR U1543 ( .A(n1376), .B(n1377), .Z(n1379) );
  XOR U1544 ( .A(n1378), .B(n1379), .Z(n1400) );
  XOR U1545 ( .A(n1401), .B(n1400), .Z(n1402) );
  XNOR U1546 ( .A(n1403), .B(n1402), .Z(n1372) );
  NAND U1547 ( .A(n1362), .B(n1361), .Z(n1366) );
  NAND U1548 ( .A(n1364), .B(n1363), .Z(n1365) );
  NAND U1549 ( .A(n1366), .B(n1365), .Z(n1373) );
  XNOR U1550 ( .A(n1372), .B(n1373), .Z(n1374) );
  XNOR U1551 ( .A(n1375), .B(n1374), .Z(n1406) );
  XNOR U1552 ( .A(n1406), .B(sreg[151]), .Z(n1408) );
  NAND U1553 ( .A(n1367), .B(sreg[150]), .Z(n1371) );
  OR U1554 ( .A(n1369), .B(n1368), .Z(n1370) );
  AND U1555 ( .A(n1371), .B(n1370), .Z(n1407) );
  XOR U1556 ( .A(n1408), .B(n1407), .Z(c[151]) );
  NANDN U1557 ( .A(n1377), .B(n1376), .Z(n1381) );
  NAND U1558 ( .A(n1379), .B(n1378), .Z(n1380) );
  NAND U1559 ( .A(n1381), .B(n1380), .Z(n1442) );
  NANDN U1560 ( .A(n1383), .B(n1382), .Z(n1387) );
  NAND U1561 ( .A(n1385), .B(n1384), .Z(n1386) );
  NAND U1562 ( .A(n1387), .B(n1386), .Z(n1440) );
  XNOR U1563 ( .A(b[7]), .B(a[26]), .Z(n1427) );
  NANDN U1564 ( .A(n1427), .B(n5293), .Z(n1390) );
  NANDN U1565 ( .A(n1388), .B(n5294), .Z(n1389) );
  NAND U1566 ( .A(n1390), .B(n1389), .Z(n1415) );
  XNOR U1567 ( .A(b[3]), .B(a[30]), .Z(n1430) );
  NANDN U1568 ( .A(n1430), .B(n5160), .Z(n1393) );
  NANDN U1569 ( .A(n1391), .B(n5161), .Z(n1392) );
  AND U1570 ( .A(n1393), .B(n1392), .Z(n1416) );
  XNOR U1571 ( .A(n1415), .B(n1416), .Z(n1417) );
  NANDN U1572 ( .A(n292), .B(a[32]), .Z(n1394) );
  XOR U1573 ( .A(n5199), .B(n1394), .Z(n1396) );
  NANDN U1574 ( .A(b[0]), .B(a[31]), .Z(n1395) );
  AND U1575 ( .A(n1396), .B(n1395), .Z(n1423) );
  XNOR U1576 ( .A(b[5]), .B(a[28]), .Z(n1436) );
  NANDN U1577 ( .A(n1436), .B(n5240), .Z(n1399) );
  NANDN U1578 ( .A(n1397), .B(n5241), .Z(n1398) );
  NAND U1579 ( .A(n1399), .B(n1398), .Z(n1421) );
  NANDN U1580 ( .A(n295), .B(a[24]), .Z(n1422) );
  XNOR U1581 ( .A(n1421), .B(n1422), .Z(n1424) );
  XOR U1582 ( .A(n1423), .B(n1424), .Z(n1418) );
  XOR U1583 ( .A(n1417), .B(n1418), .Z(n1439) );
  XOR U1584 ( .A(n1440), .B(n1439), .Z(n1441) );
  XNOR U1585 ( .A(n1442), .B(n1441), .Z(n1411) );
  NAND U1586 ( .A(n1401), .B(n1400), .Z(n1405) );
  NAND U1587 ( .A(n1403), .B(n1402), .Z(n1404) );
  NAND U1588 ( .A(n1405), .B(n1404), .Z(n1412) );
  XNOR U1589 ( .A(n1411), .B(n1412), .Z(n1413) );
  XNOR U1590 ( .A(n1414), .B(n1413), .Z(n1445) );
  XNOR U1591 ( .A(n1445), .B(sreg[152]), .Z(n1447) );
  NAND U1592 ( .A(n1406), .B(sreg[151]), .Z(n1410) );
  OR U1593 ( .A(n1408), .B(n1407), .Z(n1409) );
  AND U1594 ( .A(n1410), .B(n1409), .Z(n1446) );
  XOR U1595 ( .A(n1447), .B(n1446), .Z(c[152]) );
  NANDN U1596 ( .A(n1416), .B(n1415), .Z(n1420) );
  NAND U1597 ( .A(n1418), .B(n1417), .Z(n1419) );
  NAND U1598 ( .A(n1420), .B(n1419), .Z(n1481) );
  NANDN U1599 ( .A(n1422), .B(n1421), .Z(n1426) );
  NAND U1600 ( .A(n1424), .B(n1423), .Z(n1425) );
  NAND U1601 ( .A(n1426), .B(n1425), .Z(n1479) );
  XNOR U1602 ( .A(b[7]), .B(a[27]), .Z(n1472) );
  NANDN U1603 ( .A(n1472), .B(n5293), .Z(n1429) );
  NANDN U1604 ( .A(n1427), .B(n5294), .Z(n1428) );
  NAND U1605 ( .A(n1429), .B(n1428), .Z(n1454) );
  XNOR U1606 ( .A(b[3]), .B(a[31]), .Z(n1475) );
  NANDN U1607 ( .A(n1475), .B(n5160), .Z(n1432) );
  NANDN U1608 ( .A(n1430), .B(n5161), .Z(n1431) );
  AND U1609 ( .A(n1432), .B(n1431), .Z(n1455) );
  XNOR U1610 ( .A(n1454), .B(n1455), .Z(n1456) );
  NANDN U1611 ( .A(n292), .B(a[33]), .Z(n1433) );
  XOR U1612 ( .A(n5199), .B(n1433), .Z(n1435) );
  NANDN U1613 ( .A(b[0]), .B(a[32]), .Z(n1434) );
  AND U1614 ( .A(n1435), .B(n1434), .Z(n1462) );
  XNOR U1615 ( .A(b[5]), .B(a[29]), .Z(n1469) );
  NANDN U1616 ( .A(n1469), .B(n5240), .Z(n1438) );
  NANDN U1617 ( .A(n1436), .B(n5241), .Z(n1437) );
  NAND U1618 ( .A(n1438), .B(n1437), .Z(n1460) );
  NANDN U1619 ( .A(n295), .B(a[25]), .Z(n1461) );
  XNOR U1620 ( .A(n1460), .B(n1461), .Z(n1463) );
  XOR U1621 ( .A(n1462), .B(n1463), .Z(n1457) );
  XOR U1622 ( .A(n1456), .B(n1457), .Z(n1478) );
  XOR U1623 ( .A(n1479), .B(n1478), .Z(n1480) );
  XNOR U1624 ( .A(n1481), .B(n1480), .Z(n1450) );
  NAND U1625 ( .A(n1440), .B(n1439), .Z(n1444) );
  NAND U1626 ( .A(n1442), .B(n1441), .Z(n1443) );
  NAND U1627 ( .A(n1444), .B(n1443), .Z(n1451) );
  XNOR U1628 ( .A(n1450), .B(n1451), .Z(n1452) );
  XNOR U1629 ( .A(n1453), .B(n1452), .Z(n1484) );
  XNOR U1630 ( .A(n1484), .B(sreg[153]), .Z(n1486) );
  NAND U1631 ( .A(n1445), .B(sreg[152]), .Z(n1449) );
  OR U1632 ( .A(n1447), .B(n1446), .Z(n1448) );
  AND U1633 ( .A(n1449), .B(n1448), .Z(n1485) );
  XOR U1634 ( .A(n1486), .B(n1485), .Z(c[153]) );
  NANDN U1635 ( .A(n1455), .B(n1454), .Z(n1459) );
  NAND U1636 ( .A(n1457), .B(n1456), .Z(n1458) );
  NAND U1637 ( .A(n1459), .B(n1458), .Z(n1520) );
  NANDN U1638 ( .A(n1461), .B(n1460), .Z(n1465) );
  NAND U1639 ( .A(n1463), .B(n1462), .Z(n1464) );
  NAND U1640 ( .A(n1465), .B(n1464), .Z(n1518) );
  NANDN U1641 ( .A(n292), .B(a[34]), .Z(n1466) );
  XOR U1642 ( .A(n5199), .B(n1466), .Z(n1468) );
  NANDN U1643 ( .A(b[0]), .B(a[33]), .Z(n1467) );
  AND U1644 ( .A(n1468), .B(n1467), .Z(n1501) );
  XNOR U1645 ( .A(b[5]), .B(a[30]), .Z(n1514) );
  NANDN U1646 ( .A(n1514), .B(n5240), .Z(n1471) );
  NANDN U1647 ( .A(n1469), .B(n5241), .Z(n1470) );
  NAND U1648 ( .A(n1471), .B(n1470), .Z(n1499) );
  NANDN U1649 ( .A(n295), .B(a[26]), .Z(n1500) );
  XNOR U1650 ( .A(n1499), .B(n1500), .Z(n1502) );
  XOR U1651 ( .A(n1501), .B(n1502), .Z(n1495) );
  XNOR U1652 ( .A(b[7]), .B(a[28]), .Z(n1505) );
  NANDN U1653 ( .A(n1505), .B(n5293), .Z(n1474) );
  NANDN U1654 ( .A(n1472), .B(n5294), .Z(n1473) );
  NAND U1655 ( .A(n1474), .B(n1473), .Z(n1493) );
  XNOR U1656 ( .A(b[3]), .B(a[32]), .Z(n1508) );
  NANDN U1657 ( .A(n1508), .B(n5160), .Z(n1477) );
  NANDN U1658 ( .A(n1475), .B(n5161), .Z(n1476) );
  AND U1659 ( .A(n1477), .B(n1476), .Z(n1494) );
  XNOR U1660 ( .A(n1493), .B(n1494), .Z(n1496) );
  XOR U1661 ( .A(n1495), .B(n1496), .Z(n1517) );
  XOR U1662 ( .A(n1518), .B(n1517), .Z(n1519) );
  XNOR U1663 ( .A(n1520), .B(n1519), .Z(n1489) );
  NAND U1664 ( .A(n1479), .B(n1478), .Z(n1483) );
  NAND U1665 ( .A(n1481), .B(n1480), .Z(n1482) );
  NAND U1666 ( .A(n1483), .B(n1482), .Z(n1490) );
  XNOR U1667 ( .A(n1489), .B(n1490), .Z(n1491) );
  XNOR U1668 ( .A(n1492), .B(n1491), .Z(n1523) );
  XNOR U1669 ( .A(n1523), .B(sreg[154]), .Z(n1525) );
  NAND U1670 ( .A(n1484), .B(sreg[153]), .Z(n1488) );
  OR U1671 ( .A(n1486), .B(n1485), .Z(n1487) );
  AND U1672 ( .A(n1488), .B(n1487), .Z(n1524) );
  XOR U1673 ( .A(n1525), .B(n1524), .Z(c[154]) );
  NANDN U1674 ( .A(n1494), .B(n1493), .Z(n1498) );
  NAND U1675 ( .A(n1496), .B(n1495), .Z(n1497) );
  NAND U1676 ( .A(n1498), .B(n1497), .Z(n1559) );
  NANDN U1677 ( .A(n1500), .B(n1499), .Z(n1504) );
  NAND U1678 ( .A(n1502), .B(n1501), .Z(n1503) );
  NAND U1679 ( .A(n1504), .B(n1503), .Z(n1557) );
  XNOR U1680 ( .A(b[7]), .B(a[29]), .Z(n1544) );
  NANDN U1681 ( .A(n1544), .B(n5293), .Z(n1507) );
  NANDN U1682 ( .A(n1505), .B(n5294), .Z(n1506) );
  NAND U1683 ( .A(n1507), .B(n1506), .Z(n1532) );
  XNOR U1684 ( .A(b[3]), .B(a[33]), .Z(n1547) );
  NANDN U1685 ( .A(n1547), .B(n5160), .Z(n1510) );
  NANDN U1686 ( .A(n1508), .B(n5161), .Z(n1509) );
  AND U1687 ( .A(n1510), .B(n1509), .Z(n1533) );
  XNOR U1688 ( .A(n1532), .B(n1533), .Z(n1534) );
  NANDN U1689 ( .A(n292), .B(a[35]), .Z(n1511) );
  XOR U1690 ( .A(n5199), .B(n1511), .Z(n1513) );
  NANDN U1691 ( .A(b[0]), .B(a[34]), .Z(n1512) );
  AND U1692 ( .A(n1513), .B(n1512), .Z(n1540) );
  XNOR U1693 ( .A(b[5]), .B(a[31]), .Z(n1553) );
  NANDN U1694 ( .A(n1553), .B(n5240), .Z(n1516) );
  NANDN U1695 ( .A(n1514), .B(n5241), .Z(n1515) );
  NAND U1696 ( .A(n1516), .B(n1515), .Z(n1538) );
  NANDN U1697 ( .A(n295), .B(a[27]), .Z(n1539) );
  XNOR U1698 ( .A(n1538), .B(n1539), .Z(n1541) );
  XOR U1699 ( .A(n1540), .B(n1541), .Z(n1535) );
  XOR U1700 ( .A(n1534), .B(n1535), .Z(n1556) );
  XOR U1701 ( .A(n1557), .B(n1556), .Z(n1558) );
  XNOR U1702 ( .A(n1559), .B(n1558), .Z(n1528) );
  NAND U1703 ( .A(n1518), .B(n1517), .Z(n1522) );
  NAND U1704 ( .A(n1520), .B(n1519), .Z(n1521) );
  NAND U1705 ( .A(n1522), .B(n1521), .Z(n1529) );
  XNOR U1706 ( .A(n1528), .B(n1529), .Z(n1530) );
  XNOR U1707 ( .A(n1531), .B(n1530), .Z(n1562) );
  XNOR U1708 ( .A(n1562), .B(sreg[155]), .Z(n1564) );
  NAND U1709 ( .A(n1523), .B(sreg[154]), .Z(n1527) );
  OR U1710 ( .A(n1525), .B(n1524), .Z(n1526) );
  AND U1711 ( .A(n1527), .B(n1526), .Z(n1563) );
  XOR U1712 ( .A(n1564), .B(n1563), .Z(c[155]) );
  NANDN U1713 ( .A(n1533), .B(n1532), .Z(n1537) );
  NAND U1714 ( .A(n1535), .B(n1534), .Z(n1536) );
  NAND U1715 ( .A(n1537), .B(n1536), .Z(n1598) );
  NANDN U1716 ( .A(n1539), .B(n1538), .Z(n1543) );
  NAND U1717 ( .A(n1541), .B(n1540), .Z(n1542) );
  NAND U1718 ( .A(n1543), .B(n1542), .Z(n1596) );
  XNOR U1719 ( .A(b[7]), .B(a[30]), .Z(n1583) );
  NANDN U1720 ( .A(n1583), .B(n5293), .Z(n1546) );
  NANDN U1721 ( .A(n1544), .B(n5294), .Z(n1545) );
  NAND U1722 ( .A(n1546), .B(n1545), .Z(n1571) );
  XNOR U1723 ( .A(b[3]), .B(a[34]), .Z(n1586) );
  NANDN U1724 ( .A(n1586), .B(n5160), .Z(n1549) );
  NANDN U1725 ( .A(n1547), .B(n5161), .Z(n1548) );
  AND U1726 ( .A(n1549), .B(n1548), .Z(n1572) );
  XNOR U1727 ( .A(n1571), .B(n1572), .Z(n1573) );
  NANDN U1728 ( .A(n292), .B(a[36]), .Z(n1550) );
  XOR U1729 ( .A(n5199), .B(n1550), .Z(n1552) );
  NANDN U1730 ( .A(b[0]), .B(a[35]), .Z(n1551) );
  AND U1731 ( .A(n1552), .B(n1551), .Z(n1579) );
  XNOR U1732 ( .A(b[5]), .B(a[32]), .Z(n1592) );
  NANDN U1733 ( .A(n1592), .B(n5240), .Z(n1555) );
  NANDN U1734 ( .A(n1553), .B(n5241), .Z(n1554) );
  NAND U1735 ( .A(n1555), .B(n1554), .Z(n1577) );
  NANDN U1736 ( .A(n295), .B(a[28]), .Z(n1578) );
  XNOR U1737 ( .A(n1577), .B(n1578), .Z(n1580) );
  XOR U1738 ( .A(n1579), .B(n1580), .Z(n1574) );
  XOR U1739 ( .A(n1573), .B(n1574), .Z(n1595) );
  XOR U1740 ( .A(n1596), .B(n1595), .Z(n1597) );
  XNOR U1741 ( .A(n1598), .B(n1597), .Z(n1567) );
  NAND U1742 ( .A(n1557), .B(n1556), .Z(n1561) );
  NAND U1743 ( .A(n1559), .B(n1558), .Z(n1560) );
  NAND U1744 ( .A(n1561), .B(n1560), .Z(n1568) );
  XNOR U1745 ( .A(n1567), .B(n1568), .Z(n1569) );
  XNOR U1746 ( .A(n1570), .B(n1569), .Z(n1601) );
  XNOR U1747 ( .A(n1601), .B(sreg[156]), .Z(n1603) );
  NAND U1748 ( .A(n1562), .B(sreg[155]), .Z(n1566) );
  OR U1749 ( .A(n1564), .B(n1563), .Z(n1565) );
  AND U1750 ( .A(n1566), .B(n1565), .Z(n1602) );
  XOR U1751 ( .A(n1603), .B(n1602), .Z(c[156]) );
  NANDN U1752 ( .A(n1572), .B(n1571), .Z(n1576) );
  NAND U1753 ( .A(n1574), .B(n1573), .Z(n1575) );
  NAND U1754 ( .A(n1576), .B(n1575), .Z(n1637) );
  NANDN U1755 ( .A(n1578), .B(n1577), .Z(n1582) );
  NAND U1756 ( .A(n1580), .B(n1579), .Z(n1581) );
  NAND U1757 ( .A(n1582), .B(n1581), .Z(n1635) );
  XNOR U1758 ( .A(b[7]), .B(a[31]), .Z(n1622) );
  NANDN U1759 ( .A(n1622), .B(n5293), .Z(n1585) );
  NANDN U1760 ( .A(n1583), .B(n5294), .Z(n1584) );
  NAND U1761 ( .A(n1585), .B(n1584), .Z(n1610) );
  XNOR U1762 ( .A(b[3]), .B(a[35]), .Z(n1625) );
  NANDN U1763 ( .A(n1625), .B(n5160), .Z(n1588) );
  NANDN U1764 ( .A(n1586), .B(n5161), .Z(n1587) );
  AND U1765 ( .A(n1588), .B(n1587), .Z(n1611) );
  XNOR U1766 ( .A(n1610), .B(n1611), .Z(n1612) );
  NANDN U1767 ( .A(n292), .B(a[37]), .Z(n1589) );
  XOR U1768 ( .A(n5199), .B(n1589), .Z(n1591) );
  NANDN U1769 ( .A(b[0]), .B(a[36]), .Z(n1590) );
  AND U1770 ( .A(n1591), .B(n1590), .Z(n1618) );
  XNOR U1771 ( .A(b[5]), .B(a[33]), .Z(n1631) );
  NANDN U1772 ( .A(n1631), .B(n5240), .Z(n1594) );
  NANDN U1773 ( .A(n1592), .B(n5241), .Z(n1593) );
  NAND U1774 ( .A(n1594), .B(n1593), .Z(n1616) );
  NANDN U1775 ( .A(n295), .B(a[29]), .Z(n1617) );
  XNOR U1776 ( .A(n1616), .B(n1617), .Z(n1619) );
  XOR U1777 ( .A(n1618), .B(n1619), .Z(n1613) );
  XOR U1778 ( .A(n1612), .B(n1613), .Z(n1634) );
  XOR U1779 ( .A(n1635), .B(n1634), .Z(n1636) );
  XNOR U1780 ( .A(n1637), .B(n1636), .Z(n1606) );
  NAND U1781 ( .A(n1596), .B(n1595), .Z(n1600) );
  NAND U1782 ( .A(n1598), .B(n1597), .Z(n1599) );
  NAND U1783 ( .A(n1600), .B(n1599), .Z(n1607) );
  XNOR U1784 ( .A(n1606), .B(n1607), .Z(n1608) );
  XNOR U1785 ( .A(n1609), .B(n1608), .Z(n1640) );
  XNOR U1786 ( .A(n1640), .B(sreg[157]), .Z(n1642) );
  NAND U1787 ( .A(n1601), .B(sreg[156]), .Z(n1605) );
  OR U1788 ( .A(n1603), .B(n1602), .Z(n1604) );
  AND U1789 ( .A(n1605), .B(n1604), .Z(n1641) );
  XOR U1790 ( .A(n1642), .B(n1641), .Z(c[157]) );
  NANDN U1791 ( .A(n1611), .B(n1610), .Z(n1615) );
  NAND U1792 ( .A(n1613), .B(n1612), .Z(n1614) );
  NAND U1793 ( .A(n1615), .B(n1614), .Z(n1676) );
  NANDN U1794 ( .A(n1617), .B(n1616), .Z(n1621) );
  NAND U1795 ( .A(n1619), .B(n1618), .Z(n1620) );
  NAND U1796 ( .A(n1621), .B(n1620), .Z(n1674) );
  XNOR U1797 ( .A(b[7]), .B(a[32]), .Z(n1661) );
  NANDN U1798 ( .A(n1661), .B(n5293), .Z(n1624) );
  NANDN U1799 ( .A(n1622), .B(n5294), .Z(n1623) );
  NAND U1800 ( .A(n1624), .B(n1623), .Z(n1649) );
  XNOR U1801 ( .A(b[3]), .B(a[36]), .Z(n1664) );
  NANDN U1802 ( .A(n1664), .B(n5160), .Z(n1627) );
  NANDN U1803 ( .A(n1625), .B(n5161), .Z(n1626) );
  AND U1804 ( .A(n1627), .B(n1626), .Z(n1650) );
  XNOR U1805 ( .A(n1649), .B(n1650), .Z(n1651) );
  NANDN U1806 ( .A(n292), .B(a[38]), .Z(n1628) );
  XOR U1807 ( .A(n5199), .B(n1628), .Z(n1630) );
  NANDN U1808 ( .A(b[0]), .B(a[37]), .Z(n1629) );
  AND U1809 ( .A(n1630), .B(n1629), .Z(n1657) );
  XNOR U1810 ( .A(b[5]), .B(a[34]), .Z(n1670) );
  NANDN U1811 ( .A(n1670), .B(n5240), .Z(n1633) );
  NANDN U1812 ( .A(n1631), .B(n5241), .Z(n1632) );
  NAND U1813 ( .A(n1633), .B(n1632), .Z(n1655) );
  NANDN U1814 ( .A(n295), .B(a[30]), .Z(n1656) );
  XNOR U1815 ( .A(n1655), .B(n1656), .Z(n1658) );
  XOR U1816 ( .A(n1657), .B(n1658), .Z(n1652) );
  XOR U1817 ( .A(n1651), .B(n1652), .Z(n1673) );
  XOR U1818 ( .A(n1674), .B(n1673), .Z(n1675) );
  XNOR U1819 ( .A(n1676), .B(n1675), .Z(n1645) );
  NAND U1820 ( .A(n1635), .B(n1634), .Z(n1639) );
  NAND U1821 ( .A(n1637), .B(n1636), .Z(n1638) );
  NAND U1822 ( .A(n1639), .B(n1638), .Z(n1646) );
  XNOR U1823 ( .A(n1645), .B(n1646), .Z(n1647) );
  XNOR U1824 ( .A(n1648), .B(n1647), .Z(n1679) );
  XNOR U1825 ( .A(n1679), .B(sreg[158]), .Z(n1681) );
  NAND U1826 ( .A(n1640), .B(sreg[157]), .Z(n1644) );
  OR U1827 ( .A(n1642), .B(n1641), .Z(n1643) );
  AND U1828 ( .A(n1644), .B(n1643), .Z(n1680) );
  XOR U1829 ( .A(n1681), .B(n1680), .Z(c[158]) );
  NANDN U1830 ( .A(n1650), .B(n1649), .Z(n1654) );
  NAND U1831 ( .A(n1652), .B(n1651), .Z(n1653) );
  NAND U1832 ( .A(n1654), .B(n1653), .Z(n1715) );
  NANDN U1833 ( .A(n1656), .B(n1655), .Z(n1660) );
  NAND U1834 ( .A(n1658), .B(n1657), .Z(n1659) );
  NAND U1835 ( .A(n1660), .B(n1659), .Z(n1713) );
  XNOR U1836 ( .A(b[7]), .B(a[33]), .Z(n1700) );
  NANDN U1837 ( .A(n1700), .B(n5293), .Z(n1663) );
  NANDN U1838 ( .A(n1661), .B(n5294), .Z(n1662) );
  NAND U1839 ( .A(n1663), .B(n1662), .Z(n1688) );
  XNOR U1840 ( .A(b[3]), .B(a[37]), .Z(n1703) );
  NANDN U1841 ( .A(n1703), .B(n5160), .Z(n1666) );
  NANDN U1842 ( .A(n1664), .B(n5161), .Z(n1665) );
  AND U1843 ( .A(n1666), .B(n1665), .Z(n1689) );
  XNOR U1844 ( .A(n1688), .B(n1689), .Z(n1690) );
  NANDN U1845 ( .A(n292), .B(a[39]), .Z(n1667) );
  XOR U1846 ( .A(n5199), .B(n1667), .Z(n1669) );
  NANDN U1847 ( .A(b[0]), .B(a[38]), .Z(n1668) );
  AND U1848 ( .A(n1669), .B(n1668), .Z(n1696) );
  XNOR U1849 ( .A(b[5]), .B(a[35]), .Z(n1709) );
  NANDN U1850 ( .A(n1709), .B(n5240), .Z(n1672) );
  NANDN U1851 ( .A(n1670), .B(n5241), .Z(n1671) );
  NAND U1852 ( .A(n1672), .B(n1671), .Z(n1694) );
  NANDN U1853 ( .A(n295), .B(a[31]), .Z(n1695) );
  XNOR U1854 ( .A(n1694), .B(n1695), .Z(n1697) );
  XOR U1855 ( .A(n1696), .B(n1697), .Z(n1691) );
  XOR U1856 ( .A(n1690), .B(n1691), .Z(n1712) );
  XOR U1857 ( .A(n1713), .B(n1712), .Z(n1714) );
  XNOR U1858 ( .A(n1715), .B(n1714), .Z(n1684) );
  NAND U1859 ( .A(n1674), .B(n1673), .Z(n1678) );
  NAND U1860 ( .A(n1676), .B(n1675), .Z(n1677) );
  NAND U1861 ( .A(n1678), .B(n1677), .Z(n1685) );
  XNOR U1862 ( .A(n1684), .B(n1685), .Z(n1686) );
  XNOR U1863 ( .A(n1687), .B(n1686), .Z(n1718) );
  XNOR U1864 ( .A(n1718), .B(sreg[159]), .Z(n1720) );
  NAND U1865 ( .A(n1679), .B(sreg[158]), .Z(n1683) );
  OR U1866 ( .A(n1681), .B(n1680), .Z(n1682) );
  AND U1867 ( .A(n1683), .B(n1682), .Z(n1719) );
  XOR U1868 ( .A(n1720), .B(n1719), .Z(c[159]) );
  NANDN U1869 ( .A(n1689), .B(n1688), .Z(n1693) );
  NAND U1870 ( .A(n1691), .B(n1690), .Z(n1692) );
  NAND U1871 ( .A(n1693), .B(n1692), .Z(n1754) );
  NANDN U1872 ( .A(n1695), .B(n1694), .Z(n1699) );
  NAND U1873 ( .A(n1697), .B(n1696), .Z(n1698) );
  NAND U1874 ( .A(n1699), .B(n1698), .Z(n1752) );
  XNOR U1875 ( .A(b[7]), .B(a[34]), .Z(n1739) );
  NANDN U1876 ( .A(n1739), .B(n5293), .Z(n1702) );
  NANDN U1877 ( .A(n1700), .B(n5294), .Z(n1701) );
  NAND U1878 ( .A(n1702), .B(n1701), .Z(n1727) );
  XNOR U1879 ( .A(b[3]), .B(a[38]), .Z(n1742) );
  NANDN U1880 ( .A(n1742), .B(n5160), .Z(n1705) );
  NANDN U1881 ( .A(n1703), .B(n5161), .Z(n1704) );
  AND U1882 ( .A(n1705), .B(n1704), .Z(n1728) );
  XNOR U1883 ( .A(n1727), .B(n1728), .Z(n1729) );
  NANDN U1884 ( .A(n292), .B(a[40]), .Z(n1706) );
  XOR U1885 ( .A(n5199), .B(n1706), .Z(n1708) );
  NANDN U1886 ( .A(b[0]), .B(a[39]), .Z(n1707) );
  AND U1887 ( .A(n1708), .B(n1707), .Z(n1735) );
  XNOR U1888 ( .A(b[5]), .B(a[36]), .Z(n1748) );
  NANDN U1889 ( .A(n1748), .B(n5240), .Z(n1711) );
  NANDN U1890 ( .A(n1709), .B(n5241), .Z(n1710) );
  NAND U1891 ( .A(n1711), .B(n1710), .Z(n1733) );
  NANDN U1892 ( .A(n295), .B(a[32]), .Z(n1734) );
  XNOR U1893 ( .A(n1733), .B(n1734), .Z(n1736) );
  XOR U1894 ( .A(n1735), .B(n1736), .Z(n1730) );
  XOR U1895 ( .A(n1729), .B(n1730), .Z(n1751) );
  XOR U1896 ( .A(n1752), .B(n1751), .Z(n1753) );
  XNOR U1897 ( .A(n1754), .B(n1753), .Z(n1723) );
  NAND U1898 ( .A(n1713), .B(n1712), .Z(n1717) );
  NAND U1899 ( .A(n1715), .B(n1714), .Z(n1716) );
  NAND U1900 ( .A(n1717), .B(n1716), .Z(n1724) );
  XNOR U1901 ( .A(n1723), .B(n1724), .Z(n1725) );
  XNOR U1902 ( .A(n1726), .B(n1725), .Z(n1757) );
  XNOR U1903 ( .A(n1757), .B(sreg[160]), .Z(n1759) );
  NAND U1904 ( .A(n1718), .B(sreg[159]), .Z(n1722) );
  OR U1905 ( .A(n1720), .B(n1719), .Z(n1721) );
  AND U1906 ( .A(n1722), .B(n1721), .Z(n1758) );
  XOR U1907 ( .A(n1759), .B(n1758), .Z(c[160]) );
  NANDN U1908 ( .A(n1728), .B(n1727), .Z(n1732) );
  NAND U1909 ( .A(n1730), .B(n1729), .Z(n1731) );
  NAND U1910 ( .A(n1732), .B(n1731), .Z(n1793) );
  NANDN U1911 ( .A(n1734), .B(n1733), .Z(n1738) );
  NAND U1912 ( .A(n1736), .B(n1735), .Z(n1737) );
  NAND U1913 ( .A(n1738), .B(n1737), .Z(n1791) );
  XNOR U1914 ( .A(b[7]), .B(a[35]), .Z(n1784) );
  NANDN U1915 ( .A(n1784), .B(n5293), .Z(n1741) );
  NANDN U1916 ( .A(n1739), .B(n5294), .Z(n1740) );
  NAND U1917 ( .A(n1741), .B(n1740), .Z(n1766) );
  XNOR U1918 ( .A(b[3]), .B(a[39]), .Z(n1787) );
  NANDN U1919 ( .A(n1787), .B(n5160), .Z(n1744) );
  NANDN U1920 ( .A(n1742), .B(n5161), .Z(n1743) );
  AND U1921 ( .A(n1744), .B(n1743), .Z(n1767) );
  XNOR U1922 ( .A(n1766), .B(n1767), .Z(n1768) );
  NANDN U1923 ( .A(n292), .B(a[41]), .Z(n1745) );
  XOR U1924 ( .A(n5199), .B(n1745), .Z(n1747) );
  NANDN U1925 ( .A(b[0]), .B(a[40]), .Z(n1746) );
  AND U1926 ( .A(n1747), .B(n1746), .Z(n1774) );
  XNOR U1927 ( .A(n294), .B(a[37]), .Z(n1778) );
  NAND U1928 ( .A(n1778), .B(n5240), .Z(n1750) );
  NANDN U1929 ( .A(n1748), .B(n5241), .Z(n1749) );
  NAND U1930 ( .A(n1750), .B(n1749), .Z(n1772) );
  NANDN U1931 ( .A(n295), .B(a[33]), .Z(n1773) );
  XNOR U1932 ( .A(n1772), .B(n1773), .Z(n1775) );
  XOR U1933 ( .A(n1774), .B(n1775), .Z(n1769) );
  XOR U1934 ( .A(n1768), .B(n1769), .Z(n1790) );
  XOR U1935 ( .A(n1791), .B(n1790), .Z(n1792) );
  XNOR U1936 ( .A(n1793), .B(n1792), .Z(n1762) );
  NAND U1937 ( .A(n1752), .B(n1751), .Z(n1756) );
  NAND U1938 ( .A(n1754), .B(n1753), .Z(n1755) );
  NAND U1939 ( .A(n1756), .B(n1755), .Z(n1763) );
  XNOR U1940 ( .A(n1762), .B(n1763), .Z(n1764) );
  XNOR U1941 ( .A(n1765), .B(n1764), .Z(n1796) );
  XNOR U1942 ( .A(n1796), .B(sreg[161]), .Z(n1798) );
  NAND U1943 ( .A(n1757), .B(sreg[160]), .Z(n1761) );
  OR U1944 ( .A(n1759), .B(n1758), .Z(n1760) );
  AND U1945 ( .A(n1761), .B(n1760), .Z(n1797) );
  XOR U1946 ( .A(n1798), .B(n1797), .Z(c[161]) );
  NANDN U1947 ( .A(n1767), .B(n1766), .Z(n1771) );
  NAND U1948 ( .A(n1769), .B(n1768), .Z(n1770) );
  NAND U1949 ( .A(n1771), .B(n1770), .Z(n1832) );
  NANDN U1950 ( .A(n1773), .B(n1772), .Z(n1777) );
  NAND U1951 ( .A(n1775), .B(n1774), .Z(n1776) );
  NAND U1952 ( .A(n1777), .B(n1776), .Z(n1830) );
  XNOR U1953 ( .A(b[5]), .B(a[38]), .Z(n1814) );
  NANDN U1954 ( .A(n1814), .B(n5240), .Z(n1780) );
  NAND U1955 ( .A(n5241), .B(n1778), .Z(n1779) );
  AND U1956 ( .A(n1780), .B(n1779), .Z(n1823) );
  NANDN U1957 ( .A(n295), .B(a[34]), .Z(n1824) );
  XOR U1958 ( .A(n1823), .B(n1824), .Z(n1826) );
  NANDN U1959 ( .A(n292), .B(a[42]), .Z(n1781) );
  XOR U1960 ( .A(n5199), .B(n1781), .Z(n1783) );
  NANDN U1961 ( .A(b[0]), .B(a[41]), .Z(n1782) );
  AND U1962 ( .A(n1783), .B(n1782), .Z(n1825) );
  XNOR U1963 ( .A(n1826), .B(n1825), .Z(n1820) );
  XNOR U1964 ( .A(b[7]), .B(a[36]), .Z(n1805) );
  NANDN U1965 ( .A(n1805), .B(n5293), .Z(n1786) );
  NANDN U1966 ( .A(n1784), .B(n5294), .Z(n1785) );
  NAND U1967 ( .A(n1786), .B(n1785), .Z(n1817) );
  XNOR U1968 ( .A(b[3]), .B(a[40]), .Z(n1808) );
  NANDN U1969 ( .A(n1808), .B(n5160), .Z(n1789) );
  NANDN U1970 ( .A(n1787), .B(n5161), .Z(n1788) );
  AND U1971 ( .A(n1789), .B(n1788), .Z(n1818) );
  XNOR U1972 ( .A(n1817), .B(n1818), .Z(n1819) );
  XNOR U1973 ( .A(n1820), .B(n1819), .Z(n1829) );
  XOR U1974 ( .A(n1830), .B(n1829), .Z(n1831) );
  XNOR U1975 ( .A(n1832), .B(n1831), .Z(n1801) );
  NAND U1976 ( .A(n1791), .B(n1790), .Z(n1795) );
  NAND U1977 ( .A(n1793), .B(n1792), .Z(n1794) );
  NAND U1978 ( .A(n1795), .B(n1794), .Z(n1802) );
  XNOR U1979 ( .A(n1801), .B(n1802), .Z(n1803) );
  XNOR U1980 ( .A(n1804), .B(n1803), .Z(n1833) );
  XNOR U1981 ( .A(n1833), .B(sreg[162]), .Z(n1835) );
  NAND U1982 ( .A(n1796), .B(sreg[161]), .Z(n1800) );
  OR U1983 ( .A(n1798), .B(n1797), .Z(n1799) );
  AND U1984 ( .A(n1800), .B(n1799), .Z(n1834) );
  XOR U1985 ( .A(n1835), .B(n1834), .Z(c[162]) );
  XNOR U1986 ( .A(b[7]), .B(a[37]), .Z(n1854) );
  NANDN U1987 ( .A(n1854), .B(n5293), .Z(n1807) );
  NANDN U1988 ( .A(n1805), .B(n5294), .Z(n1806) );
  NAND U1989 ( .A(n1807), .B(n1806), .Z(n1842) );
  XNOR U1990 ( .A(b[3]), .B(a[41]), .Z(n1857) );
  NANDN U1991 ( .A(n1857), .B(n5160), .Z(n1810) );
  NANDN U1992 ( .A(n1808), .B(n5161), .Z(n1809) );
  AND U1993 ( .A(n1810), .B(n1809), .Z(n1843) );
  XNOR U1994 ( .A(n1842), .B(n1843), .Z(n1844) );
  NANDN U1995 ( .A(n292), .B(a[43]), .Z(n1811) );
  XOR U1996 ( .A(n5199), .B(n1811), .Z(n1813) );
  NANDN U1997 ( .A(b[0]), .B(a[42]), .Z(n1812) );
  AND U1998 ( .A(n1813), .B(n1812), .Z(n1850) );
  XNOR U1999 ( .A(b[5]), .B(a[39]), .Z(n1863) );
  NANDN U2000 ( .A(n1863), .B(n5240), .Z(n1816) );
  NANDN U2001 ( .A(n1814), .B(n5241), .Z(n1815) );
  NAND U2002 ( .A(n1816), .B(n1815), .Z(n1848) );
  NANDN U2003 ( .A(n295), .B(a[35]), .Z(n1849) );
  XNOR U2004 ( .A(n1848), .B(n1849), .Z(n1851) );
  XOR U2005 ( .A(n1850), .B(n1851), .Z(n1845) );
  XOR U2006 ( .A(n1844), .B(n1845), .Z(n1868) );
  NANDN U2007 ( .A(n1818), .B(n1817), .Z(n1822) );
  NANDN U2008 ( .A(n1820), .B(n1819), .Z(n1821) );
  NAND U2009 ( .A(n1822), .B(n1821), .Z(n1866) );
  OR U2010 ( .A(n1824), .B(n1823), .Z(n1828) );
  NAND U2011 ( .A(n1826), .B(n1825), .Z(n1827) );
  AND U2012 ( .A(n1828), .B(n1827), .Z(n1867) );
  XNOR U2013 ( .A(n1866), .B(n1867), .Z(n1869) );
  XNOR U2014 ( .A(n1868), .B(n1869), .Z(n1838) );
  XNOR U2015 ( .A(n1838), .B(n1839), .Z(n1840) );
  XNOR U2016 ( .A(n1841), .B(n1840), .Z(n1872) );
  XNOR U2017 ( .A(n1872), .B(sreg[163]), .Z(n1874) );
  NAND U2018 ( .A(n1833), .B(sreg[162]), .Z(n1837) );
  OR U2019 ( .A(n1835), .B(n1834), .Z(n1836) );
  AND U2020 ( .A(n1837), .B(n1836), .Z(n1873) );
  XOR U2021 ( .A(n1874), .B(n1873), .Z(c[163]) );
  NANDN U2022 ( .A(n1843), .B(n1842), .Z(n1847) );
  NAND U2023 ( .A(n1845), .B(n1844), .Z(n1846) );
  NAND U2024 ( .A(n1847), .B(n1846), .Z(n1908) );
  NANDN U2025 ( .A(n1849), .B(n1848), .Z(n1853) );
  NAND U2026 ( .A(n1851), .B(n1850), .Z(n1852) );
  NAND U2027 ( .A(n1853), .B(n1852), .Z(n1906) );
  XNOR U2028 ( .A(b[7]), .B(a[38]), .Z(n1893) );
  NANDN U2029 ( .A(n1893), .B(n5293), .Z(n1856) );
  NANDN U2030 ( .A(n1854), .B(n5294), .Z(n1855) );
  NAND U2031 ( .A(n1856), .B(n1855), .Z(n1881) );
  XNOR U2032 ( .A(b[3]), .B(a[42]), .Z(n1896) );
  NANDN U2033 ( .A(n1896), .B(n5160), .Z(n1859) );
  NANDN U2034 ( .A(n1857), .B(n5161), .Z(n1858) );
  AND U2035 ( .A(n1859), .B(n1858), .Z(n1882) );
  XNOR U2036 ( .A(n1881), .B(n1882), .Z(n1883) );
  NANDN U2037 ( .A(n292), .B(a[44]), .Z(n1860) );
  XOR U2038 ( .A(n5199), .B(n1860), .Z(n1862) );
  NANDN U2039 ( .A(b[0]), .B(a[43]), .Z(n1861) );
  AND U2040 ( .A(n1862), .B(n1861), .Z(n1889) );
  XNOR U2041 ( .A(b[5]), .B(a[40]), .Z(n1902) );
  NANDN U2042 ( .A(n1902), .B(n5240), .Z(n1865) );
  NANDN U2043 ( .A(n1863), .B(n5241), .Z(n1864) );
  NAND U2044 ( .A(n1865), .B(n1864), .Z(n1887) );
  NANDN U2045 ( .A(n295), .B(a[36]), .Z(n1888) );
  XNOR U2046 ( .A(n1887), .B(n1888), .Z(n1890) );
  XOR U2047 ( .A(n1889), .B(n1890), .Z(n1884) );
  XOR U2048 ( .A(n1883), .B(n1884), .Z(n1905) );
  XOR U2049 ( .A(n1906), .B(n1905), .Z(n1907) );
  XNOR U2050 ( .A(n1908), .B(n1907), .Z(n1877) );
  NANDN U2051 ( .A(n1867), .B(n1866), .Z(n1871) );
  NAND U2052 ( .A(n1869), .B(n1868), .Z(n1870) );
  NAND U2053 ( .A(n1871), .B(n1870), .Z(n1878) );
  XNOR U2054 ( .A(n1877), .B(n1878), .Z(n1879) );
  XNOR U2055 ( .A(n1880), .B(n1879), .Z(n1911) );
  XNOR U2056 ( .A(n1911), .B(sreg[164]), .Z(n1913) );
  NAND U2057 ( .A(n1872), .B(sreg[163]), .Z(n1876) );
  OR U2058 ( .A(n1874), .B(n1873), .Z(n1875) );
  AND U2059 ( .A(n1876), .B(n1875), .Z(n1912) );
  XOR U2060 ( .A(n1913), .B(n1912), .Z(c[164]) );
  NANDN U2061 ( .A(n1882), .B(n1881), .Z(n1886) );
  NAND U2062 ( .A(n1884), .B(n1883), .Z(n1885) );
  NAND U2063 ( .A(n1886), .B(n1885), .Z(n1947) );
  NANDN U2064 ( .A(n1888), .B(n1887), .Z(n1892) );
  NAND U2065 ( .A(n1890), .B(n1889), .Z(n1891) );
  NAND U2066 ( .A(n1892), .B(n1891), .Z(n1945) );
  XNOR U2067 ( .A(b[7]), .B(a[39]), .Z(n1932) );
  NANDN U2068 ( .A(n1932), .B(n5293), .Z(n1895) );
  NANDN U2069 ( .A(n1893), .B(n5294), .Z(n1894) );
  NAND U2070 ( .A(n1895), .B(n1894), .Z(n1920) );
  XNOR U2071 ( .A(b[3]), .B(a[43]), .Z(n1935) );
  NANDN U2072 ( .A(n1935), .B(n5160), .Z(n1898) );
  NANDN U2073 ( .A(n1896), .B(n5161), .Z(n1897) );
  AND U2074 ( .A(n1898), .B(n1897), .Z(n1921) );
  XNOR U2075 ( .A(n1920), .B(n1921), .Z(n1922) );
  NANDN U2076 ( .A(n292), .B(a[45]), .Z(n1899) );
  XOR U2077 ( .A(n5199), .B(n1899), .Z(n1901) );
  NANDN U2078 ( .A(b[0]), .B(a[44]), .Z(n1900) );
  AND U2079 ( .A(n1901), .B(n1900), .Z(n1928) );
  XNOR U2080 ( .A(b[5]), .B(a[41]), .Z(n1941) );
  NANDN U2081 ( .A(n1941), .B(n5240), .Z(n1904) );
  NANDN U2082 ( .A(n1902), .B(n5241), .Z(n1903) );
  NAND U2083 ( .A(n1904), .B(n1903), .Z(n1926) );
  NANDN U2084 ( .A(n295), .B(a[37]), .Z(n1927) );
  XNOR U2085 ( .A(n1926), .B(n1927), .Z(n1929) );
  XOR U2086 ( .A(n1928), .B(n1929), .Z(n1923) );
  XOR U2087 ( .A(n1922), .B(n1923), .Z(n1944) );
  XOR U2088 ( .A(n1945), .B(n1944), .Z(n1946) );
  XNOR U2089 ( .A(n1947), .B(n1946), .Z(n1916) );
  NAND U2090 ( .A(n1906), .B(n1905), .Z(n1910) );
  NAND U2091 ( .A(n1908), .B(n1907), .Z(n1909) );
  NAND U2092 ( .A(n1910), .B(n1909), .Z(n1917) );
  XNOR U2093 ( .A(n1916), .B(n1917), .Z(n1918) );
  XNOR U2094 ( .A(n1919), .B(n1918), .Z(n1950) );
  XNOR U2095 ( .A(n1950), .B(sreg[165]), .Z(n1952) );
  NAND U2096 ( .A(n1911), .B(sreg[164]), .Z(n1915) );
  OR U2097 ( .A(n1913), .B(n1912), .Z(n1914) );
  AND U2098 ( .A(n1915), .B(n1914), .Z(n1951) );
  XOR U2099 ( .A(n1952), .B(n1951), .Z(c[165]) );
  NANDN U2100 ( .A(n1921), .B(n1920), .Z(n1925) );
  NAND U2101 ( .A(n1923), .B(n1922), .Z(n1924) );
  NAND U2102 ( .A(n1925), .B(n1924), .Z(n1986) );
  NANDN U2103 ( .A(n1927), .B(n1926), .Z(n1931) );
  NAND U2104 ( .A(n1929), .B(n1928), .Z(n1930) );
  NAND U2105 ( .A(n1931), .B(n1930), .Z(n1984) );
  XNOR U2106 ( .A(b[7]), .B(a[40]), .Z(n1965) );
  NANDN U2107 ( .A(n1965), .B(n5293), .Z(n1934) );
  NANDN U2108 ( .A(n1932), .B(n5294), .Z(n1933) );
  NAND U2109 ( .A(n1934), .B(n1933), .Z(n1977) );
  XNOR U2110 ( .A(b[3]), .B(a[44]), .Z(n1968) );
  NANDN U2111 ( .A(n1968), .B(n5160), .Z(n1937) );
  NANDN U2112 ( .A(n1935), .B(n5161), .Z(n1936) );
  AND U2113 ( .A(n1937), .B(n1936), .Z(n1978) );
  XNOR U2114 ( .A(n1977), .B(n1978), .Z(n1979) );
  NANDN U2115 ( .A(n292), .B(a[46]), .Z(n1938) );
  XOR U2116 ( .A(n5199), .B(n1938), .Z(n1940) );
  NANDN U2117 ( .A(b[0]), .B(a[45]), .Z(n1939) );
  AND U2118 ( .A(n1940), .B(n1939), .Z(n1973) );
  XNOR U2119 ( .A(n294), .B(a[42]), .Z(n1959) );
  NAND U2120 ( .A(n1959), .B(n5240), .Z(n1943) );
  NANDN U2121 ( .A(n1941), .B(n5241), .Z(n1942) );
  NAND U2122 ( .A(n1943), .B(n1942), .Z(n1971) );
  NANDN U2123 ( .A(n295), .B(a[38]), .Z(n1972) );
  XNOR U2124 ( .A(n1971), .B(n1972), .Z(n1974) );
  XOR U2125 ( .A(n1973), .B(n1974), .Z(n1980) );
  XOR U2126 ( .A(n1979), .B(n1980), .Z(n1983) );
  XOR U2127 ( .A(n1984), .B(n1983), .Z(n1985) );
  XNOR U2128 ( .A(n1986), .B(n1985), .Z(n1955) );
  NAND U2129 ( .A(n1945), .B(n1944), .Z(n1949) );
  NAND U2130 ( .A(n1947), .B(n1946), .Z(n1948) );
  NAND U2131 ( .A(n1949), .B(n1948), .Z(n1956) );
  XNOR U2132 ( .A(n1955), .B(n1956), .Z(n1957) );
  XNOR U2133 ( .A(n1958), .B(n1957), .Z(n1989) );
  XNOR U2134 ( .A(n1989), .B(sreg[166]), .Z(n1991) );
  NAND U2135 ( .A(n1950), .B(sreg[165]), .Z(n1954) );
  OR U2136 ( .A(n1952), .B(n1951), .Z(n1953) );
  AND U2137 ( .A(n1954), .B(n1953), .Z(n1990) );
  XOR U2138 ( .A(n1991), .B(n1990), .Z(c[166]) );
  XNOR U2139 ( .A(b[5]), .B(a[43]), .Z(n2009) );
  NANDN U2140 ( .A(n2009), .B(n5240), .Z(n1961) );
  NAND U2141 ( .A(n5241), .B(n1959), .Z(n1960) );
  AND U2142 ( .A(n1961), .B(n1960), .Z(n2018) );
  NANDN U2143 ( .A(n295), .B(a[39]), .Z(n2019) );
  XOR U2144 ( .A(n2018), .B(n2019), .Z(n2021) );
  NANDN U2145 ( .A(n292), .B(a[47]), .Z(n1962) );
  XOR U2146 ( .A(n5199), .B(n1962), .Z(n1964) );
  NANDN U2147 ( .A(b[0]), .B(a[46]), .Z(n1963) );
  AND U2148 ( .A(n1964), .B(n1963), .Z(n2020) );
  XNOR U2149 ( .A(n2021), .B(n2020), .Z(n2015) );
  XNOR U2150 ( .A(b[7]), .B(a[41]), .Z(n2000) );
  NANDN U2151 ( .A(n2000), .B(n5293), .Z(n1967) );
  NANDN U2152 ( .A(n1965), .B(n5294), .Z(n1966) );
  NAND U2153 ( .A(n1967), .B(n1966), .Z(n2012) );
  XNOR U2154 ( .A(b[3]), .B(a[45]), .Z(n2003) );
  NANDN U2155 ( .A(n2003), .B(n5160), .Z(n1970) );
  NANDN U2156 ( .A(n1968), .B(n5161), .Z(n1969) );
  AND U2157 ( .A(n1970), .B(n1969), .Z(n2013) );
  XNOR U2158 ( .A(n2012), .B(n2013), .Z(n2014) );
  XNOR U2159 ( .A(n2015), .B(n2014), .Z(n2026) );
  NANDN U2160 ( .A(n1972), .B(n1971), .Z(n1976) );
  NAND U2161 ( .A(n1974), .B(n1973), .Z(n1975) );
  NAND U2162 ( .A(n1976), .B(n1975), .Z(n2024) );
  NANDN U2163 ( .A(n1978), .B(n1977), .Z(n1982) );
  NAND U2164 ( .A(n1980), .B(n1979), .Z(n1981) );
  AND U2165 ( .A(n1982), .B(n1981), .Z(n2025) );
  XNOR U2166 ( .A(n2024), .B(n2025), .Z(n2027) );
  XOR U2167 ( .A(n2026), .B(n2027), .Z(n1994) );
  NAND U2168 ( .A(n1984), .B(n1983), .Z(n1988) );
  NAND U2169 ( .A(n1986), .B(n1985), .Z(n1987) );
  NAND U2170 ( .A(n1988), .B(n1987), .Z(n1995) );
  XOR U2171 ( .A(n1994), .B(n1995), .Z(n1996) );
  XNOR U2172 ( .A(n1997), .B(n1996), .Z(n2028) );
  XNOR U2173 ( .A(n2028), .B(sreg[167]), .Z(n2030) );
  NAND U2174 ( .A(n1989), .B(sreg[166]), .Z(n1993) );
  OR U2175 ( .A(n1991), .B(n1990), .Z(n1992) );
  AND U2176 ( .A(n1993), .B(n1992), .Z(n2029) );
  XOR U2177 ( .A(n2030), .B(n2029), .Z(c[167]) );
  OR U2178 ( .A(n1995), .B(n1994), .Z(n1999) );
  NAND U2179 ( .A(n1997), .B(n1996), .Z(n1998) );
  NAND U2180 ( .A(n1999), .B(n1998), .Z(n2036) );
  XNOR U2181 ( .A(b[7]), .B(a[42]), .Z(n2049) );
  NANDN U2182 ( .A(n2049), .B(n5293), .Z(n2002) );
  NANDN U2183 ( .A(n2000), .B(n5294), .Z(n2001) );
  NAND U2184 ( .A(n2002), .B(n2001), .Z(n2037) );
  XNOR U2185 ( .A(b[3]), .B(a[46]), .Z(n2052) );
  NANDN U2186 ( .A(n2052), .B(n5160), .Z(n2005) );
  NANDN U2187 ( .A(n2003), .B(n5161), .Z(n2004) );
  AND U2188 ( .A(n2005), .B(n2004), .Z(n2038) );
  XNOR U2189 ( .A(n2037), .B(n2038), .Z(n2039) );
  NANDN U2190 ( .A(n292), .B(a[48]), .Z(n2006) );
  XOR U2191 ( .A(n5199), .B(n2006), .Z(n2008) );
  NANDN U2192 ( .A(b[0]), .B(a[47]), .Z(n2007) );
  AND U2193 ( .A(n2008), .B(n2007), .Z(n2045) );
  XNOR U2194 ( .A(b[5]), .B(a[44]), .Z(n2058) );
  NANDN U2195 ( .A(n2058), .B(n5240), .Z(n2011) );
  NANDN U2196 ( .A(n2009), .B(n5241), .Z(n2010) );
  NAND U2197 ( .A(n2011), .B(n2010), .Z(n2043) );
  NANDN U2198 ( .A(n295), .B(a[40]), .Z(n2044) );
  XNOR U2199 ( .A(n2043), .B(n2044), .Z(n2046) );
  XOR U2200 ( .A(n2045), .B(n2046), .Z(n2040) );
  XOR U2201 ( .A(n2039), .B(n2040), .Z(n2063) );
  NANDN U2202 ( .A(n2013), .B(n2012), .Z(n2017) );
  NANDN U2203 ( .A(n2015), .B(n2014), .Z(n2016) );
  NAND U2204 ( .A(n2017), .B(n2016), .Z(n2061) );
  OR U2205 ( .A(n2019), .B(n2018), .Z(n2023) );
  NAND U2206 ( .A(n2021), .B(n2020), .Z(n2022) );
  AND U2207 ( .A(n2023), .B(n2022), .Z(n2062) );
  XNOR U2208 ( .A(n2061), .B(n2062), .Z(n2064) );
  XNOR U2209 ( .A(n2063), .B(n2064), .Z(n2033) );
  XNOR U2210 ( .A(n2033), .B(n2034), .Z(n2035) );
  XNOR U2211 ( .A(n2036), .B(n2035), .Z(n2067) );
  XNOR U2212 ( .A(n2067), .B(sreg[168]), .Z(n2069) );
  NAND U2213 ( .A(n2028), .B(sreg[167]), .Z(n2032) );
  OR U2214 ( .A(n2030), .B(n2029), .Z(n2031) );
  AND U2215 ( .A(n2032), .B(n2031), .Z(n2068) );
  XOR U2216 ( .A(n2069), .B(n2068), .Z(c[168]) );
  NANDN U2217 ( .A(n2038), .B(n2037), .Z(n2042) );
  NAND U2218 ( .A(n2040), .B(n2039), .Z(n2041) );
  NAND U2219 ( .A(n2042), .B(n2041), .Z(n2103) );
  NANDN U2220 ( .A(n2044), .B(n2043), .Z(n2048) );
  NAND U2221 ( .A(n2046), .B(n2045), .Z(n2047) );
  NAND U2222 ( .A(n2048), .B(n2047), .Z(n2101) );
  XNOR U2223 ( .A(b[7]), .B(a[43]), .Z(n2088) );
  NANDN U2224 ( .A(n2088), .B(n5293), .Z(n2051) );
  NANDN U2225 ( .A(n2049), .B(n5294), .Z(n2050) );
  NAND U2226 ( .A(n2051), .B(n2050), .Z(n2076) );
  XNOR U2227 ( .A(b[3]), .B(a[47]), .Z(n2091) );
  NANDN U2228 ( .A(n2091), .B(n5160), .Z(n2054) );
  NANDN U2229 ( .A(n2052), .B(n5161), .Z(n2053) );
  AND U2230 ( .A(n2054), .B(n2053), .Z(n2077) );
  XNOR U2231 ( .A(n2076), .B(n2077), .Z(n2078) );
  NANDN U2232 ( .A(n292), .B(a[49]), .Z(n2055) );
  XOR U2233 ( .A(n5199), .B(n2055), .Z(n2057) );
  NANDN U2234 ( .A(b[0]), .B(a[48]), .Z(n2056) );
  AND U2235 ( .A(n2057), .B(n2056), .Z(n2084) );
  XNOR U2236 ( .A(b[5]), .B(a[45]), .Z(n2097) );
  NANDN U2237 ( .A(n2097), .B(n5240), .Z(n2060) );
  NANDN U2238 ( .A(n2058), .B(n5241), .Z(n2059) );
  NAND U2239 ( .A(n2060), .B(n2059), .Z(n2082) );
  NANDN U2240 ( .A(n295), .B(a[41]), .Z(n2083) );
  XNOR U2241 ( .A(n2082), .B(n2083), .Z(n2085) );
  XOR U2242 ( .A(n2084), .B(n2085), .Z(n2079) );
  XOR U2243 ( .A(n2078), .B(n2079), .Z(n2100) );
  XOR U2244 ( .A(n2101), .B(n2100), .Z(n2102) );
  XNOR U2245 ( .A(n2103), .B(n2102), .Z(n2072) );
  NANDN U2246 ( .A(n2062), .B(n2061), .Z(n2066) );
  NAND U2247 ( .A(n2064), .B(n2063), .Z(n2065) );
  NAND U2248 ( .A(n2066), .B(n2065), .Z(n2073) );
  XNOR U2249 ( .A(n2072), .B(n2073), .Z(n2074) );
  XNOR U2250 ( .A(n2075), .B(n2074), .Z(n2106) );
  XNOR U2251 ( .A(n2106), .B(sreg[169]), .Z(n2108) );
  NAND U2252 ( .A(n2067), .B(sreg[168]), .Z(n2071) );
  OR U2253 ( .A(n2069), .B(n2068), .Z(n2070) );
  AND U2254 ( .A(n2071), .B(n2070), .Z(n2107) );
  XOR U2255 ( .A(n2108), .B(n2107), .Z(c[169]) );
  NANDN U2256 ( .A(n2077), .B(n2076), .Z(n2081) );
  NAND U2257 ( .A(n2079), .B(n2078), .Z(n2080) );
  NAND U2258 ( .A(n2081), .B(n2080), .Z(n2142) );
  NANDN U2259 ( .A(n2083), .B(n2082), .Z(n2087) );
  NAND U2260 ( .A(n2085), .B(n2084), .Z(n2086) );
  NAND U2261 ( .A(n2087), .B(n2086), .Z(n2140) );
  XNOR U2262 ( .A(b[7]), .B(a[44]), .Z(n2127) );
  NANDN U2263 ( .A(n2127), .B(n5293), .Z(n2090) );
  NANDN U2264 ( .A(n2088), .B(n5294), .Z(n2089) );
  NAND U2265 ( .A(n2090), .B(n2089), .Z(n2115) );
  XNOR U2266 ( .A(b[3]), .B(a[48]), .Z(n2130) );
  NANDN U2267 ( .A(n2130), .B(n5160), .Z(n2093) );
  NANDN U2268 ( .A(n2091), .B(n5161), .Z(n2092) );
  AND U2269 ( .A(n2093), .B(n2092), .Z(n2116) );
  XNOR U2270 ( .A(n2115), .B(n2116), .Z(n2117) );
  NANDN U2271 ( .A(n292), .B(a[50]), .Z(n2094) );
  XOR U2272 ( .A(n5199), .B(n2094), .Z(n2096) );
  NANDN U2273 ( .A(b[0]), .B(a[49]), .Z(n2095) );
  AND U2274 ( .A(n2096), .B(n2095), .Z(n2123) );
  XNOR U2275 ( .A(b[5]), .B(a[46]), .Z(n2136) );
  NANDN U2276 ( .A(n2136), .B(n5240), .Z(n2099) );
  NANDN U2277 ( .A(n2097), .B(n5241), .Z(n2098) );
  NAND U2278 ( .A(n2099), .B(n2098), .Z(n2121) );
  NANDN U2279 ( .A(n295), .B(a[42]), .Z(n2122) );
  XNOR U2280 ( .A(n2121), .B(n2122), .Z(n2124) );
  XOR U2281 ( .A(n2123), .B(n2124), .Z(n2118) );
  XOR U2282 ( .A(n2117), .B(n2118), .Z(n2139) );
  XOR U2283 ( .A(n2140), .B(n2139), .Z(n2141) );
  XNOR U2284 ( .A(n2142), .B(n2141), .Z(n2111) );
  NAND U2285 ( .A(n2101), .B(n2100), .Z(n2105) );
  NAND U2286 ( .A(n2103), .B(n2102), .Z(n2104) );
  NAND U2287 ( .A(n2105), .B(n2104), .Z(n2112) );
  XNOR U2288 ( .A(n2111), .B(n2112), .Z(n2113) );
  XNOR U2289 ( .A(n2114), .B(n2113), .Z(n2145) );
  XNOR U2290 ( .A(n2145), .B(sreg[170]), .Z(n2147) );
  NAND U2291 ( .A(n2106), .B(sreg[169]), .Z(n2110) );
  OR U2292 ( .A(n2108), .B(n2107), .Z(n2109) );
  AND U2293 ( .A(n2110), .B(n2109), .Z(n2146) );
  XOR U2294 ( .A(n2147), .B(n2146), .Z(c[170]) );
  NANDN U2295 ( .A(n2116), .B(n2115), .Z(n2120) );
  NAND U2296 ( .A(n2118), .B(n2117), .Z(n2119) );
  NAND U2297 ( .A(n2120), .B(n2119), .Z(n2181) );
  NANDN U2298 ( .A(n2122), .B(n2121), .Z(n2126) );
  NAND U2299 ( .A(n2124), .B(n2123), .Z(n2125) );
  NAND U2300 ( .A(n2126), .B(n2125), .Z(n2179) );
  XNOR U2301 ( .A(b[7]), .B(a[45]), .Z(n2166) );
  NANDN U2302 ( .A(n2166), .B(n5293), .Z(n2129) );
  NANDN U2303 ( .A(n2127), .B(n5294), .Z(n2128) );
  NAND U2304 ( .A(n2129), .B(n2128), .Z(n2154) );
  XNOR U2305 ( .A(b[3]), .B(a[49]), .Z(n2169) );
  NANDN U2306 ( .A(n2169), .B(n5160), .Z(n2132) );
  NANDN U2307 ( .A(n2130), .B(n5161), .Z(n2131) );
  AND U2308 ( .A(n2132), .B(n2131), .Z(n2155) );
  XNOR U2309 ( .A(n2154), .B(n2155), .Z(n2156) );
  NANDN U2310 ( .A(n292), .B(a[51]), .Z(n2133) );
  XOR U2311 ( .A(n5199), .B(n2133), .Z(n2135) );
  NANDN U2312 ( .A(b[0]), .B(a[50]), .Z(n2134) );
  AND U2313 ( .A(n2135), .B(n2134), .Z(n2162) );
  XNOR U2314 ( .A(b[5]), .B(a[47]), .Z(n2175) );
  NANDN U2315 ( .A(n2175), .B(n5240), .Z(n2138) );
  NANDN U2316 ( .A(n2136), .B(n5241), .Z(n2137) );
  NAND U2317 ( .A(n2138), .B(n2137), .Z(n2160) );
  NANDN U2318 ( .A(n295), .B(a[43]), .Z(n2161) );
  XNOR U2319 ( .A(n2160), .B(n2161), .Z(n2163) );
  XOR U2320 ( .A(n2162), .B(n2163), .Z(n2157) );
  XOR U2321 ( .A(n2156), .B(n2157), .Z(n2178) );
  XOR U2322 ( .A(n2179), .B(n2178), .Z(n2180) );
  XNOR U2323 ( .A(n2181), .B(n2180), .Z(n2150) );
  NAND U2324 ( .A(n2140), .B(n2139), .Z(n2144) );
  NAND U2325 ( .A(n2142), .B(n2141), .Z(n2143) );
  NAND U2326 ( .A(n2144), .B(n2143), .Z(n2151) );
  XNOR U2327 ( .A(n2150), .B(n2151), .Z(n2152) );
  XNOR U2328 ( .A(n2153), .B(n2152), .Z(n2184) );
  XNOR U2329 ( .A(n2184), .B(sreg[171]), .Z(n2186) );
  NAND U2330 ( .A(n2145), .B(sreg[170]), .Z(n2149) );
  OR U2331 ( .A(n2147), .B(n2146), .Z(n2148) );
  AND U2332 ( .A(n2149), .B(n2148), .Z(n2185) );
  XOR U2333 ( .A(n2186), .B(n2185), .Z(c[171]) );
  NANDN U2334 ( .A(n2155), .B(n2154), .Z(n2159) );
  NAND U2335 ( .A(n2157), .B(n2156), .Z(n2158) );
  NAND U2336 ( .A(n2159), .B(n2158), .Z(n2220) );
  NANDN U2337 ( .A(n2161), .B(n2160), .Z(n2165) );
  NAND U2338 ( .A(n2163), .B(n2162), .Z(n2164) );
  NAND U2339 ( .A(n2165), .B(n2164), .Z(n2218) );
  XNOR U2340 ( .A(b[7]), .B(a[46]), .Z(n2205) );
  NANDN U2341 ( .A(n2205), .B(n5293), .Z(n2168) );
  NANDN U2342 ( .A(n2166), .B(n5294), .Z(n2167) );
  NAND U2343 ( .A(n2168), .B(n2167), .Z(n2193) );
  XNOR U2344 ( .A(b[3]), .B(a[50]), .Z(n2208) );
  NANDN U2345 ( .A(n2208), .B(n5160), .Z(n2171) );
  NANDN U2346 ( .A(n2169), .B(n5161), .Z(n2170) );
  AND U2347 ( .A(n2171), .B(n2170), .Z(n2194) );
  XNOR U2348 ( .A(n2193), .B(n2194), .Z(n2195) );
  NANDN U2349 ( .A(n292), .B(a[52]), .Z(n2172) );
  XOR U2350 ( .A(n5199), .B(n2172), .Z(n2174) );
  NANDN U2351 ( .A(b[0]), .B(a[51]), .Z(n2173) );
  AND U2352 ( .A(n2174), .B(n2173), .Z(n2201) );
  XNOR U2353 ( .A(b[5]), .B(a[48]), .Z(n2214) );
  NANDN U2354 ( .A(n2214), .B(n5240), .Z(n2177) );
  NANDN U2355 ( .A(n2175), .B(n5241), .Z(n2176) );
  NAND U2356 ( .A(n2177), .B(n2176), .Z(n2199) );
  NANDN U2357 ( .A(n295), .B(a[44]), .Z(n2200) );
  XNOR U2358 ( .A(n2199), .B(n2200), .Z(n2202) );
  XOR U2359 ( .A(n2201), .B(n2202), .Z(n2196) );
  XOR U2360 ( .A(n2195), .B(n2196), .Z(n2217) );
  XOR U2361 ( .A(n2218), .B(n2217), .Z(n2219) );
  XNOR U2362 ( .A(n2220), .B(n2219), .Z(n2189) );
  NAND U2363 ( .A(n2179), .B(n2178), .Z(n2183) );
  NAND U2364 ( .A(n2181), .B(n2180), .Z(n2182) );
  NAND U2365 ( .A(n2183), .B(n2182), .Z(n2190) );
  XNOR U2366 ( .A(n2189), .B(n2190), .Z(n2191) );
  XNOR U2367 ( .A(n2192), .B(n2191), .Z(n2223) );
  XNOR U2368 ( .A(n2223), .B(sreg[172]), .Z(n2225) );
  NAND U2369 ( .A(n2184), .B(sreg[171]), .Z(n2188) );
  OR U2370 ( .A(n2186), .B(n2185), .Z(n2187) );
  AND U2371 ( .A(n2188), .B(n2187), .Z(n2224) );
  XOR U2372 ( .A(n2225), .B(n2224), .Z(c[172]) );
  NANDN U2373 ( .A(n2194), .B(n2193), .Z(n2198) );
  NAND U2374 ( .A(n2196), .B(n2195), .Z(n2197) );
  NAND U2375 ( .A(n2198), .B(n2197), .Z(n2259) );
  NANDN U2376 ( .A(n2200), .B(n2199), .Z(n2204) );
  NAND U2377 ( .A(n2202), .B(n2201), .Z(n2203) );
  NAND U2378 ( .A(n2204), .B(n2203), .Z(n2257) );
  XNOR U2379 ( .A(b[7]), .B(a[47]), .Z(n2244) );
  NANDN U2380 ( .A(n2244), .B(n5293), .Z(n2207) );
  NANDN U2381 ( .A(n2205), .B(n5294), .Z(n2206) );
  NAND U2382 ( .A(n2207), .B(n2206), .Z(n2232) );
  XNOR U2383 ( .A(b[3]), .B(a[51]), .Z(n2247) );
  NANDN U2384 ( .A(n2247), .B(n5160), .Z(n2210) );
  NANDN U2385 ( .A(n2208), .B(n5161), .Z(n2209) );
  AND U2386 ( .A(n2210), .B(n2209), .Z(n2233) );
  XNOR U2387 ( .A(n2232), .B(n2233), .Z(n2234) );
  NANDN U2388 ( .A(n292), .B(a[53]), .Z(n2211) );
  XOR U2389 ( .A(n5199), .B(n2211), .Z(n2213) );
  NANDN U2390 ( .A(b[0]), .B(a[52]), .Z(n2212) );
  AND U2391 ( .A(n2213), .B(n2212), .Z(n2240) );
  XNOR U2392 ( .A(b[5]), .B(a[49]), .Z(n2253) );
  NANDN U2393 ( .A(n2253), .B(n5240), .Z(n2216) );
  NANDN U2394 ( .A(n2214), .B(n5241), .Z(n2215) );
  NAND U2395 ( .A(n2216), .B(n2215), .Z(n2238) );
  NANDN U2396 ( .A(n295), .B(a[45]), .Z(n2239) );
  XNOR U2397 ( .A(n2238), .B(n2239), .Z(n2241) );
  XOR U2398 ( .A(n2240), .B(n2241), .Z(n2235) );
  XOR U2399 ( .A(n2234), .B(n2235), .Z(n2256) );
  XOR U2400 ( .A(n2257), .B(n2256), .Z(n2258) );
  XNOR U2401 ( .A(n2259), .B(n2258), .Z(n2228) );
  NAND U2402 ( .A(n2218), .B(n2217), .Z(n2222) );
  NAND U2403 ( .A(n2220), .B(n2219), .Z(n2221) );
  NAND U2404 ( .A(n2222), .B(n2221), .Z(n2229) );
  XNOR U2405 ( .A(n2228), .B(n2229), .Z(n2230) );
  XNOR U2406 ( .A(n2231), .B(n2230), .Z(n2262) );
  XNOR U2407 ( .A(n2262), .B(sreg[173]), .Z(n2264) );
  NAND U2408 ( .A(n2223), .B(sreg[172]), .Z(n2227) );
  OR U2409 ( .A(n2225), .B(n2224), .Z(n2226) );
  AND U2410 ( .A(n2227), .B(n2226), .Z(n2263) );
  XOR U2411 ( .A(n2264), .B(n2263), .Z(c[173]) );
  NANDN U2412 ( .A(n2233), .B(n2232), .Z(n2237) );
  NAND U2413 ( .A(n2235), .B(n2234), .Z(n2236) );
  NAND U2414 ( .A(n2237), .B(n2236), .Z(n2298) );
  NANDN U2415 ( .A(n2239), .B(n2238), .Z(n2243) );
  NAND U2416 ( .A(n2241), .B(n2240), .Z(n2242) );
  NAND U2417 ( .A(n2243), .B(n2242), .Z(n2296) );
  XNOR U2418 ( .A(b[7]), .B(a[48]), .Z(n2283) );
  NANDN U2419 ( .A(n2283), .B(n5293), .Z(n2246) );
  NANDN U2420 ( .A(n2244), .B(n5294), .Z(n2245) );
  NAND U2421 ( .A(n2246), .B(n2245), .Z(n2271) );
  XNOR U2422 ( .A(b[3]), .B(a[52]), .Z(n2286) );
  NANDN U2423 ( .A(n2286), .B(n5160), .Z(n2249) );
  NANDN U2424 ( .A(n2247), .B(n5161), .Z(n2248) );
  AND U2425 ( .A(n2249), .B(n2248), .Z(n2272) );
  XNOR U2426 ( .A(n2271), .B(n2272), .Z(n2273) );
  NANDN U2427 ( .A(n292), .B(a[54]), .Z(n2250) );
  XOR U2428 ( .A(n5199), .B(n2250), .Z(n2252) );
  NANDN U2429 ( .A(b[0]), .B(a[53]), .Z(n2251) );
  AND U2430 ( .A(n2252), .B(n2251), .Z(n2279) );
  XNOR U2431 ( .A(b[5]), .B(a[50]), .Z(n2292) );
  NANDN U2432 ( .A(n2292), .B(n5240), .Z(n2255) );
  NANDN U2433 ( .A(n2253), .B(n5241), .Z(n2254) );
  NAND U2434 ( .A(n2255), .B(n2254), .Z(n2277) );
  NANDN U2435 ( .A(n295), .B(a[46]), .Z(n2278) );
  XNOR U2436 ( .A(n2277), .B(n2278), .Z(n2280) );
  XOR U2437 ( .A(n2279), .B(n2280), .Z(n2274) );
  XOR U2438 ( .A(n2273), .B(n2274), .Z(n2295) );
  XOR U2439 ( .A(n2296), .B(n2295), .Z(n2297) );
  XNOR U2440 ( .A(n2298), .B(n2297), .Z(n2267) );
  NAND U2441 ( .A(n2257), .B(n2256), .Z(n2261) );
  NAND U2442 ( .A(n2259), .B(n2258), .Z(n2260) );
  NAND U2443 ( .A(n2261), .B(n2260), .Z(n2268) );
  XNOR U2444 ( .A(n2267), .B(n2268), .Z(n2269) );
  XNOR U2445 ( .A(n2270), .B(n2269), .Z(n2301) );
  XNOR U2446 ( .A(n2301), .B(sreg[174]), .Z(n2303) );
  NAND U2447 ( .A(n2262), .B(sreg[173]), .Z(n2266) );
  OR U2448 ( .A(n2264), .B(n2263), .Z(n2265) );
  AND U2449 ( .A(n2266), .B(n2265), .Z(n2302) );
  XOR U2450 ( .A(n2303), .B(n2302), .Z(c[174]) );
  NANDN U2451 ( .A(n2272), .B(n2271), .Z(n2276) );
  NAND U2452 ( .A(n2274), .B(n2273), .Z(n2275) );
  NAND U2453 ( .A(n2276), .B(n2275), .Z(n2337) );
  NANDN U2454 ( .A(n2278), .B(n2277), .Z(n2282) );
  NAND U2455 ( .A(n2280), .B(n2279), .Z(n2281) );
  NAND U2456 ( .A(n2282), .B(n2281), .Z(n2335) );
  XNOR U2457 ( .A(b[7]), .B(a[49]), .Z(n2328) );
  NANDN U2458 ( .A(n2328), .B(n5293), .Z(n2285) );
  NANDN U2459 ( .A(n2283), .B(n5294), .Z(n2284) );
  NAND U2460 ( .A(n2285), .B(n2284), .Z(n2310) );
  XNOR U2461 ( .A(b[3]), .B(a[53]), .Z(n2331) );
  NANDN U2462 ( .A(n2331), .B(n5160), .Z(n2288) );
  NANDN U2463 ( .A(n2286), .B(n5161), .Z(n2287) );
  AND U2464 ( .A(n2288), .B(n2287), .Z(n2311) );
  XNOR U2465 ( .A(n2310), .B(n2311), .Z(n2312) );
  NANDN U2466 ( .A(n292), .B(a[55]), .Z(n2289) );
  XOR U2467 ( .A(n5199), .B(n2289), .Z(n2291) );
  IV U2468 ( .A(a[54]), .Z(n2554) );
  NANDN U2469 ( .A(n2554), .B(n292), .Z(n2290) );
  AND U2470 ( .A(n2291), .B(n2290), .Z(n2318) );
  XNOR U2471 ( .A(b[5]), .B(a[51]), .Z(n2325) );
  NANDN U2472 ( .A(n2325), .B(n5240), .Z(n2294) );
  NANDN U2473 ( .A(n2292), .B(n5241), .Z(n2293) );
  NAND U2474 ( .A(n2294), .B(n2293), .Z(n2316) );
  NANDN U2475 ( .A(n295), .B(a[47]), .Z(n2317) );
  XNOR U2476 ( .A(n2316), .B(n2317), .Z(n2319) );
  XOR U2477 ( .A(n2318), .B(n2319), .Z(n2313) );
  XOR U2478 ( .A(n2312), .B(n2313), .Z(n2334) );
  XOR U2479 ( .A(n2335), .B(n2334), .Z(n2336) );
  XNOR U2480 ( .A(n2337), .B(n2336), .Z(n2306) );
  NAND U2481 ( .A(n2296), .B(n2295), .Z(n2300) );
  NAND U2482 ( .A(n2298), .B(n2297), .Z(n2299) );
  NAND U2483 ( .A(n2300), .B(n2299), .Z(n2307) );
  XNOR U2484 ( .A(n2306), .B(n2307), .Z(n2308) );
  XNOR U2485 ( .A(n2309), .B(n2308), .Z(n2340) );
  XNOR U2486 ( .A(n2340), .B(sreg[175]), .Z(n2342) );
  NAND U2487 ( .A(n2301), .B(sreg[174]), .Z(n2305) );
  OR U2488 ( .A(n2303), .B(n2302), .Z(n2304) );
  AND U2489 ( .A(n2305), .B(n2304), .Z(n2341) );
  XOR U2490 ( .A(n2342), .B(n2341), .Z(c[175]) );
  NANDN U2491 ( .A(n2311), .B(n2310), .Z(n2315) );
  NAND U2492 ( .A(n2313), .B(n2312), .Z(n2314) );
  NAND U2493 ( .A(n2315), .B(n2314), .Z(n2376) );
  NANDN U2494 ( .A(n2317), .B(n2316), .Z(n2321) );
  NAND U2495 ( .A(n2319), .B(n2318), .Z(n2320) );
  NAND U2496 ( .A(n2321), .B(n2320), .Z(n2374) );
  NANDN U2497 ( .A(n292), .B(a[56]), .Z(n2322) );
  XOR U2498 ( .A(n5199), .B(n2322), .Z(n2324) );
  NANDN U2499 ( .A(b[0]), .B(a[55]), .Z(n2323) );
  AND U2500 ( .A(n2324), .B(n2323), .Z(n2357) );
  XNOR U2501 ( .A(b[5]), .B(a[52]), .Z(n2370) );
  NANDN U2502 ( .A(n2370), .B(n5240), .Z(n2327) );
  NANDN U2503 ( .A(n2325), .B(n5241), .Z(n2326) );
  NAND U2504 ( .A(n2327), .B(n2326), .Z(n2355) );
  NANDN U2505 ( .A(n295), .B(a[48]), .Z(n2356) );
  XNOR U2506 ( .A(n2355), .B(n2356), .Z(n2358) );
  XOR U2507 ( .A(n2357), .B(n2358), .Z(n2351) );
  XNOR U2508 ( .A(b[7]), .B(a[50]), .Z(n2361) );
  NANDN U2509 ( .A(n2361), .B(n5293), .Z(n2330) );
  NANDN U2510 ( .A(n2328), .B(n5294), .Z(n2329) );
  NAND U2511 ( .A(n2330), .B(n2329), .Z(n2349) );
  XOR U2512 ( .A(b[3]), .B(n2554), .Z(n2364) );
  NANDN U2513 ( .A(n2364), .B(n5160), .Z(n2333) );
  NANDN U2514 ( .A(n2331), .B(n5161), .Z(n2332) );
  AND U2515 ( .A(n2333), .B(n2332), .Z(n2350) );
  XNOR U2516 ( .A(n2349), .B(n2350), .Z(n2352) );
  XOR U2517 ( .A(n2351), .B(n2352), .Z(n2373) );
  XOR U2518 ( .A(n2374), .B(n2373), .Z(n2375) );
  XNOR U2519 ( .A(n2376), .B(n2375), .Z(n2345) );
  NAND U2520 ( .A(n2335), .B(n2334), .Z(n2339) );
  NAND U2521 ( .A(n2337), .B(n2336), .Z(n2338) );
  NAND U2522 ( .A(n2339), .B(n2338), .Z(n2346) );
  XNOR U2523 ( .A(n2345), .B(n2346), .Z(n2347) );
  XNOR U2524 ( .A(n2348), .B(n2347), .Z(n2379) );
  XNOR U2525 ( .A(n2379), .B(sreg[176]), .Z(n2381) );
  NAND U2526 ( .A(n2340), .B(sreg[175]), .Z(n2344) );
  OR U2527 ( .A(n2342), .B(n2341), .Z(n2343) );
  AND U2528 ( .A(n2344), .B(n2343), .Z(n2380) );
  XOR U2529 ( .A(n2381), .B(n2380), .Z(c[176]) );
  NANDN U2530 ( .A(n2350), .B(n2349), .Z(n2354) );
  NAND U2531 ( .A(n2352), .B(n2351), .Z(n2353) );
  NAND U2532 ( .A(n2354), .B(n2353), .Z(n2415) );
  NANDN U2533 ( .A(n2356), .B(n2355), .Z(n2360) );
  NAND U2534 ( .A(n2358), .B(n2357), .Z(n2359) );
  NAND U2535 ( .A(n2360), .B(n2359), .Z(n2413) );
  XNOR U2536 ( .A(b[7]), .B(a[51]), .Z(n2400) );
  NANDN U2537 ( .A(n2400), .B(n5293), .Z(n2363) );
  NANDN U2538 ( .A(n2361), .B(n5294), .Z(n2362) );
  NAND U2539 ( .A(n2363), .B(n2362), .Z(n2388) );
  XNOR U2540 ( .A(b[3]), .B(a[55]), .Z(n2403) );
  NANDN U2541 ( .A(n2403), .B(n5160), .Z(n2366) );
  NANDN U2542 ( .A(n2364), .B(n5161), .Z(n2365) );
  AND U2543 ( .A(n2366), .B(n2365), .Z(n2389) );
  XNOR U2544 ( .A(n2388), .B(n2389), .Z(n2390) );
  NANDN U2545 ( .A(n292), .B(a[57]), .Z(n2367) );
  XOR U2546 ( .A(n5199), .B(n2367), .Z(n2369) );
  NANDN U2547 ( .A(b[0]), .B(a[56]), .Z(n2368) );
  AND U2548 ( .A(n2369), .B(n2368), .Z(n2396) );
  XNOR U2549 ( .A(n294), .B(a[53]), .Z(n2406) );
  NAND U2550 ( .A(n2406), .B(n5240), .Z(n2372) );
  NANDN U2551 ( .A(n2370), .B(n5241), .Z(n2371) );
  NAND U2552 ( .A(n2372), .B(n2371), .Z(n2394) );
  NANDN U2553 ( .A(n295), .B(a[49]), .Z(n2395) );
  XNOR U2554 ( .A(n2394), .B(n2395), .Z(n2397) );
  XOR U2555 ( .A(n2396), .B(n2397), .Z(n2391) );
  XOR U2556 ( .A(n2390), .B(n2391), .Z(n2412) );
  XOR U2557 ( .A(n2413), .B(n2412), .Z(n2414) );
  XNOR U2558 ( .A(n2415), .B(n2414), .Z(n2384) );
  NAND U2559 ( .A(n2374), .B(n2373), .Z(n2378) );
  NAND U2560 ( .A(n2376), .B(n2375), .Z(n2377) );
  NAND U2561 ( .A(n2378), .B(n2377), .Z(n2385) );
  XNOR U2562 ( .A(n2384), .B(n2385), .Z(n2386) );
  XNOR U2563 ( .A(n2387), .B(n2386), .Z(n2418) );
  XNOR U2564 ( .A(n2418), .B(sreg[177]), .Z(n2420) );
  NAND U2565 ( .A(n2379), .B(sreg[176]), .Z(n2383) );
  OR U2566 ( .A(n2381), .B(n2380), .Z(n2382) );
  AND U2567 ( .A(n2383), .B(n2382), .Z(n2419) );
  XOR U2568 ( .A(n2420), .B(n2419), .Z(c[177]) );
  NANDN U2569 ( .A(n2389), .B(n2388), .Z(n2393) );
  NAND U2570 ( .A(n2391), .B(n2390), .Z(n2392) );
  NAND U2571 ( .A(n2393), .B(n2392), .Z(n2454) );
  NANDN U2572 ( .A(n2395), .B(n2394), .Z(n2399) );
  NAND U2573 ( .A(n2397), .B(n2396), .Z(n2398) );
  NAND U2574 ( .A(n2399), .B(n2398), .Z(n2452) );
  XNOR U2575 ( .A(b[7]), .B(a[52]), .Z(n2427) );
  NANDN U2576 ( .A(n2427), .B(n5293), .Z(n2402) );
  NANDN U2577 ( .A(n2400), .B(n5294), .Z(n2401) );
  NAND U2578 ( .A(n2402), .B(n2401), .Z(n2439) );
  XNOR U2579 ( .A(b[3]), .B(a[56]), .Z(n2430) );
  NANDN U2580 ( .A(n2430), .B(n5160), .Z(n2405) );
  NANDN U2581 ( .A(n2403), .B(n5161), .Z(n2404) );
  AND U2582 ( .A(n2405), .B(n2404), .Z(n2440) );
  XNOR U2583 ( .A(n2439), .B(n2440), .Z(n2441) );
  NANDN U2584 ( .A(n295), .B(a[50]), .Z(n2446) );
  XOR U2585 ( .A(b[5]), .B(n2554), .Z(n2436) );
  NANDN U2586 ( .A(n2436), .B(n5240), .Z(n2408) );
  NAND U2587 ( .A(n5241), .B(n2406), .Z(n2407) );
  AND U2588 ( .A(n2408), .B(n2407), .Z(n2445) );
  XOR U2589 ( .A(n2446), .B(n2445), .Z(n2448) );
  NANDN U2590 ( .A(n292), .B(a[58]), .Z(n2409) );
  XOR U2591 ( .A(n5199), .B(n2409), .Z(n2411) );
  NANDN U2592 ( .A(b[0]), .B(a[57]), .Z(n2410) );
  AND U2593 ( .A(n2411), .B(n2410), .Z(n2447) );
  XNOR U2594 ( .A(n2448), .B(n2447), .Z(n2442) );
  XNOR U2595 ( .A(n2441), .B(n2442), .Z(n2451) );
  XOR U2596 ( .A(n2452), .B(n2451), .Z(n2453) );
  XNOR U2597 ( .A(n2454), .B(n2453), .Z(n2423) );
  NAND U2598 ( .A(n2413), .B(n2412), .Z(n2417) );
  NAND U2599 ( .A(n2415), .B(n2414), .Z(n2416) );
  NAND U2600 ( .A(n2417), .B(n2416), .Z(n2424) );
  XNOR U2601 ( .A(n2423), .B(n2424), .Z(n2425) );
  XNOR U2602 ( .A(n2426), .B(n2425), .Z(n2455) );
  XNOR U2603 ( .A(n2455), .B(sreg[178]), .Z(n2457) );
  NAND U2604 ( .A(n2418), .B(sreg[177]), .Z(n2422) );
  OR U2605 ( .A(n2420), .B(n2419), .Z(n2421) );
  AND U2606 ( .A(n2422), .B(n2421), .Z(n2456) );
  XOR U2607 ( .A(n2457), .B(n2456), .Z(c[178]) );
  XNOR U2608 ( .A(b[7]), .B(a[53]), .Z(n2476) );
  NANDN U2609 ( .A(n2476), .B(n5293), .Z(n2429) );
  NANDN U2610 ( .A(n2427), .B(n5294), .Z(n2428) );
  NAND U2611 ( .A(n2429), .B(n2428), .Z(n2464) );
  XNOR U2612 ( .A(b[3]), .B(a[57]), .Z(n2479) );
  NANDN U2613 ( .A(n2479), .B(n5160), .Z(n2432) );
  NANDN U2614 ( .A(n2430), .B(n5161), .Z(n2431) );
  AND U2615 ( .A(n2432), .B(n2431), .Z(n2465) );
  XNOR U2616 ( .A(n2464), .B(n2465), .Z(n2466) );
  NANDN U2617 ( .A(n292), .B(a[59]), .Z(n2433) );
  XOR U2618 ( .A(n5199), .B(n2433), .Z(n2435) );
  NANDN U2619 ( .A(b[0]), .B(a[58]), .Z(n2434) );
  AND U2620 ( .A(n2435), .B(n2434), .Z(n2472) );
  XNOR U2621 ( .A(b[5]), .B(a[55]), .Z(n2485) );
  NANDN U2622 ( .A(n2485), .B(n5240), .Z(n2438) );
  NANDN U2623 ( .A(n2436), .B(n5241), .Z(n2437) );
  NAND U2624 ( .A(n2438), .B(n2437), .Z(n2470) );
  NANDN U2625 ( .A(n295), .B(a[51]), .Z(n2471) );
  XNOR U2626 ( .A(n2470), .B(n2471), .Z(n2473) );
  XOR U2627 ( .A(n2472), .B(n2473), .Z(n2467) );
  XOR U2628 ( .A(n2466), .B(n2467), .Z(n2490) );
  NANDN U2629 ( .A(n2440), .B(n2439), .Z(n2444) );
  NANDN U2630 ( .A(n2442), .B(n2441), .Z(n2443) );
  NAND U2631 ( .A(n2444), .B(n2443), .Z(n2488) );
  OR U2632 ( .A(n2446), .B(n2445), .Z(n2450) );
  NAND U2633 ( .A(n2448), .B(n2447), .Z(n2449) );
  AND U2634 ( .A(n2450), .B(n2449), .Z(n2489) );
  XNOR U2635 ( .A(n2488), .B(n2489), .Z(n2491) );
  XNOR U2636 ( .A(n2490), .B(n2491), .Z(n2460) );
  XNOR U2637 ( .A(n2460), .B(n2461), .Z(n2462) );
  XNOR U2638 ( .A(n2463), .B(n2462), .Z(n2494) );
  XNOR U2639 ( .A(n2494), .B(sreg[179]), .Z(n2496) );
  NAND U2640 ( .A(n2455), .B(sreg[178]), .Z(n2459) );
  OR U2641 ( .A(n2457), .B(n2456), .Z(n2458) );
  AND U2642 ( .A(n2459), .B(n2458), .Z(n2495) );
  XOR U2643 ( .A(n2496), .B(n2495), .Z(c[179]) );
  NANDN U2644 ( .A(n2465), .B(n2464), .Z(n2469) );
  NAND U2645 ( .A(n2467), .B(n2466), .Z(n2468) );
  NAND U2646 ( .A(n2469), .B(n2468), .Z(n2530) );
  NANDN U2647 ( .A(n2471), .B(n2470), .Z(n2475) );
  NAND U2648 ( .A(n2473), .B(n2472), .Z(n2474) );
  NAND U2649 ( .A(n2475), .B(n2474), .Z(n2528) );
  XOR U2650 ( .A(b[7]), .B(n2554), .Z(n2515) );
  NANDN U2651 ( .A(n2515), .B(n5293), .Z(n2478) );
  NANDN U2652 ( .A(n2476), .B(n5294), .Z(n2477) );
  NAND U2653 ( .A(n2478), .B(n2477), .Z(n2503) );
  XNOR U2654 ( .A(b[3]), .B(a[58]), .Z(n2518) );
  NANDN U2655 ( .A(n2518), .B(n5160), .Z(n2481) );
  NANDN U2656 ( .A(n2479), .B(n5161), .Z(n2480) );
  AND U2657 ( .A(n2481), .B(n2480), .Z(n2504) );
  XNOR U2658 ( .A(n2503), .B(n2504), .Z(n2505) );
  NANDN U2659 ( .A(n292), .B(a[60]), .Z(n2482) );
  XOR U2660 ( .A(n5199), .B(n2482), .Z(n2484) );
  NANDN U2661 ( .A(b[0]), .B(a[59]), .Z(n2483) );
  AND U2662 ( .A(n2484), .B(n2483), .Z(n2511) );
  XNOR U2663 ( .A(b[5]), .B(a[56]), .Z(n2524) );
  NANDN U2664 ( .A(n2524), .B(n5240), .Z(n2487) );
  NANDN U2665 ( .A(n2485), .B(n5241), .Z(n2486) );
  NAND U2666 ( .A(n2487), .B(n2486), .Z(n2509) );
  NANDN U2667 ( .A(n295), .B(a[52]), .Z(n2510) );
  XNOR U2668 ( .A(n2509), .B(n2510), .Z(n2512) );
  XOR U2669 ( .A(n2511), .B(n2512), .Z(n2506) );
  XOR U2670 ( .A(n2505), .B(n2506), .Z(n2527) );
  XOR U2671 ( .A(n2528), .B(n2527), .Z(n2529) );
  XNOR U2672 ( .A(n2530), .B(n2529), .Z(n2499) );
  NANDN U2673 ( .A(n2489), .B(n2488), .Z(n2493) );
  NAND U2674 ( .A(n2491), .B(n2490), .Z(n2492) );
  NAND U2675 ( .A(n2493), .B(n2492), .Z(n2500) );
  XNOR U2676 ( .A(n2499), .B(n2500), .Z(n2501) );
  XNOR U2677 ( .A(n2502), .B(n2501), .Z(n2533) );
  XNOR U2678 ( .A(n2533), .B(sreg[180]), .Z(n2535) );
  NAND U2679 ( .A(n2494), .B(sreg[179]), .Z(n2498) );
  OR U2680 ( .A(n2496), .B(n2495), .Z(n2497) );
  AND U2681 ( .A(n2498), .B(n2497), .Z(n2534) );
  XOR U2682 ( .A(n2535), .B(n2534), .Z(c[180]) );
  NANDN U2683 ( .A(n2504), .B(n2503), .Z(n2508) );
  NAND U2684 ( .A(n2506), .B(n2505), .Z(n2507) );
  NAND U2685 ( .A(n2508), .B(n2507), .Z(n2570) );
  NANDN U2686 ( .A(n2510), .B(n2509), .Z(n2514) );
  NAND U2687 ( .A(n2512), .B(n2511), .Z(n2513) );
  NAND U2688 ( .A(n2514), .B(n2513), .Z(n2568) );
  XNOR U2689 ( .A(b[7]), .B(a[55]), .Z(n2561) );
  NANDN U2690 ( .A(n2561), .B(n5293), .Z(n2517) );
  NANDN U2691 ( .A(n2515), .B(n5294), .Z(n2516) );
  NAND U2692 ( .A(n2517), .B(n2516), .Z(n2542) );
  XNOR U2693 ( .A(b[3]), .B(a[59]), .Z(n2564) );
  NANDN U2694 ( .A(n2564), .B(n5160), .Z(n2520) );
  NANDN U2695 ( .A(n2518), .B(n5161), .Z(n2519) );
  AND U2696 ( .A(n2520), .B(n2519), .Z(n2543) );
  XNOR U2697 ( .A(n2542), .B(n2543), .Z(n2544) );
  NANDN U2698 ( .A(n292), .B(a[61]), .Z(n2521) );
  XOR U2699 ( .A(n5199), .B(n2521), .Z(n2523) );
  NANDN U2700 ( .A(b[0]), .B(a[60]), .Z(n2522) );
  AND U2701 ( .A(n2523), .B(n2522), .Z(n2550) );
  XNOR U2702 ( .A(n294), .B(a[57]), .Z(n2555) );
  NAND U2703 ( .A(n2555), .B(n5240), .Z(n2526) );
  NANDN U2704 ( .A(n2524), .B(n5241), .Z(n2525) );
  NAND U2705 ( .A(n2526), .B(n2525), .Z(n2548) );
  NANDN U2706 ( .A(n295), .B(a[53]), .Z(n2549) );
  XNOR U2707 ( .A(n2548), .B(n2549), .Z(n2551) );
  XOR U2708 ( .A(n2550), .B(n2551), .Z(n2545) );
  XOR U2709 ( .A(n2544), .B(n2545), .Z(n2567) );
  XOR U2710 ( .A(n2568), .B(n2567), .Z(n2569) );
  XNOR U2711 ( .A(n2570), .B(n2569), .Z(n2538) );
  NAND U2712 ( .A(n2528), .B(n2527), .Z(n2532) );
  NAND U2713 ( .A(n2530), .B(n2529), .Z(n2531) );
  NAND U2714 ( .A(n2532), .B(n2531), .Z(n2539) );
  XNOR U2715 ( .A(n2538), .B(n2539), .Z(n2540) );
  XNOR U2716 ( .A(n2541), .B(n2540), .Z(n2573) );
  XNOR U2717 ( .A(n2573), .B(sreg[181]), .Z(n2575) );
  NAND U2718 ( .A(n2533), .B(sreg[180]), .Z(n2537) );
  OR U2719 ( .A(n2535), .B(n2534), .Z(n2536) );
  AND U2720 ( .A(n2537), .B(n2536), .Z(n2574) );
  XOR U2721 ( .A(n2575), .B(n2574), .Z(c[181]) );
  NANDN U2722 ( .A(n2543), .B(n2542), .Z(n2547) );
  NAND U2723 ( .A(n2545), .B(n2544), .Z(n2546) );
  NAND U2724 ( .A(n2547), .B(n2546), .Z(n2609) );
  NANDN U2725 ( .A(n2549), .B(n2548), .Z(n2553) );
  NAND U2726 ( .A(n2551), .B(n2550), .Z(n2552) );
  NAND U2727 ( .A(n2553), .B(n2552), .Z(n2606) );
  ANDN U2728 ( .B(b[7]), .A(n2554), .Z(n2588) );
  XNOR U2729 ( .A(b[5]), .B(a[58]), .Z(n2603) );
  NANDN U2730 ( .A(n2603), .B(n5240), .Z(n2557) );
  NAND U2731 ( .A(n5241), .B(n2555), .Z(n2556) );
  NAND U2732 ( .A(n2557), .B(n2556), .Z(n2589) );
  XOR U2733 ( .A(n2588), .B(n2589), .Z(n2590) );
  NANDN U2734 ( .A(n292), .B(a[62]), .Z(n2558) );
  XOR U2735 ( .A(n5199), .B(n2558), .Z(n2560) );
  NANDN U2736 ( .A(b[0]), .B(a[61]), .Z(n2559) );
  AND U2737 ( .A(n2560), .B(n2559), .Z(n2591) );
  XOR U2738 ( .A(n2590), .B(n2591), .Z(n2585) );
  XNOR U2739 ( .A(b[7]), .B(a[56]), .Z(n2594) );
  NANDN U2740 ( .A(n2594), .B(n5293), .Z(n2563) );
  NANDN U2741 ( .A(n2561), .B(n5294), .Z(n2562) );
  NAND U2742 ( .A(n2563), .B(n2562), .Z(n2582) );
  XNOR U2743 ( .A(b[3]), .B(a[60]), .Z(n2597) );
  NANDN U2744 ( .A(n2597), .B(n5160), .Z(n2566) );
  NANDN U2745 ( .A(n2564), .B(n5161), .Z(n2565) );
  AND U2746 ( .A(n2566), .B(n2565), .Z(n2583) );
  XNOR U2747 ( .A(n2582), .B(n2583), .Z(n2584) );
  XNOR U2748 ( .A(n2585), .B(n2584), .Z(n2607) );
  XNOR U2749 ( .A(n2606), .B(n2607), .Z(n2608) );
  XNOR U2750 ( .A(n2609), .B(n2608), .Z(n2578) );
  NAND U2751 ( .A(n2568), .B(n2567), .Z(n2572) );
  NAND U2752 ( .A(n2570), .B(n2569), .Z(n2571) );
  NAND U2753 ( .A(n2572), .B(n2571), .Z(n2579) );
  XNOR U2754 ( .A(n2578), .B(n2579), .Z(n2580) );
  XNOR U2755 ( .A(n2581), .B(n2580), .Z(n2612) );
  XNOR U2756 ( .A(n2612), .B(sreg[182]), .Z(n2614) );
  NAND U2757 ( .A(n2573), .B(sreg[181]), .Z(n2577) );
  OR U2758 ( .A(n2575), .B(n2574), .Z(n2576) );
  AND U2759 ( .A(n2577), .B(n2576), .Z(n2613) );
  XOR U2760 ( .A(n2614), .B(n2613), .Z(c[182]) );
  NANDN U2761 ( .A(n2583), .B(n2582), .Z(n2587) );
  NAND U2762 ( .A(n2585), .B(n2584), .Z(n2586) );
  NAND U2763 ( .A(n2587), .B(n2586), .Z(n2648) );
  OR U2764 ( .A(n2589), .B(n2588), .Z(n2593) );
  NANDN U2765 ( .A(n2591), .B(n2590), .Z(n2592) );
  NAND U2766 ( .A(n2593), .B(n2592), .Z(n2646) );
  XNOR U2767 ( .A(b[7]), .B(a[57]), .Z(n2633) );
  NANDN U2768 ( .A(n2633), .B(n5293), .Z(n2596) );
  NANDN U2769 ( .A(n2594), .B(n5294), .Z(n2595) );
  NAND U2770 ( .A(n2596), .B(n2595), .Z(n2621) );
  XNOR U2771 ( .A(b[3]), .B(a[61]), .Z(n2636) );
  NANDN U2772 ( .A(n2636), .B(n5160), .Z(n2599) );
  NANDN U2773 ( .A(n2597), .B(n5161), .Z(n2598) );
  AND U2774 ( .A(n2599), .B(n2598), .Z(n2622) );
  XNOR U2775 ( .A(n2621), .B(n2622), .Z(n2623) );
  NANDN U2776 ( .A(n292), .B(a[63]), .Z(n2600) );
  XOR U2777 ( .A(n5199), .B(n2600), .Z(n2602) );
  NANDN U2778 ( .A(b[0]), .B(a[62]), .Z(n2601) );
  AND U2779 ( .A(n2602), .B(n2601), .Z(n2629) );
  XNOR U2780 ( .A(b[5]), .B(a[59]), .Z(n2642) );
  NANDN U2781 ( .A(n2642), .B(n5240), .Z(n2605) );
  NANDN U2782 ( .A(n2603), .B(n5241), .Z(n2604) );
  NAND U2783 ( .A(n2605), .B(n2604), .Z(n2627) );
  NANDN U2784 ( .A(n295), .B(a[55]), .Z(n2628) );
  XNOR U2785 ( .A(n2627), .B(n2628), .Z(n2630) );
  XOR U2786 ( .A(n2629), .B(n2630), .Z(n2624) );
  XOR U2787 ( .A(n2623), .B(n2624), .Z(n2645) );
  XNOR U2788 ( .A(n2646), .B(n2645), .Z(n2647) );
  XNOR U2789 ( .A(n2648), .B(n2647), .Z(n2617) );
  NANDN U2790 ( .A(n2607), .B(n2606), .Z(n2611) );
  NAND U2791 ( .A(n2609), .B(n2608), .Z(n2610) );
  NAND U2792 ( .A(n2611), .B(n2610), .Z(n2618) );
  XNOR U2793 ( .A(n2617), .B(n2618), .Z(n2619) );
  XNOR U2794 ( .A(n2620), .B(n2619), .Z(n2649) );
  XNOR U2795 ( .A(n2649), .B(sreg[183]), .Z(n2651) );
  NAND U2796 ( .A(n2612), .B(sreg[182]), .Z(n2616) );
  OR U2797 ( .A(n2614), .B(n2613), .Z(n2615) );
  AND U2798 ( .A(n2616), .B(n2615), .Z(n2650) );
  XOR U2799 ( .A(n2651), .B(n2650), .Z(c[183]) );
  NANDN U2800 ( .A(n2622), .B(n2621), .Z(n2626) );
  NAND U2801 ( .A(n2624), .B(n2623), .Z(n2625) );
  NAND U2802 ( .A(n2626), .B(n2625), .Z(n2685) );
  NANDN U2803 ( .A(n2628), .B(n2627), .Z(n2632) );
  NAND U2804 ( .A(n2630), .B(n2629), .Z(n2631) );
  NAND U2805 ( .A(n2632), .B(n2631), .Z(n2683) );
  XNOR U2806 ( .A(b[7]), .B(a[58]), .Z(n2670) );
  NANDN U2807 ( .A(n2670), .B(n5293), .Z(n2635) );
  NANDN U2808 ( .A(n2633), .B(n5294), .Z(n2634) );
  NAND U2809 ( .A(n2635), .B(n2634), .Z(n2658) );
  XNOR U2810 ( .A(b[3]), .B(a[62]), .Z(n2673) );
  NANDN U2811 ( .A(n2673), .B(n5160), .Z(n2638) );
  NANDN U2812 ( .A(n2636), .B(n5161), .Z(n2637) );
  AND U2813 ( .A(n2638), .B(n2637), .Z(n2659) );
  XNOR U2814 ( .A(n2658), .B(n2659), .Z(n2660) );
  NANDN U2815 ( .A(n292), .B(a[64]), .Z(n2639) );
  XOR U2816 ( .A(n5199), .B(n2639), .Z(n2641) );
  NANDN U2817 ( .A(b[0]), .B(a[63]), .Z(n2640) );
  AND U2818 ( .A(n2641), .B(n2640), .Z(n2666) );
  XNOR U2819 ( .A(b[5]), .B(a[60]), .Z(n2679) );
  NANDN U2820 ( .A(n2679), .B(n5240), .Z(n2644) );
  NANDN U2821 ( .A(n2642), .B(n5241), .Z(n2643) );
  NAND U2822 ( .A(n2644), .B(n2643), .Z(n2664) );
  NANDN U2823 ( .A(n295), .B(a[56]), .Z(n2665) );
  XNOR U2824 ( .A(n2664), .B(n2665), .Z(n2667) );
  XOR U2825 ( .A(n2666), .B(n2667), .Z(n2661) );
  XOR U2826 ( .A(n2660), .B(n2661), .Z(n2682) );
  XOR U2827 ( .A(n2683), .B(n2682), .Z(n2684) );
  XNOR U2828 ( .A(n2685), .B(n2684), .Z(n2654) );
  XNOR U2829 ( .A(n2654), .B(n2655), .Z(n2656) );
  XNOR U2830 ( .A(n2657), .B(n2656), .Z(n2688) );
  XNOR U2831 ( .A(n2688), .B(sreg[184]), .Z(n2690) );
  NAND U2832 ( .A(n2649), .B(sreg[183]), .Z(n2653) );
  OR U2833 ( .A(n2651), .B(n2650), .Z(n2652) );
  AND U2834 ( .A(n2653), .B(n2652), .Z(n2689) );
  XOR U2835 ( .A(n2690), .B(n2689), .Z(c[184]) );
  NANDN U2836 ( .A(n2659), .B(n2658), .Z(n2663) );
  NAND U2837 ( .A(n2661), .B(n2660), .Z(n2662) );
  NAND U2838 ( .A(n2663), .B(n2662), .Z(n2724) );
  NANDN U2839 ( .A(n2665), .B(n2664), .Z(n2669) );
  NAND U2840 ( .A(n2667), .B(n2666), .Z(n2668) );
  NAND U2841 ( .A(n2669), .B(n2668), .Z(n2722) );
  XNOR U2842 ( .A(b[7]), .B(a[59]), .Z(n2709) );
  NANDN U2843 ( .A(n2709), .B(n5293), .Z(n2672) );
  NANDN U2844 ( .A(n2670), .B(n5294), .Z(n2671) );
  NAND U2845 ( .A(n2672), .B(n2671), .Z(n2697) );
  XNOR U2846 ( .A(b[3]), .B(a[63]), .Z(n2712) );
  NANDN U2847 ( .A(n2712), .B(n5160), .Z(n2675) );
  NANDN U2848 ( .A(n2673), .B(n5161), .Z(n2674) );
  AND U2849 ( .A(n2675), .B(n2674), .Z(n2698) );
  XNOR U2850 ( .A(n2697), .B(n2698), .Z(n2699) );
  NANDN U2851 ( .A(n292), .B(a[65]), .Z(n2676) );
  XOR U2852 ( .A(n5199), .B(n2676), .Z(n2678) );
  NANDN U2853 ( .A(b[0]), .B(a[64]), .Z(n2677) );
  AND U2854 ( .A(n2678), .B(n2677), .Z(n2705) );
  XNOR U2855 ( .A(b[5]), .B(a[61]), .Z(n2718) );
  NANDN U2856 ( .A(n2718), .B(n5240), .Z(n2681) );
  NANDN U2857 ( .A(n2679), .B(n5241), .Z(n2680) );
  NAND U2858 ( .A(n2681), .B(n2680), .Z(n2703) );
  NANDN U2859 ( .A(n295), .B(a[57]), .Z(n2704) );
  XNOR U2860 ( .A(n2703), .B(n2704), .Z(n2706) );
  XOR U2861 ( .A(n2705), .B(n2706), .Z(n2700) );
  XOR U2862 ( .A(n2699), .B(n2700), .Z(n2721) );
  XOR U2863 ( .A(n2722), .B(n2721), .Z(n2723) );
  XNOR U2864 ( .A(n2724), .B(n2723), .Z(n2693) );
  NAND U2865 ( .A(n2683), .B(n2682), .Z(n2687) );
  NAND U2866 ( .A(n2685), .B(n2684), .Z(n2686) );
  NAND U2867 ( .A(n2687), .B(n2686), .Z(n2694) );
  XNOR U2868 ( .A(n2693), .B(n2694), .Z(n2695) );
  XNOR U2869 ( .A(n2696), .B(n2695), .Z(n2727) );
  XNOR U2870 ( .A(n2727), .B(sreg[185]), .Z(n2729) );
  NAND U2871 ( .A(n2688), .B(sreg[184]), .Z(n2692) );
  OR U2872 ( .A(n2690), .B(n2689), .Z(n2691) );
  AND U2873 ( .A(n2692), .B(n2691), .Z(n2728) );
  XOR U2874 ( .A(n2729), .B(n2728), .Z(c[185]) );
  NANDN U2875 ( .A(n2698), .B(n2697), .Z(n2702) );
  NAND U2876 ( .A(n2700), .B(n2699), .Z(n2701) );
  NAND U2877 ( .A(n2702), .B(n2701), .Z(n2763) );
  NANDN U2878 ( .A(n2704), .B(n2703), .Z(n2708) );
  NAND U2879 ( .A(n2706), .B(n2705), .Z(n2707) );
  NAND U2880 ( .A(n2708), .B(n2707), .Z(n2761) );
  XNOR U2881 ( .A(b[7]), .B(a[60]), .Z(n2748) );
  NANDN U2882 ( .A(n2748), .B(n5293), .Z(n2711) );
  NANDN U2883 ( .A(n2709), .B(n5294), .Z(n2710) );
  NAND U2884 ( .A(n2711), .B(n2710), .Z(n2736) );
  XNOR U2885 ( .A(b[3]), .B(a[64]), .Z(n2751) );
  NANDN U2886 ( .A(n2751), .B(n5160), .Z(n2714) );
  NANDN U2887 ( .A(n2712), .B(n5161), .Z(n2713) );
  AND U2888 ( .A(n2714), .B(n2713), .Z(n2737) );
  XNOR U2889 ( .A(n2736), .B(n2737), .Z(n2738) );
  NANDN U2890 ( .A(n292), .B(a[66]), .Z(n2715) );
  XOR U2891 ( .A(n5199), .B(n2715), .Z(n2717) );
  NANDN U2892 ( .A(b[0]), .B(a[65]), .Z(n2716) );
  AND U2893 ( .A(n2717), .B(n2716), .Z(n2744) );
  XNOR U2894 ( .A(b[5]), .B(a[62]), .Z(n2757) );
  NANDN U2895 ( .A(n2757), .B(n5240), .Z(n2720) );
  NANDN U2896 ( .A(n2718), .B(n5241), .Z(n2719) );
  NAND U2897 ( .A(n2720), .B(n2719), .Z(n2742) );
  NANDN U2898 ( .A(n295), .B(a[58]), .Z(n2743) );
  XNOR U2899 ( .A(n2742), .B(n2743), .Z(n2745) );
  XOR U2900 ( .A(n2744), .B(n2745), .Z(n2739) );
  XOR U2901 ( .A(n2738), .B(n2739), .Z(n2760) );
  XOR U2902 ( .A(n2761), .B(n2760), .Z(n2762) );
  XNOR U2903 ( .A(n2763), .B(n2762), .Z(n2732) );
  NAND U2904 ( .A(n2722), .B(n2721), .Z(n2726) );
  NAND U2905 ( .A(n2724), .B(n2723), .Z(n2725) );
  NAND U2906 ( .A(n2726), .B(n2725), .Z(n2733) );
  XNOR U2907 ( .A(n2732), .B(n2733), .Z(n2734) );
  XNOR U2908 ( .A(n2735), .B(n2734), .Z(n2766) );
  XNOR U2909 ( .A(n2766), .B(sreg[186]), .Z(n2768) );
  NAND U2910 ( .A(n2727), .B(sreg[185]), .Z(n2731) );
  OR U2911 ( .A(n2729), .B(n2728), .Z(n2730) );
  AND U2912 ( .A(n2731), .B(n2730), .Z(n2767) );
  XOR U2913 ( .A(n2768), .B(n2767), .Z(c[186]) );
  NANDN U2914 ( .A(n2737), .B(n2736), .Z(n2741) );
  NAND U2915 ( .A(n2739), .B(n2738), .Z(n2740) );
  NAND U2916 ( .A(n2741), .B(n2740), .Z(n2802) );
  NANDN U2917 ( .A(n2743), .B(n2742), .Z(n2747) );
  NAND U2918 ( .A(n2745), .B(n2744), .Z(n2746) );
  NAND U2919 ( .A(n2747), .B(n2746), .Z(n2800) );
  XNOR U2920 ( .A(b[7]), .B(a[61]), .Z(n2787) );
  NANDN U2921 ( .A(n2787), .B(n5293), .Z(n2750) );
  NANDN U2922 ( .A(n2748), .B(n5294), .Z(n2749) );
  NAND U2923 ( .A(n2750), .B(n2749), .Z(n2775) );
  XNOR U2924 ( .A(b[3]), .B(a[65]), .Z(n2790) );
  NANDN U2925 ( .A(n2790), .B(n5160), .Z(n2753) );
  NANDN U2926 ( .A(n2751), .B(n5161), .Z(n2752) );
  AND U2927 ( .A(n2753), .B(n2752), .Z(n2776) );
  XNOR U2928 ( .A(n2775), .B(n2776), .Z(n2777) );
  NANDN U2929 ( .A(n292), .B(a[67]), .Z(n2754) );
  XOR U2930 ( .A(n5199), .B(n2754), .Z(n2756) );
  NANDN U2931 ( .A(b[0]), .B(a[66]), .Z(n2755) );
  AND U2932 ( .A(n2756), .B(n2755), .Z(n2783) );
  XNOR U2933 ( .A(b[5]), .B(a[63]), .Z(n2796) );
  NANDN U2934 ( .A(n2796), .B(n5240), .Z(n2759) );
  NANDN U2935 ( .A(n2757), .B(n5241), .Z(n2758) );
  NAND U2936 ( .A(n2759), .B(n2758), .Z(n2781) );
  NANDN U2937 ( .A(n295), .B(a[59]), .Z(n2782) );
  XNOR U2938 ( .A(n2781), .B(n2782), .Z(n2784) );
  XOR U2939 ( .A(n2783), .B(n2784), .Z(n2778) );
  XOR U2940 ( .A(n2777), .B(n2778), .Z(n2799) );
  XOR U2941 ( .A(n2800), .B(n2799), .Z(n2801) );
  XNOR U2942 ( .A(n2802), .B(n2801), .Z(n2771) );
  NAND U2943 ( .A(n2761), .B(n2760), .Z(n2765) );
  NAND U2944 ( .A(n2763), .B(n2762), .Z(n2764) );
  NAND U2945 ( .A(n2765), .B(n2764), .Z(n2772) );
  XNOR U2946 ( .A(n2771), .B(n2772), .Z(n2773) );
  XNOR U2947 ( .A(n2774), .B(n2773), .Z(n2805) );
  XNOR U2948 ( .A(n2805), .B(sreg[187]), .Z(n2807) );
  NAND U2949 ( .A(n2766), .B(sreg[186]), .Z(n2770) );
  OR U2950 ( .A(n2768), .B(n2767), .Z(n2769) );
  AND U2951 ( .A(n2770), .B(n2769), .Z(n2806) );
  XOR U2952 ( .A(n2807), .B(n2806), .Z(c[187]) );
  NANDN U2953 ( .A(n2776), .B(n2775), .Z(n2780) );
  NAND U2954 ( .A(n2778), .B(n2777), .Z(n2779) );
  NAND U2955 ( .A(n2780), .B(n2779), .Z(n2841) );
  NANDN U2956 ( .A(n2782), .B(n2781), .Z(n2786) );
  NAND U2957 ( .A(n2784), .B(n2783), .Z(n2785) );
  NAND U2958 ( .A(n2786), .B(n2785), .Z(n2839) );
  XNOR U2959 ( .A(b[7]), .B(a[62]), .Z(n2826) );
  NANDN U2960 ( .A(n2826), .B(n5293), .Z(n2789) );
  NANDN U2961 ( .A(n2787), .B(n5294), .Z(n2788) );
  NAND U2962 ( .A(n2789), .B(n2788), .Z(n2814) );
  XNOR U2963 ( .A(b[3]), .B(a[66]), .Z(n2829) );
  NANDN U2964 ( .A(n2829), .B(n5160), .Z(n2792) );
  NANDN U2965 ( .A(n2790), .B(n5161), .Z(n2791) );
  AND U2966 ( .A(n2792), .B(n2791), .Z(n2815) );
  XNOR U2967 ( .A(n2814), .B(n2815), .Z(n2816) );
  NANDN U2968 ( .A(n292), .B(a[68]), .Z(n2793) );
  XOR U2969 ( .A(n5199), .B(n2793), .Z(n2795) );
  NANDN U2970 ( .A(b[0]), .B(a[67]), .Z(n2794) );
  AND U2971 ( .A(n2795), .B(n2794), .Z(n2822) );
  XNOR U2972 ( .A(b[5]), .B(a[64]), .Z(n2835) );
  NANDN U2973 ( .A(n2835), .B(n5240), .Z(n2798) );
  NANDN U2974 ( .A(n2796), .B(n5241), .Z(n2797) );
  NAND U2975 ( .A(n2798), .B(n2797), .Z(n2820) );
  NANDN U2976 ( .A(n295), .B(a[60]), .Z(n2821) );
  XNOR U2977 ( .A(n2820), .B(n2821), .Z(n2823) );
  XOR U2978 ( .A(n2822), .B(n2823), .Z(n2817) );
  XOR U2979 ( .A(n2816), .B(n2817), .Z(n2838) );
  XOR U2980 ( .A(n2839), .B(n2838), .Z(n2840) );
  XNOR U2981 ( .A(n2841), .B(n2840), .Z(n2810) );
  NAND U2982 ( .A(n2800), .B(n2799), .Z(n2804) );
  NAND U2983 ( .A(n2802), .B(n2801), .Z(n2803) );
  NAND U2984 ( .A(n2804), .B(n2803), .Z(n2811) );
  XNOR U2985 ( .A(n2810), .B(n2811), .Z(n2812) );
  XNOR U2986 ( .A(n2813), .B(n2812), .Z(n2844) );
  XNOR U2987 ( .A(n2844), .B(sreg[188]), .Z(n2846) );
  NAND U2988 ( .A(n2805), .B(sreg[187]), .Z(n2809) );
  OR U2989 ( .A(n2807), .B(n2806), .Z(n2808) );
  AND U2990 ( .A(n2809), .B(n2808), .Z(n2845) );
  XOR U2991 ( .A(n2846), .B(n2845), .Z(c[188]) );
  NANDN U2992 ( .A(n2815), .B(n2814), .Z(n2819) );
  NAND U2993 ( .A(n2817), .B(n2816), .Z(n2818) );
  NAND U2994 ( .A(n2819), .B(n2818), .Z(n2880) );
  NANDN U2995 ( .A(n2821), .B(n2820), .Z(n2825) );
  NAND U2996 ( .A(n2823), .B(n2822), .Z(n2824) );
  NAND U2997 ( .A(n2825), .B(n2824), .Z(n2878) );
  XNOR U2998 ( .A(b[7]), .B(a[63]), .Z(n2865) );
  NANDN U2999 ( .A(n2865), .B(n5293), .Z(n2828) );
  NANDN U3000 ( .A(n2826), .B(n5294), .Z(n2827) );
  NAND U3001 ( .A(n2828), .B(n2827), .Z(n2853) );
  XNOR U3002 ( .A(b[3]), .B(a[67]), .Z(n2868) );
  NANDN U3003 ( .A(n2868), .B(n5160), .Z(n2831) );
  NANDN U3004 ( .A(n2829), .B(n5161), .Z(n2830) );
  AND U3005 ( .A(n2831), .B(n2830), .Z(n2854) );
  XNOR U3006 ( .A(n2853), .B(n2854), .Z(n2855) );
  NANDN U3007 ( .A(n292), .B(a[69]), .Z(n2832) );
  XOR U3008 ( .A(n5199), .B(n2832), .Z(n2834) );
  NANDN U3009 ( .A(b[0]), .B(a[68]), .Z(n2833) );
  AND U3010 ( .A(n2834), .B(n2833), .Z(n2861) );
  XNOR U3011 ( .A(b[5]), .B(a[65]), .Z(n2874) );
  NANDN U3012 ( .A(n2874), .B(n5240), .Z(n2837) );
  NANDN U3013 ( .A(n2835), .B(n5241), .Z(n2836) );
  NAND U3014 ( .A(n2837), .B(n2836), .Z(n2859) );
  NANDN U3015 ( .A(n295), .B(a[61]), .Z(n2860) );
  XNOR U3016 ( .A(n2859), .B(n2860), .Z(n2862) );
  XOR U3017 ( .A(n2861), .B(n2862), .Z(n2856) );
  XOR U3018 ( .A(n2855), .B(n2856), .Z(n2877) );
  XOR U3019 ( .A(n2878), .B(n2877), .Z(n2879) );
  XNOR U3020 ( .A(n2880), .B(n2879), .Z(n2849) );
  NAND U3021 ( .A(n2839), .B(n2838), .Z(n2843) );
  NAND U3022 ( .A(n2841), .B(n2840), .Z(n2842) );
  NAND U3023 ( .A(n2843), .B(n2842), .Z(n2850) );
  XNOR U3024 ( .A(n2849), .B(n2850), .Z(n2851) );
  XNOR U3025 ( .A(n2852), .B(n2851), .Z(n2883) );
  XNOR U3026 ( .A(n2883), .B(sreg[189]), .Z(n2885) );
  NAND U3027 ( .A(n2844), .B(sreg[188]), .Z(n2848) );
  OR U3028 ( .A(n2846), .B(n2845), .Z(n2847) );
  AND U3029 ( .A(n2848), .B(n2847), .Z(n2884) );
  XOR U3030 ( .A(n2885), .B(n2884), .Z(c[189]) );
  NANDN U3031 ( .A(n2854), .B(n2853), .Z(n2858) );
  NAND U3032 ( .A(n2856), .B(n2855), .Z(n2857) );
  NAND U3033 ( .A(n2858), .B(n2857), .Z(n2919) );
  NANDN U3034 ( .A(n2860), .B(n2859), .Z(n2864) );
  NAND U3035 ( .A(n2862), .B(n2861), .Z(n2863) );
  NAND U3036 ( .A(n2864), .B(n2863), .Z(n2917) );
  XNOR U3037 ( .A(b[7]), .B(a[64]), .Z(n2904) );
  NANDN U3038 ( .A(n2904), .B(n5293), .Z(n2867) );
  NANDN U3039 ( .A(n2865), .B(n5294), .Z(n2866) );
  NAND U3040 ( .A(n2867), .B(n2866), .Z(n2892) );
  XNOR U3041 ( .A(b[3]), .B(a[68]), .Z(n2907) );
  NANDN U3042 ( .A(n2907), .B(n5160), .Z(n2870) );
  NANDN U3043 ( .A(n2868), .B(n5161), .Z(n2869) );
  AND U3044 ( .A(n2870), .B(n2869), .Z(n2893) );
  XNOR U3045 ( .A(n2892), .B(n2893), .Z(n2894) );
  NANDN U3046 ( .A(n292), .B(a[70]), .Z(n2871) );
  XOR U3047 ( .A(n5199), .B(n2871), .Z(n2873) );
  NANDN U3048 ( .A(b[0]), .B(a[69]), .Z(n2872) );
  AND U3049 ( .A(n2873), .B(n2872), .Z(n2900) );
  XNOR U3050 ( .A(b[5]), .B(a[66]), .Z(n2913) );
  NANDN U3051 ( .A(n2913), .B(n5240), .Z(n2876) );
  NANDN U3052 ( .A(n2874), .B(n5241), .Z(n2875) );
  NAND U3053 ( .A(n2876), .B(n2875), .Z(n2898) );
  NANDN U3054 ( .A(n295), .B(a[62]), .Z(n2899) );
  XNOR U3055 ( .A(n2898), .B(n2899), .Z(n2901) );
  XOR U3056 ( .A(n2900), .B(n2901), .Z(n2895) );
  XOR U3057 ( .A(n2894), .B(n2895), .Z(n2916) );
  XOR U3058 ( .A(n2917), .B(n2916), .Z(n2918) );
  XNOR U3059 ( .A(n2919), .B(n2918), .Z(n2888) );
  NAND U3060 ( .A(n2878), .B(n2877), .Z(n2882) );
  NAND U3061 ( .A(n2880), .B(n2879), .Z(n2881) );
  NAND U3062 ( .A(n2882), .B(n2881), .Z(n2889) );
  XNOR U3063 ( .A(n2888), .B(n2889), .Z(n2890) );
  XNOR U3064 ( .A(n2891), .B(n2890), .Z(n2922) );
  XNOR U3065 ( .A(n2922), .B(sreg[190]), .Z(n2924) );
  NAND U3066 ( .A(n2883), .B(sreg[189]), .Z(n2887) );
  OR U3067 ( .A(n2885), .B(n2884), .Z(n2886) );
  AND U3068 ( .A(n2887), .B(n2886), .Z(n2923) );
  XOR U3069 ( .A(n2924), .B(n2923), .Z(c[190]) );
  NANDN U3070 ( .A(n2893), .B(n2892), .Z(n2897) );
  NAND U3071 ( .A(n2895), .B(n2894), .Z(n2896) );
  NAND U3072 ( .A(n2897), .B(n2896), .Z(n2958) );
  NANDN U3073 ( .A(n2899), .B(n2898), .Z(n2903) );
  NAND U3074 ( .A(n2901), .B(n2900), .Z(n2902) );
  NAND U3075 ( .A(n2903), .B(n2902), .Z(n2956) );
  XNOR U3076 ( .A(b[7]), .B(a[65]), .Z(n2949) );
  NANDN U3077 ( .A(n2949), .B(n5293), .Z(n2906) );
  NANDN U3078 ( .A(n2904), .B(n5294), .Z(n2905) );
  NAND U3079 ( .A(n2906), .B(n2905), .Z(n2931) );
  XNOR U3080 ( .A(b[3]), .B(a[69]), .Z(n2952) );
  NANDN U3081 ( .A(n2952), .B(n5160), .Z(n2909) );
  NANDN U3082 ( .A(n2907), .B(n5161), .Z(n2908) );
  AND U3083 ( .A(n2909), .B(n2908), .Z(n2932) );
  XNOR U3084 ( .A(n2931), .B(n2932), .Z(n2933) );
  NANDN U3085 ( .A(n292), .B(a[71]), .Z(n2910) );
  XOR U3086 ( .A(n5199), .B(n2910), .Z(n2912) );
  NANDN U3087 ( .A(b[0]), .B(a[70]), .Z(n2911) );
  AND U3088 ( .A(n2912), .B(n2911), .Z(n2939) );
  XNOR U3089 ( .A(b[5]), .B(a[67]), .Z(n2946) );
  NANDN U3090 ( .A(n2946), .B(n5240), .Z(n2915) );
  NANDN U3091 ( .A(n2913), .B(n5241), .Z(n2914) );
  NAND U3092 ( .A(n2915), .B(n2914), .Z(n2937) );
  NANDN U3093 ( .A(n295), .B(a[63]), .Z(n2938) );
  XNOR U3094 ( .A(n2937), .B(n2938), .Z(n2940) );
  XOR U3095 ( .A(n2939), .B(n2940), .Z(n2934) );
  XOR U3096 ( .A(n2933), .B(n2934), .Z(n2955) );
  XOR U3097 ( .A(n2956), .B(n2955), .Z(n2957) );
  XNOR U3098 ( .A(n2958), .B(n2957), .Z(n2927) );
  NAND U3099 ( .A(n2917), .B(n2916), .Z(n2921) );
  NAND U3100 ( .A(n2919), .B(n2918), .Z(n2920) );
  NAND U3101 ( .A(n2921), .B(n2920), .Z(n2928) );
  XNOR U3102 ( .A(n2927), .B(n2928), .Z(n2929) );
  XNOR U3103 ( .A(n2930), .B(n2929), .Z(n2961) );
  XNOR U3104 ( .A(n2961), .B(sreg[191]), .Z(n2963) );
  NAND U3105 ( .A(n2922), .B(sreg[190]), .Z(n2926) );
  OR U3106 ( .A(n2924), .B(n2923), .Z(n2925) );
  AND U3107 ( .A(n2926), .B(n2925), .Z(n2962) );
  XOR U3108 ( .A(n2963), .B(n2962), .Z(c[191]) );
  NANDN U3109 ( .A(n2932), .B(n2931), .Z(n2936) );
  NAND U3110 ( .A(n2934), .B(n2933), .Z(n2935) );
  NAND U3111 ( .A(n2936), .B(n2935), .Z(n2997) );
  NANDN U3112 ( .A(n2938), .B(n2937), .Z(n2942) );
  NAND U3113 ( .A(n2940), .B(n2939), .Z(n2941) );
  NAND U3114 ( .A(n2942), .B(n2941), .Z(n2995) );
  NANDN U3115 ( .A(n292), .B(a[72]), .Z(n2943) );
  XOR U3116 ( .A(n5199), .B(n2943), .Z(n2945) );
  NANDN U3117 ( .A(b[0]), .B(a[71]), .Z(n2944) );
  AND U3118 ( .A(n2945), .B(n2944), .Z(n2978) );
  XNOR U3119 ( .A(b[5]), .B(a[68]), .Z(n2991) );
  NANDN U3120 ( .A(n2991), .B(n5240), .Z(n2948) );
  NANDN U3121 ( .A(n2946), .B(n5241), .Z(n2947) );
  NAND U3122 ( .A(n2948), .B(n2947), .Z(n2976) );
  NANDN U3123 ( .A(n295), .B(a[64]), .Z(n2977) );
  XNOR U3124 ( .A(n2976), .B(n2977), .Z(n2979) );
  XOR U3125 ( .A(n2978), .B(n2979), .Z(n2972) );
  XNOR U3126 ( .A(b[7]), .B(a[66]), .Z(n2982) );
  NANDN U3127 ( .A(n2982), .B(n5293), .Z(n2951) );
  NANDN U3128 ( .A(n2949), .B(n5294), .Z(n2950) );
  NAND U3129 ( .A(n2951), .B(n2950), .Z(n2970) );
  XNOR U3130 ( .A(b[3]), .B(a[70]), .Z(n2985) );
  NANDN U3131 ( .A(n2985), .B(n5160), .Z(n2954) );
  NANDN U3132 ( .A(n2952), .B(n5161), .Z(n2953) );
  AND U3133 ( .A(n2954), .B(n2953), .Z(n2971) );
  XNOR U3134 ( .A(n2970), .B(n2971), .Z(n2973) );
  XOR U3135 ( .A(n2972), .B(n2973), .Z(n2994) );
  XOR U3136 ( .A(n2995), .B(n2994), .Z(n2996) );
  XNOR U3137 ( .A(n2997), .B(n2996), .Z(n2966) );
  NAND U3138 ( .A(n2956), .B(n2955), .Z(n2960) );
  NAND U3139 ( .A(n2958), .B(n2957), .Z(n2959) );
  NAND U3140 ( .A(n2960), .B(n2959), .Z(n2967) );
  XNOR U3141 ( .A(n2966), .B(n2967), .Z(n2968) );
  XNOR U3142 ( .A(n2969), .B(n2968), .Z(n3000) );
  XNOR U3143 ( .A(n3000), .B(sreg[192]), .Z(n3002) );
  NAND U3144 ( .A(n2961), .B(sreg[191]), .Z(n2965) );
  OR U3145 ( .A(n2963), .B(n2962), .Z(n2964) );
  AND U3146 ( .A(n2965), .B(n2964), .Z(n3001) );
  XOR U3147 ( .A(n3002), .B(n3001), .Z(c[192]) );
  NANDN U3148 ( .A(n2971), .B(n2970), .Z(n2975) );
  NAND U3149 ( .A(n2973), .B(n2972), .Z(n2974) );
  NAND U3150 ( .A(n2975), .B(n2974), .Z(n3036) );
  NANDN U3151 ( .A(n2977), .B(n2976), .Z(n2981) );
  NAND U3152 ( .A(n2979), .B(n2978), .Z(n2980) );
  NAND U3153 ( .A(n2981), .B(n2980), .Z(n3034) );
  XNOR U3154 ( .A(b[7]), .B(a[67]), .Z(n3021) );
  NANDN U3155 ( .A(n3021), .B(n5293), .Z(n2984) );
  NANDN U3156 ( .A(n2982), .B(n5294), .Z(n2983) );
  NAND U3157 ( .A(n2984), .B(n2983), .Z(n3009) );
  XNOR U3158 ( .A(b[3]), .B(a[71]), .Z(n3024) );
  NANDN U3159 ( .A(n3024), .B(n5160), .Z(n2987) );
  NANDN U3160 ( .A(n2985), .B(n5161), .Z(n2986) );
  AND U3161 ( .A(n2987), .B(n2986), .Z(n3010) );
  XNOR U3162 ( .A(n3009), .B(n3010), .Z(n3011) );
  NANDN U3163 ( .A(n292), .B(a[73]), .Z(n2988) );
  XOR U3164 ( .A(n5199), .B(n2988), .Z(n2990) );
  NANDN U3165 ( .A(b[0]), .B(a[72]), .Z(n2989) );
  AND U3166 ( .A(n2990), .B(n2989), .Z(n3017) );
  XNOR U3167 ( .A(b[5]), .B(a[69]), .Z(n3030) );
  NANDN U3168 ( .A(n3030), .B(n5240), .Z(n2993) );
  NANDN U3169 ( .A(n2991), .B(n5241), .Z(n2992) );
  NAND U3170 ( .A(n2993), .B(n2992), .Z(n3015) );
  NANDN U3171 ( .A(n295), .B(a[65]), .Z(n3016) );
  XNOR U3172 ( .A(n3015), .B(n3016), .Z(n3018) );
  XOR U3173 ( .A(n3017), .B(n3018), .Z(n3012) );
  XOR U3174 ( .A(n3011), .B(n3012), .Z(n3033) );
  XOR U3175 ( .A(n3034), .B(n3033), .Z(n3035) );
  XNOR U3176 ( .A(n3036), .B(n3035), .Z(n3005) );
  NAND U3177 ( .A(n2995), .B(n2994), .Z(n2999) );
  NAND U3178 ( .A(n2997), .B(n2996), .Z(n2998) );
  NAND U3179 ( .A(n2999), .B(n2998), .Z(n3006) );
  XNOR U3180 ( .A(n3005), .B(n3006), .Z(n3007) );
  XNOR U3181 ( .A(n3008), .B(n3007), .Z(n3039) );
  XNOR U3182 ( .A(n3039), .B(sreg[193]), .Z(n3041) );
  NAND U3183 ( .A(n3000), .B(sreg[192]), .Z(n3004) );
  OR U3184 ( .A(n3002), .B(n3001), .Z(n3003) );
  AND U3185 ( .A(n3004), .B(n3003), .Z(n3040) );
  XOR U3186 ( .A(n3041), .B(n3040), .Z(c[193]) );
  NANDN U3187 ( .A(n3010), .B(n3009), .Z(n3014) );
  NAND U3188 ( .A(n3012), .B(n3011), .Z(n3013) );
  NAND U3189 ( .A(n3014), .B(n3013), .Z(n3075) );
  NANDN U3190 ( .A(n3016), .B(n3015), .Z(n3020) );
  NAND U3191 ( .A(n3018), .B(n3017), .Z(n3019) );
  NAND U3192 ( .A(n3020), .B(n3019), .Z(n3073) );
  XNOR U3193 ( .A(b[7]), .B(a[68]), .Z(n3060) );
  NANDN U3194 ( .A(n3060), .B(n5293), .Z(n3023) );
  NANDN U3195 ( .A(n3021), .B(n5294), .Z(n3022) );
  NAND U3196 ( .A(n3023), .B(n3022), .Z(n3048) );
  XNOR U3197 ( .A(b[3]), .B(a[72]), .Z(n3063) );
  NANDN U3198 ( .A(n3063), .B(n5160), .Z(n3026) );
  NANDN U3199 ( .A(n3024), .B(n5161), .Z(n3025) );
  AND U3200 ( .A(n3026), .B(n3025), .Z(n3049) );
  XNOR U3201 ( .A(n3048), .B(n3049), .Z(n3050) );
  NANDN U3202 ( .A(n292), .B(a[74]), .Z(n3027) );
  XOR U3203 ( .A(n5199), .B(n3027), .Z(n3029) );
  NANDN U3204 ( .A(b[0]), .B(a[73]), .Z(n3028) );
  AND U3205 ( .A(n3029), .B(n3028), .Z(n3056) );
  XNOR U3206 ( .A(b[5]), .B(a[70]), .Z(n3069) );
  NANDN U3207 ( .A(n3069), .B(n5240), .Z(n3032) );
  NANDN U3208 ( .A(n3030), .B(n5241), .Z(n3031) );
  NAND U3209 ( .A(n3032), .B(n3031), .Z(n3054) );
  NANDN U3210 ( .A(n295), .B(a[66]), .Z(n3055) );
  XNOR U3211 ( .A(n3054), .B(n3055), .Z(n3057) );
  XOR U3212 ( .A(n3056), .B(n3057), .Z(n3051) );
  XOR U3213 ( .A(n3050), .B(n3051), .Z(n3072) );
  XOR U3214 ( .A(n3073), .B(n3072), .Z(n3074) );
  XNOR U3215 ( .A(n3075), .B(n3074), .Z(n3044) );
  NAND U3216 ( .A(n3034), .B(n3033), .Z(n3038) );
  NAND U3217 ( .A(n3036), .B(n3035), .Z(n3037) );
  NAND U3218 ( .A(n3038), .B(n3037), .Z(n3045) );
  XNOR U3219 ( .A(n3044), .B(n3045), .Z(n3046) );
  XNOR U3220 ( .A(n3047), .B(n3046), .Z(n3078) );
  XNOR U3221 ( .A(n3078), .B(sreg[194]), .Z(n3080) );
  NAND U3222 ( .A(n3039), .B(sreg[193]), .Z(n3043) );
  OR U3223 ( .A(n3041), .B(n3040), .Z(n3042) );
  AND U3224 ( .A(n3043), .B(n3042), .Z(n3079) );
  XOR U3225 ( .A(n3080), .B(n3079), .Z(c[194]) );
  NANDN U3226 ( .A(n3049), .B(n3048), .Z(n3053) );
  NAND U3227 ( .A(n3051), .B(n3050), .Z(n3052) );
  NAND U3228 ( .A(n3053), .B(n3052), .Z(n3114) );
  NANDN U3229 ( .A(n3055), .B(n3054), .Z(n3059) );
  NAND U3230 ( .A(n3057), .B(n3056), .Z(n3058) );
  NAND U3231 ( .A(n3059), .B(n3058), .Z(n3112) );
  XNOR U3232 ( .A(b[7]), .B(a[69]), .Z(n3099) );
  NANDN U3233 ( .A(n3099), .B(n5293), .Z(n3062) );
  NANDN U3234 ( .A(n3060), .B(n5294), .Z(n3061) );
  NAND U3235 ( .A(n3062), .B(n3061), .Z(n3087) );
  XNOR U3236 ( .A(b[3]), .B(a[73]), .Z(n3102) );
  NANDN U3237 ( .A(n3102), .B(n5160), .Z(n3065) );
  NANDN U3238 ( .A(n3063), .B(n5161), .Z(n3064) );
  AND U3239 ( .A(n3065), .B(n3064), .Z(n3088) );
  XNOR U3240 ( .A(n3087), .B(n3088), .Z(n3089) );
  NANDN U3241 ( .A(n292), .B(a[75]), .Z(n3066) );
  XOR U3242 ( .A(n5199), .B(n3066), .Z(n3068) );
  NANDN U3243 ( .A(b[0]), .B(a[74]), .Z(n3067) );
  AND U3244 ( .A(n3068), .B(n3067), .Z(n3095) );
  XNOR U3245 ( .A(b[5]), .B(a[71]), .Z(n3108) );
  NANDN U3246 ( .A(n3108), .B(n5240), .Z(n3071) );
  NANDN U3247 ( .A(n3069), .B(n5241), .Z(n3070) );
  NAND U3248 ( .A(n3071), .B(n3070), .Z(n3093) );
  NANDN U3249 ( .A(n295), .B(a[67]), .Z(n3094) );
  XNOR U3250 ( .A(n3093), .B(n3094), .Z(n3096) );
  XOR U3251 ( .A(n3095), .B(n3096), .Z(n3090) );
  XOR U3252 ( .A(n3089), .B(n3090), .Z(n3111) );
  XOR U3253 ( .A(n3112), .B(n3111), .Z(n3113) );
  XNOR U3254 ( .A(n3114), .B(n3113), .Z(n3083) );
  NAND U3255 ( .A(n3073), .B(n3072), .Z(n3077) );
  NAND U3256 ( .A(n3075), .B(n3074), .Z(n3076) );
  NAND U3257 ( .A(n3077), .B(n3076), .Z(n3084) );
  XNOR U3258 ( .A(n3083), .B(n3084), .Z(n3085) );
  XNOR U3259 ( .A(n3086), .B(n3085), .Z(n3117) );
  XNOR U3260 ( .A(n3117), .B(sreg[195]), .Z(n3119) );
  NAND U3261 ( .A(n3078), .B(sreg[194]), .Z(n3082) );
  OR U3262 ( .A(n3080), .B(n3079), .Z(n3081) );
  AND U3263 ( .A(n3082), .B(n3081), .Z(n3118) );
  XOR U3264 ( .A(n3119), .B(n3118), .Z(c[195]) );
  NANDN U3265 ( .A(n3088), .B(n3087), .Z(n3092) );
  NAND U3266 ( .A(n3090), .B(n3089), .Z(n3091) );
  NAND U3267 ( .A(n3092), .B(n3091), .Z(n3153) );
  NANDN U3268 ( .A(n3094), .B(n3093), .Z(n3098) );
  NAND U3269 ( .A(n3096), .B(n3095), .Z(n3097) );
  NAND U3270 ( .A(n3098), .B(n3097), .Z(n3151) );
  XNOR U3271 ( .A(b[7]), .B(a[70]), .Z(n3138) );
  NANDN U3272 ( .A(n3138), .B(n5293), .Z(n3101) );
  NANDN U3273 ( .A(n3099), .B(n5294), .Z(n3100) );
  NAND U3274 ( .A(n3101), .B(n3100), .Z(n3126) );
  XNOR U3275 ( .A(b[3]), .B(a[74]), .Z(n3141) );
  NANDN U3276 ( .A(n3141), .B(n5160), .Z(n3104) );
  NANDN U3277 ( .A(n3102), .B(n5161), .Z(n3103) );
  AND U3278 ( .A(n3104), .B(n3103), .Z(n3127) );
  XNOR U3279 ( .A(n3126), .B(n3127), .Z(n3128) );
  NANDN U3280 ( .A(n292), .B(a[76]), .Z(n3105) );
  XOR U3281 ( .A(n5199), .B(n3105), .Z(n3107) );
  NANDN U3282 ( .A(b[0]), .B(a[75]), .Z(n3106) );
  AND U3283 ( .A(n3107), .B(n3106), .Z(n3134) );
  XNOR U3284 ( .A(b[5]), .B(a[72]), .Z(n3147) );
  NANDN U3285 ( .A(n3147), .B(n5240), .Z(n3110) );
  NANDN U3286 ( .A(n3108), .B(n5241), .Z(n3109) );
  NAND U3287 ( .A(n3110), .B(n3109), .Z(n3132) );
  NANDN U3288 ( .A(n295), .B(a[68]), .Z(n3133) );
  XNOR U3289 ( .A(n3132), .B(n3133), .Z(n3135) );
  XOR U3290 ( .A(n3134), .B(n3135), .Z(n3129) );
  XOR U3291 ( .A(n3128), .B(n3129), .Z(n3150) );
  XOR U3292 ( .A(n3151), .B(n3150), .Z(n3152) );
  XNOR U3293 ( .A(n3153), .B(n3152), .Z(n3122) );
  NAND U3294 ( .A(n3112), .B(n3111), .Z(n3116) );
  NAND U3295 ( .A(n3114), .B(n3113), .Z(n3115) );
  NAND U3296 ( .A(n3116), .B(n3115), .Z(n3123) );
  XNOR U3297 ( .A(n3122), .B(n3123), .Z(n3124) );
  XNOR U3298 ( .A(n3125), .B(n3124), .Z(n3156) );
  XNOR U3299 ( .A(n3156), .B(sreg[196]), .Z(n3158) );
  NAND U3300 ( .A(n3117), .B(sreg[195]), .Z(n3121) );
  OR U3301 ( .A(n3119), .B(n3118), .Z(n3120) );
  AND U3302 ( .A(n3121), .B(n3120), .Z(n3157) );
  XOR U3303 ( .A(n3158), .B(n3157), .Z(c[196]) );
  NANDN U3304 ( .A(n3127), .B(n3126), .Z(n3131) );
  NAND U3305 ( .A(n3129), .B(n3128), .Z(n3130) );
  NAND U3306 ( .A(n3131), .B(n3130), .Z(n3192) );
  NANDN U3307 ( .A(n3133), .B(n3132), .Z(n3137) );
  NAND U3308 ( .A(n3135), .B(n3134), .Z(n3136) );
  NAND U3309 ( .A(n3137), .B(n3136), .Z(n3190) );
  XNOR U3310 ( .A(b[7]), .B(a[71]), .Z(n3177) );
  NANDN U3311 ( .A(n3177), .B(n5293), .Z(n3140) );
  NANDN U3312 ( .A(n3138), .B(n5294), .Z(n3139) );
  NAND U3313 ( .A(n3140), .B(n3139), .Z(n3165) );
  XNOR U3314 ( .A(b[3]), .B(a[75]), .Z(n3180) );
  NANDN U3315 ( .A(n3180), .B(n5160), .Z(n3143) );
  NANDN U3316 ( .A(n3141), .B(n5161), .Z(n3142) );
  AND U3317 ( .A(n3143), .B(n3142), .Z(n3166) );
  XNOR U3318 ( .A(n3165), .B(n3166), .Z(n3167) );
  NANDN U3319 ( .A(n292), .B(a[77]), .Z(n3144) );
  XOR U3320 ( .A(n5199), .B(n3144), .Z(n3146) );
  NANDN U3321 ( .A(b[0]), .B(a[76]), .Z(n3145) );
  AND U3322 ( .A(n3146), .B(n3145), .Z(n3173) );
  XNOR U3323 ( .A(n294), .B(a[73]), .Z(n3186) );
  NAND U3324 ( .A(n3186), .B(n5240), .Z(n3149) );
  NANDN U3325 ( .A(n3147), .B(n5241), .Z(n3148) );
  NAND U3326 ( .A(n3149), .B(n3148), .Z(n3171) );
  NANDN U3327 ( .A(n295), .B(a[69]), .Z(n3172) );
  XNOR U3328 ( .A(n3171), .B(n3172), .Z(n3174) );
  XOR U3329 ( .A(n3173), .B(n3174), .Z(n3168) );
  XOR U3330 ( .A(n3167), .B(n3168), .Z(n3189) );
  XOR U3331 ( .A(n3190), .B(n3189), .Z(n3191) );
  XNOR U3332 ( .A(n3192), .B(n3191), .Z(n3161) );
  NAND U3333 ( .A(n3151), .B(n3150), .Z(n3155) );
  NAND U3334 ( .A(n3153), .B(n3152), .Z(n3154) );
  NAND U3335 ( .A(n3155), .B(n3154), .Z(n3162) );
  XNOR U3336 ( .A(n3161), .B(n3162), .Z(n3163) );
  XNOR U3337 ( .A(n3164), .B(n3163), .Z(n3195) );
  XNOR U3338 ( .A(n3195), .B(sreg[197]), .Z(n3197) );
  NAND U3339 ( .A(n3156), .B(sreg[196]), .Z(n3160) );
  OR U3340 ( .A(n3158), .B(n3157), .Z(n3159) );
  AND U3341 ( .A(n3160), .B(n3159), .Z(n3196) );
  XOR U3342 ( .A(n3197), .B(n3196), .Z(c[197]) );
  NANDN U3343 ( .A(n3166), .B(n3165), .Z(n3170) );
  NAND U3344 ( .A(n3168), .B(n3167), .Z(n3169) );
  NAND U3345 ( .A(n3170), .B(n3169), .Z(n3231) );
  NANDN U3346 ( .A(n3172), .B(n3171), .Z(n3176) );
  NAND U3347 ( .A(n3174), .B(n3173), .Z(n3175) );
  NAND U3348 ( .A(n3176), .B(n3175), .Z(n3229) );
  XNOR U3349 ( .A(b[7]), .B(a[72]), .Z(n3204) );
  NANDN U3350 ( .A(n3204), .B(n5293), .Z(n3179) );
  NANDN U3351 ( .A(n3177), .B(n5294), .Z(n3178) );
  NAND U3352 ( .A(n3179), .B(n3178), .Z(n3216) );
  XNOR U3353 ( .A(b[3]), .B(a[76]), .Z(n3207) );
  NANDN U3354 ( .A(n3207), .B(n5160), .Z(n3182) );
  NANDN U3355 ( .A(n3180), .B(n5161), .Z(n3181) );
  AND U3356 ( .A(n3182), .B(n3181), .Z(n3217) );
  XNOR U3357 ( .A(n3216), .B(n3217), .Z(n3218) );
  NANDN U3358 ( .A(n292), .B(a[78]), .Z(n3183) );
  XOR U3359 ( .A(n5199), .B(n3183), .Z(n3185) );
  NANDN U3360 ( .A(b[0]), .B(a[77]), .Z(n3184) );
  AND U3361 ( .A(n3185), .B(n3184), .Z(n3224) );
  XNOR U3362 ( .A(b[5]), .B(a[74]), .Z(n3213) );
  NANDN U3363 ( .A(n3213), .B(n5240), .Z(n3188) );
  NAND U3364 ( .A(n5241), .B(n3186), .Z(n3187) );
  AND U3365 ( .A(n3188), .B(n3187), .Z(n3222) );
  NANDN U3366 ( .A(n295), .B(a[70]), .Z(n3223) );
  XOR U3367 ( .A(n3222), .B(n3223), .Z(n3225) );
  XNOR U3368 ( .A(n3224), .B(n3225), .Z(n3219) );
  XNOR U3369 ( .A(n3218), .B(n3219), .Z(n3228) );
  XOR U3370 ( .A(n3229), .B(n3228), .Z(n3230) );
  XNOR U3371 ( .A(n3231), .B(n3230), .Z(n3200) );
  NAND U3372 ( .A(n3190), .B(n3189), .Z(n3194) );
  NAND U3373 ( .A(n3192), .B(n3191), .Z(n3193) );
  NAND U3374 ( .A(n3194), .B(n3193), .Z(n3201) );
  XNOR U3375 ( .A(n3200), .B(n3201), .Z(n3202) );
  XNOR U3376 ( .A(n3203), .B(n3202), .Z(n3232) );
  XNOR U3377 ( .A(n3232), .B(sreg[198]), .Z(n3234) );
  NAND U3378 ( .A(n3195), .B(sreg[197]), .Z(n3199) );
  OR U3379 ( .A(n3197), .B(n3196), .Z(n3198) );
  AND U3380 ( .A(n3199), .B(n3198), .Z(n3233) );
  XOR U3381 ( .A(n3234), .B(n3233), .Z(c[198]) );
  XNOR U3382 ( .A(b[7]), .B(a[73]), .Z(n3253) );
  NANDN U3383 ( .A(n3253), .B(n5293), .Z(n3206) );
  NANDN U3384 ( .A(n3204), .B(n5294), .Z(n3205) );
  NAND U3385 ( .A(n3206), .B(n3205), .Z(n3241) );
  XNOR U3386 ( .A(b[3]), .B(a[77]), .Z(n3256) );
  NANDN U3387 ( .A(n3256), .B(n5160), .Z(n3209) );
  NANDN U3388 ( .A(n3207), .B(n5161), .Z(n3208) );
  AND U3389 ( .A(n3209), .B(n3208), .Z(n3242) );
  XNOR U3390 ( .A(n3241), .B(n3242), .Z(n3243) );
  NANDN U3391 ( .A(n292), .B(a[79]), .Z(n3210) );
  XOR U3392 ( .A(n5199), .B(n3210), .Z(n3212) );
  NANDN U3393 ( .A(b[0]), .B(a[78]), .Z(n3211) );
  AND U3394 ( .A(n3212), .B(n3211), .Z(n3249) );
  XNOR U3395 ( .A(b[5]), .B(a[75]), .Z(n3262) );
  NANDN U3396 ( .A(n3262), .B(n5240), .Z(n3215) );
  NANDN U3397 ( .A(n3213), .B(n5241), .Z(n3214) );
  NAND U3398 ( .A(n3215), .B(n3214), .Z(n3247) );
  NANDN U3399 ( .A(n295), .B(a[71]), .Z(n3248) );
  XNOR U3400 ( .A(n3247), .B(n3248), .Z(n3250) );
  XOR U3401 ( .A(n3249), .B(n3250), .Z(n3244) );
  XOR U3402 ( .A(n3243), .B(n3244), .Z(n3267) );
  NANDN U3403 ( .A(n3217), .B(n3216), .Z(n3221) );
  NANDN U3404 ( .A(n3219), .B(n3218), .Z(n3220) );
  NAND U3405 ( .A(n3221), .B(n3220), .Z(n3265) );
  OR U3406 ( .A(n3223), .B(n3222), .Z(n3227) );
  NAND U3407 ( .A(n3225), .B(n3224), .Z(n3226) );
  AND U3408 ( .A(n3227), .B(n3226), .Z(n3266) );
  XNOR U3409 ( .A(n3265), .B(n3266), .Z(n3268) );
  XNOR U3410 ( .A(n3267), .B(n3268), .Z(n3237) );
  XNOR U3411 ( .A(n3237), .B(n3238), .Z(n3239) );
  XNOR U3412 ( .A(n3240), .B(n3239), .Z(n3271) );
  XNOR U3413 ( .A(n3271), .B(sreg[199]), .Z(n3273) );
  NAND U3414 ( .A(n3232), .B(sreg[198]), .Z(n3236) );
  OR U3415 ( .A(n3234), .B(n3233), .Z(n3235) );
  AND U3416 ( .A(n3236), .B(n3235), .Z(n3272) );
  XOR U3417 ( .A(n3273), .B(n3272), .Z(c[199]) );
  NANDN U3418 ( .A(n3242), .B(n3241), .Z(n3246) );
  NAND U3419 ( .A(n3244), .B(n3243), .Z(n3245) );
  NAND U3420 ( .A(n3246), .B(n3245), .Z(n3307) );
  NANDN U3421 ( .A(n3248), .B(n3247), .Z(n3252) );
  NAND U3422 ( .A(n3250), .B(n3249), .Z(n3251) );
  NAND U3423 ( .A(n3252), .B(n3251), .Z(n3305) );
  XNOR U3424 ( .A(b[7]), .B(a[74]), .Z(n3292) );
  NANDN U3425 ( .A(n3292), .B(n5293), .Z(n3255) );
  NANDN U3426 ( .A(n3253), .B(n5294), .Z(n3254) );
  NAND U3427 ( .A(n3255), .B(n3254), .Z(n3280) );
  XNOR U3428 ( .A(b[3]), .B(a[78]), .Z(n3295) );
  NANDN U3429 ( .A(n3295), .B(n5160), .Z(n3258) );
  NANDN U3430 ( .A(n3256), .B(n5161), .Z(n3257) );
  AND U3431 ( .A(n3258), .B(n3257), .Z(n3281) );
  XNOR U3432 ( .A(n3280), .B(n3281), .Z(n3282) );
  NANDN U3433 ( .A(n292), .B(a[80]), .Z(n3259) );
  XOR U3434 ( .A(n5199), .B(n3259), .Z(n3261) );
  NANDN U3435 ( .A(b[0]), .B(a[79]), .Z(n3260) );
  AND U3436 ( .A(n3261), .B(n3260), .Z(n3288) );
  XNOR U3437 ( .A(b[5]), .B(a[76]), .Z(n3301) );
  NANDN U3438 ( .A(n3301), .B(n5240), .Z(n3264) );
  NANDN U3439 ( .A(n3262), .B(n5241), .Z(n3263) );
  NAND U3440 ( .A(n3264), .B(n3263), .Z(n3286) );
  NANDN U3441 ( .A(n295), .B(a[72]), .Z(n3287) );
  XNOR U3442 ( .A(n3286), .B(n3287), .Z(n3289) );
  XOR U3443 ( .A(n3288), .B(n3289), .Z(n3283) );
  XOR U3444 ( .A(n3282), .B(n3283), .Z(n3304) );
  XOR U3445 ( .A(n3305), .B(n3304), .Z(n3306) );
  XNOR U3446 ( .A(n3307), .B(n3306), .Z(n3276) );
  NANDN U3447 ( .A(n3266), .B(n3265), .Z(n3270) );
  NAND U3448 ( .A(n3268), .B(n3267), .Z(n3269) );
  NAND U3449 ( .A(n3270), .B(n3269), .Z(n3277) );
  XNOR U3450 ( .A(n3276), .B(n3277), .Z(n3278) );
  XNOR U3451 ( .A(n3279), .B(n3278), .Z(n3310) );
  XNOR U3452 ( .A(n3310), .B(sreg[200]), .Z(n3312) );
  NAND U3453 ( .A(n3271), .B(sreg[199]), .Z(n3275) );
  OR U3454 ( .A(n3273), .B(n3272), .Z(n3274) );
  AND U3455 ( .A(n3275), .B(n3274), .Z(n3311) );
  XOR U3456 ( .A(n3312), .B(n3311), .Z(c[200]) );
  NANDN U3457 ( .A(n3281), .B(n3280), .Z(n3285) );
  NAND U3458 ( .A(n3283), .B(n3282), .Z(n3284) );
  NAND U3459 ( .A(n3285), .B(n3284), .Z(n3346) );
  NANDN U3460 ( .A(n3287), .B(n3286), .Z(n3291) );
  NAND U3461 ( .A(n3289), .B(n3288), .Z(n3290) );
  NAND U3462 ( .A(n3291), .B(n3290), .Z(n3344) );
  XNOR U3463 ( .A(b[7]), .B(a[75]), .Z(n3331) );
  NANDN U3464 ( .A(n3331), .B(n5293), .Z(n3294) );
  NANDN U3465 ( .A(n3292), .B(n5294), .Z(n3293) );
  NAND U3466 ( .A(n3294), .B(n3293), .Z(n3319) );
  XNOR U3467 ( .A(b[3]), .B(a[79]), .Z(n3334) );
  NANDN U3468 ( .A(n3334), .B(n5160), .Z(n3297) );
  NANDN U3469 ( .A(n3295), .B(n5161), .Z(n3296) );
  AND U3470 ( .A(n3297), .B(n3296), .Z(n3320) );
  XNOR U3471 ( .A(n3319), .B(n3320), .Z(n3321) );
  NANDN U3472 ( .A(n292), .B(a[81]), .Z(n3298) );
  XOR U3473 ( .A(n5199), .B(n3298), .Z(n3300) );
  NANDN U3474 ( .A(b[0]), .B(a[80]), .Z(n3299) );
  AND U3475 ( .A(n3300), .B(n3299), .Z(n3327) );
  XNOR U3476 ( .A(b[5]), .B(a[77]), .Z(n3340) );
  NANDN U3477 ( .A(n3340), .B(n5240), .Z(n3303) );
  NANDN U3478 ( .A(n3301), .B(n5241), .Z(n3302) );
  NAND U3479 ( .A(n3303), .B(n3302), .Z(n3325) );
  NANDN U3480 ( .A(n295), .B(a[73]), .Z(n3326) );
  XNOR U3481 ( .A(n3325), .B(n3326), .Z(n3328) );
  XOR U3482 ( .A(n3327), .B(n3328), .Z(n3322) );
  XOR U3483 ( .A(n3321), .B(n3322), .Z(n3343) );
  XOR U3484 ( .A(n3344), .B(n3343), .Z(n3345) );
  XNOR U3485 ( .A(n3346), .B(n3345), .Z(n3315) );
  NAND U3486 ( .A(n3305), .B(n3304), .Z(n3309) );
  NAND U3487 ( .A(n3307), .B(n3306), .Z(n3308) );
  NAND U3488 ( .A(n3309), .B(n3308), .Z(n3316) );
  XNOR U3489 ( .A(n3315), .B(n3316), .Z(n3317) );
  XNOR U3490 ( .A(n3318), .B(n3317), .Z(n3349) );
  XNOR U3491 ( .A(n3349), .B(sreg[201]), .Z(n3351) );
  NAND U3492 ( .A(n3310), .B(sreg[200]), .Z(n3314) );
  OR U3493 ( .A(n3312), .B(n3311), .Z(n3313) );
  AND U3494 ( .A(n3314), .B(n3313), .Z(n3350) );
  XOR U3495 ( .A(n3351), .B(n3350), .Z(c[201]) );
  NANDN U3496 ( .A(n3320), .B(n3319), .Z(n3324) );
  NAND U3497 ( .A(n3322), .B(n3321), .Z(n3323) );
  NAND U3498 ( .A(n3324), .B(n3323), .Z(n3385) );
  NANDN U3499 ( .A(n3326), .B(n3325), .Z(n3330) );
  NAND U3500 ( .A(n3328), .B(n3327), .Z(n3329) );
  NAND U3501 ( .A(n3330), .B(n3329), .Z(n3383) );
  XNOR U3502 ( .A(b[7]), .B(a[76]), .Z(n3370) );
  NANDN U3503 ( .A(n3370), .B(n5293), .Z(n3333) );
  NANDN U3504 ( .A(n3331), .B(n5294), .Z(n3332) );
  NAND U3505 ( .A(n3333), .B(n3332), .Z(n3358) );
  XNOR U3506 ( .A(b[3]), .B(a[80]), .Z(n3373) );
  NANDN U3507 ( .A(n3373), .B(n5160), .Z(n3336) );
  NANDN U3508 ( .A(n3334), .B(n5161), .Z(n3335) );
  AND U3509 ( .A(n3336), .B(n3335), .Z(n3359) );
  XNOR U3510 ( .A(n3358), .B(n3359), .Z(n3360) );
  NANDN U3511 ( .A(n292), .B(a[82]), .Z(n3337) );
  XOR U3512 ( .A(n5199), .B(n3337), .Z(n3339) );
  NANDN U3513 ( .A(b[0]), .B(a[81]), .Z(n3338) );
  AND U3514 ( .A(n3339), .B(n3338), .Z(n3366) );
  XNOR U3515 ( .A(b[5]), .B(a[78]), .Z(n3379) );
  NANDN U3516 ( .A(n3379), .B(n5240), .Z(n3342) );
  NANDN U3517 ( .A(n3340), .B(n5241), .Z(n3341) );
  NAND U3518 ( .A(n3342), .B(n3341), .Z(n3364) );
  NANDN U3519 ( .A(n295), .B(a[74]), .Z(n3365) );
  XNOR U3520 ( .A(n3364), .B(n3365), .Z(n3367) );
  XOR U3521 ( .A(n3366), .B(n3367), .Z(n3361) );
  XOR U3522 ( .A(n3360), .B(n3361), .Z(n3382) );
  XOR U3523 ( .A(n3383), .B(n3382), .Z(n3384) );
  XNOR U3524 ( .A(n3385), .B(n3384), .Z(n3354) );
  NAND U3525 ( .A(n3344), .B(n3343), .Z(n3348) );
  NAND U3526 ( .A(n3346), .B(n3345), .Z(n3347) );
  NAND U3527 ( .A(n3348), .B(n3347), .Z(n3355) );
  XNOR U3528 ( .A(n3354), .B(n3355), .Z(n3356) );
  XNOR U3529 ( .A(n3357), .B(n3356), .Z(n3388) );
  XNOR U3530 ( .A(n3388), .B(sreg[202]), .Z(n3390) );
  NAND U3531 ( .A(n3349), .B(sreg[201]), .Z(n3353) );
  OR U3532 ( .A(n3351), .B(n3350), .Z(n3352) );
  AND U3533 ( .A(n3353), .B(n3352), .Z(n3389) );
  XOR U3534 ( .A(n3390), .B(n3389), .Z(c[202]) );
  NANDN U3535 ( .A(n3359), .B(n3358), .Z(n3363) );
  NAND U3536 ( .A(n3361), .B(n3360), .Z(n3362) );
  NAND U3537 ( .A(n3363), .B(n3362), .Z(n3424) );
  NANDN U3538 ( .A(n3365), .B(n3364), .Z(n3369) );
  NAND U3539 ( .A(n3367), .B(n3366), .Z(n3368) );
  NAND U3540 ( .A(n3369), .B(n3368), .Z(n3422) );
  XNOR U3541 ( .A(b[7]), .B(a[77]), .Z(n3409) );
  NANDN U3542 ( .A(n3409), .B(n5293), .Z(n3372) );
  NANDN U3543 ( .A(n3370), .B(n5294), .Z(n3371) );
  NAND U3544 ( .A(n3372), .B(n3371), .Z(n3397) );
  XNOR U3545 ( .A(b[3]), .B(a[81]), .Z(n3412) );
  NANDN U3546 ( .A(n3412), .B(n5160), .Z(n3375) );
  NANDN U3547 ( .A(n3373), .B(n5161), .Z(n3374) );
  AND U3548 ( .A(n3375), .B(n3374), .Z(n3398) );
  XNOR U3549 ( .A(n3397), .B(n3398), .Z(n3399) );
  NANDN U3550 ( .A(n292), .B(a[83]), .Z(n3376) );
  XOR U3551 ( .A(n5199), .B(n3376), .Z(n3378) );
  NANDN U3552 ( .A(b[0]), .B(a[82]), .Z(n3377) );
  AND U3553 ( .A(n3378), .B(n3377), .Z(n3405) );
  XNOR U3554 ( .A(b[5]), .B(a[79]), .Z(n3418) );
  NANDN U3555 ( .A(n3418), .B(n5240), .Z(n3381) );
  NANDN U3556 ( .A(n3379), .B(n5241), .Z(n3380) );
  NAND U3557 ( .A(n3381), .B(n3380), .Z(n3403) );
  NANDN U3558 ( .A(n295), .B(a[75]), .Z(n3404) );
  XNOR U3559 ( .A(n3403), .B(n3404), .Z(n3406) );
  XOR U3560 ( .A(n3405), .B(n3406), .Z(n3400) );
  XOR U3561 ( .A(n3399), .B(n3400), .Z(n3421) );
  XOR U3562 ( .A(n3422), .B(n3421), .Z(n3423) );
  XNOR U3563 ( .A(n3424), .B(n3423), .Z(n3393) );
  NAND U3564 ( .A(n3383), .B(n3382), .Z(n3387) );
  NAND U3565 ( .A(n3385), .B(n3384), .Z(n3386) );
  NAND U3566 ( .A(n3387), .B(n3386), .Z(n3394) );
  XNOR U3567 ( .A(n3393), .B(n3394), .Z(n3395) );
  XNOR U3568 ( .A(n3396), .B(n3395), .Z(n3427) );
  XNOR U3569 ( .A(n3427), .B(sreg[203]), .Z(n3429) );
  NAND U3570 ( .A(n3388), .B(sreg[202]), .Z(n3392) );
  OR U3571 ( .A(n3390), .B(n3389), .Z(n3391) );
  AND U3572 ( .A(n3392), .B(n3391), .Z(n3428) );
  XOR U3573 ( .A(n3429), .B(n3428), .Z(c[203]) );
  NANDN U3574 ( .A(n3398), .B(n3397), .Z(n3402) );
  NAND U3575 ( .A(n3400), .B(n3399), .Z(n3401) );
  NAND U3576 ( .A(n3402), .B(n3401), .Z(n3463) );
  NANDN U3577 ( .A(n3404), .B(n3403), .Z(n3408) );
  NAND U3578 ( .A(n3406), .B(n3405), .Z(n3407) );
  NAND U3579 ( .A(n3408), .B(n3407), .Z(n3461) );
  XNOR U3580 ( .A(b[7]), .B(a[78]), .Z(n3448) );
  NANDN U3581 ( .A(n3448), .B(n5293), .Z(n3411) );
  NANDN U3582 ( .A(n3409), .B(n5294), .Z(n3410) );
  NAND U3583 ( .A(n3411), .B(n3410), .Z(n3436) );
  XNOR U3584 ( .A(b[3]), .B(a[82]), .Z(n3451) );
  NANDN U3585 ( .A(n3451), .B(n5160), .Z(n3414) );
  NANDN U3586 ( .A(n3412), .B(n5161), .Z(n3413) );
  AND U3587 ( .A(n3414), .B(n3413), .Z(n3437) );
  XNOR U3588 ( .A(n3436), .B(n3437), .Z(n3438) );
  NANDN U3589 ( .A(n292), .B(a[84]), .Z(n3415) );
  XOR U3590 ( .A(n5199), .B(n3415), .Z(n3417) );
  NANDN U3591 ( .A(b[0]), .B(a[83]), .Z(n3416) );
  AND U3592 ( .A(n3417), .B(n3416), .Z(n3444) );
  XNOR U3593 ( .A(b[5]), .B(a[80]), .Z(n3457) );
  NANDN U3594 ( .A(n3457), .B(n5240), .Z(n3420) );
  NANDN U3595 ( .A(n3418), .B(n5241), .Z(n3419) );
  NAND U3596 ( .A(n3420), .B(n3419), .Z(n3442) );
  NANDN U3597 ( .A(n295), .B(a[76]), .Z(n3443) );
  XNOR U3598 ( .A(n3442), .B(n3443), .Z(n3445) );
  XOR U3599 ( .A(n3444), .B(n3445), .Z(n3439) );
  XOR U3600 ( .A(n3438), .B(n3439), .Z(n3460) );
  XOR U3601 ( .A(n3461), .B(n3460), .Z(n3462) );
  XNOR U3602 ( .A(n3463), .B(n3462), .Z(n3432) );
  NAND U3603 ( .A(n3422), .B(n3421), .Z(n3426) );
  NAND U3604 ( .A(n3424), .B(n3423), .Z(n3425) );
  NAND U3605 ( .A(n3426), .B(n3425), .Z(n3433) );
  XNOR U3606 ( .A(n3432), .B(n3433), .Z(n3434) );
  XNOR U3607 ( .A(n3435), .B(n3434), .Z(n3466) );
  XNOR U3608 ( .A(n3466), .B(sreg[204]), .Z(n3468) );
  NAND U3609 ( .A(n3427), .B(sreg[203]), .Z(n3431) );
  OR U3610 ( .A(n3429), .B(n3428), .Z(n3430) );
  AND U3611 ( .A(n3431), .B(n3430), .Z(n3467) );
  XOR U3612 ( .A(n3468), .B(n3467), .Z(c[204]) );
  NANDN U3613 ( .A(n3437), .B(n3436), .Z(n3441) );
  NAND U3614 ( .A(n3439), .B(n3438), .Z(n3440) );
  NAND U3615 ( .A(n3441), .B(n3440), .Z(n3502) );
  NANDN U3616 ( .A(n3443), .B(n3442), .Z(n3447) );
  NAND U3617 ( .A(n3445), .B(n3444), .Z(n3446) );
  NAND U3618 ( .A(n3447), .B(n3446), .Z(n3500) );
  XNOR U3619 ( .A(b[7]), .B(a[79]), .Z(n3487) );
  NANDN U3620 ( .A(n3487), .B(n5293), .Z(n3450) );
  NANDN U3621 ( .A(n3448), .B(n5294), .Z(n3449) );
  NAND U3622 ( .A(n3450), .B(n3449), .Z(n3475) );
  XNOR U3623 ( .A(b[3]), .B(a[83]), .Z(n3490) );
  NANDN U3624 ( .A(n3490), .B(n5160), .Z(n3453) );
  NANDN U3625 ( .A(n3451), .B(n5161), .Z(n3452) );
  AND U3626 ( .A(n3453), .B(n3452), .Z(n3476) );
  XNOR U3627 ( .A(n3475), .B(n3476), .Z(n3477) );
  NANDN U3628 ( .A(n292), .B(a[85]), .Z(n3454) );
  XOR U3629 ( .A(n5199), .B(n3454), .Z(n3456) );
  NANDN U3630 ( .A(b[0]), .B(a[84]), .Z(n3455) );
  AND U3631 ( .A(n3456), .B(n3455), .Z(n3483) );
  XNOR U3632 ( .A(b[5]), .B(a[81]), .Z(n3496) );
  NANDN U3633 ( .A(n3496), .B(n5240), .Z(n3459) );
  NANDN U3634 ( .A(n3457), .B(n5241), .Z(n3458) );
  NAND U3635 ( .A(n3459), .B(n3458), .Z(n3481) );
  NANDN U3636 ( .A(n295), .B(a[77]), .Z(n3482) );
  XNOR U3637 ( .A(n3481), .B(n3482), .Z(n3484) );
  XOR U3638 ( .A(n3483), .B(n3484), .Z(n3478) );
  XOR U3639 ( .A(n3477), .B(n3478), .Z(n3499) );
  XOR U3640 ( .A(n3500), .B(n3499), .Z(n3501) );
  XNOR U3641 ( .A(n3502), .B(n3501), .Z(n3471) );
  NAND U3642 ( .A(n3461), .B(n3460), .Z(n3465) );
  NAND U3643 ( .A(n3463), .B(n3462), .Z(n3464) );
  NAND U3644 ( .A(n3465), .B(n3464), .Z(n3472) );
  XNOR U3645 ( .A(n3471), .B(n3472), .Z(n3473) );
  XNOR U3646 ( .A(n3474), .B(n3473), .Z(n3505) );
  XNOR U3647 ( .A(n3505), .B(sreg[205]), .Z(n3507) );
  NAND U3648 ( .A(n3466), .B(sreg[204]), .Z(n3470) );
  OR U3649 ( .A(n3468), .B(n3467), .Z(n3469) );
  AND U3650 ( .A(n3470), .B(n3469), .Z(n3506) );
  XOR U3651 ( .A(n3507), .B(n3506), .Z(c[205]) );
  NANDN U3652 ( .A(n3476), .B(n3475), .Z(n3480) );
  NAND U3653 ( .A(n3478), .B(n3477), .Z(n3479) );
  NAND U3654 ( .A(n3480), .B(n3479), .Z(n3541) );
  NANDN U3655 ( .A(n3482), .B(n3481), .Z(n3486) );
  NAND U3656 ( .A(n3484), .B(n3483), .Z(n3485) );
  NAND U3657 ( .A(n3486), .B(n3485), .Z(n3539) );
  XNOR U3658 ( .A(b[7]), .B(a[80]), .Z(n3526) );
  NANDN U3659 ( .A(n3526), .B(n5293), .Z(n3489) );
  NANDN U3660 ( .A(n3487), .B(n5294), .Z(n3488) );
  NAND U3661 ( .A(n3489), .B(n3488), .Z(n3514) );
  XNOR U3662 ( .A(b[3]), .B(a[84]), .Z(n3529) );
  NANDN U3663 ( .A(n3529), .B(n5160), .Z(n3492) );
  NANDN U3664 ( .A(n3490), .B(n5161), .Z(n3491) );
  AND U3665 ( .A(n3492), .B(n3491), .Z(n3515) );
  XNOR U3666 ( .A(n3514), .B(n3515), .Z(n3516) );
  NANDN U3667 ( .A(n292), .B(a[86]), .Z(n3493) );
  XOR U3668 ( .A(n5199), .B(n3493), .Z(n3495) );
  NANDN U3669 ( .A(b[0]), .B(a[85]), .Z(n3494) );
  AND U3670 ( .A(n3495), .B(n3494), .Z(n3522) );
  XNOR U3671 ( .A(b[5]), .B(a[82]), .Z(n3535) );
  NANDN U3672 ( .A(n3535), .B(n5240), .Z(n3498) );
  NANDN U3673 ( .A(n3496), .B(n5241), .Z(n3497) );
  NAND U3674 ( .A(n3498), .B(n3497), .Z(n3520) );
  NANDN U3675 ( .A(n295), .B(a[78]), .Z(n3521) );
  XNOR U3676 ( .A(n3520), .B(n3521), .Z(n3523) );
  XOR U3677 ( .A(n3522), .B(n3523), .Z(n3517) );
  XOR U3678 ( .A(n3516), .B(n3517), .Z(n3538) );
  XOR U3679 ( .A(n3539), .B(n3538), .Z(n3540) );
  XNOR U3680 ( .A(n3541), .B(n3540), .Z(n3510) );
  NAND U3681 ( .A(n3500), .B(n3499), .Z(n3504) );
  NAND U3682 ( .A(n3502), .B(n3501), .Z(n3503) );
  NAND U3683 ( .A(n3504), .B(n3503), .Z(n3511) );
  XNOR U3684 ( .A(n3510), .B(n3511), .Z(n3512) );
  XNOR U3685 ( .A(n3513), .B(n3512), .Z(n3544) );
  XNOR U3686 ( .A(n3544), .B(sreg[206]), .Z(n3546) );
  NAND U3687 ( .A(n3505), .B(sreg[205]), .Z(n3509) );
  OR U3688 ( .A(n3507), .B(n3506), .Z(n3508) );
  AND U3689 ( .A(n3509), .B(n3508), .Z(n3545) );
  XOR U3690 ( .A(n3546), .B(n3545), .Z(c[206]) );
  NANDN U3691 ( .A(n3515), .B(n3514), .Z(n3519) );
  NAND U3692 ( .A(n3517), .B(n3516), .Z(n3518) );
  NAND U3693 ( .A(n3519), .B(n3518), .Z(n3580) );
  NANDN U3694 ( .A(n3521), .B(n3520), .Z(n3525) );
  NAND U3695 ( .A(n3523), .B(n3522), .Z(n3524) );
  NAND U3696 ( .A(n3525), .B(n3524), .Z(n3578) );
  XNOR U3697 ( .A(b[7]), .B(a[81]), .Z(n3565) );
  NANDN U3698 ( .A(n3565), .B(n5293), .Z(n3528) );
  NANDN U3699 ( .A(n3526), .B(n5294), .Z(n3527) );
  NAND U3700 ( .A(n3528), .B(n3527), .Z(n3553) );
  XNOR U3701 ( .A(b[3]), .B(a[85]), .Z(n3568) );
  NANDN U3702 ( .A(n3568), .B(n5160), .Z(n3531) );
  NANDN U3703 ( .A(n3529), .B(n5161), .Z(n3530) );
  AND U3704 ( .A(n3531), .B(n3530), .Z(n3554) );
  XNOR U3705 ( .A(n3553), .B(n3554), .Z(n3555) );
  NANDN U3706 ( .A(n292), .B(a[87]), .Z(n3532) );
  XOR U3707 ( .A(n5199), .B(n3532), .Z(n3534) );
  NANDN U3708 ( .A(b[0]), .B(a[86]), .Z(n3533) );
  AND U3709 ( .A(n3534), .B(n3533), .Z(n3561) );
  XNOR U3710 ( .A(b[5]), .B(a[83]), .Z(n3574) );
  NANDN U3711 ( .A(n3574), .B(n5240), .Z(n3537) );
  NANDN U3712 ( .A(n3535), .B(n5241), .Z(n3536) );
  NAND U3713 ( .A(n3537), .B(n3536), .Z(n3559) );
  NANDN U3714 ( .A(n295), .B(a[79]), .Z(n3560) );
  XNOR U3715 ( .A(n3559), .B(n3560), .Z(n3562) );
  XOR U3716 ( .A(n3561), .B(n3562), .Z(n3556) );
  XOR U3717 ( .A(n3555), .B(n3556), .Z(n3577) );
  XOR U3718 ( .A(n3578), .B(n3577), .Z(n3579) );
  XNOR U3719 ( .A(n3580), .B(n3579), .Z(n3549) );
  NAND U3720 ( .A(n3539), .B(n3538), .Z(n3543) );
  NAND U3721 ( .A(n3541), .B(n3540), .Z(n3542) );
  NAND U3722 ( .A(n3543), .B(n3542), .Z(n3550) );
  XNOR U3723 ( .A(n3549), .B(n3550), .Z(n3551) );
  XNOR U3724 ( .A(n3552), .B(n3551), .Z(n3583) );
  XNOR U3725 ( .A(n3583), .B(sreg[207]), .Z(n3585) );
  NAND U3726 ( .A(n3544), .B(sreg[206]), .Z(n3548) );
  OR U3727 ( .A(n3546), .B(n3545), .Z(n3547) );
  AND U3728 ( .A(n3548), .B(n3547), .Z(n3584) );
  XOR U3729 ( .A(n3585), .B(n3584), .Z(c[207]) );
  NANDN U3730 ( .A(n3554), .B(n3553), .Z(n3558) );
  NAND U3731 ( .A(n3556), .B(n3555), .Z(n3557) );
  NAND U3732 ( .A(n3558), .B(n3557), .Z(n3619) );
  NANDN U3733 ( .A(n3560), .B(n3559), .Z(n3564) );
  NAND U3734 ( .A(n3562), .B(n3561), .Z(n3563) );
  NAND U3735 ( .A(n3564), .B(n3563), .Z(n3617) );
  XNOR U3736 ( .A(b[7]), .B(a[82]), .Z(n3604) );
  NANDN U3737 ( .A(n3604), .B(n5293), .Z(n3567) );
  NANDN U3738 ( .A(n3565), .B(n5294), .Z(n3566) );
  NAND U3739 ( .A(n3567), .B(n3566), .Z(n3592) );
  XNOR U3740 ( .A(b[3]), .B(a[86]), .Z(n3607) );
  NANDN U3741 ( .A(n3607), .B(n5160), .Z(n3570) );
  NANDN U3742 ( .A(n3568), .B(n5161), .Z(n3569) );
  AND U3743 ( .A(n3570), .B(n3569), .Z(n3593) );
  XNOR U3744 ( .A(n3592), .B(n3593), .Z(n3594) );
  NANDN U3745 ( .A(n292), .B(a[88]), .Z(n3571) );
  XOR U3746 ( .A(n5199), .B(n3571), .Z(n3573) );
  NANDN U3747 ( .A(b[0]), .B(a[87]), .Z(n3572) );
  AND U3748 ( .A(n3573), .B(n3572), .Z(n3600) );
  XNOR U3749 ( .A(b[5]), .B(a[84]), .Z(n3613) );
  NANDN U3750 ( .A(n3613), .B(n5240), .Z(n3576) );
  NANDN U3751 ( .A(n3574), .B(n5241), .Z(n3575) );
  NAND U3752 ( .A(n3576), .B(n3575), .Z(n3598) );
  NANDN U3753 ( .A(n295), .B(a[80]), .Z(n3599) );
  XNOR U3754 ( .A(n3598), .B(n3599), .Z(n3601) );
  XOR U3755 ( .A(n3600), .B(n3601), .Z(n3595) );
  XOR U3756 ( .A(n3594), .B(n3595), .Z(n3616) );
  XOR U3757 ( .A(n3617), .B(n3616), .Z(n3618) );
  XNOR U3758 ( .A(n3619), .B(n3618), .Z(n3588) );
  NAND U3759 ( .A(n3578), .B(n3577), .Z(n3582) );
  NAND U3760 ( .A(n3580), .B(n3579), .Z(n3581) );
  NAND U3761 ( .A(n3582), .B(n3581), .Z(n3589) );
  XNOR U3762 ( .A(n3588), .B(n3589), .Z(n3590) );
  XNOR U3763 ( .A(n3591), .B(n3590), .Z(n3622) );
  XNOR U3764 ( .A(n3622), .B(sreg[208]), .Z(n3624) );
  NAND U3765 ( .A(n3583), .B(sreg[207]), .Z(n3587) );
  OR U3766 ( .A(n3585), .B(n3584), .Z(n3586) );
  AND U3767 ( .A(n3587), .B(n3586), .Z(n3623) );
  XOR U3768 ( .A(n3624), .B(n3623), .Z(c[208]) );
  NANDN U3769 ( .A(n3593), .B(n3592), .Z(n3597) );
  NAND U3770 ( .A(n3595), .B(n3594), .Z(n3596) );
  NAND U3771 ( .A(n3597), .B(n3596), .Z(n3658) );
  NANDN U3772 ( .A(n3599), .B(n3598), .Z(n3603) );
  NAND U3773 ( .A(n3601), .B(n3600), .Z(n3602) );
  NAND U3774 ( .A(n3603), .B(n3602), .Z(n3656) );
  XNOR U3775 ( .A(b[7]), .B(a[83]), .Z(n3643) );
  NANDN U3776 ( .A(n3643), .B(n5293), .Z(n3606) );
  NANDN U3777 ( .A(n3604), .B(n5294), .Z(n3605) );
  NAND U3778 ( .A(n3606), .B(n3605), .Z(n3631) );
  XNOR U3779 ( .A(b[3]), .B(a[87]), .Z(n3646) );
  NANDN U3780 ( .A(n3646), .B(n5160), .Z(n3609) );
  NANDN U3781 ( .A(n3607), .B(n5161), .Z(n3608) );
  AND U3782 ( .A(n3609), .B(n3608), .Z(n3632) );
  XNOR U3783 ( .A(n3631), .B(n3632), .Z(n3633) );
  NANDN U3784 ( .A(n292), .B(a[89]), .Z(n3610) );
  XOR U3785 ( .A(n5199), .B(n3610), .Z(n3612) );
  NANDN U3786 ( .A(b[0]), .B(a[88]), .Z(n3611) );
  AND U3787 ( .A(n3612), .B(n3611), .Z(n3639) );
  XNOR U3788 ( .A(b[5]), .B(a[85]), .Z(n3652) );
  NANDN U3789 ( .A(n3652), .B(n5240), .Z(n3615) );
  NANDN U3790 ( .A(n3613), .B(n5241), .Z(n3614) );
  NAND U3791 ( .A(n3615), .B(n3614), .Z(n3637) );
  NANDN U3792 ( .A(n295), .B(a[81]), .Z(n3638) );
  XNOR U3793 ( .A(n3637), .B(n3638), .Z(n3640) );
  XOR U3794 ( .A(n3639), .B(n3640), .Z(n3634) );
  XOR U3795 ( .A(n3633), .B(n3634), .Z(n3655) );
  XOR U3796 ( .A(n3656), .B(n3655), .Z(n3657) );
  XNOR U3797 ( .A(n3658), .B(n3657), .Z(n3627) );
  NAND U3798 ( .A(n3617), .B(n3616), .Z(n3621) );
  NAND U3799 ( .A(n3619), .B(n3618), .Z(n3620) );
  NAND U3800 ( .A(n3621), .B(n3620), .Z(n3628) );
  XNOR U3801 ( .A(n3627), .B(n3628), .Z(n3629) );
  XNOR U3802 ( .A(n3630), .B(n3629), .Z(n3661) );
  XNOR U3803 ( .A(n3661), .B(sreg[209]), .Z(n3663) );
  NAND U3804 ( .A(n3622), .B(sreg[208]), .Z(n3626) );
  OR U3805 ( .A(n3624), .B(n3623), .Z(n3625) );
  AND U3806 ( .A(n3626), .B(n3625), .Z(n3662) );
  XOR U3807 ( .A(n3663), .B(n3662), .Z(c[209]) );
  NANDN U3808 ( .A(n3632), .B(n3631), .Z(n3636) );
  NAND U3809 ( .A(n3634), .B(n3633), .Z(n3635) );
  NAND U3810 ( .A(n3636), .B(n3635), .Z(n3697) );
  NANDN U3811 ( .A(n3638), .B(n3637), .Z(n3642) );
  NAND U3812 ( .A(n3640), .B(n3639), .Z(n3641) );
  NAND U3813 ( .A(n3642), .B(n3641), .Z(n3695) );
  XNOR U3814 ( .A(b[7]), .B(a[84]), .Z(n3682) );
  NANDN U3815 ( .A(n3682), .B(n5293), .Z(n3645) );
  NANDN U3816 ( .A(n3643), .B(n5294), .Z(n3644) );
  NAND U3817 ( .A(n3645), .B(n3644), .Z(n3670) );
  XNOR U3818 ( .A(b[3]), .B(a[88]), .Z(n3685) );
  NANDN U3819 ( .A(n3685), .B(n5160), .Z(n3648) );
  NANDN U3820 ( .A(n3646), .B(n5161), .Z(n3647) );
  AND U3821 ( .A(n3648), .B(n3647), .Z(n3671) );
  XNOR U3822 ( .A(n3670), .B(n3671), .Z(n3672) );
  NANDN U3823 ( .A(n292), .B(a[90]), .Z(n3649) );
  XOR U3824 ( .A(n5199), .B(n3649), .Z(n3651) );
  NANDN U3825 ( .A(b[0]), .B(a[89]), .Z(n3650) );
  AND U3826 ( .A(n3651), .B(n3650), .Z(n3678) );
  XNOR U3827 ( .A(b[5]), .B(a[86]), .Z(n3691) );
  NANDN U3828 ( .A(n3691), .B(n5240), .Z(n3654) );
  NANDN U3829 ( .A(n3652), .B(n5241), .Z(n3653) );
  NAND U3830 ( .A(n3654), .B(n3653), .Z(n3676) );
  NANDN U3831 ( .A(n295), .B(a[82]), .Z(n3677) );
  XNOR U3832 ( .A(n3676), .B(n3677), .Z(n3679) );
  XOR U3833 ( .A(n3678), .B(n3679), .Z(n3673) );
  XOR U3834 ( .A(n3672), .B(n3673), .Z(n3694) );
  XOR U3835 ( .A(n3695), .B(n3694), .Z(n3696) );
  XNOR U3836 ( .A(n3697), .B(n3696), .Z(n3666) );
  NAND U3837 ( .A(n3656), .B(n3655), .Z(n3660) );
  NAND U3838 ( .A(n3658), .B(n3657), .Z(n3659) );
  NAND U3839 ( .A(n3660), .B(n3659), .Z(n3667) );
  XNOR U3840 ( .A(n3666), .B(n3667), .Z(n3668) );
  XNOR U3841 ( .A(n3669), .B(n3668), .Z(n3700) );
  XNOR U3842 ( .A(n3700), .B(sreg[210]), .Z(n3702) );
  NAND U3843 ( .A(n3661), .B(sreg[209]), .Z(n3665) );
  OR U3844 ( .A(n3663), .B(n3662), .Z(n3664) );
  AND U3845 ( .A(n3665), .B(n3664), .Z(n3701) );
  XOR U3846 ( .A(n3702), .B(n3701), .Z(c[210]) );
  NANDN U3847 ( .A(n3671), .B(n3670), .Z(n3675) );
  NAND U3848 ( .A(n3673), .B(n3672), .Z(n3674) );
  NAND U3849 ( .A(n3675), .B(n3674), .Z(n3736) );
  NANDN U3850 ( .A(n3677), .B(n3676), .Z(n3681) );
  NAND U3851 ( .A(n3679), .B(n3678), .Z(n3680) );
  NAND U3852 ( .A(n3681), .B(n3680), .Z(n3734) );
  XNOR U3853 ( .A(b[7]), .B(a[85]), .Z(n3721) );
  NANDN U3854 ( .A(n3721), .B(n5293), .Z(n3684) );
  NANDN U3855 ( .A(n3682), .B(n5294), .Z(n3683) );
  NAND U3856 ( .A(n3684), .B(n3683), .Z(n3709) );
  XNOR U3857 ( .A(b[3]), .B(a[89]), .Z(n3724) );
  NANDN U3858 ( .A(n3724), .B(n5160), .Z(n3687) );
  NANDN U3859 ( .A(n3685), .B(n5161), .Z(n3686) );
  AND U3860 ( .A(n3687), .B(n3686), .Z(n3710) );
  XNOR U3861 ( .A(n3709), .B(n3710), .Z(n3711) );
  NANDN U3862 ( .A(n292), .B(a[91]), .Z(n3688) );
  XOR U3863 ( .A(n5199), .B(n3688), .Z(n3690) );
  NANDN U3864 ( .A(b[0]), .B(a[90]), .Z(n3689) );
  AND U3865 ( .A(n3690), .B(n3689), .Z(n3717) );
  XNOR U3866 ( .A(b[5]), .B(a[87]), .Z(n3730) );
  NANDN U3867 ( .A(n3730), .B(n5240), .Z(n3693) );
  NANDN U3868 ( .A(n3691), .B(n5241), .Z(n3692) );
  NAND U3869 ( .A(n3693), .B(n3692), .Z(n3715) );
  NANDN U3870 ( .A(n295), .B(a[83]), .Z(n3716) );
  XNOR U3871 ( .A(n3715), .B(n3716), .Z(n3718) );
  XOR U3872 ( .A(n3717), .B(n3718), .Z(n3712) );
  XOR U3873 ( .A(n3711), .B(n3712), .Z(n3733) );
  XOR U3874 ( .A(n3734), .B(n3733), .Z(n3735) );
  XNOR U3875 ( .A(n3736), .B(n3735), .Z(n3705) );
  NAND U3876 ( .A(n3695), .B(n3694), .Z(n3699) );
  NAND U3877 ( .A(n3697), .B(n3696), .Z(n3698) );
  NAND U3878 ( .A(n3699), .B(n3698), .Z(n3706) );
  XNOR U3879 ( .A(n3705), .B(n3706), .Z(n3707) );
  XNOR U3880 ( .A(n3708), .B(n3707), .Z(n3739) );
  XNOR U3881 ( .A(n3739), .B(sreg[211]), .Z(n3741) );
  NAND U3882 ( .A(n3700), .B(sreg[210]), .Z(n3704) );
  OR U3883 ( .A(n3702), .B(n3701), .Z(n3703) );
  AND U3884 ( .A(n3704), .B(n3703), .Z(n3740) );
  XOR U3885 ( .A(n3741), .B(n3740), .Z(c[211]) );
  NANDN U3886 ( .A(n3710), .B(n3709), .Z(n3714) );
  NAND U3887 ( .A(n3712), .B(n3711), .Z(n3713) );
  NAND U3888 ( .A(n3714), .B(n3713), .Z(n3775) );
  NANDN U3889 ( .A(n3716), .B(n3715), .Z(n3720) );
  NAND U3890 ( .A(n3718), .B(n3717), .Z(n3719) );
  NAND U3891 ( .A(n3720), .B(n3719), .Z(n3773) );
  XNOR U3892 ( .A(b[7]), .B(a[86]), .Z(n3760) );
  NANDN U3893 ( .A(n3760), .B(n5293), .Z(n3723) );
  NANDN U3894 ( .A(n3721), .B(n5294), .Z(n3722) );
  NAND U3895 ( .A(n3723), .B(n3722), .Z(n3748) );
  XNOR U3896 ( .A(b[3]), .B(a[90]), .Z(n3763) );
  NANDN U3897 ( .A(n3763), .B(n5160), .Z(n3726) );
  NANDN U3898 ( .A(n3724), .B(n5161), .Z(n3725) );
  AND U3899 ( .A(n3726), .B(n3725), .Z(n3749) );
  XNOR U3900 ( .A(n3748), .B(n3749), .Z(n3750) );
  NANDN U3901 ( .A(n292), .B(a[92]), .Z(n3727) );
  XOR U3902 ( .A(n5199), .B(n3727), .Z(n3729) );
  NANDN U3903 ( .A(b[0]), .B(a[91]), .Z(n3728) );
  AND U3904 ( .A(n3729), .B(n3728), .Z(n3756) );
  XNOR U3905 ( .A(b[5]), .B(a[88]), .Z(n3769) );
  NANDN U3906 ( .A(n3769), .B(n5240), .Z(n3732) );
  NANDN U3907 ( .A(n3730), .B(n5241), .Z(n3731) );
  NAND U3908 ( .A(n3732), .B(n3731), .Z(n3754) );
  NANDN U3909 ( .A(n295), .B(a[84]), .Z(n3755) );
  XNOR U3910 ( .A(n3754), .B(n3755), .Z(n3757) );
  XOR U3911 ( .A(n3756), .B(n3757), .Z(n3751) );
  XOR U3912 ( .A(n3750), .B(n3751), .Z(n3772) );
  XOR U3913 ( .A(n3773), .B(n3772), .Z(n3774) );
  XNOR U3914 ( .A(n3775), .B(n3774), .Z(n3744) );
  NAND U3915 ( .A(n3734), .B(n3733), .Z(n3738) );
  NAND U3916 ( .A(n3736), .B(n3735), .Z(n3737) );
  NAND U3917 ( .A(n3738), .B(n3737), .Z(n3745) );
  XNOR U3918 ( .A(n3744), .B(n3745), .Z(n3746) );
  XNOR U3919 ( .A(n3747), .B(n3746), .Z(n3778) );
  XNOR U3920 ( .A(n3778), .B(sreg[212]), .Z(n3780) );
  NAND U3921 ( .A(n3739), .B(sreg[211]), .Z(n3743) );
  OR U3922 ( .A(n3741), .B(n3740), .Z(n3742) );
  AND U3923 ( .A(n3743), .B(n3742), .Z(n3779) );
  XOR U3924 ( .A(n3780), .B(n3779), .Z(c[212]) );
  NANDN U3925 ( .A(n3749), .B(n3748), .Z(n3753) );
  NAND U3926 ( .A(n3751), .B(n3750), .Z(n3752) );
  NAND U3927 ( .A(n3753), .B(n3752), .Z(n3814) );
  NANDN U3928 ( .A(n3755), .B(n3754), .Z(n3759) );
  NAND U3929 ( .A(n3757), .B(n3756), .Z(n3758) );
  NAND U3930 ( .A(n3759), .B(n3758), .Z(n3812) );
  XNOR U3931 ( .A(b[7]), .B(a[87]), .Z(n3799) );
  NANDN U3932 ( .A(n3799), .B(n5293), .Z(n3762) );
  NANDN U3933 ( .A(n3760), .B(n5294), .Z(n3761) );
  NAND U3934 ( .A(n3762), .B(n3761), .Z(n3787) );
  XNOR U3935 ( .A(b[3]), .B(a[91]), .Z(n3802) );
  NANDN U3936 ( .A(n3802), .B(n5160), .Z(n3765) );
  NANDN U3937 ( .A(n3763), .B(n5161), .Z(n3764) );
  AND U3938 ( .A(n3765), .B(n3764), .Z(n3788) );
  XNOR U3939 ( .A(n3787), .B(n3788), .Z(n3789) );
  NANDN U3940 ( .A(n292), .B(a[93]), .Z(n3766) );
  XOR U3941 ( .A(n5199), .B(n3766), .Z(n3768) );
  NANDN U3942 ( .A(b[0]), .B(a[92]), .Z(n3767) );
  AND U3943 ( .A(n3768), .B(n3767), .Z(n3795) );
  XNOR U3944 ( .A(b[5]), .B(a[89]), .Z(n3808) );
  NANDN U3945 ( .A(n3808), .B(n5240), .Z(n3771) );
  NANDN U3946 ( .A(n3769), .B(n5241), .Z(n3770) );
  NAND U3947 ( .A(n3771), .B(n3770), .Z(n3793) );
  NANDN U3948 ( .A(n295), .B(a[85]), .Z(n3794) );
  XNOR U3949 ( .A(n3793), .B(n3794), .Z(n3796) );
  XOR U3950 ( .A(n3795), .B(n3796), .Z(n3790) );
  XOR U3951 ( .A(n3789), .B(n3790), .Z(n3811) );
  XOR U3952 ( .A(n3812), .B(n3811), .Z(n3813) );
  XNOR U3953 ( .A(n3814), .B(n3813), .Z(n3783) );
  NAND U3954 ( .A(n3773), .B(n3772), .Z(n3777) );
  NAND U3955 ( .A(n3775), .B(n3774), .Z(n3776) );
  NAND U3956 ( .A(n3777), .B(n3776), .Z(n3784) );
  XNOR U3957 ( .A(n3783), .B(n3784), .Z(n3785) );
  XNOR U3958 ( .A(n3786), .B(n3785), .Z(n3817) );
  XNOR U3959 ( .A(n3817), .B(sreg[213]), .Z(n3819) );
  NAND U3960 ( .A(n3778), .B(sreg[212]), .Z(n3782) );
  OR U3961 ( .A(n3780), .B(n3779), .Z(n3781) );
  AND U3962 ( .A(n3782), .B(n3781), .Z(n3818) );
  XOR U3963 ( .A(n3819), .B(n3818), .Z(c[213]) );
  NANDN U3964 ( .A(n3788), .B(n3787), .Z(n3792) );
  NAND U3965 ( .A(n3790), .B(n3789), .Z(n3791) );
  NAND U3966 ( .A(n3792), .B(n3791), .Z(n3853) );
  NANDN U3967 ( .A(n3794), .B(n3793), .Z(n3798) );
  NAND U3968 ( .A(n3796), .B(n3795), .Z(n3797) );
  NAND U3969 ( .A(n3798), .B(n3797), .Z(n3851) );
  XNOR U3970 ( .A(b[7]), .B(a[88]), .Z(n3838) );
  NANDN U3971 ( .A(n3838), .B(n5293), .Z(n3801) );
  NANDN U3972 ( .A(n3799), .B(n5294), .Z(n3800) );
  NAND U3973 ( .A(n3801), .B(n3800), .Z(n3826) );
  XNOR U3974 ( .A(b[3]), .B(a[92]), .Z(n3841) );
  NANDN U3975 ( .A(n3841), .B(n5160), .Z(n3804) );
  NANDN U3976 ( .A(n3802), .B(n5161), .Z(n3803) );
  AND U3977 ( .A(n3804), .B(n3803), .Z(n3827) );
  XNOR U3978 ( .A(n3826), .B(n3827), .Z(n3828) );
  NANDN U3979 ( .A(n292), .B(a[94]), .Z(n3805) );
  XOR U3980 ( .A(n5199), .B(n3805), .Z(n3807) );
  NANDN U3981 ( .A(b[0]), .B(a[93]), .Z(n3806) );
  AND U3982 ( .A(n3807), .B(n3806), .Z(n3834) );
  XNOR U3983 ( .A(b[5]), .B(a[90]), .Z(n3847) );
  NANDN U3984 ( .A(n3847), .B(n5240), .Z(n3810) );
  NANDN U3985 ( .A(n3808), .B(n5241), .Z(n3809) );
  NAND U3986 ( .A(n3810), .B(n3809), .Z(n3832) );
  NANDN U3987 ( .A(n295), .B(a[86]), .Z(n3833) );
  XNOR U3988 ( .A(n3832), .B(n3833), .Z(n3835) );
  XOR U3989 ( .A(n3834), .B(n3835), .Z(n3829) );
  XOR U3990 ( .A(n3828), .B(n3829), .Z(n3850) );
  XOR U3991 ( .A(n3851), .B(n3850), .Z(n3852) );
  XNOR U3992 ( .A(n3853), .B(n3852), .Z(n3822) );
  NAND U3993 ( .A(n3812), .B(n3811), .Z(n3816) );
  NAND U3994 ( .A(n3814), .B(n3813), .Z(n3815) );
  NAND U3995 ( .A(n3816), .B(n3815), .Z(n3823) );
  XNOR U3996 ( .A(n3822), .B(n3823), .Z(n3824) );
  XNOR U3997 ( .A(n3825), .B(n3824), .Z(n3856) );
  XNOR U3998 ( .A(n3856), .B(sreg[214]), .Z(n3858) );
  NAND U3999 ( .A(n3817), .B(sreg[213]), .Z(n3821) );
  OR U4000 ( .A(n3819), .B(n3818), .Z(n3820) );
  AND U4001 ( .A(n3821), .B(n3820), .Z(n3857) );
  XOR U4002 ( .A(n3858), .B(n3857), .Z(c[214]) );
  NANDN U4003 ( .A(n3827), .B(n3826), .Z(n3831) );
  NAND U4004 ( .A(n3829), .B(n3828), .Z(n3830) );
  NAND U4005 ( .A(n3831), .B(n3830), .Z(n3892) );
  NANDN U4006 ( .A(n3833), .B(n3832), .Z(n3837) );
  NAND U4007 ( .A(n3835), .B(n3834), .Z(n3836) );
  NAND U4008 ( .A(n3837), .B(n3836), .Z(n3890) );
  XNOR U4009 ( .A(b[7]), .B(a[89]), .Z(n3877) );
  NANDN U4010 ( .A(n3877), .B(n5293), .Z(n3840) );
  NANDN U4011 ( .A(n3838), .B(n5294), .Z(n3839) );
  NAND U4012 ( .A(n3840), .B(n3839), .Z(n3865) );
  XNOR U4013 ( .A(b[3]), .B(a[93]), .Z(n3880) );
  NANDN U4014 ( .A(n3880), .B(n5160), .Z(n3843) );
  NANDN U4015 ( .A(n3841), .B(n5161), .Z(n3842) );
  AND U4016 ( .A(n3843), .B(n3842), .Z(n3866) );
  XNOR U4017 ( .A(n3865), .B(n3866), .Z(n3867) );
  NANDN U4018 ( .A(n292), .B(a[95]), .Z(n3844) );
  XOR U4019 ( .A(n5199), .B(n3844), .Z(n3846) );
  IV U4020 ( .A(a[94]), .Z(n4111) );
  NANDN U4021 ( .A(n4111), .B(n292), .Z(n3845) );
  AND U4022 ( .A(n3846), .B(n3845), .Z(n3873) );
  XNOR U4023 ( .A(b[5]), .B(a[91]), .Z(n3886) );
  NANDN U4024 ( .A(n3886), .B(n5240), .Z(n3849) );
  NANDN U4025 ( .A(n3847), .B(n5241), .Z(n3848) );
  NAND U4026 ( .A(n3849), .B(n3848), .Z(n3871) );
  NANDN U4027 ( .A(n295), .B(a[87]), .Z(n3872) );
  XNOR U4028 ( .A(n3871), .B(n3872), .Z(n3874) );
  XOR U4029 ( .A(n3873), .B(n3874), .Z(n3868) );
  XOR U4030 ( .A(n3867), .B(n3868), .Z(n3889) );
  XOR U4031 ( .A(n3890), .B(n3889), .Z(n3891) );
  XNOR U4032 ( .A(n3892), .B(n3891), .Z(n3861) );
  NAND U4033 ( .A(n3851), .B(n3850), .Z(n3855) );
  NAND U4034 ( .A(n3853), .B(n3852), .Z(n3854) );
  NAND U4035 ( .A(n3855), .B(n3854), .Z(n3862) );
  XNOR U4036 ( .A(n3861), .B(n3862), .Z(n3863) );
  XNOR U4037 ( .A(n3864), .B(n3863), .Z(n3895) );
  XNOR U4038 ( .A(n3895), .B(sreg[215]), .Z(n3897) );
  NAND U4039 ( .A(n3856), .B(sreg[214]), .Z(n3860) );
  OR U4040 ( .A(n3858), .B(n3857), .Z(n3859) );
  AND U4041 ( .A(n3860), .B(n3859), .Z(n3896) );
  XOR U4042 ( .A(n3897), .B(n3896), .Z(c[215]) );
  NANDN U4043 ( .A(n3866), .B(n3865), .Z(n3870) );
  NAND U4044 ( .A(n3868), .B(n3867), .Z(n3869) );
  NAND U4045 ( .A(n3870), .B(n3869), .Z(n3931) );
  NANDN U4046 ( .A(n3872), .B(n3871), .Z(n3876) );
  NAND U4047 ( .A(n3874), .B(n3873), .Z(n3875) );
  NAND U4048 ( .A(n3876), .B(n3875), .Z(n3929) );
  XNOR U4049 ( .A(b[7]), .B(a[90]), .Z(n3916) );
  NANDN U4050 ( .A(n3916), .B(n5293), .Z(n3879) );
  NANDN U4051 ( .A(n3877), .B(n5294), .Z(n3878) );
  NAND U4052 ( .A(n3879), .B(n3878), .Z(n3904) );
  XOR U4053 ( .A(b[3]), .B(n4111), .Z(n3919) );
  NANDN U4054 ( .A(n3919), .B(n5160), .Z(n3882) );
  NANDN U4055 ( .A(n3880), .B(n5161), .Z(n3881) );
  AND U4056 ( .A(n3882), .B(n3881), .Z(n3905) );
  XNOR U4057 ( .A(n3904), .B(n3905), .Z(n3906) );
  NANDN U4058 ( .A(n292), .B(a[96]), .Z(n3883) );
  XOR U4059 ( .A(n5199), .B(n3883), .Z(n3885) );
  NANDN U4060 ( .A(b[0]), .B(a[95]), .Z(n3884) );
  AND U4061 ( .A(n3885), .B(n3884), .Z(n3912) );
  XNOR U4062 ( .A(b[5]), .B(a[92]), .Z(n3925) );
  NANDN U4063 ( .A(n3925), .B(n5240), .Z(n3888) );
  NANDN U4064 ( .A(n3886), .B(n5241), .Z(n3887) );
  NAND U4065 ( .A(n3888), .B(n3887), .Z(n3910) );
  NANDN U4066 ( .A(n295), .B(a[88]), .Z(n3911) );
  XNOR U4067 ( .A(n3910), .B(n3911), .Z(n3913) );
  XOR U4068 ( .A(n3912), .B(n3913), .Z(n3907) );
  XOR U4069 ( .A(n3906), .B(n3907), .Z(n3928) );
  XOR U4070 ( .A(n3929), .B(n3928), .Z(n3930) );
  XNOR U4071 ( .A(n3931), .B(n3930), .Z(n3900) );
  NAND U4072 ( .A(n3890), .B(n3889), .Z(n3894) );
  NAND U4073 ( .A(n3892), .B(n3891), .Z(n3893) );
  NAND U4074 ( .A(n3894), .B(n3893), .Z(n3901) );
  XNOR U4075 ( .A(n3900), .B(n3901), .Z(n3902) );
  XNOR U4076 ( .A(n3903), .B(n3902), .Z(n3934) );
  XNOR U4077 ( .A(n3934), .B(sreg[216]), .Z(n3936) );
  NAND U4078 ( .A(n3895), .B(sreg[215]), .Z(n3899) );
  OR U4079 ( .A(n3897), .B(n3896), .Z(n3898) );
  AND U4080 ( .A(n3899), .B(n3898), .Z(n3935) );
  XOR U4081 ( .A(n3936), .B(n3935), .Z(c[216]) );
  NANDN U4082 ( .A(n3905), .B(n3904), .Z(n3909) );
  NAND U4083 ( .A(n3907), .B(n3906), .Z(n3908) );
  NAND U4084 ( .A(n3909), .B(n3908), .Z(n3970) );
  NANDN U4085 ( .A(n3911), .B(n3910), .Z(n3915) );
  NAND U4086 ( .A(n3913), .B(n3912), .Z(n3914) );
  NAND U4087 ( .A(n3915), .B(n3914), .Z(n3968) );
  XNOR U4088 ( .A(b[7]), .B(a[91]), .Z(n3955) );
  NANDN U4089 ( .A(n3955), .B(n5293), .Z(n3918) );
  NANDN U4090 ( .A(n3916), .B(n5294), .Z(n3917) );
  NAND U4091 ( .A(n3918), .B(n3917), .Z(n3943) );
  XNOR U4092 ( .A(b[3]), .B(a[95]), .Z(n3958) );
  NANDN U4093 ( .A(n3958), .B(n5160), .Z(n3921) );
  NANDN U4094 ( .A(n3919), .B(n5161), .Z(n3920) );
  AND U4095 ( .A(n3921), .B(n3920), .Z(n3944) );
  XNOR U4096 ( .A(n3943), .B(n3944), .Z(n3945) );
  NANDN U4097 ( .A(n292), .B(a[97]), .Z(n3922) );
  XOR U4098 ( .A(n5199), .B(n3922), .Z(n3924) );
  NANDN U4099 ( .A(b[0]), .B(a[96]), .Z(n3923) );
  AND U4100 ( .A(n3924), .B(n3923), .Z(n3951) );
  XNOR U4101 ( .A(b[5]), .B(a[93]), .Z(n3964) );
  NANDN U4102 ( .A(n3964), .B(n5240), .Z(n3927) );
  NANDN U4103 ( .A(n3925), .B(n5241), .Z(n3926) );
  NAND U4104 ( .A(n3927), .B(n3926), .Z(n3949) );
  NANDN U4105 ( .A(n295), .B(a[89]), .Z(n3950) );
  XNOR U4106 ( .A(n3949), .B(n3950), .Z(n3952) );
  XOR U4107 ( .A(n3951), .B(n3952), .Z(n3946) );
  XOR U4108 ( .A(n3945), .B(n3946), .Z(n3967) );
  XOR U4109 ( .A(n3968), .B(n3967), .Z(n3969) );
  XNOR U4110 ( .A(n3970), .B(n3969), .Z(n3939) );
  NAND U4111 ( .A(n3929), .B(n3928), .Z(n3933) );
  NAND U4112 ( .A(n3931), .B(n3930), .Z(n3932) );
  NAND U4113 ( .A(n3933), .B(n3932), .Z(n3940) );
  XNOR U4114 ( .A(n3939), .B(n3940), .Z(n3941) );
  XNOR U4115 ( .A(n3942), .B(n3941), .Z(n3973) );
  XNOR U4116 ( .A(n3973), .B(sreg[217]), .Z(n3975) );
  NAND U4117 ( .A(n3934), .B(sreg[216]), .Z(n3938) );
  OR U4118 ( .A(n3936), .B(n3935), .Z(n3937) );
  AND U4119 ( .A(n3938), .B(n3937), .Z(n3974) );
  XOR U4120 ( .A(n3975), .B(n3974), .Z(c[217]) );
  NANDN U4121 ( .A(n3944), .B(n3943), .Z(n3948) );
  NAND U4122 ( .A(n3946), .B(n3945), .Z(n3947) );
  NAND U4123 ( .A(n3948), .B(n3947), .Z(n4009) );
  NANDN U4124 ( .A(n3950), .B(n3949), .Z(n3954) );
  NAND U4125 ( .A(n3952), .B(n3951), .Z(n3953) );
  NAND U4126 ( .A(n3954), .B(n3953), .Z(n4007) );
  XNOR U4127 ( .A(b[7]), .B(a[92]), .Z(n3994) );
  NANDN U4128 ( .A(n3994), .B(n5293), .Z(n3957) );
  NANDN U4129 ( .A(n3955), .B(n5294), .Z(n3956) );
  NAND U4130 ( .A(n3957), .B(n3956), .Z(n3982) );
  XNOR U4131 ( .A(b[3]), .B(a[96]), .Z(n3997) );
  NANDN U4132 ( .A(n3997), .B(n5160), .Z(n3960) );
  NANDN U4133 ( .A(n3958), .B(n5161), .Z(n3959) );
  AND U4134 ( .A(n3960), .B(n3959), .Z(n3983) );
  XNOR U4135 ( .A(n3982), .B(n3983), .Z(n3984) );
  NANDN U4136 ( .A(n292), .B(a[98]), .Z(n3961) );
  XOR U4137 ( .A(n5199), .B(n3961), .Z(n3963) );
  NANDN U4138 ( .A(b[0]), .B(a[97]), .Z(n3962) );
  AND U4139 ( .A(n3963), .B(n3962), .Z(n3990) );
  XOR U4140 ( .A(b[5]), .B(n4111), .Z(n4003) );
  NANDN U4141 ( .A(n4003), .B(n5240), .Z(n3966) );
  NANDN U4142 ( .A(n3964), .B(n5241), .Z(n3965) );
  NAND U4143 ( .A(n3966), .B(n3965), .Z(n3988) );
  NANDN U4144 ( .A(n295), .B(a[90]), .Z(n3989) );
  XNOR U4145 ( .A(n3988), .B(n3989), .Z(n3991) );
  XOR U4146 ( .A(n3990), .B(n3991), .Z(n3985) );
  XOR U4147 ( .A(n3984), .B(n3985), .Z(n4006) );
  XOR U4148 ( .A(n4007), .B(n4006), .Z(n4008) );
  XNOR U4149 ( .A(n4009), .B(n4008), .Z(n3978) );
  NAND U4150 ( .A(n3968), .B(n3967), .Z(n3972) );
  NAND U4151 ( .A(n3970), .B(n3969), .Z(n3971) );
  NAND U4152 ( .A(n3972), .B(n3971), .Z(n3979) );
  XNOR U4153 ( .A(n3978), .B(n3979), .Z(n3980) );
  XNOR U4154 ( .A(n3981), .B(n3980), .Z(n4012) );
  XNOR U4155 ( .A(n4012), .B(sreg[218]), .Z(n4014) );
  NAND U4156 ( .A(n3973), .B(sreg[217]), .Z(n3977) );
  OR U4157 ( .A(n3975), .B(n3974), .Z(n3976) );
  AND U4158 ( .A(n3977), .B(n3976), .Z(n4013) );
  XOR U4159 ( .A(n4014), .B(n4013), .Z(c[218]) );
  NANDN U4160 ( .A(n3983), .B(n3982), .Z(n3987) );
  NAND U4161 ( .A(n3985), .B(n3984), .Z(n3986) );
  NAND U4162 ( .A(n3987), .B(n3986), .Z(n4048) );
  NANDN U4163 ( .A(n3989), .B(n3988), .Z(n3993) );
  NAND U4164 ( .A(n3991), .B(n3990), .Z(n3992) );
  NAND U4165 ( .A(n3993), .B(n3992), .Z(n4046) );
  XNOR U4166 ( .A(b[7]), .B(a[93]), .Z(n4033) );
  NANDN U4167 ( .A(n4033), .B(n5293), .Z(n3996) );
  NANDN U4168 ( .A(n3994), .B(n5294), .Z(n3995) );
  NAND U4169 ( .A(n3996), .B(n3995), .Z(n4021) );
  XNOR U4170 ( .A(b[3]), .B(a[97]), .Z(n4036) );
  NANDN U4171 ( .A(n4036), .B(n5160), .Z(n3999) );
  NANDN U4172 ( .A(n3997), .B(n5161), .Z(n3998) );
  AND U4173 ( .A(n3999), .B(n3998), .Z(n4022) );
  XNOR U4174 ( .A(n4021), .B(n4022), .Z(n4023) );
  NANDN U4175 ( .A(n292), .B(a[99]), .Z(n4000) );
  XOR U4176 ( .A(n5199), .B(n4000), .Z(n4002) );
  NANDN U4177 ( .A(b[0]), .B(a[98]), .Z(n4001) );
  AND U4178 ( .A(n4002), .B(n4001), .Z(n4029) );
  XNOR U4179 ( .A(b[5]), .B(a[95]), .Z(n4042) );
  NANDN U4180 ( .A(n4042), .B(n5240), .Z(n4005) );
  NANDN U4181 ( .A(n4003), .B(n5241), .Z(n4004) );
  NAND U4182 ( .A(n4005), .B(n4004), .Z(n4027) );
  NANDN U4183 ( .A(n295), .B(a[91]), .Z(n4028) );
  XNOR U4184 ( .A(n4027), .B(n4028), .Z(n4030) );
  XOR U4185 ( .A(n4029), .B(n4030), .Z(n4024) );
  XOR U4186 ( .A(n4023), .B(n4024), .Z(n4045) );
  XOR U4187 ( .A(n4046), .B(n4045), .Z(n4047) );
  XNOR U4188 ( .A(n4048), .B(n4047), .Z(n4017) );
  NAND U4189 ( .A(n4007), .B(n4006), .Z(n4011) );
  NAND U4190 ( .A(n4009), .B(n4008), .Z(n4010) );
  NAND U4191 ( .A(n4011), .B(n4010), .Z(n4018) );
  XNOR U4192 ( .A(n4017), .B(n4018), .Z(n4019) );
  XNOR U4193 ( .A(n4020), .B(n4019), .Z(n4051) );
  XNOR U4194 ( .A(n4051), .B(sreg[219]), .Z(n4053) );
  NAND U4195 ( .A(n4012), .B(sreg[218]), .Z(n4016) );
  OR U4196 ( .A(n4014), .B(n4013), .Z(n4015) );
  AND U4197 ( .A(n4016), .B(n4015), .Z(n4052) );
  XOR U4198 ( .A(n4053), .B(n4052), .Z(c[219]) );
  NANDN U4199 ( .A(n4022), .B(n4021), .Z(n4026) );
  NAND U4200 ( .A(n4024), .B(n4023), .Z(n4025) );
  NAND U4201 ( .A(n4026), .B(n4025), .Z(n4087) );
  NANDN U4202 ( .A(n4028), .B(n4027), .Z(n4032) );
  NAND U4203 ( .A(n4030), .B(n4029), .Z(n4031) );
  NAND U4204 ( .A(n4032), .B(n4031), .Z(n4085) );
  XOR U4205 ( .A(b[7]), .B(n4111), .Z(n4072) );
  NANDN U4206 ( .A(n4072), .B(n5293), .Z(n4035) );
  NANDN U4207 ( .A(n4033), .B(n5294), .Z(n4034) );
  NAND U4208 ( .A(n4035), .B(n4034), .Z(n4060) );
  XNOR U4209 ( .A(b[3]), .B(a[98]), .Z(n4075) );
  NANDN U4210 ( .A(n4075), .B(n5160), .Z(n4038) );
  NANDN U4211 ( .A(n4036), .B(n5161), .Z(n4037) );
  AND U4212 ( .A(n4038), .B(n4037), .Z(n4061) );
  XNOR U4213 ( .A(n4060), .B(n4061), .Z(n4062) );
  NANDN U4214 ( .A(n292), .B(a[100]), .Z(n4039) );
  XOR U4215 ( .A(n5199), .B(n4039), .Z(n4041) );
  NANDN U4216 ( .A(b[0]), .B(a[99]), .Z(n4040) );
  AND U4217 ( .A(n4041), .B(n4040), .Z(n4068) );
  XNOR U4218 ( .A(b[5]), .B(a[96]), .Z(n4081) );
  NANDN U4219 ( .A(n4081), .B(n5240), .Z(n4044) );
  NANDN U4220 ( .A(n4042), .B(n5241), .Z(n4043) );
  NAND U4221 ( .A(n4044), .B(n4043), .Z(n4066) );
  NANDN U4222 ( .A(n295), .B(a[92]), .Z(n4067) );
  XNOR U4223 ( .A(n4066), .B(n4067), .Z(n4069) );
  XOR U4224 ( .A(n4068), .B(n4069), .Z(n4063) );
  XOR U4225 ( .A(n4062), .B(n4063), .Z(n4084) );
  XOR U4226 ( .A(n4085), .B(n4084), .Z(n4086) );
  XNOR U4227 ( .A(n4087), .B(n4086), .Z(n4056) );
  NAND U4228 ( .A(n4046), .B(n4045), .Z(n4050) );
  NAND U4229 ( .A(n4048), .B(n4047), .Z(n4049) );
  NAND U4230 ( .A(n4050), .B(n4049), .Z(n4057) );
  XNOR U4231 ( .A(n4056), .B(n4057), .Z(n4058) );
  XNOR U4232 ( .A(n4059), .B(n4058), .Z(n4090) );
  XNOR U4233 ( .A(n4090), .B(sreg[220]), .Z(n4092) );
  NAND U4234 ( .A(n4051), .B(sreg[219]), .Z(n4055) );
  OR U4235 ( .A(n4053), .B(n4052), .Z(n4054) );
  AND U4236 ( .A(n4055), .B(n4054), .Z(n4091) );
  XOR U4237 ( .A(n4092), .B(n4091), .Z(c[220]) );
  NANDN U4238 ( .A(n4061), .B(n4060), .Z(n4065) );
  NAND U4239 ( .A(n4063), .B(n4062), .Z(n4064) );
  NAND U4240 ( .A(n4065), .B(n4064), .Z(n4127) );
  NANDN U4241 ( .A(n4067), .B(n4066), .Z(n4071) );
  NAND U4242 ( .A(n4069), .B(n4068), .Z(n4070) );
  NAND U4243 ( .A(n4071), .B(n4070), .Z(n4125) );
  XNOR U4244 ( .A(b[7]), .B(a[95]), .Z(n4118) );
  NANDN U4245 ( .A(n4118), .B(n5293), .Z(n4074) );
  NANDN U4246 ( .A(n4072), .B(n5294), .Z(n4073) );
  NAND U4247 ( .A(n4074), .B(n4073), .Z(n4099) );
  XNOR U4248 ( .A(b[3]), .B(a[99]), .Z(n4121) );
  NANDN U4249 ( .A(n4121), .B(n5160), .Z(n4077) );
  NANDN U4250 ( .A(n4075), .B(n5161), .Z(n4076) );
  AND U4251 ( .A(n4077), .B(n4076), .Z(n4100) );
  XNOR U4252 ( .A(n4099), .B(n4100), .Z(n4101) );
  NANDN U4253 ( .A(n292), .B(a[101]), .Z(n4078) );
  XOR U4254 ( .A(n5199), .B(n4078), .Z(n4080) );
  NANDN U4255 ( .A(b[0]), .B(a[100]), .Z(n4079) );
  AND U4256 ( .A(n4080), .B(n4079), .Z(n4107) );
  XNOR U4257 ( .A(n294), .B(a[97]), .Z(n4112) );
  NAND U4258 ( .A(n4112), .B(n5240), .Z(n4083) );
  NANDN U4259 ( .A(n4081), .B(n5241), .Z(n4082) );
  NAND U4260 ( .A(n4083), .B(n4082), .Z(n4105) );
  NANDN U4261 ( .A(n295), .B(a[93]), .Z(n4106) );
  XNOR U4262 ( .A(n4105), .B(n4106), .Z(n4108) );
  XOR U4263 ( .A(n4107), .B(n4108), .Z(n4102) );
  XOR U4264 ( .A(n4101), .B(n4102), .Z(n4124) );
  XOR U4265 ( .A(n4125), .B(n4124), .Z(n4126) );
  XNOR U4266 ( .A(n4127), .B(n4126), .Z(n4095) );
  NAND U4267 ( .A(n4085), .B(n4084), .Z(n4089) );
  NAND U4268 ( .A(n4087), .B(n4086), .Z(n4088) );
  NAND U4269 ( .A(n4089), .B(n4088), .Z(n4096) );
  XNOR U4270 ( .A(n4095), .B(n4096), .Z(n4097) );
  XNOR U4271 ( .A(n4098), .B(n4097), .Z(n4130) );
  XNOR U4272 ( .A(n4130), .B(sreg[221]), .Z(n4132) );
  NAND U4273 ( .A(n4090), .B(sreg[220]), .Z(n4094) );
  OR U4274 ( .A(n4092), .B(n4091), .Z(n4093) );
  AND U4275 ( .A(n4094), .B(n4093), .Z(n4131) );
  XOR U4276 ( .A(n4132), .B(n4131), .Z(c[221]) );
  NANDN U4277 ( .A(n4100), .B(n4099), .Z(n4104) );
  NAND U4278 ( .A(n4102), .B(n4101), .Z(n4103) );
  NAND U4279 ( .A(n4104), .B(n4103), .Z(n4166) );
  NANDN U4280 ( .A(n4106), .B(n4105), .Z(n4110) );
  NAND U4281 ( .A(n4108), .B(n4107), .Z(n4109) );
  NAND U4282 ( .A(n4110), .B(n4109), .Z(n4163) );
  ANDN U4283 ( .B(b[7]), .A(n4111), .Z(n4145) );
  XNOR U4284 ( .A(b[5]), .B(a[98]), .Z(n4160) );
  NANDN U4285 ( .A(n4160), .B(n5240), .Z(n4114) );
  NAND U4286 ( .A(n5241), .B(n4112), .Z(n4113) );
  NAND U4287 ( .A(n4114), .B(n4113), .Z(n4146) );
  XOR U4288 ( .A(n4145), .B(n4146), .Z(n4147) );
  NANDN U4289 ( .A(n292), .B(a[102]), .Z(n4115) );
  XOR U4290 ( .A(n5199), .B(n4115), .Z(n4117) );
  NANDN U4291 ( .A(b[0]), .B(a[101]), .Z(n4116) );
  AND U4292 ( .A(n4117), .B(n4116), .Z(n4148) );
  XOR U4293 ( .A(n4147), .B(n4148), .Z(n4142) );
  XNOR U4294 ( .A(b[7]), .B(a[96]), .Z(n4151) );
  NANDN U4295 ( .A(n4151), .B(n5293), .Z(n4120) );
  NANDN U4296 ( .A(n4118), .B(n5294), .Z(n4119) );
  NAND U4297 ( .A(n4120), .B(n4119), .Z(n4139) );
  XNOR U4298 ( .A(b[3]), .B(a[100]), .Z(n4154) );
  NANDN U4299 ( .A(n4154), .B(n5160), .Z(n4123) );
  NANDN U4300 ( .A(n4121), .B(n5161), .Z(n4122) );
  AND U4301 ( .A(n4123), .B(n4122), .Z(n4140) );
  XNOR U4302 ( .A(n4139), .B(n4140), .Z(n4141) );
  XNOR U4303 ( .A(n4142), .B(n4141), .Z(n4164) );
  XNOR U4304 ( .A(n4163), .B(n4164), .Z(n4165) );
  XNOR U4305 ( .A(n4166), .B(n4165), .Z(n4135) );
  NAND U4306 ( .A(n4125), .B(n4124), .Z(n4129) );
  NAND U4307 ( .A(n4127), .B(n4126), .Z(n4128) );
  NAND U4308 ( .A(n4129), .B(n4128), .Z(n4136) );
  XNOR U4309 ( .A(n4135), .B(n4136), .Z(n4137) );
  XNOR U4310 ( .A(n4138), .B(n4137), .Z(n4169) );
  XNOR U4311 ( .A(n4169), .B(sreg[222]), .Z(n4171) );
  NAND U4312 ( .A(n4130), .B(sreg[221]), .Z(n4134) );
  OR U4313 ( .A(n4132), .B(n4131), .Z(n4133) );
  AND U4314 ( .A(n4134), .B(n4133), .Z(n4170) );
  XOR U4315 ( .A(n4171), .B(n4170), .Z(c[222]) );
  NANDN U4316 ( .A(n4140), .B(n4139), .Z(n4144) );
  NAND U4317 ( .A(n4142), .B(n4141), .Z(n4143) );
  NAND U4318 ( .A(n4144), .B(n4143), .Z(n4205) );
  OR U4319 ( .A(n4146), .B(n4145), .Z(n4150) );
  NANDN U4320 ( .A(n4148), .B(n4147), .Z(n4149) );
  NAND U4321 ( .A(n4150), .B(n4149), .Z(n4203) );
  XNOR U4322 ( .A(b[7]), .B(a[97]), .Z(n4190) );
  NANDN U4323 ( .A(n4190), .B(n5293), .Z(n4153) );
  NANDN U4324 ( .A(n4151), .B(n5294), .Z(n4152) );
  NAND U4325 ( .A(n4153), .B(n4152), .Z(n4178) );
  XNOR U4326 ( .A(b[3]), .B(a[101]), .Z(n4193) );
  NANDN U4327 ( .A(n4193), .B(n5160), .Z(n4156) );
  NANDN U4328 ( .A(n4154), .B(n5161), .Z(n4155) );
  AND U4329 ( .A(n4156), .B(n4155), .Z(n4179) );
  XNOR U4330 ( .A(n4178), .B(n4179), .Z(n4180) );
  NANDN U4331 ( .A(n292), .B(a[103]), .Z(n4157) );
  XOR U4332 ( .A(n5199), .B(n4157), .Z(n4159) );
  NANDN U4333 ( .A(b[0]), .B(a[102]), .Z(n4158) );
  AND U4334 ( .A(n4159), .B(n4158), .Z(n4186) );
  XNOR U4335 ( .A(b[5]), .B(a[99]), .Z(n4199) );
  NANDN U4336 ( .A(n4199), .B(n5240), .Z(n4162) );
  NANDN U4337 ( .A(n4160), .B(n5241), .Z(n4161) );
  NAND U4338 ( .A(n4162), .B(n4161), .Z(n4184) );
  NANDN U4339 ( .A(n295), .B(a[95]), .Z(n4185) );
  XNOR U4340 ( .A(n4184), .B(n4185), .Z(n4187) );
  XOR U4341 ( .A(n4186), .B(n4187), .Z(n4181) );
  XOR U4342 ( .A(n4180), .B(n4181), .Z(n4202) );
  XNOR U4343 ( .A(n4203), .B(n4202), .Z(n4204) );
  XNOR U4344 ( .A(n4205), .B(n4204), .Z(n4174) );
  NANDN U4345 ( .A(n4164), .B(n4163), .Z(n4168) );
  NAND U4346 ( .A(n4166), .B(n4165), .Z(n4167) );
  NAND U4347 ( .A(n4168), .B(n4167), .Z(n4175) );
  XNOR U4348 ( .A(n4174), .B(n4175), .Z(n4176) );
  XNOR U4349 ( .A(n4177), .B(n4176), .Z(n4206) );
  XNOR U4350 ( .A(n4206), .B(sreg[223]), .Z(n4208) );
  NAND U4351 ( .A(n4169), .B(sreg[222]), .Z(n4173) );
  OR U4352 ( .A(n4171), .B(n4170), .Z(n4172) );
  AND U4353 ( .A(n4173), .B(n4172), .Z(n4207) );
  XOR U4354 ( .A(n4208), .B(n4207), .Z(c[223]) );
  NANDN U4355 ( .A(n4179), .B(n4178), .Z(n4183) );
  NAND U4356 ( .A(n4181), .B(n4180), .Z(n4182) );
  NAND U4357 ( .A(n4183), .B(n4182), .Z(n4242) );
  NANDN U4358 ( .A(n4185), .B(n4184), .Z(n4189) );
  NAND U4359 ( .A(n4187), .B(n4186), .Z(n4188) );
  NAND U4360 ( .A(n4189), .B(n4188), .Z(n4240) );
  XNOR U4361 ( .A(b[7]), .B(a[98]), .Z(n4227) );
  NANDN U4362 ( .A(n4227), .B(n5293), .Z(n4192) );
  NANDN U4363 ( .A(n4190), .B(n5294), .Z(n4191) );
  NAND U4364 ( .A(n4192), .B(n4191), .Z(n4215) );
  XNOR U4365 ( .A(b[3]), .B(a[102]), .Z(n4230) );
  NANDN U4366 ( .A(n4230), .B(n5160), .Z(n4195) );
  NANDN U4367 ( .A(n4193), .B(n5161), .Z(n4194) );
  AND U4368 ( .A(n4195), .B(n4194), .Z(n4216) );
  XNOR U4369 ( .A(n4215), .B(n4216), .Z(n4217) );
  NANDN U4370 ( .A(n292), .B(a[104]), .Z(n4196) );
  XOR U4371 ( .A(n5199), .B(n4196), .Z(n4198) );
  NANDN U4372 ( .A(b[0]), .B(a[103]), .Z(n4197) );
  AND U4373 ( .A(n4198), .B(n4197), .Z(n4223) );
  XNOR U4374 ( .A(b[5]), .B(a[100]), .Z(n4236) );
  NANDN U4375 ( .A(n4236), .B(n5240), .Z(n4201) );
  NANDN U4376 ( .A(n4199), .B(n5241), .Z(n4200) );
  NAND U4377 ( .A(n4201), .B(n4200), .Z(n4221) );
  NANDN U4378 ( .A(n295), .B(a[96]), .Z(n4222) );
  XNOR U4379 ( .A(n4221), .B(n4222), .Z(n4224) );
  XOR U4380 ( .A(n4223), .B(n4224), .Z(n4218) );
  XOR U4381 ( .A(n4217), .B(n4218), .Z(n4239) );
  XOR U4382 ( .A(n4240), .B(n4239), .Z(n4241) );
  XNOR U4383 ( .A(n4242), .B(n4241), .Z(n4211) );
  XNOR U4384 ( .A(n4211), .B(n4212), .Z(n4213) );
  XNOR U4385 ( .A(n4214), .B(n4213), .Z(n4245) );
  XNOR U4386 ( .A(n4245), .B(sreg[224]), .Z(n4247) );
  NAND U4387 ( .A(n4206), .B(sreg[223]), .Z(n4210) );
  OR U4388 ( .A(n4208), .B(n4207), .Z(n4209) );
  AND U4389 ( .A(n4210), .B(n4209), .Z(n4246) );
  XOR U4390 ( .A(n4247), .B(n4246), .Z(c[224]) );
  NANDN U4391 ( .A(n4216), .B(n4215), .Z(n4220) );
  NAND U4392 ( .A(n4218), .B(n4217), .Z(n4219) );
  NAND U4393 ( .A(n4220), .B(n4219), .Z(n4281) );
  NANDN U4394 ( .A(n4222), .B(n4221), .Z(n4226) );
  NAND U4395 ( .A(n4224), .B(n4223), .Z(n4225) );
  NAND U4396 ( .A(n4226), .B(n4225), .Z(n4279) );
  XNOR U4397 ( .A(b[7]), .B(a[99]), .Z(n4266) );
  NANDN U4398 ( .A(n4266), .B(n5293), .Z(n4229) );
  NANDN U4399 ( .A(n4227), .B(n5294), .Z(n4228) );
  NAND U4400 ( .A(n4229), .B(n4228), .Z(n4254) );
  XNOR U4401 ( .A(b[3]), .B(a[103]), .Z(n4269) );
  NANDN U4402 ( .A(n4269), .B(n5160), .Z(n4232) );
  NANDN U4403 ( .A(n4230), .B(n5161), .Z(n4231) );
  AND U4404 ( .A(n4232), .B(n4231), .Z(n4255) );
  XNOR U4405 ( .A(n4254), .B(n4255), .Z(n4256) );
  NANDN U4406 ( .A(n292), .B(a[105]), .Z(n4233) );
  XOR U4407 ( .A(n5199), .B(n4233), .Z(n4235) );
  NANDN U4408 ( .A(b[0]), .B(a[104]), .Z(n4234) );
  AND U4409 ( .A(n4235), .B(n4234), .Z(n4262) );
  XNOR U4410 ( .A(b[5]), .B(a[101]), .Z(n4275) );
  NANDN U4411 ( .A(n4275), .B(n5240), .Z(n4238) );
  NANDN U4412 ( .A(n4236), .B(n5241), .Z(n4237) );
  NAND U4413 ( .A(n4238), .B(n4237), .Z(n4260) );
  NANDN U4414 ( .A(n295), .B(a[97]), .Z(n4261) );
  XNOR U4415 ( .A(n4260), .B(n4261), .Z(n4263) );
  XOR U4416 ( .A(n4262), .B(n4263), .Z(n4257) );
  XOR U4417 ( .A(n4256), .B(n4257), .Z(n4278) );
  XOR U4418 ( .A(n4279), .B(n4278), .Z(n4280) );
  XNOR U4419 ( .A(n4281), .B(n4280), .Z(n4250) );
  NAND U4420 ( .A(n4240), .B(n4239), .Z(n4244) );
  NAND U4421 ( .A(n4242), .B(n4241), .Z(n4243) );
  NAND U4422 ( .A(n4244), .B(n4243), .Z(n4251) );
  XNOR U4423 ( .A(n4250), .B(n4251), .Z(n4252) );
  XNOR U4424 ( .A(n4253), .B(n4252), .Z(n4284) );
  XNOR U4425 ( .A(n4284), .B(sreg[225]), .Z(n4286) );
  NAND U4426 ( .A(n4245), .B(sreg[224]), .Z(n4249) );
  OR U4427 ( .A(n4247), .B(n4246), .Z(n4248) );
  AND U4428 ( .A(n4249), .B(n4248), .Z(n4285) );
  XOR U4429 ( .A(n4286), .B(n4285), .Z(c[225]) );
  NANDN U4430 ( .A(n4255), .B(n4254), .Z(n4259) );
  NAND U4431 ( .A(n4257), .B(n4256), .Z(n4258) );
  NAND U4432 ( .A(n4259), .B(n4258), .Z(n4320) );
  NANDN U4433 ( .A(n4261), .B(n4260), .Z(n4265) );
  NAND U4434 ( .A(n4263), .B(n4262), .Z(n4264) );
  NAND U4435 ( .A(n4265), .B(n4264), .Z(n4318) );
  XNOR U4436 ( .A(b[7]), .B(a[100]), .Z(n4305) );
  NANDN U4437 ( .A(n4305), .B(n5293), .Z(n4268) );
  NANDN U4438 ( .A(n4266), .B(n5294), .Z(n4267) );
  NAND U4439 ( .A(n4268), .B(n4267), .Z(n4293) );
  XNOR U4440 ( .A(b[3]), .B(a[104]), .Z(n4308) );
  NANDN U4441 ( .A(n4308), .B(n5160), .Z(n4271) );
  NANDN U4442 ( .A(n4269), .B(n5161), .Z(n4270) );
  AND U4443 ( .A(n4271), .B(n4270), .Z(n4294) );
  XNOR U4444 ( .A(n4293), .B(n4294), .Z(n4295) );
  NANDN U4445 ( .A(n292), .B(a[106]), .Z(n4272) );
  XOR U4446 ( .A(n5199), .B(n4272), .Z(n4274) );
  NANDN U4447 ( .A(b[0]), .B(a[105]), .Z(n4273) );
  AND U4448 ( .A(n4274), .B(n4273), .Z(n4301) );
  XNOR U4449 ( .A(b[5]), .B(a[102]), .Z(n4314) );
  NANDN U4450 ( .A(n4314), .B(n5240), .Z(n4277) );
  NANDN U4451 ( .A(n4275), .B(n5241), .Z(n4276) );
  NAND U4452 ( .A(n4277), .B(n4276), .Z(n4299) );
  NANDN U4453 ( .A(n295), .B(a[98]), .Z(n4300) );
  XNOR U4454 ( .A(n4299), .B(n4300), .Z(n4302) );
  XOR U4455 ( .A(n4301), .B(n4302), .Z(n4296) );
  XOR U4456 ( .A(n4295), .B(n4296), .Z(n4317) );
  XOR U4457 ( .A(n4318), .B(n4317), .Z(n4319) );
  XNOR U4458 ( .A(n4320), .B(n4319), .Z(n4289) );
  NAND U4459 ( .A(n4279), .B(n4278), .Z(n4283) );
  NAND U4460 ( .A(n4281), .B(n4280), .Z(n4282) );
  NAND U4461 ( .A(n4283), .B(n4282), .Z(n4290) );
  XNOR U4462 ( .A(n4289), .B(n4290), .Z(n4291) );
  XNOR U4463 ( .A(n4292), .B(n4291), .Z(n4323) );
  XNOR U4464 ( .A(n4323), .B(sreg[226]), .Z(n4325) );
  NAND U4465 ( .A(n4284), .B(sreg[225]), .Z(n4288) );
  OR U4466 ( .A(n4286), .B(n4285), .Z(n4287) );
  AND U4467 ( .A(n4288), .B(n4287), .Z(n4324) );
  XOR U4468 ( .A(n4325), .B(n4324), .Z(c[226]) );
  NANDN U4469 ( .A(n4294), .B(n4293), .Z(n4298) );
  NAND U4470 ( .A(n4296), .B(n4295), .Z(n4297) );
  NAND U4471 ( .A(n4298), .B(n4297), .Z(n4359) );
  NANDN U4472 ( .A(n4300), .B(n4299), .Z(n4304) );
  NAND U4473 ( .A(n4302), .B(n4301), .Z(n4303) );
  NAND U4474 ( .A(n4304), .B(n4303), .Z(n4357) );
  XNOR U4475 ( .A(b[7]), .B(a[101]), .Z(n4350) );
  NANDN U4476 ( .A(n4350), .B(n5293), .Z(n4307) );
  NANDN U4477 ( .A(n4305), .B(n5294), .Z(n4306) );
  NAND U4478 ( .A(n4307), .B(n4306), .Z(n4332) );
  XNOR U4479 ( .A(b[3]), .B(a[105]), .Z(n4353) );
  NANDN U4480 ( .A(n4353), .B(n5160), .Z(n4310) );
  NANDN U4481 ( .A(n4308), .B(n5161), .Z(n4309) );
  AND U4482 ( .A(n4310), .B(n4309), .Z(n4333) );
  XNOR U4483 ( .A(n4332), .B(n4333), .Z(n4334) );
  NANDN U4484 ( .A(n292), .B(a[107]), .Z(n4311) );
  XOR U4485 ( .A(n5199), .B(n4311), .Z(n4313) );
  NANDN U4486 ( .A(b[0]), .B(a[106]), .Z(n4312) );
  AND U4487 ( .A(n4313), .B(n4312), .Z(n4340) );
  XNOR U4488 ( .A(b[5]), .B(a[103]), .Z(n4347) );
  NANDN U4489 ( .A(n4347), .B(n5240), .Z(n4316) );
  NANDN U4490 ( .A(n4314), .B(n5241), .Z(n4315) );
  NAND U4491 ( .A(n4316), .B(n4315), .Z(n4338) );
  NANDN U4492 ( .A(n295), .B(a[99]), .Z(n4339) );
  XNOR U4493 ( .A(n4338), .B(n4339), .Z(n4341) );
  XOR U4494 ( .A(n4340), .B(n4341), .Z(n4335) );
  XOR U4495 ( .A(n4334), .B(n4335), .Z(n4356) );
  XOR U4496 ( .A(n4357), .B(n4356), .Z(n4358) );
  XNOR U4497 ( .A(n4359), .B(n4358), .Z(n4328) );
  NAND U4498 ( .A(n4318), .B(n4317), .Z(n4322) );
  NAND U4499 ( .A(n4320), .B(n4319), .Z(n4321) );
  NAND U4500 ( .A(n4322), .B(n4321), .Z(n4329) );
  XNOR U4501 ( .A(n4328), .B(n4329), .Z(n4330) );
  XNOR U4502 ( .A(n4331), .B(n4330), .Z(n4362) );
  XNOR U4503 ( .A(n4362), .B(sreg[227]), .Z(n4364) );
  NAND U4504 ( .A(n4323), .B(sreg[226]), .Z(n4327) );
  OR U4505 ( .A(n4325), .B(n4324), .Z(n4326) );
  AND U4506 ( .A(n4327), .B(n4326), .Z(n4363) );
  XOR U4507 ( .A(n4364), .B(n4363), .Z(c[227]) );
  NANDN U4508 ( .A(n4333), .B(n4332), .Z(n4337) );
  NAND U4509 ( .A(n4335), .B(n4334), .Z(n4336) );
  NAND U4510 ( .A(n4337), .B(n4336), .Z(n4398) );
  NANDN U4511 ( .A(n4339), .B(n4338), .Z(n4343) );
  NAND U4512 ( .A(n4341), .B(n4340), .Z(n4342) );
  NAND U4513 ( .A(n4343), .B(n4342), .Z(n4396) );
  NANDN U4514 ( .A(n292), .B(a[108]), .Z(n4344) );
  XOR U4515 ( .A(n5199), .B(n4344), .Z(n4346) );
  NANDN U4516 ( .A(b[0]), .B(a[107]), .Z(n4345) );
  AND U4517 ( .A(n4346), .B(n4345), .Z(n4379) );
  XNOR U4518 ( .A(b[5]), .B(a[104]), .Z(n4392) );
  NANDN U4519 ( .A(n4392), .B(n5240), .Z(n4349) );
  NANDN U4520 ( .A(n4347), .B(n5241), .Z(n4348) );
  NAND U4521 ( .A(n4349), .B(n4348), .Z(n4377) );
  NANDN U4522 ( .A(n295), .B(a[100]), .Z(n4378) );
  XNOR U4523 ( .A(n4377), .B(n4378), .Z(n4380) );
  XOR U4524 ( .A(n4379), .B(n4380), .Z(n4373) );
  XNOR U4525 ( .A(b[7]), .B(a[102]), .Z(n4383) );
  NANDN U4526 ( .A(n4383), .B(n5293), .Z(n4352) );
  NANDN U4527 ( .A(n4350), .B(n5294), .Z(n4351) );
  NAND U4528 ( .A(n4352), .B(n4351), .Z(n4371) );
  XNOR U4529 ( .A(b[3]), .B(a[106]), .Z(n4386) );
  NANDN U4530 ( .A(n4386), .B(n5160), .Z(n4355) );
  NANDN U4531 ( .A(n4353), .B(n5161), .Z(n4354) );
  AND U4532 ( .A(n4355), .B(n4354), .Z(n4372) );
  XNOR U4533 ( .A(n4371), .B(n4372), .Z(n4374) );
  XOR U4534 ( .A(n4373), .B(n4374), .Z(n4395) );
  XOR U4535 ( .A(n4396), .B(n4395), .Z(n4397) );
  XNOR U4536 ( .A(n4398), .B(n4397), .Z(n4367) );
  NAND U4537 ( .A(n4357), .B(n4356), .Z(n4361) );
  NAND U4538 ( .A(n4359), .B(n4358), .Z(n4360) );
  NAND U4539 ( .A(n4361), .B(n4360), .Z(n4368) );
  XNOR U4540 ( .A(n4367), .B(n4368), .Z(n4369) );
  XNOR U4541 ( .A(n4370), .B(n4369), .Z(n4401) );
  XNOR U4542 ( .A(n4401), .B(sreg[228]), .Z(n4403) );
  NAND U4543 ( .A(n4362), .B(sreg[227]), .Z(n4366) );
  OR U4544 ( .A(n4364), .B(n4363), .Z(n4365) );
  AND U4545 ( .A(n4366), .B(n4365), .Z(n4402) );
  XOR U4546 ( .A(n4403), .B(n4402), .Z(c[228]) );
  NANDN U4547 ( .A(n4372), .B(n4371), .Z(n4376) );
  NAND U4548 ( .A(n4374), .B(n4373), .Z(n4375) );
  NAND U4549 ( .A(n4376), .B(n4375), .Z(n4437) );
  NANDN U4550 ( .A(n4378), .B(n4377), .Z(n4382) );
  NAND U4551 ( .A(n4380), .B(n4379), .Z(n4381) );
  NAND U4552 ( .A(n4382), .B(n4381), .Z(n4435) );
  XNOR U4553 ( .A(b[7]), .B(a[103]), .Z(n4428) );
  NANDN U4554 ( .A(n4428), .B(n5293), .Z(n4385) );
  NANDN U4555 ( .A(n4383), .B(n5294), .Z(n4384) );
  NAND U4556 ( .A(n4385), .B(n4384), .Z(n4410) );
  XNOR U4557 ( .A(b[3]), .B(a[107]), .Z(n4431) );
  NANDN U4558 ( .A(n4431), .B(n5160), .Z(n4388) );
  NANDN U4559 ( .A(n4386), .B(n5161), .Z(n4387) );
  AND U4560 ( .A(n4388), .B(n4387), .Z(n4411) );
  XNOR U4561 ( .A(n4410), .B(n4411), .Z(n4412) );
  NANDN U4562 ( .A(n292), .B(a[109]), .Z(n4389) );
  XOR U4563 ( .A(n5199), .B(n4389), .Z(n4391) );
  NANDN U4564 ( .A(b[0]), .B(a[108]), .Z(n4390) );
  AND U4565 ( .A(n4391), .B(n4390), .Z(n4418) );
  XNOR U4566 ( .A(n294), .B(a[105]), .Z(n4422) );
  NAND U4567 ( .A(n4422), .B(n5240), .Z(n4394) );
  NANDN U4568 ( .A(n4392), .B(n5241), .Z(n4393) );
  NAND U4569 ( .A(n4394), .B(n4393), .Z(n4416) );
  NANDN U4570 ( .A(n295), .B(a[101]), .Z(n4417) );
  XNOR U4571 ( .A(n4416), .B(n4417), .Z(n4419) );
  XOR U4572 ( .A(n4418), .B(n4419), .Z(n4413) );
  XOR U4573 ( .A(n4412), .B(n4413), .Z(n4434) );
  XOR U4574 ( .A(n4435), .B(n4434), .Z(n4436) );
  XNOR U4575 ( .A(n4437), .B(n4436), .Z(n4406) );
  NAND U4576 ( .A(n4396), .B(n4395), .Z(n4400) );
  NAND U4577 ( .A(n4398), .B(n4397), .Z(n4399) );
  NAND U4578 ( .A(n4400), .B(n4399), .Z(n4407) );
  XNOR U4579 ( .A(n4406), .B(n4407), .Z(n4408) );
  XNOR U4580 ( .A(n4409), .B(n4408), .Z(n4440) );
  XNOR U4581 ( .A(n4440), .B(sreg[229]), .Z(n4442) );
  NAND U4582 ( .A(n4401), .B(sreg[228]), .Z(n4405) );
  OR U4583 ( .A(n4403), .B(n4402), .Z(n4404) );
  AND U4584 ( .A(n4405), .B(n4404), .Z(n4441) );
  XOR U4585 ( .A(n4442), .B(n4441), .Z(c[229]) );
  NANDN U4586 ( .A(n4411), .B(n4410), .Z(n4415) );
  NAND U4587 ( .A(n4413), .B(n4412), .Z(n4414) );
  NAND U4588 ( .A(n4415), .B(n4414), .Z(n4476) );
  NANDN U4589 ( .A(n4417), .B(n4416), .Z(n4421) );
  NAND U4590 ( .A(n4419), .B(n4418), .Z(n4420) );
  NAND U4591 ( .A(n4421), .B(n4420), .Z(n4474) );
  XNOR U4592 ( .A(b[5]), .B(a[106]), .Z(n4458) );
  NANDN U4593 ( .A(n4458), .B(n5240), .Z(n4424) );
  NAND U4594 ( .A(n5241), .B(n4422), .Z(n4423) );
  AND U4595 ( .A(n4424), .B(n4423), .Z(n4467) );
  NANDN U4596 ( .A(n295), .B(a[102]), .Z(n4468) );
  XOR U4597 ( .A(n4467), .B(n4468), .Z(n4470) );
  NANDN U4598 ( .A(n292), .B(a[110]), .Z(n4425) );
  XOR U4599 ( .A(n5199), .B(n4425), .Z(n4427) );
  NANDN U4600 ( .A(b[0]), .B(a[109]), .Z(n4426) );
  AND U4601 ( .A(n4427), .B(n4426), .Z(n4469) );
  XNOR U4602 ( .A(n4470), .B(n4469), .Z(n4464) );
  XNOR U4603 ( .A(b[7]), .B(a[104]), .Z(n4449) );
  NANDN U4604 ( .A(n4449), .B(n5293), .Z(n4430) );
  NANDN U4605 ( .A(n4428), .B(n5294), .Z(n4429) );
  NAND U4606 ( .A(n4430), .B(n4429), .Z(n4461) );
  XNOR U4607 ( .A(b[3]), .B(a[108]), .Z(n4452) );
  NANDN U4608 ( .A(n4452), .B(n5160), .Z(n4433) );
  NANDN U4609 ( .A(n4431), .B(n5161), .Z(n4432) );
  AND U4610 ( .A(n4433), .B(n4432), .Z(n4462) );
  XNOR U4611 ( .A(n4461), .B(n4462), .Z(n4463) );
  XNOR U4612 ( .A(n4464), .B(n4463), .Z(n4473) );
  XOR U4613 ( .A(n4474), .B(n4473), .Z(n4475) );
  XNOR U4614 ( .A(n4476), .B(n4475), .Z(n4445) );
  NAND U4615 ( .A(n4435), .B(n4434), .Z(n4439) );
  NAND U4616 ( .A(n4437), .B(n4436), .Z(n4438) );
  NAND U4617 ( .A(n4439), .B(n4438), .Z(n4446) );
  XNOR U4618 ( .A(n4445), .B(n4446), .Z(n4447) );
  XNOR U4619 ( .A(n4448), .B(n4447), .Z(n4477) );
  XNOR U4620 ( .A(n4477), .B(sreg[230]), .Z(n4479) );
  NAND U4621 ( .A(n4440), .B(sreg[229]), .Z(n4444) );
  OR U4622 ( .A(n4442), .B(n4441), .Z(n4443) );
  AND U4623 ( .A(n4444), .B(n4443), .Z(n4478) );
  XOR U4624 ( .A(n4479), .B(n4478), .Z(c[230]) );
  XNOR U4625 ( .A(b[7]), .B(a[105]), .Z(n4498) );
  NANDN U4626 ( .A(n4498), .B(n5293), .Z(n4451) );
  NANDN U4627 ( .A(n4449), .B(n5294), .Z(n4450) );
  NAND U4628 ( .A(n4451), .B(n4450), .Z(n4486) );
  XNOR U4629 ( .A(b[3]), .B(a[109]), .Z(n4501) );
  NANDN U4630 ( .A(n4501), .B(n5160), .Z(n4454) );
  NANDN U4631 ( .A(n4452), .B(n5161), .Z(n4453) );
  AND U4632 ( .A(n4454), .B(n4453), .Z(n4487) );
  XNOR U4633 ( .A(n4486), .B(n4487), .Z(n4488) );
  NANDN U4634 ( .A(n292), .B(a[111]), .Z(n4455) );
  XOR U4635 ( .A(n5199), .B(n4455), .Z(n4457) );
  NANDN U4636 ( .A(b[0]), .B(a[110]), .Z(n4456) );
  AND U4637 ( .A(n4457), .B(n4456), .Z(n4494) );
  XNOR U4638 ( .A(b[5]), .B(a[107]), .Z(n4507) );
  NANDN U4639 ( .A(n4507), .B(n5240), .Z(n4460) );
  NANDN U4640 ( .A(n4458), .B(n5241), .Z(n4459) );
  NAND U4641 ( .A(n4460), .B(n4459), .Z(n4492) );
  NANDN U4642 ( .A(n295), .B(a[103]), .Z(n4493) );
  XNOR U4643 ( .A(n4492), .B(n4493), .Z(n4495) );
  XOR U4644 ( .A(n4494), .B(n4495), .Z(n4489) );
  XOR U4645 ( .A(n4488), .B(n4489), .Z(n4512) );
  NANDN U4646 ( .A(n4462), .B(n4461), .Z(n4466) );
  NANDN U4647 ( .A(n4464), .B(n4463), .Z(n4465) );
  NAND U4648 ( .A(n4466), .B(n4465), .Z(n4510) );
  OR U4649 ( .A(n4468), .B(n4467), .Z(n4472) );
  NAND U4650 ( .A(n4470), .B(n4469), .Z(n4471) );
  AND U4651 ( .A(n4472), .B(n4471), .Z(n4511) );
  XNOR U4652 ( .A(n4510), .B(n4511), .Z(n4513) );
  XNOR U4653 ( .A(n4512), .B(n4513), .Z(n4482) );
  XNOR U4654 ( .A(n4482), .B(n4483), .Z(n4484) );
  XNOR U4655 ( .A(n4485), .B(n4484), .Z(n4516) );
  XNOR U4656 ( .A(n4516), .B(sreg[231]), .Z(n4518) );
  NAND U4657 ( .A(n4477), .B(sreg[230]), .Z(n4481) );
  OR U4658 ( .A(n4479), .B(n4478), .Z(n4480) );
  AND U4659 ( .A(n4481), .B(n4480), .Z(n4517) );
  XOR U4660 ( .A(n4518), .B(n4517), .Z(c[231]) );
  NANDN U4661 ( .A(n4487), .B(n4486), .Z(n4491) );
  NAND U4662 ( .A(n4489), .B(n4488), .Z(n4490) );
  NAND U4663 ( .A(n4491), .B(n4490), .Z(n4552) );
  NANDN U4664 ( .A(n4493), .B(n4492), .Z(n4497) );
  NAND U4665 ( .A(n4495), .B(n4494), .Z(n4496) );
  NAND U4666 ( .A(n4497), .B(n4496), .Z(n4550) );
  XNOR U4667 ( .A(b[7]), .B(a[106]), .Z(n4537) );
  NANDN U4668 ( .A(n4537), .B(n5293), .Z(n4500) );
  NANDN U4669 ( .A(n4498), .B(n5294), .Z(n4499) );
  NAND U4670 ( .A(n4500), .B(n4499), .Z(n4525) );
  XNOR U4671 ( .A(b[3]), .B(a[110]), .Z(n4540) );
  NANDN U4672 ( .A(n4540), .B(n5160), .Z(n4503) );
  NANDN U4673 ( .A(n4501), .B(n5161), .Z(n4502) );
  AND U4674 ( .A(n4503), .B(n4502), .Z(n4526) );
  XNOR U4675 ( .A(n4525), .B(n4526), .Z(n4527) );
  NANDN U4676 ( .A(n292), .B(a[112]), .Z(n4504) );
  XOR U4677 ( .A(n5199), .B(n4504), .Z(n4506) );
  NANDN U4678 ( .A(b[0]), .B(a[111]), .Z(n4505) );
  AND U4679 ( .A(n4506), .B(n4505), .Z(n4533) );
  XNOR U4680 ( .A(b[5]), .B(a[108]), .Z(n4546) );
  NANDN U4681 ( .A(n4546), .B(n5240), .Z(n4509) );
  NANDN U4682 ( .A(n4507), .B(n5241), .Z(n4508) );
  NAND U4683 ( .A(n4509), .B(n4508), .Z(n4531) );
  NANDN U4684 ( .A(n295), .B(a[104]), .Z(n4532) );
  XNOR U4685 ( .A(n4531), .B(n4532), .Z(n4534) );
  XOR U4686 ( .A(n4533), .B(n4534), .Z(n4528) );
  XOR U4687 ( .A(n4527), .B(n4528), .Z(n4549) );
  XOR U4688 ( .A(n4550), .B(n4549), .Z(n4551) );
  XNOR U4689 ( .A(n4552), .B(n4551), .Z(n4521) );
  NANDN U4690 ( .A(n4511), .B(n4510), .Z(n4515) );
  NAND U4691 ( .A(n4513), .B(n4512), .Z(n4514) );
  NAND U4692 ( .A(n4515), .B(n4514), .Z(n4522) );
  XNOR U4693 ( .A(n4521), .B(n4522), .Z(n4523) );
  XNOR U4694 ( .A(n4524), .B(n4523), .Z(n4555) );
  XNOR U4695 ( .A(n4555), .B(sreg[232]), .Z(n4557) );
  NAND U4696 ( .A(n4516), .B(sreg[231]), .Z(n4520) );
  OR U4697 ( .A(n4518), .B(n4517), .Z(n4519) );
  AND U4698 ( .A(n4520), .B(n4519), .Z(n4556) );
  XOR U4699 ( .A(n4557), .B(n4556), .Z(c[232]) );
  NANDN U4700 ( .A(n4526), .B(n4525), .Z(n4530) );
  NAND U4701 ( .A(n4528), .B(n4527), .Z(n4529) );
  NAND U4702 ( .A(n4530), .B(n4529), .Z(n4591) );
  NANDN U4703 ( .A(n4532), .B(n4531), .Z(n4536) );
  NAND U4704 ( .A(n4534), .B(n4533), .Z(n4535) );
  NAND U4705 ( .A(n4536), .B(n4535), .Z(n4589) );
  XNOR U4706 ( .A(b[7]), .B(a[107]), .Z(n4576) );
  NANDN U4707 ( .A(n4576), .B(n5293), .Z(n4539) );
  NANDN U4708 ( .A(n4537), .B(n5294), .Z(n4538) );
  NAND U4709 ( .A(n4539), .B(n4538), .Z(n4564) );
  XNOR U4710 ( .A(b[3]), .B(a[111]), .Z(n4579) );
  NANDN U4711 ( .A(n4579), .B(n5160), .Z(n4542) );
  NANDN U4712 ( .A(n4540), .B(n5161), .Z(n4541) );
  AND U4713 ( .A(n4542), .B(n4541), .Z(n4565) );
  XNOR U4714 ( .A(n4564), .B(n4565), .Z(n4566) );
  NANDN U4715 ( .A(n292), .B(a[113]), .Z(n4543) );
  XOR U4716 ( .A(n5199), .B(n4543), .Z(n4545) );
  NANDN U4717 ( .A(b[0]), .B(a[112]), .Z(n4544) );
  AND U4718 ( .A(n4545), .B(n4544), .Z(n4572) );
  XNOR U4719 ( .A(b[5]), .B(a[109]), .Z(n4585) );
  NANDN U4720 ( .A(n4585), .B(n5240), .Z(n4548) );
  NANDN U4721 ( .A(n4546), .B(n5241), .Z(n4547) );
  NAND U4722 ( .A(n4548), .B(n4547), .Z(n4570) );
  NANDN U4723 ( .A(n295), .B(a[105]), .Z(n4571) );
  XNOR U4724 ( .A(n4570), .B(n4571), .Z(n4573) );
  XOR U4725 ( .A(n4572), .B(n4573), .Z(n4567) );
  XOR U4726 ( .A(n4566), .B(n4567), .Z(n4588) );
  XOR U4727 ( .A(n4589), .B(n4588), .Z(n4590) );
  XNOR U4728 ( .A(n4591), .B(n4590), .Z(n4560) );
  NAND U4729 ( .A(n4550), .B(n4549), .Z(n4554) );
  NAND U4730 ( .A(n4552), .B(n4551), .Z(n4553) );
  NAND U4731 ( .A(n4554), .B(n4553), .Z(n4561) );
  XNOR U4732 ( .A(n4560), .B(n4561), .Z(n4562) );
  XNOR U4733 ( .A(n4563), .B(n4562), .Z(n4594) );
  XNOR U4734 ( .A(n4594), .B(sreg[233]), .Z(n4596) );
  NAND U4735 ( .A(n4555), .B(sreg[232]), .Z(n4559) );
  OR U4736 ( .A(n4557), .B(n4556), .Z(n4558) );
  AND U4737 ( .A(n4559), .B(n4558), .Z(n4595) );
  XOR U4738 ( .A(n4596), .B(n4595), .Z(c[233]) );
  NANDN U4739 ( .A(n4565), .B(n4564), .Z(n4569) );
  NAND U4740 ( .A(n4567), .B(n4566), .Z(n4568) );
  NAND U4741 ( .A(n4569), .B(n4568), .Z(n4630) );
  NANDN U4742 ( .A(n4571), .B(n4570), .Z(n4575) );
  NAND U4743 ( .A(n4573), .B(n4572), .Z(n4574) );
  NAND U4744 ( .A(n4575), .B(n4574), .Z(n4628) );
  XNOR U4745 ( .A(b[7]), .B(a[108]), .Z(n4615) );
  NANDN U4746 ( .A(n4615), .B(n5293), .Z(n4578) );
  NANDN U4747 ( .A(n4576), .B(n5294), .Z(n4577) );
  NAND U4748 ( .A(n4578), .B(n4577), .Z(n4603) );
  XNOR U4749 ( .A(b[3]), .B(a[112]), .Z(n4618) );
  NANDN U4750 ( .A(n4618), .B(n5160), .Z(n4581) );
  NANDN U4751 ( .A(n4579), .B(n5161), .Z(n4580) );
  AND U4752 ( .A(n4581), .B(n4580), .Z(n4604) );
  XNOR U4753 ( .A(n4603), .B(n4604), .Z(n4605) );
  NANDN U4754 ( .A(n292), .B(a[114]), .Z(n4582) );
  XOR U4755 ( .A(n5199), .B(n4582), .Z(n4584) );
  NANDN U4756 ( .A(b[0]), .B(a[113]), .Z(n4583) );
  AND U4757 ( .A(n4584), .B(n4583), .Z(n4611) );
  XNOR U4758 ( .A(b[5]), .B(a[110]), .Z(n4624) );
  NANDN U4759 ( .A(n4624), .B(n5240), .Z(n4587) );
  NANDN U4760 ( .A(n4585), .B(n5241), .Z(n4586) );
  NAND U4761 ( .A(n4587), .B(n4586), .Z(n4609) );
  NANDN U4762 ( .A(n295), .B(a[106]), .Z(n4610) );
  XNOR U4763 ( .A(n4609), .B(n4610), .Z(n4612) );
  XOR U4764 ( .A(n4611), .B(n4612), .Z(n4606) );
  XOR U4765 ( .A(n4605), .B(n4606), .Z(n4627) );
  XOR U4766 ( .A(n4628), .B(n4627), .Z(n4629) );
  XNOR U4767 ( .A(n4630), .B(n4629), .Z(n4599) );
  NAND U4768 ( .A(n4589), .B(n4588), .Z(n4593) );
  NAND U4769 ( .A(n4591), .B(n4590), .Z(n4592) );
  NAND U4770 ( .A(n4593), .B(n4592), .Z(n4600) );
  XNOR U4771 ( .A(n4599), .B(n4600), .Z(n4601) );
  XNOR U4772 ( .A(n4602), .B(n4601), .Z(n4633) );
  XNOR U4773 ( .A(n4633), .B(sreg[234]), .Z(n4635) );
  NAND U4774 ( .A(n4594), .B(sreg[233]), .Z(n4598) );
  OR U4775 ( .A(n4596), .B(n4595), .Z(n4597) );
  AND U4776 ( .A(n4598), .B(n4597), .Z(n4634) );
  XOR U4777 ( .A(n4635), .B(n4634), .Z(c[234]) );
  NANDN U4778 ( .A(n4604), .B(n4603), .Z(n4608) );
  NAND U4779 ( .A(n4606), .B(n4605), .Z(n4607) );
  NAND U4780 ( .A(n4608), .B(n4607), .Z(n4669) );
  NANDN U4781 ( .A(n4610), .B(n4609), .Z(n4614) );
  NAND U4782 ( .A(n4612), .B(n4611), .Z(n4613) );
  NAND U4783 ( .A(n4614), .B(n4613), .Z(n4667) );
  XNOR U4784 ( .A(b[7]), .B(a[109]), .Z(n4654) );
  NANDN U4785 ( .A(n4654), .B(n5293), .Z(n4617) );
  NANDN U4786 ( .A(n4615), .B(n5294), .Z(n4616) );
  NAND U4787 ( .A(n4617), .B(n4616), .Z(n4642) );
  XNOR U4788 ( .A(b[3]), .B(a[113]), .Z(n4657) );
  NANDN U4789 ( .A(n4657), .B(n5160), .Z(n4620) );
  NANDN U4790 ( .A(n4618), .B(n5161), .Z(n4619) );
  AND U4791 ( .A(n4620), .B(n4619), .Z(n4643) );
  XNOR U4792 ( .A(n4642), .B(n4643), .Z(n4644) );
  NANDN U4793 ( .A(n292), .B(a[115]), .Z(n4621) );
  XOR U4794 ( .A(n5199), .B(n4621), .Z(n4623) );
  NANDN U4795 ( .A(b[0]), .B(a[114]), .Z(n4622) );
  AND U4796 ( .A(n4623), .B(n4622), .Z(n4650) );
  XNOR U4797 ( .A(b[5]), .B(a[111]), .Z(n4663) );
  NANDN U4798 ( .A(n4663), .B(n5240), .Z(n4626) );
  NANDN U4799 ( .A(n4624), .B(n5241), .Z(n4625) );
  NAND U4800 ( .A(n4626), .B(n4625), .Z(n4648) );
  NANDN U4801 ( .A(n295), .B(a[107]), .Z(n4649) );
  XNOR U4802 ( .A(n4648), .B(n4649), .Z(n4651) );
  XOR U4803 ( .A(n4650), .B(n4651), .Z(n4645) );
  XOR U4804 ( .A(n4644), .B(n4645), .Z(n4666) );
  XOR U4805 ( .A(n4667), .B(n4666), .Z(n4668) );
  XNOR U4806 ( .A(n4669), .B(n4668), .Z(n4638) );
  NAND U4807 ( .A(n4628), .B(n4627), .Z(n4632) );
  NAND U4808 ( .A(n4630), .B(n4629), .Z(n4631) );
  NAND U4809 ( .A(n4632), .B(n4631), .Z(n4639) );
  XNOR U4810 ( .A(n4638), .B(n4639), .Z(n4640) );
  XNOR U4811 ( .A(n4641), .B(n4640), .Z(n4672) );
  XNOR U4812 ( .A(n4672), .B(sreg[235]), .Z(n4674) );
  NAND U4813 ( .A(n4633), .B(sreg[234]), .Z(n4637) );
  OR U4814 ( .A(n4635), .B(n4634), .Z(n4636) );
  AND U4815 ( .A(n4637), .B(n4636), .Z(n4673) );
  XOR U4816 ( .A(n4674), .B(n4673), .Z(c[235]) );
  NANDN U4817 ( .A(n4643), .B(n4642), .Z(n4647) );
  NAND U4818 ( .A(n4645), .B(n4644), .Z(n4646) );
  NAND U4819 ( .A(n4647), .B(n4646), .Z(n4708) );
  NANDN U4820 ( .A(n4649), .B(n4648), .Z(n4653) );
  NAND U4821 ( .A(n4651), .B(n4650), .Z(n4652) );
  NAND U4822 ( .A(n4653), .B(n4652), .Z(n4706) );
  XNOR U4823 ( .A(b[7]), .B(a[110]), .Z(n4693) );
  NANDN U4824 ( .A(n4693), .B(n5293), .Z(n4656) );
  NANDN U4825 ( .A(n4654), .B(n5294), .Z(n4655) );
  NAND U4826 ( .A(n4656), .B(n4655), .Z(n4681) );
  XNOR U4827 ( .A(b[3]), .B(a[114]), .Z(n4696) );
  NANDN U4828 ( .A(n4696), .B(n5160), .Z(n4659) );
  NANDN U4829 ( .A(n4657), .B(n5161), .Z(n4658) );
  AND U4830 ( .A(n4659), .B(n4658), .Z(n4682) );
  XNOR U4831 ( .A(n4681), .B(n4682), .Z(n4683) );
  NANDN U4832 ( .A(n292), .B(a[116]), .Z(n4660) );
  XOR U4833 ( .A(n5199), .B(n4660), .Z(n4662) );
  NANDN U4834 ( .A(b[0]), .B(a[115]), .Z(n4661) );
  AND U4835 ( .A(n4662), .B(n4661), .Z(n4689) );
  XNOR U4836 ( .A(b[5]), .B(a[112]), .Z(n4702) );
  NANDN U4837 ( .A(n4702), .B(n5240), .Z(n4665) );
  NANDN U4838 ( .A(n4663), .B(n5241), .Z(n4664) );
  NAND U4839 ( .A(n4665), .B(n4664), .Z(n4687) );
  NANDN U4840 ( .A(n295), .B(a[108]), .Z(n4688) );
  XNOR U4841 ( .A(n4687), .B(n4688), .Z(n4690) );
  XOR U4842 ( .A(n4689), .B(n4690), .Z(n4684) );
  XOR U4843 ( .A(n4683), .B(n4684), .Z(n4705) );
  XOR U4844 ( .A(n4706), .B(n4705), .Z(n4707) );
  XNOR U4845 ( .A(n4708), .B(n4707), .Z(n4677) );
  NAND U4846 ( .A(n4667), .B(n4666), .Z(n4671) );
  NAND U4847 ( .A(n4669), .B(n4668), .Z(n4670) );
  NAND U4848 ( .A(n4671), .B(n4670), .Z(n4678) );
  XNOR U4849 ( .A(n4677), .B(n4678), .Z(n4679) );
  XNOR U4850 ( .A(n4680), .B(n4679), .Z(n4711) );
  XNOR U4851 ( .A(n4711), .B(sreg[236]), .Z(n4713) );
  NAND U4852 ( .A(n4672), .B(sreg[235]), .Z(n4676) );
  OR U4853 ( .A(n4674), .B(n4673), .Z(n4675) );
  AND U4854 ( .A(n4676), .B(n4675), .Z(n4712) );
  XOR U4855 ( .A(n4713), .B(n4712), .Z(c[236]) );
  NANDN U4856 ( .A(n4682), .B(n4681), .Z(n4686) );
  NAND U4857 ( .A(n4684), .B(n4683), .Z(n4685) );
  NAND U4858 ( .A(n4686), .B(n4685), .Z(n4747) );
  NANDN U4859 ( .A(n4688), .B(n4687), .Z(n4692) );
  NAND U4860 ( .A(n4690), .B(n4689), .Z(n4691) );
  NAND U4861 ( .A(n4692), .B(n4691), .Z(n4745) );
  XNOR U4862 ( .A(b[7]), .B(a[111]), .Z(n4732) );
  NANDN U4863 ( .A(n4732), .B(n5293), .Z(n4695) );
  NANDN U4864 ( .A(n4693), .B(n5294), .Z(n4694) );
  NAND U4865 ( .A(n4695), .B(n4694), .Z(n4720) );
  XNOR U4866 ( .A(b[3]), .B(a[115]), .Z(n4735) );
  NANDN U4867 ( .A(n4735), .B(n5160), .Z(n4698) );
  NANDN U4868 ( .A(n4696), .B(n5161), .Z(n4697) );
  AND U4869 ( .A(n4698), .B(n4697), .Z(n4721) );
  XNOR U4870 ( .A(n4720), .B(n4721), .Z(n4722) );
  NANDN U4871 ( .A(n292), .B(a[117]), .Z(n4699) );
  XOR U4872 ( .A(n5199), .B(n4699), .Z(n4701) );
  NANDN U4873 ( .A(b[0]), .B(a[116]), .Z(n4700) );
  AND U4874 ( .A(n4701), .B(n4700), .Z(n4728) );
  XNOR U4875 ( .A(b[5]), .B(a[113]), .Z(n4741) );
  NANDN U4876 ( .A(n4741), .B(n5240), .Z(n4704) );
  NANDN U4877 ( .A(n4702), .B(n5241), .Z(n4703) );
  NAND U4878 ( .A(n4704), .B(n4703), .Z(n4726) );
  NANDN U4879 ( .A(n295), .B(a[109]), .Z(n4727) );
  XNOR U4880 ( .A(n4726), .B(n4727), .Z(n4729) );
  XOR U4881 ( .A(n4728), .B(n4729), .Z(n4723) );
  XOR U4882 ( .A(n4722), .B(n4723), .Z(n4744) );
  XOR U4883 ( .A(n4745), .B(n4744), .Z(n4746) );
  XNOR U4884 ( .A(n4747), .B(n4746), .Z(n4716) );
  NAND U4885 ( .A(n4706), .B(n4705), .Z(n4710) );
  NAND U4886 ( .A(n4708), .B(n4707), .Z(n4709) );
  NAND U4887 ( .A(n4710), .B(n4709), .Z(n4717) );
  XNOR U4888 ( .A(n4716), .B(n4717), .Z(n4718) );
  XNOR U4889 ( .A(n4719), .B(n4718), .Z(n4750) );
  XNOR U4890 ( .A(n4750), .B(sreg[237]), .Z(n4752) );
  NAND U4891 ( .A(n4711), .B(sreg[236]), .Z(n4715) );
  OR U4892 ( .A(n4713), .B(n4712), .Z(n4714) );
  AND U4893 ( .A(n4715), .B(n4714), .Z(n4751) );
  XOR U4894 ( .A(n4752), .B(n4751), .Z(c[237]) );
  NANDN U4895 ( .A(n4721), .B(n4720), .Z(n4725) );
  NAND U4896 ( .A(n4723), .B(n4722), .Z(n4724) );
  NAND U4897 ( .A(n4725), .B(n4724), .Z(n4786) );
  NANDN U4898 ( .A(n4727), .B(n4726), .Z(n4731) );
  NAND U4899 ( .A(n4729), .B(n4728), .Z(n4730) );
  NAND U4900 ( .A(n4731), .B(n4730), .Z(n4784) );
  XNOR U4901 ( .A(b[7]), .B(a[112]), .Z(n4771) );
  NANDN U4902 ( .A(n4771), .B(n5293), .Z(n4734) );
  NANDN U4903 ( .A(n4732), .B(n5294), .Z(n4733) );
  NAND U4904 ( .A(n4734), .B(n4733), .Z(n4759) );
  XNOR U4905 ( .A(b[3]), .B(a[116]), .Z(n4774) );
  NANDN U4906 ( .A(n4774), .B(n5160), .Z(n4737) );
  NANDN U4907 ( .A(n4735), .B(n5161), .Z(n4736) );
  AND U4908 ( .A(n4737), .B(n4736), .Z(n4760) );
  XNOR U4909 ( .A(n4759), .B(n4760), .Z(n4761) );
  NANDN U4910 ( .A(n292), .B(a[118]), .Z(n4738) );
  XOR U4911 ( .A(n5199), .B(n4738), .Z(n4740) );
  NANDN U4912 ( .A(b[0]), .B(a[117]), .Z(n4739) );
  AND U4913 ( .A(n4740), .B(n4739), .Z(n4767) );
  XNOR U4914 ( .A(b[5]), .B(a[114]), .Z(n4780) );
  NANDN U4915 ( .A(n4780), .B(n5240), .Z(n4743) );
  NANDN U4916 ( .A(n4741), .B(n5241), .Z(n4742) );
  NAND U4917 ( .A(n4743), .B(n4742), .Z(n4765) );
  NANDN U4918 ( .A(n295), .B(a[110]), .Z(n4766) );
  XNOR U4919 ( .A(n4765), .B(n4766), .Z(n4768) );
  XOR U4920 ( .A(n4767), .B(n4768), .Z(n4762) );
  XOR U4921 ( .A(n4761), .B(n4762), .Z(n4783) );
  XOR U4922 ( .A(n4784), .B(n4783), .Z(n4785) );
  XNOR U4923 ( .A(n4786), .B(n4785), .Z(n4755) );
  NAND U4924 ( .A(n4745), .B(n4744), .Z(n4749) );
  NAND U4925 ( .A(n4747), .B(n4746), .Z(n4748) );
  NAND U4926 ( .A(n4749), .B(n4748), .Z(n4756) );
  XNOR U4927 ( .A(n4755), .B(n4756), .Z(n4757) );
  XNOR U4928 ( .A(n4758), .B(n4757), .Z(n4789) );
  XNOR U4929 ( .A(n4789), .B(sreg[238]), .Z(n4791) );
  NAND U4930 ( .A(n4750), .B(sreg[237]), .Z(n4754) );
  OR U4931 ( .A(n4752), .B(n4751), .Z(n4753) );
  AND U4932 ( .A(n4754), .B(n4753), .Z(n4790) );
  XOR U4933 ( .A(n4791), .B(n4790), .Z(c[238]) );
  NANDN U4934 ( .A(n4760), .B(n4759), .Z(n4764) );
  NAND U4935 ( .A(n4762), .B(n4761), .Z(n4763) );
  NAND U4936 ( .A(n4764), .B(n4763), .Z(n4825) );
  NANDN U4937 ( .A(n4766), .B(n4765), .Z(n4770) );
  NAND U4938 ( .A(n4768), .B(n4767), .Z(n4769) );
  NAND U4939 ( .A(n4770), .B(n4769), .Z(n4823) );
  XNOR U4940 ( .A(b[7]), .B(a[113]), .Z(n4810) );
  NANDN U4941 ( .A(n4810), .B(n5293), .Z(n4773) );
  NANDN U4942 ( .A(n4771), .B(n5294), .Z(n4772) );
  NAND U4943 ( .A(n4773), .B(n4772), .Z(n4798) );
  XNOR U4944 ( .A(b[3]), .B(a[117]), .Z(n4813) );
  NANDN U4945 ( .A(n4813), .B(n5160), .Z(n4776) );
  NANDN U4946 ( .A(n4774), .B(n5161), .Z(n4775) );
  AND U4947 ( .A(n4776), .B(n4775), .Z(n4799) );
  XNOR U4948 ( .A(n4798), .B(n4799), .Z(n4800) );
  NANDN U4949 ( .A(n292), .B(a[119]), .Z(n4777) );
  XOR U4950 ( .A(n5199), .B(n4777), .Z(n4779) );
  NANDN U4951 ( .A(b[0]), .B(a[118]), .Z(n4778) );
  AND U4952 ( .A(n4779), .B(n4778), .Z(n4806) );
  XNOR U4953 ( .A(b[5]), .B(a[115]), .Z(n4819) );
  NANDN U4954 ( .A(n4819), .B(n5240), .Z(n4782) );
  NANDN U4955 ( .A(n4780), .B(n5241), .Z(n4781) );
  NAND U4956 ( .A(n4782), .B(n4781), .Z(n4804) );
  NANDN U4957 ( .A(n295), .B(a[111]), .Z(n4805) );
  XNOR U4958 ( .A(n4804), .B(n4805), .Z(n4807) );
  XOR U4959 ( .A(n4806), .B(n4807), .Z(n4801) );
  XOR U4960 ( .A(n4800), .B(n4801), .Z(n4822) );
  XOR U4961 ( .A(n4823), .B(n4822), .Z(n4824) );
  XNOR U4962 ( .A(n4825), .B(n4824), .Z(n4794) );
  NAND U4963 ( .A(n4784), .B(n4783), .Z(n4788) );
  NAND U4964 ( .A(n4786), .B(n4785), .Z(n4787) );
  NAND U4965 ( .A(n4788), .B(n4787), .Z(n4795) );
  XNOR U4966 ( .A(n4794), .B(n4795), .Z(n4796) );
  XNOR U4967 ( .A(n4797), .B(n4796), .Z(n4828) );
  XNOR U4968 ( .A(n4828), .B(sreg[239]), .Z(n4830) );
  NAND U4969 ( .A(n4789), .B(sreg[238]), .Z(n4793) );
  OR U4970 ( .A(n4791), .B(n4790), .Z(n4792) );
  AND U4971 ( .A(n4793), .B(n4792), .Z(n4829) );
  XOR U4972 ( .A(n4830), .B(n4829), .Z(c[239]) );
  NANDN U4973 ( .A(n4799), .B(n4798), .Z(n4803) );
  NAND U4974 ( .A(n4801), .B(n4800), .Z(n4802) );
  NAND U4975 ( .A(n4803), .B(n4802), .Z(n4864) );
  NANDN U4976 ( .A(n4805), .B(n4804), .Z(n4809) );
  NAND U4977 ( .A(n4807), .B(n4806), .Z(n4808) );
  NAND U4978 ( .A(n4809), .B(n4808), .Z(n4862) );
  XNOR U4979 ( .A(b[7]), .B(a[114]), .Z(n4849) );
  NANDN U4980 ( .A(n4849), .B(n5293), .Z(n4812) );
  NANDN U4981 ( .A(n4810), .B(n5294), .Z(n4811) );
  NAND U4982 ( .A(n4812), .B(n4811), .Z(n4837) );
  XNOR U4983 ( .A(b[3]), .B(a[118]), .Z(n4852) );
  NANDN U4984 ( .A(n4852), .B(n5160), .Z(n4815) );
  NANDN U4985 ( .A(n4813), .B(n5161), .Z(n4814) );
  AND U4986 ( .A(n4815), .B(n4814), .Z(n4838) );
  XNOR U4987 ( .A(n4837), .B(n4838), .Z(n4839) );
  NANDN U4988 ( .A(n292), .B(a[120]), .Z(n4816) );
  XOR U4989 ( .A(n5199), .B(n4816), .Z(n4818) );
  IV U4990 ( .A(a[119]), .Z(n5083) );
  NANDN U4991 ( .A(n5083), .B(n292), .Z(n4817) );
  AND U4992 ( .A(n4818), .B(n4817), .Z(n4845) );
  XNOR U4993 ( .A(b[5]), .B(a[116]), .Z(n4858) );
  NANDN U4994 ( .A(n4858), .B(n5240), .Z(n4821) );
  NANDN U4995 ( .A(n4819), .B(n5241), .Z(n4820) );
  NAND U4996 ( .A(n4821), .B(n4820), .Z(n4843) );
  NANDN U4997 ( .A(n295), .B(a[112]), .Z(n4844) );
  XNOR U4998 ( .A(n4843), .B(n4844), .Z(n4846) );
  XOR U4999 ( .A(n4845), .B(n4846), .Z(n4840) );
  XOR U5000 ( .A(n4839), .B(n4840), .Z(n4861) );
  XOR U5001 ( .A(n4862), .B(n4861), .Z(n4863) );
  XNOR U5002 ( .A(n4864), .B(n4863), .Z(n4833) );
  NAND U5003 ( .A(n4823), .B(n4822), .Z(n4827) );
  NAND U5004 ( .A(n4825), .B(n4824), .Z(n4826) );
  NAND U5005 ( .A(n4827), .B(n4826), .Z(n4834) );
  XNOR U5006 ( .A(n4833), .B(n4834), .Z(n4835) );
  XNOR U5007 ( .A(n4836), .B(n4835), .Z(n4867) );
  XNOR U5008 ( .A(n4867), .B(sreg[240]), .Z(n4869) );
  NAND U5009 ( .A(n4828), .B(sreg[239]), .Z(n4832) );
  OR U5010 ( .A(n4830), .B(n4829), .Z(n4831) );
  AND U5011 ( .A(n4832), .B(n4831), .Z(n4868) );
  XOR U5012 ( .A(n4869), .B(n4868), .Z(c[240]) );
  NANDN U5013 ( .A(n4838), .B(n4837), .Z(n4842) );
  NAND U5014 ( .A(n4840), .B(n4839), .Z(n4841) );
  NAND U5015 ( .A(n4842), .B(n4841), .Z(n4903) );
  NANDN U5016 ( .A(n4844), .B(n4843), .Z(n4848) );
  NAND U5017 ( .A(n4846), .B(n4845), .Z(n4847) );
  NAND U5018 ( .A(n4848), .B(n4847), .Z(n4901) );
  XNOR U5019 ( .A(b[7]), .B(a[115]), .Z(n4888) );
  NANDN U5020 ( .A(n4888), .B(n5293), .Z(n4851) );
  NANDN U5021 ( .A(n4849), .B(n5294), .Z(n4850) );
  NAND U5022 ( .A(n4851), .B(n4850), .Z(n4876) );
  XOR U5023 ( .A(b[3]), .B(n5083), .Z(n4891) );
  NANDN U5024 ( .A(n4891), .B(n5160), .Z(n4854) );
  NANDN U5025 ( .A(n4852), .B(n5161), .Z(n4853) );
  AND U5026 ( .A(n4854), .B(n4853), .Z(n4877) );
  XNOR U5027 ( .A(n4876), .B(n4877), .Z(n4878) );
  NANDN U5028 ( .A(n292), .B(a[121]), .Z(n4855) );
  XOR U5029 ( .A(n5199), .B(n4855), .Z(n4857) );
  NANDN U5030 ( .A(b[0]), .B(a[120]), .Z(n4856) );
  AND U5031 ( .A(n4857), .B(n4856), .Z(n4884) );
  XNOR U5032 ( .A(b[5]), .B(a[117]), .Z(n4897) );
  NANDN U5033 ( .A(n4897), .B(n5240), .Z(n4860) );
  NANDN U5034 ( .A(n4858), .B(n5241), .Z(n4859) );
  NAND U5035 ( .A(n4860), .B(n4859), .Z(n4882) );
  NANDN U5036 ( .A(n295), .B(a[113]), .Z(n4883) );
  XNOR U5037 ( .A(n4882), .B(n4883), .Z(n4885) );
  XOR U5038 ( .A(n4884), .B(n4885), .Z(n4879) );
  XOR U5039 ( .A(n4878), .B(n4879), .Z(n4900) );
  XOR U5040 ( .A(n4901), .B(n4900), .Z(n4902) );
  XNOR U5041 ( .A(n4903), .B(n4902), .Z(n4872) );
  NAND U5042 ( .A(n4862), .B(n4861), .Z(n4866) );
  NAND U5043 ( .A(n4864), .B(n4863), .Z(n4865) );
  NAND U5044 ( .A(n4866), .B(n4865), .Z(n4873) );
  XNOR U5045 ( .A(n4872), .B(n4873), .Z(n4874) );
  XNOR U5046 ( .A(n4875), .B(n4874), .Z(n4906) );
  XNOR U5047 ( .A(n4906), .B(sreg[241]), .Z(n4908) );
  NAND U5048 ( .A(n4867), .B(sreg[240]), .Z(n4871) );
  OR U5049 ( .A(n4869), .B(n4868), .Z(n4870) );
  AND U5050 ( .A(n4871), .B(n4870), .Z(n4907) );
  XOR U5051 ( .A(n4908), .B(n4907), .Z(c[241]) );
  NANDN U5052 ( .A(n4877), .B(n4876), .Z(n4881) );
  NAND U5053 ( .A(n4879), .B(n4878), .Z(n4880) );
  NAND U5054 ( .A(n4881), .B(n4880), .Z(n4942) );
  NANDN U5055 ( .A(n4883), .B(n4882), .Z(n4887) );
  NAND U5056 ( .A(n4885), .B(n4884), .Z(n4886) );
  NAND U5057 ( .A(n4887), .B(n4886), .Z(n4940) );
  XNOR U5058 ( .A(b[7]), .B(a[116]), .Z(n4927) );
  NANDN U5059 ( .A(n4927), .B(n5293), .Z(n4890) );
  NANDN U5060 ( .A(n4888), .B(n5294), .Z(n4889) );
  NAND U5061 ( .A(n4890), .B(n4889), .Z(n4915) );
  XNOR U5062 ( .A(b[3]), .B(a[120]), .Z(n4930) );
  NANDN U5063 ( .A(n4930), .B(n5160), .Z(n4893) );
  NANDN U5064 ( .A(n4891), .B(n5161), .Z(n4892) );
  AND U5065 ( .A(n4893), .B(n4892), .Z(n4916) );
  XNOR U5066 ( .A(n4915), .B(n4916), .Z(n4917) );
  NANDN U5067 ( .A(n292), .B(a[122]), .Z(n4894) );
  XOR U5068 ( .A(n5199), .B(n4894), .Z(n4896) );
  IV U5069 ( .A(a[121]), .Z(n5093) );
  NANDN U5070 ( .A(n5093), .B(n292), .Z(n4895) );
  AND U5071 ( .A(n4896), .B(n4895), .Z(n4923) );
  XNOR U5072 ( .A(b[5]), .B(a[118]), .Z(n4936) );
  NANDN U5073 ( .A(n4936), .B(n5240), .Z(n4899) );
  NANDN U5074 ( .A(n4897), .B(n5241), .Z(n4898) );
  NAND U5075 ( .A(n4899), .B(n4898), .Z(n4921) );
  NANDN U5076 ( .A(n295), .B(a[114]), .Z(n4922) );
  XNOR U5077 ( .A(n4921), .B(n4922), .Z(n4924) );
  XOR U5078 ( .A(n4923), .B(n4924), .Z(n4918) );
  XOR U5079 ( .A(n4917), .B(n4918), .Z(n4939) );
  XOR U5080 ( .A(n4940), .B(n4939), .Z(n4941) );
  XNOR U5081 ( .A(n4942), .B(n4941), .Z(n4911) );
  NAND U5082 ( .A(n4901), .B(n4900), .Z(n4905) );
  NAND U5083 ( .A(n4903), .B(n4902), .Z(n4904) );
  NAND U5084 ( .A(n4905), .B(n4904), .Z(n4912) );
  XNOR U5085 ( .A(n4911), .B(n4912), .Z(n4913) );
  XNOR U5086 ( .A(n4914), .B(n4913), .Z(n4945) );
  XNOR U5087 ( .A(n4945), .B(sreg[242]), .Z(n4947) );
  NAND U5088 ( .A(n4906), .B(sreg[241]), .Z(n4910) );
  OR U5089 ( .A(n4908), .B(n4907), .Z(n4909) );
  AND U5090 ( .A(n4910), .B(n4909), .Z(n4946) );
  XOR U5091 ( .A(n4947), .B(n4946), .Z(c[242]) );
  NANDN U5092 ( .A(n4916), .B(n4915), .Z(n4920) );
  NAND U5093 ( .A(n4918), .B(n4917), .Z(n4919) );
  NAND U5094 ( .A(n4920), .B(n4919), .Z(n4981) );
  NANDN U5095 ( .A(n4922), .B(n4921), .Z(n4926) );
  NAND U5096 ( .A(n4924), .B(n4923), .Z(n4925) );
  NAND U5097 ( .A(n4926), .B(n4925), .Z(n4979) );
  XNOR U5098 ( .A(b[7]), .B(a[117]), .Z(n4972) );
  NANDN U5099 ( .A(n4972), .B(n5293), .Z(n4929) );
  NANDN U5100 ( .A(n4927), .B(n5294), .Z(n4928) );
  NAND U5101 ( .A(n4929), .B(n4928), .Z(n4954) );
  XOR U5102 ( .A(b[3]), .B(n5093), .Z(n4975) );
  NANDN U5103 ( .A(n4975), .B(n5160), .Z(n4932) );
  NANDN U5104 ( .A(n4930), .B(n5161), .Z(n4931) );
  AND U5105 ( .A(n4932), .B(n4931), .Z(n4955) );
  XNOR U5106 ( .A(n4954), .B(n4955), .Z(n4956) );
  NANDN U5107 ( .A(n292), .B(a[123]), .Z(n4933) );
  XOR U5108 ( .A(n5199), .B(n4933), .Z(n4935) );
  NANDN U5109 ( .A(b[0]), .B(a[122]), .Z(n4934) );
  AND U5110 ( .A(n4935), .B(n4934), .Z(n4962) );
  XOR U5111 ( .A(b[5]), .B(n5083), .Z(n4969) );
  NANDN U5112 ( .A(n4969), .B(n5240), .Z(n4938) );
  NANDN U5113 ( .A(n4936), .B(n5241), .Z(n4937) );
  NAND U5114 ( .A(n4938), .B(n4937), .Z(n4960) );
  NANDN U5115 ( .A(n295), .B(a[115]), .Z(n4961) );
  XNOR U5116 ( .A(n4960), .B(n4961), .Z(n4963) );
  XOR U5117 ( .A(n4962), .B(n4963), .Z(n4957) );
  XOR U5118 ( .A(n4956), .B(n4957), .Z(n4978) );
  XOR U5119 ( .A(n4979), .B(n4978), .Z(n4980) );
  XNOR U5120 ( .A(n4981), .B(n4980), .Z(n4950) );
  NAND U5121 ( .A(n4940), .B(n4939), .Z(n4944) );
  NAND U5122 ( .A(n4942), .B(n4941), .Z(n4943) );
  NAND U5123 ( .A(n4944), .B(n4943), .Z(n4951) );
  XNOR U5124 ( .A(n4950), .B(n4951), .Z(n4952) );
  XNOR U5125 ( .A(n4953), .B(n4952), .Z(n4984) );
  XNOR U5126 ( .A(n4984), .B(sreg[243]), .Z(n4986) );
  NAND U5127 ( .A(n4945), .B(sreg[242]), .Z(n4949) );
  OR U5128 ( .A(n4947), .B(n4946), .Z(n4948) );
  AND U5129 ( .A(n4949), .B(n4948), .Z(n4985) );
  XOR U5130 ( .A(n4986), .B(n4985), .Z(c[243]) );
  NANDN U5131 ( .A(n4955), .B(n4954), .Z(n4959) );
  NAND U5132 ( .A(n4957), .B(n4956), .Z(n4958) );
  NAND U5133 ( .A(n4959), .B(n4958), .Z(n5020) );
  NANDN U5134 ( .A(n4961), .B(n4960), .Z(n4965) );
  NAND U5135 ( .A(n4963), .B(n4962), .Z(n4964) );
  NAND U5136 ( .A(n4965), .B(n4964), .Z(n5018) );
  NANDN U5137 ( .A(n292), .B(a[124]), .Z(n4966) );
  XOR U5138 ( .A(n5199), .B(n4966), .Z(n4968) );
  NANDN U5139 ( .A(b[0]), .B(a[123]), .Z(n4967) );
  AND U5140 ( .A(n4968), .B(n4967), .Z(n5001) );
  XNOR U5141 ( .A(b[5]), .B(a[120]), .Z(n5014) );
  NANDN U5142 ( .A(n5014), .B(n5240), .Z(n4971) );
  NANDN U5143 ( .A(n4969), .B(n5241), .Z(n4970) );
  NAND U5144 ( .A(n4971), .B(n4970), .Z(n4999) );
  NANDN U5145 ( .A(n295), .B(a[116]), .Z(n5000) );
  XNOR U5146 ( .A(n4999), .B(n5000), .Z(n5002) );
  XOR U5147 ( .A(n5001), .B(n5002), .Z(n4995) );
  XNOR U5148 ( .A(b[7]), .B(a[118]), .Z(n5005) );
  NANDN U5149 ( .A(n5005), .B(n5293), .Z(n4974) );
  NANDN U5150 ( .A(n4972), .B(n5294), .Z(n4973) );
  NAND U5151 ( .A(n4974), .B(n4973), .Z(n4993) );
  XNOR U5152 ( .A(b[3]), .B(a[122]), .Z(n5008) );
  NANDN U5153 ( .A(n5008), .B(n5160), .Z(n4977) );
  NANDN U5154 ( .A(n4975), .B(n5161), .Z(n4976) );
  AND U5155 ( .A(n4977), .B(n4976), .Z(n4994) );
  XNOR U5156 ( .A(n4993), .B(n4994), .Z(n4996) );
  XOR U5157 ( .A(n4995), .B(n4996), .Z(n5017) );
  XOR U5158 ( .A(n5018), .B(n5017), .Z(n5019) );
  XNOR U5159 ( .A(n5020), .B(n5019), .Z(n4989) );
  NAND U5160 ( .A(n4979), .B(n4978), .Z(n4983) );
  NAND U5161 ( .A(n4981), .B(n4980), .Z(n4982) );
  NAND U5162 ( .A(n4983), .B(n4982), .Z(n4990) );
  XNOR U5163 ( .A(n4989), .B(n4990), .Z(n4991) );
  XNOR U5164 ( .A(n4992), .B(n4991), .Z(n5023) );
  XNOR U5165 ( .A(n5023), .B(sreg[244]), .Z(n5025) );
  NAND U5166 ( .A(n4984), .B(sreg[243]), .Z(n4988) );
  OR U5167 ( .A(n4986), .B(n4985), .Z(n4987) );
  AND U5168 ( .A(n4988), .B(n4987), .Z(n5024) );
  XOR U5169 ( .A(n5025), .B(n5024), .Z(c[244]) );
  NANDN U5170 ( .A(n4994), .B(n4993), .Z(n4998) );
  NAND U5171 ( .A(n4996), .B(n4995), .Z(n4997) );
  NAND U5172 ( .A(n4998), .B(n4997), .Z(n5059) );
  NANDN U5173 ( .A(n5000), .B(n4999), .Z(n5004) );
  NAND U5174 ( .A(n5002), .B(n5001), .Z(n5003) );
  NAND U5175 ( .A(n5004), .B(n5003), .Z(n5057) );
  XOR U5176 ( .A(b[7]), .B(n5083), .Z(n5050) );
  NANDN U5177 ( .A(n5050), .B(n5293), .Z(n5007) );
  NANDN U5178 ( .A(n5005), .B(n5294), .Z(n5006) );
  NAND U5179 ( .A(n5007), .B(n5006), .Z(n5032) );
  XNOR U5180 ( .A(b[3]), .B(a[123]), .Z(n5053) );
  NANDN U5181 ( .A(n5053), .B(n5160), .Z(n5010) );
  NANDN U5182 ( .A(n5008), .B(n5161), .Z(n5009) );
  AND U5183 ( .A(n5010), .B(n5009), .Z(n5033) );
  XNOR U5184 ( .A(n5032), .B(n5033), .Z(n5034) );
  IV U5185 ( .A(a[125]), .Z(n5236) );
  NANDN U5186 ( .A(n5236), .B(b[0]), .Z(n5011) );
  XOR U5187 ( .A(n5199), .B(n5011), .Z(n5013) );
  IV U5188 ( .A(a[124]), .Z(n5204) );
  NANDN U5189 ( .A(n5204), .B(n292), .Z(n5012) );
  AND U5190 ( .A(n5013), .B(n5012), .Z(n5040) );
  XOR U5191 ( .A(b[5]), .B(n5093), .Z(n5047) );
  NANDN U5192 ( .A(n5047), .B(n5240), .Z(n5016) );
  NANDN U5193 ( .A(n5014), .B(n5241), .Z(n5015) );
  NAND U5194 ( .A(n5016), .B(n5015), .Z(n5038) );
  NANDN U5195 ( .A(n295), .B(a[117]), .Z(n5039) );
  XNOR U5196 ( .A(n5038), .B(n5039), .Z(n5041) );
  XOR U5197 ( .A(n5040), .B(n5041), .Z(n5035) );
  XOR U5198 ( .A(n5034), .B(n5035), .Z(n5056) );
  XOR U5199 ( .A(n5057), .B(n5056), .Z(n5058) );
  XNOR U5200 ( .A(n5059), .B(n5058), .Z(n5028) );
  NAND U5201 ( .A(n5018), .B(n5017), .Z(n5022) );
  NAND U5202 ( .A(n5020), .B(n5019), .Z(n5021) );
  NAND U5203 ( .A(n5022), .B(n5021), .Z(n5029) );
  XNOR U5204 ( .A(n5028), .B(n5029), .Z(n5030) );
  XNOR U5205 ( .A(n5031), .B(n5030), .Z(n5062) );
  XNOR U5206 ( .A(n5062), .B(sreg[245]), .Z(n5064) );
  NAND U5207 ( .A(n5023), .B(sreg[244]), .Z(n5027) );
  OR U5208 ( .A(n5025), .B(n5024), .Z(n5026) );
  AND U5209 ( .A(n5027), .B(n5026), .Z(n5063) );
  XOR U5210 ( .A(n5064), .B(n5063), .Z(c[245]) );
  NANDN U5211 ( .A(n5033), .B(n5032), .Z(n5037) );
  NAND U5212 ( .A(n5035), .B(n5034), .Z(n5036) );
  NAND U5213 ( .A(n5037), .B(n5036), .Z(n5100) );
  NANDN U5214 ( .A(n5039), .B(n5038), .Z(n5043) );
  NAND U5215 ( .A(n5041), .B(n5040), .Z(n5042) );
  NAND U5216 ( .A(n5043), .B(n5042), .Z(n5098) );
  IV U5217 ( .A(a[126]), .Z(n5208) );
  NANDN U5218 ( .A(n5208), .B(b[0]), .Z(n5044) );
  XOR U5219 ( .A(n5199), .B(n5044), .Z(n5046) );
  NANDN U5220 ( .A(n5236), .B(n292), .Z(n5045) );
  AND U5221 ( .A(n5046), .B(n5045), .Z(n5079) );
  XNOR U5222 ( .A(n294), .B(a[122]), .Z(n5087) );
  NAND U5223 ( .A(n5087), .B(n5240), .Z(n5049) );
  NANDN U5224 ( .A(n5047), .B(n5241), .Z(n5048) );
  NAND U5225 ( .A(n5049), .B(n5048), .Z(n5077) );
  NANDN U5226 ( .A(n295), .B(a[118]), .Z(n5078) );
  XNOR U5227 ( .A(n5077), .B(n5078), .Z(n5080) );
  XOR U5228 ( .A(n5079), .B(n5080), .Z(n5073) );
  XNOR U5229 ( .A(b[7]), .B(a[120]), .Z(n5094) );
  NANDN U5230 ( .A(n5094), .B(n5293), .Z(n5052) );
  NANDN U5231 ( .A(n5050), .B(n5294), .Z(n5051) );
  NAND U5232 ( .A(n5052), .B(n5051), .Z(n5071) );
  XOR U5233 ( .A(b[3]), .B(n5204), .Z(n5090) );
  NANDN U5234 ( .A(n5090), .B(n5160), .Z(n5055) );
  NANDN U5235 ( .A(n5053), .B(n5161), .Z(n5054) );
  AND U5236 ( .A(n5055), .B(n5054), .Z(n5072) );
  XNOR U5237 ( .A(n5071), .B(n5072), .Z(n5074) );
  XOR U5238 ( .A(n5073), .B(n5074), .Z(n5097) );
  XOR U5239 ( .A(n5098), .B(n5097), .Z(n5099) );
  XNOR U5240 ( .A(n5100), .B(n5099), .Z(n5067) );
  NAND U5241 ( .A(n5057), .B(n5056), .Z(n5061) );
  NAND U5242 ( .A(n5059), .B(n5058), .Z(n5060) );
  NAND U5243 ( .A(n5061), .B(n5060), .Z(n5068) );
  XNOR U5244 ( .A(n5067), .B(n5068), .Z(n5069) );
  XNOR U5245 ( .A(n5070), .B(n5069), .Z(n5103) );
  XNOR U5246 ( .A(n5103), .B(sreg[246]), .Z(n5105) );
  NAND U5247 ( .A(n5062), .B(sreg[245]), .Z(n5066) );
  OR U5248 ( .A(n5064), .B(n5063), .Z(n5065) );
  AND U5249 ( .A(n5066), .B(n5065), .Z(n5104) );
  XOR U5250 ( .A(n5105), .B(n5104), .Z(c[246]) );
  NANDN U5251 ( .A(n5072), .B(n5071), .Z(n5076) );
  NAND U5252 ( .A(n5074), .B(n5073), .Z(n5075) );
  NAND U5253 ( .A(n5076), .B(n5075), .Z(n5120) );
  NANDN U5254 ( .A(n5078), .B(n5077), .Z(n5082) );
  NAND U5255 ( .A(n5080), .B(n5079), .Z(n5081) );
  NAND U5256 ( .A(n5082), .B(n5081), .Z(n5118) );
  ANDN U5257 ( .B(b[7]), .A(n5083), .Z(n5132) );
  NANDN U5258 ( .A(n292), .B(a[127]), .Z(n5084) );
  XOR U5259 ( .A(n5199), .B(n5084), .Z(n5086) );
  NANDN U5260 ( .A(n5208), .B(n292), .Z(n5085) );
  AND U5261 ( .A(n5086), .B(n5085), .Z(n5130) );
  XOR U5262 ( .A(n294), .B(a[123]), .Z(n5143) );
  NANDN U5263 ( .A(n5143), .B(n5240), .Z(n5089) );
  NAND U5264 ( .A(n5241), .B(n5087), .Z(n5088) );
  AND U5265 ( .A(n5089), .B(n5088), .Z(n5129) );
  XNOR U5266 ( .A(n5130), .B(n5129), .Z(n5131) );
  XOR U5267 ( .A(n5132), .B(n5131), .Z(n5126) );
  XOR U5268 ( .A(b[3]), .B(n5236), .Z(n5138) );
  NANDN U5269 ( .A(n5138), .B(n5160), .Z(n5092) );
  NANDN U5270 ( .A(n5090), .B(n5161), .Z(n5091) );
  NAND U5271 ( .A(n5092), .B(n5091), .Z(n5123) );
  XOR U5272 ( .A(b[7]), .B(n5093), .Z(n5135) );
  NANDN U5273 ( .A(n5135), .B(n5293), .Z(n5096) );
  NANDN U5274 ( .A(n5094), .B(n5294), .Z(n5095) );
  AND U5275 ( .A(n5096), .B(n5095), .Z(n5124) );
  XNOR U5276 ( .A(n5123), .B(n5124), .Z(n5125) );
  XOR U5277 ( .A(n5126), .B(n5125), .Z(n5117) );
  XOR U5278 ( .A(n5118), .B(n5117), .Z(n5119) );
  XNOR U5279 ( .A(n5120), .B(n5119), .Z(n5113) );
  NAND U5280 ( .A(n5098), .B(n5097), .Z(n5102) );
  NAND U5281 ( .A(n5100), .B(n5099), .Z(n5101) );
  NAND U5282 ( .A(n5102), .B(n5101), .Z(n5114) );
  XNOR U5283 ( .A(n5113), .B(n5114), .Z(n5115) );
  XNOR U5284 ( .A(n5116), .B(n5115), .Z(n5108) );
  XNOR U5285 ( .A(n5108), .B(sreg[247]), .Z(n5110) );
  NAND U5286 ( .A(n5103), .B(sreg[246]), .Z(n5107) );
  OR U5287 ( .A(n5105), .B(n5104), .Z(n5106) );
  AND U5288 ( .A(n5107), .B(n5106), .Z(n5109) );
  XOR U5289 ( .A(n5110), .B(n5109), .Z(c[247]) );
  NAND U5290 ( .A(n5108), .B(sreg[247]), .Z(n5112) );
  OR U5291 ( .A(n5110), .B(n5109), .Z(n5111) );
  AND U5292 ( .A(n5112), .B(n5111), .Z(n5147) );
  NAND U5293 ( .A(n5118), .B(n5117), .Z(n5122) );
  NAND U5294 ( .A(n5120), .B(n5119), .Z(n5121) );
  NAND U5295 ( .A(n5122), .B(n5121), .Z(n5148) );
  NANDN U5296 ( .A(n5124), .B(n5123), .Z(n5128) );
  NAND U5297 ( .A(n5126), .B(n5125), .Z(n5127) );
  NAND U5298 ( .A(n5128), .B(n5127), .Z(n5180) );
  NANDN U5299 ( .A(n5130), .B(n5129), .Z(n5134) );
  NANDN U5300 ( .A(n5132), .B(n5131), .Z(n5133) );
  NAND U5301 ( .A(n5134), .B(n5133), .Z(n5177) );
  XNOR U5302 ( .A(b[7]), .B(a[122]), .Z(n5154) );
  NANDN U5303 ( .A(n5154), .B(n5293), .Z(n5137) );
  NANDN U5304 ( .A(n5135), .B(n5294), .Z(n5136) );
  NAND U5305 ( .A(n5137), .B(n5136), .Z(n5168) );
  XOR U5306 ( .A(b[3]), .B(n5208), .Z(n5162) );
  NANDN U5307 ( .A(n5162), .B(n5160), .Z(n5140) );
  NANDN U5308 ( .A(n5138), .B(n5161), .Z(n5139) );
  NAND U5309 ( .A(n5140), .B(n5139), .Z(n5165) );
  NANDN U5310 ( .A(n292), .B(b[1]), .Z(n5142) );
  OR U5311 ( .A(a[127]), .B(n5199), .Z(n5141) );
  AND U5312 ( .A(n5142), .B(n5141), .Z(n5171) );
  NANDN U5313 ( .A(n295), .B(a[120]), .Z(n5172) );
  XNOR U5314 ( .A(n5171), .B(n5172), .Z(n5173) );
  XOR U5315 ( .A(b[5]), .B(n5204), .Z(n5157) );
  NANDN U5316 ( .A(n5157), .B(n5240), .Z(n5145) );
  NANDN U5317 ( .A(n5143), .B(n5241), .Z(n5144) );
  AND U5318 ( .A(n5145), .B(n5144), .Z(n5174) );
  XNOR U5319 ( .A(n5165), .B(n5166), .Z(n5167) );
  XOR U5320 ( .A(n5168), .B(n5167), .Z(n5178) );
  XNOR U5321 ( .A(n5177), .B(n5178), .Z(n5179) );
  XOR U5322 ( .A(n5180), .B(n5179), .Z(n5149) );
  XOR U5323 ( .A(n5148), .B(n5149), .Z(n5150) );
  XOR U5324 ( .A(n5151), .B(n5150), .Z(n5146) );
  XOR U5325 ( .A(n5147), .B(n5146), .Z(c[248]) );
  OR U5326 ( .A(n5147), .B(n5146), .Z(n5220) );
  OR U5327 ( .A(n5149), .B(n5148), .Z(n5153) );
  NAND U5328 ( .A(n5151), .B(n5150), .Z(n5152) );
  NAND U5329 ( .A(n5153), .B(n5152), .Z(n5215) );
  ANDN U5330 ( .B(a[121]), .A(n295), .Z(n5249) );
  IV U5331 ( .A(n5249), .Z(n5280) );
  XNOR U5332 ( .A(b[7]), .B(a[123]), .Z(n5205) );
  NANDN U5333 ( .A(n5205), .B(n5293), .Z(n5156) );
  NANDN U5334 ( .A(n5154), .B(n5294), .Z(n5155) );
  AND U5335 ( .A(n5156), .B(n5155), .Z(n5194) );
  XOR U5336 ( .A(n5280), .B(n5194), .Z(n5196) );
  XOR U5337 ( .A(b[5]), .B(n5236), .Z(n5209) );
  NANDN U5338 ( .A(n5209), .B(n5240), .Z(n5159) );
  NANDN U5339 ( .A(n5157), .B(n5241), .Z(n5158) );
  AND U5340 ( .A(n5159), .B(n5158), .Z(n5195) );
  XOR U5341 ( .A(n5196), .B(n5195), .Z(n5191) );
  XNOR U5342 ( .A(a[127]), .B(n293), .Z(n5201) );
  NAND U5343 ( .A(n5201), .B(n5160), .Z(n5164) );
  NANDN U5344 ( .A(n5162), .B(n5161), .Z(n5163) );
  AND U5345 ( .A(n5164), .B(n5163), .Z(n5189) );
  XNOR U5346 ( .A(n5199), .B(n5189), .Z(n5190) );
  XNOR U5347 ( .A(n5191), .B(n5190), .Z(n5186) );
  NANDN U5348 ( .A(n5166), .B(n5165), .Z(n5170) );
  NAND U5349 ( .A(n5168), .B(n5167), .Z(n5169) );
  NAND U5350 ( .A(n5170), .B(n5169), .Z(n5183) );
  OR U5351 ( .A(n5172), .B(n5171), .Z(n5176) );
  OR U5352 ( .A(n5174), .B(n5173), .Z(n5175) );
  AND U5353 ( .A(n5176), .B(n5175), .Z(n5184) );
  XNOR U5354 ( .A(n5183), .B(n5184), .Z(n5185) );
  XOR U5355 ( .A(n5186), .B(n5185), .Z(n5212) );
  NANDN U5356 ( .A(n5178), .B(n5177), .Z(n5182) );
  NANDN U5357 ( .A(n5180), .B(n5179), .Z(n5181) );
  AND U5358 ( .A(n5182), .B(n5181), .Z(n5213) );
  XNOR U5359 ( .A(n5212), .B(n5213), .Z(n5214) );
  XOR U5360 ( .A(n5215), .B(n5214), .Z(n5219) );
  XOR U5361 ( .A(n5220), .B(n5219), .Z(c[249]) );
  NANDN U5362 ( .A(n5184), .B(n5183), .Z(n5188) );
  NANDN U5363 ( .A(n5186), .B(n5185), .Z(n5187) );
  NAND U5364 ( .A(n5188), .B(n5187), .Z(n5223) );
  OR U5365 ( .A(n5189), .B(b[1]), .Z(n5193) );
  NAND U5366 ( .A(n5191), .B(n5190), .Z(n5192) );
  NAND U5367 ( .A(n5193), .B(n5192), .Z(n5229) );
  NANDN U5368 ( .A(n5280), .B(n5194), .Z(n5198) );
  NANDN U5369 ( .A(n5196), .B(n5195), .Z(n5197) );
  NAND U5370 ( .A(n5198), .B(n5197), .Z(n5227) );
  NANDN U5371 ( .A(n5199), .B(b[2]), .Z(n5245) );
  XOR U5372 ( .A(n293), .B(n5245), .Z(n5203) );
  XOR U5373 ( .A(b[2]), .B(n5199), .Z(n5200) );
  NANDN U5374 ( .A(n5201), .B(n5200), .Z(n5202) );
  AND U5375 ( .A(n5203), .B(n5202), .Z(n5246) );
  NANDN U5376 ( .A(n295), .B(a[122]), .Z(n5247) );
  XNOR U5377 ( .A(n5246), .B(n5247), .Z(n5248) );
  XOR U5378 ( .A(n5280), .B(n5248), .Z(n5232) );
  XOR U5379 ( .A(b[7]), .B(n5204), .Z(n5237) );
  NANDN U5380 ( .A(n5237), .B(n5293), .Z(n5207) );
  NANDN U5381 ( .A(n5205), .B(n5294), .Z(n5206) );
  NAND U5382 ( .A(n5207), .B(n5206), .Z(n5230) );
  XOR U5383 ( .A(b[5]), .B(n5208), .Z(n5242) );
  NANDN U5384 ( .A(n5242), .B(n5240), .Z(n5211) );
  NANDN U5385 ( .A(n5209), .B(n5241), .Z(n5210) );
  AND U5386 ( .A(n5211), .B(n5210), .Z(n5231) );
  XNOR U5387 ( .A(n5230), .B(n5231), .Z(n5233) );
  XNOR U5388 ( .A(n5232), .B(n5233), .Z(n5226) );
  XOR U5389 ( .A(n5227), .B(n5226), .Z(n5228) );
  XOR U5390 ( .A(n5229), .B(n5228), .Z(n5224) );
  NANDN U5391 ( .A(n5213), .B(n5212), .Z(n5217) );
  NAND U5392 ( .A(n5215), .B(n5214), .Z(n5216) );
  AND U5393 ( .A(n5217), .B(n5216), .Z(n5225) );
  XOR U5394 ( .A(n5224), .B(n5225), .Z(n5218) );
  XNOR U5395 ( .A(n5223), .B(n5218), .Z(n5222) );
  OR U5396 ( .A(n5220), .B(n5219), .Z(n5221) );
  XOR U5397 ( .A(n5222), .B(n5221), .Z(c[250]) );
  OR U5398 ( .A(n5222), .B(n5221), .Z(n5285) );
  NANDN U5399 ( .A(n5231), .B(n5230), .Z(n5235) );
  NAND U5400 ( .A(n5233), .B(n5232), .Z(n5234) );
  NAND U5401 ( .A(n5235), .B(n5234), .Z(n5259) );
  XOR U5402 ( .A(n295), .B(n5236), .Z(n5274) );
  NAND U5403 ( .A(n5274), .B(n5293), .Z(n5239) );
  NANDN U5404 ( .A(n5237), .B(n5294), .Z(n5238) );
  NAND U5405 ( .A(n5239), .B(n5238), .Z(n5262) );
  XNOR U5406 ( .A(n294), .B(a[127]), .Z(n5271) );
  NAND U5407 ( .A(n5271), .B(n5240), .Z(n5244) );
  NANDN U5408 ( .A(n5242), .B(n5241), .Z(n5243) );
  AND U5409 ( .A(n5244), .B(n5243), .Z(n5263) );
  XNOR U5410 ( .A(n5262), .B(n5263), .Z(n5264) );
  ANDN U5411 ( .B(n5245), .A(n293), .Z(n5278) );
  NANDN U5412 ( .A(n295), .B(a[123]), .Z(n5277) );
  XOR U5413 ( .A(n5278), .B(n5277), .Z(n5279) );
  XOR U5414 ( .A(n5280), .B(n5279), .Z(n5265) );
  XOR U5415 ( .A(n5264), .B(n5265), .Z(n5256) );
  NANDN U5416 ( .A(n5247), .B(n5246), .Z(n5251) );
  NANDN U5417 ( .A(n5249), .B(n5248), .Z(n5250) );
  NAND U5418 ( .A(n5251), .B(n5250), .Z(n5257) );
  XNOR U5419 ( .A(n5256), .B(n5257), .Z(n5258) );
  XNOR U5420 ( .A(n5259), .B(n5258), .Z(n5253) );
  XNOR U5421 ( .A(n5254), .B(n5253), .Z(n5252) );
  XNOR U5422 ( .A(n5255), .B(n5252), .Z(n5284) );
  XOR U5423 ( .A(n5285), .B(n5284), .Z(c[251]) );
  NANDN U5424 ( .A(n5257), .B(n5256), .Z(n5261) );
  NANDN U5425 ( .A(n5259), .B(n5258), .Z(n5260) );
  AND U5426 ( .A(n5261), .B(n5260), .Z(n5300) );
  NANDN U5427 ( .A(n5263), .B(n5262), .Z(n5267) );
  NANDN U5428 ( .A(n5265), .B(n5264), .Z(n5266) );
  NAND U5429 ( .A(n5267), .B(n5266), .Z(n5308) );
  XOR U5430 ( .A(n294), .B(n5268), .Z(n5273) );
  XOR U5431 ( .A(n5269), .B(b[3]), .Z(n5270) );
  NANDN U5432 ( .A(n5271), .B(n5270), .Z(n5272) );
  AND U5433 ( .A(n5273), .B(n5272), .Z(n5288) );
  AND U5434 ( .A(a[124]), .B(b[7]), .Z(n5319) );
  XNOR U5435 ( .A(n5288), .B(n5319), .Z(n5289) );
  XOR U5436 ( .A(n295), .B(a[126]), .Z(n5295) );
  NANDN U5437 ( .A(n5295), .B(n5293), .Z(n5276) );
  NAND U5438 ( .A(n5294), .B(n5274), .Z(n5275) );
  NAND U5439 ( .A(n5276), .B(n5275), .Z(n5290) );
  XOR U5440 ( .A(n5289), .B(n5290), .Z(n5305) );
  OR U5441 ( .A(n5278), .B(n5277), .Z(n5282) );
  NANDN U5442 ( .A(n5280), .B(n5279), .Z(n5281) );
  AND U5443 ( .A(n5282), .B(n5281), .Z(n5306) );
  XNOR U5444 ( .A(n5305), .B(n5306), .Z(n5307) );
  XOR U5445 ( .A(n5308), .B(n5307), .Z(n5299) );
  IV U5446 ( .A(n5299), .Z(n5298) );
  XOR U5447 ( .A(n5300), .B(n5298), .Z(n5283) );
  XNOR U5448 ( .A(n5302), .B(n5283), .Z(n5287) );
  OR U5449 ( .A(n5285), .B(n5284), .Z(n5286) );
  XOR U5450 ( .A(n5287), .B(n5286), .Z(c[252]) );
  OR U5451 ( .A(n5287), .B(n5286), .Z(n5335) );
  NANDN U5452 ( .A(n295), .B(a[125]), .Z(n5318) );
  XNOR U5453 ( .A(n5317), .B(n5318), .Z(n5320) );
  NANDN U5454 ( .A(n5288), .B(n5319), .Z(n5292) );
  NANDN U5455 ( .A(n5290), .B(n5289), .Z(n5291) );
  NAND U5456 ( .A(n5292), .B(n5291), .Z(n5328) );
  XNOR U5457 ( .A(b[7]), .B(a[127]), .Z(n5313) );
  NANDN U5458 ( .A(n5313), .B(n5293), .Z(n5297) );
  NANDN U5459 ( .A(n5295), .B(n5294), .Z(n5296) );
  NAND U5460 ( .A(n5297), .B(n5296), .Z(n5327) );
  XNOR U5461 ( .A(n5328), .B(n5327), .Z(n5329) );
  XOR U5462 ( .A(n5330), .B(n5329), .Z(n5324) );
  NANDN U5463 ( .A(n5298), .B(n5300), .Z(n5304) );
  OR U5464 ( .A(n5300), .B(n5299), .Z(n5301) );
  NANDN U5465 ( .A(n5302), .B(n5301), .Z(n5303) );
  NAND U5466 ( .A(n5304), .B(n5303), .Z(n5326) );
  NANDN U5467 ( .A(n5306), .B(n5305), .Z(n5310) );
  NAND U5468 ( .A(n5308), .B(n5307), .Z(n5309) );
  NAND U5469 ( .A(n5310), .B(n5309), .Z(n5325) );
  XOR U5470 ( .A(n5326), .B(n5325), .Z(n5311) );
  XNOR U5471 ( .A(n5324), .B(n5311), .Z(n5334) );
  XNOR U5472 ( .A(n5335), .B(n5334), .Z(c[253]) );
  NANDN U5473 ( .A(n294), .B(b[6]), .Z(n5312) );
  XOR U5474 ( .A(n295), .B(n5312), .Z(n5316) );
  XOR U5475 ( .A(n5336), .B(b[5]), .Z(n5314) );
  NAND U5476 ( .A(n5314), .B(n5313), .Z(n5315) );
  AND U5477 ( .A(n5316), .B(n5315), .Z(n5342) );
  IV U5478 ( .A(n5342), .Z(n5340) );
  OR U5479 ( .A(n5318), .B(n5317), .Z(n5322) );
  NANDN U5480 ( .A(n5320), .B(n5319), .Z(n5321) );
  NAND U5481 ( .A(n5322), .B(n5321), .Z(n5343) );
  AND U5482 ( .A(b[7]), .B(a[126]), .Z(n5341) );
  XNOR U5483 ( .A(n5343), .B(n5341), .Z(n5323) );
  XOR U5484 ( .A(n5340), .B(n5323), .Z(n5339) );
  NANDN U5485 ( .A(n5328), .B(n5327), .Z(n5332) );
  NANDN U5486 ( .A(n5330), .B(n5329), .Z(n5331) );
  NAND U5487 ( .A(n5332), .B(n5331), .Z(n5337) );
  XOR U5488 ( .A(n5338), .B(n5337), .Z(n5333) );
  XNOR U5489 ( .A(n5339), .B(n5333), .Z(n5344) );
  NANDN U5490 ( .A(n5335), .B(n5334), .Z(n5345) );
  XNOR U5491 ( .A(n5344), .B(n5345), .Z(c[254]) );
endmodule

