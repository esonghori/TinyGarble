
module aes_seq_CC10 ( clk, rst, msg, key, out );
  input [127:0] msg;
  input [127:0] key;
  output [127:0] out;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460;
  wire   [127:0] state;

  DFF \state_reg[127]  ( .D(state[127]), .CLK(clk), .RST(rst), .I(msg[127]), 
        .Q(state[127]) );
  DFF \state_reg[126]  ( .D(state[126]), .CLK(clk), .RST(rst), .I(msg[126]), 
        .Q(state[126]) );
  DFF \state_reg[125]  ( .D(state[125]), .CLK(clk), .RST(rst), .I(msg[125]), 
        .Q(state[125]) );
  DFF \state_reg[124]  ( .D(state[124]), .CLK(clk), .RST(rst), .I(msg[124]), 
        .Q(state[124]) );
  DFF \state_reg[123]  ( .D(state[123]), .CLK(clk), .RST(rst), .I(msg[123]), 
        .Q(state[123]) );
  DFF \state_reg[122]  ( .D(state[122]), .CLK(clk), .RST(rst), .I(msg[122]), 
        .Q(state[122]) );
  DFF \state_reg[121]  ( .D(state[121]), .CLK(clk), .RST(rst), .I(msg[121]), 
        .Q(state[121]) );
  DFF \state_reg[120]  ( .D(state[120]), .CLK(clk), .RST(rst), .I(msg[120]), 
        .Q(state[120]) );
  DFF \state_reg[119]  ( .D(state[119]), .CLK(clk), .RST(rst), .I(msg[119]), 
        .Q(state[119]) );
  DFF \state_reg[118]  ( .D(state[118]), .CLK(clk), .RST(rst), .I(msg[118]), 
        .Q(state[118]) );
  DFF \state_reg[117]  ( .D(state[117]), .CLK(clk), .RST(rst), .I(msg[117]), 
        .Q(state[117]) );
  DFF \state_reg[116]  ( .D(state[116]), .CLK(clk), .RST(rst), .I(msg[116]), 
        .Q(state[116]) );
  DFF \state_reg[115]  ( .D(state[115]), .CLK(clk), .RST(rst), .I(msg[115]), 
        .Q(state[115]) );
  DFF \state_reg[114]  ( .D(state[114]), .CLK(clk), .RST(rst), .I(msg[114]), 
        .Q(state[114]) );
  DFF \state_reg[113]  ( .D(state[113]), .CLK(clk), .RST(rst), .I(msg[113]), 
        .Q(state[113]) );
  DFF \state_reg[112]  ( .D(state[112]), .CLK(clk), .RST(rst), .I(msg[112]), 
        .Q(state[112]) );
  DFF \state_reg[111]  ( .D(state[111]), .CLK(clk), .RST(rst), .I(msg[111]), 
        .Q(state[111]) );
  DFF \state_reg[110]  ( .D(state[110]), .CLK(clk), .RST(rst), .I(msg[110]), 
        .Q(state[110]) );
  DFF \state_reg[109]  ( .D(state[109]), .CLK(clk), .RST(rst), .I(msg[109]), 
        .Q(state[109]) );
  DFF \state_reg[108]  ( .D(state[108]), .CLK(clk), .RST(rst), .I(msg[108]), 
        .Q(state[108]) );
  DFF \state_reg[107]  ( .D(state[107]), .CLK(clk), .RST(rst), .I(msg[107]), 
        .Q(state[107]) );
  DFF \state_reg[106]  ( .D(state[106]), .CLK(clk), .RST(rst), .I(msg[106]), 
        .Q(state[106]) );
  DFF \state_reg[105]  ( .D(state[105]), .CLK(clk), .RST(rst), .I(msg[105]), 
        .Q(state[105]) );
  DFF \state_reg[104]  ( .D(state[104]), .CLK(clk), .RST(rst), .I(msg[104]), 
        .Q(state[104]) );
  DFF \state_reg[103]  ( .D(state[103]), .CLK(clk), .RST(rst), .I(msg[103]), 
        .Q(state[103]) );
  DFF \state_reg[102]  ( .D(state[102]), .CLK(clk), .RST(rst), .I(msg[102]), 
        .Q(state[102]) );
  DFF \state_reg[101]  ( .D(state[101]), .CLK(clk), .RST(rst), .I(msg[101]), 
        .Q(state[101]) );
  DFF \state_reg[100]  ( .D(state[100]), .CLK(clk), .RST(rst), .I(msg[100]), 
        .Q(state[100]) );
  DFF \state_reg[99]  ( .D(state[99]), .CLK(clk), .RST(rst), .I(msg[99]), .Q(
        state[99]) );
  DFF \state_reg[98]  ( .D(state[98]), .CLK(clk), .RST(rst), .I(msg[98]), .Q(
        state[98]) );
  DFF \state_reg[97]  ( .D(state[97]), .CLK(clk), .RST(rst), .I(msg[97]), .Q(
        state[97]) );
  DFF \state_reg[96]  ( .D(state[96]), .CLK(clk), .RST(rst), .I(msg[96]), .Q(
        state[96]) );
  DFF \state_reg[95]  ( .D(state[95]), .CLK(clk), .RST(rst), .I(msg[95]), .Q(
        state[95]) );
  DFF \state_reg[94]  ( .D(state[94]), .CLK(clk), .RST(rst), .I(msg[94]), .Q(
        state[94]) );
  DFF \state_reg[93]  ( .D(state[93]), .CLK(clk), .RST(rst), .I(msg[93]), .Q(
        state[93]) );
  DFF \state_reg[92]  ( .D(state[92]), .CLK(clk), .RST(rst), .I(msg[92]), .Q(
        state[92]) );
  DFF \state_reg[91]  ( .D(state[91]), .CLK(clk), .RST(rst), .I(msg[91]), .Q(
        state[91]) );
  DFF \state_reg[90]  ( .D(state[90]), .CLK(clk), .RST(rst), .I(msg[90]), .Q(
        state[90]) );
  DFF \state_reg[89]  ( .D(state[89]), .CLK(clk), .RST(rst), .I(msg[89]), .Q(
        state[89]) );
  DFF \state_reg[88]  ( .D(state[88]), .CLK(clk), .RST(rst), .I(msg[88]), .Q(
        state[88]) );
  DFF \state_reg[87]  ( .D(state[87]), .CLK(clk), .RST(rst), .I(msg[87]), .Q(
        state[87]) );
  DFF \state_reg[86]  ( .D(state[86]), .CLK(clk), .RST(rst), .I(msg[86]), .Q(
        state[86]) );
  DFF \state_reg[85]  ( .D(state[85]), .CLK(clk), .RST(rst), .I(msg[85]), .Q(
        state[85]) );
  DFF \state_reg[84]  ( .D(state[84]), .CLK(clk), .RST(rst), .I(msg[84]), .Q(
        state[84]) );
  DFF \state_reg[83]  ( .D(state[83]), .CLK(clk), .RST(rst), .I(msg[83]), .Q(
        state[83]) );
  DFF \state_reg[82]  ( .D(state[82]), .CLK(clk), .RST(rst), .I(msg[82]), .Q(
        state[82]) );
  DFF \state_reg[81]  ( .D(state[81]), .CLK(clk), .RST(rst), .I(msg[81]), .Q(
        state[81]) );
  DFF \state_reg[80]  ( .D(state[80]), .CLK(clk), .RST(rst), .I(msg[80]), .Q(
        state[80]) );
  DFF \state_reg[79]  ( .D(state[79]), .CLK(clk), .RST(rst), .I(msg[79]), .Q(
        state[79]) );
  DFF \state_reg[78]  ( .D(state[78]), .CLK(clk), .RST(rst), .I(msg[78]), .Q(
        state[78]) );
  DFF \state_reg[77]  ( .D(state[77]), .CLK(clk), .RST(rst), .I(msg[77]), .Q(
        state[77]) );
  DFF \state_reg[76]  ( .D(state[76]), .CLK(clk), .RST(rst), .I(msg[76]), .Q(
        state[76]) );
  DFF \state_reg[75]  ( .D(state[75]), .CLK(clk), .RST(rst), .I(msg[75]), .Q(
        state[75]) );
  DFF \state_reg[74]  ( .D(state[74]), .CLK(clk), .RST(rst), .I(msg[74]), .Q(
        state[74]) );
  DFF \state_reg[73]  ( .D(state[73]), .CLK(clk), .RST(rst), .I(msg[73]), .Q(
        state[73]) );
  DFF \state_reg[72]  ( .D(state[72]), .CLK(clk), .RST(rst), .I(msg[72]), .Q(
        state[72]) );
  DFF \state_reg[71]  ( .D(state[71]), .CLK(clk), .RST(rst), .I(msg[71]), .Q(
        state[71]) );
  DFF \state_reg[70]  ( .D(state[70]), .CLK(clk), .RST(rst), .I(msg[70]), .Q(
        state[70]) );
  DFF \state_reg[69]  ( .D(state[69]), .CLK(clk), .RST(rst), .I(msg[69]), .Q(
        state[69]) );
  DFF \state_reg[68]  ( .D(state[68]), .CLK(clk), .RST(rst), .I(msg[68]), .Q(
        state[68]) );
  DFF \state_reg[67]  ( .D(state[67]), .CLK(clk), .RST(rst), .I(msg[67]), .Q(
        state[67]) );
  DFF \state_reg[66]  ( .D(state[66]), .CLK(clk), .RST(rst), .I(msg[66]), .Q(
        state[66]) );
  DFF \state_reg[65]  ( .D(state[65]), .CLK(clk), .RST(rst), .I(msg[65]), .Q(
        state[65]) );
  DFF \state_reg[64]  ( .D(state[64]), .CLK(clk), .RST(rst), .I(msg[64]), .Q(
        state[64]) );
  DFF \state_reg[63]  ( .D(state[63]), .CLK(clk), .RST(rst), .I(msg[63]), .Q(
        state[63]) );
  DFF \state_reg[62]  ( .D(state[62]), .CLK(clk), .RST(rst), .I(msg[62]), .Q(
        state[62]) );
  DFF \state_reg[61]  ( .D(state[61]), .CLK(clk), .RST(rst), .I(msg[61]), .Q(
        state[61]) );
  DFF \state_reg[60]  ( .D(state[60]), .CLK(clk), .RST(rst), .I(msg[60]), .Q(
        state[60]) );
  DFF \state_reg[59]  ( .D(state[59]), .CLK(clk), .RST(rst), .I(msg[59]), .Q(
        state[59]) );
  DFF \state_reg[58]  ( .D(state[58]), .CLK(clk), .RST(rst), .I(msg[58]), .Q(
        state[58]) );
  DFF \state_reg[57]  ( .D(state[57]), .CLK(clk), .RST(rst), .I(msg[57]), .Q(
        state[57]) );
  DFF \state_reg[56]  ( .D(state[56]), .CLK(clk), .RST(rst), .I(msg[56]), .Q(
        state[56]) );
  DFF \state_reg[55]  ( .D(state[55]), .CLK(clk), .RST(rst), .I(msg[55]), .Q(
        state[55]) );
  DFF \state_reg[54]  ( .D(state[54]), .CLK(clk), .RST(rst), .I(msg[54]), .Q(
        state[54]) );
  DFF \state_reg[53]  ( .D(state[53]), .CLK(clk), .RST(rst), .I(msg[53]), .Q(
        state[53]) );
  DFF \state_reg[52]  ( .D(state[52]), .CLK(clk), .RST(rst), .I(msg[52]), .Q(
        state[52]) );
  DFF \state_reg[51]  ( .D(state[51]), .CLK(clk), .RST(rst), .I(msg[51]), .Q(
        state[51]) );
  DFF \state_reg[50]  ( .D(state[50]), .CLK(clk), .RST(rst), .I(msg[50]), .Q(
        state[50]) );
  DFF \state_reg[49]  ( .D(state[49]), .CLK(clk), .RST(rst), .I(msg[49]), .Q(
        state[49]) );
  DFF \state_reg[48]  ( .D(state[48]), .CLK(clk), .RST(rst), .I(msg[48]), .Q(
        state[48]) );
  DFF \state_reg[47]  ( .D(state[47]), .CLK(clk), .RST(rst), .I(msg[47]), .Q(
        state[47]) );
  DFF \state_reg[46]  ( .D(state[46]), .CLK(clk), .RST(rst), .I(msg[46]), .Q(
        state[46]) );
  DFF \state_reg[45]  ( .D(state[45]), .CLK(clk), .RST(rst), .I(msg[45]), .Q(
        state[45]) );
  DFF \state_reg[44]  ( .D(state[44]), .CLK(clk), .RST(rst), .I(msg[44]), .Q(
        state[44]) );
  DFF \state_reg[43]  ( .D(state[43]), .CLK(clk), .RST(rst), .I(msg[43]), .Q(
        state[43]) );
  DFF \state_reg[42]  ( .D(state[42]), .CLK(clk), .RST(rst), .I(msg[42]), .Q(
        state[42]) );
  DFF \state_reg[41]  ( .D(state[41]), .CLK(clk), .RST(rst), .I(msg[41]), .Q(
        state[41]) );
  DFF \state_reg[40]  ( .D(state[40]), .CLK(clk), .RST(rst), .I(msg[40]), .Q(
        state[40]) );
  DFF \state_reg[39]  ( .D(state[39]), .CLK(clk), .RST(rst), .I(msg[39]), .Q(
        state[39]) );
  DFF \state_reg[38]  ( .D(state[38]), .CLK(clk), .RST(rst), .I(msg[38]), .Q(
        state[38]) );
  DFF \state_reg[37]  ( .D(state[37]), .CLK(clk), .RST(rst), .I(msg[37]), .Q(
        state[37]) );
  DFF \state_reg[36]  ( .D(state[36]), .CLK(clk), .RST(rst), .I(msg[36]), .Q(
        state[36]) );
  DFF \state_reg[35]  ( .D(state[35]), .CLK(clk), .RST(rst), .I(msg[35]), .Q(
        state[35]) );
  DFF \state_reg[34]  ( .D(state[34]), .CLK(clk), .RST(rst), .I(msg[34]), .Q(
        state[34]) );
  DFF \state_reg[33]  ( .D(state[33]), .CLK(clk), .RST(rst), .I(msg[33]), .Q(
        state[33]) );
  DFF \state_reg[32]  ( .D(state[32]), .CLK(clk), .RST(rst), .I(msg[32]), .Q(
        state[32]) );
  DFF \state_reg[31]  ( .D(state[31]), .CLK(clk), .RST(rst), .I(msg[31]), .Q(
        state[31]) );
  DFF \state_reg[30]  ( .D(state[30]), .CLK(clk), .RST(rst), .I(msg[30]), .Q(
        state[30]) );
  DFF \state_reg[29]  ( .D(state[29]), .CLK(clk), .RST(rst), .I(msg[29]), .Q(
        state[29]) );
  DFF \state_reg[28]  ( .D(state[28]), .CLK(clk), .RST(rst), .I(msg[28]), .Q(
        state[28]) );
  DFF \state_reg[27]  ( .D(state[27]), .CLK(clk), .RST(rst), .I(msg[27]), .Q(
        state[27]) );
  DFF \state_reg[26]  ( .D(state[26]), .CLK(clk), .RST(rst), .I(msg[26]), .Q(
        state[26]) );
  DFF \state_reg[25]  ( .D(state[25]), .CLK(clk), .RST(rst), .I(msg[25]), .Q(
        state[25]) );
  DFF \state_reg[24]  ( .D(state[24]), .CLK(clk), .RST(rst), .I(msg[24]), .Q(
        state[24]) );
  DFF \state_reg[23]  ( .D(state[23]), .CLK(clk), .RST(rst), .I(msg[23]), .Q(
        state[23]) );
  DFF \state_reg[22]  ( .D(state[22]), .CLK(clk), .RST(rst), .I(msg[22]), .Q(
        state[22]) );
  DFF \state_reg[21]  ( .D(state[21]), .CLK(clk), .RST(rst), .I(msg[21]), .Q(
        state[21]) );
  DFF \state_reg[20]  ( .D(state[20]), .CLK(clk), .RST(rst), .I(msg[20]), .Q(
        state[20]) );
  DFF \state_reg[19]  ( .D(state[19]), .CLK(clk), .RST(rst), .I(msg[19]), .Q(
        state[19]) );
  DFF \state_reg[18]  ( .D(state[18]), .CLK(clk), .RST(rst), .I(msg[18]), .Q(
        state[18]) );
  DFF \state_reg[17]  ( .D(state[17]), .CLK(clk), .RST(rst), .I(msg[17]), .Q(
        state[17]) );
  DFF \state_reg[16]  ( .D(state[16]), .CLK(clk), .RST(rst), .I(msg[16]), .Q(
        state[16]) );
  DFF \state_reg[15]  ( .D(state[15]), .CLK(clk), .RST(rst), .I(msg[15]), .Q(
        state[15]) );
  DFF \state_reg[14]  ( .D(state[14]), .CLK(clk), .RST(rst), .I(msg[14]), .Q(
        state[14]) );
  DFF \state_reg[13]  ( .D(state[13]), .CLK(clk), .RST(rst), .I(msg[13]), .Q(
        state[13]) );
  DFF \state_reg[12]  ( .D(state[12]), .CLK(clk), .RST(rst), .I(msg[12]), .Q(
        state[12]) );
  DFF \state_reg[11]  ( .D(state[11]), .CLK(clk), .RST(rst), .I(msg[11]), .Q(
        state[11]) );
  DFF \state_reg[10]  ( .D(state[10]), .CLK(clk), .RST(rst), .I(msg[10]), .Q(
        state[10]) );
  DFF \state_reg[9]  ( .D(state[9]), .CLK(clk), .RST(rst), .I(msg[9]), .Q(
        state[9]) );
  DFF \state_reg[8]  ( .D(state[8]), .CLK(clk), .RST(rst), .I(msg[8]), .Q(
        state[8]) );
  DFF \state_reg[7]  ( .D(state[7]), .CLK(clk), .RST(rst), .I(msg[7]), .Q(
        state[7]) );
  DFF \state_reg[6]  ( .D(state[6]), .CLK(clk), .RST(rst), .I(msg[6]), .Q(
        state[6]) );
  DFF \state_reg[5]  ( .D(state[5]), .CLK(clk), .RST(rst), .I(msg[5]), .Q(
        state[5]) );
  DFF \state_reg[4]  ( .D(state[4]), .CLK(clk), .RST(rst), .I(msg[4]), .Q(
        state[4]) );
  DFF \state_reg[3]  ( .D(state[3]), .CLK(clk), .RST(rst), .I(msg[3]), .Q(
        state[3]) );
  DFF \state_reg[2]  ( .D(state[2]), .CLK(clk), .RST(rst), .I(msg[2]), .Q(
        state[2]) );
  DFF \state_reg[1]  ( .D(state[1]), .CLK(clk), .RST(rst), .I(msg[1]), .Q(
        state[1]) );
  DFF \state_reg[0]  ( .D(state[0]), .CLK(clk), .RST(rst), .I(msg[0]), .Q(
        state[0]) );
  XOR U4 ( .A(n1498), .B(n691), .Z(n2424) );
  XOR U5 ( .A(n1538), .B(n1469), .Z(n1589) );
  XOR U6 ( .A(n1359), .B(n1316), .Z(n1410) );
  XOR U7 ( .A(n1039), .B(n997), .Z(n1090) );
  XOR U8 ( .A(n887), .B(n842), .Z(n938) );
  XOR U9 ( .A(n732), .B(n673), .Z(n783) );
  XOR U10 ( .A(n591), .B(n580), .Z(n587) );
  XOR U11 ( .A(n240), .B(n198), .Z(n291) );
  XOR U12 ( .A(n88), .B(n42), .Z(n139) );
  XOR U13 ( .A(n1726), .B(n1683), .Z(n1777) );
  XOR U14 ( .A(n644), .B(n642), .Z(n615) );
  XOR U15 ( .A(n2267), .B(n2254), .Z(n2266) );
  XOR U16 ( .A(n2402), .B(n2392), .Z(n2399) );
  XOR U17 ( .A(n1477), .B(n1135), .Z(n1493) );
  XOR U18 ( .A(n1567), .B(n1557), .Z(n1564) );
  XOR U19 ( .A(n1517), .B(n1507), .Z(n1533) );
  XOR U20 ( .A(n1388), .B(n1378), .Z(n1385) );
  XOR U21 ( .A(n1338), .B(n1328), .Z(n1354) );
  XOR U22 ( .A(n1233), .B(n1223), .Z(n1230) );
  XOR U23 ( .A(n1068), .B(n1058), .Z(n1065) );
  XOR U24 ( .A(n1018), .B(n1009), .Z(n1034) );
  XOR U25 ( .A(n916), .B(n906), .Z(n913) );
  XOR U26 ( .A(n866), .B(n854), .Z(n882) );
  XOR U27 ( .A(n761), .B(n751), .Z(n758) );
  XOR U28 ( .A(n711), .B(n701), .Z(n727) );
  XNOR U29 ( .A(n614), .B(n622), .Z(n621) );
  XOR U30 ( .A(n269), .B(n259), .Z(n266) );
  XOR U31 ( .A(n219), .B(n210), .Z(n235) );
  XOR U32 ( .A(n117), .B(n107), .Z(n114) );
  XOR U33 ( .A(n67), .B(n54), .Z(n83) );
  XOR U34 ( .A(n2314), .B(n2304), .Z(n2311) );
  XOR U35 ( .A(n2172), .B(n2162), .Z(n2169) );
  XOR U36 ( .A(n1936), .B(n1926), .Z(n1933) );
  XOR U37 ( .A(n1755), .B(n1745), .Z(n1752) );
  XOR U38 ( .A(n1705), .B(n1695), .Z(n1721) );
  XOR U39 ( .A(n2309), .B(n2298), .Z(n2300) );
  XOR U40 ( .A(n2379), .B(n1498), .Z(n2387) );
  XOR U41 ( .A(n2027), .B(n2016), .Z(n2023) );
  XOR U42 ( .A(n2011), .B(n2005), .Z(n1660) );
  XOR U43 ( .A(n1544), .B(n1538), .Z(n1552) );
  XOR U44 ( .A(n1365), .B(n1359), .Z(n1373) );
  XOR U45 ( .A(n1183), .B(n1173), .Z(n1199) );
  XOR U46 ( .A(n1045), .B(n1039), .Z(n1053) );
  XOR U47 ( .A(n893), .B(n887), .Z(n901) );
  XOR U48 ( .A(n738), .B(n732), .Z(n746) );
  XOR U49 ( .A(n565), .B(n519), .Z(n548) );
  XOR U50 ( .A(n246), .B(n240), .Z(n254) );
  XOR U51 ( .A(n94), .B(n88), .Z(n102) );
  XOR U52 ( .A(n2122), .B(n2112), .Z(n2138) );
  XOR U53 ( .A(n1886), .B(n1876), .Z(n1902) );
  XOR U54 ( .A(n1732), .B(n1726), .Z(n1740) );
  XOR U55 ( .A(n2445), .B(n2448), .Z(n2452) );
  XOR U56 ( .A(n2407), .B(n2401), .Z(n2406) );
  ANDN U57 ( .B(n1840), .A(n1841), .Z(n1837) );
  XOR U58 ( .A(n1610), .B(n1613), .Z(n1617) );
  XOR U59 ( .A(n1572), .B(n1566), .Z(n1571) );
  XOR U60 ( .A(n1431), .B(n1434), .Z(n1438) );
  XOR U61 ( .A(n1393), .B(n1387), .Z(n1392) );
  XOR U62 ( .A(n1238), .B(n1232), .Z(n1237) );
  XOR U63 ( .A(n1111), .B(n1114), .Z(n1118) );
  XOR U64 ( .A(n1073), .B(n1067), .Z(n1072) );
  XOR U65 ( .A(n959), .B(n962), .Z(n966) );
  XOR U66 ( .A(n921), .B(n915), .Z(n920) );
  XOR U67 ( .A(n804), .B(n807), .Z(n811) );
  XOR U68 ( .A(n766), .B(n760), .Z(n765) );
  XNOR U69 ( .A(n644), .B(n647), .Z(n570) );
  XNOR U70 ( .A(n430), .B(n421), .Z(n352) );
  XOR U71 ( .A(n312), .B(n315), .Z(n319) );
  XOR U72 ( .A(n274), .B(n268), .Z(n273) );
  XOR U73 ( .A(n160), .B(n163), .Z(n167) );
  XOR U74 ( .A(n122), .B(n116), .Z(n121) );
  XNOR U75 ( .A(n2248), .B(n2366), .Z(n2258) );
  XNOR U76 ( .A(n2315), .B(n2302), .Z(n2247) );
  XOR U77 ( .A(n2177), .B(n2171), .Z(n2176) );
  XOR U78 ( .A(n1941), .B(n1935), .Z(n1940) );
  XOR U79 ( .A(n1798), .B(n1801), .Z(n1805) );
  XOR U80 ( .A(n1760), .B(n1754), .Z(n1759) );
  XOR U81 ( .A(n1493), .B(n1482), .Z(n1491) );
  XOR U82 ( .A(n1533), .B(n1522), .Z(n1531) );
  XOR U83 ( .A(n1354), .B(n1343), .Z(n1352) );
  XOR U84 ( .A(n1199), .B(n1188), .Z(n1197) );
  XOR U85 ( .A(n1034), .B(n1023), .Z(n1032) );
  XOR U86 ( .A(n882), .B(n871), .Z(n880) );
  XOR U87 ( .A(n727), .B(n716), .Z(n725) );
  XOR U88 ( .A(n436), .B(n423), .Z(n431) );
  XOR U89 ( .A(n235), .B(n224), .Z(n233) );
  XOR U90 ( .A(n83), .B(n72), .Z(n81) );
  XOR U91 ( .A(n2138), .B(n2127), .Z(n2136) );
  XOR U92 ( .A(n1902), .B(n1891), .Z(n1900) );
  XOR U93 ( .A(n1721), .B(n1710), .Z(n1719) );
  XNOR U94 ( .A(n1210), .B(n1204), .Z(n1218) );
  XOR U95 ( .A(n544), .B(n528), .Z(n559) );
  XNOR U96 ( .A(n566), .B(n615), .Z(n574) );
  XNOR U97 ( .A(n483), .B(n481), .Z(n468) );
  XNOR U98 ( .A(n2149), .B(n2143), .Z(n2157) );
  XNOR U99 ( .A(n1913), .B(n1907), .Z(n1921) );
  XNOR U100 ( .A(n2403), .B(n2390), .Z(n1136) );
  XNOR U101 ( .A(n2444), .B(n2442), .Z(n1498) );
  XOR U102 ( .A(n2080), .B(n2081), .Z(n2082) );
  XNOR U103 ( .A(n2028), .B(n2018), .Z(n1641) );
  XNOR U104 ( .A(n1609), .B(n1607), .Z(n1538) );
  XNOR U105 ( .A(n1568), .B(n1555), .Z(n1508) );
  XNOR U106 ( .A(n1430), .B(n1428), .Z(n1359) );
  XNOR U107 ( .A(n1389), .B(n1376), .Z(n1329) );
  XNOR U108 ( .A(n1234), .B(n1221), .Z(n1174) );
  XNOR U109 ( .A(n1069), .B(n1056), .Z(n1010) );
  XNOR U110 ( .A(n1110), .B(n1108), .Z(n1039) );
  XNOR U111 ( .A(n958), .B(n956), .Z(n887) );
  XNOR U112 ( .A(n917), .B(n904), .Z(n855) );
  XNOR U113 ( .A(n803), .B(n801), .Z(n732) );
  XNOR U114 ( .A(n762), .B(n749), .Z(n702) );
  XNOR U115 ( .A(n592), .B(n582), .Z(n513) );
  XNOR U116 ( .A(n270), .B(n257), .Z(n211) );
  XNOR U117 ( .A(n311), .B(n309), .Z(n240) );
  XNOR U118 ( .A(n159), .B(n157), .Z(n88) );
  XNOR U119 ( .A(n118), .B(n105), .Z(n55) );
  XOR U120 ( .A(n2319), .B(n2313), .Z(n2318) );
  XNOR U121 ( .A(n2357), .B(n2355), .Z(n2290) );
  XNOR U122 ( .A(n2173), .B(n2160), .Z(n2113) );
  XNOR U123 ( .A(n1937), .B(n1924), .Z(n1877) );
  XNOR U124 ( .A(n1797), .B(n1795), .Z(n1726) );
  XNOR U125 ( .A(n1756), .B(n1743), .Z(n1696) );
  XNOR U126 ( .A(n503), .B(n1129), .Z(n329) );
  XOR U127 ( .A(n62), .B(n1632), .Z(n3) );
  XNOR U128 ( .A(n1454), .B(n1501), .Z(n1448) );
  XNOR U129 ( .A(n1299), .B(n1322), .Z(n1293) );
  XNOR U130 ( .A(n1146), .B(n1167), .Z(n1140) );
  XNOR U131 ( .A(n982), .B(n1003), .Z(n976) );
  XNOR U132 ( .A(n827), .B(n848), .Z(n821) );
  XNOR U133 ( .A(n658), .B(n695), .Z(n652) );
  XOR U134 ( .A(n375), .B(n363), .Z(n334) );
  XNOR U135 ( .A(n183), .B(n204), .Z(n177) );
  XNOR U136 ( .A(n27), .B(n48), .Z(n21) );
  XNOR U137 ( .A(n2237), .B(n2244), .Z(n10) );
  XNOR U138 ( .A(n2002), .B(n2106), .Z(n1996) );
  XNOR U139 ( .A(n1849), .B(n1870), .Z(n1843) );
  XNOR U140 ( .A(n1668), .B(n1689), .Z(n1662) );
  XOR U141 ( .A(n1), .B(n2), .Z(out[9]) );
  XNOR U142 ( .A(n3), .B(n4), .Z(n2) );
  XOR U143 ( .A(key[9]), .B(n5), .Z(n1) );
  XOR U144 ( .A(n6), .B(n7), .Z(out[99]) );
  XNOR U145 ( .A(n8), .B(n9), .Z(n7) );
  XOR U146 ( .A(n10), .B(n11), .Z(n6) );
  XNOR U147 ( .A(key[99]), .B(n12), .Z(n11) );
  XNOR U148 ( .A(key[98]), .B(n13), .Z(out[98]) );
  XOR U149 ( .A(n14), .B(n15), .Z(out[97]) );
  XOR U150 ( .A(n8), .B(n16), .Z(n15) );
  XNOR U151 ( .A(key[97]), .B(n12), .Z(n14) );
  XOR U152 ( .A(n17), .B(n18), .Z(out[96]) );
  XNOR U153 ( .A(key[96]), .B(n19), .Z(n18) );
  XOR U154 ( .A(n20), .B(n21), .Z(out[95]) );
  XOR U155 ( .A(n22), .B(n23), .Z(n20) );
  XOR U156 ( .A(key[95]), .B(n24), .Z(n23) );
  XNOR U157 ( .A(n25), .B(n26), .Z(out[94]) );
  XNOR U158 ( .A(key[94]), .B(n27), .Z(n26) );
  XOR U159 ( .A(n28), .B(n29), .Z(out[93]) );
  XNOR U160 ( .A(n30), .B(n31), .Z(n29) );
  XOR U161 ( .A(n22), .B(n32), .Z(n31) );
  XOR U162 ( .A(n33), .B(n34), .Z(n22) );
  XNOR U163 ( .A(n35), .B(n36), .Z(n34) );
  NANDN U164 ( .A(n37), .B(n38), .Z(n36) );
  XOR U165 ( .A(n39), .B(n40), .Z(n28) );
  XOR U166 ( .A(key[93]), .B(n41), .Z(n40) );
  ANDN U167 ( .B(n42), .A(n43), .Z(n39) );
  XNOR U168 ( .A(n44), .B(n45), .Z(out[92]) );
  XOR U169 ( .A(key[92]), .B(n30), .Z(n45) );
  XOR U170 ( .A(n46), .B(n47), .Z(out[91]) );
  XOR U171 ( .A(n48), .B(n25), .Z(n47) );
  XNOR U172 ( .A(n49), .B(n50), .Z(n25) );
  XNOR U173 ( .A(n51), .B(n41), .Z(n50) );
  NOR U174 ( .A(n52), .B(n53), .Z(n41) );
  ANDN U175 ( .B(n54), .A(n55), .Z(n51) );
  XNOR U176 ( .A(n56), .B(n57), .Z(n46) );
  XNOR U177 ( .A(key[91]), .B(n58), .Z(n57) );
  XOR U178 ( .A(key[90]), .B(n44), .Z(out[90]) );
  XOR U179 ( .A(n24), .B(n59), .Z(n44) );
  XNOR U180 ( .A(n60), .B(n61), .Z(out[8]) );
  XNOR U181 ( .A(key[8]), .B(n62), .Z(n61) );
  XOR U182 ( .A(n63), .B(n21), .Z(out[89]) );
  XOR U183 ( .A(n49), .B(n64), .Z(n48) );
  XNOR U184 ( .A(n65), .B(n66), .Z(n64) );
  NANDN U185 ( .A(n37), .B(n67), .Z(n66) );
  XNOR U186 ( .A(n32), .B(n68), .Z(n49) );
  XNOR U187 ( .A(n69), .B(n70), .Z(n68) );
  NANDN U188 ( .A(n71), .B(n72), .Z(n70) );
  XOR U189 ( .A(n59), .B(n56), .Z(n27) );
  XNOR U190 ( .A(n32), .B(n73), .Z(n56) );
  XNOR U191 ( .A(n65), .B(n74), .Z(n73) );
  NAND U192 ( .A(n75), .B(n76), .Z(n74) );
  OR U193 ( .A(n77), .B(n78), .Z(n65) );
  XOR U194 ( .A(n79), .B(n69), .Z(n32) );
  NANDN U195 ( .A(n80), .B(n81), .Z(n69) );
  AND U196 ( .A(n82), .B(n83), .Z(n79) );
  XOR U197 ( .A(key[89]), .B(n24), .Z(n63) );
  IV U198 ( .A(n58), .Z(n24) );
  XNOR U199 ( .A(n84), .B(n85), .Z(n58) );
  XNOR U200 ( .A(n86), .B(n87), .Z(n85) );
  NANDN U201 ( .A(n43), .B(n88), .Z(n87) );
  XNOR U202 ( .A(n30), .B(n89), .Z(out[88]) );
  XOR U203 ( .A(key[88]), .B(n59), .Z(n89) );
  XNOR U204 ( .A(n84), .B(n90), .Z(n59) );
  XOR U205 ( .A(n91), .B(n35), .Z(n90) );
  OR U206 ( .A(n92), .B(n77), .Z(n35) );
  XNOR U207 ( .A(n37), .B(n93), .Z(n77) );
  AND U208 ( .A(n94), .B(n75), .Z(n91) );
  XNOR U209 ( .A(n33), .B(n95), .Z(n30) );
  XOR U210 ( .A(n96), .B(n86), .Z(n95) );
  OR U211 ( .A(n97), .B(n52), .Z(n86) );
  XNOR U212 ( .A(n55), .B(n43), .Z(n52) );
  NOR U213 ( .A(n98), .B(n55), .Z(n96) );
  XNOR U214 ( .A(n84), .B(n99), .Z(n33) );
  XNOR U215 ( .A(n100), .B(n101), .Z(n99) );
  NANDN U216 ( .A(n71), .B(n102), .Z(n101) );
  XOR U217 ( .A(n103), .B(n100), .Z(n84) );
  OR U218 ( .A(n80), .B(n104), .Z(n100) );
  XOR U219 ( .A(n82), .B(n71), .Z(n80) );
  XNOR U220 ( .A(n93), .B(n43), .Z(n71) );
  XOR U221 ( .A(n105), .B(n106), .Z(n43) );
  NANDN U222 ( .A(n107), .B(n108), .Z(n106) );
  IV U223 ( .A(n75), .Z(n93) );
  XOR U224 ( .A(n109), .B(n110), .Z(n75) );
  NANDN U225 ( .A(n107), .B(n111), .Z(n110) );
  ANDN U226 ( .B(n82), .A(n112), .Z(n103) );
  XOR U227 ( .A(n55), .B(n37), .Z(n82) );
  XOR U228 ( .A(n113), .B(n109), .Z(n37) );
  NANDN U229 ( .A(n114), .B(n115), .Z(n109) );
  AND U230 ( .A(n116), .B(n117), .Z(n113) );
  ANDN U231 ( .B(n119), .A(n114), .Z(n105) );
  XOR U232 ( .A(n120), .B(n121), .Z(n107) );
  XNOR U233 ( .A(n123), .B(n124), .Z(n120) );
  XNOR U234 ( .A(n125), .B(n126), .Z(n124) );
  AND U235 ( .A(n127), .B(n116), .Z(n125) );
  AND U236 ( .A(n127), .B(n117), .Z(n118) );
  XOR U237 ( .A(n123), .B(n128), .Z(n117) );
  XOR U238 ( .A(n129), .B(n126), .Z(n128) );
  NAND U239 ( .A(n115), .B(n119), .Z(n126) );
  XOR U240 ( .A(n108), .B(n127), .Z(n119) );
  XOR U241 ( .A(n111), .B(n116), .Z(n115) );
  XNOR U242 ( .A(n130), .B(n131), .Z(n116) );
  XOR U243 ( .A(n132), .B(n133), .Z(n131) );
  XNOR U244 ( .A(n134), .B(n135), .Z(n130) );
  ANDN U245 ( .B(n54), .A(n98), .Z(n134) );
  AND U246 ( .A(n108), .B(n111), .Z(n129) );
  XNOR U247 ( .A(n108), .B(n111), .Z(n123) );
  XNOR U248 ( .A(n136), .B(n137), .Z(n111) );
  XOR U249 ( .A(n138), .B(n139), .Z(n137) );
  XOR U250 ( .A(n132), .B(n140), .Z(n136) );
  XNOR U251 ( .A(n141), .B(n135), .Z(n140) );
  OR U252 ( .A(n53), .B(n97), .Z(n135) );
  XOR U253 ( .A(n98), .B(n88), .Z(n97) );
  XOR U254 ( .A(n142), .B(n42), .Z(n53) );
  AND U255 ( .A(n42), .B(n88), .Z(n141) );
  XNOR U256 ( .A(n143), .B(n144), .Z(n108) );
  XOR U257 ( .A(n145), .B(n146), .Z(n144) );
  XNOR U258 ( .A(n67), .B(n132), .Z(n146) );
  XNOR U259 ( .A(n98), .B(n54), .Z(n132) );
  XOR U260 ( .A(n38), .B(n147), .Z(n143) );
  XNOR U261 ( .A(n148), .B(n149), .Z(n147) );
  AND U262 ( .A(n76), .B(n94), .Z(n148) );
  IV U263 ( .A(n122), .Z(n127) );
  XOR U264 ( .A(n150), .B(n151), .Z(n122) );
  XNOR U265 ( .A(n133), .B(n152), .Z(n151) );
  XNOR U266 ( .A(n76), .B(n139), .Z(n152) );
  XOR U267 ( .A(n145), .B(n153), .Z(n133) );
  XNOR U268 ( .A(n154), .B(n155), .Z(n153) );
  NAND U269 ( .A(n72), .B(n102), .Z(n155) );
  IV U270 ( .A(n138), .Z(n145) );
  XOR U271 ( .A(n156), .B(n154), .Z(n138) );
  NANDN U272 ( .A(n104), .B(n81), .Z(n154) );
  XOR U273 ( .A(n76), .B(n42), .Z(n72) );
  XOR U274 ( .A(n157), .B(n158), .Z(n42) );
  XOR U275 ( .A(n159), .B(n160), .Z(n158) );
  XOR U276 ( .A(n112), .B(n102), .Z(n104) );
  ANDN U277 ( .B(n83), .A(n112), .Z(n156) );
  XNOR U278 ( .A(n161), .B(n98), .Z(n112) );
  XNOR U279 ( .A(n162), .B(n163), .Z(n98) );
  XOR U280 ( .A(n164), .B(n159), .Z(n162) );
  XOR U281 ( .A(n94), .B(n165), .Z(n150) );
  XNOR U282 ( .A(n166), .B(n149), .Z(n165) );
  OR U283 ( .A(n78), .B(n92), .Z(n149) );
  XNOR U284 ( .A(n38), .B(n94), .Z(n92) );
  XNOR U285 ( .A(n67), .B(n76), .Z(n78) );
  XOR U286 ( .A(n142), .B(n167), .Z(n76) );
  XOR U287 ( .A(state[90]), .B(key[90]), .Z(n163) );
  IV U288 ( .A(n54), .Z(n142) );
  XOR U289 ( .A(n157), .B(n168), .Z(n54) );
  XNOR U290 ( .A(n159), .B(n169), .Z(n168) );
  AND U291 ( .A(n38), .B(n67), .Z(n166) );
  XOR U292 ( .A(n157), .B(n170), .Z(n67) );
  XNOR U293 ( .A(n159), .B(n171), .Z(n170) );
  XOR U294 ( .A(n161), .B(n172), .Z(n159) );
  XNOR U295 ( .A(state[94]), .B(key[94]), .Z(n172) );
  XNOR U296 ( .A(state[93]), .B(key[93]), .Z(n157) );
  XNOR U297 ( .A(n173), .B(n174), .Z(n94) );
  XNOR U298 ( .A(n171), .B(n169), .Z(n174) );
  XOR U299 ( .A(state[95]), .B(key[95]), .Z(n169) );
  XOR U300 ( .A(state[92]), .B(key[92]), .Z(n171) );
  XOR U301 ( .A(n38), .B(n164), .Z(n173) );
  XOR U302 ( .A(n160), .B(n175), .Z(n164) );
  XNOR U303 ( .A(state[91]), .B(key[91]), .Z(n175) );
  XNOR U304 ( .A(state[89]), .B(key[89]), .Z(n160) );
  IV U305 ( .A(n161), .Z(n38) );
  XNOR U306 ( .A(state[88]), .B(key[88]), .Z(n161) );
  XOR U307 ( .A(n176), .B(n177), .Z(out[87]) );
  XOR U308 ( .A(n178), .B(n179), .Z(n176) );
  XNOR U309 ( .A(key[87]), .B(n180), .Z(n179) );
  XNOR U310 ( .A(n181), .B(n182), .Z(out[86]) );
  XNOR U311 ( .A(key[86]), .B(n183), .Z(n182) );
  XOR U312 ( .A(n184), .B(n185), .Z(out[85]) );
  XNOR U313 ( .A(n186), .B(n187), .Z(n185) );
  XOR U314 ( .A(n178), .B(n188), .Z(n187) );
  XOR U315 ( .A(n189), .B(n190), .Z(n178) );
  XNOR U316 ( .A(n191), .B(n192), .Z(n190) );
  NANDN U317 ( .A(n193), .B(n194), .Z(n192) );
  XOR U318 ( .A(n195), .B(n196), .Z(n184) );
  XOR U319 ( .A(key[85]), .B(n197), .Z(n196) );
  ANDN U320 ( .B(n198), .A(n199), .Z(n195) );
  XNOR U321 ( .A(n200), .B(n201), .Z(out[84]) );
  XOR U322 ( .A(key[84]), .B(n186), .Z(n201) );
  XOR U323 ( .A(n202), .B(n203), .Z(out[83]) );
  XOR U324 ( .A(n204), .B(n181), .Z(n203) );
  XNOR U325 ( .A(n205), .B(n206), .Z(n181) );
  XNOR U326 ( .A(n207), .B(n197), .Z(n206) );
  NOR U327 ( .A(n208), .B(n209), .Z(n197) );
  ANDN U328 ( .B(n210), .A(n211), .Z(n207) );
  XNOR U329 ( .A(n212), .B(n213), .Z(n202) );
  XNOR U330 ( .A(key[83]), .B(n180), .Z(n213) );
  XOR U331 ( .A(key[82]), .B(n200), .Z(out[82]) );
  XNOR U332 ( .A(n180), .B(n214), .Z(n200) );
  XOR U333 ( .A(n215), .B(n177), .Z(out[81]) );
  XOR U334 ( .A(n205), .B(n216), .Z(n204) );
  XNOR U335 ( .A(n217), .B(n218), .Z(n216) );
  NANDN U336 ( .A(n193), .B(n219), .Z(n218) );
  XNOR U337 ( .A(n188), .B(n220), .Z(n205) );
  XNOR U338 ( .A(n221), .B(n222), .Z(n220) );
  NANDN U339 ( .A(n223), .B(n224), .Z(n222) );
  XOR U340 ( .A(n214), .B(n212), .Z(n183) );
  XNOR U341 ( .A(n188), .B(n225), .Z(n212) );
  XNOR U342 ( .A(n217), .B(n226), .Z(n225) );
  NAND U343 ( .A(n227), .B(n228), .Z(n226) );
  OR U344 ( .A(n229), .B(n230), .Z(n217) );
  XOR U345 ( .A(n231), .B(n221), .Z(n188) );
  NANDN U346 ( .A(n232), .B(n233), .Z(n221) );
  AND U347 ( .A(n234), .B(n235), .Z(n231) );
  XNOR U348 ( .A(key[81]), .B(n180), .Z(n215) );
  XNOR U349 ( .A(n236), .B(n237), .Z(n180) );
  XNOR U350 ( .A(n238), .B(n239), .Z(n237) );
  NANDN U351 ( .A(n199), .B(n240), .Z(n239) );
  XNOR U352 ( .A(n186), .B(n241), .Z(out[80]) );
  XOR U353 ( .A(key[80]), .B(n214), .Z(n241) );
  XNOR U354 ( .A(n236), .B(n242), .Z(n214) );
  XOR U355 ( .A(n243), .B(n191), .Z(n242) );
  OR U356 ( .A(n244), .B(n229), .Z(n191) );
  XNOR U357 ( .A(n193), .B(n245), .Z(n229) );
  AND U358 ( .A(n246), .B(n227), .Z(n243) );
  XNOR U359 ( .A(n189), .B(n247), .Z(n186) );
  XOR U360 ( .A(n248), .B(n238), .Z(n247) );
  OR U361 ( .A(n249), .B(n208), .Z(n238) );
  XNOR U362 ( .A(n211), .B(n199), .Z(n208) );
  NOR U363 ( .A(n250), .B(n211), .Z(n248) );
  XNOR U364 ( .A(n236), .B(n251), .Z(n189) );
  XNOR U365 ( .A(n252), .B(n253), .Z(n251) );
  NANDN U366 ( .A(n223), .B(n254), .Z(n253) );
  XOR U367 ( .A(n255), .B(n252), .Z(n236) );
  OR U368 ( .A(n232), .B(n256), .Z(n252) );
  XOR U369 ( .A(n234), .B(n223), .Z(n232) );
  XNOR U370 ( .A(n245), .B(n199), .Z(n223) );
  XOR U371 ( .A(n257), .B(n258), .Z(n199) );
  NANDN U372 ( .A(n259), .B(n260), .Z(n258) );
  IV U373 ( .A(n227), .Z(n245) );
  XOR U374 ( .A(n261), .B(n262), .Z(n227) );
  NANDN U375 ( .A(n259), .B(n263), .Z(n262) );
  ANDN U376 ( .B(n234), .A(n264), .Z(n255) );
  XOR U377 ( .A(n211), .B(n193), .Z(n234) );
  XOR U378 ( .A(n265), .B(n261), .Z(n193) );
  NANDN U379 ( .A(n266), .B(n267), .Z(n261) );
  AND U380 ( .A(n268), .B(n269), .Z(n265) );
  ANDN U381 ( .B(n271), .A(n266), .Z(n257) );
  XOR U382 ( .A(n272), .B(n273), .Z(n259) );
  XNOR U383 ( .A(n275), .B(n276), .Z(n272) );
  XNOR U384 ( .A(n277), .B(n278), .Z(n276) );
  AND U385 ( .A(n279), .B(n268), .Z(n277) );
  AND U386 ( .A(n279), .B(n269), .Z(n270) );
  XOR U387 ( .A(n275), .B(n280), .Z(n269) );
  XOR U388 ( .A(n281), .B(n278), .Z(n280) );
  NAND U389 ( .A(n267), .B(n271), .Z(n278) );
  XOR U390 ( .A(n260), .B(n279), .Z(n271) );
  XOR U391 ( .A(n263), .B(n268), .Z(n267) );
  XNOR U392 ( .A(n282), .B(n283), .Z(n268) );
  XOR U393 ( .A(n284), .B(n285), .Z(n283) );
  XNOR U394 ( .A(n286), .B(n287), .Z(n282) );
  ANDN U395 ( .B(n210), .A(n250), .Z(n286) );
  AND U396 ( .A(n260), .B(n263), .Z(n281) );
  XNOR U397 ( .A(n260), .B(n263), .Z(n275) );
  XNOR U398 ( .A(n288), .B(n289), .Z(n263) );
  XOR U399 ( .A(n290), .B(n291), .Z(n289) );
  XOR U400 ( .A(n284), .B(n292), .Z(n288) );
  XNOR U401 ( .A(n293), .B(n287), .Z(n292) );
  OR U402 ( .A(n209), .B(n249), .Z(n287) );
  XOR U403 ( .A(n250), .B(n240), .Z(n249) );
  XOR U404 ( .A(n294), .B(n198), .Z(n209) );
  AND U405 ( .A(n198), .B(n240), .Z(n293) );
  XNOR U406 ( .A(n295), .B(n296), .Z(n260) );
  XOR U407 ( .A(n297), .B(n298), .Z(n296) );
  XNOR U408 ( .A(n219), .B(n284), .Z(n298) );
  XNOR U409 ( .A(n250), .B(n210), .Z(n284) );
  XOR U410 ( .A(n194), .B(n299), .Z(n295) );
  XNOR U411 ( .A(n300), .B(n301), .Z(n299) );
  AND U412 ( .A(n228), .B(n246), .Z(n300) );
  IV U413 ( .A(n274), .Z(n279) );
  XOR U414 ( .A(n302), .B(n303), .Z(n274) );
  XNOR U415 ( .A(n285), .B(n304), .Z(n303) );
  XNOR U416 ( .A(n228), .B(n291), .Z(n304) );
  XOR U417 ( .A(n297), .B(n305), .Z(n285) );
  XNOR U418 ( .A(n306), .B(n307), .Z(n305) );
  NAND U419 ( .A(n224), .B(n254), .Z(n307) );
  IV U420 ( .A(n290), .Z(n297) );
  XOR U421 ( .A(n308), .B(n306), .Z(n290) );
  NANDN U422 ( .A(n256), .B(n233), .Z(n306) );
  XOR U423 ( .A(n228), .B(n198), .Z(n224) );
  XOR U424 ( .A(n309), .B(n310), .Z(n198) );
  XOR U425 ( .A(n311), .B(n312), .Z(n310) );
  XOR U426 ( .A(n264), .B(n254), .Z(n256) );
  ANDN U427 ( .B(n235), .A(n264), .Z(n308) );
  XNOR U428 ( .A(n313), .B(n250), .Z(n264) );
  XNOR U429 ( .A(n314), .B(n315), .Z(n250) );
  XOR U430 ( .A(n316), .B(n311), .Z(n314) );
  XOR U431 ( .A(n246), .B(n317), .Z(n302) );
  XNOR U432 ( .A(n318), .B(n301), .Z(n317) );
  OR U433 ( .A(n230), .B(n244), .Z(n301) );
  XNOR U434 ( .A(n194), .B(n246), .Z(n244) );
  XNOR U435 ( .A(n219), .B(n228), .Z(n230) );
  XOR U436 ( .A(n294), .B(n319), .Z(n228) );
  XOR U437 ( .A(state[50]), .B(key[50]), .Z(n315) );
  IV U438 ( .A(n210), .Z(n294) );
  XOR U439 ( .A(n309), .B(n320), .Z(n210) );
  XNOR U440 ( .A(n311), .B(n321), .Z(n320) );
  AND U441 ( .A(n194), .B(n219), .Z(n318) );
  XOR U442 ( .A(n309), .B(n322), .Z(n219) );
  XNOR U443 ( .A(n311), .B(n323), .Z(n322) );
  XOR U444 ( .A(n313), .B(n324), .Z(n311) );
  XNOR U445 ( .A(state[54]), .B(key[54]), .Z(n324) );
  XNOR U446 ( .A(state[53]), .B(key[53]), .Z(n309) );
  XNOR U447 ( .A(n325), .B(n326), .Z(n246) );
  XNOR U448 ( .A(n323), .B(n321), .Z(n326) );
  XOR U449 ( .A(state[55]), .B(key[55]), .Z(n321) );
  XOR U450 ( .A(state[52]), .B(key[52]), .Z(n323) );
  XOR U451 ( .A(n194), .B(n316), .Z(n325) );
  XOR U452 ( .A(n312), .B(n327), .Z(n316) );
  XNOR U453 ( .A(state[51]), .B(key[51]), .Z(n327) );
  XNOR U454 ( .A(state[49]), .B(key[49]), .Z(n312) );
  IV U455 ( .A(n313), .Z(n194) );
  XNOR U456 ( .A(state[48]), .B(key[48]), .Z(n313) );
  XOR U457 ( .A(n328), .B(n329), .Z(out[7]) );
  XOR U458 ( .A(n330), .B(n331), .Z(n328) );
  XNOR U459 ( .A(key[7]), .B(n332), .Z(n331) );
  XOR U460 ( .A(n333), .B(n334), .Z(out[79]) );
  XOR U461 ( .A(n335), .B(n336), .Z(n333) );
  XNOR U462 ( .A(key[79]), .B(n337), .Z(n336) );
  XOR U463 ( .A(n338), .B(n339), .Z(out[78]) );
  XOR U464 ( .A(n340), .B(n341), .Z(n339) );
  XNOR U465 ( .A(key[78]), .B(n342), .Z(n338) );
  XOR U466 ( .A(n343), .B(n344), .Z(out[77]) );
  XNOR U467 ( .A(n345), .B(n346), .Z(n344) );
  XOR U468 ( .A(n335), .B(n347), .Z(n346) );
  XOR U469 ( .A(n348), .B(n349), .Z(n335) );
  XNOR U470 ( .A(n350), .B(n351), .Z(n349) );
  NANDN U471 ( .A(n352), .B(n353), .Z(n351) );
  XOR U472 ( .A(n354), .B(n355), .Z(n343) );
  XOR U473 ( .A(key[77]), .B(n356), .Z(n355) );
  AND U474 ( .A(n357), .B(n358), .Z(n354) );
  XNOR U475 ( .A(n359), .B(n360), .Z(out[76]) );
  XOR U476 ( .A(key[76]), .B(n345), .Z(n360) );
  XOR U477 ( .A(n361), .B(n362), .Z(out[75]) );
  XOR U478 ( .A(n363), .B(n341), .Z(n362) );
  XNOR U479 ( .A(n364), .B(n365), .Z(n341) );
  XNOR U480 ( .A(n366), .B(n356), .Z(n365) );
  NOR U481 ( .A(n367), .B(n368), .Z(n356) );
  ANDN U482 ( .B(n369), .A(n370), .Z(n366) );
  XNOR U483 ( .A(n371), .B(n372), .Z(n361) );
  XNOR U484 ( .A(key[75]), .B(n337), .Z(n372) );
  XOR U485 ( .A(key[74]), .B(n359), .Z(out[74]) );
  XOR U486 ( .A(n373), .B(n342), .Z(n359) );
  XOR U487 ( .A(n374), .B(n334), .Z(out[73]) );
  XOR U488 ( .A(n364), .B(n376), .Z(n363) );
  XOR U489 ( .A(n377), .B(n378), .Z(n376) );
  ANDN U490 ( .B(n379), .A(n352), .Z(n377) );
  XNOR U491 ( .A(n347), .B(n380), .Z(n364) );
  XNOR U492 ( .A(n381), .B(n382), .Z(n380) );
  NAND U493 ( .A(n383), .B(n384), .Z(n382) );
  XNOR U494 ( .A(n342), .B(n371), .Z(n375) );
  IV U495 ( .A(n340), .Z(n371) );
  XOR U496 ( .A(n347), .B(n385), .Z(n340) );
  XNOR U497 ( .A(n378), .B(n386), .Z(n385) );
  NANDN U498 ( .A(n387), .B(n388), .Z(n386) );
  OR U499 ( .A(n389), .B(n390), .Z(n378) );
  XOR U500 ( .A(n391), .B(n381), .Z(n347) );
  NANDN U501 ( .A(n392), .B(n393), .Z(n381) );
  AND U502 ( .A(n394), .B(n395), .Z(n391) );
  XOR U503 ( .A(key[73]), .B(n373), .Z(n374) );
  IV U504 ( .A(n337), .Z(n373) );
  XNOR U505 ( .A(n396), .B(n397), .Z(n337) );
  XNOR U506 ( .A(n398), .B(n399), .Z(n397) );
  NAND U507 ( .A(n400), .B(n358), .Z(n399) );
  XNOR U508 ( .A(n345), .B(n401), .Z(out[72]) );
  XOR U509 ( .A(key[72]), .B(n342), .Z(n401) );
  XNOR U510 ( .A(n396), .B(n402), .Z(n342) );
  XOR U511 ( .A(n403), .B(n350), .Z(n402) );
  OR U512 ( .A(n404), .B(n389), .Z(n350) );
  XNOR U513 ( .A(n352), .B(n387), .Z(n389) );
  ANDN U514 ( .B(n405), .A(n387), .Z(n403) );
  XNOR U515 ( .A(n348), .B(n406), .Z(n345) );
  XNOR U516 ( .A(n398), .B(n407), .Z(n406) );
  NANDN U517 ( .A(n370), .B(n408), .Z(n407) );
  OR U518 ( .A(n409), .B(n367), .Z(n398) );
  XNOR U519 ( .A(n370), .B(n410), .Z(n367) );
  XNOR U520 ( .A(n396), .B(n411), .Z(n348) );
  XNOR U521 ( .A(n412), .B(n413), .Z(n411) );
  NAND U522 ( .A(n384), .B(n414), .Z(n413) );
  XOR U523 ( .A(n415), .B(n412), .Z(n396) );
  OR U524 ( .A(n392), .B(n416), .Z(n412) );
  XNOR U525 ( .A(n394), .B(n384), .Z(n392) );
  XNOR U526 ( .A(n387), .B(n358), .Z(n384) );
  IV U527 ( .A(n410), .Z(n358) );
  XNOR U528 ( .A(n417), .B(n418), .Z(n410) );
  NAND U529 ( .A(n419), .B(n420), .Z(n418) );
  XOR U530 ( .A(n421), .B(n422), .Z(n387) );
  NAND U531 ( .A(n423), .B(n419), .Z(n422) );
  ANDN U532 ( .B(n394), .A(n424), .Z(n415) );
  XOR U533 ( .A(n352), .B(n370), .Z(n394) );
  XNOR U534 ( .A(n417), .B(n425), .Z(n370) );
  OR U535 ( .A(n426), .B(n427), .Z(n425) );
  NAND U536 ( .A(n428), .B(n429), .Z(n417) );
  ANDN U537 ( .B(n429), .A(n431), .Z(n421) );
  XNOR U538 ( .A(n426), .B(n419), .Z(n429) );
  XNOR U539 ( .A(n432), .B(n433), .Z(n419) );
  XNOR U540 ( .A(n434), .B(n427), .Z(n433) );
  IV U541 ( .A(n435), .Z(n427) );
  XNOR U542 ( .A(n436), .B(n437), .Z(n432) );
  XNOR U543 ( .A(n438), .B(n439), .Z(n437) );
  ANDN U544 ( .B(n435), .A(n436), .Z(n438) );
  NOR U545 ( .A(n426), .B(n436), .Z(n430) );
  XNOR U546 ( .A(n434), .B(n440), .Z(n426) );
  XNOR U547 ( .A(n439), .B(n441), .Z(n440) );
  NAND U548 ( .A(n423), .B(n420), .Z(n441) );
  NANDN U549 ( .A(n431), .B(n428), .Z(n439) );
  XOR U550 ( .A(n420), .B(n435), .Z(n428) );
  XNOR U551 ( .A(n442), .B(n443), .Z(n435) );
  XOR U552 ( .A(n444), .B(n445), .Z(n443) );
  XOR U553 ( .A(n388), .B(n446), .Z(n445) );
  XOR U554 ( .A(n405), .B(n447), .Z(n442) );
  XNOR U555 ( .A(n448), .B(n449), .Z(n447) );
  AND U556 ( .A(n353), .B(n379), .Z(n448) );
  XOR U557 ( .A(n450), .B(n451), .Z(n436) );
  XNOR U558 ( .A(n452), .B(n446), .Z(n451) );
  XOR U559 ( .A(n453), .B(n454), .Z(n446) );
  XNOR U560 ( .A(n455), .B(n456), .Z(n454) );
  NAND U561 ( .A(n414), .B(n383), .Z(n456) );
  XNOR U562 ( .A(n457), .B(n458), .Z(n450) );
  AND U563 ( .A(n408), .B(n369), .Z(n457) );
  XNOR U564 ( .A(n423), .B(n420), .Z(n434) );
  XNOR U565 ( .A(n459), .B(n460), .Z(n420) );
  XNOR U566 ( .A(n461), .B(n462), .Z(n460) );
  XOR U567 ( .A(n452), .B(n379), .Z(n462) );
  XOR U568 ( .A(n353), .B(n463), .Z(n459) );
  XNOR U569 ( .A(n464), .B(n449), .Z(n463) );
  OR U570 ( .A(n390), .B(n404), .Z(n449) );
  XOR U571 ( .A(n353), .B(n465), .Z(n404) );
  XNOR U572 ( .A(n379), .B(n388), .Z(n390) );
  AND U573 ( .A(n388), .B(n405), .Z(n464) );
  XNOR U574 ( .A(n466), .B(n467), .Z(n423) );
  XNOR U575 ( .A(n453), .B(n444), .Z(n467) );
  XNOR U576 ( .A(n468), .B(n357), .Z(n444) );
  IV U577 ( .A(n461), .Z(n453) );
  XOR U578 ( .A(n469), .B(n455), .Z(n461) );
  NANDN U579 ( .A(n416), .B(n393), .Z(n455) );
  XOR U580 ( .A(n395), .B(n383), .Z(n393) );
  XNOR U581 ( .A(n470), .B(n388), .Z(n383) );
  XOR U582 ( .A(n471), .B(n472), .Z(n388) );
  XOR U583 ( .A(n473), .B(n474), .Z(n472) );
  XOR U584 ( .A(n424), .B(n414), .Z(n416) );
  XOR U585 ( .A(n465), .B(n468), .Z(n414) );
  IV U586 ( .A(n405), .Z(n465) );
  XNOR U587 ( .A(n475), .B(n476), .Z(n405) );
  XNOR U588 ( .A(n477), .B(n478), .Z(n476) );
  XOR U589 ( .A(n353), .B(n479), .Z(n475) );
  ANDN U590 ( .B(n395), .A(n424), .Z(n469) );
  XOR U591 ( .A(n353), .B(n480), .Z(n424) );
  XNOR U592 ( .A(n471), .B(n379), .Z(n395) );
  XOR U593 ( .A(n481), .B(n482), .Z(n379) );
  XOR U594 ( .A(n483), .B(n478), .Z(n482) );
  XOR U595 ( .A(state[12]), .B(key[12]), .Z(n478) );
  XNOR U596 ( .A(n452), .B(n484), .Z(n466) );
  XNOR U597 ( .A(n485), .B(n458), .Z(n484) );
  OR U598 ( .A(n368), .B(n409), .Z(n458) );
  XOR U599 ( .A(n408), .B(n468), .Z(n409) );
  XOR U600 ( .A(n369), .B(n470), .Z(n368) );
  IV U601 ( .A(n357), .Z(n470) );
  AND U602 ( .A(n400), .B(n357), .Z(n485) );
  XOR U603 ( .A(n481), .B(n486), .Z(n357) );
  XNOR U604 ( .A(n483), .B(n473), .Z(n486) );
  IV U605 ( .A(n468), .Z(n400) );
  XNOR U606 ( .A(n480), .B(n471), .Z(n452) );
  IV U607 ( .A(n369), .Z(n471) );
  XOR U608 ( .A(n481), .B(n487), .Z(n369) );
  XOR U609 ( .A(n483), .B(n477), .Z(n487) );
  XOR U610 ( .A(state[15]), .B(key[15]), .Z(n477) );
  XNOR U611 ( .A(state[13]), .B(key[13]), .Z(n481) );
  IV U612 ( .A(n408), .Z(n480) );
  XOR U613 ( .A(n488), .B(n474), .Z(n408) );
  XOR U614 ( .A(state[10]), .B(key[10]), .Z(n474) );
  XNOR U615 ( .A(n479), .B(n483), .Z(n488) );
  XOR U616 ( .A(n353), .B(n489), .Z(n483) );
  XNOR U617 ( .A(state[14]), .B(key[14]), .Z(n489) );
  XOR U618 ( .A(state[8]), .B(key[8]), .Z(n353) );
  XOR U619 ( .A(n473), .B(n490), .Z(n479) );
  XNOR U620 ( .A(state[11]), .B(key[11]), .Z(n490) );
  XNOR U621 ( .A(state[9]), .B(key[9]), .Z(n473) );
  XOR U622 ( .A(n491), .B(n492), .Z(out[71]) );
  XNOR U623 ( .A(n493), .B(n494), .Z(n491) );
  XNOR U624 ( .A(key[71]), .B(n495), .Z(n494) );
  XOR U625 ( .A(n496), .B(n497), .Z(out[70]) );
  XNOR U626 ( .A(n498), .B(n499), .Z(n497) );
  XNOR U627 ( .A(key[70]), .B(n500), .Z(n496) );
  XNOR U628 ( .A(n501), .B(n502), .Z(out[6]) );
  XNOR U629 ( .A(key[6]), .B(n503), .Z(n502) );
  XOR U630 ( .A(n504), .B(n505), .Z(out[69]) );
  XNOR U631 ( .A(n506), .B(n507), .Z(n505) );
  XNOR U632 ( .A(n495), .B(n508), .Z(n507) );
  XNOR U633 ( .A(n509), .B(n510), .Z(n495) );
  XNOR U634 ( .A(n511), .B(n512), .Z(n510) );
  NANDN U635 ( .A(n513), .B(n514), .Z(n512) );
  XNOR U636 ( .A(n515), .B(n516), .Z(n504) );
  XOR U637 ( .A(key[69]), .B(n517), .Z(n516) );
  AND U638 ( .A(n518), .B(n519), .Z(n517) );
  XNOR U639 ( .A(n520), .B(n521), .Z(out[68]) );
  XOR U640 ( .A(key[68]), .B(n506), .Z(n521) );
  XOR U641 ( .A(n522), .B(n523), .Z(out[67]) );
  XNOR U642 ( .A(n524), .B(n499), .Z(n523) );
  XNOR U643 ( .A(n525), .B(n526), .Z(n499) );
  XNOR U644 ( .A(n515), .B(n527), .Z(n526) );
  NAND U645 ( .A(n528), .B(n529), .Z(n527) );
  NANDN U646 ( .A(n530), .B(n531), .Z(n515) );
  XNOR U647 ( .A(n532), .B(n533), .Z(n522) );
  XNOR U648 ( .A(key[67]), .B(n498), .Z(n533) );
  XOR U649 ( .A(key[66]), .B(n520), .Z(out[66]) );
  XOR U650 ( .A(n534), .B(n524), .Z(n520) );
  XOR U651 ( .A(n535), .B(n492), .Z(out[65]) );
  XNOR U652 ( .A(n532), .B(n524), .Z(n492) );
  XNOR U653 ( .A(n536), .B(n537), .Z(n524) );
  XNOR U654 ( .A(n538), .B(n539), .Z(n537) );
  NAND U655 ( .A(n540), .B(n519), .Z(n539) );
  XNOR U656 ( .A(n525), .B(n541), .Z(n532) );
  XNOR U657 ( .A(n542), .B(n543), .Z(n541) );
  NANDN U658 ( .A(n513), .B(n544), .Z(n543) );
  XNOR U659 ( .A(n508), .B(n545), .Z(n525) );
  XNOR U660 ( .A(n546), .B(n547), .Z(n545) );
  NANDN U661 ( .A(n548), .B(n549), .Z(n547) );
  XNOR U662 ( .A(key[65]), .B(n493), .Z(n535) );
  XNOR U663 ( .A(n500), .B(n498), .Z(n493) );
  XNOR U664 ( .A(n508), .B(n550), .Z(n498) );
  XOR U665 ( .A(n551), .B(n542), .Z(n550) );
  OR U666 ( .A(n552), .B(n553), .Z(n542) );
  AND U667 ( .A(n554), .B(n555), .Z(n551) );
  XOR U668 ( .A(n556), .B(n546), .Z(n508) );
  NANDN U669 ( .A(n557), .B(n558), .Z(n546) );
  AND U670 ( .A(n559), .B(n560), .Z(n556) );
  IV U671 ( .A(n534), .Z(n500) );
  XNOR U672 ( .A(n506), .B(n561), .Z(out[64]) );
  XNOR U673 ( .A(key[64]), .B(n534), .Z(n561) );
  XOR U674 ( .A(n536), .B(n562), .Z(n534) );
  XOR U675 ( .A(n563), .B(n511), .Z(n562) );
  OR U676 ( .A(n564), .B(n552), .Z(n511) );
  XNOR U677 ( .A(n513), .B(n565), .Z(n552) );
  AND U678 ( .A(n566), .B(n555), .Z(n563) );
  IV U679 ( .A(n565), .Z(n555) );
  XNOR U680 ( .A(n509), .B(n567), .Z(n506) );
  XOR U681 ( .A(n568), .B(n538), .Z(n567) );
  NANDN U682 ( .A(n569), .B(n531), .Z(n538) );
  XOR U683 ( .A(n529), .B(n519), .Z(n531) );
  AND U684 ( .A(n529), .B(n570), .Z(n568) );
  XNOR U685 ( .A(n536), .B(n571), .Z(n509) );
  XNOR U686 ( .A(n572), .B(n573), .Z(n571) );
  NANDN U687 ( .A(n548), .B(n574), .Z(n573) );
  XOR U688 ( .A(n575), .B(n572), .Z(n536) );
  OR U689 ( .A(n557), .B(n576), .Z(n572) );
  XNOR U690 ( .A(n577), .B(n548), .Z(n557) );
  XOR U691 ( .A(n578), .B(n579), .Z(n519) );
  NANDN U692 ( .A(n580), .B(n581), .Z(n579) );
  XOR U693 ( .A(n582), .B(n583), .Z(n565) );
  NANDN U694 ( .A(n580), .B(n584), .Z(n583) );
  NOR U695 ( .A(n577), .B(n585), .Z(n575) );
  IV U696 ( .A(n560), .Z(n577) );
  XNOR U697 ( .A(n513), .B(n529), .Z(n560) );
  XNOR U698 ( .A(n586), .B(n578), .Z(n529) );
  NANDN U699 ( .A(n587), .B(n588), .Z(n578) );
  XNOR U700 ( .A(n581), .B(n589), .Z(n588) );
  AND U701 ( .A(n590), .B(n591), .Z(n586) );
  ANDN U702 ( .B(n593), .A(n587), .Z(n582) );
  XOR U703 ( .A(n594), .B(n595), .Z(n580) );
  XNOR U704 ( .A(n590), .B(n596), .Z(n595) );
  XNOR U705 ( .A(n597), .B(n598), .Z(n594) );
  XNOR U706 ( .A(n599), .B(n600), .Z(n598) );
  AND U707 ( .A(n596), .B(n590), .Z(n599) );
  AND U708 ( .A(n596), .B(n591), .Z(n592) );
  XOR U709 ( .A(n597), .B(n601), .Z(n591) );
  XOR U710 ( .A(n602), .B(n600), .Z(n601) );
  NAND U711 ( .A(n593), .B(n603), .Z(n600) );
  XOR U712 ( .A(n581), .B(n590), .Z(n603) );
  IV U713 ( .A(n589), .Z(n590) );
  XOR U714 ( .A(n604), .B(n605), .Z(n589) );
  XNOR U715 ( .A(n606), .B(n607), .Z(n605) );
  XNOR U716 ( .A(n554), .B(n608), .Z(n607) );
  XOR U717 ( .A(n566), .B(n609), .Z(n604) );
  XNOR U718 ( .A(n610), .B(n611), .Z(n609) );
  AND U719 ( .A(n514), .B(n544), .Z(n610) );
  XOR U720 ( .A(n584), .B(n596), .Z(n593) );
  AND U721 ( .A(n581), .B(n584), .Z(n602) );
  XNOR U722 ( .A(n581), .B(n584), .Z(n597) );
  XNOR U723 ( .A(n612), .B(n613), .Z(n584) );
  XOR U724 ( .A(n614), .B(n608), .Z(n613) );
  XNOR U725 ( .A(n615), .B(n518), .Z(n608) );
  XOR U726 ( .A(n616), .B(n617), .Z(n612) );
  XNOR U727 ( .A(n618), .B(n619), .Z(n617) );
  AND U728 ( .A(n540), .B(n518), .Z(n618) );
  XNOR U729 ( .A(n620), .B(n621), .Z(n581) );
  XNOR U730 ( .A(n544), .B(n616), .Z(n622) );
  XOR U731 ( .A(n514), .B(n623), .Z(n620) );
  XNOR U732 ( .A(n624), .B(n611), .Z(n623) );
  OR U733 ( .A(n553), .B(n564), .Z(n611) );
  XNOR U734 ( .A(n514), .B(n566), .Z(n564) );
  XOR U735 ( .A(n544), .B(n625), .Z(n553) );
  AND U736 ( .A(n566), .B(n554), .Z(n624) );
  XNOR U737 ( .A(n626), .B(n627), .Z(n596) );
  XNOR U738 ( .A(n614), .B(n606), .Z(n627) );
  XOR U739 ( .A(n616), .B(n628), .Z(n606) );
  XNOR U740 ( .A(n629), .B(n630), .Z(n628) );
  NAND U741 ( .A(n574), .B(n549), .Z(n630) );
  XNOR U742 ( .A(n631), .B(n629), .Z(n616) );
  NANDN U743 ( .A(n576), .B(n558), .Z(n629) );
  XOR U744 ( .A(n559), .B(n549), .Z(n558) );
  XOR U745 ( .A(n625), .B(n632), .Z(n549) );
  IV U746 ( .A(n554), .Z(n625) );
  XNOR U747 ( .A(n528), .B(n633), .Z(n554) );
  XNOR U748 ( .A(n634), .B(n635), .Z(n633) );
  XOR U749 ( .A(n585), .B(n574), .Z(n576) );
  XNOR U750 ( .A(n636), .B(n637), .Z(n566) );
  XNOR U751 ( .A(n638), .B(n639), .Z(n637) );
  XOR U752 ( .A(n514), .B(n640), .Z(n636) );
  ANDN U753 ( .B(n559), .A(n585), .Z(n631) );
  XOR U754 ( .A(n514), .B(n641), .Z(n585) );
  XOR U755 ( .A(n642), .B(n643), .Z(n544) );
  XNOR U756 ( .A(n644), .B(n639), .Z(n643) );
  XOR U757 ( .A(state[100]), .B(key[100]), .Z(n639) );
  XOR U758 ( .A(n641), .B(n528), .Z(n614) );
  IV U759 ( .A(n570), .Z(n641) );
  XNOR U760 ( .A(n645), .B(n619), .Z(n626) );
  OR U761 ( .A(n530), .B(n569), .Z(n619) );
  XNOR U762 ( .A(n570), .B(n540), .Z(n569) );
  IV U763 ( .A(n615), .Z(n540) );
  XOR U764 ( .A(n528), .B(n632), .Z(n530) );
  IV U765 ( .A(n518), .Z(n632) );
  XOR U766 ( .A(n642), .B(n646), .Z(n518) );
  XOR U767 ( .A(n644), .B(n635), .Z(n646) );
  AND U768 ( .A(n528), .B(n570), .Z(n645) );
  XOR U769 ( .A(n640), .B(n634), .Z(n647) );
  XNOR U770 ( .A(state[98]), .B(key[98]), .Z(n634) );
  XOR U771 ( .A(n635), .B(n648), .Z(n640) );
  XNOR U772 ( .A(state[99]), .B(key[99]), .Z(n648) );
  XNOR U773 ( .A(state[97]), .B(key[97]), .Z(n635) );
  XOR U774 ( .A(n642), .B(n649), .Z(n528) );
  XNOR U775 ( .A(n644), .B(n638), .Z(n649) );
  XOR U776 ( .A(state[103]), .B(key[103]), .Z(n638) );
  XNOR U777 ( .A(n514), .B(n650), .Z(n644) );
  XNOR U778 ( .A(state[102]), .B(key[102]), .Z(n650) );
  XOR U779 ( .A(state[96]), .B(key[96]), .Z(n514) );
  XNOR U780 ( .A(state[101]), .B(key[101]), .Z(n642) );
  XOR U781 ( .A(n651), .B(n652), .Z(out[63]) );
  XOR U782 ( .A(n653), .B(n654), .Z(n651) );
  XOR U783 ( .A(key[63]), .B(n655), .Z(n654) );
  XNOR U784 ( .A(n656), .B(n657), .Z(out[62]) );
  XNOR U785 ( .A(key[62]), .B(n658), .Z(n657) );
  XOR U786 ( .A(n659), .B(n660), .Z(out[61]) );
  XNOR U787 ( .A(n661), .B(n662), .Z(n660) );
  XOR U788 ( .A(n653), .B(n663), .Z(n662) );
  XOR U789 ( .A(n664), .B(n665), .Z(n653) );
  XNOR U790 ( .A(n666), .B(n667), .Z(n665) );
  NANDN U791 ( .A(n668), .B(n669), .Z(n667) );
  XOR U792 ( .A(n670), .B(n671), .Z(n659) );
  XOR U793 ( .A(key[61]), .B(n672), .Z(n671) );
  ANDN U794 ( .B(n673), .A(n674), .Z(n670) );
  XNOR U795 ( .A(n675), .B(n676), .Z(out[60]) );
  XOR U796 ( .A(key[60]), .B(n661), .Z(n676) );
  XOR U797 ( .A(n677), .B(n678), .Z(out[5]) );
  XNOR U798 ( .A(n679), .B(n680), .Z(n678) );
  XOR U799 ( .A(n330), .B(n681), .Z(n680) );
  XOR U800 ( .A(n682), .B(n683), .Z(n330) );
  XNOR U801 ( .A(n684), .B(n685), .Z(n683) );
  NANDN U802 ( .A(n686), .B(n687), .Z(n685) );
  XOR U803 ( .A(n688), .B(n689), .Z(n677) );
  XOR U804 ( .A(key[5]), .B(n690), .Z(n689) );
  ANDN U805 ( .B(n691), .A(n692), .Z(n688) );
  XOR U806 ( .A(n693), .B(n694), .Z(out[59]) );
  XOR U807 ( .A(n695), .B(n656), .Z(n694) );
  XNOR U808 ( .A(n696), .B(n697), .Z(n656) );
  XNOR U809 ( .A(n698), .B(n672), .Z(n697) );
  NOR U810 ( .A(n699), .B(n700), .Z(n672) );
  ANDN U811 ( .B(n701), .A(n702), .Z(n698) );
  XNOR U812 ( .A(n703), .B(n704), .Z(n693) );
  XNOR U813 ( .A(key[59]), .B(n705), .Z(n704) );
  XOR U814 ( .A(key[58]), .B(n675), .Z(out[58]) );
  XOR U815 ( .A(n655), .B(n706), .Z(n675) );
  XOR U816 ( .A(n707), .B(n652), .Z(out[57]) );
  XOR U817 ( .A(n696), .B(n708), .Z(n695) );
  XNOR U818 ( .A(n709), .B(n710), .Z(n708) );
  NANDN U819 ( .A(n668), .B(n711), .Z(n710) );
  XNOR U820 ( .A(n663), .B(n712), .Z(n696) );
  XNOR U821 ( .A(n713), .B(n714), .Z(n712) );
  NANDN U822 ( .A(n715), .B(n716), .Z(n714) );
  XOR U823 ( .A(n706), .B(n703), .Z(n658) );
  XNOR U824 ( .A(n663), .B(n717), .Z(n703) );
  XNOR U825 ( .A(n709), .B(n718), .Z(n717) );
  NAND U826 ( .A(n719), .B(n720), .Z(n718) );
  OR U827 ( .A(n721), .B(n722), .Z(n709) );
  XOR U828 ( .A(n723), .B(n713), .Z(n663) );
  NANDN U829 ( .A(n724), .B(n725), .Z(n713) );
  AND U830 ( .A(n726), .B(n727), .Z(n723) );
  XOR U831 ( .A(key[57]), .B(n655), .Z(n707) );
  IV U832 ( .A(n705), .Z(n655) );
  XNOR U833 ( .A(n728), .B(n729), .Z(n705) );
  XNOR U834 ( .A(n730), .B(n731), .Z(n729) );
  NANDN U835 ( .A(n674), .B(n732), .Z(n731) );
  XNOR U836 ( .A(n661), .B(n733), .Z(out[56]) );
  XOR U837 ( .A(key[56]), .B(n706), .Z(n733) );
  XNOR U838 ( .A(n728), .B(n734), .Z(n706) );
  XOR U839 ( .A(n735), .B(n666), .Z(n734) );
  OR U840 ( .A(n736), .B(n721), .Z(n666) );
  XNOR U841 ( .A(n668), .B(n737), .Z(n721) );
  AND U842 ( .A(n738), .B(n719), .Z(n735) );
  XNOR U843 ( .A(n664), .B(n739), .Z(n661) );
  XOR U844 ( .A(n740), .B(n730), .Z(n739) );
  OR U845 ( .A(n741), .B(n699), .Z(n730) );
  XNOR U846 ( .A(n702), .B(n674), .Z(n699) );
  NOR U847 ( .A(n742), .B(n702), .Z(n740) );
  XNOR U848 ( .A(n728), .B(n743), .Z(n664) );
  XNOR U849 ( .A(n744), .B(n745), .Z(n743) );
  NANDN U850 ( .A(n715), .B(n746), .Z(n745) );
  XOR U851 ( .A(n747), .B(n744), .Z(n728) );
  OR U852 ( .A(n724), .B(n748), .Z(n744) );
  XOR U853 ( .A(n726), .B(n715), .Z(n724) );
  XNOR U854 ( .A(n737), .B(n674), .Z(n715) );
  XOR U855 ( .A(n749), .B(n750), .Z(n674) );
  NANDN U856 ( .A(n751), .B(n752), .Z(n750) );
  IV U857 ( .A(n719), .Z(n737) );
  XOR U858 ( .A(n753), .B(n754), .Z(n719) );
  NANDN U859 ( .A(n751), .B(n755), .Z(n754) );
  ANDN U860 ( .B(n726), .A(n756), .Z(n747) );
  XOR U861 ( .A(n702), .B(n668), .Z(n726) );
  XOR U862 ( .A(n757), .B(n753), .Z(n668) );
  NANDN U863 ( .A(n758), .B(n759), .Z(n753) );
  AND U864 ( .A(n760), .B(n761), .Z(n757) );
  ANDN U865 ( .B(n763), .A(n758), .Z(n749) );
  XOR U866 ( .A(n764), .B(n765), .Z(n751) );
  XNOR U867 ( .A(n767), .B(n768), .Z(n764) );
  XNOR U868 ( .A(n769), .B(n770), .Z(n768) );
  AND U869 ( .A(n771), .B(n760), .Z(n769) );
  AND U870 ( .A(n771), .B(n761), .Z(n762) );
  XOR U871 ( .A(n767), .B(n772), .Z(n761) );
  XOR U872 ( .A(n773), .B(n770), .Z(n772) );
  NAND U873 ( .A(n759), .B(n763), .Z(n770) );
  XOR U874 ( .A(n752), .B(n771), .Z(n763) );
  XOR U875 ( .A(n755), .B(n760), .Z(n759) );
  XNOR U876 ( .A(n774), .B(n775), .Z(n760) );
  XOR U877 ( .A(n776), .B(n777), .Z(n775) );
  XNOR U878 ( .A(n778), .B(n779), .Z(n774) );
  ANDN U879 ( .B(n701), .A(n742), .Z(n778) );
  AND U880 ( .A(n752), .B(n755), .Z(n773) );
  XNOR U881 ( .A(n752), .B(n755), .Z(n767) );
  XNOR U882 ( .A(n780), .B(n781), .Z(n755) );
  XOR U883 ( .A(n782), .B(n783), .Z(n781) );
  XOR U884 ( .A(n776), .B(n784), .Z(n780) );
  XNOR U885 ( .A(n785), .B(n779), .Z(n784) );
  OR U886 ( .A(n700), .B(n741), .Z(n779) );
  XOR U887 ( .A(n742), .B(n732), .Z(n741) );
  XOR U888 ( .A(n786), .B(n673), .Z(n700) );
  AND U889 ( .A(n673), .B(n732), .Z(n785) );
  XNOR U890 ( .A(n787), .B(n788), .Z(n752) );
  XOR U891 ( .A(n789), .B(n790), .Z(n788) );
  XNOR U892 ( .A(n711), .B(n776), .Z(n790) );
  XNOR U893 ( .A(n742), .B(n701), .Z(n776) );
  XOR U894 ( .A(n669), .B(n791), .Z(n787) );
  XNOR U895 ( .A(n792), .B(n793), .Z(n791) );
  AND U896 ( .A(n720), .B(n738), .Z(n792) );
  IV U897 ( .A(n766), .Z(n771) );
  XOR U898 ( .A(n794), .B(n795), .Z(n766) );
  XNOR U899 ( .A(n777), .B(n796), .Z(n795) );
  XNOR U900 ( .A(n720), .B(n783), .Z(n796) );
  XOR U901 ( .A(n789), .B(n797), .Z(n777) );
  XNOR U902 ( .A(n798), .B(n799), .Z(n797) );
  NAND U903 ( .A(n716), .B(n746), .Z(n799) );
  IV U904 ( .A(n782), .Z(n789) );
  XOR U905 ( .A(n800), .B(n798), .Z(n782) );
  NANDN U906 ( .A(n748), .B(n725), .Z(n798) );
  XOR U907 ( .A(n720), .B(n673), .Z(n716) );
  XOR U908 ( .A(n801), .B(n802), .Z(n673) );
  XOR U909 ( .A(n803), .B(n804), .Z(n802) );
  XOR U910 ( .A(n756), .B(n746), .Z(n748) );
  ANDN U911 ( .B(n727), .A(n756), .Z(n800) );
  XNOR U912 ( .A(n805), .B(n742), .Z(n756) );
  XNOR U913 ( .A(n806), .B(n807), .Z(n742) );
  XOR U914 ( .A(n808), .B(n803), .Z(n806) );
  XOR U915 ( .A(n738), .B(n809), .Z(n794) );
  XNOR U916 ( .A(n810), .B(n793), .Z(n809) );
  OR U917 ( .A(n722), .B(n736), .Z(n793) );
  XNOR U918 ( .A(n669), .B(n738), .Z(n736) );
  XNOR U919 ( .A(n711), .B(n720), .Z(n722) );
  XOR U920 ( .A(n786), .B(n811), .Z(n720) );
  XOR U921 ( .A(state[58]), .B(key[58]), .Z(n807) );
  IV U922 ( .A(n701), .Z(n786) );
  XOR U923 ( .A(n801), .B(n812), .Z(n701) );
  XNOR U924 ( .A(n803), .B(n813), .Z(n812) );
  AND U925 ( .A(n669), .B(n711), .Z(n810) );
  XOR U926 ( .A(n801), .B(n814), .Z(n711) );
  XNOR U927 ( .A(n803), .B(n815), .Z(n814) );
  XOR U928 ( .A(n805), .B(n816), .Z(n803) );
  XNOR U929 ( .A(state[62]), .B(key[62]), .Z(n816) );
  XNOR U930 ( .A(state[61]), .B(key[61]), .Z(n801) );
  XNOR U931 ( .A(n817), .B(n818), .Z(n738) );
  XNOR U932 ( .A(n815), .B(n813), .Z(n818) );
  XOR U933 ( .A(state[63]), .B(key[63]), .Z(n813) );
  XOR U934 ( .A(state[60]), .B(key[60]), .Z(n815) );
  XOR U935 ( .A(n669), .B(n808), .Z(n817) );
  XOR U936 ( .A(n804), .B(n819), .Z(n808) );
  XNOR U937 ( .A(state[59]), .B(key[59]), .Z(n819) );
  XNOR U938 ( .A(state[57]), .B(key[57]), .Z(n804) );
  IV U939 ( .A(n805), .Z(n669) );
  XNOR U940 ( .A(state[56]), .B(key[56]), .Z(n805) );
  XOR U941 ( .A(n820), .B(n821), .Z(out[55]) );
  XOR U942 ( .A(n822), .B(n823), .Z(n820) );
  XOR U943 ( .A(key[55]), .B(n824), .Z(n823) );
  XNOR U944 ( .A(n825), .B(n826), .Z(out[54]) );
  XNOR U945 ( .A(key[54]), .B(n827), .Z(n826) );
  XOR U946 ( .A(n828), .B(n829), .Z(out[53]) );
  XNOR U947 ( .A(n830), .B(n831), .Z(n829) );
  XOR U948 ( .A(n822), .B(n832), .Z(n831) );
  XOR U949 ( .A(n833), .B(n834), .Z(n822) );
  XNOR U950 ( .A(n835), .B(n836), .Z(n834) );
  NANDN U951 ( .A(n837), .B(n838), .Z(n836) );
  XOR U952 ( .A(n839), .B(n840), .Z(n828) );
  XOR U953 ( .A(key[53]), .B(n841), .Z(n840) );
  ANDN U954 ( .B(n842), .A(n843), .Z(n839) );
  XNOR U955 ( .A(n844), .B(n845), .Z(out[52]) );
  XOR U956 ( .A(key[52]), .B(n830), .Z(n845) );
  XOR U957 ( .A(n846), .B(n847), .Z(out[51]) );
  XOR U958 ( .A(n848), .B(n825), .Z(n847) );
  XNOR U959 ( .A(n849), .B(n850), .Z(n825) );
  XNOR U960 ( .A(n851), .B(n841), .Z(n850) );
  NOR U961 ( .A(n852), .B(n853), .Z(n841) );
  ANDN U962 ( .B(n854), .A(n855), .Z(n851) );
  XNOR U963 ( .A(n856), .B(n857), .Z(n846) );
  XNOR U964 ( .A(key[51]), .B(n858), .Z(n857) );
  XOR U965 ( .A(key[50]), .B(n844), .Z(out[50]) );
  XOR U966 ( .A(n824), .B(n859), .Z(n844) );
  XNOR U967 ( .A(n860), .B(n861), .Z(out[4]) );
  XOR U968 ( .A(key[4]), .B(n679), .Z(n861) );
  XOR U969 ( .A(n862), .B(n821), .Z(out[49]) );
  XOR U970 ( .A(n849), .B(n863), .Z(n848) );
  XNOR U971 ( .A(n864), .B(n865), .Z(n863) );
  NANDN U972 ( .A(n837), .B(n866), .Z(n865) );
  XNOR U973 ( .A(n832), .B(n867), .Z(n849) );
  XNOR U974 ( .A(n868), .B(n869), .Z(n867) );
  NANDN U975 ( .A(n870), .B(n871), .Z(n869) );
  XOR U976 ( .A(n859), .B(n856), .Z(n827) );
  XNOR U977 ( .A(n832), .B(n872), .Z(n856) );
  XNOR U978 ( .A(n864), .B(n873), .Z(n872) );
  NAND U979 ( .A(n874), .B(n875), .Z(n873) );
  OR U980 ( .A(n876), .B(n877), .Z(n864) );
  XOR U981 ( .A(n878), .B(n868), .Z(n832) );
  NANDN U982 ( .A(n879), .B(n880), .Z(n868) );
  AND U983 ( .A(n881), .B(n882), .Z(n878) );
  XOR U984 ( .A(key[49]), .B(n824), .Z(n862) );
  IV U985 ( .A(n858), .Z(n824) );
  XNOR U986 ( .A(n883), .B(n884), .Z(n858) );
  XNOR U987 ( .A(n885), .B(n886), .Z(n884) );
  NANDN U988 ( .A(n843), .B(n887), .Z(n886) );
  XNOR U989 ( .A(n830), .B(n888), .Z(out[48]) );
  XOR U990 ( .A(key[48]), .B(n859), .Z(n888) );
  XNOR U991 ( .A(n883), .B(n889), .Z(n859) );
  XOR U992 ( .A(n890), .B(n835), .Z(n889) );
  OR U993 ( .A(n891), .B(n876), .Z(n835) );
  XNOR U994 ( .A(n837), .B(n892), .Z(n876) );
  AND U995 ( .A(n893), .B(n874), .Z(n890) );
  XNOR U996 ( .A(n833), .B(n894), .Z(n830) );
  XOR U997 ( .A(n895), .B(n885), .Z(n894) );
  OR U998 ( .A(n896), .B(n852), .Z(n885) );
  XNOR U999 ( .A(n855), .B(n843), .Z(n852) );
  NOR U1000 ( .A(n897), .B(n855), .Z(n895) );
  XNOR U1001 ( .A(n883), .B(n898), .Z(n833) );
  XNOR U1002 ( .A(n899), .B(n900), .Z(n898) );
  NANDN U1003 ( .A(n870), .B(n901), .Z(n900) );
  XOR U1004 ( .A(n902), .B(n899), .Z(n883) );
  OR U1005 ( .A(n879), .B(n903), .Z(n899) );
  XOR U1006 ( .A(n881), .B(n870), .Z(n879) );
  XNOR U1007 ( .A(n892), .B(n843), .Z(n870) );
  XOR U1008 ( .A(n904), .B(n905), .Z(n843) );
  NANDN U1009 ( .A(n906), .B(n907), .Z(n905) );
  IV U1010 ( .A(n874), .Z(n892) );
  XOR U1011 ( .A(n908), .B(n909), .Z(n874) );
  NANDN U1012 ( .A(n906), .B(n910), .Z(n909) );
  ANDN U1013 ( .B(n881), .A(n911), .Z(n902) );
  XOR U1014 ( .A(n855), .B(n837), .Z(n881) );
  XOR U1015 ( .A(n912), .B(n908), .Z(n837) );
  NANDN U1016 ( .A(n913), .B(n914), .Z(n908) );
  AND U1017 ( .A(n915), .B(n916), .Z(n912) );
  ANDN U1018 ( .B(n918), .A(n913), .Z(n904) );
  XOR U1019 ( .A(n919), .B(n920), .Z(n906) );
  XNOR U1020 ( .A(n922), .B(n923), .Z(n919) );
  XNOR U1021 ( .A(n924), .B(n925), .Z(n923) );
  AND U1022 ( .A(n926), .B(n915), .Z(n924) );
  AND U1023 ( .A(n926), .B(n916), .Z(n917) );
  XOR U1024 ( .A(n922), .B(n927), .Z(n916) );
  XOR U1025 ( .A(n928), .B(n925), .Z(n927) );
  NAND U1026 ( .A(n914), .B(n918), .Z(n925) );
  XOR U1027 ( .A(n907), .B(n926), .Z(n918) );
  XOR U1028 ( .A(n910), .B(n915), .Z(n914) );
  XNOR U1029 ( .A(n929), .B(n930), .Z(n915) );
  XOR U1030 ( .A(n931), .B(n932), .Z(n930) );
  XNOR U1031 ( .A(n933), .B(n934), .Z(n929) );
  ANDN U1032 ( .B(n854), .A(n897), .Z(n933) );
  AND U1033 ( .A(n907), .B(n910), .Z(n928) );
  XNOR U1034 ( .A(n907), .B(n910), .Z(n922) );
  XNOR U1035 ( .A(n935), .B(n936), .Z(n910) );
  XOR U1036 ( .A(n937), .B(n938), .Z(n936) );
  XOR U1037 ( .A(n931), .B(n939), .Z(n935) );
  XNOR U1038 ( .A(n940), .B(n934), .Z(n939) );
  OR U1039 ( .A(n853), .B(n896), .Z(n934) );
  XOR U1040 ( .A(n897), .B(n887), .Z(n896) );
  XOR U1041 ( .A(n941), .B(n842), .Z(n853) );
  AND U1042 ( .A(n842), .B(n887), .Z(n940) );
  XNOR U1043 ( .A(n942), .B(n943), .Z(n907) );
  XOR U1044 ( .A(n944), .B(n945), .Z(n943) );
  XNOR U1045 ( .A(n866), .B(n931), .Z(n945) );
  XNOR U1046 ( .A(n897), .B(n854), .Z(n931) );
  XOR U1047 ( .A(n838), .B(n946), .Z(n942) );
  XNOR U1048 ( .A(n947), .B(n948), .Z(n946) );
  AND U1049 ( .A(n875), .B(n893), .Z(n947) );
  IV U1050 ( .A(n921), .Z(n926) );
  XOR U1051 ( .A(n949), .B(n950), .Z(n921) );
  XNOR U1052 ( .A(n932), .B(n951), .Z(n950) );
  XNOR U1053 ( .A(n875), .B(n938), .Z(n951) );
  XOR U1054 ( .A(n944), .B(n952), .Z(n932) );
  XNOR U1055 ( .A(n953), .B(n954), .Z(n952) );
  NAND U1056 ( .A(n871), .B(n901), .Z(n954) );
  IV U1057 ( .A(n937), .Z(n944) );
  XOR U1058 ( .A(n955), .B(n953), .Z(n937) );
  NANDN U1059 ( .A(n903), .B(n880), .Z(n953) );
  XOR U1060 ( .A(n875), .B(n842), .Z(n871) );
  XOR U1061 ( .A(n956), .B(n957), .Z(n842) );
  XOR U1062 ( .A(n958), .B(n959), .Z(n957) );
  XOR U1063 ( .A(n911), .B(n901), .Z(n903) );
  ANDN U1064 ( .B(n882), .A(n911), .Z(n955) );
  XNOR U1065 ( .A(n960), .B(n897), .Z(n911) );
  XNOR U1066 ( .A(n961), .B(n962), .Z(n897) );
  XOR U1067 ( .A(n963), .B(n958), .Z(n961) );
  XOR U1068 ( .A(n893), .B(n964), .Z(n949) );
  XNOR U1069 ( .A(n965), .B(n948), .Z(n964) );
  OR U1070 ( .A(n877), .B(n891), .Z(n948) );
  XNOR U1071 ( .A(n838), .B(n893), .Z(n891) );
  XNOR U1072 ( .A(n866), .B(n875), .Z(n877) );
  XOR U1073 ( .A(n941), .B(n966), .Z(n875) );
  XOR U1074 ( .A(state[18]), .B(key[18]), .Z(n962) );
  IV U1075 ( .A(n854), .Z(n941) );
  XOR U1076 ( .A(n956), .B(n967), .Z(n854) );
  XNOR U1077 ( .A(n958), .B(n968), .Z(n967) );
  AND U1078 ( .A(n838), .B(n866), .Z(n965) );
  XOR U1079 ( .A(n956), .B(n969), .Z(n866) );
  XNOR U1080 ( .A(n958), .B(n970), .Z(n969) );
  XOR U1081 ( .A(n960), .B(n971), .Z(n958) );
  XNOR U1082 ( .A(state[22]), .B(key[22]), .Z(n971) );
  XNOR U1083 ( .A(state[21]), .B(key[21]), .Z(n956) );
  XNOR U1084 ( .A(n972), .B(n973), .Z(n893) );
  XNOR U1085 ( .A(n970), .B(n968), .Z(n973) );
  XOR U1086 ( .A(state[23]), .B(key[23]), .Z(n968) );
  XOR U1087 ( .A(state[20]), .B(key[20]), .Z(n970) );
  XOR U1088 ( .A(n838), .B(n963), .Z(n972) );
  XOR U1089 ( .A(n959), .B(n974), .Z(n963) );
  XNOR U1090 ( .A(state[19]), .B(key[19]), .Z(n974) );
  XNOR U1091 ( .A(state[17]), .B(key[17]), .Z(n959) );
  IV U1092 ( .A(n960), .Z(n838) );
  XNOR U1093 ( .A(state[16]), .B(key[16]), .Z(n960) );
  XOR U1094 ( .A(n975), .B(n976), .Z(out[47]) );
  XOR U1095 ( .A(n977), .B(n978), .Z(n975) );
  XNOR U1096 ( .A(key[47]), .B(n979), .Z(n978) );
  XNOR U1097 ( .A(n980), .B(n981), .Z(out[46]) );
  XNOR U1098 ( .A(key[46]), .B(n982), .Z(n981) );
  XOR U1099 ( .A(n983), .B(n984), .Z(out[45]) );
  XNOR U1100 ( .A(n985), .B(n986), .Z(n984) );
  XOR U1101 ( .A(n977), .B(n987), .Z(n986) );
  XOR U1102 ( .A(n988), .B(n989), .Z(n977) );
  XNOR U1103 ( .A(n990), .B(n991), .Z(n989) );
  NANDN U1104 ( .A(n992), .B(n993), .Z(n991) );
  XOR U1105 ( .A(n994), .B(n995), .Z(n983) );
  XOR U1106 ( .A(key[45]), .B(n996), .Z(n995) );
  ANDN U1107 ( .B(n997), .A(n998), .Z(n994) );
  XNOR U1108 ( .A(n999), .B(n1000), .Z(out[44]) );
  XOR U1109 ( .A(key[44]), .B(n985), .Z(n1000) );
  XOR U1110 ( .A(n1001), .B(n1002), .Z(out[43]) );
  XOR U1111 ( .A(n1003), .B(n980), .Z(n1002) );
  XNOR U1112 ( .A(n1004), .B(n1005), .Z(n980) );
  XNOR U1113 ( .A(n1006), .B(n996), .Z(n1005) );
  NOR U1114 ( .A(n1007), .B(n1008), .Z(n996) );
  ANDN U1115 ( .B(n1009), .A(n1010), .Z(n1006) );
  XNOR U1116 ( .A(n1011), .B(n1012), .Z(n1001) );
  XNOR U1117 ( .A(key[43]), .B(n979), .Z(n1012) );
  XOR U1118 ( .A(key[42]), .B(n999), .Z(out[42]) );
  XNOR U1119 ( .A(n979), .B(n1013), .Z(n999) );
  XOR U1120 ( .A(n1014), .B(n976), .Z(out[41]) );
  XOR U1121 ( .A(n1004), .B(n1015), .Z(n1003) );
  XNOR U1122 ( .A(n1016), .B(n1017), .Z(n1015) );
  NANDN U1123 ( .A(n992), .B(n1018), .Z(n1017) );
  XNOR U1124 ( .A(n987), .B(n1019), .Z(n1004) );
  XNOR U1125 ( .A(n1020), .B(n1021), .Z(n1019) );
  NANDN U1126 ( .A(n1022), .B(n1023), .Z(n1021) );
  XOR U1127 ( .A(n1013), .B(n1011), .Z(n982) );
  XNOR U1128 ( .A(n987), .B(n1024), .Z(n1011) );
  XNOR U1129 ( .A(n1016), .B(n1025), .Z(n1024) );
  NAND U1130 ( .A(n1026), .B(n1027), .Z(n1025) );
  OR U1131 ( .A(n1028), .B(n1029), .Z(n1016) );
  XOR U1132 ( .A(n1030), .B(n1020), .Z(n987) );
  NANDN U1133 ( .A(n1031), .B(n1032), .Z(n1020) );
  AND U1134 ( .A(n1033), .B(n1034), .Z(n1030) );
  XNOR U1135 ( .A(key[41]), .B(n979), .Z(n1014) );
  XNOR U1136 ( .A(n1035), .B(n1036), .Z(n979) );
  XNOR U1137 ( .A(n1037), .B(n1038), .Z(n1036) );
  NANDN U1138 ( .A(n998), .B(n1039), .Z(n1038) );
  XNOR U1139 ( .A(n985), .B(n1040), .Z(out[40]) );
  XOR U1140 ( .A(key[40]), .B(n1013), .Z(n1040) );
  XNOR U1141 ( .A(n1035), .B(n1041), .Z(n1013) );
  XOR U1142 ( .A(n1042), .B(n990), .Z(n1041) );
  OR U1143 ( .A(n1043), .B(n1028), .Z(n990) );
  XNOR U1144 ( .A(n992), .B(n1044), .Z(n1028) );
  AND U1145 ( .A(n1045), .B(n1026), .Z(n1042) );
  XNOR U1146 ( .A(n988), .B(n1046), .Z(n985) );
  XOR U1147 ( .A(n1047), .B(n1037), .Z(n1046) );
  OR U1148 ( .A(n1048), .B(n1007), .Z(n1037) );
  XNOR U1149 ( .A(n1010), .B(n998), .Z(n1007) );
  NOR U1150 ( .A(n1049), .B(n1010), .Z(n1047) );
  XNOR U1151 ( .A(n1035), .B(n1050), .Z(n988) );
  XNOR U1152 ( .A(n1051), .B(n1052), .Z(n1050) );
  NANDN U1153 ( .A(n1022), .B(n1053), .Z(n1052) );
  XOR U1154 ( .A(n1054), .B(n1051), .Z(n1035) );
  OR U1155 ( .A(n1031), .B(n1055), .Z(n1051) );
  XOR U1156 ( .A(n1033), .B(n1022), .Z(n1031) );
  XNOR U1157 ( .A(n1044), .B(n998), .Z(n1022) );
  XOR U1158 ( .A(n1056), .B(n1057), .Z(n998) );
  NANDN U1159 ( .A(n1058), .B(n1059), .Z(n1057) );
  IV U1160 ( .A(n1026), .Z(n1044) );
  XOR U1161 ( .A(n1060), .B(n1061), .Z(n1026) );
  NANDN U1162 ( .A(n1058), .B(n1062), .Z(n1061) );
  ANDN U1163 ( .B(n1033), .A(n1063), .Z(n1054) );
  XOR U1164 ( .A(n1010), .B(n992), .Z(n1033) );
  XOR U1165 ( .A(n1064), .B(n1060), .Z(n992) );
  NANDN U1166 ( .A(n1065), .B(n1066), .Z(n1060) );
  AND U1167 ( .A(n1067), .B(n1068), .Z(n1064) );
  ANDN U1168 ( .B(n1070), .A(n1065), .Z(n1056) );
  XOR U1169 ( .A(n1071), .B(n1072), .Z(n1058) );
  XNOR U1170 ( .A(n1074), .B(n1075), .Z(n1071) );
  XNOR U1171 ( .A(n1076), .B(n1077), .Z(n1075) );
  AND U1172 ( .A(n1078), .B(n1067), .Z(n1076) );
  AND U1173 ( .A(n1078), .B(n1068), .Z(n1069) );
  XOR U1174 ( .A(n1074), .B(n1079), .Z(n1068) );
  XOR U1175 ( .A(n1080), .B(n1077), .Z(n1079) );
  NAND U1176 ( .A(n1066), .B(n1070), .Z(n1077) );
  XOR U1177 ( .A(n1059), .B(n1078), .Z(n1070) );
  XOR U1178 ( .A(n1062), .B(n1067), .Z(n1066) );
  XNOR U1179 ( .A(n1081), .B(n1082), .Z(n1067) );
  XOR U1180 ( .A(n1083), .B(n1084), .Z(n1082) );
  XNOR U1181 ( .A(n1085), .B(n1086), .Z(n1081) );
  ANDN U1182 ( .B(n1009), .A(n1049), .Z(n1085) );
  AND U1183 ( .A(n1059), .B(n1062), .Z(n1080) );
  XNOR U1184 ( .A(n1059), .B(n1062), .Z(n1074) );
  XNOR U1185 ( .A(n1087), .B(n1088), .Z(n1062) );
  XOR U1186 ( .A(n1089), .B(n1090), .Z(n1088) );
  XOR U1187 ( .A(n1083), .B(n1091), .Z(n1087) );
  XNOR U1188 ( .A(n1092), .B(n1086), .Z(n1091) );
  OR U1189 ( .A(n1008), .B(n1048), .Z(n1086) );
  XOR U1190 ( .A(n1049), .B(n1039), .Z(n1048) );
  XOR U1191 ( .A(n1093), .B(n997), .Z(n1008) );
  AND U1192 ( .A(n997), .B(n1039), .Z(n1092) );
  XNOR U1193 ( .A(n1094), .B(n1095), .Z(n1059) );
  XOR U1194 ( .A(n1096), .B(n1097), .Z(n1095) );
  XNOR U1195 ( .A(n1018), .B(n1083), .Z(n1097) );
  XNOR U1196 ( .A(n1049), .B(n1009), .Z(n1083) );
  XOR U1197 ( .A(n993), .B(n1098), .Z(n1094) );
  XNOR U1198 ( .A(n1099), .B(n1100), .Z(n1098) );
  AND U1199 ( .A(n1027), .B(n1045), .Z(n1099) );
  IV U1200 ( .A(n1073), .Z(n1078) );
  XOR U1201 ( .A(n1101), .B(n1102), .Z(n1073) );
  XNOR U1202 ( .A(n1084), .B(n1103), .Z(n1102) );
  XNOR U1203 ( .A(n1027), .B(n1090), .Z(n1103) );
  XOR U1204 ( .A(n1096), .B(n1104), .Z(n1084) );
  XNOR U1205 ( .A(n1105), .B(n1106), .Z(n1104) );
  NAND U1206 ( .A(n1023), .B(n1053), .Z(n1106) );
  IV U1207 ( .A(n1089), .Z(n1096) );
  XOR U1208 ( .A(n1107), .B(n1105), .Z(n1089) );
  NANDN U1209 ( .A(n1055), .B(n1032), .Z(n1105) );
  XOR U1210 ( .A(n1027), .B(n997), .Z(n1023) );
  XOR U1211 ( .A(n1108), .B(n1109), .Z(n997) );
  XOR U1212 ( .A(n1110), .B(n1111), .Z(n1109) );
  XOR U1213 ( .A(n1063), .B(n1053), .Z(n1055) );
  ANDN U1214 ( .B(n1034), .A(n1063), .Z(n1107) );
  XNOR U1215 ( .A(n1112), .B(n1049), .Z(n1063) );
  XNOR U1216 ( .A(n1113), .B(n1114), .Z(n1049) );
  XOR U1217 ( .A(n1115), .B(n1110), .Z(n1113) );
  XOR U1218 ( .A(n1045), .B(n1116), .Z(n1101) );
  XNOR U1219 ( .A(n1117), .B(n1100), .Z(n1116) );
  OR U1220 ( .A(n1029), .B(n1043), .Z(n1100) );
  XNOR U1221 ( .A(n993), .B(n1045), .Z(n1043) );
  XNOR U1222 ( .A(n1018), .B(n1027), .Z(n1029) );
  XOR U1223 ( .A(n1093), .B(n1118), .Z(n1027) );
  XOR U1224 ( .A(state[106]), .B(key[106]), .Z(n1114) );
  IV U1225 ( .A(n1009), .Z(n1093) );
  XOR U1226 ( .A(n1108), .B(n1119), .Z(n1009) );
  XNOR U1227 ( .A(n1110), .B(n1120), .Z(n1119) );
  AND U1228 ( .A(n993), .B(n1018), .Z(n1117) );
  XOR U1229 ( .A(n1108), .B(n1121), .Z(n1018) );
  XNOR U1230 ( .A(n1110), .B(n1122), .Z(n1121) );
  XOR U1231 ( .A(n1112), .B(n1123), .Z(n1110) );
  XNOR U1232 ( .A(state[110]), .B(key[110]), .Z(n1123) );
  XNOR U1233 ( .A(state[109]), .B(key[109]), .Z(n1108) );
  XNOR U1234 ( .A(n1124), .B(n1125), .Z(n1045) );
  XNOR U1235 ( .A(n1122), .B(n1120), .Z(n1125) );
  XOR U1236 ( .A(state[111]), .B(key[111]), .Z(n1120) );
  XOR U1237 ( .A(state[108]), .B(key[108]), .Z(n1122) );
  XOR U1238 ( .A(n993), .B(n1115), .Z(n1124) );
  XOR U1239 ( .A(n1111), .B(n1126), .Z(n1115) );
  XNOR U1240 ( .A(state[107]), .B(key[107]), .Z(n1126) );
  XNOR U1241 ( .A(state[105]), .B(key[105]), .Z(n1111) );
  IV U1242 ( .A(n1112), .Z(n993) );
  XNOR U1243 ( .A(state[104]), .B(key[104]), .Z(n1112) );
  XOR U1244 ( .A(n1127), .B(n1128), .Z(out[3]) );
  XOR U1245 ( .A(n1129), .B(n501), .Z(n1128) );
  XNOR U1246 ( .A(n1130), .B(n1131), .Z(n501) );
  XNOR U1247 ( .A(n1132), .B(n690), .Z(n1131) );
  NOR U1248 ( .A(n1133), .B(n1134), .Z(n690) );
  ANDN U1249 ( .B(n1135), .A(n1136), .Z(n1132) );
  XNOR U1250 ( .A(n1137), .B(n1138), .Z(n1127) );
  XNOR U1251 ( .A(key[3]), .B(n332), .Z(n1138) );
  XOR U1252 ( .A(n1139), .B(n1140), .Z(out[39]) );
  XOR U1253 ( .A(n1141), .B(n1142), .Z(n1139) );
  XOR U1254 ( .A(key[39]), .B(n1143), .Z(n1142) );
  XNOR U1255 ( .A(n1144), .B(n1145), .Z(out[38]) );
  XNOR U1256 ( .A(key[38]), .B(n1146), .Z(n1145) );
  XOR U1257 ( .A(n1147), .B(n1148), .Z(out[37]) );
  XNOR U1258 ( .A(n1149), .B(n1150), .Z(n1148) );
  XOR U1259 ( .A(n1141), .B(n1151), .Z(n1150) );
  XOR U1260 ( .A(n1152), .B(n1153), .Z(n1141) );
  XNOR U1261 ( .A(n1154), .B(n1155), .Z(n1153) );
  NANDN U1262 ( .A(n1156), .B(n1157), .Z(n1155) );
  XOR U1263 ( .A(n1158), .B(n1159), .Z(n1147) );
  XOR U1264 ( .A(key[37]), .B(n1160), .Z(n1159) );
  ANDN U1265 ( .B(n1161), .A(n1162), .Z(n1158) );
  XNOR U1266 ( .A(n1163), .B(n1164), .Z(out[36]) );
  XOR U1267 ( .A(key[36]), .B(n1149), .Z(n1164) );
  XOR U1268 ( .A(n1165), .B(n1166), .Z(out[35]) );
  XOR U1269 ( .A(n1167), .B(n1144), .Z(n1166) );
  XNOR U1270 ( .A(n1168), .B(n1169), .Z(n1144) );
  XNOR U1271 ( .A(n1170), .B(n1160), .Z(n1169) );
  NOR U1272 ( .A(n1171), .B(n1172), .Z(n1160) );
  ANDN U1273 ( .B(n1173), .A(n1174), .Z(n1170) );
  XNOR U1274 ( .A(n1175), .B(n1176), .Z(n1165) );
  XNOR U1275 ( .A(key[35]), .B(n1177), .Z(n1176) );
  XOR U1276 ( .A(key[34]), .B(n1163), .Z(out[34]) );
  XOR U1277 ( .A(n1143), .B(n1178), .Z(n1163) );
  XOR U1278 ( .A(n1179), .B(n1140), .Z(out[33]) );
  XOR U1279 ( .A(n1168), .B(n1180), .Z(n1167) );
  XNOR U1280 ( .A(n1181), .B(n1182), .Z(n1180) );
  NANDN U1281 ( .A(n1156), .B(n1183), .Z(n1182) );
  XNOR U1282 ( .A(n1151), .B(n1184), .Z(n1168) );
  XNOR U1283 ( .A(n1185), .B(n1186), .Z(n1184) );
  NANDN U1284 ( .A(n1187), .B(n1188), .Z(n1186) );
  XOR U1285 ( .A(n1178), .B(n1175), .Z(n1146) );
  XNOR U1286 ( .A(n1151), .B(n1189), .Z(n1175) );
  XNOR U1287 ( .A(n1181), .B(n1190), .Z(n1189) );
  NAND U1288 ( .A(n1191), .B(n1192), .Z(n1190) );
  OR U1289 ( .A(n1193), .B(n1194), .Z(n1181) );
  XOR U1290 ( .A(n1195), .B(n1185), .Z(n1151) );
  NANDN U1291 ( .A(n1196), .B(n1197), .Z(n1185) );
  AND U1292 ( .A(n1198), .B(n1199), .Z(n1195) );
  XOR U1293 ( .A(key[33]), .B(n1143), .Z(n1179) );
  IV U1294 ( .A(n1177), .Z(n1143) );
  XNOR U1295 ( .A(n1200), .B(n1201), .Z(n1177) );
  XNOR U1296 ( .A(n1202), .B(n1203), .Z(n1201) );
  OR U1297 ( .A(n1204), .B(n1162), .Z(n1203) );
  XNOR U1298 ( .A(n1149), .B(n1205), .Z(out[32]) );
  XOR U1299 ( .A(key[32]), .B(n1178), .Z(n1205) );
  XNOR U1300 ( .A(n1200), .B(n1206), .Z(n1178) );
  XOR U1301 ( .A(n1207), .B(n1154), .Z(n1206) );
  OR U1302 ( .A(n1208), .B(n1193), .Z(n1154) );
  XNOR U1303 ( .A(n1156), .B(n1209), .Z(n1193) );
  AND U1304 ( .A(n1210), .B(n1191), .Z(n1207) );
  XNOR U1305 ( .A(n1152), .B(n1211), .Z(n1149) );
  XOR U1306 ( .A(n1212), .B(n1202), .Z(n1211) );
  OR U1307 ( .A(n1213), .B(n1171), .Z(n1202) );
  XNOR U1308 ( .A(n1174), .B(n1162), .Z(n1171) );
  NOR U1309 ( .A(n1214), .B(n1174), .Z(n1212) );
  XNOR U1310 ( .A(n1200), .B(n1215), .Z(n1152) );
  XNOR U1311 ( .A(n1216), .B(n1217), .Z(n1215) );
  NANDN U1312 ( .A(n1187), .B(n1218), .Z(n1217) );
  XOR U1313 ( .A(n1219), .B(n1216), .Z(n1200) );
  OR U1314 ( .A(n1196), .B(n1220), .Z(n1216) );
  XOR U1315 ( .A(n1198), .B(n1187), .Z(n1196) );
  XNOR U1316 ( .A(n1209), .B(n1162), .Z(n1187) );
  XOR U1317 ( .A(n1221), .B(n1222), .Z(n1162) );
  NANDN U1318 ( .A(n1223), .B(n1224), .Z(n1222) );
  IV U1319 ( .A(n1191), .Z(n1209) );
  XOR U1320 ( .A(n1225), .B(n1226), .Z(n1191) );
  NANDN U1321 ( .A(n1223), .B(n1227), .Z(n1226) );
  ANDN U1322 ( .B(n1198), .A(n1228), .Z(n1219) );
  XOR U1323 ( .A(n1174), .B(n1156), .Z(n1198) );
  XOR U1324 ( .A(n1229), .B(n1225), .Z(n1156) );
  NANDN U1325 ( .A(n1230), .B(n1231), .Z(n1225) );
  AND U1326 ( .A(n1232), .B(n1233), .Z(n1229) );
  ANDN U1327 ( .B(n1235), .A(n1230), .Z(n1221) );
  XOR U1328 ( .A(n1236), .B(n1237), .Z(n1223) );
  XNOR U1329 ( .A(n1239), .B(n1240), .Z(n1236) );
  XNOR U1330 ( .A(n1241), .B(n1242), .Z(n1240) );
  AND U1331 ( .A(n1243), .B(n1232), .Z(n1241) );
  AND U1332 ( .A(n1243), .B(n1233), .Z(n1234) );
  XOR U1333 ( .A(n1239), .B(n1244), .Z(n1233) );
  XOR U1334 ( .A(n1245), .B(n1242), .Z(n1244) );
  NAND U1335 ( .A(n1231), .B(n1235), .Z(n1242) );
  XOR U1336 ( .A(n1224), .B(n1243), .Z(n1235) );
  XOR U1337 ( .A(n1227), .B(n1232), .Z(n1231) );
  XNOR U1338 ( .A(n1246), .B(n1247), .Z(n1232) );
  XOR U1339 ( .A(n1248), .B(n1249), .Z(n1247) );
  XNOR U1340 ( .A(n1250), .B(n1251), .Z(n1246) );
  ANDN U1341 ( .B(n1173), .A(n1214), .Z(n1250) );
  AND U1342 ( .A(n1224), .B(n1227), .Z(n1245) );
  XNOR U1343 ( .A(n1224), .B(n1227), .Z(n1239) );
  XNOR U1344 ( .A(n1252), .B(n1253), .Z(n1227) );
  XOR U1345 ( .A(n1254), .B(n1255), .Z(n1253) );
  XOR U1346 ( .A(n1248), .B(n1256), .Z(n1252) );
  XNOR U1347 ( .A(n1257), .B(n1251), .Z(n1256) );
  OR U1348 ( .A(n1172), .B(n1213), .Z(n1251) );
  XNOR U1349 ( .A(n1214), .B(n1204), .Z(n1213) );
  XOR U1350 ( .A(n1258), .B(n1161), .Z(n1172) );
  ANDN U1351 ( .B(n1161), .A(n1204), .Z(n1257) );
  XNOR U1352 ( .A(n1259), .B(n1260), .Z(n1224) );
  XOR U1353 ( .A(n1261), .B(n1262), .Z(n1260) );
  XNOR U1354 ( .A(n1183), .B(n1248), .Z(n1262) );
  XNOR U1355 ( .A(n1214), .B(n1173), .Z(n1248) );
  XOR U1356 ( .A(n1157), .B(n1263), .Z(n1259) );
  XNOR U1357 ( .A(n1264), .B(n1265), .Z(n1263) );
  AND U1358 ( .A(n1192), .B(n1210), .Z(n1264) );
  IV U1359 ( .A(n1238), .Z(n1243) );
  XOR U1360 ( .A(n1266), .B(n1267), .Z(n1238) );
  XNOR U1361 ( .A(n1249), .B(n1268), .Z(n1267) );
  XNOR U1362 ( .A(n1192), .B(n1255), .Z(n1268) );
  XNOR U1363 ( .A(n1204), .B(n1161), .Z(n1255) );
  XOR U1364 ( .A(n1261), .B(n1269), .Z(n1249) );
  XNOR U1365 ( .A(n1270), .B(n1271), .Z(n1269) );
  NAND U1366 ( .A(n1188), .B(n1218), .Z(n1271) );
  IV U1367 ( .A(n1254), .Z(n1261) );
  XOR U1368 ( .A(n1272), .B(n1270), .Z(n1254) );
  NANDN U1369 ( .A(n1220), .B(n1197), .Z(n1270) );
  XOR U1370 ( .A(n1192), .B(n1161), .Z(n1188) );
  XOR U1371 ( .A(n1273), .B(n1274), .Z(n1161) );
  XOR U1372 ( .A(n1275), .B(n1276), .Z(n1274) );
  XOR U1373 ( .A(n1228), .B(n1218), .Z(n1220) );
  XOR U1374 ( .A(n1275), .B(n1273), .Z(n1204) );
  ANDN U1375 ( .B(n1199), .A(n1228), .Z(n1272) );
  XNOR U1376 ( .A(n1277), .B(n1214), .Z(n1228) );
  XOR U1377 ( .A(n1278), .B(n1279), .Z(n1214) );
  XNOR U1378 ( .A(n1280), .B(n1275), .Z(n1278) );
  XOR U1379 ( .A(n1210), .B(n1281), .Z(n1266) );
  XNOR U1380 ( .A(n1282), .B(n1265), .Z(n1281) );
  OR U1381 ( .A(n1194), .B(n1208), .Z(n1265) );
  XNOR U1382 ( .A(n1157), .B(n1210), .Z(n1208) );
  XNOR U1383 ( .A(n1183), .B(n1192), .Z(n1194) );
  XOR U1384 ( .A(n1258), .B(n1283), .Z(n1192) );
  XNOR U1385 ( .A(n1276), .B(n1279), .Z(n1283) );
  XNOR U1386 ( .A(state[66]), .B(key[66]), .Z(n1279) );
  IV U1387 ( .A(n1173), .Z(n1258) );
  XOR U1388 ( .A(n1273), .B(n1284), .Z(n1173) );
  XOR U1389 ( .A(n1275), .B(n1285), .Z(n1284) );
  AND U1390 ( .A(n1157), .B(n1183), .Z(n1282) );
  XOR U1391 ( .A(n1273), .B(n1286), .Z(n1183) );
  XOR U1392 ( .A(n1275), .B(n1287), .Z(n1286) );
  XOR U1393 ( .A(n1277), .B(n1288), .Z(n1275) );
  XNOR U1394 ( .A(state[70]), .B(key[70]), .Z(n1288) );
  XNOR U1395 ( .A(state[69]), .B(key[69]), .Z(n1273) );
  XNOR U1396 ( .A(n1289), .B(n1290), .Z(n1210) );
  XNOR U1397 ( .A(n1287), .B(n1285), .Z(n1290) );
  XNOR U1398 ( .A(state[71]), .B(key[71]), .Z(n1285) );
  XNOR U1399 ( .A(state[68]), .B(key[68]), .Z(n1287) );
  XNOR U1400 ( .A(n1157), .B(n1280), .Z(n1289) );
  XNOR U1401 ( .A(n1276), .B(n1291), .Z(n1280) );
  XNOR U1402 ( .A(state[67]), .B(key[67]), .Z(n1291) );
  XNOR U1403 ( .A(state[65]), .B(key[65]), .Z(n1276) );
  IV U1404 ( .A(n1277), .Z(n1157) );
  XNOR U1405 ( .A(state[64]), .B(key[64]), .Z(n1277) );
  XOR U1406 ( .A(n1292), .B(n1293), .Z(out[31]) );
  XOR U1407 ( .A(n1294), .B(n1295), .Z(n1292) );
  XOR U1408 ( .A(key[31]), .B(n1296), .Z(n1295) );
  XNOR U1409 ( .A(n1297), .B(n1298), .Z(out[30]) );
  XNOR U1410 ( .A(key[30]), .B(n1299), .Z(n1298) );
  XOR U1411 ( .A(key[2]), .B(n860), .Z(out[2]) );
  XOR U1412 ( .A(n1300), .B(n1301), .Z(n860) );
  XOR U1413 ( .A(n1302), .B(n1303), .Z(out[29]) );
  XNOR U1414 ( .A(n1304), .B(n1305), .Z(n1303) );
  XOR U1415 ( .A(n1294), .B(n1306), .Z(n1305) );
  XOR U1416 ( .A(n1307), .B(n1308), .Z(n1294) );
  XNOR U1417 ( .A(n1309), .B(n1310), .Z(n1308) );
  NANDN U1418 ( .A(n1311), .B(n1312), .Z(n1310) );
  XOR U1419 ( .A(n1313), .B(n1314), .Z(n1302) );
  XOR U1420 ( .A(key[29]), .B(n1315), .Z(n1314) );
  ANDN U1421 ( .B(n1316), .A(n1317), .Z(n1313) );
  XNOR U1422 ( .A(n1318), .B(n1319), .Z(out[28]) );
  XOR U1423 ( .A(key[28]), .B(n1304), .Z(n1319) );
  XOR U1424 ( .A(n1320), .B(n1321), .Z(out[27]) );
  XOR U1425 ( .A(n1322), .B(n1297), .Z(n1321) );
  XNOR U1426 ( .A(n1323), .B(n1324), .Z(n1297) );
  XNOR U1427 ( .A(n1325), .B(n1315), .Z(n1324) );
  NOR U1428 ( .A(n1326), .B(n1327), .Z(n1315) );
  ANDN U1429 ( .B(n1328), .A(n1329), .Z(n1325) );
  XNOR U1430 ( .A(n1330), .B(n1331), .Z(n1320) );
  XNOR U1431 ( .A(key[27]), .B(n1332), .Z(n1331) );
  XOR U1432 ( .A(key[26]), .B(n1318), .Z(out[26]) );
  XOR U1433 ( .A(n1296), .B(n1333), .Z(n1318) );
  XOR U1434 ( .A(n1334), .B(n1293), .Z(out[25]) );
  XOR U1435 ( .A(n1323), .B(n1335), .Z(n1322) );
  XNOR U1436 ( .A(n1336), .B(n1337), .Z(n1335) );
  NANDN U1437 ( .A(n1311), .B(n1338), .Z(n1337) );
  XNOR U1438 ( .A(n1306), .B(n1339), .Z(n1323) );
  XNOR U1439 ( .A(n1340), .B(n1341), .Z(n1339) );
  NANDN U1440 ( .A(n1342), .B(n1343), .Z(n1341) );
  XOR U1441 ( .A(n1333), .B(n1330), .Z(n1299) );
  XNOR U1442 ( .A(n1306), .B(n1344), .Z(n1330) );
  XNOR U1443 ( .A(n1336), .B(n1345), .Z(n1344) );
  NAND U1444 ( .A(n1346), .B(n1347), .Z(n1345) );
  OR U1445 ( .A(n1348), .B(n1349), .Z(n1336) );
  XOR U1446 ( .A(n1350), .B(n1340), .Z(n1306) );
  NANDN U1447 ( .A(n1351), .B(n1352), .Z(n1340) );
  AND U1448 ( .A(n1353), .B(n1354), .Z(n1350) );
  XOR U1449 ( .A(key[25]), .B(n1296), .Z(n1334) );
  IV U1450 ( .A(n1332), .Z(n1296) );
  XNOR U1451 ( .A(n1355), .B(n1356), .Z(n1332) );
  XNOR U1452 ( .A(n1357), .B(n1358), .Z(n1356) );
  NANDN U1453 ( .A(n1317), .B(n1359), .Z(n1358) );
  XNOR U1454 ( .A(n1304), .B(n1360), .Z(out[24]) );
  XOR U1455 ( .A(key[24]), .B(n1333), .Z(n1360) );
  XNOR U1456 ( .A(n1355), .B(n1361), .Z(n1333) );
  XOR U1457 ( .A(n1362), .B(n1309), .Z(n1361) );
  OR U1458 ( .A(n1363), .B(n1348), .Z(n1309) );
  XNOR U1459 ( .A(n1311), .B(n1364), .Z(n1348) );
  AND U1460 ( .A(n1365), .B(n1346), .Z(n1362) );
  XNOR U1461 ( .A(n1307), .B(n1366), .Z(n1304) );
  XOR U1462 ( .A(n1367), .B(n1357), .Z(n1366) );
  OR U1463 ( .A(n1368), .B(n1326), .Z(n1357) );
  XNOR U1464 ( .A(n1329), .B(n1317), .Z(n1326) );
  NOR U1465 ( .A(n1369), .B(n1329), .Z(n1367) );
  XNOR U1466 ( .A(n1355), .B(n1370), .Z(n1307) );
  XNOR U1467 ( .A(n1371), .B(n1372), .Z(n1370) );
  NANDN U1468 ( .A(n1342), .B(n1373), .Z(n1372) );
  XOR U1469 ( .A(n1374), .B(n1371), .Z(n1355) );
  OR U1470 ( .A(n1351), .B(n1375), .Z(n1371) );
  XOR U1471 ( .A(n1353), .B(n1342), .Z(n1351) );
  XNOR U1472 ( .A(n1364), .B(n1317), .Z(n1342) );
  XOR U1473 ( .A(n1376), .B(n1377), .Z(n1317) );
  NANDN U1474 ( .A(n1378), .B(n1379), .Z(n1377) );
  IV U1475 ( .A(n1346), .Z(n1364) );
  XOR U1476 ( .A(n1380), .B(n1381), .Z(n1346) );
  NANDN U1477 ( .A(n1378), .B(n1382), .Z(n1381) );
  ANDN U1478 ( .B(n1353), .A(n1383), .Z(n1374) );
  XOR U1479 ( .A(n1329), .B(n1311), .Z(n1353) );
  XOR U1480 ( .A(n1384), .B(n1380), .Z(n1311) );
  NANDN U1481 ( .A(n1385), .B(n1386), .Z(n1380) );
  AND U1482 ( .A(n1387), .B(n1388), .Z(n1384) );
  ANDN U1483 ( .B(n1390), .A(n1385), .Z(n1376) );
  XOR U1484 ( .A(n1391), .B(n1392), .Z(n1378) );
  XNOR U1485 ( .A(n1394), .B(n1395), .Z(n1391) );
  XNOR U1486 ( .A(n1396), .B(n1397), .Z(n1395) );
  AND U1487 ( .A(n1398), .B(n1387), .Z(n1396) );
  AND U1488 ( .A(n1398), .B(n1388), .Z(n1389) );
  XOR U1489 ( .A(n1394), .B(n1399), .Z(n1388) );
  XOR U1490 ( .A(n1400), .B(n1397), .Z(n1399) );
  NAND U1491 ( .A(n1386), .B(n1390), .Z(n1397) );
  XOR U1492 ( .A(n1379), .B(n1398), .Z(n1390) );
  XOR U1493 ( .A(n1382), .B(n1387), .Z(n1386) );
  XNOR U1494 ( .A(n1401), .B(n1402), .Z(n1387) );
  XOR U1495 ( .A(n1403), .B(n1404), .Z(n1402) );
  XNOR U1496 ( .A(n1405), .B(n1406), .Z(n1401) );
  ANDN U1497 ( .B(n1328), .A(n1369), .Z(n1405) );
  AND U1498 ( .A(n1379), .B(n1382), .Z(n1400) );
  XNOR U1499 ( .A(n1379), .B(n1382), .Z(n1394) );
  XNOR U1500 ( .A(n1407), .B(n1408), .Z(n1382) );
  XOR U1501 ( .A(n1409), .B(n1410), .Z(n1408) );
  XOR U1502 ( .A(n1403), .B(n1411), .Z(n1407) );
  XNOR U1503 ( .A(n1412), .B(n1406), .Z(n1411) );
  OR U1504 ( .A(n1327), .B(n1368), .Z(n1406) );
  XOR U1505 ( .A(n1369), .B(n1359), .Z(n1368) );
  XOR U1506 ( .A(n1413), .B(n1316), .Z(n1327) );
  AND U1507 ( .A(n1316), .B(n1359), .Z(n1412) );
  XNOR U1508 ( .A(n1414), .B(n1415), .Z(n1379) );
  XOR U1509 ( .A(n1416), .B(n1417), .Z(n1415) );
  XNOR U1510 ( .A(n1338), .B(n1403), .Z(n1417) );
  XNOR U1511 ( .A(n1369), .B(n1328), .Z(n1403) );
  XOR U1512 ( .A(n1312), .B(n1418), .Z(n1414) );
  XNOR U1513 ( .A(n1419), .B(n1420), .Z(n1418) );
  AND U1514 ( .A(n1347), .B(n1365), .Z(n1419) );
  IV U1515 ( .A(n1393), .Z(n1398) );
  XOR U1516 ( .A(n1421), .B(n1422), .Z(n1393) );
  XNOR U1517 ( .A(n1404), .B(n1423), .Z(n1422) );
  XNOR U1518 ( .A(n1347), .B(n1410), .Z(n1423) );
  XOR U1519 ( .A(n1416), .B(n1424), .Z(n1404) );
  XNOR U1520 ( .A(n1425), .B(n1426), .Z(n1424) );
  NAND U1521 ( .A(n1343), .B(n1373), .Z(n1426) );
  IV U1522 ( .A(n1409), .Z(n1416) );
  XOR U1523 ( .A(n1427), .B(n1425), .Z(n1409) );
  NANDN U1524 ( .A(n1375), .B(n1352), .Z(n1425) );
  XOR U1525 ( .A(n1347), .B(n1316), .Z(n1343) );
  XOR U1526 ( .A(n1428), .B(n1429), .Z(n1316) );
  XOR U1527 ( .A(n1430), .B(n1431), .Z(n1429) );
  XOR U1528 ( .A(n1383), .B(n1373), .Z(n1375) );
  ANDN U1529 ( .B(n1354), .A(n1383), .Z(n1427) );
  XNOR U1530 ( .A(n1432), .B(n1369), .Z(n1383) );
  XNOR U1531 ( .A(n1433), .B(n1434), .Z(n1369) );
  XOR U1532 ( .A(n1435), .B(n1430), .Z(n1433) );
  XOR U1533 ( .A(n1365), .B(n1436), .Z(n1421) );
  XNOR U1534 ( .A(n1437), .B(n1420), .Z(n1436) );
  OR U1535 ( .A(n1349), .B(n1363), .Z(n1420) );
  XNOR U1536 ( .A(n1312), .B(n1365), .Z(n1363) );
  XNOR U1537 ( .A(n1338), .B(n1347), .Z(n1349) );
  XOR U1538 ( .A(n1413), .B(n1438), .Z(n1347) );
  XOR U1539 ( .A(state[26]), .B(key[26]), .Z(n1434) );
  IV U1540 ( .A(n1328), .Z(n1413) );
  XOR U1541 ( .A(n1428), .B(n1439), .Z(n1328) );
  XNOR U1542 ( .A(n1430), .B(n1440), .Z(n1439) );
  AND U1543 ( .A(n1312), .B(n1338), .Z(n1437) );
  XOR U1544 ( .A(n1428), .B(n1441), .Z(n1338) );
  XNOR U1545 ( .A(n1430), .B(n1442), .Z(n1441) );
  XOR U1546 ( .A(n1432), .B(n1443), .Z(n1430) );
  XNOR U1547 ( .A(state[30]), .B(key[30]), .Z(n1443) );
  XNOR U1548 ( .A(state[29]), .B(key[29]), .Z(n1428) );
  XNOR U1549 ( .A(n1444), .B(n1445), .Z(n1365) );
  XNOR U1550 ( .A(n1442), .B(n1440), .Z(n1445) );
  XOR U1551 ( .A(state[31]), .B(key[31]), .Z(n1440) );
  XOR U1552 ( .A(state[28]), .B(key[28]), .Z(n1442) );
  XOR U1553 ( .A(n1312), .B(n1435), .Z(n1444) );
  XOR U1554 ( .A(n1431), .B(n1446), .Z(n1435) );
  XNOR U1555 ( .A(state[27]), .B(key[27]), .Z(n1446) );
  XNOR U1556 ( .A(state[25]), .B(key[25]), .Z(n1431) );
  IV U1557 ( .A(n1432), .Z(n1312) );
  XNOR U1558 ( .A(state[24]), .B(key[24]), .Z(n1432) );
  XOR U1559 ( .A(n1447), .B(n1448), .Z(out[23]) );
  XOR U1560 ( .A(n1449), .B(n1450), .Z(n1447) );
  XOR U1561 ( .A(key[23]), .B(n1451), .Z(n1450) );
  XNOR U1562 ( .A(n1452), .B(n1453), .Z(out[22]) );
  XNOR U1563 ( .A(key[22]), .B(n1454), .Z(n1453) );
  XOR U1564 ( .A(n1455), .B(n1456), .Z(out[21]) );
  XNOR U1565 ( .A(n1457), .B(n1458), .Z(n1456) );
  XOR U1566 ( .A(n1449), .B(n1459), .Z(n1458) );
  XOR U1567 ( .A(n1460), .B(n1461), .Z(n1449) );
  XNOR U1568 ( .A(n1462), .B(n1463), .Z(n1461) );
  NANDN U1569 ( .A(n1464), .B(n1465), .Z(n1463) );
  XOR U1570 ( .A(n1466), .B(n1467), .Z(n1455) );
  XOR U1571 ( .A(key[21]), .B(n1468), .Z(n1467) );
  ANDN U1572 ( .B(n1469), .A(n1470), .Z(n1466) );
  XNOR U1573 ( .A(n1471), .B(n1472), .Z(out[20]) );
  XOR U1574 ( .A(key[20]), .B(n1457), .Z(n1472) );
  XOR U1575 ( .A(n1473), .B(n329), .Z(out[1]) );
  XOR U1576 ( .A(n1130), .B(n1474), .Z(n1129) );
  XNOR U1577 ( .A(n1475), .B(n1476), .Z(n1474) );
  NANDN U1578 ( .A(n686), .B(n1477), .Z(n1476) );
  XNOR U1579 ( .A(n681), .B(n1478), .Z(n1130) );
  XNOR U1580 ( .A(n1479), .B(n1480), .Z(n1478) );
  NANDN U1581 ( .A(n1481), .B(n1482), .Z(n1480) );
  XOR U1582 ( .A(n1301), .B(n1137), .Z(n503) );
  XNOR U1583 ( .A(n681), .B(n1483), .Z(n1137) );
  XNOR U1584 ( .A(n1475), .B(n1484), .Z(n1483) );
  NAND U1585 ( .A(n1485), .B(n1486), .Z(n1484) );
  OR U1586 ( .A(n1487), .B(n1488), .Z(n1475) );
  XOR U1587 ( .A(n1489), .B(n1479), .Z(n681) );
  NANDN U1588 ( .A(n1490), .B(n1491), .Z(n1479) );
  AND U1589 ( .A(n1492), .B(n1493), .Z(n1489) );
  XOR U1590 ( .A(key[1]), .B(n1300), .Z(n1473) );
  IV U1591 ( .A(n332), .Z(n1300) );
  XNOR U1592 ( .A(n1494), .B(n1495), .Z(n332) );
  XNOR U1593 ( .A(n1496), .B(n1497), .Z(n1495) );
  NANDN U1594 ( .A(n692), .B(n1498), .Z(n1497) );
  XOR U1595 ( .A(n1499), .B(n1500), .Z(out[19]) );
  XOR U1596 ( .A(n1501), .B(n1452), .Z(n1500) );
  XNOR U1597 ( .A(n1502), .B(n1503), .Z(n1452) );
  XNOR U1598 ( .A(n1504), .B(n1468), .Z(n1503) );
  NOR U1599 ( .A(n1505), .B(n1506), .Z(n1468) );
  ANDN U1600 ( .B(n1507), .A(n1508), .Z(n1504) );
  XNOR U1601 ( .A(n1509), .B(n1510), .Z(n1499) );
  XNOR U1602 ( .A(key[19]), .B(n1511), .Z(n1510) );
  XOR U1603 ( .A(key[18]), .B(n1471), .Z(out[18]) );
  XOR U1604 ( .A(n1451), .B(n1512), .Z(n1471) );
  XOR U1605 ( .A(n1513), .B(n1448), .Z(out[17]) );
  XOR U1606 ( .A(n1502), .B(n1514), .Z(n1501) );
  XNOR U1607 ( .A(n1515), .B(n1516), .Z(n1514) );
  NANDN U1608 ( .A(n1464), .B(n1517), .Z(n1516) );
  XNOR U1609 ( .A(n1459), .B(n1518), .Z(n1502) );
  XNOR U1610 ( .A(n1519), .B(n1520), .Z(n1518) );
  NANDN U1611 ( .A(n1521), .B(n1522), .Z(n1520) );
  XOR U1612 ( .A(n1512), .B(n1509), .Z(n1454) );
  XNOR U1613 ( .A(n1459), .B(n1523), .Z(n1509) );
  XNOR U1614 ( .A(n1515), .B(n1524), .Z(n1523) );
  NAND U1615 ( .A(n1525), .B(n1526), .Z(n1524) );
  OR U1616 ( .A(n1527), .B(n1528), .Z(n1515) );
  XOR U1617 ( .A(n1529), .B(n1519), .Z(n1459) );
  NANDN U1618 ( .A(n1530), .B(n1531), .Z(n1519) );
  AND U1619 ( .A(n1532), .B(n1533), .Z(n1529) );
  XOR U1620 ( .A(key[17]), .B(n1451), .Z(n1513) );
  IV U1621 ( .A(n1511), .Z(n1451) );
  XNOR U1622 ( .A(n1534), .B(n1535), .Z(n1511) );
  XNOR U1623 ( .A(n1536), .B(n1537), .Z(n1535) );
  NANDN U1624 ( .A(n1470), .B(n1538), .Z(n1537) );
  XNOR U1625 ( .A(n1457), .B(n1539), .Z(out[16]) );
  XOR U1626 ( .A(key[16]), .B(n1512), .Z(n1539) );
  XNOR U1627 ( .A(n1534), .B(n1540), .Z(n1512) );
  XOR U1628 ( .A(n1541), .B(n1462), .Z(n1540) );
  OR U1629 ( .A(n1542), .B(n1527), .Z(n1462) );
  XNOR U1630 ( .A(n1464), .B(n1543), .Z(n1527) );
  AND U1631 ( .A(n1544), .B(n1525), .Z(n1541) );
  XNOR U1632 ( .A(n1460), .B(n1545), .Z(n1457) );
  XOR U1633 ( .A(n1546), .B(n1536), .Z(n1545) );
  OR U1634 ( .A(n1547), .B(n1505), .Z(n1536) );
  XNOR U1635 ( .A(n1508), .B(n1470), .Z(n1505) );
  NOR U1636 ( .A(n1548), .B(n1508), .Z(n1546) );
  XNOR U1637 ( .A(n1534), .B(n1549), .Z(n1460) );
  XNOR U1638 ( .A(n1550), .B(n1551), .Z(n1549) );
  NANDN U1639 ( .A(n1521), .B(n1552), .Z(n1551) );
  XOR U1640 ( .A(n1553), .B(n1550), .Z(n1534) );
  OR U1641 ( .A(n1530), .B(n1554), .Z(n1550) );
  XOR U1642 ( .A(n1532), .B(n1521), .Z(n1530) );
  XNOR U1643 ( .A(n1543), .B(n1470), .Z(n1521) );
  XOR U1644 ( .A(n1555), .B(n1556), .Z(n1470) );
  NANDN U1645 ( .A(n1557), .B(n1558), .Z(n1556) );
  IV U1646 ( .A(n1525), .Z(n1543) );
  XOR U1647 ( .A(n1559), .B(n1560), .Z(n1525) );
  NANDN U1648 ( .A(n1557), .B(n1561), .Z(n1560) );
  ANDN U1649 ( .B(n1532), .A(n1562), .Z(n1553) );
  XOR U1650 ( .A(n1508), .B(n1464), .Z(n1532) );
  XOR U1651 ( .A(n1563), .B(n1559), .Z(n1464) );
  NANDN U1652 ( .A(n1564), .B(n1565), .Z(n1559) );
  AND U1653 ( .A(n1566), .B(n1567), .Z(n1563) );
  ANDN U1654 ( .B(n1569), .A(n1564), .Z(n1555) );
  XOR U1655 ( .A(n1570), .B(n1571), .Z(n1557) );
  XNOR U1656 ( .A(n1573), .B(n1574), .Z(n1570) );
  XNOR U1657 ( .A(n1575), .B(n1576), .Z(n1574) );
  AND U1658 ( .A(n1577), .B(n1566), .Z(n1575) );
  AND U1659 ( .A(n1577), .B(n1567), .Z(n1568) );
  XOR U1660 ( .A(n1573), .B(n1578), .Z(n1567) );
  XOR U1661 ( .A(n1579), .B(n1576), .Z(n1578) );
  NAND U1662 ( .A(n1565), .B(n1569), .Z(n1576) );
  XOR U1663 ( .A(n1558), .B(n1577), .Z(n1569) );
  XOR U1664 ( .A(n1561), .B(n1566), .Z(n1565) );
  XNOR U1665 ( .A(n1580), .B(n1581), .Z(n1566) );
  XOR U1666 ( .A(n1582), .B(n1583), .Z(n1581) );
  XNOR U1667 ( .A(n1584), .B(n1585), .Z(n1580) );
  ANDN U1668 ( .B(n1507), .A(n1548), .Z(n1584) );
  AND U1669 ( .A(n1558), .B(n1561), .Z(n1579) );
  XNOR U1670 ( .A(n1558), .B(n1561), .Z(n1573) );
  XNOR U1671 ( .A(n1586), .B(n1587), .Z(n1561) );
  XOR U1672 ( .A(n1588), .B(n1589), .Z(n1587) );
  XOR U1673 ( .A(n1582), .B(n1590), .Z(n1586) );
  XNOR U1674 ( .A(n1591), .B(n1585), .Z(n1590) );
  OR U1675 ( .A(n1506), .B(n1547), .Z(n1585) );
  XOR U1676 ( .A(n1548), .B(n1538), .Z(n1547) );
  XOR U1677 ( .A(n1592), .B(n1469), .Z(n1506) );
  AND U1678 ( .A(n1469), .B(n1538), .Z(n1591) );
  XNOR U1679 ( .A(n1593), .B(n1594), .Z(n1558) );
  XOR U1680 ( .A(n1595), .B(n1596), .Z(n1594) );
  XNOR U1681 ( .A(n1517), .B(n1582), .Z(n1596) );
  XNOR U1682 ( .A(n1548), .B(n1507), .Z(n1582) );
  XOR U1683 ( .A(n1465), .B(n1597), .Z(n1593) );
  XNOR U1684 ( .A(n1598), .B(n1599), .Z(n1597) );
  AND U1685 ( .A(n1526), .B(n1544), .Z(n1598) );
  IV U1686 ( .A(n1572), .Z(n1577) );
  XOR U1687 ( .A(n1600), .B(n1601), .Z(n1572) );
  XNOR U1688 ( .A(n1583), .B(n1602), .Z(n1601) );
  XNOR U1689 ( .A(n1526), .B(n1589), .Z(n1602) );
  XOR U1690 ( .A(n1595), .B(n1603), .Z(n1583) );
  XNOR U1691 ( .A(n1604), .B(n1605), .Z(n1603) );
  NAND U1692 ( .A(n1522), .B(n1552), .Z(n1605) );
  IV U1693 ( .A(n1588), .Z(n1595) );
  XOR U1694 ( .A(n1606), .B(n1604), .Z(n1588) );
  NANDN U1695 ( .A(n1554), .B(n1531), .Z(n1604) );
  XOR U1696 ( .A(n1526), .B(n1469), .Z(n1522) );
  XOR U1697 ( .A(n1607), .B(n1608), .Z(n1469) );
  XOR U1698 ( .A(n1609), .B(n1610), .Z(n1608) );
  XOR U1699 ( .A(n1562), .B(n1552), .Z(n1554) );
  ANDN U1700 ( .B(n1533), .A(n1562), .Z(n1606) );
  XNOR U1701 ( .A(n1611), .B(n1548), .Z(n1562) );
  XNOR U1702 ( .A(n1612), .B(n1613), .Z(n1548) );
  XOR U1703 ( .A(n1614), .B(n1609), .Z(n1612) );
  XOR U1704 ( .A(n1544), .B(n1615), .Z(n1600) );
  XNOR U1705 ( .A(n1616), .B(n1599), .Z(n1615) );
  OR U1706 ( .A(n1528), .B(n1542), .Z(n1599) );
  XNOR U1707 ( .A(n1465), .B(n1544), .Z(n1542) );
  XNOR U1708 ( .A(n1517), .B(n1526), .Z(n1528) );
  XOR U1709 ( .A(n1592), .B(n1617), .Z(n1526) );
  XOR U1710 ( .A(state[114]), .B(key[114]), .Z(n1613) );
  IV U1711 ( .A(n1507), .Z(n1592) );
  XOR U1712 ( .A(n1607), .B(n1618), .Z(n1507) );
  XNOR U1713 ( .A(n1609), .B(n1619), .Z(n1618) );
  AND U1714 ( .A(n1465), .B(n1517), .Z(n1616) );
  XOR U1715 ( .A(n1607), .B(n1620), .Z(n1517) );
  XNOR U1716 ( .A(n1609), .B(n1621), .Z(n1620) );
  XOR U1717 ( .A(n1611), .B(n1622), .Z(n1609) );
  XNOR U1718 ( .A(state[118]), .B(key[118]), .Z(n1622) );
  XNOR U1719 ( .A(state[117]), .B(key[117]), .Z(n1607) );
  XNOR U1720 ( .A(n1623), .B(n1624), .Z(n1544) );
  XNOR U1721 ( .A(n1621), .B(n1619), .Z(n1624) );
  XOR U1722 ( .A(state[119]), .B(key[119]), .Z(n1619) );
  XOR U1723 ( .A(state[116]), .B(key[116]), .Z(n1621) );
  XOR U1724 ( .A(n1465), .B(n1614), .Z(n1623) );
  XOR U1725 ( .A(n1610), .B(n1625), .Z(n1614) );
  XNOR U1726 ( .A(state[115]), .B(key[115]), .Z(n1625) );
  XNOR U1727 ( .A(state[113]), .B(key[113]), .Z(n1610) );
  IV U1728 ( .A(n1611), .Z(n1465) );
  XNOR U1729 ( .A(state[112]), .B(key[112]), .Z(n1611) );
  XOR U1730 ( .A(n1626), .B(n1627), .Z(out[15]) );
  XNOR U1731 ( .A(n4), .B(n1628), .Z(n1627) );
  XNOR U1732 ( .A(n3), .B(n1629), .Z(n1626) );
  XOR U1733 ( .A(key[15]), .B(n5), .Z(n1629) );
  XNOR U1734 ( .A(n1630), .B(n1631), .Z(out[14]) );
  XOR U1735 ( .A(key[14]), .B(n3), .Z(n1631) );
  XOR U1736 ( .A(n1633), .B(n1634), .Z(out[13]) );
  XNOR U1737 ( .A(n1628), .B(n1635), .Z(n1634) );
  XNOR U1738 ( .A(n1636), .B(n60), .Z(n1635) );
  XNOR U1739 ( .A(n1637), .B(n1638), .Z(n1628) );
  XNOR U1740 ( .A(n1639), .B(n1640), .Z(n1638) );
  NANDN U1741 ( .A(n1641), .B(n1642), .Z(n1640) );
  XOR U1742 ( .A(n1643), .B(n1644), .Z(n1633) );
  XOR U1743 ( .A(key[13]), .B(n1645), .Z(n1644) );
  AND U1744 ( .A(n1646), .B(n1647), .Z(n1643) );
  XNOR U1745 ( .A(n1648), .B(n1649), .Z(out[12]) );
  XOR U1746 ( .A(key[12]), .B(n60), .Z(n1649) );
  XNOR U1747 ( .A(n1637), .B(n1650), .Z(n60) );
  XOR U1748 ( .A(n1651), .B(n1652), .Z(n1650) );
  ANDN U1749 ( .B(n1653), .A(n1654), .Z(n1651) );
  XNOR U1750 ( .A(n1655), .B(n1656), .Z(n1637) );
  XNOR U1751 ( .A(n1657), .B(n1658), .Z(n1656) );
  NANDN U1752 ( .A(n1659), .B(n1660), .Z(n1658) );
  XOR U1753 ( .A(n1661), .B(n1662), .Z(out[127]) );
  XOR U1754 ( .A(n1663), .B(n1664), .Z(n1661) );
  XOR U1755 ( .A(key[127]), .B(n1665), .Z(n1664) );
  XNOR U1756 ( .A(n1666), .B(n1667), .Z(out[126]) );
  XNOR U1757 ( .A(key[126]), .B(n1668), .Z(n1667) );
  XOR U1758 ( .A(n1669), .B(n1670), .Z(out[125]) );
  XNOR U1759 ( .A(n1671), .B(n1672), .Z(n1670) );
  XOR U1760 ( .A(n1663), .B(n1673), .Z(n1672) );
  XOR U1761 ( .A(n1674), .B(n1675), .Z(n1663) );
  XNOR U1762 ( .A(n1676), .B(n1677), .Z(n1675) );
  NANDN U1763 ( .A(n1678), .B(n1679), .Z(n1677) );
  XOR U1764 ( .A(n1680), .B(n1681), .Z(n1669) );
  XOR U1765 ( .A(key[125]), .B(n1682), .Z(n1681) );
  ANDN U1766 ( .B(n1683), .A(n1684), .Z(n1680) );
  XNOR U1767 ( .A(n1685), .B(n1686), .Z(out[124]) );
  XOR U1768 ( .A(key[124]), .B(n1671), .Z(n1686) );
  XOR U1769 ( .A(n1687), .B(n1688), .Z(out[123]) );
  XOR U1770 ( .A(n1689), .B(n1666), .Z(n1688) );
  XNOR U1771 ( .A(n1690), .B(n1691), .Z(n1666) );
  XNOR U1772 ( .A(n1692), .B(n1682), .Z(n1691) );
  NOR U1773 ( .A(n1693), .B(n1694), .Z(n1682) );
  ANDN U1774 ( .B(n1695), .A(n1696), .Z(n1692) );
  XNOR U1775 ( .A(n1697), .B(n1698), .Z(n1687) );
  XNOR U1776 ( .A(key[123]), .B(n1699), .Z(n1698) );
  XOR U1777 ( .A(key[122]), .B(n1685), .Z(out[122]) );
  XOR U1778 ( .A(n1665), .B(n1700), .Z(n1685) );
  XOR U1779 ( .A(n1701), .B(n1662), .Z(out[121]) );
  XOR U1780 ( .A(n1690), .B(n1702), .Z(n1689) );
  XNOR U1781 ( .A(n1703), .B(n1704), .Z(n1702) );
  NANDN U1782 ( .A(n1678), .B(n1705), .Z(n1704) );
  XNOR U1783 ( .A(n1673), .B(n1706), .Z(n1690) );
  XNOR U1784 ( .A(n1707), .B(n1708), .Z(n1706) );
  NANDN U1785 ( .A(n1709), .B(n1710), .Z(n1708) );
  XOR U1786 ( .A(n1700), .B(n1697), .Z(n1668) );
  XNOR U1787 ( .A(n1673), .B(n1711), .Z(n1697) );
  XNOR U1788 ( .A(n1703), .B(n1712), .Z(n1711) );
  NAND U1789 ( .A(n1713), .B(n1714), .Z(n1712) );
  OR U1790 ( .A(n1715), .B(n1716), .Z(n1703) );
  XOR U1791 ( .A(n1717), .B(n1707), .Z(n1673) );
  NANDN U1792 ( .A(n1718), .B(n1719), .Z(n1707) );
  AND U1793 ( .A(n1720), .B(n1721), .Z(n1717) );
  XOR U1794 ( .A(key[121]), .B(n1665), .Z(n1701) );
  IV U1795 ( .A(n1699), .Z(n1665) );
  XNOR U1796 ( .A(n1722), .B(n1723), .Z(n1699) );
  XNOR U1797 ( .A(n1724), .B(n1725), .Z(n1723) );
  NANDN U1798 ( .A(n1684), .B(n1726), .Z(n1725) );
  XNOR U1799 ( .A(n1671), .B(n1727), .Z(out[120]) );
  XOR U1800 ( .A(key[120]), .B(n1700), .Z(n1727) );
  XNOR U1801 ( .A(n1722), .B(n1728), .Z(n1700) );
  XOR U1802 ( .A(n1729), .B(n1676), .Z(n1728) );
  OR U1803 ( .A(n1730), .B(n1715), .Z(n1676) );
  XNOR U1804 ( .A(n1678), .B(n1731), .Z(n1715) );
  AND U1805 ( .A(n1732), .B(n1713), .Z(n1729) );
  XNOR U1806 ( .A(n1674), .B(n1733), .Z(n1671) );
  XOR U1807 ( .A(n1734), .B(n1724), .Z(n1733) );
  OR U1808 ( .A(n1735), .B(n1693), .Z(n1724) );
  XNOR U1809 ( .A(n1696), .B(n1684), .Z(n1693) );
  NOR U1810 ( .A(n1736), .B(n1696), .Z(n1734) );
  XNOR U1811 ( .A(n1722), .B(n1737), .Z(n1674) );
  XNOR U1812 ( .A(n1738), .B(n1739), .Z(n1737) );
  NANDN U1813 ( .A(n1709), .B(n1740), .Z(n1739) );
  XOR U1814 ( .A(n1741), .B(n1738), .Z(n1722) );
  OR U1815 ( .A(n1718), .B(n1742), .Z(n1738) );
  XOR U1816 ( .A(n1720), .B(n1709), .Z(n1718) );
  XNOR U1817 ( .A(n1731), .B(n1684), .Z(n1709) );
  XOR U1818 ( .A(n1743), .B(n1744), .Z(n1684) );
  NANDN U1819 ( .A(n1745), .B(n1746), .Z(n1744) );
  IV U1820 ( .A(n1713), .Z(n1731) );
  XOR U1821 ( .A(n1747), .B(n1748), .Z(n1713) );
  NANDN U1822 ( .A(n1745), .B(n1749), .Z(n1748) );
  ANDN U1823 ( .B(n1720), .A(n1750), .Z(n1741) );
  XOR U1824 ( .A(n1696), .B(n1678), .Z(n1720) );
  XOR U1825 ( .A(n1751), .B(n1747), .Z(n1678) );
  NANDN U1826 ( .A(n1752), .B(n1753), .Z(n1747) );
  AND U1827 ( .A(n1754), .B(n1755), .Z(n1751) );
  ANDN U1828 ( .B(n1757), .A(n1752), .Z(n1743) );
  XOR U1829 ( .A(n1758), .B(n1759), .Z(n1745) );
  XNOR U1830 ( .A(n1761), .B(n1762), .Z(n1758) );
  XNOR U1831 ( .A(n1763), .B(n1764), .Z(n1762) );
  AND U1832 ( .A(n1765), .B(n1754), .Z(n1763) );
  AND U1833 ( .A(n1765), .B(n1755), .Z(n1756) );
  XOR U1834 ( .A(n1761), .B(n1766), .Z(n1755) );
  XOR U1835 ( .A(n1767), .B(n1764), .Z(n1766) );
  NAND U1836 ( .A(n1753), .B(n1757), .Z(n1764) );
  XOR U1837 ( .A(n1746), .B(n1765), .Z(n1757) );
  XOR U1838 ( .A(n1749), .B(n1754), .Z(n1753) );
  XNOR U1839 ( .A(n1768), .B(n1769), .Z(n1754) );
  XOR U1840 ( .A(n1770), .B(n1771), .Z(n1769) );
  XNOR U1841 ( .A(n1772), .B(n1773), .Z(n1768) );
  ANDN U1842 ( .B(n1695), .A(n1736), .Z(n1772) );
  AND U1843 ( .A(n1746), .B(n1749), .Z(n1767) );
  XNOR U1844 ( .A(n1746), .B(n1749), .Z(n1761) );
  XNOR U1845 ( .A(n1774), .B(n1775), .Z(n1749) );
  XOR U1846 ( .A(n1776), .B(n1777), .Z(n1775) );
  XOR U1847 ( .A(n1770), .B(n1778), .Z(n1774) );
  XNOR U1848 ( .A(n1779), .B(n1773), .Z(n1778) );
  OR U1849 ( .A(n1694), .B(n1735), .Z(n1773) );
  XOR U1850 ( .A(n1736), .B(n1726), .Z(n1735) );
  XOR U1851 ( .A(n1780), .B(n1683), .Z(n1694) );
  AND U1852 ( .A(n1683), .B(n1726), .Z(n1779) );
  XNOR U1853 ( .A(n1781), .B(n1782), .Z(n1746) );
  XOR U1854 ( .A(n1783), .B(n1784), .Z(n1782) );
  XNOR U1855 ( .A(n1705), .B(n1770), .Z(n1784) );
  XNOR U1856 ( .A(n1736), .B(n1695), .Z(n1770) );
  XOR U1857 ( .A(n1679), .B(n1785), .Z(n1781) );
  XNOR U1858 ( .A(n1786), .B(n1787), .Z(n1785) );
  AND U1859 ( .A(n1714), .B(n1732), .Z(n1786) );
  IV U1860 ( .A(n1760), .Z(n1765) );
  XOR U1861 ( .A(n1788), .B(n1789), .Z(n1760) );
  XNOR U1862 ( .A(n1771), .B(n1790), .Z(n1789) );
  XNOR U1863 ( .A(n1714), .B(n1777), .Z(n1790) );
  XOR U1864 ( .A(n1783), .B(n1791), .Z(n1771) );
  XNOR U1865 ( .A(n1792), .B(n1793), .Z(n1791) );
  NAND U1866 ( .A(n1710), .B(n1740), .Z(n1793) );
  IV U1867 ( .A(n1776), .Z(n1783) );
  XOR U1868 ( .A(n1794), .B(n1792), .Z(n1776) );
  NANDN U1869 ( .A(n1742), .B(n1719), .Z(n1792) );
  XOR U1870 ( .A(n1714), .B(n1683), .Z(n1710) );
  XOR U1871 ( .A(n1795), .B(n1796), .Z(n1683) );
  XOR U1872 ( .A(n1797), .B(n1798), .Z(n1796) );
  XOR U1873 ( .A(n1750), .B(n1740), .Z(n1742) );
  ANDN U1874 ( .B(n1721), .A(n1750), .Z(n1794) );
  XNOR U1875 ( .A(n1799), .B(n1736), .Z(n1750) );
  XNOR U1876 ( .A(n1800), .B(n1801), .Z(n1736) );
  XOR U1877 ( .A(n1802), .B(n1797), .Z(n1800) );
  XOR U1878 ( .A(n1732), .B(n1803), .Z(n1788) );
  XNOR U1879 ( .A(n1804), .B(n1787), .Z(n1803) );
  OR U1880 ( .A(n1716), .B(n1730), .Z(n1787) );
  XNOR U1881 ( .A(n1679), .B(n1732), .Z(n1730) );
  XNOR U1882 ( .A(n1705), .B(n1714), .Z(n1716) );
  XOR U1883 ( .A(n1780), .B(n1805), .Z(n1714) );
  XOR U1884 ( .A(state[122]), .B(key[122]), .Z(n1801) );
  IV U1885 ( .A(n1695), .Z(n1780) );
  XOR U1886 ( .A(n1795), .B(n1806), .Z(n1695) );
  XNOR U1887 ( .A(n1797), .B(n1807), .Z(n1806) );
  AND U1888 ( .A(n1679), .B(n1705), .Z(n1804) );
  XOR U1889 ( .A(n1795), .B(n1808), .Z(n1705) );
  XNOR U1890 ( .A(n1797), .B(n1809), .Z(n1808) );
  XOR U1891 ( .A(n1799), .B(n1810), .Z(n1797) );
  XNOR U1892 ( .A(state[126]), .B(key[126]), .Z(n1810) );
  XNOR U1893 ( .A(state[125]), .B(key[125]), .Z(n1795) );
  XNOR U1894 ( .A(n1811), .B(n1812), .Z(n1732) );
  XNOR U1895 ( .A(n1809), .B(n1807), .Z(n1812) );
  XOR U1896 ( .A(state[127]), .B(key[127]), .Z(n1807) );
  XOR U1897 ( .A(state[124]), .B(key[124]), .Z(n1809) );
  XOR U1898 ( .A(n1679), .B(n1802), .Z(n1811) );
  XOR U1899 ( .A(n1798), .B(n1813), .Z(n1802) );
  XNOR U1900 ( .A(state[123]), .B(key[123]), .Z(n1813) );
  XNOR U1901 ( .A(state[121]), .B(key[121]), .Z(n1798) );
  IV U1902 ( .A(n1799), .Z(n1679) );
  XNOR U1903 ( .A(state[120]), .B(key[120]), .Z(n1799) );
  XOR U1904 ( .A(n1814), .B(n1815), .Z(out[11]) );
  XNOR U1905 ( .A(n4), .B(n1630), .Z(n1815) );
  XNOR U1906 ( .A(n1816), .B(n1817), .Z(n1630) );
  XNOR U1907 ( .A(n1818), .B(n1645), .Z(n1817) );
  NOR U1908 ( .A(n1819), .B(n1820), .Z(n1645) );
  ANDN U1909 ( .B(n1821), .A(n1654), .Z(n1818) );
  XNOR U1910 ( .A(n1632), .B(n1822), .Z(n1814) );
  XOR U1911 ( .A(key[11]), .B(n5), .Z(n1822) );
  XOR U1912 ( .A(n1816), .B(n1823), .Z(n5) );
  XNOR U1913 ( .A(n1824), .B(n1825), .Z(n1823) );
  NANDN U1914 ( .A(n1641), .B(n1826), .Z(n1825) );
  XNOR U1915 ( .A(n1636), .B(n1827), .Z(n1816) );
  XNOR U1916 ( .A(n1828), .B(n1829), .Z(n1827) );
  NANDN U1917 ( .A(n1659), .B(n1830), .Z(n1829) );
  XNOR U1918 ( .A(n1636), .B(n1831), .Z(n1632) );
  XNOR U1919 ( .A(n1824), .B(n1832), .Z(n1831) );
  NANDN U1920 ( .A(n1833), .B(n1834), .Z(n1832) );
  OR U1921 ( .A(n1835), .B(n1836), .Z(n1824) );
  XOR U1922 ( .A(n1837), .B(n1828), .Z(n1636) );
  OR U1923 ( .A(n1838), .B(n1839), .Z(n1828) );
  XOR U1924 ( .A(n1842), .B(n1843), .Z(out[119]) );
  XOR U1925 ( .A(n1844), .B(n1845), .Z(n1842) );
  XOR U1926 ( .A(key[119]), .B(n1846), .Z(n1845) );
  XNOR U1927 ( .A(n1847), .B(n1848), .Z(out[118]) );
  XNOR U1928 ( .A(key[118]), .B(n1849), .Z(n1848) );
  XOR U1929 ( .A(n1850), .B(n1851), .Z(out[117]) );
  XNOR U1930 ( .A(n1852), .B(n1853), .Z(n1851) );
  XOR U1931 ( .A(n1844), .B(n1854), .Z(n1853) );
  XOR U1932 ( .A(n1855), .B(n1856), .Z(n1844) );
  XNOR U1933 ( .A(n1857), .B(n1858), .Z(n1856) );
  NANDN U1934 ( .A(n1859), .B(n1860), .Z(n1858) );
  XOR U1935 ( .A(n1861), .B(n1862), .Z(n1850) );
  XOR U1936 ( .A(key[117]), .B(n1863), .Z(n1862) );
  ANDN U1937 ( .B(n1864), .A(n1865), .Z(n1861) );
  XNOR U1938 ( .A(n1866), .B(n1867), .Z(out[116]) );
  XOR U1939 ( .A(key[116]), .B(n1852), .Z(n1867) );
  XOR U1940 ( .A(n1868), .B(n1869), .Z(out[115]) );
  XOR U1941 ( .A(n1870), .B(n1847), .Z(n1869) );
  XNOR U1942 ( .A(n1871), .B(n1872), .Z(n1847) );
  XNOR U1943 ( .A(n1873), .B(n1863), .Z(n1872) );
  NOR U1944 ( .A(n1874), .B(n1875), .Z(n1863) );
  ANDN U1945 ( .B(n1876), .A(n1877), .Z(n1873) );
  XNOR U1946 ( .A(n1878), .B(n1879), .Z(n1868) );
  XNOR U1947 ( .A(key[115]), .B(n1880), .Z(n1879) );
  XOR U1948 ( .A(key[114]), .B(n1866), .Z(out[114]) );
  XOR U1949 ( .A(n1846), .B(n1881), .Z(n1866) );
  XOR U1950 ( .A(n1882), .B(n1843), .Z(out[113]) );
  XOR U1951 ( .A(n1871), .B(n1883), .Z(n1870) );
  XNOR U1952 ( .A(n1884), .B(n1885), .Z(n1883) );
  NANDN U1953 ( .A(n1859), .B(n1886), .Z(n1885) );
  XNOR U1954 ( .A(n1854), .B(n1887), .Z(n1871) );
  XNOR U1955 ( .A(n1888), .B(n1889), .Z(n1887) );
  NANDN U1956 ( .A(n1890), .B(n1891), .Z(n1889) );
  XOR U1957 ( .A(n1881), .B(n1878), .Z(n1849) );
  XNOR U1958 ( .A(n1854), .B(n1892), .Z(n1878) );
  XNOR U1959 ( .A(n1884), .B(n1893), .Z(n1892) );
  NAND U1960 ( .A(n1894), .B(n1895), .Z(n1893) );
  OR U1961 ( .A(n1896), .B(n1897), .Z(n1884) );
  XOR U1962 ( .A(n1898), .B(n1888), .Z(n1854) );
  NANDN U1963 ( .A(n1899), .B(n1900), .Z(n1888) );
  AND U1964 ( .A(n1901), .B(n1902), .Z(n1898) );
  XOR U1965 ( .A(key[113]), .B(n1846), .Z(n1882) );
  IV U1966 ( .A(n1880), .Z(n1846) );
  XNOR U1967 ( .A(n1903), .B(n1904), .Z(n1880) );
  XNOR U1968 ( .A(n1905), .B(n1906), .Z(n1904) );
  OR U1969 ( .A(n1907), .B(n1865), .Z(n1906) );
  XNOR U1970 ( .A(n1852), .B(n1908), .Z(out[112]) );
  XOR U1971 ( .A(key[112]), .B(n1881), .Z(n1908) );
  XNOR U1972 ( .A(n1903), .B(n1909), .Z(n1881) );
  XOR U1973 ( .A(n1910), .B(n1857), .Z(n1909) );
  OR U1974 ( .A(n1911), .B(n1896), .Z(n1857) );
  XNOR U1975 ( .A(n1859), .B(n1912), .Z(n1896) );
  AND U1976 ( .A(n1913), .B(n1894), .Z(n1910) );
  XNOR U1977 ( .A(n1855), .B(n1914), .Z(n1852) );
  XOR U1978 ( .A(n1915), .B(n1905), .Z(n1914) );
  OR U1979 ( .A(n1916), .B(n1874), .Z(n1905) );
  XNOR U1980 ( .A(n1877), .B(n1865), .Z(n1874) );
  NOR U1981 ( .A(n1917), .B(n1877), .Z(n1915) );
  XNOR U1982 ( .A(n1903), .B(n1918), .Z(n1855) );
  XNOR U1983 ( .A(n1919), .B(n1920), .Z(n1918) );
  NANDN U1984 ( .A(n1890), .B(n1921), .Z(n1920) );
  XOR U1985 ( .A(n1922), .B(n1919), .Z(n1903) );
  OR U1986 ( .A(n1899), .B(n1923), .Z(n1919) );
  XOR U1987 ( .A(n1901), .B(n1890), .Z(n1899) );
  XNOR U1988 ( .A(n1912), .B(n1865), .Z(n1890) );
  XOR U1989 ( .A(n1924), .B(n1925), .Z(n1865) );
  NANDN U1990 ( .A(n1926), .B(n1927), .Z(n1925) );
  IV U1991 ( .A(n1894), .Z(n1912) );
  XOR U1992 ( .A(n1928), .B(n1929), .Z(n1894) );
  NANDN U1993 ( .A(n1926), .B(n1930), .Z(n1929) );
  ANDN U1994 ( .B(n1901), .A(n1931), .Z(n1922) );
  XOR U1995 ( .A(n1877), .B(n1859), .Z(n1901) );
  XOR U1996 ( .A(n1932), .B(n1928), .Z(n1859) );
  NANDN U1997 ( .A(n1933), .B(n1934), .Z(n1928) );
  AND U1998 ( .A(n1935), .B(n1936), .Z(n1932) );
  ANDN U1999 ( .B(n1938), .A(n1933), .Z(n1924) );
  XOR U2000 ( .A(n1939), .B(n1940), .Z(n1926) );
  XNOR U2001 ( .A(n1942), .B(n1943), .Z(n1939) );
  XNOR U2002 ( .A(n1944), .B(n1945), .Z(n1943) );
  AND U2003 ( .A(n1946), .B(n1935), .Z(n1944) );
  AND U2004 ( .A(n1946), .B(n1936), .Z(n1937) );
  XOR U2005 ( .A(n1942), .B(n1947), .Z(n1936) );
  XOR U2006 ( .A(n1948), .B(n1945), .Z(n1947) );
  NAND U2007 ( .A(n1934), .B(n1938), .Z(n1945) );
  XOR U2008 ( .A(n1927), .B(n1946), .Z(n1938) );
  XOR U2009 ( .A(n1930), .B(n1935), .Z(n1934) );
  XNOR U2010 ( .A(n1949), .B(n1950), .Z(n1935) );
  XOR U2011 ( .A(n1951), .B(n1952), .Z(n1950) );
  XNOR U2012 ( .A(n1953), .B(n1954), .Z(n1949) );
  ANDN U2013 ( .B(n1876), .A(n1917), .Z(n1953) );
  AND U2014 ( .A(n1927), .B(n1930), .Z(n1948) );
  XNOR U2015 ( .A(n1927), .B(n1930), .Z(n1942) );
  XNOR U2016 ( .A(n1955), .B(n1956), .Z(n1930) );
  XOR U2017 ( .A(n1957), .B(n1958), .Z(n1956) );
  XOR U2018 ( .A(n1951), .B(n1959), .Z(n1955) );
  XNOR U2019 ( .A(n1960), .B(n1954), .Z(n1959) );
  OR U2020 ( .A(n1875), .B(n1916), .Z(n1954) );
  XNOR U2021 ( .A(n1917), .B(n1907), .Z(n1916) );
  XOR U2022 ( .A(n1961), .B(n1864), .Z(n1875) );
  ANDN U2023 ( .B(n1864), .A(n1907), .Z(n1960) );
  XNOR U2024 ( .A(n1962), .B(n1963), .Z(n1927) );
  XOR U2025 ( .A(n1964), .B(n1965), .Z(n1963) );
  XNOR U2026 ( .A(n1886), .B(n1951), .Z(n1965) );
  XNOR U2027 ( .A(n1917), .B(n1876), .Z(n1951) );
  XOR U2028 ( .A(n1860), .B(n1966), .Z(n1962) );
  XNOR U2029 ( .A(n1967), .B(n1968), .Z(n1966) );
  AND U2030 ( .A(n1895), .B(n1913), .Z(n1967) );
  IV U2031 ( .A(n1941), .Z(n1946) );
  XOR U2032 ( .A(n1969), .B(n1970), .Z(n1941) );
  XNOR U2033 ( .A(n1952), .B(n1971), .Z(n1970) );
  XNOR U2034 ( .A(n1895), .B(n1958), .Z(n1971) );
  XNOR U2035 ( .A(n1907), .B(n1864), .Z(n1958) );
  XOR U2036 ( .A(n1964), .B(n1972), .Z(n1952) );
  XNOR U2037 ( .A(n1973), .B(n1974), .Z(n1972) );
  NAND U2038 ( .A(n1891), .B(n1921), .Z(n1974) );
  IV U2039 ( .A(n1957), .Z(n1964) );
  XOR U2040 ( .A(n1975), .B(n1973), .Z(n1957) );
  NANDN U2041 ( .A(n1923), .B(n1900), .Z(n1973) );
  XOR U2042 ( .A(n1895), .B(n1864), .Z(n1891) );
  XOR U2043 ( .A(n1976), .B(n1977), .Z(n1864) );
  XOR U2044 ( .A(n1978), .B(n1979), .Z(n1977) );
  XOR U2045 ( .A(n1931), .B(n1921), .Z(n1923) );
  XOR U2046 ( .A(n1978), .B(n1976), .Z(n1907) );
  ANDN U2047 ( .B(n1902), .A(n1931), .Z(n1975) );
  XNOR U2048 ( .A(n1980), .B(n1917), .Z(n1931) );
  XOR U2049 ( .A(n1981), .B(n1982), .Z(n1917) );
  XNOR U2050 ( .A(n1983), .B(n1978), .Z(n1981) );
  XOR U2051 ( .A(n1913), .B(n1984), .Z(n1969) );
  XNOR U2052 ( .A(n1985), .B(n1968), .Z(n1984) );
  OR U2053 ( .A(n1897), .B(n1911), .Z(n1968) );
  XNOR U2054 ( .A(n1860), .B(n1913), .Z(n1911) );
  XNOR U2055 ( .A(n1886), .B(n1895), .Z(n1897) );
  XOR U2056 ( .A(n1961), .B(n1986), .Z(n1895) );
  XNOR U2057 ( .A(n1979), .B(n1982), .Z(n1986) );
  XNOR U2058 ( .A(state[82]), .B(key[82]), .Z(n1982) );
  IV U2059 ( .A(n1876), .Z(n1961) );
  XOR U2060 ( .A(n1976), .B(n1987), .Z(n1876) );
  XOR U2061 ( .A(n1978), .B(n1988), .Z(n1987) );
  AND U2062 ( .A(n1860), .B(n1886), .Z(n1985) );
  XOR U2063 ( .A(n1976), .B(n1989), .Z(n1886) );
  XOR U2064 ( .A(n1978), .B(n1990), .Z(n1989) );
  XOR U2065 ( .A(n1980), .B(n1991), .Z(n1978) );
  XNOR U2066 ( .A(state[86]), .B(key[86]), .Z(n1991) );
  XNOR U2067 ( .A(state[85]), .B(key[85]), .Z(n1976) );
  XNOR U2068 ( .A(n1992), .B(n1993), .Z(n1913) );
  XNOR U2069 ( .A(n1990), .B(n1988), .Z(n1993) );
  XNOR U2070 ( .A(state[87]), .B(key[87]), .Z(n1988) );
  XNOR U2071 ( .A(state[84]), .B(key[84]), .Z(n1990) );
  XNOR U2072 ( .A(n1860), .B(n1983), .Z(n1992) );
  XNOR U2073 ( .A(n1979), .B(n1994), .Z(n1983) );
  XNOR U2074 ( .A(state[83]), .B(key[83]), .Z(n1994) );
  XNOR U2075 ( .A(state[81]), .B(key[81]), .Z(n1979) );
  IV U2076 ( .A(n1980), .Z(n1860) );
  XNOR U2077 ( .A(state[80]), .B(key[80]), .Z(n1980) );
  XOR U2078 ( .A(n1995), .B(n1996), .Z(out[111]) );
  XOR U2079 ( .A(n1997), .B(n1998), .Z(n1995) );
  XOR U2080 ( .A(key[111]), .B(n1999), .Z(n1998) );
  XNOR U2081 ( .A(n2000), .B(n2001), .Z(out[110]) );
  XNOR U2082 ( .A(key[110]), .B(n2002), .Z(n2001) );
  XOR U2083 ( .A(key[10]), .B(n1648), .Z(out[10]) );
  XOR U2084 ( .A(n62), .B(n4), .Z(n1648) );
  XNOR U2085 ( .A(n1655), .B(n2003), .Z(n4) );
  XNOR U2086 ( .A(n1652), .B(n2004), .Z(n2003) );
  NAND U2087 ( .A(n1647), .B(n2005), .Z(n2004) );
  OR U2088 ( .A(n2006), .B(n1819), .Z(n1652) );
  XNOR U2089 ( .A(n1654), .B(n2007), .Z(n1819) );
  XOR U2090 ( .A(n1655), .B(n2008), .Z(n62) );
  XOR U2091 ( .A(n2009), .B(n1639), .Z(n2008) );
  OR U2092 ( .A(n1835), .B(n2010), .Z(n1639) );
  XNOR U2093 ( .A(n1641), .B(n1833), .Z(n1835) );
  ANDN U2094 ( .B(n2011), .A(n1833), .Z(n2009) );
  XOR U2095 ( .A(n2012), .B(n1657), .Z(n1655) );
  OR U2096 ( .A(n1839), .B(n2013), .Z(n1657) );
  XNOR U2097 ( .A(n1841), .B(n1659), .Z(n1839) );
  XNOR U2098 ( .A(n1833), .B(n2007), .Z(n1659) );
  IV U2099 ( .A(n1647), .Z(n2007) );
  XOR U2100 ( .A(n2014), .B(n2015), .Z(n1647) );
  NANDN U2101 ( .A(n2016), .B(n2017), .Z(n2015) );
  XOR U2102 ( .A(n2018), .B(n2019), .Z(n1833) );
  NANDN U2103 ( .A(n2016), .B(n2020), .Z(n2019) );
  NOR U2104 ( .A(n1841), .B(n2021), .Z(n2012) );
  XNOR U2105 ( .A(n1641), .B(n1654), .Z(n1841) );
  XOR U2106 ( .A(n2022), .B(n2014), .Z(n1654) );
  NANDN U2107 ( .A(n2023), .B(n2024), .Z(n2014) );
  XNOR U2108 ( .A(n2017), .B(n2025), .Z(n2024) );
  AND U2109 ( .A(n2026), .B(n2027), .Z(n2022) );
  ANDN U2110 ( .B(n2029), .A(n2023), .Z(n2018) );
  XOR U2111 ( .A(n2030), .B(n2031), .Z(n2016) );
  XNOR U2112 ( .A(n2026), .B(n2032), .Z(n2031) );
  XNOR U2113 ( .A(n2033), .B(n2034), .Z(n2030) );
  XNOR U2114 ( .A(n2035), .B(n2036), .Z(n2034) );
  AND U2115 ( .A(n2032), .B(n2026), .Z(n2035) );
  AND U2116 ( .A(n2032), .B(n2027), .Z(n2028) );
  XOR U2117 ( .A(n2033), .B(n2037), .Z(n2027) );
  XOR U2118 ( .A(n2038), .B(n2036), .Z(n2037) );
  NAND U2119 ( .A(n2029), .B(n2039), .Z(n2036) );
  XOR U2120 ( .A(n2017), .B(n2026), .Z(n2039) );
  IV U2121 ( .A(n2025), .Z(n2026) );
  XOR U2122 ( .A(n2040), .B(n2041), .Z(n2025) );
  XNOR U2123 ( .A(n2042), .B(n2043), .Z(n2041) );
  XNOR U2124 ( .A(n2011), .B(n2044), .Z(n2043) );
  XOR U2125 ( .A(n1834), .B(n2045), .Z(n2040) );
  XNOR U2126 ( .A(n2046), .B(n2047), .Z(n2045) );
  AND U2127 ( .A(n1642), .B(n1826), .Z(n2046) );
  XOR U2128 ( .A(n2020), .B(n2032), .Z(n2029) );
  AND U2129 ( .A(n2017), .B(n2020), .Z(n2038) );
  XNOR U2130 ( .A(n2017), .B(n2020), .Z(n2033) );
  XNOR U2131 ( .A(n2048), .B(n2049), .Z(n2020) );
  XOR U2132 ( .A(n2050), .B(n2044), .Z(n2049) );
  XNOR U2133 ( .A(n2051), .B(n2005), .Z(n2044) );
  XOR U2134 ( .A(n2052), .B(n2053), .Z(n2048) );
  XNOR U2135 ( .A(n2054), .B(n2055), .Z(n2053) );
  AND U2136 ( .A(n2005), .B(n1646), .Z(n2054) );
  IV U2137 ( .A(n2051), .Z(n1646) );
  XNOR U2138 ( .A(n2056), .B(n2057), .Z(n2017) );
  XOR U2139 ( .A(n2058), .B(n2059), .Z(n2057) );
  XNOR U2140 ( .A(n1826), .B(n2052), .Z(n2059) );
  XOR U2141 ( .A(n1642), .B(n2060), .Z(n2056) );
  XNOR U2142 ( .A(n2061), .B(n2047), .Z(n2060) );
  OR U2143 ( .A(n1836), .B(n2010), .Z(n2047) );
  XNOR U2144 ( .A(n1642), .B(n2011), .Z(n2010) );
  XNOR U2145 ( .A(n1826), .B(n1834), .Z(n1836) );
  AND U2146 ( .A(n1834), .B(n2011), .Z(n2061) );
  XNOR U2147 ( .A(n2062), .B(n2063), .Z(n2032) );
  XNOR U2148 ( .A(n2050), .B(n2042), .Z(n2063) );
  XOR U2149 ( .A(n2052), .B(n2064), .Z(n2042) );
  XNOR U2150 ( .A(n2065), .B(n2066), .Z(n2064) );
  NAND U2151 ( .A(n1660), .B(n1830), .Z(n2066) );
  XNOR U2152 ( .A(n2067), .B(n2065), .Z(n2052) );
  OR U2153 ( .A(n2013), .B(n1838), .Z(n2065) );
  XNOR U2154 ( .A(n1840), .B(n1830), .Z(n1838) );
  XNOR U2155 ( .A(n2051), .B(n1834), .Z(n1830) );
  XNOR U2156 ( .A(n2068), .B(n2069), .Z(n1834) );
  XNOR U2157 ( .A(n1821), .B(n2070), .Z(n2069) );
  XOR U2158 ( .A(n2021), .B(n1660), .Z(n2013) );
  XNOR U2159 ( .A(n2071), .B(n2072), .Z(n2011) );
  XNOR U2160 ( .A(n2073), .B(n2074), .Z(n2072) );
  XNOR U2161 ( .A(n1642), .B(n2075), .Z(n2071) );
  ANDN U2162 ( .B(n1840), .A(n2021), .Z(n2067) );
  XOR U2163 ( .A(n1642), .B(n2076), .Z(n2021) );
  XNOR U2164 ( .A(n2077), .B(n1826), .Z(n1840) );
  XNOR U2165 ( .A(n2074), .B(n2078), .Z(n1826) );
  XOR U2166 ( .A(state[76]), .B(key[76]), .Z(n2074) );
  IV U2167 ( .A(n2058), .Z(n2050) );
  XNOR U2168 ( .A(n2077), .B(n1653), .Z(n2058) );
  IV U2169 ( .A(n1821), .Z(n2077) );
  XNOR U2170 ( .A(n2079), .B(n2055), .Z(n2062) );
  OR U2171 ( .A(n1820), .B(n2006), .Z(n2055) );
  XOR U2172 ( .A(n2076), .B(n2005), .Z(n2006) );
  XNOR U2173 ( .A(n2080), .B(n2081), .Z(n2005) );
  XOR U2174 ( .A(n1821), .B(n2051), .Z(n1820) );
  XOR U2175 ( .A(n2070), .B(n2082), .Z(n2051) );
  AND U2176 ( .A(n1821), .B(n1653), .Z(n2079) );
  IV U2177 ( .A(n2076), .Z(n1653) );
  XOR U2178 ( .A(n2073), .B(n2083), .Z(n2076) );
  XNOR U2179 ( .A(n2080), .B(n2068), .Z(n2083) );
  XOR U2180 ( .A(state[74]), .B(key[74]), .Z(n2068) );
  XNOR U2181 ( .A(n2070), .B(n2084), .Z(n2073) );
  XNOR U2182 ( .A(state[75]), .B(key[75]), .Z(n2084) );
  XOR U2183 ( .A(state[73]), .B(key[73]), .Z(n2070) );
  XOR U2184 ( .A(n2075), .B(n2078), .Z(n1821) );
  XOR U2185 ( .A(n2080), .B(n2081), .Z(n2078) );
  XNOR U2186 ( .A(state[77]), .B(key[77]), .Z(n2081) );
  XNOR U2187 ( .A(n1642), .B(n2085), .Z(n2080) );
  XNOR U2188 ( .A(state[78]), .B(key[78]), .Z(n2085) );
  XOR U2189 ( .A(state[72]), .B(key[72]), .Z(n1642) );
  XNOR U2190 ( .A(state[79]), .B(key[79]), .Z(n2075) );
  XOR U2191 ( .A(n2086), .B(n2087), .Z(out[109]) );
  XNOR U2192 ( .A(n2088), .B(n2089), .Z(n2087) );
  XOR U2193 ( .A(n1997), .B(n2090), .Z(n2089) );
  XOR U2194 ( .A(n2091), .B(n2092), .Z(n1997) );
  XNOR U2195 ( .A(n2093), .B(n2094), .Z(n2092) );
  NANDN U2196 ( .A(n2095), .B(n2096), .Z(n2094) );
  XOR U2197 ( .A(n2097), .B(n2098), .Z(n2086) );
  XOR U2198 ( .A(key[109]), .B(n2099), .Z(n2098) );
  ANDN U2199 ( .B(n2100), .A(n2101), .Z(n2097) );
  XNOR U2200 ( .A(n2102), .B(n2103), .Z(out[108]) );
  XOR U2201 ( .A(key[108]), .B(n2088), .Z(n2103) );
  XOR U2202 ( .A(n2104), .B(n2105), .Z(out[107]) );
  XOR U2203 ( .A(n2106), .B(n2000), .Z(n2105) );
  XNOR U2204 ( .A(n2107), .B(n2108), .Z(n2000) );
  XNOR U2205 ( .A(n2109), .B(n2099), .Z(n2108) );
  NOR U2206 ( .A(n2110), .B(n2111), .Z(n2099) );
  ANDN U2207 ( .B(n2112), .A(n2113), .Z(n2109) );
  XNOR U2208 ( .A(n2114), .B(n2115), .Z(n2104) );
  XNOR U2209 ( .A(key[107]), .B(n2116), .Z(n2115) );
  XOR U2210 ( .A(key[106]), .B(n2102), .Z(out[106]) );
  XOR U2211 ( .A(n1999), .B(n2117), .Z(n2102) );
  XOR U2212 ( .A(n2118), .B(n1996), .Z(out[105]) );
  XOR U2213 ( .A(n2107), .B(n2119), .Z(n2106) );
  XNOR U2214 ( .A(n2120), .B(n2121), .Z(n2119) );
  NANDN U2215 ( .A(n2095), .B(n2122), .Z(n2121) );
  XNOR U2216 ( .A(n2090), .B(n2123), .Z(n2107) );
  XNOR U2217 ( .A(n2124), .B(n2125), .Z(n2123) );
  NANDN U2218 ( .A(n2126), .B(n2127), .Z(n2125) );
  XOR U2219 ( .A(n2117), .B(n2114), .Z(n2002) );
  XNOR U2220 ( .A(n2090), .B(n2128), .Z(n2114) );
  XNOR U2221 ( .A(n2120), .B(n2129), .Z(n2128) );
  NAND U2222 ( .A(n2130), .B(n2131), .Z(n2129) );
  OR U2223 ( .A(n2132), .B(n2133), .Z(n2120) );
  XOR U2224 ( .A(n2134), .B(n2124), .Z(n2090) );
  NANDN U2225 ( .A(n2135), .B(n2136), .Z(n2124) );
  AND U2226 ( .A(n2137), .B(n2138), .Z(n2134) );
  XOR U2227 ( .A(key[105]), .B(n1999), .Z(n2118) );
  IV U2228 ( .A(n2116), .Z(n1999) );
  XNOR U2229 ( .A(n2139), .B(n2140), .Z(n2116) );
  XNOR U2230 ( .A(n2141), .B(n2142), .Z(n2140) );
  OR U2231 ( .A(n2143), .B(n2101), .Z(n2142) );
  XNOR U2232 ( .A(n2088), .B(n2144), .Z(out[104]) );
  XOR U2233 ( .A(key[104]), .B(n2117), .Z(n2144) );
  XNOR U2234 ( .A(n2139), .B(n2145), .Z(n2117) );
  XOR U2235 ( .A(n2146), .B(n2093), .Z(n2145) );
  OR U2236 ( .A(n2147), .B(n2132), .Z(n2093) );
  XNOR U2237 ( .A(n2095), .B(n2148), .Z(n2132) );
  AND U2238 ( .A(n2149), .B(n2130), .Z(n2146) );
  XNOR U2239 ( .A(n2091), .B(n2150), .Z(n2088) );
  XOR U2240 ( .A(n2151), .B(n2141), .Z(n2150) );
  OR U2241 ( .A(n2152), .B(n2110), .Z(n2141) );
  XNOR U2242 ( .A(n2113), .B(n2101), .Z(n2110) );
  NOR U2243 ( .A(n2153), .B(n2113), .Z(n2151) );
  XNOR U2244 ( .A(n2139), .B(n2154), .Z(n2091) );
  XNOR U2245 ( .A(n2155), .B(n2156), .Z(n2154) );
  NANDN U2246 ( .A(n2126), .B(n2157), .Z(n2156) );
  XOR U2247 ( .A(n2158), .B(n2155), .Z(n2139) );
  OR U2248 ( .A(n2135), .B(n2159), .Z(n2155) );
  XOR U2249 ( .A(n2137), .B(n2126), .Z(n2135) );
  XNOR U2250 ( .A(n2148), .B(n2101), .Z(n2126) );
  XOR U2251 ( .A(n2160), .B(n2161), .Z(n2101) );
  NANDN U2252 ( .A(n2162), .B(n2163), .Z(n2161) );
  IV U2253 ( .A(n2130), .Z(n2148) );
  XOR U2254 ( .A(n2164), .B(n2165), .Z(n2130) );
  NANDN U2255 ( .A(n2162), .B(n2166), .Z(n2165) );
  ANDN U2256 ( .B(n2137), .A(n2167), .Z(n2158) );
  XOR U2257 ( .A(n2113), .B(n2095), .Z(n2137) );
  XOR U2258 ( .A(n2168), .B(n2164), .Z(n2095) );
  NANDN U2259 ( .A(n2169), .B(n2170), .Z(n2164) );
  AND U2260 ( .A(n2171), .B(n2172), .Z(n2168) );
  ANDN U2261 ( .B(n2174), .A(n2169), .Z(n2160) );
  XOR U2262 ( .A(n2175), .B(n2176), .Z(n2162) );
  XNOR U2263 ( .A(n2178), .B(n2179), .Z(n2175) );
  XNOR U2264 ( .A(n2180), .B(n2181), .Z(n2179) );
  AND U2265 ( .A(n2182), .B(n2171), .Z(n2180) );
  AND U2266 ( .A(n2182), .B(n2172), .Z(n2173) );
  XOR U2267 ( .A(n2178), .B(n2183), .Z(n2172) );
  XOR U2268 ( .A(n2184), .B(n2181), .Z(n2183) );
  NAND U2269 ( .A(n2170), .B(n2174), .Z(n2181) );
  XOR U2270 ( .A(n2163), .B(n2182), .Z(n2174) );
  XOR U2271 ( .A(n2166), .B(n2171), .Z(n2170) );
  XNOR U2272 ( .A(n2185), .B(n2186), .Z(n2171) );
  XOR U2273 ( .A(n2187), .B(n2188), .Z(n2186) );
  XNOR U2274 ( .A(n2189), .B(n2190), .Z(n2185) );
  ANDN U2275 ( .B(n2112), .A(n2153), .Z(n2189) );
  AND U2276 ( .A(n2163), .B(n2166), .Z(n2184) );
  XNOR U2277 ( .A(n2163), .B(n2166), .Z(n2178) );
  XNOR U2278 ( .A(n2191), .B(n2192), .Z(n2166) );
  XOR U2279 ( .A(n2193), .B(n2194), .Z(n2192) );
  XOR U2280 ( .A(n2187), .B(n2195), .Z(n2191) );
  XNOR U2281 ( .A(n2196), .B(n2190), .Z(n2195) );
  OR U2282 ( .A(n2111), .B(n2152), .Z(n2190) );
  XNOR U2283 ( .A(n2153), .B(n2143), .Z(n2152) );
  XOR U2284 ( .A(n2197), .B(n2100), .Z(n2111) );
  ANDN U2285 ( .B(n2100), .A(n2143), .Z(n2196) );
  XNOR U2286 ( .A(n2198), .B(n2199), .Z(n2163) );
  XOR U2287 ( .A(n2200), .B(n2201), .Z(n2199) );
  XNOR U2288 ( .A(n2122), .B(n2187), .Z(n2201) );
  XNOR U2289 ( .A(n2153), .B(n2112), .Z(n2187) );
  XOR U2290 ( .A(n2096), .B(n2202), .Z(n2198) );
  XNOR U2291 ( .A(n2203), .B(n2204), .Z(n2202) );
  AND U2292 ( .A(n2131), .B(n2149), .Z(n2203) );
  IV U2293 ( .A(n2177), .Z(n2182) );
  XOR U2294 ( .A(n2205), .B(n2206), .Z(n2177) );
  XNOR U2295 ( .A(n2188), .B(n2207), .Z(n2206) );
  XNOR U2296 ( .A(n2131), .B(n2194), .Z(n2207) );
  XNOR U2297 ( .A(n2143), .B(n2100), .Z(n2194) );
  XOR U2298 ( .A(n2200), .B(n2208), .Z(n2188) );
  XNOR U2299 ( .A(n2209), .B(n2210), .Z(n2208) );
  NAND U2300 ( .A(n2127), .B(n2157), .Z(n2210) );
  IV U2301 ( .A(n2193), .Z(n2200) );
  XOR U2302 ( .A(n2211), .B(n2209), .Z(n2193) );
  NANDN U2303 ( .A(n2159), .B(n2136), .Z(n2209) );
  XOR U2304 ( .A(n2131), .B(n2100), .Z(n2127) );
  XOR U2305 ( .A(n2212), .B(n2213), .Z(n2100) );
  XOR U2306 ( .A(n2214), .B(n2215), .Z(n2213) );
  XOR U2307 ( .A(n2167), .B(n2157), .Z(n2159) );
  XOR U2308 ( .A(n2214), .B(n2212), .Z(n2143) );
  ANDN U2309 ( .B(n2138), .A(n2167), .Z(n2211) );
  XNOR U2310 ( .A(n2216), .B(n2153), .Z(n2167) );
  XOR U2311 ( .A(n2217), .B(n2218), .Z(n2153) );
  XNOR U2312 ( .A(n2219), .B(n2214), .Z(n2217) );
  XOR U2313 ( .A(n2149), .B(n2220), .Z(n2205) );
  XNOR U2314 ( .A(n2221), .B(n2204), .Z(n2220) );
  OR U2315 ( .A(n2133), .B(n2147), .Z(n2204) );
  XNOR U2316 ( .A(n2096), .B(n2149), .Z(n2147) );
  XNOR U2317 ( .A(n2122), .B(n2131), .Z(n2133) );
  XOR U2318 ( .A(n2197), .B(n2222), .Z(n2131) );
  XNOR U2319 ( .A(n2215), .B(n2218), .Z(n2222) );
  XNOR U2320 ( .A(state[42]), .B(key[42]), .Z(n2218) );
  IV U2321 ( .A(n2112), .Z(n2197) );
  XOR U2322 ( .A(n2212), .B(n2223), .Z(n2112) );
  XOR U2323 ( .A(n2214), .B(n2224), .Z(n2223) );
  AND U2324 ( .A(n2096), .B(n2122), .Z(n2221) );
  XOR U2325 ( .A(n2212), .B(n2225), .Z(n2122) );
  XOR U2326 ( .A(n2214), .B(n2226), .Z(n2225) );
  XOR U2327 ( .A(n2216), .B(n2227), .Z(n2214) );
  XNOR U2328 ( .A(state[46]), .B(key[46]), .Z(n2227) );
  XNOR U2329 ( .A(state[45]), .B(key[45]), .Z(n2212) );
  XNOR U2330 ( .A(n2228), .B(n2229), .Z(n2149) );
  XNOR U2331 ( .A(n2226), .B(n2224), .Z(n2229) );
  XNOR U2332 ( .A(state[47]), .B(key[47]), .Z(n2224) );
  XNOR U2333 ( .A(state[44]), .B(key[44]), .Z(n2226) );
  XNOR U2334 ( .A(n2096), .B(n2219), .Z(n2228) );
  XNOR U2335 ( .A(n2215), .B(n2230), .Z(n2219) );
  XNOR U2336 ( .A(state[43]), .B(key[43]), .Z(n2230) );
  XNOR U2337 ( .A(state[41]), .B(key[41]), .Z(n2215) );
  IV U2338 ( .A(n2216), .Z(n2096) );
  XNOR U2339 ( .A(state[40]), .B(key[40]), .Z(n2216) );
  XOR U2340 ( .A(n2231), .B(n2232), .Z(out[103]) );
  XOR U2341 ( .A(n16), .B(n2233), .Z(n2232) );
  IV U2342 ( .A(n2234), .Z(n16) );
  XNOR U2343 ( .A(n8), .B(n2235), .Z(n2231) );
  XOR U2344 ( .A(key[103]), .B(n2236), .Z(n2235) );
  XOR U2345 ( .A(n2237), .B(n2238), .Z(n8) );
  XNOR U2346 ( .A(n2239), .B(n2240), .Z(n2238) );
  NANDN U2347 ( .A(n2241), .B(n2242), .Z(n2240) );
  XNOR U2348 ( .A(n2234), .B(n2243), .Z(out[102]) );
  XNOR U2349 ( .A(key[102]), .B(n10), .Z(n2243) );
  XNOR U2350 ( .A(n2245), .B(n2246), .Z(n2244) );
  NANDN U2351 ( .A(n2247), .B(n2248), .Z(n2246) );
  XOR U2352 ( .A(n2249), .B(n2250), .Z(n2237) );
  XNOR U2353 ( .A(n2251), .B(n2252), .Z(n2250) );
  NANDN U2354 ( .A(n2253), .B(n2254), .Z(n2252) );
  XOR U2355 ( .A(n9), .B(n19), .Z(n2234) );
  XNOR U2356 ( .A(n2249), .B(n2255), .Z(n9) );
  XNOR U2357 ( .A(n2239), .B(n2256), .Z(n2255) );
  NAND U2358 ( .A(n2257), .B(n2258), .Z(n2256) );
  OR U2359 ( .A(n2259), .B(n2260), .Z(n2239) );
  XOR U2360 ( .A(n2261), .B(n2262), .Z(out[101]) );
  XNOR U2361 ( .A(n2233), .B(n2263), .Z(n2262) );
  XOR U2362 ( .A(n2249), .B(n17), .Z(n2263) );
  XOR U2363 ( .A(n2264), .B(n2251), .Z(n2249) );
  NANDN U2364 ( .A(n2265), .B(n2266), .Z(n2251) );
  AND U2365 ( .A(n2267), .B(n2268), .Z(n2264) );
  XNOR U2366 ( .A(n2269), .B(n2270), .Z(n2233) );
  XNOR U2367 ( .A(n2271), .B(n2272), .Z(n2270) );
  NANDN U2368 ( .A(n2241), .B(n2273), .Z(n2272) );
  XOR U2369 ( .A(n2274), .B(n2275), .Z(n2261) );
  XNOR U2370 ( .A(key[101]), .B(n2245), .Z(n2275) );
  NANDN U2371 ( .A(n2276), .B(n2277), .Z(n2245) );
  AND U2372 ( .A(n2278), .B(n2279), .Z(n2274) );
  XOR U2373 ( .A(n17), .B(n2280), .Z(out[100]) );
  XNOR U2374 ( .A(key[100]), .B(n13), .Z(n2280) );
  XNOR U2375 ( .A(n12), .B(n19), .Z(n13) );
  XOR U2376 ( .A(n2281), .B(n2282), .Z(n19) );
  XOR U2377 ( .A(n2283), .B(n2271), .Z(n2282) );
  OR U2378 ( .A(n2259), .B(n2284), .Z(n2271) );
  XNOR U2379 ( .A(n2241), .B(n2285), .Z(n2259) );
  NOR U2380 ( .A(n2285), .B(n2286), .Z(n2283) );
  IV U2381 ( .A(n2236), .Z(n12) );
  XOR U2382 ( .A(n2281), .B(n2287), .Z(n2236) );
  XNOR U2383 ( .A(n2288), .B(n2289), .Z(n2287) );
  NAND U2384 ( .A(n2290), .B(n2278), .Z(n2289) );
  XOR U2385 ( .A(n2269), .B(n2291), .Z(n17) );
  XOR U2386 ( .A(n2292), .B(n2288), .Z(n2291) );
  NANDN U2387 ( .A(n2293), .B(n2277), .Z(n2288) );
  XNOR U2388 ( .A(n2247), .B(n2278), .Z(n2277) );
  NOR U2389 ( .A(n2294), .B(n2247), .Z(n2292) );
  XNOR U2390 ( .A(n2281), .B(n2295), .Z(n2269) );
  XNOR U2391 ( .A(n2296), .B(n2297), .Z(n2295) );
  OR U2392 ( .A(n2298), .B(n2253), .Z(n2297) );
  XOR U2393 ( .A(n2299), .B(n2296), .Z(n2281) );
  OR U2394 ( .A(n2265), .B(n2300), .Z(n2296) );
  XNOR U2395 ( .A(n2301), .B(n2253), .Z(n2265) );
  XOR U2396 ( .A(n2285), .B(n2278), .Z(n2253) );
  XNOR U2397 ( .A(n2302), .B(n2303), .Z(n2278) );
  NANDN U2398 ( .A(n2304), .B(n2305), .Z(n2303) );
  IV U2399 ( .A(n2257), .Z(n2285) );
  XOR U2400 ( .A(n2306), .B(n2307), .Z(n2257) );
  NANDN U2401 ( .A(n2304), .B(n2308), .Z(n2307) );
  AND U2402 ( .A(n2268), .B(n2309), .Z(n2299) );
  IV U2403 ( .A(n2301), .Z(n2268) );
  XNOR U2404 ( .A(n2247), .B(n2241), .Z(n2301) );
  XOR U2405 ( .A(n2310), .B(n2306), .Z(n2241) );
  NANDN U2406 ( .A(n2311), .B(n2312), .Z(n2306) );
  AND U2407 ( .A(n2313), .B(n2314), .Z(n2310) );
  ANDN U2408 ( .B(n2316), .A(n2311), .Z(n2302) );
  XOR U2409 ( .A(n2317), .B(n2318), .Z(n2304) );
  XNOR U2410 ( .A(n2320), .B(n2321), .Z(n2317) );
  XNOR U2411 ( .A(n2322), .B(n2323), .Z(n2321) );
  AND U2412 ( .A(n2324), .B(n2313), .Z(n2322) );
  AND U2413 ( .A(n2324), .B(n2314), .Z(n2315) );
  XOR U2414 ( .A(n2320), .B(n2325), .Z(n2314) );
  XOR U2415 ( .A(n2326), .B(n2323), .Z(n2325) );
  NAND U2416 ( .A(n2312), .B(n2316), .Z(n2323) );
  XOR U2417 ( .A(n2305), .B(n2324), .Z(n2316) );
  XOR U2418 ( .A(n2308), .B(n2313), .Z(n2312) );
  XNOR U2419 ( .A(n2327), .B(n2328), .Z(n2313) );
  XOR U2420 ( .A(n2329), .B(n2330), .Z(n2328) );
  XNOR U2421 ( .A(n2331), .B(n2332), .Z(n2327) );
  ANDN U2422 ( .B(n2248), .A(n2294), .Z(n2331) );
  AND U2423 ( .A(n2305), .B(n2308), .Z(n2326) );
  XNOR U2424 ( .A(n2305), .B(n2308), .Z(n2320) );
  XNOR U2425 ( .A(n2333), .B(n2334), .Z(n2308) );
  XNOR U2426 ( .A(n2335), .B(n2336), .Z(n2334) );
  XOR U2427 ( .A(n2329), .B(n2337), .Z(n2333) );
  XNOR U2428 ( .A(n2338), .B(n2332), .Z(n2337) );
  OR U2429 ( .A(n2276), .B(n2293), .Z(n2332) );
  XNOR U2430 ( .A(n2294), .B(n2339), .Z(n2293) );
  XOR U2431 ( .A(n2248), .B(n2340), .Z(n2276) );
  AND U2432 ( .A(n2279), .B(n2290), .Z(n2338) );
  XNOR U2433 ( .A(n2341), .B(n2342), .Z(n2305) );
  XOR U2434 ( .A(n2343), .B(n2344), .Z(n2342) );
  XNOR U2435 ( .A(n2242), .B(n2329), .Z(n2344) );
  XNOR U2436 ( .A(n2294), .B(n2248), .Z(n2329) );
  XOR U2437 ( .A(n2273), .B(n2345), .Z(n2341) );
  XNOR U2438 ( .A(n2346), .B(n2347), .Z(n2345) );
  ANDN U2439 ( .B(n2258), .A(n2286), .Z(n2346) );
  IV U2440 ( .A(n2319), .Z(n2324) );
  XOR U2441 ( .A(n2348), .B(n2349), .Z(n2319) );
  XNOR U2442 ( .A(n2330), .B(n2350), .Z(n2349) );
  XOR U2443 ( .A(n2258), .B(n2336), .Z(n2350) );
  XNOR U2444 ( .A(n2339), .B(n2340), .Z(n2336) );
  IV U2445 ( .A(n2279), .Z(n2340) );
  XOR U2446 ( .A(n2343), .B(n2351), .Z(n2330) );
  XNOR U2447 ( .A(n2352), .B(n2353), .Z(n2351) );
  NANDN U2448 ( .A(n2298), .B(n2254), .Z(n2353) );
  IV U2449 ( .A(n2335), .Z(n2343) );
  XOR U2450 ( .A(n2354), .B(n2352), .Z(n2335) );
  NANDN U2451 ( .A(n2300), .B(n2266), .Z(n2352) );
  XOR U2452 ( .A(n2258), .B(n2279), .Z(n2254) );
  XOR U2453 ( .A(n2355), .B(n2356), .Z(n2279) );
  XOR U2454 ( .A(n2357), .B(n2358), .Z(n2356) );
  XNOR U2455 ( .A(n2339), .B(n2286), .Z(n2298) );
  IV U2456 ( .A(n2290), .Z(n2339) );
  AND U2457 ( .A(n2267), .B(n2309), .Z(n2354) );
  XOR U2458 ( .A(n2359), .B(n2294), .Z(n2309) );
  XOR U2459 ( .A(n2360), .B(n2361), .Z(n2294) );
  XNOR U2460 ( .A(n2357), .B(n2362), .Z(n2361) );
  XNOR U2461 ( .A(n2363), .B(n2248), .Z(n2267) );
  XNOR U2462 ( .A(n2286), .B(n2364), .Z(n2348) );
  XNOR U2463 ( .A(n2365), .B(n2347), .Z(n2364) );
  OR U2464 ( .A(n2260), .B(n2284), .Z(n2347) );
  XOR U2465 ( .A(n2273), .B(n2286), .Z(n2284) );
  XNOR U2466 ( .A(n2242), .B(n2258), .Z(n2260) );
  XOR U2467 ( .A(n2362), .B(n2358), .Z(n2366) );
  XOR U2468 ( .A(state[2]), .B(key[2]), .Z(n2362) );
  XNOR U2469 ( .A(n2367), .B(n2368), .Z(n2248) );
  AND U2470 ( .A(n2242), .B(n2273), .Z(n2365) );
  IV U2471 ( .A(n2363), .Z(n2242) );
  XOR U2472 ( .A(n2369), .B(n2368), .Z(n2363) );
  XOR U2473 ( .A(n2357), .B(n2355), .Z(n2368) );
  XNOR U2474 ( .A(state[5]), .B(key[5]), .Z(n2355) );
  XOR U2475 ( .A(n2359), .B(n2370), .Z(n2357) );
  XNOR U2476 ( .A(state[6]), .B(key[6]), .Z(n2370) );
  XOR U2477 ( .A(n2371), .B(n2372), .Z(n2286) );
  XNOR U2478 ( .A(n2369), .B(n2367), .Z(n2372) );
  XOR U2479 ( .A(state[7]), .B(key[7]), .Z(n2367) );
  XOR U2480 ( .A(state[4]), .B(key[4]), .Z(n2369) );
  XOR U2481 ( .A(n2273), .B(n2360), .Z(n2371) );
  XOR U2482 ( .A(n2358), .B(n2373), .Z(n2360) );
  XNOR U2483 ( .A(state[3]), .B(key[3]), .Z(n2373) );
  XNOR U2484 ( .A(state[1]), .B(key[1]), .Z(n2358) );
  IV U2485 ( .A(n2359), .Z(n2273) );
  XNOR U2486 ( .A(state[0]), .B(key[0]), .Z(n2359) );
  XNOR U2487 ( .A(n679), .B(n2374), .Z(out[0]) );
  XOR U2488 ( .A(key[0]), .B(n1301), .Z(n2374) );
  XNOR U2489 ( .A(n1494), .B(n2375), .Z(n1301) );
  XOR U2490 ( .A(n2376), .B(n684), .Z(n2375) );
  OR U2491 ( .A(n2377), .B(n1487), .Z(n684) );
  XNOR U2492 ( .A(n686), .B(n2378), .Z(n1487) );
  AND U2493 ( .A(n2379), .B(n1485), .Z(n2376) );
  XNOR U2494 ( .A(n682), .B(n2380), .Z(n679) );
  XOR U2495 ( .A(n2381), .B(n1496), .Z(n2380) );
  OR U2496 ( .A(n2382), .B(n1133), .Z(n1496) );
  XNOR U2497 ( .A(n1136), .B(n692), .Z(n1133) );
  NOR U2498 ( .A(n2383), .B(n1136), .Z(n2381) );
  XNOR U2499 ( .A(n1494), .B(n2384), .Z(n682) );
  XNOR U2500 ( .A(n2385), .B(n2386), .Z(n2384) );
  NANDN U2501 ( .A(n1481), .B(n2387), .Z(n2386) );
  XOR U2502 ( .A(n2388), .B(n2385), .Z(n1494) );
  OR U2503 ( .A(n1490), .B(n2389), .Z(n2385) );
  XOR U2504 ( .A(n1492), .B(n1481), .Z(n1490) );
  XNOR U2505 ( .A(n2378), .B(n692), .Z(n1481) );
  XOR U2506 ( .A(n2390), .B(n2391), .Z(n692) );
  NANDN U2507 ( .A(n2392), .B(n2393), .Z(n2391) );
  IV U2508 ( .A(n1485), .Z(n2378) );
  XOR U2509 ( .A(n2394), .B(n2395), .Z(n1485) );
  NANDN U2510 ( .A(n2392), .B(n2396), .Z(n2395) );
  ANDN U2511 ( .B(n1492), .A(n2397), .Z(n2388) );
  XOR U2512 ( .A(n1136), .B(n686), .Z(n1492) );
  XOR U2513 ( .A(n2398), .B(n2394), .Z(n686) );
  NANDN U2514 ( .A(n2399), .B(n2400), .Z(n2394) );
  AND U2515 ( .A(n2401), .B(n2402), .Z(n2398) );
  ANDN U2516 ( .B(n2404), .A(n2399), .Z(n2390) );
  XOR U2517 ( .A(n2405), .B(n2406), .Z(n2392) );
  XNOR U2518 ( .A(n2408), .B(n2409), .Z(n2405) );
  XNOR U2519 ( .A(n2410), .B(n2411), .Z(n2409) );
  AND U2520 ( .A(n2412), .B(n2401), .Z(n2410) );
  AND U2521 ( .A(n2412), .B(n2402), .Z(n2403) );
  XOR U2522 ( .A(n2408), .B(n2413), .Z(n2402) );
  XOR U2523 ( .A(n2414), .B(n2411), .Z(n2413) );
  NAND U2524 ( .A(n2400), .B(n2404), .Z(n2411) );
  XOR U2525 ( .A(n2393), .B(n2412), .Z(n2404) );
  XOR U2526 ( .A(n2396), .B(n2401), .Z(n2400) );
  XNOR U2527 ( .A(n2415), .B(n2416), .Z(n2401) );
  XOR U2528 ( .A(n2417), .B(n2418), .Z(n2416) );
  XNOR U2529 ( .A(n2419), .B(n2420), .Z(n2415) );
  ANDN U2530 ( .B(n1135), .A(n2383), .Z(n2419) );
  AND U2531 ( .A(n2393), .B(n2396), .Z(n2414) );
  XNOR U2532 ( .A(n2393), .B(n2396), .Z(n2408) );
  XNOR U2533 ( .A(n2421), .B(n2422), .Z(n2396) );
  XOR U2534 ( .A(n2423), .B(n2424), .Z(n2422) );
  XOR U2535 ( .A(n2417), .B(n2425), .Z(n2421) );
  XNOR U2536 ( .A(n2426), .B(n2420), .Z(n2425) );
  OR U2537 ( .A(n1134), .B(n2382), .Z(n2420) );
  XOR U2538 ( .A(n2383), .B(n1498), .Z(n2382) );
  XOR U2539 ( .A(n2427), .B(n691), .Z(n1134) );
  AND U2540 ( .A(n691), .B(n1498), .Z(n2426) );
  XNOR U2541 ( .A(n2428), .B(n2429), .Z(n2393) );
  XOR U2542 ( .A(n2430), .B(n2431), .Z(n2429) );
  XNOR U2543 ( .A(n1477), .B(n2417), .Z(n2431) );
  XNOR U2544 ( .A(n2383), .B(n1135), .Z(n2417) );
  XOR U2545 ( .A(n687), .B(n2432), .Z(n2428) );
  XNOR U2546 ( .A(n2433), .B(n2434), .Z(n2432) );
  AND U2547 ( .A(n1486), .B(n2379), .Z(n2433) );
  IV U2548 ( .A(n2407), .Z(n2412) );
  XOR U2549 ( .A(n2435), .B(n2436), .Z(n2407) );
  XNOR U2550 ( .A(n2418), .B(n2437), .Z(n2436) );
  XNOR U2551 ( .A(n1486), .B(n2424), .Z(n2437) );
  XOR U2552 ( .A(n2430), .B(n2438), .Z(n2418) );
  XNOR U2553 ( .A(n2439), .B(n2440), .Z(n2438) );
  NAND U2554 ( .A(n1482), .B(n2387), .Z(n2440) );
  IV U2555 ( .A(n2423), .Z(n2430) );
  XOR U2556 ( .A(n2441), .B(n2439), .Z(n2423) );
  NANDN U2557 ( .A(n2389), .B(n1491), .Z(n2439) );
  XOR U2558 ( .A(n1486), .B(n691), .Z(n1482) );
  XOR U2559 ( .A(n2442), .B(n2443), .Z(n691) );
  XOR U2560 ( .A(n2444), .B(n2445), .Z(n2443) );
  XOR U2561 ( .A(n2397), .B(n2387), .Z(n2389) );
  ANDN U2562 ( .B(n1493), .A(n2397), .Z(n2441) );
  XNOR U2563 ( .A(n2446), .B(n2383), .Z(n2397) );
  XNOR U2564 ( .A(n2447), .B(n2448), .Z(n2383) );
  XOR U2565 ( .A(n2449), .B(n2444), .Z(n2447) );
  XOR U2566 ( .A(n2379), .B(n2450), .Z(n2435) );
  XNOR U2567 ( .A(n2451), .B(n2434), .Z(n2450) );
  OR U2568 ( .A(n1488), .B(n2377), .Z(n2434) );
  XNOR U2569 ( .A(n687), .B(n2379), .Z(n2377) );
  XNOR U2570 ( .A(n1477), .B(n1486), .Z(n1488) );
  XOR U2571 ( .A(n2427), .B(n2452), .Z(n1486) );
  XOR U2572 ( .A(state[34]), .B(key[34]), .Z(n2448) );
  IV U2573 ( .A(n1135), .Z(n2427) );
  XOR U2574 ( .A(n2442), .B(n2453), .Z(n1135) );
  XNOR U2575 ( .A(n2444), .B(n2454), .Z(n2453) );
  AND U2576 ( .A(n687), .B(n1477), .Z(n2451) );
  XOR U2577 ( .A(n2442), .B(n2455), .Z(n1477) );
  XNOR U2578 ( .A(n2444), .B(n2456), .Z(n2455) );
  XOR U2579 ( .A(n2446), .B(n2457), .Z(n2444) );
  XNOR U2580 ( .A(state[38]), .B(key[38]), .Z(n2457) );
  XNOR U2581 ( .A(state[37]), .B(key[37]), .Z(n2442) );
  XNOR U2582 ( .A(n2458), .B(n2459), .Z(n2379) );
  XNOR U2583 ( .A(n2456), .B(n2454), .Z(n2459) );
  XOR U2584 ( .A(state[39]), .B(key[39]), .Z(n2454) );
  XOR U2585 ( .A(state[36]), .B(key[36]), .Z(n2456) );
  XOR U2586 ( .A(n687), .B(n2449), .Z(n2458) );
  XOR U2587 ( .A(n2445), .B(n2460), .Z(n2449) );
  XNOR U2588 ( .A(state[35]), .B(key[35]), .Z(n2460) );
  XNOR U2589 ( .A(state[33]), .B(key[33]), .Z(n2445) );
  IV U2590 ( .A(n2446), .Z(n687) );
  XNOR U2591 ( .A(state[32]), .B(key[32]), .Z(n2446) );
endmodule

