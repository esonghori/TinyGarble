
module compare_N16384_CC512 ( clk, rst, x, y, g, e );
  input [31:0] x;
  input [31:0] y;
  input clk, rst;
  output g, e;
  wire   ebreg, n4, n5, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169;

  DFF ebreg_reg ( .D(n5), .CLK(clk), .RST(rst), .Q(ebreg) );
  DFF greg_reg ( .D(n4), .CLK(clk), .RST(rst), .Q(g) );
  IV U10 ( .A(ebreg), .Z(e) );
  XNOR U11 ( .A(y[23]), .B(x[23]), .Z(n9) );
  NANDN U12 ( .A(x[22]), .B(y[22]), .Z(n8) );
  NAND U13 ( .A(n9), .B(n8), .Z(n139) );
  XNOR U14 ( .A(y[17]), .B(x[17]), .Z(n11) );
  NANDN U15 ( .A(x[16]), .B(y[16]), .Z(n10) );
  NAND U16 ( .A(n11), .B(n10), .Z(n121) );
  NOR U17 ( .A(n139), .B(n121), .Z(n17) );
  XNOR U18 ( .A(y[21]), .B(x[21]), .Z(n13) );
  NANDN U19 ( .A(x[20]), .B(y[20]), .Z(n12) );
  NAND U20 ( .A(n13), .B(n12), .Z(n133) );
  XNOR U21 ( .A(y[19]), .B(x[19]), .Z(n15) );
  NANDN U22 ( .A(x[18]), .B(y[18]), .Z(n14) );
  NAND U23 ( .A(n15), .B(n14), .Z(n127) );
  NOR U24 ( .A(n133), .B(n127), .Z(n16) );
  AND U25 ( .A(n17), .B(n16), .Z(n70) );
  XNOR U26 ( .A(y[11]), .B(x[11]), .Z(n19) );
  NANDN U27 ( .A(x[10]), .B(y[10]), .Z(n18) );
  NAND U28 ( .A(n19), .B(n18), .Z(n105) );
  XNOR U29 ( .A(y[5]), .B(x[5]), .Z(n21) );
  NANDN U30 ( .A(x[4]), .B(y[4]), .Z(n20) );
  NAND U31 ( .A(n21), .B(n20), .Z(n93) );
  NOR U32 ( .A(n105), .B(n93), .Z(n27) );
  XNOR U33 ( .A(y[9]), .B(x[9]), .Z(n23) );
  NANDN U34 ( .A(x[8]), .B(y[8]), .Z(n22) );
  NAND U35 ( .A(n23), .B(n22), .Z(n101) );
  XNOR U36 ( .A(y[7]), .B(x[7]), .Z(n25) );
  NANDN U37 ( .A(x[6]), .B(y[6]), .Z(n24) );
  NAND U38 ( .A(n25), .B(n24), .Z(n97) );
  NOR U39 ( .A(n101), .B(n97), .Z(n26) );
  AND U40 ( .A(n27), .B(n26), .Z(n39) );
  XNOR U41 ( .A(y[31]), .B(x[31]), .Z(n29) );
  NANDN U42 ( .A(x[30]), .B(y[30]), .Z(n28) );
  NAND U43 ( .A(n29), .B(n28), .Z(n163) );
  XNOR U44 ( .A(y[25]), .B(x[25]), .Z(n31) );
  NANDN U45 ( .A(x[24]), .B(y[24]), .Z(n30) );
  NAND U46 ( .A(n31), .B(n30), .Z(n145) );
  NOR U47 ( .A(n163), .B(n145), .Z(n37) );
  XNOR U48 ( .A(y[29]), .B(x[29]), .Z(n33) );
  NANDN U49 ( .A(x[28]), .B(y[28]), .Z(n32) );
  NAND U50 ( .A(n33), .B(n32), .Z(n157) );
  XNOR U51 ( .A(y[27]), .B(x[27]), .Z(n35) );
  NANDN U52 ( .A(x[26]), .B(y[26]), .Z(n34) );
  NAND U53 ( .A(n35), .B(n34), .Z(n151) );
  NOR U54 ( .A(n157), .B(n151), .Z(n36) );
  AND U55 ( .A(n37), .B(n36), .Z(n38) );
  AND U56 ( .A(n39), .B(n38), .Z(n68) );
  XNOR U57 ( .A(y[1]), .B(x[1]), .Z(n41) );
  NANDN U58 ( .A(x[0]), .B(y[0]), .Z(n40) );
  AND U59 ( .A(n41), .B(n40), .Z(n44) );
  XNOR U60 ( .A(y[13]), .B(x[13]), .Z(n43) );
  NANDN U61 ( .A(x[12]), .B(y[12]), .Z(n42) );
  NAND U62 ( .A(n43), .B(n42), .Z(n108) );
  ANDN U63 ( .B(n44), .A(n108), .Z(n50) );
  XNOR U64 ( .A(x[3]), .B(y[3]), .Z(n46) );
  NANDN U65 ( .A(x[2]), .B(y[2]), .Z(n45) );
  NAND U66 ( .A(n46), .B(n45), .Z(n89) );
  XNOR U67 ( .A(y[15]), .B(x[15]), .Z(n48) );
  NANDN U68 ( .A(x[14]), .B(y[14]), .Z(n47) );
  NAND U69 ( .A(n48), .B(n47), .Z(n115) );
  NOR U70 ( .A(n89), .B(n115), .Z(n49) );
  AND U71 ( .A(n50), .B(n49), .Z(n66) );
  ANDN U72 ( .B(x[30]), .A(y[30]), .Z(n159) );
  ANDN U73 ( .B(x[24]), .A(y[24]), .Z(n141) );
  NOR U74 ( .A(n159), .B(n141), .Z(n52) );
  ANDN U75 ( .B(x[28]), .A(y[28]), .Z(n153) );
  ANDN U76 ( .B(x[26]), .A(y[26]), .Z(n147) );
  NOR U77 ( .A(n153), .B(n147), .Z(n51) );
  AND U78 ( .A(n52), .B(n51), .Z(n56) );
  ANDN U79 ( .B(x[6]), .A(y[6]), .Z(n78) );
  ANDN U80 ( .B(x[4]), .A(y[4]), .Z(n80) );
  NOR U81 ( .A(n78), .B(n80), .Z(n54) );
  NANDN U82 ( .A(y[0]), .B(x[0]), .Z(n82) );
  ANDN U83 ( .B(x[2]), .A(y[2]), .Z(n86) );
  ANDN U84 ( .B(n82), .A(n86), .Z(n53) );
  AND U85 ( .A(n54), .B(n53), .Z(n55) );
  AND U86 ( .A(n56), .B(n55), .Z(n64) );
  ANDN U87 ( .B(x[22]), .A(y[22]), .Z(n135) );
  ANDN U88 ( .B(x[16]), .A(y[16]), .Z(n119) );
  NOR U89 ( .A(n135), .B(n119), .Z(n58) );
  ANDN U90 ( .B(x[20]), .A(y[20]), .Z(n129) );
  ANDN U91 ( .B(x[18]), .A(y[18]), .Z(n123) );
  NOR U92 ( .A(n129), .B(n123), .Z(n57) );
  AND U93 ( .A(n58), .B(n57), .Z(n62) );
  ANDN U94 ( .B(x[14]), .A(y[14]), .Z(n113) );
  ANDN U95 ( .B(x[8]), .A(y[8]), .Z(n76) );
  NOR U96 ( .A(n113), .B(n76), .Z(n60) );
  ANDN U97 ( .B(x[12]), .A(y[12]), .Z(n72) );
  ANDN U98 ( .B(x[10]), .A(y[10]), .Z(n74) );
  NOR U99 ( .A(n72), .B(n74), .Z(n59) );
  AND U100 ( .A(n60), .B(n59), .Z(n61) );
  AND U101 ( .A(n62), .B(n61), .Z(n63) );
  AND U102 ( .A(n64), .B(n63), .Z(n65) );
  AND U103 ( .A(n66), .B(n65), .Z(n67) );
  AND U104 ( .A(n68), .B(n67), .Z(n69) );
  AND U105 ( .A(n70), .B(n69), .Z(n71) );
  NAND U106 ( .A(e), .B(n71), .Z(n5) );
  NANDN U107 ( .A(n71), .B(e), .Z(n167) );
  ANDN U108 ( .B(x[31]), .A(y[31]), .Z(n165) );
  ANDN U109 ( .B(x[15]), .A(y[15]), .Z(n117) );
  NANDN U110 ( .A(y[13]), .B(x[13]), .Z(n111) );
  NANDN U111 ( .A(y[11]), .B(x[11]), .Z(n73) );
  ANDN U112 ( .B(n73), .A(n72), .Z(n107) );
  NANDN U113 ( .A(y[9]), .B(x[9]), .Z(n75) );
  ANDN U114 ( .B(n75), .A(n74), .Z(n103) );
  NANDN U115 ( .A(y[7]), .B(x[7]), .Z(n77) );
  ANDN U116 ( .B(n77), .A(n76), .Z(n99) );
  NANDN U117 ( .A(y[5]), .B(x[5]), .Z(n79) );
  ANDN U118 ( .B(n79), .A(n78), .Z(n95) );
  NANDN U119 ( .A(y[3]), .B(x[3]), .Z(n81) );
  ANDN U120 ( .B(n81), .A(n80), .Z(n91) );
  NANDN U121 ( .A(x[1]), .B(n82), .Z(n85) );
  XNOR U122 ( .A(n82), .B(x[1]), .Z(n83) );
  NAND U123 ( .A(n83), .B(y[1]), .Z(n84) );
  NAND U124 ( .A(n85), .B(n84), .Z(n87) );
  ANDN U125 ( .B(n87), .A(n86), .Z(n88) );
  OR U126 ( .A(n89), .B(n88), .Z(n90) );
  AND U127 ( .A(n91), .B(n90), .Z(n92) );
  OR U128 ( .A(n93), .B(n92), .Z(n94) );
  AND U129 ( .A(n95), .B(n94), .Z(n96) );
  OR U130 ( .A(n97), .B(n96), .Z(n98) );
  AND U131 ( .A(n99), .B(n98), .Z(n100) );
  OR U132 ( .A(n101), .B(n100), .Z(n102) );
  AND U133 ( .A(n103), .B(n102), .Z(n104) );
  OR U134 ( .A(n105), .B(n104), .Z(n106) );
  AND U135 ( .A(n107), .B(n106), .Z(n109) );
  OR U136 ( .A(n109), .B(n108), .Z(n110) );
  AND U137 ( .A(n111), .B(n110), .Z(n112) );
  NANDN U138 ( .A(n113), .B(n112), .Z(n114) );
  NANDN U139 ( .A(n115), .B(n114), .Z(n116) );
  NANDN U140 ( .A(n117), .B(n116), .Z(n118) );
  OR U141 ( .A(n119), .B(n118), .Z(n120) );
  NANDN U142 ( .A(n121), .B(n120), .Z(n122) );
  NANDN U143 ( .A(n123), .B(n122), .Z(n125) );
  ANDN U144 ( .B(x[17]), .A(y[17]), .Z(n124) );
  OR U145 ( .A(n125), .B(n124), .Z(n126) );
  NANDN U146 ( .A(n127), .B(n126), .Z(n128) );
  NANDN U147 ( .A(n129), .B(n128), .Z(n131) );
  ANDN U148 ( .B(x[19]), .A(y[19]), .Z(n130) );
  OR U149 ( .A(n131), .B(n130), .Z(n132) );
  NANDN U150 ( .A(n133), .B(n132), .Z(n134) );
  NANDN U151 ( .A(n135), .B(n134), .Z(n137) );
  ANDN U152 ( .B(x[21]), .A(y[21]), .Z(n136) );
  OR U153 ( .A(n137), .B(n136), .Z(n138) );
  NANDN U154 ( .A(n139), .B(n138), .Z(n140) );
  NANDN U155 ( .A(n141), .B(n140), .Z(n143) );
  ANDN U156 ( .B(x[23]), .A(y[23]), .Z(n142) );
  OR U157 ( .A(n143), .B(n142), .Z(n144) );
  NANDN U158 ( .A(n145), .B(n144), .Z(n146) );
  NANDN U159 ( .A(n147), .B(n146), .Z(n149) );
  ANDN U160 ( .B(x[25]), .A(y[25]), .Z(n148) );
  OR U161 ( .A(n149), .B(n148), .Z(n150) );
  NANDN U162 ( .A(n151), .B(n150), .Z(n152) );
  NANDN U163 ( .A(n153), .B(n152), .Z(n155) );
  ANDN U164 ( .B(x[27]), .A(y[27]), .Z(n154) );
  OR U165 ( .A(n155), .B(n154), .Z(n156) );
  NANDN U166 ( .A(n157), .B(n156), .Z(n158) );
  NANDN U167 ( .A(n159), .B(n158), .Z(n161) );
  ANDN U168 ( .B(x[29]), .A(y[29]), .Z(n160) );
  OR U169 ( .A(n161), .B(n160), .Z(n162) );
  NANDN U170 ( .A(n163), .B(n162), .Z(n164) );
  NANDN U171 ( .A(n165), .B(n164), .Z(n166) );
  NANDN U172 ( .A(n167), .B(n166), .Z(n169) );
  NAND U173 ( .A(n167), .B(g), .Z(n168) );
  NAND U174 ( .A(n169), .B(n168), .Z(n4) );
endmodule

