
module mult_N64_CC1 ( clk, rst, a, b, c );
  input [63:0] a;
  input [63:0] b;
  output [127:0] c;
  input clk, rst;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
         n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
         n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345,
         n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
         n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
         n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369,
         n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
         n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
         n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
         n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
         n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
         n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417,
         n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
         n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
         n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441,
         n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
         n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
         n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
         n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
         n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
         n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489,
         n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
         n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
         n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
         n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537,
         n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
         n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
         n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561,
         n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569,
         n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
         n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585,
         n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593,
         n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601,
         n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609,
         n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617,
         n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625,
         n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633,
         n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
         n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
         n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657,
         n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665,
         n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673,
         n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681,
         n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
         n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697,
         n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705,
         n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
         n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
         n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729,
         n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737,
         n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745,
         n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753,
         n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761,
         n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769,
         n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777,
         n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785,
         n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
         n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801,
         n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809,
         n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817,
         n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825,
         n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833,
         n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841,
         n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849,
         n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857,
         n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865,
         n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873,
         n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881,
         n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889,
         n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897,
         n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905,
         n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913,
         n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921,
         n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929,
         n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
         n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945,
         n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953,
         n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961,
         n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969,
         n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977,
         n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985,
         n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993,
         n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001,
         n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
         n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017,
         n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025,
         n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
         n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041,
         n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049,
         n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057,
         n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065,
         n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073,
         n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
         n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089,
         n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097,
         n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
         n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113,
         n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121,
         n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129,
         n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137,
         n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145,
         n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153,
         n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161,
         n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169,
         n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
         n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185,
         n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193,
         n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201,
         n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209,
         n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217,
         n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225,
         n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233,
         n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241,
         n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249,
         n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257,
         n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265,
         n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273,
         n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281,
         n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289,
         n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297,
         n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305,
         n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313,
         n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321,
         n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329,
         n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337,
         n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345,
         n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353,
         n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361,
         n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369,
         n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377,
         n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385,
         n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393,
         n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401,
         n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409,
         n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417,
         n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425,
         n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433,
         n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441,
         n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449,
         n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457,
         n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465,
         n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473,
         n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481,
         n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489,
         n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497,
         n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505,
         n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513,
         n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521,
         n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529,
         n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537,
         n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545,
         n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553,
         n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561,
         n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569,
         n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577,
         n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585,
         n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593,
         n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601,
         n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609,
         n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617,
         n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625,
         n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633,
         n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641,
         n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649,
         n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657,
         n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665,
         n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673,
         n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681,
         n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689,
         n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697,
         n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705,
         n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713,
         n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721,
         n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729,
         n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737,
         n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745,
         n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753,
         n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761,
         n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769,
         n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777,
         n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785,
         n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793,
         n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801,
         n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809,
         n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817,
         n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825,
         n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833,
         n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841,
         n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849,
         n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857,
         n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865,
         n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873,
         n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881,
         n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889,
         n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897,
         n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905,
         n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913,
         n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921,
         n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929,
         n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937,
         n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945,
         n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953,
         n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961,
         n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969,
         n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977,
         n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985,
         n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993,
         n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001,
         n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009,
         n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017,
         n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025,
         n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033,
         n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041,
         n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049,
         n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057,
         n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065,
         n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073,
         n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081,
         n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089,
         n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097,
         n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105,
         n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113,
         n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121,
         n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129,
         n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137,
         n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145,
         n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153,
         n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161,
         n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169,
         n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177,
         n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185,
         n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193,
         n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201,
         n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209,
         n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217,
         n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225,
         n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233,
         n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241,
         n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249,
         n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257,
         n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265,
         n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273,
         n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281,
         n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289,
         n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297,
         n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305,
         n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313,
         n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321,
         n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329,
         n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337,
         n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345,
         n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353,
         n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361,
         n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369,
         n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377,
         n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385,
         n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393,
         n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401,
         n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409,
         n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417,
         n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425,
         n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433,
         n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441,
         n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449,
         n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457,
         n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465,
         n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473,
         n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481,
         n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489,
         n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497,
         n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505,
         n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513,
         n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521,
         n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529,
         n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537,
         n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545,
         n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553,
         n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561,
         n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569,
         n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577,
         n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585,
         n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593,
         n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601,
         n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609,
         n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617,
         n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625,
         n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633,
         n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641,
         n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649,
         n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657,
         n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665,
         n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673,
         n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681,
         n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689,
         n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697,
         n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705,
         n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713,
         n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721,
         n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729,
         n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737,
         n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745,
         n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753,
         n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761,
         n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769,
         n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777,
         n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785,
         n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793,
         n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801,
         n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809,
         n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817,
         n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825,
         n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833,
         n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841,
         n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849,
         n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857,
         n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865,
         n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873,
         n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881,
         n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889,
         n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897,
         n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905,
         n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913,
         n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921,
         n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929,
         n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937,
         n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945,
         n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953,
         n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961,
         n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969,
         n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977,
         n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985,
         n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993,
         n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001,
         n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009,
         n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017,
         n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025,
         n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033,
         n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041,
         n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049,
         n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057,
         n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065,
         n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073,
         n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081,
         n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089,
         n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097,
         n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105,
         n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113,
         n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121,
         n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129,
         n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137,
         n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145,
         n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153,
         n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161,
         n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169,
         n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177,
         n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185,
         n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193,
         n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201,
         n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209,
         n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217,
         n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225,
         n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233,
         n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241,
         n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249,
         n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257,
         n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265,
         n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273,
         n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281,
         n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289,
         n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297,
         n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305,
         n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313,
         n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321,
         n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329,
         n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337,
         n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345,
         n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353,
         n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361,
         n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369,
         n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377,
         n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385,
         n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393,
         n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401,
         n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409,
         n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417,
         n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425,
         n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433,
         n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441,
         n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449,
         n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457,
         n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465,
         n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473,
         n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481,
         n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489,
         n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497,
         n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505,
         n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513,
         n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521,
         n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529,
         n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537,
         n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545,
         n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553,
         n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561,
         n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569,
         n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577,
         n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585,
         n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593,
         n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601,
         n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609,
         n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617,
         n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625,
         n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633,
         n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641,
         n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649,
         n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657,
         n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665,
         n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673,
         n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681,
         n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689,
         n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697,
         n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705,
         n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713,
         n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721,
         n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729,
         n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737,
         n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745,
         n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753,
         n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761,
         n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769,
         n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777,
         n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785,
         n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793,
         n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801,
         n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809,
         n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817,
         n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825,
         n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833,
         n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841,
         n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849,
         n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857,
         n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865,
         n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873,
         n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881,
         n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889,
         n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897,
         n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905,
         n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913,
         n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921,
         n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929,
         n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937,
         n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945,
         n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953,
         n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961,
         n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969,
         n24970, n24971, n24972;

  XNOR U2 ( .A(n6149), .B(n6150), .Z(n6426) );
  XNOR U3 ( .A(n8448), .B(n8449), .Z(n8451) );
  XNOR U4 ( .A(n9147), .B(n9148), .Z(n9150) );
  NAND U5 ( .A(n11080), .B(n11083), .Z(n2) );
  XOR U6 ( .A(n11080), .B(n11083), .Z(n3) );
  NANDN U7 ( .A(n11081), .B(n3), .Z(n4) );
  NAND U8 ( .A(n2), .B(n4), .Z(n10782) );
  NAND U9 ( .A(n11534), .B(n11537), .Z(n5) );
  XOR U10 ( .A(n11534), .B(n11537), .Z(n6) );
  NANDN U11 ( .A(n11535), .B(n6), .Z(n7) );
  NAND U12 ( .A(n5), .B(n7), .Z(n11124) );
  XOR U13 ( .A(n12246), .B(n12248), .Z(n8) );
  NANDN U14 ( .A(n12247), .B(n8), .Z(n9) );
  NAND U15 ( .A(n12246), .B(n12248), .Z(n10) );
  AND U16 ( .A(n9), .B(n10), .Z(n11837) );
  NAND U17 ( .A(n12219), .B(n12222), .Z(n11) );
  XOR U18 ( .A(n12219), .B(n12222), .Z(n12) );
  NANDN U19 ( .A(n12220), .B(n12), .Z(n13) );
  NAND U20 ( .A(n11), .B(n13), .Z(n11812) );
  NAND U21 ( .A(n12547), .B(n12550), .Z(n14) );
  XOR U22 ( .A(n12547), .B(n12550), .Z(n15) );
  NANDN U23 ( .A(n12548), .B(n15), .Z(n16) );
  NAND U24 ( .A(n14), .B(n16), .Z(n12245) );
  NAND U25 ( .A(n13159), .B(n13162), .Z(n17) );
  XOR U26 ( .A(n13159), .B(n13162), .Z(n18) );
  NANDN U27 ( .A(n13160), .B(n18), .Z(n19) );
  NAND U28 ( .A(n17), .B(n19), .Z(n12929) );
  XOR U29 ( .A(n13866), .B(n13868), .Z(n20) );
  NANDN U30 ( .A(n13867), .B(n20), .Z(n21) );
  NAND U31 ( .A(n13866), .B(n13868), .Z(n22) );
  AND U32 ( .A(n21), .B(n22), .Z(n13517) );
  NAND U33 ( .A(n13848), .B(n13851), .Z(n23) );
  XOR U34 ( .A(n13848), .B(n13851), .Z(n24) );
  NANDN U35 ( .A(n13849), .B(n24), .Z(n25) );
  NAND U36 ( .A(n23), .B(n25), .Z(n13499) );
  NAND U37 ( .A(n14233), .B(n14236), .Z(n26) );
  XOR U38 ( .A(n14233), .B(n14236), .Z(n27) );
  NANDN U39 ( .A(n14234), .B(n27), .Z(n28) );
  NAND U40 ( .A(n26), .B(n28), .Z(n13865) );
  NAND U41 ( .A(n14254), .B(n14256), .Z(n29) );
  XOR U42 ( .A(n14254), .B(n14256), .Z(n30) );
  NANDN U43 ( .A(n14253), .B(n30), .Z(n31) );
  NAND U44 ( .A(n29), .B(n31), .Z(n13890) );
  NAND U45 ( .A(n14940), .B(n14943), .Z(n32) );
  XOR U46 ( .A(n14940), .B(n14943), .Z(n33) );
  NANDN U47 ( .A(n14941), .B(n33), .Z(n34) );
  NAND U48 ( .A(n32), .B(n34), .Z(n14568) );
  NAND U49 ( .A(n14776), .B(n14779), .Z(n35) );
  XOR U50 ( .A(n14776), .B(n14779), .Z(n36) );
  NAND U51 ( .A(n36), .B(n14777), .Z(n37) );
  NAND U52 ( .A(n35), .B(n37), .Z(n14873) );
  NANDN U53 ( .A(n15994), .B(n15996), .Z(n38) );
  OR U54 ( .A(n15996), .B(n15667), .Z(n39) );
  NANDN U55 ( .A(n15993), .B(n39), .Z(n40) );
  NAND U56 ( .A(n38), .B(n40), .Z(n15669) );
  XOR U57 ( .A(n16362), .B(n16360), .Z(n41) );
  NANDN U58 ( .A(n16359), .B(n41), .Z(n42) );
  NAND U59 ( .A(n16362), .B(n16360), .Z(n43) );
  AND U60 ( .A(n42), .B(n43), .Z(n15998) );
  XOR U61 ( .A(n15787), .B(n15788), .Z(n44) );
  NANDN U62 ( .A(n15790), .B(n44), .Z(n45) );
  NAND U63 ( .A(n15787), .B(n15788), .Z(n46) );
  AND U64 ( .A(n45), .B(n46), .Z(n15914) );
  NAND U65 ( .A(n17392), .B(n17395), .Z(n47) );
  XOR U66 ( .A(n17392), .B(n17395), .Z(n48) );
  NANDN U67 ( .A(n17393), .B(n48), .Z(n49) );
  NAND U68 ( .A(n47), .B(n49), .Z(n17062) );
  NAND U69 ( .A(n18059), .B(n18062), .Z(n50) );
  XOR U70 ( .A(n18059), .B(n18062), .Z(n51) );
  NANDN U71 ( .A(n18060), .B(n51), .Z(n52) );
  NAND U72 ( .A(n50), .B(n52), .Z(n17743) );
  XOR U73 ( .A(n20173), .B(n20172), .Z(n53) );
  NANDN U74 ( .A(n20175), .B(n53), .Z(n54) );
  NAND U75 ( .A(n20173), .B(n20172), .Z(n55) );
  AND U76 ( .A(n54), .B(n55), .Z(n20425) );
  NAND U77 ( .A(n22728), .B(n22727), .Z(n56) );
  NAND U78 ( .A(n22725), .B(n22726), .Z(n57) );
  NAND U79 ( .A(n56), .B(n57), .Z(n22870) );
  NAND U80 ( .A(n18792), .B(n18793), .Z(n58) );
  NAND U81 ( .A(n18473), .B(n18474), .Z(n59) );
  NAND U82 ( .A(n58), .B(n59), .Z(n18478) );
  NANDN U83 ( .A(n3885), .B(n3394), .Z(n60) );
  XNOR U84 ( .A(n3392), .B(n60), .Z(n61) );
  NANDN U85 ( .A(n3394), .B(n3393), .Z(n62) );
  NAND U86 ( .A(n61), .B(n62), .Z(n3648) );
  XNOR U87 ( .A(n4417), .B(n4418), .Z(n4693) );
  NANDN U88 ( .A(n6733), .B(n6128), .Z(n63) );
  XNOR U89 ( .A(n6126), .B(n63), .Z(n64) );
  NANDN U90 ( .A(n6128), .B(n6127), .Z(n65) );
  NAND U91 ( .A(n64), .B(n65), .Z(n6432) );
  XNOR U92 ( .A(n6462), .B(n6463), .Z(n6726) );
  XNOR U93 ( .A(n4182), .B(n4183), .Z(n4406) );
  XNOR U94 ( .A(n4445), .B(n4446), .Z(n4677) );
  XNOR U95 ( .A(n5272), .B(n5273), .Z(n5526) );
  XNOR U96 ( .A(n6452), .B(n6453), .Z(n6729) );
  XNOR U97 ( .A(n7074), .B(n7075), .Z(n7077) );
  XNOR U98 ( .A(n6185), .B(n6186), .Z(n6422) );
  XNOR U99 ( .A(n5599), .B(n5600), .Z(n5813) );
  NANDN U100 ( .A(n8390), .B(n7729), .Z(n66) );
  XNOR U101 ( .A(n7727), .B(n66), .Z(n67) );
  NANDN U102 ( .A(n7729), .B(n7728), .Z(n68) );
  NAND U103 ( .A(n67), .B(n68), .Z(n8065) );
  XNOR U104 ( .A(n7784), .B(n7785), .Z(n8047) );
  XNOR U105 ( .A(n8127), .B(n8128), .Z(n8377) );
  XNOR U106 ( .A(n7457), .B(n7458), .Z(n7711) );
  XNOR U107 ( .A(n6504), .B(n6505), .Z(n6809) );
  XNOR U108 ( .A(n8464), .B(n8465), .Z(n8826) );
  XNOR U109 ( .A(n8450), .B(n8451), .Z(n8739) );
  NANDN U110 ( .A(n9431), .B(n8752), .Z(n69) );
  XNOR U111 ( .A(n8750), .B(n69), .Z(n70) );
  NANDN U112 ( .A(n8752), .B(n8751), .Z(n71) );
  NAND U113 ( .A(n70), .B(n71), .Z(n9055) );
  XNOR U114 ( .A(n8807), .B(n8808), .Z(n9116) );
  XNOR U115 ( .A(n9455), .B(n9456), .Z(n9458) );
  XNOR U116 ( .A(n9093), .B(n9094), .Z(n9419) );
  XNOR U117 ( .A(n9157), .B(n9158), .Z(n9160) );
  NAND U118 ( .A(n9892), .B(n9894), .Z(n72) );
  XOR U119 ( .A(n9892), .B(n9894), .Z(n73) );
  NANDN U120 ( .A(n9893), .B(n73), .Z(n74) );
  NAND U121 ( .A(n72), .B(n74), .Z(n9528) );
  XNOR U122 ( .A(n9818), .B(n9819), .Z(n10325) );
  XNOR U123 ( .A(n9499), .B(n9500), .Z(n9770) );
  XNOR U124 ( .A(n10300), .B(n10301), .Z(n10303) );
  XNOR U125 ( .A(n9800), .B(n9801), .Z(n10306) );
  XNOR U126 ( .A(n9854), .B(n9855), .Z(n10360) );
  NAND U127 ( .A(n11041), .B(n11044), .Z(n75) );
  XOR U128 ( .A(n11041), .B(n11044), .Z(n76) );
  NANDN U129 ( .A(n11042), .B(n76), .Z(n77) );
  NAND U130 ( .A(n75), .B(n77), .Z(n10762) );
  XNOR U131 ( .A(n10356), .B(n10357), .Z(n10785) );
  XOR U132 ( .A(n9767), .B(n9768), .Z(n78) );
  NANDN U133 ( .A(n9769), .B(n78), .Z(n79) );
  NAND U134 ( .A(n9767), .B(n9768), .Z(n80) );
  AND U135 ( .A(n79), .B(n80), .Z(n9542) );
  NAND U136 ( .A(n11463), .B(n11466), .Z(n81) );
  XOR U137 ( .A(n11463), .B(n11466), .Z(n82) );
  NANDN U138 ( .A(n11464), .B(n82), .Z(n83) );
  NAND U139 ( .A(n81), .B(n83), .Z(n11027) );
  XOR U140 ( .A(n11071), .B(n11069), .Z(n84) );
  NANDN U141 ( .A(n11070), .B(n84), .Z(n85) );
  NAND U142 ( .A(n11071), .B(n11069), .Z(n86) );
  AND U143 ( .A(n85), .B(n86), .Z(n10779) );
  XOR U144 ( .A(n11770), .B(n11772), .Z(n87) );
  NANDN U145 ( .A(n11771), .B(n87), .Z(n88) );
  NAND U146 ( .A(n11770), .B(n11772), .Z(n89) );
  AND U147 ( .A(n88), .B(n89), .Z(n11483) );
  NAND U148 ( .A(n11794), .B(n11797), .Z(n90) );
  XOR U149 ( .A(n11794), .B(n11797), .Z(n91) );
  NANDN U150 ( .A(n11795), .B(n91), .Z(n92) );
  NAND U151 ( .A(n90), .B(n92), .Z(n11498) );
  XNOR U152 ( .A(n11139), .B(n11140), .Z(n11407) );
  XNOR U153 ( .A(n11734), .B(n11735), .Z(n11737) );
  NAND U154 ( .A(n11847), .B(n11846), .Z(n93) );
  XOR U155 ( .A(n11847), .B(n11846), .Z(n94) );
  NANDN U156 ( .A(n11845), .B(n94), .Z(n95) );
  NAND U157 ( .A(n93), .B(n95), .Z(n11543) );
  XNOR U158 ( .A(n11811), .B(n11812), .Z(n12227) );
  NANDN U159 ( .A(n12558), .B(n12560), .Z(n96) );
  OR U160 ( .A(n12560), .B(n12253), .Z(n97) );
  NANDN U161 ( .A(n12557), .B(n97), .Z(n98) );
  NAND U162 ( .A(n96), .B(n98), .Z(n12257) );
  NAND U163 ( .A(n12948), .B(n12946), .Z(n99) );
  XOR U164 ( .A(n12948), .B(n12946), .Z(n100) );
  NANDN U165 ( .A(n12947), .B(n100), .Z(n101) );
  NAND U166 ( .A(n99), .B(n101), .Z(n12562) );
  XNOR U167 ( .A(n13084), .B(n13085), .Z(n13087) );
  XOR U168 ( .A(n12900), .B(n12901), .Z(n102) );
  NANDN U169 ( .A(n12902), .B(n102), .Z(n103) );
  NAND U170 ( .A(n12900), .B(n12901), .Z(n104) );
  AND U171 ( .A(n103), .B(n104), .Z(n12509) );
  XNOR U172 ( .A(n2988), .B(n2987), .Z(n2979) );
  XOR U173 ( .A(n13126), .B(n13128), .Z(n105) );
  NANDN U174 ( .A(n13127), .B(n105), .Z(n106) );
  NAND U175 ( .A(n13126), .B(n13128), .Z(n107) );
  AND U176 ( .A(n106), .B(n107), .Z(n12903) );
  XOR U177 ( .A(n13141), .B(n13143), .Z(n108) );
  NANDN U178 ( .A(n13142), .B(n108), .Z(n109) );
  NAND U179 ( .A(n13141), .B(n13143), .Z(n110) );
  AND U180 ( .A(n109), .B(n110), .Z(n12914) );
  NAND U181 ( .A(n12962), .B(n12961), .Z(n111) );
  XOR U182 ( .A(n12962), .B(n12961), .Z(n112) );
  NANDN U183 ( .A(n12963), .B(n112), .Z(n113) );
  NAND U184 ( .A(n111), .B(n113), .Z(n12576) );
  XNOR U185 ( .A(n13413), .B(n13414), .Z(n13726) );
  NAND U186 ( .A(n13509), .B(n13511), .Z(n114) );
  XOR U187 ( .A(n13509), .B(n13511), .Z(n115) );
  NANDN U188 ( .A(n13508), .B(n115), .Z(n116) );
  NAND U189 ( .A(n114), .B(n116), .Z(n13177) );
  XNOR U190 ( .A(n14118), .B(n14119), .Z(n14121) );
  XNOR U191 ( .A(n12931), .B(n12932), .Z(n117) );
  XNOR U192 ( .A(n12930), .B(n117), .Z(n13168) );
  NANDN U193 ( .A(n13844), .B(n13489), .Z(n118) );
  NAND U194 ( .A(n13844), .B(n13845), .Z(n119) );
  NANDN U195 ( .A(n13843), .B(n119), .Z(n120) );
  NAND U196 ( .A(n118), .B(n120), .Z(n13495) );
  XNOR U197 ( .A(n14132), .B(n14133), .Z(n14411) );
  NANDN U198 ( .A(n13857), .B(n13859), .Z(n121) );
  OR U199 ( .A(n13859), .B(n13507), .Z(n122) );
  NANDN U200 ( .A(n13856), .B(n122), .Z(n123) );
  NAND U201 ( .A(n121), .B(n123), .Z(n13513) );
  XNOR U202 ( .A(n13864), .B(n13865), .Z(n14076) );
  XOR U203 ( .A(n14565), .B(n14566), .Z(n124) );
  XNOR U204 ( .A(n14564), .B(n124), .Z(n14949) );
  XNOR U205 ( .A(n14156), .B(n14157), .Z(n14478) );
  NAND U206 ( .A(n14528), .B(n14527), .Z(n125) );
  XOR U207 ( .A(n14528), .B(n14527), .Z(n126) );
  NANDN U208 ( .A(n14529), .B(n126), .Z(n127) );
  NAND U209 ( .A(n125), .B(n127), .Z(n14214) );
  NAND U210 ( .A(n14551), .B(n14554), .Z(n128) );
  XOR U211 ( .A(n14551), .B(n14554), .Z(n129) );
  NANDN U212 ( .A(n14552), .B(n129), .Z(n130) );
  NAND U213 ( .A(n128), .B(n130), .Z(n14238) );
  NAND U214 ( .A(n14571), .B(n14574), .Z(n131) );
  XOR U215 ( .A(n14571), .B(n14574), .Z(n132) );
  NANDN U216 ( .A(n14572), .B(n132), .Z(n133) );
  NAND U217 ( .A(n131), .B(n133), .Z(n14260) );
  NAND U218 ( .A(n14270), .B(n14273), .Z(n134) );
  XOR U219 ( .A(n14270), .B(n14273), .Z(n135) );
  NANDN U220 ( .A(n14271), .B(n135), .Z(n136) );
  NAND U221 ( .A(n134), .B(n136), .Z(n13902) );
  XNOR U222 ( .A(n14462), .B(n14463), .Z(n14836) );
  NANDN U223 ( .A(n15948), .B(n15613), .Z(n137) );
  NAND U224 ( .A(n15948), .B(n15949), .Z(n138) );
  NANDN U225 ( .A(n15947), .B(n138), .Z(n139) );
  NAND U226 ( .A(n137), .B(n139), .Z(n15619) );
  NANDN U227 ( .A(n15979), .B(n15648), .Z(n140) );
  NAND U228 ( .A(n15979), .B(n15980), .Z(n141) );
  NANDN U229 ( .A(n15978), .B(n141), .Z(n142) );
  NAND U230 ( .A(n140), .B(n142), .Z(n15650) );
  NAND U231 ( .A(n15196), .B(n15197), .Z(n143) );
  XOR U232 ( .A(n15196), .B(n15197), .Z(n144) );
  NANDN U233 ( .A(n15195), .B(n144), .Z(n145) );
  NAND U234 ( .A(n143), .B(n145), .Z(n15097) );
  NAND U235 ( .A(n16340), .B(n16343), .Z(n146) );
  XOR U236 ( .A(n16340), .B(n16343), .Z(n147) );
  NANDN U237 ( .A(n16341), .B(n147), .Z(n148) );
  NAND U238 ( .A(n146), .B(n148), .Z(n15977) );
  NAND U239 ( .A(n16647), .B(n16649), .Z(n149) );
  XOR U240 ( .A(n16647), .B(n16649), .Z(n150) );
  NANDN U241 ( .A(n16648), .B(n150), .Z(n151) );
  NAND U242 ( .A(n149), .B(n151), .Z(n16319) );
  XNOR U243 ( .A(n15997), .B(n15998), .Z(n16368) );
  XOR U244 ( .A(n15671), .B(n15672), .Z(n152) );
  XNOR U245 ( .A(n15670), .B(n152), .Z(n15771) );
  XNOR U246 ( .A(n4362), .B(n4363), .Z(n4627) );
  NAND U247 ( .A(n16615), .B(n16618), .Z(n153) );
  XOR U248 ( .A(n16615), .B(n16618), .Z(n154) );
  NANDN U249 ( .A(n16616), .B(n154), .Z(n155) );
  NAND U250 ( .A(n153), .B(n155), .Z(n16279) );
  XOR U251 ( .A(n16280), .B(n16282), .Z(n156) );
  NANDN U252 ( .A(n16281), .B(n156), .Z(n157) );
  NAND U253 ( .A(n16280), .B(n16282), .Z(n158) );
  AND U254 ( .A(n157), .B(n158), .Z(n16152) );
  XOR U255 ( .A(n18067), .B(n18068), .Z(n159) );
  NANDN U256 ( .A(n18069), .B(n159), .Z(n160) );
  NAND U257 ( .A(n18067), .B(n18068), .Z(n161) );
  AND U258 ( .A(n160), .B(n161), .Z(n17749) );
  XNOR U259 ( .A(n17059), .B(n17058), .Z(n162) );
  XNOR U260 ( .A(n17060), .B(n162), .Z(n17157) );
  NAND U261 ( .A(n18415), .B(n18418), .Z(n163) );
  XOR U262 ( .A(n18415), .B(n18418), .Z(n164) );
  NANDN U263 ( .A(n18416), .B(n164), .Z(n165) );
  NAND U264 ( .A(n163), .B(n165), .Z(n18071) );
  XNOR U265 ( .A(n5470), .B(n5471), .Z(n5764) );
  XOR U266 ( .A(n17850), .B(n17851), .Z(n166) );
  NANDN U267 ( .A(n17853), .B(n166), .Z(n167) );
  NAND U268 ( .A(n17850), .B(n17851), .Z(n168) );
  AND U269 ( .A(n167), .B(n168), .Z(n18049) );
  XOR U270 ( .A(n18199), .B(n18198), .Z(n169) );
  NANDN U271 ( .A(n18201), .B(n169), .Z(n170) );
  NAND U272 ( .A(n18199), .B(n18198), .Z(n171) );
  AND U273 ( .A(n170), .B(n171), .Z(n18394) );
  NAND U274 ( .A(n19085), .B(n19087), .Z(n172) );
  XOR U275 ( .A(n19085), .B(n19087), .Z(n173) );
  NANDN U276 ( .A(n19084), .B(n173), .Z(n174) );
  NAND U277 ( .A(n172), .B(n174), .Z(n18746) );
  NANDN U278 ( .A(n18448), .B(n18771), .Z(n175) );
  OR U279 ( .A(n18771), .B(n18770), .Z(n176) );
  NANDN U280 ( .A(n18773), .B(n176), .Z(n177) );
  NAND U281 ( .A(n175), .B(n177), .Z(n18452) );
  XOR U282 ( .A(n19753), .B(n19752), .Z(n178) );
  NANDN U283 ( .A(n19755), .B(n178), .Z(n179) );
  NAND U284 ( .A(n19753), .B(n19752), .Z(n180) );
  AND U285 ( .A(n179), .B(n180), .Z(n19762) );
  NAND U286 ( .A(n18780), .B(n18781), .Z(n181) );
  NAND U287 ( .A(n18462), .B(n18461), .Z(n182) );
  NAND U288 ( .A(n181), .B(n182), .Z(n18466) );
  XNOR U289 ( .A(n20890), .B(n20891), .Z(n20893) );
  XOR U290 ( .A(n20489), .B(n20490), .Z(n183) );
  NANDN U291 ( .A(n20492), .B(n183), .Z(n184) );
  NAND U292 ( .A(n20489), .B(n20490), .Z(n185) );
  AND U293 ( .A(n184), .B(n185), .Z(n20756) );
  NAND U294 ( .A(n19459), .B(n19460), .Z(n186) );
  NAND U295 ( .A(n19141), .B(n19140), .Z(n187) );
  NAND U296 ( .A(n186), .B(n187), .Z(n19145) );
  NAND U297 ( .A(n9363), .B(n9364), .Z(n188) );
  NANDN U298 ( .A(n9388), .B(n9387), .Z(n189) );
  NAND U299 ( .A(n188), .B(n189), .Z(n9367) );
  NAND U300 ( .A(n22873), .B(n22872), .Z(n190) );
  NAND U301 ( .A(n22871), .B(n22870), .Z(n191) );
  NAND U302 ( .A(n190), .B(n191), .Z(n22999) );
  XNOR U303 ( .A(n21222), .B(n21223), .Z(n21225) );
  NAND U304 ( .A(n18797), .B(n18796), .Z(n192) );
  NAND U305 ( .A(n18477), .B(n18478), .Z(n193) );
  NAND U306 ( .A(n192), .B(n193), .Z(n18801) );
  XNOR U307 ( .A(n9377), .B(n9378), .Z(n9380) );
  NAND U308 ( .A(n22724), .B(n22723), .Z(n194) );
  NAND U309 ( .A(n22721), .B(n22722), .Z(n195) );
  NAND U310 ( .A(n194), .B(n195), .Z(n22862) );
  NAND U311 ( .A(n19153), .B(n19152), .Z(n196) );
  NAND U312 ( .A(n18807), .B(n18806), .Z(n197) );
  AND U313 ( .A(n196), .B(n197), .Z(n18808) );
  XOR U314 ( .A(n13696), .B(n13695), .Z(n13689) );
  NANDN U315 ( .A(n4411), .B(n3886), .Z(n198) );
  XNOR U316 ( .A(n3884), .B(n198), .Z(n199) );
  NANDN U317 ( .A(n3886), .B(n3885), .Z(n200) );
  NAND U318 ( .A(n199), .B(n200), .Z(n4152) );
  NANDN U319 ( .A(n5531), .B(n4952), .Z(n201) );
  XNOR U320 ( .A(n4950), .B(n201), .Z(n202) );
  NANDN U321 ( .A(n4952), .B(n4951), .Z(n203) );
  NAND U322 ( .A(n202), .B(n203), .Z(n5242) );
  XNOR U323 ( .A(n4154), .B(n4155), .Z(n4422) );
  XNOR U324 ( .A(n5244), .B(n5245), .Z(n5542) );
  XNOR U325 ( .A(n3403), .B(n3404), .Z(n3406) );
  XNOR U326 ( .A(n4694), .B(n4695), .Z(n4970) );
  XNOR U327 ( .A(n6438), .B(n6439), .Z(n6441) );
  XNOR U328 ( .A(n3641), .B(n3642), .Z(n3673) );
  XNOR U329 ( .A(n3417), .B(n3418), .Z(n3677) );
  XNOR U330 ( .A(n6145), .B(n6146), .Z(n6450) );
  XNOR U331 ( .A(n3917), .B(n3918), .Z(n4143) );
  XNOR U332 ( .A(n6460), .B(n6461), .Z(n6727) );
  XNOR U333 ( .A(n6159), .B(n6160), .Z(n6423) );
  XNOR U334 ( .A(n4180), .B(n4181), .Z(n4407) );
  XNOR U335 ( .A(n4443), .B(n4444), .Z(n4678) );
  XNOR U336 ( .A(n4716), .B(n4717), .Z(n4946) );
  XNOR U337 ( .A(n4985), .B(n4986), .Z(n5233) );
  XNOR U338 ( .A(n5270), .B(n5271), .Z(n5527) );
  XNOR U339 ( .A(n5565), .B(n5566), .Z(n5823) );
  XNOR U340 ( .A(n5862), .B(n5863), .Z(n6120) );
  XNOR U341 ( .A(n6765), .B(n6766), .Z(n7055) );
  XNOR U342 ( .A(n7057), .B(n7058), .Z(n7060) );
  XNOR U343 ( .A(n7407), .B(n7408), .Z(n7410) );
  XNOR U344 ( .A(n5003), .B(n5004), .Z(n5006) );
  XNOR U345 ( .A(n4736), .B(n4737), .Z(n5010) );
  XNOR U346 ( .A(n5585), .B(n5586), .Z(n5588) );
  XNOR U347 ( .A(n7397), .B(n7398), .Z(n7739) );
  XNOR U348 ( .A(n7386), .B(n7387), .Z(n7720) );
  XNOR U349 ( .A(n7126), .B(n7127), .Z(n7373) );
  XNOR U350 ( .A(n6795), .B(n6796), .Z(n7052) );
  XNOR U351 ( .A(n6494), .B(n6495), .Z(n6721) );
  XNOR U352 ( .A(n7746), .B(n7747), .Z(n8083) );
  XNOR U353 ( .A(n7431), .B(n7432), .Z(n7773) );
  XNOR U354 ( .A(n8056), .B(n8057), .Z(n8384) );
  XNOR U355 ( .A(n7774), .B(n7775), .Z(n8048) );
  XNOR U356 ( .A(n8042), .B(n8043), .Z(n8045) );
  XNOR U357 ( .A(n7136), .B(n7137), .Z(n7370) );
  XNOR U358 ( .A(n6502), .B(n6503), .Z(n6810) );
  XNOR U359 ( .A(n6199), .B(n6200), .Z(n6417) );
  XNOR U360 ( .A(n8079), .B(n8080), .Z(n8412) );
  XNOR U361 ( .A(n8400), .B(n8401), .Z(n8403) );
  XNOR U362 ( .A(n8101), .B(n8102), .Z(n8439) );
  XNOR U363 ( .A(n8131), .B(n8132), .Z(n8473) );
  XNOR U364 ( .A(n8385), .B(n8386), .Z(n8423) );
  XNOR U365 ( .A(n8115), .B(n8116), .Z(n8382) );
  XNOR U366 ( .A(n8119), .B(n8120), .Z(n8380) );
  XNOR U367 ( .A(n8135), .B(n8136), .Z(n8138) );
  XNOR U368 ( .A(n8761), .B(n8762), .Z(n8764) );
  XOR U369 ( .A(n9429), .B(n9430), .Z(n204) );
  NANDN U370 ( .A(n9432), .B(n9431), .Z(n205) );
  NAND U371 ( .A(n204), .B(n205), .Z(n9780) );
  XOR U372 ( .A(n9043), .B(n9044), .Z(n9105) );
  XNOR U373 ( .A(n8817), .B(n8818), .Z(n9127) );
  XNOR U374 ( .A(n9109), .B(n9110), .Z(n9112) );
  XOR U375 ( .A(n9137), .B(n9138), .Z(n9140) );
  XNOR U376 ( .A(n9457), .B(n9458), .Z(n9811) );
  XNOR U377 ( .A(n9115), .B(n9116), .Z(n9118) );
  XNOR U378 ( .A(n9149), .B(n9150), .Z(n9412) );
  XNOR U379 ( .A(n9788), .B(n9789), .Z(n10294) );
  XNOR U380 ( .A(n9417), .B(n9418), .Z(n9480) );
  XNOR U381 ( .A(n9159), .B(n9160), .Z(n9410) );
  XNOR U382 ( .A(n9521), .B(n9522), .Z(n9886) );
  XNOR U383 ( .A(n10290), .B(n10291), .Z(n10721) );
  XNOR U384 ( .A(n8855), .B(n8856), .Z(n9034) );
  XNOR U385 ( .A(n9798), .B(n9799), .Z(n10307) );
  XNOR U386 ( .A(n10320), .B(n10321), .Z(n10765) );
  XNOR U387 ( .A(n11002), .B(n11003), .Z(n11005) );
  XNOR U388 ( .A(n11435), .B(n11436), .Z(n11438) );
  XNOR U389 ( .A(n10362), .B(n10363), .Z(n10789) );
  XNOR U390 ( .A(n9864), .B(n9865), .Z(n10375) );
  XOR U391 ( .A(n9768), .B(n9769), .Z(n206) );
  XNOR U392 ( .A(n9767), .B(n206), .Z(n10423) );
  XNOR U393 ( .A(n9541), .B(n9542), .Z(n9918) );
  XNOR U394 ( .A(n11716), .B(n11717), .Z(n11719) );
  XNOR U395 ( .A(n12136), .B(n12137), .Z(n12139) );
  XNOR U396 ( .A(n10332), .B(n10333), .Z(n10770) );
  XNOR U397 ( .A(n10784), .B(n10785), .Z(n11089) );
  XNOR U398 ( .A(n10372), .B(n10373), .Z(n10713) );
  XNOR U399 ( .A(n10425), .B(n10426), .Z(n10826) );
  XNOR U400 ( .A(n12439), .B(n12440), .Z(n12442) );
  NANDN U401 ( .A(n11029), .B(n10755), .Z(n207) );
  NAND U402 ( .A(n11029), .B(n11030), .Z(n208) );
  NANDN U403 ( .A(n11028), .B(n208), .Z(n209) );
  NAND U404 ( .A(n207), .B(n209), .Z(n10759) );
  XNOR U405 ( .A(n11076), .B(n11077), .Z(n11501) );
  XNOR U406 ( .A(n12834), .B(n12835), .Z(n12837) );
  XNOR U407 ( .A(n11485), .B(n11486), .Z(n11774) );
  XOR U408 ( .A(n11838), .B(n11840), .Z(n210) );
  NANDN U409 ( .A(n11839), .B(n210), .Z(n211) );
  NAND U410 ( .A(n11838), .B(n11840), .Z(n212) );
  AND U411 ( .A(n211), .B(n212), .Z(n11538) );
  XNOR U412 ( .A(n11123), .B(n11124), .Z(n11409) );
  XNOR U413 ( .A(n11836), .B(n11837), .Z(n12251) );
  XNOR U414 ( .A(n13066), .B(n13067), .Z(n13069) );
  XNOR U415 ( .A(n11479), .B(n11480), .Z(n11764) );
  XNOR U416 ( .A(n11782), .B(n11783), .Z(n12200) );
  XNOR U417 ( .A(n11494), .B(n11495), .Z(n11786) );
  XNOR U418 ( .A(n13383), .B(n13384), .Z(n13386) );
  XNOR U419 ( .A(n12158), .B(n12159), .Z(n12161) );
  XNOR U420 ( .A(n12850), .B(n12851), .Z(n12853) );
  XOR U421 ( .A(n12499), .B(n12501), .Z(n213) );
  NANDN U422 ( .A(n12500), .B(n213), .Z(n214) );
  NAND U423 ( .A(n12499), .B(n12501), .Z(n215) );
  AND U424 ( .A(n214), .B(n215), .Z(n12196) );
  XOR U425 ( .A(n12517), .B(n12519), .Z(n216) );
  NANDN U426 ( .A(n12518), .B(n216), .Z(n217) );
  NAND U427 ( .A(n12517), .B(n12519), .Z(n218) );
  AND U428 ( .A(n217), .B(n218), .Z(n12212) );
  XNOR U429 ( .A(n11814), .B(n11815), .Z(n219) );
  XNOR U430 ( .A(n11813), .B(n219), .Z(n12228) );
  NAND U431 ( .A(n11854), .B(n11857), .Z(n220) );
  XOR U432 ( .A(n11854), .B(n11857), .Z(n221) );
  NANDN U433 ( .A(n11855), .B(n221), .Z(n222) );
  NAND U434 ( .A(n220), .B(n222), .Z(n11548) );
  NAND U435 ( .A(n12263), .B(n12261), .Z(n223) );
  XOR U436 ( .A(n12263), .B(n12261), .Z(n224) );
  NANDN U437 ( .A(n12262), .B(n224), .Z(n225) );
  NAND U438 ( .A(n223), .B(n225), .Z(n11859) );
  XNOR U439 ( .A(n13735), .B(n13736), .Z(n13738) );
  XNOR U440 ( .A(n12856), .B(n12857), .Z(n12859) );
  NAND U441 ( .A(n12541), .B(n12544), .Z(n226) );
  XOR U442 ( .A(n12541), .B(n12544), .Z(n227) );
  NANDN U443 ( .A(n12542), .B(n227), .Z(n228) );
  NAND U444 ( .A(n226), .B(n228), .Z(n12236) );
  NAND U445 ( .A(n12565), .B(n12568), .Z(n229) );
  XOR U446 ( .A(n12565), .B(n12568), .Z(n230) );
  NANDN U447 ( .A(n12566), .B(n230), .Z(n231) );
  NAND U448 ( .A(n229), .B(n231), .Z(n12264) );
  XNOR U449 ( .A(n13399), .B(n13400), .Z(n13402) );
  XNOR U450 ( .A(n12481), .B(n12482), .Z(n12880) );
  NAND U451 ( .A(n12894), .B(n12897), .Z(n232) );
  XOR U452 ( .A(n12894), .B(n12897), .Z(n233) );
  NANDN U453 ( .A(n12895), .B(n233), .Z(n234) );
  NAND U454 ( .A(n232), .B(n234), .Z(n12498) );
  NANDN U455 ( .A(n12908), .B(n12514), .Z(n235) );
  NAND U456 ( .A(n12908), .B(n12909), .Z(n236) );
  NANDN U457 ( .A(n12907), .B(n236), .Z(n237) );
  NAND U458 ( .A(n235), .B(n237), .Z(n12516) );
  XNOR U459 ( .A(n12530), .B(n12531), .Z(n12922) );
  NAND U460 ( .A(n13151), .B(n13154), .Z(n238) );
  XOR U461 ( .A(n13151), .B(n13154), .Z(n239) );
  NANDN U462 ( .A(n13152), .B(n239), .Z(n240) );
  NAND U463 ( .A(n238), .B(n240), .Z(n12924) );
  NAND U464 ( .A(n13178), .B(n13181), .Z(n241) );
  XOR U465 ( .A(n13178), .B(n13181), .Z(n242) );
  NANDN U466 ( .A(n13179), .B(n242), .Z(n243) );
  NAND U467 ( .A(n241), .B(n243), .Z(n12944) );
  NAND U468 ( .A(n12953), .B(n12956), .Z(n244) );
  XOR U469 ( .A(n12953), .B(n12956), .Z(n245) );
  NANDN U470 ( .A(n12954), .B(n245), .Z(n246) );
  NAND U471 ( .A(n244), .B(n246), .Z(n12570) );
  XNOR U472 ( .A(n12576), .B(n12577), .Z(n12804) );
  XNOR U473 ( .A(n2982), .B(n2981), .Z(n2975) );
  XNOR U474 ( .A(n3000), .B(n2999), .Z(n3003) );
  XNOR U475 ( .A(n13753), .B(n13754), .Z(n13756) );
  XNOR U476 ( .A(n13405), .B(n13406), .Z(n13408) );
  NAND U477 ( .A(n13135), .B(n13138), .Z(n247) );
  XOR U478 ( .A(n13135), .B(n13138), .Z(n248) );
  NANDN U479 ( .A(n13136), .B(n248), .Z(n249) );
  NAND U480 ( .A(n247), .B(n249), .Z(n12910) );
  NANDN U481 ( .A(n13483), .B(n13150), .Z(n250) );
  NAND U482 ( .A(n13483), .B(n13484), .Z(n251) );
  NANDN U483 ( .A(n13482), .B(n251), .Z(n252) );
  NAND U484 ( .A(n250), .B(n252), .Z(n13156) );
  XNOR U485 ( .A(n2951), .B(n2952), .Z(n3319) );
  XOR U486 ( .A(n13436), .B(n13438), .Z(n253) );
  NANDN U487 ( .A(n13437), .B(n253), .Z(n254) );
  NAND U488 ( .A(n13436), .B(n13438), .Z(n255) );
  AND U489 ( .A(n254), .B(n255), .Z(n13113) );
  NAND U490 ( .A(n13458), .B(n13461), .Z(n256) );
  XOR U491 ( .A(n13458), .B(n13461), .Z(n257) );
  NANDN U492 ( .A(n13459), .B(n257), .Z(n258) );
  NAND U493 ( .A(n256), .B(n258), .Z(n13130) );
  NAND U494 ( .A(n13501), .B(n13500), .Z(n259) );
  XOR U495 ( .A(n13501), .B(n13500), .Z(n260) );
  NANDN U496 ( .A(n13502), .B(n260), .Z(n261) );
  NAND U497 ( .A(n259), .B(n261), .Z(n13170) );
  NANDN U498 ( .A(n13524), .B(n13526), .Z(n262) );
  OR U499 ( .A(n13526), .B(n13194), .Z(n263) );
  NANDN U500 ( .A(n13523), .B(n263), .Z(n264) );
  NAND U501 ( .A(n262), .B(n264), .Z(n13200) );
  NAND U502 ( .A(n13878), .B(n13881), .Z(n265) );
  XOR U503 ( .A(n13878), .B(n13881), .Z(n266) );
  NANDN U504 ( .A(n13879), .B(n266), .Z(n267) );
  NAND U505 ( .A(n265), .B(n267), .Z(n13528) );
  XNOR U506 ( .A(n14444), .B(n14445), .Z(n14447) );
  NAND U507 ( .A(n13833), .B(n13836), .Z(n268) );
  XOR U508 ( .A(n13833), .B(n13836), .Z(n269) );
  NANDN U509 ( .A(n13834), .B(n269), .Z(n270) );
  NAND U510 ( .A(n268), .B(n270), .Z(n13480) );
  XNOR U511 ( .A(n3324), .B(n3325), .Z(n3567) );
  XNOR U512 ( .A(n3044), .B(n3043), .Z(n3055) );
  XNOR U513 ( .A(n13777), .B(n13778), .Z(n14148) );
  XNOR U514 ( .A(n14144), .B(n14145), .Z(n14466) );
  XOR U515 ( .A(n14173), .B(n14175), .Z(n271) );
  NAND U516 ( .A(n271), .B(n14174), .Z(n272) );
  NAND U517 ( .A(n14173), .B(n14175), .Z(n273) );
  AND U518 ( .A(n272), .B(n273), .Z(n13800) );
  XNOR U519 ( .A(n13498), .B(n13499), .Z(n13711) );
  NAND U520 ( .A(n14218), .B(n14221), .Z(n274) );
  XOR U521 ( .A(n14218), .B(n14221), .Z(n275) );
  NANDN U522 ( .A(n14219), .B(n275), .Z(n276) );
  NAND U523 ( .A(n274), .B(n276), .Z(n13853) );
  NAND U524 ( .A(n14535), .B(n14534), .Z(n277) );
  XOR U525 ( .A(n14535), .B(n14534), .Z(n278) );
  NANDN U526 ( .A(n14536), .B(n278), .Z(n279) );
  NAND U527 ( .A(n277), .B(n279), .Z(n14222) );
  XOR U528 ( .A(n13868), .B(n13867), .Z(n280) );
  XNOR U529 ( .A(n13866), .B(n280), .Z(n14077) );
  NANDN U530 ( .A(n14565), .B(n14250), .Z(n281) );
  NAND U531 ( .A(n14565), .B(n14566), .Z(n282) );
  NANDN U532 ( .A(n14564), .B(n282), .Z(n283) );
  NAND U533 ( .A(n281), .B(n283), .Z(n14252) );
  XOR U534 ( .A(n14261), .B(n14263), .Z(n284) );
  NANDN U535 ( .A(n14262), .B(n284), .Z(n285) );
  NAND U536 ( .A(n14261), .B(n14263), .Z(n286) );
  AND U537 ( .A(n285), .B(n286), .Z(n13898) );
  XNOR U538 ( .A(n14452), .B(n14453), .Z(n14824) );
  XNOR U539 ( .A(n14154), .B(n14155), .Z(n14479) );
  XOR U540 ( .A(n14933), .B(n14935), .Z(n287) );
  NANDN U541 ( .A(n14934), .B(n287), .Z(n288) );
  NAND U542 ( .A(n14933), .B(n14935), .Z(n289) );
  AND U543 ( .A(n288), .B(n289), .Z(n14561) );
  XNOR U544 ( .A(n4326), .B(n4327), .Z(n4594) );
  XNOR U545 ( .A(n4069), .B(n4070), .Z(n4330) );
  XNOR U546 ( .A(n3338), .B(n3339), .Z(n3580) );
  XNOR U547 ( .A(n14460), .B(n14461), .Z(n14837) );
  NAND U548 ( .A(n14909), .B(n14912), .Z(n290) );
  XOR U549 ( .A(n14909), .B(n14912), .Z(n291) );
  NANDN U550 ( .A(n14910), .B(n291), .Z(n292) );
  NAND U551 ( .A(n290), .B(n292), .Z(n14538) );
  XNOR U552 ( .A(n14259), .B(n14260), .Z(n14386) );
  XNOR U553 ( .A(n13901), .B(n13902), .Z(n14072) );
  NAND U554 ( .A(n13225), .B(n13226), .Z(n293) );
  NAND U555 ( .A(n12987), .B(n12986), .Z(n294) );
  NAND U556 ( .A(n293), .B(n294), .Z(n12991) );
  XNOR U557 ( .A(n3114), .B(n3113), .Z(n3119) );
  XNOR U558 ( .A(n14474), .B(n14475), .Z(n14848) );
  NAND U559 ( .A(n15290), .B(n15293), .Z(n295) );
  XOR U560 ( .A(n15290), .B(n15293), .Z(n296) );
  NANDN U561 ( .A(n15291), .B(n296), .Z(n297) );
  NAND U562 ( .A(n295), .B(n297), .Z(n14973) );
  NAND U563 ( .A(n15659), .B(n15662), .Z(n298) );
  XOR U564 ( .A(n15659), .B(n15662), .Z(n299) );
  NANDN U565 ( .A(n15660), .B(n299), .Z(n300) );
  NAND U566 ( .A(n298), .B(n300), .Z(n15289) );
  NAND U567 ( .A(n13240), .B(n13239), .Z(n301) );
  NAND U568 ( .A(n12994), .B(n12995), .Z(n302) );
  NAND U569 ( .A(n301), .B(n302), .Z(n13246) );
  XNOR U570 ( .A(n5153), .B(n5154), .Z(n5438) );
  XNOR U571 ( .A(n10155), .B(n10154), .Z(n10156) );
  XOR U572 ( .A(n15097), .B(n15098), .Z(n303) );
  NANDN U573 ( .A(n15100), .B(n303), .Z(n304) );
  NAND U574 ( .A(n15097), .B(n15098), .Z(n305) );
  AND U575 ( .A(n304), .B(n305), .Z(n15204) );
  NAND U576 ( .A(n15578), .B(n15581), .Z(n306) );
  XOR U577 ( .A(n15578), .B(n15581), .Z(n307) );
  NANDN U578 ( .A(n15579), .B(n307), .Z(n308) );
  NAND U579 ( .A(n306), .B(n308), .Z(n15459) );
  NAND U580 ( .A(n15937), .B(n15940), .Z(n309) );
  XOR U581 ( .A(n15937), .B(n15940), .Z(n310) );
  NANDN U582 ( .A(n15938), .B(n310), .Z(n311) );
  NAND U583 ( .A(n309), .B(n311), .Z(n15607) );
  NAND U584 ( .A(n16314), .B(n16317), .Z(n312) );
  XOR U585 ( .A(n16314), .B(n16317), .Z(n313) );
  NANDN U586 ( .A(n16315), .B(n313), .Z(n314) );
  NAND U587 ( .A(n312), .B(n314), .Z(n15957) );
  XOR U588 ( .A(n16347), .B(n16348), .Z(n315) );
  XNOR U589 ( .A(n16346), .B(n315), .Z(n16684) );
  XNOR U590 ( .A(n4617), .B(n4618), .Z(n4890) );
  NAND U591 ( .A(n17034), .B(n17037), .Z(n316) );
  XOR U592 ( .A(n17034), .B(n17037), .Z(n317) );
  NANDN U593 ( .A(n17035), .B(n317), .Z(n318) );
  NAND U594 ( .A(n316), .B(n318), .Z(n16673) );
  XOR U595 ( .A(n16372), .B(n16373), .Z(n319) );
  NANDN U596 ( .A(n16374), .B(n319), .Z(n320) );
  NAND U597 ( .A(n16372), .B(n16373), .Z(n321) );
  AND U598 ( .A(n320), .B(n321), .Z(n16006) );
  XNOR U599 ( .A(n4360), .B(n4361), .Z(n4628) );
  XNOR U600 ( .A(n4105), .B(n4106), .Z(n4366) );
  XNOR U601 ( .A(n16307), .B(n16308), .Z(n16479) );
  NAND U602 ( .A(n17386), .B(n17389), .Z(n322) );
  XOR U603 ( .A(n17386), .B(n17389), .Z(n323) );
  NANDN U604 ( .A(n17387), .B(n323), .Z(n324) );
  NAND U605 ( .A(n322), .B(n324), .Z(n17054) );
  NANDN U606 ( .A(n16698), .B(n16700), .Z(n325) );
  OR U607 ( .A(n16700), .B(n16369), .Z(n326) );
  NANDN U608 ( .A(n16697), .B(n326), .Z(n327) );
  NAND U609 ( .A(n325), .B(n327), .Z(n16370) );
  XNOR U610 ( .A(n6329), .B(n6330), .Z(n6375) );
  XNOR U611 ( .A(n16281), .B(n16282), .Z(n328) );
  XNOR U612 ( .A(n16280), .B(n328), .Z(n16490) );
  XOR U613 ( .A(n17744), .B(n17746), .Z(n329) );
  NANDN U614 ( .A(n17745), .B(n329), .Z(n330) );
  NAND U615 ( .A(n17744), .B(n17746), .Z(n331) );
  AND U616 ( .A(n330), .B(n331), .Z(n17385) );
  NAND U617 ( .A(n13260), .B(n13259), .Z(n332) );
  NAND U618 ( .A(n13002), .B(n13003), .Z(n333) );
  NAND U619 ( .A(n332), .B(n333), .Z(n13266) );
  XNOR U620 ( .A(n6335), .B(n6336), .Z(n6644) );
  NAND U621 ( .A(n16981), .B(n16983), .Z(n334) );
  XOR U622 ( .A(n16981), .B(n16983), .Z(n335) );
  NANDN U623 ( .A(n16982), .B(n335), .Z(n336) );
  NAND U624 ( .A(n334), .B(n336), .Z(n16990) );
  NAND U625 ( .A(n17400), .B(n17402), .Z(n337) );
  XOR U626 ( .A(n17400), .B(n17402), .Z(n338) );
  NANDN U627 ( .A(n17401), .B(n338), .Z(n339) );
  NAND U628 ( .A(n337), .B(n339), .Z(n17066) );
  XOR U629 ( .A(n17757), .B(n17759), .Z(n340) );
  NANDN U630 ( .A(n17758), .B(n340), .Z(n341) );
  NAND U631 ( .A(n17757), .B(n17759), .Z(n342) );
  AND U632 ( .A(n341), .B(n342), .Z(n17404) );
  NAND U633 ( .A(n17317), .B(n17320), .Z(n343) );
  XOR U634 ( .A(n17317), .B(n17320), .Z(n344) );
  NANDN U635 ( .A(n17318), .B(n344), .Z(n345) );
  NAND U636 ( .A(n343), .B(n345), .Z(n16984) );
  NAND U637 ( .A(n18052), .B(n18054), .Z(n346) );
  XOR U638 ( .A(n18052), .B(n18054), .Z(n347) );
  NANDN U639 ( .A(n18053), .B(n347), .Z(n348) );
  NAND U640 ( .A(n346), .B(n348), .Z(n17735) );
  XNOR U641 ( .A(n5189), .B(n5190), .Z(n5474) );
  NAND U642 ( .A(n18039), .B(n18042), .Z(n349) );
  XOR U643 ( .A(n18039), .B(n18042), .Z(n350) );
  NAND U644 ( .A(n350), .B(n18040), .Z(n351) );
  NAND U645 ( .A(n349), .B(n351), .Z(n17850) );
  NAND U646 ( .A(n18402), .B(n18401), .Z(n352) );
  XOR U647 ( .A(n18402), .B(n18401), .Z(n353) );
  NANDN U648 ( .A(n18400), .B(n353), .Z(n354) );
  NAND U649 ( .A(n352), .B(n354), .Z(n18056) );
  NAND U650 ( .A(n18734), .B(n18737), .Z(n355) );
  XOR U651 ( .A(n18734), .B(n18737), .Z(n356) );
  NANDN U652 ( .A(n18735), .B(n356), .Z(n357) );
  NAND U653 ( .A(n355), .B(n357), .Z(n18420) );
  NAND U654 ( .A(n18425), .B(n18428), .Z(n358) );
  XOR U655 ( .A(n18425), .B(n18428), .Z(n359) );
  NANDN U656 ( .A(n18426), .B(n359), .Z(n360) );
  NAND U657 ( .A(n358), .B(n360), .Z(n18079) );
  XNOR U658 ( .A(n7005), .B(n7006), .Z(n7289) );
  XNOR U659 ( .A(n5763), .B(n5764), .Z(n6060) );
  XOR U660 ( .A(n6353), .B(n6354), .Z(n6663) );
  NAND U661 ( .A(n17701), .B(n17704), .Z(n361) );
  XOR U662 ( .A(n17701), .B(n17704), .Z(n362) );
  NANDN U663 ( .A(n17702), .B(n362), .Z(n363) );
  NAND U664 ( .A(n361), .B(n363), .Z(n17534) );
  NANDN U665 ( .A(n18440), .B(n18763), .Z(n364) );
  OR U666 ( .A(n18763), .B(n18762), .Z(n365) );
  NANDN U667 ( .A(n18765), .B(n365), .Z(n366) );
  NAND U668 ( .A(n364), .B(n366), .Z(n18444) );
  NAND U669 ( .A(n13280), .B(n13279), .Z(n367) );
  NAND U670 ( .A(n13010), .B(n13011), .Z(n368) );
  NAND U671 ( .A(n367), .B(n368), .Z(n13286) );
  NANDN U672 ( .A(n19099), .B(n18751), .Z(n369) );
  NAND U673 ( .A(n19099), .B(n19100), .Z(n370) );
  NANDN U674 ( .A(n19098), .B(n370), .Z(n371) );
  NAND U675 ( .A(n369), .B(n371), .Z(n18757) );
  XOR U676 ( .A(n18098), .B(n18099), .Z(n18100) );
  XNOR U677 ( .A(n6981), .B(n6982), .Z(n7305) );
  NAND U678 ( .A(n18386), .B(n18388), .Z(n372) );
  XOR U679 ( .A(n18386), .B(n18388), .Z(n373) );
  NANDN U680 ( .A(n18387), .B(n373), .Z(n374) );
  NAND U681 ( .A(n372), .B(n374), .Z(n18199) );
  NAND U682 ( .A(n18693), .B(n18696), .Z(n375) );
  XOR U683 ( .A(n18693), .B(n18696), .Z(n376) );
  NANDN U684 ( .A(n18694), .B(n376), .Z(n377) );
  NAND U685 ( .A(n375), .B(n377), .Z(n18390) );
  XOR U686 ( .A(n18503), .B(n18504), .Z(n378) );
  NANDN U687 ( .A(n18506), .B(n378), .Z(n379) );
  NAND U688 ( .A(n18503), .B(n18504), .Z(n380) );
  AND U689 ( .A(n379), .B(n380), .Z(n18710) );
  XNOR U690 ( .A(n6371), .B(n6372), .Z(n6680) );
  XNOR U691 ( .A(n19881), .B(n19882), .Z(n19884) );
  XOR U692 ( .A(n7657), .B(n7658), .Z(n7965) );
  XNOR U693 ( .A(n6682), .B(n6683), .Z(n6998) );
  XNOR U694 ( .A(n19889), .B(n19890), .Z(n20206) );
  XNOR U695 ( .A(n19122), .B(n19123), .Z(n19441) );
  NAND U696 ( .A(n13300), .B(n13299), .Z(n381) );
  NAND U697 ( .A(n13018), .B(n13019), .Z(n382) );
  NAND U698 ( .A(n381), .B(n382), .Z(n13306) );
  XNOR U699 ( .A(n6999), .B(n7000), .Z(n7320) );
  XNOR U700 ( .A(n20224), .B(n20225), .Z(n20549) );
  NAND U701 ( .A(n19746), .B(n19748), .Z(n383) );
  XOR U702 ( .A(n19746), .B(n19748), .Z(n384) );
  NANDN U703 ( .A(n19745), .B(n384), .Z(n385) );
  NAND U704 ( .A(n383), .B(n385), .Z(n19753) );
  XNOR U705 ( .A(n8309), .B(n8310), .Z(n8652) );
  XNOR U706 ( .A(n20537), .B(n20538), .Z(n20540) );
  NAND U707 ( .A(n20447), .B(n20449), .Z(n386) );
  XOR U708 ( .A(n20447), .B(n20449), .Z(n387) );
  NANDN U709 ( .A(n20446), .B(n387), .Z(n388) );
  NAND U710 ( .A(n386), .B(n388), .Z(n20118) );
  XOR U711 ( .A(n20169), .B(n20168), .Z(n389) );
  NANDN U712 ( .A(n20171), .B(n389), .Z(n390) );
  NAND U713 ( .A(n20169), .B(n20168), .Z(n391) );
  AND U714 ( .A(n390), .B(n391), .Z(n20433) );
  NAND U715 ( .A(n19452), .B(n19451), .Z(n392) );
  NAND U716 ( .A(n18832), .B(n18833), .Z(n393) );
  NAND U717 ( .A(n392), .B(n393), .Z(n19139) );
  NAND U718 ( .A(n18786), .B(n18787), .Z(n394) );
  NAND U719 ( .A(n18467), .B(n18468), .Z(n395) );
  NAND U720 ( .A(n394), .B(n395), .Z(n18472) );
  XNOR U721 ( .A(n10223), .B(n10222), .Z(n10228) );
  NAND U722 ( .A(n20749), .B(n20752), .Z(n396) );
  XOR U723 ( .A(n20749), .B(n20752), .Z(n397) );
  NANDN U724 ( .A(n20750), .B(n397), .Z(n398) );
  NAND U725 ( .A(n396), .B(n398), .Z(n20489) );
  NAND U726 ( .A(n13320), .B(n13319), .Z(n399) );
  NAND U727 ( .A(n13026), .B(n13027), .Z(n400) );
  NAND U728 ( .A(n399), .B(n400), .Z(n13326) );
  NAND U729 ( .A(n9361), .B(n9362), .Z(n401) );
  NANDN U730 ( .A(n9714), .B(n9713), .Z(n402) );
  NAND U731 ( .A(n401), .B(n402), .Z(n9363) );
  NAND U732 ( .A(n21549), .B(n21548), .Z(n403) );
  NANDN U733 ( .A(n21215), .B(n21214), .Z(n404) );
  AND U734 ( .A(n403), .B(n404), .Z(n21218) );
  XOR U735 ( .A(n20827), .B(n20826), .Z(n405) );
  NANDN U736 ( .A(n20829), .B(n405), .Z(n406) );
  NAND U737 ( .A(n20827), .B(n20826), .Z(n407) );
  AND U738 ( .A(n406), .B(n407), .Z(n21101) );
  XNOR U739 ( .A(n9365), .B(n9366), .Z(n9368) );
  XNOR U740 ( .A(n9015), .B(n9016), .Z(n9371) );
  NAND U741 ( .A(n22838), .B(n22837), .Z(n408) );
  NANDN U742 ( .A(n22840), .B(n22839), .Z(n409) );
  NAND U743 ( .A(n408), .B(n409), .Z(n22866) );
  NAND U744 ( .A(n19147), .B(n19146), .Z(n410) );
  NAND U745 ( .A(n18799), .B(n18798), .Z(n411) );
  AND U746 ( .A(n410), .B(n411), .Z(n18802) );
  XNOR U747 ( .A(n21236), .B(n21237), .Z(n21570) );
  XNOR U748 ( .A(n21474), .B(n21475), .Z(n21477) );
  NAND U749 ( .A(n18823), .B(n18822), .Z(n412) );
  NANDN U750 ( .A(n19467), .B(n19468), .Z(n413) );
  NAND U751 ( .A(n412), .B(n413), .Z(n19149) );
  NAND U752 ( .A(n20136), .B(n20135), .Z(n414) );
  NANDN U753 ( .A(n20153), .B(n20152), .Z(n415) );
  AND U754 ( .A(n414), .B(n415), .Z(n20140) );
  NAND U755 ( .A(n17823), .B(n17822), .Z(n416) );
  NANDN U756 ( .A(n18149), .B(n18148), .Z(n417) );
  AND U757 ( .A(n416), .B(n417), .Z(n17827) );
  XNOR U758 ( .A(n9379), .B(n9380), .Z(n9384) );
  XNOR U759 ( .A(n21566), .B(n21567), .Z(n21888) );
  NAND U760 ( .A(n23124), .B(n23123), .Z(n418) );
  NANDN U761 ( .A(n23126), .B(n23125), .Z(n419) );
  NAND U762 ( .A(n418), .B(n419), .Z(n23363) );
  NAND U763 ( .A(n23115), .B(n23114), .Z(n420) );
  NAND U764 ( .A(n23112), .B(n23113), .Z(n421) );
  NAND U765 ( .A(n420), .B(n421), .Z(n23120) );
  NAND U766 ( .A(n23359), .B(n23360), .Z(n422) );
  NANDN U767 ( .A(n23362), .B(n23361), .Z(n423) );
  AND U768 ( .A(n422), .B(n423), .Z(n23478) );
  XOR U769 ( .A(n21483), .B(n21480), .Z(n424) );
  NANDN U770 ( .A(n21481), .B(n424), .Z(n425) );
  NAND U771 ( .A(n21483), .B(n21480), .Z(n426) );
  AND U772 ( .A(n425), .B(n426), .Z(n21149) );
  NAND U773 ( .A(n21147), .B(n21146), .Z(n427) );
  NANDN U774 ( .A(n20807), .B(n20806), .Z(n428) );
  AND U775 ( .A(n427), .B(n428), .Z(n20808) );
  NAND U776 ( .A(n18811), .B(n18810), .Z(n429) );
  XOR U777 ( .A(n18811), .B(n18810), .Z(n430) );
  NANDN U778 ( .A(n18813), .B(n430), .Z(n431) );
  NAND U779 ( .A(n429), .B(n431), .Z(n18486) );
  NAND U780 ( .A(n13654), .B(n13653), .Z(n432) );
  NANDN U781 ( .A(n14045), .B(n14044), .Z(n433) );
  AND U782 ( .A(n432), .B(n433), .Z(n13670) );
  XNOR U783 ( .A(n13688), .B(n13687), .Z(n13690) );
  XNOR U784 ( .A(n10102), .B(n10103), .Z(n10263) );
  XNOR U785 ( .A(n10257), .B(n10256), .Z(n10259) );
  NAND U786 ( .A(n19159), .B(n19158), .Z(n434) );
  NAND U787 ( .A(n19154), .B(n19155), .Z(n435) );
  NAND U788 ( .A(n434), .B(n435), .Z(n19479) );
  AND U789 ( .A(n20484), .B(n20483), .Z(n24682) );
  NAND U790 ( .A(n24663), .B(n24666), .Z(n436) );
  XOR U791 ( .A(n24663), .B(n24666), .Z(n437) );
  NAND U792 ( .A(n437), .B(n24664), .Z(n438) );
  NAND U793 ( .A(n436), .B(n438), .Z(n24670) );
  OR U794 ( .A(n24737), .B(n24738), .Z(n439) );
  NAND U795 ( .A(n24740), .B(n24739), .Z(n440) );
  NAND U796 ( .A(n439), .B(n440), .Z(n441) );
  NANDN U797 ( .A(n24750), .B(n441), .Z(n442) );
  NANDN U798 ( .A(n24745), .B(n14727), .Z(n443) );
  NAND U799 ( .A(n442), .B(n443), .Z(n444) );
  NOR U800 ( .A(n24741), .B(n24750), .Z(n445) );
  NAND U801 ( .A(n24744), .B(n445), .Z(n446) );
  NANDN U802 ( .A(n444), .B(n446), .Z(n447) );
  AND U803 ( .A(n24753), .B(n447), .Z(n448) );
  XOR U804 ( .A(n448), .B(n24756), .Z(n449) );
  NAND U805 ( .A(n449), .B(n24755), .Z(n450) );
  NAND U806 ( .A(n448), .B(n24756), .Z(n451) );
  AND U807 ( .A(n450), .B(n451), .Z(n24759) );
  NANDN U808 ( .A(n3644), .B(n3157), .Z(n452) );
  XNOR U809 ( .A(n3155), .B(n452), .Z(n453) );
  NANDN U810 ( .A(n3157), .B(n3156), .Z(n454) );
  NAND U811 ( .A(n453), .B(n454), .Z(n3397) );
  NANDN U812 ( .A(n4682), .B(n4149), .Z(n455) );
  XNOR U813 ( .A(n4147), .B(n455), .Z(n456) );
  NANDN U814 ( .A(n4149), .B(n4148), .Z(n457) );
  NAND U815 ( .A(n456), .B(n457), .Z(n4415) );
  NANDN U816 ( .A(n5828), .B(n5239), .Z(n458) );
  XNOR U817 ( .A(n5237), .B(n458), .Z(n459) );
  NANDN U818 ( .A(n5239), .B(n5238), .Z(n460) );
  NAND U819 ( .A(n459), .B(n460), .Z(n5535) );
  XNOR U820 ( .A(n2595), .B(n2596), .Z(n3153) );
  XNOR U821 ( .A(n3168), .B(n3169), .Z(n3390) );
  XNOR U822 ( .A(n3405), .B(n3406), .Z(n3661) );
  XNOR U823 ( .A(n3895), .B(n3896), .Z(n3898) );
  XNOR U824 ( .A(n4158), .B(n4159), .Z(n4161) );
  XNOR U825 ( .A(n5248), .B(n5249), .Z(n5251) );
  XNOR U826 ( .A(n4963), .B(n4964), .Z(n5256) );
  XNOR U827 ( .A(n5537), .B(n5538), .Z(n5839) );
  XNOR U828 ( .A(n5834), .B(n5835), .Z(n6138) );
  XNOR U829 ( .A(n4427), .B(n4428), .Z(n4705) );
  XNOR U830 ( .A(n4700), .B(n4701), .Z(n4973) );
  XNOR U831 ( .A(n4969), .B(n4970), .Z(n5260) );
  XNOR U832 ( .A(n5547), .B(n5548), .Z(n5851) );
  XNOR U833 ( .A(n5844), .B(n5845), .Z(n6125) );
  XNOR U834 ( .A(n3668), .B(n3669), .Z(n3881) );
  XNOR U835 ( .A(n6440), .B(n6441), .Z(n6730) );
  XNOR U836 ( .A(n6743), .B(n6744), .Z(n6746) );
  XNOR U837 ( .A(n5856), .B(n5857), .Z(n6160) );
  XNOR U838 ( .A(n5559), .B(n5560), .Z(n5863) );
  XNOR U839 ( .A(n6143), .B(n6144), .Z(n6451) );
  XNOR U840 ( .A(n3678), .B(n3679), .Z(n3879) );
  XNOR U841 ( .A(n4714), .B(n4715), .Z(n4947) );
  XNOR U842 ( .A(n4983), .B(n4984), .Z(n5234) );
  XNOR U843 ( .A(n4186), .B(n4187), .Z(n4454) );
  NANDN U844 ( .A(n7391), .B(n6734), .Z(n461) );
  XNOR U845 ( .A(n6732), .B(n461), .Z(n462) );
  NANDN U846 ( .A(n6734), .B(n6733), .Z(n463) );
  NAND U847 ( .A(n462), .B(n463), .Z(n7068) );
  XOR U848 ( .A(n6773), .B(n6774), .Z(n6775) );
  XOR U849 ( .A(n6470), .B(n6471), .Z(n6473) );
  XOR U850 ( .A(n6167), .B(n6168), .Z(n6169) );
  XOR U851 ( .A(n4724), .B(n4725), .Z(n4726) );
  XOR U852 ( .A(n5870), .B(n5871), .Z(n5873) );
  XNOR U853 ( .A(n7070), .B(n7071), .Z(n7402) );
  XNOR U854 ( .A(n6763), .B(n6764), .Z(n7056) );
  XNOR U855 ( .A(n5286), .B(n5287), .Z(n5586) );
  XNOR U856 ( .A(n5579), .B(n5580), .Z(n5822) );
  XNOR U857 ( .A(n7059), .B(n7060), .Z(n7383) );
  XNOR U858 ( .A(n7384), .B(n7385), .Z(n7387) );
  XNOR U859 ( .A(n7419), .B(n7420), .Z(n7722) );
  XNOR U860 ( .A(n5005), .B(n5006), .Z(n5228) );
  XNOR U861 ( .A(n7409), .B(n7410), .Z(n7751) );
  XNOR U862 ( .A(n7122), .B(n7123), .Z(n7374) );
  XNOR U863 ( .A(n6791), .B(n6792), .Z(n7053) );
  XNOR U864 ( .A(n6490), .B(n6491), .Z(n6722) );
  XNOR U865 ( .A(n5009), .B(n5010), .Z(n5012) );
  XNOR U866 ( .A(n5593), .B(n5594), .Z(n5815) );
  XNOR U867 ( .A(n7738), .B(n7739), .Z(n7741) );
  XNOR U868 ( .A(n6421), .B(n6422), .Z(n6495) );
  XNOR U869 ( .A(n6189), .B(n6190), .Z(n6420) );
  XNOR U870 ( .A(n8054), .B(n8055), .Z(n8057) );
  XNOR U871 ( .A(n7792), .B(n7793), .Z(n8128) );
  XNOR U872 ( .A(n6193), .B(n6194), .Z(n6505) );
  XNOR U873 ( .A(n5892), .B(n5893), .Z(n6200) );
  XNOR U874 ( .A(n8071), .B(n8072), .Z(n8074) );
  XNOR U875 ( .A(n7772), .B(n7773), .Z(n8049) );
  XNOR U876 ( .A(n8099), .B(n8100), .Z(n8102) );
  XNOR U877 ( .A(n8125), .B(n8126), .Z(n8378) );
  XNOR U878 ( .A(n7798), .B(n7799), .Z(n8040) );
  XNOR U879 ( .A(n7455), .B(n7456), .Z(n7712) );
  XNOR U880 ( .A(n7134), .B(n7135), .Z(n7371) );
  XNOR U881 ( .A(n6803), .B(n6804), .Z(n7141) );
  XNOR U882 ( .A(n8085), .B(n8086), .Z(n8388) );
  XNOR U883 ( .A(n8089), .B(n8090), .Z(n8386) );
  XNOR U884 ( .A(n8105), .B(n8106), .Z(n8443) );
  XNOR U885 ( .A(n6205), .B(n6206), .Z(n6513) );
  XNOR U886 ( .A(n8402), .B(n8403), .Z(n8748) );
  XOR U887 ( .A(n6815), .B(n6816), .Z(n6818) );
  XNOR U888 ( .A(n8414), .B(n8415), .Z(n8747) );
  XOR U889 ( .A(n8791), .B(n8792), .Z(n8794) );
  XNOR U890 ( .A(n8381), .B(n8382), .Z(n8455) );
  XNOR U891 ( .A(n8379), .B(n8380), .Z(n8458) );
  XNOR U892 ( .A(n8375), .B(n8376), .Z(n8479) );
  XNOR U893 ( .A(n8141), .B(n8142), .Z(n8484) );
  XNOR U894 ( .A(n7812), .B(n7813), .Z(n8145) );
  XNOR U895 ( .A(n8801), .B(n8802), .Z(n9110) );
  XNOR U896 ( .A(n8837), .B(n8838), .Z(n9148) );
  XNOR U897 ( .A(n7818), .B(n7819), .Z(n8151) );
  XNOR U898 ( .A(n7477), .B(n7478), .Z(n7822) );
  XOR U899 ( .A(n9049), .B(n9050), .Z(n464) );
  NANDN U900 ( .A(n9052), .B(n9051), .Z(n465) );
  NAND U901 ( .A(n464), .B(n465), .Z(n9427) );
  XNOR U902 ( .A(n9075), .B(n9076), .Z(n9456) );
  XNOR U903 ( .A(n8811), .B(n8812), .Z(n9042) );
  XNOR U904 ( .A(n8763), .B(n8764), .Z(n9068) );
  XNOR U905 ( .A(n9063), .B(n9064), .Z(n9425) );
  XOR U906 ( .A(n9095), .B(n9096), .Z(n9420) );
  XOR U907 ( .A(n8726), .B(n8727), .Z(n8729) );
  XNOR U908 ( .A(n9047), .B(n9048), .Z(n9422) );
  XNOR U909 ( .A(n9812), .B(n9813), .Z(n10319) );
  XNOR U910 ( .A(n9415), .B(n9416), .Z(n9484) );
  XNOR U911 ( .A(n9117), .B(n9118), .Z(n9492) );
  XOR U912 ( .A(n9523), .B(n9524), .Z(n9887) );
  XNOR U913 ( .A(n8500), .B(n8501), .Z(n8722) );
  XNOR U914 ( .A(n8163), .B(n8164), .Z(n8372) );
  XNOR U915 ( .A(n9794), .B(n9795), .Z(n10301) );
  XOR U916 ( .A(n9423), .B(n9424), .Z(n9468) );
  XNOR U917 ( .A(n9479), .B(n9480), .Z(n9841) );
  XNOR U918 ( .A(n9846), .B(n9847), .Z(n10355) );
  XNOR U919 ( .A(n9517), .B(n9518), .Z(n9880) );
  XOR U920 ( .A(n9529), .B(n9530), .Z(n9900) );
  XNOR U921 ( .A(n9409), .B(n9410), .Z(n9905) );
  XNOR U922 ( .A(n10731), .B(n10732), .Z(n10734) );
  XNOR U923 ( .A(n10296), .B(n10297), .Z(n10748) );
  XNOR U924 ( .A(n10324), .B(n10325), .Z(n10327) );
  XNOR U925 ( .A(n9836), .B(n9837), .Z(n10342) );
  XNOR U926 ( .A(n9868), .B(n9869), .Z(n9870) );
  XNOR U927 ( .A(n10743), .B(n10744), .Z(n11023) );
  XOR U928 ( .A(n10709), .B(n10710), .Z(n11115) );
  XNOR U929 ( .A(n9177), .B(n9178), .Z(n9180) );
  XNOR U930 ( .A(n2850), .B(n2849), .Z(n2851) );
  XNOR U931 ( .A(n11004), .B(n11005), .Z(n11444) );
  XNOR U932 ( .A(n11437), .B(n11438), .Z(n11723) );
  XNOR U933 ( .A(n11020), .B(n11021), .Z(n11457) );
  XNOR U934 ( .A(n10308), .B(n10309), .Z(n10757) );
  XNOR U935 ( .A(n10788), .B(n10789), .Z(n10791) );
  XNOR U936 ( .A(n10386), .B(n10387), .Z(n10711) );
  XNOR U937 ( .A(n10414), .B(n10415), .Z(n10820) );
  NAND U938 ( .A(n11526), .B(n11529), .Z(n466) );
  XOR U939 ( .A(n11526), .B(n11529), .Z(n467) );
  NANDN U940 ( .A(n11527), .B(n467), .Z(n468) );
  NAND U941 ( .A(n466), .B(n468), .Z(n11120) );
  XOR U942 ( .A(n11125), .B(n11127), .Z(n469) );
  NANDN U943 ( .A(n11126), .B(n469), .Z(n470) );
  NAND U944 ( .A(n11125), .B(n11127), .Z(n471) );
  AND U945 ( .A(n470), .B(n471), .Z(n10818) );
  XNOR U946 ( .A(n10418), .B(n10419), .Z(n10705) );
  XOR U947 ( .A(n10264), .B(n10265), .Z(n10430) );
  XNOR U948 ( .A(n9549), .B(n9550), .Z(n9927) );
  XNOR U949 ( .A(n11718), .B(n11719), .Z(n12145) );
  XNOR U950 ( .A(n12138), .B(n12139), .Z(n12446) );
  XOR U951 ( .A(n11029), .B(n11030), .Z(n472) );
  XNOR U952 ( .A(n11028), .B(n472), .Z(n11472) );
  XNOR U953 ( .A(n10758), .B(n10759), .Z(n11033) );
  XNOR U954 ( .A(n11467), .B(n11468), .Z(n11753) );
  XNOR U955 ( .A(n11049), .B(n11050), .Z(n11486) );
  XNOR U956 ( .A(n10338), .B(n10339), .Z(n10775) );
  XNOR U957 ( .A(n11088), .B(n11089), .Z(n11091) );
  NAND U958 ( .A(n11100), .B(n11102), .Z(n473) );
  XOR U959 ( .A(n11100), .B(n11102), .Z(n474) );
  NANDN U960 ( .A(n11101), .B(n474), .Z(n475) );
  NAND U961 ( .A(n473), .B(n475), .Z(n10802) );
  XNOR U962 ( .A(n9924), .B(n9925), .Z(n10433) );
  XNOR U963 ( .A(n2894), .B(n2893), .Z(n2895) );
  XNOR U964 ( .A(n12441), .B(n12442), .Z(n12843) );
  XNOR U965 ( .A(n11063), .B(n11064), .Z(n11493) );
  NAND U966 ( .A(n11512), .B(n11515), .Z(n476) );
  XOR U967 ( .A(n11512), .B(n11515), .Z(n477) );
  NANDN U968 ( .A(n11513), .B(n477), .Z(n478) );
  NAND U969 ( .A(n476), .B(n478), .Z(n11104) );
  NAND U970 ( .A(n11828), .B(n11831), .Z(n479) );
  XOR U971 ( .A(n11828), .B(n11831), .Z(n480) );
  NANDN U972 ( .A(n11829), .B(n480), .Z(n481) );
  NAND U973 ( .A(n479), .B(n481), .Z(n11530) );
  XNOR U974 ( .A(n12836), .B(n12837), .Z(n13073) );
  XNOR U975 ( .A(n11746), .B(n11747), .Z(n12170) );
  XNOR U976 ( .A(n11477), .B(n11478), .Z(n11765) );
  NAND U977 ( .A(n12122), .B(n12125), .Z(n482) );
  XOR U978 ( .A(n12122), .B(n12125), .Z(n483) );
  NANDN U979 ( .A(n12123), .B(n483), .Z(n484) );
  NAND U980 ( .A(n482), .B(n484), .Z(n11776) );
  NANDN U981 ( .A(n11780), .B(n11491), .Z(n485) );
  NAND U982 ( .A(n11780), .B(n11781), .Z(n486) );
  NANDN U983 ( .A(n11779), .B(n486), .Z(n487) );
  NAND U984 ( .A(n485), .B(n487), .Z(n11495) );
  NANDN U985 ( .A(n12215), .B(n11802), .Z(n488) );
  NAND U986 ( .A(n12215), .B(n12216), .Z(n489) );
  NANDN U987 ( .A(n12214), .B(n489), .Z(n490) );
  NAND U988 ( .A(n488), .B(n490), .Z(n11808) );
  XOR U989 ( .A(n11813), .B(n11815), .Z(n491) );
  NANDN U990 ( .A(n11814), .B(n491), .Z(n492) );
  NAND U991 ( .A(n11813), .B(n11815), .Z(n493) );
  AND U992 ( .A(n492), .B(n493), .Z(n11510) );
  NAND U993 ( .A(n12238), .B(n12241), .Z(n494) );
  XOR U994 ( .A(n12238), .B(n12241), .Z(n495) );
  NANDN U995 ( .A(n12239), .B(n495), .Z(n496) );
  NAND U996 ( .A(n494), .B(n496), .Z(n11833) );
  XNOR U997 ( .A(n11145), .B(n11146), .Z(n11551) );
  XNOR U998 ( .A(n10838), .B(n10839), .Z(n11155) );
  XNOR U999 ( .A(n2932), .B(n2931), .Z(n2933) );
  XNOR U1000 ( .A(n13068), .B(n13069), .Z(n13392) );
  XNOR U1001 ( .A(n12457), .B(n12458), .Z(n12460) );
  XNOR U1002 ( .A(n11760), .B(n11761), .Z(n12182) );
  XOR U1003 ( .A(n12254), .B(n12255), .Z(n497) );
  NANDN U1004 ( .A(n12256), .B(n497), .Z(n498) );
  NAND U1005 ( .A(n12254), .B(n12255), .Z(n499) );
  AND U1006 ( .A(n498), .B(n499), .Z(n11849) );
  XOR U1007 ( .A(n11544), .B(n11545), .Z(n11852) );
  XNOR U1008 ( .A(n11157), .B(n11158), .Z(n11557) );
  XNOR U1009 ( .A(n2966), .B(n2965), .Z(n2968) );
  XNOR U1010 ( .A(n13385), .B(n13386), .Z(n13742) );
  XNOR U1011 ( .A(n12463), .B(n12464), .Z(n12466) );
  XNOR U1012 ( .A(n12160), .B(n12161), .Z(n12472) );
  XNOR U1013 ( .A(n12202), .B(n12203), .Z(n12506) );
  XNOR U1014 ( .A(n12208), .B(n12209), .Z(n12512) );
  NAND U1015 ( .A(n12535), .B(n12536), .Z(n500) );
  XOR U1016 ( .A(n12535), .B(n12536), .Z(n501) );
  NANDN U1017 ( .A(n12534), .B(n501), .Z(n502) );
  NAND U1018 ( .A(n500), .B(n502), .Z(n12229) );
  XNOR U1019 ( .A(n12244), .B(n12245), .Z(n12555) );
  NAND U1020 ( .A(n12940), .B(n12939), .Z(n503) );
  XOR U1021 ( .A(n12940), .B(n12939), .Z(n504) );
  NANDN U1022 ( .A(n12941), .B(n504), .Z(n505) );
  NAND U1023 ( .A(n503), .B(n505), .Z(n12551) );
  NAND U1024 ( .A(n11862), .B(n11865), .Z(n506) );
  XOR U1025 ( .A(n11862), .B(n11865), .Z(n507) );
  NANDN U1026 ( .A(n11863), .B(n507), .Z(n508) );
  NAND U1027 ( .A(n506), .B(n508), .Z(n11555) );
  XOR U1028 ( .A(n2946), .B(n2945), .Z(n3309) );
  XNOR U1029 ( .A(n14102), .B(n14103), .Z(n14105) );
  XNOR U1030 ( .A(n13743), .B(n13744), .Z(n14093) );
  XNOR U1031 ( .A(n13090), .B(n13091), .Z(n13093) );
  XNOR U1032 ( .A(n12487), .B(n12488), .Z(n12886) );
  XNOR U1033 ( .A(n12190), .B(n12191), .Z(n12427) );
  NAND U1034 ( .A(n12923), .B(n12921), .Z(n509) );
  XOR U1035 ( .A(n12923), .B(n12921), .Z(n510) );
  NANDN U1036 ( .A(n12922), .B(n510), .Z(n511) );
  NAND U1037 ( .A(n509), .B(n511), .Z(n12533) );
  NANDN U1038 ( .A(n12574), .B(n12270), .Z(n512) );
  NAND U1039 ( .A(n12574), .B(n12575), .Z(n513) );
  NANDN U1040 ( .A(n12573), .B(n513), .Z(n514) );
  NAND U1041 ( .A(n512), .B(n514), .Z(n12276) );
  XNOR U1042 ( .A(n14110), .B(n14111), .Z(n14432) );
  XNOR U1043 ( .A(n13759), .B(n13760), .Z(n13762) );
  XNOR U1044 ( .A(n13098), .B(n13099), .Z(n13417) );
  XNOR U1045 ( .A(n12864), .B(n12865), .Z(n13057) );
  XNOR U1046 ( .A(n12497), .B(n12498), .Z(n12820) );
  XOR U1047 ( .A(n12917), .B(n12918), .Z(n515) );
  XNOR U1048 ( .A(n12916), .B(n515), .Z(n13149) );
  NAND U1049 ( .A(n13173), .B(n13171), .Z(n516) );
  XOR U1050 ( .A(n13173), .B(n13171), .Z(n517) );
  NANDN U1051 ( .A(n13172), .B(n517), .Z(n518) );
  NAND U1052 ( .A(n516), .B(n518), .Z(n12937) );
  XOR U1053 ( .A(n12417), .B(n12418), .Z(n12962) );
  NAND U1054 ( .A(n13195), .B(n13198), .Z(n519) );
  XOR U1055 ( .A(n13195), .B(n13198), .Z(n520) );
  NANDN U1056 ( .A(n13196), .B(n520), .Z(n521) );
  NAND U1057 ( .A(n519), .B(n521), .Z(n12959) );
  XNOR U1058 ( .A(n3006), .B(n3005), .Z(n3011) );
  XOR U1059 ( .A(n3028), .B(n3027), .Z(n3033) );
  XNOR U1060 ( .A(n13407), .B(n13408), .Z(n13768) );
  NAND U1061 ( .A(n13811), .B(n13814), .Z(n522) );
  XOR U1062 ( .A(n13811), .B(n13814), .Z(n523) );
  NANDN U1063 ( .A(n13812), .B(n523), .Z(n524) );
  NAND U1064 ( .A(n522), .B(n524), .Z(n13468) );
  NAND U1065 ( .A(n13474), .B(n13477), .Z(n525) );
  XOR U1066 ( .A(n13474), .B(n13477), .Z(n526) );
  NANDN U1067 ( .A(n13475), .B(n526), .Z(n527) );
  NAND U1068 ( .A(n525), .B(n527), .Z(n13145) );
  XNOR U1069 ( .A(n13199), .B(n13200), .Z(n13531) );
  XNOR U1070 ( .A(n13527), .B(n13528), .Z(n13884) );
  XOR U1071 ( .A(n12588), .B(n12589), .Z(n12590) );
  XOR U1072 ( .A(n3555), .B(n3556), .Z(n3805) );
  XNOR U1073 ( .A(n3048), .B(n3047), .Z(n3049) );
  XNOR U1074 ( .A(n14124), .B(n14125), .Z(n14127) );
  XNOR U1075 ( .A(n13425), .B(n13426), .Z(n13781) );
  XNOR U1076 ( .A(n13108), .B(n13109), .Z(n13429) );
  XNOR U1077 ( .A(n13519), .B(n13520), .Z(n528) );
  XNOR U1078 ( .A(n13518), .B(n528), .Z(n13871) );
  NAND U1079 ( .A(n13541), .B(n13544), .Z(n529) );
  XOR U1080 ( .A(n13541), .B(n13544), .Z(n530) );
  NANDN U1081 ( .A(n13542), .B(n530), .Z(n531) );
  NAND U1082 ( .A(n529), .B(n531), .Z(n13216) );
  XNOR U1083 ( .A(n3806), .B(n3807), .Z(n4063) );
  XNOR U1084 ( .A(n3561), .B(n3562), .Z(n3810) );
  XNOR U1085 ( .A(n14446), .B(n14447), .Z(n14819) );
  XNOR U1086 ( .A(n13797), .B(n13798), .Z(n13799) );
  NAND U1087 ( .A(n14186), .B(n14189), .Z(n532) );
  XOR U1088 ( .A(n14186), .B(n14189), .Z(n533) );
  NANDN U1089 ( .A(n14187), .B(n533), .Z(n534) );
  NAND U1090 ( .A(n532), .B(n534), .Z(n13816) );
  XOR U1091 ( .A(n13501), .B(n13502), .Z(n535) );
  XNOR U1092 ( .A(n13500), .B(n535), .Z(n13712) );
  XOR U1093 ( .A(n14557), .B(n14559), .Z(n536) );
  NANDN U1094 ( .A(n14558), .B(n536), .Z(n537) );
  NAND U1095 ( .A(n14557), .B(n14559), .Z(n538) );
  AND U1096 ( .A(n537), .B(n538), .Z(n14242) );
  NAND U1097 ( .A(n13893), .B(n13896), .Z(n539) );
  XOR U1098 ( .A(n13893), .B(n13896), .Z(n540) );
  NANDN U1099 ( .A(n13894), .B(n540), .Z(n541) );
  NAND U1100 ( .A(n539), .B(n541), .Z(n13545) );
  XNOR U1101 ( .A(n4061), .B(n4062), .Z(n4325) );
  XNOR U1102 ( .A(n3074), .B(n3073), .Z(n3075) );
  XOR U1103 ( .A(n3094), .B(n3093), .Z(n3099) );
  XOR U1104 ( .A(n13844), .B(n13845), .Z(n542) );
  XNOR U1105 ( .A(n13843), .B(n542), .Z(n14083) );
  NAND U1106 ( .A(n14541), .B(n14544), .Z(n543) );
  XOR U1107 ( .A(n14541), .B(n14544), .Z(n544) );
  NANDN U1108 ( .A(n14542), .B(n544), .Z(n545) );
  NAND U1109 ( .A(n543), .B(n545), .Z(n14226) );
  XOR U1110 ( .A(n3573), .B(n3574), .Z(n3825) );
  XNOR U1111 ( .A(n3039), .B(n3040), .Z(n3344) );
  XNOR U1112 ( .A(n3108), .B(n3107), .Z(n3111) );
  XNOR U1113 ( .A(n14832), .B(n14833), .Z(n15159) );
  XOR U1114 ( .A(n14167), .B(n14169), .Z(n546) );
  NANDN U1115 ( .A(n14168), .B(n546), .Z(n547) );
  NAND U1116 ( .A(n14167), .B(n14169), .Z(n548) );
  AND U1117 ( .A(n547), .B(n548), .Z(n14175) );
  XOR U1118 ( .A(n14084), .B(n14085), .Z(n14528) );
  NAND U1119 ( .A(n14903), .B(n14906), .Z(n549) );
  XOR U1120 ( .A(n14903), .B(n14906), .Z(n550) );
  NANDN U1121 ( .A(n14904), .B(n550), .Z(n551) );
  NAND U1122 ( .A(n549), .B(n551), .Z(n14531) );
  NAND U1123 ( .A(n14919), .B(n14922), .Z(n552) );
  XOR U1124 ( .A(n14919), .B(n14922), .Z(n553) );
  NANDN U1125 ( .A(n14920), .B(n553), .Z(n554) );
  NAND U1126 ( .A(n552), .B(n554), .Z(n14546) );
  NAND U1127 ( .A(n15242), .B(n15245), .Z(n555) );
  XOR U1128 ( .A(n15242), .B(n15245), .Z(n556) );
  NANDN U1129 ( .A(n15243), .B(n556), .Z(n557) );
  NAND U1130 ( .A(n555), .B(n557), .Z(n14917) );
  NAND U1131 ( .A(n14954), .B(n14957), .Z(n558) );
  XOR U1132 ( .A(n14954), .B(n14957), .Z(n559) );
  NANDN U1133 ( .A(n14955), .B(n559), .Z(n560) );
  NAND U1134 ( .A(n558), .B(n560), .Z(n14576) );
  XNOR U1135 ( .A(n14262), .B(n14263), .Z(n561) );
  XNOR U1136 ( .A(n14261), .B(n561), .Z(n14387) );
  NAND U1137 ( .A(n15640), .B(n15643), .Z(n562) );
  XOR U1138 ( .A(n15640), .B(n15643), .Z(n563) );
  NANDN U1139 ( .A(n15641), .B(n563), .Z(n564) );
  NAND U1140 ( .A(n562), .B(n564), .Z(n15273) );
  XNOR U1141 ( .A(n13910), .B(n13911), .Z(n14279) );
  NAND U1142 ( .A(n13558), .B(n13560), .Z(n565) );
  XOR U1143 ( .A(n13558), .B(n13560), .Z(n566) );
  NANDN U1144 ( .A(n13557), .B(n566), .Z(n567) );
  NAND U1145 ( .A(n565), .B(n567), .Z(n13228) );
  XNOR U1146 ( .A(n4591), .B(n4592), .Z(n4866) );
  XNOR U1147 ( .A(n3579), .B(n3580), .Z(n3828) );
  XOR U1148 ( .A(n10139), .B(n10138), .Z(n10132) );
  XNOR U1149 ( .A(n14472), .B(n14473), .Z(n14849) );
  XNOR U1150 ( .A(n14844), .B(n14845), .Z(n15171) );
  XNOR U1151 ( .A(n14162), .B(n14163), .Z(n14485) );
  NAND U1152 ( .A(n15256), .B(n15259), .Z(n568) );
  XOR U1153 ( .A(n15256), .B(n15259), .Z(n569) );
  NANDN U1154 ( .A(n15257), .B(n569), .Z(n570) );
  NAND U1155 ( .A(n568), .B(n570), .Z(n14936) );
  XNOR U1156 ( .A(n14392), .B(n14393), .Z(n14934) );
  NAND U1157 ( .A(n14969), .B(n14972), .Z(n571) );
  XOR U1158 ( .A(n14969), .B(n14972), .Z(n572) );
  NANDN U1159 ( .A(n14970), .B(n572), .Z(n573) );
  NAND U1160 ( .A(n571), .B(n573), .Z(n14590) );
  XOR U1161 ( .A(n14586), .B(n14588), .Z(n574) );
  NANDN U1162 ( .A(n14587), .B(n574), .Z(n575) );
  NAND U1163 ( .A(n14586), .B(n14588), .Z(n576) );
  AND U1164 ( .A(n575), .B(n576), .Z(n14277) );
  NAND U1165 ( .A(n13230), .B(n13229), .Z(n577) );
  NAND U1166 ( .A(n12990), .B(n12991), .Z(n578) );
  NAND U1167 ( .A(n577), .B(n578), .Z(n13236) );
  XNOR U1168 ( .A(n4599), .B(n4600), .Z(n4872) );
  XNOR U1169 ( .A(n3830), .B(n3831), .Z(n4086) );
  XNOR U1170 ( .A(n14486), .B(n14487), .Z(n14860) );
  XNOR U1171 ( .A(n14856), .B(n14857), .Z(n15183) );
  XOR U1172 ( .A(n14505), .B(n14506), .Z(n579) );
  XNOR U1173 ( .A(n14504), .B(n579), .Z(n14775) );
  XNOR U1174 ( .A(n15228), .B(n15229), .Z(n15589) );
  NAND U1175 ( .A(n15603), .B(n15606), .Z(n580) );
  XOR U1176 ( .A(n15603), .B(n15606), .Z(n581) );
  NANDN U1177 ( .A(n15604), .B(n581), .Z(n582) );
  NAND U1178 ( .A(n580), .B(n582), .Z(n15241) );
  XNOR U1179 ( .A(n15649), .B(n15650), .Z(n15984) );
  XOR U1180 ( .A(n3591), .B(n3592), .Z(n3841) );
  XNOR U1181 ( .A(n4087), .B(n4088), .Z(n4348) );
  XNOR U1182 ( .A(n22677), .B(n22676), .Z(n22678) );
  XNOR U1183 ( .A(n14866), .B(n14867), .Z(n15102) );
  NANDN U1184 ( .A(n15671), .B(n15298), .Z(n583) );
  NAND U1185 ( .A(n15671), .B(n15672), .Z(n584) );
  NANDN U1186 ( .A(n15670), .B(n584), .Z(n585) );
  NAND U1187 ( .A(n583), .B(n585), .Z(n15304) );
  XNOR U1188 ( .A(n3597), .B(n3598), .Z(n3846) );
  XNOR U1189 ( .A(n22671), .B(n22670), .Z(n22672) );
  XOR U1190 ( .A(n15921), .B(n15922), .Z(n586) );
  NANDN U1191 ( .A(n15924), .B(n586), .Z(n587) );
  NAND U1192 ( .A(n15921), .B(n15922), .Z(n588) );
  AND U1193 ( .A(n587), .B(n588), .Z(n15929) );
  XOR U1194 ( .A(n15979), .B(n15980), .Z(n589) );
  XNOR U1195 ( .A(n15978), .B(n589), .Z(n16139) );
  XNOR U1196 ( .A(n15307), .B(n15308), .Z(n15310) );
  XNOR U1197 ( .A(n4099), .B(n4100), .Z(n4363) );
  XNOR U1198 ( .A(n5727), .B(n5728), .Z(n6024) );
  XOR U1199 ( .A(n10157), .B(n10156), .Z(n10162) );
  NAND U1200 ( .A(n15897), .B(n15900), .Z(n590) );
  XOR U1201 ( .A(n15897), .B(n15900), .Z(n591) );
  NANDN U1202 ( .A(n15898), .B(n591), .Z(n592) );
  NAND U1203 ( .A(n590), .B(n592), .Z(n15570) );
  NAND U1204 ( .A(n15572), .B(n15575), .Z(n593) );
  XOR U1205 ( .A(n15572), .B(n15575), .Z(n594) );
  NANDN U1206 ( .A(n15573), .B(n594), .Z(n595) );
  NAND U1207 ( .A(n593), .B(n595), .Z(n15463) );
  NAND U1208 ( .A(n16652), .B(n16655), .Z(n596) );
  XOR U1209 ( .A(n16652), .B(n16655), .Z(n597) );
  NANDN U1210 ( .A(n16653), .B(n597), .Z(n598) );
  NAND U1211 ( .A(n596), .B(n598), .Z(n16326) );
  NAND U1212 ( .A(n17045), .B(n17048), .Z(n599) );
  XOR U1213 ( .A(n17045), .B(n17048), .Z(n600) );
  NANDN U1214 ( .A(n17046), .B(n600), .Z(n601) );
  NAND U1215 ( .A(n599), .B(n601), .Z(n16681) );
  XNOR U1216 ( .A(n16684), .B(n16685), .Z(n16686) );
  NAND U1217 ( .A(n13250), .B(n13249), .Z(n602) );
  NAND U1218 ( .A(n12998), .B(n12999), .Z(n603) );
  NAND U1219 ( .A(n602), .B(n603), .Z(n13256) );
  XNOR U1220 ( .A(n6026), .B(n6027), .Z(n6330) );
  XNOR U1221 ( .A(n5733), .B(n5734), .Z(n6030) );
  NAND U1222 ( .A(n16262), .B(n16265), .Z(n604) );
  XOR U1223 ( .A(n16262), .B(n16265), .Z(n605) );
  NANDN U1224 ( .A(n16263), .B(n605), .Z(n606) );
  NAND U1225 ( .A(n604), .B(n606), .Z(n15902) );
  XOR U1226 ( .A(n15948), .B(n15949), .Z(n607) );
  XNOR U1227 ( .A(n15947), .B(n607), .Z(n16148) );
  NAND U1228 ( .A(n17016), .B(n17019), .Z(n608) );
  XOR U1229 ( .A(n17016), .B(n17019), .Z(n609) );
  NANDN U1230 ( .A(n17017), .B(n609), .Z(n610) );
  NAND U1231 ( .A(n608), .B(n610), .Z(n16657) );
  NANDN U1232 ( .A(n17378), .B(n17042), .Z(n611) );
  NAND U1233 ( .A(n17378), .B(n17379), .Z(n612) );
  NANDN U1234 ( .A(n17377), .B(n612), .Z(n613) );
  NAND U1235 ( .A(n611), .B(n613), .Z(n17044) );
  XOR U1236 ( .A(n16373), .B(n16374), .Z(n614) );
  XNOR U1237 ( .A(n16372), .B(n614), .Z(n16467) );
  NAND U1238 ( .A(n17058), .B(n17060), .Z(n615) );
  XOR U1239 ( .A(n17058), .B(n17060), .Z(n616) );
  NANDN U1240 ( .A(n17059), .B(n616), .Z(n617) );
  NAND U1241 ( .A(n615), .B(n617), .Z(n16696) );
  XNOR U1242 ( .A(n4629), .B(n4630), .Z(n4903) );
  XNOR U1243 ( .A(n6327), .B(n6328), .Z(n6376) );
  XOR U1244 ( .A(n5171), .B(n5172), .Z(n5457) );
  XOR U1245 ( .A(n16625), .B(n16626), .Z(n618) );
  NANDN U1246 ( .A(n16627), .B(n618), .Z(n619) );
  NAND U1247 ( .A(n16625), .B(n16626), .Z(n620) );
  AND U1248 ( .A(n619), .B(n620), .Z(n16485) );
  XOR U1249 ( .A(n16481), .B(n16482), .Z(n621) );
  NANDN U1250 ( .A(n16484), .B(n621), .Z(n622) );
  NAND U1251 ( .A(n16481), .B(n16482), .Z(n623) );
  AND U1252 ( .A(n622), .B(n623), .Z(n16639) );
  XNOR U1253 ( .A(n4904), .B(n4905), .Z(n5183) );
  XNOR U1254 ( .A(n4635), .B(n4636), .Z(n4908) );
  XOR U1255 ( .A(n16978), .B(n16976), .Z(n624) );
  NANDN U1256 ( .A(n16975), .B(n624), .Z(n625) );
  NAND U1257 ( .A(n16978), .B(n16976), .Z(n626) );
  AND U1258 ( .A(n625), .B(n626), .Z(n16624) );
  NAND U1259 ( .A(n17736), .B(n17739), .Z(n627) );
  XOR U1260 ( .A(n17736), .B(n17739), .Z(n628) );
  NANDN U1261 ( .A(n17737), .B(n628), .Z(n629) );
  NAND U1262 ( .A(n627), .B(n629), .Z(n17381) );
  NAND U1263 ( .A(n17751), .B(n17754), .Z(n630) );
  XOR U1264 ( .A(n17751), .B(n17754), .Z(n631) );
  NANDN U1265 ( .A(n17752), .B(n631), .Z(n632) );
  NAND U1266 ( .A(n630), .B(n632), .Z(n17397) );
  XNOR U1267 ( .A(n17061), .B(n17062), .Z(n17158) );
  XNOR U1268 ( .A(n17065), .B(n17066), .Z(n17156) );
  XOR U1269 ( .A(n16711), .B(n16712), .Z(n16713) );
  NANDN U1270 ( .A(n17326), .B(n16991), .Z(n633) );
  NAND U1271 ( .A(n17326), .B(n17327), .Z(n634) );
  NANDN U1272 ( .A(n17325), .B(n634), .Z(n635) );
  NAND U1273 ( .A(n633), .B(n635), .Z(n17167) );
  XNOR U1274 ( .A(n17742), .B(n17743), .Z(n17846) );
  NAND U1275 ( .A(n13270), .B(n13269), .Z(n636) );
  NAND U1276 ( .A(n13006), .B(n13007), .Z(n637) );
  NAND U1277 ( .A(n636), .B(n637), .Z(n13276) );
  XNOR U1278 ( .A(n6686), .B(n6687), .Z(n6963) );
  NAND U1279 ( .A(n17693), .B(n17696), .Z(n638) );
  XOR U1280 ( .A(n17693), .B(n17696), .Z(n639) );
  NANDN U1281 ( .A(n17694), .B(n639), .Z(n640) );
  NAND U1282 ( .A(n638), .B(n640), .Z(n17329) );
  XNOR U1283 ( .A(n17730), .B(n17731), .Z(n641) );
  XNOR U1284 ( .A(n17729), .B(n641), .Z(n18051) );
  XOR U1285 ( .A(n18742), .B(n18743), .Z(n642) );
  NANDN U1286 ( .A(n18744), .B(n642), .Z(n643) );
  NAND U1287 ( .A(n18742), .B(n18743), .Z(n644) );
  AND U1288 ( .A(n643), .B(n644), .Z(n18424) );
  NAND U1289 ( .A(n18082), .B(n18085), .Z(n645) );
  XOR U1290 ( .A(n18082), .B(n18085), .Z(n646) );
  NANDN U1291 ( .A(n18083), .B(n646), .Z(n647) );
  NAND U1292 ( .A(n645), .B(n647), .Z(n17768) );
  NAND U1293 ( .A(n18432), .B(n18435), .Z(n648) );
  XOR U1294 ( .A(n18432), .B(n18435), .Z(n649) );
  NANDN U1295 ( .A(n18433), .B(n649), .Z(n650) );
  NAND U1296 ( .A(n648), .B(n650), .Z(n18087) );
  XNOR U1297 ( .A(n5761), .B(n5762), .Z(n6061) );
  XNOR U1298 ( .A(n6054), .B(n6055), .Z(n6359) );
  NAND U1299 ( .A(n18034), .B(n18036), .Z(n651) );
  XOR U1300 ( .A(n18034), .B(n18036), .Z(n652) );
  NANDN U1301 ( .A(n18035), .B(n652), .Z(n653) );
  NAND U1302 ( .A(n651), .B(n653), .Z(n17854) );
  XOR U1303 ( .A(n18048), .B(n18049), .Z(n654) );
  XNOR U1304 ( .A(n18047), .B(n654), .Z(n18197) );
  XNOR U1305 ( .A(n18055), .B(n18056), .Z(n18192) );
  XNOR U1306 ( .A(n5769), .B(n5770), .Z(n6066) );
  NAND U1307 ( .A(n18378), .B(n18381), .Z(n655) );
  XOR U1308 ( .A(n18378), .B(n18381), .Z(n656) );
  NANDN U1309 ( .A(n18379), .B(n656), .Z(n657) );
  NAND U1310 ( .A(n655), .B(n657), .Z(n18033) );
  XNOR U1311 ( .A(n18745), .B(n18746), .Z(n19090) );
  XNOR U1312 ( .A(n7296), .B(n7297), .Z(n7326) );
  XNOR U1313 ( .A(n7623), .B(n7624), .Z(n7660) );
  XOR U1314 ( .A(n7661), .B(n7662), .Z(n7957) );
  XNOR U1315 ( .A(n6068), .B(n6069), .Z(n6372) );
  NAND U1316 ( .A(n18703), .B(n18706), .Z(n658) );
  XOR U1317 ( .A(n18703), .B(n18706), .Z(n659) );
  NANDN U1318 ( .A(n18704), .B(n659), .Z(n660) );
  NAND U1319 ( .A(n658), .B(n660), .Z(n18503) );
  XOR U1320 ( .A(n18717), .B(n18718), .Z(n661) );
  NANDN U1321 ( .A(n18720), .B(n661), .Z(n662) );
  NAND U1322 ( .A(n18717), .B(n18718), .Z(n663) );
  AND U1323 ( .A(n662), .B(n663), .Z(n18727) );
  NANDN U1324 ( .A(n19425), .B(n19105), .Z(n664) );
  NAND U1325 ( .A(n19425), .B(n19426), .Z(n665) );
  NANDN U1326 ( .A(n19424), .B(n665), .Z(n666) );
  NAND U1327 ( .A(n664), .B(n666), .Z(n19107) );
  XOR U1328 ( .A(n18497), .B(n18498), .Z(n19116) );
  XNOR U1329 ( .A(n18449), .B(n18450), .Z(n18495) );
  NAND U1330 ( .A(n13290), .B(n13289), .Z(n667) );
  NAND U1331 ( .A(n13014), .B(n13015), .Z(n668) );
  NAND U1332 ( .A(n667), .B(n668), .Z(n13296) );
  XNOR U1333 ( .A(n7304), .B(n7305), .Z(n7631) );
  XNOR U1334 ( .A(n6369), .B(n6370), .Z(n6681) );
  NAND U1335 ( .A(n19767), .B(n19770), .Z(n669) );
  XOR U1336 ( .A(n19767), .B(n19770), .Z(n670) );
  NANDN U1337 ( .A(n19768), .B(n670), .Z(n671) );
  NAND U1338 ( .A(n669), .B(n671), .Z(n19428) );
  NAND U1339 ( .A(n16412), .B(n16411), .Z(n672) );
  NANDN U1340 ( .A(n16742), .B(n16741), .Z(n673) );
  AND U1341 ( .A(n672), .B(n673), .Z(n16416) );
  XOR U1342 ( .A(n6993), .B(n6994), .Z(n7315) );
  XNOR U1343 ( .A(n19883), .B(n19884), .Z(n20223) );
  XNOR U1344 ( .A(n20216), .B(n20217), .Z(n20219) );
  NAND U1345 ( .A(n19730), .B(n19733), .Z(n674) );
  XOR U1346 ( .A(n19730), .B(n19733), .Z(n675) );
  NANDN U1347 ( .A(n19731), .B(n675), .Z(n676) );
  NAND U1348 ( .A(n674), .B(n676), .Z(n19394) );
  XOR U1349 ( .A(n19761), .B(n19762), .Z(n677) );
  XNOR U1350 ( .A(n19760), .B(n677), .Z(n19836) );
  XNOR U1351 ( .A(n19162), .B(n19163), .Z(n19447) );
  XOR U1352 ( .A(n19132), .B(n19135), .Z(n678) );
  NANDN U1353 ( .A(n19133), .B(n678), .Z(n679) );
  NAND U1354 ( .A(n19132), .B(n19135), .Z(n680) );
  AND U1355 ( .A(n679), .B(n680), .Z(n18831) );
  XOR U1356 ( .A(n8329), .B(n8330), .Z(n8649) );
  XNOR U1357 ( .A(n8307), .B(n8308), .Z(n8653) );
  NAND U1358 ( .A(n20115), .B(n20116), .Z(n681) );
  XOR U1359 ( .A(n20115), .B(n20116), .Z(n682) );
  NANDN U1360 ( .A(n20114), .B(n682), .Z(n683) );
  NAND U1361 ( .A(n681), .B(n683), .Z(n19794) );
  NAND U1362 ( .A(n13310), .B(n13309), .Z(n684) );
  NAND U1363 ( .A(n13022), .B(n13023), .Z(n685) );
  NAND U1364 ( .A(n684), .B(n685), .Z(n13316) );
  XOR U1365 ( .A(n7990), .B(n7991), .Z(n8314) );
  XNOR U1366 ( .A(n7649), .B(n7650), .Z(n7984) );
  XNOR U1367 ( .A(n20545), .B(n20546), .Z(n20865) );
  XNOR U1368 ( .A(n20555), .B(n20556), .Z(n20558) );
  XOR U1369 ( .A(n20758), .B(n20759), .Z(n686) );
  NANDN U1370 ( .A(n20761), .B(n686), .Z(n687) );
  NAND U1371 ( .A(n20758), .B(n20759), .Z(n688) );
  AND U1372 ( .A(n687), .B(n688), .Z(n20764) );
  NAND U1373 ( .A(n20778), .B(n20781), .Z(n689) );
  XOR U1374 ( .A(n20778), .B(n20781), .Z(n690) );
  NANDN U1375 ( .A(n20779), .B(n690), .Z(n691) );
  NAND U1376 ( .A(n689), .B(n691), .Z(n20450) );
  XNOR U1377 ( .A(n20117), .B(n20118), .Z(n20162) );
  XOR U1378 ( .A(n18827), .B(n18824), .Z(n692) );
  NANDN U1379 ( .A(n18825), .B(n692), .Z(n693) );
  NAND U1380 ( .A(n18827), .B(n18824), .Z(n694) );
  AND U1381 ( .A(n693), .B(n694), .Z(n18791) );
  NAND U1382 ( .A(n17116), .B(n17115), .Z(n695) );
  NANDN U1383 ( .A(n17458), .B(n17457), .Z(n696) );
  AND U1384 ( .A(n695), .B(n696), .Z(n17120) );
  XNOR U1385 ( .A(n20874), .B(n20875), .Z(n20877) );
  XNOR U1386 ( .A(n20882), .B(n20883), .Z(n21216) );
  NAND U1387 ( .A(n19454), .B(n19453), .Z(n697) );
  NANDN U1388 ( .A(n19498), .B(n19499), .Z(n698) );
  NAND U1389 ( .A(n697), .B(n698), .Z(n19458) );
  NAND U1390 ( .A(n19456), .B(n19455), .Z(n699) );
  NAND U1391 ( .A(n19138), .B(n19139), .Z(n700) );
  NAND U1392 ( .A(n699), .B(n700), .Z(n19460) );
  NAND U1393 ( .A(n18789), .B(n18788), .Z(n701) );
  NAND U1394 ( .A(n18471), .B(n18472), .Z(n702) );
  NAND U1395 ( .A(n701), .B(n702), .Z(n18793) );
  XNOR U1396 ( .A(n8325), .B(n8326), .Z(n8671) );
  XNOR U1397 ( .A(n20892), .B(n20893), .Z(n21229) );
  XNOR U1398 ( .A(n20794), .B(n20795), .Z(n21134) );
  NAND U1399 ( .A(n20159), .B(n20157), .Z(n703) );
  XOR U1400 ( .A(n20159), .B(n20157), .Z(n704) );
  NANDN U1401 ( .A(n20156), .B(n704), .Z(n705) );
  NAND U1402 ( .A(n703), .B(n705), .Z(n20132) );
  NAND U1403 ( .A(n12763), .B(n12762), .Z(n706) );
  NANDN U1404 ( .A(n13325), .B(n13326), .Z(n707) );
  NAND U1405 ( .A(n706), .B(n707), .Z(n13031) );
  XOR U1406 ( .A(n9017), .B(n9018), .Z(n9372) );
  XNOR U1407 ( .A(n22583), .B(n22582), .Z(n22577) );
  NAND U1408 ( .A(n21092), .B(n21095), .Z(n708) );
  XOR U1409 ( .A(n21092), .B(n21095), .Z(n709) );
  NANDN U1410 ( .A(n21093), .B(n709), .Z(n710) );
  NAND U1411 ( .A(n708), .B(n710), .Z(n20827) );
  XNOR U1412 ( .A(n21460), .B(n21461), .Z(n21462) );
  NAND U1413 ( .A(n20461), .B(n20460), .Z(n711) );
  NANDN U1414 ( .A(n20485), .B(n20486), .Z(n712) );
  NAND U1415 ( .A(n711), .B(n712), .Z(n20800) );
  XNOR U1416 ( .A(n9385), .B(n9386), .Z(n9720) );
  XNOR U1417 ( .A(n10239), .B(n10238), .Z(n10241) );
  XNOR U1418 ( .A(n22569), .B(n22568), .Z(n22570) );
  NAND U1419 ( .A(n22869), .B(n22868), .Z(n713) );
  NAND U1420 ( .A(n22867), .B(n22866), .Z(n714) );
  NAND U1421 ( .A(n713), .B(n714), .Z(n23108) );
  XNOR U1422 ( .A(n21224), .B(n21225), .Z(n21559) );
  XNOR U1423 ( .A(n21234), .B(n21235), .Z(n21571) );
  NAND U1424 ( .A(n19491), .B(n19490), .Z(n715) );
  NAND U1425 ( .A(n19466), .B(n19465), .Z(n716) );
  NAND U1426 ( .A(n715), .B(n716), .Z(n19470) );
  NAND U1427 ( .A(n18803), .B(n18802), .Z(n717) );
  NANDN U1428 ( .A(n18819), .B(n18818), .Z(n718) );
  AND U1429 ( .A(n717), .B(n718), .Z(n18807) );
  XNOR U1430 ( .A(n10245), .B(n10244), .Z(n10247) );
  XNOR U1431 ( .A(n21554), .B(n21555), .Z(n21845) );
  XNOR U1432 ( .A(n21564), .B(n21565), .Z(n21889) );
  NAND U1433 ( .A(n17140), .B(n17139), .Z(n719) );
  NANDN U1434 ( .A(n17492), .B(n17491), .Z(n720) );
  AND U1435 ( .A(n719), .B(n720), .Z(n17144) );
  NAND U1436 ( .A(n14050), .B(n14051), .Z(n721) );
  NANDN U1437 ( .A(n14037), .B(n14036), .Z(n722) );
  AND U1438 ( .A(n721), .B(n722), .Z(n14039) );
  XNOR U1439 ( .A(n9729), .B(n9730), .Z(n10101) );
  XOR U1440 ( .A(n22283), .B(n22284), .Z(n723) );
  NANDN U1441 ( .A(n22286), .B(n723), .Z(n724) );
  NAND U1442 ( .A(n22283), .B(n22284), .Z(n725) );
  AND U1443 ( .A(n724), .B(n725), .Z(n21967) );
  XOR U1444 ( .A(n22363), .B(n22364), .Z(n726) );
  NANDN U1445 ( .A(n22366), .B(n726), .Z(n727) );
  NAND U1446 ( .A(n22363), .B(n22364), .Z(n728) );
  AND U1447 ( .A(n727), .B(n728), .Z(n22043) );
  NAND U1448 ( .A(n21823), .B(n21825), .Z(n729) );
  XOR U1449 ( .A(n21823), .B(n21825), .Z(n730) );
  NANDN U1450 ( .A(n21822), .B(n730), .Z(n731) );
  NAND U1451 ( .A(n729), .B(n731), .Z(n21485) );
  NAND U1452 ( .A(n20155), .B(n20154), .Z(n732) );
  NANDN U1453 ( .A(n20810), .B(n20811), .Z(n733) );
  NAND U1454 ( .A(n732), .B(n733), .Z(n20475) );
  NAND U1455 ( .A(n23364), .B(n23363), .Z(n734) );
  NANDN U1456 ( .A(n23366), .B(n23365), .Z(n735) );
  NAND U1457 ( .A(n734), .B(n735), .Z(n23367) );
  NAND U1458 ( .A(n23119), .B(n23120), .Z(n736) );
  NANDN U1459 ( .A(n23122), .B(n23121), .Z(n737) );
  AND U1460 ( .A(n736), .B(n737), .Z(n23249) );
  NAND U1461 ( .A(n23480), .B(n23479), .Z(n738) );
  NAND U1462 ( .A(n23478), .B(n23477), .Z(n739) );
  AND U1463 ( .A(n738), .B(n739), .Z(n23596) );
  XOR U1464 ( .A(n22464), .B(n22461), .Z(n740) );
  NAND U1465 ( .A(n740), .B(n22462), .Z(n741) );
  NAND U1466 ( .A(n22464), .B(n22461), .Z(n742) );
  AND U1467 ( .A(n741), .B(n742), .Z(n22469) );
  NAND U1468 ( .A(n22146), .B(n22147), .Z(n743) );
  NANDN U1469 ( .A(n22164), .B(n22163), .Z(n744) );
  NAND U1470 ( .A(n743), .B(n744), .Z(n22484) );
  NAND U1471 ( .A(n19478), .B(n19477), .Z(n745) );
  NANDN U1472 ( .A(n19483), .B(n19482), .Z(n746) );
  AND U1473 ( .A(n745), .B(n746), .Z(n20150) );
  AND U1474 ( .A(n20478), .B(n20479), .Z(n24684) );
  NAND U1475 ( .A(n18487), .B(n18488), .Z(n747) );
  NANDN U1476 ( .A(n18159), .B(n18158), .Z(n748) );
  AND U1477 ( .A(n747), .B(n748), .Z(n18490) );
  NAND U1478 ( .A(n18815), .B(n18814), .Z(n749) );
  NAND U1479 ( .A(n18486), .B(n18485), .Z(n750) );
  NAND U1480 ( .A(n749), .B(n750), .Z(n18491) );
  AND U1481 ( .A(n19479), .B(n19480), .Z(n24702) );
  NAND U1482 ( .A(n22993), .B(n22992), .Z(n751) );
  NANDN U1483 ( .A(n22995), .B(n22994), .Z(n752) );
  NAND U1484 ( .A(n751), .B(n752), .Z(n23117) );
  ANDN U1485 ( .B(n22496), .A(n22495), .Z(n24674) );
  NAND U1486 ( .A(n24722), .B(n24724), .Z(n753) );
  XOR U1487 ( .A(n24722), .B(n24724), .Z(n754) );
  NANDN U1488 ( .A(n24721), .B(n754), .Z(n755) );
  NAND U1489 ( .A(n753), .B(n755), .Z(n24726) );
  ANDN U1490 ( .B(n13701), .A(n13702), .Z(n24764) );
  NAND U1491 ( .A(n24784), .B(n24786), .Z(n756) );
  XOR U1492 ( .A(n24784), .B(n24786), .Z(n757) );
  NANDN U1493 ( .A(n24783), .B(n757), .Z(n758) );
  NAND U1494 ( .A(n756), .B(n758), .Z(n24788) );
  NAND U1495 ( .A(n24793), .B(n24796), .Z(n759) );
  XOR U1496 ( .A(n24793), .B(n24796), .Z(n760) );
  NANDN U1497 ( .A(n24794), .B(n760), .Z(n761) );
  NAND U1498 ( .A(n759), .B(n761), .Z(n22847) );
  NAND U1499 ( .A(n23818), .B(n23817), .Z(n762) );
  NAND U1500 ( .A(n23816), .B(n23815), .Z(n763) );
  NAND U1501 ( .A(n762), .B(n763), .Z(n23913) );
  NAND U1502 ( .A(n24643), .B(n24644), .Z(n764) );
  NANDN U1503 ( .A(n24646), .B(n24645), .Z(n765) );
  AND U1504 ( .A(n764), .B(n765), .Z(n24654) );
  NANDN U1505 ( .A(n4148), .B(n3645), .Z(n766) );
  XNOR U1506 ( .A(n3643), .B(n766), .Z(n767) );
  NANDN U1507 ( .A(n3645), .B(n3644), .Z(n768) );
  NAND U1508 ( .A(n767), .B(n768), .Z(n3889) );
  NANDN U1509 ( .A(n4951), .B(n4412), .Z(n769) );
  XNOR U1510 ( .A(n4410), .B(n769), .Z(n770) );
  NANDN U1511 ( .A(n4412), .B(n4411), .Z(n771) );
  NAND U1512 ( .A(n770), .B(n771), .Z(n4686) );
  XNOR U1513 ( .A(n4688), .B(n4689), .Z(n4962) );
  XNOR U1514 ( .A(n4957), .B(n4958), .Z(n5249) );
  NANDN U1515 ( .A(n2473), .B(n2374), .Z(n772) );
  XNOR U1516 ( .A(n2372), .B(n772), .Z(n2376) );
  XNOR U1517 ( .A(n3656), .B(n3657), .Z(n3882) );
  XNOR U1518 ( .A(n3897), .B(n3898), .Z(n4164) );
  XNOR U1519 ( .A(n4160), .B(n4161), .Z(n4429) );
  XNOR U1520 ( .A(n4423), .B(n4424), .Z(n4701) );
  XNOR U1521 ( .A(n5541), .B(n5542), .Z(n5544) );
  NANDN U1522 ( .A(n6428), .B(n5829), .Z(n773) );
  XNOR U1523 ( .A(n5827), .B(n773), .Z(n774) );
  NANDN U1524 ( .A(n5829), .B(n5828), .Z(n775) );
  NAND U1525 ( .A(n774), .B(n775), .Z(n6131) );
  XNOR U1526 ( .A(n2599), .B(n2600), .Z(n3177) );
  XNOR U1527 ( .A(n3172), .B(n3173), .Z(n3389) );
  XNOR U1528 ( .A(n3660), .B(n3661), .Z(n3663) );
  XNOR U1529 ( .A(n3409), .B(n3410), .Z(n3666) );
  XNOR U1530 ( .A(n4698), .B(n4699), .Z(n4974) );
  XNOR U1531 ( .A(n4967), .B(n4968), .Z(n5261) );
  XNOR U1532 ( .A(n5254), .B(n5255), .Z(n5554) );
  XNOR U1533 ( .A(n6133), .B(n6134), .Z(n6439) );
  XNOR U1534 ( .A(n5838), .B(n5839), .Z(n5841) );
  XNOR U1535 ( .A(n6137), .B(n6138), .Z(n6140) );
  XNOR U1536 ( .A(n6434), .B(n6435), .Z(n6744) );
  XNOR U1537 ( .A(n4172), .B(n4173), .Z(n4408) );
  XNOR U1538 ( .A(n4435), .B(n4436), .Z(n4679) );
  XNOR U1539 ( .A(n5852), .B(n5853), .Z(n6122) );
  XNOR U1540 ( .A(n3672), .B(n3673), .Z(n3916) );
  XNOR U1541 ( .A(n3911), .B(n3912), .Z(n4181) );
  XNOR U1542 ( .A(n4979), .B(n4980), .Z(n5273) );
  XNOR U1543 ( .A(n5266), .B(n5267), .Z(n5566) );
  XNOR U1544 ( .A(n3676), .B(n3677), .Z(n3679) );
  XNOR U1545 ( .A(n6157), .B(n6158), .Z(n6424) );
  XNOR U1546 ( .A(n5563), .B(n5564), .Z(n5824) );
  XNOR U1547 ( .A(n5860), .B(n5861), .Z(n6121) );
  XNOR U1548 ( .A(n6739), .B(n6740), .Z(n7075) );
  XNOR U1549 ( .A(n6728), .B(n6729), .Z(n6760) );
  XNOR U1550 ( .A(n6749), .B(n6750), .Z(n7087) );
  XNOR U1551 ( .A(n4720), .B(n4721), .Z(n4994) );
  XNOR U1552 ( .A(n5276), .B(n5277), .Z(n5574) );
  XNOR U1553 ( .A(n4989), .B(n4990), .Z(n5281) );
  XNOR U1554 ( .A(n6456), .B(n6457), .Z(n6764) );
  XNOR U1555 ( .A(n6769), .B(n6770), .Z(n7103) );
  XNOR U1556 ( .A(n7082), .B(n7083), .Z(n7413) );
  XOR U1557 ( .A(n4141), .B(n4142), .Z(n4191) );
  XOR U1558 ( .A(n4453), .B(n4454), .Z(n4455) );
  XNOR U1559 ( .A(n6781), .B(n6782), .Z(n7115) );
  XNOR U1560 ( .A(n6476), .B(n6477), .Z(n6725) );
  XNOR U1561 ( .A(n6175), .B(n6176), .Z(n6483) );
  XNOR U1562 ( .A(n4999), .B(n5000), .Z(n5230) );
  XNOR U1563 ( .A(n5876), .B(n5877), .Z(n6119) );
  NANDN U1564 ( .A(n7728), .B(n7065), .Z(n776) );
  XNOR U1565 ( .A(n7063), .B(n776), .Z(n777) );
  NANDN U1566 ( .A(n7065), .B(n7064), .Z(n778) );
  NAND U1567 ( .A(n777), .B(n778), .Z(n7395) );
  XNOR U1568 ( .A(n7401), .B(n7402), .Z(n7404) );
  XNOR U1569 ( .A(n7108), .B(n7109), .Z(n7377) );
  XNOR U1570 ( .A(n5587), .B(n5588), .Z(n5820) );
  XNOR U1571 ( .A(n7721), .B(n7722), .Z(n7723) );
  XNOR U1572 ( .A(n7425), .B(n7426), .Z(n7767) );
  XNOR U1573 ( .A(n7443), .B(n7444), .Z(n7715) );
  XOR U1574 ( .A(n5227), .B(n5228), .Z(n5295) );
  XNOR U1575 ( .A(n7750), .B(n7751), .Z(n7753) );
  XNOR U1576 ( .A(n7756), .B(n7757), .Z(n8055) );
  XNOR U1577 ( .A(n7429), .B(n7430), .Z(n7432) );
  XNOR U1578 ( .A(n7380), .B(n7381), .Z(n7718) );
  XNOR U1579 ( .A(n7447), .B(n7448), .Z(n7714) );
  XNOR U1580 ( .A(n5597), .B(n5598), .Z(n5814) );
  XOR U1581 ( .A(n5300), .B(n5301), .Z(n5606) );
  XNOR U1582 ( .A(n7740), .B(n7741), .Z(n8078) );
  XNOR U1583 ( .A(n7372), .B(n7373), .Z(n7452) );
  XNOR U1584 ( .A(n7130), .B(n7131), .Z(n7458) );
  XNOR U1585 ( .A(n6799), .B(n6800), .Z(n7135) );
  XNOR U1586 ( .A(n6419), .B(n6420), .Z(n6499) );
  XNOR U1587 ( .A(n7796), .B(n7797), .Z(n8041) );
  NAND U1588 ( .A(n3214), .B(n3215), .Z(n779) );
  NANDN U1589 ( .A(n3371), .B(n3370), .Z(n780) );
  NAND U1590 ( .A(n779), .B(n780), .Z(n3368) );
  XNOR U1591 ( .A(n8073), .B(n8074), .Z(n8406) );
  XOR U1592 ( .A(n8430), .B(n8431), .Z(n8432) );
  XNOR U1593 ( .A(n8046), .B(n8047), .Z(n8120) );
  XNOR U1594 ( .A(n8044), .B(n8045), .Z(n8463) );
  XNOR U1595 ( .A(n6811), .B(n6812), .Z(n7147) );
  XNOR U1596 ( .A(n6508), .B(n6509), .Z(n6816) );
  XNOR U1597 ( .A(n8387), .B(n8388), .Z(n8418) );
  XNOR U1598 ( .A(n8109), .B(n8110), .Z(n8449) );
  XNOR U1599 ( .A(n8438), .B(n8439), .Z(n8740) );
  XNOR U1600 ( .A(n8137), .B(n8138), .Z(n8376) );
  XOR U1601 ( .A(n7806), .B(n7807), .Z(n7809) );
  XNOR U1602 ( .A(n6512), .B(n6513), .Z(n6515) );
  NANDN U1603 ( .A(n8751), .B(n8062), .Z(n781) );
  XNOR U1604 ( .A(n8060), .B(n781), .Z(n782) );
  NANDN U1605 ( .A(n8062), .B(n8061), .Z(n783) );
  NAND U1606 ( .A(n782), .B(n783), .Z(n8394) );
  XNOR U1607 ( .A(n8422), .B(n8423), .Z(n8786) );
  XOR U1608 ( .A(n8831), .B(n8832), .Z(n8834) );
  XNOR U1609 ( .A(n7471), .B(n7472), .Z(n7819) );
  XNOR U1610 ( .A(n7152), .B(n7153), .Z(n7478) );
  XNOR U1611 ( .A(n8396), .B(n8397), .Z(n8762) );
  XNOR U1612 ( .A(n8482), .B(n8483), .Z(n8731) );
  XNOR U1613 ( .A(n8147), .B(n8148), .Z(n8489) );
  XNOR U1614 ( .A(n7816), .B(n7817), .Z(n8152) );
  XNOR U1615 ( .A(n9099), .B(n9100), .Z(n9102) );
  XNOR U1616 ( .A(n8815), .B(n8816), .Z(n8818) );
  XNOR U1617 ( .A(n8736), .B(n8737), .Z(n8821) );
  XNOR U1618 ( .A(n8841), .B(n8842), .Z(n9037) );
  XNOR U1619 ( .A(n7483), .B(n7484), .Z(n7828) );
  XNOR U1620 ( .A(n9057), .B(n9058), .Z(n9440) );
  XNOR U1621 ( .A(n9782), .B(n9783), .Z(n10289) );
  XOR U1622 ( .A(n9085), .B(n9086), .Z(n9088) );
  XNOR U1623 ( .A(n9081), .B(n9082), .Z(n9463) );
  XNOR U1624 ( .A(n9111), .B(n9112), .Z(n9414) );
  XNOR U1625 ( .A(n9041), .B(n9042), .Z(n9121) );
  XNOR U1626 ( .A(n9441), .B(n9442), .Z(n9792) );
  XNOR U1627 ( .A(n9786), .B(n9787), .Z(n10295) );
  XNOR U1628 ( .A(n9810), .B(n9811), .Z(n9813) );
  XNOR U1629 ( .A(n9515), .B(n9516), .Z(n9518) );
  XNOR U1630 ( .A(n9411), .B(n9412), .Z(n9892) );
  XNOR U1631 ( .A(n9165), .B(n9166), .Z(n9536) );
  XNOR U1632 ( .A(n8724), .B(n8725), .Z(n8851) );
  XNOR U1633 ( .A(n8498), .B(n8499), .Z(n8723) );
  XNOR U1634 ( .A(n9069), .B(n9070), .Z(n9449) );
  XNOR U1635 ( .A(n9848), .B(n9849), .Z(n10354) );
  XNOR U1636 ( .A(n9505), .B(n9506), .Z(n9869) );
  XNOR U1637 ( .A(n9888), .B(n9889), .Z(n10272) );
  NAND U1638 ( .A(n9905), .B(n9907), .Z(n784) );
  XOR U1639 ( .A(n9905), .B(n9907), .Z(n785) );
  NANDN U1640 ( .A(n9906), .B(n785), .Z(n786) );
  NAND U1641 ( .A(n784), .B(n786), .Z(n9534) );
  XNOR U1642 ( .A(n8371), .B(n8372), .Z(n8504) );
  XNOR U1643 ( .A(n10284), .B(n10285), .Z(n10737) );
  XNOR U1644 ( .A(n9451), .B(n9452), .Z(n9804) );
  XNOR U1645 ( .A(n9822), .B(n9823), .Z(n9825) );
  XNOR U1646 ( .A(n9840), .B(n9841), .Z(n9843) );
  XNOR U1647 ( .A(n9834), .B(n9835), .Z(n10343) );
  XNOR U1648 ( .A(n9493), .B(n9494), .Z(n9860) );
  XOR U1649 ( .A(n9511), .B(n9512), .Z(n9875) );
  XNOR U1650 ( .A(n10739), .B(n10740), .Z(n11014) );
  XNOR U1651 ( .A(n10302), .B(n10303), .Z(n10754) );
  XNOR U1652 ( .A(n10749), .B(n10750), .Z(n10992) );
  XOR U1653 ( .A(n9828), .B(n9829), .Z(n9830) );
  XNOR U1654 ( .A(n10326), .B(n10327), .Z(n10718) );
  XNOR U1655 ( .A(n10764), .B(n10765), .Z(n11047) );
  XNOR U1656 ( .A(n10344), .B(n10345), .Z(n10776) );
  XNOR U1657 ( .A(n9858), .B(n9859), .Z(n10367) );
  XNOR U1658 ( .A(n9876), .B(n9877), .Z(n10384) );
  XNOR U1659 ( .A(n10268), .B(n10269), .Z(n10270) );
  XNOR U1660 ( .A(n10404), .B(n10405), .Z(n10814) );
  XOR U1661 ( .A(n9543), .B(n9544), .Z(n9919) );
  XNOR U1662 ( .A(n9179), .B(n9180), .Z(n9547) );
  XNOR U1663 ( .A(n10778), .B(n10779), .Z(n11074) );
  NAND U1664 ( .A(n11115), .B(n11118), .Z(n787) );
  XOR U1665 ( .A(n11115), .B(n11118), .Z(n788) );
  NANDN U1666 ( .A(n11116), .B(n788), .Z(n789) );
  NAND U1667 ( .A(n787), .B(n789), .Z(n10812) );
  XNOR U1668 ( .A(n10422), .B(n10423), .Z(n790) );
  XNOR U1669 ( .A(n10424), .B(n790), .Z(n10827) );
  XNOR U1670 ( .A(n2866), .B(n2865), .Z(n2867) );
  XNOR U1671 ( .A(n11443), .B(n11444), .Z(n11728) );
  XOR U1672 ( .A(n11425), .B(n11426), .Z(n11448) );
  XNOR U1673 ( .A(n10756), .B(n10757), .Z(n11034) );
  XNOR U1674 ( .A(n11057), .B(n11058), .Z(n11489) );
  XNOR U1675 ( .A(n11061), .B(n11062), .Z(n11064) );
  XNOR U1676 ( .A(n10790), .B(n10791), .Z(n11096) );
  XNOR U1677 ( .A(n10380), .B(n10381), .Z(n10800) );
  XOR U1678 ( .A(n11136), .B(n11138), .Z(n791) );
  NANDN U1679 ( .A(n11137), .B(n791), .Z(n792) );
  NAND U1680 ( .A(n11136), .B(n11138), .Z(n793) );
  AND U1681 ( .A(n792), .B(n793), .Z(n10824) );
  XNOR U1682 ( .A(n12144), .B(n12145), .Z(n12451) );
  XOR U1683 ( .A(n12126), .B(n12127), .Z(n12149) );
  XNOR U1684 ( .A(n11752), .B(n11753), .Z(n11755) );
  XNOR U1685 ( .A(n11090), .B(n11091), .Z(n11505) );
  NAND U1686 ( .A(n11803), .B(n11806), .Z(n794) );
  XOR U1687 ( .A(n11803), .B(n11806), .Z(n795) );
  NANDN U1688 ( .A(n11804), .B(n795), .Z(n796) );
  NAND U1689 ( .A(n794), .B(n796), .Z(n11506) );
  XNOR U1690 ( .A(n11100), .B(n11101), .Z(n797) );
  XNOR U1691 ( .A(n11102), .B(n797), .Z(n11416) );
  XNOR U1692 ( .A(n11839), .B(n11840), .Z(n798) );
  XNOR U1693 ( .A(n11838), .B(n798), .Z(n12252) );
  XNOR U1694 ( .A(n10435), .B(n10436), .Z(n10836) );
  XNOR U1695 ( .A(n2916), .B(n2915), .Z(n2917) );
  XNOR U1696 ( .A(n12842), .B(n12843), .Z(n13078) );
  XOR U1697 ( .A(n12824), .B(n12825), .Z(n12847) );
  XOR U1698 ( .A(n11748), .B(n11749), .Z(n12171) );
  XNOR U1699 ( .A(n11473), .B(n11474), .Z(n11758) );
  XNOR U1700 ( .A(n11039), .B(n11040), .Z(n11424) );
  XNOR U1701 ( .A(n11070), .B(n11071), .Z(n799) );
  XNOR U1702 ( .A(n11069), .B(n799), .Z(n11421) );
  XNOR U1703 ( .A(n11132), .B(n11133), .Z(n11545) );
  XNOR U1704 ( .A(n12178), .B(n12179), .Z(n12485) );
  XNOR U1705 ( .A(n11788), .B(n11789), .Z(n12209) );
  XNOR U1706 ( .A(n11807), .B(n11808), .Z(n12118) );
  XNOR U1707 ( .A(n11542), .B(n11543), .Z(n11853) );
  XOR U1708 ( .A(n11846), .B(n11845), .Z(n800) );
  XNOR U1709 ( .A(n11847), .B(n800), .Z(n12113) );
  XNOR U1710 ( .A(n11149), .B(n11150), .Z(n11406) );
  XNOR U1711 ( .A(n2944), .B(n2943), .Z(n2945) );
  XNOR U1712 ( .A(n2960), .B(n2959), .Z(n2961) );
  XNOR U1713 ( .A(n13391), .B(n13392), .Z(n13747) );
  XOR U1714 ( .A(n13373), .B(n13374), .Z(n13396) );
  XNOR U1715 ( .A(n11742), .B(n11743), .Z(n12165) );
  XNOR U1716 ( .A(n11766), .B(n11767), .Z(n12189) );
  XNOR U1717 ( .A(n12194), .B(n12195), .Z(n12505) );
  XOR U1718 ( .A(n12215), .B(n12216), .Z(n801) );
  XNOR U1719 ( .A(n12214), .B(n801), .Z(n12425) );
  XNOR U1720 ( .A(n12247), .B(n12248), .Z(n802) );
  XNOR U1721 ( .A(n12246), .B(n802), .Z(n12556) );
  NAND U1722 ( .A(n12271), .B(n12274), .Z(n803) );
  XOR U1723 ( .A(n12271), .B(n12274), .Z(n804) );
  NANDN U1724 ( .A(n12272), .B(n804), .Z(n805) );
  NAND U1725 ( .A(n803), .B(n805), .Z(n11867) );
  XNOR U1726 ( .A(n2907), .B(n2908), .Z(n3308) );
  XNOR U1727 ( .A(n2980), .B(n2979), .Z(n2981) );
  XNOR U1728 ( .A(n12166), .B(n12167), .Z(n12430) );
  XNOR U1729 ( .A(n13092), .B(n13093), .Z(n13412) );
  XNOR U1730 ( .A(n12858), .B(n12859), .Z(n13099) );
  XNOR U1731 ( .A(n12465), .B(n12466), .Z(n12863) );
  XNOR U1732 ( .A(n12471), .B(n12472), .Z(n12868) );
  XOR U1733 ( .A(n12232), .B(n12233), .Z(n806) );
  XNOR U1734 ( .A(n12231), .B(n806), .Z(n12423) );
  XNOR U1735 ( .A(n12535), .B(n12536), .Z(n807) );
  XNOR U1736 ( .A(n12534), .B(n807), .Z(n12812) );
  XNOR U1737 ( .A(n12551), .B(n12552), .Z(n12810) );
  NAND U1738 ( .A(n13184), .B(n13187), .Z(n808) );
  XOR U1739 ( .A(n13184), .B(n13187), .Z(n809) );
  NANDN U1740 ( .A(n13185), .B(n809), .Z(n810) );
  NAND U1741 ( .A(n808), .B(n810), .Z(n12951) );
  NAND U1742 ( .A(n13519), .B(n13518), .Z(n811) );
  XOR U1743 ( .A(n13519), .B(n13518), .Z(n812) );
  NANDN U1744 ( .A(n13520), .B(n812), .Z(n813) );
  NAND U1745 ( .A(n811), .B(n813), .Z(n13188) );
  XNOR U1746 ( .A(n12275), .B(n12276), .Z(n12415) );
  XOR U1747 ( .A(n12574), .B(n12575), .Z(n814) );
  XNOR U1748 ( .A(n12573), .B(n814), .Z(n12805) );
  XOR U1749 ( .A(n11870), .B(n11871), .Z(n11872) );
  XNOR U1750 ( .A(n2974), .B(n2973), .Z(n2976) );
  XNOR U1751 ( .A(n2998), .B(n2997), .Z(n2999) );
  XNOR U1752 ( .A(n14108), .B(n14109), .Z(n14433) );
  XOR U1753 ( .A(n14092), .B(n14093), .Z(n14115) );
  XNOR U1754 ( .A(n12500), .B(n12501), .Z(n815) );
  XNOR U1755 ( .A(n12499), .B(n815), .Z(n12821) );
  NAND U1756 ( .A(n13118), .B(n13121), .Z(n816) );
  XOR U1757 ( .A(n13118), .B(n13121), .Z(n817) );
  NANDN U1758 ( .A(n13119), .B(n817), .Z(n818) );
  NAND U1759 ( .A(n816), .B(n818), .Z(n12892) );
  NAND U1760 ( .A(n13464), .B(n13467), .Z(n819) );
  XOR U1761 ( .A(n13464), .B(n13467), .Z(n820) );
  NANDN U1762 ( .A(n13465), .B(n820), .Z(n821) );
  NAND U1763 ( .A(n819), .B(n821), .Z(n13134) );
  XOR U1764 ( .A(n12908), .B(n12909), .Z(n822) );
  XNOR U1765 ( .A(n12907), .B(n822), .Z(n13047) );
  XNOR U1766 ( .A(n12518), .B(n12519), .Z(n823) );
  XNOR U1767 ( .A(n12517), .B(n823), .Z(n12817) );
  XNOR U1768 ( .A(n12921), .B(n12922), .Z(n824) );
  XNOR U1769 ( .A(n12923), .B(n824), .Z(n13045) );
  XNOR U1770 ( .A(n12935), .B(n12936), .Z(n13172) );
  XNOR U1771 ( .A(n3547), .B(n3548), .Z(n3800) );
  XNOR U1772 ( .A(n3314), .B(n3315), .Z(n3556) );
  XNOR U1773 ( .A(n3032), .B(n3031), .Z(n3034) );
  XNOR U1774 ( .A(n13761), .B(n13762), .Z(n14131) );
  XNOR U1775 ( .A(n12882), .B(n12883), .Z(n13114) );
  NAND U1776 ( .A(n13448), .B(n13451), .Z(n825) );
  XOR U1777 ( .A(n13448), .B(n13451), .Z(n826) );
  NANDN U1778 ( .A(n13449), .B(n826), .Z(n827) );
  NAND U1779 ( .A(n825), .B(n827), .Z(n13123) );
  XNOR U1780 ( .A(n13155), .B(n13156), .Z(n13487) );
  XNOR U1781 ( .A(n12928), .B(n12929), .Z(n13167) );
  XNOR U1782 ( .A(n13169), .B(n13170), .Z(n13505) );
  XNOR U1783 ( .A(n12940), .B(n12941), .Z(n828) );
  XNOR U1784 ( .A(n12939), .B(n828), .Z(n13042) );
  XNOR U1785 ( .A(n12962), .B(n12963), .Z(n829) );
  XNOR U1786 ( .A(n12961), .B(n829), .Z(n13038) );
  XNOR U1787 ( .A(n3020), .B(n3019), .Z(n3021) );
  XNOR U1788 ( .A(n3050), .B(n3049), .Z(n3041) );
  XNOR U1789 ( .A(n13767), .B(n13768), .Z(n14136) );
  XNOR U1790 ( .A(n13423), .B(n13424), .Z(n13782) );
  NAND U1791 ( .A(n14196), .B(n14199), .Z(n830) );
  XOR U1792 ( .A(n14196), .B(n14199), .Z(n831) );
  NANDN U1793 ( .A(n14197), .B(n831), .Z(n832) );
  NAND U1794 ( .A(n830), .B(n832), .Z(n13824) );
  XNOR U1795 ( .A(n13361), .B(n13362), .Z(n13867) );
  XOR U1796 ( .A(n13886), .B(n13887), .Z(n833) );
  NANDN U1797 ( .A(n13888), .B(n833), .Z(n834) );
  NAND U1798 ( .A(n13886), .B(n13887), .Z(n835) );
  AND U1799 ( .A(n834), .B(n835), .Z(n13537) );
  XNOR U1800 ( .A(n14248), .B(n14249), .Z(n14250) );
  NAND U1801 ( .A(n13211), .B(n13214), .Z(n836) );
  XOR U1802 ( .A(n13211), .B(n13214), .Z(n837) );
  NANDN U1803 ( .A(n13212), .B(n837), .Z(n838) );
  NAND U1804 ( .A(n836), .B(n838), .Z(n12975) );
  XOR U1805 ( .A(n11179), .B(n11180), .Z(n839) );
  NANDN U1806 ( .A(n11182), .B(n839), .Z(n840) );
  NAND U1807 ( .A(n11179), .B(n11180), .Z(n841) );
  AND U1808 ( .A(n840), .B(n841), .Z(n11184) );
  XNOR U1809 ( .A(n3559), .B(n3560), .Z(n3811) );
  XOR U1810 ( .A(n3326), .B(n3327), .Z(n3568) );
  XNOR U1811 ( .A(n2995), .B(n2996), .Z(n3331) );
  XNOR U1812 ( .A(n3062), .B(n3061), .Z(n3063) );
  XNOR U1813 ( .A(n14126), .B(n14127), .Z(n14453) );
  XNOR U1814 ( .A(n13775), .B(n13776), .Z(n14149) );
  XNOR U1815 ( .A(n14142), .B(n14143), .Z(n14467) );
  NAND U1816 ( .A(n14511), .B(n14514), .Z(n842) );
  XOR U1817 ( .A(n14511), .B(n14514), .Z(n843) );
  NANDN U1818 ( .A(n14512), .B(n843), .Z(n844) );
  NAND U1819 ( .A(n842), .B(n844), .Z(n14194) );
  XOR U1820 ( .A(n13483), .B(n13484), .Z(n845) );
  XNOR U1821 ( .A(n13482), .B(n845), .Z(n13715) );
  XOR U1822 ( .A(n14228), .B(n14230), .Z(n846) );
  NANDN U1823 ( .A(n14229), .B(n846), .Z(n847) );
  NAND U1824 ( .A(n14228), .B(n14230), .Z(n848) );
  AND U1825 ( .A(n847), .B(n848), .Z(n13861) );
  XNOR U1826 ( .A(n13512), .B(n13513), .Z(n13710) );
  XNOR U1827 ( .A(n13889), .B(n13890), .Z(n14074) );
  NAND U1828 ( .A(n12983), .B(n12985), .Z(n849) );
  XOR U1829 ( .A(n12983), .B(n12985), .Z(n850) );
  NANDN U1830 ( .A(n12982), .B(n850), .Z(n851) );
  NAND U1831 ( .A(n849), .B(n851), .Z(n12597) );
  XNOR U1832 ( .A(n3098), .B(n3097), .Z(n3100) );
  XNOR U1833 ( .A(n14450), .B(n14451), .Z(n14825) );
  XNOR U1834 ( .A(n14820), .B(n14821), .Z(n15104) );
  XNOR U1835 ( .A(n13789), .B(n13790), .Z(n14160) );
  XNOR U1836 ( .A(n13437), .B(n13438), .Z(n852) );
  XNOR U1837 ( .A(n13436), .B(n852), .Z(n13724) );
  XOR U1838 ( .A(n14244), .B(n14245), .Z(n853) );
  XNOR U1839 ( .A(n14243), .B(n853), .Z(n14390) );
  XNOR U1840 ( .A(n3816), .B(n3817), .Z(n4075) );
  XNOR U1841 ( .A(n3571), .B(n3572), .Z(n3824) );
  XOR U1842 ( .A(n3076), .B(n3075), .Z(n3345) );
  XNOR U1843 ( .A(n3106), .B(n3105), .Z(n3107) );
  XNOR U1844 ( .A(n14214), .B(n14215), .Z(n14398) );
  XOR U1845 ( .A(n14082), .B(n14083), .Z(n14535) );
  NAND U1846 ( .A(n14927), .B(n14930), .Z(n854) );
  XOR U1847 ( .A(n14927), .B(n14930), .Z(n855) );
  NANDN U1848 ( .A(n14928), .B(n855), .Z(n856) );
  NAND U1849 ( .A(n854), .B(n856), .Z(n14550) );
  XNOR U1850 ( .A(n14237), .B(n14238), .Z(n14393) );
  NAND U1851 ( .A(n15264), .B(n15267), .Z(n857) );
  XOR U1852 ( .A(n15264), .B(n15267), .Z(n858) );
  NANDN U1853 ( .A(n15265), .B(n858), .Z(n859) );
  NAND U1854 ( .A(n857), .B(n859), .Z(n14944) );
  XOR U1855 ( .A(n14579), .B(n14580), .Z(n860) );
  NANDN U1856 ( .A(n14581), .B(n860), .Z(n861) );
  NAND U1857 ( .A(n14579), .B(n14580), .Z(n862) );
  AND U1858 ( .A(n861), .B(n862), .Z(n14268) );
  XNOR U1859 ( .A(n13904), .B(n13905), .Z(n863) );
  XNOR U1860 ( .A(n13903), .B(n863), .Z(n14073) );
  XOR U1861 ( .A(n14964), .B(n14966), .Z(n864) );
  NANDN U1862 ( .A(n14965), .B(n864), .Z(n865) );
  NAND U1863 ( .A(n14964), .B(n14966), .Z(n866) );
  AND U1864 ( .A(n865), .B(n866), .Z(n14583) );
  XOR U1865 ( .A(n4593), .B(n4594), .Z(n4867) );
  XNOR U1866 ( .A(n4073), .B(n4074), .Z(n4338) );
  XNOR U1867 ( .A(n3118), .B(n3117), .Z(n3120) );
  XNOR U1868 ( .A(n10131), .B(n10130), .Z(n10133) );
  XNOR U1869 ( .A(n14480), .B(n14481), .Z(n14855) );
  NAND U1870 ( .A(n14406), .B(n14409), .Z(n867) );
  XOR U1871 ( .A(n14406), .B(n14409), .Z(n868) );
  NANDN U1872 ( .A(n14407), .B(n868), .Z(n869) );
  NAND U1873 ( .A(n867), .B(n869), .Z(n14506) );
  XNOR U1874 ( .A(n14528), .B(n14529), .Z(n870) );
  XNOR U1875 ( .A(n14527), .B(n870), .Z(n14769) );
  NAND U1876 ( .A(n15224), .B(n15227), .Z(n871) );
  XOR U1877 ( .A(n15224), .B(n15227), .Z(n872) );
  NANDN U1878 ( .A(n15225), .B(n872), .Z(n873) );
  NAND U1879 ( .A(n871), .B(n873), .Z(n14901) );
  NAND U1880 ( .A(n15248), .B(n15251), .Z(n874) );
  XOR U1881 ( .A(n15248), .B(n15251), .Z(n875) );
  NANDN U1882 ( .A(n15249), .B(n875), .Z(n876) );
  NAND U1883 ( .A(n874), .B(n876), .Z(n14925) );
  NAND U1884 ( .A(n15630), .B(n15633), .Z(n877) );
  XOR U1885 ( .A(n15630), .B(n15633), .Z(n878) );
  NANDN U1886 ( .A(n15631), .B(n878), .Z(n879) );
  NAND U1887 ( .A(n877), .B(n879), .Z(n15269) );
  NAND U1888 ( .A(n15282), .B(n15285), .Z(n880) );
  XOR U1889 ( .A(n15282), .B(n15285), .Z(n881) );
  NANDN U1890 ( .A(n15283), .B(n881), .Z(n882) );
  NAND U1891 ( .A(n880), .B(n882), .Z(n14962) );
  NAND U1892 ( .A(n13354), .B(n13353), .Z(n883) );
  NANDN U1893 ( .A(n13227), .B(n13228), .Z(n884) );
  AND U1894 ( .A(n883), .B(n884), .Z(n13232) );
  XNOR U1895 ( .A(n3350), .B(n3351), .Z(n3592) );
  XNOR U1896 ( .A(n4868), .B(n4869), .Z(n5147) );
  XNOR U1897 ( .A(n4336), .B(n4337), .Z(n4605) );
  XNOR U1898 ( .A(n3583), .B(n3584), .Z(n3836) );
  XNOR U1899 ( .A(n3083), .B(n3084), .Z(n3355) );
  XNOR U1900 ( .A(n22689), .B(n22688), .Z(n22690) );
  XNOR U1901 ( .A(n14838), .B(n14839), .Z(n15166) );
  XNOR U1902 ( .A(n15095), .B(n15096), .Z(n15220) );
  NAND U1903 ( .A(n15614), .B(n15617), .Z(n885) );
  XOR U1904 ( .A(n15614), .B(n15617), .Z(n886) );
  NANDN U1905 ( .A(n15615), .B(n886), .Z(n887) );
  NAND U1906 ( .A(n885), .B(n887), .Z(n15253) );
  NAND U1907 ( .A(n15651), .B(n15654), .Z(n888) );
  XOR U1908 ( .A(n15651), .B(n15654), .Z(n889) );
  NANDN U1909 ( .A(n15652), .B(n889), .Z(n890) );
  NAND U1910 ( .A(n888), .B(n890), .Z(n15281) );
  XOR U1911 ( .A(n14593), .B(n14594), .Z(n14595) );
  XNOR U1912 ( .A(n5145), .B(n5146), .Z(n5433) );
  XNOR U1913 ( .A(n4603), .B(n4604), .Z(n4880) );
  XNOR U1914 ( .A(n4085), .B(n4086), .Z(n4349) );
  XNOR U1915 ( .A(n14850), .B(n14851), .Z(n15178) );
  XNOR U1916 ( .A(n14498), .B(n14499), .Z(n14779) );
  XNOR U1917 ( .A(n15599), .B(n15600), .Z(n15785) );
  XNOR U1918 ( .A(n15618), .B(n15619), .Z(n15781) );
  NAND U1919 ( .A(n15962), .B(n15965), .Z(n891) );
  XOR U1920 ( .A(n15962), .B(n15965), .Z(n892) );
  NANDN U1921 ( .A(n15963), .B(n892), .Z(n893) );
  NAND U1922 ( .A(n891), .B(n893), .Z(n15634) );
  NAND U1923 ( .A(n15299), .B(n15302), .Z(n894) );
  XOR U1924 ( .A(n15299), .B(n15302), .Z(n895) );
  NANDN U1925 ( .A(n15300), .B(n895), .Z(n896) );
  NAND U1926 ( .A(n894), .B(n896), .Z(n14980) );
  XNOR U1927 ( .A(n3842), .B(n3843), .Z(n4097) );
  XNOR U1928 ( .A(n5434), .B(n5435), .Z(n5728) );
  XNOR U1929 ( .A(n4878), .B(n4879), .Z(n5159) );
  XNOR U1930 ( .A(n4350), .B(n4351), .Z(n4618) );
  XNOR U1931 ( .A(n3595), .B(n3596), .Z(n3847) );
  XNOR U1932 ( .A(n22679), .B(n22678), .Z(n22673) );
  XNOR U1933 ( .A(n14862), .B(n14863), .Z(n15189) );
  NAND U1934 ( .A(n15562), .B(n15565), .Z(n897) );
  XOR U1935 ( .A(n15562), .B(n15565), .Z(n898) );
  NANDN U1936 ( .A(n15563), .B(n898), .Z(n899) );
  NAND U1937 ( .A(n897), .B(n899), .Z(n15199) );
  XOR U1938 ( .A(n15215), .B(n15216), .Z(n900) );
  XNOR U1939 ( .A(n15214), .B(n900), .Z(n15461) );
  NAND U1940 ( .A(n16322), .B(n16325), .Z(n901) );
  XOR U1941 ( .A(n16322), .B(n16325), .Z(n902) );
  NANDN U1942 ( .A(n16323), .B(n902), .Z(n903) );
  NAND U1943 ( .A(n901), .B(n903), .Z(n15961) );
  NAND U1944 ( .A(n16668), .B(n16671), .Z(n904) );
  XOR U1945 ( .A(n16668), .B(n16671), .Z(n905) );
  NANDN U1946 ( .A(n16669), .B(n905), .Z(n906) );
  NAND U1947 ( .A(n904), .B(n906), .Z(n16338) );
  XOR U1948 ( .A(n16348), .B(n16347), .Z(n907) );
  NANDN U1949 ( .A(n16346), .B(n907), .Z(n908) );
  NAND U1950 ( .A(n16348), .B(n16347), .Z(n909) );
  AND U1951 ( .A(n908), .B(n909), .Z(n15990) );
  XNOR U1952 ( .A(n15303), .B(n15304), .Z(n15446) );
  XNOR U1953 ( .A(n15668), .B(n15669), .Z(n15772) );
  NAND U1954 ( .A(n13576), .B(n13575), .Z(n910) );
  NANDN U1955 ( .A(n13241), .B(n13242), .Z(n911) );
  AND U1956 ( .A(n910), .B(n911), .Z(n13243) );
  NAND U1957 ( .A(n13574), .B(n13573), .Z(n912) );
  NANDN U1958 ( .A(n13929), .B(n13928), .Z(n913) );
  AND U1959 ( .A(n912), .B(n913), .Z(n13578) );
  NAND U1960 ( .A(n12795), .B(n12794), .Z(n914) );
  NANDN U1961 ( .A(n13245), .B(n13246), .Z(n915) );
  NAND U1962 ( .A(n914), .B(n915), .Z(n12999) );
  XNOR U1963 ( .A(n5725), .B(n5726), .Z(n6025) );
  XNOR U1964 ( .A(n5157), .B(n5158), .Z(n5446) );
  XNOR U1965 ( .A(n4615), .B(n4616), .Z(n4891) );
  XNOR U1966 ( .A(n22665), .B(n22664), .Z(n22666) );
  XOR U1967 ( .A(n15204), .B(n15205), .Z(n916) );
  XNOR U1968 ( .A(n15203), .B(n916), .Z(n15465) );
  XOR U1969 ( .A(n16292), .B(n16293), .Z(n917) );
  NANDN U1970 ( .A(n16295), .B(n917), .Z(n918) );
  NAND U1971 ( .A(n16292), .B(n16293), .Z(n919) );
  AND U1972 ( .A(n918), .B(n919), .Z(n16302) );
  XOR U1973 ( .A(n15773), .B(n15774), .Z(n16359) );
  XNOR U1974 ( .A(n5444), .B(n5445), .Z(n5739) );
  XNOR U1975 ( .A(n4892), .B(n4893), .Z(n5172) );
  XNOR U1976 ( .A(n10167), .B(n10166), .Z(n10169) );
  XNOR U1977 ( .A(n22659), .B(n22658), .Z(n22660) );
  NAND U1978 ( .A(n16256), .B(n16259), .Z(n920) );
  XOR U1979 ( .A(n16256), .B(n16259), .Z(n921) );
  NANDN U1980 ( .A(n16257), .B(n921), .Z(n922) );
  NAND U1981 ( .A(n920), .B(n922), .Z(n15890) );
  XNOR U1982 ( .A(n15791), .B(n15792), .Z(n16273) );
  XNOR U1983 ( .A(n16310), .B(n16311), .Z(n923) );
  XNOR U1984 ( .A(n16309), .B(n923), .Z(n16480) );
  NAND U1985 ( .A(n17024), .B(n17027), .Z(n924) );
  XOR U1986 ( .A(n17024), .B(n17027), .Z(n925) );
  NANDN U1987 ( .A(n17025), .B(n925), .Z(n926) );
  NAND U1988 ( .A(n924), .B(n926), .Z(n16665) );
  NANDN U1989 ( .A(n17052), .B(n16686), .Z(n927) );
  NAND U1990 ( .A(n17052), .B(n17053), .Z(n928) );
  NANDN U1991 ( .A(n17051), .B(n928), .Z(n929) );
  NAND U1992 ( .A(n927), .B(n929), .Z(n16692) );
  XNOR U1993 ( .A(n16363), .B(n16364), .Z(n16470) );
  XOR U1994 ( .A(n15684), .B(n15681), .Z(n930) );
  NANDN U1995 ( .A(n15682), .B(n930), .Z(n931) );
  NAND U1996 ( .A(n15684), .B(n15681), .Z(n932) );
  AND U1997 ( .A(n931), .B(n932), .Z(n15442) );
  XNOR U1998 ( .A(n16009), .B(n16010), .Z(n16380) );
  XNOR U1999 ( .A(n6032), .B(n6033), .Z(n6336) );
  XNOR U2000 ( .A(n5737), .B(n5738), .Z(n6038) );
  XNOR U2001 ( .A(n5169), .B(n5170), .Z(n5456) );
  XNOR U2002 ( .A(n10173), .B(n10172), .Z(n10175) );
  NAND U2003 ( .A(n16593), .B(n16596), .Z(n933) );
  XOR U2004 ( .A(n16593), .B(n16596), .Z(n934) );
  NANDN U2005 ( .A(n16594), .B(n934), .Z(n935) );
  NAND U2006 ( .A(n933), .B(n935), .Z(n16255) );
  NAND U2007 ( .A(n16607), .B(n16610), .Z(n936) );
  XOR U2008 ( .A(n16607), .B(n16610), .Z(n937) );
  NANDN U2009 ( .A(n16608), .B(n937), .Z(n938) );
  NAND U2010 ( .A(n936), .B(n938), .Z(n16271) );
  XOR U2011 ( .A(n16287), .B(n16288), .Z(n939) );
  XNOR U2012 ( .A(n16286), .B(n939), .Z(n16488) );
  XNOR U2013 ( .A(n16147), .B(n16148), .Z(n16647) );
  NAND U2014 ( .A(n17363), .B(n17366), .Z(n940) );
  XOR U2015 ( .A(n17363), .B(n17366), .Z(n941) );
  NANDN U2016 ( .A(n17364), .B(n941), .Z(n942) );
  NAND U2017 ( .A(n940), .B(n942), .Z(n17028) );
  XNOR U2018 ( .A(n17043), .B(n17044), .Z(n17162) );
  NAND U2019 ( .A(n17067), .B(n17070), .Z(n943) );
  XOR U2020 ( .A(n17067), .B(n17070), .Z(n944) );
  NANDN U2021 ( .A(n17068), .B(n944), .Z(n945) );
  NAND U2022 ( .A(n943), .B(n945), .Z(n16708) );
  XNOR U2023 ( .A(n4902), .B(n4903), .Z(n5184) );
  XNOR U2024 ( .A(n6333), .B(n6334), .Z(n6645) );
  XNOR U2025 ( .A(n5458), .B(n5459), .Z(n5749) );
  XNOR U2026 ( .A(n10125), .B(n10124), .Z(n10127) );
  NAND U2027 ( .A(n16941), .B(n16944), .Z(n946) );
  XOR U2028 ( .A(n16941), .B(n16944), .Z(n947) );
  NANDN U2029 ( .A(n16942), .B(n947), .Z(n948) );
  NAND U2030 ( .A(n946), .B(n948), .Z(n16592) );
  NAND U2031 ( .A(n16959), .B(n16962), .Z(n949) );
  XOR U2032 ( .A(n16959), .B(n16962), .Z(n950) );
  NANDN U2033 ( .A(n16960), .B(n950), .Z(n951) );
  NAND U2034 ( .A(n949), .B(n951), .Z(n16612) );
  XOR U2035 ( .A(n16639), .B(n16640), .Z(n952) );
  XNOR U2036 ( .A(n16638), .B(n952), .Z(n17003) );
  XOR U2037 ( .A(n16988), .B(n16990), .Z(n953) );
  NAND U2038 ( .A(n953), .B(n16989), .Z(n954) );
  NAND U2039 ( .A(n16988), .B(n16990), .Z(n955) );
  AND U2040 ( .A(n954), .B(n955), .Z(n16993) );
  XNOR U2041 ( .A(n16825), .B(n16826), .Z(n17400) );
  NAND U2042 ( .A(n15002), .B(n15001), .Z(n956) );
  NANDN U2043 ( .A(n15324), .B(n15323), .Z(n957) );
  AND U2044 ( .A(n956), .B(n957), .Z(n15006) );
  NAND U2045 ( .A(n14309), .B(n14308), .Z(n958) );
  NANDN U2046 ( .A(n14626), .B(n14625), .Z(n959) );
  AND U2047 ( .A(n958), .B(n959), .Z(n14313) );
  NAND U2048 ( .A(n13592), .B(n13591), .Z(n960) );
  NANDN U2049 ( .A(n13261), .B(n13262), .Z(n961) );
  AND U2050 ( .A(n960), .B(n961), .Z(n13263) );
  NAND U2051 ( .A(n13590), .B(n13589), .Z(n962) );
  NANDN U2052 ( .A(n13953), .B(n13952), .Z(n963) );
  AND U2053 ( .A(n962), .B(n963), .Z(n13594) );
  NAND U2054 ( .A(n12787), .B(n12786), .Z(n964) );
  NANDN U2055 ( .A(n13265), .B(n13266), .Z(n965) );
  NAND U2056 ( .A(n964), .B(n965), .Z(n13007) );
  XOR U2057 ( .A(n6959), .B(n6960), .Z(n7008) );
  XNOR U2058 ( .A(n5181), .B(n5182), .Z(n5469) );
  XNOR U2059 ( .A(n6646), .B(n6647), .Z(n6687) );
  XNOR U2060 ( .A(n6042), .B(n6043), .Z(n6347) );
  XNOR U2061 ( .A(n5751), .B(n5752), .Z(n6048) );
  XNOR U2062 ( .A(n10179), .B(n10178), .Z(n10181) );
  NAND U2063 ( .A(n17275), .B(n17278), .Z(n966) );
  XOR U2064 ( .A(n17275), .B(n17278), .Z(n967) );
  NANDN U2065 ( .A(n17276), .B(n967), .Z(n968) );
  NAND U2066 ( .A(n966), .B(n968), .Z(n16946) );
  NAND U2067 ( .A(n17291), .B(n17294), .Z(n969) );
  XOR U2068 ( .A(n17291), .B(n17294), .Z(n970) );
  NANDN U2069 ( .A(n17292), .B(n970), .Z(n971) );
  NAND U2070 ( .A(n969), .B(n971), .Z(n16958) );
  NAND U2071 ( .A(n17309), .B(n17312), .Z(n972) );
  XOR U2072 ( .A(n17309), .B(n17312), .Z(n973) );
  NANDN U2073 ( .A(n17310), .B(n973), .Z(n974) );
  NAND U2074 ( .A(n972), .B(n974), .Z(n16974) );
  XOR U2075 ( .A(n16626), .B(n16627), .Z(n975) );
  XNOR U2076 ( .A(n16625), .B(n975), .Z(n16837) );
  XOR U2077 ( .A(n17378), .B(n17379), .Z(n976) );
  XNOR U2078 ( .A(n17377), .B(n976), .Z(n17528) );
  XNOR U2079 ( .A(n17157), .B(n17158), .Z(n17758) );
  NAND U2080 ( .A(n18074), .B(n18077), .Z(n977) );
  XOR U2081 ( .A(n18074), .B(n18077), .Z(n978) );
  NANDN U2082 ( .A(n18075), .B(n978), .Z(n979) );
  NAND U2083 ( .A(n977), .B(n979), .Z(n17760) );
  NAND U2084 ( .A(n17764), .B(n17767), .Z(n980) );
  XOR U2085 ( .A(n17764), .B(n17767), .Z(n981) );
  NANDN U2086 ( .A(n17765), .B(n981), .Z(n982) );
  NAND U2087 ( .A(n980), .B(n982), .Z(n17412) );
  XNOR U2088 ( .A(n6345), .B(n6346), .Z(n6658) );
  XNOR U2089 ( .A(n10185), .B(n10184), .Z(n10187) );
  NAND U2090 ( .A(n17645), .B(n17648), .Z(n983) );
  XOR U2091 ( .A(n17645), .B(n17648), .Z(n984) );
  NANDN U2092 ( .A(n17646), .B(n984), .Z(n985) );
  NAND U2093 ( .A(n983), .B(n985), .Z(n17280) );
  NAND U2094 ( .A(n17661), .B(n17664), .Z(n986) );
  XOR U2095 ( .A(n17661), .B(n17664), .Z(n987) );
  NANDN U2096 ( .A(n17662), .B(n987), .Z(n988) );
  NAND U2097 ( .A(n986), .B(n988), .Z(n17296) );
  NAND U2098 ( .A(n17679), .B(n17682), .Z(n989) );
  XOR U2099 ( .A(n17679), .B(n17682), .Z(n990) );
  NANDN U2100 ( .A(n17680), .B(n990), .Z(n991) );
  NAND U2101 ( .A(n989), .B(n991), .Z(n17314) );
  XOR U2102 ( .A(n17339), .B(n17340), .Z(n992) );
  NANDN U2103 ( .A(n17342), .B(n992), .Z(n993) );
  NAND U2104 ( .A(n17339), .B(n17340), .Z(n994) );
  AND U2105 ( .A(n993), .B(n994), .Z(n17349) );
  XNOR U2106 ( .A(n17529), .B(n17530), .Z(n18052) );
  XNOR U2107 ( .A(n17727), .B(n17728), .Z(n18050) );
  NAND U2108 ( .A(n18409), .B(n18412), .Z(n995) );
  XOR U2109 ( .A(n18409), .B(n18412), .Z(n996) );
  NANDN U2110 ( .A(n18410), .B(n996), .Z(n997) );
  NAND U2111 ( .A(n995), .B(n997), .Z(n18064) );
  XOR U2112 ( .A(n18068), .B(n18069), .Z(n998) );
  XNOR U2113 ( .A(n18067), .B(n998), .Z(n18189) );
  XOR U2114 ( .A(n17415), .B(n17416), .Z(n17417) );
  NAND U2115 ( .A(n15700), .B(n15699), .Z(n999) );
  NANDN U2116 ( .A(n16026), .B(n16025), .Z(n1000) );
  AND U2117 ( .A(n999), .B(n1000), .Z(n15704) );
  XNOR U2118 ( .A(n7288), .B(n7289), .Z(n7616) );
  XNOR U2119 ( .A(n6656), .B(n6657), .Z(n6975) );
  XNOR U2120 ( .A(n10191), .B(n10190), .Z(n10193) );
  NAND U2121 ( .A(n17968), .B(n17971), .Z(n1001) );
  XOR U2122 ( .A(n17968), .B(n17971), .Z(n1002) );
  NANDN U2123 ( .A(n17969), .B(n1002), .Z(n1003) );
  NAND U2124 ( .A(n1001), .B(n1003), .Z(n17650) );
  NAND U2125 ( .A(n17984), .B(n17987), .Z(n1004) );
  XOR U2126 ( .A(n17984), .B(n17987), .Z(n1005) );
  NANDN U2127 ( .A(n17985), .B(n1005), .Z(n1006) );
  NAND U2128 ( .A(n1004), .B(n1006), .Z(n17666) );
  NAND U2129 ( .A(n18000), .B(n18003), .Z(n1007) );
  XOR U2130 ( .A(n18000), .B(n18003), .Z(n1008) );
  NANDN U2131 ( .A(n18001), .B(n1008), .Z(n1009) );
  NAND U2132 ( .A(n1007), .B(n1009), .Z(n17678) );
  NAND U2133 ( .A(n18016), .B(n18019), .Z(n1010) );
  XOR U2134 ( .A(n18016), .B(n18019), .Z(n1011) );
  NANDN U2135 ( .A(n18017), .B(n1011), .Z(n1012) );
  NAND U2136 ( .A(n1010), .B(n1012), .Z(n17698) );
  XOR U2137 ( .A(n17326), .B(n17327), .Z(n1013) );
  XNOR U2138 ( .A(n17325), .B(n1013), .Z(n17538) );
  XOR U2139 ( .A(n17711), .B(n17712), .Z(n1014) );
  XNOR U2140 ( .A(n17710), .B(n1014), .Z(n17857) );
  XOR U2141 ( .A(n18195), .B(n18194), .Z(n1015) );
  NANDN U2142 ( .A(n18197), .B(n1015), .Z(n1016) );
  NAND U2143 ( .A(n18195), .B(n18194), .Z(n1017) );
  AND U2144 ( .A(n1016), .B(n1017), .Z(n18402) );
  XNOR U2145 ( .A(n18419), .B(n18420), .Z(n18740) );
  NANDN U2146 ( .A(n18431), .B(n18753), .Z(n1018) );
  OR U2147 ( .A(n18753), .B(n18752), .Z(n1019) );
  NANDN U2148 ( .A(n18755), .B(n1019), .Z(n1020) );
  NAND U2149 ( .A(n1018), .B(n1020), .Z(n18436) );
  XOR U2150 ( .A(n18441), .B(n18443), .Z(n1021) );
  NANDN U2151 ( .A(n18442), .B(n1021), .Z(n1022) );
  NAND U2152 ( .A(n18441), .B(n18443), .Z(n1023) );
  AND U2153 ( .A(n1022), .B(n1023), .Z(n18091) );
  NAND U2154 ( .A(n15018), .B(n15017), .Z(n1024) );
  NANDN U2155 ( .A(n15348), .B(n15347), .Z(n1025) );
  AND U2156 ( .A(n1024), .B(n1025), .Z(n15022) );
  XNOR U2157 ( .A(n7292), .B(n7293), .Z(n7621) );
  XNOR U2158 ( .A(n6973), .B(n6974), .Z(n7298) );
  XNOR U2159 ( .A(n6357), .B(n6358), .Z(n6670) );
  XNOR U2160 ( .A(n10119), .B(n10118), .Z(n10121) );
  NAND U2161 ( .A(n18312), .B(n18315), .Z(n1026) );
  XOR U2162 ( .A(n18312), .B(n18315), .Z(n1027) );
  NANDN U2163 ( .A(n18313), .B(n1027), .Z(n1028) );
  NAND U2164 ( .A(n1026), .B(n1028), .Z(n17973) );
  XOR U2165 ( .A(n18333), .B(n18330), .Z(n1029) );
  NANDN U2166 ( .A(n18331), .B(n1029), .Z(n1030) );
  NAND U2167 ( .A(n18333), .B(n18330), .Z(n1031) );
  AND U2168 ( .A(n1030), .B(n1031), .Z(n17989) );
  NAND U2169 ( .A(n18346), .B(n18349), .Z(n1032) );
  XOR U2170 ( .A(n18346), .B(n18349), .Z(n1033) );
  NANDN U2171 ( .A(n18347), .B(n1033), .Z(n1034) );
  NAND U2172 ( .A(n1032), .B(n1034), .Z(n18005) );
  NAND U2173 ( .A(n18362), .B(n18365), .Z(n1035) );
  XOR U2174 ( .A(n18362), .B(n18365), .Z(n1036) );
  NANDN U2175 ( .A(n18363), .B(n1036), .Z(n1037) );
  NAND U2176 ( .A(n1035), .B(n1037), .Z(n18021) );
  XNOR U2177 ( .A(n18756), .B(n18757), .Z(n19103) );
  NAND U2178 ( .A(n14325), .B(n14324), .Z(n1038) );
  NANDN U2179 ( .A(n14650), .B(n14649), .Z(n1039) );
  AND U2180 ( .A(n1038), .B(n1039), .Z(n14329) );
  NAND U2181 ( .A(n13608), .B(n13607), .Z(n1040) );
  NANDN U2182 ( .A(n13281), .B(n13282), .Z(n1041) );
  AND U2183 ( .A(n1040), .B(n1041), .Z(n13283) );
  NAND U2184 ( .A(n13606), .B(n13605), .Z(n1042) );
  NANDN U2185 ( .A(n13977), .B(n13976), .Z(n1043) );
  AND U2186 ( .A(n1042), .B(n1043), .Z(n13610) );
  NAND U2187 ( .A(n12779), .B(n12778), .Z(n1044) );
  NANDN U2188 ( .A(n13285), .B(n13286), .Z(n1045) );
  NAND U2189 ( .A(n1044), .B(n1045), .Z(n13015) );
  XNOR U2190 ( .A(n6365), .B(n6366), .Z(n6674) );
  XNOR U2191 ( .A(n6668), .B(n6669), .Z(n6987) );
  XNOR U2192 ( .A(n10197), .B(n10196), .Z(n10199) );
  XOR U2193 ( .A(n18624), .B(n18621), .Z(n1046) );
  NANDN U2194 ( .A(n18622), .B(n1046), .Z(n1047) );
  NAND U2195 ( .A(n18624), .B(n18621), .Z(n1048) );
  AND U2196 ( .A(n1047), .B(n1048), .Z(n18317) );
  XOR U2197 ( .A(n18640), .B(n18637), .Z(n1049) );
  NANDN U2198 ( .A(n18638), .B(n1049), .Z(n1050) );
  NAND U2199 ( .A(n18640), .B(n18637), .Z(n1051) );
  AND U2200 ( .A(n1050), .B(n1051), .Z(n18335) );
  NAND U2201 ( .A(n18653), .B(n18656), .Z(n1052) );
  XOR U2202 ( .A(n18653), .B(n18656), .Z(n1053) );
  NANDN U2203 ( .A(n18654), .B(n1053), .Z(n1054) );
  NAND U2204 ( .A(n1052), .B(n1054), .Z(n18351) );
  NAND U2205 ( .A(n18669), .B(n18672), .Z(n1055) );
  XOR U2206 ( .A(n18669), .B(n18672), .Z(n1056) );
  NANDN U2207 ( .A(n18670), .B(n1056), .Z(n1057) );
  NAND U2208 ( .A(n1055), .B(n1057), .Z(n18367) );
  XNOR U2209 ( .A(n18034), .B(n18035), .Z(n1058) );
  XNOR U2210 ( .A(n18036), .B(n1058), .Z(n18202) );
  NAND U2211 ( .A(n18685), .B(n18688), .Z(n1059) );
  XOR U2212 ( .A(n18685), .B(n18688), .Z(n1060) );
  NANDN U2213 ( .A(n18686), .B(n1060), .Z(n1061) );
  NAND U2214 ( .A(n1059), .B(n1061), .Z(n18383) );
  XOR U2215 ( .A(n18394), .B(n18395), .Z(n1062) );
  XNOR U2216 ( .A(n18393), .B(n1062), .Z(n18506) );
  NAND U2217 ( .A(n19116), .B(n19119), .Z(n1063) );
  XOR U2218 ( .A(n19116), .B(n19119), .Z(n1064) );
  NANDN U2219 ( .A(n19117), .B(n1064), .Z(n1065) );
  NAND U2220 ( .A(n1063), .B(n1065), .Z(n18769) );
  XNOR U2221 ( .A(n7302), .B(n7303), .Z(n7632) );
  XNOR U2222 ( .A(n6985), .B(n6986), .Z(n7308) );
  XNOR U2223 ( .A(n10203), .B(n10202), .Z(n10205) );
  XNOR U2224 ( .A(n19550), .B(n19551), .Z(n19890) );
  NAND U2225 ( .A(n18954), .B(n18957), .Z(n1066) );
  XOR U2226 ( .A(n18954), .B(n18957), .Z(n1067) );
  NANDN U2227 ( .A(n18955), .B(n1067), .Z(n1068) );
  NAND U2228 ( .A(n1066), .B(n1068), .Z(n18626) );
  NAND U2229 ( .A(n18971), .B(n18973), .Z(n1069) );
  XOR U2230 ( .A(n18971), .B(n18973), .Z(n1070) );
  NANDN U2231 ( .A(n18970), .B(n1070), .Z(n1071) );
  NAND U2232 ( .A(n1069), .B(n1071), .Z(n18642) );
  NAND U2233 ( .A(n18989), .B(n18991), .Z(n1072) );
  XOR U2234 ( .A(n18989), .B(n18991), .Z(n1073) );
  NANDN U2235 ( .A(n18988), .B(n1073), .Z(n1074) );
  NAND U2236 ( .A(n1072), .B(n1074), .Z(n18658) );
  NAND U2237 ( .A(n19004), .B(n19007), .Z(n1075) );
  XOR U2238 ( .A(n19004), .B(n19007), .Z(n1076) );
  NANDN U2239 ( .A(n19005), .B(n1076), .Z(n1077) );
  NAND U2240 ( .A(n1075), .B(n1077), .Z(n18674) );
  NAND U2241 ( .A(n19022), .B(n19025), .Z(n1078) );
  XOR U2242 ( .A(n19022), .B(n19025), .Z(n1079) );
  NANDN U2243 ( .A(n19023), .B(n1079), .Z(n1080) );
  NAND U2244 ( .A(n1078), .B(n1080), .Z(n18690) );
  NAND U2245 ( .A(n19040), .B(n19043), .Z(n1081) );
  XOR U2246 ( .A(n19040), .B(n19043), .Z(n1082) );
  NANDN U2247 ( .A(n19041), .B(n1082), .Z(n1083) );
  NAND U2248 ( .A(n1081), .B(n1083), .Z(n18702) );
  XOR U2249 ( .A(n18726), .B(n18727), .Z(n1084) );
  XNOR U2250 ( .A(n18725), .B(n1084), .Z(n18841) );
  XNOR U2251 ( .A(n18836), .B(n18837), .Z(n19078) );
  XOR U2252 ( .A(n19099), .B(n19100), .Z(n1085) );
  XNOR U2253 ( .A(n19098), .B(n1085), .Z(n19168) );
  NAND U2254 ( .A(n19431), .B(n19434), .Z(n1086) );
  XOR U2255 ( .A(n19431), .B(n19434), .Z(n1087) );
  NANDN U2256 ( .A(n19432), .B(n1087), .Z(n1088) );
  NAND U2257 ( .A(n1086), .B(n1088), .Z(n19114) );
  NAND U2258 ( .A(n19775), .B(n19778), .Z(n1089) );
  XOR U2259 ( .A(n19775), .B(n19778), .Z(n1090) );
  NANDN U2260 ( .A(n19776), .B(n1090), .Z(n1091) );
  NAND U2261 ( .A(n1089), .B(n1091), .Z(n19436) );
  XNOR U2262 ( .A(n18495), .B(n18496), .Z(n18776) );
  XOR U2263 ( .A(n18460), .B(n18457), .Z(n1092) );
  NANDN U2264 ( .A(n18458), .B(n1092), .Z(n1093) );
  NAND U2265 ( .A(n18460), .B(n18457), .Z(n1094) );
  AND U2266 ( .A(n1093), .B(n1094), .Z(n18178) );
  NAND U2267 ( .A(n15716), .B(n15715), .Z(n1095) );
  NANDN U2268 ( .A(n16048), .B(n16047), .Z(n1096) );
  AND U2269 ( .A(n1095), .B(n1096), .Z(n15720) );
  XNOR U2270 ( .A(n7994), .B(n7995), .Z(n8299) );
  XNOR U2271 ( .A(n7633), .B(n7634), .Z(n7656) );
  XNOR U2272 ( .A(n10209), .B(n10208), .Z(n10211) );
  XNOR U2273 ( .A(n19887), .B(n19888), .Z(n20207) );
  NAND U2274 ( .A(n19293), .B(n19296), .Z(n1097) );
  XOR U2275 ( .A(n19293), .B(n19296), .Z(n1098) );
  NANDN U2276 ( .A(n19294), .B(n1098), .Z(n1099) );
  NAND U2277 ( .A(n1097), .B(n1099), .Z(n18959) );
  NAND U2278 ( .A(n19309), .B(n19312), .Z(n1100) );
  XOR U2279 ( .A(n19309), .B(n19312), .Z(n1101) );
  NANDN U2280 ( .A(n19310), .B(n1101), .Z(n1102) );
  NAND U2281 ( .A(n1100), .B(n1102), .Z(n18975) );
  XOR U2282 ( .A(n19330), .B(n19327), .Z(n1103) );
  NANDN U2283 ( .A(n19328), .B(n1103), .Z(n1104) );
  NAND U2284 ( .A(n19330), .B(n19327), .Z(n1105) );
  AND U2285 ( .A(n1104), .B(n1105), .Z(n18992) );
  NAND U2286 ( .A(n19343), .B(n19346), .Z(n1106) );
  XOR U2287 ( .A(n19343), .B(n19346), .Z(n1107) );
  NANDN U2288 ( .A(n19344), .B(n1107), .Z(n1108) );
  NAND U2289 ( .A(n1106), .B(n1108), .Z(n19009) );
  XOR U2290 ( .A(n19362), .B(n19359), .Z(n1109) );
  NANDN U2291 ( .A(n19360), .B(n1109), .Z(n1110) );
  NAND U2292 ( .A(n19362), .B(n19359), .Z(n1111) );
  AND U2293 ( .A(n1110), .B(n1111), .Z(n19027) );
  NAND U2294 ( .A(n19375), .B(n19378), .Z(n1112) );
  XOR U2295 ( .A(n19375), .B(n19378), .Z(n1113) );
  NANDN U2296 ( .A(n19376), .B(n1113), .Z(n1114) );
  NAND U2297 ( .A(n1112), .B(n1114), .Z(n19039) );
  NAND U2298 ( .A(n20100), .B(n20103), .Z(n1115) );
  XOR U2299 ( .A(n20100), .B(n20103), .Z(n1116) );
  NANDN U2300 ( .A(n20101), .B(n1116), .Z(n1117) );
  NAND U2301 ( .A(n1115), .B(n1117), .Z(n19779) );
  NAND U2302 ( .A(n15034), .B(n15033), .Z(n1118) );
  NANDN U2303 ( .A(n15372), .B(n15371), .Z(n1119) );
  AND U2304 ( .A(n1118), .B(n1119), .Z(n15038) );
  XNOR U2305 ( .A(n7992), .B(n7993), .Z(n8304) );
  XNOR U2306 ( .A(n10113), .B(n10112), .Z(n10115) );
  NAND U2307 ( .A(n20236), .B(n20237), .Z(n1120) );
  NANDN U2308 ( .A(n20567), .B(n20568), .Z(n1121) );
  AND U2309 ( .A(n1120), .B(n1121), .Z(n20241) );
  NAND U2310 ( .A(n19632), .B(n19635), .Z(n1122) );
  XOR U2311 ( .A(n19632), .B(n19635), .Z(n1123) );
  NANDN U2312 ( .A(n19633), .B(n1123), .Z(n1124) );
  NAND U2313 ( .A(n1122), .B(n1124), .Z(n19298) );
  NAND U2314 ( .A(n19648), .B(n19651), .Z(n1125) );
  XOR U2315 ( .A(n19648), .B(n19651), .Z(n1126) );
  NANDN U2316 ( .A(n19649), .B(n1126), .Z(n1127) );
  NAND U2317 ( .A(n1125), .B(n1127), .Z(n19314) );
  NAND U2318 ( .A(n19662), .B(n19665), .Z(n1128) );
  XOR U2319 ( .A(n19662), .B(n19665), .Z(n1129) );
  NANDN U2320 ( .A(n19663), .B(n1129), .Z(n1130) );
  NAND U2321 ( .A(n1128), .B(n1130), .Z(n19326) );
  XOR U2322 ( .A(n19683), .B(n19681), .Z(n1131) );
  NANDN U2323 ( .A(n19680), .B(n1131), .Z(n1132) );
  NAND U2324 ( .A(n19683), .B(n19681), .Z(n1133) );
  AND U2325 ( .A(n1132), .B(n1133), .Z(n19348) );
  XOR U2326 ( .A(n19699), .B(n19696), .Z(n1134) );
  NANDN U2327 ( .A(n19697), .B(n1134), .Z(n1135) );
  NAND U2328 ( .A(n19699), .B(n19696), .Z(n1136) );
  AND U2329 ( .A(n1135), .B(n1136), .Z(n19364) );
  NAND U2330 ( .A(n19712), .B(n19715), .Z(n1137) );
  XOR U2331 ( .A(n19712), .B(n19715), .Z(n1138) );
  NANDN U2332 ( .A(n19713), .B(n1138), .Z(n1139) );
  NAND U2333 ( .A(n1137), .B(n1139), .Z(n19380) );
  NAND U2334 ( .A(n19736), .B(n19739), .Z(n1140) );
  XOR U2335 ( .A(n19736), .B(n19739), .Z(n1141) );
  NANDN U2336 ( .A(n19737), .B(n1141), .Z(n1142) );
  NAND U2337 ( .A(n1140), .B(n1142), .Z(n19401) );
  XOR U2338 ( .A(n19173), .B(n19174), .Z(n1143) );
  XNOR U2339 ( .A(n19172), .B(n1143), .Z(n19746) );
  XNOR U2340 ( .A(n19447), .B(n19448), .Z(n19796) );
  NAND U2341 ( .A(n16420), .B(n16419), .Z(n1144) );
  NANDN U2342 ( .A(n16752), .B(n16751), .Z(n1145) );
  AND U2343 ( .A(n1144), .B(n1145), .Z(n16424) );
  NAND U2344 ( .A(n14341), .B(n14340), .Z(n1146) );
  NANDN U2345 ( .A(n14674), .B(n14673), .Z(n1147) );
  AND U2346 ( .A(n1146), .B(n1147), .Z(n14345) );
  NAND U2347 ( .A(n13624), .B(n13623), .Z(n1148) );
  NANDN U2348 ( .A(n13301), .B(n13302), .Z(n1149) );
  AND U2349 ( .A(n1148), .B(n1149), .Z(n13303) );
  NAND U2350 ( .A(n13622), .B(n13621), .Z(n1150) );
  NANDN U2351 ( .A(n14001), .B(n14000), .Z(n1151) );
  AND U2352 ( .A(n1150), .B(n1151), .Z(n13626) );
  NAND U2353 ( .A(n12771), .B(n12770), .Z(n1152) );
  NANDN U2354 ( .A(n13305), .B(n13306), .Z(n1153) );
  NAND U2355 ( .A(n1152), .B(n1153), .Z(n13023) );
  XNOR U2356 ( .A(n10215), .B(n10214), .Z(n10217) );
  XNOR U2357 ( .A(n20218), .B(n20219), .Z(n20544) );
  NAND U2358 ( .A(n19963), .B(n19966), .Z(n1154) );
  XOR U2359 ( .A(n19963), .B(n19966), .Z(n1155) );
  NANDN U2360 ( .A(n19964), .B(n1155), .Z(n1156) );
  NAND U2361 ( .A(n1154), .B(n1156), .Z(n19631) );
  NAND U2362 ( .A(n19981), .B(n19984), .Z(n1157) );
  XOR U2363 ( .A(n19981), .B(n19984), .Z(n1158) );
  NANDN U2364 ( .A(n19982), .B(n1158), .Z(n1159) );
  NAND U2365 ( .A(n1157), .B(n1159), .Z(n19647) );
  NAND U2366 ( .A(n19995), .B(n19998), .Z(n1160) );
  XOR U2367 ( .A(n19995), .B(n19998), .Z(n1161) );
  NANDN U2368 ( .A(n19996), .B(n1161), .Z(n1162) );
  NAND U2369 ( .A(n1160), .B(n1162), .Z(n19666) );
  NAND U2370 ( .A(n20011), .B(n20014), .Z(n1163) );
  XOR U2371 ( .A(n20011), .B(n20014), .Z(n1164) );
  NANDN U2372 ( .A(n20012), .B(n1164), .Z(n1165) );
  NAND U2373 ( .A(n1163), .B(n1165), .Z(n19678) );
  NAND U2374 ( .A(n20027), .B(n20030), .Z(n1166) );
  XOR U2375 ( .A(n20027), .B(n20030), .Z(n1167) );
  NANDN U2376 ( .A(n20028), .B(n1167), .Z(n1168) );
  NAND U2377 ( .A(n1166), .B(n1168), .Z(n19701) );
  NAND U2378 ( .A(n20043), .B(n20046), .Z(n1169) );
  XOR U2379 ( .A(n20043), .B(n20046), .Z(n1170) );
  NANDN U2380 ( .A(n20044), .B(n1170), .Z(n1171) );
  NAND U2381 ( .A(n1169), .B(n1171), .Z(n19717) );
  NAND U2382 ( .A(n20059), .B(n20062), .Z(n1172) );
  XOR U2383 ( .A(n20059), .B(n20062), .Z(n1173) );
  NANDN U2384 ( .A(n20060), .B(n1173), .Z(n1174) );
  NAND U2385 ( .A(n1172), .B(n1174), .Z(n19729) );
  NAND U2386 ( .A(n20075), .B(n20078), .Z(n1175) );
  XOR U2387 ( .A(n20075), .B(n20078), .Z(n1176) );
  NANDN U2388 ( .A(n20076), .B(n1176), .Z(n1177) );
  NAND U2389 ( .A(n1175), .B(n1177), .Z(n19838) );
  NAND U2390 ( .A(n18831), .B(n18829), .Z(n1178) );
  XOR U2391 ( .A(n18831), .B(n18829), .Z(n1179) );
  NANDN U2392 ( .A(n18828), .B(n1179), .Z(n1180) );
  NAND U2393 ( .A(n1178), .B(n1180), .Z(n18785) );
  NAND U2394 ( .A(n19131), .B(n19130), .Z(n1181) );
  NANDN U2395 ( .A(n19160), .B(n19161), .Z(n1182) );
  NAND U2396 ( .A(n1181), .B(n1182), .Z(n19452) );
  NAND U2397 ( .A(n18783), .B(n18782), .Z(n1183) );
  NAND U2398 ( .A(n18465), .B(n18466), .Z(n1184) );
  NAND U2399 ( .A(n1183), .B(n1184), .Z(n18787) );
  NAND U2400 ( .A(n15732), .B(n15731), .Z(n1185) );
  NANDN U2401 ( .A(n16072), .B(n16071), .Z(n1186) );
  AND U2402 ( .A(n1185), .B(n1186), .Z(n15736) );
  XNOR U2403 ( .A(n7978), .B(n7979), .Z(n8318) );
  XNOR U2404 ( .A(n20539), .B(n20540), .Z(n20883) );
  NAND U2405 ( .A(n20290), .B(n20293), .Z(n1187) );
  XOR U2406 ( .A(n20290), .B(n20293), .Z(n1188) );
  NANDN U2407 ( .A(n20291), .B(n1188), .Z(n1189) );
  NAND U2408 ( .A(n1187), .B(n1189), .Z(n19968) );
  XOR U2409 ( .A(n20311), .B(n20309), .Z(n1190) );
  NANDN U2410 ( .A(n20308), .B(n1190), .Z(n1191) );
  NAND U2411 ( .A(n20311), .B(n20309), .Z(n1192) );
  AND U2412 ( .A(n1191), .B(n1192), .Z(n19980) );
  NAND U2413 ( .A(n20322), .B(n20325), .Z(n1193) );
  XOR U2414 ( .A(n20322), .B(n20325), .Z(n1194) );
  NANDN U2415 ( .A(n20323), .B(n1194), .Z(n1195) );
  NAND U2416 ( .A(n1193), .B(n1195), .Z(n20000) );
  NAND U2417 ( .A(n20340), .B(n20343), .Z(n1196) );
  XOR U2418 ( .A(n20340), .B(n20343), .Z(n1197) );
  NANDN U2419 ( .A(n20341), .B(n1197), .Z(n1198) );
  NAND U2420 ( .A(n1196), .B(n1198), .Z(n20016) );
  NAND U2421 ( .A(n20360), .B(n20363), .Z(n1199) );
  XOR U2422 ( .A(n20360), .B(n20363), .Z(n1200) );
  NANDN U2423 ( .A(n20361), .B(n1200), .Z(n1201) );
  NAND U2424 ( .A(n1199), .B(n1201), .Z(n20032) );
  NAND U2425 ( .A(n20374), .B(n20377), .Z(n1202) );
  XOR U2426 ( .A(n20374), .B(n20377), .Z(n1203) );
  NANDN U2427 ( .A(n20375), .B(n1203), .Z(n1204) );
  NAND U2428 ( .A(n1202), .B(n1204), .Z(n20048) );
  NAND U2429 ( .A(n20390), .B(n20393), .Z(n1205) );
  XOR U2430 ( .A(n20390), .B(n20393), .Z(n1206) );
  NANDN U2431 ( .A(n20391), .B(n1206), .Z(n1207) );
  NAND U2432 ( .A(n1205), .B(n1207), .Z(n20064) );
  NAND U2433 ( .A(n20408), .B(n20411), .Z(n1208) );
  XOR U2434 ( .A(n20408), .B(n20411), .Z(n1209) );
  NANDN U2435 ( .A(n20409), .B(n1209), .Z(n1210) );
  NAND U2436 ( .A(n1208), .B(n1210), .Z(n20080) );
  XOR U2437 ( .A(n20092), .B(n20093), .Z(n1211) );
  XNOR U2438 ( .A(n20091), .B(n1211), .Z(n20171) );
  XNOR U2439 ( .A(n20115), .B(n20116), .Z(n1212) );
  XNOR U2440 ( .A(n20114), .B(n1212), .Z(n20163) );
  XOR U2441 ( .A(n8678), .B(n8679), .Z(n9008) );
  XNOR U2442 ( .A(n8319), .B(n8320), .Z(n8665) );
  XNOR U2443 ( .A(n7984), .B(n7985), .Z(n8324) );
  XNOR U2444 ( .A(n20880), .B(n20881), .Z(n21217) );
  XNOR U2445 ( .A(n20557), .B(n20558), .Z(n20896) );
  NAND U2446 ( .A(n20619), .B(n20622), .Z(n1213) );
  XOR U2447 ( .A(n20619), .B(n20622), .Z(n1214) );
  NANDN U2448 ( .A(n20620), .B(n1214), .Z(n1215) );
  NAND U2449 ( .A(n1213), .B(n1215), .Z(n20295) );
  NAND U2450 ( .A(n20635), .B(n20638), .Z(n1216) );
  XOR U2451 ( .A(n20635), .B(n20638), .Z(n1217) );
  NANDN U2452 ( .A(n20636), .B(n1217), .Z(n1218) );
  NAND U2453 ( .A(n1216), .B(n1218), .Z(n20306) );
  NAND U2454 ( .A(n20651), .B(n20654), .Z(n1219) );
  XOR U2455 ( .A(n20651), .B(n20654), .Z(n1220) );
  NANDN U2456 ( .A(n20652), .B(n1220), .Z(n1221) );
  NAND U2457 ( .A(n1219), .B(n1221), .Z(n20327) );
  XOR U2458 ( .A(n20670), .B(n20667), .Z(n1222) );
  NANDN U2459 ( .A(n20668), .B(n1222), .Z(n1223) );
  NAND U2460 ( .A(n20670), .B(n20667), .Z(n1224) );
  AND U2461 ( .A(n1223), .B(n1224), .Z(n20345) );
  XOR U2462 ( .A(n20688), .B(n20685), .Z(n1225) );
  NANDN U2463 ( .A(n20686), .B(n1225), .Z(n1226) );
  NAND U2464 ( .A(n20688), .B(n20685), .Z(n1227) );
  AND U2465 ( .A(n1226), .B(n1227), .Z(n20359) );
  NAND U2466 ( .A(n20699), .B(n20702), .Z(n1228) );
  XOR U2467 ( .A(n20699), .B(n20702), .Z(n1229) );
  NANDN U2468 ( .A(n20700), .B(n1229), .Z(n1230) );
  NAND U2469 ( .A(n1228), .B(n1230), .Z(n20379) );
  NAND U2470 ( .A(n20715), .B(n20718), .Z(n1231) );
  XOR U2471 ( .A(n20715), .B(n20718), .Z(n1232) );
  NANDN U2472 ( .A(n20716), .B(n1232), .Z(n1233) );
  NAND U2473 ( .A(n1231), .B(n1233), .Z(n20395) );
  NAND U2474 ( .A(n20734), .B(n20732), .Z(n1234) );
  XOR U2475 ( .A(n20734), .B(n20732), .Z(n1235) );
  NANDN U2476 ( .A(n20731), .B(n1235), .Z(n1236) );
  NAND U2477 ( .A(n1234), .B(n1236), .Z(n20413) );
  XOR U2478 ( .A(n20425), .B(n20426), .Z(n1237) );
  XNOR U2479 ( .A(n20424), .B(n1237), .Z(n20492) );
  NAND U2480 ( .A(n21101), .B(n21102), .Z(n1238) );
  XOR U2481 ( .A(n21101), .B(n21102), .Z(n1239) );
  NANDN U2482 ( .A(n21104), .B(n1239), .Z(n1240) );
  NAND U2483 ( .A(n1238), .B(n1240), .Z(n21109) );
  NAND U2484 ( .A(n21126), .B(n21129), .Z(n1241) );
  XOR U2485 ( .A(n21126), .B(n21129), .Z(n1242) );
  NANDN U2486 ( .A(n21127), .B(n1242), .Z(n1243) );
  NAND U2487 ( .A(n1241), .B(n1243), .Z(n20789) );
  NAND U2488 ( .A(n19143), .B(n19142), .Z(n1244) );
  NAND U2489 ( .A(n18791), .B(n18790), .Z(n1245) );
  AND U2490 ( .A(n1244), .B(n1245), .Z(n18794) );
  NAND U2491 ( .A(n16436), .B(n16435), .Z(n1246) );
  NANDN U2492 ( .A(n16776), .B(n16775), .Z(n1247) );
  AND U2493 ( .A(n1246), .B(n1247), .Z(n16440) );
  NAND U2494 ( .A(n15050), .B(n15049), .Z(n1248) );
  NANDN U2495 ( .A(n15396), .B(n15395), .Z(n1249) );
  AND U2496 ( .A(n1248), .B(n1249), .Z(n15054) );
  XNOR U2497 ( .A(n8676), .B(n8677), .Z(n9011) );
  XNOR U2498 ( .A(n10229), .B(n10228), .Z(n10109) );
  NAND U2499 ( .A(n20952), .B(n20955), .Z(n1250) );
  XOR U2500 ( .A(n20952), .B(n20955), .Z(n1251) );
  NANDN U2501 ( .A(n20953), .B(n1251), .Z(n1252) );
  NAND U2502 ( .A(n1250), .B(n1252), .Z(n20624) );
  NAND U2503 ( .A(n20968), .B(n20971), .Z(n1253) );
  XOR U2504 ( .A(n20968), .B(n20971), .Z(n1254) );
  NANDN U2505 ( .A(n20969), .B(n1254), .Z(n1255) );
  NAND U2506 ( .A(n1253), .B(n1255), .Z(n20640) );
  NAND U2507 ( .A(n20986), .B(n20989), .Z(n1256) );
  XOR U2508 ( .A(n20986), .B(n20989), .Z(n1257) );
  NANDN U2509 ( .A(n20987), .B(n1257), .Z(n1258) );
  NAND U2510 ( .A(n1256), .B(n1258), .Z(n20656) );
  NAND U2511 ( .A(n21003), .B(n21005), .Z(n1259) );
  XOR U2512 ( .A(n21003), .B(n21005), .Z(n1260) );
  NANDN U2513 ( .A(n21002), .B(n1260), .Z(n1261) );
  NAND U2514 ( .A(n1259), .B(n1261), .Z(n20672) );
  XOR U2515 ( .A(n21023), .B(n21021), .Z(n1262) );
  NANDN U2516 ( .A(n21020), .B(n1262), .Z(n1263) );
  NAND U2517 ( .A(n21023), .B(n21021), .Z(n1264) );
  AND U2518 ( .A(n1263), .B(n1264), .Z(n20684) );
  NAND U2519 ( .A(n21036), .B(n21039), .Z(n1265) );
  XOR U2520 ( .A(n21036), .B(n21039), .Z(n1266) );
  NANDN U2521 ( .A(n21037), .B(n1266), .Z(n1267) );
  NAND U2522 ( .A(n1265), .B(n1267), .Z(n20704) );
  NAND U2523 ( .A(n21052), .B(n21055), .Z(n1268) );
  XOR U2524 ( .A(n21052), .B(n21055), .Z(n1269) );
  NANDN U2525 ( .A(n21053), .B(n1269), .Z(n1270) );
  NAND U2526 ( .A(n1268), .B(n1270), .Z(n20720) );
  NAND U2527 ( .A(n21070), .B(n21073), .Z(n1271) );
  XOR U2528 ( .A(n21070), .B(n21073), .Z(n1272) );
  NANDN U2529 ( .A(n21071), .B(n1272), .Z(n1273) );
  NAND U2530 ( .A(n1271), .B(n1273), .Z(n20736) );
  NAND U2531 ( .A(n21084), .B(n21087), .Z(n1274) );
  XOR U2532 ( .A(n21084), .B(n21087), .Z(n1275) );
  NANDN U2533 ( .A(n21085), .B(n1275), .Z(n1276) );
  NAND U2534 ( .A(n1274), .B(n1276), .Z(n20748) );
  XNOR U2535 ( .A(n20792), .B(n20793), .Z(n20795) );
  NAND U2536 ( .A(n20465), .B(n20463), .Z(n1277) );
  XOR U2537 ( .A(n20465), .B(n20463), .Z(n1278) );
  NANDN U2538 ( .A(n20462), .B(n1278), .Z(n1279) );
  NAND U2539 ( .A(n1277), .B(n1279), .Z(n20156) );
  NAND U2540 ( .A(n19497), .B(n19496), .Z(n1280) );
  NAND U2541 ( .A(n19457), .B(n19458), .Z(n1281) );
  AND U2542 ( .A(n1280), .B(n1281), .Z(n19461) );
  NAND U2543 ( .A(n17124), .B(n17123), .Z(n1282) );
  NANDN U2544 ( .A(n17468), .B(n17467), .Z(n1283) );
  AND U2545 ( .A(n1282), .B(n1283), .Z(n17128) );
  NAND U2546 ( .A(n14357), .B(n14356), .Z(n1284) );
  NANDN U2547 ( .A(n14698), .B(n14697), .Z(n1285) );
  AND U2548 ( .A(n1284), .B(n1285), .Z(n14361) );
  NAND U2549 ( .A(n13640), .B(n13639), .Z(n1286) );
  NANDN U2550 ( .A(n13321), .B(n13322), .Z(n1287) );
  AND U2551 ( .A(n1286), .B(n1287), .Z(n13323) );
  NAND U2552 ( .A(n13638), .B(n13637), .Z(n1288) );
  NANDN U2553 ( .A(n14025), .B(n14024), .Z(n1289) );
  AND U2554 ( .A(n1288), .B(n1289), .Z(n13642) );
  XNOR U2555 ( .A(n8672), .B(n8673), .Z(n9021) );
  XNOR U2556 ( .A(n10233), .B(n10232), .Z(n10234) );
  XNOR U2557 ( .A(n21212), .B(n21213), .Z(n21548) );
  NAND U2558 ( .A(n21288), .B(n21291), .Z(n1290) );
  XOR U2559 ( .A(n21288), .B(n21291), .Z(n1291) );
  NANDN U2560 ( .A(n21289), .B(n1291), .Z(n1292) );
  NAND U2561 ( .A(n1290), .B(n1292), .Z(n20957) );
  NAND U2562 ( .A(n21304), .B(n21307), .Z(n1293) );
  XOR U2563 ( .A(n21304), .B(n21307), .Z(n1294) );
  NANDN U2564 ( .A(n21305), .B(n1294), .Z(n1295) );
  NAND U2565 ( .A(n1293), .B(n1295), .Z(n20973) );
  XOR U2566 ( .A(n21323), .B(n21320), .Z(n1296) );
  NANDN U2567 ( .A(n21321), .B(n1296), .Z(n1297) );
  NAND U2568 ( .A(n21323), .B(n21320), .Z(n1298) );
  AND U2569 ( .A(n1297), .B(n1298), .Z(n20991) );
  NAND U2570 ( .A(n21336), .B(n21339), .Z(n1299) );
  XOR U2571 ( .A(n21336), .B(n21339), .Z(n1300) );
  NANDN U2572 ( .A(n21337), .B(n1300), .Z(n1301) );
  NAND U2573 ( .A(n1299), .B(n1301), .Z(n21007) );
  XOR U2574 ( .A(n21355), .B(n21352), .Z(n1302) );
  NANDN U2575 ( .A(n21353), .B(n1302), .Z(n1303) );
  NAND U2576 ( .A(n21355), .B(n21352), .Z(n1304) );
  AND U2577 ( .A(n1303), .B(n1304), .Z(n21025) );
  NAND U2578 ( .A(n21368), .B(n21371), .Z(n1305) );
  XOR U2579 ( .A(n21368), .B(n21371), .Z(n1306) );
  NANDN U2580 ( .A(n21369), .B(n1306), .Z(n1307) );
  NAND U2581 ( .A(n1305), .B(n1307), .Z(n21041) );
  NAND U2582 ( .A(n21384), .B(n21387), .Z(n1308) );
  XOR U2583 ( .A(n21384), .B(n21387), .Z(n1309) );
  NANDN U2584 ( .A(n21385), .B(n1309), .Z(n1310) );
  NAND U2585 ( .A(n1308), .B(n1310), .Z(n21057) );
  NAND U2586 ( .A(n21400), .B(n21403), .Z(n1311) );
  XOR U2587 ( .A(n21400), .B(n21403), .Z(n1312) );
  NANDN U2588 ( .A(n21401), .B(n1312), .Z(n1313) );
  NAND U2589 ( .A(n1311), .B(n1313), .Z(n21069) );
  NAND U2590 ( .A(n21416), .B(n21419), .Z(n1314) );
  XOR U2591 ( .A(n21416), .B(n21419), .Z(n1315) );
  NANDN U2592 ( .A(n21417), .B(n1315), .Z(n1316) );
  NAND U2593 ( .A(n1314), .B(n1316), .Z(n21089) );
  XOR U2594 ( .A(n21435), .B(n21432), .Z(n1317) );
  NANDN U2595 ( .A(n21433), .B(n1317), .Z(n1318) );
  NAND U2596 ( .A(n21435), .B(n21432), .Z(n1319) );
  AND U2597 ( .A(n1318), .B(n1319), .Z(n21157) );
  NAND U2598 ( .A(n15748), .B(n15747), .Z(n1320) );
  NANDN U2599 ( .A(n16096), .B(n16095), .Z(n1321) );
  AND U2600 ( .A(n1320), .B(n1321), .Z(n15752) );
  NAND U2601 ( .A(n13330), .B(n13329), .Z(n1322) );
  NAND U2602 ( .A(n13030), .B(n13031), .Z(n1323) );
  NAND U2603 ( .A(n1322), .B(n1323), .Z(n13663) );
  NAND U2604 ( .A(n9718), .B(n9717), .Z(n1324) );
  NANDN U2605 ( .A(n10084), .B(n10085), .Z(n1325) );
  AND U2606 ( .A(n1324), .B(n1325), .Z(n10093) );
  NAND U2607 ( .A(n22999), .B(n22998), .Z(n1326) );
  NAND U2608 ( .A(n22996), .B(n22997), .Z(n1327) );
  NAND U2609 ( .A(n1326), .B(n1327), .Z(n23127) );
  XNOR U2610 ( .A(n21230), .B(n21231), .Z(n21567) );
  NAND U2611 ( .A(n21620), .B(n21623), .Z(n1328) );
  XOR U2612 ( .A(n21620), .B(n21623), .Z(n1329) );
  NANDN U2613 ( .A(n21621), .B(n1329), .Z(n1330) );
  NAND U2614 ( .A(n1328), .B(n1330), .Z(n21293) );
  NAND U2615 ( .A(n21636), .B(n21639), .Z(n1331) );
  XOR U2616 ( .A(n21636), .B(n21639), .Z(n1332) );
  NANDN U2617 ( .A(n21637), .B(n1332), .Z(n1333) );
  NAND U2618 ( .A(n1331), .B(n1333), .Z(n21309) );
  XOR U2619 ( .A(n21655), .B(n21653), .Z(n1334) );
  NANDN U2620 ( .A(n21652), .B(n1334), .Z(n1335) );
  NAND U2621 ( .A(n21655), .B(n21653), .Z(n1336) );
  AND U2622 ( .A(n1335), .B(n1336), .Z(n21325) );
  NAND U2623 ( .A(n21670), .B(n21673), .Z(n1337) );
  XOR U2624 ( .A(n21670), .B(n21673), .Z(n1338) );
  NANDN U2625 ( .A(n21671), .B(n1338), .Z(n1339) );
  NAND U2626 ( .A(n1337), .B(n1339), .Z(n21341) );
  XOR U2627 ( .A(n21689), .B(n21686), .Z(n1340) );
  NANDN U2628 ( .A(n21687), .B(n1340), .Z(n1341) );
  NAND U2629 ( .A(n21689), .B(n21686), .Z(n1342) );
  AND U2630 ( .A(n1341), .B(n1342), .Z(n21357) );
  NAND U2631 ( .A(n21702), .B(n21705), .Z(n1343) );
  XOR U2632 ( .A(n21702), .B(n21705), .Z(n1344) );
  NANDN U2633 ( .A(n21703), .B(n1344), .Z(n1345) );
  NAND U2634 ( .A(n1343), .B(n1345), .Z(n21373) );
  NAND U2635 ( .A(n21720), .B(n21723), .Z(n1346) );
  XOR U2636 ( .A(n21720), .B(n21723), .Z(n1347) );
  NANDN U2637 ( .A(n21721), .B(n1347), .Z(n1348) );
  NAND U2638 ( .A(n1346), .B(n1348), .Z(n21389) );
  NAND U2639 ( .A(n21736), .B(n21739), .Z(n1349) );
  XOR U2640 ( .A(n21736), .B(n21739), .Z(n1350) );
  NANDN U2641 ( .A(n21737), .B(n1350), .Z(n1351) );
  NAND U2642 ( .A(n1349), .B(n1351), .Z(n21405) );
  NAND U2643 ( .A(n21752), .B(n21755), .Z(n1352) );
  XOR U2644 ( .A(n21752), .B(n21755), .Z(n1353) );
  NANDN U2645 ( .A(n21753), .B(n1353), .Z(n1354) );
  NAND U2646 ( .A(n1352), .B(n1354), .Z(n21421) );
  NAND U2647 ( .A(n21770), .B(n21773), .Z(n1355) );
  XOR U2648 ( .A(n21770), .B(n21773), .Z(n1356) );
  NANDN U2649 ( .A(n21771), .B(n1356), .Z(n1357) );
  NAND U2650 ( .A(n1355), .B(n1357), .Z(n21437) );
  XOR U2651 ( .A(n21796), .B(n21795), .Z(n1358) );
  NANDN U2652 ( .A(n21798), .B(n1358), .Z(n1359) );
  NAND U2653 ( .A(n21796), .B(n21795), .Z(n1360) );
  AND U2654 ( .A(n1359), .B(n1360), .Z(n21805) );
  XNOR U2655 ( .A(n21476), .B(n21477), .Z(n21817) );
  NAND U2656 ( .A(n18800), .B(n18801), .Z(n1361) );
  NAND U2657 ( .A(n18480), .B(n18479), .Z(n1362) );
  NAND U2658 ( .A(n1361), .B(n1362), .Z(n18484) );
  XNOR U2659 ( .A(n9723), .B(n9724), .Z(n9725) );
  XNOR U2660 ( .A(n22563), .B(n22562), .Z(n22564) );
  XOR U2661 ( .A(n21945), .B(n21943), .Z(n1363) );
  NANDN U2662 ( .A(n21942), .B(n1363), .Z(n1364) );
  NAND U2663 ( .A(n21945), .B(n21943), .Z(n1365) );
  AND U2664 ( .A(n1364), .B(n1365), .Z(n21619) );
  NAND U2665 ( .A(n21962), .B(n21965), .Z(n1366) );
  XOR U2666 ( .A(n21962), .B(n21965), .Z(n1367) );
  NANDN U2667 ( .A(n21963), .B(n1367), .Z(n1368) );
  NAND U2668 ( .A(n1366), .B(n1368), .Z(n21635) );
  XOR U2669 ( .A(n21981), .B(n21979), .Z(n1369) );
  NANDN U2670 ( .A(n21978), .B(n1369), .Z(n1370) );
  NAND U2671 ( .A(n21981), .B(n21979), .Z(n1371) );
  AND U2672 ( .A(n1370), .B(n1371), .Z(n21651) );
  NAND U2673 ( .A(n21999), .B(n22001), .Z(n1372) );
  XOR U2674 ( .A(n21999), .B(n22001), .Z(n1373) );
  NANDN U2675 ( .A(n21998), .B(n1373), .Z(n1374) );
  NAND U2676 ( .A(n1372), .B(n1374), .Z(n21669) );
  XOR U2677 ( .A(n22021), .B(n22019), .Z(n1375) );
  NANDN U2678 ( .A(n22018), .B(n1375), .Z(n1376) );
  NAND U2679 ( .A(n22021), .B(n22019), .Z(n1377) );
  AND U2680 ( .A(n1376), .B(n1377), .Z(n21684) );
  XOR U2681 ( .A(n22041), .B(n22038), .Z(n1378) );
  NANDN U2682 ( .A(n22039), .B(n1378), .Z(n1379) );
  NAND U2683 ( .A(n22041), .B(n22038), .Z(n1380) );
  AND U2684 ( .A(n1379), .B(n1380), .Z(n21707) );
  XOR U2685 ( .A(n22057), .B(n22055), .Z(n1381) );
  NANDN U2686 ( .A(n22054), .B(n1381), .Z(n1382) );
  NAND U2687 ( .A(n22057), .B(n22055), .Z(n1383) );
  AND U2688 ( .A(n1382), .B(n1383), .Z(n21719) );
  XOR U2689 ( .A(n22077), .B(n22075), .Z(n1384) );
  NANDN U2690 ( .A(n22074), .B(n1384), .Z(n1385) );
  NAND U2691 ( .A(n22077), .B(n22075), .Z(n1386) );
  AND U2692 ( .A(n1385), .B(n1386), .Z(n21735) );
  XOR U2693 ( .A(n22097), .B(n22095), .Z(n1387) );
  NANDN U2694 ( .A(n22094), .B(n1387), .Z(n1388) );
  NAND U2695 ( .A(n22097), .B(n22095), .Z(n1389) );
  AND U2696 ( .A(n1388), .B(n1389), .Z(n21751) );
  NAND U2697 ( .A(n22115), .B(n22117), .Z(n1390) );
  XOR U2698 ( .A(n22115), .B(n22117), .Z(n1391) );
  NANDN U2699 ( .A(n22114), .B(n1391), .Z(n1392) );
  NAND U2700 ( .A(n1390), .B(n1392), .Z(n21769) );
  NAND U2701 ( .A(n20805), .B(n20804), .Z(n1393) );
  NAND U2702 ( .A(n20470), .B(n20471), .Z(n1394) );
  NAND U2703 ( .A(n1393), .B(n1394), .Z(n20811) );
  NAND U2704 ( .A(n19469), .B(n19470), .Z(n1395) );
  NANDN U2705 ( .A(n19486), .B(n19487), .Z(n1396) );
  NAND U2706 ( .A(n1395), .B(n1396), .Z(n19474) );
  NAND U2707 ( .A(n19472), .B(n19471), .Z(n1397) );
  NAND U2708 ( .A(n19148), .B(n19149), .Z(n1398) );
  NAND U2709 ( .A(n1397), .B(n1398), .Z(n19476) );
  NAND U2710 ( .A(n20473), .B(n20472), .Z(n1399) );
  NAND U2711 ( .A(n20140), .B(n20139), .Z(n1400) );
  AND U2712 ( .A(n1399), .B(n1400), .Z(n20143) );
  NAND U2713 ( .A(n16800), .B(n16799), .Z(n1401) );
  NAND U2714 ( .A(n16452), .B(n16451), .Z(n1402) );
  AND U2715 ( .A(n1401), .B(n1402), .Z(n16456) );
  XNOR U2716 ( .A(n9383), .B(n9384), .Z(n9730) );
  XNOR U2717 ( .A(n22557), .B(n22556), .Z(n22558) );
  NAND U2718 ( .A(n22842), .B(n22841), .Z(n1403) );
  NANDN U2719 ( .A(n22844), .B(n22843), .Z(n1404) );
  NAND U2720 ( .A(n1403), .B(n1404), .Z(n22859) );
  NAND U2721 ( .A(n22865), .B(n22864), .Z(n1405) );
  NAND U2722 ( .A(n22863), .B(n22862), .Z(n1406) );
  NAND U2723 ( .A(n1405), .B(n1406), .Z(n23115) );
  XNOR U2724 ( .A(n21572), .B(n21573), .Z(n21895) );
  XOR U2725 ( .A(n22273), .B(n22274), .Z(n1407) );
  NANDN U2726 ( .A(n22276), .B(n1407), .Z(n1408) );
  NAND U2727 ( .A(n22273), .B(n22274), .Z(n1409) );
  AND U2728 ( .A(n1408), .B(n1409), .Z(n21959) );
  XOR U2729 ( .A(n22293), .B(n22294), .Z(n1410) );
  NANDN U2730 ( .A(n22296), .B(n1410), .Z(n1411) );
  NAND U2731 ( .A(n22293), .B(n22294), .Z(n1412) );
  AND U2732 ( .A(n1411), .B(n1412), .Z(n21975) );
  XOR U2733 ( .A(n22313), .B(n22314), .Z(n1413) );
  NANDN U2734 ( .A(n22316), .B(n1413), .Z(n1414) );
  NAND U2735 ( .A(n22313), .B(n22314), .Z(n1415) );
  AND U2736 ( .A(n1414), .B(n1415), .Z(n21995) );
  XOR U2737 ( .A(n22333), .B(n22334), .Z(n1416) );
  NANDN U2738 ( .A(n22336), .B(n1416), .Z(n1417) );
  NAND U2739 ( .A(n22333), .B(n22334), .Z(n1418) );
  AND U2740 ( .A(n1417), .B(n1418), .Z(n22015) );
  XOR U2741 ( .A(n22356), .B(n22353), .Z(n1419) );
  NAND U2742 ( .A(n1419), .B(n22354), .Z(n1420) );
  NAND U2743 ( .A(n22356), .B(n22353), .Z(n1421) );
  AND U2744 ( .A(n1420), .B(n1421), .Z(n22035) );
  XOR U2745 ( .A(n22373), .B(n22374), .Z(n1422) );
  NANDN U2746 ( .A(n22376), .B(n1422), .Z(n1423) );
  NAND U2747 ( .A(n22373), .B(n22374), .Z(n1424) );
  AND U2748 ( .A(n1423), .B(n1424), .Z(n22051) );
  XOR U2749 ( .A(n22393), .B(n22394), .Z(n1425) );
  NANDN U2750 ( .A(n22396), .B(n1425), .Z(n1426) );
  NAND U2751 ( .A(n22393), .B(n22394), .Z(n1427) );
  AND U2752 ( .A(n1426), .B(n1427), .Z(n22071) );
  XOR U2753 ( .A(n22413), .B(n22414), .Z(n1428) );
  NANDN U2754 ( .A(n22416), .B(n1428), .Z(n1429) );
  NAND U2755 ( .A(n22413), .B(n22414), .Z(n1430) );
  AND U2756 ( .A(n1429), .B(n1430), .Z(n22091) );
  XOR U2757 ( .A(n22433), .B(n22434), .Z(n1431) );
  NANDN U2758 ( .A(n22436), .B(n1431), .Z(n1432) );
  NAND U2759 ( .A(n22433), .B(n22434), .Z(n1433) );
  AND U2760 ( .A(n1432), .B(n1433), .Z(n22111) );
  XOR U2761 ( .A(n22453), .B(n22454), .Z(n1434) );
  NANDN U2762 ( .A(n22456), .B(n1434), .Z(n1435) );
  NAND U2763 ( .A(n22453), .B(n22454), .Z(n1436) );
  AND U2764 ( .A(n1435), .B(n1436), .Z(n22131) );
  NAND U2765 ( .A(n21837), .B(n21839), .Z(n1437) );
  XOR U2766 ( .A(n21837), .B(n21839), .Z(n1438) );
  NANDN U2767 ( .A(n21836), .B(n1438), .Z(n1439) );
  NAND U2768 ( .A(n1437), .B(n1439), .Z(n22140) );
  NAND U2769 ( .A(n18808), .B(n18809), .Z(n1440) );
  NANDN U2770 ( .A(n18816), .B(n18817), .Z(n1441) );
  AND U2771 ( .A(n1440), .B(n1441), .Z(n19157) );
  NAND U2772 ( .A(n17831), .B(n17830), .Z(n1442) );
  NANDN U2773 ( .A(n18157), .B(n18156), .Z(n1443) );
  AND U2774 ( .A(n1442), .B(n1443), .Z(n17835) );
  NAND U2775 ( .A(n14722), .B(n14721), .Z(n1444) );
  NANDN U2776 ( .A(n14373), .B(n14372), .Z(n1445) );
  NAND U2777 ( .A(n1444), .B(n1445), .Z(n14377) );
  XNOR U2778 ( .A(n10262), .B(n10263), .Z(n10978) );
  XNOR U2779 ( .A(n21884), .B(n21885), .Z(n22213) );
  XNOR U2780 ( .A(n21896), .B(n21897), .Z(n22219) );
  XOR U2781 ( .A(n24966), .B(n24965), .Z(n1446) );
  NANDN U2782 ( .A(n24968), .B(n1446), .Z(n1447) );
  NAND U2783 ( .A(n24966), .B(n24965), .Z(n1448) );
  AND U2784 ( .A(n1447), .B(n1448), .Z(n22218) );
  NAND U2785 ( .A(n24818), .B(n24820), .Z(n1449) );
  XOR U2786 ( .A(n24818), .B(n24820), .Z(n1450) );
  NANDN U2787 ( .A(n24817), .B(n1450), .Z(n1451) );
  NAND U2788 ( .A(n1449), .B(n1451), .Z(n22272) );
  XOR U2789 ( .A(n24834), .B(n24831), .Z(n1452) );
  NANDN U2790 ( .A(n24832), .B(n1452), .Z(n1453) );
  NAND U2791 ( .A(n24834), .B(n24831), .Z(n1454) );
  AND U2792 ( .A(n1453), .B(n1454), .Z(n22291) );
  XOR U2793 ( .A(n24846), .B(n24843), .Z(n1455) );
  NANDN U2794 ( .A(n24844), .B(n1455), .Z(n1456) );
  NAND U2795 ( .A(n24846), .B(n24843), .Z(n1457) );
  AND U2796 ( .A(n1456), .B(n1457), .Z(n22311) );
  XOR U2797 ( .A(n24858), .B(n24857), .Z(n1458) );
  NANDN U2798 ( .A(n24860), .B(n1458), .Z(n1459) );
  NAND U2799 ( .A(n24858), .B(n24857), .Z(n1460) );
  AND U2800 ( .A(n1459), .B(n1460), .Z(n22331) );
  NAND U2801 ( .A(n24870), .B(n24872), .Z(n1461) );
  XOR U2802 ( .A(n24870), .B(n24872), .Z(n1462) );
  NANDN U2803 ( .A(n24869), .B(n1462), .Z(n1463) );
  NAND U2804 ( .A(n1461), .B(n1463), .Z(n22352) );
  NAND U2805 ( .A(n24882), .B(n24884), .Z(n1464) );
  XOR U2806 ( .A(n24882), .B(n24884), .Z(n1465) );
  NANDN U2807 ( .A(n24881), .B(n1465), .Z(n1466) );
  NAND U2808 ( .A(n1464), .B(n1466), .Z(n22372) );
  XOR U2809 ( .A(n24896), .B(n24895), .Z(n1467) );
  NANDN U2810 ( .A(n24898), .B(n1467), .Z(n1468) );
  NAND U2811 ( .A(n24896), .B(n24895), .Z(n1469) );
  AND U2812 ( .A(n1468), .B(n1469), .Z(n22391) );
  NAND U2813 ( .A(n24908), .B(n24910), .Z(n1470) );
  XOR U2814 ( .A(n24908), .B(n24910), .Z(n1471) );
  NANDN U2815 ( .A(n24907), .B(n1471), .Z(n1472) );
  NAND U2816 ( .A(n1470), .B(n1472), .Z(n22412) );
  XOR U2817 ( .A(n24922), .B(n24921), .Z(n1473) );
  NANDN U2818 ( .A(n24924), .B(n1473), .Z(n1474) );
  NAND U2819 ( .A(n24922), .B(n24921), .Z(n1475) );
  AND U2820 ( .A(n1474), .B(n1475), .Z(n22431) );
  XOR U2821 ( .A(n24934), .B(n24933), .Z(n1476) );
  NANDN U2822 ( .A(n24936), .B(n1476), .Z(n1477) );
  NAND U2823 ( .A(n24934), .B(n24933), .Z(n1478) );
  AND U2824 ( .A(n1477), .B(n1478), .Z(n22451) );
  NAND U2825 ( .A(n24946), .B(n24948), .Z(n1479) );
  XOR U2826 ( .A(n24946), .B(n24948), .Z(n1480) );
  NANDN U2827 ( .A(n24945), .B(n1480), .Z(n1481) );
  NAND U2828 ( .A(n1479), .B(n1481), .Z(n22474) );
  XOR U2829 ( .A(n22149), .B(n22150), .Z(n1482) );
  XNOR U2830 ( .A(n22148), .B(n1482), .Z(n22486) );
  NAND U2831 ( .A(n14378), .B(n14379), .Z(n1483) );
  NANDN U2832 ( .A(n14047), .B(n14046), .Z(n1484) );
  AND U2833 ( .A(n1483), .B(n1484), .Z(n14381) );
  ANDN U2834 ( .B(n23367), .A(n23368), .Z(n23486) );
  AND U2835 ( .A(n23117), .B(n23118), .Z(n23715) );
  XNOR U2836 ( .A(n22493), .B(n22494), .Z(n24664) );
  NAND U2837 ( .A(n24677), .B(n24680), .Z(n1485) );
  XOR U2838 ( .A(n24677), .B(n24680), .Z(n1486) );
  NANDN U2839 ( .A(n24678), .B(n1486), .Z(n1487) );
  NAND U2840 ( .A(n1485), .B(n1487), .Z(n24686) );
  NAND U2841 ( .A(n20149), .B(n20150), .Z(n24698) );
  ANDN U2842 ( .B(n18491), .A(n18492), .Z(n24715) );
  NAND U2843 ( .A(n24726), .B(n24725), .Z(n1488) );
  NAND U2844 ( .A(n22509), .B(n22508), .Z(n1489) );
  NAND U2845 ( .A(n1488), .B(n1489), .Z(n24727) );
  NAND U2846 ( .A(n24764), .B(n24766), .Z(n1490) );
  XOR U2847 ( .A(n24764), .B(n24766), .Z(n1491) );
  NANDN U2848 ( .A(n24763), .B(n1491), .Z(n1492) );
  NAND U2849 ( .A(n1490), .B(n1492), .Z(n24770) );
  NAND U2850 ( .A(n24788), .B(n24787), .Z(n1493) );
  NAND U2851 ( .A(n22549), .B(n22548), .Z(n1494) );
  NAND U2852 ( .A(n1493), .B(n1494), .Z(n24789) );
  XOR U2853 ( .A(n22847), .B(n22845), .Z(n1495) );
  NANDN U2854 ( .A(n22846), .B(n1495), .Z(n1496) );
  NAND U2855 ( .A(n22847), .B(n22845), .Z(n1497) );
  AND U2856 ( .A(n1496), .B(n1497), .Z(n22850) );
  NAND U2857 ( .A(n23914), .B(n23913), .Z(n1498) );
  NAND U2858 ( .A(n23912), .B(n23911), .Z(n1499) );
  NAND U2859 ( .A(n1498), .B(n1499), .Z(n23917) );
  ANDN U2860 ( .B(n24641), .A(n24642), .Z(n24658) );
  NANDN U2861 ( .A(n5238), .B(n4683), .Z(n1500) );
  XNOR U2862 ( .A(n4681), .B(n1500), .Z(n1501) );
  NANDN U2863 ( .A(n4683), .B(n4682), .Z(n1502) );
  NAND U2864 ( .A(n1501), .B(n1502), .Z(n4955) );
  XNOR U2865 ( .A(n2589), .B(n2590), .Z(n3166) );
  XNOR U2866 ( .A(n3162), .B(n3163), .Z(n3404) );
  XNOR U2867 ( .A(n3399), .B(n3400), .Z(n3654) );
  XNOR U2868 ( .A(n3650), .B(n3651), .Z(n3896) );
  XNOR U2869 ( .A(n3891), .B(n3892), .Z(n4159) );
  XNOR U2870 ( .A(n2479), .B(n2480), .Z(n2593) );
  NANDN U2871 ( .A(n6127), .B(n5532), .Z(n1503) );
  XNOR U2872 ( .A(n5530), .B(n1503), .Z(n1504) );
  NANDN U2873 ( .A(n5532), .B(n5531), .Z(n1505) );
  NAND U2874 ( .A(n1504), .B(n1505), .Z(n5832) );
  XNOR U2875 ( .A(n4421), .B(n4422), .Z(n4424) );
  XNOR U2876 ( .A(n4692), .B(n4693), .Z(n4695) );
  XNOR U2877 ( .A(n4961), .B(n4962), .Z(n4964) );
  XNOR U2878 ( .A(n5250), .B(n5251), .Z(n5549) );
  XOR U2879 ( .A(n2483), .B(n2484), .Z(n2485) );
  XNOR U2880 ( .A(n5543), .B(n5544), .Z(n5846) );
  XNOR U2881 ( .A(n3662), .B(n3663), .Z(n3905) );
  XNOR U2882 ( .A(n3901), .B(n3902), .Z(n4170) );
  XNOR U2883 ( .A(n4166), .B(n4167), .Z(n4433) );
  XOR U2884 ( .A(n3176), .B(n3177), .Z(n3178) );
  XOR U2885 ( .A(n3388), .B(n3389), .Z(n3414) );
  XNOR U2886 ( .A(n4706), .B(n4707), .Z(n4948) );
  XNOR U2887 ( .A(n4975), .B(n4976), .Z(n5235) );
  XNOR U2888 ( .A(n5262), .B(n5263), .Z(n5528) );
  XNOR U2889 ( .A(n5555), .B(n5556), .Z(n5825) );
  XNOR U2890 ( .A(n5840), .B(n5841), .Z(n6146) );
  XNOR U2891 ( .A(n6139), .B(n6140), .Z(n6444) );
  XNOR U2892 ( .A(n3880), .B(n3881), .Z(n3912) );
  XNOR U2893 ( .A(n6153), .B(n6154), .Z(n6463) );
  XNOR U2894 ( .A(n4176), .B(n4177), .Z(n4446) );
  XNOR U2895 ( .A(n4439), .B(n4440), .Z(n4717) );
  XNOR U2896 ( .A(n4710), .B(n4711), .Z(n4986) );
  NANDN U2897 ( .A(n7064), .B(n6429), .Z(n1506) );
  XNOR U2898 ( .A(n6427), .B(n1506), .Z(n1507) );
  NANDN U2899 ( .A(n6429), .B(n6428), .Z(n1508) );
  NAND U2900 ( .A(n1507), .B(n1508), .Z(n6737) );
  XNOR U2901 ( .A(n6446), .B(n6447), .Z(n6753) );
  XNOR U2902 ( .A(n6745), .B(n6746), .Z(n7080) );
  XNOR U2903 ( .A(n3915), .B(n3916), .Z(n4144) );
  XNOR U2904 ( .A(n6425), .B(n6426), .Z(n6457) );
  XNOR U2905 ( .A(n3878), .B(n3879), .Z(n3921) );
  XNOR U2906 ( .A(n6466), .B(n6467), .Z(n6774) );
  XNOR U2907 ( .A(n6163), .B(n6164), .Z(n6471) );
  XNOR U2908 ( .A(n4449), .B(n4450), .Z(n4725) );
  XNOR U2909 ( .A(n5866), .B(n5867), .Z(n6168) );
  XNOR U2910 ( .A(n5569), .B(n5570), .Z(n5871) );
  XNOR U2911 ( .A(n6759), .B(n6760), .Z(n7058) );
  XOR U2912 ( .A(n4993), .B(n4994), .Z(n4996) );
  XOR U2913 ( .A(n5573), .B(n5574), .Z(n5576) );
  XOR U2914 ( .A(n5280), .B(n5281), .Z(n5283) );
  XNOR U2915 ( .A(n7076), .B(n7077), .Z(n7408) );
  XOR U2916 ( .A(n7102), .B(n7103), .Z(n7105) );
  XNOR U2917 ( .A(n7088), .B(n7089), .Z(n7388) );
  XNOR U2918 ( .A(n7092), .B(n7093), .Z(n7385) );
  XOR U2919 ( .A(n4404), .B(n4405), .Z(n4460) );
  XNOR U2920 ( .A(n4730), .B(n4731), .Z(n5004) );
  XNOR U2921 ( .A(n7415), .B(n7416), .Z(n7725) );
  XOR U2922 ( .A(n7114), .B(n7115), .Z(n7116) );
  XNOR U2923 ( .A(n6785), .B(n6786), .Z(n7120) );
  XOR U2924 ( .A(n6482), .B(n6483), .Z(n6484) );
  XNOR U2925 ( .A(n6179), .B(n6180), .Z(n6488) );
  XNOR U2926 ( .A(n5290), .B(n5291), .Z(n5591) );
  XNOR U2927 ( .A(n5882), .B(n5883), .Z(n6183) );
  XNOR U2928 ( .A(n7403), .B(n7404), .Z(n7744) );
  XNOR U2929 ( .A(n7098), .B(n7099), .Z(n7430) );
  XOR U2930 ( .A(n5819), .B(n5820), .Z(n5887) );
  XNOR U2931 ( .A(n5011), .B(n5012), .Z(n5301) );
  NANDN U2932 ( .A(n8061), .B(n7392), .Z(n1509) );
  XNOR U2933 ( .A(n7390), .B(n1509), .Z(n1510) );
  NANDN U2934 ( .A(n7392), .B(n7391), .Z(n1511) );
  NAND U2935 ( .A(n1510), .B(n1511), .Z(n7732) );
  XNOR U2936 ( .A(n7437), .B(n7438), .Z(n7782) );
  XOR U2937 ( .A(n7766), .B(n7767), .Z(n7768) );
  XNOR U2938 ( .A(n5817), .B(n5818), .Z(n6115) );
  XNOR U2939 ( .A(n5298), .B(n5299), .Z(n5605) );
  XNOR U2940 ( .A(n7734), .B(n7735), .Z(n8072) );
  XNOR U2941 ( .A(n7752), .B(n7753), .Z(n8058) );
  XNOR U2942 ( .A(n7762), .B(n7763), .Z(n8100) );
  XNOR U2943 ( .A(n7788), .B(n7789), .Z(n8043) );
  XNOR U2944 ( .A(n7713), .B(n7714), .Z(n7793) );
  XNOR U2945 ( .A(n7451), .B(n7452), .Z(n7799) );
  XNOR U2946 ( .A(n7051), .B(n7052), .Z(n7131) );
  XNOR U2947 ( .A(n6720), .B(n6721), .Z(n6800) );
  XNOR U2948 ( .A(n6498), .B(n6499), .Z(n6805) );
  XNOR U2949 ( .A(n5603), .B(n5604), .Z(n5899) );
  XNOR U2950 ( .A(n8077), .B(n8078), .Z(n8080) );
  XNOR U2951 ( .A(n8067), .B(n8068), .Z(n8401) );
  XNOR U2952 ( .A(n8095), .B(n8096), .Z(n8431) );
  XNOR U2953 ( .A(n7778), .B(n7779), .Z(n8113) );
  XNOR U2954 ( .A(n6197), .B(n6198), .Z(n6418) );
  XNOR U2955 ( .A(n5896), .B(n5897), .Z(n6204) );
  XNOR U2956 ( .A(n7802), .B(n7803), .Z(n8136) );
  XNOR U2957 ( .A(n7461), .B(n7462), .Z(n7807) );
  NAND U2958 ( .A(n3456), .B(n3455), .Z(n1512) );
  NANDN U2959 ( .A(n3619), .B(n3620), .Z(n1513) );
  AND U2960 ( .A(n1512), .B(n1513), .Z(n3616) );
  XNOR U2961 ( .A(n8426), .B(n8427), .Z(n8792) );
  XNOR U2962 ( .A(n8436), .B(n8437), .Z(n8741) );
  XOR U2963 ( .A(n8442), .B(n8443), .Z(n8444) );
  XNOR U2964 ( .A(n8468), .B(n8469), .Z(n8832) );
  XOR U2965 ( .A(n8472), .B(n8473), .Z(n8475) );
  XOR U2966 ( .A(n7465), .B(n7466), .Z(n7468) );
  XOR U2967 ( .A(n7146), .B(n7147), .Z(n7148) );
  XNOR U2968 ( .A(n6514), .B(n6515), .Z(n6823) );
  XNOR U2969 ( .A(n8408), .B(n8409), .Z(n8771) );
  XNOR U2970 ( .A(n8825), .B(n8826), .Z(n8827) );
  XNOR U2971 ( .A(n8478), .B(n8479), .Z(n8732) );
  XNOR U2972 ( .A(n6821), .B(n6822), .Z(n7159) );
  NANDN U2973 ( .A(n9051), .B(n8391), .Z(n1514) );
  XNOR U2974 ( .A(n8389), .B(n1514), .Z(n1515) );
  NANDN U2975 ( .A(n8391), .B(n8390), .Z(n1516) );
  NAND U2976 ( .A(n1515), .B(n1516), .Z(n8755) );
  XNOR U2977 ( .A(n8767), .B(n8768), .Z(n9074) );
  XNOR U2978 ( .A(n8744), .B(n8745), .Z(n8781) );
  XNOR U2979 ( .A(n8746), .B(n8747), .Z(n8777) );
  XOR U2980 ( .A(n8785), .B(n8786), .Z(n8788) );
  XNOR U2981 ( .A(n8797), .B(n8798), .Z(n9044) );
  XNOR U2982 ( .A(n8454), .B(n8455), .Z(n8816) );
  XNOR U2983 ( .A(n8738), .B(n8739), .Z(n8812) );
  XNOR U2984 ( .A(n7475), .B(n7476), .Z(n7823) );
  XNOR U2985 ( .A(n7156), .B(n7157), .Z(n7482) );
  XNOR U2986 ( .A(n8757), .B(n8758), .Z(n9061) );
  XNOR U2987 ( .A(n8845), .B(n8846), .Z(n9158) );
  XOR U2988 ( .A(n8488), .B(n8489), .Z(n8491) );
  NAND U2989 ( .A(n3608), .B(n3607), .Z(n1517) );
  NANDN U2990 ( .A(n3473), .B(n3474), .Z(n1518) );
  AND U2991 ( .A(n1517), .B(n1518), .Z(n3478) );
  XNOR U2992 ( .A(n9435), .B(n9436), .Z(n9787) );
  XNOR U2993 ( .A(n9079), .B(n9080), .Z(n9464) );
  XNOR U2994 ( .A(n9101), .B(n9102), .Z(n9418) );
  XNOR U2995 ( .A(n9125), .B(n9126), .Z(n9504) );
  XNOR U2996 ( .A(n9143), .B(n9144), .Z(n9524) );
  XOR U2997 ( .A(n8373), .B(n8374), .Z(n8495) );
  XNOR U2998 ( .A(n8159), .B(n8160), .Z(n8501) );
  XNOR U2999 ( .A(n7830), .B(n7831), .Z(n8036) );
  XNOR U3000 ( .A(n9067), .B(n9068), .Z(n9070) );
  XNOR U3001 ( .A(n9439), .B(n9440), .Z(n9793) );
  XNOR U3002 ( .A(n10288), .B(n10289), .Z(n10291) );
  XNOR U3003 ( .A(n9461), .B(n9462), .Z(n9817) );
  XNOR U3004 ( .A(n9413), .B(n9414), .Z(n9487) );
  XNOR U3005 ( .A(n9483), .B(n9484), .Z(n9849) );
  XOR U3006 ( .A(n9131), .B(n9132), .Z(n9134) );
  XNOR U3007 ( .A(n9153), .B(n9154), .Z(n9530) );
  XNOR U3008 ( .A(n9445), .B(n9446), .Z(n9799) );
  XNOR U3009 ( .A(n10318), .B(n10319), .Z(n10321) );
  XNOR U3010 ( .A(n9475), .B(n9476), .Z(n9835) );
  XNOR U3011 ( .A(n9491), .B(n9492), .Z(n9494) );
  XNOR U3012 ( .A(n9497), .B(n9498), .Z(n9771) );
  XNOR U3013 ( .A(n9893), .B(n9892), .Z(n1519) );
  XNOR U3014 ( .A(n9894), .B(n1519), .Z(n9895) );
  XOR U3015 ( .A(n9535), .B(n9536), .Z(n9913) );
  XOR U3016 ( .A(n9035), .B(n9036), .Z(n9170) );
  XNOR U3017 ( .A(n10282), .B(n10283), .Z(n10738) );
  XNOR U3018 ( .A(n9471), .B(n9472), .Z(n9829) );
  XNOR U3019 ( .A(n9852), .B(n9853), .Z(n10361) );
  XNOR U3020 ( .A(n9509), .B(n9510), .Z(n9874) );
  XNOR U3021 ( .A(n9906), .B(n9905), .Z(n1520) );
  XNOR U3022 ( .A(n9907), .B(n1520), .Z(n9908) );
  XOR U3023 ( .A(n9033), .B(n9034), .Z(n9174) );
  XNOR U3024 ( .A(n8720), .B(n8721), .Z(n8859) );
  XNOR U3025 ( .A(n10733), .B(n10734), .Z(n11008) );
  XNOR U3026 ( .A(n10747), .B(n10748), .Z(n10993) );
  XNOR U3027 ( .A(n9824), .B(n9825), .Z(n10333) );
  XNOR U3028 ( .A(n9842), .B(n9843), .Z(n10348) );
  XNOR U3029 ( .A(n9882), .B(n9883), .Z(n10390) );
  XOR U3030 ( .A(n2852), .B(n2851), .Z(n2844) );
  XNOR U3031 ( .A(n11010), .B(n11011), .Z(n11426) );
  XOR U3032 ( .A(n11022), .B(n11023), .Z(n11458) );
  XNOR U3033 ( .A(n9806), .B(n9807), .Z(n10312) );
  XNOR U3034 ( .A(n10753), .B(n10754), .Z(n10755) );
  XNOR U3035 ( .A(n10330), .B(n10331), .Z(n10771) );
  XNOR U3036 ( .A(n10350), .B(n10351), .Z(n10715) );
  XNOR U3037 ( .A(n10378), .B(n10379), .Z(n10381) );
  XOR U3038 ( .A(n10374), .B(n10375), .Z(n10714) );
  XNOR U3039 ( .A(n10392), .B(n10393), .Z(n10808) );
  NAND U3040 ( .A(n11109), .B(n11112), .Z(n1521) );
  XOR U3041 ( .A(n11109), .B(n11112), .Z(n1522) );
  NANDN U3042 ( .A(n11110), .B(n1522), .Z(n1523) );
  NAND U3043 ( .A(n1521), .B(n1523), .Z(n10806) );
  NAND U3044 ( .A(n10423), .B(n10424), .Z(n1524) );
  XOR U3045 ( .A(n10423), .B(n10424), .Z(n1525) );
  NANDN U3046 ( .A(n10422), .B(n1525), .Z(n1526) );
  NAND U3047 ( .A(n1524), .B(n1526), .Z(n9920) );
  XNOR U3048 ( .A(n11441), .B(n11442), .Z(n11729) );
  XNOR U3049 ( .A(n11724), .B(n11725), .Z(n12127) );
  XNOR U3050 ( .A(n10314), .B(n10315), .Z(n10719) );
  NAND U3051 ( .A(n11053), .B(n11056), .Z(n1527) );
  XOR U3052 ( .A(n11053), .B(n11056), .Z(n1528) );
  NANDN U3053 ( .A(n11054), .B(n1528), .Z(n1529) );
  NAND U3054 ( .A(n1527), .B(n1529), .Z(n10768) );
  XNOR U3055 ( .A(n10368), .B(n10369), .Z(n10794) );
  NAND U3056 ( .A(n11518), .B(n11521), .Z(n1530) );
  XOR U3057 ( .A(n11518), .B(n11521), .Z(n1531) );
  NANDN U3058 ( .A(n11519), .B(n1531), .Z(n1532) );
  NAND U3059 ( .A(n1530), .B(n1532), .Z(n11108) );
  XOR U3060 ( .A(n9926), .B(n9927), .Z(n10434) );
  XOR U3061 ( .A(n2896), .B(n2895), .Z(n2901) );
  XNOR U3062 ( .A(n12142), .B(n12143), .Z(n12452) );
  XNOR U3063 ( .A(n12447), .B(n12448), .Z(n12825) );
  XNOR U3064 ( .A(n11471), .B(n11472), .Z(n11474) );
  XNOR U3065 ( .A(n11035), .B(n11036), .Z(n11480) );
  XOR U3066 ( .A(n10774), .B(n10775), .Z(n11071) );
  XNOR U3067 ( .A(n11084), .B(n11085), .Z(n11419) );
  XNOR U3068 ( .A(n11500), .B(n11501), .Z(n11800) );
  XNOR U3069 ( .A(n10796), .B(n10797), .Z(n10990) );
  XNOR U3070 ( .A(n11094), .B(n11095), .Z(n11418) );
  XNOR U3071 ( .A(n11126), .B(n11127), .Z(n1533) );
  XNOR U3072 ( .A(n11125), .B(n1533), .Z(n11410) );
  XOR U3073 ( .A(n11138), .B(n11137), .Z(n1534) );
  XNOR U3074 ( .A(n11136), .B(n1534), .Z(n11408) );
  XOR U3075 ( .A(n10830), .B(n10831), .Z(n10832) );
  NAND U3076 ( .A(n4648), .B(n4647), .Z(n1535) );
  NANDN U3077 ( .A(n4536), .B(n4535), .Z(n1536) );
  AND U3078 ( .A(n1535), .B(n1536), .Z(n4646) );
  XNOR U3079 ( .A(n2918), .B(n2917), .Z(n2909) );
  XNOR U3080 ( .A(n11453), .B(n11454), .Z(n11740) );
  XNOR U3081 ( .A(n12840), .B(n12841), .Z(n13079) );
  XNOR U3082 ( .A(n11736), .B(n11737), .Z(n12159) );
  XNOR U3083 ( .A(n11754), .B(n11755), .Z(n12176) );
  XNOR U3084 ( .A(n11773), .B(n11774), .Z(n11775) );
  XOR U3085 ( .A(n11780), .B(n11781), .Z(n1537) );
  XNOR U3086 ( .A(n11779), .B(n1537), .Z(n12201) );
  XNOR U3087 ( .A(n11067), .B(n11068), .Z(n11422) );
  XNOR U3088 ( .A(n11492), .B(n11493), .Z(n11787) );
  XNOR U3089 ( .A(n11504), .B(n11505), .Z(n11707) );
  NAND U3090 ( .A(n11820), .B(n11823), .Z(n1538) );
  XOR U3091 ( .A(n11820), .B(n11823), .Z(n1539) );
  NANDN U3092 ( .A(n11821), .B(n1539), .Z(n1540) );
  NAND U3093 ( .A(n1538), .B(n1540), .Z(n11522) );
  XOR U3094 ( .A(n2934), .B(n2933), .Z(n2937) );
  XNOR U3095 ( .A(n13074), .B(n13075), .Z(n13374) );
  XNOR U3096 ( .A(n12154), .B(n12155), .Z(n12464) );
  XNOR U3097 ( .A(n12459), .B(n12460), .Z(n12857) );
  NAND U3098 ( .A(n12522), .B(n12525), .Z(n1541) );
  XOR U3099 ( .A(n12522), .B(n12525), .Z(n1542) );
  NANDN U3100 ( .A(n12523), .B(n1542), .Z(n1543) );
  NAND U3101 ( .A(n1541), .B(n1543), .Z(n12223) );
  XOR U3102 ( .A(n12231), .B(n12232), .Z(n1544) );
  NANDN U3103 ( .A(n12233), .B(n1544), .Z(n1545) );
  NAND U3104 ( .A(n12231), .B(n12232), .Z(n1546) );
  AND U3105 ( .A(n1545), .B(n1546), .Z(n11825) );
  XOR U3106 ( .A(n12255), .B(n12256), .Z(n1547) );
  XNOR U3107 ( .A(n12254), .B(n1547), .Z(n12420) );
  XNOR U3108 ( .A(n12561), .B(n12562), .Z(n12808) );
  XNOR U3109 ( .A(n11550), .B(n11551), .Z(n11700) );
  XOR U3110 ( .A(n2962), .B(n2961), .Z(n2967) );
  XNOR U3111 ( .A(n13389), .B(n13390), .Z(n13748) );
  XNOR U3112 ( .A(n12852), .B(n12853), .Z(n13091) );
  XNOR U3113 ( .A(n11771), .B(n11772), .Z(n1548) );
  XNOR U3114 ( .A(n11770), .B(n1548), .Z(n12125) );
  XNOR U3115 ( .A(n12206), .B(n12207), .Z(n12513) );
  XNOR U3116 ( .A(n11792), .B(n11793), .Z(n12121) );
  XOR U3117 ( .A(n12916), .B(n12917), .Z(n1549) );
  NANDN U3118 ( .A(n12918), .B(n1549), .Z(n1550) );
  NAND U3119 ( .A(n12916), .B(n12917), .Z(n1551) );
  AND U3120 ( .A(n1550), .B(n1551), .Z(n12527) );
  XNOR U3121 ( .A(n12268), .B(n12269), .Z(n12270) );
  XOR U3122 ( .A(n11556), .B(n11557), .Z(n11871) );
  XNOR U3123 ( .A(n2954), .B(n2953), .Z(n2955) );
  XNOR U3124 ( .A(n2986), .B(n2985), .Z(n2987) );
  XNOR U3125 ( .A(n13737), .B(n13738), .Z(n14111) );
  XNOR U3126 ( .A(n13086), .B(n13087), .Z(n13406) );
  XNOR U3127 ( .A(n13401), .B(n13402), .Z(n13760) );
  XNOR U3128 ( .A(n12469), .B(n12470), .Z(n12869) );
  XNOR U3129 ( .A(n12184), .B(n12185), .Z(n12491) );
  XNOR U3130 ( .A(n12188), .B(n12189), .Z(n12428) );
  XOR U3131 ( .A(n12930), .B(n12932), .Z(n1552) );
  NANDN U3132 ( .A(n12931), .B(n1552), .Z(n1553) );
  NAND U3133 ( .A(n12930), .B(n12932), .Z(n1554) );
  AND U3134 ( .A(n1553), .B(n1554), .Z(n12540) );
  XOR U3135 ( .A(n12261), .B(n12262), .Z(n1555) );
  XNOR U3136 ( .A(n12263), .B(n1555), .Z(n12417) );
  XNOR U3137 ( .A(n13188), .B(n13189), .Z(n13359) );
  NAND U3138 ( .A(n11563), .B(n11565), .Z(n1556) );
  XOR U3139 ( .A(n11563), .B(n11565), .Z(n1557) );
  NANDN U3140 ( .A(n11562), .B(n1557), .Z(n1558) );
  NAND U3141 ( .A(n1556), .B(n1558), .Z(n11164) );
  XNOR U3142 ( .A(n3306), .B(n3307), .Z(n3549) );
  XNOR U3143 ( .A(n2929), .B(n2930), .Z(n3313) );
  XNOR U3144 ( .A(n3004), .B(n3003), .Z(n3005) );
  XNOR U3145 ( .A(n14420), .B(n14421), .Z(n14422) );
  XNOR U3146 ( .A(n14104), .B(n14105), .Z(n14427) );
  XOR U3147 ( .A(n12429), .B(n12430), .Z(n12476) );
  XNOR U3148 ( .A(n13096), .B(n13097), .Z(n13418) );
  XNOR U3149 ( .A(n12493), .B(n12494), .Z(n12822) );
  XNOR U3150 ( .A(n12888), .B(n12889), .Z(n13052) );
  XOR U3151 ( .A(n12901), .B(n12902), .Z(n1559) );
  XNOR U3152 ( .A(n12900), .B(n1559), .Z(n13049) );
  XOR U3153 ( .A(n12421), .B(n12422), .Z(n12940) );
  XOR U3154 ( .A(n12947), .B(n12948), .Z(n1560) );
  XNOR U3155 ( .A(n12946), .B(n1560), .Z(n13041) );
  XNOR U3156 ( .A(n13192), .B(n13193), .Z(n13194) );
  NAND U3157 ( .A(n12968), .B(n12971), .Z(n1561) );
  XOR U3158 ( .A(n12968), .B(n12971), .Z(n1562) );
  NANDN U3159 ( .A(n12969), .B(n1562), .Z(n1563) );
  NAND U3160 ( .A(n1561), .B(n1563), .Z(n12581) );
  NAND U3161 ( .A(n12582), .B(n12585), .Z(n1564) );
  XOR U3162 ( .A(n12582), .B(n12585), .Z(n1565) );
  NANDN U3163 ( .A(n12583), .B(n1565), .Z(n1566) );
  NAND U3164 ( .A(n1564), .B(n1566), .Z(n12280) );
  XOR U3165 ( .A(n12290), .B(n12287), .Z(n1567) );
  NAND U3166 ( .A(n1567), .B(n12288), .Z(n1568) );
  NAND U3167 ( .A(n12290), .B(n12287), .Z(n1569) );
  AND U3168 ( .A(n1568), .B(n1569), .Z(n11879) );
  XNOR U3169 ( .A(n3010), .B(n3009), .Z(n3012) );
  XNOR U3170 ( .A(n3026), .B(n3025), .Z(n3027) );
  XNOR U3171 ( .A(n13755), .B(n13756), .Z(n14125) );
  XNOR U3172 ( .A(n14120), .B(n14121), .Z(n14445) );
  XOR U3173 ( .A(n13725), .B(n13726), .Z(n13772) );
  XOR U3174 ( .A(n13056), .B(n13057), .Z(n13103) );
  XNOR U3175 ( .A(n13148), .B(n13149), .Z(n13150) );
  NAND U3176 ( .A(n13490), .B(n13493), .Z(n1570) );
  XOR U3177 ( .A(n13490), .B(n13493), .Z(n1571) );
  NANDN U3178 ( .A(n13491), .B(n1571), .Z(n1572) );
  NAND U3179 ( .A(n1570), .B(n1572), .Z(n13164) );
  XOR U3180 ( .A(n13172), .B(n13173), .Z(n1573) );
  XNOR U3181 ( .A(n13171), .B(n1573), .Z(n13506) );
  XNOR U3182 ( .A(n12937), .B(n12938), .Z(n13043) );
  NAND U3183 ( .A(n13205), .B(n13208), .Z(n1574) );
  XOR U3184 ( .A(n13205), .B(n13208), .Z(n1575) );
  NANDN U3185 ( .A(n13206), .B(n1575), .Z(n1576) );
  NAND U3186 ( .A(n1574), .B(n1576), .Z(n12966) );
  NAND U3187 ( .A(n13533), .B(n13536), .Z(n1577) );
  XOR U3188 ( .A(n13533), .B(n13536), .Z(n1578) );
  NANDN U3189 ( .A(n13534), .B(n1578), .Z(n1579) );
  NAND U3190 ( .A(n1577), .B(n1579), .Z(n13204) );
  NAND U3191 ( .A(n5200), .B(n5199), .Z(n1580) );
  NAND U3192 ( .A(n5109), .B(n5110), .Z(n1581) );
  AND U3193 ( .A(n1580), .B(n1581), .Z(n5112) );
  XNOR U3194 ( .A(n3798), .B(n3799), .Z(n4057) );
  XNOR U3195 ( .A(n3553), .B(n3554), .Z(n3804) );
  XNOR U3196 ( .A(n3320), .B(n3321), .Z(n3562) );
  XNOR U3197 ( .A(n2991), .B(n2992), .Z(n3327) );
  XNOR U3198 ( .A(n3042), .B(n3041), .Z(n3043) );
  XNOR U3199 ( .A(n14438), .B(n14439), .Z(n14440) );
  XNOR U3200 ( .A(n13765), .B(n13766), .Z(n14137) );
  XNOR U3201 ( .A(n12874), .B(n12875), .Z(n13055) );
  XOR U3202 ( .A(n13128), .B(n13127), .Z(n1582) );
  XNOR U3203 ( .A(n13126), .B(n1582), .Z(n13370) );
  NAND U3204 ( .A(n13805), .B(n13808), .Z(n1583) );
  XOR U3205 ( .A(n13805), .B(n13808), .Z(n1584) );
  NANDN U3206 ( .A(n13806), .B(n1584), .Z(n1585) );
  NAND U3207 ( .A(n1583), .B(n1585), .Z(n13456) );
  NAND U3208 ( .A(n13819), .B(n13822), .Z(n1586) );
  XOR U3209 ( .A(n13819), .B(n13822), .Z(n1587) );
  NANDN U3210 ( .A(n13820), .B(n1587), .Z(n1588) );
  NAND U3211 ( .A(n1586), .B(n1588), .Z(n13472) );
  XOR U3212 ( .A(n13143), .B(n13142), .Z(n1589) );
  XNOR U3213 ( .A(n13141), .B(n1589), .Z(n13366) );
  XNOR U3214 ( .A(n13494), .B(n13495), .Z(n13713) );
  XNOR U3215 ( .A(n13516), .B(n13517), .Z(n13872) );
  XNOR U3216 ( .A(n4055), .B(n4056), .Z(n4320) );
  XNOR U3217 ( .A(n3054), .B(n3053), .Z(n3056) );
  XOR U3218 ( .A(n3064), .B(n3063), .Z(n3067) );
  XOR U3219 ( .A(n14410), .B(n14411), .Z(n14457) );
  XNOR U3220 ( .A(n13431), .B(n13432), .Z(n13787) );
  XNOR U3221 ( .A(n13783), .B(n13784), .Z(n14157) );
  NAND U3222 ( .A(n14210), .B(n14213), .Z(n1590) );
  XOR U3223 ( .A(n14210), .B(n14213), .Z(n1591) );
  NANDN U3224 ( .A(n14211), .B(n1591), .Z(n1592) );
  NAND U3225 ( .A(n1590), .B(n1592), .Z(n13842) );
  XOR U3226 ( .A(n13887), .B(n13888), .Z(n1593) );
  XNOR U3227 ( .A(n13886), .B(n1593), .Z(n14075) );
  XNOR U3228 ( .A(n14251), .B(n14252), .Z(n14389) );
  XOR U3229 ( .A(n13219), .B(n13220), .Z(n13221) );
  NAND U3230 ( .A(n11581), .B(n11583), .Z(n1594) );
  XOR U3231 ( .A(n11581), .B(n11583), .Z(n1595) );
  NANDN U3232 ( .A(n11580), .B(n1595), .Z(n1596) );
  NAND U3233 ( .A(n1594), .B(n1596), .Z(n11186) );
  XNOR U3234 ( .A(n4318), .B(n4319), .Z(n4587) );
  XNOR U3235 ( .A(n3812), .B(n3813), .Z(n4070) );
  XNOR U3236 ( .A(n3565), .B(n3566), .Z(n3818) );
  XNOR U3237 ( .A(n3332), .B(n3333), .Z(n3574) );
  XNOR U3238 ( .A(n3017), .B(n3018), .Z(n3337) );
  XNOR U3239 ( .A(n3092), .B(n3091), .Z(n3093) );
  XNOR U3240 ( .A(n13803), .B(n13804), .Z(n14091) );
  NAND U3241 ( .A(n14519), .B(n14522), .Z(n1597) );
  XOR U3242 ( .A(n14519), .B(n14522), .Z(n1598) );
  NANDN U3243 ( .A(n14520), .B(n1598), .Z(n1599) );
  NAND U3244 ( .A(n1597), .B(n1599), .Z(n14206) );
  NAND U3245 ( .A(n14895), .B(n14898), .Z(n1600) );
  XOR U3246 ( .A(n14895), .B(n14898), .Z(n1601) );
  NANDN U3247 ( .A(n14896), .B(n1601), .Z(n1602) );
  NAND U3248 ( .A(n1600), .B(n1602), .Z(n14524) );
  XNOR U3249 ( .A(n14222), .B(n14223), .Z(n14396) );
  XNOR U3250 ( .A(n13709), .B(n13710), .Z(n14233) );
  XNOR U3251 ( .A(n14241), .B(n14242), .Z(n14391) );
  XOR U3252 ( .A(n13903), .B(n13905), .Z(n1603) );
  NANDN U3253 ( .A(n13904), .B(n1603), .Z(n1604) );
  NAND U3254 ( .A(n13903), .B(n13905), .Z(n1605) );
  AND U3255 ( .A(n1604), .B(n1605), .Z(n13550) );
  NAND U3256 ( .A(n12981), .B(n12980), .Z(n1606) );
  NANDN U3257 ( .A(n13034), .B(n13035), .Z(n1607) );
  NAND U3258 ( .A(n1606), .B(n1607), .Z(n13226) );
  XNOR U3259 ( .A(n4585), .B(n4586), .Z(n4862) );
  XNOR U3260 ( .A(n4067), .B(n4068), .Z(n4331) );
  XNOR U3261 ( .A(n3086), .B(n3085), .Z(n3087) );
  XNOR U3262 ( .A(n3112), .B(n3111), .Z(n3113) );
  XOR U3263 ( .A(n15103), .B(n15104), .Z(n15150) );
  XNOR U3264 ( .A(n14830), .B(n14831), .Z(n15160) );
  XNOR U3265 ( .A(n14150), .B(n14151), .Z(n14473) );
  XNOR U3266 ( .A(n14468), .B(n14469), .Z(n14845) );
  XOR U3267 ( .A(n14229), .B(n14230), .Z(n1608) );
  XNOR U3268 ( .A(n14228), .B(n1608), .Z(n14394) );
  XNOR U3269 ( .A(n14558), .B(n14559), .Z(n1609) );
  XNOR U3270 ( .A(n14557), .B(n1609), .Z(n14761) );
  XOR U3271 ( .A(n14580), .B(n14581), .Z(n1610) );
  XNOR U3272 ( .A(n14579), .B(n1610), .Z(n14757) );
  XNOR U3273 ( .A(n4860), .B(n4861), .Z(n5141) );
  XNOR U3274 ( .A(n3079), .B(n3080), .Z(n3348) );
  XNOR U3275 ( .A(n4332), .B(n4333), .Z(n4600) );
  XNOR U3276 ( .A(n3822), .B(n3823), .Z(n4081) );
  XNOR U3277 ( .A(n3577), .B(n3578), .Z(n3829) );
  XNOR U3278 ( .A(n3342), .B(n3343), .Z(n3585) );
  XNOR U3279 ( .A(n10137), .B(n10136), .Z(n10138) );
  XNOR U3280 ( .A(n14842), .B(n14843), .Z(n15172) );
  XNOR U3281 ( .A(n14168), .B(n14169), .Z(n1611) );
  XNOR U3282 ( .A(n14167), .B(n1611), .Z(n14493) );
  XOR U3283 ( .A(n14174), .B(n14175), .Z(n1612) );
  XNOR U3284 ( .A(n14173), .B(n1612), .Z(n14176) );
  XNOR U3285 ( .A(n14535), .B(n14536), .Z(n1613) );
  XNOR U3286 ( .A(n14534), .B(n1613), .Z(n14767) );
  NAND U3287 ( .A(n15232), .B(n15235), .Z(n1614) );
  XOR U3288 ( .A(n15232), .B(n15235), .Z(n1615) );
  NANDN U3289 ( .A(n15233), .B(n1615), .Z(n1616) );
  NAND U3290 ( .A(n1614), .B(n1616), .Z(n14913) );
  XNOR U3291 ( .A(n5139), .B(n5140), .Z(n5428) );
  NAND U3292 ( .A(n6301), .B(n6302), .Z(n1617) );
  NANDN U3293 ( .A(n6382), .B(n6381), .Z(n1618) );
  NAND U3294 ( .A(n1617), .B(n1618), .Z(n6303) );
  XNOR U3295 ( .A(n4597), .B(n4598), .Z(n4873) );
  XNOR U3296 ( .A(n4079), .B(n4080), .Z(n4344) );
  XNOR U3297 ( .A(n10143), .B(n10142), .Z(n10144) );
  XNOR U3298 ( .A(n22683), .B(n22682), .Z(n22685) );
  XNOR U3299 ( .A(n15153), .B(n15154), .Z(n15527) );
  XNOR U3300 ( .A(n14484), .B(n14485), .Z(n14861) );
  XNOR U3301 ( .A(n14854), .B(n14855), .Z(n15184) );
  XOR U3302 ( .A(n14773), .B(n14772), .Z(n1619) );
  NANDN U3303 ( .A(n14775), .B(n1619), .Z(n1620) );
  NAND U3304 ( .A(n14773), .B(n14772), .Z(n1621) );
  AND U3305 ( .A(n1620), .B(n1621), .Z(n14881) );
  NAND U3306 ( .A(n15595), .B(n15598), .Z(n1622) );
  XOR U3307 ( .A(n15595), .B(n15598), .Z(n1623) );
  NANDN U3308 ( .A(n15596), .B(n1623), .Z(n1624) );
  NAND U3309 ( .A(n1622), .B(n1624), .Z(n15237) );
  NAND U3310 ( .A(n15624), .B(n15627), .Z(n1625) );
  XOR U3311 ( .A(n15624), .B(n15627), .Z(n1626) );
  NANDN U3312 ( .A(n15625), .B(n1626), .Z(n1627) );
  NAND U3313 ( .A(n1625), .B(n1627), .Z(n15261) );
  XOR U3314 ( .A(n14934), .B(n14935), .Z(n1628) );
  XNOR U3315 ( .A(n14933), .B(n1628), .Z(n15086) );
  NAND U3316 ( .A(n15968), .B(n15971), .Z(n1629) );
  XOR U3317 ( .A(n15968), .B(n15971), .Z(n1630) );
  NANDN U3318 ( .A(n15969), .B(n1630), .Z(n1631) );
  NAND U3319 ( .A(n1629), .B(n1631), .Z(n15638) );
  XNOR U3320 ( .A(n15646), .B(n15647), .Z(n15648) );
  XOR U3321 ( .A(n14966), .B(n14965), .Z(n1632) );
  XNOR U3322 ( .A(n14964), .B(n1632), .Z(n15079) );
  XOR U3323 ( .A(n14588), .B(n14587), .Z(n1633) );
  XNOR U3324 ( .A(n14586), .B(n1633), .Z(n14755) );
  XNOR U3325 ( .A(n15296), .B(n15297), .Z(n15298) );
  NAND U3326 ( .A(n14285), .B(n14287), .Z(n1634) );
  XOR U3327 ( .A(n14285), .B(n14287), .Z(n1635) );
  NANDN U3328 ( .A(n14284), .B(n1635), .Z(n1636) );
  NAND U3329 ( .A(n1634), .B(n1636), .Z(n13917) );
  NAND U3330 ( .A(n13568), .B(n13567), .Z(n1637) );
  NANDN U3331 ( .A(n13232), .B(n13231), .Z(n1638) );
  AND U3332 ( .A(n1637), .B(n1638), .Z(n13233) );
  NAND U3333 ( .A(n12799), .B(n12798), .Z(n1639) );
  NANDN U3334 ( .A(n13235), .B(n13236), .Z(n1640) );
  NAND U3335 ( .A(n1639), .B(n1640), .Z(n12995) );
  XNOR U3336 ( .A(n5426), .B(n5427), .Z(n5721) );
  XNOR U3337 ( .A(n3589), .B(n3590), .Z(n3840) );
  XNOR U3338 ( .A(n4874), .B(n4875), .Z(n5154) );
  XNOR U3339 ( .A(n4342), .B(n4343), .Z(n4611) );
  XNOR U3340 ( .A(n3834), .B(n3835), .Z(n4093) );
  XNOR U3341 ( .A(n3356), .B(n3357), .Z(n3598) );
  XNOR U3342 ( .A(n10149), .B(n10148), .Z(n10151) );
  XNOR U3343 ( .A(n15165), .B(n15166), .Z(n15539) );
  XOR U3344 ( .A(n14873), .B(n14874), .Z(n1641) );
  XNOR U3345 ( .A(n14872), .B(n1641), .Z(n15100) );
  NAND U3346 ( .A(n15952), .B(n15955), .Z(n1642) );
  XOR U3347 ( .A(n15952), .B(n15955), .Z(n1643) );
  NANDN U3348 ( .A(n15953), .B(n1643), .Z(n1644) );
  NAND U3349 ( .A(n1642), .B(n1644), .Z(n15622) );
  NAND U3350 ( .A(n16330), .B(n16333), .Z(n1645) );
  XOR U3351 ( .A(n16330), .B(n16333), .Z(n1646) );
  NANDN U3352 ( .A(n16331), .B(n1646), .Z(n1647) );
  NAND U3353 ( .A(n1645), .B(n1647), .Z(n15973) );
  NAND U3354 ( .A(n15985), .B(n15988), .Z(n1648) );
  XOR U3355 ( .A(n15985), .B(n15988), .Z(n1649) );
  NANDN U3356 ( .A(n15986), .B(n1649), .Z(n1650) );
  NAND U3357 ( .A(n1648), .B(n1650), .Z(n15657) );
  XNOR U3358 ( .A(n15665), .B(n15666), .Z(n15667) );
  NAND U3359 ( .A(n14984), .B(n14986), .Z(n1651) );
  XOR U3360 ( .A(n14984), .B(n14986), .Z(n1652) );
  NANDN U3361 ( .A(n14983), .B(n1652), .Z(n1653) );
  NAND U3362 ( .A(n1651), .B(n1653), .Z(n14602) );
  XNOR U3363 ( .A(n5719), .B(n5720), .Z(n6020) );
  XNOR U3364 ( .A(n5151), .B(n5152), .Z(n5439) );
  XNOR U3365 ( .A(n4609), .B(n4610), .Z(n4886) );
  XNOR U3366 ( .A(n4091), .B(n4092), .Z(n4356) );
  XNOR U3367 ( .A(n15177), .B(n15178), .Z(n15551) );
  XOR U3368 ( .A(n15587), .B(n15588), .Z(n1654) );
  XNOR U3369 ( .A(n15586), .B(n1654), .Z(n15924) );
  XNOR U3370 ( .A(n15611), .B(n15612), .Z(n15613) );
  NAND U3371 ( .A(n16676), .B(n16679), .Z(n1655) );
  XOR U3372 ( .A(n16676), .B(n16679), .Z(n1656) );
  NANDN U3373 ( .A(n16677), .B(n1656), .Z(n1657) );
  NAND U3374 ( .A(n1655), .B(n1657), .Z(n16349) );
  XNOR U3375 ( .A(n15989), .B(n15990), .Z(n16353) );
  XNOR U3376 ( .A(n15309), .B(n15310), .Z(n15675) );
  XNOR U3377 ( .A(n6018), .B(n6019), .Z(n6072) );
  XNOR U3378 ( .A(n5440), .B(n5441), .Z(n5734) );
  XNOR U3379 ( .A(n4884), .B(n4885), .Z(n5165) );
  XNOR U3380 ( .A(n4354), .B(n4355), .Z(n4623) );
  XNOR U3381 ( .A(n3848), .B(n3849), .Z(n4106) );
  XNOR U3382 ( .A(n10161), .B(n10160), .Z(n10163) );
  NAND U3383 ( .A(n15891), .B(n15894), .Z(n1658) );
  XOR U3384 ( .A(n15891), .B(n15894), .Z(n1659) );
  NANDN U3385 ( .A(n15892), .B(n1659), .Z(n1660) );
  NAND U3386 ( .A(n1658), .B(n1660), .Z(n15566) );
  XNOR U3387 ( .A(n15195), .B(n15196), .Z(n1661) );
  XNOR U3388 ( .A(n15197), .B(n1661), .Z(n15467) );
  NAND U3389 ( .A(n15905), .B(n15908), .Z(n1662) );
  XOR U3390 ( .A(n15905), .B(n15908), .Z(n1663) );
  NANDN U3391 ( .A(n15906), .B(n1663), .Z(n1664) );
  NAND U3392 ( .A(n1662), .B(n1664), .Z(n15787) );
  XOR U3393 ( .A(n16309), .B(n16311), .Z(n1665) );
  NANDN U3394 ( .A(n16310), .B(n1665), .Z(n1666) );
  NAND U3395 ( .A(n16309), .B(n16311), .Z(n1667) );
  AND U3396 ( .A(n1666), .B(n1667), .Z(n15946) );
  XNOR U3397 ( .A(n16318), .B(n16319), .Z(n16477) );
  NAND U3398 ( .A(n16660), .B(n16663), .Z(n1668) );
  XOR U3399 ( .A(n16660), .B(n16663), .Z(n1669) );
  NANDN U3400 ( .A(n16661), .B(n1669), .Z(n1670) );
  NAND U3401 ( .A(n1668), .B(n1670), .Z(n16334) );
  XNOR U3402 ( .A(n16367), .B(n16368), .Z(n16369) );
  NAND U3403 ( .A(n16001), .B(n16004), .Z(n1671) );
  XOR U3404 ( .A(n16001), .B(n16004), .Z(n1672) );
  NANDN U3405 ( .A(n16002), .B(n1672), .Z(n1673) );
  NAND U3406 ( .A(n1671), .B(n1673), .Z(n15678) );
  XNOR U3407 ( .A(n5731), .B(n5732), .Z(n6031) );
  XNOR U3408 ( .A(n5163), .B(n5164), .Z(n5452) );
  XNOR U3409 ( .A(n4621), .B(n4622), .Z(n4898) );
  XNOR U3410 ( .A(n4103), .B(n4104), .Z(n4367) );
  XNOR U3411 ( .A(n22667), .B(n22666), .Z(n22661) );
  XOR U3412 ( .A(n16275), .B(n16272), .Z(n1674) );
  NANDN U3413 ( .A(n16273), .B(n1674), .Z(n1675) );
  NAND U3414 ( .A(n16275), .B(n16272), .Z(n1676) );
  AND U3415 ( .A(n1675), .B(n1676), .Z(n15910) );
  XOR U3416 ( .A(n16301), .B(n16302), .Z(n1677) );
  XNOR U3417 ( .A(n16300), .B(n1677), .Z(n16484) );
  XNOR U3418 ( .A(n16691), .B(n16692), .Z(n16827) );
  XOR U3419 ( .A(n15445), .B(n15442), .Z(n1678) );
  NAND U3420 ( .A(n1678), .B(n15443), .Z(n1679) );
  NAND U3421 ( .A(n15445), .B(n15442), .Z(n1680) );
  AND U3422 ( .A(n1679), .B(n1680), .Z(n15318) );
  NAND U3423 ( .A(n14301), .B(n14300), .Z(n1681) );
  NANDN U3424 ( .A(n14614), .B(n14613), .Z(n1682) );
  AND U3425 ( .A(n1681), .B(n1682), .Z(n14305) );
  NAND U3426 ( .A(n13584), .B(n13583), .Z(n1683) );
  NANDN U3427 ( .A(n13251), .B(n13252), .Z(n1684) );
  AND U3428 ( .A(n1683), .B(n1684), .Z(n13253) );
  NAND U3429 ( .A(n13582), .B(n13581), .Z(n1685) );
  NANDN U3430 ( .A(n13941), .B(n13940), .Z(n1686) );
  AND U3431 ( .A(n1685), .B(n1686), .Z(n13586) );
  NAND U3432 ( .A(n12791), .B(n12790), .Z(n1687) );
  NANDN U3433 ( .A(n13255), .B(n13256), .Z(n1688) );
  NAND U3434 ( .A(n1687), .B(n1688), .Z(n13003) );
  XNOR U3435 ( .A(n5450), .B(n5451), .Z(n5745) );
  XNOR U3436 ( .A(n4896), .B(n4897), .Z(n5177) );
  XNOR U3437 ( .A(n4368), .B(n4369), .Z(n4636) );
  XNOR U3438 ( .A(n22653), .B(n22652), .Z(n22654) );
  XOR U3439 ( .A(n16602), .B(n16599), .Z(n1689) );
  NANDN U3440 ( .A(n16600), .B(n1689), .Z(n1690) );
  NAND U3441 ( .A(n16602), .B(n16599), .Z(n1691) );
  AND U3442 ( .A(n1690), .B(n1691), .Z(n16267) );
  XNOR U3443 ( .A(n16278), .B(n16279), .Z(n16489) );
  XNOR U3444 ( .A(n17040), .B(n17041), .Z(n17042) );
  NAND U3445 ( .A(n17371), .B(n17374), .Z(n1692) );
  XOR U3446 ( .A(n17371), .B(n17374), .Z(n1693) );
  NANDN U3447 ( .A(n17372), .B(n1693), .Z(n1694) );
  NAND U3448 ( .A(n1692), .B(n1694), .Z(n17032) );
  XOR U3449 ( .A(n17052), .B(n17053), .Z(n1695) );
  XNOR U3450 ( .A(n17051), .B(n1695), .Z(n17160) );
  XNOR U3451 ( .A(n16469), .B(n16470), .Z(n17058) );
  NAND U3452 ( .A(n16703), .B(n16706), .Z(n1696) );
  XOR U3453 ( .A(n16703), .B(n16706), .Z(n1697) );
  NANDN U3454 ( .A(n16704), .B(n1697), .Z(n1698) );
  NAND U3455 ( .A(n1696), .B(n1698), .Z(n16378) );
  XNOR U3456 ( .A(n6640), .B(n6641), .Z(n6960) );
  XNOR U3457 ( .A(n6036), .B(n6037), .Z(n6341) );
  XNOR U3458 ( .A(n5743), .B(n5744), .Z(n6044) );
  XNOR U3459 ( .A(n5175), .B(n5176), .Z(n5464) );
  XNOR U3460 ( .A(n4633), .B(n4634), .Z(n4909) );
  XNOR U3461 ( .A(n22647), .B(n22646), .Z(n22648) );
  XOR U3462 ( .A(n16952), .B(n16949), .Z(n1699) );
  NANDN U3463 ( .A(n16950), .B(n1699), .Z(n1700) );
  NAND U3464 ( .A(n16952), .B(n16949), .Z(n1701) );
  AND U3465 ( .A(n1700), .B(n1701), .Z(n16604) );
  XOR U3466 ( .A(n16968), .B(n16965), .Z(n1702) );
  NANDN U3467 ( .A(n16966), .B(n1702), .Z(n1703) );
  NAND U3468 ( .A(n16968), .B(n16965), .Z(n1704) );
  AND U3469 ( .A(n1703), .B(n1704), .Z(n16620) );
  XOR U3470 ( .A(n16152), .B(n16153), .Z(n1705) );
  XNOR U3471 ( .A(n16151), .B(n1705), .Z(n16627) );
  XOR U3472 ( .A(n17001), .B(n17000), .Z(n1706) );
  NANDN U3473 ( .A(n17003), .B(n1706), .Z(n1707) );
  NAND U3474 ( .A(n17001), .B(n17000), .Z(n1708) );
  AND U3475 ( .A(n1707), .B(n1708), .Z(n17008) );
  XOR U3476 ( .A(n16648), .B(n16647), .Z(n1709) );
  XNOR U3477 ( .A(n16649), .B(n1709), .Z(n16835) );
  XOR U3478 ( .A(n17729), .B(n17731), .Z(n1710) );
  NANDN U3479 ( .A(n17730), .B(n1710), .Z(n1711) );
  NAND U3480 ( .A(n17729), .B(n17731), .Z(n1712) );
  AND U3481 ( .A(n1711), .B(n1712), .Z(n17370) );
  NAND U3482 ( .A(n16386), .B(n16388), .Z(n1713) );
  XOR U3483 ( .A(n16386), .B(n16388), .Z(n1714) );
  NANDN U3484 ( .A(n16385), .B(n1714), .Z(n1715) );
  NAND U3485 ( .A(n1713), .B(n1715), .Z(n16016) );
  XNOR U3486 ( .A(n6957), .B(n6958), .Z(n7007) );
  XNOR U3487 ( .A(n6339), .B(n6340), .Z(n6652) );
  XNOR U3488 ( .A(n5462), .B(n5463), .Z(n5757) );
  XNOR U3489 ( .A(n4910), .B(n4911), .Z(n5190) );
  XNOR U3490 ( .A(n22641), .B(n22640), .Z(n22643) );
  XOR U3491 ( .A(n17286), .B(n17283), .Z(n1716) );
  NANDN U3492 ( .A(n17284), .B(n1716), .Z(n1717) );
  NAND U3493 ( .A(n17286), .B(n17283), .Z(n1718) );
  AND U3494 ( .A(n1717), .B(n1718), .Z(n16954) );
  NAND U3495 ( .A(n17301), .B(n17304), .Z(n1719) );
  XOR U3496 ( .A(n17301), .B(n17304), .Z(n1720) );
  NANDN U3497 ( .A(n17302), .B(n1720), .Z(n1721) );
  NAND U3498 ( .A(n1719), .B(n1721), .Z(n16970) );
  XOR U3499 ( .A(n16989), .B(n16990), .Z(n1722) );
  XNOR U3500 ( .A(n16988), .B(n1722), .Z(n16991) );
  XNOR U3501 ( .A(n16981), .B(n16982), .Z(n1723) );
  XNOR U3502 ( .A(n16983), .B(n1723), .Z(n17172) );
  XNOR U3503 ( .A(n17745), .B(n17746), .Z(n1724) );
  XNOR U3504 ( .A(n17744), .B(n1724), .Z(n17847) );
  XOR U3505 ( .A(n17401), .B(n17400), .Z(n1725) );
  XNOR U3506 ( .A(n17402), .B(n1725), .Z(n17522) );
  NAND U3507 ( .A(n17407), .B(n17410), .Z(n1726) );
  XOR U3508 ( .A(n17407), .B(n17410), .Z(n1727) );
  NANDN U3509 ( .A(n17408), .B(n1727), .Z(n1728) );
  NAND U3510 ( .A(n1726), .B(n1728), .Z(n17074) );
  XNOR U3511 ( .A(n6650), .B(n6651), .Z(n6969) );
  XNOR U3512 ( .A(n6050), .B(n6051), .Z(n6354) );
  XNOR U3513 ( .A(n5755), .B(n5756), .Z(n6056) );
  XNOR U3514 ( .A(n5187), .B(n5188), .Z(n5475) );
  XNOR U3515 ( .A(n22695), .B(n22694), .Z(n22696) );
  NAND U3516 ( .A(n17655), .B(n17658), .Z(n1729) );
  XOR U3517 ( .A(n17655), .B(n17658), .Z(n1730) );
  NANDN U3518 ( .A(n17656), .B(n1730), .Z(n1731) );
  NAND U3519 ( .A(n1729), .B(n1731), .Z(n17288) );
  NAND U3520 ( .A(n17672), .B(n17670), .Z(n1732) );
  XOR U3521 ( .A(n17672), .B(n17670), .Z(n1733) );
  NANDN U3522 ( .A(n17669), .B(n1733), .Z(n1734) );
  NAND U3523 ( .A(n1732), .B(n1734), .Z(n17306) );
  XOR U3524 ( .A(n17688), .B(n17685), .Z(n1735) );
  NANDN U3525 ( .A(n17686), .B(n1735), .Z(n1736) );
  NAND U3526 ( .A(n17688), .B(n17685), .Z(n1737) );
  AND U3527 ( .A(n1736), .B(n1737), .Z(n17322) );
  XNOR U3528 ( .A(n17734), .B(n17735), .Z(n17849) );
  XOR U3529 ( .A(n17758), .B(n17759), .Z(n1738) );
  XNOR U3530 ( .A(n17757), .B(n1738), .Z(n17843) );
  NAND U3531 ( .A(n15010), .B(n15009), .Z(n1739) );
  NANDN U3532 ( .A(n15336), .B(n15335), .Z(n1740) );
  AND U3533 ( .A(n1739), .B(n1740), .Z(n15014) );
  NAND U3534 ( .A(n17082), .B(n17084), .Z(n1741) );
  XOR U3535 ( .A(n17082), .B(n17084), .Z(n1742) );
  NANDN U3536 ( .A(n17081), .B(n1742), .Z(n1743) );
  NAND U3537 ( .A(n1741), .B(n1743), .Z(n16720) );
  NAND U3538 ( .A(n16132), .B(n16131), .Z(n1744) );
  XOR U3539 ( .A(n16132), .B(n16131), .Z(n1745) );
  NAND U3540 ( .A(n1745), .B(n16134), .Z(n1746) );
  NAND U3541 ( .A(n1744), .B(n1746), .Z(n16030) );
  NAND U3542 ( .A(n14317), .B(n14316), .Z(n1747) );
  NANDN U3543 ( .A(n14638), .B(n14637), .Z(n1748) );
  AND U3544 ( .A(n1747), .B(n1748), .Z(n14321) );
  NAND U3545 ( .A(n13600), .B(n13599), .Z(n1749) );
  NANDN U3546 ( .A(n13271), .B(n13272), .Z(n1750) );
  AND U3547 ( .A(n1749), .B(n1750), .Z(n13273) );
  NAND U3548 ( .A(n13598), .B(n13597), .Z(n1751) );
  NANDN U3549 ( .A(n13965), .B(n13964), .Z(n1752) );
  AND U3550 ( .A(n1751), .B(n1752), .Z(n13602) );
  NAND U3551 ( .A(n12783), .B(n12782), .Z(n1753) );
  NANDN U3552 ( .A(n13275), .B(n13276), .Z(n1754) );
  NAND U3553 ( .A(n1753), .B(n1754), .Z(n13011) );
  XNOR U3554 ( .A(n6967), .B(n6968), .Z(n7003) );
  XNOR U3555 ( .A(n6351), .B(n6352), .Z(n6662) );
  XNOR U3556 ( .A(n5476), .B(n5477), .Z(n5770) );
  XNOR U3557 ( .A(n22635), .B(n22634), .Z(n22636) );
  NAND U3558 ( .A(n17976), .B(n17979), .Z(n1755) );
  XOR U3559 ( .A(n17976), .B(n17979), .Z(n1756) );
  NANDN U3560 ( .A(n17977), .B(n1756), .Z(n1757) );
  NAND U3561 ( .A(n1755), .B(n1757), .Z(n17654) );
  NAND U3562 ( .A(n17992), .B(n17995), .Z(n1758) );
  XOR U3563 ( .A(n17992), .B(n17995), .Z(n1759) );
  NANDN U3564 ( .A(n17993), .B(n1759), .Z(n1760) );
  NAND U3565 ( .A(n1758), .B(n1760), .Z(n17674) );
  NAND U3566 ( .A(n18008), .B(n18011), .Z(n1761) );
  XOR U3567 ( .A(n18008), .B(n18011), .Z(n1762) );
  NANDN U3568 ( .A(n18009), .B(n1762), .Z(n1763) );
  NAND U3569 ( .A(n1761), .B(n1763), .Z(n17690) );
  NAND U3570 ( .A(n18024), .B(n18027), .Z(n1764) );
  XOR U3571 ( .A(n18024), .B(n18027), .Z(n1765) );
  NANDN U3572 ( .A(n18025), .B(n1765), .Z(n1766) );
  NAND U3573 ( .A(n1764), .B(n1766), .Z(n17706) );
  XOR U3574 ( .A(n17334), .B(n17335), .Z(n1767) );
  XNOR U3575 ( .A(n17333), .B(n1767), .Z(n17536) );
  XOR U3576 ( .A(n18053), .B(n18052), .Z(n1768) );
  XNOR U3577 ( .A(n18054), .B(n1768), .Z(n18193) );
  NAND U3578 ( .A(n18092), .B(n18095), .Z(n1769) );
  XOR U3579 ( .A(n18092), .B(n18095), .Z(n1770) );
  NANDN U3580 ( .A(n18093), .B(n1770), .Z(n1771) );
  NAND U3581 ( .A(n1769), .B(n1771), .Z(n17773) );
  XOR U3582 ( .A(n7615), .B(n7616), .Z(n7618) );
  XNOR U3583 ( .A(n6062), .B(n6063), .Z(n6366) );
  XNOR U3584 ( .A(n6664), .B(n6665), .Z(n6979) );
  XNOR U3585 ( .A(n5767), .B(n5768), .Z(n6067) );
  XNOR U3586 ( .A(n22629), .B(n22628), .Z(n22630) );
  XOR U3587 ( .A(n18325), .B(n18323), .Z(n1772) );
  NANDN U3588 ( .A(n18322), .B(n1772), .Z(n1773) );
  NAND U3589 ( .A(n18325), .B(n18323), .Z(n1774) );
  AND U3590 ( .A(n1773), .B(n1774), .Z(n17981) );
  NAND U3591 ( .A(n18340), .B(n18343), .Z(n1775) );
  XOR U3592 ( .A(n18340), .B(n18343), .Z(n1776) );
  NANDN U3593 ( .A(n18341), .B(n1776), .Z(n1777) );
  NAND U3594 ( .A(n1775), .B(n1777), .Z(n17997) );
  XOR U3595 ( .A(n18357), .B(n18354), .Z(n1778) );
  NANDN U3596 ( .A(n18355), .B(n1778), .Z(n1779) );
  NAND U3597 ( .A(n18357), .B(n18354), .Z(n1780) );
  AND U3598 ( .A(n1779), .B(n1780), .Z(n18013) );
  NAND U3599 ( .A(n18370), .B(n18373), .Z(n1781) );
  XOR U3600 ( .A(n18370), .B(n18373), .Z(n1782) );
  NANDN U3601 ( .A(n18371), .B(n1782), .Z(n1783) );
  NAND U3602 ( .A(n1781), .B(n1783), .Z(n18029) );
  XOR U3603 ( .A(n17717), .B(n17718), .Z(n1784) );
  XNOR U3604 ( .A(n17716), .B(n1784), .Z(n18039) );
  XOR U3605 ( .A(n18401), .B(n18402), .Z(n1785) );
  XNOR U3606 ( .A(n18400), .B(n1785), .Z(n18720) );
  XOR U3607 ( .A(n18743), .B(n18744), .Z(n1786) );
  XNOR U3608 ( .A(n18742), .B(n1786), .Z(n19091) );
  XNOR U3609 ( .A(n18749), .B(n18750), .Z(n18751) );
  XNOR U3610 ( .A(n18442), .B(n18443), .Z(n1787) );
  XNOR U3611 ( .A(n18441), .B(n1787), .Z(n18497) );
  NAND U3612 ( .A(n19108), .B(n19111), .Z(n1788) );
  XOR U3613 ( .A(n19108), .B(n19111), .Z(n1789) );
  NANDN U3614 ( .A(n19109), .B(n1789), .Z(n1790) );
  NAND U3615 ( .A(n1788), .B(n1790), .Z(n18761) );
  NAND U3616 ( .A(n17779), .B(n17781), .Z(n1791) );
  XOR U3617 ( .A(n17779), .B(n17781), .Z(n1792) );
  NANDN U3618 ( .A(n17778), .B(n1792), .Z(n1793) );
  NAND U3619 ( .A(n1791), .B(n1793), .Z(n17424) );
  NAND U3620 ( .A(n15708), .B(n15707), .Z(n1794) );
  NANDN U3621 ( .A(n16036), .B(n16035), .Z(n1795) );
  AND U3622 ( .A(n1794), .B(n1795), .Z(n15712) );
  XNOR U3623 ( .A(n6363), .B(n6364), .Z(n6675) );
  XNOR U3624 ( .A(n22623), .B(n22622), .Z(n22625) );
  XNOR U3625 ( .A(n19548), .B(n19549), .Z(n19551) );
  NAND U3626 ( .A(n18629), .B(n18632), .Z(n1796) );
  XOR U3627 ( .A(n18629), .B(n18632), .Z(n1797) );
  NANDN U3628 ( .A(n18630), .B(n1797), .Z(n1798) );
  NAND U3629 ( .A(n1796), .B(n1798), .Z(n18320) );
  NAND U3630 ( .A(n18645), .B(n18648), .Z(n1799) );
  XOR U3631 ( .A(n18645), .B(n18648), .Z(n1800) );
  NANDN U3632 ( .A(n18646), .B(n1800), .Z(n1801) );
  NAND U3633 ( .A(n1799), .B(n1801), .Z(n18339) );
  NAND U3634 ( .A(n18661), .B(n18664), .Z(n1802) );
  XOR U3635 ( .A(n18661), .B(n18664), .Z(n1803) );
  NANDN U3636 ( .A(n18662), .B(n1803), .Z(n1804) );
  NAND U3637 ( .A(n1802), .B(n1804), .Z(n18359) );
  NAND U3638 ( .A(n18677), .B(n18680), .Z(n1805) );
  XOR U3639 ( .A(n18677), .B(n18680), .Z(n1806) );
  NANDN U3640 ( .A(n18678), .B(n1806), .Z(n1807) );
  NAND U3641 ( .A(n1805), .B(n1807), .Z(n18375) );
  XNOR U3642 ( .A(n18386), .B(n18387), .Z(n1808) );
  XNOR U3643 ( .A(n18388), .B(n1808), .Z(n18508) );
  XNOR U3644 ( .A(n19082), .B(n19083), .Z(n19171) );
  NAND U3645 ( .A(n15026), .B(n15025), .Z(n1809) );
  NANDN U3646 ( .A(n15360), .B(n15359), .Z(n1810) );
  AND U3647 ( .A(n1809), .B(n1810), .Z(n15030) );
  XNOR U3648 ( .A(n7627), .B(n7628), .Z(n7658) );
  XOR U3649 ( .A(n7659), .B(n7660), .Z(n7961) );
  XNOR U3650 ( .A(n6676), .B(n6677), .Z(n6994) );
  XNOR U3651 ( .A(n22617), .B(n22616), .Z(n22618) );
  NAND U3652 ( .A(n18962), .B(n18965), .Z(n1811) );
  XOR U3653 ( .A(n18962), .B(n18965), .Z(n1812) );
  NANDN U3654 ( .A(n18963), .B(n1812), .Z(n1813) );
  NAND U3655 ( .A(n1811), .B(n1813), .Z(n18634) );
  XOR U3656 ( .A(n18983), .B(n18981), .Z(n1814) );
  NANDN U3657 ( .A(n18980), .B(n1814), .Z(n1815) );
  NAND U3658 ( .A(n18983), .B(n18981), .Z(n1816) );
  AND U3659 ( .A(n1815), .B(n1816), .Z(n18650) );
  NAND U3660 ( .A(n18996), .B(n18999), .Z(n1817) );
  XOR U3661 ( .A(n18996), .B(n18999), .Z(n1818) );
  NANDN U3662 ( .A(n18997), .B(n1818), .Z(n1819) );
  NAND U3663 ( .A(n1817), .B(n1819), .Z(n18666) );
  XOR U3664 ( .A(n19017), .B(n19015), .Z(n1820) );
  NANDN U3665 ( .A(n19014), .B(n1820), .Z(n1821) );
  NAND U3666 ( .A(n19017), .B(n19015), .Z(n1822) );
  AND U3667 ( .A(n1821), .B(n1822), .Z(n18682) );
  NAND U3668 ( .A(n19030), .B(n19033), .Z(n1823) );
  XOR U3669 ( .A(n19030), .B(n19033), .Z(n1824) );
  NANDN U3670 ( .A(n19031), .B(n1824), .Z(n1825) );
  NAND U3671 ( .A(n1823), .B(n1825), .Z(n18698) );
  XOR U3672 ( .A(n19049), .B(n19046), .Z(n1826) );
  NANDN U3673 ( .A(n19047), .B(n1826), .Z(n1827) );
  NAND U3674 ( .A(n19049), .B(n19046), .Z(n1828) );
  AND U3675 ( .A(n1827), .B(n1828), .Z(n19055) );
  XOR U3676 ( .A(n18839), .B(n18838), .Z(n1829) );
  NANDN U3677 ( .A(n18841), .B(n1829), .Z(n1830) );
  NAND U3678 ( .A(n18839), .B(n18838), .Z(n1831) );
  AND U3679 ( .A(n1830), .B(n1831), .Z(n19072) );
  XOR U3680 ( .A(n19425), .B(n19426), .Z(n1832) );
  XNOR U3681 ( .A(n19424), .B(n1832), .Z(n19505) );
  XNOR U3682 ( .A(n19106), .B(n19107), .Z(n19167) );
  XNOR U3683 ( .A(n18776), .B(n18777), .Z(n19125) );
  NAND U3684 ( .A(n16814), .B(n16813), .Z(n1833) );
  XOR U3685 ( .A(n16814), .B(n16813), .Z(n1834) );
  NANDN U3686 ( .A(n16816), .B(n1834), .Z(n1835) );
  NAND U3687 ( .A(n1833), .B(n1835), .Z(n16746) );
  NAND U3688 ( .A(n14333), .B(n14332), .Z(n1836) );
  NANDN U3689 ( .A(n14662), .B(n14661), .Z(n1837) );
  AND U3690 ( .A(n1836), .B(n1837), .Z(n14337) );
  NAND U3691 ( .A(n13616), .B(n13615), .Z(n1838) );
  NANDN U3692 ( .A(n13291), .B(n13292), .Z(n1839) );
  AND U3693 ( .A(n1838), .B(n1839), .Z(n13293) );
  NAND U3694 ( .A(n13614), .B(n13613), .Z(n1840) );
  NANDN U3695 ( .A(n13989), .B(n13988), .Z(n1841) );
  AND U3696 ( .A(n1840), .B(n1841), .Z(n13618) );
  NAND U3697 ( .A(n12775), .B(n12774), .Z(n1842) );
  NANDN U3698 ( .A(n13295), .B(n13296), .Z(n1843) );
  NAND U3699 ( .A(n1842), .B(n1843), .Z(n13019) );
  NAND U3700 ( .A(n8297), .B(n8298), .Z(n1844) );
  NANDN U3701 ( .A(n8334), .B(n8333), .Z(n1845) );
  AND U3702 ( .A(n1844), .B(n1845), .Z(n8332) );
  XNOR U3703 ( .A(n6991), .B(n6992), .Z(n7314) );
  XNOR U3704 ( .A(n22611), .B(n22610), .Z(n22612) );
  NAND U3705 ( .A(n19301), .B(n19304), .Z(n1846) );
  XOR U3706 ( .A(n19301), .B(n19304), .Z(n1847) );
  NANDN U3707 ( .A(n19302), .B(n1847), .Z(n1848) );
  NAND U3708 ( .A(n1846), .B(n1848), .Z(n18967) );
  NAND U3709 ( .A(n19317), .B(n19320), .Z(n1849) );
  XOR U3710 ( .A(n19317), .B(n19320), .Z(n1850) );
  NANDN U3711 ( .A(n19318), .B(n1850), .Z(n1851) );
  NAND U3712 ( .A(n1849), .B(n1851), .Z(n18978) );
  NAND U3713 ( .A(n19336), .B(n19338), .Z(n1852) );
  XOR U3714 ( .A(n19336), .B(n19338), .Z(n1853) );
  NANDN U3715 ( .A(n19335), .B(n1853), .Z(n1854) );
  NAND U3716 ( .A(n1852), .B(n1854), .Z(n19001) );
  NAND U3717 ( .A(n19351), .B(n19354), .Z(n1855) );
  XOR U3718 ( .A(n19351), .B(n19354), .Z(n1856) );
  NANDN U3719 ( .A(n19352), .B(n1856), .Z(n1857) );
  NAND U3720 ( .A(n1855), .B(n1857), .Z(n19012) );
  NAND U3721 ( .A(n19367), .B(n19370), .Z(n1858) );
  XOR U3722 ( .A(n19367), .B(n19370), .Z(n1859) );
  NANDN U3723 ( .A(n19368), .B(n1859), .Z(n1860) );
  NAND U3724 ( .A(n1858), .B(n1860), .Z(n19035) );
  NAND U3725 ( .A(n19385), .B(n19388), .Z(n1861) );
  XOR U3726 ( .A(n19385), .B(n19388), .Z(n1862) );
  NANDN U3727 ( .A(n19386), .B(n1862), .Z(n1863) );
  NAND U3728 ( .A(n1861), .B(n1863), .Z(n19051) );
  NAND U3729 ( .A(n19786), .B(n19788), .Z(n1864) );
  XOR U3730 ( .A(n19786), .B(n19788), .Z(n1865) );
  NANDN U3731 ( .A(n19785), .B(n1865), .Z(n1866) );
  NAND U3732 ( .A(n1864), .B(n1866), .Z(n19440) );
  NAND U3733 ( .A(n19442), .B(n19444), .Z(n1867) );
  XOR U3734 ( .A(n19442), .B(n19444), .Z(n1868) );
  NANDN U3735 ( .A(n19441), .B(n1868), .Z(n1869) );
  NAND U3736 ( .A(n1867), .B(n1869), .Z(n19127) );
  XOR U3737 ( .A(n18181), .B(n18178), .Z(n1870) );
  NAND U3738 ( .A(n1870), .B(n18179), .Z(n1871) );
  NAND U3739 ( .A(n18181), .B(n18178), .Z(n1872) );
  AND U3740 ( .A(n1871), .B(n1872), .Z(n18109) );
  NAND U3741 ( .A(n18456), .B(n18455), .Z(n1873) );
  NANDN U3742 ( .A(n18493), .B(n18494), .Z(n1874) );
  NAND U3743 ( .A(n1873), .B(n1874), .Z(n18781) );
  NAND U3744 ( .A(n15724), .B(n15723), .Z(n1875) );
  NANDN U3745 ( .A(n16060), .B(n16059), .Z(n1876) );
  AND U3746 ( .A(n1875), .B(n1876), .Z(n15728) );
  XNOR U3747 ( .A(n8303), .B(n8304), .Z(n8330) );
  XNOR U3748 ( .A(n7655), .B(n7656), .Z(n7968) );
  XOR U3749 ( .A(n7637), .B(n7638), .Z(n7975) );
  XNOR U3750 ( .A(n6997), .B(n6998), .Z(n7321) );
  XNOR U3751 ( .A(n22605), .B(n22604), .Z(n22606) );
  XNOR U3752 ( .A(n20222), .B(n20223), .Z(n20550) );
  NAND U3753 ( .A(n19638), .B(n19641), .Z(n1877) );
  XOR U3754 ( .A(n19638), .B(n19641), .Z(n1878) );
  NANDN U3755 ( .A(n19639), .B(n1878), .Z(n1879) );
  NAND U3756 ( .A(n1877), .B(n1879), .Z(n19306) );
  NAND U3757 ( .A(n19654), .B(n19657), .Z(n1880) );
  XOR U3758 ( .A(n19654), .B(n19657), .Z(n1881) );
  NANDN U3759 ( .A(n19655), .B(n1881), .Z(n1882) );
  NAND U3760 ( .A(n1880), .B(n1882), .Z(n19322) );
  NAND U3761 ( .A(n19671), .B(n19673), .Z(n1883) );
  XOR U3762 ( .A(n19671), .B(n19673), .Z(n1884) );
  NANDN U3763 ( .A(n19670), .B(n1884), .Z(n1885) );
  NAND U3764 ( .A(n1883), .B(n1885), .Z(n19340) );
  NAND U3765 ( .A(n19688), .B(n19691), .Z(n1886) );
  XOR U3766 ( .A(n19688), .B(n19691), .Z(n1887) );
  NANDN U3767 ( .A(n19689), .B(n1887), .Z(n1888) );
  NAND U3768 ( .A(n1886), .B(n1888), .Z(n19356) );
  NAND U3769 ( .A(n19704), .B(n19707), .Z(n1889) );
  XOR U3770 ( .A(n19704), .B(n19707), .Z(n1890) );
  NANDN U3771 ( .A(n19705), .B(n1890), .Z(n1891) );
  NAND U3772 ( .A(n1889), .B(n1891), .Z(n19372) );
  NAND U3773 ( .A(n19723), .B(n19721), .Z(n1892) );
  XOR U3774 ( .A(n19723), .B(n19721), .Z(n1893) );
  NANDN U3775 ( .A(n19720), .B(n1893), .Z(n1894) );
  NAND U3776 ( .A(n1892), .B(n1894), .Z(n19390) );
  XOR U3777 ( .A(n19178), .B(n19175), .Z(n1895) );
  NAND U3778 ( .A(n1895), .B(n19176), .Z(n1896) );
  NAND U3779 ( .A(n19178), .B(n19175), .Z(n1897) );
  AND U3780 ( .A(n1896), .B(n1897), .Z(n19402) );
  XOR U3781 ( .A(n19410), .B(n19411), .Z(n1898) );
  XNOR U3782 ( .A(n19409), .B(n1898), .Z(n19755) );
  NAND U3783 ( .A(n20106), .B(n20109), .Z(n1899) );
  XOR U3784 ( .A(n20106), .B(n20109), .Z(n1900) );
  NANDN U3785 ( .A(n20107), .B(n1900), .Z(n1901) );
  NAND U3786 ( .A(n1899), .B(n1901), .Z(n19784) );
  NAND U3787 ( .A(n20440), .B(n20443), .Z(n1902) );
  XOR U3788 ( .A(n20440), .B(n20443), .Z(n1903) );
  NANDN U3789 ( .A(n20441), .B(n1903), .Z(n1904) );
  NAND U3790 ( .A(n1902), .B(n1904), .Z(n20111) );
  XNOR U3791 ( .A(n22599), .B(n22598), .Z(n22601) );
  XNOR U3792 ( .A(n20228), .B(n20229), .Z(n20556) );
  NAND U3793 ( .A(n20572), .B(n20571), .Z(n1905) );
  NANDN U3794 ( .A(n20241), .B(n20240), .Z(n1906) );
  AND U3795 ( .A(n1905), .B(n1906), .Z(n20245) );
  NAND U3796 ( .A(n19971), .B(n19974), .Z(n1907) );
  XOR U3797 ( .A(n19971), .B(n19974), .Z(n1908) );
  NANDN U3798 ( .A(n19972), .B(n1908), .Z(n1909) );
  NAND U3799 ( .A(n1907), .B(n1909), .Z(n19643) );
  NAND U3800 ( .A(n19987), .B(n19990), .Z(n1910) );
  XOR U3801 ( .A(n19987), .B(n19990), .Z(n1911) );
  NANDN U3802 ( .A(n19988), .B(n1911), .Z(n1912) );
  NAND U3803 ( .A(n1910), .B(n1912), .Z(n19659) );
  NAND U3804 ( .A(n20004), .B(n20006), .Z(n1913) );
  XOR U3805 ( .A(n20004), .B(n20006), .Z(n1914) );
  NANDN U3806 ( .A(n20003), .B(n1914), .Z(n1915) );
  NAND U3807 ( .A(n1913), .B(n1915), .Z(n19675) );
  XOR U3808 ( .A(n20022), .B(n20019), .Z(n1916) );
  NANDN U3809 ( .A(n20020), .B(n1916), .Z(n1917) );
  NAND U3810 ( .A(n20022), .B(n20019), .Z(n1918) );
  AND U3811 ( .A(n1917), .B(n1918), .Z(n19693) );
  NAND U3812 ( .A(n20035), .B(n20038), .Z(n1919) );
  XOR U3813 ( .A(n20035), .B(n20038), .Z(n1920) );
  NANDN U3814 ( .A(n20036), .B(n1920), .Z(n1921) );
  NAND U3815 ( .A(n1919), .B(n1921), .Z(n19709) );
  NAND U3816 ( .A(n20051), .B(n20054), .Z(n1922) );
  XOR U3817 ( .A(n20051), .B(n20054), .Z(n1923) );
  NANDN U3818 ( .A(n20052), .B(n1923), .Z(n1924) );
  NAND U3819 ( .A(n1922), .B(n1924), .Z(n19725) );
  NAND U3820 ( .A(n20067), .B(n20070), .Z(n1925) );
  XOR U3821 ( .A(n20067), .B(n20070), .Z(n1926) );
  NANDN U3822 ( .A(n20068), .B(n1926), .Z(n1927) );
  NAND U3823 ( .A(n1925), .B(n1927), .Z(n19740) );
  XOR U3824 ( .A(n19833), .B(n19834), .Z(n1928) );
  NANDN U3825 ( .A(n19836), .B(n1928), .Z(n1929) );
  NAND U3826 ( .A(n19833), .B(n19834), .Z(n1930) );
  AND U3827 ( .A(n1929), .B(n1930), .Z(n20093) );
  NAND U3828 ( .A(n15042), .B(n15041), .Z(n1931) );
  NANDN U3829 ( .A(n15384), .B(n15383), .Z(n1932) );
  AND U3830 ( .A(n1931), .B(n1932), .Z(n15046) );
  XNOR U3831 ( .A(n8654), .B(n8655), .Z(n8679) );
  XNOR U3832 ( .A(n22593), .B(n22592), .Z(n22594) );
  XOR U3833 ( .A(n20301), .B(n20298), .Z(n1933) );
  NANDN U3834 ( .A(n20299), .B(n1933), .Z(n1934) );
  NAND U3835 ( .A(n20301), .B(n20298), .Z(n1935) );
  AND U3836 ( .A(n1934), .B(n1935), .Z(n19976) );
  XOR U3837 ( .A(n20317), .B(n20314), .Z(n1936) );
  NANDN U3838 ( .A(n20315), .B(n1936), .Z(n1937) );
  NAND U3839 ( .A(n20317), .B(n20314), .Z(n1938) );
  AND U3840 ( .A(n1937), .B(n1938), .Z(n19992) );
  NAND U3841 ( .A(n20330), .B(n20333), .Z(n1939) );
  XOR U3842 ( .A(n20330), .B(n20333), .Z(n1940) );
  NANDN U3843 ( .A(n20331), .B(n1940), .Z(n1941) );
  NAND U3844 ( .A(n1939), .B(n1941), .Z(n20008) );
  NAND U3845 ( .A(n20349), .B(n20351), .Z(n1942) );
  XOR U3846 ( .A(n20349), .B(n20351), .Z(n1943) );
  NANDN U3847 ( .A(n20348), .B(n1943), .Z(n1944) );
  NAND U3848 ( .A(n1942), .B(n1944), .Z(n20024) );
  NAND U3849 ( .A(n20366), .B(n20369), .Z(n1945) );
  XOR U3850 ( .A(n20366), .B(n20369), .Z(n1946) );
  NANDN U3851 ( .A(n20367), .B(n1946), .Z(n1947) );
  NAND U3852 ( .A(n1945), .B(n1947), .Z(n20040) );
  NAND U3853 ( .A(n20382), .B(n20385), .Z(n1948) );
  XOR U3854 ( .A(n20382), .B(n20385), .Z(n1949) );
  NANDN U3855 ( .A(n20383), .B(n1949), .Z(n1950) );
  NAND U3856 ( .A(n1948), .B(n1950), .Z(n20056) );
  XOR U3857 ( .A(n20401), .B(n20398), .Z(n1951) );
  NANDN U3858 ( .A(n20399), .B(n1951), .Z(n1952) );
  NAND U3859 ( .A(n20401), .B(n20398), .Z(n1953) );
  AND U3860 ( .A(n1952), .B(n1953), .Z(n20072) );
  XOR U3861 ( .A(n20121), .B(n20122), .Z(n20123) );
  NAND U3862 ( .A(n19802), .B(n19804), .Z(n1954) );
  XOR U3863 ( .A(n19802), .B(n19804), .Z(n1955) );
  NANDN U3864 ( .A(n19801), .B(n1955), .Z(n1956) );
  NAND U3865 ( .A(n1954), .B(n1956), .Z(n19454) );
  NAND U3866 ( .A(n19137), .B(n19136), .Z(n1957) );
  NAND U3867 ( .A(n18785), .B(n18784), .Z(n1958) );
  AND U3868 ( .A(n1957), .B(n1958), .Z(n18827) );
  NAND U3869 ( .A(n16428), .B(n16427), .Z(n1959) );
  NANDN U3870 ( .A(n16764), .B(n16763), .Z(n1960) );
  AND U3871 ( .A(n1959), .B(n1960), .Z(n16432) );
  NAND U3872 ( .A(n14349), .B(n14348), .Z(n1961) );
  NANDN U3873 ( .A(n14686), .B(n14685), .Z(n1962) );
  AND U3874 ( .A(n1961), .B(n1962), .Z(n14353) );
  NAND U3875 ( .A(n13632), .B(n13631), .Z(n1963) );
  NANDN U3876 ( .A(n13311), .B(n13312), .Z(n1964) );
  AND U3877 ( .A(n1963), .B(n1964), .Z(n13313) );
  NAND U3878 ( .A(n13630), .B(n13629), .Z(n1965) );
  NANDN U3879 ( .A(n14013), .B(n14012), .Z(n1966) );
  AND U3880 ( .A(n1965), .B(n1966), .Z(n13634) );
  NAND U3881 ( .A(n12767), .B(n12766), .Z(n1967) );
  NANDN U3882 ( .A(n13315), .B(n13316), .Z(n1968) );
  NAND U3883 ( .A(n1967), .B(n1968), .Z(n13027) );
  NAND U3884 ( .A(n9006), .B(n9005), .Z(n1969) );
  NANDN U3885 ( .A(n9030), .B(n9029), .Z(n1970) );
  AND U3886 ( .A(n1969), .B(n1970), .Z(n9028) );
  XNOR U3887 ( .A(n8658), .B(n8659), .Z(n8660) );
  XOR U3888 ( .A(n20864), .B(n20865), .Z(n20887) );
  NAND U3889 ( .A(n20627), .B(n20630), .Z(n1971) );
  XOR U3890 ( .A(n20627), .B(n20630), .Z(n1972) );
  NANDN U3891 ( .A(n20628), .B(n1972), .Z(n1973) );
  NAND U3892 ( .A(n1971), .B(n1973), .Z(n20303) );
  NAND U3893 ( .A(n20644), .B(n20646), .Z(n1974) );
  XOR U3894 ( .A(n20644), .B(n20646), .Z(n1975) );
  NANDN U3895 ( .A(n20643), .B(n1975), .Z(n1976) );
  NAND U3896 ( .A(n1974), .B(n1976), .Z(n20319) );
  NAND U3897 ( .A(n20659), .B(n20662), .Z(n1977) );
  XOR U3898 ( .A(n20659), .B(n20662), .Z(n1978) );
  NANDN U3899 ( .A(n20660), .B(n1978), .Z(n1979) );
  NAND U3900 ( .A(n1977), .B(n1979), .Z(n20334) );
  NAND U3901 ( .A(n20675), .B(n20678), .Z(n1980) );
  XOR U3902 ( .A(n20675), .B(n20678), .Z(n1981) );
  NANDN U3903 ( .A(n20676), .B(n1981), .Z(n1982) );
  NAND U3904 ( .A(n1980), .B(n1982), .Z(n20352) );
  NAND U3905 ( .A(n20691), .B(n20694), .Z(n1983) );
  XOR U3906 ( .A(n20691), .B(n20694), .Z(n1984) );
  NANDN U3907 ( .A(n20692), .B(n1984), .Z(n1985) );
  NAND U3908 ( .A(n1983), .B(n1985), .Z(n20371) );
  NAND U3909 ( .A(n20707), .B(n20710), .Z(n1986) );
  XOR U3910 ( .A(n20707), .B(n20710), .Z(n1987) );
  NANDN U3911 ( .A(n20708), .B(n1987), .Z(n1988) );
  NAND U3912 ( .A(n1986), .B(n1988), .Z(n20387) );
  NAND U3913 ( .A(n20723), .B(n20726), .Z(n1989) );
  XOR U3914 ( .A(n20723), .B(n20726), .Z(n1990) );
  NANDN U3915 ( .A(n20724), .B(n1990), .Z(n1991) );
  NAND U3916 ( .A(n1989), .B(n1991), .Z(n20403) );
  NAND U3917 ( .A(n20739), .B(n20742), .Z(n1992) );
  XOR U3918 ( .A(n20739), .B(n20742), .Z(n1993) );
  NANDN U3919 ( .A(n20740), .B(n1993), .Z(n1994) );
  NAND U3920 ( .A(n1992), .B(n1994), .Z(n20421) );
  NAND U3921 ( .A(n20416), .B(n20419), .Z(n1995) );
  XOR U3922 ( .A(n20416), .B(n20419), .Z(n1996) );
  NANDN U3923 ( .A(n20417), .B(n1996), .Z(n1997) );
  NAND U3924 ( .A(n1995), .B(n1997), .Z(n20173) );
  XOR U3925 ( .A(n20432), .B(n20433), .Z(n1998) );
  XNOR U3926 ( .A(n20431), .B(n1998), .Z(n20761) );
  NAND U3927 ( .A(n20784), .B(n20787), .Z(n1999) );
  XOR U3928 ( .A(n20784), .B(n20787), .Z(n2000) );
  NANDN U3929 ( .A(n20785), .B(n2000), .Z(n2001) );
  NAND U3930 ( .A(n1999), .B(n2001), .Z(n20457) );
  XOR U3931 ( .A(n17508), .B(n17505), .Z(n2002) );
  NAND U3932 ( .A(n2002), .B(n17506), .Z(n2003) );
  NAND U3933 ( .A(n17508), .B(n17505), .Z(n2004) );
  AND U3934 ( .A(n2003), .B(n2004), .Z(n17462) );
  NAND U3935 ( .A(n15740), .B(n15739), .Z(n2005) );
  NANDN U3936 ( .A(n16084), .B(n16083), .Z(n2006) );
  AND U3937 ( .A(n2005), .B(n2006), .Z(n15744) );
  XOR U3938 ( .A(n8664), .B(n8665), .Z(n8667) );
  XNOR U3939 ( .A(n20876), .B(n20877), .Z(n21213) );
  NAND U3940 ( .A(n21265), .B(n21264), .Z(n2007) );
  NANDN U3941 ( .A(n20927), .B(n20926), .Z(n2008) );
  AND U3942 ( .A(n2007), .B(n2008), .Z(n20931) );
  NAND U3943 ( .A(n20960), .B(n20963), .Z(n2009) );
  XOR U3944 ( .A(n20960), .B(n20963), .Z(n2010) );
  NANDN U3945 ( .A(n20961), .B(n2010), .Z(n2011) );
  NAND U3946 ( .A(n2009), .B(n2011), .Z(n20632) );
  NAND U3947 ( .A(n20977), .B(n20979), .Z(n2012) );
  XOR U3948 ( .A(n20977), .B(n20979), .Z(n2013) );
  NANDN U3949 ( .A(n20976), .B(n2013), .Z(n2014) );
  NAND U3950 ( .A(n2012), .B(n2014), .Z(n20648) );
  NAND U3951 ( .A(n20994), .B(n20997), .Z(n2015) );
  XOR U3952 ( .A(n20994), .B(n20997), .Z(n2016) );
  NANDN U3953 ( .A(n20995), .B(n2016), .Z(n2017) );
  NAND U3954 ( .A(n2015), .B(n2017), .Z(n20664) );
  XOR U3955 ( .A(n21015), .B(n21013), .Z(n2018) );
  NANDN U3956 ( .A(n21012), .B(n2018), .Z(n2019) );
  NAND U3957 ( .A(n21015), .B(n21013), .Z(n2020) );
  AND U3958 ( .A(n2019), .B(n2020), .Z(n20680) );
  XOR U3959 ( .A(n21031), .B(n21028), .Z(n2021) );
  NANDN U3960 ( .A(n21029), .B(n2021), .Z(n2022) );
  NAND U3961 ( .A(n21031), .B(n21028), .Z(n2023) );
  AND U3962 ( .A(n2022), .B(n2023), .Z(n20696) );
  NAND U3963 ( .A(n21044), .B(n21047), .Z(n2024) );
  XOR U3964 ( .A(n21044), .B(n21047), .Z(n2025) );
  NANDN U3965 ( .A(n21045), .B(n2025), .Z(n2026) );
  NAND U3966 ( .A(n2024), .B(n2026), .Z(n20712) );
  NAND U3967 ( .A(n21060), .B(n21063), .Z(n2027) );
  XOR U3968 ( .A(n21060), .B(n21063), .Z(n2028) );
  NANDN U3969 ( .A(n21061), .B(n2028), .Z(n2029) );
  NAND U3970 ( .A(n2027), .B(n2029), .Z(n20728) );
  NAND U3971 ( .A(n21076), .B(n21079), .Z(n2030) );
  XOR U3972 ( .A(n21076), .B(n21079), .Z(n2031) );
  NANDN U3973 ( .A(n21077), .B(n2031), .Z(n2032) );
  NAND U3974 ( .A(n2030), .B(n2032), .Z(n20744) );
  NAND U3975 ( .A(n18795), .B(n18794), .Z(n2033) );
  NANDN U3976 ( .A(n18821), .B(n18820), .Z(n2034) );
  AND U3977 ( .A(n2033), .B(n2034), .Z(n18799) );
  NAND U3978 ( .A(n10078), .B(n10079), .Z(n2035) );
  NANDN U3979 ( .A(n9716), .B(n9715), .Z(n2036) );
  NAND U3980 ( .A(n2035), .B(n2036), .Z(n9717) );
  XNOR U3981 ( .A(n9367), .B(n9368), .Z(n9386) );
  XNOR U3982 ( .A(n8670), .B(n8671), .Z(n9022) );
  XNOR U3983 ( .A(n21206), .B(n21207), .Z(n21208) );
  XNOR U3984 ( .A(n21218), .B(n21219), .Z(n21527) );
  XNOR U3985 ( .A(n21228), .B(n21229), .Z(n21231) );
  XNOR U3986 ( .A(n20898), .B(n20899), .Z(n21237) );
  NAND U3987 ( .A(n21296), .B(n21299), .Z(n2037) );
  XOR U3988 ( .A(n21296), .B(n21299), .Z(n2038) );
  NANDN U3989 ( .A(n21297), .B(n2038), .Z(n2039) );
  NAND U3990 ( .A(n2037), .B(n2039), .Z(n20965) );
  NAND U3991 ( .A(n21312), .B(n21315), .Z(n2040) );
  XOR U3992 ( .A(n21312), .B(n21315), .Z(n2041) );
  NANDN U3993 ( .A(n21313), .B(n2041), .Z(n2042) );
  NAND U3994 ( .A(n2040), .B(n2042), .Z(n20980) );
  NAND U3995 ( .A(n21328), .B(n21331), .Z(n2043) );
  XOR U3996 ( .A(n21328), .B(n21331), .Z(n2044) );
  NANDN U3997 ( .A(n21329), .B(n2044), .Z(n2045) );
  NAND U3998 ( .A(n2043), .B(n2045), .Z(n20999) );
  NAND U3999 ( .A(n21344), .B(n21347), .Z(n2046) );
  XOR U4000 ( .A(n21344), .B(n21347), .Z(n2047) );
  NANDN U4001 ( .A(n21345), .B(n2047), .Z(n2048) );
  NAND U4002 ( .A(n2046), .B(n2048), .Z(n21010) );
  XOR U4003 ( .A(n21365), .B(n21362), .Z(n2049) );
  NANDN U4004 ( .A(n21363), .B(n2049), .Z(n2050) );
  NAND U4005 ( .A(n21365), .B(n21362), .Z(n2051) );
  AND U4006 ( .A(n2050), .B(n2051), .Z(n21033) );
  NAND U4007 ( .A(n21376), .B(n21379), .Z(n2052) );
  XOR U4008 ( .A(n21376), .B(n21379), .Z(n2053) );
  NANDN U4009 ( .A(n21377), .B(n2053), .Z(n2054) );
  NAND U4010 ( .A(n2052), .B(n2054), .Z(n21049) );
  NAND U4011 ( .A(n21392), .B(n21395), .Z(n2055) );
  XOR U4012 ( .A(n21392), .B(n21395), .Z(n2056) );
  NANDN U4013 ( .A(n21393), .B(n2056), .Z(n2057) );
  NAND U4014 ( .A(n2055), .B(n2057), .Z(n21065) );
  NAND U4015 ( .A(n21408), .B(n21411), .Z(n2058) );
  XOR U4016 ( .A(n21408), .B(n21411), .Z(n2059) );
  NANDN U4017 ( .A(n21409), .B(n2059), .Z(n2060) );
  NAND U4018 ( .A(n2058), .B(n2060), .Z(n21081) );
  NAND U4019 ( .A(n21424), .B(n21427), .Z(n2061) );
  XOR U4020 ( .A(n21424), .B(n21427), .Z(n2062) );
  NANDN U4021 ( .A(n21425), .B(n2062), .Z(n2063) );
  NAND U4022 ( .A(n2061), .B(n2063), .Z(n21097) );
  XOR U4023 ( .A(n20756), .B(n20757), .Z(n2064) );
  XNOR U4024 ( .A(n20755), .B(n2064), .Z(n20829) );
  XOR U4025 ( .A(n21449), .B(n21448), .Z(n2065) );
  NANDN U4026 ( .A(n21451), .B(n2065), .Z(n2066) );
  NAND U4027 ( .A(n21449), .B(n21448), .Z(n2067) );
  AND U4028 ( .A(n2066), .B(n2067), .Z(n21457) );
  NAND U4029 ( .A(n21468), .B(n21471), .Z(n2068) );
  XOR U4030 ( .A(n21468), .B(n21471), .Z(n2069) );
  NANDN U4031 ( .A(n21469), .B(n2069), .Z(n2070) );
  NAND U4032 ( .A(n2068), .B(n2070), .Z(n21133) );
  NAND U4033 ( .A(n19462), .B(n19461), .Z(n2071) );
  NANDN U4034 ( .A(n19493), .B(n19492), .Z(n2072) );
  AND U4035 ( .A(n2071), .B(n2072), .Z(n19466) );
  NAND U4036 ( .A(n19464), .B(n19463), .Z(n2073) );
  NAND U4037 ( .A(n19144), .B(n19145), .Z(n2074) );
  NAND U4038 ( .A(n2073), .B(n2074), .Z(n19468) );
  NAND U4039 ( .A(n20469), .B(n20468), .Z(n2075) );
  NAND U4040 ( .A(n20132), .B(n20131), .Z(n2076) );
  AND U4041 ( .A(n2075), .B(n2076), .Z(n20135) );
  NAND U4042 ( .A(n16444), .B(n16443), .Z(n2077) );
  NANDN U4043 ( .A(n16788), .B(n16787), .Z(n2078) );
  AND U4044 ( .A(n2077), .B(n2078), .Z(n16448) );
  NAND U4045 ( .A(n15058), .B(n15057), .Z(n2079) );
  NANDN U4046 ( .A(n15408), .B(n15407), .Z(n2080) );
  AND U4047 ( .A(n2079), .B(n2080), .Z(n15062) );
  XNOR U4048 ( .A(n9023), .B(n9024), .Z(n9378) );
  XOR U4049 ( .A(n10235), .B(n10234), .Z(n10240) );
  XNOR U4050 ( .A(n22577), .B(n22576), .Z(n22571) );
  NAND U4051 ( .A(n21628), .B(n21631), .Z(n2081) );
  XOR U4052 ( .A(n21628), .B(n21631), .Z(n2082) );
  NANDN U4053 ( .A(n21629), .B(n2082), .Z(n2083) );
  NAND U4054 ( .A(n2081), .B(n2083), .Z(n21301) );
  NAND U4055 ( .A(n21644), .B(n21647), .Z(n2084) );
  XOR U4056 ( .A(n21644), .B(n21647), .Z(n2085) );
  NANDN U4057 ( .A(n21645), .B(n2085), .Z(n2086) );
  NAND U4058 ( .A(n2084), .B(n2086), .Z(n21317) );
  XOR U4059 ( .A(n21663), .B(n21661), .Z(n2087) );
  NANDN U4060 ( .A(n21660), .B(n2087), .Z(n2088) );
  NAND U4061 ( .A(n21663), .B(n21661), .Z(n2089) );
  AND U4062 ( .A(n2088), .B(n2089), .Z(n21333) );
  NAND U4063 ( .A(n21678), .B(n21681), .Z(n2090) );
  XOR U4064 ( .A(n21678), .B(n21681), .Z(n2091) );
  NANDN U4065 ( .A(n21679), .B(n2091), .Z(n2092) );
  NAND U4066 ( .A(n2090), .B(n2092), .Z(n21349) );
  NAND U4067 ( .A(n21696), .B(n21699), .Z(n2093) );
  XOR U4068 ( .A(n21696), .B(n21699), .Z(n2094) );
  NANDN U4069 ( .A(n21697), .B(n2094), .Z(n2095) );
  NAND U4070 ( .A(n2093), .B(n2095), .Z(n21361) );
  NAND U4071 ( .A(n21712), .B(n21715), .Z(n2096) );
  XOR U4072 ( .A(n21712), .B(n21715), .Z(n2097) );
  NANDN U4073 ( .A(n21713), .B(n2097), .Z(n2098) );
  NAND U4074 ( .A(n2096), .B(n2098), .Z(n21381) );
  NAND U4075 ( .A(n21728), .B(n21731), .Z(n2099) );
  XOR U4076 ( .A(n21728), .B(n21731), .Z(n2100) );
  NANDN U4077 ( .A(n21729), .B(n2100), .Z(n2101) );
  NAND U4078 ( .A(n2099), .B(n2101), .Z(n21397) );
  XOR U4079 ( .A(n21747), .B(n21744), .Z(n2102) );
  NANDN U4080 ( .A(n21745), .B(n2102), .Z(n2103) );
  NAND U4081 ( .A(n21747), .B(n21744), .Z(n2104) );
  AND U4082 ( .A(n2103), .B(n2104), .Z(n21413) );
  XOR U4083 ( .A(n21763), .B(n21761), .Z(n2105) );
  NANDN U4084 ( .A(n21760), .B(n2105), .Z(n2106) );
  NAND U4085 ( .A(n21763), .B(n21761), .Z(n2107) );
  AND U4086 ( .A(n2106), .B(n2107), .Z(n21429) );
  XOR U4087 ( .A(n22127), .B(n22125), .Z(n2108) );
  NANDN U4088 ( .A(n22124), .B(n2108), .Z(n2109) );
  NAND U4089 ( .A(n22127), .B(n22125), .Z(n2110) );
  AND U4090 ( .A(n2109), .B(n2110), .Z(n21777) );
  NAND U4091 ( .A(n21778), .B(n21781), .Z(n2111) );
  XOR U4092 ( .A(n21778), .B(n21781), .Z(n2112) );
  NANDN U4093 ( .A(n21779), .B(n2112), .Z(n2113) );
  NAND U4094 ( .A(n2111), .B(n2113), .Z(n21784) );
  XNOR U4095 ( .A(n21466), .B(n21467), .Z(n21811) );
  NAND U4096 ( .A(n21139), .B(n21141), .Z(n2114) );
  XOR U4097 ( .A(n21139), .B(n21141), .Z(n2115) );
  NANDN U4098 ( .A(n21138), .B(n2115), .Z(n2116) );
  NAND U4099 ( .A(n2114), .B(n2116), .Z(n20819) );
  NAND U4100 ( .A(n17132), .B(n17131), .Z(n2117) );
  NANDN U4101 ( .A(n17480), .B(n17479), .Z(n2118) );
  AND U4102 ( .A(n2117), .B(n2118), .Z(n17136) );
  NAND U4103 ( .A(n14710), .B(n14709), .Z(n2119) );
  NAND U4104 ( .A(n14365), .B(n14364), .Z(n2120) );
  AND U4105 ( .A(n2119), .B(n2120), .Z(n14369) );
  NAND U4106 ( .A(n13648), .B(n13647), .Z(n2121) );
  NANDN U4107 ( .A(n13331), .B(n13332), .Z(n2122) );
  AND U4108 ( .A(n2121), .B(n2122), .Z(n13655) );
  NAND U4109 ( .A(n13646), .B(n13645), .Z(n2123) );
  NANDN U4110 ( .A(n14035), .B(n14034), .Z(n2124) );
  AND U4111 ( .A(n2123), .B(n2124), .Z(n13650) );
  NAND U4112 ( .A(n23109), .B(n23108), .Z(n2125) );
  NANDN U4113 ( .A(n23111), .B(n23110), .Z(n2126) );
  NAND U4114 ( .A(n2125), .B(n2126), .Z(n23124) );
  NAND U4115 ( .A(n23130), .B(n23129), .Z(n2127) );
  NAND U4116 ( .A(n23128), .B(n23127), .Z(n2128) );
  NAND U4117 ( .A(n2127), .B(n2128), .Z(n23361) );
  XNOR U4118 ( .A(n21558), .B(n21559), .Z(n21560) );
  XOR U4119 ( .A(n21955), .B(n21953), .Z(n2129) );
  NANDN U4120 ( .A(n21952), .B(n2129), .Z(n2130) );
  NAND U4121 ( .A(n21955), .B(n21953), .Z(n2131) );
  AND U4122 ( .A(n2130), .B(n2131), .Z(n21627) );
  XOR U4123 ( .A(n21971), .B(n21969), .Z(n2132) );
  NANDN U4124 ( .A(n21968), .B(n2132), .Z(n2133) );
  NAND U4125 ( .A(n21971), .B(n21969), .Z(n2134) );
  AND U4126 ( .A(n2133), .B(n2134), .Z(n21643) );
  XOR U4127 ( .A(n21991), .B(n21989), .Z(n2135) );
  NANDN U4128 ( .A(n21988), .B(n2135), .Z(n2136) );
  NAND U4129 ( .A(n21991), .B(n21989), .Z(n2137) );
  AND U4130 ( .A(n2136), .B(n2137), .Z(n21658) );
  XOR U4131 ( .A(n22011), .B(n22009), .Z(n2138) );
  NANDN U4132 ( .A(n22008), .B(n2138), .Z(n2139) );
  NAND U4133 ( .A(n22011), .B(n22009), .Z(n2140) );
  AND U4134 ( .A(n2139), .B(n2140), .Z(n21677) );
  NAND U4135 ( .A(n22029), .B(n22031), .Z(n2141) );
  XOR U4136 ( .A(n22029), .B(n22031), .Z(n2142) );
  NANDN U4137 ( .A(n22028), .B(n2142), .Z(n2143) );
  NAND U4138 ( .A(n2141), .B(n2143), .Z(n21695) );
  XOR U4139 ( .A(n22047), .B(n22045), .Z(n2144) );
  NANDN U4140 ( .A(n22044), .B(n2144), .Z(n2145) );
  NAND U4141 ( .A(n22047), .B(n22045), .Z(n2146) );
  AND U4142 ( .A(n2145), .B(n2146), .Z(n21711) );
  XOR U4143 ( .A(n22067), .B(n22065), .Z(n2147) );
  NANDN U4144 ( .A(n22064), .B(n2147), .Z(n2148) );
  NAND U4145 ( .A(n22067), .B(n22065), .Z(n2149) );
  AND U4146 ( .A(n2148), .B(n2149), .Z(n21727) );
  XOR U4147 ( .A(n22087), .B(n22085), .Z(n2150) );
  NANDN U4148 ( .A(n22084), .B(n2150), .Z(n2151) );
  NAND U4149 ( .A(n22087), .B(n22085), .Z(n2152) );
  AND U4150 ( .A(n2151), .B(n2152), .Z(n21743) );
  XOR U4151 ( .A(n22107), .B(n22105), .Z(n2153) );
  NANDN U4152 ( .A(n22104), .B(n2153), .Z(n2154) );
  NAND U4153 ( .A(n22107), .B(n22105), .Z(n2155) );
  AND U4154 ( .A(n2154), .B(n2155), .Z(n21758) );
  XOR U4155 ( .A(n21805), .B(n21806), .Z(n2156) );
  XNOR U4156 ( .A(n21804), .B(n2156), .Z(n21835) );
  XNOR U4157 ( .A(n21816), .B(n21817), .Z(n22152) );
  XOR U4158 ( .A(n18171), .B(n18168), .Z(n2157) );
  NAND U4159 ( .A(n2157), .B(n18169), .Z(n2158) );
  NAND U4160 ( .A(n18171), .B(n18168), .Z(n2159) );
  AND U4161 ( .A(n2158), .B(n2159), .Z(n18151) );
  NAND U4162 ( .A(n18805), .B(n18804), .Z(n2160) );
  NAND U4163 ( .A(n18483), .B(n18484), .Z(n2161) );
  NAND U4164 ( .A(n2160), .B(n2161), .Z(n18811) );
  NAND U4165 ( .A(n15756), .B(n15755), .Z(n2162) );
  NANDN U4166 ( .A(n16108), .B(n16107), .Z(n2163) );
  AND U4167 ( .A(n2162), .B(n2163), .Z(n15760) );
  XOR U4168 ( .A(n9733), .B(n9734), .Z(n10097) );
  XOR U4169 ( .A(n21844), .B(n21845), .Z(n21879) );
  XOR U4170 ( .A(n22263), .B(n22264), .Z(n2164) );
  NANDN U4171 ( .A(n22266), .B(n2164), .Z(n2165) );
  NAND U4172 ( .A(n22263), .B(n22264), .Z(n2166) );
  AND U4173 ( .A(n2165), .B(n2166), .Z(n21949) );
  XOR U4174 ( .A(n22303), .B(n22304), .Z(n2167) );
  NANDN U4175 ( .A(n22306), .B(n2167), .Z(n2168) );
  NAND U4176 ( .A(n22303), .B(n22304), .Z(n2169) );
  AND U4177 ( .A(n2168), .B(n2169), .Z(n21985) );
  XOR U4178 ( .A(n22326), .B(n22323), .Z(n2170) );
  NAND U4179 ( .A(n2170), .B(n22324), .Z(n2171) );
  NAND U4180 ( .A(n22326), .B(n22323), .Z(n2172) );
  AND U4181 ( .A(n2171), .B(n2172), .Z(n22005) );
  XOR U4182 ( .A(n22343), .B(n22344), .Z(n2173) );
  NANDN U4183 ( .A(n22346), .B(n2173), .Z(n2174) );
  NAND U4184 ( .A(n22343), .B(n22344), .Z(n2175) );
  AND U4185 ( .A(n2174), .B(n2175), .Z(n22025) );
  XOR U4186 ( .A(n22383), .B(n22384), .Z(n2176) );
  NANDN U4187 ( .A(n22386), .B(n2176), .Z(n2177) );
  NAND U4188 ( .A(n22383), .B(n22384), .Z(n2178) );
  AND U4189 ( .A(n2177), .B(n2178), .Z(n22061) );
  XOR U4190 ( .A(n22403), .B(n22404), .Z(n2179) );
  NANDN U4191 ( .A(n22406), .B(n2179), .Z(n2180) );
  NAND U4192 ( .A(n22403), .B(n22404), .Z(n2181) );
  AND U4193 ( .A(n2180), .B(n2181), .Z(n22081) );
  XOR U4194 ( .A(n22423), .B(n22424), .Z(n2182) );
  NANDN U4195 ( .A(n22426), .B(n2182), .Z(n2183) );
  NAND U4196 ( .A(n22423), .B(n22424), .Z(n2184) );
  AND U4197 ( .A(n2183), .B(n2184), .Z(n22101) );
  XOR U4198 ( .A(n22446), .B(n22443), .Z(n2185) );
  NAND U4199 ( .A(n2185), .B(n22444), .Z(n2186) );
  NAND U4200 ( .A(n22446), .B(n22443), .Z(n2187) );
  AND U4201 ( .A(n2186), .B(n2187), .Z(n22121) );
  NAND U4202 ( .A(n19475), .B(n19476), .Z(n2188) );
  NAND U4203 ( .A(n19150), .B(n19151), .Z(n2189) );
  NAND U4204 ( .A(n2188), .B(n2189), .Z(n19155) );
  NAND U4205 ( .A(n19485), .B(n19484), .Z(n2190) );
  NAND U4206 ( .A(n19473), .B(n19474), .Z(n2191) );
  AND U4207 ( .A(n2190), .B(n2191), .Z(n19477) );
  NAND U4208 ( .A(n20144), .B(n20143), .Z(n2192) );
  NANDN U4209 ( .A(n20477), .B(n20476), .Z(n2193) );
  AND U4210 ( .A(n2192), .B(n2193), .Z(n20479) );
  OR U4211 ( .A(n14731), .B(n14730), .Z(n2194) );
  NAND U4212 ( .A(n14719), .B(n14720), .Z(n2195) );
  AND U4213 ( .A(n2194), .B(n2195), .Z(n14729) );
  XNOR U4214 ( .A(n10100), .B(n10101), .Z(n10103) );
  XOR U4215 ( .A(n10253), .B(n10252), .Z(n10258) );
  NAND U4216 ( .A(n22859), .B(n22858), .Z(n2196) );
  NANDN U4217 ( .A(n22861), .B(n22860), .Z(n2197) );
  NAND U4218 ( .A(n2196), .B(n2197), .Z(n22992) );
  XNOR U4219 ( .A(n21890), .B(n21891), .Z(n22166) );
  XNOR U4220 ( .A(n21894), .B(n21895), .Z(n22220) );
  XOR U4221 ( .A(n24814), .B(n24811), .Z(n2198) );
  NANDN U4222 ( .A(n24812), .B(n2198), .Z(n2199) );
  NAND U4223 ( .A(n24814), .B(n24811), .Z(n2200) );
  AND U4224 ( .A(n2199), .B(n2200), .Z(n22261) );
  NAND U4225 ( .A(n24826), .B(n24828), .Z(n2201) );
  XOR U4226 ( .A(n24826), .B(n24828), .Z(n2202) );
  NANDN U4227 ( .A(n24825), .B(n2202), .Z(n2203) );
  NAND U4228 ( .A(n2201), .B(n2203), .Z(n22282) );
  NAND U4229 ( .A(n21967), .B(n21966), .Z(n2204) );
  NANDN U4230 ( .A(n22289), .B(n22290), .Z(n2205) );
  NAND U4231 ( .A(n2204), .B(n2205), .Z(n22294) );
  XOR U4232 ( .A(n24838), .B(n24837), .Z(n2206) );
  NANDN U4233 ( .A(n24840), .B(n2206), .Z(n2207) );
  NAND U4234 ( .A(n24838), .B(n24837), .Z(n2208) );
  AND U4235 ( .A(n2207), .B(n2208), .Z(n22301) );
  NAND U4236 ( .A(n24850), .B(n24852), .Z(n2209) );
  XOR U4237 ( .A(n24850), .B(n24852), .Z(n2210) );
  NANDN U4238 ( .A(n24849), .B(n2210), .Z(n2211) );
  NAND U4239 ( .A(n2209), .B(n2211), .Z(n22322) );
  NAND U4240 ( .A(n24864), .B(n24866), .Z(n2212) );
  XOR U4241 ( .A(n24864), .B(n24866), .Z(n2213) );
  NANDN U4242 ( .A(n24863), .B(n2213), .Z(n2214) );
  NAND U4243 ( .A(n2212), .B(n2214), .Z(n22342) );
  NAND U4244 ( .A(n24876), .B(n24878), .Z(n2215) );
  XOR U4245 ( .A(n24876), .B(n24878), .Z(n2216) );
  NANDN U4246 ( .A(n24875), .B(n2216), .Z(n2217) );
  NAND U4247 ( .A(n2215), .B(n2217), .Z(n22362) );
  NAND U4248 ( .A(n22043), .B(n22042), .Z(n2218) );
  NANDN U4249 ( .A(n22369), .B(n22370), .Z(n2219) );
  NAND U4250 ( .A(n2218), .B(n2219), .Z(n22374) );
  NAND U4251 ( .A(n24890), .B(n24892), .Z(n2220) );
  XOR U4252 ( .A(n24890), .B(n24892), .Z(n2221) );
  NANDN U4253 ( .A(n24889), .B(n2221), .Z(n2222) );
  NAND U4254 ( .A(n2220), .B(n2222), .Z(n22382) );
  NAND U4255 ( .A(n24902), .B(n24904), .Z(n2223) );
  XOR U4256 ( .A(n24902), .B(n24904), .Z(n2224) );
  NANDN U4257 ( .A(n24901), .B(n2224), .Z(n2225) );
  NAND U4258 ( .A(n2223), .B(n2225), .Z(n22402) );
  NAND U4259 ( .A(n24914), .B(n24916), .Z(n2226) );
  XOR U4260 ( .A(n24914), .B(n24916), .Z(n2227) );
  NANDN U4261 ( .A(n24913), .B(n2227), .Z(n2228) );
  NAND U4262 ( .A(n2226), .B(n2228), .Z(n22422) );
  NAND U4263 ( .A(n24928), .B(n24930), .Z(n2229) );
  XOR U4264 ( .A(n24928), .B(n24930), .Z(n2230) );
  NANDN U4265 ( .A(n24927), .B(n2230), .Z(n2231) );
  NAND U4266 ( .A(n2229), .B(n2231), .Z(n22442) );
  XOR U4267 ( .A(n24942), .B(n24939), .Z(n2232) );
  NANDN U4268 ( .A(n24940), .B(n2232), .Z(n2233) );
  NAND U4269 ( .A(n24942), .B(n24939), .Z(n2234) );
  AND U4270 ( .A(n2233), .B(n2234), .Z(n22465) );
  XOR U4271 ( .A(n22472), .B(n22469), .Z(n2235) );
  NANDN U4272 ( .A(n22470), .B(n2235), .Z(n2236) );
  NAND U4273 ( .A(n22472), .B(n22469), .Z(n2237) );
  AND U4274 ( .A(n2236), .B(n2237), .Z(n22476) );
  NAND U4275 ( .A(n24956), .B(n24953), .Z(n2238) );
  XOR U4276 ( .A(n24956), .B(n24953), .Z(n2239) );
  NANDN U4277 ( .A(n24954), .B(n2239), .Z(n2240) );
  NAND U4278 ( .A(n2238), .B(n2240), .Z(n22482) );
  NAND U4279 ( .A(n22484), .B(n22486), .Z(n2241) );
  XOR U4280 ( .A(n22484), .B(n22486), .Z(n2242) );
  NANDN U4281 ( .A(n22483), .B(n2242), .Z(n2243) );
  NAND U4282 ( .A(n2241), .B(n2243), .Z(n22160) );
  NAND U4283 ( .A(n20815), .B(n20814), .Z(n2244) );
  NAND U4284 ( .A(n20474), .B(n20475), .Z(n2245) );
  NAND U4285 ( .A(n2244), .B(n2245), .Z(n20483) );
  ANDN U4286 ( .B(n16804), .A(n16803), .Z(n16462) );
  NAND U4287 ( .A(n14724), .B(n14723), .Z(n2246) );
  NAND U4288 ( .A(n14376), .B(n14377), .Z(n2247) );
  NAND U4289 ( .A(n2246), .B(n2247), .Z(n14725) );
  XOR U4290 ( .A(n22703), .B(n22702), .Z(n22554) );
  XNOR U4291 ( .A(n22217), .B(n22218), .Z(n24970) );
  NANDN U4292 ( .A(n24668), .B(n24667), .Z(n2248) );
  NAND U4293 ( .A(n24670), .B(n2248), .Z(n2249) );
  NANDN U4294 ( .A(n24672), .B(n2249), .Z(n2250) );
  XOR U4295 ( .A(n24673), .B(n24674), .Z(n2251) );
  NAND U4296 ( .A(n2251), .B(n2250), .Z(n2252) );
  NAND U4297 ( .A(n24673), .B(n24674), .Z(n2253) );
  AND U4298 ( .A(n2252), .B(n2253), .Z(n24680) );
  NANDN U4299 ( .A(n19481), .B(n24702), .Z(n2254) );
  AND U4300 ( .A(n24703), .B(n2254), .Z(n2255) );
  AND U4301 ( .A(n24710), .B(n24713), .Z(n2256) );
  ANDN U4302 ( .B(n24706), .A(n24705), .Z(n2257) );
  NAND U4303 ( .A(n24704), .B(n2255), .Z(n2258) );
  NAND U4304 ( .A(n2256), .B(n2258), .Z(n2259) );
  NANDN U4305 ( .A(n2257), .B(n2259), .Z(n2260) );
  XOR U4306 ( .A(n24715), .B(n24716), .Z(n2261) );
  NAND U4307 ( .A(n2261), .B(n2260), .Z(n2262) );
  NAND U4308 ( .A(n24715), .B(n24716), .Z(n2263) );
  AND U4309 ( .A(n2262), .B(n2263), .Z(n24719) );
  ANDN U4310 ( .B(n18163), .A(n18162), .Z(n24722) );
  NAND U4311 ( .A(n24728), .B(n24727), .Z(n2264) );
  NAND U4312 ( .A(n17151), .B(n17152), .Z(n2265) );
  AND U4313 ( .A(n2264), .B(n2265), .Z(n24730) );
  NAND U4314 ( .A(n24760), .B(n24759), .Z(n2266) );
  XOR U4315 ( .A(n24760), .B(n24759), .Z(n2267) );
  NANDN U4316 ( .A(n24762), .B(n2267), .Z(n2268) );
  NAND U4317 ( .A(n2266), .B(n2268), .Z(n24763) );
  NAND U4318 ( .A(n24768), .B(n24767), .Z(n24772) );
  NAND U4319 ( .A(n24790), .B(n24789), .Z(n2269) );
  NAND U4320 ( .A(n10980), .B(n10981), .Z(n2270) );
  AND U4321 ( .A(n2269), .B(n2270), .Z(n24792) );
  XOR U4322 ( .A(n22849), .B(n22851), .Z(n2271) );
  NAND U4323 ( .A(n2271), .B(n22850), .Z(n2272) );
  NAND U4324 ( .A(n22849), .B(n22851), .Z(n2273) );
  AND U4325 ( .A(n2272), .B(n2273), .Z(n22988) );
  NANDN U4326 ( .A(n23710), .B(n23709), .Z(n2274) );
  AND U4327 ( .A(n23711), .B(n2274), .Z(n2275) );
  AND U4328 ( .A(n23707), .B(n23708), .Z(n2276) );
  OR U4329 ( .A(n23706), .B(n23705), .Z(n2277) );
  NANDN U4330 ( .A(n2275), .B(n2276), .Z(n2278) );
  NAND U4331 ( .A(n2277), .B(n2278), .Z(n2279) );
  AND U4332 ( .A(n23716), .B(n2276), .Z(n2280) );
  NANDN U4333 ( .A(n23715), .B(n23714), .Z(n2281) );
  AND U4334 ( .A(n2280), .B(n2281), .Z(n2282) );
  NOR U4335 ( .A(n2282), .B(n2279), .Z(n2283) );
  OR U4336 ( .A(n23713), .B(n23712), .Z(n2284) );
  NAND U4337 ( .A(n2283), .B(n2284), .Z(n2285) );
  NANDN U4338 ( .A(n23704), .B(n23712), .Z(n2286) );
  AND U4339 ( .A(n2285), .B(n2286), .Z(n23817) );
  NAND U4340 ( .A(n23918), .B(n23917), .Z(n2287) );
  NAND U4341 ( .A(n23915), .B(n23916), .Z(n2288) );
  AND U4342 ( .A(n2287), .B(n2288), .Z(n24088) );
  NAND U4343 ( .A(n24655), .B(n24656), .Z(n2289) );
  NANDN U4344 ( .A(n24658), .B(n24657), .Z(n2290) );
  AND U4345 ( .A(n2289), .B(n2290), .Z(n2291) );
  NAND U4346 ( .A(a[63]), .B(n24654), .Z(n2292) );
  XNOR U4347 ( .A(n2291), .B(n2292), .Z(c[127]) );
  AND U4348 ( .A(a[62]), .B(b[38]), .Z(n10253) );
  AND U4349 ( .A(a[41]), .B(b[59]), .Z(n10148) );
  AND U4350 ( .A(a[40]), .B(b[59]), .Z(n3083) );
  AND U4351 ( .A(a[37]), .B(b[59]), .Z(n3017) );
  AND U4352 ( .A(a[34]), .B(b[59]), .Z(n2951) );
  NAND U4353 ( .A(a[32]), .B(b[59]), .Z(n2907) );
  AND U4354 ( .A(a[31]), .B(b[59]), .Z(n2886) );
  AND U4355 ( .A(b[63]), .B(a[14]), .Z(n2434) );
  AND U4356 ( .A(b[62]), .B(a[15]), .Z(n2432) );
  AND U4357 ( .A(b[63]), .B(a[13]), .Z(n2339) );
  AND U4358 ( .A(b[63]), .B(a[12]), .Z(n2335) );
  AND U4359 ( .A(b[63]), .B(a[11]), .Z(n2331) );
  AND U4360 ( .A(b[63]), .B(a[10]), .Z(n2327) );
  AND U4361 ( .A(b[63]), .B(a[9]), .Z(n2323) );
  AND U4362 ( .A(b[63]), .B(a[8]), .Z(n2319) );
  AND U4363 ( .A(b[63]), .B(a[7]), .Z(n2315) );
  AND U4364 ( .A(b[63]), .B(a[6]), .Z(n2311) );
  AND U4365 ( .A(b[63]), .B(a[5]), .Z(n2307) );
  AND U4366 ( .A(b[63]), .B(a[4]), .Z(n2303) );
  AND U4367 ( .A(b[63]), .B(a[3]), .Z(n2299) );
  NAND U4368 ( .A(b[62]), .B(a[2]), .Z(n2372) );
  AND U4369 ( .A(b[63]), .B(a[1]), .Z(n2374) );
  NANDN U4370 ( .A(n2372), .B(n2374), .Z(n2297) );
  NAND U4371 ( .A(b[62]), .B(a[0]), .Z(n2373) );
  NANDN U4372 ( .A(n2373), .B(a[1]), .Z(n2293) );
  NANDN U4373 ( .A(a[2]), .B(n2293), .Z(n2294) );
  AND U4374 ( .A(b[63]), .B(n2294), .Z(n2295) );
  AND U4375 ( .A(n2297), .B(n2295), .Z(n2365) );
  AND U4376 ( .A(b[62]), .B(a[3]), .Z(n2364) );
  NAND U4377 ( .A(n2365), .B(n2364), .Z(n2296) );
  AND U4378 ( .A(n2297), .B(n2296), .Z(n2298) );
  NANDN U4379 ( .A(n2299), .B(n2298), .Z(n2301) );
  XOR U4380 ( .A(n2299), .B(n2298), .Z(n2362) );
  AND U4381 ( .A(b[62]), .B(a[4]), .Z(n2363) );
  OR U4382 ( .A(n2362), .B(n2363), .Z(n2300) );
  NAND U4383 ( .A(n2301), .B(n2300), .Z(n2302) );
  NANDN U4384 ( .A(n2303), .B(n2302), .Z(n2305) );
  AND U4385 ( .A(b[62]), .B(a[5]), .Z(n2361) );
  XNOR U4386 ( .A(n2303), .B(n2302), .Z(n2360) );
  NANDN U4387 ( .A(n2361), .B(n2360), .Z(n2304) );
  NAND U4388 ( .A(n2305), .B(n2304), .Z(n2306) );
  NANDN U4389 ( .A(n2307), .B(n2306), .Z(n2309) );
  XOR U4390 ( .A(n2307), .B(n2306), .Z(n2358) );
  AND U4391 ( .A(b[62]), .B(a[6]), .Z(n2359) );
  OR U4392 ( .A(n2358), .B(n2359), .Z(n2308) );
  NAND U4393 ( .A(n2309), .B(n2308), .Z(n2310) );
  NANDN U4394 ( .A(n2311), .B(n2310), .Z(n2313) );
  XOR U4395 ( .A(n2311), .B(n2310), .Z(n2356) );
  AND U4396 ( .A(b[62]), .B(a[7]), .Z(n2357) );
  OR U4397 ( .A(n2356), .B(n2357), .Z(n2312) );
  NAND U4398 ( .A(n2313), .B(n2312), .Z(n2314) );
  NANDN U4399 ( .A(n2315), .B(n2314), .Z(n2317) );
  XOR U4400 ( .A(n2315), .B(n2314), .Z(n2354) );
  AND U4401 ( .A(b[62]), .B(a[8]), .Z(n2355) );
  OR U4402 ( .A(n2354), .B(n2355), .Z(n2316) );
  NAND U4403 ( .A(n2317), .B(n2316), .Z(n2318) );
  NANDN U4404 ( .A(n2319), .B(n2318), .Z(n2321) );
  XOR U4405 ( .A(n2319), .B(n2318), .Z(n2352) );
  AND U4406 ( .A(b[62]), .B(a[9]), .Z(n2353) );
  OR U4407 ( .A(n2352), .B(n2353), .Z(n2320) );
  NAND U4408 ( .A(n2321), .B(n2320), .Z(n2322) );
  NANDN U4409 ( .A(n2323), .B(n2322), .Z(n2325) );
  XOR U4410 ( .A(n2323), .B(n2322), .Z(n2350) );
  AND U4411 ( .A(b[62]), .B(a[10]), .Z(n2351) );
  OR U4412 ( .A(n2350), .B(n2351), .Z(n2324) );
  NAND U4413 ( .A(n2325), .B(n2324), .Z(n2326) );
  NANDN U4414 ( .A(n2327), .B(n2326), .Z(n2329) );
  AND U4415 ( .A(b[62]), .B(a[11]), .Z(n2349) );
  XNOR U4416 ( .A(n2327), .B(n2326), .Z(n2348) );
  NANDN U4417 ( .A(n2349), .B(n2348), .Z(n2328) );
  NAND U4418 ( .A(n2329), .B(n2328), .Z(n2330) );
  NANDN U4419 ( .A(n2331), .B(n2330), .Z(n2333) );
  AND U4420 ( .A(b[62]), .B(a[12]), .Z(n2347) );
  XNOR U4421 ( .A(n2331), .B(n2330), .Z(n2346) );
  NANDN U4422 ( .A(n2347), .B(n2346), .Z(n2332) );
  NAND U4423 ( .A(n2333), .B(n2332), .Z(n2334) );
  NANDN U4424 ( .A(n2335), .B(n2334), .Z(n2337) );
  AND U4425 ( .A(b[62]), .B(a[13]), .Z(n2345) );
  XNOR U4426 ( .A(n2335), .B(n2334), .Z(n2344) );
  NANDN U4427 ( .A(n2345), .B(n2344), .Z(n2336) );
  NAND U4428 ( .A(n2337), .B(n2336), .Z(n2338) );
  NANDN U4429 ( .A(n2339), .B(n2338), .Z(n2341) );
  AND U4430 ( .A(b[62]), .B(a[14]), .Z(n2343) );
  XNOR U4431 ( .A(n2339), .B(n2338), .Z(n2342) );
  NANDN U4432 ( .A(n2343), .B(n2342), .Z(n2340) );
  NAND U4433 ( .A(n2341), .B(n2340), .Z(n2431) );
  XNOR U4434 ( .A(n2432), .B(n2431), .Z(n2433) );
  XOR U4435 ( .A(n2434), .B(n2433), .Z(n2428) );
  XOR U4436 ( .A(n2343), .B(n2342), .Z(n2424) );
  XOR U4437 ( .A(n2345), .B(n2344), .Z(n2420) );
  XOR U4438 ( .A(n2347), .B(n2346), .Z(n2416) );
  XOR U4439 ( .A(n2349), .B(n2348), .Z(n2412) );
  XOR U4440 ( .A(n2351), .B(n2350), .Z(n2408) );
  XOR U4441 ( .A(n2353), .B(n2352), .Z(n2404) );
  XOR U4442 ( .A(n2355), .B(n2354), .Z(n2400) );
  XOR U4443 ( .A(n2357), .B(n2356), .Z(n2396) );
  XOR U4444 ( .A(n2359), .B(n2358), .Z(n2392) );
  XOR U4445 ( .A(n2361), .B(n2360), .Z(n2387) );
  XOR U4446 ( .A(n2363), .B(n2362), .Z(n2384) );
  XOR U4447 ( .A(n2365), .B(n2364), .Z(n2380) );
  AND U4448 ( .A(a[2]), .B(b[61]), .Z(n2470) );
  AND U4449 ( .A(b[63]), .B(a[0]), .Z(n2367) );
  NAND U4450 ( .A(a[0]), .B(b[61]), .Z(n2368) );
  IV U4451 ( .A(n2368), .Z(n2581) );
  AND U4452 ( .A(b[62]), .B(a[1]), .Z(n2369) );
  NANDN U4453 ( .A(n2581), .B(n2369), .Z(n2366) );
  XNOR U4454 ( .A(n2367), .B(n2366), .Z(n2469) );
  NAND U4455 ( .A(n2470), .B(n2469), .Z(n2371) );
  ANDN U4456 ( .B(n2369), .A(n2368), .Z(n2471) );
  NANDN U4457 ( .A(b[63]), .B(n2471), .Z(n2370) );
  AND U4458 ( .A(n2371), .B(n2370), .Z(n2375) );
  IV U4459 ( .A(n2373), .Z(n2473) );
  NAND U4460 ( .A(n2375), .B(n2376), .Z(n2378) );
  AND U4461 ( .A(a[3]), .B(b[61]), .Z(n2483) );
  XOR U4462 ( .A(n2376), .B(n2375), .Z(n2484) );
  NANDN U4463 ( .A(n2483), .B(n2484), .Z(n2377) );
  NAND U4464 ( .A(n2378), .B(n2377), .Z(n2379) );
  NANDN U4465 ( .A(n2380), .B(n2379), .Z(n2382) );
  XOR U4466 ( .A(n2380), .B(n2379), .Z(n2467) );
  AND U4467 ( .A(a[4]), .B(b[61]), .Z(n2468) );
  OR U4468 ( .A(n2467), .B(n2468), .Z(n2381) );
  AND U4469 ( .A(n2382), .B(n2381), .Z(n2383) );
  NANDN U4470 ( .A(n2384), .B(n2383), .Z(n2386) );
  NAND U4471 ( .A(a[5]), .B(b[61]), .Z(n2493) );
  XNOR U4472 ( .A(n2384), .B(n2383), .Z(n2494) );
  NANDN U4473 ( .A(n2493), .B(n2494), .Z(n2385) );
  AND U4474 ( .A(n2386), .B(n2385), .Z(n2388) );
  NANDN U4475 ( .A(n2387), .B(n2388), .Z(n2390) );
  AND U4476 ( .A(a[6]), .B(b[61]), .Z(n2500) );
  XNOR U4477 ( .A(n2388), .B(n2387), .Z(n2499) );
  NANDN U4478 ( .A(n2500), .B(n2499), .Z(n2389) );
  AND U4479 ( .A(n2390), .B(n2389), .Z(n2391) );
  NANDN U4480 ( .A(n2392), .B(n2391), .Z(n2394) );
  XNOR U4481 ( .A(n2392), .B(n2391), .Z(n2466) );
  AND U4482 ( .A(a[7]), .B(b[61]), .Z(n2465) );
  NAND U4483 ( .A(n2466), .B(n2465), .Z(n2393) );
  NAND U4484 ( .A(n2394), .B(n2393), .Z(n2395) );
  NANDN U4485 ( .A(n2396), .B(n2395), .Z(n2398) );
  XNOR U4486 ( .A(n2396), .B(n2395), .Z(n2464) );
  AND U4487 ( .A(a[8]), .B(b[61]), .Z(n2463) );
  NAND U4488 ( .A(n2464), .B(n2463), .Z(n2397) );
  NAND U4489 ( .A(n2398), .B(n2397), .Z(n2399) );
  NANDN U4490 ( .A(n2400), .B(n2399), .Z(n2402) );
  XNOR U4491 ( .A(n2400), .B(n2399), .Z(n2462) );
  AND U4492 ( .A(a[9]), .B(b[61]), .Z(n2461) );
  NAND U4493 ( .A(n2462), .B(n2461), .Z(n2401) );
  NAND U4494 ( .A(n2402), .B(n2401), .Z(n2403) );
  NANDN U4495 ( .A(n2404), .B(n2403), .Z(n2406) );
  XNOR U4496 ( .A(n2404), .B(n2403), .Z(n2518) );
  AND U4497 ( .A(a[10]), .B(b[61]), .Z(n2517) );
  NAND U4498 ( .A(n2518), .B(n2517), .Z(n2405) );
  NAND U4499 ( .A(n2406), .B(n2405), .Z(n2407) );
  NANDN U4500 ( .A(n2408), .B(n2407), .Z(n2410) );
  XNOR U4501 ( .A(n2408), .B(n2407), .Z(n2460) );
  AND U4502 ( .A(a[11]), .B(b[61]), .Z(n2459) );
  NAND U4503 ( .A(n2460), .B(n2459), .Z(n2409) );
  NAND U4504 ( .A(n2410), .B(n2409), .Z(n2411) );
  NAND U4505 ( .A(n2412), .B(n2411), .Z(n2414) );
  XOR U4506 ( .A(n2412), .B(n2411), .Z(n2458) );
  AND U4507 ( .A(a[12]), .B(b[61]), .Z(n2457) );
  NAND U4508 ( .A(n2458), .B(n2457), .Z(n2413) );
  NAND U4509 ( .A(n2414), .B(n2413), .Z(n2415) );
  NAND U4510 ( .A(n2416), .B(n2415), .Z(n2418) );
  XOR U4511 ( .A(n2416), .B(n2415), .Z(n2456) );
  AND U4512 ( .A(a[13]), .B(b[61]), .Z(n2455) );
  NAND U4513 ( .A(n2456), .B(n2455), .Z(n2417) );
  NAND U4514 ( .A(n2418), .B(n2417), .Z(n2419) );
  NAND U4515 ( .A(n2420), .B(n2419), .Z(n2422) );
  XOR U4516 ( .A(n2420), .B(n2419), .Z(n2454) );
  AND U4517 ( .A(a[14]), .B(b[61]), .Z(n2453) );
  NAND U4518 ( .A(n2454), .B(n2453), .Z(n2421) );
  NAND U4519 ( .A(n2422), .B(n2421), .Z(n2423) );
  NAND U4520 ( .A(n2424), .B(n2423), .Z(n2426) );
  NAND U4521 ( .A(a[15]), .B(b[61]), .Z(n2449) );
  XOR U4522 ( .A(n2424), .B(n2423), .Z(n2450) );
  NANDN U4523 ( .A(n2449), .B(n2450), .Z(n2425) );
  NAND U4524 ( .A(n2426), .B(n2425), .Z(n2427) );
  NAND U4525 ( .A(n2428), .B(n2427), .Z(n2430) );
  NAND U4526 ( .A(a[16]), .B(b[61]), .Z(n2543) );
  XOR U4527 ( .A(n2428), .B(n2427), .Z(n2544) );
  NANDN U4528 ( .A(n2543), .B(n2544), .Z(n2429) );
  AND U4529 ( .A(n2430), .B(n2429), .Z(n2438) );
  AND U4530 ( .A(a[17]), .B(b[61]), .Z(n2437) );
  NANDN U4531 ( .A(n2438), .B(n2437), .Z(n2440) );
  AND U4532 ( .A(b[62]), .B(a[16]), .Z(n2441) );
  NAND U4533 ( .A(b[63]), .B(a[15]), .Z(n2442) );
  XNOR U4534 ( .A(n2441), .B(n2442), .Z(n2443) );
  NANDN U4535 ( .A(n2432), .B(n2431), .Z(n2436) );
  NANDN U4536 ( .A(n2434), .B(n2433), .Z(n2435) );
  NAND U4537 ( .A(n2436), .B(n2435), .Z(n2444) );
  XNOR U4538 ( .A(n2443), .B(n2444), .Z(n2448) );
  XNOR U4539 ( .A(n2438), .B(n2437), .Z(n2447) );
  NAND U4540 ( .A(n2448), .B(n2447), .Z(n2439) );
  AND U4541 ( .A(n2440), .B(n2439), .Z(n2674) );
  NANDN U4542 ( .A(n2442), .B(n2441), .Z(n2446) );
  NANDN U4543 ( .A(n2444), .B(n2443), .Z(n2445) );
  AND U4544 ( .A(n2446), .B(n2445), .Z(n2668) );
  AND U4545 ( .A(b[62]), .B(a[17]), .Z(n2667) );
  XNOR U4546 ( .A(n2668), .B(n2667), .Z(n2669) );
  NAND U4547 ( .A(b[63]), .B(a[16]), .Z(n2670) );
  XNOR U4548 ( .A(n2669), .B(n2670), .Z(n2673) );
  XNOR U4549 ( .A(n2674), .B(n2673), .Z(n2676) );
  AND U4550 ( .A(a[18]), .B(b[61]), .Z(n2675) );
  XOR U4551 ( .A(n2676), .B(n2675), .Z(n2682) );
  AND U4552 ( .A(a[19]), .B(b[60]), .Z(n2680) );
  XOR U4553 ( .A(n2448), .B(n2447), .Z(n2548) );
  NAND U4554 ( .A(a[16]), .B(b[60]), .Z(n2451) );
  XNOR U4555 ( .A(n2450), .B(n2449), .Z(n2452) );
  NANDN U4556 ( .A(n2451), .B(n2452), .Z(n2540) );
  XNOR U4557 ( .A(n2452), .B(n2451), .Z(n2554) );
  XOR U4558 ( .A(n2454), .B(n2453), .Z(n2536) );
  XOR U4559 ( .A(n2456), .B(n2455), .Z(n2532) );
  XOR U4560 ( .A(n2458), .B(n2457), .Z(n2528) );
  XOR U4561 ( .A(n2460), .B(n2459), .Z(n2524) );
  XOR U4562 ( .A(n2462), .B(n2461), .Z(n2514) );
  XOR U4563 ( .A(n2464), .B(n2463), .Z(n2510) );
  XOR U4564 ( .A(n2466), .B(n2465), .Z(n2506) );
  XOR U4565 ( .A(n2468), .B(n2467), .Z(n2490) );
  XOR U4566 ( .A(n2470), .B(n2469), .Z(n2479) );
  NAND U4567 ( .A(a[0]), .B(b[60]), .Z(n3156) );
  AND U4568 ( .A(a[1]), .B(b[61]), .Z(n2474) );
  NANDN U4569 ( .A(n3156), .B(n2474), .Z(n2579) );
  OR U4570 ( .A(n2579), .B(n2471), .Z(n2478) );
  ANDN U4571 ( .B(n2474), .A(n3156), .Z(n2472) );
  XNOR U4572 ( .A(n2472), .B(n2471), .Z(n2476) );
  OR U4573 ( .A(n2474), .B(n2473), .Z(n2475) );
  NAND U4574 ( .A(n2476), .B(n2475), .Z(n2587) );
  AND U4575 ( .A(a[2]), .B(b[60]), .Z(n2588) );
  NANDN U4576 ( .A(n2587), .B(n2588), .Z(n2477) );
  AND U4577 ( .A(n2478), .B(n2477), .Z(n2480) );
  NANDN U4578 ( .A(n2479), .B(n2480), .Z(n2482) );
  AND U4579 ( .A(a[3]), .B(b[60]), .Z(n2594) );
  NANDN U4580 ( .A(n2594), .B(n2593), .Z(n2481) );
  AND U4581 ( .A(n2482), .B(n2481), .Z(n2486) );
  NAND U4582 ( .A(n2486), .B(n2485), .Z(n2488) );
  AND U4583 ( .A(a[4]), .B(b[60]), .Z(n2578) );
  XOR U4584 ( .A(n2486), .B(n2485), .Z(n2577) );
  NAND U4585 ( .A(n2578), .B(n2577), .Z(n2487) );
  NAND U4586 ( .A(n2488), .B(n2487), .Z(n2489) );
  NANDN U4587 ( .A(n2490), .B(n2489), .Z(n2492) );
  XNOR U4588 ( .A(n2490), .B(n2489), .Z(n2604) );
  AND U4589 ( .A(a[5]), .B(b[60]), .Z(n2603) );
  NAND U4590 ( .A(n2604), .B(n2603), .Z(n2491) );
  AND U4591 ( .A(n2492), .B(n2491), .Z(n2496) );
  AND U4592 ( .A(a[6]), .B(b[60]), .Z(n2495) );
  NANDN U4593 ( .A(n2496), .B(n2495), .Z(n2498) );
  XOR U4594 ( .A(n2494), .B(n2493), .Z(n2573) );
  XNOR U4595 ( .A(n2496), .B(n2495), .Z(n2574) );
  NANDN U4596 ( .A(n2573), .B(n2574), .Z(n2497) );
  NAND U4597 ( .A(n2498), .B(n2497), .Z(n2501) );
  XNOR U4598 ( .A(n2500), .B(n2499), .Z(n2502) );
  NANDN U4599 ( .A(n2501), .B(n2502), .Z(n2504) );
  XOR U4600 ( .A(n2502), .B(n2501), .Z(n2571) );
  AND U4601 ( .A(a[7]), .B(b[60]), .Z(n2572) );
  OR U4602 ( .A(n2571), .B(n2572), .Z(n2503) );
  NAND U4603 ( .A(n2504), .B(n2503), .Z(n2505) );
  NANDN U4604 ( .A(n2506), .B(n2505), .Z(n2508) );
  XOR U4605 ( .A(n2506), .B(n2505), .Z(n2569) );
  AND U4606 ( .A(a[8]), .B(b[60]), .Z(n2570) );
  OR U4607 ( .A(n2569), .B(n2570), .Z(n2507) );
  NAND U4608 ( .A(n2508), .B(n2507), .Z(n2509) );
  NANDN U4609 ( .A(n2510), .B(n2509), .Z(n2512) );
  XOR U4610 ( .A(n2510), .B(n2509), .Z(n2567) );
  AND U4611 ( .A(a[9]), .B(b[60]), .Z(n2568) );
  OR U4612 ( .A(n2567), .B(n2568), .Z(n2511) );
  NAND U4613 ( .A(n2512), .B(n2511), .Z(n2513) );
  NANDN U4614 ( .A(n2514), .B(n2513), .Z(n2516) );
  AND U4615 ( .A(a[10]), .B(b[60]), .Z(n2566) );
  XNOR U4616 ( .A(n2514), .B(n2513), .Z(n2565) );
  NANDN U4617 ( .A(n2566), .B(n2565), .Z(n2515) );
  AND U4618 ( .A(n2516), .B(n2515), .Z(n2520) );
  XNOR U4619 ( .A(n2518), .B(n2517), .Z(n2519) );
  NANDN U4620 ( .A(n2520), .B(n2519), .Z(n2522) );
  XOR U4621 ( .A(n2520), .B(n2519), .Z(n2563) );
  AND U4622 ( .A(a[11]), .B(b[60]), .Z(n2564) );
  OR U4623 ( .A(n2563), .B(n2564), .Z(n2521) );
  NAND U4624 ( .A(n2522), .B(n2521), .Z(n2523) );
  NANDN U4625 ( .A(n2524), .B(n2523), .Z(n2526) );
  XOR U4626 ( .A(n2524), .B(n2523), .Z(n2559) );
  AND U4627 ( .A(a[12]), .B(b[60]), .Z(n2560) );
  OR U4628 ( .A(n2559), .B(n2560), .Z(n2525) );
  NAND U4629 ( .A(n2526), .B(n2525), .Z(n2527) );
  NANDN U4630 ( .A(n2528), .B(n2527), .Z(n2530) );
  AND U4631 ( .A(a[13]), .B(b[60]), .Z(n2558) );
  XNOR U4632 ( .A(n2528), .B(n2527), .Z(n2557) );
  NANDN U4633 ( .A(n2558), .B(n2557), .Z(n2529) );
  NAND U4634 ( .A(n2530), .B(n2529), .Z(n2531) );
  NANDN U4635 ( .A(n2532), .B(n2531), .Z(n2534) );
  AND U4636 ( .A(a[14]), .B(b[60]), .Z(n2638) );
  XNOR U4637 ( .A(n2532), .B(n2531), .Z(n2637) );
  NANDN U4638 ( .A(n2638), .B(n2637), .Z(n2533) );
  NAND U4639 ( .A(n2534), .B(n2533), .Z(n2535) );
  NANDN U4640 ( .A(n2536), .B(n2535), .Z(n2538) );
  AND U4641 ( .A(a[15]), .B(b[60]), .Z(n2556) );
  XNOR U4642 ( .A(n2536), .B(n2535), .Z(n2555) );
  NANDN U4643 ( .A(n2556), .B(n2555), .Z(n2537) );
  AND U4644 ( .A(n2538), .B(n2537), .Z(n2553) );
  NAND U4645 ( .A(n2554), .B(n2553), .Z(n2539) );
  AND U4646 ( .A(n2540), .B(n2539), .Z(n2542) );
  AND U4647 ( .A(a[17]), .B(b[60]), .Z(n2541) );
  NANDN U4648 ( .A(n2542), .B(n2541), .Z(n2546) );
  XNOR U4649 ( .A(n2542), .B(n2541), .Z(n2652) );
  XNOR U4650 ( .A(n2544), .B(n2543), .Z(n2651) );
  NAND U4651 ( .A(n2652), .B(n2651), .Z(n2545) );
  AND U4652 ( .A(n2546), .B(n2545), .Z(n2547) );
  NANDN U4653 ( .A(n2548), .B(n2547), .Z(n2550) );
  AND U4654 ( .A(a[18]), .B(b[60]), .Z(n2552) );
  XNOR U4655 ( .A(n2548), .B(n2547), .Z(n2551) );
  NANDN U4656 ( .A(n2552), .B(n2551), .Z(n2549) );
  NAND U4657 ( .A(n2550), .B(n2549), .Z(n2679) );
  XNOR U4658 ( .A(n2680), .B(n2679), .Z(n2681) );
  XOR U4659 ( .A(n2682), .B(n2681), .Z(n2662) );
  AND U4660 ( .A(a[19]), .B(b[59]), .Z(n2657) );
  XOR U4661 ( .A(n2552), .B(n2551), .Z(n2658) );
  NAND U4662 ( .A(n2657), .B(n2658), .Z(n2660) );
  XOR U4663 ( .A(n2554), .B(n2553), .Z(n2648) );
  AND U4664 ( .A(a[16]), .B(b[59]), .Z(n2643) );
  XOR U4665 ( .A(n2556), .B(n2555), .Z(n2644) );
  NAND U4666 ( .A(n2643), .B(n2644), .Z(n2646) );
  XOR U4667 ( .A(n2558), .B(n2557), .Z(n2634) );
  AND U4668 ( .A(a[14]), .B(b[59]), .Z(n2633) );
  NAND U4669 ( .A(n2634), .B(n2633), .Z(n2636) );
  XOR U4670 ( .A(n2560), .B(n2559), .Z(n2562) );
  AND U4671 ( .A(a[13]), .B(b[59]), .Z(n2561) );
  NANDN U4672 ( .A(n2562), .B(n2561), .Z(n2632) );
  XOR U4673 ( .A(n2562), .B(n2561), .Z(n3137) );
  XOR U4674 ( .A(n2564), .B(n2563), .Z(n2628) );
  XOR U4675 ( .A(n2566), .B(n2565), .Z(n2623) );
  XOR U4676 ( .A(n2568), .B(n2567), .Z(n2620) );
  XOR U4677 ( .A(n2570), .B(n2569), .Z(n2616) );
  XOR U4678 ( .A(n2572), .B(n2571), .Z(n2612) );
  AND U4679 ( .A(a[8]), .B(b[59]), .Z(n2611) );
  NANDN U4680 ( .A(n2612), .B(n2611), .Z(n2614) );
  NAND U4681 ( .A(a[7]), .B(b[59]), .Z(n2575) );
  XNOR U4682 ( .A(n2574), .B(n2573), .Z(n2576) );
  NANDN U4683 ( .A(n2575), .B(n2576), .Z(n2610) );
  XOR U4684 ( .A(n2576), .B(n2575), .Z(n3186) );
  XOR U4685 ( .A(n2578), .B(n2577), .Z(n2599) );
  NAND U4686 ( .A(a[0]), .B(b[59]), .Z(n3393) );
  AND U4687 ( .A(a[1]), .B(b[60]), .Z(n2582) );
  NANDN U4688 ( .A(n3393), .B(n2582), .Z(n3155) );
  NANDN U4689 ( .A(n3155), .B(n2579), .Z(n2586) );
  ANDN U4690 ( .B(n2582), .A(n3393), .Z(n2580) );
  XOR U4691 ( .A(n2580), .B(n2579), .Z(n2584) );
  OR U4692 ( .A(n2582), .B(n2581), .Z(n2583) );
  NAND U4693 ( .A(n2584), .B(n2583), .Z(n3160) );
  AND U4694 ( .A(a[2]), .B(b[59]), .Z(n3161) );
  NANDN U4695 ( .A(n3160), .B(n3161), .Z(n2585) );
  AND U4696 ( .A(n2586), .B(n2585), .Z(n2589) );
  AND U4697 ( .A(a[3]), .B(b[59]), .Z(n2590) );
  NANDN U4698 ( .A(n2589), .B(n2590), .Z(n2592) );
  XNOR U4699 ( .A(n2588), .B(n2587), .Z(n3167) );
  NAND U4700 ( .A(n3167), .B(n3166), .Z(n2591) );
  AND U4701 ( .A(n2592), .B(n2591), .Z(n2595) );
  XOR U4702 ( .A(n2594), .B(n2593), .Z(n2596) );
  NANDN U4703 ( .A(n2595), .B(n2596), .Z(n2598) );
  AND U4704 ( .A(a[4]), .B(b[59]), .Z(n3154) );
  NAND U4705 ( .A(n3154), .B(n3153), .Z(n2597) );
  AND U4706 ( .A(n2598), .B(n2597), .Z(n2600) );
  NANDN U4707 ( .A(n2599), .B(n2600), .Z(n2602) );
  AND U4708 ( .A(a[5]), .B(b[59]), .Z(n3176) );
  NANDN U4709 ( .A(n3176), .B(n3177), .Z(n2601) );
  AND U4710 ( .A(n2602), .B(n2601), .Z(n2606) );
  XNOR U4711 ( .A(n2604), .B(n2603), .Z(n2605) );
  NANDN U4712 ( .A(n2606), .B(n2605), .Z(n2608) );
  XOR U4713 ( .A(n2606), .B(n2605), .Z(n3151) );
  AND U4714 ( .A(a[6]), .B(b[59]), .Z(n3152) );
  OR U4715 ( .A(n3151), .B(n3152), .Z(n2607) );
  AND U4716 ( .A(n2608), .B(n2607), .Z(n3187) );
  NANDN U4717 ( .A(n3186), .B(n3187), .Z(n2609) );
  AND U4718 ( .A(n2610), .B(n2609), .Z(n3148) );
  XNOR U4719 ( .A(n2612), .B(n2611), .Z(n3147) );
  NANDN U4720 ( .A(n3148), .B(n3147), .Z(n2613) );
  NAND U4721 ( .A(n2614), .B(n2613), .Z(n2615) );
  NANDN U4722 ( .A(n2616), .B(n2615), .Z(n2618) );
  NAND U4723 ( .A(a[9]), .B(b[59]), .Z(n3145) );
  XNOR U4724 ( .A(n2616), .B(n2615), .Z(n3146) );
  NANDN U4725 ( .A(n3145), .B(n3146), .Z(n2617) );
  NAND U4726 ( .A(n2618), .B(n2617), .Z(n2619) );
  NANDN U4727 ( .A(n2620), .B(n2619), .Z(n2622) );
  NAND U4728 ( .A(a[10]), .B(b[59]), .Z(n3198) );
  XNOR U4729 ( .A(n2620), .B(n2619), .Z(n3199) );
  NANDN U4730 ( .A(n3198), .B(n3199), .Z(n2621) );
  AND U4731 ( .A(n2622), .B(n2621), .Z(n2624) );
  NANDN U4732 ( .A(n2623), .B(n2624), .Z(n2626) );
  AND U4733 ( .A(a[11]), .B(b[59]), .Z(n3144) );
  XNOR U4734 ( .A(n2624), .B(n2623), .Z(n3143) );
  NANDN U4735 ( .A(n3144), .B(n3143), .Z(n2625) );
  AND U4736 ( .A(n2626), .B(n2625), .Z(n2627) );
  NANDN U4737 ( .A(n2628), .B(n2627), .Z(n2630) );
  XNOR U4738 ( .A(n2628), .B(n2627), .Z(n3140) );
  AND U4739 ( .A(a[12]), .B(b[59]), .Z(n3139) );
  NAND U4740 ( .A(n3140), .B(n3139), .Z(n2629) );
  AND U4741 ( .A(n2630), .B(n2629), .Z(n3138) );
  OR U4742 ( .A(n3137), .B(n3138), .Z(n2631) );
  AND U4743 ( .A(n2632), .B(n2631), .Z(n3136) );
  XOR U4744 ( .A(n2634), .B(n2633), .Z(n3135) );
  NANDN U4745 ( .A(n3136), .B(n3135), .Z(n2635) );
  AND U4746 ( .A(n2636), .B(n2635), .Z(n2640) );
  AND U4747 ( .A(a[15]), .B(b[59]), .Z(n2639) );
  NANDN U4748 ( .A(n2640), .B(n2639), .Z(n2642) );
  XOR U4749 ( .A(n2638), .B(n2637), .Z(n3134) );
  XNOR U4750 ( .A(n2640), .B(n2639), .Z(n3133) );
  NAND U4751 ( .A(n3134), .B(n3133), .Z(n2641) );
  AND U4752 ( .A(n2642), .B(n2641), .Z(n3132) );
  XOR U4753 ( .A(n2644), .B(n2643), .Z(n3131) );
  NANDN U4754 ( .A(n3132), .B(n3131), .Z(n2645) );
  AND U4755 ( .A(n2646), .B(n2645), .Z(n2647) );
  NANDN U4756 ( .A(n2648), .B(n2647), .Z(n2650) );
  AND U4757 ( .A(a[17]), .B(b[59]), .Z(n3130) );
  XNOR U4758 ( .A(n2648), .B(n2647), .Z(n3129) );
  NANDN U4759 ( .A(n3130), .B(n3129), .Z(n2649) );
  NAND U4760 ( .A(n2650), .B(n2649), .Z(n2653) );
  XOR U4761 ( .A(n2652), .B(n2651), .Z(n2654) );
  NANDN U4762 ( .A(n2653), .B(n2654), .Z(n2656) );
  NAND U4763 ( .A(a[18]), .B(b[59]), .Z(n3127) );
  XNOR U4764 ( .A(n2654), .B(n2653), .Z(n3128) );
  NANDN U4765 ( .A(n3127), .B(n3128), .Z(n2655) );
  AND U4766 ( .A(n2656), .B(n2655), .Z(n3233) );
  XOR U4767 ( .A(n2658), .B(n2657), .Z(n3232) );
  NANDN U4768 ( .A(n3233), .B(n3232), .Z(n2659) );
  NAND U4769 ( .A(n2660), .B(n2659), .Z(n2661) );
  NAND U4770 ( .A(n2662), .B(n2661), .Z(n2664) );
  XOR U4771 ( .A(n2662), .B(n2661), .Z(n3126) );
  AND U4772 ( .A(a[20]), .B(b[59]), .Z(n3125) );
  NAND U4773 ( .A(n3126), .B(n3125), .Z(n2663) );
  AND U4774 ( .A(n2664), .B(n2663), .Z(n2666) );
  AND U4775 ( .A(a[21]), .B(b[59]), .Z(n2665) );
  NANDN U4776 ( .A(n2666), .B(n2665), .Z(n2686) );
  XNOR U4777 ( .A(n2666), .B(n2665), .Z(n3123) );
  AND U4778 ( .A(b[63]), .B(a[17]), .Z(n2698) );
  AND U4779 ( .A(b[62]), .B(a[18]), .Z(n2696) );
  NANDN U4780 ( .A(n2668), .B(n2667), .Z(n2672) );
  NANDN U4781 ( .A(n2670), .B(n2669), .Z(n2671) );
  AND U4782 ( .A(n2672), .B(n2671), .Z(n2695) );
  XNOR U4783 ( .A(n2696), .B(n2695), .Z(n2697) );
  XOR U4784 ( .A(n2698), .B(n2697), .Z(n2691) );
  NANDN U4785 ( .A(n2674), .B(n2673), .Z(n2678) );
  NAND U4786 ( .A(n2676), .B(n2675), .Z(n2677) );
  AND U4787 ( .A(n2678), .B(n2677), .Z(n2690) );
  AND U4788 ( .A(a[19]), .B(b[61]), .Z(n2689) );
  XNOR U4789 ( .A(n2690), .B(n2689), .Z(n2692) );
  XNOR U4790 ( .A(n2691), .B(n2692), .Z(n2703) );
  AND U4791 ( .A(a[20]), .B(b[60]), .Z(n2702) );
  NANDN U4792 ( .A(n2680), .B(n2679), .Z(n2684) );
  NANDN U4793 ( .A(n2682), .B(n2681), .Z(n2683) );
  NAND U4794 ( .A(n2684), .B(n2683), .Z(n2701) );
  XNOR U4795 ( .A(n2702), .B(n2701), .Z(n2704) );
  XNOR U4796 ( .A(n2703), .B(n2704), .Z(n3124) );
  NAND U4797 ( .A(n3123), .B(n3124), .Z(n2685) );
  AND U4798 ( .A(n2686), .B(n2685), .Z(n2688) );
  AND U4799 ( .A(a[22]), .B(b[59]), .Z(n2687) );
  NANDN U4800 ( .A(n2688), .B(n2687), .Z(n2708) );
  XNOR U4801 ( .A(n2688), .B(n2687), .Z(n3247) );
  AND U4802 ( .A(a[20]), .B(b[61]), .Z(n2722) );
  NANDN U4803 ( .A(n2690), .B(n2689), .Z(n2694) );
  NAND U4804 ( .A(n2692), .B(n2691), .Z(n2693) );
  AND U4805 ( .A(n2694), .B(n2693), .Z(n2721) );
  XNOR U4806 ( .A(n2722), .B(n2721), .Z(n2724) );
  AND U4807 ( .A(b[63]), .B(a[18]), .Z(n2718) );
  AND U4808 ( .A(b[62]), .B(a[19]), .Z(n2716) );
  NANDN U4809 ( .A(n2696), .B(n2695), .Z(n2700) );
  NANDN U4810 ( .A(n2698), .B(n2697), .Z(n2699) );
  NAND U4811 ( .A(n2700), .B(n2699), .Z(n2715) );
  XNOR U4812 ( .A(n2716), .B(n2715), .Z(n2717) );
  XNOR U4813 ( .A(n2718), .B(n2717), .Z(n2723) );
  XOR U4814 ( .A(n2724), .B(n2723), .Z(n2712) );
  NANDN U4815 ( .A(n2702), .B(n2701), .Z(n2706) );
  NAND U4816 ( .A(n2704), .B(n2703), .Z(n2705) );
  AND U4817 ( .A(n2706), .B(n2705), .Z(n2709) );
  NAND U4818 ( .A(a[21]), .B(b[60]), .Z(n2710) );
  XNOR U4819 ( .A(n2709), .B(n2710), .Z(n2711) );
  XNOR U4820 ( .A(n2712), .B(n2711), .Z(n3246) );
  NAND U4821 ( .A(n3247), .B(n3246), .Z(n2707) );
  AND U4822 ( .A(n2708), .B(n2707), .Z(n2728) );
  AND U4823 ( .A(a[23]), .B(b[59]), .Z(n2727) );
  NANDN U4824 ( .A(n2728), .B(n2727), .Z(n2730) );
  NANDN U4825 ( .A(n2710), .B(n2709), .Z(n2714) );
  NANDN U4826 ( .A(n2712), .B(n2711), .Z(n2713) );
  AND U4827 ( .A(n2714), .B(n2713), .Z(n2746) );
  AND U4828 ( .A(a[22]), .B(b[60]), .Z(n2745) );
  XNOR U4829 ( .A(n2746), .B(n2745), .Z(n2748) );
  AND U4830 ( .A(b[63]), .B(a[19]), .Z(n2736) );
  AND U4831 ( .A(b[62]), .B(a[20]), .Z(n2734) );
  NANDN U4832 ( .A(n2716), .B(n2715), .Z(n2720) );
  NANDN U4833 ( .A(n2718), .B(n2717), .Z(n2719) );
  NAND U4834 ( .A(n2720), .B(n2719), .Z(n2733) );
  XNOR U4835 ( .A(n2734), .B(n2733), .Z(n2735) );
  XOR U4836 ( .A(n2736), .B(n2735), .Z(n2739) );
  NANDN U4837 ( .A(n2722), .B(n2721), .Z(n2726) );
  NAND U4838 ( .A(n2724), .B(n2723), .Z(n2725) );
  AND U4839 ( .A(n2726), .B(n2725), .Z(n2740) );
  XOR U4840 ( .A(n2739), .B(n2740), .Z(n2741) );
  NAND U4841 ( .A(a[21]), .B(b[61]), .Z(n2742) );
  XNOR U4842 ( .A(n2741), .B(n2742), .Z(n2747) );
  XOR U4843 ( .A(n2748), .B(n2747), .Z(n3253) );
  XNOR U4844 ( .A(n2728), .B(n2727), .Z(n3252) );
  NAND U4845 ( .A(n3253), .B(n3252), .Z(n2729) );
  AND U4846 ( .A(n2730), .B(n2729), .Z(n2732) );
  AND U4847 ( .A(a[24]), .B(b[59]), .Z(n2731) );
  NANDN U4848 ( .A(n2732), .B(n2731), .Z(n2752) );
  XNOR U4849 ( .A(n2732), .B(n2731), .Z(n3259) );
  AND U4850 ( .A(b[63]), .B(a[20]), .Z(n2768) );
  AND U4851 ( .A(b[62]), .B(a[21]), .Z(n2766) );
  NANDN U4852 ( .A(n2734), .B(n2733), .Z(n2738) );
  NANDN U4853 ( .A(n2736), .B(n2735), .Z(n2737) );
  NAND U4854 ( .A(n2738), .B(n2737), .Z(n2765) );
  XNOR U4855 ( .A(n2766), .B(n2765), .Z(n2767) );
  XOR U4856 ( .A(n2768), .B(n2767), .Z(n2760) );
  NAND U4857 ( .A(n2740), .B(n2739), .Z(n2744) );
  NANDN U4858 ( .A(n2742), .B(n2741), .Z(n2743) );
  NAND U4859 ( .A(n2744), .B(n2743), .Z(n2759) );
  XOR U4860 ( .A(n2760), .B(n2759), .Z(n2761) );
  NAND U4861 ( .A(a[22]), .B(b[61]), .Z(n2762) );
  XNOR U4862 ( .A(n2761), .B(n2762), .Z(n2756) );
  NANDN U4863 ( .A(n2746), .B(n2745), .Z(n2750) );
  NAND U4864 ( .A(n2748), .B(n2747), .Z(n2749) );
  AND U4865 ( .A(n2750), .B(n2749), .Z(n2754) );
  AND U4866 ( .A(a[23]), .B(b[60]), .Z(n2753) );
  XNOR U4867 ( .A(n2754), .B(n2753), .Z(n2755) );
  XOR U4868 ( .A(n2756), .B(n2755), .Z(n3258) );
  NAND U4869 ( .A(n3259), .B(n3258), .Z(n2751) );
  AND U4870 ( .A(n2752), .B(n2751), .Z(n2772) );
  AND U4871 ( .A(a[25]), .B(b[59]), .Z(n2771) );
  NANDN U4872 ( .A(n2772), .B(n2771), .Z(n2774) );
  AND U4873 ( .A(a[24]), .B(b[60]), .Z(n2778) );
  NANDN U4874 ( .A(n2754), .B(n2753), .Z(n2758) );
  NAND U4875 ( .A(n2756), .B(n2755), .Z(n2757) );
  AND U4876 ( .A(n2758), .B(n2757), .Z(n2777) );
  XNOR U4877 ( .A(n2778), .B(n2777), .Z(n2780) );
  AND U4878 ( .A(a[23]), .B(b[61]), .Z(n2792) );
  NAND U4879 ( .A(n2760), .B(n2759), .Z(n2764) );
  NANDN U4880 ( .A(n2762), .B(n2761), .Z(n2763) );
  AND U4881 ( .A(n2764), .B(n2763), .Z(n2790) );
  AND U4882 ( .A(b[63]), .B(a[21]), .Z(n2786) );
  AND U4883 ( .A(b[62]), .B(a[22]), .Z(n2784) );
  NANDN U4884 ( .A(n2766), .B(n2765), .Z(n2770) );
  NANDN U4885 ( .A(n2768), .B(n2767), .Z(n2769) );
  NAND U4886 ( .A(n2770), .B(n2769), .Z(n2783) );
  XNOR U4887 ( .A(n2784), .B(n2783), .Z(n2785) );
  XNOR U4888 ( .A(n2786), .B(n2785), .Z(n2789) );
  XOR U4889 ( .A(n2790), .B(n2789), .Z(n2791) );
  XNOR U4890 ( .A(n2792), .B(n2791), .Z(n2779) );
  XOR U4891 ( .A(n2780), .B(n2779), .Z(n3267) );
  XNOR U4892 ( .A(n2772), .B(n2771), .Z(n3266) );
  NANDN U4893 ( .A(n3267), .B(n3266), .Z(n2773) );
  AND U4894 ( .A(n2774), .B(n2773), .Z(n2776) );
  AND U4895 ( .A(a[26]), .B(b[59]), .Z(n2775) );
  NANDN U4896 ( .A(n2776), .B(n2775), .Z(n2796) );
  XNOR U4897 ( .A(n2776), .B(n2775), .Z(n3271) );
  NANDN U4898 ( .A(n2778), .B(n2777), .Z(n2782) );
  NAND U4899 ( .A(n2780), .B(n2779), .Z(n2781) );
  AND U4900 ( .A(n2782), .B(n2781), .Z(n2811) );
  NAND U4901 ( .A(a[25]), .B(b[60]), .Z(n2812) );
  XNOR U4902 ( .A(n2811), .B(n2812), .Z(n2814) );
  AND U4903 ( .A(b[63]), .B(a[22]), .Z(n2802) );
  AND U4904 ( .A(b[62]), .B(a[23]), .Z(n2800) );
  NANDN U4905 ( .A(n2784), .B(n2783), .Z(n2788) );
  NANDN U4906 ( .A(n2786), .B(n2785), .Z(n2787) );
  NAND U4907 ( .A(n2788), .B(n2787), .Z(n2799) );
  XNOR U4908 ( .A(n2800), .B(n2799), .Z(n2801) );
  XOR U4909 ( .A(n2802), .B(n2801), .Z(n2805) );
  NAND U4910 ( .A(n2790), .B(n2789), .Z(n2794) );
  NANDN U4911 ( .A(n2792), .B(n2791), .Z(n2793) );
  AND U4912 ( .A(n2794), .B(n2793), .Z(n2806) );
  XOR U4913 ( .A(n2805), .B(n2806), .Z(n2807) );
  NAND U4914 ( .A(a[24]), .B(b[61]), .Z(n2808) );
  XNOR U4915 ( .A(n2807), .B(n2808), .Z(n2813) );
  XOR U4916 ( .A(n2814), .B(n2813), .Z(n3270) );
  NAND U4917 ( .A(n3271), .B(n3270), .Z(n2795) );
  AND U4918 ( .A(n2796), .B(n2795), .Z(n2798) );
  AND U4919 ( .A(a[27]), .B(b[59]), .Z(n2797) );
  NANDN U4920 ( .A(n2798), .B(n2797), .Z(n2818) );
  XNOR U4921 ( .A(n2798), .B(n2797), .Z(n3276) );
  AND U4922 ( .A(a[25]), .B(b[61]), .Z(n2830) );
  AND U4923 ( .A(b[63]), .B(a[23]), .Z(n2824) );
  AND U4924 ( .A(b[62]), .B(a[24]), .Z(n2822) );
  NANDN U4925 ( .A(n2800), .B(n2799), .Z(n2804) );
  NANDN U4926 ( .A(n2802), .B(n2801), .Z(n2803) );
  NAND U4927 ( .A(n2804), .B(n2803), .Z(n2821) );
  XNOR U4928 ( .A(n2822), .B(n2821), .Z(n2823) );
  XOR U4929 ( .A(n2824), .B(n2823), .Z(n2828) );
  NAND U4930 ( .A(n2806), .B(n2805), .Z(n2810) );
  NANDN U4931 ( .A(n2808), .B(n2807), .Z(n2809) );
  NAND U4932 ( .A(n2810), .B(n2809), .Z(n2827) );
  XOR U4933 ( .A(n2828), .B(n2827), .Z(n2829) );
  XOR U4934 ( .A(n2830), .B(n2829), .Z(n2836) );
  AND U4935 ( .A(a[26]), .B(b[60]), .Z(n2834) );
  NANDN U4936 ( .A(n2812), .B(n2811), .Z(n2816) );
  NAND U4937 ( .A(n2814), .B(n2813), .Z(n2815) );
  AND U4938 ( .A(n2816), .B(n2815), .Z(n2833) );
  XNOR U4939 ( .A(n2834), .B(n2833), .Z(n2835) );
  XOR U4940 ( .A(n2836), .B(n2835), .Z(n3277) );
  NAND U4941 ( .A(n3276), .B(n3277), .Z(n2817) );
  AND U4942 ( .A(n2818), .B(n2817), .Z(n2820) );
  AND U4943 ( .A(a[28]), .B(b[59]), .Z(n2819) );
  NANDN U4944 ( .A(n2820), .B(n2819), .Z(n2840) );
  XNOR U4945 ( .A(n2820), .B(n2819), .Z(n3282) );
  AND U4946 ( .A(a[26]), .B(b[61]), .Z(n2846) );
  AND U4947 ( .A(b[63]), .B(a[24]), .Z(n2852) );
  AND U4948 ( .A(b[62]), .B(a[25]), .Z(n2850) );
  NANDN U4949 ( .A(n2822), .B(n2821), .Z(n2826) );
  NANDN U4950 ( .A(n2824), .B(n2823), .Z(n2825) );
  NAND U4951 ( .A(n2826), .B(n2825), .Z(n2849) );
  NAND U4952 ( .A(n2828), .B(n2827), .Z(n2832) );
  NAND U4953 ( .A(n2830), .B(n2829), .Z(n2831) );
  NAND U4954 ( .A(n2832), .B(n2831), .Z(n2843) );
  XOR U4955 ( .A(n2844), .B(n2843), .Z(n2845) );
  XOR U4956 ( .A(n2846), .B(n2845), .Z(n2858) );
  AND U4957 ( .A(a[27]), .B(b[60]), .Z(n2856) );
  NANDN U4958 ( .A(n2834), .B(n2833), .Z(n2838) );
  NANDN U4959 ( .A(n2836), .B(n2835), .Z(n2837) );
  NAND U4960 ( .A(n2838), .B(n2837), .Z(n2855) );
  XNOR U4961 ( .A(n2856), .B(n2855), .Z(n2857) );
  XOR U4962 ( .A(n2858), .B(n2857), .Z(n3283) );
  NAND U4963 ( .A(n3282), .B(n3283), .Z(n2839) );
  AND U4964 ( .A(n2840), .B(n2839), .Z(n2842) );
  AND U4965 ( .A(a[29]), .B(b[59]), .Z(n2841) );
  NANDN U4966 ( .A(n2842), .B(n2841), .Z(n2862) );
  XNOR U4967 ( .A(n2842), .B(n2841), .Z(n3288) );
  AND U4968 ( .A(a[27]), .B(b[61]), .Z(n2874) );
  NAND U4969 ( .A(n2844), .B(n2843), .Z(n2848) );
  NAND U4970 ( .A(n2846), .B(n2845), .Z(n2847) );
  AND U4971 ( .A(n2848), .B(n2847), .Z(n2872) );
  AND U4972 ( .A(b[63]), .B(a[25]), .Z(n2868) );
  AND U4973 ( .A(b[62]), .B(a[26]), .Z(n2866) );
  NANDN U4974 ( .A(n2850), .B(n2849), .Z(n2854) );
  NANDN U4975 ( .A(n2852), .B(n2851), .Z(n2853) );
  NAND U4976 ( .A(n2854), .B(n2853), .Z(n2865) );
  XOR U4977 ( .A(n2868), .B(n2867), .Z(n2871) );
  XNOR U4978 ( .A(n2872), .B(n2871), .Z(n2873) );
  XOR U4979 ( .A(n2874), .B(n2873), .Z(n2880) );
  AND U4980 ( .A(a[28]), .B(b[60]), .Z(n2878) );
  NANDN U4981 ( .A(n2856), .B(n2855), .Z(n2860) );
  NANDN U4982 ( .A(n2858), .B(n2857), .Z(n2859) );
  NAND U4983 ( .A(n2860), .B(n2859), .Z(n2877) );
  XNOR U4984 ( .A(n2878), .B(n2877), .Z(n2879) );
  XOR U4985 ( .A(n2880), .B(n2879), .Z(n3289) );
  NAND U4986 ( .A(n3288), .B(n3289), .Z(n2861) );
  AND U4987 ( .A(n2862), .B(n2861), .Z(n2864) );
  AND U4988 ( .A(a[30]), .B(b[59]), .Z(n2863) );
  NANDN U4989 ( .A(n2864), .B(n2863), .Z(n2884) );
  XNOR U4990 ( .A(n2864), .B(n2863), .Z(n3295) );
  AND U4991 ( .A(b[63]), .B(a[26]), .Z(n2896) );
  AND U4992 ( .A(b[62]), .B(a[27]), .Z(n2894) );
  NANDN U4993 ( .A(n2866), .B(n2865), .Z(n2870) );
  NANDN U4994 ( .A(n2868), .B(n2867), .Z(n2869) );
  NAND U4995 ( .A(n2870), .B(n2869), .Z(n2893) );
  NANDN U4996 ( .A(n2872), .B(n2871), .Z(n2876) );
  NAND U4997 ( .A(n2874), .B(n2873), .Z(n2875) );
  AND U4998 ( .A(n2876), .B(n2875), .Z(n2900) );
  AND U4999 ( .A(a[28]), .B(b[61]), .Z(n2899) );
  XNOR U5000 ( .A(n2900), .B(n2899), .Z(n2902) );
  XOR U5001 ( .A(n2901), .B(n2902), .Z(n2890) );
  NANDN U5002 ( .A(n2878), .B(n2877), .Z(n2882) );
  NANDN U5003 ( .A(n2880), .B(n2879), .Z(n2881) );
  AND U5004 ( .A(n2882), .B(n2881), .Z(n2887) );
  NAND U5005 ( .A(a[29]), .B(b[60]), .Z(n2888) );
  XNOR U5006 ( .A(n2887), .B(n2888), .Z(n2889) );
  XOR U5007 ( .A(n2890), .B(n2889), .Z(n3294) );
  NAND U5008 ( .A(n3295), .B(n3294), .Z(n2883) );
  AND U5009 ( .A(n2884), .B(n2883), .Z(n2885) );
  NANDN U5010 ( .A(n2886), .B(n2885), .Z(n2906) );
  XNOR U5011 ( .A(n2886), .B(n2885), .Z(n3303) );
  AND U5012 ( .A(a[30]), .B(b[60]), .Z(n2922) );
  NANDN U5013 ( .A(n2888), .B(n2887), .Z(n2892) );
  NAND U5014 ( .A(n2890), .B(n2889), .Z(n2891) );
  AND U5015 ( .A(n2892), .B(n2891), .Z(n2921) );
  XNOR U5016 ( .A(n2922), .B(n2921), .Z(n2924) );
  AND U5017 ( .A(a[29]), .B(b[61]), .Z(n2912) );
  AND U5018 ( .A(b[63]), .B(a[27]), .Z(n2918) );
  AND U5019 ( .A(b[62]), .B(a[28]), .Z(n2916) );
  NANDN U5020 ( .A(n2894), .B(n2893), .Z(n2898) );
  NANDN U5021 ( .A(n2896), .B(n2895), .Z(n2897) );
  NAND U5022 ( .A(n2898), .B(n2897), .Z(n2915) );
  NANDN U5023 ( .A(n2900), .B(n2899), .Z(n2904) );
  NAND U5024 ( .A(n2902), .B(n2901), .Z(n2903) );
  NAND U5025 ( .A(n2904), .B(n2903), .Z(n2910) );
  XNOR U5026 ( .A(n2909), .B(n2910), .Z(n2911) );
  XNOR U5027 ( .A(n2912), .B(n2911), .Z(n2923) );
  XOR U5028 ( .A(n2924), .B(n2923), .Z(n3302) );
  NAND U5029 ( .A(n3303), .B(n3302), .Z(n2905) );
  AND U5030 ( .A(n2906), .B(n2905), .Z(n2908) );
  NANDN U5031 ( .A(n2907), .B(n2908), .Z(n2928) );
  AND U5032 ( .A(a[30]), .B(b[61]), .Z(n2940) );
  NANDN U5033 ( .A(n2910), .B(n2909), .Z(n2914) );
  NANDN U5034 ( .A(n2912), .B(n2911), .Z(n2913) );
  AND U5035 ( .A(n2914), .B(n2913), .Z(n2938) );
  AND U5036 ( .A(b[63]), .B(a[28]), .Z(n2934) );
  AND U5037 ( .A(b[62]), .B(a[29]), .Z(n2932) );
  NANDN U5038 ( .A(n2916), .B(n2915), .Z(n2920) );
  NANDN U5039 ( .A(n2918), .B(n2917), .Z(n2919) );
  NAND U5040 ( .A(n2920), .B(n2919), .Z(n2931) );
  XOR U5041 ( .A(n2938), .B(n2937), .Z(n2939) );
  XOR U5042 ( .A(n2940), .B(n2939), .Z(n2946) );
  AND U5043 ( .A(a[31]), .B(b[60]), .Z(n2944) );
  NANDN U5044 ( .A(n2922), .B(n2921), .Z(n2926) );
  NAND U5045 ( .A(n2924), .B(n2923), .Z(n2925) );
  NAND U5046 ( .A(n2926), .B(n2925), .Z(n2943) );
  NAND U5047 ( .A(n3308), .B(n3309), .Z(n2927) );
  AND U5048 ( .A(n2928), .B(n2927), .Z(n2929) );
  AND U5049 ( .A(a[33]), .B(b[59]), .Z(n2930) );
  NANDN U5050 ( .A(n2929), .B(n2930), .Z(n2950) );
  AND U5051 ( .A(b[63]), .B(a[29]), .Z(n2962) );
  AND U5052 ( .A(b[62]), .B(a[30]), .Z(n2960) );
  NANDN U5053 ( .A(n2932), .B(n2931), .Z(n2936) );
  NANDN U5054 ( .A(n2934), .B(n2933), .Z(n2935) );
  NAND U5055 ( .A(n2936), .B(n2935), .Z(n2959) );
  NAND U5056 ( .A(n2938), .B(n2937), .Z(n2942) );
  NAND U5057 ( .A(n2940), .B(n2939), .Z(n2941) );
  AND U5058 ( .A(n2942), .B(n2941), .Z(n2966) );
  AND U5059 ( .A(a[31]), .B(b[61]), .Z(n2965) );
  XOR U5060 ( .A(n2967), .B(n2968), .Z(n2956) );
  NANDN U5061 ( .A(n2944), .B(n2943), .Z(n2948) );
  NANDN U5062 ( .A(n2946), .B(n2945), .Z(n2947) );
  AND U5063 ( .A(n2948), .B(n2947), .Z(n2953) );
  NAND U5064 ( .A(a[32]), .B(b[60]), .Z(n2954) );
  XOR U5065 ( .A(n2956), .B(n2955), .Z(n3312) );
  NAND U5066 ( .A(n3313), .B(n3312), .Z(n2949) );
  AND U5067 ( .A(n2950), .B(n2949), .Z(n2952) );
  NANDN U5068 ( .A(n2951), .B(n2952), .Z(n2972) );
  AND U5069 ( .A(a[33]), .B(b[60]), .Z(n2974) );
  NANDN U5070 ( .A(n2954), .B(n2953), .Z(n2958) );
  NAND U5071 ( .A(n2956), .B(n2955), .Z(n2957) );
  AND U5072 ( .A(n2958), .B(n2957), .Z(n2973) );
  AND U5073 ( .A(a[32]), .B(b[61]), .Z(n2982) );
  AND U5074 ( .A(b[63]), .B(a[30]), .Z(n2988) );
  AND U5075 ( .A(b[62]), .B(a[31]), .Z(n2986) );
  NANDN U5076 ( .A(n2960), .B(n2959), .Z(n2964) );
  NANDN U5077 ( .A(n2962), .B(n2961), .Z(n2963) );
  NAND U5078 ( .A(n2964), .B(n2963), .Z(n2985) );
  NANDN U5079 ( .A(n2966), .B(n2965), .Z(n2970) );
  NAND U5080 ( .A(n2968), .B(n2967), .Z(n2969) );
  NAND U5081 ( .A(n2970), .B(n2969), .Z(n2980) );
  XOR U5082 ( .A(n2976), .B(n2975), .Z(n3318) );
  NAND U5083 ( .A(n3319), .B(n3318), .Z(n2971) );
  NAND U5084 ( .A(n2972), .B(n2971), .Z(n2991) );
  AND U5085 ( .A(a[35]), .B(b[59]), .Z(n2992) );
  NANDN U5086 ( .A(n2991), .B(n2992), .Z(n2994) );
  AND U5087 ( .A(a[34]), .B(b[60]), .Z(n3010) );
  NANDN U5088 ( .A(n2974), .B(n2973), .Z(n2978) );
  NAND U5089 ( .A(n2976), .B(n2975), .Z(n2977) );
  NAND U5090 ( .A(n2978), .B(n2977), .Z(n3009) );
  AND U5091 ( .A(a[33]), .B(b[61]), .Z(n3006) );
  NANDN U5092 ( .A(n2980), .B(n2979), .Z(n2984) );
  NANDN U5093 ( .A(n2982), .B(n2981), .Z(n2983) );
  AND U5094 ( .A(n2984), .B(n2983), .Z(n3004) );
  AND U5095 ( .A(b[63]), .B(a[31]), .Z(n3000) );
  AND U5096 ( .A(b[62]), .B(a[32]), .Z(n2998) );
  NANDN U5097 ( .A(n2986), .B(n2985), .Z(n2990) );
  NANDN U5098 ( .A(n2988), .B(n2987), .Z(n2989) );
  NAND U5099 ( .A(n2990), .B(n2989), .Z(n2997) );
  XOR U5100 ( .A(n3012), .B(n3011), .Z(n3326) );
  NANDN U5101 ( .A(n3326), .B(n3327), .Z(n2993) );
  AND U5102 ( .A(n2994), .B(n2993), .Z(n2995) );
  AND U5103 ( .A(a[36]), .B(b[59]), .Z(n2996) );
  NANDN U5104 ( .A(n2995), .B(n2996), .Z(n3016) );
  AND U5105 ( .A(b[63]), .B(a[32]), .Z(n3028) );
  AND U5106 ( .A(b[62]), .B(a[33]), .Z(n3026) );
  NANDN U5107 ( .A(n2998), .B(n2997), .Z(n3002) );
  NANDN U5108 ( .A(n3000), .B(n2999), .Z(n3001) );
  NAND U5109 ( .A(n3002), .B(n3001), .Z(n3025) );
  NANDN U5110 ( .A(n3004), .B(n3003), .Z(n3008) );
  NANDN U5111 ( .A(n3006), .B(n3005), .Z(n3007) );
  AND U5112 ( .A(n3008), .B(n3007), .Z(n3031) );
  NAND U5113 ( .A(a[34]), .B(b[61]), .Z(n3032) );
  XOR U5114 ( .A(n3033), .B(n3034), .Z(n3022) );
  AND U5115 ( .A(a[35]), .B(b[60]), .Z(n3019) );
  NANDN U5116 ( .A(n3010), .B(n3009), .Z(n3014) );
  NAND U5117 ( .A(n3012), .B(n3011), .Z(n3013) );
  NAND U5118 ( .A(n3014), .B(n3013), .Z(n3020) );
  XOR U5119 ( .A(n3022), .B(n3021), .Z(n3330) );
  NAND U5120 ( .A(n3331), .B(n3330), .Z(n3015) );
  AND U5121 ( .A(n3016), .B(n3015), .Z(n3018) );
  NANDN U5122 ( .A(n3017), .B(n3018), .Z(n3038) );
  AND U5123 ( .A(a[36]), .B(b[60]), .Z(n3054) );
  NANDN U5124 ( .A(n3020), .B(n3019), .Z(n3024) );
  NAND U5125 ( .A(n3022), .B(n3021), .Z(n3023) );
  AND U5126 ( .A(n3024), .B(n3023), .Z(n3053) );
  AND U5127 ( .A(a[35]), .B(b[61]), .Z(n3044) );
  AND U5128 ( .A(b[63]), .B(a[33]), .Z(n3050) );
  AND U5129 ( .A(b[62]), .B(a[34]), .Z(n3048) );
  NANDN U5130 ( .A(n3026), .B(n3025), .Z(n3030) );
  NANDN U5131 ( .A(n3028), .B(n3027), .Z(n3029) );
  NAND U5132 ( .A(n3030), .B(n3029), .Z(n3047) );
  NANDN U5133 ( .A(n3032), .B(n3031), .Z(n3036) );
  NAND U5134 ( .A(n3034), .B(n3033), .Z(n3035) );
  NAND U5135 ( .A(n3036), .B(n3035), .Z(n3042) );
  XOR U5136 ( .A(n3056), .B(n3055), .Z(n3336) );
  NAND U5137 ( .A(n3337), .B(n3336), .Z(n3037) );
  NAND U5138 ( .A(n3038), .B(n3037), .Z(n3039) );
  AND U5139 ( .A(a[38]), .B(b[59]), .Z(n3040) );
  NANDN U5140 ( .A(n3039), .B(n3040), .Z(n3060) );
  AND U5141 ( .A(a[36]), .B(b[61]), .Z(n3070) );
  NANDN U5142 ( .A(n3042), .B(n3041), .Z(n3046) );
  NANDN U5143 ( .A(n3044), .B(n3043), .Z(n3045) );
  AND U5144 ( .A(n3046), .B(n3045), .Z(n3068) );
  AND U5145 ( .A(b[63]), .B(a[34]), .Z(n3064) );
  AND U5146 ( .A(b[62]), .B(a[35]), .Z(n3062) );
  NANDN U5147 ( .A(n3048), .B(n3047), .Z(n3052) );
  NANDN U5148 ( .A(n3050), .B(n3049), .Z(n3051) );
  NAND U5149 ( .A(n3052), .B(n3051), .Z(n3061) );
  XOR U5150 ( .A(n3068), .B(n3067), .Z(n3069) );
  XOR U5151 ( .A(n3070), .B(n3069), .Z(n3076) );
  AND U5152 ( .A(a[37]), .B(b[60]), .Z(n3074) );
  NANDN U5153 ( .A(n3054), .B(n3053), .Z(n3058) );
  NAND U5154 ( .A(n3056), .B(n3055), .Z(n3057) );
  NAND U5155 ( .A(n3058), .B(n3057), .Z(n3073) );
  NAND U5156 ( .A(n3344), .B(n3345), .Z(n3059) );
  AND U5157 ( .A(n3060), .B(n3059), .Z(n3079) );
  AND U5158 ( .A(a[39]), .B(b[59]), .Z(n3080) );
  NANDN U5159 ( .A(n3079), .B(n3080), .Z(n3082) );
  AND U5160 ( .A(b[63]), .B(a[35]), .Z(n3094) );
  AND U5161 ( .A(b[62]), .B(a[36]), .Z(n3092) );
  NANDN U5162 ( .A(n3062), .B(n3061), .Z(n3066) );
  NANDN U5163 ( .A(n3064), .B(n3063), .Z(n3065) );
  NAND U5164 ( .A(n3066), .B(n3065), .Z(n3091) );
  NAND U5165 ( .A(n3068), .B(n3067), .Z(n3072) );
  NAND U5166 ( .A(n3070), .B(n3069), .Z(n3071) );
  AND U5167 ( .A(n3072), .B(n3071), .Z(n3098) );
  AND U5168 ( .A(a[37]), .B(b[61]), .Z(n3097) );
  XOR U5169 ( .A(n3099), .B(n3100), .Z(n3088) );
  AND U5170 ( .A(a[38]), .B(b[60]), .Z(n3085) );
  NANDN U5171 ( .A(n3074), .B(n3073), .Z(n3078) );
  NANDN U5172 ( .A(n3076), .B(n3075), .Z(n3077) );
  NAND U5173 ( .A(n3078), .B(n3077), .Z(n3086) );
  XOR U5174 ( .A(n3088), .B(n3087), .Z(n3349) );
  NAND U5175 ( .A(n3349), .B(n3348), .Z(n3081) );
  AND U5176 ( .A(n3082), .B(n3081), .Z(n3084) );
  NANDN U5177 ( .A(n3083), .B(n3084), .Z(n3104) );
  AND U5178 ( .A(a[39]), .B(b[60]), .Z(n3118) );
  NANDN U5179 ( .A(n3086), .B(n3085), .Z(n3090) );
  NAND U5180 ( .A(n3088), .B(n3087), .Z(n3089) );
  AND U5181 ( .A(n3090), .B(n3089), .Z(n3117) );
  AND U5182 ( .A(a[38]), .B(b[61]), .Z(n3114) );
  AND U5183 ( .A(b[63]), .B(a[36]), .Z(n3108) );
  AND U5184 ( .A(b[62]), .B(a[37]), .Z(n3106) );
  NANDN U5185 ( .A(n3092), .B(n3091), .Z(n3096) );
  NANDN U5186 ( .A(n3094), .B(n3093), .Z(n3095) );
  NAND U5187 ( .A(n3096), .B(n3095), .Z(n3105) );
  NANDN U5188 ( .A(n3098), .B(n3097), .Z(n3102) );
  NAND U5189 ( .A(n3100), .B(n3099), .Z(n3101) );
  NAND U5190 ( .A(n3102), .B(n3101), .Z(n3112) );
  XOR U5191 ( .A(n3120), .B(n3119), .Z(n3354) );
  NAND U5192 ( .A(n3355), .B(n3354), .Z(n3103) );
  NAND U5193 ( .A(n3104), .B(n3103), .Z(n10149) );
  AND U5194 ( .A(b[63]), .B(a[37]), .Z(n10139) );
  AND U5195 ( .A(b[62]), .B(a[38]), .Z(n10137) );
  NANDN U5196 ( .A(n3106), .B(n3105), .Z(n3110) );
  NANDN U5197 ( .A(n3108), .B(n3107), .Z(n3109) );
  NAND U5198 ( .A(n3110), .B(n3109), .Z(n10136) );
  NANDN U5199 ( .A(n3112), .B(n3111), .Z(n3116) );
  NANDN U5200 ( .A(n3114), .B(n3113), .Z(n3115) );
  AND U5201 ( .A(n3116), .B(n3115), .Z(n10130) );
  NAND U5202 ( .A(a[39]), .B(b[61]), .Z(n10131) );
  XOR U5203 ( .A(n10132), .B(n10133), .Z(n10145) );
  NANDN U5204 ( .A(n3118), .B(n3117), .Z(n3122) );
  NAND U5205 ( .A(n3120), .B(n3119), .Z(n3121) );
  AND U5206 ( .A(n3122), .B(n3121), .Z(n10142) );
  NAND U5207 ( .A(a[40]), .B(b[60]), .Z(n10143) );
  XOR U5208 ( .A(n10145), .B(n10144), .Z(n10150) );
  XOR U5209 ( .A(n10151), .B(n10150), .Z(n10157) );
  AND U5210 ( .A(a[42]), .B(b[58]), .Z(n10155) );
  AND U5211 ( .A(a[40]), .B(b[58]), .Z(n3350) );
  AND U5212 ( .A(a[39]), .B(b[58]), .Z(n3342) );
  AND U5213 ( .A(a[37]), .B(b[58]), .Z(n3332) );
  AND U5214 ( .A(a[36]), .B(b[58]), .Z(n3324) );
  NAND U5215 ( .A(a[35]), .B(b[58]), .Z(n3320) );
  AND U5216 ( .A(a[34]), .B(b[58]), .Z(n3314) );
  AND U5217 ( .A(a[33]), .B(b[58]), .Z(n3306) );
  AND U5218 ( .A(a[32]), .B(b[58]), .Z(n3301) );
  AND U5219 ( .A(a[31]), .B(b[58]), .Z(n3297) );
  NAND U5220 ( .A(a[28]), .B(b[58]), .Z(n3278) );
  AND U5221 ( .A(a[27]), .B(b[58]), .Z(n3273) );
  AND U5222 ( .A(a[26]), .B(b[58]), .Z(n3265) );
  AND U5223 ( .A(a[25]), .B(b[58]), .Z(n3261) );
  AND U5224 ( .A(a[24]), .B(b[58]), .Z(n3255) );
  AND U5225 ( .A(a[23]), .B(b[58]), .Z(n3249) );
  XNOR U5226 ( .A(n3124), .B(n3123), .Z(n3243) );
  XOR U5227 ( .A(n3126), .B(n3125), .Z(n3239) );
  NAND U5228 ( .A(a[19]), .B(b[58]), .Z(n3228) );
  XNOR U5229 ( .A(n3128), .B(n3127), .Z(n3229) );
  NANDN U5230 ( .A(n3228), .B(n3229), .Z(n3231) );
  AND U5231 ( .A(a[18]), .B(b[58]), .Z(n3224) );
  XOR U5232 ( .A(n3130), .B(n3129), .Z(n3225) );
  NAND U5233 ( .A(n3224), .B(n3225), .Z(n3227) );
  NAND U5234 ( .A(a[17]), .B(b[58]), .Z(n3220) );
  XNOR U5235 ( .A(n3132), .B(n3131), .Z(n3221) );
  NANDN U5236 ( .A(n3220), .B(n3221), .Z(n3223) );
  NAND U5237 ( .A(a[16]), .B(b[58]), .Z(n3216) );
  XOR U5238 ( .A(n3134), .B(n3133), .Z(n3217) );
  NANDN U5239 ( .A(n3216), .B(n3217), .Z(n3219) );
  XOR U5240 ( .A(n3136), .B(n3135), .Z(n3215) );
  XOR U5241 ( .A(n3138), .B(n3137), .Z(n3211) );
  XOR U5242 ( .A(n3140), .B(n3139), .Z(n3142) );
  NAND U5243 ( .A(a[13]), .B(b[58]), .Z(n3141) );
  NANDN U5244 ( .A(n3142), .B(n3141), .Z(n3209) );
  XOR U5245 ( .A(n3142), .B(n3141), .Z(n3374) );
  XOR U5246 ( .A(n3144), .B(n3143), .Z(n3204) );
  XOR U5247 ( .A(n3146), .B(n3145), .Z(n3194) );
  AND U5248 ( .A(a[10]), .B(b[58]), .Z(n3195) );
  NANDN U5249 ( .A(n3194), .B(n3195), .Z(n3197) );
  XOR U5250 ( .A(n3148), .B(n3147), .Z(n3149) );
  AND U5251 ( .A(a[9]), .B(b[58]), .Z(n3150) );
  NANDN U5252 ( .A(n3149), .B(n3150), .Z(n3193) );
  XOR U5253 ( .A(n3150), .B(n3149), .Z(n3382) );
  XOR U5254 ( .A(n3152), .B(n3151), .Z(n3183) );
  XOR U5255 ( .A(n3154), .B(n3153), .Z(n3172) );
  NAND U5256 ( .A(a[0]), .B(b[58]), .Z(n3644) );
  AND U5257 ( .A(a[1]), .B(b[59]), .Z(n3157) );
  NANDN U5258 ( .A(n3644), .B(n3157), .Z(n3392) );
  NANDN U5259 ( .A(n3392), .B(n3155), .Z(n3159) );
  AND U5260 ( .A(a[2]), .B(b[58]), .Z(n3398) );
  NANDN U5261 ( .A(n3397), .B(n3398), .Z(n3158) );
  AND U5262 ( .A(n3159), .B(n3158), .Z(n3162) );
  AND U5263 ( .A(a[3]), .B(b[58]), .Z(n3163) );
  NANDN U5264 ( .A(n3162), .B(n3163), .Z(n3165) );
  XOR U5265 ( .A(n3161), .B(n3160), .Z(n3403) );
  NANDN U5266 ( .A(n3403), .B(n3404), .Z(n3164) );
  AND U5267 ( .A(n3165), .B(n3164), .Z(n3168) );
  XOR U5268 ( .A(n3167), .B(n3166), .Z(n3169) );
  NANDN U5269 ( .A(n3168), .B(n3169), .Z(n3171) );
  AND U5270 ( .A(a[4]), .B(b[58]), .Z(n3391) );
  NAND U5271 ( .A(n3391), .B(n3390), .Z(n3170) );
  AND U5272 ( .A(n3171), .B(n3170), .Z(n3173) );
  NANDN U5273 ( .A(n3172), .B(n3173), .Z(n3175) );
  AND U5274 ( .A(a[5]), .B(b[58]), .Z(n3388) );
  NANDN U5275 ( .A(n3388), .B(n3389), .Z(n3174) );
  AND U5276 ( .A(n3175), .B(n3174), .Z(n3179) );
  NAND U5277 ( .A(n3179), .B(n3178), .Z(n3181) );
  AND U5278 ( .A(a[6]), .B(b[58]), .Z(n3387) );
  XOR U5279 ( .A(n3179), .B(n3178), .Z(n3386) );
  NAND U5280 ( .A(n3387), .B(n3386), .Z(n3180) );
  NAND U5281 ( .A(n3181), .B(n3180), .Z(n3182) );
  NANDN U5282 ( .A(n3183), .B(n3182), .Z(n3185) );
  NAND U5283 ( .A(a[7]), .B(b[58]), .Z(n3384) );
  XNOR U5284 ( .A(n3183), .B(n3182), .Z(n3385) );
  NANDN U5285 ( .A(n3384), .B(n3385), .Z(n3184) );
  AND U5286 ( .A(n3185), .B(n3184), .Z(n3189) );
  XNOR U5287 ( .A(n3187), .B(n3186), .Z(n3188) );
  NANDN U5288 ( .A(n3189), .B(n3188), .Z(n3191) );
  NAND U5289 ( .A(a[8]), .B(b[58]), .Z(n3425) );
  XNOR U5290 ( .A(n3189), .B(n3188), .Z(n3426) );
  NANDN U5291 ( .A(n3425), .B(n3426), .Z(n3190) );
  AND U5292 ( .A(n3191), .B(n3190), .Z(n3383) );
  OR U5293 ( .A(n3382), .B(n3383), .Z(n3192) );
  AND U5294 ( .A(n3193), .B(n3192), .Z(n3436) );
  XNOR U5295 ( .A(n3195), .B(n3194), .Z(n3435) );
  NANDN U5296 ( .A(n3436), .B(n3435), .Z(n3196) );
  AND U5297 ( .A(n3197), .B(n3196), .Z(n3201) );
  XNOR U5298 ( .A(n3199), .B(n3198), .Z(n3200) );
  NANDN U5299 ( .A(n3201), .B(n3200), .Z(n3203) );
  NAND U5300 ( .A(a[11]), .B(b[58]), .Z(n3380) );
  XNOR U5301 ( .A(n3201), .B(n3200), .Z(n3381) );
  NANDN U5302 ( .A(n3380), .B(n3381), .Z(n3202) );
  AND U5303 ( .A(n3203), .B(n3202), .Z(n3205) );
  NANDN U5304 ( .A(n3204), .B(n3205), .Z(n3207) );
  XOR U5305 ( .A(n3205), .B(n3204), .Z(n3378) );
  AND U5306 ( .A(a[12]), .B(b[58]), .Z(n3379) );
  OR U5307 ( .A(n3378), .B(n3379), .Z(n3206) );
  AND U5308 ( .A(n3207), .B(n3206), .Z(n3375) );
  OR U5309 ( .A(n3374), .B(n3375), .Z(n3208) );
  NAND U5310 ( .A(n3209), .B(n3208), .Z(n3210) );
  NANDN U5311 ( .A(n3211), .B(n3210), .Z(n3213) );
  XOR U5312 ( .A(n3211), .B(n3210), .Z(n3372) );
  AND U5313 ( .A(a[14]), .B(b[58]), .Z(n3373) );
  OR U5314 ( .A(n3372), .B(n3373), .Z(n3212) );
  NAND U5315 ( .A(n3213), .B(n3212), .Z(n3214) );
  AND U5316 ( .A(a[15]), .B(b[58]), .Z(n3371) );
  XOR U5317 ( .A(n3215), .B(n3214), .Z(n3370) );
  XNOR U5318 ( .A(n3217), .B(n3216), .Z(n3369) );
  NANDN U5319 ( .A(n3368), .B(n3369), .Z(n3218) );
  AND U5320 ( .A(n3219), .B(n3218), .Z(n3462) );
  XNOR U5321 ( .A(n3221), .B(n3220), .Z(n3461) );
  NANDN U5322 ( .A(n3462), .B(n3461), .Z(n3222) );
  AND U5323 ( .A(n3223), .B(n3222), .Z(n3367) );
  XOR U5324 ( .A(n3225), .B(n3224), .Z(n3366) );
  NANDN U5325 ( .A(n3367), .B(n3366), .Z(n3226) );
  AND U5326 ( .A(n3227), .B(n3226), .Z(n3472) );
  XNOR U5327 ( .A(n3229), .B(n3228), .Z(n3471) );
  NANDN U5328 ( .A(n3472), .B(n3471), .Z(n3230) );
  AND U5329 ( .A(n3231), .B(n3230), .Z(n3235) );
  XNOR U5330 ( .A(n3233), .B(n3232), .Z(n3234) );
  NANDN U5331 ( .A(n3235), .B(n3234), .Z(n3237) );
  NAND U5332 ( .A(a[20]), .B(b[58]), .Z(n3475) );
  XNOR U5333 ( .A(n3235), .B(n3234), .Z(n3476) );
  NANDN U5334 ( .A(n3475), .B(n3476), .Z(n3236) );
  AND U5335 ( .A(n3237), .B(n3236), .Z(n3238) );
  NANDN U5336 ( .A(n3239), .B(n3238), .Z(n3241) );
  AND U5337 ( .A(a[21]), .B(b[58]), .Z(n3365) );
  XNOR U5338 ( .A(n3239), .B(n3238), .Z(n3364) );
  NANDN U5339 ( .A(n3365), .B(n3364), .Z(n3240) );
  NAND U5340 ( .A(n3241), .B(n3240), .Z(n3242) );
  NAND U5341 ( .A(n3243), .B(n3242), .Z(n3245) );
  AND U5342 ( .A(a[22]), .B(b[58]), .Z(n3363) );
  XOR U5343 ( .A(n3243), .B(n3242), .Z(n3362) );
  NANDN U5344 ( .A(n3363), .B(n3362), .Z(n3244) );
  NAND U5345 ( .A(n3245), .B(n3244), .Z(n3248) );
  NANDN U5346 ( .A(n3249), .B(n3248), .Z(n3251) );
  XOR U5347 ( .A(n3247), .B(n3246), .Z(n3361) );
  XNOR U5348 ( .A(n3249), .B(n3248), .Z(n3360) );
  NANDN U5349 ( .A(n3361), .B(n3360), .Z(n3250) );
  NAND U5350 ( .A(n3251), .B(n3250), .Z(n3254) );
  NANDN U5351 ( .A(n3255), .B(n3254), .Z(n3257) );
  XOR U5352 ( .A(n3253), .B(n3252), .Z(n3496) );
  XNOR U5353 ( .A(n3255), .B(n3254), .Z(n3495) );
  NANDN U5354 ( .A(n3496), .B(n3495), .Z(n3256) );
  NAND U5355 ( .A(n3257), .B(n3256), .Z(n3260) );
  NANDN U5356 ( .A(n3261), .B(n3260), .Z(n3263) );
  XOR U5357 ( .A(n3259), .B(n3258), .Z(n3502) );
  XNOR U5358 ( .A(n3261), .B(n3260), .Z(n3501) );
  NANDN U5359 ( .A(n3502), .B(n3501), .Z(n3262) );
  NAND U5360 ( .A(n3263), .B(n3262), .Z(n3264) );
  NANDN U5361 ( .A(n3265), .B(n3264), .Z(n3269) );
  XNOR U5362 ( .A(n3265), .B(n3264), .Z(n3507) );
  XOR U5363 ( .A(n3267), .B(n3266), .Z(n3508) );
  NAND U5364 ( .A(n3507), .B(n3508), .Z(n3268) );
  NAND U5365 ( .A(n3269), .B(n3268), .Z(n3272) );
  NANDN U5366 ( .A(n3273), .B(n3272), .Z(n3275) );
  XOR U5367 ( .A(n3271), .B(n3270), .Z(n3514) );
  XNOR U5368 ( .A(n3273), .B(n3272), .Z(n3513) );
  NANDN U5369 ( .A(n3514), .B(n3513), .Z(n3274) );
  AND U5370 ( .A(n3275), .B(n3274), .Z(n3279) );
  NANDN U5371 ( .A(n3278), .B(n3279), .Z(n3281) );
  XOR U5372 ( .A(n3277), .B(n3276), .Z(n3520) );
  XNOR U5373 ( .A(n3279), .B(n3278), .Z(n3519) );
  NAND U5374 ( .A(n3520), .B(n3519), .Z(n3280) );
  AND U5375 ( .A(n3281), .B(n3280), .Z(n3285) );
  AND U5376 ( .A(a[29]), .B(b[58]), .Z(n3284) );
  NANDN U5377 ( .A(n3285), .B(n3284), .Z(n3287) );
  XOR U5378 ( .A(n3283), .B(n3282), .Z(n3524) );
  XNOR U5379 ( .A(n3285), .B(n3284), .Z(n3523) );
  NAND U5380 ( .A(n3524), .B(n3523), .Z(n3286) );
  AND U5381 ( .A(n3287), .B(n3286), .Z(n3291) );
  AND U5382 ( .A(a[30]), .B(b[58]), .Z(n3290) );
  NANDN U5383 ( .A(n3291), .B(n3290), .Z(n3293) );
  XOR U5384 ( .A(n3289), .B(n3288), .Z(n3530) );
  XNOR U5385 ( .A(n3291), .B(n3290), .Z(n3529) );
  NAND U5386 ( .A(n3530), .B(n3529), .Z(n3292) );
  AND U5387 ( .A(n3293), .B(n3292), .Z(n3296) );
  NANDN U5388 ( .A(n3297), .B(n3296), .Z(n3299) );
  XOR U5389 ( .A(n3295), .B(n3294), .Z(n3538) );
  XNOR U5390 ( .A(n3297), .B(n3296), .Z(n3537) );
  NANDN U5391 ( .A(n3538), .B(n3537), .Z(n3298) );
  NAND U5392 ( .A(n3299), .B(n3298), .Z(n3300) );
  NANDN U5393 ( .A(n3301), .B(n3300), .Z(n3305) );
  XNOR U5394 ( .A(n3301), .B(n3300), .Z(n3542) );
  XOR U5395 ( .A(n3303), .B(n3302), .Z(n3541) );
  NAND U5396 ( .A(n3542), .B(n3541), .Z(n3304) );
  NAND U5397 ( .A(n3305), .B(n3304), .Z(n3307) );
  NANDN U5398 ( .A(n3306), .B(n3307), .Z(n3311) );
  XNOR U5399 ( .A(n3309), .B(n3308), .Z(n3550) );
  NAND U5400 ( .A(n3549), .B(n3550), .Z(n3310) );
  NAND U5401 ( .A(n3311), .B(n3310), .Z(n3315) );
  NANDN U5402 ( .A(n3314), .B(n3315), .Z(n3317) );
  XOR U5403 ( .A(n3313), .B(n3312), .Z(n3555) );
  NANDN U5404 ( .A(n3555), .B(n3556), .Z(n3316) );
  AND U5405 ( .A(n3317), .B(n3316), .Z(n3321) );
  NANDN U5406 ( .A(n3320), .B(n3321), .Z(n3323) );
  XOR U5407 ( .A(n3319), .B(n3318), .Z(n3561) );
  NANDN U5408 ( .A(n3561), .B(n3562), .Z(n3322) );
  AND U5409 ( .A(n3323), .B(n3322), .Z(n3325) );
  NANDN U5410 ( .A(n3324), .B(n3325), .Z(n3329) );
  NAND U5411 ( .A(n3567), .B(n3568), .Z(n3328) );
  NAND U5412 ( .A(n3329), .B(n3328), .Z(n3333) );
  NANDN U5413 ( .A(n3332), .B(n3333), .Z(n3335) );
  XOR U5414 ( .A(n3331), .B(n3330), .Z(n3573) );
  NANDN U5415 ( .A(n3573), .B(n3574), .Z(n3334) );
  NAND U5416 ( .A(n3335), .B(n3334), .Z(n3338) );
  AND U5417 ( .A(a[38]), .B(b[58]), .Z(n3339) );
  NANDN U5418 ( .A(n3338), .B(n3339), .Z(n3341) );
  XOR U5419 ( .A(n3337), .B(n3336), .Z(n3579) );
  NANDN U5420 ( .A(n3579), .B(n3580), .Z(n3340) );
  AND U5421 ( .A(n3341), .B(n3340), .Z(n3343) );
  NANDN U5422 ( .A(n3342), .B(n3343), .Z(n3347) );
  XNOR U5423 ( .A(n3345), .B(n3344), .Z(n3586) );
  NAND U5424 ( .A(n3585), .B(n3586), .Z(n3346) );
  NAND U5425 ( .A(n3347), .B(n3346), .Z(n3351) );
  NANDN U5426 ( .A(n3350), .B(n3351), .Z(n3353) );
  XOR U5427 ( .A(n3349), .B(n3348), .Z(n3591) );
  NANDN U5428 ( .A(n3591), .B(n3592), .Z(n3352) );
  NAND U5429 ( .A(n3353), .B(n3352), .Z(n3356) );
  AND U5430 ( .A(a[41]), .B(b[58]), .Z(n3357) );
  NANDN U5431 ( .A(n3356), .B(n3357), .Z(n3359) );
  XOR U5432 ( .A(n3355), .B(n3354), .Z(n3597) );
  NANDN U5433 ( .A(n3597), .B(n3598), .Z(n3358) );
  AND U5434 ( .A(n3359), .B(n3358), .Z(n10154) );
  AND U5435 ( .A(a[43]), .B(b[57]), .Z(n10160) );
  NAND U5436 ( .A(a[33]), .B(b[57]), .Z(n3543) );
  AND U5437 ( .A(a[32]), .B(b[57]), .Z(n3536) );
  AND U5438 ( .A(a[31]), .B(b[57]), .Z(n3532) );
  AND U5439 ( .A(a[30]), .B(b[57]), .Z(n3526) );
  XOR U5440 ( .A(n3361), .B(n3360), .Z(n3490) );
  AND U5441 ( .A(a[23]), .B(b[57]), .Z(n3485) );
  XOR U5442 ( .A(n3363), .B(n3362), .Z(n3486) );
  NAND U5443 ( .A(n3485), .B(n3486), .Z(n3488) );
  XOR U5444 ( .A(n3365), .B(n3364), .Z(n3482) );
  NAND U5445 ( .A(a[20]), .B(b[57]), .Z(n3473) );
  AND U5446 ( .A(a[19]), .B(b[57]), .Z(n3468) );
  XOR U5447 ( .A(n3367), .B(n3366), .Z(n3467) );
  NANDN U5448 ( .A(n3468), .B(n3467), .Z(n3470) );
  XOR U5449 ( .A(n3369), .B(n3368), .Z(n3457) );
  AND U5450 ( .A(a[17]), .B(b[57]), .Z(n3458) );
  NANDN U5451 ( .A(n3457), .B(n3458), .Z(n3460) );
  XOR U5452 ( .A(n3371), .B(n3370), .Z(n3456) );
  XOR U5453 ( .A(n3373), .B(n3372), .Z(n3452) );
  XOR U5454 ( .A(n3375), .B(n3374), .Z(n3377) );
  AND U5455 ( .A(a[14]), .B(b[57]), .Z(n3376) );
  NANDN U5456 ( .A(n3377), .B(n3376), .Z(n3450) );
  XOR U5457 ( .A(n3377), .B(n3376), .Z(n3623) );
  XOR U5458 ( .A(n3379), .B(n3378), .Z(n3446) );
  NAND U5459 ( .A(a[12]), .B(b[57]), .Z(n3441) );
  XNOR U5460 ( .A(n3381), .B(n3380), .Z(n3442) );
  NANDN U5461 ( .A(n3441), .B(n3442), .Z(n3444) );
  XOR U5462 ( .A(n3383), .B(n3382), .Z(n3432) );
  XOR U5463 ( .A(n3385), .B(n3384), .Z(n3421) );
  AND U5464 ( .A(a[8]), .B(b[57]), .Z(n3422) );
  NANDN U5465 ( .A(n3421), .B(n3422), .Z(n3424) );
  NAND U5466 ( .A(a[7]), .B(b[57]), .Z(n3417) );
  XOR U5467 ( .A(n3387), .B(n3386), .Z(n3418) );
  NANDN U5468 ( .A(n3417), .B(n3418), .Z(n3420) );
  AND U5469 ( .A(a[6]), .B(b[57]), .Z(n3413) );
  NAND U5470 ( .A(n3413), .B(n3414), .Z(n3416) );
  XOR U5471 ( .A(n3391), .B(n3390), .Z(n3409) );
  NAND U5472 ( .A(a[0]), .B(b[57]), .Z(n3885) );
  AND U5473 ( .A(a[1]), .B(b[58]), .Z(n3394) );
  NANDN U5474 ( .A(n3885), .B(n3394), .Z(n3643) );
  NANDN U5475 ( .A(n3643), .B(n3392), .Z(n3396) );
  AND U5476 ( .A(a[2]), .B(b[57]), .Z(n3649) );
  NANDN U5477 ( .A(n3648), .B(n3649), .Z(n3395) );
  AND U5478 ( .A(n3396), .B(n3395), .Z(n3399) );
  XNOR U5479 ( .A(n3398), .B(n3397), .Z(n3400) );
  NANDN U5480 ( .A(n3399), .B(n3400), .Z(n3402) );
  AND U5481 ( .A(a[3]), .B(b[57]), .Z(n3655) );
  NAND U5482 ( .A(n3655), .B(n3654), .Z(n3401) );
  AND U5483 ( .A(n3402), .B(n3401), .Z(n3405) );
  NANDN U5484 ( .A(n3405), .B(n3406), .Z(n3408) );
  NAND U5485 ( .A(a[4]), .B(b[57]), .Z(n3660) );
  NANDN U5486 ( .A(n3660), .B(n3661), .Z(n3407) );
  AND U5487 ( .A(n3408), .B(n3407), .Z(n3410) );
  NANDN U5488 ( .A(n3409), .B(n3410), .Z(n3412) );
  AND U5489 ( .A(a[5]), .B(b[57]), .Z(n3667) );
  NANDN U5490 ( .A(n3667), .B(n3666), .Z(n3411) );
  NAND U5491 ( .A(n3412), .B(n3411), .Z(n3641) );
  XOR U5492 ( .A(n3414), .B(n3413), .Z(n3642) );
  NANDN U5493 ( .A(n3641), .B(n3642), .Z(n3415) );
  AND U5494 ( .A(n3416), .B(n3415), .Z(n3676) );
  NANDN U5495 ( .A(n3676), .B(n3677), .Z(n3419) );
  AND U5496 ( .A(n3420), .B(n3419), .Z(n3683) );
  XNOR U5497 ( .A(n3422), .B(n3421), .Z(n3682) );
  NANDN U5498 ( .A(n3683), .B(n3682), .Z(n3423) );
  AND U5499 ( .A(n3424), .B(n3423), .Z(n3428) );
  XNOR U5500 ( .A(n3426), .B(n3425), .Z(n3427) );
  NANDN U5501 ( .A(n3428), .B(n3427), .Z(n3430) );
  NAND U5502 ( .A(a[9]), .B(b[57]), .Z(n3639) );
  XNOR U5503 ( .A(n3428), .B(n3427), .Z(n3640) );
  NANDN U5504 ( .A(n3639), .B(n3640), .Z(n3429) );
  AND U5505 ( .A(n3430), .B(n3429), .Z(n3431) );
  NANDN U5506 ( .A(n3432), .B(n3431), .Z(n3434) );
  XOR U5507 ( .A(n3432), .B(n3431), .Z(n3635) );
  AND U5508 ( .A(a[10]), .B(b[57]), .Z(n3636) );
  OR U5509 ( .A(n3635), .B(n3636), .Z(n3433) );
  NAND U5510 ( .A(n3434), .B(n3433), .Z(n3437) );
  XNOR U5511 ( .A(n3436), .B(n3435), .Z(n3438) );
  NANDN U5512 ( .A(n3437), .B(n3438), .Z(n3440) );
  NAND U5513 ( .A(a[11]), .B(b[57]), .Z(n3633) );
  XNOR U5514 ( .A(n3438), .B(n3437), .Z(n3634) );
  NANDN U5515 ( .A(n3633), .B(n3634), .Z(n3439) );
  AND U5516 ( .A(n3440), .B(n3439), .Z(n3630) );
  XNOR U5517 ( .A(n3442), .B(n3441), .Z(n3629) );
  NANDN U5518 ( .A(n3630), .B(n3629), .Z(n3443) );
  NAND U5519 ( .A(n3444), .B(n3443), .Z(n3445) );
  NANDN U5520 ( .A(n3446), .B(n3445), .Z(n3448) );
  NAND U5521 ( .A(a[13]), .B(b[57]), .Z(n3625) );
  XNOR U5522 ( .A(n3446), .B(n3445), .Z(n3626) );
  NANDN U5523 ( .A(n3625), .B(n3626), .Z(n3447) );
  AND U5524 ( .A(n3448), .B(n3447), .Z(n3624) );
  OR U5525 ( .A(n3623), .B(n3624), .Z(n3449) );
  NAND U5526 ( .A(n3450), .B(n3449), .Z(n3451) );
  NANDN U5527 ( .A(n3452), .B(n3451), .Z(n3454) );
  XNOR U5528 ( .A(n3452), .B(n3451), .Z(n3622) );
  AND U5529 ( .A(a[15]), .B(b[57]), .Z(n3621) );
  NAND U5530 ( .A(n3622), .B(n3621), .Z(n3453) );
  NAND U5531 ( .A(n3454), .B(n3453), .Z(n3455) );
  NAND U5532 ( .A(a[16]), .B(b[57]), .Z(n3619) );
  XOR U5533 ( .A(n3456), .B(n3455), .Z(n3620) );
  XNOR U5534 ( .A(n3458), .B(n3457), .Z(n3615) );
  NANDN U5535 ( .A(n3616), .B(n3615), .Z(n3459) );
  AND U5536 ( .A(n3460), .B(n3459), .Z(n3464) );
  XNOR U5537 ( .A(n3462), .B(n3461), .Z(n3463) );
  NANDN U5538 ( .A(n3464), .B(n3463), .Z(n3466) );
  XNOR U5539 ( .A(n3464), .B(n3463), .Z(n3614) );
  AND U5540 ( .A(a[18]), .B(b[57]), .Z(n3613) );
  NAND U5541 ( .A(n3614), .B(n3613), .Z(n3465) );
  AND U5542 ( .A(n3466), .B(n3465), .Z(n3612) );
  XNOR U5543 ( .A(n3468), .B(n3467), .Z(n3611) );
  NAND U5544 ( .A(n3612), .B(n3611), .Z(n3469) );
  AND U5545 ( .A(n3470), .B(n3469), .Z(n3474) );
  XNOR U5546 ( .A(n3472), .B(n3471), .Z(n3607) );
  XNOR U5547 ( .A(n3474), .B(n3473), .Z(n3608) );
  XNOR U5548 ( .A(n3476), .B(n3475), .Z(n3477) );
  NANDN U5549 ( .A(n3478), .B(n3477), .Z(n3480) );
  NAND U5550 ( .A(a[21]), .B(b[57]), .Z(n3605) );
  XNOR U5551 ( .A(n3478), .B(n3477), .Z(n3606) );
  NANDN U5552 ( .A(n3605), .B(n3606), .Z(n3479) );
  NAND U5553 ( .A(n3480), .B(n3479), .Z(n3481) );
  NAND U5554 ( .A(n3482), .B(n3481), .Z(n3484) );
  NAND U5555 ( .A(a[22]), .B(b[57]), .Z(n3730) );
  XOR U5556 ( .A(n3482), .B(n3481), .Z(n3731) );
  NANDN U5557 ( .A(n3730), .B(n3731), .Z(n3483) );
  AND U5558 ( .A(n3484), .B(n3483), .Z(n3737) );
  XOR U5559 ( .A(n3486), .B(n3485), .Z(n3736) );
  NANDN U5560 ( .A(n3737), .B(n3736), .Z(n3487) );
  NAND U5561 ( .A(n3488), .B(n3487), .Z(n3489) );
  NAND U5562 ( .A(n3490), .B(n3489), .Z(n3492) );
  NAND U5563 ( .A(a[24]), .B(b[57]), .Z(n3603) );
  XOR U5564 ( .A(n3490), .B(n3489), .Z(n3604) );
  NANDN U5565 ( .A(n3603), .B(n3604), .Z(n3491) );
  AND U5566 ( .A(n3492), .B(n3491), .Z(n3494) );
  AND U5567 ( .A(a[25]), .B(b[57]), .Z(n3493) );
  NANDN U5568 ( .A(n3494), .B(n3493), .Z(n3498) );
  XNOR U5569 ( .A(n3494), .B(n3493), .Z(n3601) );
  XOR U5570 ( .A(n3496), .B(n3495), .Z(n3602) );
  NAND U5571 ( .A(n3601), .B(n3602), .Z(n3497) );
  AND U5572 ( .A(n3498), .B(n3497), .Z(n3500) );
  AND U5573 ( .A(a[26]), .B(b[57]), .Z(n3499) );
  NANDN U5574 ( .A(n3500), .B(n3499), .Z(n3504) );
  XNOR U5575 ( .A(n3500), .B(n3499), .Z(n3752) );
  XOR U5576 ( .A(n3502), .B(n3501), .Z(n3753) );
  NAND U5577 ( .A(n3752), .B(n3753), .Z(n3503) );
  AND U5578 ( .A(n3504), .B(n3503), .Z(n3506) );
  AND U5579 ( .A(a[27]), .B(b[57]), .Z(n3505) );
  NANDN U5580 ( .A(n3506), .B(n3505), .Z(n3510) );
  XNOR U5581 ( .A(n3506), .B(n3505), .Z(n3758) );
  XNOR U5582 ( .A(n3508), .B(n3507), .Z(n3759) );
  NAND U5583 ( .A(n3758), .B(n3759), .Z(n3509) );
  AND U5584 ( .A(n3510), .B(n3509), .Z(n3512) );
  AND U5585 ( .A(a[28]), .B(b[57]), .Z(n3511) );
  NANDN U5586 ( .A(n3512), .B(n3511), .Z(n3516) );
  XNOR U5587 ( .A(n3512), .B(n3511), .Z(n3764) );
  XOR U5588 ( .A(n3514), .B(n3513), .Z(n3765) );
  NAND U5589 ( .A(n3764), .B(n3765), .Z(n3515) );
  AND U5590 ( .A(n3516), .B(n3515), .Z(n3518) );
  AND U5591 ( .A(a[29]), .B(b[57]), .Z(n3517) );
  NANDN U5592 ( .A(n3518), .B(n3517), .Z(n3522) );
  XNOR U5593 ( .A(n3518), .B(n3517), .Z(n3769) );
  XOR U5594 ( .A(n3520), .B(n3519), .Z(n3768) );
  NAND U5595 ( .A(n3769), .B(n3768), .Z(n3521) );
  AND U5596 ( .A(n3522), .B(n3521), .Z(n3525) );
  NANDN U5597 ( .A(n3526), .B(n3525), .Z(n3528) );
  XOR U5598 ( .A(n3524), .B(n3523), .Z(n3777) );
  XNOR U5599 ( .A(n3526), .B(n3525), .Z(n3776) );
  NANDN U5600 ( .A(n3777), .B(n3776), .Z(n3527) );
  NAND U5601 ( .A(n3528), .B(n3527), .Z(n3531) );
  NANDN U5602 ( .A(n3532), .B(n3531), .Z(n3534) );
  XOR U5603 ( .A(n3530), .B(n3529), .Z(n3783) );
  XNOR U5604 ( .A(n3532), .B(n3531), .Z(n3782) );
  NANDN U5605 ( .A(n3783), .B(n3782), .Z(n3533) );
  NAND U5606 ( .A(n3534), .B(n3533), .Z(n3535) );
  NANDN U5607 ( .A(n3536), .B(n3535), .Z(n3540) );
  XNOR U5608 ( .A(n3536), .B(n3535), .Z(n3787) );
  XNOR U5609 ( .A(n3538), .B(n3537), .Z(n3786) );
  NAND U5610 ( .A(n3787), .B(n3786), .Z(n3539) );
  AND U5611 ( .A(n3540), .B(n3539), .Z(n3544) );
  NANDN U5612 ( .A(n3543), .B(n3544), .Z(n3546) );
  XOR U5613 ( .A(n3542), .B(n3541), .Z(n3795) );
  XNOR U5614 ( .A(n3544), .B(n3543), .Z(n3794) );
  NANDN U5615 ( .A(n3795), .B(n3794), .Z(n3545) );
  AND U5616 ( .A(n3546), .B(n3545), .Z(n3547) );
  AND U5617 ( .A(a[34]), .B(b[57]), .Z(n3548) );
  NANDN U5618 ( .A(n3547), .B(n3548), .Z(n3552) );
  XNOR U5619 ( .A(n3550), .B(n3549), .Z(n3801) );
  NAND U5620 ( .A(n3800), .B(n3801), .Z(n3551) );
  AND U5621 ( .A(n3552), .B(n3551), .Z(n3553) );
  AND U5622 ( .A(a[35]), .B(b[57]), .Z(n3554) );
  NANDN U5623 ( .A(n3553), .B(n3554), .Z(n3558) );
  NAND U5624 ( .A(n3804), .B(n3805), .Z(n3557) );
  AND U5625 ( .A(n3558), .B(n3557), .Z(n3559) );
  AND U5626 ( .A(a[36]), .B(b[57]), .Z(n3560) );
  NANDN U5627 ( .A(n3559), .B(n3560), .Z(n3564) );
  NAND U5628 ( .A(n3811), .B(n3810), .Z(n3563) );
  AND U5629 ( .A(n3564), .B(n3563), .Z(n3565) );
  AND U5630 ( .A(a[37]), .B(b[57]), .Z(n3566) );
  NANDN U5631 ( .A(n3565), .B(n3566), .Z(n3570) );
  XNOR U5632 ( .A(n3568), .B(n3567), .Z(n3819) );
  NAND U5633 ( .A(n3818), .B(n3819), .Z(n3569) );
  AND U5634 ( .A(n3570), .B(n3569), .Z(n3571) );
  AND U5635 ( .A(a[38]), .B(b[57]), .Z(n3572) );
  NANDN U5636 ( .A(n3571), .B(n3572), .Z(n3576) );
  NAND U5637 ( .A(n3824), .B(n3825), .Z(n3575) );
  AND U5638 ( .A(n3576), .B(n3575), .Z(n3577) );
  AND U5639 ( .A(a[39]), .B(b[57]), .Z(n3578) );
  NANDN U5640 ( .A(n3577), .B(n3578), .Z(n3582) );
  NAND U5641 ( .A(n3829), .B(n3828), .Z(n3581) );
  AND U5642 ( .A(n3582), .B(n3581), .Z(n3583) );
  AND U5643 ( .A(a[40]), .B(b[57]), .Z(n3584) );
  NANDN U5644 ( .A(n3583), .B(n3584), .Z(n3588) );
  XNOR U5645 ( .A(n3586), .B(n3585), .Z(n3837) );
  NAND U5646 ( .A(n3836), .B(n3837), .Z(n3587) );
  AND U5647 ( .A(n3588), .B(n3587), .Z(n3589) );
  AND U5648 ( .A(a[41]), .B(b[57]), .Z(n3590) );
  NANDN U5649 ( .A(n3589), .B(n3590), .Z(n3594) );
  NAND U5650 ( .A(n3840), .B(n3841), .Z(n3593) );
  AND U5651 ( .A(n3594), .B(n3593), .Z(n3595) );
  AND U5652 ( .A(a[42]), .B(b[57]), .Z(n3596) );
  NANDN U5653 ( .A(n3595), .B(n3596), .Z(n3600) );
  NAND U5654 ( .A(n3847), .B(n3846), .Z(n3599) );
  AND U5655 ( .A(n3600), .B(n3599), .Z(n10161) );
  XNOR U5656 ( .A(n10162), .B(n10163), .Z(n10168) );
  AND U5657 ( .A(a[44]), .B(b[56]), .Z(n10167) );
  AND U5658 ( .A(a[43]), .B(b[56]), .Z(n3848) );
  AND U5659 ( .A(a[41]), .B(b[56]), .Z(n3834) );
  AND U5660 ( .A(a[40]), .B(b[56]), .Z(n3830) );
  AND U5661 ( .A(a[39]), .B(b[56]), .Z(n3822) );
  AND U5662 ( .A(a[38]), .B(b[56]), .Z(n3816) );
  AND U5663 ( .A(a[37]), .B(b[56]), .Z(n3812) );
  NAND U5664 ( .A(a[36]), .B(b[56]), .Z(n3806) );
  AND U5665 ( .A(a[35]), .B(b[56]), .Z(n3798) );
  AND U5666 ( .A(a[34]), .B(b[56]), .Z(n3793) );
  NAND U5667 ( .A(a[33]), .B(b[56]), .Z(n3788) );
  AND U5668 ( .A(a[32]), .B(b[56]), .Z(n3781) );
  AND U5669 ( .A(a[31]), .B(b[56]), .Z(n3775) );
  AND U5670 ( .A(a[30]), .B(b[56]), .Z(n3771) );
  AND U5671 ( .A(a[29]), .B(b[56]), .Z(n3763) );
  AND U5672 ( .A(a[28]), .B(b[56]), .Z(n3757) );
  AND U5673 ( .A(a[27]), .B(b[56]), .Z(n3751) );
  NAND U5674 ( .A(a[26]), .B(b[56]), .Z(n3746) );
  XOR U5675 ( .A(n3602), .B(n3601), .Z(n3747) );
  NANDN U5676 ( .A(n3746), .B(n3747), .Z(n3749) );
  NAND U5677 ( .A(a[25]), .B(b[56]), .Z(n3742) );
  XNOR U5678 ( .A(n3604), .B(n3603), .Z(n3743) );
  NANDN U5679 ( .A(n3742), .B(n3743), .Z(n3745) );
  NAND U5680 ( .A(a[22]), .B(b[56]), .Z(n3726) );
  XNOR U5681 ( .A(n3606), .B(n3605), .Z(n3727) );
  NANDN U5682 ( .A(n3726), .B(n3727), .Z(n3729) );
  NAND U5683 ( .A(a[21]), .B(b[56]), .Z(n3609) );
  XOR U5684 ( .A(n3608), .B(n3607), .Z(n3610) );
  NANDN U5685 ( .A(n3609), .B(n3610), .Z(n3725) );
  XOR U5686 ( .A(n3610), .B(n3609), .Z(n3858) );
  XOR U5687 ( .A(n3612), .B(n3611), .Z(n3721) );
  XOR U5688 ( .A(n3614), .B(n3613), .Z(n3717) );
  NAND U5689 ( .A(a[18]), .B(b[56]), .Z(n3617) );
  XNOR U5690 ( .A(n3616), .B(n3615), .Z(n3618) );
  NANDN U5691 ( .A(n3617), .B(n3618), .Z(n3715) );
  XOR U5692 ( .A(n3618), .B(n3617), .Z(n3862) );
  NAND U5693 ( .A(a[17]), .B(b[56]), .Z(n3710) );
  XNOR U5694 ( .A(n3620), .B(n3619), .Z(n3711) );
  NANDN U5695 ( .A(n3710), .B(n3711), .Z(n3713) );
  XOR U5696 ( .A(n3622), .B(n3621), .Z(n3707) );
  XOR U5697 ( .A(n3624), .B(n3623), .Z(n3703) );
  XOR U5698 ( .A(n3626), .B(n3625), .Z(n3627) );
  AND U5699 ( .A(a[14]), .B(b[56]), .Z(n3628) );
  NANDN U5700 ( .A(n3627), .B(n3628), .Z(n3701) );
  XOR U5701 ( .A(n3628), .B(n3627), .Z(n3870) );
  NAND U5702 ( .A(a[13]), .B(b[56]), .Z(n3631) );
  XNOR U5703 ( .A(n3630), .B(n3629), .Z(n3632) );
  NANDN U5704 ( .A(n3631), .B(n3632), .Z(n3699) );
  XOR U5705 ( .A(n3632), .B(n3631), .Z(n3872) );
  NAND U5706 ( .A(a[12]), .B(b[56]), .Z(n3694) );
  XNOR U5707 ( .A(n3634), .B(n3633), .Z(n3695) );
  NANDN U5708 ( .A(n3694), .B(n3695), .Z(n3697) );
  XOR U5709 ( .A(n3636), .B(n3635), .Z(n3638) );
  AND U5710 ( .A(a[11]), .B(b[56]), .Z(n3637) );
  NANDN U5711 ( .A(n3638), .B(n3637), .Z(n3693) );
  XOR U5712 ( .A(n3638), .B(n3637), .Z(n3876) );
  XOR U5713 ( .A(n3640), .B(n3639), .Z(n3688) );
  AND U5714 ( .A(a[10]), .B(b[56]), .Z(n3689) );
  NANDN U5715 ( .A(n3688), .B(n3689), .Z(n3691) );
  NAND U5716 ( .A(a[7]), .B(b[56]), .Z(n3672) );
  NANDN U5717 ( .A(n3672), .B(n3673), .Z(n3675) );
  NAND U5718 ( .A(a[0]), .B(b[56]), .Z(n4148) );
  AND U5719 ( .A(a[1]), .B(b[57]), .Z(n3645) );
  NANDN U5720 ( .A(n4148), .B(n3645), .Z(n3884) );
  NANDN U5721 ( .A(n3884), .B(n3643), .Z(n3647) );
  AND U5722 ( .A(a[2]), .B(b[56]), .Z(n3890) );
  NANDN U5723 ( .A(n3889), .B(n3890), .Z(n3646) );
  AND U5724 ( .A(n3647), .B(n3646), .Z(n3650) );
  AND U5725 ( .A(a[3]), .B(b[56]), .Z(n3651) );
  NANDN U5726 ( .A(n3650), .B(n3651), .Z(n3653) );
  XOR U5727 ( .A(n3649), .B(n3648), .Z(n3895) );
  NANDN U5728 ( .A(n3895), .B(n3896), .Z(n3652) );
  AND U5729 ( .A(n3653), .B(n3652), .Z(n3656) );
  XOR U5730 ( .A(n3655), .B(n3654), .Z(n3657) );
  NANDN U5731 ( .A(n3656), .B(n3657), .Z(n3659) );
  AND U5732 ( .A(a[4]), .B(b[56]), .Z(n3883) );
  NAND U5733 ( .A(n3883), .B(n3882), .Z(n3658) );
  AND U5734 ( .A(n3659), .B(n3658), .Z(n3662) );
  NANDN U5735 ( .A(n3662), .B(n3663), .Z(n3665) );
  AND U5736 ( .A(a[5]), .B(b[56]), .Z(n3906) );
  NAND U5737 ( .A(n3906), .B(n3905), .Z(n3664) );
  AND U5738 ( .A(n3665), .B(n3664), .Z(n3668) );
  XOR U5739 ( .A(n3667), .B(n3666), .Z(n3669) );
  NANDN U5740 ( .A(n3668), .B(n3669), .Z(n3671) );
  NAND U5741 ( .A(a[6]), .B(b[56]), .Z(n3880) );
  NANDN U5742 ( .A(n3880), .B(n3881), .Z(n3670) );
  AND U5743 ( .A(n3671), .B(n3670), .Z(n3915) );
  NANDN U5744 ( .A(n3915), .B(n3916), .Z(n3674) );
  AND U5745 ( .A(n3675), .B(n3674), .Z(n3678) );
  NANDN U5746 ( .A(n3678), .B(n3679), .Z(n3681) );
  NAND U5747 ( .A(a[8]), .B(b[56]), .Z(n3878) );
  NANDN U5748 ( .A(n3878), .B(n3879), .Z(n3680) );
  AND U5749 ( .A(n3681), .B(n3680), .Z(n3685) );
  XNOR U5750 ( .A(n3683), .B(n3682), .Z(n3684) );
  NANDN U5751 ( .A(n3685), .B(n3684), .Z(n3687) );
  NAND U5752 ( .A(a[9]), .B(b[56]), .Z(n3925) );
  XNOR U5753 ( .A(n3685), .B(n3684), .Z(n3926) );
  NANDN U5754 ( .A(n3925), .B(n3926), .Z(n3686) );
  AND U5755 ( .A(n3687), .B(n3686), .Z(n3932) );
  XNOR U5756 ( .A(n3689), .B(n3688), .Z(n3931) );
  NANDN U5757 ( .A(n3932), .B(n3931), .Z(n3690) );
  AND U5758 ( .A(n3691), .B(n3690), .Z(n3877) );
  OR U5759 ( .A(n3876), .B(n3877), .Z(n3692) );
  AND U5760 ( .A(n3693), .B(n3692), .Z(n3875) );
  XNOR U5761 ( .A(n3695), .B(n3694), .Z(n3874) );
  NANDN U5762 ( .A(n3875), .B(n3874), .Z(n3696) );
  AND U5763 ( .A(n3697), .B(n3696), .Z(n3873) );
  OR U5764 ( .A(n3872), .B(n3873), .Z(n3698) );
  AND U5765 ( .A(n3699), .B(n3698), .Z(n3871) );
  OR U5766 ( .A(n3870), .B(n3871), .Z(n3700) );
  AND U5767 ( .A(n3701), .B(n3700), .Z(n3702) );
  NANDN U5768 ( .A(n3703), .B(n3702), .Z(n3705) );
  XOR U5769 ( .A(n3703), .B(n3702), .Z(n3868) );
  AND U5770 ( .A(a[15]), .B(b[56]), .Z(n3869) );
  OR U5771 ( .A(n3868), .B(n3869), .Z(n3704) );
  NAND U5772 ( .A(n3705), .B(n3704), .Z(n3706) );
  NANDN U5773 ( .A(n3707), .B(n3706), .Z(n3709) );
  XOR U5774 ( .A(n3707), .B(n3706), .Z(n3864) );
  AND U5775 ( .A(a[16]), .B(b[56]), .Z(n3865) );
  OR U5776 ( .A(n3864), .B(n3865), .Z(n3708) );
  NAND U5777 ( .A(n3709), .B(n3708), .Z(n3959) );
  XNOR U5778 ( .A(n3711), .B(n3710), .Z(n3960) );
  NANDN U5779 ( .A(n3959), .B(n3960), .Z(n3712) );
  AND U5780 ( .A(n3713), .B(n3712), .Z(n3863) );
  OR U5781 ( .A(n3862), .B(n3863), .Z(n3714) );
  AND U5782 ( .A(n3715), .B(n3714), .Z(n3716) );
  NANDN U5783 ( .A(n3717), .B(n3716), .Z(n3719) );
  XOR U5784 ( .A(n3717), .B(n3716), .Z(n3969) );
  AND U5785 ( .A(a[19]), .B(b[56]), .Z(n3970) );
  OR U5786 ( .A(n3969), .B(n3970), .Z(n3718) );
  AND U5787 ( .A(n3719), .B(n3718), .Z(n3720) );
  NANDN U5788 ( .A(n3721), .B(n3720), .Z(n3723) );
  NAND U5789 ( .A(a[20]), .B(b[56]), .Z(n3860) );
  XNOR U5790 ( .A(n3721), .B(n3720), .Z(n3861) );
  NANDN U5791 ( .A(n3860), .B(n3861), .Z(n3722) );
  AND U5792 ( .A(n3723), .B(n3722), .Z(n3859) );
  OR U5793 ( .A(n3858), .B(n3859), .Z(n3724) );
  AND U5794 ( .A(n3725), .B(n3724), .Z(n3857) );
  XNOR U5795 ( .A(n3727), .B(n3726), .Z(n3856) );
  NANDN U5796 ( .A(n3857), .B(n3856), .Z(n3728) );
  AND U5797 ( .A(n3729), .B(n3728), .Z(n3733) );
  XNOR U5798 ( .A(n3731), .B(n3730), .Z(n3732) );
  NANDN U5799 ( .A(n3733), .B(n3732), .Z(n3735) );
  NAND U5800 ( .A(a[23]), .B(b[56]), .Z(n3987) );
  XNOR U5801 ( .A(n3733), .B(n3732), .Z(n3988) );
  NANDN U5802 ( .A(n3987), .B(n3988), .Z(n3734) );
  AND U5803 ( .A(n3735), .B(n3734), .Z(n3738) );
  XOR U5804 ( .A(n3737), .B(n3736), .Z(n3739) );
  NAND U5805 ( .A(n3738), .B(n3739), .Z(n3741) );
  AND U5806 ( .A(a[24]), .B(b[56]), .Z(n3855) );
  XOR U5807 ( .A(n3739), .B(n3738), .Z(n3854) );
  NANDN U5808 ( .A(n3855), .B(n3854), .Z(n3740) );
  AND U5809 ( .A(n3741), .B(n3740), .Z(n3998) );
  XNOR U5810 ( .A(n3743), .B(n3742), .Z(n3997) );
  NAND U5811 ( .A(n3998), .B(n3997), .Z(n3744) );
  AND U5812 ( .A(n3745), .B(n3744), .Z(n4004) );
  XNOR U5813 ( .A(n3747), .B(n3746), .Z(n4003) );
  NANDN U5814 ( .A(n4004), .B(n4003), .Z(n3748) );
  AND U5815 ( .A(n3749), .B(n3748), .Z(n3750) );
  NANDN U5816 ( .A(n3751), .B(n3750), .Z(n3755) );
  XNOR U5817 ( .A(n3751), .B(n3750), .Z(n3852) );
  XNOR U5818 ( .A(n3753), .B(n3752), .Z(n3853) );
  NAND U5819 ( .A(n3852), .B(n3853), .Z(n3754) );
  NAND U5820 ( .A(n3755), .B(n3754), .Z(n3756) );
  NANDN U5821 ( .A(n3757), .B(n3756), .Z(n3761) );
  XNOR U5822 ( .A(n3757), .B(n3756), .Z(n4015) );
  XNOR U5823 ( .A(n3759), .B(n3758), .Z(n4016) );
  NAND U5824 ( .A(n4015), .B(n4016), .Z(n3760) );
  NAND U5825 ( .A(n3761), .B(n3760), .Z(n3762) );
  NANDN U5826 ( .A(n3763), .B(n3762), .Z(n3767) );
  XNOR U5827 ( .A(n3763), .B(n3762), .Z(n4021) );
  XNOR U5828 ( .A(n3765), .B(n3764), .Z(n4022) );
  NAND U5829 ( .A(n4021), .B(n4022), .Z(n3766) );
  NAND U5830 ( .A(n3767), .B(n3766), .Z(n3770) );
  NANDN U5831 ( .A(n3771), .B(n3770), .Z(n3773) );
  XOR U5832 ( .A(n3769), .B(n3768), .Z(n4028) );
  XNOR U5833 ( .A(n3771), .B(n3770), .Z(n4027) );
  NANDN U5834 ( .A(n4028), .B(n4027), .Z(n3772) );
  NAND U5835 ( .A(n3773), .B(n3772), .Z(n3774) );
  NANDN U5836 ( .A(n3775), .B(n3774), .Z(n3779) );
  XNOR U5837 ( .A(n3775), .B(n3774), .Z(n4032) );
  XNOR U5838 ( .A(n3777), .B(n3776), .Z(n4031) );
  NAND U5839 ( .A(n4032), .B(n4031), .Z(n3778) );
  NAND U5840 ( .A(n3779), .B(n3778), .Z(n3780) );
  NANDN U5841 ( .A(n3781), .B(n3780), .Z(n3785) );
  XNOR U5842 ( .A(n3781), .B(n3780), .Z(n4038) );
  XNOR U5843 ( .A(n3783), .B(n3782), .Z(n4037) );
  NAND U5844 ( .A(n4038), .B(n4037), .Z(n3784) );
  AND U5845 ( .A(n3785), .B(n3784), .Z(n3789) );
  NANDN U5846 ( .A(n3788), .B(n3789), .Z(n3791) );
  XOR U5847 ( .A(n3787), .B(n3786), .Z(n4046) );
  XNOR U5848 ( .A(n3789), .B(n3788), .Z(n4045) );
  NANDN U5849 ( .A(n4046), .B(n4045), .Z(n3790) );
  AND U5850 ( .A(n3791), .B(n3790), .Z(n3792) );
  NANDN U5851 ( .A(n3793), .B(n3792), .Z(n3797) );
  XNOR U5852 ( .A(n3793), .B(n3792), .Z(n4051) );
  XOR U5853 ( .A(n3795), .B(n3794), .Z(n4052) );
  NAND U5854 ( .A(n4051), .B(n4052), .Z(n3796) );
  NAND U5855 ( .A(n3797), .B(n3796), .Z(n3799) );
  NANDN U5856 ( .A(n3798), .B(n3799), .Z(n3803) );
  XNOR U5857 ( .A(n3801), .B(n3800), .Z(n4058) );
  NAND U5858 ( .A(n4057), .B(n4058), .Z(n3802) );
  AND U5859 ( .A(n3803), .B(n3802), .Z(n3807) );
  NANDN U5860 ( .A(n3806), .B(n3807), .Z(n3809) );
  XOR U5861 ( .A(n3805), .B(n3804), .Z(n4064) );
  NAND U5862 ( .A(n4064), .B(n4063), .Z(n3808) );
  AND U5863 ( .A(n3809), .B(n3808), .Z(n3813) );
  NANDN U5864 ( .A(n3812), .B(n3813), .Z(n3815) );
  XOR U5865 ( .A(n3811), .B(n3810), .Z(n4069) );
  NANDN U5866 ( .A(n4069), .B(n4070), .Z(n3814) );
  NAND U5867 ( .A(n3815), .B(n3814), .Z(n3817) );
  NANDN U5868 ( .A(n3816), .B(n3817), .Z(n3821) );
  XNOR U5869 ( .A(n3819), .B(n3818), .Z(n4076) );
  NAND U5870 ( .A(n4075), .B(n4076), .Z(n3820) );
  NAND U5871 ( .A(n3821), .B(n3820), .Z(n3823) );
  NANDN U5872 ( .A(n3822), .B(n3823), .Z(n3827) );
  XNOR U5873 ( .A(n3825), .B(n3824), .Z(n4082) );
  NAND U5874 ( .A(n4081), .B(n4082), .Z(n3826) );
  NAND U5875 ( .A(n3827), .B(n3826), .Z(n3831) );
  NANDN U5876 ( .A(n3830), .B(n3831), .Z(n3833) );
  XOR U5877 ( .A(n3829), .B(n3828), .Z(n4085) );
  NANDN U5878 ( .A(n4085), .B(n4086), .Z(n3832) );
  NAND U5879 ( .A(n3833), .B(n3832), .Z(n3835) );
  NANDN U5880 ( .A(n3834), .B(n3835), .Z(n3839) );
  XNOR U5881 ( .A(n3837), .B(n3836), .Z(n4094) );
  NAND U5882 ( .A(n4093), .B(n4094), .Z(n3838) );
  NAND U5883 ( .A(n3839), .B(n3838), .Z(n3842) );
  AND U5884 ( .A(a[42]), .B(b[56]), .Z(n3843) );
  NANDN U5885 ( .A(n3842), .B(n3843), .Z(n3845) );
  XOR U5886 ( .A(n3841), .B(n3840), .Z(n4098) );
  NAND U5887 ( .A(n4098), .B(n4097), .Z(n3844) );
  AND U5888 ( .A(n3845), .B(n3844), .Z(n3849) );
  NANDN U5889 ( .A(n3848), .B(n3849), .Z(n3851) );
  XOR U5890 ( .A(n3847), .B(n3846), .Z(n4105) );
  NANDN U5891 ( .A(n4105), .B(n4106), .Z(n3850) );
  NAND U5892 ( .A(n3851), .B(n3850), .Z(n10166) );
  XNOR U5893 ( .A(n10168), .B(n10169), .Z(n10174) );
  AND U5894 ( .A(a[45]), .B(b[55]), .Z(n10172) );
  AND U5895 ( .A(a[44]), .B(b[55]), .Z(n4103) );
  AND U5896 ( .A(a[43]), .B(b[55]), .Z(n4099) );
  AND U5897 ( .A(a[41]), .B(b[55]), .Z(n4087) );
  AND U5898 ( .A(a[38]), .B(b[55]), .Z(n4067) );
  NAND U5899 ( .A(a[36]), .B(b[55]), .Z(n4055) );
  AND U5900 ( .A(a[35]), .B(b[55]), .Z(n4050) );
  NAND U5901 ( .A(a[32]), .B(b[55]), .Z(n4033) );
  AND U5902 ( .A(a[31]), .B(b[55]), .Z(n4026) );
  AND U5903 ( .A(a[28]), .B(b[55]), .Z(n4009) );
  XNOR U5904 ( .A(n3853), .B(n3852), .Z(n4010) );
  NAND U5905 ( .A(n4009), .B(n4010), .Z(n4012) );
  AND U5906 ( .A(a[25]), .B(b[55]), .Z(n3993) );
  XOR U5907 ( .A(n3855), .B(n3854), .Z(n3994) );
  NAND U5908 ( .A(n3993), .B(n3994), .Z(n3996) );
  XOR U5909 ( .A(n3857), .B(n3856), .Z(n3983) );
  XOR U5910 ( .A(n3859), .B(n3858), .Z(n3980) );
  NAND U5911 ( .A(a[21]), .B(b[55]), .Z(n3975) );
  XNOR U5912 ( .A(n3861), .B(n3860), .Z(n3976) );
  NANDN U5913 ( .A(n3975), .B(n3976), .Z(n3978) );
  NAND U5914 ( .A(a[20]), .B(b[55]), .Z(n3971) );
  AND U5915 ( .A(a[19]), .B(b[55]), .Z(n3966) );
  XNOR U5916 ( .A(n3863), .B(n3862), .Z(n3965) );
  NANDN U5917 ( .A(n3966), .B(n3965), .Z(n3968) );
  XOR U5918 ( .A(n3865), .B(n3864), .Z(n3867) );
  AND U5919 ( .A(a[17]), .B(b[55]), .Z(n3866) );
  NANDN U5920 ( .A(n3867), .B(n3866), .Z(n3958) );
  XOR U5921 ( .A(n3867), .B(n3866), .Z(n4127) );
  XOR U5922 ( .A(n3869), .B(n3868), .Z(n3954) );
  XOR U5923 ( .A(n3871), .B(n3870), .Z(n3950) );
  XOR U5924 ( .A(n3873), .B(n3872), .Z(n3946) );
  NAND U5925 ( .A(a[13]), .B(b[55]), .Z(n3941) );
  XNOR U5926 ( .A(n3875), .B(n3874), .Z(n3942) );
  NANDN U5927 ( .A(n3941), .B(n3942), .Z(n3944) );
  XOR U5928 ( .A(n3877), .B(n3876), .Z(n3938) );
  AND U5929 ( .A(a[9]), .B(b[55]), .Z(n3922) );
  NAND U5930 ( .A(n3922), .B(n3921), .Z(n3924) );
  NAND U5931 ( .A(a[7]), .B(b[55]), .Z(n3911) );
  NANDN U5932 ( .A(n3911), .B(n3912), .Z(n3914) );
  XOR U5933 ( .A(n3883), .B(n3882), .Z(n3901) );
  NAND U5934 ( .A(a[0]), .B(b[55]), .Z(n4411) );
  AND U5935 ( .A(a[1]), .B(b[56]), .Z(n3886) );
  NANDN U5936 ( .A(n4411), .B(n3886), .Z(n4147) );
  NANDN U5937 ( .A(n4147), .B(n3884), .Z(n3888) );
  AND U5938 ( .A(a[2]), .B(b[55]), .Z(n4153) );
  NANDN U5939 ( .A(n4152), .B(n4153), .Z(n3887) );
  AND U5940 ( .A(n3888), .B(n3887), .Z(n3891) );
  AND U5941 ( .A(a[3]), .B(b[55]), .Z(n3892) );
  NANDN U5942 ( .A(n3891), .B(n3892), .Z(n3894) );
  XOR U5943 ( .A(n3890), .B(n3889), .Z(n4158) );
  NANDN U5944 ( .A(n4158), .B(n4159), .Z(n3893) );
  AND U5945 ( .A(n3894), .B(n3893), .Z(n3897) );
  NANDN U5946 ( .A(n3897), .B(n3898), .Z(n3900) );
  AND U5947 ( .A(a[4]), .B(b[55]), .Z(n4165) );
  NAND U5948 ( .A(n4165), .B(n4164), .Z(n3899) );
  AND U5949 ( .A(n3900), .B(n3899), .Z(n3902) );
  NANDN U5950 ( .A(n3901), .B(n3902), .Z(n3904) );
  AND U5951 ( .A(a[5]), .B(b[55]), .Z(n4171) );
  NANDN U5952 ( .A(n4171), .B(n4170), .Z(n3903) );
  AND U5953 ( .A(n3904), .B(n3903), .Z(n3908) );
  XOR U5954 ( .A(n3906), .B(n3905), .Z(n3907) );
  NAND U5955 ( .A(n3908), .B(n3907), .Z(n3910) );
  AND U5956 ( .A(a[6]), .B(b[55]), .Z(n4146) );
  XOR U5957 ( .A(n3908), .B(n3907), .Z(n4145) );
  NAND U5958 ( .A(n4146), .B(n4145), .Z(n3909) );
  AND U5959 ( .A(n3910), .B(n3909), .Z(n4180) );
  NANDN U5960 ( .A(n4180), .B(n4181), .Z(n3913) );
  AND U5961 ( .A(n3914), .B(n3913), .Z(n3917) );
  AND U5962 ( .A(a[8]), .B(b[55]), .Z(n3918) );
  NANDN U5963 ( .A(n3917), .B(n3918), .Z(n3920) );
  NAND U5964 ( .A(n4144), .B(n4143), .Z(n3919) );
  AND U5965 ( .A(n3920), .B(n3919), .Z(n4141) );
  XOR U5966 ( .A(n3922), .B(n3921), .Z(n4142) );
  NANDN U5967 ( .A(n4141), .B(n4142), .Z(n3923) );
  AND U5968 ( .A(n3924), .B(n3923), .Z(n3928) );
  AND U5969 ( .A(a[10]), .B(b[55]), .Z(n3927) );
  NANDN U5970 ( .A(n3928), .B(n3927), .Z(n3930) );
  XOR U5971 ( .A(n3926), .B(n3925), .Z(n4139) );
  XNOR U5972 ( .A(n3928), .B(n3927), .Z(n4140) );
  NANDN U5973 ( .A(n4139), .B(n4140), .Z(n3929) );
  AND U5974 ( .A(n3930), .B(n3929), .Z(n3934) );
  XNOR U5975 ( .A(n3932), .B(n3931), .Z(n3933) );
  NANDN U5976 ( .A(n3934), .B(n3933), .Z(n3936) );
  NAND U5977 ( .A(a[11]), .B(b[55]), .Z(n4198) );
  XNOR U5978 ( .A(n3934), .B(n3933), .Z(n4199) );
  NANDN U5979 ( .A(n4198), .B(n4199), .Z(n3935) );
  AND U5980 ( .A(n3936), .B(n3935), .Z(n3937) );
  NANDN U5981 ( .A(n3938), .B(n3937), .Z(n3940) );
  XOR U5982 ( .A(n3938), .B(n3937), .Z(n4137) );
  AND U5983 ( .A(a[12]), .B(b[55]), .Z(n4138) );
  OR U5984 ( .A(n4137), .B(n4138), .Z(n3939) );
  NAND U5985 ( .A(n3940), .B(n3939), .Z(n4208) );
  XNOR U5986 ( .A(n3942), .B(n3941), .Z(n4209) );
  NANDN U5987 ( .A(n4208), .B(n4209), .Z(n3943) );
  AND U5988 ( .A(n3944), .B(n3943), .Z(n3945) );
  NANDN U5989 ( .A(n3946), .B(n3945), .Z(n3948) );
  XOR U5990 ( .A(n3946), .B(n3945), .Z(n4135) );
  AND U5991 ( .A(a[14]), .B(b[55]), .Z(n4136) );
  OR U5992 ( .A(n4135), .B(n4136), .Z(n3947) );
  NAND U5993 ( .A(n3948), .B(n3947), .Z(n3949) );
  NANDN U5994 ( .A(n3950), .B(n3949), .Z(n3952) );
  XOR U5995 ( .A(n3950), .B(n3949), .Z(n4133) );
  AND U5996 ( .A(a[15]), .B(b[55]), .Z(n4134) );
  OR U5997 ( .A(n4133), .B(n4134), .Z(n3951) );
  AND U5998 ( .A(n3952), .B(n3951), .Z(n3953) );
  NANDN U5999 ( .A(n3954), .B(n3953), .Z(n3956) );
  XNOR U6000 ( .A(n3954), .B(n3953), .Z(n4132) );
  AND U6001 ( .A(a[16]), .B(b[55]), .Z(n4131) );
  NAND U6002 ( .A(n4132), .B(n4131), .Z(n3955) );
  AND U6003 ( .A(n3956), .B(n3955), .Z(n4128) );
  OR U6004 ( .A(n4127), .B(n4128), .Z(n3957) );
  AND U6005 ( .A(n3958), .B(n3957), .Z(n3962) );
  XNOR U6006 ( .A(n3960), .B(n3959), .Z(n3961) );
  NANDN U6007 ( .A(n3962), .B(n3961), .Z(n3964) );
  NAND U6008 ( .A(a[18]), .B(b[55]), .Z(n4125) );
  XNOR U6009 ( .A(n3962), .B(n3961), .Z(n4126) );
  NANDN U6010 ( .A(n4125), .B(n4126), .Z(n3963) );
  AND U6011 ( .A(n3964), .B(n3963), .Z(n4124) );
  XNOR U6012 ( .A(n3966), .B(n3965), .Z(n4123) );
  NAND U6013 ( .A(n4124), .B(n4123), .Z(n3967) );
  AND U6014 ( .A(n3968), .B(n3967), .Z(n3972) );
  NANDN U6015 ( .A(n3971), .B(n3972), .Z(n3974) );
  XOR U6016 ( .A(n3970), .B(n3969), .Z(n4239) );
  XNOR U6017 ( .A(n3972), .B(n3971), .Z(n4238) );
  NANDN U6018 ( .A(n4239), .B(n4238), .Z(n3973) );
  AND U6019 ( .A(n3974), .B(n3973), .Z(n4243) );
  XNOR U6020 ( .A(n3976), .B(n3975), .Z(n4242) );
  NANDN U6021 ( .A(n4243), .B(n4242), .Z(n3977) );
  AND U6022 ( .A(n3978), .B(n3977), .Z(n3979) );
  NANDN U6023 ( .A(n3980), .B(n3979), .Z(n3982) );
  XOR U6024 ( .A(n3980), .B(n3979), .Z(n4121) );
  AND U6025 ( .A(a[22]), .B(b[55]), .Z(n4122) );
  OR U6026 ( .A(n4121), .B(n4122), .Z(n3981) );
  AND U6027 ( .A(n3982), .B(n3981), .Z(n3984) );
  NANDN U6028 ( .A(n3983), .B(n3984), .Z(n3986) );
  NAND U6029 ( .A(a[23]), .B(b[55]), .Z(n4119) );
  XNOR U6030 ( .A(n3984), .B(n3983), .Z(n4120) );
  NANDN U6031 ( .A(n4119), .B(n4120), .Z(n3985) );
  AND U6032 ( .A(n3986), .B(n3985), .Z(n3990) );
  XNOR U6033 ( .A(n3988), .B(n3987), .Z(n3989) );
  NANDN U6034 ( .A(n3990), .B(n3989), .Z(n3992) );
  NAND U6035 ( .A(a[24]), .B(b[55]), .Z(n4117) );
  XNOR U6036 ( .A(n3990), .B(n3989), .Z(n4118) );
  NANDN U6037 ( .A(n4117), .B(n4118), .Z(n3991) );
  AND U6038 ( .A(n3992), .B(n3991), .Z(n4261) );
  XOR U6039 ( .A(n3994), .B(n3993), .Z(n4260) );
  NANDN U6040 ( .A(n4261), .B(n4260), .Z(n3995) );
  AND U6041 ( .A(n3996), .B(n3995), .Z(n4000) );
  XOR U6042 ( .A(n3998), .B(n3997), .Z(n3999) );
  NANDN U6043 ( .A(n4000), .B(n3999), .Z(n4002) );
  NAND U6044 ( .A(a[26]), .B(b[55]), .Z(n4115) );
  XNOR U6045 ( .A(n4000), .B(n3999), .Z(n4116) );
  NANDN U6046 ( .A(n4115), .B(n4116), .Z(n4001) );
  AND U6047 ( .A(n4002), .B(n4001), .Z(n4006) );
  XNOR U6048 ( .A(n4004), .B(n4003), .Z(n4005) );
  NANDN U6049 ( .A(n4006), .B(n4005), .Z(n4008) );
  NAND U6050 ( .A(a[27]), .B(b[55]), .Z(n4113) );
  XNOR U6051 ( .A(n4006), .B(n4005), .Z(n4114) );
  NANDN U6052 ( .A(n4113), .B(n4114), .Z(n4007) );
  AND U6053 ( .A(n4008), .B(n4007), .Z(n4112) );
  XOR U6054 ( .A(n4010), .B(n4009), .Z(n4111) );
  NANDN U6055 ( .A(n4112), .B(n4111), .Z(n4011) );
  AND U6056 ( .A(n4012), .B(n4011), .Z(n4014) );
  AND U6057 ( .A(a[29]), .B(b[55]), .Z(n4013) );
  NANDN U6058 ( .A(n4014), .B(n4013), .Z(n4018) );
  XNOR U6059 ( .A(n4014), .B(n4013), .Z(n4109) );
  XNOR U6060 ( .A(n4016), .B(n4015), .Z(n4110) );
  NAND U6061 ( .A(n4109), .B(n4110), .Z(n4017) );
  AND U6062 ( .A(n4018), .B(n4017), .Z(n4020) );
  AND U6063 ( .A(a[30]), .B(b[55]), .Z(n4019) );
  NANDN U6064 ( .A(n4020), .B(n4019), .Z(n4024) );
  XNOR U6065 ( .A(n4020), .B(n4019), .Z(n4284) );
  XNOR U6066 ( .A(n4022), .B(n4021), .Z(n4285) );
  NAND U6067 ( .A(n4284), .B(n4285), .Z(n4023) );
  AND U6068 ( .A(n4024), .B(n4023), .Z(n4025) );
  NANDN U6069 ( .A(n4026), .B(n4025), .Z(n4030) );
  XNOR U6070 ( .A(n4026), .B(n4025), .Z(n4289) );
  XNOR U6071 ( .A(n4028), .B(n4027), .Z(n4288) );
  NAND U6072 ( .A(n4289), .B(n4288), .Z(n4029) );
  AND U6073 ( .A(n4030), .B(n4029), .Z(n4034) );
  NANDN U6074 ( .A(n4033), .B(n4034), .Z(n4036) );
  XOR U6075 ( .A(n4032), .B(n4031), .Z(n4295) );
  XNOR U6076 ( .A(n4034), .B(n4033), .Z(n4294) );
  NANDN U6077 ( .A(n4295), .B(n4294), .Z(n4035) );
  AND U6078 ( .A(n4036), .B(n4035), .Z(n4040) );
  AND U6079 ( .A(a[33]), .B(b[55]), .Z(n4039) );
  NANDN U6080 ( .A(n4040), .B(n4039), .Z(n4042) );
  XOR U6081 ( .A(n4038), .B(n4037), .Z(n4301) );
  XNOR U6082 ( .A(n4040), .B(n4039), .Z(n4300) );
  NANDN U6083 ( .A(n4301), .B(n4300), .Z(n4041) );
  AND U6084 ( .A(n4042), .B(n4041), .Z(n4044) );
  AND U6085 ( .A(a[34]), .B(b[55]), .Z(n4043) );
  NANDN U6086 ( .A(n4044), .B(n4043), .Z(n4048) );
  XNOR U6087 ( .A(n4044), .B(n4043), .Z(n4307) );
  XNOR U6088 ( .A(n4046), .B(n4045), .Z(n4306) );
  NAND U6089 ( .A(n4307), .B(n4306), .Z(n4047) );
  AND U6090 ( .A(n4048), .B(n4047), .Z(n4049) );
  NANDN U6091 ( .A(n4050), .B(n4049), .Z(n4054) );
  XNOR U6092 ( .A(n4050), .B(n4049), .Z(n4313) );
  XOR U6093 ( .A(n4052), .B(n4051), .Z(n4312) );
  NAND U6094 ( .A(n4313), .B(n4312), .Z(n4053) );
  AND U6095 ( .A(n4054), .B(n4053), .Z(n4056) );
  NANDN U6096 ( .A(n4055), .B(n4056), .Z(n4060) );
  XNOR U6097 ( .A(n4058), .B(n4057), .Z(n4321) );
  NAND U6098 ( .A(n4320), .B(n4321), .Z(n4059) );
  AND U6099 ( .A(n4060), .B(n4059), .Z(n4061) );
  AND U6100 ( .A(a[37]), .B(b[55]), .Z(n4062) );
  NANDN U6101 ( .A(n4061), .B(n4062), .Z(n4066) );
  XOR U6102 ( .A(n4064), .B(n4063), .Z(n4324) );
  NAND U6103 ( .A(n4325), .B(n4324), .Z(n4065) );
  AND U6104 ( .A(n4066), .B(n4065), .Z(n4068) );
  NANDN U6105 ( .A(n4067), .B(n4068), .Z(n4072) );
  NAND U6106 ( .A(n4331), .B(n4330), .Z(n4071) );
  NAND U6107 ( .A(n4072), .B(n4071), .Z(n4073) );
  AND U6108 ( .A(a[39]), .B(b[55]), .Z(n4074) );
  NANDN U6109 ( .A(n4073), .B(n4074), .Z(n4078) );
  XNOR U6110 ( .A(n4076), .B(n4075), .Z(n4339) );
  NAND U6111 ( .A(n4338), .B(n4339), .Z(n4077) );
  AND U6112 ( .A(n4078), .B(n4077), .Z(n4079) );
  AND U6113 ( .A(a[40]), .B(b[55]), .Z(n4080) );
  NANDN U6114 ( .A(n4079), .B(n4080), .Z(n4084) );
  XNOR U6115 ( .A(n4082), .B(n4081), .Z(n4345) );
  NAND U6116 ( .A(n4344), .B(n4345), .Z(n4083) );
  AND U6117 ( .A(n4084), .B(n4083), .Z(n4088) );
  NANDN U6118 ( .A(n4087), .B(n4088), .Z(n4090) );
  NAND U6119 ( .A(n4349), .B(n4348), .Z(n4089) );
  NAND U6120 ( .A(n4090), .B(n4089), .Z(n4091) );
  AND U6121 ( .A(a[42]), .B(b[55]), .Z(n4092) );
  NANDN U6122 ( .A(n4091), .B(n4092), .Z(n4096) );
  XNOR U6123 ( .A(n4094), .B(n4093), .Z(n4357) );
  NAND U6124 ( .A(n4356), .B(n4357), .Z(n4095) );
  AND U6125 ( .A(n4096), .B(n4095), .Z(n4100) );
  NANDN U6126 ( .A(n4099), .B(n4100), .Z(n4102) );
  XOR U6127 ( .A(n4098), .B(n4097), .Z(n4362) );
  NANDN U6128 ( .A(n4362), .B(n4363), .Z(n4101) );
  NAND U6129 ( .A(n4102), .B(n4101), .Z(n4104) );
  NANDN U6130 ( .A(n4103), .B(n4104), .Z(n4108) );
  NAND U6131 ( .A(n4367), .B(n4366), .Z(n4107) );
  NAND U6132 ( .A(n4108), .B(n4107), .Z(n10173) );
  XNOR U6133 ( .A(n10174), .B(n10175), .Z(n10126) );
  AND U6134 ( .A(a[46]), .B(b[54]), .Z(n10125) );
  AND U6135 ( .A(a[44]), .B(b[54]), .Z(n4360) );
  AND U6136 ( .A(a[43]), .B(b[54]), .Z(n4354) );
  AND U6137 ( .A(a[41]), .B(b[54]), .Z(n4342) );
  AND U6138 ( .A(a[40]), .B(b[54]), .Z(n4336) );
  NAND U6139 ( .A(a[39]), .B(b[54]), .Z(n4332) );
  AND U6140 ( .A(a[38]), .B(b[54]), .Z(n4326) );
  AND U6141 ( .A(a[37]), .B(b[54]), .Z(n4318) );
  NAND U6142 ( .A(a[36]), .B(b[54]), .Z(n4314) );
  AND U6143 ( .A(a[35]), .B(b[54]), .Z(n4309) );
  NAND U6144 ( .A(a[32]), .B(b[54]), .Z(n4290) );
  AND U6145 ( .A(a[31]), .B(b[54]), .Z(n4283) );
  NAND U6146 ( .A(a[30]), .B(b[54]), .Z(n4278) );
  XOR U6147 ( .A(n4110), .B(n4109), .Z(n4279) );
  NANDN U6148 ( .A(n4278), .B(n4279), .Z(n4281) );
  NAND U6149 ( .A(a[29]), .B(b[54]), .Z(n4274) );
  XNOR U6150 ( .A(n4112), .B(n4111), .Z(n4275) );
  NANDN U6151 ( .A(n4274), .B(n4275), .Z(n4277) );
  NAND U6152 ( .A(a[28]), .B(b[54]), .Z(n4270) );
  XNOR U6153 ( .A(n4114), .B(n4113), .Z(n4271) );
  NANDN U6154 ( .A(n4270), .B(n4271), .Z(n4273) );
  NAND U6155 ( .A(a[27]), .B(b[54]), .Z(n4266) );
  XNOR U6156 ( .A(n4116), .B(n4115), .Z(n4267) );
  NANDN U6157 ( .A(n4266), .B(n4267), .Z(n4269) );
  NAND U6158 ( .A(a[25]), .B(b[54]), .Z(n4256) );
  XNOR U6159 ( .A(n4118), .B(n4117), .Z(n4257) );
  NANDN U6160 ( .A(n4256), .B(n4257), .Z(n4259) );
  NAND U6161 ( .A(a[24]), .B(b[54]), .Z(n4252) );
  XNOR U6162 ( .A(n4120), .B(n4119), .Z(n4253) );
  NANDN U6163 ( .A(n4252), .B(n4253), .Z(n4255) );
  XOR U6164 ( .A(n4122), .B(n4121), .Z(n4249) );
  XOR U6165 ( .A(n4124), .B(n4123), .Z(n4233) );
  AND U6166 ( .A(a[20]), .B(b[54]), .Z(n4232) );
  NANDN U6167 ( .A(n4233), .B(n4232), .Z(n4235) );
  XOR U6168 ( .A(n4126), .B(n4125), .Z(n4228) );
  AND U6169 ( .A(a[18]), .B(b[54]), .Z(n4130) );
  XNOR U6170 ( .A(n4128), .B(n4127), .Z(n4129) );
  NANDN U6171 ( .A(n4130), .B(n4129), .Z(n4227) );
  XOR U6172 ( .A(n4130), .B(n4129), .Z(n4394) );
  XOR U6173 ( .A(n4132), .B(n4131), .Z(n4223) );
  XOR U6174 ( .A(n4134), .B(n4133), .Z(n4219) );
  AND U6175 ( .A(a[16]), .B(b[54]), .Z(n4218) );
  NANDN U6176 ( .A(n4219), .B(n4218), .Z(n4221) );
  XOR U6177 ( .A(n4136), .B(n4135), .Z(n4215) );
  AND U6178 ( .A(a[15]), .B(b[54]), .Z(n4214) );
  NANDN U6179 ( .A(n4215), .B(n4214), .Z(n4217) );
  XOR U6180 ( .A(n4138), .B(n4137), .Z(n4205) );
  AND U6181 ( .A(a[13]), .B(b[54]), .Z(n4204) );
  NANDN U6182 ( .A(n4205), .B(n4204), .Z(n4207) );
  XOR U6183 ( .A(n4140), .B(n4139), .Z(n4194) );
  XOR U6184 ( .A(n4144), .B(n4143), .Z(n4186) );
  NAND U6185 ( .A(a[7]), .B(b[54]), .Z(n4176) );
  XOR U6186 ( .A(n4146), .B(n4145), .Z(n4177) );
  NANDN U6187 ( .A(n4176), .B(n4177), .Z(n4179) );
  NAND U6188 ( .A(a[0]), .B(b[54]), .Z(n4682) );
  AND U6189 ( .A(a[1]), .B(b[55]), .Z(n4149) );
  NANDN U6190 ( .A(n4682), .B(n4149), .Z(n4410) );
  NANDN U6191 ( .A(n4410), .B(n4147), .Z(n4151) );
  AND U6192 ( .A(a[2]), .B(b[54]), .Z(n4416) );
  NANDN U6193 ( .A(n4415), .B(n4416), .Z(n4150) );
  AND U6194 ( .A(n4151), .B(n4150), .Z(n4154) );
  AND U6195 ( .A(a[3]), .B(b[54]), .Z(n4155) );
  NANDN U6196 ( .A(n4154), .B(n4155), .Z(n4157) );
  XOR U6197 ( .A(n4153), .B(n4152), .Z(n4421) );
  NANDN U6198 ( .A(n4421), .B(n4422), .Z(n4156) );
  AND U6199 ( .A(n4157), .B(n4156), .Z(n4160) );
  NANDN U6200 ( .A(n4160), .B(n4161), .Z(n4163) );
  AND U6201 ( .A(a[4]), .B(b[54]), .Z(n4430) );
  NAND U6202 ( .A(n4430), .B(n4429), .Z(n4162) );
  AND U6203 ( .A(n4163), .B(n4162), .Z(n4166) );
  XOR U6204 ( .A(n4165), .B(n4164), .Z(n4167) );
  NANDN U6205 ( .A(n4166), .B(n4167), .Z(n4169) );
  AND U6206 ( .A(a[5]), .B(b[54]), .Z(n4434) );
  NAND U6207 ( .A(n4434), .B(n4433), .Z(n4168) );
  AND U6208 ( .A(n4169), .B(n4168), .Z(n4172) );
  XOR U6209 ( .A(n4171), .B(n4170), .Z(n4173) );
  NANDN U6210 ( .A(n4172), .B(n4173), .Z(n4175) );
  AND U6211 ( .A(a[6]), .B(b[54]), .Z(n4409) );
  NAND U6212 ( .A(n4409), .B(n4408), .Z(n4174) );
  AND U6213 ( .A(n4175), .B(n4174), .Z(n4445) );
  NANDN U6214 ( .A(n4445), .B(n4446), .Z(n4178) );
  AND U6215 ( .A(n4179), .B(n4178), .Z(n4182) );
  AND U6216 ( .A(a[8]), .B(b[54]), .Z(n4183) );
  NANDN U6217 ( .A(n4182), .B(n4183), .Z(n4185) );
  NAND U6218 ( .A(n4407), .B(n4406), .Z(n4184) );
  AND U6219 ( .A(n4185), .B(n4184), .Z(n4187) );
  NANDN U6220 ( .A(n4186), .B(n4187), .Z(n4189) );
  AND U6221 ( .A(a[9]), .B(b[54]), .Z(n4453) );
  NANDN U6222 ( .A(n4453), .B(n4454), .Z(n4188) );
  NAND U6223 ( .A(n4189), .B(n4188), .Z(n4190) );
  NAND U6224 ( .A(n4191), .B(n4190), .Z(n4193) );
  AND U6225 ( .A(a[10]), .B(b[54]), .Z(n4404) );
  XOR U6226 ( .A(n4191), .B(n4190), .Z(n4405) );
  NANDN U6227 ( .A(n4404), .B(n4405), .Z(n4192) );
  AND U6228 ( .A(n4193), .B(n4192), .Z(n4195) );
  NANDN U6229 ( .A(n4194), .B(n4195), .Z(n4197) );
  NAND U6230 ( .A(a[11]), .B(b[54]), .Z(n4402) );
  XNOR U6231 ( .A(n4195), .B(n4194), .Z(n4403) );
  NANDN U6232 ( .A(n4402), .B(n4403), .Z(n4196) );
  AND U6233 ( .A(n4197), .B(n4196), .Z(n4201) );
  XNOR U6234 ( .A(n4199), .B(n4198), .Z(n4200) );
  NANDN U6235 ( .A(n4201), .B(n4200), .Z(n4203) );
  NAND U6236 ( .A(a[12]), .B(b[54]), .Z(n4400) );
  XNOR U6237 ( .A(n4201), .B(n4200), .Z(n4401) );
  NANDN U6238 ( .A(n4400), .B(n4401), .Z(n4202) );
  AND U6239 ( .A(n4203), .B(n4202), .Z(n4472) );
  XNOR U6240 ( .A(n4205), .B(n4204), .Z(n4471) );
  NANDN U6241 ( .A(n4472), .B(n4471), .Z(n4206) );
  AND U6242 ( .A(n4207), .B(n4206), .Z(n4211) );
  XNOR U6243 ( .A(n4209), .B(n4208), .Z(n4210) );
  NANDN U6244 ( .A(n4211), .B(n4210), .Z(n4213) );
  NAND U6245 ( .A(a[14]), .B(b[54]), .Z(n4477) );
  XNOR U6246 ( .A(n4211), .B(n4210), .Z(n4478) );
  NANDN U6247 ( .A(n4477), .B(n4478), .Z(n4212) );
  AND U6248 ( .A(n4213), .B(n4212), .Z(n4399) );
  XNOR U6249 ( .A(n4215), .B(n4214), .Z(n4398) );
  NANDN U6250 ( .A(n4399), .B(n4398), .Z(n4216) );
  AND U6251 ( .A(n4217), .B(n4216), .Z(n4488) );
  XNOR U6252 ( .A(n4219), .B(n4218), .Z(n4487) );
  NANDN U6253 ( .A(n4488), .B(n4487), .Z(n4220) );
  AND U6254 ( .A(n4221), .B(n4220), .Z(n4222) );
  NANDN U6255 ( .A(n4223), .B(n4222), .Z(n4225) );
  AND U6256 ( .A(a[17]), .B(b[54]), .Z(n4397) );
  XNOR U6257 ( .A(n4223), .B(n4222), .Z(n4396) );
  NANDN U6258 ( .A(n4397), .B(n4396), .Z(n4224) );
  AND U6259 ( .A(n4225), .B(n4224), .Z(n4395) );
  OR U6260 ( .A(n4394), .B(n4395), .Z(n4226) );
  AND U6261 ( .A(n4227), .B(n4226), .Z(n4229) );
  NANDN U6262 ( .A(n4228), .B(n4229), .Z(n4231) );
  NAND U6263 ( .A(a[19]), .B(b[54]), .Z(n4390) );
  XNOR U6264 ( .A(n4229), .B(n4228), .Z(n4391) );
  NANDN U6265 ( .A(n4390), .B(n4391), .Z(n4230) );
  AND U6266 ( .A(n4231), .B(n4230), .Z(n4504) );
  XNOR U6267 ( .A(n4233), .B(n4232), .Z(n4503) );
  NANDN U6268 ( .A(n4504), .B(n4503), .Z(n4234) );
  AND U6269 ( .A(n4235), .B(n4234), .Z(n4237) );
  AND U6270 ( .A(a[21]), .B(b[54]), .Z(n4236) );
  NANDN U6271 ( .A(n4237), .B(n4236), .Z(n4241) );
  XOR U6272 ( .A(n4237), .B(n4236), .Z(n4509) );
  XNOR U6273 ( .A(n4239), .B(n4238), .Z(n4510) );
  NANDN U6274 ( .A(n4509), .B(n4510), .Z(n4240) );
  AND U6275 ( .A(n4241), .B(n4240), .Z(n4245) );
  XNOR U6276 ( .A(n4243), .B(n4242), .Z(n4244) );
  NANDN U6277 ( .A(n4245), .B(n4244), .Z(n4247) );
  XNOR U6278 ( .A(n4245), .B(n4244), .Z(n4389) );
  AND U6279 ( .A(a[22]), .B(b[54]), .Z(n4388) );
  NAND U6280 ( .A(n4389), .B(n4388), .Z(n4246) );
  NAND U6281 ( .A(n4247), .B(n4246), .Z(n4248) );
  NANDN U6282 ( .A(n4249), .B(n4248), .Z(n4251) );
  XNOR U6283 ( .A(n4249), .B(n4248), .Z(n4387) );
  AND U6284 ( .A(a[23]), .B(b[54]), .Z(n4386) );
  NAND U6285 ( .A(n4387), .B(n4386), .Z(n4250) );
  AND U6286 ( .A(n4251), .B(n4250), .Z(n4383) );
  XNOR U6287 ( .A(n4253), .B(n4252), .Z(n4382) );
  NANDN U6288 ( .A(n4383), .B(n4382), .Z(n4254) );
  AND U6289 ( .A(n4255), .B(n4254), .Z(n4381) );
  XNOR U6290 ( .A(n4257), .B(n4256), .Z(n4380) );
  NANDN U6291 ( .A(n4381), .B(n4380), .Z(n4258) );
  AND U6292 ( .A(n4259), .B(n4258), .Z(n4262) );
  XOR U6293 ( .A(n4261), .B(n4260), .Z(n4263) );
  NAND U6294 ( .A(n4262), .B(n4263), .Z(n4265) );
  AND U6295 ( .A(a[26]), .B(b[54]), .Z(n4379) );
  XOR U6296 ( .A(n4263), .B(n4262), .Z(n4378) );
  NANDN U6297 ( .A(n4379), .B(n4378), .Z(n4264) );
  AND U6298 ( .A(n4265), .B(n4264), .Z(n4534) );
  XNOR U6299 ( .A(n4267), .B(n4266), .Z(n4533) );
  NAND U6300 ( .A(n4534), .B(n4533), .Z(n4268) );
  AND U6301 ( .A(n4269), .B(n4268), .Z(n4377) );
  XNOR U6302 ( .A(n4271), .B(n4270), .Z(n4376) );
  NANDN U6303 ( .A(n4377), .B(n4376), .Z(n4272) );
  AND U6304 ( .A(n4273), .B(n4272), .Z(n4375) );
  XNOR U6305 ( .A(n4275), .B(n4274), .Z(n4374) );
  NANDN U6306 ( .A(n4375), .B(n4374), .Z(n4276) );
  AND U6307 ( .A(n4277), .B(n4276), .Z(n4546) );
  XNOR U6308 ( .A(n4279), .B(n4278), .Z(n4545) );
  NANDN U6309 ( .A(n4546), .B(n4545), .Z(n4280) );
  AND U6310 ( .A(n4281), .B(n4280), .Z(n4282) );
  NANDN U6311 ( .A(n4283), .B(n4282), .Z(n4287) );
  XNOR U6312 ( .A(n4283), .B(n4282), .Z(n4372) );
  XNOR U6313 ( .A(n4285), .B(n4284), .Z(n4373) );
  NAND U6314 ( .A(n4372), .B(n4373), .Z(n4286) );
  AND U6315 ( .A(n4287), .B(n4286), .Z(n4291) );
  NANDN U6316 ( .A(n4290), .B(n4291), .Z(n4293) );
  XOR U6317 ( .A(n4289), .B(n4288), .Z(n4558) );
  XNOR U6318 ( .A(n4291), .B(n4290), .Z(n4557) );
  NANDN U6319 ( .A(n4558), .B(n4557), .Z(n4292) );
  AND U6320 ( .A(n4293), .B(n4292), .Z(n4297) );
  AND U6321 ( .A(a[33]), .B(b[54]), .Z(n4296) );
  NANDN U6322 ( .A(n4297), .B(n4296), .Z(n4299) );
  XNOR U6323 ( .A(n4295), .B(n4294), .Z(n4564) );
  XNOR U6324 ( .A(n4297), .B(n4296), .Z(n4563) );
  NAND U6325 ( .A(n4564), .B(n4563), .Z(n4298) );
  AND U6326 ( .A(n4299), .B(n4298), .Z(n4303) );
  AND U6327 ( .A(a[34]), .B(b[54]), .Z(n4302) );
  NANDN U6328 ( .A(n4303), .B(n4302), .Z(n4305) );
  XNOR U6329 ( .A(n4301), .B(n4300), .Z(n4568) );
  XNOR U6330 ( .A(n4303), .B(n4302), .Z(n4567) );
  NAND U6331 ( .A(n4568), .B(n4567), .Z(n4304) );
  AND U6332 ( .A(n4305), .B(n4304), .Z(n4308) );
  NANDN U6333 ( .A(n4309), .B(n4308), .Z(n4311) );
  XOR U6334 ( .A(n4307), .B(n4306), .Z(n4576) );
  XNOR U6335 ( .A(n4309), .B(n4308), .Z(n4575) );
  NANDN U6336 ( .A(n4576), .B(n4575), .Z(n4310) );
  AND U6337 ( .A(n4311), .B(n4310), .Z(n4315) );
  NANDN U6338 ( .A(n4314), .B(n4315), .Z(n4317) );
  XOR U6339 ( .A(n4313), .B(n4312), .Z(n4582) );
  XNOR U6340 ( .A(n4315), .B(n4314), .Z(n4581) );
  NANDN U6341 ( .A(n4582), .B(n4581), .Z(n4316) );
  AND U6342 ( .A(n4317), .B(n4316), .Z(n4319) );
  NANDN U6343 ( .A(n4318), .B(n4319), .Z(n4323) );
  XNOR U6344 ( .A(n4321), .B(n4320), .Z(n4588) );
  NAND U6345 ( .A(n4587), .B(n4588), .Z(n4322) );
  NAND U6346 ( .A(n4323), .B(n4322), .Z(n4327) );
  NANDN U6347 ( .A(n4326), .B(n4327), .Z(n4329) );
  XOR U6348 ( .A(n4325), .B(n4324), .Z(n4593) );
  NANDN U6349 ( .A(n4593), .B(n4594), .Z(n4328) );
  AND U6350 ( .A(n4329), .B(n4328), .Z(n4333) );
  NANDN U6351 ( .A(n4332), .B(n4333), .Z(n4335) );
  XOR U6352 ( .A(n4331), .B(n4330), .Z(n4599) );
  NANDN U6353 ( .A(n4599), .B(n4600), .Z(n4334) );
  AND U6354 ( .A(n4335), .B(n4334), .Z(n4337) );
  NANDN U6355 ( .A(n4336), .B(n4337), .Z(n4341) );
  XNOR U6356 ( .A(n4339), .B(n4338), .Z(n4606) );
  NAND U6357 ( .A(n4605), .B(n4606), .Z(n4340) );
  NAND U6358 ( .A(n4341), .B(n4340), .Z(n4343) );
  NANDN U6359 ( .A(n4342), .B(n4343), .Z(n4347) );
  XNOR U6360 ( .A(n4345), .B(n4344), .Z(n4612) );
  NAND U6361 ( .A(n4611), .B(n4612), .Z(n4346) );
  NAND U6362 ( .A(n4347), .B(n4346), .Z(n4350) );
  AND U6363 ( .A(a[42]), .B(b[54]), .Z(n4351) );
  NANDN U6364 ( .A(n4350), .B(n4351), .Z(n4353) );
  XOR U6365 ( .A(n4349), .B(n4348), .Z(n4617) );
  NANDN U6366 ( .A(n4617), .B(n4618), .Z(n4352) );
  AND U6367 ( .A(n4353), .B(n4352), .Z(n4355) );
  NANDN U6368 ( .A(n4354), .B(n4355), .Z(n4359) );
  XNOR U6369 ( .A(n4357), .B(n4356), .Z(n4624) );
  NAND U6370 ( .A(n4623), .B(n4624), .Z(n4358) );
  NAND U6371 ( .A(n4359), .B(n4358), .Z(n4361) );
  NANDN U6372 ( .A(n4360), .B(n4361), .Z(n4365) );
  NAND U6373 ( .A(n4628), .B(n4627), .Z(n4364) );
  NAND U6374 ( .A(n4365), .B(n4364), .Z(n4368) );
  AND U6375 ( .A(a[45]), .B(b[54]), .Z(n4369) );
  NANDN U6376 ( .A(n4368), .B(n4369), .Z(n4371) );
  XOR U6377 ( .A(n4367), .B(n4366), .Z(n4635) );
  NANDN U6378 ( .A(n4635), .B(n4636), .Z(n4370) );
  AND U6379 ( .A(n4371), .B(n4370), .Z(n10124) );
  XNOR U6380 ( .A(n10126), .B(n10127), .Z(n10180) );
  AND U6381 ( .A(a[47]), .B(b[53]), .Z(n10178) );
  NAND U6382 ( .A(a[36]), .B(b[53]), .Z(n4573) );
  AND U6383 ( .A(a[35]), .B(b[53]), .Z(n4570) );
  AND U6384 ( .A(a[32]), .B(b[53]), .Z(n4551) );
  XNOR U6385 ( .A(n4373), .B(n4372), .Z(n4552) );
  NAND U6386 ( .A(n4551), .B(n4552), .Z(n4554) );
  XOR U6387 ( .A(n4375), .B(n4374), .Z(n4542) );
  AND U6388 ( .A(a[29]), .B(b[53]), .Z(n4538) );
  XOR U6389 ( .A(n4377), .B(n4376), .Z(n4537) );
  NANDN U6390 ( .A(n4538), .B(n4537), .Z(n4540) );
  XOR U6391 ( .A(n4379), .B(n4378), .Z(n4530) );
  AND U6392 ( .A(a[27]), .B(b[53]), .Z(n4529) );
  NAND U6393 ( .A(n4530), .B(n4529), .Z(n4532) );
  NAND U6394 ( .A(a[26]), .B(b[53]), .Z(n4525) );
  XNOR U6395 ( .A(n4381), .B(n4380), .Z(n4526) );
  NANDN U6396 ( .A(n4525), .B(n4526), .Z(n4528) );
  NAND U6397 ( .A(a[25]), .B(b[53]), .Z(n4384) );
  XNOR U6398 ( .A(n4383), .B(n4382), .Z(n4385) );
  NANDN U6399 ( .A(n4384), .B(n4385), .Z(n4524) );
  XOR U6400 ( .A(n4385), .B(n4384), .Z(n4798) );
  XOR U6401 ( .A(n4387), .B(n4386), .Z(n4520) );
  XOR U6402 ( .A(n4389), .B(n4388), .Z(n4516) );
  NAND U6403 ( .A(a[20]), .B(b[53]), .Z(n4392) );
  XNOR U6404 ( .A(n4391), .B(n4390), .Z(n4393) );
  NANDN U6405 ( .A(n4392), .B(n4393), .Z(n4502) );
  XOR U6406 ( .A(n4393), .B(n4392), .Z(n4661) );
  XOR U6407 ( .A(n4395), .B(n4394), .Z(n4498) );
  XOR U6408 ( .A(n4397), .B(n4396), .Z(n4493) );
  XOR U6409 ( .A(n4399), .B(n4398), .Z(n4483) );
  AND U6410 ( .A(a[16]), .B(b[53]), .Z(n4484) );
  NANDN U6411 ( .A(n4483), .B(n4484), .Z(n4486) );
  XOR U6412 ( .A(n4401), .B(n4400), .Z(n4467) );
  AND U6413 ( .A(a[13]), .B(b[53]), .Z(n4468) );
  NANDN U6414 ( .A(n4467), .B(n4468), .Z(n4470) );
  XOR U6415 ( .A(n4403), .B(n4402), .Z(n4463) );
  AND U6416 ( .A(a[12]), .B(b[53]), .Z(n4464) );
  NANDN U6417 ( .A(n4463), .B(n4464), .Z(n4466) );
  XOR U6418 ( .A(n4407), .B(n4406), .Z(n4449) );
  NAND U6419 ( .A(a[7]), .B(b[53]), .Z(n4439) );
  XOR U6420 ( .A(n4409), .B(n4408), .Z(n4440) );
  NANDN U6421 ( .A(n4439), .B(n4440), .Z(n4442) );
  NAND U6422 ( .A(a[0]), .B(b[53]), .Z(n4951) );
  AND U6423 ( .A(a[1]), .B(b[54]), .Z(n4412) );
  NANDN U6424 ( .A(n4951), .B(n4412), .Z(n4681) );
  NANDN U6425 ( .A(n4681), .B(n4410), .Z(n4414) );
  AND U6426 ( .A(a[2]), .B(b[53]), .Z(n4687) );
  NANDN U6427 ( .A(n4686), .B(n4687), .Z(n4413) );
  AND U6428 ( .A(n4414), .B(n4413), .Z(n4417) );
  AND U6429 ( .A(a[3]), .B(b[53]), .Z(n4418) );
  NANDN U6430 ( .A(n4417), .B(n4418), .Z(n4420) );
  XOR U6431 ( .A(n4416), .B(n4415), .Z(n4692) );
  NANDN U6432 ( .A(n4692), .B(n4693), .Z(n4419) );
  AND U6433 ( .A(n4420), .B(n4419), .Z(n4423) );
  NANDN U6434 ( .A(n4423), .B(n4424), .Z(n4426) );
  NAND U6435 ( .A(a[4]), .B(b[53]), .Z(n4700) );
  NANDN U6436 ( .A(n4700), .B(n4701), .Z(n4425) );
  AND U6437 ( .A(n4426), .B(n4425), .Z(n4427) );
  AND U6438 ( .A(a[5]), .B(b[53]), .Z(n4428) );
  NANDN U6439 ( .A(n4427), .B(n4428), .Z(n4432) );
  XOR U6440 ( .A(n4430), .B(n4429), .Z(n4704) );
  NAND U6441 ( .A(n4705), .B(n4704), .Z(n4431) );
  AND U6442 ( .A(n4432), .B(n4431), .Z(n4435) );
  XOR U6443 ( .A(n4434), .B(n4433), .Z(n4436) );
  NANDN U6444 ( .A(n4435), .B(n4436), .Z(n4438) );
  AND U6445 ( .A(a[6]), .B(b[53]), .Z(n4680) );
  NAND U6446 ( .A(n4680), .B(n4679), .Z(n4437) );
  AND U6447 ( .A(n4438), .B(n4437), .Z(n4716) );
  NANDN U6448 ( .A(n4716), .B(n4717), .Z(n4441) );
  AND U6449 ( .A(n4442), .B(n4441), .Z(n4443) );
  AND U6450 ( .A(a[8]), .B(b[53]), .Z(n4444) );
  NANDN U6451 ( .A(n4443), .B(n4444), .Z(n4448) );
  NAND U6452 ( .A(n4678), .B(n4677), .Z(n4447) );
  AND U6453 ( .A(n4448), .B(n4447), .Z(n4450) );
  NANDN U6454 ( .A(n4449), .B(n4450), .Z(n4452) );
  AND U6455 ( .A(a[9]), .B(b[53]), .Z(n4724) );
  NANDN U6456 ( .A(n4724), .B(n4725), .Z(n4451) );
  AND U6457 ( .A(n4452), .B(n4451), .Z(n4456) );
  NAND U6458 ( .A(n4456), .B(n4455), .Z(n4458) );
  AND U6459 ( .A(a[10]), .B(b[53]), .Z(n4676) );
  XOR U6460 ( .A(n4456), .B(n4455), .Z(n4675) );
  NAND U6461 ( .A(n4676), .B(n4675), .Z(n4457) );
  NAND U6462 ( .A(n4458), .B(n4457), .Z(n4459) );
  NAND U6463 ( .A(n4460), .B(n4459), .Z(n4462) );
  XOR U6464 ( .A(n4460), .B(n4459), .Z(n4735) );
  AND U6465 ( .A(a[11]), .B(b[53]), .Z(n4734) );
  NAND U6466 ( .A(n4735), .B(n4734), .Z(n4461) );
  AND U6467 ( .A(n4462), .B(n4461), .Z(n4741) );
  XNOR U6468 ( .A(n4464), .B(n4463), .Z(n4740) );
  NANDN U6469 ( .A(n4741), .B(n4740), .Z(n4465) );
  AND U6470 ( .A(n4466), .B(n4465), .Z(n4749) );
  XNOR U6471 ( .A(n4468), .B(n4467), .Z(n4748) );
  NANDN U6472 ( .A(n4749), .B(n4748), .Z(n4469) );
  AND U6473 ( .A(n4470), .B(n4469), .Z(n4474) );
  XNOR U6474 ( .A(n4472), .B(n4471), .Z(n4473) );
  NANDN U6475 ( .A(n4474), .B(n4473), .Z(n4476) );
  XNOR U6476 ( .A(n4474), .B(n4473), .Z(n4674) );
  AND U6477 ( .A(a[14]), .B(b[53]), .Z(n4673) );
  NAND U6478 ( .A(n4674), .B(n4673), .Z(n4475) );
  AND U6479 ( .A(n4476), .B(n4475), .Z(n4480) );
  XNOR U6480 ( .A(n4478), .B(n4477), .Z(n4479) );
  NANDN U6481 ( .A(n4480), .B(n4479), .Z(n4482) );
  XNOR U6482 ( .A(n4480), .B(n4479), .Z(n4670) );
  AND U6483 ( .A(a[15]), .B(b[53]), .Z(n4669) );
  NAND U6484 ( .A(n4670), .B(n4669), .Z(n4481) );
  AND U6485 ( .A(n4482), .B(n4481), .Z(n4666) );
  XNOR U6486 ( .A(n4484), .B(n4483), .Z(n4665) );
  NANDN U6487 ( .A(n4666), .B(n4665), .Z(n4485) );
  AND U6488 ( .A(n4486), .B(n4485), .Z(n4490) );
  XNOR U6489 ( .A(n4488), .B(n4487), .Z(n4489) );
  NANDN U6490 ( .A(n4490), .B(n4489), .Z(n4492) );
  NAND U6491 ( .A(a[17]), .B(b[53]), .Z(n4760) );
  XNOR U6492 ( .A(n4490), .B(n4489), .Z(n4761) );
  NANDN U6493 ( .A(n4760), .B(n4761), .Z(n4491) );
  AND U6494 ( .A(n4492), .B(n4491), .Z(n4494) );
  NANDN U6495 ( .A(n4493), .B(n4494), .Z(n4496) );
  XOR U6496 ( .A(n4494), .B(n4493), .Z(n4663) );
  AND U6497 ( .A(a[18]), .B(b[53]), .Z(n4664) );
  OR U6498 ( .A(n4663), .B(n4664), .Z(n4495) );
  AND U6499 ( .A(n4496), .B(n4495), .Z(n4497) );
  NANDN U6500 ( .A(n4498), .B(n4497), .Z(n4500) );
  NAND U6501 ( .A(a[19]), .B(b[53]), .Z(n4770) );
  XNOR U6502 ( .A(n4498), .B(n4497), .Z(n4771) );
  NANDN U6503 ( .A(n4770), .B(n4771), .Z(n4499) );
  AND U6504 ( .A(n4500), .B(n4499), .Z(n4662) );
  OR U6505 ( .A(n4661), .B(n4662), .Z(n4501) );
  AND U6506 ( .A(n4502), .B(n4501), .Z(n4506) );
  XNOR U6507 ( .A(n4504), .B(n4503), .Z(n4505) );
  NANDN U6508 ( .A(n4506), .B(n4505), .Z(n4508) );
  NAND U6509 ( .A(a[21]), .B(b[53]), .Z(n4657) );
  XNOR U6510 ( .A(n4506), .B(n4505), .Z(n4658) );
  NANDN U6511 ( .A(n4657), .B(n4658), .Z(n4507) );
  AND U6512 ( .A(n4508), .B(n4507), .Z(n4512) );
  XNOR U6513 ( .A(n4510), .B(n4509), .Z(n4511) );
  NANDN U6514 ( .A(n4512), .B(n4511), .Z(n4514) );
  NAND U6515 ( .A(a[22]), .B(b[53]), .Z(n4782) );
  XNOR U6516 ( .A(n4512), .B(n4511), .Z(n4783) );
  NANDN U6517 ( .A(n4782), .B(n4783), .Z(n4513) );
  AND U6518 ( .A(n4514), .B(n4513), .Z(n4515) );
  NANDN U6519 ( .A(n4516), .B(n4515), .Z(n4518) );
  XOR U6520 ( .A(n4516), .B(n4515), .Z(n4655) );
  AND U6521 ( .A(a[23]), .B(b[53]), .Z(n4656) );
  OR U6522 ( .A(n4655), .B(n4656), .Z(n4517) );
  NAND U6523 ( .A(n4518), .B(n4517), .Z(n4519) );
  NANDN U6524 ( .A(n4520), .B(n4519), .Z(n4522) );
  XOR U6525 ( .A(n4520), .B(n4519), .Z(n4792) );
  AND U6526 ( .A(a[24]), .B(b[53]), .Z(n4793) );
  OR U6527 ( .A(n4792), .B(n4793), .Z(n4521) );
  AND U6528 ( .A(n4522), .B(n4521), .Z(n4799) );
  NANDN U6529 ( .A(n4798), .B(n4799), .Z(n4523) );
  AND U6530 ( .A(n4524), .B(n4523), .Z(n4654) );
  XNOR U6531 ( .A(n4526), .B(n4525), .Z(n4653) );
  NANDN U6532 ( .A(n4654), .B(n4653), .Z(n4527) );
  AND U6533 ( .A(n4528), .B(n4527), .Z(n4652) );
  XOR U6534 ( .A(n4530), .B(n4529), .Z(n4651) );
  NANDN U6535 ( .A(n4652), .B(n4651), .Z(n4531) );
  AND U6536 ( .A(n4532), .B(n4531), .Z(n4536) );
  AND U6537 ( .A(a[28]), .B(b[53]), .Z(n4535) );
  XOR U6538 ( .A(n4534), .B(n4533), .Z(n4647) );
  XNOR U6539 ( .A(n4536), .B(n4535), .Z(n4648) );
  XNOR U6540 ( .A(n4538), .B(n4537), .Z(n4645) );
  NAND U6541 ( .A(n4646), .B(n4645), .Z(n4539) );
  NAND U6542 ( .A(n4540), .B(n4539), .Z(n4541) );
  NAND U6543 ( .A(n4542), .B(n4541), .Z(n4544) );
  AND U6544 ( .A(a[30]), .B(b[53]), .Z(n4644) );
  XOR U6545 ( .A(n4542), .B(n4541), .Z(n4643) );
  NANDN U6546 ( .A(n4644), .B(n4643), .Z(n4543) );
  NAND U6547 ( .A(n4544), .B(n4543), .Z(n4547) );
  XNOR U6548 ( .A(n4546), .B(n4545), .Z(n4548) );
  NANDN U6549 ( .A(n4547), .B(n4548), .Z(n4550) );
  NAND U6550 ( .A(a[31]), .B(b[53]), .Z(n4822) );
  XNOR U6551 ( .A(n4548), .B(n4547), .Z(n4823) );
  NANDN U6552 ( .A(n4822), .B(n4823), .Z(n4549) );
  AND U6553 ( .A(n4550), .B(n4549), .Z(n4642) );
  XOR U6554 ( .A(n4552), .B(n4551), .Z(n4641) );
  NANDN U6555 ( .A(n4642), .B(n4641), .Z(n4553) );
  AND U6556 ( .A(n4554), .B(n4553), .Z(n4556) );
  AND U6557 ( .A(a[33]), .B(b[53]), .Z(n4555) );
  NANDN U6558 ( .A(n4556), .B(n4555), .Z(n4560) );
  XNOR U6559 ( .A(n4556), .B(n4555), .Z(n4640) );
  XNOR U6560 ( .A(n4558), .B(n4557), .Z(n4639) );
  NAND U6561 ( .A(n4640), .B(n4639), .Z(n4559) );
  AND U6562 ( .A(n4560), .B(n4559), .Z(n4562) );
  AND U6563 ( .A(a[34]), .B(b[53]), .Z(n4561) );
  NANDN U6564 ( .A(n4562), .B(n4561), .Z(n4566) );
  XNOR U6565 ( .A(n4562), .B(n4561), .Z(n4837) );
  XOR U6566 ( .A(n4564), .B(n4563), .Z(n4836) );
  NAND U6567 ( .A(n4837), .B(n4836), .Z(n4565) );
  AND U6568 ( .A(n4566), .B(n4565), .Z(n4569) );
  NANDN U6569 ( .A(n4570), .B(n4569), .Z(n4572) );
  XOR U6570 ( .A(n4568), .B(n4567), .Z(n4845) );
  XNOR U6571 ( .A(n4570), .B(n4569), .Z(n4844) );
  NANDN U6572 ( .A(n4845), .B(n4844), .Z(n4571) );
  AND U6573 ( .A(n4572), .B(n4571), .Z(n4574) );
  NANDN U6574 ( .A(n4573), .B(n4574), .Z(n4578) );
  XNOR U6575 ( .A(n4574), .B(n4573), .Z(n4848) );
  XOR U6576 ( .A(n4576), .B(n4575), .Z(n4849) );
  NAND U6577 ( .A(n4848), .B(n4849), .Z(n4577) );
  AND U6578 ( .A(n4578), .B(n4577), .Z(n4580) );
  AND U6579 ( .A(a[37]), .B(b[53]), .Z(n4579) );
  NANDN U6580 ( .A(n4580), .B(n4579), .Z(n4584) );
  XNOR U6581 ( .A(n4580), .B(n4579), .Z(n4855) );
  XNOR U6582 ( .A(n4582), .B(n4581), .Z(n4854) );
  NAND U6583 ( .A(n4855), .B(n4854), .Z(n4583) );
  AND U6584 ( .A(n4584), .B(n4583), .Z(n4585) );
  AND U6585 ( .A(a[38]), .B(b[53]), .Z(n4586) );
  NANDN U6586 ( .A(n4585), .B(n4586), .Z(n4590) );
  XNOR U6587 ( .A(n4588), .B(n4587), .Z(n4863) );
  NAND U6588 ( .A(n4862), .B(n4863), .Z(n4589) );
  AND U6589 ( .A(n4590), .B(n4589), .Z(n4591) );
  AND U6590 ( .A(a[39]), .B(b[53]), .Z(n4592) );
  NANDN U6591 ( .A(n4591), .B(n4592), .Z(n4596) );
  NAND U6592 ( .A(n4866), .B(n4867), .Z(n4595) );
  AND U6593 ( .A(n4596), .B(n4595), .Z(n4597) );
  AND U6594 ( .A(a[40]), .B(b[53]), .Z(n4598) );
  NANDN U6595 ( .A(n4597), .B(n4598), .Z(n4602) );
  NAND U6596 ( .A(n4873), .B(n4872), .Z(n4601) );
  AND U6597 ( .A(n4602), .B(n4601), .Z(n4603) );
  AND U6598 ( .A(a[41]), .B(b[53]), .Z(n4604) );
  NANDN U6599 ( .A(n4603), .B(n4604), .Z(n4608) );
  XNOR U6600 ( .A(n4606), .B(n4605), .Z(n4881) );
  NAND U6601 ( .A(n4880), .B(n4881), .Z(n4607) );
  AND U6602 ( .A(n4608), .B(n4607), .Z(n4609) );
  AND U6603 ( .A(a[42]), .B(b[53]), .Z(n4610) );
  NANDN U6604 ( .A(n4609), .B(n4610), .Z(n4614) );
  XNOR U6605 ( .A(n4612), .B(n4611), .Z(n4887) );
  NAND U6606 ( .A(n4886), .B(n4887), .Z(n4613) );
  AND U6607 ( .A(n4614), .B(n4613), .Z(n4615) );
  AND U6608 ( .A(a[43]), .B(b[53]), .Z(n4616) );
  NANDN U6609 ( .A(n4615), .B(n4616), .Z(n4620) );
  NAND U6610 ( .A(n4891), .B(n4890), .Z(n4619) );
  AND U6611 ( .A(n4620), .B(n4619), .Z(n4621) );
  AND U6612 ( .A(a[44]), .B(b[53]), .Z(n4622) );
  NANDN U6613 ( .A(n4621), .B(n4622), .Z(n4626) );
  XNOR U6614 ( .A(n4624), .B(n4623), .Z(n4899) );
  NAND U6615 ( .A(n4898), .B(n4899), .Z(n4625) );
  AND U6616 ( .A(n4626), .B(n4625), .Z(n4629) );
  AND U6617 ( .A(a[45]), .B(b[53]), .Z(n4630) );
  NANDN U6618 ( .A(n4629), .B(n4630), .Z(n4632) );
  XOR U6619 ( .A(n4628), .B(n4627), .Z(n4902) );
  NANDN U6620 ( .A(n4902), .B(n4903), .Z(n4631) );
  AND U6621 ( .A(n4632), .B(n4631), .Z(n4633) );
  AND U6622 ( .A(a[46]), .B(b[53]), .Z(n4634) );
  NANDN U6623 ( .A(n4633), .B(n4634), .Z(n4638) );
  NAND U6624 ( .A(n4909), .B(n4908), .Z(n4637) );
  AND U6625 ( .A(n4638), .B(n4637), .Z(n10179) );
  XNOR U6626 ( .A(n10180), .B(n10181), .Z(n10186) );
  AND U6627 ( .A(a[48]), .B(b[52]), .Z(n10185) );
  AND U6628 ( .A(a[47]), .B(b[52]), .Z(n4910) );
  AND U6629 ( .A(a[45]), .B(b[52]), .Z(n4896) );
  AND U6630 ( .A(a[44]), .B(b[52]), .Z(n4892) );
  AND U6631 ( .A(a[43]), .B(b[52]), .Z(n4884) );
  AND U6632 ( .A(a[42]), .B(b[52]), .Z(n4878) );
  AND U6633 ( .A(a[41]), .B(b[52]), .Z(n4874) );
  NAND U6634 ( .A(a[40]), .B(b[52]), .Z(n4868) );
  AND U6635 ( .A(a[39]), .B(b[52]), .Z(n4860) );
  AND U6636 ( .A(a[38]), .B(b[52]), .Z(n4857) );
  NAND U6637 ( .A(a[37]), .B(b[52]), .Z(n4850) );
  AND U6638 ( .A(a[36]), .B(b[52]), .Z(n4843) );
  AND U6639 ( .A(a[35]), .B(b[52]), .Z(n4839) );
  AND U6640 ( .A(a[34]), .B(b[52]), .Z(n4833) );
  XOR U6641 ( .A(n4640), .B(n4639), .Z(n4832) );
  NAND U6642 ( .A(n4833), .B(n4832), .Z(n4835) );
  NAND U6643 ( .A(a[33]), .B(b[52]), .Z(n4828) );
  XNOR U6644 ( .A(n4642), .B(n4641), .Z(n4829) );
  NANDN U6645 ( .A(n4828), .B(n4829), .Z(n4831) );
  AND U6646 ( .A(a[31]), .B(b[52]), .Z(n4818) );
  XOR U6647 ( .A(n4644), .B(n4643), .Z(n4819) );
  NAND U6648 ( .A(n4818), .B(n4819), .Z(n4821) );
  XOR U6649 ( .A(n4646), .B(n4645), .Z(n4815) );
  AND U6650 ( .A(a[30]), .B(b[52]), .Z(n4814) );
  NANDN U6651 ( .A(n4815), .B(n4814), .Z(n4817) );
  NAND U6652 ( .A(a[29]), .B(b[52]), .Z(n4649) );
  XOR U6653 ( .A(n4648), .B(n4647), .Z(n4650) );
  NANDN U6654 ( .A(n4649), .B(n4650), .Z(n4813) );
  XOR U6655 ( .A(n4650), .B(n4649), .Z(n4922) );
  NAND U6656 ( .A(a[28]), .B(b[52]), .Z(n4808) );
  XNOR U6657 ( .A(n4652), .B(n4651), .Z(n4809) );
  NANDN U6658 ( .A(n4808), .B(n4809), .Z(n4811) );
  NAND U6659 ( .A(a[27]), .B(b[52]), .Z(n4804) );
  XNOR U6660 ( .A(n4654), .B(n4653), .Z(n4805) );
  NANDN U6661 ( .A(n4804), .B(n4805), .Z(n4807) );
  XOR U6662 ( .A(n4656), .B(n4655), .Z(n4789) );
  AND U6663 ( .A(a[24]), .B(b[52]), .Z(n4788) );
  NANDN U6664 ( .A(n4789), .B(n4788), .Z(n4791) );
  NAND U6665 ( .A(a[22]), .B(b[52]), .Z(n4659) );
  XNOR U6666 ( .A(n4658), .B(n4657), .Z(n4660) );
  NANDN U6667 ( .A(n4659), .B(n4660), .Z(n4781) );
  XOR U6668 ( .A(n4660), .B(n4659), .Z(n5053) );
  XOR U6669 ( .A(n4662), .B(n4661), .Z(n4777) );
  XOR U6670 ( .A(n4664), .B(n4663), .Z(n4767) );
  AND U6671 ( .A(a[19]), .B(b[52]), .Z(n4766) );
  NANDN U6672 ( .A(n4767), .B(n4766), .Z(n4769) );
  XOR U6673 ( .A(n4666), .B(n4665), .Z(n4667) );
  AND U6674 ( .A(a[17]), .B(b[52]), .Z(n4668) );
  NANDN U6675 ( .A(n4667), .B(n4668), .Z(n4759) );
  XNOR U6676 ( .A(n4668), .B(n4667), .Z(n4935) );
  AND U6677 ( .A(a[16]), .B(b[52]), .Z(n4672) );
  XNOR U6678 ( .A(n4670), .B(n4669), .Z(n4671) );
  NANDN U6679 ( .A(n4672), .B(n4671), .Z(n4757) );
  XOR U6680 ( .A(n4672), .B(n4671), .Z(n4936) );
  XOR U6681 ( .A(n4674), .B(n4673), .Z(n4753) );
  NAND U6682 ( .A(a[13]), .B(b[52]), .Z(n4742) );
  XOR U6683 ( .A(n4676), .B(n4675), .Z(n4730) );
  XOR U6684 ( .A(n4678), .B(n4677), .Z(n4720) );
  NAND U6685 ( .A(a[7]), .B(b[52]), .Z(n4710) );
  XOR U6686 ( .A(n4680), .B(n4679), .Z(n4711) );
  NANDN U6687 ( .A(n4710), .B(n4711), .Z(n4713) );
  NAND U6688 ( .A(a[0]), .B(b[52]), .Z(n5238) );
  AND U6689 ( .A(a[1]), .B(b[53]), .Z(n4683) );
  NANDN U6690 ( .A(n5238), .B(n4683), .Z(n4950) );
  NANDN U6691 ( .A(n4950), .B(n4681), .Z(n4685) );
  AND U6692 ( .A(a[2]), .B(b[52]), .Z(n4956) );
  NANDN U6693 ( .A(n4955), .B(n4956), .Z(n4684) );
  AND U6694 ( .A(n4685), .B(n4684), .Z(n4688) );
  AND U6695 ( .A(a[3]), .B(b[52]), .Z(n4689) );
  NANDN U6696 ( .A(n4688), .B(n4689), .Z(n4691) );
  XOR U6697 ( .A(n4687), .B(n4686), .Z(n4961) );
  NANDN U6698 ( .A(n4961), .B(n4962), .Z(n4690) );
  AND U6699 ( .A(n4691), .B(n4690), .Z(n4694) );
  NANDN U6700 ( .A(n4694), .B(n4695), .Z(n4697) );
  NAND U6701 ( .A(a[4]), .B(b[52]), .Z(n4969) );
  NANDN U6702 ( .A(n4969), .B(n4970), .Z(n4696) );
  AND U6703 ( .A(n4697), .B(n4696), .Z(n4698) );
  AND U6704 ( .A(a[5]), .B(b[52]), .Z(n4699) );
  NANDN U6705 ( .A(n4698), .B(n4699), .Z(n4703) );
  NAND U6706 ( .A(n4974), .B(n4973), .Z(n4702) );
  AND U6707 ( .A(n4703), .B(n4702), .Z(n4706) );
  XOR U6708 ( .A(n4705), .B(n4704), .Z(n4707) );
  NANDN U6709 ( .A(n4706), .B(n4707), .Z(n4709) );
  AND U6710 ( .A(a[6]), .B(b[52]), .Z(n4949) );
  NAND U6711 ( .A(n4949), .B(n4948), .Z(n4708) );
  AND U6712 ( .A(n4709), .B(n4708), .Z(n4985) );
  NANDN U6713 ( .A(n4985), .B(n4986), .Z(n4712) );
  AND U6714 ( .A(n4713), .B(n4712), .Z(n4714) );
  AND U6715 ( .A(a[8]), .B(b[52]), .Z(n4715) );
  NANDN U6716 ( .A(n4714), .B(n4715), .Z(n4719) );
  NAND U6717 ( .A(n4947), .B(n4946), .Z(n4718) );
  AND U6718 ( .A(n4719), .B(n4718), .Z(n4721) );
  NANDN U6719 ( .A(n4720), .B(n4721), .Z(n4723) );
  AND U6720 ( .A(a[9]), .B(b[52]), .Z(n4993) );
  NANDN U6721 ( .A(n4993), .B(n4994), .Z(n4722) );
  AND U6722 ( .A(n4723), .B(n4722), .Z(n4727) );
  NAND U6723 ( .A(n4727), .B(n4726), .Z(n4729) );
  XOR U6724 ( .A(n4727), .B(n4726), .Z(n4945) );
  AND U6725 ( .A(a[10]), .B(b[52]), .Z(n4944) );
  NAND U6726 ( .A(n4945), .B(n4944), .Z(n4728) );
  AND U6727 ( .A(n4729), .B(n4728), .Z(n4731) );
  NANDN U6728 ( .A(n4730), .B(n4731), .Z(n4733) );
  AND U6729 ( .A(a[11]), .B(b[52]), .Z(n5003) );
  NANDN U6730 ( .A(n5003), .B(n5004), .Z(n4732) );
  AND U6731 ( .A(n4733), .B(n4732), .Z(n4736) );
  XNOR U6732 ( .A(n4735), .B(n4734), .Z(n4737) );
  NANDN U6733 ( .A(n4736), .B(n4737), .Z(n4739) );
  AND U6734 ( .A(a[12]), .B(b[52]), .Z(n5009) );
  NANDN U6735 ( .A(n5009), .B(n5010), .Z(n4738) );
  AND U6736 ( .A(n4739), .B(n4738), .Z(n4743) );
  NANDN U6737 ( .A(n4742), .B(n4743), .Z(n4745) );
  XOR U6738 ( .A(n4741), .B(n4740), .Z(n4940) );
  XNOR U6739 ( .A(n4743), .B(n4742), .Z(n4941) );
  NANDN U6740 ( .A(n4940), .B(n4941), .Z(n4744) );
  AND U6741 ( .A(n4745), .B(n4744), .Z(n4747) );
  AND U6742 ( .A(a[14]), .B(b[52]), .Z(n4746) );
  NANDN U6743 ( .A(n4747), .B(n4746), .Z(n4751) );
  XNOR U6744 ( .A(n4747), .B(n4746), .Z(n4939) );
  XNOR U6745 ( .A(n4749), .B(n4748), .Z(n4938) );
  NAND U6746 ( .A(n4939), .B(n4938), .Z(n4750) );
  AND U6747 ( .A(n4751), .B(n4750), .Z(n4752) );
  NANDN U6748 ( .A(n4753), .B(n4752), .Z(n4755) );
  AND U6749 ( .A(a[15]), .B(b[52]), .Z(n5022) );
  XNOR U6750 ( .A(n4753), .B(n4752), .Z(n5021) );
  NANDN U6751 ( .A(n5022), .B(n5021), .Z(n4754) );
  AND U6752 ( .A(n4755), .B(n4754), .Z(n4937) );
  OR U6753 ( .A(n4936), .B(n4937), .Z(n4756) );
  AND U6754 ( .A(n4757), .B(n4756), .Z(n4934) );
  NAND U6755 ( .A(n4935), .B(n4934), .Z(n4758) );
  AND U6756 ( .A(n4759), .B(n4758), .Z(n4763) );
  XNOR U6757 ( .A(n4761), .B(n4760), .Z(n4762) );
  NANDN U6758 ( .A(n4763), .B(n4762), .Z(n4765) );
  NAND U6759 ( .A(a[18]), .B(b[52]), .Z(n5035) );
  XNOR U6760 ( .A(n4763), .B(n4762), .Z(n5036) );
  NANDN U6761 ( .A(n5035), .B(n5036), .Z(n4764) );
  AND U6762 ( .A(n4765), .B(n4764), .Z(n4931) );
  XNOR U6763 ( .A(n4767), .B(n4766), .Z(n4930) );
  NANDN U6764 ( .A(n4931), .B(n4930), .Z(n4768) );
  AND U6765 ( .A(n4769), .B(n4768), .Z(n4773) );
  XNOR U6766 ( .A(n4771), .B(n4770), .Z(n4772) );
  NANDN U6767 ( .A(n4773), .B(n4772), .Z(n4775) );
  NAND U6768 ( .A(a[20]), .B(b[52]), .Z(n5043) );
  XNOR U6769 ( .A(n4773), .B(n4772), .Z(n5044) );
  NANDN U6770 ( .A(n5043), .B(n5044), .Z(n4774) );
  AND U6771 ( .A(n4775), .B(n4774), .Z(n4776) );
  NANDN U6772 ( .A(n4777), .B(n4776), .Z(n4779) );
  AND U6773 ( .A(a[21]), .B(b[52]), .Z(n4929) );
  XNOR U6774 ( .A(n4777), .B(n4776), .Z(n4928) );
  NANDN U6775 ( .A(n4929), .B(n4928), .Z(n4778) );
  AND U6776 ( .A(n4779), .B(n4778), .Z(n5054) );
  NANDN U6777 ( .A(n5053), .B(n5054), .Z(n4780) );
  AND U6778 ( .A(n4781), .B(n4780), .Z(n4785) );
  AND U6779 ( .A(a[23]), .B(b[52]), .Z(n4784) );
  NANDN U6780 ( .A(n4785), .B(n4784), .Z(n4787) );
  XOR U6781 ( .A(n4783), .B(n4782), .Z(n5059) );
  XNOR U6782 ( .A(n4785), .B(n4784), .Z(n5060) );
  NANDN U6783 ( .A(n5059), .B(n5060), .Z(n4786) );
  AND U6784 ( .A(n4787), .B(n4786), .Z(n5066) );
  XNOR U6785 ( .A(n4789), .B(n4788), .Z(n5065) );
  NANDN U6786 ( .A(n5066), .B(n5065), .Z(n4790) );
  AND U6787 ( .A(n4791), .B(n4790), .Z(n4795) );
  AND U6788 ( .A(a[25]), .B(b[52]), .Z(n4794) );
  NANDN U6789 ( .A(n4795), .B(n4794), .Z(n4797) );
  XOR U6790 ( .A(n4793), .B(n4792), .Z(n5072) );
  XNOR U6791 ( .A(n4795), .B(n4794), .Z(n5071) );
  NANDN U6792 ( .A(n5072), .B(n5071), .Z(n4796) );
  AND U6793 ( .A(n4797), .B(n4796), .Z(n4801) );
  XNOR U6794 ( .A(n4799), .B(n4798), .Z(n4800) );
  NANDN U6795 ( .A(n4801), .B(n4800), .Z(n4803) );
  XNOR U6796 ( .A(n4801), .B(n4800), .Z(n4927) );
  AND U6797 ( .A(a[26]), .B(b[52]), .Z(n4926) );
  NAND U6798 ( .A(n4927), .B(n4926), .Z(n4802) );
  AND U6799 ( .A(n4803), .B(n4802), .Z(n4925) );
  XNOR U6800 ( .A(n4805), .B(n4804), .Z(n4924) );
  NANDN U6801 ( .A(n4925), .B(n4924), .Z(n4806) );
  AND U6802 ( .A(n4807), .B(n4806), .Z(n5086) );
  XNOR U6803 ( .A(n4809), .B(n4808), .Z(n5085) );
  NANDN U6804 ( .A(n5086), .B(n5085), .Z(n4810) );
  AND U6805 ( .A(n4811), .B(n4810), .Z(n4923) );
  OR U6806 ( .A(n4922), .B(n4923), .Z(n4812) );
  AND U6807 ( .A(n4813), .B(n4812), .Z(n5096) );
  XNOR U6808 ( .A(n4815), .B(n4814), .Z(n5095) );
  NANDN U6809 ( .A(n5096), .B(n5095), .Z(n4816) );
  AND U6810 ( .A(n4817), .B(n4816), .Z(n4921) );
  XOR U6811 ( .A(n4819), .B(n4818), .Z(n4920) );
  NANDN U6812 ( .A(n4921), .B(n4920), .Z(n4820) );
  AND U6813 ( .A(n4821), .B(n4820), .Z(n4825) );
  XNOR U6814 ( .A(n4823), .B(n4822), .Z(n4824) );
  NANDN U6815 ( .A(n4825), .B(n4824), .Z(n4827) );
  XNOR U6816 ( .A(n4825), .B(n4824), .Z(n4919) );
  AND U6817 ( .A(a[32]), .B(b[52]), .Z(n4918) );
  NAND U6818 ( .A(n4919), .B(n4918), .Z(n4826) );
  AND U6819 ( .A(n4827), .B(n4826), .Z(n4917) );
  XNOR U6820 ( .A(n4829), .B(n4828), .Z(n4916) );
  NANDN U6821 ( .A(n4917), .B(n4916), .Z(n4830) );
  AND U6822 ( .A(n4831), .B(n4830), .Z(n5114) );
  XOR U6823 ( .A(n4833), .B(n4832), .Z(n5113) );
  NANDN U6824 ( .A(n5114), .B(n5113), .Z(n4834) );
  AND U6825 ( .A(n4835), .B(n4834), .Z(n4838) );
  NANDN U6826 ( .A(n4839), .B(n4838), .Z(n4841) );
  XOR U6827 ( .A(n4837), .B(n4836), .Z(n4915) );
  XNOR U6828 ( .A(n4839), .B(n4838), .Z(n4914) );
  NANDN U6829 ( .A(n4915), .B(n4914), .Z(n4840) );
  NAND U6830 ( .A(n4841), .B(n4840), .Z(n4842) );
  NANDN U6831 ( .A(n4843), .B(n4842), .Z(n4847) );
  XNOR U6832 ( .A(n4843), .B(n4842), .Z(n5122) );
  XNOR U6833 ( .A(n4845), .B(n4844), .Z(n5121) );
  NAND U6834 ( .A(n5122), .B(n5121), .Z(n4846) );
  AND U6835 ( .A(n4847), .B(n4846), .Z(n4851) );
  NANDN U6836 ( .A(n4850), .B(n4851), .Z(n4853) );
  XOR U6837 ( .A(n4849), .B(n4848), .Z(n5130) );
  XNOR U6838 ( .A(n4851), .B(n4850), .Z(n5129) );
  NAND U6839 ( .A(n5130), .B(n5129), .Z(n4852) );
  AND U6840 ( .A(n4853), .B(n4852), .Z(n4856) );
  NANDN U6841 ( .A(n4857), .B(n4856), .Z(n4859) );
  XOR U6842 ( .A(n4855), .B(n4854), .Z(n5136) );
  XNOR U6843 ( .A(n4857), .B(n4856), .Z(n5135) );
  NANDN U6844 ( .A(n5136), .B(n5135), .Z(n4858) );
  NAND U6845 ( .A(n4859), .B(n4858), .Z(n4861) );
  NANDN U6846 ( .A(n4860), .B(n4861), .Z(n4865) );
  XNOR U6847 ( .A(n4863), .B(n4862), .Z(n5142) );
  NAND U6848 ( .A(n5141), .B(n5142), .Z(n4864) );
  AND U6849 ( .A(n4865), .B(n4864), .Z(n4869) );
  NANDN U6850 ( .A(n4868), .B(n4869), .Z(n4871) );
  XOR U6851 ( .A(n4867), .B(n4866), .Z(n5148) );
  NAND U6852 ( .A(n5148), .B(n5147), .Z(n4870) );
  AND U6853 ( .A(n4871), .B(n4870), .Z(n4875) );
  NANDN U6854 ( .A(n4874), .B(n4875), .Z(n4877) );
  XOR U6855 ( .A(n4873), .B(n4872), .Z(n5153) );
  NANDN U6856 ( .A(n5153), .B(n5154), .Z(n4876) );
  NAND U6857 ( .A(n4877), .B(n4876), .Z(n4879) );
  NANDN U6858 ( .A(n4878), .B(n4879), .Z(n4883) );
  XNOR U6859 ( .A(n4881), .B(n4880), .Z(n5160) );
  NAND U6860 ( .A(n5159), .B(n5160), .Z(n4882) );
  NAND U6861 ( .A(n4883), .B(n4882), .Z(n4885) );
  NANDN U6862 ( .A(n4884), .B(n4885), .Z(n4889) );
  XNOR U6863 ( .A(n4887), .B(n4886), .Z(n5166) );
  NAND U6864 ( .A(n5165), .B(n5166), .Z(n4888) );
  NAND U6865 ( .A(n4889), .B(n4888), .Z(n4893) );
  NANDN U6866 ( .A(n4892), .B(n4893), .Z(n4895) );
  XOR U6867 ( .A(n4891), .B(n4890), .Z(n5171) );
  NANDN U6868 ( .A(n5171), .B(n5172), .Z(n4894) );
  NAND U6869 ( .A(n4895), .B(n4894), .Z(n4897) );
  NANDN U6870 ( .A(n4896), .B(n4897), .Z(n4901) );
  XNOR U6871 ( .A(n4899), .B(n4898), .Z(n5178) );
  NAND U6872 ( .A(n5177), .B(n5178), .Z(n4900) );
  NAND U6873 ( .A(n4901), .B(n4900), .Z(n4904) );
  AND U6874 ( .A(a[46]), .B(b[52]), .Z(n4905) );
  NANDN U6875 ( .A(n4904), .B(n4905), .Z(n4907) );
  NAND U6876 ( .A(n5184), .B(n5183), .Z(n4906) );
  AND U6877 ( .A(n4907), .B(n4906), .Z(n4911) );
  NANDN U6878 ( .A(n4910), .B(n4911), .Z(n4913) );
  XOR U6879 ( .A(n4909), .B(n4908), .Z(n5189) );
  NANDN U6880 ( .A(n5189), .B(n5190), .Z(n4912) );
  NAND U6881 ( .A(n4913), .B(n4912), .Z(n10184) );
  XNOR U6882 ( .A(n10186), .B(n10187), .Z(n10192) );
  AND U6883 ( .A(a[49]), .B(b[51]), .Z(n10190) );
  AND U6884 ( .A(a[48]), .B(b[51]), .Z(n5187) );
  AND U6885 ( .A(a[42]), .B(b[51]), .Z(n5151) );
  AND U6886 ( .A(a[36]), .B(b[51]), .Z(n5117) );
  XOR U6887 ( .A(n4915), .B(n4914), .Z(n5118) );
  NAND U6888 ( .A(n5117), .B(n5118), .Z(n5120) );
  XNOR U6889 ( .A(n4917), .B(n4916), .Z(n5109) );
  XOR U6890 ( .A(n4919), .B(n4918), .Z(n5106) );
  NAND U6891 ( .A(a[32]), .B(b[51]), .Z(n5101) );
  XNOR U6892 ( .A(n4921), .B(n4920), .Z(n5102) );
  NANDN U6893 ( .A(n5101), .B(n5102), .Z(n5104) );
  XOR U6894 ( .A(n4923), .B(n4922), .Z(n5092) );
  XOR U6895 ( .A(n4925), .B(n4924), .Z(n5081) );
  XOR U6896 ( .A(n4927), .B(n4926), .Z(n5078) );
  XOR U6897 ( .A(n4929), .B(n4928), .Z(n5049) );
  NAND U6898 ( .A(a[20]), .B(b[51]), .Z(n4932) );
  XNOR U6899 ( .A(n4931), .B(n4930), .Z(n4933) );
  NANDN U6900 ( .A(n4932), .B(n4933), .Z(n5042) );
  XOR U6901 ( .A(n4933), .B(n4932), .Z(n5332) );
  XOR U6902 ( .A(n4935), .B(n4934), .Z(n5032) );
  XOR U6903 ( .A(n4937), .B(n4936), .Z(n5028) );
  AND U6904 ( .A(a[15]), .B(b[51]), .Z(n5018) );
  XNOR U6905 ( .A(n4939), .B(n4938), .Z(n5017) );
  NANDN U6906 ( .A(n5018), .B(n5017), .Z(n5020) );
  NAND U6907 ( .A(a[14]), .B(b[51]), .Z(n4942) );
  XNOR U6908 ( .A(n4941), .B(n4940), .Z(n4943) );
  NANDN U6909 ( .A(n4942), .B(n4943), .Z(n5016) );
  XOR U6910 ( .A(n4943), .B(n4942), .Z(n5304) );
  XOR U6911 ( .A(n4945), .B(n4944), .Z(n4999) );
  XOR U6912 ( .A(n4947), .B(n4946), .Z(n4989) );
  NAND U6913 ( .A(a[7]), .B(b[51]), .Z(n4979) );
  XOR U6914 ( .A(n4949), .B(n4948), .Z(n4980) );
  NANDN U6915 ( .A(n4979), .B(n4980), .Z(n4982) );
  NAND U6916 ( .A(a[0]), .B(b[51]), .Z(n5531) );
  AND U6917 ( .A(a[1]), .B(b[52]), .Z(n4952) );
  NANDN U6918 ( .A(n5531), .B(n4952), .Z(n5237) );
  NANDN U6919 ( .A(n5237), .B(n4950), .Z(n4954) );
  AND U6920 ( .A(a[2]), .B(b[51]), .Z(n5243) );
  NANDN U6921 ( .A(n5242), .B(n5243), .Z(n4953) );
  AND U6922 ( .A(n4954), .B(n4953), .Z(n4957) );
  AND U6923 ( .A(a[3]), .B(b[51]), .Z(n4958) );
  NANDN U6924 ( .A(n4957), .B(n4958), .Z(n4960) );
  XOR U6925 ( .A(n4956), .B(n4955), .Z(n5248) );
  NANDN U6926 ( .A(n5248), .B(n5249), .Z(n4959) );
  AND U6927 ( .A(n4960), .B(n4959), .Z(n4963) );
  NANDN U6928 ( .A(n4963), .B(n4964), .Z(n4966) );
  AND U6929 ( .A(a[4]), .B(b[51]), .Z(n5257) );
  NAND U6930 ( .A(n5257), .B(n5256), .Z(n4965) );
  AND U6931 ( .A(n4966), .B(n4965), .Z(n4967) );
  AND U6932 ( .A(a[5]), .B(b[51]), .Z(n4968) );
  NANDN U6933 ( .A(n4967), .B(n4968), .Z(n4972) );
  NAND U6934 ( .A(n5261), .B(n5260), .Z(n4971) );
  AND U6935 ( .A(n4972), .B(n4971), .Z(n4975) );
  XOR U6936 ( .A(n4974), .B(n4973), .Z(n4976) );
  NANDN U6937 ( .A(n4975), .B(n4976), .Z(n4978) );
  AND U6938 ( .A(a[6]), .B(b[51]), .Z(n5236) );
  NAND U6939 ( .A(n5236), .B(n5235), .Z(n4977) );
  AND U6940 ( .A(n4978), .B(n4977), .Z(n5272) );
  NANDN U6941 ( .A(n5272), .B(n5273), .Z(n4981) );
  AND U6942 ( .A(n4982), .B(n4981), .Z(n4983) );
  AND U6943 ( .A(a[8]), .B(b[51]), .Z(n4984) );
  NANDN U6944 ( .A(n4983), .B(n4984), .Z(n4988) );
  NAND U6945 ( .A(n5234), .B(n5233), .Z(n4987) );
  AND U6946 ( .A(n4988), .B(n4987), .Z(n4990) );
  NANDN U6947 ( .A(n4989), .B(n4990), .Z(n4992) );
  AND U6948 ( .A(a[9]), .B(b[51]), .Z(n5280) );
  NANDN U6949 ( .A(n5280), .B(n5281), .Z(n4991) );
  AND U6950 ( .A(n4992), .B(n4991), .Z(n4995) );
  NAND U6951 ( .A(n4995), .B(n4996), .Z(n4998) );
  XOR U6952 ( .A(n4996), .B(n4995), .Z(n5232) );
  AND U6953 ( .A(a[10]), .B(b[51]), .Z(n5231) );
  NAND U6954 ( .A(n5232), .B(n5231), .Z(n4997) );
  AND U6955 ( .A(n4998), .B(n4997), .Z(n5000) );
  NANDN U6956 ( .A(n4999), .B(n5000), .Z(n5002) );
  NAND U6957 ( .A(a[11]), .B(b[51]), .Z(n5229) );
  NAND U6958 ( .A(n5230), .B(n5229), .Z(n5001) );
  AND U6959 ( .A(n5002), .B(n5001), .Z(n5005) );
  NANDN U6960 ( .A(n5005), .B(n5006), .Z(n5008) );
  AND U6961 ( .A(a[12]), .B(b[51]), .Z(n5227) );
  NANDN U6962 ( .A(n5227), .B(n5228), .Z(n5007) );
  AND U6963 ( .A(n5008), .B(n5007), .Z(n5011) );
  NANDN U6964 ( .A(n5011), .B(n5012), .Z(n5014) );
  AND U6965 ( .A(a[13]), .B(b[51]), .Z(n5300) );
  NANDN U6966 ( .A(n5300), .B(n5301), .Z(n5013) );
  AND U6967 ( .A(n5014), .B(n5013), .Z(n5305) );
  NANDN U6968 ( .A(n5304), .B(n5305), .Z(n5015) );
  NAND U6969 ( .A(n5016), .B(n5015), .Z(n5225) );
  XNOR U6970 ( .A(n5018), .B(n5017), .Z(n5226) );
  NANDN U6971 ( .A(n5225), .B(n5226), .Z(n5019) );
  AND U6972 ( .A(n5020), .B(n5019), .Z(n5024) );
  XNOR U6973 ( .A(n5022), .B(n5021), .Z(n5023) );
  NANDN U6974 ( .A(n5024), .B(n5023), .Z(n5026) );
  AND U6975 ( .A(a[16]), .B(b[51]), .Z(n5315) );
  XNOR U6976 ( .A(n5024), .B(n5023), .Z(n5314) );
  NANDN U6977 ( .A(n5315), .B(n5314), .Z(n5025) );
  AND U6978 ( .A(n5026), .B(n5025), .Z(n5027) );
  NANDN U6979 ( .A(n5028), .B(n5027), .Z(n5030) );
  XNOR U6980 ( .A(n5028), .B(n5027), .Z(n5224) );
  AND U6981 ( .A(a[17]), .B(b[51]), .Z(n5223) );
  NAND U6982 ( .A(n5224), .B(n5223), .Z(n5029) );
  AND U6983 ( .A(n5030), .B(n5029), .Z(n5031) );
  NANDN U6984 ( .A(n5032), .B(n5031), .Z(n5034) );
  XOR U6985 ( .A(n5032), .B(n5031), .Z(n5221) );
  AND U6986 ( .A(a[18]), .B(b[51]), .Z(n5222) );
  OR U6987 ( .A(n5221), .B(n5222), .Z(n5033) );
  NAND U6988 ( .A(n5034), .B(n5033), .Z(n5037) );
  XNOR U6989 ( .A(n5036), .B(n5035), .Z(n5038) );
  NANDN U6990 ( .A(n5037), .B(n5038), .Z(n5040) );
  XNOR U6991 ( .A(n5038), .B(n5037), .Z(n5220) );
  AND U6992 ( .A(a[19]), .B(b[51]), .Z(n5219) );
  NAND U6993 ( .A(n5220), .B(n5219), .Z(n5039) );
  AND U6994 ( .A(n5040), .B(n5039), .Z(n5333) );
  OR U6995 ( .A(n5332), .B(n5333), .Z(n5041) );
  AND U6996 ( .A(n5042), .B(n5041), .Z(n5046) );
  XNOR U6997 ( .A(n5044), .B(n5043), .Z(n5045) );
  NANDN U6998 ( .A(n5046), .B(n5045), .Z(n5048) );
  NAND U6999 ( .A(a[21]), .B(b[51]), .Z(n5338) );
  XNOR U7000 ( .A(n5046), .B(n5045), .Z(n5339) );
  NANDN U7001 ( .A(n5338), .B(n5339), .Z(n5047) );
  AND U7002 ( .A(n5048), .B(n5047), .Z(n5050) );
  NANDN U7003 ( .A(n5049), .B(n5050), .Z(n5052) );
  XOR U7004 ( .A(n5050), .B(n5049), .Z(n5217) );
  AND U7005 ( .A(a[22]), .B(b[51]), .Z(n5218) );
  OR U7006 ( .A(n5217), .B(n5218), .Z(n5051) );
  NAND U7007 ( .A(n5052), .B(n5051), .Z(n5055) );
  XNOR U7008 ( .A(n5054), .B(n5053), .Z(n5056) );
  NANDN U7009 ( .A(n5055), .B(n5056), .Z(n5058) );
  NAND U7010 ( .A(a[23]), .B(b[51]), .Z(n5213) );
  XNOR U7011 ( .A(n5056), .B(n5055), .Z(n5214) );
  NANDN U7012 ( .A(n5213), .B(n5214), .Z(n5057) );
  AND U7013 ( .A(n5058), .B(n5057), .Z(n5062) );
  AND U7014 ( .A(a[24]), .B(b[51]), .Z(n5061) );
  NANDN U7015 ( .A(n5062), .B(n5061), .Z(n5064) );
  XOR U7016 ( .A(n5060), .B(n5059), .Z(n5350) );
  XNOR U7017 ( .A(n5062), .B(n5061), .Z(n5351) );
  NANDN U7018 ( .A(n5350), .B(n5351), .Z(n5063) );
  AND U7019 ( .A(n5064), .B(n5063), .Z(n5068) );
  XNOR U7020 ( .A(n5066), .B(n5065), .Z(n5067) );
  NANDN U7021 ( .A(n5068), .B(n5067), .Z(n5070) );
  NAND U7022 ( .A(a[25]), .B(b[51]), .Z(n5356) );
  XNOR U7023 ( .A(n5068), .B(n5067), .Z(n5357) );
  NANDN U7024 ( .A(n5356), .B(n5357), .Z(n5069) );
  AND U7025 ( .A(n5070), .B(n5069), .Z(n5074) );
  XNOR U7026 ( .A(n5072), .B(n5071), .Z(n5073) );
  NANDN U7027 ( .A(n5074), .B(n5073), .Z(n5076) );
  NAND U7028 ( .A(a[26]), .B(b[51]), .Z(n5362) );
  XNOR U7029 ( .A(n5074), .B(n5073), .Z(n5363) );
  NANDN U7030 ( .A(n5362), .B(n5363), .Z(n5075) );
  AND U7031 ( .A(n5076), .B(n5075), .Z(n5077) );
  NANDN U7032 ( .A(n5078), .B(n5077), .Z(n5080) );
  XOR U7033 ( .A(n5078), .B(n5077), .Z(n5209) );
  AND U7034 ( .A(a[27]), .B(b[51]), .Z(n5210) );
  OR U7035 ( .A(n5209), .B(n5210), .Z(n5079) );
  AND U7036 ( .A(n5080), .B(n5079), .Z(n5082) );
  NANDN U7037 ( .A(n5081), .B(n5082), .Z(n5084) );
  NAND U7038 ( .A(a[28]), .B(b[51]), .Z(n5372) );
  XNOR U7039 ( .A(n5082), .B(n5081), .Z(n5373) );
  NANDN U7040 ( .A(n5372), .B(n5373), .Z(n5083) );
  AND U7041 ( .A(n5084), .B(n5083), .Z(n5088) );
  XNOR U7042 ( .A(n5086), .B(n5085), .Z(n5087) );
  NANDN U7043 ( .A(n5088), .B(n5087), .Z(n5090) );
  XNOR U7044 ( .A(n5088), .B(n5087), .Z(n5208) );
  AND U7045 ( .A(a[29]), .B(b[51]), .Z(n5207) );
  NAND U7046 ( .A(n5208), .B(n5207), .Z(n5089) );
  AND U7047 ( .A(n5090), .B(n5089), .Z(n5091) );
  NANDN U7048 ( .A(n5092), .B(n5091), .Z(n5094) );
  XOR U7049 ( .A(n5092), .B(n5091), .Z(n5205) );
  AND U7050 ( .A(a[30]), .B(b[51]), .Z(n5206) );
  OR U7051 ( .A(n5205), .B(n5206), .Z(n5093) );
  NAND U7052 ( .A(n5094), .B(n5093), .Z(n5097) );
  XNOR U7053 ( .A(n5096), .B(n5095), .Z(n5098) );
  NANDN U7054 ( .A(n5097), .B(n5098), .Z(n5100) );
  NAND U7055 ( .A(a[31]), .B(b[51]), .Z(n5384) );
  XNOR U7056 ( .A(n5098), .B(n5097), .Z(n5385) );
  NANDN U7057 ( .A(n5384), .B(n5385), .Z(n5099) );
  AND U7058 ( .A(n5100), .B(n5099), .Z(n5204) );
  XNOR U7059 ( .A(n5102), .B(n5101), .Z(n5203) );
  NANDN U7060 ( .A(n5204), .B(n5203), .Z(n5103) );
  AND U7061 ( .A(n5104), .B(n5103), .Z(n5105) );
  NANDN U7062 ( .A(n5106), .B(n5105), .Z(n5108) );
  AND U7063 ( .A(a[33]), .B(b[51]), .Z(n5202) );
  XNOR U7064 ( .A(n5106), .B(n5105), .Z(n5201) );
  NANDN U7065 ( .A(n5202), .B(n5201), .Z(n5107) );
  AND U7066 ( .A(n5108), .B(n5107), .Z(n5110) );
  XOR U7067 ( .A(n5110), .B(n5109), .Z(n5200) );
  AND U7068 ( .A(a[34]), .B(b[51]), .Z(n5199) );
  AND U7069 ( .A(a[35]), .B(b[51]), .Z(n5111) );
  NANDN U7070 ( .A(n5112), .B(n5111), .Z(n5116) );
  XNOR U7071 ( .A(n5112), .B(n5111), .Z(n5196) );
  XNOR U7072 ( .A(n5114), .B(n5113), .Z(n5195) );
  NAND U7073 ( .A(n5196), .B(n5195), .Z(n5115) );
  AND U7074 ( .A(n5116), .B(n5115), .Z(n5194) );
  XOR U7075 ( .A(n5118), .B(n5117), .Z(n5193) );
  NANDN U7076 ( .A(n5194), .B(n5193), .Z(n5119) );
  AND U7077 ( .A(n5120), .B(n5119), .Z(n5124) );
  AND U7078 ( .A(a[37]), .B(b[51]), .Z(n5123) );
  NANDN U7079 ( .A(n5124), .B(n5123), .Z(n5126) );
  XOR U7080 ( .A(n5122), .B(n5121), .Z(n5409) );
  XNOR U7081 ( .A(n5124), .B(n5123), .Z(n5408) );
  NANDN U7082 ( .A(n5409), .B(n5408), .Z(n5125) );
  AND U7083 ( .A(n5126), .B(n5125), .Z(n5128) );
  AND U7084 ( .A(a[38]), .B(b[51]), .Z(n5127) );
  NANDN U7085 ( .A(n5128), .B(n5127), .Z(n5132) );
  XNOR U7086 ( .A(n5128), .B(n5127), .Z(n5415) );
  XOR U7087 ( .A(n5130), .B(n5129), .Z(n5414) );
  NAND U7088 ( .A(n5415), .B(n5414), .Z(n5131) );
  AND U7089 ( .A(n5132), .B(n5131), .Z(n5134) );
  AND U7090 ( .A(a[39]), .B(b[51]), .Z(n5133) );
  NANDN U7091 ( .A(n5134), .B(n5133), .Z(n5138) );
  XNOR U7092 ( .A(n5134), .B(n5133), .Z(n5420) );
  XOR U7093 ( .A(n5136), .B(n5135), .Z(n5421) );
  NAND U7094 ( .A(n5420), .B(n5421), .Z(n5137) );
  AND U7095 ( .A(n5138), .B(n5137), .Z(n5139) );
  AND U7096 ( .A(a[40]), .B(b[51]), .Z(n5140) );
  NANDN U7097 ( .A(n5139), .B(n5140), .Z(n5144) );
  XNOR U7098 ( .A(n5142), .B(n5141), .Z(n5429) );
  NAND U7099 ( .A(n5428), .B(n5429), .Z(n5143) );
  AND U7100 ( .A(n5144), .B(n5143), .Z(n5145) );
  AND U7101 ( .A(a[41]), .B(b[51]), .Z(n5146) );
  NANDN U7102 ( .A(n5145), .B(n5146), .Z(n5150) );
  XOR U7103 ( .A(n5148), .B(n5147), .Z(n5432) );
  NAND U7104 ( .A(n5433), .B(n5432), .Z(n5149) );
  AND U7105 ( .A(n5150), .B(n5149), .Z(n5152) );
  NANDN U7106 ( .A(n5151), .B(n5152), .Z(n5156) );
  NAND U7107 ( .A(n5439), .B(n5438), .Z(n5155) );
  NAND U7108 ( .A(n5156), .B(n5155), .Z(n5157) );
  AND U7109 ( .A(a[43]), .B(b[51]), .Z(n5158) );
  NANDN U7110 ( .A(n5157), .B(n5158), .Z(n5162) );
  XNOR U7111 ( .A(n5160), .B(n5159), .Z(n5447) );
  NAND U7112 ( .A(n5446), .B(n5447), .Z(n5161) );
  AND U7113 ( .A(n5162), .B(n5161), .Z(n5163) );
  AND U7114 ( .A(a[44]), .B(b[51]), .Z(n5164) );
  NANDN U7115 ( .A(n5163), .B(n5164), .Z(n5168) );
  XNOR U7116 ( .A(n5166), .B(n5165), .Z(n5453) );
  NAND U7117 ( .A(n5452), .B(n5453), .Z(n5167) );
  AND U7118 ( .A(n5168), .B(n5167), .Z(n5169) );
  AND U7119 ( .A(a[45]), .B(b[51]), .Z(n5170) );
  NANDN U7120 ( .A(n5169), .B(n5170), .Z(n5174) );
  NAND U7121 ( .A(n5456), .B(n5457), .Z(n5173) );
  AND U7122 ( .A(n5174), .B(n5173), .Z(n5175) );
  AND U7123 ( .A(a[46]), .B(b[51]), .Z(n5176) );
  NANDN U7124 ( .A(n5175), .B(n5176), .Z(n5180) );
  XNOR U7125 ( .A(n5178), .B(n5177), .Z(n5465) );
  NAND U7126 ( .A(n5464), .B(n5465), .Z(n5179) );
  AND U7127 ( .A(n5180), .B(n5179), .Z(n5181) );
  AND U7128 ( .A(a[47]), .B(b[51]), .Z(n5182) );
  NANDN U7129 ( .A(n5181), .B(n5182), .Z(n5186) );
  XOR U7130 ( .A(n5184), .B(n5183), .Z(n5468) );
  NAND U7131 ( .A(n5469), .B(n5468), .Z(n5185) );
  AND U7132 ( .A(n5186), .B(n5185), .Z(n5188) );
  NANDN U7133 ( .A(n5187), .B(n5188), .Z(n5192) );
  NAND U7134 ( .A(n5475), .B(n5474), .Z(n5191) );
  NAND U7135 ( .A(n5192), .B(n5191), .Z(n10191) );
  XNOR U7136 ( .A(n10192), .B(n10193), .Z(n10120) );
  AND U7137 ( .A(a[50]), .B(b[50]), .Z(n10119) );
  AND U7138 ( .A(a[48]), .B(b[50]), .Z(n5470) );
  AND U7139 ( .A(a[47]), .B(b[50]), .Z(n5462) );
  AND U7140 ( .A(a[45]), .B(b[50]), .Z(n5450) );
  AND U7141 ( .A(a[44]), .B(b[50]), .Z(n5444) );
  NAND U7142 ( .A(a[43]), .B(b[50]), .Z(n5440) );
  AND U7143 ( .A(a[42]), .B(b[50]), .Z(n5434) );
  AND U7144 ( .A(a[41]), .B(b[50]), .Z(n5426) );
  NAND U7145 ( .A(a[40]), .B(b[50]), .Z(n5422) );
  AND U7146 ( .A(a[39]), .B(b[50]), .Z(n5417) );
  NAND U7147 ( .A(a[37]), .B(b[50]), .Z(n5404) );
  XNOR U7148 ( .A(n5194), .B(n5193), .Z(n5405) );
  NANDN U7149 ( .A(n5404), .B(n5405), .Z(n5407) );
  NAND U7150 ( .A(a[36]), .B(b[50]), .Z(n5197) );
  XOR U7151 ( .A(n5196), .B(n5195), .Z(n5198) );
  NANDN U7152 ( .A(n5197), .B(n5198), .Z(n5403) );
  XNOR U7153 ( .A(n5198), .B(n5197), .Z(n5485) );
  XOR U7154 ( .A(n5200), .B(n5199), .Z(n5399) );
  XOR U7155 ( .A(n5202), .B(n5201), .Z(n5394) );
  XOR U7156 ( .A(n5204), .B(n5203), .Z(n5390) );
  AND U7157 ( .A(a[33]), .B(b[50]), .Z(n5391) );
  NANDN U7158 ( .A(n5390), .B(n5391), .Z(n5393) );
  XOR U7159 ( .A(n5206), .B(n5205), .Z(n5381) );
  XOR U7160 ( .A(n5208), .B(n5207), .Z(n5377) );
  XOR U7161 ( .A(n5210), .B(n5209), .Z(n5212) );
  AND U7162 ( .A(a[28]), .B(b[50]), .Z(n5211) );
  NANDN U7163 ( .A(n5212), .B(n5211), .Z(n5369) );
  XOR U7164 ( .A(n5212), .B(n5211), .Z(n5498) );
  NAND U7165 ( .A(a[24]), .B(b[50]), .Z(n5215) );
  XNOR U7166 ( .A(n5214), .B(n5213), .Z(n5216) );
  NANDN U7167 ( .A(n5215), .B(n5216), .Z(n5349) );
  XOR U7168 ( .A(n5216), .B(n5215), .Z(n5504) );
  XOR U7169 ( .A(n5218), .B(n5217), .Z(n5345) );
  AND U7170 ( .A(a[23]), .B(b[50]), .Z(n5344) );
  NANDN U7171 ( .A(n5345), .B(n5344), .Z(n5347) );
  XOR U7172 ( .A(n5220), .B(n5219), .Z(n5329) );
  XOR U7173 ( .A(n5222), .B(n5221), .Z(n5325) );
  AND U7174 ( .A(a[19]), .B(b[50]), .Z(n5324) );
  NANDN U7175 ( .A(n5325), .B(n5324), .Z(n5327) );
  XOR U7176 ( .A(n5224), .B(n5223), .Z(n5321) );
  XOR U7177 ( .A(n5226), .B(n5225), .Z(n5310) );
  AND U7178 ( .A(a[13]), .B(b[50]), .Z(n5294) );
  NAND U7179 ( .A(n5294), .B(n5295), .Z(n5297) );
  XOR U7180 ( .A(n5230), .B(n5229), .Z(n5290) );
  XOR U7181 ( .A(n5232), .B(n5231), .Z(n5286) );
  XOR U7182 ( .A(n5234), .B(n5233), .Z(n5276) );
  NAND U7183 ( .A(a[7]), .B(b[50]), .Z(n5266) );
  XOR U7184 ( .A(n5236), .B(n5235), .Z(n5267) );
  NANDN U7185 ( .A(n5266), .B(n5267), .Z(n5269) );
  NAND U7186 ( .A(a[0]), .B(b[50]), .Z(n5828) );
  AND U7187 ( .A(a[1]), .B(b[51]), .Z(n5239) );
  NANDN U7188 ( .A(n5828), .B(n5239), .Z(n5530) );
  NANDN U7189 ( .A(n5530), .B(n5237), .Z(n5241) );
  AND U7190 ( .A(a[2]), .B(b[50]), .Z(n5536) );
  NANDN U7191 ( .A(n5535), .B(n5536), .Z(n5240) );
  AND U7192 ( .A(n5241), .B(n5240), .Z(n5244) );
  AND U7193 ( .A(a[3]), .B(b[50]), .Z(n5245) );
  NANDN U7194 ( .A(n5244), .B(n5245), .Z(n5247) );
  XOR U7195 ( .A(n5243), .B(n5242), .Z(n5541) );
  NANDN U7196 ( .A(n5541), .B(n5542), .Z(n5246) );
  AND U7197 ( .A(n5247), .B(n5246), .Z(n5250) );
  NANDN U7198 ( .A(n5250), .B(n5251), .Z(n5253) );
  AND U7199 ( .A(a[4]), .B(b[50]), .Z(n5550) );
  NAND U7200 ( .A(n5550), .B(n5549), .Z(n5252) );
  AND U7201 ( .A(n5253), .B(n5252), .Z(n5254) );
  AND U7202 ( .A(a[5]), .B(b[50]), .Z(n5255) );
  NANDN U7203 ( .A(n5254), .B(n5255), .Z(n5259) );
  XOR U7204 ( .A(n5257), .B(n5256), .Z(n5553) );
  NAND U7205 ( .A(n5554), .B(n5553), .Z(n5258) );
  AND U7206 ( .A(n5259), .B(n5258), .Z(n5262) );
  XOR U7207 ( .A(n5261), .B(n5260), .Z(n5263) );
  NANDN U7208 ( .A(n5262), .B(n5263), .Z(n5265) );
  AND U7209 ( .A(a[6]), .B(b[50]), .Z(n5529) );
  NAND U7210 ( .A(n5529), .B(n5528), .Z(n5264) );
  AND U7211 ( .A(n5265), .B(n5264), .Z(n5565) );
  NANDN U7212 ( .A(n5565), .B(n5566), .Z(n5268) );
  AND U7213 ( .A(n5269), .B(n5268), .Z(n5270) );
  AND U7214 ( .A(a[8]), .B(b[50]), .Z(n5271) );
  NANDN U7215 ( .A(n5270), .B(n5271), .Z(n5275) );
  NAND U7216 ( .A(n5527), .B(n5526), .Z(n5274) );
  AND U7217 ( .A(n5275), .B(n5274), .Z(n5277) );
  NANDN U7218 ( .A(n5276), .B(n5277), .Z(n5279) );
  AND U7219 ( .A(a[9]), .B(b[50]), .Z(n5573) );
  NANDN U7220 ( .A(n5573), .B(n5574), .Z(n5278) );
  AND U7221 ( .A(n5279), .B(n5278), .Z(n5282) );
  NAND U7222 ( .A(n5282), .B(n5283), .Z(n5285) );
  AND U7223 ( .A(a[10]), .B(b[50]), .Z(n5582) );
  XOR U7224 ( .A(n5283), .B(n5282), .Z(n5581) );
  NAND U7225 ( .A(n5582), .B(n5581), .Z(n5284) );
  AND U7226 ( .A(n5285), .B(n5284), .Z(n5287) );
  NANDN U7227 ( .A(n5286), .B(n5287), .Z(n5289) );
  AND U7228 ( .A(a[11]), .B(b[50]), .Z(n5585) );
  NANDN U7229 ( .A(n5585), .B(n5586), .Z(n5288) );
  AND U7230 ( .A(n5289), .B(n5288), .Z(n5291) );
  NANDN U7231 ( .A(n5290), .B(n5291), .Z(n5293) );
  AND U7232 ( .A(a[12]), .B(b[50]), .Z(n5592) );
  NAND U7233 ( .A(n5592), .B(n5591), .Z(n5292) );
  AND U7234 ( .A(n5293), .B(n5292), .Z(n5599) );
  XOR U7235 ( .A(n5295), .B(n5294), .Z(n5600) );
  NANDN U7236 ( .A(n5599), .B(n5600), .Z(n5296) );
  AND U7237 ( .A(n5297), .B(n5296), .Z(n5298) );
  AND U7238 ( .A(a[14]), .B(b[50]), .Z(n5299) );
  NANDN U7239 ( .A(n5298), .B(n5299), .Z(n5303) );
  NAND U7240 ( .A(n5605), .B(n5606), .Z(n5302) );
  AND U7241 ( .A(n5303), .B(n5302), .Z(n5307) );
  XNOR U7242 ( .A(n5305), .B(n5304), .Z(n5306) );
  NANDN U7243 ( .A(n5307), .B(n5306), .Z(n5309) );
  XNOR U7244 ( .A(n5307), .B(n5306), .Z(n5525) );
  AND U7245 ( .A(a[15]), .B(b[50]), .Z(n5524) );
  NAND U7246 ( .A(n5525), .B(n5524), .Z(n5308) );
  AND U7247 ( .A(n5309), .B(n5308), .Z(n5311) );
  NANDN U7248 ( .A(n5310), .B(n5311), .Z(n5313) );
  XOR U7249 ( .A(n5311), .B(n5310), .Z(n5520) );
  AND U7250 ( .A(a[16]), .B(b[50]), .Z(n5521) );
  OR U7251 ( .A(n5520), .B(n5521), .Z(n5312) );
  AND U7252 ( .A(n5313), .B(n5312), .Z(n5317) );
  XNOR U7253 ( .A(n5315), .B(n5314), .Z(n5316) );
  NANDN U7254 ( .A(n5317), .B(n5316), .Z(n5319) );
  AND U7255 ( .A(a[17]), .B(b[50]), .Z(n5517) );
  XNOR U7256 ( .A(n5317), .B(n5316), .Z(n5516) );
  NANDN U7257 ( .A(n5517), .B(n5516), .Z(n5318) );
  NAND U7258 ( .A(n5319), .B(n5318), .Z(n5320) );
  NANDN U7259 ( .A(n5321), .B(n5320), .Z(n5323) );
  XOR U7260 ( .A(n5321), .B(n5320), .Z(n5514) );
  AND U7261 ( .A(a[18]), .B(b[50]), .Z(n5515) );
  OR U7262 ( .A(n5514), .B(n5515), .Z(n5322) );
  NAND U7263 ( .A(n5323), .B(n5322), .Z(n5512) );
  XNOR U7264 ( .A(n5325), .B(n5324), .Z(n5513) );
  NANDN U7265 ( .A(n5512), .B(n5513), .Z(n5326) );
  AND U7266 ( .A(n5327), .B(n5326), .Z(n5328) );
  NANDN U7267 ( .A(n5329), .B(n5328), .Z(n5331) );
  XOR U7268 ( .A(n5329), .B(n5328), .Z(n5510) );
  AND U7269 ( .A(a[20]), .B(b[50]), .Z(n5511) );
  OR U7270 ( .A(n5510), .B(n5511), .Z(n5330) );
  AND U7271 ( .A(n5331), .B(n5330), .Z(n5335) );
  XNOR U7272 ( .A(n5333), .B(n5332), .Z(n5334) );
  NANDN U7273 ( .A(n5335), .B(n5334), .Z(n5337) );
  XOR U7274 ( .A(n5335), .B(n5334), .Z(n5508) );
  AND U7275 ( .A(a[21]), .B(b[50]), .Z(n5509) );
  OR U7276 ( .A(n5508), .B(n5509), .Z(n5336) );
  NAND U7277 ( .A(n5337), .B(n5336), .Z(n5340) );
  XNOR U7278 ( .A(n5339), .B(n5338), .Z(n5341) );
  NANDN U7279 ( .A(n5340), .B(n5341), .Z(n5343) );
  NAND U7280 ( .A(a[22]), .B(b[50]), .Z(n5506) );
  XNOR U7281 ( .A(n5341), .B(n5340), .Z(n5507) );
  NANDN U7282 ( .A(n5506), .B(n5507), .Z(n5342) );
  AND U7283 ( .A(n5343), .B(n5342), .Z(n5638) );
  XNOR U7284 ( .A(n5345), .B(n5344), .Z(n5637) );
  NANDN U7285 ( .A(n5638), .B(n5637), .Z(n5346) );
  AND U7286 ( .A(n5347), .B(n5346), .Z(n5505) );
  OR U7287 ( .A(n5504), .B(n5505), .Z(n5348) );
  AND U7288 ( .A(n5349), .B(n5348), .Z(n5353) );
  AND U7289 ( .A(a[25]), .B(b[50]), .Z(n5352) );
  NANDN U7290 ( .A(n5353), .B(n5352), .Z(n5355) );
  XOR U7291 ( .A(n5351), .B(n5350), .Z(n5647) );
  XNOR U7292 ( .A(n5353), .B(n5352), .Z(n5648) );
  NANDN U7293 ( .A(n5647), .B(n5648), .Z(n5354) );
  AND U7294 ( .A(n5355), .B(n5354), .Z(n5359) );
  AND U7295 ( .A(a[26]), .B(b[50]), .Z(n5358) );
  NANDN U7296 ( .A(n5359), .B(n5358), .Z(n5361) );
  XOR U7297 ( .A(n5357), .B(n5356), .Z(n5502) );
  XNOR U7298 ( .A(n5359), .B(n5358), .Z(n5503) );
  NANDN U7299 ( .A(n5502), .B(n5503), .Z(n5360) );
  AND U7300 ( .A(n5361), .B(n5360), .Z(n5365) );
  XNOR U7301 ( .A(n5363), .B(n5362), .Z(n5364) );
  NANDN U7302 ( .A(n5365), .B(n5364), .Z(n5367) );
  NAND U7303 ( .A(a[27]), .B(b[50]), .Z(n5500) );
  XNOR U7304 ( .A(n5365), .B(n5364), .Z(n5501) );
  NANDN U7305 ( .A(n5500), .B(n5501), .Z(n5366) );
  AND U7306 ( .A(n5367), .B(n5366), .Z(n5499) );
  OR U7307 ( .A(n5498), .B(n5499), .Z(n5368) );
  AND U7308 ( .A(n5369), .B(n5368), .Z(n5371) );
  AND U7309 ( .A(a[29]), .B(b[50]), .Z(n5370) );
  NANDN U7310 ( .A(n5371), .B(n5370), .Z(n5375) );
  XNOR U7311 ( .A(n5371), .B(n5370), .Z(n5497) );
  XNOR U7312 ( .A(n5373), .B(n5372), .Z(n5496) );
  NAND U7313 ( .A(n5497), .B(n5496), .Z(n5374) );
  AND U7314 ( .A(n5375), .B(n5374), .Z(n5376) );
  NANDN U7315 ( .A(n5377), .B(n5376), .Z(n5379) );
  XOR U7316 ( .A(n5377), .B(n5376), .Z(n5494) );
  AND U7317 ( .A(a[30]), .B(b[50]), .Z(n5495) );
  OR U7318 ( .A(n5494), .B(n5495), .Z(n5378) );
  AND U7319 ( .A(n5379), .B(n5378), .Z(n5380) );
  NANDN U7320 ( .A(n5381), .B(n5380), .Z(n5383) );
  XNOR U7321 ( .A(n5381), .B(n5380), .Z(n5493) );
  AND U7322 ( .A(a[31]), .B(b[50]), .Z(n5492) );
  NAND U7323 ( .A(n5493), .B(n5492), .Z(n5382) );
  AND U7324 ( .A(n5383), .B(n5382), .Z(n5387) );
  XNOR U7325 ( .A(n5385), .B(n5384), .Z(n5386) );
  NANDN U7326 ( .A(n5387), .B(n5386), .Z(n5389) );
  NAND U7327 ( .A(a[32]), .B(b[50]), .Z(n5490) );
  XNOR U7328 ( .A(n5387), .B(n5386), .Z(n5491) );
  NANDN U7329 ( .A(n5490), .B(n5491), .Z(n5388) );
  AND U7330 ( .A(n5389), .B(n5388), .Z(n5489) );
  XNOR U7331 ( .A(n5391), .B(n5390), .Z(n5488) );
  NANDN U7332 ( .A(n5489), .B(n5488), .Z(n5392) );
  AND U7333 ( .A(n5393), .B(n5392), .Z(n5395) );
  NANDN U7334 ( .A(n5394), .B(n5395), .Z(n5397) );
  AND U7335 ( .A(a[34]), .B(b[50]), .Z(n5688) );
  XNOR U7336 ( .A(n5395), .B(n5394), .Z(n5687) );
  NANDN U7337 ( .A(n5688), .B(n5687), .Z(n5396) );
  NAND U7338 ( .A(n5397), .B(n5396), .Z(n5398) );
  NANDN U7339 ( .A(n5399), .B(n5398), .Z(n5401) );
  XOR U7340 ( .A(n5399), .B(n5398), .Z(n5486) );
  AND U7341 ( .A(a[35]), .B(b[50]), .Z(n5487) );
  OR U7342 ( .A(n5486), .B(n5487), .Z(n5400) );
  AND U7343 ( .A(n5401), .B(n5400), .Z(n5484) );
  NAND U7344 ( .A(n5485), .B(n5484), .Z(n5402) );
  AND U7345 ( .A(n5403), .B(n5402), .Z(n5700) );
  XNOR U7346 ( .A(n5405), .B(n5404), .Z(n5699) );
  NANDN U7347 ( .A(n5700), .B(n5699), .Z(n5406) );
  AND U7348 ( .A(n5407), .B(n5406), .Z(n5410) );
  XOR U7349 ( .A(n5409), .B(n5408), .Z(n5411) );
  NAND U7350 ( .A(n5410), .B(n5411), .Z(n5413) );
  AND U7351 ( .A(a[38]), .B(b[50]), .Z(n5483) );
  XOR U7352 ( .A(n5411), .B(n5410), .Z(n5482) );
  NANDN U7353 ( .A(n5483), .B(n5482), .Z(n5412) );
  NAND U7354 ( .A(n5413), .B(n5412), .Z(n5416) );
  NANDN U7355 ( .A(n5417), .B(n5416), .Z(n5419) );
  XOR U7356 ( .A(n5415), .B(n5414), .Z(n5481) );
  XNOR U7357 ( .A(n5417), .B(n5416), .Z(n5480) );
  NANDN U7358 ( .A(n5481), .B(n5480), .Z(n5418) );
  AND U7359 ( .A(n5419), .B(n5418), .Z(n5423) );
  NANDN U7360 ( .A(n5422), .B(n5423), .Z(n5425) );
  XOR U7361 ( .A(n5421), .B(n5420), .Z(n5716) );
  XNOR U7362 ( .A(n5423), .B(n5422), .Z(n5715) );
  NAND U7363 ( .A(n5716), .B(n5715), .Z(n5424) );
  AND U7364 ( .A(n5425), .B(n5424), .Z(n5427) );
  NANDN U7365 ( .A(n5426), .B(n5427), .Z(n5431) );
  XNOR U7366 ( .A(n5429), .B(n5428), .Z(n5722) );
  NAND U7367 ( .A(n5721), .B(n5722), .Z(n5430) );
  NAND U7368 ( .A(n5431), .B(n5430), .Z(n5435) );
  NANDN U7369 ( .A(n5434), .B(n5435), .Z(n5437) );
  XOR U7370 ( .A(n5433), .B(n5432), .Z(n5727) );
  NANDN U7371 ( .A(n5727), .B(n5728), .Z(n5436) );
  AND U7372 ( .A(n5437), .B(n5436), .Z(n5441) );
  NANDN U7373 ( .A(n5440), .B(n5441), .Z(n5443) );
  XOR U7374 ( .A(n5439), .B(n5438), .Z(n5733) );
  NANDN U7375 ( .A(n5733), .B(n5734), .Z(n5442) );
  AND U7376 ( .A(n5443), .B(n5442), .Z(n5445) );
  NANDN U7377 ( .A(n5444), .B(n5445), .Z(n5449) );
  XNOR U7378 ( .A(n5447), .B(n5446), .Z(n5740) );
  NAND U7379 ( .A(n5739), .B(n5740), .Z(n5448) );
  NAND U7380 ( .A(n5449), .B(n5448), .Z(n5451) );
  NANDN U7381 ( .A(n5450), .B(n5451), .Z(n5455) );
  XNOR U7382 ( .A(n5453), .B(n5452), .Z(n5746) );
  NAND U7383 ( .A(n5745), .B(n5746), .Z(n5454) );
  NAND U7384 ( .A(n5455), .B(n5454), .Z(n5458) );
  AND U7385 ( .A(a[46]), .B(b[50]), .Z(n5459) );
  NANDN U7386 ( .A(n5458), .B(n5459), .Z(n5461) );
  XOR U7387 ( .A(n5457), .B(n5456), .Z(n5750) );
  NAND U7388 ( .A(n5750), .B(n5749), .Z(n5460) );
  AND U7389 ( .A(n5461), .B(n5460), .Z(n5463) );
  NANDN U7390 ( .A(n5462), .B(n5463), .Z(n5467) );
  XNOR U7391 ( .A(n5465), .B(n5464), .Z(n5758) );
  NAND U7392 ( .A(n5757), .B(n5758), .Z(n5466) );
  NAND U7393 ( .A(n5467), .B(n5466), .Z(n5471) );
  NANDN U7394 ( .A(n5470), .B(n5471), .Z(n5473) );
  XOR U7395 ( .A(n5469), .B(n5468), .Z(n5763) );
  NANDN U7396 ( .A(n5763), .B(n5764), .Z(n5472) );
  NAND U7397 ( .A(n5473), .B(n5472), .Z(n5476) );
  AND U7398 ( .A(a[49]), .B(b[50]), .Z(n5477) );
  NANDN U7399 ( .A(n5476), .B(n5477), .Z(n5479) );
  XOR U7400 ( .A(n5475), .B(n5474), .Z(n5769) );
  NANDN U7401 ( .A(n5769), .B(n5770), .Z(n5478) );
  AND U7402 ( .A(n5479), .B(n5478), .Z(n10118) );
  XNOR U7403 ( .A(n10120), .B(n10121), .Z(n10198) );
  AND U7404 ( .A(a[51]), .B(b[49]), .Z(n10196) );
  AND U7405 ( .A(a[49]), .B(b[49]), .Z(n5761) );
  NAND U7406 ( .A(a[44]), .B(b[49]), .Z(n5731) );
  AND U7407 ( .A(a[43]), .B(b[49]), .Z(n5725) );
  XOR U7408 ( .A(n5481), .B(n5480), .Z(n5710) );
  AND U7409 ( .A(a[39]), .B(b[49]), .Z(n5705) );
  XOR U7410 ( .A(n5483), .B(n5482), .Z(n5706) );
  NAND U7411 ( .A(n5705), .B(n5706), .Z(n5708) );
  XOR U7412 ( .A(n5485), .B(n5484), .Z(n5696) );
  XOR U7413 ( .A(n5487), .B(n5486), .Z(n5692) );
  AND U7414 ( .A(a[36]), .B(b[49]), .Z(n5691) );
  NANDN U7415 ( .A(n5692), .B(n5691), .Z(n5694) );
  AND U7416 ( .A(a[35]), .B(b[49]), .Z(n5686) );
  NAND U7417 ( .A(a[34]), .B(b[49]), .Z(n5681) );
  XNOR U7418 ( .A(n5489), .B(n5488), .Z(n5682) );
  NANDN U7419 ( .A(n5681), .B(n5682), .Z(n5684) );
  XOR U7420 ( .A(n5491), .B(n5490), .Z(n5677) );
  XOR U7421 ( .A(n5493), .B(n5492), .Z(n5674) );
  XOR U7422 ( .A(n5495), .B(n5494), .Z(n5670) );
  XOR U7423 ( .A(n5497), .B(n5496), .Z(n5666) );
  XOR U7424 ( .A(n5499), .B(n5498), .Z(n5662) );
  XOR U7425 ( .A(n5501), .B(n5500), .Z(n5657) );
  AND U7426 ( .A(a[28]), .B(b[49]), .Z(n5658) );
  NANDN U7427 ( .A(n5657), .B(n5658), .Z(n5660) );
  NAND U7428 ( .A(a[27]), .B(b[49]), .Z(n5653) );
  XNOR U7429 ( .A(n5503), .B(n5502), .Z(n5654) );
  NANDN U7430 ( .A(n5653), .B(n5654), .Z(n5656) );
  XOR U7431 ( .A(n5505), .B(n5504), .Z(n5644) );
  NAND U7432 ( .A(a[23]), .B(b[49]), .Z(n5633) );
  XNOR U7433 ( .A(n5507), .B(n5506), .Z(n5634) );
  NANDN U7434 ( .A(n5633), .B(n5634), .Z(n5636) );
  XOR U7435 ( .A(n5509), .B(n5508), .Z(n5630) );
  XOR U7436 ( .A(n5511), .B(n5510), .Z(n5626) );
  AND U7437 ( .A(a[21]), .B(b[49]), .Z(n5625) );
  NANDN U7438 ( .A(n5626), .B(n5625), .Z(n5628) );
  NAND U7439 ( .A(a[20]), .B(b[49]), .Z(n5621) );
  XNOR U7440 ( .A(n5513), .B(n5512), .Z(n5622) );
  NANDN U7441 ( .A(n5621), .B(n5622), .Z(n5624) );
  XOR U7442 ( .A(n5515), .B(n5514), .Z(n5618) );
  AND U7443 ( .A(a[18]), .B(b[49]), .Z(n5519) );
  XNOR U7444 ( .A(n5517), .B(n5516), .Z(n5518) );
  NANDN U7445 ( .A(n5519), .B(n5518), .Z(n5616) );
  XNOR U7446 ( .A(n5519), .B(n5518), .Z(n5806) );
  XOR U7447 ( .A(n5521), .B(n5520), .Z(n5523) );
  AND U7448 ( .A(a[17]), .B(b[49]), .Z(n5522) );
  NANDN U7449 ( .A(n5523), .B(n5522), .Z(n5614) );
  XOR U7450 ( .A(n5523), .B(n5522), .Z(n5809) );
  XOR U7451 ( .A(n5525), .B(n5524), .Z(n5610) );
  AND U7452 ( .A(a[11]), .B(b[49]), .Z(n5579) );
  XOR U7453 ( .A(n5527), .B(n5526), .Z(n5569) );
  NAND U7454 ( .A(a[7]), .B(b[49]), .Z(n5559) );
  XOR U7455 ( .A(n5529), .B(n5528), .Z(n5560) );
  NANDN U7456 ( .A(n5559), .B(n5560), .Z(n5562) );
  NAND U7457 ( .A(a[0]), .B(b[49]), .Z(n6127) );
  AND U7458 ( .A(a[1]), .B(b[50]), .Z(n5532) );
  NANDN U7459 ( .A(n6127), .B(n5532), .Z(n5827) );
  NANDN U7460 ( .A(n5827), .B(n5530), .Z(n5534) );
  AND U7461 ( .A(a[2]), .B(b[49]), .Z(n5833) );
  NANDN U7462 ( .A(n5832), .B(n5833), .Z(n5533) );
  AND U7463 ( .A(n5534), .B(n5533), .Z(n5537) );
  AND U7464 ( .A(a[3]), .B(b[49]), .Z(n5538) );
  NANDN U7465 ( .A(n5537), .B(n5538), .Z(n5540) );
  XOR U7466 ( .A(n5536), .B(n5535), .Z(n5838) );
  NANDN U7467 ( .A(n5838), .B(n5839), .Z(n5539) );
  AND U7468 ( .A(n5540), .B(n5539), .Z(n5543) );
  NANDN U7469 ( .A(n5543), .B(n5544), .Z(n5546) );
  AND U7470 ( .A(a[4]), .B(b[49]), .Z(n5847) );
  NAND U7471 ( .A(n5847), .B(n5846), .Z(n5545) );
  AND U7472 ( .A(n5546), .B(n5545), .Z(n5547) );
  AND U7473 ( .A(a[5]), .B(b[49]), .Z(n5548) );
  NANDN U7474 ( .A(n5547), .B(n5548), .Z(n5552) );
  XOR U7475 ( .A(n5550), .B(n5549), .Z(n5850) );
  NAND U7476 ( .A(n5851), .B(n5850), .Z(n5551) );
  AND U7477 ( .A(n5552), .B(n5551), .Z(n5555) );
  XOR U7478 ( .A(n5554), .B(n5553), .Z(n5556) );
  NANDN U7479 ( .A(n5555), .B(n5556), .Z(n5558) );
  AND U7480 ( .A(a[6]), .B(b[49]), .Z(n5826) );
  NAND U7481 ( .A(n5826), .B(n5825), .Z(n5557) );
  AND U7482 ( .A(n5558), .B(n5557), .Z(n5862) );
  NANDN U7483 ( .A(n5862), .B(n5863), .Z(n5561) );
  AND U7484 ( .A(n5562), .B(n5561), .Z(n5563) );
  AND U7485 ( .A(a[8]), .B(b[49]), .Z(n5564) );
  NANDN U7486 ( .A(n5563), .B(n5564), .Z(n5568) );
  NAND U7487 ( .A(n5824), .B(n5823), .Z(n5567) );
  AND U7488 ( .A(n5568), .B(n5567), .Z(n5570) );
  NANDN U7489 ( .A(n5569), .B(n5570), .Z(n5572) );
  AND U7490 ( .A(a[9]), .B(b[49]), .Z(n5870) );
  NANDN U7491 ( .A(n5870), .B(n5871), .Z(n5571) );
  AND U7492 ( .A(n5572), .B(n5571), .Z(n5575) );
  NAND U7493 ( .A(n5575), .B(n5576), .Z(n5578) );
  AND U7494 ( .A(a[10]), .B(b[49]), .Z(n5879) );
  XOR U7495 ( .A(n5576), .B(n5575), .Z(n5878) );
  NAND U7496 ( .A(n5879), .B(n5878), .Z(n5577) );
  AND U7497 ( .A(n5578), .B(n5577), .Z(n5580) );
  NANDN U7498 ( .A(n5579), .B(n5580), .Z(n5584) );
  XNOR U7499 ( .A(n5582), .B(n5581), .Z(n5821) );
  NAND U7500 ( .A(n5822), .B(n5821), .Z(n5583) );
  AND U7501 ( .A(n5584), .B(n5583), .Z(n5587) );
  NANDN U7502 ( .A(n5587), .B(n5588), .Z(n5590) );
  AND U7503 ( .A(a[12]), .B(b[49]), .Z(n5819) );
  NANDN U7504 ( .A(n5819), .B(n5820), .Z(n5589) );
  NAND U7505 ( .A(n5590), .B(n5589), .Z(n5593) );
  XOR U7506 ( .A(n5592), .B(n5591), .Z(n5594) );
  NANDN U7507 ( .A(n5593), .B(n5594), .Z(n5596) );
  AND U7508 ( .A(a[13]), .B(b[49]), .Z(n5816) );
  NAND U7509 ( .A(n5816), .B(n5815), .Z(n5595) );
  AND U7510 ( .A(n5596), .B(n5595), .Z(n5597) );
  AND U7511 ( .A(a[14]), .B(b[49]), .Z(n5598) );
  NANDN U7512 ( .A(n5597), .B(n5598), .Z(n5602) );
  NAND U7513 ( .A(n5814), .B(n5813), .Z(n5601) );
  AND U7514 ( .A(n5602), .B(n5601), .Z(n5603) );
  AND U7515 ( .A(a[15]), .B(b[49]), .Z(n5604) );
  NANDN U7516 ( .A(n5603), .B(n5604), .Z(n5608) );
  XOR U7517 ( .A(n5606), .B(n5605), .Z(n5898) );
  NAND U7518 ( .A(n5899), .B(n5898), .Z(n5607) );
  AND U7519 ( .A(n5608), .B(n5607), .Z(n5609) );
  NANDN U7520 ( .A(n5610), .B(n5609), .Z(n5612) );
  XOR U7521 ( .A(n5610), .B(n5609), .Z(n5811) );
  AND U7522 ( .A(a[16]), .B(b[49]), .Z(n5812) );
  OR U7523 ( .A(n5811), .B(n5812), .Z(n5611) );
  AND U7524 ( .A(n5612), .B(n5611), .Z(n5810) );
  NANDN U7525 ( .A(n5809), .B(n5810), .Z(n5613) );
  AND U7526 ( .A(n5614), .B(n5613), .Z(n5805) );
  NAND U7527 ( .A(n5806), .B(n5805), .Z(n5615) );
  AND U7528 ( .A(n5616), .B(n5615), .Z(n5617) );
  NANDN U7529 ( .A(n5618), .B(n5617), .Z(n5620) );
  XNOR U7530 ( .A(n5618), .B(n5617), .Z(n5804) );
  AND U7531 ( .A(a[19]), .B(b[49]), .Z(n5803) );
  NAND U7532 ( .A(n5804), .B(n5803), .Z(n5619) );
  AND U7533 ( .A(n5620), .B(n5619), .Z(n5802) );
  XNOR U7534 ( .A(n5622), .B(n5621), .Z(n5801) );
  NANDN U7535 ( .A(n5802), .B(n5801), .Z(n5623) );
  AND U7536 ( .A(n5624), .B(n5623), .Z(n5800) );
  XNOR U7537 ( .A(n5626), .B(n5625), .Z(n5799) );
  NANDN U7538 ( .A(n5800), .B(n5799), .Z(n5627) );
  NAND U7539 ( .A(n5628), .B(n5627), .Z(n5629) );
  NANDN U7540 ( .A(n5630), .B(n5629), .Z(n5632) );
  NAND U7541 ( .A(a[22]), .B(b[49]), .Z(n5924) );
  XNOR U7542 ( .A(n5630), .B(n5629), .Z(n5925) );
  NANDN U7543 ( .A(n5924), .B(n5925), .Z(n5631) );
  AND U7544 ( .A(n5632), .B(n5631), .Z(n5931) );
  XNOR U7545 ( .A(n5634), .B(n5633), .Z(n5930) );
  NANDN U7546 ( .A(n5931), .B(n5930), .Z(n5635) );
  AND U7547 ( .A(n5636), .B(n5635), .Z(n5640) );
  AND U7548 ( .A(a[24]), .B(b[49]), .Z(n5639) );
  NANDN U7549 ( .A(n5640), .B(n5639), .Z(n5642) );
  XOR U7550 ( .A(n5638), .B(n5637), .Z(n5797) );
  XNOR U7551 ( .A(n5640), .B(n5639), .Z(n5798) );
  NANDN U7552 ( .A(n5797), .B(n5798), .Z(n5641) );
  AND U7553 ( .A(n5642), .B(n5641), .Z(n5643) );
  NANDN U7554 ( .A(n5644), .B(n5643), .Z(n5646) );
  XOR U7555 ( .A(n5644), .B(n5643), .Z(n5795) );
  AND U7556 ( .A(a[25]), .B(b[49]), .Z(n5796) );
  OR U7557 ( .A(n5795), .B(n5796), .Z(n5645) );
  NAND U7558 ( .A(n5646), .B(n5645), .Z(n5649) );
  XNOR U7559 ( .A(n5648), .B(n5647), .Z(n5650) );
  NANDN U7560 ( .A(n5649), .B(n5650), .Z(n5652) );
  XNOR U7561 ( .A(n5650), .B(n5649), .Z(n5794) );
  AND U7562 ( .A(a[26]), .B(b[49]), .Z(n5793) );
  NAND U7563 ( .A(n5794), .B(n5793), .Z(n5651) );
  AND U7564 ( .A(n5652), .B(n5651), .Z(n5792) );
  XNOR U7565 ( .A(n5654), .B(n5653), .Z(n5791) );
  NANDN U7566 ( .A(n5792), .B(n5791), .Z(n5655) );
  AND U7567 ( .A(n5656), .B(n5655), .Z(n5953) );
  XNOR U7568 ( .A(n5658), .B(n5657), .Z(n5952) );
  NANDN U7569 ( .A(n5953), .B(n5952), .Z(n5659) );
  AND U7570 ( .A(n5660), .B(n5659), .Z(n5661) );
  NANDN U7571 ( .A(n5662), .B(n5661), .Z(n5664) );
  AND U7572 ( .A(a[29]), .B(b[49]), .Z(n5790) );
  XNOR U7573 ( .A(n5662), .B(n5661), .Z(n5789) );
  NANDN U7574 ( .A(n5790), .B(n5789), .Z(n5663) );
  NAND U7575 ( .A(n5664), .B(n5663), .Z(n5665) );
  NANDN U7576 ( .A(n5666), .B(n5665), .Z(n5668) );
  XOR U7577 ( .A(n5666), .B(n5665), .Z(n5787) );
  AND U7578 ( .A(a[30]), .B(b[49]), .Z(n5788) );
  OR U7579 ( .A(n5787), .B(n5788), .Z(n5667) );
  AND U7580 ( .A(n5668), .B(n5667), .Z(n5669) );
  NANDN U7581 ( .A(n5670), .B(n5669), .Z(n5672) );
  NAND U7582 ( .A(a[31]), .B(b[49]), .Z(n5785) );
  XNOR U7583 ( .A(n5670), .B(n5669), .Z(n5786) );
  NANDN U7584 ( .A(n5785), .B(n5786), .Z(n5671) );
  AND U7585 ( .A(n5672), .B(n5671), .Z(n5673) );
  NANDN U7586 ( .A(n5674), .B(n5673), .Z(n5676) );
  XOR U7587 ( .A(n5674), .B(n5673), .Z(n5972) );
  AND U7588 ( .A(a[32]), .B(b[49]), .Z(n5973) );
  OR U7589 ( .A(n5972), .B(n5973), .Z(n5675) );
  AND U7590 ( .A(n5676), .B(n5675), .Z(n5678) );
  NANDN U7591 ( .A(n5677), .B(n5678), .Z(n5680) );
  NAND U7592 ( .A(a[33]), .B(b[49]), .Z(n5976) );
  XNOR U7593 ( .A(n5678), .B(n5677), .Z(n5977) );
  NANDN U7594 ( .A(n5976), .B(n5977), .Z(n5679) );
  AND U7595 ( .A(n5680), .B(n5679), .Z(n5784) );
  XNOR U7596 ( .A(n5682), .B(n5681), .Z(n5783) );
  NANDN U7597 ( .A(n5784), .B(n5783), .Z(n5683) );
  AND U7598 ( .A(n5684), .B(n5683), .Z(n5685) );
  NANDN U7599 ( .A(n5686), .B(n5685), .Z(n5690) );
  XNOR U7600 ( .A(n5686), .B(n5685), .Z(n5987) );
  XNOR U7601 ( .A(n5688), .B(n5687), .Z(n5986) );
  NAND U7602 ( .A(n5987), .B(n5986), .Z(n5689) );
  NAND U7603 ( .A(n5690), .B(n5689), .Z(n5992) );
  XNOR U7604 ( .A(n5692), .B(n5691), .Z(n5993) );
  NANDN U7605 ( .A(n5992), .B(n5993), .Z(n5693) );
  AND U7606 ( .A(n5694), .B(n5693), .Z(n5695) );
  NANDN U7607 ( .A(n5696), .B(n5695), .Z(n5698) );
  AND U7608 ( .A(a[37]), .B(b[49]), .Z(n5782) );
  XNOR U7609 ( .A(n5696), .B(n5695), .Z(n5781) );
  NANDN U7610 ( .A(n5782), .B(n5781), .Z(n5697) );
  AND U7611 ( .A(n5698), .B(n5697), .Z(n5702) );
  XNOR U7612 ( .A(n5700), .B(n5699), .Z(n5701) );
  NAND U7613 ( .A(n5702), .B(n5701), .Z(n5704) );
  NAND U7614 ( .A(a[38]), .B(b[49]), .Z(n5779) );
  XOR U7615 ( .A(n5702), .B(n5701), .Z(n5780) );
  NANDN U7616 ( .A(n5779), .B(n5780), .Z(n5703) );
  AND U7617 ( .A(n5704), .B(n5703), .Z(n5778) );
  XOR U7618 ( .A(n5706), .B(n5705), .Z(n5777) );
  NANDN U7619 ( .A(n5778), .B(n5777), .Z(n5707) );
  NAND U7620 ( .A(n5708), .B(n5707), .Z(n5709) );
  NAND U7621 ( .A(n5710), .B(n5709), .Z(n5712) );
  XOR U7622 ( .A(n5710), .B(n5709), .Z(n5776) );
  AND U7623 ( .A(a[40]), .B(b[49]), .Z(n5775) );
  NAND U7624 ( .A(n5776), .B(n5775), .Z(n5711) );
  AND U7625 ( .A(n5712), .B(n5711), .Z(n5714) );
  AND U7626 ( .A(a[41]), .B(b[49]), .Z(n5713) );
  NANDN U7627 ( .A(n5714), .B(n5713), .Z(n5718) );
  XNOR U7628 ( .A(n5714), .B(n5713), .Z(n5774) );
  XOR U7629 ( .A(n5716), .B(n5715), .Z(n5773) );
  NAND U7630 ( .A(n5774), .B(n5773), .Z(n5717) );
  AND U7631 ( .A(n5718), .B(n5717), .Z(n5719) );
  AND U7632 ( .A(a[42]), .B(b[49]), .Z(n5720) );
  NANDN U7633 ( .A(n5719), .B(n5720), .Z(n5724) );
  XNOR U7634 ( .A(n5722), .B(n5721), .Z(n6021) );
  NAND U7635 ( .A(n6020), .B(n6021), .Z(n5723) );
  AND U7636 ( .A(n5724), .B(n5723), .Z(n5726) );
  NANDN U7637 ( .A(n5725), .B(n5726), .Z(n5730) );
  NAND U7638 ( .A(n6025), .B(n6024), .Z(n5729) );
  AND U7639 ( .A(n5730), .B(n5729), .Z(n5732) );
  NANDN U7640 ( .A(n5731), .B(n5732), .Z(n5736) );
  NAND U7641 ( .A(n6031), .B(n6030), .Z(n5735) );
  AND U7642 ( .A(n5736), .B(n5735), .Z(n5737) );
  AND U7643 ( .A(a[45]), .B(b[49]), .Z(n5738) );
  NANDN U7644 ( .A(n5737), .B(n5738), .Z(n5742) );
  XNOR U7645 ( .A(n5740), .B(n5739), .Z(n6039) );
  NAND U7646 ( .A(n6038), .B(n6039), .Z(n5741) );
  AND U7647 ( .A(n5742), .B(n5741), .Z(n5743) );
  AND U7648 ( .A(a[46]), .B(b[49]), .Z(n5744) );
  NANDN U7649 ( .A(n5743), .B(n5744), .Z(n5748) );
  XNOR U7650 ( .A(n5746), .B(n5745), .Z(n6045) );
  NAND U7651 ( .A(n6044), .B(n6045), .Z(n5747) );
  AND U7652 ( .A(n5748), .B(n5747), .Z(n5751) );
  AND U7653 ( .A(a[47]), .B(b[49]), .Z(n5752) );
  NANDN U7654 ( .A(n5751), .B(n5752), .Z(n5754) );
  XOR U7655 ( .A(n5750), .B(n5749), .Z(n6049) );
  NAND U7656 ( .A(n6049), .B(n6048), .Z(n5753) );
  AND U7657 ( .A(n5754), .B(n5753), .Z(n5755) );
  AND U7658 ( .A(a[48]), .B(b[49]), .Z(n5756) );
  NANDN U7659 ( .A(n5755), .B(n5756), .Z(n5760) );
  XNOR U7660 ( .A(n5758), .B(n5757), .Z(n6057) );
  NAND U7661 ( .A(n6056), .B(n6057), .Z(n5759) );
  AND U7662 ( .A(n5760), .B(n5759), .Z(n5762) );
  NANDN U7663 ( .A(n5761), .B(n5762), .Z(n5766) );
  NAND U7664 ( .A(n6061), .B(n6060), .Z(n5765) );
  NAND U7665 ( .A(n5766), .B(n5765), .Z(n5767) );
  AND U7666 ( .A(a[50]), .B(b[49]), .Z(n5768) );
  NANDN U7667 ( .A(n5767), .B(n5768), .Z(n5772) );
  NAND U7668 ( .A(n6067), .B(n6066), .Z(n5771) );
  AND U7669 ( .A(n5772), .B(n5771), .Z(n10197) );
  XNOR U7670 ( .A(n10198), .B(n10199), .Z(n10204) );
  AND U7671 ( .A(a[52]), .B(b[48]), .Z(n10203) );
  AND U7672 ( .A(a[51]), .B(b[48]), .Z(n6068) );
  AND U7673 ( .A(a[49]), .B(b[48]), .Z(n6054) );
  AND U7674 ( .A(a[48]), .B(b[48]), .Z(n6050) );
  AND U7675 ( .A(a[47]), .B(b[48]), .Z(n6042) );
  AND U7676 ( .A(a[46]), .B(b[48]), .Z(n6036) );
  AND U7677 ( .A(a[45]), .B(b[48]), .Z(n6032) );
  NAND U7678 ( .A(a[44]), .B(b[48]), .Z(n6026) );
  AND U7679 ( .A(a[43]), .B(b[48]), .Z(n6018) );
  XOR U7680 ( .A(n5774), .B(n5773), .Z(n6015) );
  XOR U7681 ( .A(n5776), .B(n5775), .Z(n6011) );
  NAND U7682 ( .A(a[40]), .B(b[48]), .Z(n6006) );
  XNOR U7683 ( .A(n5778), .B(n5777), .Z(n6007) );
  NANDN U7684 ( .A(n6006), .B(n6007), .Z(n6009) );
  NAND U7685 ( .A(a[39]), .B(b[48]), .Z(n6002) );
  XNOR U7686 ( .A(n5780), .B(n5779), .Z(n6003) );
  NANDN U7687 ( .A(n6002), .B(n6003), .Z(n6005) );
  XOR U7688 ( .A(n5782), .B(n5781), .Z(n5999) );
  AND U7689 ( .A(a[38]), .B(b[48]), .Z(n5998) );
  NAND U7690 ( .A(n5999), .B(n5998), .Z(n6001) );
  NAND U7691 ( .A(a[35]), .B(b[48]), .Z(n5982) );
  XNOR U7692 ( .A(n5784), .B(n5783), .Z(n5983) );
  NANDN U7693 ( .A(n5982), .B(n5983), .Z(n5985) );
  XOR U7694 ( .A(n5786), .B(n5785), .Z(n5966) );
  AND U7695 ( .A(a[32]), .B(b[48]), .Z(n5967) );
  NANDN U7696 ( .A(n5966), .B(n5967), .Z(n5969) );
  XOR U7697 ( .A(n5788), .B(n5787), .Z(n5963) );
  AND U7698 ( .A(a[31]), .B(b[48]), .Z(n5962) );
  NANDN U7699 ( .A(n5963), .B(n5962), .Z(n5965) );
  XOR U7700 ( .A(n5790), .B(n5789), .Z(n5958) );
  XOR U7701 ( .A(n5792), .B(n5791), .Z(n5948) );
  AND U7702 ( .A(a[28]), .B(b[48]), .Z(n5949) );
  NANDN U7703 ( .A(n5948), .B(n5949), .Z(n5951) );
  XOR U7704 ( .A(n5794), .B(n5793), .Z(n5945) );
  XOR U7705 ( .A(n5796), .B(n5795), .Z(n5941) );
  AND U7706 ( .A(a[26]), .B(b[48]), .Z(n5940) );
  NANDN U7707 ( .A(n5941), .B(n5940), .Z(n5943) );
  XOR U7708 ( .A(n5798), .B(n5797), .Z(n5936) );
  AND U7709 ( .A(a[25]), .B(b[48]), .Z(n5937) );
  NANDN U7710 ( .A(n5936), .B(n5937), .Z(n5939) );
  XOR U7711 ( .A(n5800), .B(n5799), .Z(n5920) );
  AND U7712 ( .A(a[22]), .B(b[48]), .Z(n5921) );
  NANDN U7713 ( .A(n5920), .B(n5921), .Z(n5923) );
  NAND U7714 ( .A(a[21]), .B(b[48]), .Z(n5916) );
  XNOR U7715 ( .A(n5802), .B(n5801), .Z(n5917) );
  NANDN U7716 ( .A(n5916), .B(n5917), .Z(n5919) );
  AND U7717 ( .A(a[20]), .B(b[48]), .Z(n5913) );
  XNOR U7718 ( .A(n5804), .B(n5803), .Z(n5912) );
  NANDN U7719 ( .A(n5913), .B(n5912), .Z(n5915) );
  XOR U7720 ( .A(n5806), .B(n5805), .Z(n5808) );
  AND U7721 ( .A(a[19]), .B(b[48]), .Z(n5807) );
  NANDN U7722 ( .A(n5808), .B(n5807), .Z(n5911) );
  XOR U7723 ( .A(n5808), .B(n5807), .Z(n6110) );
  XOR U7724 ( .A(n5810), .B(n5809), .Z(n5906) );
  AND U7725 ( .A(a[18]), .B(b[48]), .Z(n5907) );
  NANDN U7726 ( .A(n5906), .B(n5907), .Z(n5909) );
  XOR U7727 ( .A(n5812), .B(n5811), .Z(n5903) );
  NAND U7728 ( .A(a[15]), .B(b[48]), .Z(n5892) );
  XOR U7729 ( .A(n5814), .B(n5813), .Z(n5893) );
  NANDN U7730 ( .A(n5892), .B(n5893), .Z(n5895) );
  NAND U7731 ( .A(a[14]), .B(b[48]), .Z(n5817) );
  XOR U7732 ( .A(n5816), .B(n5815), .Z(n5818) );
  NANDN U7733 ( .A(n5817), .B(n5818), .Z(n5891) );
  XOR U7734 ( .A(n5822), .B(n5821), .Z(n5882) );
  AND U7735 ( .A(a[11]), .B(b[48]), .Z(n5876) );
  XOR U7736 ( .A(n5824), .B(n5823), .Z(n5866) );
  NAND U7737 ( .A(a[7]), .B(b[48]), .Z(n5856) );
  XOR U7738 ( .A(n5826), .B(n5825), .Z(n5857) );
  NANDN U7739 ( .A(n5856), .B(n5857), .Z(n5859) );
  AND U7740 ( .A(a[5]), .B(b[48]), .Z(n5844) );
  NAND U7741 ( .A(a[0]), .B(b[48]), .Z(n6428) );
  AND U7742 ( .A(a[1]), .B(b[49]), .Z(n5829) );
  NANDN U7743 ( .A(n6428), .B(n5829), .Z(n6126) );
  NANDN U7744 ( .A(n6126), .B(n5827), .Z(n5831) );
  AND U7745 ( .A(a[2]), .B(b[48]), .Z(n6132) );
  NANDN U7746 ( .A(n6131), .B(n6132), .Z(n5830) );
  AND U7747 ( .A(n5831), .B(n5830), .Z(n5834) );
  AND U7748 ( .A(a[3]), .B(b[48]), .Z(n5835) );
  NANDN U7749 ( .A(n5834), .B(n5835), .Z(n5837) );
  XOR U7750 ( .A(n5833), .B(n5832), .Z(n6137) );
  NANDN U7751 ( .A(n6137), .B(n6138), .Z(n5836) );
  AND U7752 ( .A(n5837), .B(n5836), .Z(n5840) );
  NANDN U7753 ( .A(n5840), .B(n5841), .Z(n5843) );
  NAND U7754 ( .A(a[4]), .B(b[48]), .Z(n6145) );
  NANDN U7755 ( .A(n6145), .B(n6146), .Z(n5842) );
  AND U7756 ( .A(n5843), .B(n5842), .Z(n5845) );
  NANDN U7757 ( .A(n5844), .B(n5845), .Z(n5849) );
  XNOR U7758 ( .A(n5847), .B(n5846), .Z(n6124) );
  NAND U7759 ( .A(n6125), .B(n6124), .Z(n5848) );
  NAND U7760 ( .A(n5849), .B(n5848), .Z(n5852) );
  XOR U7761 ( .A(n5851), .B(n5850), .Z(n5853) );
  NANDN U7762 ( .A(n5852), .B(n5853), .Z(n5855) );
  AND U7763 ( .A(a[6]), .B(b[48]), .Z(n6123) );
  NAND U7764 ( .A(n6123), .B(n6122), .Z(n5854) );
  AND U7765 ( .A(n5855), .B(n5854), .Z(n6159) );
  NANDN U7766 ( .A(n6159), .B(n6160), .Z(n5858) );
  AND U7767 ( .A(n5859), .B(n5858), .Z(n5860) );
  AND U7768 ( .A(a[8]), .B(b[48]), .Z(n5861) );
  NANDN U7769 ( .A(n5860), .B(n5861), .Z(n5865) );
  NAND U7770 ( .A(n6121), .B(n6120), .Z(n5864) );
  AND U7771 ( .A(n5865), .B(n5864), .Z(n5867) );
  NANDN U7772 ( .A(n5866), .B(n5867), .Z(n5869) );
  AND U7773 ( .A(a[9]), .B(b[48]), .Z(n6167) );
  NANDN U7774 ( .A(n6167), .B(n6168), .Z(n5868) );
  AND U7775 ( .A(n5869), .B(n5868), .Z(n5872) );
  NAND U7776 ( .A(n5872), .B(n5873), .Z(n5875) );
  AND U7777 ( .A(a[10]), .B(b[48]), .Z(n6174) );
  XOR U7778 ( .A(n5873), .B(n5872), .Z(n6173) );
  NAND U7779 ( .A(n6174), .B(n6173), .Z(n5874) );
  AND U7780 ( .A(n5875), .B(n5874), .Z(n5877) );
  NANDN U7781 ( .A(n5876), .B(n5877), .Z(n5881) );
  XNOR U7782 ( .A(n5879), .B(n5878), .Z(n6118) );
  NAND U7783 ( .A(n6119), .B(n6118), .Z(n5880) );
  AND U7784 ( .A(n5881), .B(n5880), .Z(n5883) );
  NANDN U7785 ( .A(n5882), .B(n5883), .Z(n5885) );
  AND U7786 ( .A(a[12]), .B(b[48]), .Z(n6184) );
  NAND U7787 ( .A(n6184), .B(n6183), .Z(n5884) );
  NAND U7788 ( .A(n5885), .B(n5884), .Z(n5886) );
  NAND U7789 ( .A(n5887), .B(n5886), .Z(n5889) );
  AND U7790 ( .A(a[13]), .B(b[48]), .Z(n6117) );
  XOR U7791 ( .A(n5887), .B(n5886), .Z(n6116) );
  NAND U7792 ( .A(n6117), .B(n6116), .Z(n5888) );
  NAND U7793 ( .A(n5889), .B(n5888), .Z(n6114) );
  NAND U7794 ( .A(n6115), .B(n6114), .Z(n5890) );
  AND U7795 ( .A(n5891), .B(n5890), .Z(n6199) );
  NANDN U7796 ( .A(n6199), .B(n6200), .Z(n5894) );
  AND U7797 ( .A(n5895), .B(n5894), .Z(n5896) );
  AND U7798 ( .A(a[16]), .B(b[48]), .Z(n5897) );
  NANDN U7799 ( .A(n5896), .B(n5897), .Z(n5901) );
  XOR U7800 ( .A(n5899), .B(n5898), .Z(n6203) );
  NAND U7801 ( .A(n6204), .B(n6203), .Z(n5900) );
  NAND U7802 ( .A(n5901), .B(n5900), .Z(n5902) );
  NANDN U7803 ( .A(n5903), .B(n5902), .Z(n5905) );
  NAND U7804 ( .A(a[17]), .B(b[48]), .Z(n6112) );
  XNOR U7805 ( .A(n5903), .B(n5902), .Z(n6113) );
  NANDN U7806 ( .A(n6112), .B(n6113), .Z(n5904) );
  AND U7807 ( .A(n5905), .B(n5904), .Z(n6214) );
  XNOR U7808 ( .A(n5907), .B(n5906), .Z(n6213) );
  NANDN U7809 ( .A(n6214), .B(n6213), .Z(n5908) );
  AND U7810 ( .A(n5909), .B(n5908), .Z(n6111) );
  OR U7811 ( .A(n6110), .B(n6111), .Z(n5910) );
  NAND U7812 ( .A(n5911), .B(n5910), .Z(n6106) );
  XNOR U7813 ( .A(n5913), .B(n5912), .Z(n6107) );
  NANDN U7814 ( .A(n6106), .B(n6107), .Z(n5914) );
  NAND U7815 ( .A(n5915), .B(n5914), .Z(n6104) );
  XNOR U7816 ( .A(n5917), .B(n5916), .Z(n6105) );
  NANDN U7817 ( .A(n6104), .B(n6105), .Z(n5918) );
  AND U7818 ( .A(n5919), .B(n5918), .Z(n6230) );
  XNOR U7819 ( .A(n5921), .B(n5920), .Z(n6229) );
  NANDN U7820 ( .A(n6230), .B(n6229), .Z(n5922) );
  AND U7821 ( .A(n5923), .B(n5922), .Z(n5927) );
  XNOR U7822 ( .A(n5925), .B(n5924), .Z(n5926) );
  NANDN U7823 ( .A(n5927), .B(n5926), .Z(n5929) );
  XNOR U7824 ( .A(n5927), .B(n5926), .Z(n6103) );
  AND U7825 ( .A(a[23]), .B(b[48]), .Z(n6102) );
  NAND U7826 ( .A(n6103), .B(n6102), .Z(n5928) );
  AND U7827 ( .A(n5929), .B(n5928), .Z(n5933) );
  XNOR U7828 ( .A(n5931), .B(n5930), .Z(n5932) );
  NANDN U7829 ( .A(n5933), .B(n5932), .Z(n5935) );
  NAND U7830 ( .A(a[24]), .B(b[48]), .Z(n6100) );
  XNOR U7831 ( .A(n5933), .B(n5932), .Z(n6101) );
  NANDN U7832 ( .A(n6100), .B(n6101), .Z(n5934) );
  AND U7833 ( .A(n5935), .B(n5934), .Z(n6244) );
  XNOR U7834 ( .A(n5937), .B(n5936), .Z(n6243) );
  NANDN U7835 ( .A(n6244), .B(n6243), .Z(n5938) );
  AND U7836 ( .A(n5939), .B(n5938), .Z(n6099) );
  XNOR U7837 ( .A(n5941), .B(n5940), .Z(n6098) );
  NANDN U7838 ( .A(n6099), .B(n6098), .Z(n5942) );
  AND U7839 ( .A(n5943), .B(n5942), .Z(n5944) );
  NANDN U7840 ( .A(n5945), .B(n5944), .Z(n5947) );
  XOR U7841 ( .A(n5945), .B(n5944), .Z(n6096) );
  AND U7842 ( .A(a[27]), .B(b[48]), .Z(n6097) );
  OR U7843 ( .A(n6096), .B(n6097), .Z(n5946) );
  NAND U7844 ( .A(n5947), .B(n5946), .Z(n6094) );
  XNOR U7845 ( .A(n5949), .B(n5948), .Z(n6095) );
  NANDN U7846 ( .A(n6094), .B(n6095), .Z(n5950) );
  AND U7847 ( .A(n5951), .B(n5950), .Z(n5955) );
  XNOR U7848 ( .A(n5953), .B(n5952), .Z(n5954) );
  NANDN U7849 ( .A(n5955), .B(n5954), .Z(n5957) );
  XNOR U7850 ( .A(n5955), .B(n5954), .Z(n6093) );
  AND U7851 ( .A(a[29]), .B(b[48]), .Z(n6092) );
  NAND U7852 ( .A(n6093), .B(n6092), .Z(n5956) );
  AND U7853 ( .A(n5957), .B(n5956), .Z(n5959) );
  NANDN U7854 ( .A(n5958), .B(n5959), .Z(n5961) );
  XOR U7855 ( .A(n5959), .B(n5958), .Z(n6090) );
  AND U7856 ( .A(a[30]), .B(b[48]), .Z(n6091) );
  OR U7857 ( .A(n6090), .B(n6091), .Z(n5960) );
  NAND U7858 ( .A(n5961), .B(n5960), .Z(n6088) );
  XNOR U7859 ( .A(n5963), .B(n5962), .Z(n6089) );
  NANDN U7860 ( .A(n6088), .B(n6089), .Z(n5964) );
  AND U7861 ( .A(n5965), .B(n5964), .Z(n6274) );
  XNOR U7862 ( .A(n5967), .B(n5966), .Z(n6273) );
  NANDN U7863 ( .A(n6274), .B(n6273), .Z(n5968) );
  AND U7864 ( .A(n5969), .B(n5968), .Z(n5971) );
  AND U7865 ( .A(a[33]), .B(b[48]), .Z(n5970) );
  NANDN U7866 ( .A(n5971), .B(n5970), .Z(n5975) );
  XOR U7867 ( .A(n5971), .B(n5970), .Z(n6086) );
  XOR U7868 ( .A(n5973), .B(n5972), .Z(n6087) );
  OR U7869 ( .A(n6086), .B(n6087), .Z(n5974) );
  AND U7870 ( .A(n5975), .B(n5974), .Z(n5979) );
  XNOR U7871 ( .A(n5977), .B(n5976), .Z(n5978) );
  NANDN U7872 ( .A(n5979), .B(n5978), .Z(n5981) );
  NAND U7873 ( .A(a[34]), .B(b[48]), .Z(n6283) );
  XNOR U7874 ( .A(n5979), .B(n5978), .Z(n6284) );
  NANDN U7875 ( .A(n6283), .B(n6284), .Z(n5980) );
  AND U7876 ( .A(n5981), .B(n5980), .Z(n6083) );
  XNOR U7877 ( .A(n5983), .B(n5982), .Z(n6082) );
  NANDN U7878 ( .A(n6083), .B(n6082), .Z(n5984) );
  AND U7879 ( .A(n5985), .B(n5984), .Z(n5989) );
  AND U7880 ( .A(a[36]), .B(b[48]), .Z(n5988) );
  NANDN U7881 ( .A(n5989), .B(n5988), .Z(n5991) );
  XOR U7882 ( .A(n5987), .B(n5986), .Z(n6292) );
  XNOR U7883 ( .A(n5989), .B(n5988), .Z(n6291) );
  NANDN U7884 ( .A(n6292), .B(n6291), .Z(n5990) );
  AND U7885 ( .A(n5991), .B(n5990), .Z(n5995) );
  XNOR U7886 ( .A(n5993), .B(n5992), .Z(n5994) );
  NANDN U7887 ( .A(n5995), .B(n5994), .Z(n5997) );
  NAND U7888 ( .A(a[37]), .B(b[48]), .Z(n6080) );
  XNOR U7889 ( .A(n5995), .B(n5994), .Z(n6081) );
  NANDN U7890 ( .A(n6080), .B(n6081), .Z(n5996) );
  AND U7891 ( .A(n5997), .B(n5996), .Z(n6079) );
  XOR U7892 ( .A(n5999), .B(n5998), .Z(n6078) );
  NANDN U7893 ( .A(n6079), .B(n6078), .Z(n6000) );
  AND U7894 ( .A(n6001), .B(n6000), .Z(n6077) );
  XNOR U7895 ( .A(n6003), .B(n6002), .Z(n6076) );
  NANDN U7896 ( .A(n6077), .B(n6076), .Z(n6004) );
  AND U7897 ( .A(n6005), .B(n6004), .Z(n6308) );
  XNOR U7898 ( .A(n6007), .B(n6006), .Z(n6307) );
  NANDN U7899 ( .A(n6308), .B(n6307), .Z(n6008) );
  AND U7900 ( .A(n6009), .B(n6008), .Z(n6010) );
  NANDN U7901 ( .A(n6011), .B(n6010), .Z(n6013) );
  AND U7902 ( .A(a[41]), .B(b[48]), .Z(n6075) );
  XNOR U7903 ( .A(n6011), .B(n6010), .Z(n6074) );
  NANDN U7904 ( .A(n6075), .B(n6074), .Z(n6012) );
  NAND U7905 ( .A(n6013), .B(n6012), .Z(n6014) );
  NANDN U7906 ( .A(n6015), .B(n6014), .Z(n6017) );
  AND U7907 ( .A(a[42]), .B(b[48]), .Z(n6320) );
  XNOR U7908 ( .A(n6015), .B(n6014), .Z(n6319) );
  NANDN U7909 ( .A(n6320), .B(n6319), .Z(n6016) );
  NAND U7910 ( .A(n6017), .B(n6016), .Z(n6019) );
  NANDN U7911 ( .A(n6018), .B(n6019), .Z(n6023) );
  XNOR U7912 ( .A(n6021), .B(n6020), .Z(n6073) );
  NAND U7913 ( .A(n6072), .B(n6073), .Z(n6022) );
  AND U7914 ( .A(n6023), .B(n6022), .Z(n6027) );
  NANDN U7915 ( .A(n6026), .B(n6027), .Z(n6029) );
  XOR U7916 ( .A(n6025), .B(n6024), .Z(n6329) );
  NANDN U7917 ( .A(n6329), .B(n6330), .Z(n6028) );
  AND U7918 ( .A(n6029), .B(n6028), .Z(n6033) );
  NANDN U7919 ( .A(n6032), .B(n6033), .Z(n6035) );
  XOR U7920 ( .A(n6031), .B(n6030), .Z(n6335) );
  NANDN U7921 ( .A(n6335), .B(n6336), .Z(n6034) );
  NAND U7922 ( .A(n6035), .B(n6034), .Z(n6037) );
  NANDN U7923 ( .A(n6036), .B(n6037), .Z(n6041) );
  XNOR U7924 ( .A(n6039), .B(n6038), .Z(n6342) );
  NAND U7925 ( .A(n6341), .B(n6342), .Z(n6040) );
  NAND U7926 ( .A(n6041), .B(n6040), .Z(n6043) );
  NANDN U7927 ( .A(n6042), .B(n6043), .Z(n6047) );
  XNOR U7928 ( .A(n6045), .B(n6044), .Z(n6348) );
  NAND U7929 ( .A(n6347), .B(n6348), .Z(n6046) );
  NAND U7930 ( .A(n6047), .B(n6046), .Z(n6051) );
  NANDN U7931 ( .A(n6050), .B(n6051), .Z(n6053) );
  XOR U7932 ( .A(n6049), .B(n6048), .Z(n6353) );
  NANDN U7933 ( .A(n6353), .B(n6354), .Z(n6052) );
  NAND U7934 ( .A(n6053), .B(n6052), .Z(n6055) );
  NANDN U7935 ( .A(n6054), .B(n6055), .Z(n6059) );
  XNOR U7936 ( .A(n6057), .B(n6056), .Z(n6360) );
  NAND U7937 ( .A(n6359), .B(n6360), .Z(n6058) );
  NAND U7938 ( .A(n6059), .B(n6058), .Z(n6062) );
  AND U7939 ( .A(a[50]), .B(b[48]), .Z(n6063) );
  NANDN U7940 ( .A(n6062), .B(n6063), .Z(n6065) );
  XOR U7941 ( .A(n6061), .B(n6060), .Z(n6365) );
  NANDN U7942 ( .A(n6365), .B(n6366), .Z(n6064) );
  AND U7943 ( .A(n6065), .B(n6064), .Z(n6069) );
  NANDN U7944 ( .A(n6068), .B(n6069), .Z(n6071) );
  XOR U7945 ( .A(n6067), .B(n6066), .Z(n6371) );
  NANDN U7946 ( .A(n6371), .B(n6372), .Z(n6070) );
  NAND U7947 ( .A(n6071), .B(n6070), .Z(n10202) );
  XNOR U7948 ( .A(n10204), .B(n10205), .Z(n10210) );
  AND U7949 ( .A(a[53]), .B(b[47]), .Z(n10208) );
  AND U7950 ( .A(a[52]), .B(b[47]), .Z(n6369) );
  AND U7951 ( .A(a[46]), .B(b[47]), .Z(n6333) );
  AND U7952 ( .A(a[44]), .B(b[47]), .Z(n6323) );
  XNOR U7953 ( .A(n6073), .B(n6072), .Z(n6324) );
  NAND U7954 ( .A(n6323), .B(n6324), .Z(n6326) );
  AND U7955 ( .A(a[42]), .B(b[47]), .Z(n6313) );
  XOR U7956 ( .A(n6075), .B(n6074), .Z(n6314) );
  NAND U7957 ( .A(n6313), .B(n6314), .Z(n6316) );
  XOR U7958 ( .A(n6077), .B(n6076), .Z(n6304) );
  XOR U7959 ( .A(n6079), .B(n6078), .Z(n6302) );
  XOR U7960 ( .A(n6081), .B(n6080), .Z(n6297) );
  AND U7961 ( .A(a[38]), .B(b[47]), .Z(n6298) );
  NANDN U7962 ( .A(n6297), .B(n6298), .Z(n6300) );
  XOR U7963 ( .A(n6083), .B(n6082), .Z(n6084) );
  AND U7964 ( .A(a[36]), .B(b[47]), .Z(n6085) );
  NANDN U7965 ( .A(n6084), .B(n6085), .Z(n6290) );
  XOR U7966 ( .A(n6085), .B(n6084), .Z(n6383) );
  XOR U7967 ( .A(n6087), .B(n6086), .Z(n6280) );
  NAND U7968 ( .A(a[32]), .B(b[47]), .Z(n6269) );
  XNOR U7969 ( .A(n6089), .B(n6088), .Z(n6270) );
  NANDN U7970 ( .A(n6269), .B(n6270), .Z(n6272) );
  XOR U7971 ( .A(n6091), .B(n6090), .Z(n6266) );
  XOR U7972 ( .A(n6093), .B(n6092), .Z(n6262) );
  NAND U7973 ( .A(a[29]), .B(b[47]), .Z(n6257) );
  XNOR U7974 ( .A(n6095), .B(n6094), .Z(n6258) );
  NANDN U7975 ( .A(n6257), .B(n6258), .Z(n6260) );
  XOR U7976 ( .A(n6097), .B(n6096), .Z(n6254) );
  NAND U7977 ( .A(a[27]), .B(b[47]), .Z(n6249) );
  XNOR U7978 ( .A(n6099), .B(n6098), .Z(n6250) );
  NANDN U7979 ( .A(n6249), .B(n6250), .Z(n6252) );
  XOR U7980 ( .A(n6101), .B(n6100), .Z(n6239) );
  XOR U7981 ( .A(n6103), .B(n6102), .Z(n6236) );
  NAND U7982 ( .A(a[22]), .B(b[47]), .Z(n6225) );
  XNOR U7983 ( .A(n6105), .B(n6104), .Z(n6226) );
  NANDN U7984 ( .A(n6225), .B(n6226), .Z(n6228) );
  AND U7985 ( .A(a[21]), .B(b[47]), .Z(n6109) );
  XNOR U7986 ( .A(n6107), .B(n6106), .Z(n6108) );
  NANDN U7987 ( .A(n6109), .B(n6108), .Z(n6224) );
  XOR U7988 ( .A(n6109), .B(n6108), .Z(n6409) );
  XOR U7989 ( .A(n6111), .B(n6110), .Z(n6220) );
  XOR U7990 ( .A(n6113), .B(n6112), .Z(n6209) );
  AND U7991 ( .A(a[18]), .B(b[47]), .Z(n6210) );
  NANDN U7992 ( .A(n6209), .B(n6210), .Z(n6212) );
  NAND U7993 ( .A(a[16]), .B(b[47]), .Z(n6197) );
  AND U7994 ( .A(a[15]), .B(b[47]), .Z(n6193) );
  XNOR U7995 ( .A(n6115), .B(n6114), .Z(n6194) );
  NANDN U7996 ( .A(n6193), .B(n6194), .Z(n6196) );
  XOR U7997 ( .A(n6117), .B(n6116), .Z(n6189) );
  NAND U7998 ( .A(a[14]), .B(b[47]), .Z(n6190) );
  NANDN U7999 ( .A(n6189), .B(n6190), .Z(n6192) );
  XOR U8000 ( .A(n6119), .B(n6118), .Z(n6179) );
  AND U8001 ( .A(a[11]), .B(b[47]), .Z(n6175) );
  XOR U8002 ( .A(n6121), .B(n6120), .Z(n6163) );
  NAND U8003 ( .A(a[7]), .B(b[47]), .Z(n6153) );
  XOR U8004 ( .A(n6123), .B(n6122), .Z(n6154) );
  NANDN U8005 ( .A(n6153), .B(n6154), .Z(n6156) );
  XOR U8006 ( .A(n6125), .B(n6124), .Z(n6149) );
  NAND U8007 ( .A(a[0]), .B(b[47]), .Z(n6733) );
  AND U8008 ( .A(a[1]), .B(b[48]), .Z(n6128) );
  NANDN U8009 ( .A(n6733), .B(n6128), .Z(n6427) );
  NANDN U8010 ( .A(n6427), .B(n6126), .Z(n6130) );
  AND U8011 ( .A(a[2]), .B(b[47]), .Z(n6433) );
  NANDN U8012 ( .A(n6432), .B(n6433), .Z(n6129) );
  AND U8013 ( .A(n6130), .B(n6129), .Z(n6133) );
  AND U8014 ( .A(a[3]), .B(b[47]), .Z(n6134) );
  NANDN U8015 ( .A(n6133), .B(n6134), .Z(n6136) );
  XOR U8016 ( .A(n6132), .B(n6131), .Z(n6438) );
  NANDN U8017 ( .A(n6438), .B(n6439), .Z(n6135) );
  AND U8018 ( .A(n6136), .B(n6135), .Z(n6139) );
  NANDN U8019 ( .A(n6139), .B(n6140), .Z(n6142) );
  AND U8020 ( .A(a[4]), .B(b[47]), .Z(n6445) );
  NAND U8021 ( .A(n6445), .B(n6444), .Z(n6141) );
  AND U8022 ( .A(n6142), .B(n6141), .Z(n6143) );
  AND U8023 ( .A(a[5]), .B(b[47]), .Z(n6144) );
  NANDN U8024 ( .A(n6143), .B(n6144), .Z(n6148) );
  NAND U8025 ( .A(n6451), .B(n6450), .Z(n6147) );
  NAND U8026 ( .A(n6148), .B(n6147), .Z(n6150) );
  NANDN U8027 ( .A(n6149), .B(n6150), .Z(n6152) );
  NAND U8028 ( .A(a[6]), .B(b[47]), .Z(n6425) );
  NANDN U8029 ( .A(n6425), .B(n6426), .Z(n6151) );
  AND U8030 ( .A(n6152), .B(n6151), .Z(n6462) );
  NANDN U8031 ( .A(n6462), .B(n6463), .Z(n6155) );
  AND U8032 ( .A(n6156), .B(n6155), .Z(n6157) );
  AND U8033 ( .A(a[8]), .B(b[47]), .Z(n6158) );
  NANDN U8034 ( .A(n6157), .B(n6158), .Z(n6162) );
  NAND U8035 ( .A(n6424), .B(n6423), .Z(n6161) );
  AND U8036 ( .A(n6162), .B(n6161), .Z(n6164) );
  NANDN U8037 ( .A(n6163), .B(n6164), .Z(n6166) );
  AND U8038 ( .A(a[9]), .B(b[47]), .Z(n6470) );
  NANDN U8039 ( .A(n6470), .B(n6471), .Z(n6165) );
  AND U8040 ( .A(n6166), .B(n6165), .Z(n6170) );
  NAND U8041 ( .A(n6170), .B(n6169), .Z(n6172) );
  XOR U8042 ( .A(n6170), .B(n6169), .Z(n6479) );
  AND U8043 ( .A(a[10]), .B(b[47]), .Z(n6478) );
  NAND U8044 ( .A(n6479), .B(n6478), .Z(n6171) );
  AND U8045 ( .A(n6172), .B(n6171), .Z(n6176) );
  NANDN U8046 ( .A(n6175), .B(n6176), .Z(n6178) );
  XOR U8047 ( .A(n6174), .B(n6173), .Z(n6482) );
  NANDN U8048 ( .A(n6482), .B(n6483), .Z(n6177) );
  AND U8049 ( .A(n6178), .B(n6177), .Z(n6180) );
  NANDN U8050 ( .A(n6179), .B(n6180), .Z(n6182) );
  AND U8051 ( .A(a[12]), .B(b[47]), .Z(n6489) );
  NAND U8052 ( .A(n6489), .B(n6488), .Z(n6181) );
  AND U8053 ( .A(n6182), .B(n6181), .Z(n6185) );
  XOR U8054 ( .A(n6184), .B(n6183), .Z(n6186) );
  NANDN U8055 ( .A(n6185), .B(n6186), .Z(n6188) );
  NAND U8056 ( .A(a[13]), .B(b[47]), .Z(n6421) );
  NANDN U8057 ( .A(n6421), .B(n6422), .Z(n6187) );
  NAND U8058 ( .A(n6188), .B(n6187), .Z(n6419) );
  NANDN U8059 ( .A(n6419), .B(n6420), .Z(n6191) );
  AND U8060 ( .A(n6192), .B(n6191), .Z(n6504) );
  NANDN U8061 ( .A(n6504), .B(n6505), .Z(n6195) );
  AND U8062 ( .A(n6196), .B(n6195), .Z(n6198) );
  NANDN U8063 ( .A(n6197), .B(n6198), .Z(n6202) );
  NAND U8064 ( .A(n6418), .B(n6417), .Z(n6201) );
  AND U8065 ( .A(n6202), .B(n6201), .Z(n6205) );
  XOR U8066 ( .A(n6204), .B(n6203), .Z(n6206) );
  NANDN U8067 ( .A(n6205), .B(n6206), .Z(n6208) );
  NAND U8068 ( .A(a[17]), .B(b[47]), .Z(n6512) );
  NANDN U8069 ( .A(n6512), .B(n6513), .Z(n6207) );
  AND U8070 ( .A(n6208), .B(n6207), .Z(n6519) );
  XNOR U8071 ( .A(n6210), .B(n6209), .Z(n6518) );
  NANDN U8072 ( .A(n6519), .B(n6518), .Z(n6211) );
  AND U8073 ( .A(n6212), .B(n6211), .Z(n6216) );
  XNOR U8074 ( .A(n6214), .B(n6213), .Z(n6215) );
  NANDN U8075 ( .A(n6216), .B(n6215), .Z(n6218) );
  NAND U8076 ( .A(a[19]), .B(b[47]), .Z(n6415) );
  XNOR U8077 ( .A(n6216), .B(n6215), .Z(n6416) );
  NANDN U8078 ( .A(n6415), .B(n6416), .Z(n6217) );
  AND U8079 ( .A(n6218), .B(n6217), .Z(n6219) );
  NANDN U8080 ( .A(n6220), .B(n6219), .Z(n6222) );
  XOR U8081 ( .A(n6220), .B(n6219), .Z(n6413) );
  AND U8082 ( .A(a[20]), .B(b[47]), .Z(n6414) );
  OR U8083 ( .A(n6413), .B(n6414), .Z(n6221) );
  AND U8084 ( .A(n6222), .B(n6221), .Z(n6410) );
  OR U8085 ( .A(n6409), .B(n6410), .Z(n6223) );
  NAND U8086 ( .A(n6224), .B(n6223), .Z(n6534) );
  XNOR U8087 ( .A(n6226), .B(n6225), .Z(n6535) );
  NANDN U8088 ( .A(n6534), .B(n6535), .Z(n6227) );
  AND U8089 ( .A(n6228), .B(n6227), .Z(n6232) );
  XNOR U8090 ( .A(n6230), .B(n6229), .Z(n6231) );
  NANDN U8091 ( .A(n6232), .B(n6231), .Z(n6234) );
  NAND U8092 ( .A(a[23]), .B(b[47]), .Z(n6542) );
  XNOR U8093 ( .A(n6232), .B(n6231), .Z(n6543) );
  NANDN U8094 ( .A(n6542), .B(n6543), .Z(n6233) );
  AND U8095 ( .A(n6234), .B(n6233), .Z(n6235) );
  NANDN U8096 ( .A(n6236), .B(n6235), .Z(n6238) );
  XOR U8097 ( .A(n6236), .B(n6235), .Z(n6407) );
  AND U8098 ( .A(a[24]), .B(b[47]), .Z(n6408) );
  OR U8099 ( .A(n6407), .B(n6408), .Z(n6237) );
  AND U8100 ( .A(n6238), .B(n6237), .Z(n6240) );
  NANDN U8101 ( .A(n6239), .B(n6240), .Z(n6242) );
  NAND U8102 ( .A(a[25]), .B(b[47]), .Z(n6405) );
  XNOR U8103 ( .A(n6240), .B(n6239), .Z(n6406) );
  NANDN U8104 ( .A(n6405), .B(n6406), .Z(n6241) );
  AND U8105 ( .A(n6242), .B(n6241), .Z(n6246) );
  XNOR U8106 ( .A(n6244), .B(n6243), .Z(n6245) );
  NANDN U8107 ( .A(n6246), .B(n6245), .Z(n6248) );
  NAND U8108 ( .A(a[26]), .B(b[47]), .Z(n6401) );
  XNOR U8109 ( .A(n6246), .B(n6245), .Z(n6402) );
  NANDN U8110 ( .A(n6401), .B(n6402), .Z(n6247) );
  AND U8111 ( .A(n6248), .B(n6247), .Z(n6557) );
  XNOR U8112 ( .A(n6250), .B(n6249), .Z(n6556) );
  NANDN U8113 ( .A(n6557), .B(n6556), .Z(n6251) );
  NAND U8114 ( .A(n6252), .B(n6251), .Z(n6253) );
  NANDN U8115 ( .A(n6254), .B(n6253), .Z(n6256) );
  NAND U8116 ( .A(a[28]), .B(b[47]), .Z(n6399) );
  XNOR U8117 ( .A(n6254), .B(n6253), .Z(n6400) );
  NANDN U8118 ( .A(n6399), .B(n6400), .Z(n6255) );
  AND U8119 ( .A(n6256), .B(n6255), .Z(n6567) );
  XNOR U8120 ( .A(n6258), .B(n6257), .Z(n6566) );
  NANDN U8121 ( .A(n6567), .B(n6566), .Z(n6259) );
  AND U8122 ( .A(n6260), .B(n6259), .Z(n6261) );
  NANDN U8123 ( .A(n6262), .B(n6261), .Z(n6264) );
  XOR U8124 ( .A(n6262), .B(n6261), .Z(n6395) );
  AND U8125 ( .A(a[30]), .B(b[47]), .Z(n6396) );
  OR U8126 ( .A(n6395), .B(n6396), .Z(n6263) );
  AND U8127 ( .A(n6264), .B(n6263), .Z(n6265) );
  NANDN U8128 ( .A(n6266), .B(n6265), .Z(n6268) );
  NAND U8129 ( .A(a[31]), .B(b[47]), .Z(n6393) );
  XNOR U8130 ( .A(n6266), .B(n6265), .Z(n6394) );
  NANDN U8131 ( .A(n6393), .B(n6394), .Z(n6267) );
  AND U8132 ( .A(n6268), .B(n6267), .Z(n6390) );
  XNOR U8133 ( .A(n6270), .B(n6269), .Z(n6389) );
  NANDN U8134 ( .A(n6390), .B(n6389), .Z(n6271) );
  AND U8135 ( .A(n6272), .B(n6271), .Z(n6276) );
  AND U8136 ( .A(a[33]), .B(b[47]), .Z(n6275) );
  NANDN U8137 ( .A(n6276), .B(n6275), .Z(n6278) );
  XOR U8138 ( .A(n6274), .B(n6273), .Z(n6580) );
  XNOR U8139 ( .A(n6276), .B(n6275), .Z(n6581) );
  NANDN U8140 ( .A(n6580), .B(n6581), .Z(n6277) );
  AND U8141 ( .A(n6278), .B(n6277), .Z(n6279) );
  NANDN U8142 ( .A(n6280), .B(n6279), .Z(n6282) );
  XOR U8143 ( .A(n6280), .B(n6279), .Z(n6586) );
  AND U8144 ( .A(a[34]), .B(b[47]), .Z(n6587) );
  OR U8145 ( .A(n6586), .B(n6587), .Z(n6281) );
  NAND U8146 ( .A(n6282), .B(n6281), .Z(n6285) );
  XNOR U8147 ( .A(n6284), .B(n6283), .Z(n6286) );
  NANDN U8148 ( .A(n6285), .B(n6286), .Z(n6288) );
  XNOR U8149 ( .A(n6286), .B(n6285), .Z(n6388) );
  AND U8150 ( .A(a[35]), .B(b[47]), .Z(n6387) );
  NAND U8151 ( .A(n6388), .B(n6387), .Z(n6287) );
  AND U8152 ( .A(n6288), .B(n6287), .Z(n6384) );
  OR U8153 ( .A(n6383), .B(n6384), .Z(n6289) );
  AND U8154 ( .A(n6290), .B(n6289), .Z(n6294) );
  XNOR U8155 ( .A(n6292), .B(n6291), .Z(n6293) );
  NANDN U8156 ( .A(n6294), .B(n6293), .Z(n6296) );
  NAND U8157 ( .A(a[37]), .B(b[47]), .Z(n6598) );
  XNOR U8158 ( .A(n6294), .B(n6293), .Z(n6599) );
  NANDN U8159 ( .A(n6598), .B(n6599), .Z(n6295) );
  AND U8160 ( .A(n6296), .B(n6295), .Z(n6605) );
  XNOR U8161 ( .A(n6298), .B(n6297), .Z(n6604) );
  NANDN U8162 ( .A(n6605), .B(n6604), .Z(n6299) );
  AND U8163 ( .A(n6300), .B(n6299), .Z(n6301) );
  AND U8164 ( .A(a[39]), .B(b[47]), .Z(n6382) );
  XOR U8165 ( .A(n6302), .B(n6301), .Z(n6381) );
  NAND U8166 ( .A(n6304), .B(n6303), .Z(n6306) );
  AND U8167 ( .A(a[40]), .B(b[47]), .Z(n6615) );
  XOR U8168 ( .A(n6304), .B(n6303), .Z(n6614) );
  NANDN U8169 ( .A(n6615), .B(n6614), .Z(n6305) );
  AND U8170 ( .A(n6306), .B(n6305), .Z(n6310) );
  XNOR U8171 ( .A(n6308), .B(n6307), .Z(n6309) );
  NAND U8172 ( .A(n6310), .B(n6309), .Z(n6312) );
  XOR U8173 ( .A(n6310), .B(n6309), .Z(n6380) );
  AND U8174 ( .A(a[41]), .B(b[47]), .Z(n6379) );
  NAND U8175 ( .A(n6380), .B(n6379), .Z(n6311) );
  AND U8176 ( .A(n6312), .B(n6311), .Z(n6378) );
  XOR U8177 ( .A(n6314), .B(n6313), .Z(n6377) );
  NANDN U8178 ( .A(n6378), .B(n6377), .Z(n6315) );
  AND U8179 ( .A(n6316), .B(n6315), .Z(n6318) );
  AND U8180 ( .A(a[43]), .B(b[47]), .Z(n6317) );
  NANDN U8181 ( .A(n6318), .B(n6317), .Z(n6322) );
  XNOR U8182 ( .A(n6318), .B(n6317), .Z(n6628) );
  XOR U8183 ( .A(n6320), .B(n6319), .Z(n6629) );
  NAND U8184 ( .A(n6628), .B(n6629), .Z(n6321) );
  AND U8185 ( .A(n6322), .B(n6321), .Z(n6635) );
  XOR U8186 ( .A(n6324), .B(n6323), .Z(n6634) );
  NANDN U8187 ( .A(n6635), .B(n6634), .Z(n6325) );
  AND U8188 ( .A(n6326), .B(n6325), .Z(n6327) );
  AND U8189 ( .A(a[45]), .B(b[47]), .Z(n6328) );
  NANDN U8190 ( .A(n6327), .B(n6328), .Z(n6332) );
  NAND U8191 ( .A(n6376), .B(n6375), .Z(n6331) );
  AND U8192 ( .A(n6332), .B(n6331), .Z(n6334) );
  NANDN U8193 ( .A(n6333), .B(n6334), .Z(n6338) );
  NAND U8194 ( .A(n6645), .B(n6644), .Z(n6337) );
  NAND U8195 ( .A(n6338), .B(n6337), .Z(n6339) );
  AND U8196 ( .A(a[47]), .B(b[47]), .Z(n6340) );
  NANDN U8197 ( .A(n6339), .B(n6340), .Z(n6344) );
  XNOR U8198 ( .A(n6342), .B(n6341), .Z(n6653) );
  NAND U8199 ( .A(n6652), .B(n6653), .Z(n6343) );
  AND U8200 ( .A(n6344), .B(n6343), .Z(n6345) );
  AND U8201 ( .A(a[48]), .B(b[47]), .Z(n6346) );
  NANDN U8202 ( .A(n6345), .B(n6346), .Z(n6350) );
  XNOR U8203 ( .A(n6348), .B(n6347), .Z(n6659) );
  NAND U8204 ( .A(n6658), .B(n6659), .Z(n6349) );
  AND U8205 ( .A(n6350), .B(n6349), .Z(n6351) );
  AND U8206 ( .A(a[49]), .B(b[47]), .Z(n6352) );
  NANDN U8207 ( .A(n6351), .B(n6352), .Z(n6356) );
  NAND U8208 ( .A(n6662), .B(n6663), .Z(n6355) );
  AND U8209 ( .A(n6356), .B(n6355), .Z(n6357) );
  AND U8210 ( .A(a[50]), .B(b[47]), .Z(n6358) );
  NANDN U8211 ( .A(n6357), .B(n6358), .Z(n6362) );
  XNOR U8212 ( .A(n6360), .B(n6359), .Z(n6671) );
  NAND U8213 ( .A(n6670), .B(n6671), .Z(n6361) );
  AND U8214 ( .A(n6362), .B(n6361), .Z(n6363) );
  AND U8215 ( .A(a[51]), .B(b[47]), .Z(n6364) );
  NANDN U8216 ( .A(n6363), .B(n6364), .Z(n6368) );
  NAND U8217 ( .A(n6675), .B(n6674), .Z(n6367) );
  AND U8218 ( .A(n6368), .B(n6367), .Z(n6370) );
  NANDN U8219 ( .A(n6369), .B(n6370), .Z(n6374) );
  NAND U8220 ( .A(n6681), .B(n6680), .Z(n6373) );
  NAND U8221 ( .A(n6374), .B(n6373), .Z(n10209) );
  XNOR U8222 ( .A(n10210), .B(n10211), .Z(n10114) );
  AND U8223 ( .A(a[54]), .B(b[46]), .Z(n10113) );
  AND U8224 ( .A(a[52]), .B(b[46]), .Z(n6676) );
  AND U8225 ( .A(a[51]), .B(b[46]), .Z(n6668) );
  AND U8226 ( .A(a[49]), .B(b[46]), .Z(n6656) );
  AND U8227 ( .A(a[48]), .B(b[46]), .Z(n6650) );
  NAND U8228 ( .A(a[47]), .B(b[46]), .Z(n6646) );
  XOR U8229 ( .A(n6376), .B(n6375), .Z(n6640) );
  XOR U8230 ( .A(n6378), .B(n6377), .Z(n6625) );
  XOR U8231 ( .A(n6380), .B(n6379), .Z(n6621) );
  XOR U8232 ( .A(n6382), .B(n6381), .Z(n6610) );
  NAND U8233 ( .A(a[38]), .B(b[46]), .Z(n6600) );
  AND U8234 ( .A(a[37]), .B(b[46]), .Z(n6386) );
  XNOR U8235 ( .A(n6384), .B(n6383), .Z(n6385) );
  NANDN U8236 ( .A(n6386), .B(n6385), .Z(n6597) );
  XOR U8237 ( .A(n6386), .B(n6385), .Z(n6911) );
  XOR U8238 ( .A(n6388), .B(n6387), .Z(n6593) );
  NAND U8239 ( .A(a[33]), .B(b[46]), .Z(n6391) );
  XNOR U8240 ( .A(n6390), .B(n6389), .Z(n6392) );
  NANDN U8241 ( .A(n6391), .B(n6392), .Z(n6579) );
  XOR U8242 ( .A(n6392), .B(n6391), .Z(n6702) );
  XOR U8243 ( .A(n6394), .B(n6393), .Z(n6574) );
  AND U8244 ( .A(a[32]), .B(b[46]), .Z(n6575) );
  NANDN U8245 ( .A(n6574), .B(n6575), .Z(n6577) );
  XOR U8246 ( .A(n6396), .B(n6395), .Z(n6398) );
  AND U8247 ( .A(a[31]), .B(b[46]), .Z(n6397) );
  NANDN U8248 ( .A(n6398), .B(n6397), .Z(n6573) );
  XOR U8249 ( .A(n6398), .B(n6397), .Z(n6887) );
  XOR U8250 ( .A(n6400), .B(n6399), .Z(n6562) );
  AND U8251 ( .A(a[29]), .B(b[46]), .Z(n6563) );
  NANDN U8252 ( .A(n6562), .B(n6563), .Z(n6565) );
  NAND U8253 ( .A(a[27]), .B(b[46]), .Z(n6403) );
  XNOR U8254 ( .A(n6402), .B(n6401), .Z(n6404) );
  NANDN U8255 ( .A(n6403), .B(n6404), .Z(n6555) );
  XOR U8256 ( .A(n6404), .B(n6403), .Z(n6714) );
  XOR U8257 ( .A(n6406), .B(n6405), .Z(n6550) );
  AND U8258 ( .A(a[26]), .B(b[46]), .Z(n6551) );
  NANDN U8259 ( .A(n6550), .B(n6551), .Z(n6553) );
  XOR U8260 ( .A(n6408), .B(n6407), .Z(n6547) );
  AND U8261 ( .A(a[25]), .B(b[46]), .Z(n6546) );
  NANDN U8262 ( .A(n6547), .B(n6546), .Z(n6549) );
  XOR U8263 ( .A(n6410), .B(n6409), .Z(n6412) );
  AND U8264 ( .A(a[22]), .B(b[46]), .Z(n6411) );
  NANDN U8265 ( .A(n6412), .B(n6411), .Z(n6533) );
  XOR U8266 ( .A(n6412), .B(n6411), .Z(n6845) );
  XOR U8267 ( .A(n6414), .B(n6413), .Z(n6529) );
  AND U8268 ( .A(a[21]), .B(b[46]), .Z(n6528) );
  NANDN U8269 ( .A(n6529), .B(n6528), .Z(n6531) );
  XOR U8270 ( .A(n6416), .B(n6415), .Z(n6524) );
  AND U8271 ( .A(a[20]), .B(b[46]), .Z(n6525) );
  NANDN U8272 ( .A(n6524), .B(n6525), .Z(n6527) );
  XOR U8273 ( .A(n6418), .B(n6417), .Z(n6508) );
  AND U8274 ( .A(a[16]), .B(b[46]), .Z(n6502) );
  AND U8275 ( .A(a[15]), .B(b[46]), .Z(n6498) );
  NANDN U8276 ( .A(n6498), .B(n6499), .Z(n6501) );
  NAND U8277 ( .A(a[14]), .B(b[46]), .Z(n6494) );
  NANDN U8278 ( .A(n6494), .B(n6495), .Z(n6497) );
  AND U8279 ( .A(a[11]), .B(b[46]), .Z(n6476) );
  XOR U8280 ( .A(n6424), .B(n6423), .Z(n6466) );
  NAND U8281 ( .A(a[7]), .B(b[46]), .Z(n6456) );
  NANDN U8282 ( .A(n6456), .B(n6457), .Z(n6459) );
  NAND U8283 ( .A(a[0]), .B(b[46]), .Z(n7064) );
  AND U8284 ( .A(a[1]), .B(b[47]), .Z(n6429) );
  NANDN U8285 ( .A(n7064), .B(n6429), .Z(n6732) );
  NANDN U8286 ( .A(n6732), .B(n6427), .Z(n6431) );
  AND U8287 ( .A(a[2]), .B(b[46]), .Z(n6738) );
  NANDN U8288 ( .A(n6737), .B(n6738), .Z(n6430) );
  AND U8289 ( .A(n6431), .B(n6430), .Z(n6434) );
  AND U8290 ( .A(a[3]), .B(b[46]), .Z(n6435) );
  NANDN U8291 ( .A(n6434), .B(n6435), .Z(n6437) );
  XOR U8292 ( .A(n6433), .B(n6432), .Z(n6743) );
  NANDN U8293 ( .A(n6743), .B(n6744), .Z(n6436) );
  AND U8294 ( .A(n6437), .B(n6436), .Z(n6440) );
  NANDN U8295 ( .A(n6440), .B(n6441), .Z(n6443) );
  AND U8296 ( .A(a[4]), .B(b[46]), .Z(n6731) );
  NAND U8297 ( .A(n6731), .B(n6730), .Z(n6442) );
  AND U8298 ( .A(n6443), .B(n6442), .Z(n6446) );
  AND U8299 ( .A(a[5]), .B(b[46]), .Z(n6447) );
  NANDN U8300 ( .A(n6446), .B(n6447), .Z(n6449) );
  XOR U8301 ( .A(n6445), .B(n6444), .Z(n6754) );
  NAND U8302 ( .A(n6754), .B(n6753), .Z(n6448) );
  AND U8303 ( .A(n6449), .B(n6448), .Z(n6452) );
  XOR U8304 ( .A(n6451), .B(n6450), .Z(n6453) );
  NANDN U8305 ( .A(n6452), .B(n6453), .Z(n6455) );
  NAND U8306 ( .A(a[6]), .B(b[46]), .Z(n6728) );
  NANDN U8307 ( .A(n6728), .B(n6729), .Z(n6454) );
  AND U8308 ( .A(n6455), .B(n6454), .Z(n6763) );
  NANDN U8309 ( .A(n6763), .B(n6764), .Z(n6458) );
  AND U8310 ( .A(n6459), .B(n6458), .Z(n6460) );
  AND U8311 ( .A(a[8]), .B(b[46]), .Z(n6461) );
  NANDN U8312 ( .A(n6460), .B(n6461), .Z(n6465) );
  NAND U8313 ( .A(n6727), .B(n6726), .Z(n6464) );
  AND U8314 ( .A(n6465), .B(n6464), .Z(n6467) );
  NANDN U8315 ( .A(n6466), .B(n6467), .Z(n6469) );
  AND U8316 ( .A(a[9]), .B(b[46]), .Z(n6773) );
  NANDN U8317 ( .A(n6773), .B(n6774), .Z(n6468) );
  AND U8318 ( .A(n6469), .B(n6468), .Z(n6472) );
  NAND U8319 ( .A(n6472), .B(n6473), .Z(n6475) );
  AND U8320 ( .A(a[10]), .B(b[46]), .Z(n6780) );
  XOR U8321 ( .A(n6473), .B(n6472), .Z(n6779) );
  NAND U8322 ( .A(n6780), .B(n6779), .Z(n6474) );
  AND U8323 ( .A(n6475), .B(n6474), .Z(n6477) );
  NANDN U8324 ( .A(n6476), .B(n6477), .Z(n6481) );
  XNOR U8325 ( .A(n6479), .B(n6478), .Z(n6724) );
  NAND U8326 ( .A(n6725), .B(n6724), .Z(n6480) );
  AND U8327 ( .A(n6481), .B(n6480), .Z(n6485) );
  NAND U8328 ( .A(n6485), .B(n6484), .Z(n6487) );
  AND U8329 ( .A(a[12]), .B(b[46]), .Z(n6790) );
  XOR U8330 ( .A(n6485), .B(n6484), .Z(n6789) );
  NAND U8331 ( .A(n6790), .B(n6789), .Z(n6486) );
  AND U8332 ( .A(n6487), .B(n6486), .Z(n6490) );
  XOR U8333 ( .A(n6489), .B(n6488), .Z(n6491) );
  NANDN U8334 ( .A(n6490), .B(n6491), .Z(n6493) );
  AND U8335 ( .A(a[13]), .B(b[46]), .Z(n6723) );
  NAND U8336 ( .A(n6723), .B(n6722), .Z(n6492) );
  AND U8337 ( .A(n6493), .B(n6492), .Z(n6720) );
  NANDN U8338 ( .A(n6720), .B(n6721), .Z(n6496) );
  AND U8339 ( .A(n6497), .B(n6496), .Z(n6806) );
  NAND U8340 ( .A(n6806), .B(n6805), .Z(n6500) );
  NAND U8341 ( .A(n6501), .B(n6500), .Z(n6503) );
  NANDN U8342 ( .A(n6502), .B(n6503), .Z(n6507) );
  NAND U8343 ( .A(n6810), .B(n6809), .Z(n6506) );
  NAND U8344 ( .A(n6507), .B(n6506), .Z(n6509) );
  NANDN U8345 ( .A(n6508), .B(n6509), .Z(n6511) );
  AND U8346 ( .A(a[17]), .B(b[46]), .Z(n6815) );
  NANDN U8347 ( .A(n6815), .B(n6816), .Z(n6510) );
  NAND U8348 ( .A(n6511), .B(n6510), .Z(n6514) );
  NANDN U8349 ( .A(n6514), .B(n6515), .Z(n6517) );
  AND U8350 ( .A(a[18]), .B(b[46]), .Z(n6824) );
  NAND U8351 ( .A(n6824), .B(n6823), .Z(n6516) );
  AND U8352 ( .A(n6517), .B(n6516), .Z(n6521) );
  XNOR U8353 ( .A(n6519), .B(n6518), .Z(n6520) );
  NANDN U8354 ( .A(n6521), .B(n6520), .Z(n6523) );
  NAND U8355 ( .A(a[19]), .B(b[46]), .Z(n6827) );
  XNOR U8356 ( .A(n6521), .B(n6520), .Z(n6828) );
  NANDN U8357 ( .A(n6827), .B(n6828), .Z(n6522) );
  AND U8358 ( .A(n6523), .B(n6522), .Z(n6719) );
  XNOR U8359 ( .A(n6525), .B(n6524), .Z(n6718) );
  NANDN U8360 ( .A(n6719), .B(n6718), .Z(n6526) );
  AND U8361 ( .A(n6527), .B(n6526), .Z(n6838) );
  XNOR U8362 ( .A(n6529), .B(n6528), .Z(n6837) );
  NANDN U8363 ( .A(n6838), .B(n6837), .Z(n6530) );
  AND U8364 ( .A(n6531), .B(n6530), .Z(n6846) );
  OR U8365 ( .A(n6845), .B(n6846), .Z(n6532) );
  AND U8366 ( .A(n6533), .B(n6532), .Z(n6537) );
  AND U8367 ( .A(a[23]), .B(b[46]), .Z(n6536) );
  NANDN U8368 ( .A(n6537), .B(n6536), .Z(n6539) );
  XOR U8369 ( .A(n6535), .B(n6534), .Z(n6849) );
  XNOR U8370 ( .A(n6537), .B(n6536), .Z(n6850) );
  NANDN U8371 ( .A(n6849), .B(n6850), .Z(n6538) );
  AND U8372 ( .A(n6539), .B(n6538), .Z(n6541) );
  AND U8373 ( .A(a[24]), .B(b[46]), .Z(n6540) );
  NANDN U8374 ( .A(n6541), .B(n6540), .Z(n6545) );
  XOR U8375 ( .A(n6541), .B(n6540), .Z(n6716) );
  XNOR U8376 ( .A(n6543), .B(n6542), .Z(n6717) );
  NANDN U8377 ( .A(n6716), .B(n6717), .Z(n6544) );
  AND U8378 ( .A(n6545), .B(n6544), .Z(n6860) );
  XNOR U8379 ( .A(n6547), .B(n6546), .Z(n6859) );
  NANDN U8380 ( .A(n6860), .B(n6859), .Z(n6548) );
  AND U8381 ( .A(n6549), .B(n6548), .Z(n6866) );
  XNOR U8382 ( .A(n6551), .B(n6550), .Z(n6865) );
  NANDN U8383 ( .A(n6866), .B(n6865), .Z(n6552) );
  AND U8384 ( .A(n6553), .B(n6552), .Z(n6715) );
  OR U8385 ( .A(n6714), .B(n6715), .Z(n6554) );
  AND U8386 ( .A(n6555), .B(n6554), .Z(n6559) );
  XNOR U8387 ( .A(n6557), .B(n6556), .Z(n6558) );
  NANDN U8388 ( .A(n6559), .B(n6558), .Z(n6561) );
  NAND U8389 ( .A(a[28]), .B(b[46]), .Z(n6710) );
  XNOR U8390 ( .A(n6559), .B(n6558), .Z(n6711) );
  NANDN U8391 ( .A(n6710), .B(n6711), .Z(n6560) );
  AND U8392 ( .A(n6561), .B(n6560), .Z(n6878) );
  XNOR U8393 ( .A(n6563), .B(n6562), .Z(n6877) );
  NANDN U8394 ( .A(n6878), .B(n6877), .Z(n6564) );
  AND U8395 ( .A(n6565), .B(n6564), .Z(n6569) );
  XNOR U8396 ( .A(n6567), .B(n6566), .Z(n6568) );
  NANDN U8397 ( .A(n6569), .B(n6568), .Z(n6571) );
  XNOR U8398 ( .A(n6569), .B(n6568), .Z(n6709) );
  AND U8399 ( .A(a[30]), .B(b[46]), .Z(n6708) );
  NAND U8400 ( .A(n6709), .B(n6708), .Z(n6570) );
  AND U8401 ( .A(n6571), .B(n6570), .Z(n6888) );
  OR U8402 ( .A(n6887), .B(n6888), .Z(n6572) );
  AND U8403 ( .A(n6573), .B(n6572), .Z(n6705) );
  XNOR U8404 ( .A(n6575), .B(n6574), .Z(n6704) );
  NANDN U8405 ( .A(n6705), .B(n6704), .Z(n6576) );
  AND U8406 ( .A(n6577), .B(n6576), .Z(n6703) );
  OR U8407 ( .A(n6702), .B(n6703), .Z(n6578) );
  AND U8408 ( .A(n6579), .B(n6578), .Z(n6583) );
  AND U8409 ( .A(a[34]), .B(b[46]), .Z(n6582) );
  NANDN U8410 ( .A(n6583), .B(n6582), .Z(n6585) );
  XOR U8411 ( .A(n6581), .B(n6580), .Z(n6700) );
  XNOR U8412 ( .A(n6583), .B(n6582), .Z(n6701) );
  NANDN U8413 ( .A(n6700), .B(n6701), .Z(n6584) );
  AND U8414 ( .A(n6585), .B(n6584), .Z(n6589) );
  AND U8415 ( .A(a[35]), .B(b[46]), .Z(n6588) );
  NANDN U8416 ( .A(n6589), .B(n6588), .Z(n6591) );
  XOR U8417 ( .A(n6587), .B(n6586), .Z(n6699) );
  XNOR U8418 ( .A(n6589), .B(n6588), .Z(n6698) );
  NANDN U8419 ( .A(n6699), .B(n6698), .Z(n6590) );
  AND U8420 ( .A(n6591), .B(n6590), .Z(n6592) );
  NANDN U8421 ( .A(n6593), .B(n6592), .Z(n6595) );
  XOR U8422 ( .A(n6593), .B(n6592), .Z(n6696) );
  AND U8423 ( .A(a[36]), .B(b[46]), .Z(n6697) );
  OR U8424 ( .A(n6696), .B(n6697), .Z(n6594) );
  AND U8425 ( .A(n6595), .B(n6594), .Z(n6912) );
  OR U8426 ( .A(n6911), .B(n6912), .Z(n6596) );
  AND U8427 ( .A(n6597), .B(n6596), .Z(n6601) );
  NANDN U8428 ( .A(n6600), .B(n6601), .Z(n6603) );
  XOR U8429 ( .A(n6599), .B(n6598), .Z(n6694) );
  XNOR U8430 ( .A(n6601), .B(n6600), .Z(n6695) );
  NANDN U8431 ( .A(n6694), .B(n6695), .Z(n6602) );
  AND U8432 ( .A(n6603), .B(n6602), .Z(n6607) );
  XNOR U8433 ( .A(n6605), .B(n6604), .Z(n6606) );
  NANDN U8434 ( .A(n6607), .B(n6606), .Z(n6609) );
  NAND U8435 ( .A(a[39]), .B(b[46]), .Z(n6921) );
  XNOR U8436 ( .A(n6607), .B(n6606), .Z(n6922) );
  NANDN U8437 ( .A(n6921), .B(n6922), .Z(n6608) );
  AND U8438 ( .A(n6609), .B(n6608), .Z(n6611) );
  NANDN U8439 ( .A(n6610), .B(n6611), .Z(n6613) );
  AND U8440 ( .A(a[40]), .B(b[46]), .Z(n6693) );
  XNOR U8441 ( .A(n6611), .B(n6610), .Z(n6692) );
  NANDN U8442 ( .A(n6693), .B(n6692), .Z(n6612) );
  AND U8443 ( .A(n6613), .B(n6612), .Z(n6617) );
  XNOR U8444 ( .A(n6615), .B(n6614), .Z(n6616) );
  NANDN U8445 ( .A(n6617), .B(n6616), .Z(n6619) );
  XOR U8446 ( .A(n6617), .B(n6616), .Z(n6690) );
  AND U8447 ( .A(a[41]), .B(b[46]), .Z(n6691) );
  OR U8448 ( .A(n6690), .B(n6691), .Z(n6618) );
  NAND U8449 ( .A(n6619), .B(n6618), .Z(n6620) );
  NANDN U8450 ( .A(n6621), .B(n6620), .Z(n6623) );
  AND U8451 ( .A(a[42]), .B(b[46]), .Z(n6689) );
  XNOR U8452 ( .A(n6621), .B(n6620), .Z(n6688) );
  NANDN U8453 ( .A(n6689), .B(n6688), .Z(n6622) );
  NAND U8454 ( .A(n6623), .B(n6622), .Z(n6624) );
  NAND U8455 ( .A(n6625), .B(n6624), .Z(n6627) );
  AND U8456 ( .A(a[43]), .B(b[46]), .Z(n6940) );
  XOR U8457 ( .A(n6625), .B(n6624), .Z(n6939) );
  NANDN U8458 ( .A(n6940), .B(n6939), .Z(n6626) );
  AND U8459 ( .A(n6627), .B(n6626), .Z(n6631) );
  XNOR U8460 ( .A(n6629), .B(n6628), .Z(n6630) );
  NANDN U8461 ( .A(n6631), .B(n6630), .Z(n6633) );
  AND U8462 ( .A(a[44]), .B(b[46]), .Z(n6946) );
  XNOR U8463 ( .A(n6631), .B(n6630), .Z(n6945) );
  NANDN U8464 ( .A(n6946), .B(n6945), .Z(n6632) );
  AND U8465 ( .A(n6633), .B(n6632), .Z(n6637) );
  XNOR U8466 ( .A(n6635), .B(n6634), .Z(n6636) );
  NAND U8467 ( .A(n6637), .B(n6636), .Z(n6639) );
  NAND U8468 ( .A(a[45]), .B(b[46]), .Z(n6951) );
  XOR U8469 ( .A(n6637), .B(n6636), .Z(n6952) );
  NANDN U8470 ( .A(n6951), .B(n6952), .Z(n6638) );
  AND U8471 ( .A(n6639), .B(n6638), .Z(n6641) );
  NANDN U8472 ( .A(n6640), .B(n6641), .Z(n6643) );
  AND U8473 ( .A(a[46]), .B(b[46]), .Z(n6959) );
  NANDN U8474 ( .A(n6959), .B(n6960), .Z(n6642) );
  AND U8475 ( .A(n6643), .B(n6642), .Z(n6647) );
  NANDN U8476 ( .A(n6646), .B(n6647), .Z(n6649) );
  XOR U8477 ( .A(n6645), .B(n6644), .Z(n6686) );
  NANDN U8478 ( .A(n6686), .B(n6687), .Z(n6648) );
  AND U8479 ( .A(n6649), .B(n6648), .Z(n6651) );
  NANDN U8480 ( .A(n6650), .B(n6651), .Z(n6655) );
  XNOR U8481 ( .A(n6653), .B(n6652), .Z(n6970) );
  NAND U8482 ( .A(n6969), .B(n6970), .Z(n6654) );
  NAND U8483 ( .A(n6655), .B(n6654), .Z(n6657) );
  NANDN U8484 ( .A(n6656), .B(n6657), .Z(n6661) );
  XNOR U8485 ( .A(n6659), .B(n6658), .Z(n6976) );
  NAND U8486 ( .A(n6975), .B(n6976), .Z(n6660) );
  NAND U8487 ( .A(n6661), .B(n6660), .Z(n6664) );
  AND U8488 ( .A(a[50]), .B(b[46]), .Z(n6665) );
  NANDN U8489 ( .A(n6664), .B(n6665), .Z(n6667) );
  XOR U8490 ( .A(n6663), .B(n6662), .Z(n6980) );
  NAND U8491 ( .A(n6980), .B(n6979), .Z(n6666) );
  AND U8492 ( .A(n6667), .B(n6666), .Z(n6669) );
  NANDN U8493 ( .A(n6668), .B(n6669), .Z(n6673) );
  XNOR U8494 ( .A(n6671), .B(n6670), .Z(n6988) );
  NAND U8495 ( .A(n6987), .B(n6988), .Z(n6672) );
  NAND U8496 ( .A(n6673), .B(n6672), .Z(n6677) );
  NANDN U8497 ( .A(n6676), .B(n6677), .Z(n6679) );
  XOR U8498 ( .A(n6675), .B(n6674), .Z(n6993) );
  NANDN U8499 ( .A(n6993), .B(n6994), .Z(n6678) );
  NAND U8500 ( .A(n6679), .B(n6678), .Z(n6682) );
  AND U8501 ( .A(a[53]), .B(b[46]), .Z(n6683) );
  NANDN U8502 ( .A(n6682), .B(n6683), .Z(n6685) );
  XOR U8503 ( .A(n6681), .B(n6680), .Z(n6997) );
  NANDN U8504 ( .A(n6997), .B(n6998), .Z(n6684) );
  AND U8505 ( .A(n6685), .B(n6684), .Z(n10112) );
  XNOR U8506 ( .A(n10114), .B(n10115), .Z(n10216) );
  AND U8507 ( .A(a[55]), .B(b[45]), .Z(n10214) );
  AND U8508 ( .A(a[51]), .B(b[45]), .Z(n6981) );
  AND U8509 ( .A(a[48]), .B(b[45]), .Z(n6964) );
  NAND U8510 ( .A(n6964), .B(n6963), .Z(n6966) );
  XOR U8511 ( .A(n6689), .B(n6688), .Z(n6936) );
  AND U8512 ( .A(a[43]), .B(b[45]), .Z(n6935) );
  NAND U8513 ( .A(n6936), .B(n6935), .Z(n6938) );
  XOR U8514 ( .A(n6691), .B(n6690), .Z(n6932) );
  XOR U8515 ( .A(n6693), .B(n6692), .Z(n6927) );
  NAND U8516 ( .A(a[39]), .B(b[45]), .Z(n6917) );
  XNOR U8517 ( .A(n6695), .B(n6694), .Z(n6918) );
  NANDN U8518 ( .A(n6917), .B(n6918), .Z(n6920) );
  XOR U8519 ( .A(n6697), .B(n6696), .Z(n6908) );
  AND U8520 ( .A(a[37]), .B(b[45]), .Z(n6907) );
  NANDN U8521 ( .A(n6908), .B(n6907), .Z(n6910) );
  NAND U8522 ( .A(a[36]), .B(b[45]), .Z(n6903) );
  XNOR U8523 ( .A(n6699), .B(n6698), .Z(n6904) );
  NANDN U8524 ( .A(n6903), .B(n6904), .Z(n6906) );
  XOR U8525 ( .A(n6701), .B(n6700), .Z(n6899) );
  XOR U8526 ( .A(n6703), .B(n6702), .Z(n6896) );
  XOR U8527 ( .A(n6705), .B(n6704), .Z(n6706) );
  AND U8528 ( .A(a[33]), .B(b[45]), .Z(n6707) );
  NANDN U8529 ( .A(n6706), .B(n6707), .Z(n6894) );
  XOR U8530 ( .A(n6707), .B(n6706), .Z(n7031) );
  XOR U8531 ( .A(n6709), .B(n6708), .Z(n6884) );
  XOR U8532 ( .A(n6711), .B(n6710), .Z(n6712) );
  AND U8533 ( .A(a[29]), .B(b[45]), .Z(n6713) );
  NANDN U8534 ( .A(n6712), .B(n6713), .Z(n6876) );
  XOR U8535 ( .A(n6713), .B(n6712), .Z(n7039) );
  XOR U8536 ( .A(n6715), .B(n6714), .Z(n6872) );
  NAND U8537 ( .A(a[25]), .B(b[45]), .Z(n6855) );
  XNOR U8538 ( .A(n6717), .B(n6716), .Z(n6856) );
  NANDN U8539 ( .A(n6855), .B(n6856), .Z(n6858) );
  AND U8540 ( .A(a[23]), .B(b[45]), .Z(n6844) );
  XOR U8541 ( .A(n6719), .B(n6718), .Z(n6833) );
  AND U8542 ( .A(a[21]), .B(b[45]), .Z(n6834) );
  NANDN U8543 ( .A(n6833), .B(n6834), .Z(n6836) );
  AND U8544 ( .A(a[16]), .B(b[45]), .Z(n6803) );
  NAND U8545 ( .A(a[15]), .B(b[45]), .Z(n6799) );
  NANDN U8546 ( .A(n6799), .B(n6800), .Z(n6802) );
  NAND U8547 ( .A(a[14]), .B(b[45]), .Z(n6795) );
  XOR U8548 ( .A(n6723), .B(n6722), .Z(n6796) );
  NANDN U8549 ( .A(n6795), .B(n6796), .Z(n6798) );
  XOR U8550 ( .A(n6725), .B(n6724), .Z(n6785) );
  AND U8551 ( .A(a[11]), .B(b[45]), .Z(n6781) );
  XOR U8552 ( .A(n6727), .B(n6726), .Z(n6769) );
  NAND U8553 ( .A(a[7]), .B(b[45]), .Z(n6759) );
  NANDN U8554 ( .A(n6759), .B(n6760), .Z(n6762) );
  XOR U8555 ( .A(n6731), .B(n6730), .Z(n6749) );
  NAND U8556 ( .A(a[0]), .B(b[45]), .Z(n7391) );
  AND U8557 ( .A(a[1]), .B(b[46]), .Z(n6734) );
  NANDN U8558 ( .A(n7391), .B(n6734), .Z(n7063) );
  NANDN U8559 ( .A(n7063), .B(n6732), .Z(n6736) );
  AND U8560 ( .A(a[2]), .B(b[45]), .Z(n7069) );
  NANDN U8561 ( .A(n7068), .B(n7069), .Z(n6735) );
  AND U8562 ( .A(n6736), .B(n6735), .Z(n6739) );
  AND U8563 ( .A(a[3]), .B(b[45]), .Z(n6740) );
  NANDN U8564 ( .A(n6739), .B(n6740), .Z(n6742) );
  XOR U8565 ( .A(n6738), .B(n6737), .Z(n7074) );
  NANDN U8566 ( .A(n7074), .B(n7075), .Z(n6741) );
  AND U8567 ( .A(n6742), .B(n6741), .Z(n6745) );
  NANDN U8568 ( .A(n6745), .B(n6746), .Z(n6748) );
  AND U8569 ( .A(a[4]), .B(b[45]), .Z(n7081) );
  NAND U8570 ( .A(n7081), .B(n7080), .Z(n6747) );
  AND U8571 ( .A(n6748), .B(n6747), .Z(n6750) );
  NANDN U8572 ( .A(n6749), .B(n6750), .Z(n6752) );
  NAND U8573 ( .A(a[5]), .B(b[45]), .Z(n7086) );
  NAND U8574 ( .A(n7087), .B(n7086), .Z(n6751) );
  AND U8575 ( .A(n6752), .B(n6751), .Z(n6756) );
  XOR U8576 ( .A(n6754), .B(n6753), .Z(n6755) );
  NAND U8577 ( .A(n6756), .B(n6755), .Z(n6758) );
  AND U8578 ( .A(a[6]), .B(b[45]), .Z(n7062) );
  XOR U8579 ( .A(n6756), .B(n6755), .Z(n7061) );
  NAND U8580 ( .A(n7062), .B(n7061), .Z(n6757) );
  AND U8581 ( .A(n6758), .B(n6757), .Z(n7057) );
  NANDN U8582 ( .A(n7057), .B(n7058), .Z(n6761) );
  AND U8583 ( .A(n6762), .B(n6761), .Z(n6765) );
  AND U8584 ( .A(a[8]), .B(b[45]), .Z(n6766) );
  NANDN U8585 ( .A(n6765), .B(n6766), .Z(n6768) );
  NAND U8586 ( .A(n7056), .B(n7055), .Z(n6767) );
  AND U8587 ( .A(n6768), .B(n6767), .Z(n6770) );
  NANDN U8588 ( .A(n6769), .B(n6770), .Z(n6772) );
  AND U8589 ( .A(a[9]), .B(b[45]), .Z(n7102) );
  NANDN U8590 ( .A(n7102), .B(n7103), .Z(n6771) );
  AND U8591 ( .A(n6772), .B(n6771), .Z(n6776) );
  NAND U8592 ( .A(n6776), .B(n6775), .Z(n6778) );
  XOR U8593 ( .A(n6776), .B(n6775), .Z(n7111) );
  AND U8594 ( .A(a[10]), .B(b[45]), .Z(n7110) );
  NAND U8595 ( .A(n7111), .B(n7110), .Z(n6777) );
  AND U8596 ( .A(n6778), .B(n6777), .Z(n6782) );
  NANDN U8597 ( .A(n6781), .B(n6782), .Z(n6784) );
  XOR U8598 ( .A(n6780), .B(n6779), .Z(n7114) );
  NANDN U8599 ( .A(n7114), .B(n7115), .Z(n6783) );
  AND U8600 ( .A(n6784), .B(n6783), .Z(n6786) );
  NANDN U8601 ( .A(n6785), .B(n6786), .Z(n6788) );
  AND U8602 ( .A(a[12]), .B(b[45]), .Z(n7121) );
  NAND U8603 ( .A(n7121), .B(n7120), .Z(n6787) );
  AND U8604 ( .A(n6788), .B(n6787), .Z(n6791) );
  XOR U8605 ( .A(n6790), .B(n6789), .Z(n6792) );
  NANDN U8606 ( .A(n6791), .B(n6792), .Z(n6794) );
  AND U8607 ( .A(a[13]), .B(b[45]), .Z(n7054) );
  NAND U8608 ( .A(n7054), .B(n7053), .Z(n6793) );
  AND U8609 ( .A(n6794), .B(n6793), .Z(n7051) );
  NANDN U8610 ( .A(n7051), .B(n7052), .Z(n6797) );
  AND U8611 ( .A(n6798), .B(n6797), .Z(n7134) );
  NANDN U8612 ( .A(n7134), .B(n7135), .Z(n6801) );
  AND U8613 ( .A(n6802), .B(n6801), .Z(n6804) );
  NANDN U8614 ( .A(n6803), .B(n6804), .Z(n6808) );
  XOR U8615 ( .A(n6806), .B(n6805), .Z(n7140) );
  NAND U8616 ( .A(n7141), .B(n7140), .Z(n6807) );
  AND U8617 ( .A(n6808), .B(n6807), .Z(n6811) );
  XOR U8618 ( .A(n6810), .B(n6809), .Z(n6812) );
  NANDN U8619 ( .A(n6811), .B(n6812), .Z(n6814) );
  AND U8620 ( .A(a[17]), .B(b[45]), .Z(n7146) );
  NANDN U8621 ( .A(n7146), .B(n7147), .Z(n6813) );
  AND U8622 ( .A(n6814), .B(n6813), .Z(n6817) );
  NAND U8623 ( .A(n6817), .B(n6818), .Z(n6820) );
  AND U8624 ( .A(a[18]), .B(b[45]), .Z(n7050) );
  XOR U8625 ( .A(n6818), .B(n6817), .Z(n7049) );
  NAND U8626 ( .A(n7050), .B(n7049), .Z(n6819) );
  AND U8627 ( .A(n6820), .B(n6819), .Z(n6821) );
  AND U8628 ( .A(a[19]), .B(b[45]), .Z(n6822) );
  NANDN U8629 ( .A(n6821), .B(n6822), .Z(n6826) );
  XOR U8630 ( .A(n6824), .B(n6823), .Z(n7158) );
  NAND U8631 ( .A(n7159), .B(n7158), .Z(n6825) );
  AND U8632 ( .A(n6826), .B(n6825), .Z(n6830) );
  XNOR U8633 ( .A(n6828), .B(n6827), .Z(n6829) );
  NANDN U8634 ( .A(n6830), .B(n6829), .Z(n6832) );
  NAND U8635 ( .A(a[20]), .B(b[45]), .Z(n7162) );
  XNOR U8636 ( .A(n6830), .B(n6829), .Z(n7163) );
  NANDN U8637 ( .A(n7162), .B(n7163), .Z(n6831) );
  AND U8638 ( .A(n6832), .B(n6831), .Z(n7169) );
  XNOR U8639 ( .A(n6834), .B(n6833), .Z(n7168) );
  NANDN U8640 ( .A(n7169), .B(n7168), .Z(n6835) );
  AND U8641 ( .A(n6836), .B(n6835), .Z(n6840) );
  XNOR U8642 ( .A(n6838), .B(n6837), .Z(n6839) );
  NANDN U8643 ( .A(n6840), .B(n6839), .Z(n6842) );
  NAND U8644 ( .A(a[22]), .B(b[45]), .Z(n7047) );
  XNOR U8645 ( .A(n6840), .B(n6839), .Z(n7048) );
  NANDN U8646 ( .A(n7047), .B(n7048), .Z(n6841) );
  AND U8647 ( .A(n6842), .B(n6841), .Z(n6843) );
  NANDN U8648 ( .A(n6844), .B(n6843), .Z(n6848) );
  XOR U8649 ( .A(n6844), .B(n6843), .Z(n7045) );
  XOR U8650 ( .A(n6846), .B(n6845), .Z(n7046) );
  OR U8651 ( .A(n7045), .B(n7046), .Z(n6847) );
  NAND U8652 ( .A(n6848), .B(n6847), .Z(n6851) );
  XNOR U8653 ( .A(n6850), .B(n6849), .Z(n6852) );
  NANDN U8654 ( .A(n6851), .B(n6852), .Z(n6854) );
  NAND U8655 ( .A(a[24]), .B(b[45]), .Z(n7182) );
  XNOR U8656 ( .A(n6852), .B(n6851), .Z(n7183) );
  NANDN U8657 ( .A(n7182), .B(n7183), .Z(n6853) );
  AND U8658 ( .A(n6854), .B(n6853), .Z(n7189) );
  XNOR U8659 ( .A(n6856), .B(n6855), .Z(n7188) );
  NANDN U8660 ( .A(n7189), .B(n7188), .Z(n6857) );
  AND U8661 ( .A(n6858), .B(n6857), .Z(n6862) );
  XNOR U8662 ( .A(n6860), .B(n6859), .Z(n6861) );
  NANDN U8663 ( .A(n6862), .B(n6861), .Z(n6864) );
  NAND U8664 ( .A(a[26]), .B(b[45]), .Z(n7043) );
  XNOR U8665 ( .A(n6862), .B(n6861), .Z(n7044) );
  NANDN U8666 ( .A(n7043), .B(n7044), .Z(n6863) );
  AND U8667 ( .A(n6864), .B(n6863), .Z(n6868) );
  XNOR U8668 ( .A(n6866), .B(n6865), .Z(n6867) );
  NANDN U8669 ( .A(n6868), .B(n6867), .Z(n6870) );
  NAND U8670 ( .A(a[27]), .B(b[45]), .Z(n7198) );
  XNOR U8671 ( .A(n6868), .B(n6867), .Z(n7199) );
  NANDN U8672 ( .A(n7198), .B(n7199), .Z(n6869) );
  AND U8673 ( .A(n6870), .B(n6869), .Z(n6871) );
  NANDN U8674 ( .A(n6872), .B(n6871), .Z(n6874) );
  XOR U8675 ( .A(n6872), .B(n6871), .Z(n7041) );
  AND U8676 ( .A(a[28]), .B(b[45]), .Z(n7042) );
  OR U8677 ( .A(n7041), .B(n7042), .Z(n6873) );
  AND U8678 ( .A(n6874), .B(n6873), .Z(n7040) );
  NANDN U8679 ( .A(n7039), .B(n7040), .Z(n6875) );
  AND U8680 ( .A(n6876), .B(n6875), .Z(n6880) );
  XNOR U8681 ( .A(n6878), .B(n6877), .Z(n6879) );
  NANDN U8682 ( .A(n6880), .B(n6879), .Z(n6882) );
  NAND U8683 ( .A(a[30]), .B(b[45]), .Z(n7037) );
  XNOR U8684 ( .A(n6880), .B(n6879), .Z(n7038) );
  NANDN U8685 ( .A(n7037), .B(n7038), .Z(n6881) );
  AND U8686 ( .A(n6882), .B(n6881), .Z(n6883) );
  NANDN U8687 ( .A(n6884), .B(n6883), .Z(n6886) );
  XOR U8688 ( .A(n6884), .B(n6883), .Z(n7035) );
  AND U8689 ( .A(a[31]), .B(b[45]), .Z(n7036) );
  OR U8690 ( .A(n7035), .B(n7036), .Z(n6885) );
  AND U8691 ( .A(n6886), .B(n6885), .Z(n6890) );
  XNOR U8692 ( .A(n6888), .B(n6887), .Z(n6889) );
  NANDN U8693 ( .A(n6890), .B(n6889), .Z(n6892) );
  XOR U8694 ( .A(n6890), .B(n6889), .Z(n7033) );
  AND U8695 ( .A(a[32]), .B(b[45]), .Z(n7034) );
  OR U8696 ( .A(n7033), .B(n7034), .Z(n6891) );
  AND U8697 ( .A(n6892), .B(n6891), .Z(n7032) );
  NANDN U8698 ( .A(n7031), .B(n7032), .Z(n6893) );
  AND U8699 ( .A(n6894), .B(n6893), .Z(n6895) );
  NANDN U8700 ( .A(n6896), .B(n6895), .Z(n6898) );
  XOR U8701 ( .A(n6896), .B(n6895), .Z(n7027) );
  AND U8702 ( .A(a[34]), .B(b[45]), .Z(n7028) );
  OR U8703 ( .A(n7027), .B(n7028), .Z(n6897) );
  AND U8704 ( .A(n6898), .B(n6897), .Z(n6900) );
  NANDN U8705 ( .A(n6899), .B(n6900), .Z(n6902) );
  NAND U8706 ( .A(a[35]), .B(b[45]), .Z(n7025) );
  XNOR U8707 ( .A(n6900), .B(n6899), .Z(n7026) );
  NANDN U8708 ( .A(n7025), .B(n7026), .Z(n6901) );
  AND U8709 ( .A(n6902), .B(n6901), .Z(n7235) );
  XNOR U8710 ( .A(n6904), .B(n6903), .Z(n7234) );
  NANDN U8711 ( .A(n7235), .B(n7234), .Z(n6905) );
  AND U8712 ( .A(n6906), .B(n6905), .Z(n7024) );
  XNOR U8713 ( .A(n6908), .B(n6907), .Z(n7023) );
  NANDN U8714 ( .A(n7024), .B(n7023), .Z(n6909) );
  AND U8715 ( .A(n6910), .B(n6909), .Z(n6914) );
  AND U8716 ( .A(a[38]), .B(b[45]), .Z(n6913) );
  NANDN U8717 ( .A(n6914), .B(n6913), .Z(n6916) );
  XOR U8718 ( .A(n6912), .B(n6911), .Z(n7020) );
  XNOR U8719 ( .A(n6914), .B(n6913), .Z(n7019) );
  NANDN U8720 ( .A(n7020), .B(n7019), .Z(n6915) );
  AND U8721 ( .A(n6916), .B(n6915), .Z(n7247) );
  XNOR U8722 ( .A(n6918), .B(n6917), .Z(n7246) );
  NANDN U8723 ( .A(n7247), .B(n7246), .Z(n6919) );
  AND U8724 ( .A(n6920), .B(n6919), .Z(n6924) );
  XNOR U8725 ( .A(n6922), .B(n6921), .Z(n6923) );
  NANDN U8726 ( .A(n6924), .B(n6923), .Z(n6926) );
  XNOR U8727 ( .A(n6924), .B(n6923), .Z(n7018) );
  AND U8728 ( .A(a[40]), .B(b[45]), .Z(n7017) );
  NAND U8729 ( .A(n7018), .B(n7017), .Z(n6925) );
  AND U8730 ( .A(n6926), .B(n6925), .Z(n6928) );
  NANDN U8731 ( .A(n6927), .B(n6928), .Z(n6930) );
  AND U8732 ( .A(a[41]), .B(b[45]), .Z(n7257) );
  XNOR U8733 ( .A(n6928), .B(n6927), .Z(n7256) );
  NANDN U8734 ( .A(n7257), .B(n7256), .Z(n6929) );
  AND U8735 ( .A(n6930), .B(n6929), .Z(n6931) );
  NANDN U8736 ( .A(n6932), .B(n6931), .Z(n6934) );
  XNOR U8737 ( .A(n6932), .B(n6931), .Z(n7014) );
  AND U8738 ( .A(a[42]), .B(b[45]), .Z(n7013) );
  NAND U8739 ( .A(n7014), .B(n7013), .Z(n6933) );
  AND U8740 ( .A(n6934), .B(n6933), .Z(n7265) );
  XOR U8741 ( .A(n6936), .B(n6935), .Z(n7264) );
  NANDN U8742 ( .A(n7265), .B(n7264), .Z(n6937) );
  AND U8743 ( .A(n6938), .B(n6937), .Z(n6942) );
  AND U8744 ( .A(a[44]), .B(b[45]), .Z(n6941) );
  NANDN U8745 ( .A(n6942), .B(n6941), .Z(n6944) );
  XOR U8746 ( .A(n6940), .B(n6939), .Z(n7271) );
  XNOR U8747 ( .A(n6942), .B(n6941), .Z(n7270) );
  NAND U8748 ( .A(n7271), .B(n7270), .Z(n6943) );
  AND U8749 ( .A(n6944), .B(n6943), .Z(n6948) );
  XNOR U8750 ( .A(n6946), .B(n6945), .Z(n6947) );
  NAND U8751 ( .A(n6948), .B(n6947), .Z(n6950) );
  AND U8752 ( .A(a[45]), .B(b[45]), .Z(n7012) );
  XOR U8753 ( .A(n6948), .B(n6947), .Z(n7011) );
  NANDN U8754 ( .A(n7012), .B(n7011), .Z(n6949) );
  AND U8755 ( .A(n6950), .B(n6949), .Z(n6954) );
  XNOR U8756 ( .A(n6952), .B(n6951), .Z(n6953) );
  NAND U8757 ( .A(n6954), .B(n6953), .Z(n6956) );
  NAND U8758 ( .A(a[46]), .B(b[45]), .Z(n7009) );
  XOR U8759 ( .A(n6954), .B(n6953), .Z(n7010) );
  NANDN U8760 ( .A(n7009), .B(n7010), .Z(n6955) );
  AND U8761 ( .A(n6956), .B(n6955), .Z(n6957) );
  AND U8762 ( .A(a[47]), .B(b[45]), .Z(n6958) );
  NANDN U8763 ( .A(n6957), .B(n6958), .Z(n6962) );
  NAND U8764 ( .A(n7007), .B(n7008), .Z(n6961) );
  AND U8765 ( .A(n6962), .B(n6961), .Z(n7005) );
  XOR U8766 ( .A(n6964), .B(n6963), .Z(n7006) );
  NANDN U8767 ( .A(n7005), .B(n7006), .Z(n6965) );
  AND U8768 ( .A(n6966), .B(n6965), .Z(n6967) );
  AND U8769 ( .A(a[49]), .B(b[45]), .Z(n6968) );
  NANDN U8770 ( .A(n6967), .B(n6968), .Z(n6972) );
  XNOR U8771 ( .A(n6970), .B(n6969), .Z(n7004) );
  NAND U8772 ( .A(n7003), .B(n7004), .Z(n6971) );
  AND U8773 ( .A(n6972), .B(n6971), .Z(n6973) );
  AND U8774 ( .A(a[50]), .B(b[45]), .Z(n6974) );
  NANDN U8775 ( .A(n6973), .B(n6974), .Z(n6978) );
  XNOR U8776 ( .A(n6976), .B(n6975), .Z(n7299) );
  NAND U8777 ( .A(n7298), .B(n7299), .Z(n6977) );
  AND U8778 ( .A(n6978), .B(n6977), .Z(n6982) );
  NANDN U8779 ( .A(n6981), .B(n6982), .Z(n6984) );
  XOR U8780 ( .A(n6980), .B(n6979), .Z(n7304) );
  NANDN U8781 ( .A(n7304), .B(n7305), .Z(n6983) );
  NAND U8782 ( .A(n6984), .B(n6983), .Z(n6985) );
  AND U8783 ( .A(a[52]), .B(b[45]), .Z(n6986) );
  NANDN U8784 ( .A(n6985), .B(n6986), .Z(n6990) );
  XNOR U8785 ( .A(n6988), .B(n6987), .Z(n7309) );
  NAND U8786 ( .A(n7308), .B(n7309), .Z(n6989) );
  AND U8787 ( .A(n6990), .B(n6989), .Z(n6991) );
  AND U8788 ( .A(a[53]), .B(b[45]), .Z(n6992) );
  NANDN U8789 ( .A(n6991), .B(n6992), .Z(n6996) );
  NAND U8790 ( .A(n7314), .B(n7315), .Z(n6995) );
  AND U8791 ( .A(n6996), .B(n6995), .Z(n6999) );
  AND U8792 ( .A(a[54]), .B(b[45]), .Z(n7000) );
  NANDN U8793 ( .A(n6999), .B(n7000), .Z(n7002) );
  NAND U8794 ( .A(n7321), .B(n7320), .Z(n7001) );
  AND U8795 ( .A(n7002), .B(n7001), .Z(n10215) );
  XOR U8796 ( .A(n10216), .B(n10217), .Z(n10223) );
  NAND U8797 ( .A(a[56]), .B(b[44]), .Z(n10221) );
  AND U8798 ( .A(a[54]), .B(b[44]), .Z(n7317) );
  NAND U8799 ( .A(a[53]), .B(b[44]), .Z(n7311) );
  AND U8800 ( .A(a[52]), .B(b[44]), .Z(n7302) );
  AND U8801 ( .A(a[51]), .B(b[44]), .Z(n7296) );
  NAND U8802 ( .A(a[50]), .B(b[44]), .Z(n7292) );
  XOR U8803 ( .A(n7004), .B(n7003), .Z(n7293) );
  NANDN U8804 ( .A(n7292), .B(n7293), .Z(n7295) );
  NAND U8805 ( .A(a[49]), .B(b[44]), .Z(n7288) );
  NANDN U8806 ( .A(n7288), .B(n7289), .Z(n7291) );
  NAND U8807 ( .A(a[48]), .B(b[44]), .Z(n7284) );
  XOR U8808 ( .A(n7008), .B(n7007), .Z(n7285) );
  NANDN U8809 ( .A(n7284), .B(n7285), .Z(n7287) );
  NAND U8810 ( .A(a[47]), .B(b[44]), .Z(n7280) );
  XNOR U8811 ( .A(n7010), .B(n7009), .Z(n7281) );
  NANDN U8812 ( .A(n7280), .B(n7281), .Z(n7283) );
  XOR U8813 ( .A(n7012), .B(n7011), .Z(n7277) );
  AND U8814 ( .A(a[46]), .B(b[44]), .Z(n7276) );
  NAND U8815 ( .A(n7277), .B(n7276), .Z(n7279) );
  NAND U8816 ( .A(a[44]), .B(b[44]), .Z(n7266) );
  AND U8817 ( .A(a[43]), .B(b[44]), .Z(n7016) );
  XNOR U8818 ( .A(n7014), .B(n7013), .Z(n7015) );
  NANDN U8819 ( .A(n7016), .B(n7015), .Z(n7263) );
  XOR U8820 ( .A(n7016), .B(n7015), .Z(n7334) );
  XOR U8821 ( .A(n7018), .B(n7017), .Z(n7253) );
  XOR U8822 ( .A(n7020), .B(n7019), .Z(n7021) );
  AND U8823 ( .A(a[39]), .B(b[44]), .Z(n7022) );
  NANDN U8824 ( .A(n7021), .B(n7022), .Z(n7245) );
  XOR U8825 ( .A(n7022), .B(n7021), .Z(n7342) );
  NAND U8826 ( .A(a[38]), .B(b[44]), .Z(n7240) );
  XNOR U8827 ( .A(n7024), .B(n7023), .Z(n7241) );
  NANDN U8828 ( .A(n7240), .B(n7241), .Z(n7243) );
  XOR U8829 ( .A(n7026), .B(n7025), .Z(n7230) );
  AND U8830 ( .A(a[36]), .B(b[44]), .Z(n7231) );
  NANDN U8831 ( .A(n7230), .B(n7231), .Z(n7233) );
  XOR U8832 ( .A(n7028), .B(n7027), .Z(n7030) );
  AND U8833 ( .A(a[35]), .B(b[44]), .Z(n7029) );
  NANDN U8834 ( .A(n7030), .B(n7029), .Z(n7229) );
  XOR U8835 ( .A(n7030), .B(n7029), .Z(n7346) );
  XOR U8836 ( .A(n7032), .B(n7031), .Z(n7224) );
  AND U8837 ( .A(a[34]), .B(b[44]), .Z(n7225) );
  NANDN U8838 ( .A(n7224), .B(n7225), .Z(n7227) );
  XOR U8839 ( .A(n7034), .B(n7033), .Z(n7221) );
  AND U8840 ( .A(a[33]), .B(b[44]), .Z(n7220) );
  NANDN U8841 ( .A(n7221), .B(n7220), .Z(n7223) );
  XOR U8842 ( .A(n7036), .B(n7035), .Z(n7217) );
  XOR U8843 ( .A(n7038), .B(n7037), .Z(n7212) );
  AND U8844 ( .A(a[31]), .B(b[44]), .Z(n7213) );
  NANDN U8845 ( .A(n7212), .B(n7213), .Z(n7215) );
  XOR U8846 ( .A(n7040), .B(n7039), .Z(n7208) );
  AND U8847 ( .A(a[30]), .B(b[44]), .Z(n7209) );
  NANDN U8848 ( .A(n7208), .B(n7209), .Z(n7211) );
  XOR U8849 ( .A(n7042), .B(n7041), .Z(n7205) );
  AND U8850 ( .A(a[29]), .B(b[44]), .Z(n7204) );
  NANDN U8851 ( .A(n7205), .B(n7204), .Z(n7207) );
  XOR U8852 ( .A(n7044), .B(n7043), .Z(n7194) );
  AND U8853 ( .A(a[27]), .B(b[44]), .Z(n7195) );
  NANDN U8854 ( .A(n7194), .B(n7195), .Z(n7197) );
  XOR U8855 ( .A(n7046), .B(n7045), .Z(n7179) );
  NAND U8856 ( .A(a[23]), .B(b[44]), .Z(n7174) );
  XNOR U8857 ( .A(n7048), .B(n7047), .Z(n7175) );
  NANDN U8858 ( .A(n7174), .B(n7175), .Z(n7177) );
  NAND U8859 ( .A(a[19]), .B(b[44]), .Z(n7152) );
  XOR U8860 ( .A(n7050), .B(n7049), .Z(n7153) );
  NANDN U8861 ( .A(n7152), .B(n7153), .Z(n7155) );
  NAND U8862 ( .A(a[15]), .B(b[44]), .Z(n7130) );
  NANDN U8863 ( .A(n7130), .B(n7131), .Z(n7133) );
  NAND U8864 ( .A(a[14]), .B(b[44]), .Z(n7126) );
  XOR U8865 ( .A(n7054), .B(n7053), .Z(n7127) );
  NANDN U8866 ( .A(n7126), .B(n7127), .Z(n7129) );
  AND U8867 ( .A(a[11]), .B(b[44]), .Z(n7108) );
  XOR U8868 ( .A(n7056), .B(n7055), .Z(n7098) );
  NAND U8869 ( .A(a[8]), .B(b[44]), .Z(n7059) );
  NANDN U8870 ( .A(n7059), .B(n7060), .Z(n7097) );
  NAND U8871 ( .A(a[7]), .B(b[44]), .Z(n7092) );
  XOR U8872 ( .A(n7062), .B(n7061), .Z(n7093) );
  NANDN U8873 ( .A(n7092), .B(n7093), .Z(n7095) );
  NAND U8874 ( .A(a[0]), .B(b[44]), .Z(n7728) );
  AND U8875 ( .A(a[1]), .B(b[45]), .Z(n7065) );
  NANDN U8876 ( .A(n7728), .B(n7065), .Z(n7390) );
  NANDN U8877 ( .A(n7390), .B(n7063), .Z(n7067) );
  AND U8878 ( .A(a[2]), .B(b[44]), .Z(n7396) );
  NANDN U8879 ( .A(n7395), .B(n7396), .Z(n7066) );
  AND U8880 ( .A(n7067), .B(n7066), .Z(n7070) );
  AND U8881 ( .A(a[3]), .B(b[44]), .Z(n7071) );
  NANDN U8882 ( .A(n7070), .B(n7071), .Z(n7073) );
  XOR U8883 ( .A(n7069), .B(n7068), .Z(n7401) );
  NANDN U8884 ( .A(n7401), .B(n7402), .Z(n7072) );
  AND U8885 ( .A(n7073), .B(n7072), .Z(n7076) );
  NANDN U8886 ( .A(n7076), .B(n7077), .Z(n7079) );
  NAND U8887 ( .A(a[4]), .B(b[44]), .Z(n7407) );
  NANDN U8888 ( .A(n7407), .B(n7408), .Z(n7078) );
  AND U8889 ( .A(n7079), .B(n7078), .Z(n7082) );
  XOR U8890 ( .A(n7081), .B(n7080), .Z(n7083) );
  NANDN U8891 ( .A(n7082), .B(n7083), .Z(n7085) );
  AND U8892 ( .A(a[5]), .B(b[44]), .Z(n7414) );
  NAND U8893 ( .A(n7414), .B(n7413), .Z(n7084) );
  AND U8894 ( .A(n7085), .B(n7084), .Z(n7088) );
  XNOR U8895 ( .A(n7087), .B(n7086), .Z(n7089) );
  NANDN U8896 ( .A(n7088), .B(n7089), .Z(n7091) );
  AND U8897 ( .A(a[6]), .B(b[44]), .Z(n7389) );
  NAND U8898 ( .A(n7389), .B(n7388), .Z(n7090) );
  AND U8899 ( .A(n7091), .B(n7090), .Z(n7384) );
  NANDN U8900 ( .A(n7384), .B(n7385), .Z(n7094) );
  NAND U8901 ( .A(n7095), .B(n7094), .Z(n7382) );
  NAND U8902 ( .A(n7383), .B(n7382), .Z(n7096) );
  AND U8903 ( .A(n7097), .B(n7096), .Z(n7099) );
  NANDN U8904 ( .A(n7098), .B(n7099), .Z(n7101) );
  AND U8905 ( .A(a[9]), .B(b[44]), .Z(n7429) );
  NANDN U8906 ( .A(n7429), .B(n7430), .Z(n7100) );
  AND U8907 ( .A(n7101), .B(n7100), .Z(n7104) );
  NAND U8908 ( .A(n7104), .B(n7105), .Z(n7107) );
  AND U8909 ( .A(a[10]), .B(b[44]), .Z(n7379) );
  XOR U8910 ( .A(n7105), .B(n7104), .Z(n7378) );
  NAND U8911 ( .A(n7379), .B(n7378), .Z(n7106) );
  AND U8912 ( .A(n7107), .B(n7106), .Z(n7109) );
  NANDN U8913 ( .A(n7108), .B(n7109), .Z(n7113) );
  XNOR U8914 ( .A(n7111), .B(n7110), .Z(n7376) );
  NAND U8915 ( .A(n7377), .B(n7376), .Z(n7112) );
  AND U8916 ( .A(n7113), .B(n7112), .Z(n7117) );
  NAND U8917 ( .A(n7117), .B(n7116), .Z(n7119) );
  AND U8918 ( .A(a[12]), .B(b[44]), .Z(n7442) );
  XOR U8919 ( .A(n7117), .B(n7116), .Z(n7441) );
  NAND U8920 ( .A(n7442), .B(n7441), .Z(n7118) );
  AND U8921 ( .A(n7119), .B(n7118), .Z(n7122) );
  XOR U8922 ( .A(n7121), .B(n7120), .Z(n7123) );
  NANDN U8923 ( .A(n7122), .B(n7123), .Z(n7125) );
  AND U8924 ( .A(a[13]), .B(b[44]), .Z(n7375) );
  NAND U8925 ( .A(n7375), .B(n7374), .Z(n7124) );
  AND U8926 ( .A(n7125), .B(n7124), .Z(n7372) );
  NANDN U8927 ( .A(n7372), .B(n7373), .Z(n7128) );
  AND U8928 ( .A(n7129), .B(n7128), .Z(n7457) );
  NANDN U8929 ( .A(n7457), .B(n7458), .Z(n7132) );
  AND U8930 ( .A(n7133), .B(n7132), .Z(n7136) );
  AND U8931 ( .A(a[16]), .B(b[44]), .Z(n7137) );
  NANDN U8932 ( .A(n7136), .B(n7137), .Z(n7139) );
  NAND U8933 ( .A(n7371), .B(n7370), .Z(n7138) );
  AND U8934 ( .A(n7139), .B(n7138), .Z(n7143) );
  XOR U8935 ( .A(n7141), .B(n7140), .Z(n7142) );
  NAND U8936 ( .A(n7143), .B(n7142), .Z(n7145) );
  AND U8937 ( .A(a[17]), .B(b[44]), .Z(n7465) );
  XOR U8938 ( .A(n7143), .B(n7142), .Z(n7466) );
  NANDN U8939 ( .A(n7465), .B(n7466), .Z(n7144) );
  AND U8940 ( .A(n7145), .B(n7144), .Z(n7149) );
  NAND U8941 ( .A(n7149), .B(n7148), .Z(n7151) );
  XOR U8942 ( .A(n7149), .B(n7148), .Z(n7369) );
  AND U8943 ( .A(a[18]), .B(b[44]), .Z(n7368) );
  NAND U8944 ( .A(n7369), .B(n7368), .Z(n7150) );
  AND U8945 ( .A(n7151), .B(n7150), .Z(n7477) );
  NANDN U8946 ( .A(n7477), .B(n7478), .Z(n7154) );
  AND U8947 ( .A(n7155), .B(n7154), .Z(n7156) );
  AND U8948 ( .A(a[20]), .B(b[44]), .Z(n7157) );
  NANDN U8949 ( .A(n7156), .B(n7157), .Z(n7161) );
  XOR U8950 ( .A(n7159), .B(n7158), .Z(n7481) );
  NAND U8951 ( .A(n7482), .B(n7481), .Z(n7160) );
  AND U8952 ( .A(n7161), .B(n7160), .Z(n7165) );
  XNOR U8953 ( .A(n7163), .B(n7162), .Z(n7164) );
  NANDN U8954 ( .A(n7165), .B(n7164), .Z(n7167) );
  XNOR U8955 ( .A(n7165), .B(n7164), .Z(n7367) );
  AND U8956 ( .A(a[21]), .B(b[44]), .Z(n7366) );
  NAND U8957 ( .A(n7367), .B(n7366), .Z(n7166) );
  AND U8958 ( .A(n7167), .B(n7166), .Z(n7171) );
  XNOR U8959 ( .A(n7169), .B(n7168), .Z(n7170) );
  NANDN U8960 ( .A(n7171), .B(n7170), .Z(n7173) );
  NAND U8961 ( .A(a[22]), .B(b[44]), .Z(n7491) );
  XNOR U8962 ( .A(n7171), .B(n7170), .Z(n7492) );
  NANDN U8963 ( .A(n7491), .B(n7492), .Z(n7172) );
  AND U8964 ( .A(n7173), .B(n7172), .Z(n7365) );
  XNOR U8965 ( .A(n7175), .B(n7174), .Z(n7364) );
  NANDN U8966 ( .A(n7365), .B(n7364), .Z(n7176) );
  NAND U8967 ( .A(n7177), .B(n7176), .Z(n7178) );
  NANDN U8968 ( .A(n7179), .B(n7178), .Z(n7181) );
  NAND U8969 ( .A(a[24]), .B(b[44]), .Z(n7501) );
  XNOR U8970 ( .A(n7179), .B(n7178), .Z(n7502) );
  NANDN U8971 ( .A(n7501), .B(n7502), .Z(n7180) );
  AND U8972 ( .A(n7181), .B(n7180), .Z(n7185) );
  XNOR U8973 ( .A(n7183), .B(n7182), .Z(n7184) );
  NANDN U8974 ( .A(n7185), .B(n7184), .Z(n7187) );
  NAND U8975 ( .A(a[25]), .B(b[44]), .Z(n7362) );
  XNOR U8976 ( .A(n7185), .B(n7184), .Z(n7363) );
  NANDN U8977 ( .A(n7362), .B(n7363), .Z(n7186) );
  AND U8978 ( .A(n7187), .B(n7186), .Z(n7191) );
  AND U8979 ( .A(a[26]), .B(b[44]), .Z(n7190) );
  NANDN U8980 ( .A(n7191), .B(n7190), .Z(n7193) );
  XOR U8981 ( .A(n7189), .B(n7188), .Z(n7511) );
  XNOR U8982 ( .A(n7191), .B(n7190), .Z(n7512) );
  NANDN U8983 ( .A(n7511), .B(n7512), .Z(n7192) );
  AND U8984 ( .A(n7193), .B(n7192), .Z(n7518) );
  XNOR U8985 ( .A(n7195), .B(n7194), .Z(n7517) );
  NANDN U8986 ( .A(n7518), .B(n7517), .Z(n7196) );
  AND U8987 ( .A(n7197), .B(n7196), .Z(n7201) );
  XNOR U8988 ( .A(n7199), .B(n7198), .Z(n7200) );
  NANDN U8989 ( .A(n7201), .B(n7200), .Z(n7203) );
  NAND U8990 ( .A(a[28]), .B(b[44]), .Z(n7360) );
  XNOR U8991 ( .A(n7201), .B(n7200), .Z(n7361) );
  NANDN U8992 ( .A(n7360), .B(n7361), .Z(n7202) );
  AND U8993 ( .A(n7203), .B(n7202), .Z(n7357) );
  XNOR U8994 ( .A(n7205), .B(n7204), .Z(n7356) );
  NANDN U8995 ( .A(n7357), .B(n7356), .Z(n7206) );
  AND U8996 ( .A(n7207), .B(n7206), .Z(n7355) );
  XNOR U8997 ( .A(n7209), .B(n7208), .Z(n7354) );
  NANDN U8998 ( .A(n7355), .B(n7354), .Z(n7210) );
  AND U8999 ( .A(n7211), .B(n7210), .Z(n7534) );
  XNOR U9000 ( .A(n7213), .B(n7212), .Z(n7533) );
  NANDN U9001 ( .A(n7534), .B(n7533), .Z(n7214) );
  NAND U9002 ( .A(n7215), .B(n7214), .Z(n7216) );
  NANDN U9003 ( .A(n7217), .B(n7216), .Z(n7219) );
  XNOR U9004 ( .A(n7217), .B(n7216), .Z(n7353) );
  AND U9005 ( .A(a[32]), .B(b[44]), .Z(n7352) );
  NAND U9006 ( .A(n7353), .B(n7352), .Z(n7218) );
  AND U9007 ( .A(n7219), .B(n7218), .Z(n7349) );
  XNOR U9008 ( .A(n7221), .B(n7220), .Z(n7348) );
  NANDN U9009 ( .A(n7349), .B(n7348), .Z(n7222) );
  AND U9010 ( .A(n7223), .B(n7222), .Z(n7546) );
  XNOR U9011 ( .A(n7225), .B(n7224), .Z(n7545) );
  NANDN U9012 ( .A(n7546), .B(n7545), .Z(n7226) );
  AND U9013 ( .A(n7227), .B(n7226), .Z(n7347) );
  OR U9014 ( .A(n7346), .B(n7347), .Z(n7228) );
  AND U9015 ( .A(n7229), .B(n7228), .Z(n7345) );
  XNOR U9016 ( .A(n7231), .B(n7230), .Z(n7344) );
  NANDN U9017 ( .A(n7345), .B(n7344), .Z(n7232) );
  AND U9018 ( .A(n7233), .B(n7232), .Z(n7237) );
  XNOR U9019 ( .A(n7235), .B(n7234), .Z(n7236) );
  NANDN U9020 ( .A(n7237), .B(n7236), .Z(n7239) );
  NAND U9021 ( .A(a[37]), .B(b[44]), .Z(n7561) );
  XNOR U9022 ( .A(n7237), .B(n7236), .Z(n7562) );
  NANDN U9023 ( .A(n7561), .B(n7562), .Z(n7238) );
  AND U9024 ( .A(n7239), .B(n7238), .Z(n7566) );
  XNOR U9025 ( .A(n7241), .B(n7240), .Z(n7565) );
  NANDN U9026 ( .A(n7566), .B(n7565), .Z(n7242) );
  AND U9027 ( .A(n7243), .B(n7242), .Z(n7343) );
  OR U9028 ( .A(n7342), .B(n7343), .Z(n7244) );
  AND U9029 ( .A(n7245), .B(n7244), .Z(n7249) );
  XNOR U9030 ( .A(n7247), .B(n7246), .Z(n7248) );
  NANDN U9031 ( .A(n7249), .B(n7248), .Z(n7251) );
  NAND U9032 ( .A(a[40]), .B(b[44]), .Z(n7575) );
  XNOR U9033 ( .A(n7249), .B(n7248), .Z(n7576) );
  NANDN U9034 ( .A(n7575), .B(n7576), .Z(n7250) );
  AND U9035 ( .A(n7251), .B(n7250), .Z(n7252) );
  NANDN U9036 ( .A(n7253), .B(n7252), .Z(n7255) );
  AND U9037 ( .A(a[41]), .B(b[44]), .Z(n7341) );
  XNOR U9038 ( .A(n7253), .B(n7252), .Z(n7340) );
  NANDN U9039 ( .A(n7341), .B(n7340), .Z(n7254) );
  AND U9040 ( .A(n7255), .B(n7254), .Z(n7259) );
  XNOR U9041 ( .A(n7257), .B(n7256), .Z(n7258) );
  NANDN U9042 ( .A(n7259), .B(n7258), .Z(n7261) );
  XOR U9043 ( .A(n7259), .B(n7258), .Z(n7338) );
  AND U9044 ( .A(a[42]), .B(b[44]), .Z(n7339) );
  OR U9045 ( .A(n7338), .B(n7339), .Z(n7260) );
  AND U9046 ( .A(n7261), .B(n7260), .Z(n7335) );
  OR U9047 ( .A(n7334), .B(n7335), .Z(n7262) );
  AND U9048 ( .A(n7263), .B(n7262), .Z(n7267) );
  NANDN U9049 ( .A(n7266), .B(n7267), .Z(n7269) );
  XOR U9050 ( .A(n7265), .B(n7264), .Z(n7591) );
  XNOR U9051 ( .A(n7267), .B(n7266), .Z(n7592) );
  NANDN U9052 ( .A(n7591), .B(n7592), .Z(n7268) );
  AND U9053 ( .A(n7269), .B(n7268), .Z(n7273) );
  XOR U9054 ( .A(n7271), .B(n7270), .Z(n7272) );
  NANDN U9055 ( .A(n7273), .B(n7272), .Z(n7275) );
  XNOR U9056 ( .A(n7273), .B(n7272), .Z(n7333) );
  AND U9057 ( .A(a[45]), .B(b[44]), .Z(n7332) );
  NAND U9058 ( .A(n7333), .B(n7332), .Z(n7274) );
  AND U9059 ( .A(n7275), .B(n7274), .Z(n7602) );
  XOR U9060 ( .A(n7277), .B(n7276), .Z(n7601) );
  NANDN U9061 ( .A(n7602), .B(n7601), .Z(n7278) );
  AND U9062 ( .A(n7279), .B(n7278), .Z(n7329) );
  XNOR U9063 ( .A(n7281), .B(n7280), .Z(n7328) );
  NANDN U9064 ( .A(n7329), .B(n7328), .Z(n7282) );
  AND U9065 ( .A(n7283), .B(n7282), .Z(n7610) );
  XNOR U9066 ( .A(n7285), .B(n7284), .Z(n7609) );
  NANDN U9067 ( .A(n7610), .B(n7609), .Z(n7286) );
  AND U9068 ( .A(n7287), .B(n7286), .Z(n7615) );
  NANDN U9069 ( .A(n7615), .B(n7616), .Z(n7290) );
  AND U9070 ( .A(n7291), .B(n7290), .Z(n7622) );
  NANDN U9071 ( .A(n7622), .B(n7621), .Z(n7294) );
  AND U9072 ( .A(n7295), .B(n7294), .Z(n7297) );
  NANDN U9073 ( .A(n7296), .B(n7297), .Z(n7301) );
  XNOR U9074 ( .A(n7299), .B(n7298), .Z(n7327) );
  NAND U9075 ( .A(n7326), .B(n7327), .Z(n7300) );
  NAND U9076 ( .A(n7301), .B(n7300), .Z(n7303) );
  NANDN U9077 ( .A(n7302), .B(n7303), .Z(n7307) );
  NAND U9078 ( .A(n7632), .B(n7631), .Z(n7306) );
  NAND U9079 ( .A(n7307), .B(n7306), .Z(n7310) );
  NAND U9080 ( .A(n7311), .B(n7310), .Z(n7313) );
  XOR U9081 ( .A(n7309), .B(n7308), .Z(n7637) );
  XOR U9082 ( .A(n7311), .B(n7310), .Z(n7638) );
  NANDN U9083 ( .A(n7637), .B(n7638), .Z(n7312) );
  AND U9084 ( .A(n7313), .B(n7312), .Z(n7316) );
  NAND U9085 ( .A(n7317), .B(n7316), .Z(n7319) );
  XOR U9086 ( .A(n7315), .B(n7314), .Z(n7644) );
  XOR U9087 ( .A(n7317), .B(n7316), .Z(n7643) );
  NAND U9088 ( .A(n7644), .B(n7643), .Z(n7318) );
  AND U9089 ( .A(n7319), .B(n7318), .Z(n7322) );
  NAND U9090 ( .A(a[55]), .B(b[44]), .Z(n7323) );
  NAND U9091 ( .A(n7322), .B(n7323), .Z(n7325) );
  XOR U9092 ( .A(n7321), .B(n7320), .Z(n7649) );
  XOR U9093 ( .A(n7323), .B(n7322), .Z(n7650) );
  NANDN U9094 ( .A(n7649), .B(n7650), .Z(n7324) );
  NAND U9095 ( .A(n7325), .B(n7324), .Z(n10220) );
  XOR U9096 ( .A(n10221), .B(n10220), .Z(n10222) );
  NAND U9097 ( .A(a[57]), .B(b[43]), .Z(n10226) );
  AND U9098 ( .A(a[56]), .B(b[43]), .Z(n7652) );
  AND U9099 ( .A(a[54]), .B(b[43]), .Z(n7640) );
  AND U9100 ( .A(a[52]), .B(b[43]), .Z(n7627) );
  XOR U9101 ( .A(n7327), .B(n7326), .Z(n7628) );
  NANDN U9102 ( .A(n7627), .B(n7628), .Z(n7630) );
  NAND U9103 ( .A(a[48]), .B(b[43]), .Z(n7330) );
  XNOR U9104 ( .A(n7329), .B(n7328), .Z(n7331) );
  NANDN U9105 ( .A(n7330), .B(n7331), .Z(n7608) );
  XOR U9106 ( .A(n7331), .B(n7330), .Z(n7665) );
  XOR U9107 ( .A(n7333), .B(n7332), .Z(n7598) );
  XOR U9108 ( .A(n7335), .B(n7334), .Z(n7337) );
  AND U9109 ( .A(a[44]), .B(b[43]), .Z(n7336) );
  NANDN U9110 ( .A(n7337), .B(n7336), .Z(n7590) );
  XOR U9111 ( .A(n7337), .B(n7336), .Z(n7673) );
  XOR U9112 ( .A(n7339), .B(n7338), .Z(n7586) );
  XOR U9113 ( .A(n7341), .B(n7340), .Z(n7581) );
  XOR U9114 ( .A(n7343), .B(n7342), .Z(n7572) );
  NAND U9115 ( .A(a[37]), .B(b[43]), .Z(n7555) );
  XNOR U9116 ( .A(n7345), .B(n7344), .Z(n7556) );
  NANDN U9117 ( .A(n7555), .B(n7556), .Z(n7558) );
  XOR U9118 ( .A(n7347), .B(n7346), .Z(n7552) );
  XOR U9119 ( .A(n7349), .B(n7348), .Z(n7350) );
  AND U9120 ( .A(a[34]), .B(b[43]), .Z(n7351) );
  NANDN U9121 ( .A(n7350), .B(n7351), .Z(n7544) );
  XOR U9122 ( .A(n7351), .B(n7350), .Z(n7691) );
  AND U9123 ( .A(a[33]), .B(b[43]), .Z(n7540) );
  XNOR U9124 ( .A(n7353), .B(n7352), .Z(n7539) );
  NANDN U9125 ( .A(n7540), .B(n7539), .Z(n7542) );
  XOR U9126 ( .A(n7355), .B(n7354), .Z(n7529) );
  AND U9127 ( .A(a[31]), .B(b[43]), .Z(n7530) );
  NANDN U9128 ( .A(n7529), .B(n7530), .Z(n7532) );
  NAND U9129 ( .A(a[30]), .B(b[43]), .Z(n7358) );
  XNOR U9130 ( .A(n7357), .B(n7356), .Z(n7359) );
  NANDN U9131 ( .A(n7358), .B(n7359), .Z(n7528) );
  XOR U9132 ( .A(n7359), .B(n7358), .Z(n7699) );
  NAND U9133 ( .A(a[29]), .B(b[43]), .Z(n7523) );
  XNOR U9134 ( .A(n7361), .B(n7360), .Z(n7524) );
  NANDN U9135 ( .A(n7523), .B(n7524), .Z(n7526) );
  XOR U9136 ( .A(n7363), .B(n7362), .Z(n7507) );
  AND U9137 ( .A(a[26]), .B(b[43]), .Z(n7508) );
  NANDN U9138 ( .A(n7507), .B(n7508), .Z(n7510) );
  NAND U9139 ( .A(a[24]), .B(b[43]), .Z(n7497) );
  XNOR U9140 ( .A(n7365), .B(n7364), .Z(n7498) );
  NANDN U9141 ( .A(n7497), .B(n7498), .Z(n7500) );
  XOR U9142 ( .A(n7367), .B(n7366), .Z(n7488) );
  NAND U9143 ( .A(a[20]), .B(b[43]), .Z(n7475) );
  XOR U9144 ( .A(n7369), .B(n7368), .Z(n7471) );
  XOR U9145 ( .A(n7371), .B(n7370), .Z(n7461) );
  NAND U9146 ( .A(a[15]), .B(b[43]), .Z(n7451) );
  NANDN U9147 ( .A(n7451), .B(n7452), .Z(n7454) );
  NAND U9148 ( .A(a[14]), .B(b[43]), .Z(n7447) );
  XOR U9149 ( .A(n7375), .B(n7374), .Z(n7448) );
  NANDN U9150 ( .A(n7447), .B(n7448), .Z(n7450) );
  XOR U9151 ( .A(n7377), .B(n7376), .Z(n7437) );
  AND U9152 ( .A(a[11]), .B(b[43]), .Z(n7380) );
  XNOR U9153 ( .A(n7379), .B(n7378), .Z(n7381) );
  NANDN U9154 ( .A(n7380), .B(n7381), .Z(n7436) );
  XOR U9155 ( .A(n7383), .B(n7382), .Z(n7425) );
  NAND U9156 ( .A(a[8]), .B(b[43]), .Z(n7386) );
  NANDN U9157 ( .A(n7386), .B(n7387), .Z(n7424) );
  NAND U9158 ( .A(a[7]), .B(b[43]), .Z(n7419) );
  XOR U9159 ( .A(n7389), .B(n7388), .Z(n7420) );
  NANDN U9160 ( .A(n7419), .B(n7420), .Z(n7422) );
  NAND U9161 ( .A(a[0]), .B(b[43]), .Z(n8061) );
  AND U9162 ( .A(a[1]), .B(b[44]), .Z(n7392) );
  NANDN U9163 ( .A(n8061), .B(n7392), .Z(n7727) );
  NANDN U9164 ( .A(n7727), .B(n7390), .Z(n7394) );
  AND U9165 ( .A(a[2]), .B(b[43]), .Z(n7733) );
  NANDN U9166 ( .A(n7732), .B(n7733), .Z(n7393) );
  AND U9167 ( .A(n7394), .B(n7393), .Z(n7397) );
  AND U9168 ( .A(a[3]), .B(b[43]), .Z(n7398) );
  NANDN U9169 ( .A(n7397), .B(n7398), .Z(n7400) );
  XOR U9170 ( .A(n7396), .B(n7395), .Z(n7738) );
  NANDN U9171 ( .A(n7738), .B(n7739), .Z(n7399) );
  AND U9172 ( .A(n7400), .B(n7399), .Z(n7403) );
  NANDN U9173 ( .A(n7403), .B(n7404), .Z(n7406) );
  AND U9174 ( .A(a[4]), .B(b[43]), .Z(n7745) );
  NAND U9175 ( .A(n7745), .B(n7744), .Z(n7405) );
  AND U9176 ( .A(n7406), .B(n7405), .Z(n7409) );
  NANDN U9177 ( .A(n7409), .B(n7410), .Z(n7412) );
  NAND U9178 ( .A(a[5]), .B(b[43]), .Z(n7750) );
  NANDN U9179 ( .A(n7750), .B(n7751), .Z(n7411) );
  AND U9180 ( .A(n7412), .B(n7411), .Z(n7415) );
  XOR U9181 ( .A(n7414), .B(n7413), .Z(n7416) );
  NANDN U9182 ( .A(n7415), .B(n7416), .Z(n7418) );
  AND U9183 ( .A(a[6]), .B(b[43]), .Z(n7726) );
  NAND U9184 ( .A(n7726), .B(n7725), .Z(n7417) );
  AND U9185 ( .A(n7418), .B(n7417), .Z(n7721) );
  NANDN U9186 ( .A(n7721), .B(n7722), .Z(n7421) );
  NAND U9187 ( .A(n7422), .B(n7421), .Z(n7719) );
  NAND U9188 ( .A(n7720), .B(n7719), .Z(n7423) );
  AND U9189 ( .A(n7424), .B(n7423), .Z(n7426) );
  NANDN U9190 ( .A(n7425), .B(n7426), .Z(n7428) );
  AND U9191 ( .A(a[9]), .B(b[43]), .Z(n7766) );
  NANDN U9192 ( .A(n7766), .B(n7767), .Z(n7427) );
  AND U9193 ( .A(n7428), .B(n7427), .Z(n7431) );
  NANDN U9194 ( .A(n7431), .B(n7432), .Z(n7434) );
  AND U9195 ( .A(a[10]), .B(b[43]), .Z(n7772) );
  NANDN U9196 ( .A(n7772), .B(n7773), .Z(n7433) );
  NAND U9197 ( .A(n7434), .B(n7433), .Z(n7717) );
  NAND U9198 ( .A(n7718), .B(n7717), .Z(n7435) );
  AND U9199 ( .A(n7436), .B(n7435), .Z(n7438) );
  NANDN U9200 ( .A(n7437), .B(n7438), .Z(n7440) );
  AND U9201 ( .A(a[12]), .B(b[43]), .Z(n7783) );
  NAND U9202 ( .A(n7783), .B(n7782), .Z(n7439) );
  AND U9203 ( .A(n7440), .B(n7439), .Z(n7443) );
  XOR U9204 ( .A(n7442), .B(n7441), .Z(n7444) );
  NANDN U9205 ( .A(n7443), .B(n7444), .Z(n7446) );
  AND U9206 ( .A(a[13]), .B(b[43]), .Z(n7716) );
  NAND U9207 ( .A(n7716), .B(n7715), .Z(n7445) );
  AND U9208 ( .A(n7446), .B(n7445), .Z(n7713) );
  NANDN U9209 ( .A(n7713), .B(n7714), .Z(n7449) );
  AND U9210 ( .A(n7450), .B(n7449), .Z(n7798) );
  NANDN U9211 ( .A(n7798), .B(n7799), .Z(n7453) );
  AND U9212 ( .A(n7454), .B(n7453), .Z(n7455) );
  AND U9213 ( .A(a[16]), .B(b[43]), .Z(n7456) );
  NANDN U9214 ( .A(n7455), .B(n7456), .Z(n7460) );
  NAND U9215 ( .A(n7712), .B(n7711), .Z(n7459) );
  AND U9216 ( .A(n7460), .B(n7459), .Z(n7462) );
  NANDN U9217 ( .A(n7461), .B(n7462), .Z(n7464) );
  AND U9218 ( .A(a[17]), .B(b[43]), .Z(n7806) );
  NANDN U9219 ( .A(n7806), .B(n7807), .Z(n7463) );
  AND U9220 ( .A(n7464), .B(n7463), .Z(n7467) );
  NAND U9221 ( .A(n7467), .B(n7468), .Z(n7470) );
  AND U9222 ( .A(a[18]), .B(b[43]), .Z(n7710) );
  XOR U9223 ( .A(n7468), .B(n7467), .Z(n7709) );
  NAND U9224 ( .A(n7710), .B(n7709), .Z(n7469) );
  AND U9225 ( .A(n7470), .B(n7469), .Z(n7472) );
  NANDN U9226 ( .A(n7471), .B(n7472), .Z(n7474) );
  AND U9227 ( .A(a[19]), .B(b[43]), .Z(n7818) );
  NANDN U9228 ( .A(n7818), .B(n7819), .Z(n7473) );
  AND U9229 ( .A(n7474), .B(n7473), .Z(n7476) );
  NANDN U9230 ( .A(n7475), .B(n7476), .Z(n7480) );
  NAND U9231 ( .A(n7823), .B(n7822), .Z(n7479) );
  AND U9232 ( .A(n7480), .B(n7479), .Z(n7483) );
  XOR U9233 ( .A(n7482), .B(n7481), .Z(n7484) );
  NANDN U9234 ( .A(n7483), .B(n7484), .Z(n7486) );
  AND U9235 ( .A(a[21]), .B(b[43]), .Z(n7829) );
  NAND U9236 ( .A(n7829), .B(n7828), .Z(n7485) );
  AND U9237 ( .A(n7486), .B(n7485), .Z(n7487) );
  NANDN U9238 ( .A(n7488), .B(n7487), .Z(n7490) );
  XOR U9239 ( .A(n7488), .B(n7487), .Z(n7834) );
  AND U9240 ( .A(a[22]), .B(b[43]), .Z(n7835) );
  OR U9241 ( .A(n7834), .B(n7835), .Z(n7489) );
  NAND U9242 ( .A(n7490), .B(n7489), .Z(n7493) );
  XNOR U9243 ( .A(n7492), .B(n7491), .Z(n7494) );
  NANDN U9244 ( .A(n7493), .B(n7494), .Z(n7496) );
  NAND U9245 ( .A(a[23]), .B(b[43]), .Z(n7707) );
  XNOR U9246 ( .A(n7494), .B(n7493), .Z(n7708) );
  NANDN U9247 ( .A(n7707), .B(n7708), .Z(n7495) );
  AND U9248 ( .A(n7496), .B(n7495), .Z(n7845) );
  XNOR U9249 ( .A(n7498), .B(n7497), .Z(n7844) );
  NANDN U9250 ( .A(n7845), .B(n7844), .Z(n7499) );
  AND U9251 ( .A(n7500), .B(n7499), .Z(n7504) );
  XNOR U9252 ( .A(n7502), .B(n7501), .Z(n7503) );
  NANDN U9253 ( .A(n7504), .B(n7503), .Z(n7506) );
  NAND U9254 ( .A(a[25]), .B(b[43]), .Z(n7850) );
  XNOR U9255 ( .A(n7504), .B(n7503), .Z(n7851) );
  NANDN U9256 ( .A(n7850), .B(n7851), .Z(n7505) );
  AND U9257 ( .A(n7506), .B(n7505), .Z(n7706) );
  XNOR U9258 ( .A(n7508), .B(n7507), .Z(n7705) );
  NANDN U9259 ( .A(n7706), .B(n7705), .Z(n7509) );
  AND U9260 ( .A(n7510), .B(n7509), .Z(n7514) );
  XNOR U9261 ( .A(n7512), .B(n7511), .Z(n7513) );
  NANDN U9262 ( .A(n7514), .B(n7513), .Z(n7516) );
  NAND U9263 ( .A(a[27]), .B(b[43]), .Z(n7703) );
  XNOR U9264 ( .A(n7514), .B(n7513), .Z(n7704) );
  NANDN U9265 ( .A(n7703), .B(n7704), .Z(n7515) );
  AND U9266 ( .A(n7516), .B(n7515), .Z(n7520) );
  XNOR U9267 ( .A(n7518), .B(n7517), .Z(n7519) );
  NANDN U9268 ( .A(n7520), .B(n7519), .Z(n7522) );
  NAND U9269 ( .A(a[28]), .B(b[43]), .Z(n7864) );
  XNOR U9270 ( .A(n7520), .B(n7519), .Z(n7865) );
  NANDN U9271 ( .A(n7864), .B(n7865), .Z(n7521) );
  AND U9272 ( .A(n7522), .B(n7521), .Z(n7702) );
  XNOR U9273 ( .A(n7524), .B(n7523), .Z(n7701) );
  NANDN U9274 ( .A(n7702), .B(n7701), .Z(n7525) );
  AND U9275 ( .A(n7526), .B(n7525), .Z(n7700) );
  OR U9276 ( .A(n7699), .B(n7700), .Z(n7527) );
  AND U9277 ( .A(n7528), .B(n7527), .Z(n7696) );
  XNOR U9278 ( .A(n7530), .B(n7529), .Z(n7695) );
  NANDN U9279 ( .A(n7696), .B(n7695), .Z(n7531) );
  AND U9280 ( .A(n7532), .B(n7531), .Z(n7536) );
  XNOR U9281 ( .A(n7534), .B(n7533), .Z(n7535) );
  NANDN U9282 ( .A(n7536), .B(n7535), .Z(n7538) );
  NAND U9283 ( .A(a[32]), .B(b[43]), .Z(n7880) );
  XNOR U9284 ( .A(n7536), .B(n7535), .Z(n7881) );
  NANDN U9285 ( .A(n7880), .B(n7881), .Z(n7537) );
  AND U9286 ( .A(n7538), .B(n7537), .Z(n7694) );
  XNOR U9287 ( .A(n7540), .B(n7539), .Z(n7693) );
  NAND U9288 ( .A(n7694), .B(n7693), .Z(n7541) );
  AND U9289 ( .A(n7542), .B(n7541), .Z(n7692) );
  NANDN U9290 ( .A(n7691), .B(n7692), .Z(n7543) );
  AND U9291 ( .A(n7544), .B(n7543), .Z(n7548) );
  XNOR U9292 ( .A(n7546), .B(n7545), .Z(n7547) );
  NANDN U9293 ( .A(n7548), .B(n7547), .Z(n7550) );
  NAND U9294 ( .A(a[35]), .B(b[43]), .Z(n7687) );
  XNOR U9295 ( .A(n7548), .B(n7547), .Z(n7688) );
  NANDN U9296 ( .A(n7687), .B(n7688), .Z(n7549) );
  AND U9297 ( .A(n7550), .B(n7549), .Z(n7551) );
  NANDN U9298 ( .A(n7552), .B(n7551), .Z(n7554) );
  XOR U9299 ( .A(n7552), .B(n7551), .Z(n7683) );
  AND U9300 ( .A(a[36]), .B(b[43]), .Z(n7684) );
  OR U9301 ( .A(n7683), .B(n7684), .Z(n7553) );
  NAND U9302 ( .A(n7554), .B(n7553), .Z(n7898) );
  XNOR U9303 ( .A(n7556), .B(n7555), .Z(n7899) );
  NANDN U9304 ( .A(n7898), .B(n7899), .Z(n7557) );
  AND U9305 ( .A(n7558), .B(n7557), .Z(n7560) );
  AND U9306 ( .A(a[38]), .B(b[43]), .Z(n7559) );
  NANDN U9307 ( .A(n7560), .B(n7559), .Z(n7564) );
  XOR U9308 ( .A(n7560), .B(n7559), .Z(n7681) );
  XNOR U9309 ( .A(n7562), .B(n7561), .Z(n7682) );
  NANDN U9310 ( .A(n7681), .B(n7682), .Z(n7563) );
  AND U9311 ( .A(n7564), .B(n7563), .Z(n7568) );
  XNOR U9312 ( .A(n7566), .B(n7565), .Z(n7567) );
  NANDN U9313 ( .A(n7568), .B(n7567), .Z(n7570) );
  NAND U9314 ( .A(a[39]), .B(b[43]), .Z(n7908) );
  XNOR U9315 ( .A(n7568), .B(n7567), .Z(n7909) );
  NANDN U9316 ( .A(n7908), .B(n7909), .Z(n7569) );
  AND U9317 ( .A(n7570), .B(n7569), .Z(n7571) );
  NANDN U9318 ( .A(n7572), .B(n7571), .Z(n7574) );
  XOR U9319 ( .A(n7572), .B(n7571), .Z(n7677) );
  AND U9320 ( .A(a[40]), .B(b[43]), .Z(n7678) );
  OR U9321 ( .A(n7677), .B(n7678), .Z(n7573) );
  NAND U9322 ( .A(n7574), .B(n7573), .Z(n7577) );
  XNOR U9323 ( .A(n7576), .B(n7575), .Z(n7578) );
  NANDN U9324 ( .A(n7577), .B(n7578), .Z(n7580) );
  NAND U9325 ( .A(a[41]), .B(b[43]), .Z(n7916) );
  XNOR U9326 ( .A(n7578), .B(n7577), .Z(n7917) );
  NANDN U9327 ( .A(n7916), .B(n7917), .Z(n7579) );
  AND U9328 ( .A(n7580), .B(n7579), .Z(n7582) );
  NANDN U9329 ( .A(n7581), .B(n7582), .Z(n7584) );
  XOR U9330 ( .A(n7582), .B(n7581), .Z(n7675) );
  AND U9331 ( .A(a[42]), .B(b[43]), .Z(n7676) );
  OR U9332 ( .A(n7675), .B(n7676), .Z(n7583) );
  AND U9333 ( .A(n7584), .B(n7583), .Z(n7585) );
  NANDN U9334 ( .A(n7586), .B(n7585), .Z(n7588) );
  NAND U9335 ( .A(a[43]), .B(b[43]), .Z(n7926) );
  XNOR U9336 ( .A(n7586), .B(n7585), .Z(n7927) );
  NANDN U9337 ( .A(n7926), .B(n7927), .Z(n7587) );
  AND U9338 ( .A(n7588), .B(n7587), .Z(n7674) );
  OR U9339 ( .A(n7673), .B(n7674), .Z(n7589) );
  AND U9340 ( .A(n7590), .B(n7589), .Z(n7594) );
  AND U9341 ( .A(a[45]), .B(b[43]), .Z(n7593) );
  NANDN U9342 ( .A(n7594), .B(n7593), .Z(n7596) );
  XOR U9343 ( .A(n7592), .B(n7591), .Z(n7671) );
  XNOR U9344 ( .A(n7594), .B(n7593), .Z(n7672) );
  NANDN U9345 ( .A(n7671), .B(n7672), .Z(n7595) );
  AND U9346 ( .A(n7596), .B(n7595), .Z(n7597) );
  NANDN U9347 ( .A(n7598), .B(n7597), .Z(n7600) );
  XOR U9348 ( .A(n7598), .B(n7597), .Z(n7669) );
  AND U9349 ( .A(a[46]), .B(b[43]), .Z(n7670) );
  OR U9350 ( .A(n7669), .B(n7670), .Z(n7599) );
  AND U9351 ( .A(n7600), .B(n7599), .Z(n7604) );
  XOR U9352 ( .A(n7602), .B(n7601), .Z(n7603) );
  NANDN U9353 ( .A(n7604), .B(n7603), .Z(n7606) );
  XOR U9354 ( .A(n7604), .B(n7603), .Z(n7944) );
  AND U9355 ( .A(a[47]), .B(b[43]), .Z(n7945) );
  OR U9356 ( .A(n7944), .B(n7945), .Z(n7605) );
  AND U9357 ( .A(n7606), .B(n7605), .Z(n7666) );
  NANDN U9358 ( .A(n7665), .B(n7666), .Z(n7607) );
  AND U9359 ( .A(n7608), .B(n7607), .Z(n7612) );
  XNOR U9360 ( .A(n7610), .B(n7609), .Z(n7611) );
  NANDN U9361 ( .A(n7612), .B(n7611), .Z(n7614) );
  NAND U9362 ( .A(a[49]), .B(b[43]), .Z(n7663) );
  XNOR U9363 ( .A(n7612), .B(n7611), .Z(n7664) );
  NANDN U9364 ( .A(n7663), .B(n7664), .Z(n7613) );
  AND U9365 ( .A(n7614), .B(n7613), .Z(n7617) );
  NAND U9366 ( .A(n7617), .B(n7618), .Z(n7620) );
  AND U9367 ( .A(a[50]), .B(b[43]), .Z(n7661) );
  XOR U9368 ( .A(n7618), .B(n7617), .Z(n7662) );
  NANDN U9369 ( .A(n7661), .B(n7662), .Z(n7619) );
  AND U9370 ( .A(n7620), .B(n7619), .Z(n7623) );
  XOR U9371 ( .A(n7622), .B(n7621), .Z(n7624) );
  NANDN U9372 ( .A(n7623), .B(n7624), .Z(n7626) );
  AND U9373 ( .A(a[51]), .B(b[43]), .Z(n7659) );
  NANDN U9374 ( .A(n7659), .B(n7660), .Z(n7625) );
  AND U9375 ( .A(n7626), .B(n7625), .Z(n7657) );
  NANDN U9376 ( .A(n7657), .B(n7658), .Z(n7629) );
  NAND U9377 ( .A(n7630), .B(n7629), .Z(n7633) );
  AND U9378 ( .A(a[53]), .B(b[43]), .Z(n7634) );
  NANDN U9379 ( .A(n7633), .B(n7634), .Z(n7636) );
  XOR U9380 ( .A(n7632), .B(n7631), .Z(n7655) );
  NANDN U9381 ( .A(n7655), .B(n7656), .Z(n7635) );
  NAND U9382 ( .A(n7636), .B(n7635), .Z(n7639) );
  NAND U9383 ( .A(n7640), .B(n7639), .Z(n7642) );
  XOR U9384 ( .A(n7640), .B(n7639), .Z(n7974) );
  NAND U9385 ( .A(n7975), .B(n7974), .Z(n7641) );
  AND U9386 ( .A(n7642), .B(n7641), .Z(n7645) );
  NAND U9387 ( .A(a[55]), .B(b[43]), .Z(n7646) );
  NAND U9388 ( .A(n7645), .B(n7646), .Z(n7648) );
  XOR U9389 ( .A(n7644), .B(n7643), .Z(n7978) );
  XOR U9390 ( .A(n7646), .B(n7645), .Z(n7979) );
  NANDN U9391 ( .A(n7978), .B(n7979), .Z(n7647) );
  AND U9392 ( .A(n7648), .B(n7647), .Z(n7651) );
  NAND U9393 ( .A(n7652), .B(n7651), .Z(n7654) );
  XOR U9394 ( .A(n7652), .B(n7651), .Z(n7985) );
  NANDN U9395 ( .A(n7984), .B(n7985), .Z(n7653) );
  AND U9396 ( .A(n7654), .B(n7653), .Z(n10227) );
  XNOR U9397 ( .A(n10226), .B(n10227), .Z(n10229) );
  NAND U9398 ( .A(a[58]), .B(b[42]), .Z(n10106) );
  NAND U9399 ( .A(a[56]), .B(b[42]), .Z(n7981) );
  AND U9400 ( .A(a[54]), .B(b[42]), .Z(n7969) );
  NAND U9401 ( .A(n7969), .B(n7968), .Z(n7971) );
  AND U9402 ( .A(a[53]), .B(b[42]), .Z(n7964) );
  NAND U9403 ( .A(n7964), .B(n7965), .Z(n7967) );
  AND U9404 ( .A(a[52]), .B(b[42]), .Z(n7960) );
  NAND U9405 ( .A(n7960), .B(n7961), .Z(n7963) );
  AND U9406 ( .A(a[51]), .B(b[42]), .Z(n7956) );
  NAND U9407 ( .A(n7956), .B(n7957), .Z(n7959) );
  NAND U9408 ( .A(a[50]), .B(b[42]), .Z(n7952) );
  XNOR U9409 ( .A(n7664), .B(n7663), .Z(n7953) );
  NANDN U9410 ( .A(n7952), .B(n7953), .Z(n7955) );
  NAND U9411 ( .A(a[49]), .B(b[42]), .Z(n7667) );
  XNOR U9412 ( .A(n7666), .B(n7665), .Z(n7668) );
  NANDN U9413 ( .A(n7667), .B(n7668), .Z(n7951) );
  XOR U9414 ( .A(n7668), .B(n7667), .Z(n8000) );
  XOR U9415 ( .A(n7670), .B(n7669), .Z(n7941) );
  AND U9416 ( .A(a[47]), .B(b[42]), .Z(n7940) );
  NANDN U9417 ( .A(n7941), .B(n7940), .Z(n7943) );
  NAND U9418 ( .A(a[46]), .B(b[42]), .Z(n7936) );
  XNOR U9419 ( .A(n7672), .B(n7671), .Z(n7937) );
  NANDN U9420 ( .A(n7936), .B(n7937), .Z(n7939) );
  XOR U9421 ( .A(n7674), .B(n7673), .Z(n7933) );
  XOR U9422 ( .A(n7676), .B(n7675), .Z(n7923) );
  AND U9423 ( .A(a[43]), .B(b[42]), .Z(n7922) );
  NANDN U9424 ( .A(n7923), .B(n7922), .Z(n7925) );
  XOR U9425 ( .A(n7678), .B(n7677), .Z(n7680) );
  AND U9426 ( .A(a[41]), .B(b[42]), .Z(n7679) );
  NANDN U9427 ( .A(n7680), .B(n7679), .Z(n7915) );
  XOR U9428 ( .A(n7680), .B(n7679), .Z(n8016) );
  NAND U9429 ( .A(a[39]), .B(b[42]), .Z(n7904) );
  XNOR U9430 ( .A(n7682), .B(n7681), .Z(n7905) );
  NANDN U9431 ( .A(n7904), .B(n7905), .Z(n7907) );
  XOR U9432 ( .A(n7684), .B(n7683), .Z(n7686) );
  AND U9433 ( .A(a[37]), .B(b[42]), .Z(n7685) );
  NANDN U9434 ( .A(n7686), .B(n7685), .Z(n7897) );
  XOR U9435 ( .A(n7686), .B(n7685), .Z(n8022) );
  NAND U9436 ( .A(a[36]), .B(b[42]), .Z(n7689) );
  XNOR U9437 ( .A(n7688), .B(n7687), .Z(n7690) );
  NANDN U9438 ( .A(n7689), .B(n7690), .Z(n7895) );
  XOR U9439 ( .A(n7690), .B(n7689), .Z(n8026) );
  XOR U9440 ( .A(n7692), .B(n7691), .Z(n7890) );
  AND U9441 ( .A(a[35]), .B(b[42]), .Z(n7891) );
  NANDN U9442 ( .A(n7890), .B(n7891), .Z(n7893) );
  XOR U9443 ( .A(n7694), .B(n7693), .Z(n7887) );
  AND U9444 ( .A(a[34]), .B(b[42]), .Z(n7886) );
  NANDN U9445 ( .A(n7887), .B(n7886), .Z(n7889) );
  XOR U9446 ( .A(n7696), .B(n7695), .Z(n7697) );
  AND U9447 ( .A(a[32]), .B(b[42]), .Z(n7698) );
  NANDN U9448 ( .A(n7697), .B(n7698), .Z(n7879) );
  XOR U9449 ( .A(n7698), .B(n7697), .Z(n8030) );
  XOR U9450 ( .A(n7700), .B(n7699), .Z(n7875) );
  XOR U9451 ( .A(n7702), .B(n7701), .Z(n7870) );
  AND U9452 ( .A(a[30]), .B(b[42]), .Z(n7871) );
  NANDN U9453 ( .A(n7870), .B(n7871), .Z(n7873) );
  NAND U9454 ( .A(a[28]), .B(b[42]), .Z(n7860) );
  XNOR U9455 ( .A(n7704), .B(n7703), .Z(n7861) );
  NANDN U9456 ( .A(n7860), .B(n7861), .Z(n7863) );
  XOR U9457 ( .A(n7706), .B(n7705), .Z(n7856) );
  AND U9458 ( .A(a[27]), .B(b[42]), .Z(n7857) );
  NANDN U9459 ( .A(n7856), .B(n7857), .Z(n7859) );
  NAND U9460 ( .A(a[24]), .B(b[42]), .Z(n7840) );
  XNOR U9461 ( .A(n7708), .B(n7707), .Z(n7841) );
  NANDN U9462 ( .A(n7840), .B(n7841), .Z(n7843) );
  AND U9463 ( .A(a[20]), .B(b[42]), .Z(n7816) );
  AND U9464 ( .A(a[19]), .B(b[42]), .Z(n7812) );
  XNOR U9465 ( .A(n7710), .B(n7709), .Z(n7813) );
  NANDN U9466 ( .A(n7812), .B(n7813), .Z(n7815) );
  XOR U9467 ( .A(n7712), .B(n7711), .Z(n7802) );
  NAND U9468 ( .A(a[15]), .B(b[42]), .Z(n7792) );
  NANDN U9469 ( .A(n7792), .B(n7793), .Z(n7795) );
  NAND U9470 ( .A(a[14]), .B(b[42]), .Z(n7788) );
  XOR U9471 ( .A(n7716), .B(n7715), .Z(n7789) );
  NANDN U9472 ( .A(n7788), .B(n7789), .Z(n7791) );
  XOR U9473 ( .A(n7718), .B(n7717), .Z(n7778) );
  AND U9474 ( .A(a[11]), .B(b[42]), .Z(n7774) );
  XOR U9475 ( .A(n7720), .B(n7719), .Z(n7762) );
  AND U9476 ( .A(a[8]), .B(b[42]), .Z(n7724) );
  NAND U9477 ( .A(n7724), .B(n7723), .Z(n7761) );
  XOR U9478 ( .A(n7724), .B(n7723), .Z(n8053) );
  NAND U9479 ( .A(a[7]), .B(b[42]), .Z(n7756) );
  XOR U9480 ( .A(n7726), .B(n7725), .Z(n7757) );
  NANDN U9481 ( .A(n7756), .B(n7757), .Z(n7759) );
  NAND U9482 ( .A(a[0]), .B(b[42]), .Z(n8390) );
  AND U9483 ( .A(a[1]), .B(b[43]), .Z(n7729) );
  NANDN U9484 ( .A(n8390), .B(n7729), .Z(n8060) );
  NANDN U9485 ( .A(n8060), .B(n7727), .Z(n7731) );
  AND U9486 ( .A(a[2]), .B(b[42]), .Z(n8066) );
  NANDN U9487 ( .A(n8065), .B(n8066), .Z(n7730) );
  AND U9488 ( .A(n7731), .B(n7730), .Z(n7734) );
  AND U9489 ( .A(a[3]), .B(b[42]), .Z(n7735) );
  NANDN U9490 ( .A(n7734), .B(n7735), .Z(n7737) );
  XOR U9491 ( .A(n7733), .B(n7732), .Z(n8071) );
  NANDN U9492 ( .A(n8071), .B(n8072), .Z(n7736) );
  AND U9493 ( .A(n7737), .B(n7736), .Z(n7740) );
  NANDN U9494 ( .A(n7740), .B(n7741), .Z(n7743) );
  NAND U9495 ( .A(a[4]), .B(b[42]), .Z(n8077) );
  NANDN U9496 ( .A(n8077), .B(n8078), .Z(n7742) );
  AND U9497 ( .A(n7743), .B(n7742), .Z(n7746) );
  XOR U9498 ( .A(n7745), .B(n7744), .Z(n7747) );
  NANDN U9499 ( .A(n7746), .B(n7747), .Z(n7749) );
  AND U9500 ( .A(a[5]), .B(b[42]), .Z(n8084) );
  NAND U9501 ( .A(n8084), .B(n8083), .Z(n7748) );
  AND U9502 ( .A(n7749), .B(n7748), .Z(n7752) );
  NANDN U9503 ( .A(n7752), .B(n7753), .Z(n7755) );
  AND U9504 ( .A(a[6]), .B(b[42]), .Z(n8059) );
  NAND U9505 ( .A(n8059), .B(n8058), .Z(n7754) );
  AND U9506 ( .A(n7755), .B(n7754), .Z(n8054) );
  NANDN U9507 ( .A(n8054), .B(n8055), .Z(n7758) );
  NAND U9508 ( .A(n7759), .B(n7758), .Z(n8052) );
  NAND U9509 ( .A(n8053), .B(n8052), .Z(n7760) );
  AND U9510 ( .A(n7761), .B(n7760), .Z(n7763) );
  NANDN U9511 ( .A(n7762), .B(n7763), .Z(n7765) );
  AND U9512 ( .A(a[9]), .B(b[42]), .Z(n8099) );
  NANDN U9513 ( .A(n8099), .B(n8100), .Z(n7764) );
  AND U9514 ( .A(n7765), .B(n7764), .Z(n7769) );
  NAND U9515 ( .A(n7769), .B(n7768), .Z(n7771) );
  XOR U9516 ( .A(n7769), .B(n7768), .Z(n8051) );
  AND U9517 ( .A(a[10]), .B(b[42]), .Z(n8050) );
  NAND U9518 ( .A(n8051), .B(n8050), .Z(n7770) );
  AND U9519 ( .A(n7771), .B(n7770), .Z(n7775) );
  NANDN U9520 ( .A(n7774), .B(n7775), .Z(n7777) );
  NAND U9521 ( .A(n8049), .B(n8048), .Z(n7776) );
  AND U9522 ( .A(n7777), .B(n7776), .Z(n7779) );
  NANDN U9523 ( .A(n7778), .B(n7779), .Z(n7781) );
  AND U9524 ( .A(a[12]), .B(b[42]), .Z(n8114) );
  NAND U9525 ( .A(n8114), .B(n8113), .Z(n7780) );
  AND U9526 ( .A(n7781), .B(n7780), .Z(n7784) );
  XOR U9527 ( .A(n7783), .B(n7782), .Z(n7785) );
  NANDN U9528 ( .A(n7784), .B(n7785), .Z(n7787) );
  NAND U9529 ( .A(a[13]), .B(b[42]), .Z(n8046) );
  NANDN U9530 ( .A(n8046), .B(n8047), .Z(n7786) );
  AND U9531 ( .A(n7787), .B(n7786), .Z(n8042) );
  NANDN U9532 ( .A(n8042), .B(n8043), .Z(n7790) );
  AND U9533 ( .A(n7791), .B(n7790), .Z(n8127) );
  NANDN U9534 ( .A(n8127), .B(n8128), .Z(n7794) );
  AND U9535 ( .A(n7795), .B(n7794), .Z(n7796) );
  AND U9536 ( .A(a[16]), .B(b[42]), .Z(n7797) );
  NANDN U9537 ( .A(n7796), .B(n7797), .Z(n7801) );
  NAND U9538 ( .A(n8041), .B(n8040), .Z(n7800) );
  AND U9539 ( .A(n7801), .B(n7800), .Z(n7803) );
  NANDN U9540 ( .A(n7802), .B(n7803), .Z(n7805) );
  AND U9541 ( .A(a[17]), .B(b[42]), .Z(n8135) );
  NANDN U9542 ( .A(n8135), .B(n8136), .Z(n7804) );
  AND U9543 ( .A(n7805), .B(n7804), .Z(n7808) );
  NAND U9544 ( .A(n7808), .B(n7809), .Z(n7811) );
  AND U9545 ( .A(a[18]), .B(b[42]), .Z(n8039) );
  XOR U9546 ( .A(n7809), .B(n7808), .Z(n8038) );
  NAND U9547 ( .A(n8039), .B(n8038), .Z(n7810) );
  AND U9548 ( .A(n7811), .B(n7810), .Z(n8146) );
  NAND U9549 ( .A(n8146), .B(n8145), .Z(n7814) );
  NAND U9550 ( .A(n7815), .B(n7814), .Z(n7817) );
  NANDN U9551 ( .A(n7816), .B(n7817), .Z(n7821) );
  NAND U9552 ( .A(n8152), .B(n8151), .Z(n7820) );
  AND U9553 ( .A(n7821), .B(n7820), .Z(n7825) );
  XOR U9554 ( .A(n7823), .B(n7822), .Z(n7824) );
  NAND U9555 ( .A(n7825), .B(n7824), .Z(n7827) );
  AND U9556 ( .A(a[21]), .B(b[42]), .Z(n8158) );
  XOR U9557 ( .A(n7825), .B(n7824), .Z(n8157) );
  NAND U9558 ( .A(n8158), .B(n8157), .Z(n7826) );
  AND U9559 ( .A(n7827), .B(n7826), .Z(n7830) );
  XOR U9560 ( .A(n7829), .B(n7828), .Z(n7831) );
  NANDN U9561 ( .A(n7830), .B(n7831), .Z(n7833) );
  AND U9562 ( .A(a[22]), .B(b[42]), .Z(n8037) );
  NAND U9563 ( .A(n8037), .B(n8036), .Z(n7832) );
  AND U9564 ( .A(n7833), .B(n7832), .Z(n7837) );
  XNOR U9565 ( .A(n7835), .B(n7834), .Z(n7836) );
  NANDN U9566 ( .A(n7837), .B(n7836), .Z(n7839) );
  NAND U9567 ( .A(a[23]), .B(b[42]), .Z(n8167) );
  XNOR U9568 ( .A(n7837), .B(n7836), .Z(n8168) );
  NANDN U9569 ( .A(n8167), .B(n8168), .Z(n7838) );
  AND U9570 ( .A(n7839), .B(n7838), .Z(n8174) );
  XNOR U9571 ( .A(n7841), .B(n7840), .Z(n8173) );
  NANDN U9572 ( .A(n8174), .B(n8173), .Z(n7842) );
  AND U9573 ( .A(n7843), .B(n7842), .Z(n7847) );
  XNOR U9574 ( .A(n7845), .B(n7844), .Z(n7846) );
  NANDN U9575 ( .A(n7847), .B(n7846), .Z(n7849) );
  NAND U9576 ( .A(a[25]), .B(b[42]), .Z(n8179) );
  XNOR U9577 ( .A(n7847), .B(n7846), .Z(n8180) );
  NANDN U9578 ( .A(n8179), .B(n8180), .Z(n7848) );
  AND U9579 ( .A(n7849), .B(n7848), .Z(n7853) );
  XNOR U9580 ( .A(n7851), .B(n7850), .Z(n7852) );
  NANDN U9581 ( .A(n7853), .B(n7852), .Z(n7855) );
  NAND U9582 ( .A(a[26]), .B(b[42]), .Z(n8185) );
  XNOR U9583 ( .A(n7853), .B(n7852), .Z(n8186) );
  NANDN U9584 ( .A(n8185), .B(n8186), .Z(n7854) );
  AND U9585 ( .A(n7855), .B(n7854), .Z(n8192) );
  XNOR U9586 ( .A(n7857), .B(n7856), .Z(n8191) );
  NANDN U9587 ( .A(n8192), .B(n8191), .Z(n7858) );
  AND U9588 ( .A(n7859), .B(n7858), .Z(n8035) );
  XNOR U9589 ( .A(n7861), .B(n7860), .Z(n8034) );
  NANDN U9590 ( .A(n8035), .B(n8034), .Z(n7862) );
  AND U9591 ( .A(n7863), .B(n7862), .Z(n7867) );
  XNOR U9592 ( .A(n7865), .B(n7864), .Z(n7866) );
  NANDN U9593 ( .A(n7867), .B(n7866), .Z(n7869) );
  NAND U9594 ( .A(a[29]), .B(b[42]), .Z(n8201) );
  XNOR U9595 ( .A(n7867), .B(n7866), .Z(n8202) );
  NANDN U9596 ( .A(n8201), .B(n8202), .Z(n7868) );
  AND U9597 ( .A(n7869), .B(n7868), .Z(n8208) );
  XNOR U9598 ( .A(n7871), .B(n7870), .Z(n8207) );
  NANDN U9599 ( .A(n8208), .B(n8207), .Z(n7872) );
  AND U9600 ( .A(n7873), .B(n7872), .Z(n7874) );
  NANDN U9601 ( .A(n7875), .B(n7874), .Z(n7877) );
  XOR U9602 ( .A(n7875), .B(n7874), .Z(n8032) );
  AND U9603 ( .A(a[31]), .B(b[42]), .Z(n8033) );
  OR U9604 ( .A(n8032), .B(n8033), .Z(n7876) );
  AND U9605 ( .A(n7877), .B(n7876), .Z(n8031) );
  NANDN U9606 ( .A(n8030), .B(n8031), .Z(n7878) );
  AND U9607 ( .A(n7879), .B(n7878), .Z(n7883) );
  XNOR U9608 ( .A(n7881), .B(n7880), .Z(n7882) );
  NANDN U9609 ( .A(n7883), .B(n7882), .Z(n7885) );
  NAND U9610 ( .A(a[33]), .B(b[42]), .Z(n8221) );
  XNOR U9611 ( .A(n7883), .B(n7882), .Z(n8222) );
  NANDN U9612 ( .A(n8221), .B(n8222), .Z(n7884) );
  AND U9613 ( .A(n7885), .B(n7884), .Z(n8228) );
  XNOR U9614 ( .A(n7887), .B(n7886), .Z(n8227) );
  NANDN U9615 ( .A(n8228), .B(n8227), .Z(n7888) );
  AND U9616 ( .A(n7889), .B(n7888), .Z(n8029) );
  XNOR U9617 ( .A(n7891), .B(n7890), .Z(n8028) );
  NANDN U9618 ( .A(n8029), .B(n8028), .Z(n7892) );
  AND U9619 ( .A(n7893), .B(n7892), .Z(n8027) );
  OR U9620 ( .A(n8026), .B(n8027), .Z(n7894) );
  AND U9621 ( .A(n7895), .B(n7894), .Z(n8023) );
  OR U9622 ( .A(n8022), .B(n8023), .Z(n7896) );
  AND U9623 ( .A(n7897), .B(n7896), .Z(n7901) );
  XNOR U9624 ( .A(n7899), .B(n7898), .Z(n7900) );
  NANDN U9625 ( .A(n7901), .B(n7900), .Z(n7903) );
  NAND U9626 ( .A(a[38]), .B(b[42]), .Z(n8020) );
  XNOR U9627 ( .A(n7901), .B(n7900), .Z(n8021) );
  NANDN U9628 ( .A(n8020), .B(n8021), .Z(n7902) );
  AND U9629 ( .A(n7903), .B(n7902), .Z(n8248) );
  XNOR U9630 ( .A(n7905), .B(n7904), .Z(n8247) );
  NANDN U9631 ( .A(n8248), .B(n8247), .Z(n7906) );
  AND U9632 ( .A(n7907), .B(n7906), .Z(n7911) );
  XNOR U9633 ( .A(n7909), .B(n7908), .Z(n7910) );
  NANDN U9634 ( .A(n7911), .B(n7910), .Z(n7913) );
  NAND U9635 ( .A(a[40]), .B(b[42]), .Z(n8253) );
  XNOR U9636 ( .A(n7911), .B(n7910), .Z(n8254) );
  NANDN U9637 ( .A(n8253), .B(n8254), .Z(n7912) );
  AND U9638 ( .A(n7913), .B(n7912), .Z(n8017) );
  OR U9639 ( .A(n8016), .B(n8017), .Z(n7914) );
  AND U9640 ( .A(n7915), .B(n7914), .Z(n7919) );
  XNOR U9641 ( .A(n7917), .B(n7916), .Z(n7918) );
  NANDN U9642 ( .A(n7919), .B(n7918), .Z(n7921) );
  NAND U9643 ( .A(a[42]), .B(b[42]), .Z(n8012) );
  XNOR U9644 ( .A(n7919), .B(n7918), .Z(n8013) );
  NANDN U9645 ( .A(n8012), .B(n8013), .Z(n7920) );
  AND U9646 ( .A(n7921), .B(n7920), .Z(n8264) );
  XNOR U9647 ( .A(n7923), .B(n7922), .Z(n8263) );
  NANDN U9648 ( .A(n8264), .B(n8263), .Z(n7924) );
  AND U9649 ( .A(n7925), .B(n7924), .Z(n7929) );
  AND U9650 ( .A(a[44]), .B(b[42]), .Z(n7928) );
  NANDN U9651 ( .A(n7929), .B(n7928), .Z(n7931) );
  XOR U9652 ( .A(n7927), .B(n7926), .Z(n8010) );
  XNOR U9653 ( .A(n7929), .B(n7928), .Z(n8011) );
  NANDN U9654 ( .A(n8010), .B(n8011), .Z(n7930) );
  AND U9655 ( .A(n7931), .B(n7930), .Z(n7932) );
  NANDN U9656 ( .A(n7933), .B(n7932), .Z(n7935) );
  XOR U9657 ( .A(n7933), .B(n7932), .Z(n8008) );
  AND U9658 ( .A(a[45]), .B(b[42]), .Z(n8009) );
  OR U9659 ( .A(n8008), .B(n8009), .Z(n7934) );
  NAND U9660 ( .A(n7935), .B(n7934), .Z(n8006) );
  XNOR U9661 ( .A(n7937), .B(n7936), .Z(n8007) );
  NANDN U9662 ( .A(n8006), .B(n8007), .Z(n7938) );
  AND U9663 ( .A(n7939), .B(n7938), .Z(n8005) );
  XNOR U9664 ( .A(n7941), .B(n7940), .Z(n8004) );
  NANDN U9665 ( .A(n8005), .B(n8004), .Z(n7942) );
  AND U9666 ( .A(n7943), .B(n7942), .Z(n7947) );
  AND U9667 ( .A(a[48]), .B(b[42]), .Z(n7946) );
  NANDN U9668 ( .A(n7947), .B(n7946), .Z(n7949) );
  XOR U9669 ( .A(n7945), .B(n7944), .Z(n8003) );
  XNOR U9670 ( .A(n7947), .B(n7946), .Z(n8002) );
  NANDN U9671 ( .A(n8003), .B(n8002), .Z(n7948) );
  AND U9672 ( .A(n7949), .B(n7948), .Z(n8001) );
  OR U9673 ( .A(n8000), .B(n8001), .Z(n7950) );
  AND U9674 ( .A(n7951), .B(n7950), .Z(n7999) );
  XNOR U9675 ( .A(n7953), .B(n7952), .Z(n7998) );
  NANDN U9676 ( .A(n7999), .B(n7998), .Z(n7954) );
  AND U9677 ( .A(n7955), .B(n7954), .Z(n7997) );
  XOR U9678 ( .A(n7957), .B(n7956), .Z(n7996) );
  NANDN U9679 ( .A(n7997), .B(n7996), .Z(n7958) );
  AND U9680 ( .A(n7959), .B(n7958), .Z(n7994) );
  XOR U9681 ( .A(n7961), .B(n7960), .Z(n7995) );
  NANDN U9682 ( .A(n7994), .B(n7995), .Z(n7962) );
  AND U9683 ( .A(n7963), .B(n7962), .Z(n7992) );
  XOR U9684 ( .A(n7965), .B(n7964), .Z(n7993) );
  NANDN U9685 ( .A(n7992), .B(n7993), .Z(n7966) );
  AND U9686 ( .A(n7967), .B(n7966), .Z(n8307) );
  XOR U9687 ( .A(n7969), .B(n7968), .Z(n8308) );
  NANDN U9688 ( .A(n8307), .B(n8308), .Z(n7970) );
  AND U9689 ( .A(n7971), .B(n7970), .Z(n7972) );
  NAND U9690 ( .A(a[55]), .B(b[42]), .Z(n7973) );
  NAND U9691 ( .A(n7972), .B(n7973), .Z(n7977) );
  XNOR U9692 ( .A(n7973), .B(n7972), .Z(n7990) );
  XNOR U9693 ( .A(n7975), .B(n7974), .Z(n7991) );
  NANDN U9694 ( .A(n7990), .B(n7991), .Z(n7976) );
  NAND U9695 ( .A(n7977), .B(n7976), .Z(n7980) );
  NAND U9696 ( .A(n7981), .B(n7980), .Z(n7983) );
  XOR U9697 ( .A(n7981), .B(n7980), .Z(n8317) );
  NAND U9698 ( .A(n8318), .B(n8317), .Z(n7982) );
  AND U9699 ( .A(n7983), .B(n7982), .Z(n7987) );
  AND U9700 ( .A(a[57]), .B(b[42]), .Z(n7986) );
  NAND U9701 ( .A(n7987), .B(n7986), .Z(n7989) );
  XOR U9702 ( .A(n7987), .B(n7986), .Z(n8323) );
  NAND U9703 ( .A(n8324), .B(n8323), .Z(n7988) );
  AND U9704 ( .A(n7989), .B(n7988), .Z(n10107) );
  XOR U9705 ( .A(n10106), .B(n10107), .Z(n10108) );
  XOR U9706 ( .A(n10109), .B(n10108), .Z(n10235) );
  AND U9707 ( .A(a[58]), .B(b[41]), .Z(n8325) );
  AND U9708 ( .A(a[56]), .B(b[41]), .Z(n8313) );
  NAND U9709 ( .A(n8313), .B(n8314), .Z(n8316) );
  NAND U9710 ( .A(a[54]), .B(b[41]), .Z(n8303) );
  NANDN U9711 ( .A(n8303), .B(n8304), .Z(n8306) );
  AND U9712 ( .A(a[53]), .B(b[41]), .Z(n8300) );
  NAND U9713 ( .A(n8300), .B(n8299), .Z(n8302) );
  XNOR U9714 ( .A(n7997), .B(n7996), .Z(n8297) );
  AND U9715 ( .A(a[52]), .B(b[41]), .Z(n8298) );
  XOR U9716 ( .A(n7999), .B(n7998), .Z(n8293) );
  AND U9717 ( .A(a[50]), .B(b[41]), .Z(n8290) );
  XNOR U9718 ( .A(n8001), .B(n8000), .Z(n8289) );
  NANDN U9719 ( .A(n8290), .B(n8289), .Z(n8292) );
  NAND U9720 ( .A(a[49]), .B(b[41]), .Z(n8285) );
  XNOR U9721 ( .A(n8003), .B(n8002), .Z(n8286) );
  NANDN U9722 ( .A(n8285), .B(n8286), .Z(n8288) );
  NAND U9723 ( .A(a[48]), .B(b[41]), .Z(n8281) );
  XNOR U9724 ( .A(n8005), .B(n8004), .Z(n8282) );
  NANDN U9725 ( .A(n8281), .B(n8282), .Z(n8284) );
  NAND U9726 ( .A(a[47]), .B(b[41]), .Z(n8277) );
  XNOR U9727 ( .A(n8007), .B(n8006), .Z(n8278) );
  NANDN U9728 ( .A(n8277), .B(n8278), .Z(n8280) );
  XOR U9729 ( .A(n8009), .B(n8008), .Z(n8274) );
  AND U9730 ( .A(a[46]), .B(b[41]), .Z(n8273) );
  NANDN U9731 ( .A(n8274), .B(n8273), .Z(n8276) );
  NAND U9732 ( .A(a[45]), .B(b[41]), .Z(n8269) );
  XNOR U9733 ( .A(n8011), .B(n8010), .Z(n8270) );
  NANDN U9734 ( .A(n8269), .B(n8270), .Z(n8272) );
  XOR U9735 ( .A(n8013), .B(n8012), .Z(n8014) );
  AND U9736 ( .A(a[43]), .B(b[41]), .Z(n8015) );
  NANDN U9737 ( .A(n8014), .B(n8015), .Z(n8262) );
  XOR U9738 ( .A(n8015), .B(n8014), .Z(n8343) );
  AND U9739 ( .A(a[42]), .B(b[41]), .Z(n8019) );
  XNOR U9740 ( .A(n8017), .B(n8016), .Z(n8018) );
  NANDN U9741 ( .A(n8019), .B(n8018), .Z(n8260) );
  XNOR U9742 ( .A(n8019), .B(n8018), .Z(n8346) );
  XOR U9743 ( .A(n8021), .B(n8020), .Z(n8243) );
  AND U9744 ( .A(a[38]), .B(b[41]), .Z(n8025) );
  XNOR U9745 ( .A(n8023), .B(n8022), .Z(n8024) );
  NANDN U9746 ( .A(n8025), .B(n8024), .Z(n8242) );
  XOR U9747 ( .A(n8025), .B(n8024), .Z(n8351) );
  XOR U9748 ( .A(n8027), .B(n8026), .Z(n8238) );
  XOR U9749 ( .A(n8029), .B(n8028), .Z(n8233) );
  AND U9750 ( .A(a[36]), .B(b[41]), .Z(n8234) );
  NANDN U9751 ( .A(n8233), .B(n8234), .Z(n8236) );
  XOR U9752 ( .A(n8031), .B(n8030), .Z(n8217) );
  AND U9753 ( .A(a[33]), .B(b[41]), .Z(n8218) );
  NANDN U9754 ( .A(n8217), .B(n8218), .Z(n8220) );
  XOR U9755 ( .A(n8033), .B(n8032), .Z(n8214) );
  NAND U9756 ( .A(a[29]), .B(b[41]), .Z(n8197) );
  XNOR U9757 ( .A(n8035), .B(n8034), .Z(n8198) );
  NANDN U9758 ( .A(n8197), .B(n8198), .Z(n8200) );
  NAND U9759 ( .A(a[23]), .B(b[41]), .Z(n8163) );
  XOR U9760 ( .A(n8037), .B(n8036), .Z(n8164) );
  NANDN U9761 ( .A(n8163), .B(n8164), .Z(n8166) );
  NAND U9762 ( .A(a[19]), .B(b[41]), .Z(n8141) );
  XOR U9763 ( .A(n8039), .B(n8038), .Z(n8142) );
  NANDN U9764 ( .A(n8141), .B(n8142), .Z(n8144) );
  XOR U9765 ( .A(n8041), .B(n8040), .Z(n8131) );
  NAND U9766 ( .A(a[15]), .B(b[41]), .Z(n8044) );
  NANDN U9767 ( .A(n8044), .B(n8045), .Z(n8124) );
  NAND U9768 ( .A(a[14]), .B(b[41]), .Z(n8119) );
  NANDN U9769 ( .A(n8119), .B(n8120), .Z(n8122) );
  XOR U9770 ( .A(n8049), .B(n8048), .Z(n8109) );
  AND U9771 ( .A(a[11]), .B(b[41]), .Z(n8105) );
  XNOR U9772 ( .A(n8051), .B(n8050), .Z(n8106) );
  NANDN U9773 ( .A(n8105), .B(n8106), .Z(n8108) );
  XOR U9774 ( .A(n8053), .B(n8052), .Z(n8095) );
  NAND U9775 ( .A(a[8]), .B(b[41]), .Z(n8056) );
  NANDN U9776 ( .A(n8056), .B(n8057), .Z(n8094) );
  NAND U9777 ( .A(a[7]), .B(b[41]), .Z(n8089) );
  XOR U9778 ( .A(n8059), .B(n8058), .Z(n8090) );
  NANDN U9779 ( .A(n8089), .B(n8090), .Z(n8092) );
  NAND U9780 ( .A(a[0]), .B(b[41]), .Z(n8751) );
  AND U9781 ( .A(a[1]), .B(b[42]), .Z(n8062) );
  NANDN U9782 ( .A(n8751), .B(n8062), .Z(n8389) );
  NANDN U9783 ( .A(n8389), .B(n8060), .Z(n8064) );
  AND U9784 ( .A(a[2]), .B(b[41]), .Z(n8395) );
  NANDN U9785 ( .A(n8394), .B(n8395), .Z(n8063) );
  AND U9786 ( .A(n8064), .B(n8063), .Z(n8067) );
  AND U9787 ( .A(a[3]), .B(b[41]), .Z(n8068) );
  NANDN U9788 ( .A(n8067), .B(n8068), .Z(n8070) );
  XOR U9789 ( .A(n8066), .B(n8065), .Z(n8400) );
  NANDN U9790 ( .A(n8400), .B(n8401), .Z(n8069) );
  AND U9791 ( .A(n8070), .B(n8069), .Z(n8073) );
  NANDN U9792 ( .A(n8073), .B(n8074), .Z(n8076) );
  AND U9793 ( .A(a[4]), .B(b[41]), .Z(n8407) );
  NAND U9794 ( .A(n8407), .B(n8406), .Z(n8075) );
  AND U9795 ( .A(n8076), .B(n8075), .Z(n8079) );
  NANDN U9796 ( .A(n8079), .B(n8080), .Z(n8082) );
  AND U9797 ( .A(a[5]), .B(b[41]), .Z(n8413) );
  NAND U9798 ( .A(n8413), .B(n8412), .Z(n8081) );
  AND U9799 ( .A(n8082), .B(n8081), .Z(n8085) );
  XOR U9800 ( .A(n8084), .B(n8083), .Z(n8086) );
  NANDN U9801 ( .A(n8085), .B(n8086), .Z(n8088) );
  NAND U9802 ( .A(a[6]), .B(b[41]), .Z(n8387) );
  NANDN U9803 ( .A(n8387), .B(n8388), .Z(n8087) );
  AND U9804 ( .A(n8088), .B(n8087), .Z(n8385) );
  NANDN U9805 ( .A(n8385), .B(n8386), .Z(n8091) );
  NAND U9806 ( .A(n8092), .B(n8091), .Z(n8383) );
  NAND U9807 ( .A(n8384), .B(n8383), .Z(n8093) );
  AND U9808 ( .A(n8094), .B(n8093), .Z(n8096) );
  NANDN U9809 ( .A(n8095), .B(n8096), .Z(n8098) );
  AND U9810 ( .A(a[9]), .B(b[41]), .Z(n8430) );
  NANDN U9811 ( .A(n8430), .B(n8431), .Z(n8097) );
  AND U9812 ( .A(n8098), .B(n8097), .Z(n8101) );
  NANDN U9813 ( .A(n8101), .B(n8102), .Z(n8104) );
  AND U9814 ( .A(a[10]), .B(b[41]), .Z(n8438) );
  NANDN U9815 ( .A(n8438), .B(n8439), .Z(n8103) );
  AND U9816 ( .A(n8104), .B(n8103), .Z(n8442) );
  NANDN U9817 ( .A(n8442), .B(n8443), .Z(n8107) );
  AND U9818 ( .A(n8108), .B(n8107), .Z(n8110) );
  NANDN U9819 ( .A(n8109), .B(n8110), .Z(n8112) );
  NAND U9820 ( .A(a[12]), .B(b[41]), .Z(n8448) );
  NANDN U9821 ( .A(n8448), .B(n8449), .Z(n8111) );
  AND U9822 ( .A(n8112), .B(n8111), .Z(n8115) );
  XOR U9823 ( .A(n8114), .B(n8113), .Z(n8116) );
  NANDN U9824 ( .A(n8115), .B(n8116), .Z(n8118) );
  NAND U9825 ( .A(a[13]), .B(b[41]), .Z(n8381) );
  NANDN U9826 ( .A(n8381), .B(n8382), .Z(n8117) );
  AND U9827 ( .A(n8118), .B(n8117), .Z(n8379) );
  NANDN U9828 ( .A(n8379), .B(n8380), .Z(n8121) );
  NAND U9829 ( .A(n8122), .B(n8121), .Z(n8462) );
  NAND U9830 ( .A(n8463), .B(n8462), .Z(n8123) );
  AND U9831 ( .A(n8124), .B(n8123), .Z(n8125) );
  AND U9832 ( .A(a[16]), .B(b[41]), .Z(n8126) );
  NANDN U9833 ( .A(n8125), .B(n8126), .Z(n8130) );
  NAND U9834 ( .A(n8378), .B(n8377), .Z(n8129) );
  AND U9835 ( .A(n8130), .B(n8129), .Z(n8132) );
  NANDN U9836 ( .A(n8131), .B(n8132), .Z(n8134) );
  AND U9837 ( .A(a[17]), .B(b[41]), .Z(n8472) );
  NANDN U9838 ( .A(n8472), .B(n8473), .Z(n8133) );
  AND U9839 ( .A(n8134), .B(n8133), .Z(n8137) );
  NANDN U9840 ( .A(n8137), .B(n8138), .Z(n8140) );
  AND U9841 ( .A(a[18]), .B(b[41]), .Z(n8375) );
  NANDN U9842 ( .A(n8375), .B(n8376), .Z(n8139) );
  AND U9843 ( .A(n8140), .B(n8139), .Z(n8485) );
  NAND U9844 ( .A(n8485), .B(n8484), .Z(n8143) );
  AND U9845 ( .A(n8144), .B(n8143), .Z(n8147) );
  AND U9846 ( .A(a[20]), .B(b[41]), .Z(n8148) );
  NANDN U9847 ( .A(n8147), .B(n8148), .Z(n8150) );
  XOR U9848 ( .A(n8146), .B(n8145), .Z(n8488) );
  NANDN U9849 ( .A(n8488), .B(n8489), .Z(n8149) );
  AND U9850 ( .A(n8150), .B(n8149), .Z(n8154) );
  XOR U9851 ( .A(n8152), .B(n8151), .Z(n8153) );
  NAND U9852 ( .A(n8154), .B(n8153), .Z(n8156) );
  AND U9853 ( .A(a[21]), .B(b[41]), .Z(n8373) );
  XOR U9854 ( .A(n8154), .B(n8153), .Z(n8374) );
  NANDN U9855 ( .A(n8373), .B(n8374), .Z(n8155) );
  NAND U9856 ( .A(n8156), .B(n8155), .Z(n8159) );
  XOR U9857 ( .A(n8158), .B(n8157), .Z(n8160) );
  NANDN U9858 ( .A(n8159), .B(n8160), .Z(n8162) );
  NAND U9859 ( .A(a[22]), .B(b[41]), .Z(n8500) );
  NANDN U9860 ( .A(n8500), .B(n8501), .Z(n8161) );
  AND U9861 ( .A(n8162), .B(n8161), .Z(n8371) );
  NANDN U9862 ( .A(n8371), .B(n8372), .Z(n8165) );
  AND U9863 ( .A(n8166), .B(n8165), .Z(n8170) );
  XNOR U9864 ( .A(n8168), .B(n8167), .Z(n8169) );
  NANDN U9865 ( .A(n8170), .B(n8169), .Z(n8172) );
  NAND U9866 ( .A(a[24]), .B(b[41]), .Z(n8508) );
  XNOR U9867 ( .A(n8170), .B(n8169), .Z(n8509) );
  NANDN U9868 ( .A(n8508), .B(n8509), .Z(n8171) );
  AND U9869 ( .A(n8172), .B(n8171), .Z(n8176) );
  AND U9870 ( .A(a[25]), .B(b[41]), .Z(n8175) );
  NANDN U9871 ( .A(n8176), .B(n8175), .Z(n8178) );
  XOR U9872 ( .A(n8174), .B(n8173), .Z(n8514) );
  XNOR U9873 ( .A(n8176), .B(n8175), .Z(n8515) );
  NANDN U9874 ( .A(n8514), .B(n8515), .Z(n8177) );
  AND U9875 ( .A(n8178), .B(n8177), .Z(n8182) );
  XNOR U9876 ( .A(n8180), .B(n8179), .Z(n8181) );
  NANDN U9877 ( .A(n8182), .B(n8181), .Z(n8184) );
  NAND U9878 ( .A(a[26]), .B(b[41]), .Z(n8369) );
  XNOR U9879 ( .A(n8182), .B(n8181), .Z(n8370) );
  NANDN U9880 ( .A(n8369), .B(n8370), .Z(n8183) );
  AND U9881 ( .A(n8184), .B(n8183), .Z(n8188) );
  XNOR U9882 ( .A(n8186), .B(n8185), .Z(n8187) );
  NANDN U9883 ( .A(n8188), .B(n8187), .Z(n8190) );
  NAND U9884 ( .A(a[27]), .B(b[41]), .Z(n8524) );
  XNOR U9885 ( .A(n8188), .B(n8187), .Z(n8525) );
  NANDN U9886 ( .A(n8524), .B(n8525), .Z(n8189) );
  AND U9887 ( .A(n8190), .B(n8189), .Z(n8194) );
  XNOR U9888 ( .A(n8192), .B(n8191), .Z(n8193) );
  NANDN U9889 ( .A(n8194), .B(n8193), .Z(n8196) );
  NAND U9890 ( .A(a[28]), .B(b[41]), .Z(n8367) );
  XNOR U9891 ( .A(n8194), .B(n8193), .Z(n8368) );
  NANDN U9892 ( .A(n8367), .B(n8368), .Z(n8195) );
  AND U9893 ( .A(n8196), .B(n8195), .Z(n8535) );
  XNOR U9894 ( .A(n8198), .B(n8197), .Z(n8534) );
  NANDN U9895 ( .A(n8535), .B(n8534), .Z(n8199) );
  AND U9896 ( .A(n8200), .B(n8199), .Z(n8204) );
  XNOR U9897 ( .A(n8202), .B(n8201), .Z(n8203) );
  NANDN U9898 ( .A(n8204), .B(n8203), .Z(n8206) );
  NAND U9899 ( .A(a[30]), .B(b[41]), .Z(n8365) );
  XNOR U9900 ( .A(n8204), .B(n8203), .Z(n8366) );
  NANDN U9901 ( .A(n8365), .B(n8366), .Z(n8205) );
  AND U9902 ( .A(n8206), .B(n8205), .Z(n8210) );
  XNOR U9903 ( .A(n8208), .B(n8207), .Z(n8209) );
  NANDN U9904 ( .A(n8210), .B(n8209), .Z(n8212) );
  NAND U9905 ( .A(a[31]), .B(b[41]), .Z(n8544) );
  XNOR U9906 ( .A(n8210), .B(n8209), .Z(n8545) );
  NANDN U9907 ( .A(n8544), .B(n8545), .Z(n8211) );
  NAND U9908 ( .A(n8212), .B(n8211), .Z(n8213) );
  NANDN U9909 ( .A(n8214), .B(n8213), .Z(n8216) );
  NAND U9910 ( .A(a[32]), .B(b[41]), .Z(n8363) );
  XNOR U9911 ( .A(n8214), .B(n8213), .Z(n8364) );
  NANDN U9912 ( .A(n8363), .B(n8364), .Z(n8215) );
  AND U9913 ( .A(n8216), .B(n8215), .Z(n8362) );
  XNOR U9914 ( .A(n8218), .B(n8217), .Z(n8361) );
  NANDN U9915 ( .A(n8362), .B(n8361), .Z(n8219) );
  AND U9916 ( .A(n8220), .B(n8219), .Z(n8224) );
  XNOR U9917 ( .A(n8222), .B(n8221), .Z(n8223) );
  NANDN U9918 ( .A(n8224), .B(n8223), .Z(n8226) );
  NAND U9919 ( .A(a[34]), .B(b[41]), .Z(n8558) );
  XNOR U9920 ( .A(n8224), .B(n8223), .Z(n8559) );
  NANDN U9921 ( .A(n8558), .B(n8559), .Z(n8225) );
  AND U9922 ( .A(n8226), .B(n8225), .Z(n8230) );
  XNOR U9923 ( .A(n8228), .B(n8227), .Z(n8229) );
  NANDN U9924 ( .A(n8230), .B(n8229), .Z(n8232) );
  XNOR U9925 ( .A(n8230), .B(n8229), .Z(n8360) );
  AND U9926 ( .A(a[35]), .B(b[41]), .Z(n8359) );
  NAND U9927 ( .A(n8360), .B(n8359), .Z(n8231) );
  AND U9928 ( .A(n8232), .B(n8231), .Z(n8358) );
  XNOR U9929 ( .A(n8234), .B(n8233), .Z(n8357) );
  NANDN U9930 ( .A(n8358), .B(n8357), .Z(n8235) );
  AND U9931 ( .A(n8236), .B(n8235), .Z(n8237) );
  NANDN U9932 ( .A(n8238), .B(n8237), .Z(n8240) );
  XOR U9933 ( .A(n8238), .B(n8237), .Z(n8353) );
  AND U9934 ( .A(a[37]), .B(b[41]), .Z(n8354) );
  OR U9935 ( .A(n8353), .B(n8354), .Z(n8239) );
  AND U9936 ( .A(n8240), .B(n8239), .Z(n8352) );
  OR U9937 ( .A(n8351), .B(n8352), .Z(n8241) );
  AND U9938 ( .A(n8242), .B(n8241), .Z(n8244) );
  NANDN U9939 ( .A(n8243), .B(n8244), .Z(n8246) );
  NAND U9940 ( .A(a[39]), .B(b[41]), .Z(n8349) );
  XNOR U9941 ( .A(n8244), .B(n8243), .Z(n8350) );
  NANDN U9942 ( .A(n8349), .B(n8350), .Z(n8245) );
  AND U9943 ( .A(n8246), .B(n8245), .Z(n8250) );
  XNOR U9944 ( .A(n8248), .B(n8247), .Z(n8249) );
  NANDN U9945 ( .A(n8250), .B(n8249), .Z(n8252) );
  NAND U9946 ( .A(a[40]), .B(b[41]), .Z(n8582) );
  XNOR U9947 ( .A(n8250), .B(n8249), .Z(n8583) );
  NANDN U9948 ( .A(n8582), .B(n8583), .Z(n8251) );
  AND U9949 ( .A(n8252), .B(n8251), .Z(n8256) );
  XNOR U9950 ( .A(n8254), .B(n8253), .Z(n8255) );
  NANDN U9951 ( .A(n8256), .B(n8255), .Z(n8258) );
  NAND U9952 ( .A(a[41]), .B(b[41]), .Z(n8347) );
  XNOR U9953 ( .A(n8256), .B(n8255), .Z(n8348) );
  NANDN U9954 ( .A(n8347), .B(n8348), .Z(n8257) );
  AND U9955 ( .A(n8258), .B(n8257), .Z(n8345) );
  NAND U9956 ( .A(n8346), .B(n8345), .Z(n8259) );
  AND U9957 ( .A(n8260), .B(n8259), .Z(n8344) );
  NANDN U9958 ( .A(n8343), .B(n8344), .Z(n8261) );
  AND U9959 ( .A(n8262), .B(n8261), .Z(n8266) );
  XNOR U9960 ( .A(n8264), .B(n8263), .Z(n8265) );
  NANDN U9961 ( .A(n8266), .B(n8265), .Z(n8268) );
  NAND U9962 ( .A(a[44]), .B(b[41]), .Z(n8600) );
  XNOR U9963 ( .A(n8266), .B(n8265), .Z(n8601) );
  NANDN U9964 ( .A(n8600), .B(n8601), .Z(n8267) );
  AND U9965 ( .A(n8268), .B(n8267), .Z(n8607) );
  XNOR U9966 ( .A(n8270), .B(n8269), .Z(n8606) );
  NANDN U9967 ( .A(n8607), .B(n8606), .Z(n8271) );
  AND U9968 ( .A(n8272), .B(n8271), .Z(n8342) );
  XNOR U9969 ( .A(n8274), .B(n8273), .Z(n8341) );
  NANDN U9970 ( .A(n8342), .B(n8341), .Z(n8275) );
  AND U9971 ( .A(n8276), .B(n8275), .Z(n8340) );
  XNOR U9972 ( .A(n8278), .B(n8277), .Z(n8339) );
  NANDN U9973 ( .A(n8340), .B(n8339), .Z(n8279) );
  AND U9974 ( .A(n8280), .B(n8279), .Z(n8621) );
  XNOR U9975 ( .A(n8282), .B(n8281), .Z(n8620) );
  NANDN U9976 ( .A(n8621), .B(n8620), .Z(n8283) );
  AND U9977 ( .A(n8284), .B(n8283), .Z(n8338) );
  XNOR U9978 ( .A(n8286), .B(n8285), .Z(n8337) );
  NANDN U9979 ( .A(n8338), .B(n8337), .Z(n8287) );
  AND U9980 ( .A(n8288), .B(n8287), .Z(n8631) );
  XNOR U9981 ( .A(n8290), .B(n8289), .Z(n8630) );
  NAND U9982 ( .A(n8631), .B(n8630), .Z(n8291) );
  AND U9983 ( .A(n8292), .B(n8291), .Z(n8294) );
  NANDN U9984 ( .A(n8293), .B(n8294), .Z(n8296) );
  NAND U9985 ( .A(a[51]), .B(b[41]), .Z(n8636) );
  XNOR U9986 ( .A(n8294), .B(n8293), .Z(n8637) );
  NANDN U9987 ( .A(n8636), .B(n8637), .Z(n8295) );
  AND U9988 ( .A(n8296), .B(n8295), .Z(n8334) );
  XOR U9989 ( .A(n8298), .B(n8297), .Z(n8333) );
  XOR U9990 ( .A(n8300), .B(n8299), .Z(n8331) );
  NANDN U9991 ( .A(n8332), .B(n8331), .Z(n8301) );
  AND U9992 ( .A(n8302), .B(n8301), .Z(n8329) );
  NANDN U9993 ( .A(n8329), .B(n8330), .Z(n8305) );
  AND U9994 ( .A(n8306), .B(n8305), .Z(n8309) );
  AND U9995 ( .A(a[55]), .B(b[41]), .Z(n8310) );
  NANDN U9996 ( .A(n8309), .B(n8310), .Z(n8312) );
  NAND U9997 ( .A(n8653), .B(n8652), .Z(n8311) );
  AND U9998 ( .A(n8312), .B(n8311), .Z(n8658) );
  XOR U9999 ( .A(n8314), .B(n8313), .Z(n8659) );
  NANDN U10000 ( .A(n8658), .B(n8659), .Z(n8315) );
  AND U10001 ( .A(n8316), .B(n8315), .Z(n8319) );
  AND U10002 ( .A(a[57]), .B(b[41]), .Z(n8320) );
  NANDN U10003 ( .A(n8319), .B(n8320), .Z(n8322) );
  XOR U10004 ( .A(n8318), .B(n8317), .Z(n8664) );
  NANDN U10005 ( .A(n8664), .B(n8665), .Z(n8321) );
  AND U10006 ( .A(n8322), .B(n8321), .Z(n8326) );
  NANDN U10007 ( .A(n8325), .B(n8326), .Z(n8328) );
  XOR U10008 ( .A(n8324), .B(n8323), .Z(n8670) );
  NANDN U10009 ( .A(n8670), .B(n8671), .Z(n8327) );
  AND U10010 ( .A(n8328), .B(n8327), .Z(n10232) );
  NAND U10011 ( .A(a[59]), .B(b[41]), .Z(n10233) );
  AND U10012 ( .A(a[60]), .B(b[40]), .Z(n10239) );
  AND U10013 ( .A(a[59]), .B(b[40]), .Z(n8672) );
  NAND U10014 ( .A(a[54]), .B(b[40]), .Z(n8644) );
  XNOR U10015 ( .A(n8332), .B(n8331), .Z(n8645) );
  NANDN U10016 ( .A(n8644), .B(n8645), .Z(n8647) );
  NAND U10017 ( .A(a[53]), .B(b[40]), .Z(n8335) );
  XNOR U10018 ( .A(n8334), .B(n8333), .Z(n8336) );
  NANDN U10019 ( .A(n8335), .B(n8336), .Z(n8643) );
  XOR U10020 ( .A(n8336), .B(n8335), .Z(n8684) );
  XOR U10021 ( .A(n8338), .B(n8337), .Z(n8626) );
  AND U10022 ( .A(a[50]), .B(b[40]), .Z(n8627) );
  NANDN U10023 ( .A(n8626), .B(n8627), .Z(n8629) );
  NAND U10024 ( .A(a[48]), .B(b[40]), .Z(n8616) );
  XNOR U10025 ( .A(n8340), .B(n8339), .Z(n8617) );
  NANDN U10026 ( .A(n8616), .B(n8617), .Z(n8619) );
  XOR U10027 ( .A(n8342), .B(n8341), .Z(n8612) );
  AND U10028 ( .A(a[47]), .B(b[40]), .Z(n8613) );
  NANDN U10029 ( .A(n8612), .B(n8613), .Z(n8615) );
  XOR U10030 ( .A(n8344), .B(n8343), .Z(n8596) );
  AND U10031 ( .A(a[44]), .B(b[40]), .Z(n8597) );
  NANDN U10032 ( .A(n8596), .B(n8597), .Z(n8599) );
  XOR U10033 ( .A(n8346), .B(n8345), .Z(n8593) );
  XOR U10034 ( .A(n8348), .B(n8347), .Z(n8588) );
  AND U10035 ( .A(a[42]), .B(b[40]), .Z(n8589) );
  NANDN U10036 ( .A(n8588), .B(n8589), .Z(n8591) );
  XOR U10037 ( .A(n8350), .B(n8349), .Z(n8578) );
  AND U10038 ( .A(a[40]), .B(b[40]), .Z(n8579) );
  NANDN U10039 ( .A(n8578), .B(n8579), .Z(n8581) );
  XOR U10040 ( .A(n8352), .B(n8351), .Z(n8575) );
  XOR U10041 ( .A(n8354), .B(n8353), .Z(n8356) );
  AND U10042 ( .A(a[38]), .B(b[40]), .Z(n8355) );
  NANDN U10043 ( .A(n8356), .B(n8355), .Z(n8573) );
  XOR U10044 ( .A(n8356), .B(n8355), .Z(n8710) );
  XOR U10045 ( .A(n8358), .B(n8357), .Z(n8568) );
  AND U10046 ( .A(a[37]), .B(b[40]), .Z(n8569) );
  NANDN U10047 ( .A(n8568), .B(n8569), .Z(n8571) );
  XOR U10048 ( .A(n8360), .B(n8359), .Z(n8565) );
  XOR U10049 ( .A(n8362), .B(n8361), .Z(n8554) );
  AND U10050 ( .A(a[34]), .B(b[40]), .Z(n8555) );
  NANDN U10051 ( .A(n8554), .B(n8555), .Z(n8557) );
  NAND U10052 ( .A(a[33]), .B(b[40]), .Z(n8550) );
  XNOR U10053 ( .A(n8364), .B(n8363), .Z(n8551) );
  NANDN U10054 ( .A(n8550), .B(n8551), .Z(n8553) );
  XOR U10055 ( .A(n8366), .B(n8365), .Z(n8540) );
  AND U10056 ( .A(a[31]), .B(b[40]), .Z(n8541) );
  NANDN U10057 ( .A(n8540), .B(n8541), .Z(n8543) );
  XOR U10058 ( .A(n8368), .B(n8367), .Z(n8530) );
  AND U10059 ( .A(a[29]), .B(b[40]), .Z(n8531) );
  NANDN U10060 ( .A(n8530), .B(n8531), .Z(n8533) );
  XOR U10061 ( .A(n8370), .B(n8369), .Z(n8520) );
  AND U10062 ( .A(a[27]), .B(b[40]), .Z(n8521) );
  NANDN U10063 ( .A(n8520), .B(n8521), .Z(n8523) );
  AND U10064 ( .A(a[24]), .B(b[40]), .Z(n8505) );
  NAND U10065 ( .A(n8505), .B(n8504), .Z(n8507) );
  AND U10066 ( .A(a[22]), .B(b[40]), .Z(n8494) );
  NAND U10067 ( .A(n8494), .B(n8495), .Z(n8497) );
  NAND U10068 ( .A(a[20]), .B(b[40]), .Z(n8482) );
  AND U10069 ( .A(a[19]), .B(b[40]), .Z(n8478) );
  NANDN U10070 ( .A(n8478), .B(n8479), .Z(n8481) );
  XOR U10071 ( .A(n8378), .B(n8377), .Z(n8468) );
  AND U10072 ( .A(a[16]), .B(b[40]), .Z(n8464) );
  AND U10073 ( .A(a[15]), .B(b[40]), .Z(n8459) );
  NAND U10074 ( .A(n8459), .B(n8458), .Z(n8461) );
  NAND U10075 ( .A(a[14]), .B(b[40]), .Z(n8454) );
  NANDN U10076 ( .A(n8454), .B(n8455), .Z(n8457) );
  AND U10077 ( .A(a[11]), .B(b[40]), .Z(n8436) );
  XOR U10078 ( .A(n8384), .B(n8383), .Z(n8426) );
  NAND U10079 ( .A(a[8]), .B(b[40]), .Z(n8422) );
  NANDN U10080 ( .A(n8422), .B(n8423), .Z(n8425) );
  AND U10081 ( .A(a[7]), .B(b[40]), .Z(n8419) );
  NAND U10082 ( .A(n8419), .B(n8418), .Z(n8421) );
  NAND U10083 ( .A(a[0]), .B(b[40]), .Z(n9051) );
  AND U10084 ( .A(a[1]), .B(b[41]), .Z(n8391) );
  NANDN U10085 ( .A(n9051), .B(n8391), .Z(n8750) );
  NANDN U10086 ( .A(n8750), .B(n8389), .Z(n8393) );
  AND U10087 ( .A(a[2]), .B(b[40]), .Z(n8756) );
  NANDN U10088 ( .A(n8755), .B(n8756), .Z(n8392) );
  AND U10089 ( .A(n8393), .B(n8392), .Z(n8396) );
  AND U10090 ( .A(a[3]), .B(b[40]), .Z(n8397) );
  NANDN U10091 ( .A(n8396), .B(n8397), .Z(n8399) );
  XOR U10092 ( .A(n8395), .B(n8394), .Z(n8761) );
  NANDN U10093 ( .A(n8761), .B(n8762), .Z(n8398) );
  AND U10094 ( .A(n8399), .B(n8398), .Z(n8402) );
  NANDN U10095 ( .A(n8402), .B(n8403), .Z(n8405) );
  AND U10096 ( .A(a[4]), .B(b[40]), .Z(n8749) );
  NAND U10097 ( .A(n8749), .B(n8748), .Z(n8404) );
  AND U10098 ( .A(n8405), .B(n8404), .Z(n8408) );
  XOR U10099 ( .A(n8407), .B(n8406), .Z(n8409) );
  NANDN U10100 ( .A(n8408), .B(n8409), .Z(n8411) );
  AND U10101 ( .A(a[5]), .B(b[40]), .Z(n8772) );
  NAND U10102 ( .A(n8772), .B(n8771), .Z(n8410) );
  AND U10103 ( .A(n8411), .B(n8410), .Z(n8414) );
  XOR U10104 ( .A(n8413), .B(n8412), .Z(n8415) );
  NANDN U10105 ( .A(n8414), .B(n8415), .Z(n8417) );
  NAND U10106 ( .A(a[6]), .B(b[40]), .Z(n8746) );
  NANDN U10107 ( .A(n8746), .B(n8747), .Z(n8416) );
  AND U10108 ( .A(n8417), .B(n8416), .Z(n8744) );
  XOR U10109 ( .A(n8419), .B(n8418), .Z(n8745) );
  NANDN U10110 ( .A(n8744), .B(n8745), .Z(n8420) );
  AND U10111 ( .A(n8421), .B(n8420), .Z(n8785) );
  NANDN U10112 ( .A(n8785), .B(n8786), .Z(n8424) );
  AND U10113 ( .A(n8425), .B(n8424), .Z(n8427) );
  NANDN U10114 ( .A(n8426), .B(n8427), .Z(n8429) );
  AND U10115 ( .A(a[9]), .B(b[40]), .Z(n8791) );
  NANDN U10116 ( .A(n8791), .B(n8792), .Z(n8428) );
  AND U10117 ( .A(n8429), .B(n8428), .Z(n8433) );
  NAND U10118 ( .A(n8433), .B(n8432), .Z(n8435) );
  XOR U10119 ( .A(n8433), .B(n8432), .Z(n8743) );
  AND U10120 ( .A(a[10]), .B(b[40]), .Z(n8742) );
  NAND U10121 ( .A(n8743), .B(n8742), .Z(n8434) );
  AND U10122 ( .A(n8435), .B(n8434), .Z(n8437) );
  NANDN U10123 ( .A(n8436), .B(n8437), .Z(n8441) );
  NAND U10124 ( .A(n8741), .B(n8740), .Z(n8440) );
  AND U10125 ( .A(n8441), .B(n8440), .Z(n8445) );
  NAND U10126 ( .A(n8445), .B(n8444), .Z(n8447) );
  AND U10127 ( .A(a[12]), .B(b[40]), .Z(n8806) );
  XOR U10128 ( .A(n8445), .B(n8444), .Z(n8805) );
  NAND U10129 ( .A(n8806), .B(n8805), .Z(n8446) );
  AND U10130 ( .A(n8447), .B(n8446), .Z(n8450) );
  NANDN U10131 ( .A(n8450), .B(n8451), .Z(n8453) );
  NAND U10132 ( .A(a[13]), .B(b[40]), .Z(n8738) );
  NANDN U10133 ( .A(n8738), .B(n8739), .Z(n8452) );
  AND U10134 ( .A(n8453), .B(n8452), .Z(n8815) );
  NANDN U10135 ( .A(n8815), .B(n8816), .Z(n8456) );
  AND U10136 ( .A(n8457), .B(n8456), .Z(n8736) );
  XOR U10137 ( .A(n8459), .B(n8458), .Z(n8737) );
  NANDN U10138 ( .A(n8736), .B(n8737), .Z(n8460) );
  AND U10139 ( .A(n8461), .B(n8460), .Z(n8465) );
  NANDN U10140 ( .A(n8464), .B(n8465), .Z(n8467) );
  XOR U10141 ( .A(n8463), .B(n8462), .Z(n8825) );
  NANDN U10142 ( .A(n8825), .B(n8826), .Z(n8466) );
  NAND U10143 ( .A(n8467), .B(n8466), .Z(n8469) );
  NANDN U10144 ( .A(n8468), .B(n8469), .Z(n8471) );
  AND U10145 ( .A(a[17]), .B(b[40]), .Z(n8831) );
  NANDN U10146 ( .A(n8831), .B(n8832), .Z(n8470) );
  AND U10147 ( .A(n8471), .B(n8470), .Z(n8474) );
  NAND U10148 ( .A(n8474), .B(n8475), .Z(n8477) );
  XOR U10149 ( .A(n8475), .B(n8474), .Z(n8735) );
  AND U10150 ( .A(a[18]), .B(b[40]), .Z(n8734) );
  NAND U10151 ( .A(n8735), .B(n8734), .Z(n8476) );
  AND U10152 ( .A(n8477), .B(n8476), .Z(n8733) );
  NAND U10153 ( .A(n8733), .B(n8732), .Z(n8480) );
  AND U10154 ( .A(n8481), .B(n8480), .Z(n8483) );
  NANDN U10155 ( .A(n8482), .B(n8483), .Z(n8487) );
  XOR U10156 ( .A(n8485), .B(n8484), .Z(n8730) );
  NAND U10157 ( .A(n8731), .B(n8730), .Z(n8486) );
  AND U10158 ( .A(n8487), .B(n8486), .Z(n8490) );
  NAND U10159 ( .A(n8490), .B(n8491), .Z(n8493) );
  AND U10160 ( .A(a[21]), .B(b[40]), .Z(n8726) );
  XOR U10161 ( .A(n8491), .B(n8490), .Z(n8727) );
  NANDN U10162 ( .A(n8726), .B(n8727), .Z(n8492) );
  NAND U10163 ( .A(n8493), .B(n8492), .Z(n8724) );
  XOR U10164 ( .A(n8495), .B(n8494), .Z(n8725) );
  NANDN U10165 ( .A(n8724), .B(n8725), .Z(n8496) );
  AND U10166 ( .A(n8497), .B(n8496), .Z(n8498) );
  AND U10167 ( .A(a[23]), .B(b[40]), .Z(n8499) );
  NANDN U10168 ( .A(n8498), .B(n8499), .Z(n8503) );
  NAND U10169 ( .A(n8723), .B(n8722), .Z(n8502) );
  AND U10170 ( .A(n8503), .B(n8502), .Z(n8720) );
  XOR U10171 ( .A(n8505), .B(n8504), .Z(n8721) );
  NANDN U10172 ( .A(n8720), .B(n8721), .Z(n8506) );
  AND U10173 ( .A(n8507), .B(n8506), .Z(n8511) );
  XNOR U10174 ( .A(n8509), .B(n8508), .Z(n8510) );
  NANDN U10175 ( .A(n8511), .B(n8510), .Z(n8513) );
  NAND U10176 ( .A(a[25]), .B(b[40]), .Z(n8718) );
  XNOR U10177 ( .A(n8511), .B(n8510), .Z(n8719) );
  NANDN U10178 ( .A(n8718), .B(n8719), .Z(n8512) );
  AND U10179 ( .A(n8513), .B(n8512), .Z(n8517) );
  XNOR U10180 ( .A(n8515), .B(n8514), .Z(n8516) );
  NANDN U10181 ( .A(n8517), .B(n8516), .Z(n8519) );
  NAND U10182 ( .A(a[26]), .B(b[40]), .Z(n8867) );
  XNOR U10183 ( .A(n8517), .B(n8516), .Z(n8868) );
  NANDN U10184 ( .A(n8867), .B(n8868), .Z(n8518) );
  AND U10185 ( .A(n8519), .B(n8518), .Z(n8874) );
  XNOR U10186 ( .A(n8521), .B(n8520), .Z(n8873) );
  NANDN U10187 ( .A(n8874), .B(n8873), .Z(n8522) );
  AND U10188 ( .A(n8523), .B(n8522), .Z(n8527) );
  XNOR U10189 ( .A(n8525), .B(n8524), .Z(n8526) );
  NANDN U10190 ( .A(n8527), .B(n8526), .Z(n8529) );
  NAND U10191 ( .A(a[28]), .B(b[40]), .Z(n8879) );
  XNOR U10192 ( .A(n8527), .B(n8526), .Z(n8880) );
  NANDN U10193 ( .A(n8879), .B(n8880), .Z(n8528) );
  AND U10194 ( .A(n8529), .B(n8528), .Z(n8886) );
  XNOR U10195 ( .A(n8531), .B(n8530), .Z(n8885) );
  NANDN U10196 ( .A(n8886), .B(n8885), .Z(n8532) );
  AND U10197 ( .A(n8533), .B(n8532), .Z(n8537) );
  XNOR U10198 ( .A(n8535), .B(n8534), .Z(n8536) );
  NANDN U10199 ( .A(n8537), .B(n8536), .Z(n8539) );
  NAND U10200 ( .A(a[30]), .B(b[40]), .Z(n8891) );
  XNOR U10201 ( .A(n8537), .B(n8536), .Z(n8892) );
  NANDN U10202 ( .A(n8891), .B(n8892), .Z(n8538) );
  AND U10203 ( .A(n8539), .B(n8538), .Z(n8717) );
  XNOR U10204 ( .A(n8541), .B(n8540), .Z(n8716) );
  NANDN U10205 ( .A(n8717), .B(n8716), .Z(n8542) );
  AND U10206 ( .A(n8543), .B(n8542), .Z(n8547) );
  XNOR U10207 ( .A(n8545), .B(n8544), .Z(n8546) );
  NANDN U10208 ( .A(n8547), .B(n8546), .Z(n8549) );
  NAND U10209 ( .A(a[32]), .B(b[40]), .Z(n8901) );
  XNOR U10210 ( .A(n8547), .B(n8546), .Z(n8902) );
  NANDN U10211 ( .A(n8901), .B(n8902), .Z(n8548) );
  AND U10212 ( .A(n8549), .B(n8548), .Z(n8908) );
  XNOR U10213 ( .A(n8551), .B(n8550), .Z(n8907) );
  NANDN U10214 ( .A(n8908), .B(n8907), .Z(n8552) );
  AND U10215 ( .A(n8553), .B(n8552), .Z(n8914) );
  XNOR U10216 ( .A(n8555), .B(n8554), .Z(n8913) );
  NANDN U10217 ( .A(n8914), .B(n8913), .Z(n8556) );
  AND U10218 ( .A(n8557), .B(n8556), .Z(n8561) );
  XNOR U10219 ( .A(n8559), .B(n8558), .Z(n8560) );
  NANDN U10220 ( .A(n8561), .B(n8560), .Z(n8563) );
  NAND U10221 ( .A(a[35]), .B(b[40]), .Z(n8714) );
  XNOR U10222 ( .A(n8561), .B(n8560), .Z(n8715) );
  NANDN U10223 ( .A(n8714), .B(n8715), .Z(n8562) );
  AND U10224 ( .A(n8563), .B(n8562), .Z(n8564) );
  NANDN U10225 ( .A(n8565), .B(n8564), .Z(n8567) );
  XOR U10226 ( .A(n8565), .B(n8564), .Z(n8712) );
  AND U10227 ( .A(a[36]), .B(b[40]), .Z(n8713) );
  OR U10228 ( .A(n8712), .B(n8713), .Z(n8566) );
  NAND U10229 ( .A(n8567), .B(n8566), .Z(n8927) );
  XNOR U10230 ( .A(n8569), .B(n8568), .Z(n8928) );
  NANDN U10231 ( .A(n8927), .B(n8928), .Z(n8570) );
  AND U10232 ( .A(n8571), .B(n8570), .Z(n8711) );
  OR U10233 ( .A(n8710), .B(n8711), .Z(n8572) );
  NAND U10234 ( .A(n8573), .B(n8572), .Z(n8574) );
  NANDN U10235 ( .A(n8575), .B(n8574), .Z(n8577) );
  NAND U10236 ( .A(a[39]), .B(b[40]), .Z(n8706) );
  XNOR U10237 ( .A(n8575), .B(n8574), .Z(n8707) );
  NANDN U10238 ( .A(n8706), .B(n8707), .Z(n8576) );
  AND U10239 ( .A(n8577), .B(n8576), .Z(n8705) );
  XNOR U10240 ( .A(n8579), .B(n8578), .Z(n8704) );
  NANDN U10241 ( .A(n8705), .B(n8704), .Z(n8580) );
  AND U10242 ( .A(n8581), .B(n8580), .Z(n8585) );
  AND U10243 ( .A(a[41]), .B(b[40]), .Z(n8584) );
  NANDN U10244 ( .A(n8585), .B(n8584), .Z(n8587) );
  XOR U10245 ( .A(n8583), .B(n8582), .Z(n8700) );
  XNOR U10246 ( .A(n8585), .B(n8584), .Z(n8701) );
  NANDN U10247 ( .A(n8700), .B(n8701), .Z(n8586) );
  AND U10248 ( .A(n8587), .B(n8586), .Z(n8946) );
  XNOR U10249 ( .A(n8589), .B(n8588), .Z(n8945) );
  NANDN U10250 ( .A(n8946), .B(n8945), .Z(n8590) );
  NAND U10251 ( .A(n8591), .B(n8590), .Z(n8592) );
  NANDN U10252 ( .A(n8593), .B(n8592), .Z(n8595) );
  XNOR U10253 ( .A(n8593), .B(n8592), .Z(n8699) );
  AND U10254 ( .A(a[43]), .B(b[40]), .Z(n8698) );
  NAND U10255 ( .A(n8699), .B(n8698), .Z(n8594) );
  AND U10256 ( .A(n8595), .B(n8594), .Z(n8697) );
  XNOR U10257 ( .A(n8597), .B(n8596), .Z(n8696) );
  NANDN U10258 ( .A(n8697), .B(n8696), .Z(n8598) );
  AND U10259 ( .A(n8599), .B(n8598), .Z(n8603) );
  XNOR U10260 ( .A(n8601), .B(n8600), .Z(n8602) );
  NANDN U10261 ( .A(n8603), .B(n8602), .Z(n8605) );
  NAND U10262 ( .A(a[45]), .B(b[40]), .Z(n8959) );
  XNOR U10263 ( .A(n8603), .B(n8602), .Z(n8960) );
  NANDN U10264 ( .A(n8959), .B(n8960), .Z(n8604) );
  AND U10265 ( .A(n8605), .B(n8604), .Z(n8609) );
  XNOR U10266 ( .A(n8607), .B(n8606), .Z(n8608) );
  NANDN U10267 ( .A(n8609), .B(n8608), .Z(n8611) );
  NAND U10268 ( .A(a[46]), .B(b[40]), .Z(n8694) );
  XNOR U10269 ( .A(n8609), .B(n8608), .Z(n8695) );
  NANDN U10270 ( .A(n8694), .B(n8695), .Z(n8610) );
  AND U10271 ( .A(n8611), .B(n8610), .Z(n8693) );
  XNOR U10272 ( .A(n8613), .B(n8612), .Z(n8692) );
  NANDN U10273 ( .A(n8693), .B(n8692), .Z(n8614) );
  AND U10274 ( .A(n8615), .B(n8614), .Z(n8974) );
  XNOR U10275 ( .A(n8617), .B(n8616), .Z(n8973) );
  NANDN U10276 ( .A(n8974), .B(n8973), .Z(n8618) );
  AND U10277 ( .A(n8619), .B(n8618), .Z(n8623) );
  XNOR U10278 ( .A(n8621), .B(n8620), .Z(n8622) );
  NANDN U10279 ( .A(n8623), .B(n8622), .Z(n8625) );
  NAND U10280 ( .A(a[49]), .B(b[40]), .Z(n8688) );
  XNOR U10281 ( .A(n8623), .B(n8622), .Z(n8689) );
  NANDN U10282 ( .A(n8688), .B(n8689), .Z(n8624) );
  AND U10283 ( .A(n8625), .B(n8624), .Z(n8982) );
  XNOR U10284 ( .A(n8627), .B(n8626), .Z(n8981) );
  NANDN U10285 ( .A(n8982), .B(n8981), .Z(n8628) );
  AND U10286 ( .A(n8629), .B(n8628), .Z(n8633) );
  XNOR U10287 ( .A(n8631), .B(n8630), .Z(n8632) );
  NANDN U10288 ( .A(n8633), .B(n8632), .Z(n8635) );
  NAND U10289 ( .A(a[51]), .B(b[40]), .Z(n8987) );
  XNOR U10290 ( .A(n8633), .B(n8632), .Z(n8988) );
  NANDN U10291 ( .A(n8987), .B(n8988), .Z(n8634) );
  AND U10292 ( .A(n8635), .B(n8634), .Z(n8639) );
  XNOR U10293 ( .A(n8637), .B(n8636), .Z(n8638) );
  NANDN U10294 ( .A(n8639), .B(n8638), .Z(n8641) );
  NAND U10295 ( .A(a[52]), .B(b[40]), .Z(n8686) );
  XNOR U10296 ( .A(n8639), .B(n8638), .Z(n8687) );
  NANDN U10297 ( .A(n8686), .B(n8687), .Z(n8640) );
  AND U10298 ( .A(n8641), .B(n8640), .Z(n8685) );
  OR U10299 ( .A(n8684), .B(n8685), .Z(n8642) );
  AND U10300 ( .A(n8643), .B(n8642), .Z(n8683) );
  XNOR U10301 ( .A(n8645), .B(n8644), .Z(n8682) );
  NANDN U10302 ( .A(n8683), .B(n8682), .Z(n8646) );
  AND U10303 ( .A(n8647), .B(n8646), .Z(n8648) );
  NAND U10304 ( .A(n8649), .B(n8648), .Z(n8651) );
  AND U10305 ( .A(a[55]), .B(b[40]), .Z(n8681) );
  XOR U10306 ( .A(n8649), .B(n8648), .Z(n8680) );
  NANDN U10307 ( .A(n8681), .B(n8680), .Z(n8650) );
  AND U10308 ( .A(n8651), .B(n8650), .Z(n8654) );
  XNOR U10309 ( .A(n8653), .B(n8652), .Z(n8655) );
  NANDN U10310 ( .A(n8654), .B(n8655), .Z(n8657) );
  AND U10311 ( .A(a[56]), .B(b[40]), .Z(n8678) );
  NANDN U10312 ( .A(n8678), .B(n8679), .Z(n8656) );
  AND U10313 ( .A(n8657), .B(n8656), .Z(n8661) );
  NAND U10314 ( .A(n8661), .B(n8660), .Z(n8663) );
  NAND U10315 ( .A(a[57]), .B(b[40]), .Z(n8676) );
  XOR U10316 ( .A(n8661), .B(n8660), .Z(n8677) );
  NANDN U10317 ( .A(n8676), .B(n8677), .Z(n8662) );
  AND U10318 ( .A(n8663), .B(n8662), .Z(n8666) );
  NAND U10319 ( .A(n8666), .B(n8667), .Z(n8669) );
  AND U10320 ( .A(a[58]), .B(b[40]), .Z(n9017) );
  XOR U10321 ( .A(n8667), .B(n8666), .Z(n9018) );
  NANDN U10322 ( .A(n9017), .B(n9018), .Z(n8668) );
  NAND U10323 ( .A(n8669), .B(n8668), .Z(n8673) );
  NANDN U10324 ( .A(n8672), .B(n8673), .Z(n8675) );
  NAND U10325 ( .A(n9022), .B(n9021), .Z(n8674) );
  NAND U10326 ( .A(n8675), .B(n8674), .Z(n10238) );
  XNOR U10327 ( .A(n10240), .B(n10241), .Z(n10246) );
  AND U10328 ( .A(a[58]), .B(b[39]), .Z(n9012) );
  NAND U10329 ( .A(n9012), .B(n9011), .Z(n9014) );
  AND U10330 ( .A(a[57]), .B(b[39]), .Z(n9007) );
  NAND U10331 ( .A(n9008), .B(n9007), .Z(n9010) );
  XOR U10332 ( .A(n8681), .B(n8680), .Z(n9006) );
  AND U10333 ( .A(a[56]), .B(b[39]), .Z(n9005) );
  XOR U10334 ( .A(n8683), .B(n8682), .Z(n9001) );
  XOR U10335 ( .A(n8685), .B(n8684), .Z(n8998) );
  NAND U10336 ( .A(a[53]), .B(b[39]), .Z(n8993) );
  XNOR U10337 ( .A(n8687), .B(n8686), .Z(n8994) );
  NANDN U10338 ( .A(n8993), .B(n8994), .Z(n8996) );
  XOR U10339 ( .A(n8689), .B(n8688), .Z(n8690) );
  AND U10340 ( .A(a[50]), .B(b[39]), .Z(n8691) );
  NANDN U10341 ( .A(n8690), .B(n8691), .Z(n8980) );
  XOR U10342 ( .A(n8691), .B(n8690), .Z(n9327) );
  XOR U10343 ( .A(n8693), .B(n8692), .Z(n8969) );
  AND U10344 ( .A(a[48]), .B(b[39]), .Z(n8970) );
  NANDN U10345 ( .A(n8969), .B(n8970), .Z(n8972) );
  NAND U10346 ( .A(a[47]), .B(b[39]), .Z(n8965) );
  XNOR U10347 ( .A(n8695), .B(n8694), .Z(n8966) );
  NANDN U10348 ( .A(n8965), .B(n8966), .Z(n8968) );
  XOR U10349 ( .A(n8697), .B(n8696), .Z(n8955) );
  AND U10350 ( .A(a[44]), .B(b[39]), .Z(n8952) );
  XNOR U10351 ( .A(n8699), .B(n8698), .Z(n8951) );
  NANDN U10352 ( .A(n8952), .B(n8951), .Z(n8954) );
  XOR U10353 ( .A(n8701), .B(n8700), .Z(n8702) );
  AND U10354 ( .A(a[42]), .B(b[39]), .Z(n8703) );
  NANDN U10355 ( .A(n8702), .B(n8703), .Z(n8944) );
  XOR U10356 ( .A(n8703), .B(n8702), .Z(n9031) );
  NAND U10357 ( .A(a[41]), .B(b[39]), .Z(n8939) );
  XNOR U10358 ( .A(n8705), .B(n8704), .Z(n8940) );
  NANDN U10359 ( .A(n8939), .B(n8940), .Z(n8942) );
  NAND U10360 ( .A(a[40]), .B(b[39]), .Z(n8708) );
  XNOR U10361 ( .A(n8707), .B(n8706), .Z(n8709) );
  NANDN U10362 ( .A(n8708), .B(n8709), .Z(n8938) );
  XOR U10363 ( .A(n8709), .B(n8708), .Z(n9267) );
  XOR U10364 ( .A(n8711), .B(n8710), .Z(n8934) );
  XOR U10365 ( .A(n8713), .B(n8712), .Z(n8924) );
  XOR U10366 ( .A(n8715), .B(n8714), .Z(n8919) );
  AND U10367 ( .A(a[36]), .B(b[39]), .Z(n8920) );
  NANDN U10368 ( .A(n8919), .B(n8920), .Z(n8922) );
  XOR U10369 ( .A(n8717), .B(n8716), .Z(n8897) );
  AND U10370 ( .A(a[32]), .B(b[39]), .Z(n8898) );
  NANDN U10371 ( .A(n8897), .B(n8898), .Z(n8900) );
  XOR U10372 ( .A(n8719), .B(n8718), .Z(n8863) );
  AND U10373 ( .A(a[26]), .B(b[39]), .Z(n8864) );
  NANDN U10374 ( .A(n8863), .B(n8864), .Z(n8866) );
  AND U10375 ( .A(a[25]), .B(b[39]), .Z(n8860) );
  NAND U10376 ( .A(n8860), .B(n8859), .Z(n8862) );
  NAND U10377 ( .A(a[24]), .B(b[39]), .Z(n8855) );
  XOR U10378 ( .A(n8723), .B(n8722), .Z(n8856) );
  NANDN U10379 ( .A(n8855), .B(n8856), .Z(n8858) );
  AND U10380 ( .A(a[23]), .B(b[39]), .Z(n8852) );
  NAND U10381 ( .A(n8852), .B(n8851), .Z(n8854) );
  AND U10382 ( .A(a[22]), .B(b[39]), .Z(n8728) );
  NAND U10383 ( .A(n8728), .B(n8729), .Z(n8850) );
  XOR U10384 ( .A(n8729), .B(n8728), .Z(n9164) );
  XOR U10385 ( .A(n8731), .B(n8730), .Z(n8845) );
  XOR U10386 ( .A(n8733), .B(n8732), .Z(n8841) );
  AND U10387 ( .A(a[20]), .B(b[39]), .Z(n8842) );
  NANDN U10388 ( .A(n8841), .B(n8842), .Z(n8844) );
  XOR U10389 ( .A(n8735), .B(n8734), .Z(n8837) );
  AND U10390 ( .A(a[16]), .B(b[39]), .Z(n8822) );
  NAND U10391 ( .A(n8822), .B(n8821), .Z(n8824) );
  NAND U10392 ( .A(a[14]), .B(b[39]), .Z(n8811) );
  NANDN U10393 ( .A(n8811), .B(n8812), .Z(n8814) );
  XOR U10394 ( .A(n8741), .B(n8740), .Z(n8801) );
  XOR U10395 ( .A(n8743), .B(n8742), .Z(n8797) );
  AND U10396 ( .A(a[8]), .B(b[39]), .Z(n8782) );
  NAND U10397 ( .A(n8782), .B(n8781), .Z(n8784) );
  AND U10398 ( .A(a[7]), .B(b[39]), .Z(n8778) );
  NAND U10399 ( .A(n8778), .B(n8777), .Z(n8780) );
  XOR U10400 ( .A(n8749), .B(n8748), .Z(n8767) );
  NAND U10401 ( .A(a[0]), .B(b[39]), .Z(n9431) );
  AND U10402 ( .A(a[1]), .B(b[40]), .Z(n8752) );
  NANDN U10403 ( .A(n9431), .B(n8752), .Z(n9049) );
  NANDN U10404 ( .A(n9049), .B(n8750), .Z(n8754) );
  AND U10405 ( .A(a[2]), .B(b[39]), .Z(n9056) );
  NANDN U10406 ( .A(n9055), .B(n9056), .Z(n8753) );
  AND U10407 ( .A(n8754), .B(n8753), .Z(n8757) );
  AND U10408 ( .A(a[3]), .B(b[39]), .Z(n8758) );
  NANDN U10409 ( .A(n8757), .B(n8758), .Z(n8760) );
  XNOR U10410 ( .A(n8756), .B(n8755), .Z(n9062) );
  NAND U10411 ( .A(n9062), .B(n9061), .Z(n8759) );
  AND U10412 ( .A(n8760), .B(n8759), .Z(n8763) );
  NANDN U10413 ( .A(n8763), .B(n8764), .Z(n8766) );
  NAND U10414 ( .A(a[4]), .B(b[39]), .Z(n9067) );
  NANDN U10415 ( .A(n9067), .B(n9068), .Z(n8765) );
  AND U10416 ( .A(n8766), .B(n8765), .Z(n8768) );
  NANDN U10417 ( .A(n8767), .B(n8768), .Z(n8770) );
  NAND U10418 ( .A(a[5]), .B(b[39]), .Z(n9073) );
  NAND U10419 ( .A(n9074), .B(n9073), .Z(n8769) );
  AND U10420 ( .A(n8770), .B(n8769), .Z(n8774) );
  XOR U10421 ( .A(n8772), .B(n8771), .Z(n8773) );
  NAND U10422 ( .A(n8774), .B(n8773), .Z(n8776) );
  NAND U10423 ( .A(a[6]), .B(b[39]), .Z(n9081) );
  XOR U10424 ( .A(n8774), .B(n8773), .Z(n9082) );
  NANDN U10425 ( .A(n9081), .B(n9082), .Z(n8775) );
  AND U10426 ( .A(n8776), .B(n8775), .Z(n9085) );
  XOR U10427 ( .A(n8778), .B(n8777), .Z(n9086) );
  NANDN U10428 ( .A(n9085), .B(n9086), .Z(n8779) );
  AND U10429 ( .A(n8780), .B(n8779), .Z(n9046) );
  XOR U10430 ( .A(n8782), .B(n8781), .Z(n9045) );
  NANDN U10431 ( .A(n9046), .B(n9045), .Z(n8783) );
  AND U10432 ( .A(n8784), .B(n8783), .Z(n8787) );
  NAND U10433 ( .A(n8787), .B(n8788), .Z(n8790) );
  AND U10434 ( .A(a[9]), .B(b[39]), .Z(n9095) );
  XOR U10435 ( .A(n8788), .B(n8787), .Z(n9096) );
  NANDN U10436 ( .A(n9095), .B(n9096), .Z(n8789) );
  AND U10437 ( .A(n8790), .B(n8789), .Z(n8793) );
  NAND U10438 ( .A(n8793), .B(n8794), .Z(n8796) );
  NAND U10439 ( .A(a[10]), .B(b[39]), .Z(n9099) );
  XOR U10440 ( .A(n8794), .B(n8793), .Z(n9100) );
  NANDN U10441 ( .A(n9099), .B(n9100), .Z(n8795) );
  AND U10442 ( .A(n8796), .B(n8795), .Z(n8798) );
  NANDN U10443 ( .A(n8797), .B(n8798), .Z(n8800) );
  AND U10444 ( .A(a[11]), .B(b[39]), .Z(n9043) );
  NANDN U10445 ( .A(n9043), .B(n9044), .Z(n8799) );
  AND U10446 ( .A(n8800), .B(n8799), .Z(n8802) );
  NANDN U10447 ( .A(n8801), .B(n8802), .Z(n8804) );
  NAND U10448 ( .A(a[12]), .B(b[39]), .Z(n9109) );
  NANDN U10449 ( .A(n9109), .B(n9110), .Z(n8803) );
  AND U10450 ( .A(n8804), .B(n8803), .Z(n8807) );
  XOR U10451 ( .A(n8806), .B(n8805), .Z(n8808) );
  NANDN U10452 ( .A(n8807), .B(n8808), .Z(n8810) );
  NAND U10453 ( .A(a[13]), .B(b[39]), .Z(n9115) );
  NANDN U10454 ( .A(n9115), .B(n9116), .Z(n8809) );
  AND U10455 ( .A(n8810), .B(n8809), .Z(n9041) );
  NANDN U10456 ( .A(n9041), .B(n9042), .Z(n8813) );
  AND U10457 ( .A(n8814), .B(n8813), .Z(n8817) );
  NANDN U10458 ( .A(n8817), .B(n8818), .Z(n8820) );
  AND U10459 ( .A(a[15]), .B(b[39]), .Z(n9128) );
  NAND U10460 ( .A(n9128), .B(n9127), .Z(n8819) );
  AND U10461 ( .A(n8820), .B(n8819), .Z(n9131) );
  XOR U10462 ( .A(n8822), .B(n8821), .Z(n9132) );
  NANDN U10463 ( .A(n9131), .B(n9132), .Z(n8823) );
  AND U10464 ( .A(n8824), .B(n8823), .Z(n8828) );
  NAND U10465 ( .A(n8828), .B(n8827), .Z(n8830) );
  AND U10466 ( .A(a[17]), .B(b[39]), .Z(n9137) );
  XOR U10467 ( .A(n8828), .B(n8827), .Z(n9138) );
  NANDN U10468 ( .A(n9137), .B(n9138), .Z(n8829) );
  AND U10469 ( .A(n8830), .B(n8829), .Z(n8833) );
  NAND U10470 ( .A(n8833), .B(n8834), .Z(n8836) );
  XOR U10471 ( .A(n8834), .B(n8833), .Z(n9040) );
  AND U10472 ( .A(a[18]), .B(b[39]), .Z(n9039) );
  NAND U10473 ( .A(n9040), .B(n9039), .Z(n8835) );
  AND U10474 ( .A(n8836), .B(n8835), .Z(n8838) );
  NANDN U10475 ( .A(n8837), .B(n8838), .Z(n8840) );
  AND U10476 ( .A(a[19]), .B(b[39]), .Z(n9147) );
  NANDN U10477 ( .A(n9147), .B(n9148), .Z(n8839) );
  AND U10478 ( .A(n8840), .B(n8839), .Z(n9038) );
  NAND U10479 ( .A(n9038), .B(n9037), .Z(n8843) );
  AND U10480 ( .A(n8844), .B(n8843), .Z(n8846) );
  NANDN U10481 ( .A(n8845), .B(n8846), .Z(n8848) );
  AND U10482 ( .A(a[21]), .B(b[39]), .Z(n9157) );
  NANDN U10483 ( .A(n9157), .B(n9158), .Z(n8847) );
  AND U10484 ( .A(n8848), .B(n8847), .Z(n9163) );
  NAND U10485 ( .A(n9164), .B(n9163), .Z(n8849) );
  AND U10486 ( .A(n8850), .B(n8849), .Z(n9035) );
  XOR U10487 ( .A(n8852), .B(n8851), .Z(n9036) );
  NANDN U10488 ( .A(n9035), .B(n9036), .Z(n8853) );
  AND U10489 ( .A(n8854), .B(n8853), .Z(n9033) );
  NANDN U10490 ( .A(n9033), .B(n9034), .Z(n8857) );
  AND U10491 ( .A(n8858), .B(n8857), .Z(n9177) );
  XOR U10492 ( .A(n8860), .B(n8859), .Z(n9178) );
  NANDN U10493 ( .A(n9177), .B(n9178), .Z(n8861) );
  AND U10494 ( .A(n8862), .B(n8861), .Z(n9184) );
  XNOR U10495 ( .A(n8864), .B(n8863), .Z(n9183) );
  NANDN U10496 ( .A(n9184), .B(n9183), .Z(n8865) );
  AND U10497 ( .A(n8866), .B(n8865), .Z(n8870) );
  XNOR U10498 ( .A(n8868), .B(n8867), .Z(n8869) );
  NANDN U10499 ( .A(n8870), .B(n8869), .Z(n8872) );
  NAND U10500 ( .A(a[27]), .B(b[39]), .Z(n9189) );
  XNOR U10501 ( .A(n8870), .B(n8869), .Z(n9190) );
  NANDN U10502 ( .A(n9189), .B(n9190), .Z(n8871) );
  AND U10503 ( .A(n8872), .B(n8871), .Z(n8876) );
  XNOR U10504 ( .A(n8874), .B(n8873), .Z(n8875) );
  NANDN U10505 ( .A(n8876), .B(n8875), .Z(n8878) );
  NAND U10506 ( .A(a[28]), .B(b[39]), .Z(n9195) );
  XNOR U10507 ( .A(n8876), .B(n8875), .Z(n9196) );
  NANDN U10508 ( .A(n9195), .B(n9196), .Z(n8877) );
  AND U10509 ( .A(n8878), .B(n8877), .Z(n8882) );
  XNOR U10510 ( .A(n8880), .B(n8879), .Z(n8881) );
  NANDN U10511 ( .A(n8882), .B(n8881), .Z(n8884) );
  NAND U10512 ( .A(a[29]), .B(b[39]), .Z(n9201) );
  XNOR U10513 ( .A(n8882), .B(n8881), .Z(n9202) );
  NANDN U10514 ( .A(n9201), .B(n9202), .Z(n8883) );
  AND U10515 ( .A(n8884), .B(n8883), .Z(n8888) );
  XNOR U10516 ( .A(n8886), .B(n8885), .Z(n8887) );
  NANDN U10517 ( .A(n8888), .B(n8887), .Z(n8890) );
  NAND U10518 ( .A(a[30]), .B(b[39]), .Z(n9207) );
  XNOR U10519 ( .A(n8888), .B(n8887), .Z(n9208) );
  NANDN U10520 ( .A(n9207), .B(n9208), .Z(n8889) );
  AND U10521 ( .A(n8890), .B(n8889), .Z(n8894) );
  XNOR U10522 ( .A(n8892), .B(n8891), .Z(n8893) );
  NANDN U10523 ( .A(n8894), .B(n8893), .Z(n8896) );
  XNOR U10524 ( .A(n8894), .B(n8893), .Z(n9216) );
  AND U10525 ( .A(a[31]), .B(b[39]), .Z(n9215) );
  NAND U10526 ( .A(n9216), .B(n9215), .Z(n8895) );
  AND U10527 ( .A(n8896), .B(n8895), .Z(n9220) );
  XNOR U10528 ( .A(n8898), .B(n8897), .Z(n9219) );
  NANDN U10529 ( .A(n9220), .B(n9219), .Z(n8899) );
  AND U10530 ( .A(n8900), .B(n8899), .Z(n8904) );
  XNOR U10531 ( .A(n8902), .B(n8901), .Z(n8903) );
  NANDN U10532 ( .A(n8904), .B(n8903), .Z(n8906) );
  NAND U10533 ( .A(a[33]), .B(b[39]), .Z(n9225) );
  XNOR U10534 ( .A(n8904), .B(n8903), .Z(n9226) );
  NANDN U10535 ( .A(n9225), .B(n9226), .Z(n8905) );
  AND U10536 ( .A(n8906), .B(n8905), .Z(n8910) );
  XNOR U10537 ( .A(n8908), .B(n8907), .Z(n8909) );
  NANDN U10538 ( .A(n8910), .B(n8909), .Z(n8912) );
  NAND U10539 ( .A(a[34]), .B(b[39]), .Z(n9231) );
  XNOR U10540 ( .A(n8910), .B(n8909), .Z(n9232) );
  NANDN U10541 ( .A(n9231), .B(n9232), .Z(n8911) );
  AND U10542 ( .A(n8912), .B(n8911), .Z(n8916) );
  XNOR U10543 ( .A(n8914), .B(n8913), .Z(n8915) );
  NANDN U10544 ( .A(n8916), .B(n8915), .Z(n8918) );
  NAND U10545 ( .A(a[35]), .B(b[39]), .Z(n9237) );
  XNOR U10546 ( .A(n8916), .B(n8915), .Z(n9238) );
  NANDN U10547 ( .A(n9237), .B(n9238), .Z(n8917) );
  AND U10548 ( .A(n8918), .B(n8917), .Z(n9244) );
  XNOR U10549 ( .A(n8920), .B(n8919), .Z(n9243) );
  NANDN U10550 ( .A(n9244), .B(n9243), .Z(n8921) );
  NAND U10551 ( .A(n8922), .B(n8921), .Z(n8923) );
  NANDN U10552 ( .A(n8924), .B(n8923), .Z(n8926) );
  XNOR U10553 ( .A(n8924), .B(n8923), .Z(n9252) );
  AND U10554 ( .A(a[37]), .B(b[39]), .Z(n9251) );
  NAND U10555 ( .A(n9252), .B(n9251), .Z(n8925) );
  AND U10556 ( .A(n8926), .B(n8925), .Z(n8930) );
  XNOR U10557 ( .A(n8928), .B(n8927), .Z(n8929) );
  NANDN U10558 ( .A(n8930), .B(n8929), .Z(n8932) );
  NAND U10559 ( .A(a[38]), .B(b[39]), .Z(n9257) );
  XNOR U10560 ( .A(n8930), .B(n8929), .Z(n9258) );
  NANDN U10561 ( .A(n9257), .B(n9258), .Z(n8931) );
  AND U10562 ( .A(n8932), .B(n8931), .Z(n8933) );
  NANDN U10563 ( .A(n8934), .B(n8933), .Z(n8936) );
  XOR U10564 ( .A(n8934), .B(n8933), .Z(n9261) );
  AND U10565 ( .A(a[39]), .B(b[39]), .Z(n9262) );
  OR U10566 ( .A(n9261), .B(n9262), .Z(n8935) );
  AND U10567 ( .A(n8936), .B(n8935), .Z(n9268) );
  NANDN U10568 ( .A(n9267), .B(n9268), .Z(n8937) );
  AND U10569 ( .A(n8938), .B(n8937), .Z(n9274) );
  XNOR U10570 ( .A(n8940), .B(n8939), .Z(n9273) );
  NANDN U10571 ( .A(n9274), .B(n9273), .Z(n8941) );
  AND U10572 ( .A(n8942), .B(n8941), .Z(n9032) );
  OR U10573 ( .A(n9031), .B(n9032), .Z(n8943) );
  AND U10574 ( .A(n8944), .B(n8943), .Z(n8948) );
  XNOR U10575 ( .A(n8946), .B(n8945), .Z(n8947) );
  NANDN U10576 ( .A(n8948), .B(n8947), .Z(n8950) );
  NAND U10577 ( .A(a[43]), .B(b[39]), .Z(n9283) );
  XNOR U10578 ( .A(n8948), .B(n8947), .Z(n9284) );
  NANDN U10579 ( .A(n9283), .B(n9284), .Z(n8949) );
  NAND U10580 ( .A(n8950), .B(n8949), .Z(n9291) );
  XNOR U10581 ( .A(n8952), .B(n8951), .Z(n9292) );
  NANDN U10582 ( .A(n9291), .B(n9292), .Z(n8953) );
  AND U10583 ( .A(n8954), .B(n8953), .Z(n8956) );
  NANDN U10584 ( .A(n8955), .B(n8956), .Z(n8958) );
  NAND U10585 ( .A(a[45]), .B(b[39]), .Z(n9295) );
  XNOR U10586 ( .A(n8956), .B(n8955), .Z(n9296) );
  NANDN U10587 ( .A(n9295), .B(n9296), .Z(n8957) );
  AND U10588 ( .A(n8958), .B(n8957), .Z(n8962) );
  XNOR U10589 ( .A(n8960), .B(n8959), .Z(n8961) );
  NANDN U10590 ( .A(n8962), .B(n8961), .Z(n8964) );
  NAND U10591 ( .A(a[46]), .B(b[39]), .Z(n9301) );
  XNOR U10592 ( .A(n8962), .B(n8961), .Z(n9302) );
  NANDN U10593 ( .A(n9301), .B(n9302), .Z(n8963) );
  AND U10594 ( .A(n8964), .B(n8963), .Z(n9308) );
  XNOR U10595 ( .A(n8966), .B(n8965), .Z(n9307) );
  NANDN U10596 ( .A(n9308), .B(n9307), .Z(n8967) );
  AND U10597 ( .A(n8968), .B(n8967), .Z(n9314) );
  XNOR U10598 ( .A(n8970), .B(n8969), .Z(n9313) );
  NANDN U10599 ( .A(n9314), .B(n9313), .Z(n8971) );
  AND U10600 ( .A(n8972), .B(n8971), .Z(n8976) );
  XNOR U10601 ( .A(n8974), .B(n8973), .Z(n8975) );
  NANDN U10602 ( .A(n8976), .B(n8975), .Z(n8978) );
  XNOR U10603 ( .A(n8976), .B(n8975), .Z(n9322) );
  AND U10604 ( .A(a[49]), .B(b[39]), .Z(n9321) );
  NAND U10605 ( .A(n9322), .B(n9321), .Z(n8977) );
  AND U10606 ( .A(n8978), .B(n8977), .Z(n9328) );
  OR U10607 ( .A(n9327), .B(n9328), .Z(n8979) );
  AND U10608 ( .A(n8980), .B(n8979), .Z(n8984) );
  XNOR U10609 ( .A(n8982), .B(n8981), .Z(n8983) );
  NANDN U10610 ( .A(n8984), .B(n8983), .Z(n8986) );
  NAND U10611 ( .A(a[51]), .B(b[39]), .Z(n9331) );
  XNOR U10612 ( .A(n8984), .B(n8983), .Z(n9332) );
  NANDN U10613 ( .A(n9331), .B(n9332), .Z(n8985) );
  AND U10614 ( .A(n8986), .B(n8985), .Z(n8990) );
  XNOR U10615 ( .A(n8988), .B(n8987), .Z(n8989) );
  NANDN U10616 ( .A(n8990), .B(n8989), .Z(n8992) );
  NAND U10617 ( .A(a[52]), .B(b[39]), .Z(n9337) );
  XNOR U10618 ( .A(n8990), .B(n8989), .Z(n9338) );
  NANDN U10619 ( .A(n9337), .B(n9338), .Z(n8991) );
  AND U10620 ( .A(n8992), .B(n8991), .Z(n9344) );
  XNOR U10621 ( .A(n8994), .B(n8993), .Z(n9343) );
  NANDN U10622 ( .A(n9344), .B(n9343), .Z(n8995) );
  AND U10623 ( .A(n8996), .B(n8995), .Z(n8997) );
  NANDN U10624 ( .A(n8998), .B(n8997), .Z(n9000) );
  XOR U10625 ( .A(n8998), .B(n8997), .Z(n9349) );
  AND U10626 ( .A(a[54]), .B(b[39]), .Z(n9350) );
  OR U10627 ( .A(n9349), .B(n9350), .Z(n8999) );
  AND U10628 ( .A(n9000), .B(n8999), .Z(n9002) );
  NANDN U10629 ( .A(n9001), .B(n9002), .Z(n9004) );
  NAND U10630 ( .A(a[55]), .B(b[39]), .Z(n9355) );
  XNOR U10631 ( .A(n9002), .B(n9001), .Z(n9356) );
  NANDN U10632 ( .A(n9355), .B(n9356), .Z(n9003) );
  AND U10633 ( .A(n9004), .B(n9003), .Z(n9030) );
  XOR U10634 ( .A(n9006), .B(n9005), .Z(n9029) );
  XOR U10635 ( .A(n9008), .B(n9007), .Z(n9027) );
  NANDN U10636 ( .A(n9028), .B(n9027), .Z(n9009) );
  AND U10637 ( .A(n9010), .B(n9009), .Z(n9365) );
  XOR U10638 ( .A(n9012), .B(n9011), .Z(n9366) );
  NANDN U10639 ( .A(n9365), .B(n9366), .Z(n9013) );
  AND U10640 ( .A(n9014), .B(n9013), .Z(n9015) );
  AND U10641 ( .A(a[59]), .B(b[39]), .Z(n9016) );
  NANDN U10642 ( .A(n9015), .B(n9016), .Z(n9020) );
  NAND U10643 ( .A(n9371), .B(n9372), .Z(n9019) );
  AND U10644 ( .A(n9020), .B(n9019), .Z(n9023) );
  AND U10645 ( .A(a[60]), .B(b[39]), .Z(n9024) );
  NANDN U10646 ( .A(n9023), .B(n9024), .Z(n9026) );
  XOR U10647 ( .A(n9022), .B(n9021), .Z(n9377) );
  NANDN U10648 ( .A(n9377), .B(n9378), .Z(n9025) );
  AND U10649 ( .A(n9026), .B(n9025), .Z(n10245) );
  AND U10650 ( .A(a[61]), .B(b[39]), .Z(n10244) );
  XNOR U10651 ( .A(n10246), .B(n10247), .Z(n10250) );
  XOR U10652 ( .A(n9028), .B(n9027), .Z(n9364) );
  XOR U10653 ( .A(n9030), .B(n9029), .Z(n9362) );
  NAND U10654 ( .A(a[52]), .B(b[38]), .Z(n9333) );
  AND U10655 ( .A(a[51]), .B(b[38]), .Z(n9326) );
  AND U10656 ( .A(a[50]), .B(b[38]), .Z(n9320) );
  NAND U10657 ( .A(a[46]), .B(b[38]), .Z(n9297) );
  AND U10658 ( .A(a[45]), .B(b[38]), .Z(n9290) );
  NAND U10659 ( .A(a[44]), .B(b[38]), .Z(n9285) );
  XOR U10660 ( .A(n9032), .B(n9031), .Z(n9280) );
  NAND U10661 ( .A(a[39]), .B(b[38]), .Z(n9255) );
  AND U10662 ( .A(a[38]), .B(b[38]), .Z(n9250) );
  AND U10663 ( .A(a[32]), .B(b[38]), .Z(n9214) );
  XOR U10664 ( .A(n9038), .B(n9037), .Z(n9153) );
  XOR U10665 ( .A(n9040), .B(n9039), .Z(n9143) );
  AND U10666 ( .A(a[15]), .B(b[38]), .Z(n9122) );
  NAND U10667 ( .A(n9122), .B(n9121), .Z(n9124) );
  AND U10668 ( .A(a[12]), .B(b[38]), .Z(n9106) );
  NAND U10669 ( .A(n9106), .B(n9105), .Z(n9108) );
  NAND U10670 ( .A(a[10]), .B(b[38]), .Z(n9093) );
  AND U10671 ( .A(a[9]), .B(b[38]), .Z(n9047) );
  XOR U10672 ( .A(n9046), .B(n9045), .Z(n9048) );
  NANDN U10673 ( .A(n9047), .B(n9048), .Z(n9092) );
  AND U10674 ( .A(a[0]), .B(b[38]), .Z(n9774) );
  AND U10675 ( .A(a[1]), .B(b[39]), .Z(n9052) );
  NAND U10676 ( .A(n9774), .B(n9052), .Z(n9429) );
  NANDN U10677 ( .A(n9429), .B(n9049), .Z(n9054) );
  AND U10678 ( .A(n9774), .B(n9052), .Z(n9050) );
  AND U10679 ( .A(a[2]), .B(b[38]), .Z(n9428) );
  NANDN U10680 ( .A(n9427), .B(n9428), .Z(n9053) );
  AND U10681 ( .A(n9054), .B(n9053), .Z(n9057) );
  XNOR U10682 ( .A(n9056), .B(n9055), .Z(n9058) );
  NANDN U10683 ( .A(n9057), .B(n9058), .Z(n9060) );
  NAND U10684 ( .A(a[3]), .B(b[38]), .Z(n9439) );
  NANDN U10685 ( .A(n9439), .B(n9440), .Z(n9059) );
  AND U10686 ( .A(n9060), .B(n9059), .Z(n9063) );
  XOR U10687 ( .A(n9062), .B(n9061), .Z(n9064) );
  NANDN U10688 ( .A(n9063), .B(n9064), .Z(n9066) );
  AND U10689 ( .A(a[4]), .B(b[38]), .Z(n9426) );
  NAND U10690 ( .A(n9426), .B(n9425), .Z(n9065) );
  AND U10691 ( .A(n9066), .B(n9065), .Z(n9069) );
  NANDN U10692 ( .A(n9069), .B(n9070), .Z(n9072) );
  AND U10693 ( .A(a[5]), .B(b[38]), .Z(n9450) );
  NAND U10694 ( .A(n9450), .B(n9449), .Z(n9071) );
  AND U10695 ( .A(n9072), .B(n9071), .Z(n9075) );
  AND U10696 ( .A(a[6]), .B(b[38]), .Z(n9076) );
  NANDN U10697 ( .A(n9075), .B(n9076), .Z(n9078) );
  XOR U10698 ( .A(n9074), .B(n9073), .Z(n9455) );
  NANDN U10699 ( .A(n9455), .B(n9456), .Z(n9077) );
  AND U10700 ( .A(n9078), .B(n9077), .Z(n9079) );
  AND U10701 ( .A(a[7]), .B(b[38]), .Z(n9080) );
  NANDN U10702 ( .A(n9079), .B(n9080), .Z(n9084) );
  NAND U10703 ( .A(n9464), .B(n9463), .Z(n9083) );
  AND U10704 ( .A(n9084), .B(n9083), .Z(n9087) );
  NAND U10705 ( .A(n9087), .B(n9088), .Z(n9090) );
  AND U10706 ( .A(a[8]), .B(b[38]), .Z(n9423) );
  XOR U10707 ( .A(n9088), .B(n9087), .Z(n9424) );
  NANDN U10708 ( .A(n9423), .B(n9424), .Z(n9089) );
  NAND U10709 ( .A(n9090), .B(n9089), .Z(n9421) );
  NAND U10710 ( .A(n9422), .B(n9421), .Z(n9091) );
  AND U10711 ( .A(n9092), .B(n9091), .Z(n9094) );
  NANDN U10712 ( .A(n9093), .B(n9094), .Z(n9098) );
  NAND U10713 ( .A(n9419), .B(n9420), .Z(n9097) );
  AND U10714 ( .A(n9098), .B(n9097), .Z(n9101) );
  NANDN U10715 ( .A(n9101), .B(n9102), .Z(n9104) );
  NAND U10716 ( .A(a[11]), .B(b[38]), .Z(n9417) );
  NANDN U10717 ( .A(n9417), .B(n9418), .Z(n9103) );
  AND U10718 ( .A(n9104), .B(n9103), .Z(n9415) );
  XOR U10719 ( .A(n9106), .B(n9105), .Z(n9416) );
  NANDN U10720 ( .A(n9415), .B(n9416), .Z(n9107) );
  AND U10721 ( .A(n9108), .B(n9107), .Z(n9111) );
  NANDN U10722 ( .A(n9111), .B(n9112), .Z(n9114) );
  NAND U10723 ( .A(a[13]), .B(b[38]), .Z(n9413) );
  NANDN U10724 ( .A(n9413), .B(n9414), .Z(n9113) );
  AND U10725 ( .A(n9114), .B(n9113), .Z(n9117) );
  NANDN U10726 ( .A(n9117), .B(n9118), .Z(n9120) );
  NAND U10727 ( .A(a[14]), .B(b[38]), .Z(n9491) );
  NANDN U10728 ( .A(n9491), .B(n9492), .Z(n9119) );
  AND U10729 ( .A(n9120), .B(n9119), .Z(n9497) );
  XOR U10730 ( .A(n9122), .B(n9121), .Z(n9498) );
  NANDN U10731 ( .A(n9497), .B(n9498), .Z(n9123) );
  AND U10732 ( .A(n9124), .B(n9123), .Z(n9125) );
  AND U10733 ( .A(a[16]), .B(b[38]), .Z(n9126) );
  NANDN U10734 ( .A(n9125), .B(n9126), .Z(n9130) );
  XOR U10735 ( .A(n9128), .B(n9127), .Z(n9503) );
  NAND U10736 ( .A(n9504), .B(n9503), .Z(n9129) );
  AND U10737 ( .A(n9130), .B(n9129), .Z(n9133) );
  NAND U10738 ( .A(n9133), .B(n9134), .Z(n9136) );
  AND U10739 ( .A(a[17]), .B(b[38]), .Z(n9511) );
  XOR U10740 ( .A(n9134), .B(n9133), .Z(n9512) );
  NANDN U10741 ( .A(n9511), .B(n9512), .Z(n9135) );
  AND U10742 ( .A(n9136), .B(n9135), .Z(n9139) );
  NAND U10743 ( .A(n9139), .B(n9140), .Z(n9142) );
  NAND U10744 ( .A(a[18]), .B(b[38]), .Z(n9515) );
  XOR U10745 ( .A(n9140), .B(n9139), .Z(n9516) );
  NANDN U10746 ( .A(n9515), .B(n9516), .Z(n9141) );
  AND U10747 ( .A(n9142), .B(n9141), .Z(n9144) );
  NANDN U10748 ( .A(n9143), .B(n9144), .Z(n9146) );
  AND U10749 ( .A(a[19]), .B(b[38]), .Z(n9523) );
  NANDN U10750 ( .A(n9523), .B(n9524), .Z(n9145) );
  AND U10751 ( .A(n9146), .B(n9145), .Z(n9149) );
  NANDN U10752 ( .A(n9149), .B(n9150), .Z(n9152) );
  AND U10753 ( .A(a[20]), .B(b[38]), .Z(n9411) );
  NANDN U10754 ( .A(n9411), .B(n9412), .Z(n9151) );
  NAND U10755 ( .A(n9152), .B(n9151), .Z(n9154) );
  NANDN U10756 ( .A(n9153), .B(n9154), .Z(n9156) );
  AND U10757 ( .A(a[21]), .B(b[38]), .Z(n9529) );
  NANDN U10758 ( .A(n9529), .B(n9530), .Z(n9155) );
  AND U10759 ( .A(n9156), .B(n9155), .Z(n9159) );
  NANDN U10760 ( .A(n9159), .B(n9160), .Z(n9162) );
  AND U10761 ( .A(a[22]), .B(b[38]), .Z(n9409) );
  NANDN U10762 ( .A(n9409), .B(n9410), .Z(n9161) );
  AND U10763 ( .A(n9162), .B(n9161), .Z(n9165) );
  XNOR U10764 ( .A(n9164), .B(n9163), .Z(n9166) );
  NANDN U10765 ( .A(n9165), .B(n9166), .Z(n9168) );
  AND U10766 ( .A(a[23]), .B(b[38]), .Z(n9535) );
  NANDN U10767 ( .A(n9535), .B(n9536), .Z(n9167) );
  NAND U10768 ( .A(n9168), .B(n9167), .Z(n9169) );
  NAND U10769 ( .A(n9170), .B(n9169), .Z(n9172) );
  NAND U10770 ( .A(a[24]), .B(b[38]), .Z(n9540) );
  XOR U10771 ( .A(n9170), .B(n9169), .Z(n9539) );
  NAND U10772 ( .A(n9540), .B(n9539), .Z(n9171) );
  NAND U10773 ( .A(n9172), .B(n9171), .Z(n9173) );
  NAND U10774 ( .A(n9174), .B(n9173), .Z(n9176) );
  AND U10775 ( .A(a[25]), .B(b[38]), .Z(n9543) );
  XOR U10776 ( .A(n9174), .B(n9173), .Z(n9544) );
  NANDN U10777 ( .A(n9543), .B(n9544), .Z(n9175) );
  NAND U10778 ( .A(n9176), .B(n9175), .Z(n9179) );
  NANDN U10779 ( .A(n9179), .B(n9180), .Z(n9182) );
  AND U10780 ( .A(a[26]), .B(b[38]), .Z(n9548) );
  NAND U10781 ( .A(n9548), .B(n9547), .Z(n9181) );
  AND U10782 ( .A(n9182), .B(n9181), .Z(n9186) );
  XNOR U10783 ( .A(n9184), .B(n9183), .Z(n9185) );
  NANDN U10784 ( .A(n9186), .B(n9185), .Z(n9188) );
  NAND U10785 ( .A(a[27]), .B(b[38]), .Z(n9407) );
  XNOR U10786 ( .A(n9186), .B(n9185), .Z(n9408) );
  NANDN U10787 ( .A(n9407), .B(n9408), .Z(n9187) );
  AND U10788 ( .A(n9188), .B(n9187), .Z(n9192) );
  XNOR U10789 ( .A(n9190), .B(n9189), .Z(n9191) );
  NANDN U10790 ( .A(n9192), .B(n9191), .Z(n9194) );
  NAND U10791 ( .A(a[28]), .B(b[38]), .Z(n9557) );
  XNOR U10792 ( .A(n9192), .B(n9191), .Z(n9558) );
  NANDN U10793 ( .A(n9557), .B(n9558), .Z(n9193) );
  AND U10794 ( .A(n9194), .B(n9193), .Z(n9198) );
  AND U10795 ( .A(a[29]), .B(b[38]), .Z(n9197) );
  NANDN U10796 ( .A(n9198), .B(n9197), .Z(n9200) );
  XOR U10797 ( .A(n9196), .B(n9195), .Z(n9563) );
  XNOR U10798 ( .A(n9198), .B(n9197), .Z(n9564) );
  NANDN U10799 ( .A(n9563), .B(n9564), .Z(n9199) );
  AND U10800 ( .A(n9200), .B(n9199), .Z(n9204) );
  AND U10801 ( .A(a[30]), .B(b[38]), .Z(n9203) );
  NANDN U10802 ( .A(n9204), .B(n9203), .Z(n9206) );
  XOR U10803 ( .A(n9202), .B(n9201), .Z(n9405) );
  XNOR U10804 ( .A(n9204), .B(n9203), .Z(n9406) );
  NANDN U10805 ( .A(n9405), .B(n9406), .Z(n9205) );
  AND U10806 ( .A(n9206), .B(n9205), .Z(n9210) );
  AND U10807 ( .A(a[31]), .B(b[38]), .Z(n9209) );
  NANDN U10808 ( .A(n9210), .B(n9209), .Z(n9212) );
  XOR U10809 ( .A(n9208), .B(n9207), .Z(n9573) );
  XNOR U10810 ( .A(n9210), .B(n9209), .Z(n9574) );
  NANDN U10811 ( .A(n9573), .B(n9574), .Z(n9211) );
  AND U10812 ( .A(n9212), .B(n9211), .Z(n9213) );
  NANDN U10813 ( .A(n9214), .B(n9213), .Z(n9218) );
  XOR U10814 ( .A(n9214), .B(n9213), .Z(n9579) );
  XOR U10815 ( .A(n9216), .B(n9215), .Z(n9580) );
  OR U10816 ( .A(n9579), .B(n9580), .Z(n9217) );
  NAND U10817 ( .A(n9218), .B(n9217), .Z(n9221) );
  XNOR U10818 ( .A(n9220), .B(n9219), .Z(n9222) );
  NANDN U10819 ( .A(n9221), .B(n9222), .Z(n9224) );
  NAND U10820 ( .A(a[33]), .B(b[38]), .Z(n9585) );
  XNOR U10821 ( .A(n9222), .B(n9221), .Z(n9586) );
  NANDN U10822 ( .A(n9585), .B(n9586), .Z(n9223) );
  AND U10823 ( .A(n9224), .B(n9223), .Z(n9228) );
  AND U10824 ( .A(a[34]), .B(b[38]), .Z(n9227) );
  NANDN U10825 ( .A(n9228), .B(n9227), .Z(n9230) );
  XOR U10826 ( .A(n9226), .B(n9225), .Z(n9403) );
  XNOR U10827 ( .A(n9228), .B(n9227), .Z(n9404) );
  NANDN U10828 ( .A(n9403), .B(n9404), .Z(n9229) );
  AND U10829 ( .A(n9230), .B(n9229), .Z(n9234) );
  AND U10830 ( .A(a[35]), .B(b[38]), .Z(n9233) );
  NANDN U10831 ( .A(n9234), .B(n9233), .Z(n9236) );
  XOR U10832 ( .A(n9232), .B(n9231), .Z(n9595) );
  XNOR U10833 ( .A(n9234), .B(n9233), .Z(n9596) );
  NANDN U10834 ( .A(n9595), .B(n9596), .Z(n9235) );
  AND U10835 ( .A(n9236), .B(n9235), .Z(n9240) );
  AND U10836 ( .A(a[36]), .B(b[38]), .Z(n9239) );
  NANDN U10837 ( .A(n9240), .B(n9239), .Z(n9242) );
  XOR U10838 ( .A(n9238), .B(n9237), .Z(n9601) );
  XNOR U10839 ( .A(n9240), .B(n9239), .Z(n9602) );
  NANDN U10840 ( .A(n9601), .B(n9602), .Z(n9241) );
  AND U10841 ( .A(n9242), .B(n9241), .Z(n9246) );
  XNOR U10842 ( .A(n9244), .B(n9243), .Z(n9245) );
  NANDN U10843 ( .A(n9246), .B(n9245), .Z(n9248) );
  NAND U10844 ( .A(a[37]), .B(b[38]), .Z(n9607) );
  XNOR U10845 ( .A(n9246), .B(n9245), .Z(n9608) );
  NANDN U10846 ( .A(n9607), .B(n9608), .Z(n9247) );
  AND U10847 ( .A(n9248), .B(n9247), .Z(n9249) );
  NANDN U10848 ( .A(n9250), .B(n9249), .Z(n9254) );
  XOR U10849 ( .A(n9250), .B(n9249), .Z(n9401) );
  XOR U10850 ( .A(n9252), .B(n9251), .Z(n9402) );
  OR U10851 ( .A(n9401), .B(n9402), .Z(n9253) );
  AND U10852 ( .A(n9254), .B(n9253), .Z(n9256) );
  NANDN U10853 ( .A(n9255), .B(n9256), .Z(n9260) );
  XNOR U10854 ( .A(n9256), .B(n9255), .Z(n9620) );
  XNOR U10855 ( .A(n9258), .B(n9257), .Z(n9619) );
  NAND U10856 ( .A(n9620), .B(n9619), .Z(n9259) );
  AND U10857 ( .A(n9260), .B(n9259), .Z(n9264) );
  AND U10858 ( .A(a[40]), .B(b[38]), .Z(n9263) );
  NANDN U10859 ( .A(n9264), .B(n9263), .Z(n9266) );
  XOR U10860 ( .A(n9262), .B(n9261), .Z(n9626) );
  XNOR U10861 ( .A(n9264), .B(n9263), .Z(n9625) );
  NANDN U10862 ( .A(n9626), .B(n9625), .Z(n9265) );
  AND U10863 ( .A(n9266), .B(n9265), .Z(n9270) );
  XNOR U10864 ( .A(n9268), .B(n9267), .Z(n9269) );
  NANDN U10865 ( .A(n9270), .B(n9269), .Z(n9272) );
  NAND U10866 ( .A(a[41]), .B(b[38]), .Z(n9629) );
  XNOR U10867 ( .A(n9270), .B(n9269), .Z(n9630) );
  NANDN U10868 ( .A(n9629), .B(n9630), .Z(n9271) );
  AND U10869 ( .A(n9272), .B(n9271), .Z(n9276) );
  XNOR U10870 ( .A(n9274), .B(n9273), .Z(n9275) );
  NANDN U10871 ( .A(n9276), .B(n9275), .Z(n9278) );
  XNOR U10872 ( .A(n9276), .B(n9275), .Z(n9638) );
  AND U10873 ( .A(a[42]), .B(b[38]), .Z(n9637) );
  NAND U10874 ( .A(n9638), .B(n9637), .Z(n9277) );
  AND U10875 ( .A(n9278), .B(n9277), .Z(n9279) );
  NANDN U10876 ( .A(n9280), .B(n9279), .Z(n9282) );
  XOR U10877 ( .A(n9280), .B(n9279), .Z(n9399) );
  AND U10878 ( .A(a[43]), .B(b[38]), .Z(n9400) );
  OR U10879 ( .A(n9399), .B(n9400), .Z(n9281) );
  AND U10880 ( .A(n9282), .B(n9281), .Z(n9286) );
  NANDN U10881 ( .A(n9285), .B(n9286), .Z(n9288) );
  XOR U10882 ( .A(n9284), .B(n9283), .Z(n9397) );
  XNOR U10883 ( .A(n9286), .B(n9285), .Z(n9398) );
  NANDN U10884 ( .A(n9397), .B(n9398), .Z(n9287) );
  AND U10885 ( .A(n9288), .B(n9287), .Z(n9289) );
  NANDN U10886 ( .A(n9290), .B(n9289), .Z(n9294) );
  XNOR U10887 ( .A(n9290), .B(n9289), .Z(n9396) );
  XNOR U10888 ( .A(n9292), .B(n9291), .Z(n9395) );
  NAND U10889 ( .A(n9396), .B(n9395), .Z(n9293) );
  AND U10890 ( .A(n9294), .B(n9293), .Z(n9298) );
  NANDN U10891 ( .A(n9297), .B(n9298), .Z(n9300) );
  XOR U10892 ( .A(n9296), .B(n9295), .Z(n9653) );
  XNOR U10893 ( .A(n9298), .B(n9297), .Z(n9654) );
  NANDN U10894 ( .A(n9653), .B(n9654), .Z(n9299) );
  AND U10895 ( .A(n9300), .B(n9299), .Z(n9304) );
  AND U10896 ( .A(a[47]), .B(b[38]), .Z(n9303) );
  NANDN U10897 ( .A(n9304), .B(n9303), .Z(n9306) );
  XOR U10898 ( .A(n9302), .B(n9301), .Z(n9659) );
  XNOR U10899 ( .A(n9304), .B(n9303), .Z(n9660) );
  NANDN U10900 ( .A(n9659), .B(n9660), .Z(n9305) );
  AND U10901 ( .A(n9306), .B(n9305), .Z(n9310) );
  XNOR U10902 ( .A(n9308), .B(n9307), .Z(n9309) );
  NANDN U10903 ( .A(n9310), .B(n9309), .Z(n9312) );
  NAND U10904 ( .A(a[48]), .B(b[38]), .Z(n9665) );
  XNOR U10905 ( .A(n9310), .B(n9309), .Z(n9666) );
  NANDN U10906 ( .A(n9665), .B(n9666), .Z(n9311) );
  AND U10907 ( .A(n9312), .B(n9311), .Z(n9316) );
  XNOR U10908 ( .A(n9314), .B(n9313), .Z(n9315) );
  NANDN U10909 ( .A(n9316), .B(n9315), .Z(n9318) );
  NAND U10910 ( .A(a[49]), .B(b[38]), .Z(n9671) );
  XNOR U10911 ( .A(n9316), .B(n9315), .Z(n9672) );
  NANDN U10912 ( .A(n9671), .B(n9672), .Z(n9317) );
  AND U10913 ( .A(n9318), .B(n9317), .Z(n9319) );
  NANDN U10914 ( .A(n9320), .B(n9319), .Z(n9324) );
  XOR U10915 ( .A(n9320), .B(n9319), .Z(n9393) );
  XOR U10916 ( .A(n9322), .B(n9321), .Z(n9394) );
  OR U10917 ( .A(n9393), .B(n9394), .Z(n9323) );
  NAND U10918 ( .A(n9324), .B(n9323), .Z(n9325) );
  NANDN U10919 ( .A(n9326), .B(n9325), .Z(n9330) );
  XOR U10920 ( .A(n9326), .B(n9325), .Z(n9391) );
  XOR U10921 ( .A(n9328), .B(n9327), .Z(n9392) );
  OR U10922 ( .A(n9391), .B(n9392), .Z(n9329) );
  AND U10923 ( .A(n9330), .B(n9329), .Z(n9334) );
  NANDN U10924 ( .A(n9333), .B(n9334), .Z(n9336) );
  XOR U10925 ( .A(n9332), .B(n9331), .Z(n9685) );
  XNOR U10926 ( .A(n9334), .B(n9333), .Z(n9686) );
  NANDN U10927 ( .A(n9685), .B(n9686), .Z(n9335) );
  AND U10928 ( .A(n9336), .B(n9335), .Z(n9340) );
  AND U10929 ( .A(a[53]), .B(b[38]), .Z(n9339) );
  NANDN U10930 ( .A(n9340), .B(n9339), .Z(n9342) );
  XOR U10931 ( .A(n9338), .B(n9337), .Z(n9691) );
  XNOR U10932 ( .A(n9340), .B(n9339), .Z(n9692) );
  NANDN U10933 ( .A(n9691), .B(n9692), .Z(n9341) );
  AND U10934 ( .A(n9342), .B(n9341), .Z(n9346) );
  XNOR U10935 ( .A(n9344), .B(n9343), .Z(n9345) );
  NANDN U10936 ( .A(n9346), .B(n9345), .Z(n9348) );
  NAND U10937 ( .A(a[54]), .B(b[38]), .Z(n9699) );
  XNOR U10938 ( .A(n9346), .B(n9345), .Z(n9700) );
  NANDN U10939 ( .A(n9699), .B(n9700), .Z(n9347) );
  AND U10940 ( .A(n9348), .B(n9347), .Z(n9352) );
  AND U10941 ( .A(a[55]), .B(b[38]), .Z(n9351) );
  NANDN U10942 ( .A(n9352), .B(n9351), .Z(n9354) );
  XOR U10943 ( .A(n9350), .B(n9349), .Z(n9706) );
  XNOR U10944 ( .A(n9352), .B(n9351), .Z(n9705) );
  NANDN U10945 ( .A(n9706), .B(n9705), .Z(n9353) );
  AND U10946 ( .A(n9354), .B(n9353), .Z(n9358) );
  AND U10947 ( .A(a[56]), .B(b[38]), .Z(n9357) );
  NANDN U10948 ( .A(n9358), .B(n9357), .Z(n9360) );
  XOR U10949 ( .A(n9356), .B(n9355), .Z(n9389) );
  XNOR U10950 ( .A(n9358), .B(n9357), .Z(n9390) );
  NANDN U10951 ( .A(n9389), .B(n9390), .Z(n9359) );
  AND U10952 ( .A(n9360), .B(n9359), .Z(n9361) );
  AND U10953 ( .A(a[57]), .B(b[38]), .Z(n9714) );
  XOR U10954 ( .A(n9362), .B(n9361), .Z(n9713) );
  AND U10955 ( .A(a[58]), .B(b[38]), .Z(n9388) );
  XOR U10956 ( .A(n9364), .B(n9363), .Z(n9387) );
  NANDN U10957 ( .A(n9367), .B(n9368), .Z(n9370) );
  NAND U10958 ( .A(a[59]), .B(b[38]), .Z(n9385) );
  NANDN U10959 ( .A(n9385), .B(n9386), .Z(n9369) );
  AND U10960 ( .A(n9370), .B(n9369), .Z(n9373) );
  XNOR U10961 ( .A(n9372), .B(n9371), .Z(n9374) );
  NAND U10962 ( .A(n9373), .B(n9374), .Z(n9376) );
  AND U10963 ( .A(a[60]), .B(b[38]), .Z(n9723) );
  XOR U10964 ( .A(n9374), .B(n9373), .Z(n9724) );
  NANDN U10965 ( .A(n9723), .B(n9724), .Z(n9375) );
  NAND U10966 ( .A(n9376), .B(n9375), .Z(n9379) );
  NANDN U10967 ( .A(n9379), .B(n9380), .Z(n9382) );
  NAND U10968 ( .A(a[61]), .B(b[38]), .Z(n9383) );
  NANDN U10969 ( .A(n9383), .B(n9384), .Z(n9381) );
  AND U10970 ( .A(n9382), .B(n9381), .Z(n10251) );
  XOR U10971 ( .A(n10250), .B(n10251), .Z(n10252) );
  NAND U10972 ( .A(a[62]), .B(b[37]), .Z(n9729) );
  NANDN U10973 ( .A(n9729), .B(n9730), .Z(n9732) );
  NAND U10974 ( .A(a[60]), .B(b[37]), .Z(n9719) );
  NANDN U10975 ( .A(n9719), .B(n9720), .Z(n9722) );
  XOR U10976 ( .A(n9388), .B(n9387), .Z(n9718) );
  NAND U10977 ( .A(a[57]), .B(b[37]), .Z(n9709) );
  XNOR U10978 ( .A(n9390), .B(n9389), .Z(n9710) );
  NANDN U10979 ( .A(n9709), .B(n9710), .Z(n9712) );
  XOR U10980 ( .A(n9392), .B(n9391), .Z(n9682) );
  AND U10981 ( .A(a[52]), .B(b[37]), .Z(n9681) );
  NANDN U10982 ( .A(n9682), .B(n9681), .Z(n9684) );
  XOR U10983 ( .A(n9394), .B(n9393), .Z(n9678) );
  AND U10984 ( .A(a[51]), .B(b[37]), .Z(n9677) );
  NANDN U10985 ( .A(n9678), .B(n9677), .Z(n9680) );
  XOR U10986 ( .A(n9396), .B(n9395), .Z(n9650) );
  AND U10987 ( .A(a[46]), .B(b[37]), .Z(n9649) );
  NANDN U10988 ( .A(n9650), .B(n9649), .Z(n9652) );
  NAND U10989 ( .A(a[45]), .B(b[37]), .Z(n9645) );
  XNOR U10990 ( .A(n9398), .B(n9397), .Z(n9646) );
  NANDN U10991 ( .A(n9645), .B(n9646), .Z(n9648) );
  XOR U10992 ( .A(n9400), .B(n9399), .Z(n9642) );
  AND U10993 ( .A(a[43]), .B(b[37]), .Z(n9636) );
  NAND U10994 ( .A(a[41]), .B(b[37]), .Z(n9623) );
  AND U10995 ( .A(a[40]), .B(b[37]), .Z(n9618) );
  XOR U10996 ( .A(n9402), .B(n9401), .Z(n9614) );
  AND U10997 ( .A(a[39]), .B(b[37]), .Z(n9613) );
  NANDN U10998 ( .A(n9614), .B(n9613), .Z(n9616) );
  NAND U10999 ( .A(a[35]), .B(b[37]), .Z(n9591) );
  XNOR U11000 ( .A(n9404), .B(n9403), .Z(n9592) );
  NANDN U11001 ( .A(n9591), .B(n9592), .Z(n9594) );
  NAND U11002 ( .A(a[31]), .B(b[37]), .Z(n9569) );
  XNOR U11003 ( .A(n9406), .B(n9405), .Z(n9570) );
  NANDN U11004 ( .A(n9569), .B(n9570), .Z(n9572) );
  NAND U11005 ( .A(a[28]), .B(b[37]), .Z(n9553) );
  XNOR U11006 ( .A(n9408), .B(n9407), .Z(n9554) );
  NANDN U11007 ( .A(n9553), .B(n9554), .Z(n9556) );
  AND U11008 ( .A(a[27]), .B(b[37]), .Z(n9549) );
  NAND U11009 ( .A(a[26]), .B(b[37]), .Z(n9541) );
  AND U11010 ( .A(a[14]), .B(b[37]), .Z(n9488) );
  NAND U11011 ( .A(n9488), .B(n9487), .Z(n9490) );
  NAND U11012 ( .A(a[13]), .B(b[37]), .Z(n9483) );
  NANDN U11013 ( .A(n9483), .B(n9484), .Z(n9486) );
  NAND U11014 ( .A(a[12]), .B(b[37]), .Z(n9479) );
  NANDN U11015 ( .A(n9479), .B(n9480), .Z(n9482) );
  NAND U11016 ( .A(a[11]), .B(b[37]), .Z(n9475) );
  XOR U11017 ( .A(n9420), .B(n9419), .Z(n9476) );
  NANDN U11018 ( .A(n9475), .B(n9476), .Z(n9478) );
  XOR U11019 ( .A(n9422), .B(n9421), .Z(n9471) );
  AND U11020 ( .A(a[10]), .B(b[37]), .Z(n9472) );
  NANDN U11021 ( .A(n9471), .B(n9472), .Z(n9474) );
  NAND U11022 ( .A(a[5]), .B(b[37]), .Z(n9445) );
  XOR U11023 ( .A(n9426), .B(n9425), .Z(n9446) );
  NANDN U11024 ( .A(n9445), .B(n9446), .Z(n9448) );
  NAND U11025 ( .A(a[3]), .B(b[37]), .Z(n9435) );
  XNOR U11026 ( .A(n9428), .B(n9427), .Z(n9436) );
  NANDN U11027 ( .A(n9435), .B(n9436), .Z(n9438) );
  AND U11028 ( .A(a[0]), .B(b[37]), .Z(n10279) );
  AND U11029 ( .A(a[1]), .B(b[38]), .Z(n9432) );
  AND U11030 ( .A(n10279), .B(n9432), .Z(n9430) );
  NANDN U11031 ( .A(n9050), .B(n9430), .Z(n9434) );
  AND U11032 ( .A(a[2]), .B(b[37]), .Z(n9781) );
  NANDN U11033 ( .A(n9780), .B(n9781), .Z(n9433) );
  AND U11034 ( .A(n9434), .B(n9433), .Z(n9786) );
  NANDN U11035 ( .A(n9786), .B(n9787), .Z(n9437) );
  AND U11036 ( .A(n9438), .B(n9437), .Z(n9441) );
  AND U11037 ( .A(a[4]), .B(b[37]), .Z(n9442) );
  NANDN U11038 ( .A(n9441), .B(n9442), .Z(n9444) );
  NAND U11039 ( .A(n9793), .B(n9792), .Z(n9443) );
  AND U11040 ( .A(n9444), .B(n9443), .Z(n9798) );
  NANDN U11041 ( .A(n9798), .B(n9799), .Z(n9447) );
  AND U11042 ( .A(n9448), .B(n9447), .Z(n9451) );
  AND U11043 ( .A(a[6]), .B(b[37]), .Z(n9452) );
  NANDN U11044 ( .A(n9451), .B(n9452), .Z(n9454) );
  XOR U11045 ( .A(n9450), .B(n9449), .Z(n9805) );
  NAND U11046 ( .A(n9805), .B(n9804), .Z(n9453) );
  AND U11047 ( .A(n9454), .B(n9453), .Z(n9457) );
  NANDN U11048 ( .A(n9457), .B(n9458), .Z(n9460) );
  NAND U11049 ( .A(a[7]), .B(b[37]), .Z(n9810) );
  NANDN U11050 ( .A(n9810), .B(n9811), .Z(n9459) );
  AND U11051 ( .A(n9460), .B(n9459), .Z(n9461) );
  AND U11052 ( .A(a[8]), .B(b[37]), .Z(n9462) );
  NANDN U11053 ( .A(n9461), .B(n9462), .Z(n9466) );
  XOR U11054 ( .A(n9464), .B(n9463), .Z(n9816) );
  NAND U11055 ( .A(n9817), .B(n9816), .Z(n9465) );
  NAND U11056 ( .A(n9466), .B(n9465), .Z(n9467) );
  NAND U11057 ( .A(n9468), .B(n9467), .Z(n9470) );
  NAND U11058 ( .A(a[9]), .B(b[37]), .Z(n9822) );
  XOR U11059 ( .A(n9468), .B(n9467), .Z(n9823) );
  NANDN U11060 ( .A(n9822), .B(n9823), .Z(n9469) );
  AND U11061 ( .A(n9470), .B(n9469), .Z(n9828) );
  NANDN U11062 ( .A(n9828), .B(n9829), .Z(n9473) );
  AND U11063 ( .A(n9474), .B(n9473), .Z(n9834) );
  NANDN U11064 ( .A(n9834), .B(n9835), .Z(n9477) );
  AND U11065 ( .A(n9478), .B(n9477), .Z(n9840) );
  NANDN U11066 ( .A(n9840), .B(n9841), .Z(n9481) );
  AND U11067 ( .A(n9482), .B(n9481), .Z(n9848) );
  NANDN U11068 ( .A(n9848), .B(n9849), .Z(n9485) );
  AND U11069 ( .A(n9486), .B(n9485), .Z(n9854) );
  XOR U11070 ( .A(n9488), .B(n9487), .Z(n9855) );
  NANDN U11071 ( .A(n9854), .B(n9855), .Z(n9489) );
  AND U11072 ( .A(n9490), .B(n9489), .Z(n9493) );
  NANDN U11073 ( .A(n9493), .B(n9494), .Z(n9496) );
  AND U11074 ( .A(a[15]), .B(b[37]), .Z(n9861) );
  NAND U11075 ( .A(n9861), .B(n9860), .Z(n9495) );
  AND U11076 ( .A(n9496), .B(n9495), .Z(n9499) );
  AND U11077 ( .A(a[16]), .B(b[37]), .Z(n9500) );
  NANDN U11078 ( .A(n9499), .B(n9500), .Z(n9502) );
  NAND U11079 ( .A(n9771), .B(n9770), .Z(n9501) );
  AND U11080 ( .A(n9502), .B(n9501), .Z(n9505) );
  XOR U11081 ( .A(n9504), .B(n9503), .Z(n9506) );
  NANDN U11082 ( .A(n9505), .B(n9506), .Z(n9508) );
  NAND U11083 ( .A(a[17]), .B(b[37]), .Z(n9868) );
  NANDN U11084 ( .A(n9868), .B(n9869), .Z(n9507) );
  AND U11085 ( .A(n9508), .B(n9507), .Z(n9509) );
  AND U11086 ( .A(a[18]), .B(b[37]), .Z(n9510) );
  NANDN U11087 ( .A(n9509), .B(n9510), .Z(n9514) );
  NAND U11088 ( .A(n9874), .B(n9875), .Z(n9513) );
  AND U11089 ( .A(n9514), .B(n9513), .Z(n9517) );
  NANDN U11090 ( .A(n9517), .B(n9518), .Z(n9520) );
  AND U11091 ( .A(a[19]), .B(b[37]), .Z(n9881) );
  NAND U11092 ( .A(n9881), .B(n9880), .Z(n9519) );
  AND U11093 ( .A(n9520), .B(n9519), .Z(n9521) );
  AND U11094 ( .A(a[20]), .B(b[37]), .Z(n9522) );
  NANDN U11095 ( .A(n9521), .B(n9522), .Z(n9526) );
  NAND U11096 ( .A(n9886), .B(n9887), .Z(n9525) );
  NAND U11097 ( .A(n9526), .B(n9525), .Z(n9893) );
  NAND U11098 ( .A(a[21]), .B(b[37]), .Z(n9894) );
  AND U11099 ( .A(a[22]), .B(b[37]), .Z(n9527) );
  NANDN U11100 ( .A(n9528), .B(n9527), .Z(n9532) );
  XNOR U11101 ( .A(n9528), .B(n9527), .Z(n9899) );
  NAND U11102 ( .A(n9899), .B(n9900), .Z(n9531) );
  NAND U11103 ( .A(n9532), .B(n9531), .Z(n9906) );
  NAND U11104 ( .A(a[23]), .B(b[37]), .Z(n9907) );
  AND U11105 ( .A(a[24]), .B(b[37]), .Z(n9533) );
  NANDN U11106 ( .A(n9534), .B(n9533), .Z(n9538) );
  XNOR U11107 ( .A(n9534), .B(n9533), .Z(n9912) );
  NAND U11108 ( .A(n9912), .B(n9913), .Z(n9537) );
  NAND U11109 ( .A(n9538), .B(n9537), .Z(n9769) );
  XOR U11110 ( .A(n9540), .B(n9539), .Z(n9768) );
  NAND U11111 ( .A(a[25]), .B(b[37]), .Z(n9767) );
  NANDN U11112 ( .A(n9541), .B(n9542), .Z(n9546) );
  NAND U11113 ( .A(n9918), .B(n9919), .Z(n9545) );
  AND U11114 ( .A(n9546), .B(n9545), .Z(n9550) );
  NANDN U11115 ( .A(n9549), .B(n9550), .Z(n9552) );
  XOR U11116 ( .A(n9548), .B(n9547), .Z(n9926) );
  NANDN U11117 ( .A(n9926), .B(n9927), .Z(n9551) );
  NAND U11118 ( .A(n9552), .B(n9551), .Z(n9932) );
  XNOR U11119 ( .A(n9554), .B(n9553), .Z(n9933) );
  NANDN U11120 ( .A(n9932), .B(n9933), .Z(n9555) );
  AND U11121 ( .A(n9556), .B(n9555), .Z(n9560) );
  AND U11122 ( .A(a[29]), .B(b[37]), .Z(n9559) );
  NANDN U11123 ( .A(n9560), .B(n9559), .Z(n9562) );
  XOR U11124 ( .A(n9558), .B(n9557), .Z(n9938) );
  XNOR U11125 ( .A(n9560), .B(n9559), .Z(n9939) );
  NANDN U11126 ( .A(n9938), .B(n9939), .Z(n9561) );
  AND U11127 ( .A(n9562), .B(n9561), .Z(n9566) );
  XNOR U11128 ( .A(n9564), .B(n9563), .Z(n9565) );
  NANDN U11129 ( .A(n9566), .B(n9565), .Z(n9568) );
  NAND U11130 ( .A(a[30]), .B(b[37]), .Z(n9942) );
  XNOR U11131 ( .A(n9566), .B(n9565), .Z(n9943) );
  NANDN U11132 ( .A(n9942), .B(n9943), .Z(n9567) );
  AND U11133 ( .A(n9568), .B(n9567), .Z(n9764) );
  XNOR U11134 ( .A(n9570), .B(n9569), .Z(n9763) );
  NANDN U11135 ( .A(n9764), .B(n9763), .Z(n9571) );
  AND U11136 ( .A(n9572), .B(n9571), .Z(n9576) );
  AND U11137 ( .A(a[32]), .B(b[37]), .Z(n9575) );
  NANDN U11138 ( .A(n9576), .B(n9575), .Z(n9578) );
  XOR U11139 ( .A(n9574), .B(n9573), .Z(n9950) );
  XNOR U11140 ( .A(n9576), .B(n9575), .Z(n9951) );
  NANDN U11141 ( .A(n9950), .B(n9951), .Z(n9577) );
  AND U11142 ( .A(n9578), .B(n9577), .Z(n9582) );
  AND U11143 ( .A(a[33]), .B(b[37]), .Z(n9581) );
  NANDN U11144 ( .A(n9582), .B(n9581), .Z(n9584) );
  XOR U11145 ( .A(n9580), .B(n9579), .Z(n9957) );
  XNOR U11146 ( .A(n9582), .B(n9581), .Z(n9956) );
  NANDN U11147 ( .A(n9957), .B(n9956), .Z(n9583) );
  AND U11148 ( .A(n9584), .B(n9583), .Z(n9588) );
  XNOR U11149 ( .A(n9586), .B(n9585), .Z(n9587) );
  NANDN U11150 ( .A(n9588), .B(n9587), .Z(n9590) );
  NAND U11151 ( .A(a[34]), .B(b[37]), .Z(n9761) );
  XNOR U11152 ( .A(n9588), .B(n9587), .Z(n9762) );
  NANDN U11153 ( .A(n9761), .B(n9762), .Z(n9589) );
  AND U11154 ( .A(n9590), .B(n9589), .Z(n9969) );
  XNOR U11155 ( .A(n9592), .B(n9591), .Z(n9968) );
  NANDN U11156 ( .A(n9969), .B(n9968), .Z(n9593) );
  AND U11157 ( .A(n9594), .B(n9593), .Z(n9598) );
  AND U11158 ( .A(a[36]), .B(b[37]), .Z(n9597) );
  NANDN U11159 ( .A(n9598), .B(n9597), .Z(n9600) );
  XOR U11160 ( .A(n9596), .B(n9595), .Z(n9972) );
  XNOR U11161 ( .A(n9598), .B(n9597), .Z(n9973) );
  NANDN U11162 ( .A(n9972), .B(n9973), .Z(n9599) );
  AND U11163 ( .A(n9600), .B(n9599), .Z(n9604) );
  AND U11164 ( .A(a[37]), .B(b[37]), .Z(n9603) );
  NANDN U11165 ( .A(n9604), .B(n9603), .Z(n9606) );
  XOR U11166 ( .A(n9602), .B(n9601), .Z(n9757) );
  XNOR U11167 ( .A(n9604), .B(n9603), .Z(n9758) );
  NANDN U11168 ( .A(n9757), .B(n9758), .Z(n9605) );
  AND U11169 ( .A(n9606), .B(n9605), .Z(n9610) );
  XNOR U11170 ( .A(n9608), .B(n9607), .Z(n9609) );
  NANDN U11171 ( .A(n9610), .B(n9609), .Z(n9612) );
  NAND U11172 ( .A(a[38]), .B(b[37]), .Z(n9982) );
  XNOR U11173 ( .A(n9610), .B(n9609), .Z(n9983) );
  NANDN U11174 ( .A(n9982), .B(n9983), .Z(n9611) );
  AND U11175 ( .A(n9612), .B(n9611), .Z(n9754) );
  XNOR U11176 ( .A(n9614), .B(n9613), .Z(n9753) );
  NANDN U11177 ( .A(n9754), .B(n9753), .Z(n9615) );
  AND U11178 ( .A(n9616), .B(n9615), .Z(n9617) );
  NANDN U11179 ( .A(n9618), .B(n9617), .Z(n9622) );
  XOR U11180 ( .A(n9618), .B(n9617), .Z(n9988) );
  XOR U11181 ( .A(n9620), .B(n9619), .Z(n9989) );
  OR U11182 ( .A(n9988), .B(n9989), .Z(n9621) );
  AND U11183 ( .A(n9622), .B(n9621), .Z(n9624) );
  NANDN U11184 ( .A(n9623), .B(n9624), .Z(n9628) );
  XOR U11185 ( .A(n9624), .B(n9623), .Z(n9994) );
  XNOR U11186 ( .A(n9626), .B(n9625), .Z(n9995) );
  NANDN U11187 ( .A(n9994), .B(n9995), .Z(n9627) );
  AND U11188 ( .A(n9628), .B(n9627), .Z(n9632) );
  XNOR U11189 ( .A(n9630), .B(n9629), .Z(n9631) );
  NANDN U11190 ( .A(n9632), .B(n9631), .Z(n9634) );
  NAND U11191 ( .A(a[42]), .B(b[37]), .Z(n10000) );
  XNOR U11192 ( .A(n9632), .B(n9631), .Z(n10001) );
  NANDN U11193 ( .A(n10000), .B(n10001), .Z(n9633) );
  AND U11194 ( .A(n9634), .B(n9633), .Z(n9635) );
  NANDN U11195 ( .A(n9636), .B(n9635), .Z(n9640) );
  XOR U11196 ( .A(n9636), .B(n9635), .Z(n9751) );
  XOR U11197 ( .A(n9638), .B(n9637), .Z(n9752) );
  OR U11198 ( .A(n9751), .B(n9752), .Z(n9639) );
  AND U11199 ( .A(n9640), .B(n9639), .Z(n9641) );
  NANDN U11200 ( .A(n9642), .B(n9641), .Z(n9644) );
  NAND U11201 ( .A(a[44]), .B(b[37]), .Z(n9747) );
  XNOR U11202 ( .A(n9642), .B(n9641), .Z(n9748) );
  NANDN U11203 ( .A(n9747), .B(n9748), .Z(n9643) );
  AND U11204 ( .A(n9644), .B(n9643), .Z(n10015) );
  XNOR U11205 ( .A(n9646), .B(n9645), .Z(n10014) );
  NANDN U11206 ( .A(n10015), .B(n10014), .Z(n9647) );
  AND U11207 ( .A(n9648), .B(n9647), .Z(n10019) );
  XNOR U11208 ( .A(n9650), .B(n9649), .Z(n10018) );
  NANDN U11209 ( .A(n10019), .B(n10018), .Z(n9651) );
  AND U11210 ( .A(n9652), .B(n9651), .Z(n9656) );
  XNOR U11211 ( .A(n9654), .B(n9653), .Z(n9655) );
  NANDN U11212 ( .A(n9656), .B(n9655), .Z(n9658) );
  NAND U11213 ( .A(a[47]), .B(b[37]), .Z(n10024) );
  XNOR U11214 ( .A(n9656), .B(n9655), .Z(n10025) );
  NANDN U11215 ( .A(n10024), .B(n10025), .Z(n9657) );
  AND U11216 ( .A(n9658), .B(n9657), .Z(n9662) );
  AND U11217 ( .A(a[48]), .B(b[37]), .Z(n9661) );
  NANDN U11218 ( .A(n9662), .B(n9661), .Z(n9664) );
  XOR U11219 ( .A(n9660), .B(n9659), .Z(n10030) );
  XNOR U11220 ( .A(n9662), .B(n9661), .Z(n10031) );
  NANDN U11221 ( .A(n10030), .B(n10031), .Z(n9663) );
  AND U11222 ( .A(n9664), .B(n9663), .Z(n9668) );
  XNOR U11223 ( .A(n9666), .B(n9665), .Z(n9667) );
  NANDN U11224 ( .A(n9668), .B(n9667), .Z(n9670) );
  NAND U11225 ( .A(a[49]), .B(b[37]), .Z(n9743) );
  XNOR U11226 ( .A(n9668), .B(n9667), .Z(n9744) );
  NANDN U11227 ( .A(n9743), .B(n9744), .Z(n9669) );
  AND U11228 ( .A(n9670), .B(n9669), .Z(n9674) );
  AND U11229 ( .A(a[50]), .B(b[37]), .Z(n9673) );
  NANDN U11230 ( .A(n9674), .B(n9673), .Z(n9676) );
  XOR U11231 ( .A(n9672), .B(n9671), .Z(n10038) );
  XNOR U11232 ( .A(n9674), .B(n9673), .Z(n10039) );
  NANDN U11233 ( .A(n10038), .B(n10039), .Z(n9675) );
  AND U11234 ( .A(n9676), .B(n9675), .Z(n10045) );
  XNOR U11235 ( .A(n9678), .B(n9677), .Z(n10044) );
  NANDN U11236 ( .A(n10045), .B(n10044), .Z(n9679) );
  AND U11237 ( .A(n9680), .B(n9679), .Z(n9742) );
  XNOR U11238 ( .A(n9682), .B(n9681), .Z(n9741) );
  NANDN U11239 ( .A(n9742), .B(n9741), .Z(n9683) );
  AND U11240 ( .A(n9684), .B(n9683), .Z(n9688) );
  XNOR U11241 ( .A(n9686), .B(n9685), .Z(n9687) );
  NANDN U11242 ( .A(n9688), .B(n9687), .Z(n9690) );
  NAND U11243 ( .A(a[53]), .B(b[37]), .Z(n10056) );
  XNOR U11244 ( .A(n9688), .B(n9687), .Z(n10057) );
  NANDN U11245 ( .A(n10056), .B(n10057), .Z(n9689) );
  AND U11246 ( .A(n9690), .B(n9689), .Z(n9694) );
  XNOR U11247 ( .A(n9692), .B(n9691), .Z(n9693) );
  NANDN U11248 ( .A(n9694), .B(n9693), .Z(n9696) );
  NAND U11249 ( .A(a[54]), .B(b[37]), .Z(n9737) );
  XNOR U11250 ( .A(n9694), .B(n9693), .Z(n9738) );
  NANDN U11251 ( .A(n9737), .B(n9738), .Z(n9695) );
  AND U11252 ( .A(n9696), .B(n9695), .Z(n9698) );
  AND U11253 ( .A(a[55]), .B(b[37]), .Z(n9697) );
  NANDN U11254 ( .A(n9698), .B(n9697), .Z(n9702) );
  XOR U11255 ( .A(n9698), .B(n9697), .Z(n10062) );
  XNOR U11256 ( .A(n9700), .B(n9699), .Z(n10063) );
  NANDN U11257 ( .A(n10062), .B(n10063), .Z(n9701) );
  AND U11258 ( .A(n9702), .B(n9701), .Z(n9704) );
  AND U11259 ( .A(a[56]), .B(b[37]), .Z(n9703) );
  NANDN U11260 ( .A(n9704), .B(n9703), .Z(n9708) );
  XOR U11261 ( .A(n9704), .B(n9703), .Z(n10068) );
  XNOR U11262 ( .A(n9706), .B(n9705), .Z(n10069) );
  NANDN U11263 ( .A(n10068), .B(n10069), .Z(n9707) );
  AND U11264 ( .A(n9708), .B(n9707), .Z(n9736) );
  XNOR U11265 ( .A(n9710), .B(n9709), .Z(n9735) );
  NANDN U11266 ( .A(n9736), .B(n9735), .Z(n9711) );
  AND U11267 ( .A(n9712), .B(n9711), .Z(n9716) );
  AND U11268 ( .A(a[58]), .B(b[37]), .Z(n9715) );
  XOR U11269 ( .A(n9714), .B(n9713), .Z(n10079) );
  XNOR U11270 ( .A(n9716), .B(n9715), .Z(n10078) );
  NAND U11271 ( .A(a[59]), .B(b[37]), .Z(n10084) );
  XOR U11272 ( .A(n9718), .B(n9717), .Z(n10085) );
  XNOR U11273 ( .A(n9720), .B(n9719), .Z(n10092) );
  NANDN U11274 ( .A(n10093), .B(n10092), .Z(n9721) );
  AND U11275 ( .A(n9722), .B(n9721), .Z(n9726) );
  NAND U11276 ( .A(n9726), .B(n9725), .Z(n9728) );
  AND U11277 ( .A(a[61]), .B(b[37]), .Z(n9733) );
  XOR U11278 ( .A(n9726), .B(n9725), .Z(n9734) );
  NANDN U11279 ( .A(n9733), .B(n9734), .Z(n9727) );
  NAND U11280 ( .A(n9728), .B(n9727), .Z(n10100) );
  NANDN U11281 ( .A(n10100), .B(n10101), .Z(n9731) );
  AND U11282 ( .A(n9732), .B(n9731), .Z(n10257) );
  AND U11283 ( .A(a[63]), .B(b[37]), .Z(n10256) );
  XOR U11284 ( .A(n10258), .B(n10259), .Z(n10643) );
  NAND U11285 ( .A(a[58]), .B(b[36]), .Z(n10074) );
  XNOR U11286 ( .A(n9736), .B(n9735), .Z(n10075) );
  NANDN U11287 ( .A(n10074), .B(n10075), .Z(n10077) );
  NAND U11288 ( .A(a[55]), .B(b[36]), .Z(n9739) );
  XNOR U11289 ( .A(n9738), .B(n9737), .Z(n9740) );
  NANDN U11290 ( .A(n9739), .B(n9740), .Z(n10061) );
  XOR U11291 ( .A(n9740), .B(n9739), .Z(n10597) );
  NAND U11292 ( .A(a[53]), .B(b[36]), .Z(n10050) );
  XNOR U11293 ( .A(n9742), .B(n9741), .Z(n10051) );
  NANDN U11294 ( .A(n10050), .B(n10051), .Z(n10053) );
  NAND U11295 ( .A(a[50]), .B(b[36]), .Z(n9745) );
  XNOR U11296 ( .A(n9744), .B(n9743), .Z(n9746) );
  NANDN U11297 ( .A(n9745), .B(n9746), .Z(n10037) );
  XOR U11298 ( .A(n9746), .B(n9745), .Z(n10567) );
  NAND U11299 ( .A(a[45]), .B(b[36]), .Z(n9749) );
  XNOR U11300 ( .A(n9748), .B(n9747), .Z(n9750) );
  NANDN U11301 ( .A(n9749), .B(n9750), .Z(n10011) );
  XOR U11302 ( .A(n9750), .B(n9749), .Z(n10537) );
  XOR U11303 ( .A(n9752), .B(n9751), .Z(n10007) );
  NAND U11304 ( .A(a[40]), .B(b[36]), .Z(n9755) );
  XNOR U11305 ( .A(n9754), .B(n9753), .Z(n9756) );
  NANDN U11306 ( .A(n9755), .B(n9756), .Z(n9987) );
  XOR U11307 ( .A(n9756), .B(n9755), .Z(n10507) );
  NAND U11308 ( .A(a[38]), .B(b[36]), .Z(n9759) );
  XNOR U11309 ( .A(n9758), .B(n9757), .Z(n9760) );
  NANDN U11310 ( .A(n9759), .B(n9760), .Z(n9979) );
  XOR U11311 ( .A(n9760), .B(n9759), .Z(n10495) );
  NAND U11312 ( .A(a[35]), .B(b[36]), .Z(n9962) );
  XNOR U11313 ( .A(n9762), .B(n9761), .Z(n9963) );
  NANDN U11314 ( .A(n9962), .B(n9963), .Z(n9965) );
  NAND U11315 ( .A(a[32]), .B(b[36]), .Z(n9765) );
  XNOR U11316 ( .A(n9764), .B(n9763), .Z(n9766) );
  NANDN U11317 ( .A(n9765), .B(n9766), .Z(n9949) );
  XOR U11318 ( .A(n9766), .B(n9765), .Z(n10459) );
  NAND U11319 ( .A(a[28]), .B(b[36]), .Z(n9924) );
  XOR U11320 ( .A(n9771), .B(n9770), .Z(n9864) );
  NAND U11321 ( .A(a[12]), .B(b[36]), .Z(n9836) );
  AND U11322 ( .A(a[0]), .B(b[36]), .Z(n10725) );
  AND U11323 ( .A(a[1]), .B(b[37]), .Z(n9775) );
  AND U11324 ( .A(n10725), .B(n9775), .Z(n9772) );
  NAND U11325 ( .A(a[2]), .B(n9772), .Z(n9779) );
  NAND U11326 ( .A(b[37]), .B(a[1]), .Z(n9773) );
  XOR U11327 ( .A(n9774), .B(n9773), .Z(n10284) );
  NAND U11328 ( .A(n9775), .B(a[0]), .Z(n9776) );
  XNOR U11329 ( .A(a[2]), .B(n9776), .Z(n9777) );
  AND U11330 ( .A(b[36]), .B(n9777), .Z(n10285) );
  NANDN U11331 ( .A(n10284), .B(n10285), .Z(n9778) );
  AND U11332 ( .A(n9779), .B(n9778), .Z(n9782) );
  XNOR U11333 ( .A(n9781), .B(n9780), .Z(n9783) );
  NANDN U11334 ( .A(n9782), .B(n9783), .Z(n9785) );
  NAND U11335 ( .A(a[3]), .B(b[36]), .Z(n10288) );
  NANDN U11336 ( .A(n10288), .B(n10289), .Z(n9784) );
  AND U11337 ( .A(n9785), .B(n9784), .Z(n9788) );
  AND U11338 ( .A(a[4]), .B(b[36]), .Z(n9789) );
  NANDN U11339 ( .A(n9788), .B(n9789), .Z(n9791) );
  NAND U11340 ( .A(n10295), .B(n10294), .Z(n9790) );
  AND U11341 ( .A(n9791), .B(n9790), .Z(n9794) );
  XOR U11342 ( .A(n9793), .B(n9792), .Z(n9795) );
  NANDN U11343 ( .A(n9794), .B(n9795), .Z(n9797) );
  NAND U11344 ( .A(a[5]), .B(b[36]), .Z(n10300) );
  NANDN U11345 ( .A(n10300), .B(n10301), .Z(n9796) );
  AND U11346 ( .A(n9797), .B(n9796), .Z(n9800) );
  AND U11347 ( .A(a[6]), .B(b[36]), .Z(n9801) );
  NANDN U11348 ( .A(n9800), .B(n9801), .Z(n9803) );
  NAND U11349 ( .A(n10307), .B(n10306), .Z(n9802) );
  AND U11350 ( .A(n9803), .B(n9802), .Z(n9806) );
  XOR U11351 ( .A(n9805), .B(n9804), .Z(n9807) );
  NANDN U11352 ( .A(n9806), .B(n9807), .Z(n9809) );
  AND U11353 ( .A(a[7]), .B(b[36]), .Z(n10313) );
  NAND U11354 ( .A(n10313), .B(n10312), .Z(n9808) );
  AND U11355 ( .A(n9809), .B(n9808), .Z(n9812) );
  NANDN U11356 ( .A(n9812), .B(n9813), .Z(n9815) );
  NAND U11357 ( .A(a[8]), .B(b[36]), .Z(n10318) );
  NANDN U11358 ( .A(n10318), .B(n10319), .Z(n9814) );
  AND U11359 ( .A(n9815), .B(n9814), .Z(n9818) );
  XOR U11360 ( .A(n9817), .B(n9816), .Z(n9819) );
  NANDN U11361 ( .A(n9818), .B(n9819), .Z(n9821) );
  NAND U11362 ( .A(a[9]), .B(b[36]), .Z(n10324) );
  NANDN U11363 ( .A(n10324), .B(n10325), .Z(n9820) );
  AND U11364 ( .A(n9821), .B(n9820), .Z(n9824) );
  NANDN U11365 ( .A(n9824), .B(n9825), .Z(n9827) );
  NAND U11366 ( .A(a[10]), .B(b[36]), .Z(n10332) );
  NANDN U11367 ( .A(n10332), .B(n10333), .Z(n9826) );
  AND U11368 ( .A(n9827), .B(n9826), .Z(n9831) );
  NAND U11369 ( .A(n9831), .B(n9830), .Z(n9833) );
  XOR U11370 ( .A(n9831), .B(n9830), .Z(n10337) );
  NAND U11371 ( .A(a[11]), .B(b[36]), .Z(n10336) );
  NAND U11372 ( .A(n10337), .B(n10336), .Z(n9832) );
  AND U11373 ( .A(n9833), .B(n9832), .Z(n9837) );
  NANDN U11374 ( .A(n9836), .B(n9837), .Z(n9839) );
  NAND U11375 ( .A(n10343), .B(n10342), .Z(n9838) );
  AND U11376 ( .A(n9839), .B(n9838), .Z(n9842) );
  NANDN U11377 ( .A(n9842), .B(n9843), .Z(n9845) );
  AND U11378 ( .A(a[13]), .B(b[36]), .Z(n10349) );
  NAND U11379 ( .A(n10349), .B(n10348), .Z(n9844) );
  AND U11380 ( .A(n9845), .B(n9844), .Z(n9846) );
  AND U11381 ( .A(a[14]), .B(b[36]), .Z(n9847) );
  NANDN U11382 ( .A(n9846), .B(n9847), .Z(n9851) );
  NAND U11383 ( .A(n10355), .B(n10354), .Z(n9850) );
  AND U11384 ( .A(n9851), .B(n9850), .Z(n9852) );
  AND U11385 ( .A(a[15]), .B(b[36]), .Z(n9853) );
  NANDN U11386 ( .A(n9852), .B(n9853), .Z(n9857) );
  NAND U11387 ( .A(n10361), .B(n10360), .Z(n9856) );
  AND U11388 ( .A(n9857), .B(n9856), .Z(n9858) );
  AND U11389 ( .A(a[16]), .B(b[36]), .Z(n9859) );
  NANDN U11390 ( .A(n9858), .B(n9859), .Z(n9863) );
  XOR U11391 ( .A(n9861), .B(n9860), .Z(n10366) );
  NAND U11392 ( .A(n10367), .B(n10366), .Z(n9862) );
  AND U11393 ( .A(n9863), .B(n9862), .Z(n9865) );
  NANDN U11394 ( .A(n9864), .B(n9865), .Z(n9867) );
  AND U11395 ( .A(a[17]), .B(b[36]), .Z(n10374) );
  NANDN U11396 ( .A(n10374), .B(n10375), .Z(n9866) );
  AND U11397 ( .A(n9867), .B(n9866), .Z(n9871) );
  NAND U11398 ( .A(n9871), .B(n9870), .Z(n9873) );
  NAND U11399 ( .A(a[18]), .B(b[36]), .Z(n10378) );
  XOR U11400 ( .A(n9871), .B(n9870), .Z(n10379) );
  NANDN U11401 ( .A(n10378), .B(n10379), .Z(n9872) );
  AND U11402 ( .A(n9873), .B(n9872), .Z(n9876) );
  AND U11403 ( .A(a[19]), .B(b[36]), .Z(n9877) );
  NANDN U11404 ( .A(n9876), .B(n9877), .Z(n9879) );
  XOR U11405 ( .A(n9875), .B(n9874), .Z(n10385) );
  NAND U11406 ( .A(n10385), .B(n10384), .Z(n9878) );
  AND U11407 ( .A(n9879), .B(n9878), .Z(n9882) );
  XOR U11408 ( .A(n9881), .B(n9880), .Z(n9883) );
  NANDN U11409 ( .A(n9882), .B(n9883), .Z(n9885) );
  AND U11410 ( .A(a[20]), .B(b[36]), .Z(n10391) );
  NAND U11411 ( .A(n10391), .B(n10390), .Z(n9884) );
  AND U11412 ( .A(n9885), .B(n9884), .Z(n9888) );
  XOR U11413 ( .A(n9887), .B(n9886), .Z(n9889) );
  NANDN U11414 ( .A(n9888), .B(n9889), .Z(n9891) );
  AND U11415 ( .A(a[21]), .B(b[36]), .Z(n10273) );
  NAND U11416 ( .A(n10273), .B(n10272), .Z(n9890) );
  AND U11417 ( .A(n9891), .B(n9890), .Z(n10400) );
  IV U11418 ( .A(n9895), .Z(n10401) );
  OR U11419 ( .A(n10400), .B(n10401), .Z(n9898) );
  ANDN U11420 ( .B(n10400), .A(n9895), .Z(n9896) );
  NAND U11421 ( .A(a[22]), .B(b[36]), .Z(n10403) );
  OR U11422 ( .A(n9896), .B(n10403), .Z(n9897) );
  AND U11423 ( .A(n9898), .B(n9897), .Z(n9902) );
  XOR U11424 ( .A(n9900), .B(n9899), .Z(n9901) );
  NANDN U11425 ( .A(n9902), .B(n9901), .Z(n9904) );
  NAND U11426 ( .A(a[23]), .B(b[36]), .Z(n10268) );
  XNOR U11427 ( .A(n9902), .B(n9901), .Z(n10269) );
  NANDN U11428 ( .A(n10268), .B(n10269), .Z(n9903) );
  AND U11429 ( .A(n9904), .B(n9903), .Z(n10410) );
  IV U11430 ( .A(n9908), .Z(n10411) );
  OR U11431 ( .A(n10410), .B(n10411), .Z(n9911) );
  ANDN U11432 ( .B(n10410), .A(n9908), .Z(n9909) );
  NAND U11433 ( .A(a[24]), .B(b[36]), .Z(n10413) );
  OR U11434 ( .A(n9909), .B(n10413), .Z(n9910) );
  AND U11435 ( .A(n9911), .B(n9910), .Z(n9915) );
  XOR U11436 ( .A(n9913), .B(n9912), .Z(n9914) );
  NANDN U11437 ( .A(n9915), .B(n9914), .Z(n9917) );
  XNOR U11438 ( .A(n9915), .B(n9914), .Z(n10267) );
  AND U11439 ( .A(a[25]), .B(b[36]), .Z(n10266) );
  NAND U11440 ( .A(n10267), .B(n10266), .Z(n9916) );
  NAND U11441 ( .A(n9917), .B(n9916), .Z(n10422) );
  NAND U11442 ( .A(a[26]), .B(b[36]), .Z(n10424) );
  XNOR U11443 ( .A(n9919), .B(n9918), .Z(n9921) );
  NAND U11444 ( .A(n9920), .B(n9921), .Z(n9923) );
  AND U11445 ( .A(a[27]), .B(b[36]), .Z(n10264) );
  XOR U11446 ( .A(n9921), .B(n9920), .Z(n10265) );
  NANDN U11447 ( .A(n10264), .B(n10265), .Z(n9922) );
  AND U11448 ( .A(n9923), .B(n9922), .Z(n9925) );
  NANDN U11449 ( .A(n9924), .B(n9925), .Z(n9929) );
  NAND U11450 ( .A(n10433), .B(n10434), .Z(n9928) );
  AND U11451 ( .A(n9929), .B(n9928), .Z(n9931) );
  AND U11452 ( .A(a[29]), .B(b[36]), .Z(n9930) );
  NANDN U11453 ( .A(n9931), .B(n9930), .Z(n9935) );
  XOR U11454 ( .A(n9931), .B(n9930), .Z(n10439) );
  XNOR U11455 ( .A(n9933), .B(n9932), .Z(n10440) );
  NANDN U11456 ( .A(n10439), .B(n10440), .Z(n9934) );
  AND U11457 ( .A(n9935), .B(n9934), .Z(n9937) );
  AND U11458 ( .A(a[30]), .B(b[36]), .Z(n9936) );
  NANDN U11459 ( .A(n9937), .B(n9936), .Z(n9941) );
  XOR U11460 ( .A(n9937), .B(n9936), .Z(n10445) );
  XNOR U11461 ( .A(n9939), .B(n9938), .Z(n10446) );
  NANDN U11462 ( .A(n10445), .B(n10446), .Z(n9940) );
  AND U11463 ( .A(n9941), .B(n9940), .Z(n9945) );
  XNOR U11464 ( .A(n9943), .B(n9942), .Z(n9944) );
  NANDN U11465 ( .A(n9945), .B(n9944), .Z(n9947) );
  NAND U11466 ( .A(a[31]), .B(b[36]), .Z(n10451) );
  XNOR U11467 ( .A(n9945), .B(n9944), .Z(n10452) );
  NANDN U11468 ( .A(n10451), .B(n10452), .Z(n9946) );
  AND U11469 ( .A(n9947), .B(n9946), .Z(n10460) );
  OR U11470 ( .A(n10459), .B(n10460), .Z(n9948) );
  AND U11471 ( .A(n9949), .B(n9948), .Z(n9953) );
  XNOR U11472 ( .A(n9951), .B(n9950), .Z(n9952) );
  NANDN U11473 ( .A(n9953), .B(n9952), .Z(n9955) );
  XNOR U11474 ( .A(n9953), .B(n9952), .Z(n10466) );
  AND U11475 ( .A(a[33]), .B(b[36]), .Z(n10465) );
  NAND U11476 ( .A(n10466), .B(n10465), .Z(n9954) );
  AND U11477 ( .A(n9955), .B(n9954), .Z(n9959) );
  AND U11478 ( .A(a[34]), .B(b[36]), .Z(n9958) );
  NANDN U11479 ( .A(n9959), .B(n9958), .Z(n9961) );
  XNOR U11480 ( .A(n9957), .B(n9956), .Z(n10472) );
  XNOR U11481 ( .A(n9959), .B(n9958), .Z(n10471) );
  NAND U11482 ( .A(n10472), .B(n10471), .Z(n9960) );
  AND U11483 ( .A(n9961), .B(n9960), .Z(n10476) );
  XNOR U11484 ( .A(n9963), .B(n9962), .Z(n10475) );
  NANDN U11485 ( .A(n10476), .B(n10475), .Z(n9964) );
  AND U11486 ( .A(n9965), .B(n9964), .Z(n9967) );
  AND U11487 ( .A(a[36]), .B(b[36]), .Z(n9966) );
  NANDN U11488 ( .A(n9967), .B(n9966), .Z(n9971) );
  XOR U11489 ( .A(n9967), .B(n9966), .Z(n10481) );
  XNOR U11490 ( .A(n9969), .B(n9968), .Z(n10482) );
  NANDN U11491 ( .A(n10481), .B(n10482), .Z(n9970) );
  AND U11492 ( .A(n9971), .B(n9970), .Z(n9975) );
  XNOR U11493 ( .A(n9973), .B(n9972), .Z(n9974) );
  NANDN U11494 ( .A(n9975), .B(n9974), .Z(n9977) );
  XNOR U11495 ( .A(n9975), .B(n9974), .Z(n10490) );
  AND U11496 ( .A(a[37]), .B(b[36]), .Z(n10489) );
  NAND U11497 ( .A(n10490), .B(n10489), .Z(n9976) );
  AND U11498 ( .A(n9977), .B(n9976), .Z(n10496) );
  OR U11499 ( .A(n10495), .B(n10496), .Z(n9978) );
  AND U11500 ( .A(n9979), .B(n9978), .Z(n9981) );
  AND U11501 ( .A(a[39]), .B(b[36]), .Z(n9980) );
  NANDN U11502 ( .A(n9981), .B(n9980), .Z(n9985) );
  XOR U11503 ( .A(n9981), .B(n9980), .Z(n10499) );
  XNOR U11504 ( .A(n9983), .B(n9982), .Z(n10500) );
  NANDN U11505 ( .A(n10499), .B(n10500), .Z(n9984) );
  AND U11506 ( .A(n9985), .B(n9984), .Z(n10508) );
  OR U11507 ( .A(n10507), .B(n10508), .Z(n9986) );
  AND U11508 ( .A(n9987), .B(n9986), .Z(n9991) );
  AND U11509 ( .A(a[41]), .B(b[36]), .Z(n9990) );
  NANDN U11510 ( .A(n9991), .B(n9990), .Z(n9993) );
  XOR U11511 ( .A(n9989), .B(n9988), .Z(n10512) );
  XNOR U11512 ( .A(n9991), .B(n9990), .Z(n10511) );
  NANDN U11513 ( .A(n10512), .B(n10511), .Z(n9992) );
  AND U11514 ( .A(n9993), .B(n9992), .Z(n9997) );
  XNOR U11515 ( .A(n9995), .B(n9994), .Z(n9996) );
  NANDN U11516 ( .A(n9997), .B(n9996), .Z(n9999) );
  XNOR U11517 ( .A(n9997), .B(n9996), .Z(n10520) );
  AND U11518 ( .A(a[42]), .B(b[36]), .Z(n10519) );
  NAND U11519 ( .A(n10520), .B(n10519), .Z(n9998) );
  AND U11520 ( .A(n9999), .B(n9998), .Z(n10003) );
  XNOR U11521 ( .A(n10001), .B(n10000), .Z(n10002) );
  NANDN U11522 ( .A(n10003), .B(n10002), .Z(n10005) );
  XNOR U11523 ( .A(n10003), .B(n10002), .Z(n10526) );
  AND U11524 ( .A(a[43]), .B(b[36]), .Z(n10525) );
  NAND U11525 ( .A(n10526), .B(n10525), .Z(n10004) );
  NAND U11526 ( .A(n10005), .B(n10004), .Z(n10006) );
  NANDN U11527 ( .A(n10007), .B(n10006), .Z(n10009) );
  XNOR U11528 ( .A(n10007), .B(n10006), .Z(n10532) );
  AND U11529 ( .A(a[44]), .B(b[36]), .Z(n10531) );
  NAND U11530 ( .A(n10532), .B(n10531), .Z(n10008) );
  AND U11531 ( .A(n10009), .B(n10008), .Z(n10538) );
  OR U11532 ( .A(n10537), .B(n10538), .Z(n10010) );
  AND U11533 ( .A(n10011), .B(n10010), .Z(n10013) );
  AND U11534 ( .A(a[46]), .B(b[36]), .Z(n10012) );
  NANDN U11535 ( .A(n10013), .B(n10012), .Z(n10017) );
  XOR U11536 ( .A(n10013), .B(n10012), .Z(n10541) );
  XNOR U11537 ( .A(n10015), .B(n10014), .Z(n10542) );
  NANDN U11538 ( .A(n10541), .B(n10542), .Z(n10016) );
  AND U11539 ( .A(n10017), .B(n10016), .Z(n10021) );
  XNOR U11540 ( .A(n10019), .B(n10018), .Z(n10020) );
  NANDN U11541 ( .A(n10021), .B(n10020), .Z(n10023) );
  NAND U11542 ( .A(a[47]), .B(b[36]), .Z(n10547) );
  XNOR U11543 ( .A(n10021), .B(n10020), .Z(n10548) );
  NANDN U11544 ( .A(n10547), .B(n10548), .Z(n10022) );
  AND U11545 ( .A(n10023), .B(n10022), .Z(n10027) );
  XNOR U11546 ( .A(n10025), .B(n10024), .Z(n10026) );
  NANDN U11547 ( .A(n10027), .B(n10026), .Z(n10029) );
  XNOR U11548 ( .A(n10027), .B(n10026), .Z(n10556) );
  AND U11549 ( .A(a[48]), .B(b[36]), .Z(n10555) );
  NAND U11550 ( .A(n10556), .B(n10555), .Z(n10028) );
  AND U11551 ( .A(n10029), .B(n10028), .Z(n10033) );
  XNOR U11552 ( .A(n10031), .B(n10030), .Z(n10032) );
  NANDN U11553 ( .A(n10033), .B(n10032), .Z(n10035) );
  XNOR U11554 ( .A(n10033), .B(n10032), .Z(n10562) );
  AND U11555 ( .A(a[49]), .B(b[36]), .Z(n10561) );
  NAND U11556 ( .A(n10562), .B(n10561), .Z(n10034) );
  AND U11557 ( .A(n10035), .B(n10034), .Z(n10568) );
  OR U11558 ( .A(n10567), .B(n10568), .Z(n10036) );
  AND U11559 ( .A(n10037), .B(n10036), .Z(n10041) );
  XNOR U11560 ( .A(n10039), .B(n10038), .Z(n10040) );
  NANDN U11561 ( .A(n10041), .B(n10040), .Z(n10043) );
  XNOR U11562 ( .A(n10041), .B(n10040), .Z(n10574) );
  AND U11563 ( .A(a[51]), .B(b[36]), .Z(n10573) );
  NAND U11564 ( .A(n10574), .B(n10573), .Z(n10042) );
  AND U11565 ( .A(n10043), .B(n10042), .Z(n10047) );
  XNOR U11566 ( .A(n10045), .B(n10044), .Z(n10046) );
  NANDN U11567 ( .A(n10047), .B(n10046), .Z(n10049) );
  NAND U11568 ( .A(a[52]), .B(b[36]), .Z(n10579) );
  XNOR U11569 ( .A(n10047), .B(n10046), .Z(n10580) );
  NANDN U11570 ( .A(n10579), .B(n10580), .Z(n10048) );
  AND U11571 ( .A(n10049), .B(n10048), .Z(n10584) );
  XNOR U11572 ( .A(n10051), .B(n10050), .Z(n10583) );
  NANDN U11573 ( .A(n10584), .B(n10583), .Z(n10052) );
  AND U11574 ( .A(n10053), .B(n10052), .Z(n10055) );
  AND U11575 ( .A(a[54]), .B(b[36]), .Z(n10054) );
  NANDN U11576 ( .A(n10055), .B(n10054), .Z(n10059) );
  XOR U11577 ( .A(n10055), .B(n10054), .Z(n10589) );
  XNOR U11578 ( .A(n10057), .B(n10056), .Z(n10590) );
  NANDN U11579 ( .A(n10589), .B(n10590), .Z(n10058) );
  AND U11580 ( .A(n10059), .B(n10058), .Z(n10598) );
  OR U11581 ( .A(n10597), .B(n10598), .Z(n10060) );
  AND U11582 ( .A(n10061), .B(n10060), .Z(n10065) );
  XNOR U11583 ( .A(n10063), .B(n10062), .Z(n10064) );
  NANDN U11584 ( .A(n10065), .B(n10064), .Z(n10067) );
  NAND U11585 ( .A(a[56]), .B(b[36]), .Z(n10601) );
  XNOR U11586 ( .A(n10065), .B(n10064), .Z(n10602) );
  NANDN U11587 ( .A(n10601), .B(n10602), .Z(n10066) );
  AND U11588 ( .A(n10067), .B(n10066), .Z(n10071) );
  AND U11589 ( .A(a[57]), .B(b[36]), .Z(n10070) );
  NANDN U11590 ( .A(n10071), .B(n10070), .Z(n10073) );
  XNOR U11591 ( .A(n10069), .B(n10068), .Z(n10610) );
  XNOR U11592 ( .A(n10071), .B(n10070), .Z(n10609) );
  NAND U11593 ( .A(n10610), .B(n10609), .Z(n10072) );
  AND U11594 ( .A(n10073), .B(n10072), .Z(n10614) );
  XNOR U11595 ( .A(n10075), .B(n10074), .Z(n10613) );
  NANDN U11596 ( .A(n10614), .B(n10613), .Z(n10076) );
  AND U11597 ( .A(n10077), .B(n10076), .Z(n10081) );
  XOR U11598 ( .A(n10079), .B(n10078), .Z(n10080) );
  NANDN U11599 ( .A(n10081), .B(n10080), .Z(n10083) );
  XNOR U11600 ( .A(n10081), .B(n10080), .Z(n10622) );
  AND U11601 ( .A(a[59]), .B(b[36]), .Z(n10621) );
  NAND U11602 ( .A(n10622), .B(n10621), .Z(n10082) );
  AND U11603 ( .A(n10083), .B(n10082), .Z(n10087) );
  AND U11604 ( .A(a[60]), .B(b[36]), .Z(n10086) );
  NANDN U11605 ( .A(n10087), .B(n10086), .Z(n10089) );
  XOR U11606 ( .A(n10085), .B(n10084), .Z(n10625) );
  XNOR U11607 ( .A(n10087), .B(n10086), .Z(n10626) );
  NANDN U11608 ( .A(n10625), .B(n10626), .Z(n10088) );
  AND U11609 ( .A(n10089), .B(n10088), .Z(n10091) );
  AND U11610 ( .A(a[61]), .B(b[36]), .Z(n10090) );
  NANDN U11611 ( .A(n10091), .B(n10090), .Z(n10095) );
  XOR U11612 ( .A(n10091), .B(n10090), .Z(n10631) );
  XNOR U11613 ( .A(n10093), .B(n10092), .Z(n10632) );
  NANDN U11614 ( .A(n10631), .B(n10632), .Z(n10094) );
  NAND U11615 ( .A(n10095), .B(n10094), .Z(n10096) );
  NAND U11616 ( .A(n10097), .B(n10096), .Z(n10099) );
  NAND U11617 ( .A(a[62]), .B(b[36]), .Z(n10637) );
  XOR U11618 ( .A(n10097), .B(n10096), .Z(n10638) );
  NANDN U11619 ( .A(n10637), .B(n10638), .Z(n10098) );
  AND U11620 ( .A(n10099), .B(n10098), .Z(n10102) );
  NANDN U11621 ( .A(n10102), .B(n10103), .Z(n10105) );
  NAND U11622 ( .A(a[63]), .B(b[36]), .Z(n10262) );
  NANDN U11623 ( .A(n10262), .B(n10263), .Z(n10104) );
  AND U11624 ( .A(n10105), .B(n10104), .Z(n10644) );
  ANDN U11625 ( .B(n10643), .A(n10644), .Z(n24793) );
  NAND U11626 ( .A(n10107), .B(n10106), .Z(n10111) );
  NAND U11627 ( .A(n10109), .B(n10108), .Z(n10110) );
  AND U11628 ( .A(n10111), .B(n10110), .Z(n22575) );
  AND U11629 ( .A(a[59]), .B(b[42]), .Z(n22574) );
  XOR U11630 ( .A(n22575), .B(n22574), .Z(n22576) );
  NANDN U11631 ( .A(n10113), .B(n10112), .Z(n10117) );
  NAND U11632 ( .A(n10115), .B(n10114), .Z(n10116) );
  AND U11633 ( .A(n10117), .B(n10116), .Z(n22598) );
  NAND U11634 ( .A(a[55]), .B(b[46]), .Z(n22599) );
  NANDN U11635 ( .A(n10119), .B(n10118), .Z(n10123) );
  NAND U11636 ( .A(n10121), .B(n10120), .Z(n10122) );
  AND U11637 ( .A(n10123), .B(n10122), .Z(n22622) );
  NAND U11638 ( .A(a[51]), .B(b[50]), .Z(n22623) );
  NANDN U11639 ( .A(n10125), .B(n10124), .Z(n10129) );
  NAND U11640 ( .A(n10127), .B(n10126), .Z(n10128) );
  AND U11641 ( .A(n10129), .B(n10128), .Z(n22640) );
  NAND U11642 ( .A(a[47]), .B(b[54]), .Z(n22641) );
  NANDN U11643 ( .A(n10131), .B(n10130), .Z(n10135) );
  NAND U11644 ( .A(n10133), .B(n10132), .Z(n10134) );
  AND U11645 ( .A(n10135), .B(n10134), .Z(n22683) );
  AND U11646 ( .A(b[63]), .B(a[38]), .Z(n22691) );
  NANDN U11647 ( .A(n10137), .B(n10136), .Z(n10141) );
  NANDN U11648 ( .A(n10139), .B(n10138), .Z(n10140) );
  AND U11649 ( .A(n10141), .B(n10140), .Z(n22688) );
  NAND U11650 ( .A(b[62]), .B(a[39]), .Z(n22689) );
  XOR U11651 ( .A(n22691), .B(n22690), .Z(n22682) );
  AND U11652 ( .A(a[40]), .B(b[61]), .Z(n22684) );
  XOR U11653 ( .A(n22685), .B(n22684), .Z(n22677) );
  NAND U11654 ( .A(a[41]), .B(b[60]), .Z(n22676) );
  NANDN U11655 ( .A(n10143), .B(n10142), .Z(n10147) );
  NAND U11656 ( .A(n10145), .B(n10144), .Z(n10146) );
  NAND U11657 ( .A(n10147), .B(n10146), .Z(n22679) );
  NANDN U11658 ( .A(n10149), .B(n10148), .Z(n10153) );
  NAND U11659 ( .A(n10151), .B(n10150), .Z(n10152) );
  AND U11660 ( .A(n10153), .B(n10152), .Z(n22670) );
  AND U11661 ( .A(a[42]), .B(b[59]), .Z(n22671) );
  XOR U11662 ( .A(n22673), .B(n22672), .Z(n22667) );
  NANDN U11663 ( .A(n10155), .B(n10154), .Z(n10159) );
  NANDN U11664 ( .A(n10157), .B(n10156), .Z(n10158) );
  AND U11665 ( .A(n10159), .B(n10158), .Z(n22664) );
  NAND U11666 ( .A(a[43]), .B(b[58]), .Z(n22665) );
  NANDN U11667 ( .A(n10161), .B(n10160), .Z(n10165) );
  NAND U11668 ( .A(n10163), .B(n10162), .Z(n10164) );
  AND U11669 ( .A(n10165), .B(n10164), .Z(n22659) );
  AND U11670 ( .A(a[44]), .B(b[57]), .Z(n22658) );
  XOR U11671 ( .A(n22661), .B(n22660), .Z(n22655) );
  NANDN U11672 ( .A(n10167), .B(n10166), .Z(n10171) );
  NAND U11673 ( .A(n10169), .B(n10168), .Z(n10170) );
  AND U11674 ( .A(n10171), .B(n10170), .Z(n22652) );
  NAND U11675 ( .A(a[45]), .B(b[56]), .Z(n22653) );
  XOR U11676 ( .A(n22655), .B(n22654), .Z(n22649) );
  NANDN U11677 ( .A(n10173), .B(n10172), .Z(n10177) );
  NAND U11678 ( .A(n10175), .B(n10174), .Z(n10176) );
  AND U11679 ( .A(n10177), .B(n10176), .Z(n22647) );
  AND U11680 ( .A(a[46]), .B(b[55]), .Z(n22646) );
  XOR U11681 ( .A(n22649), .B(n22648), .Z(n22642) );
  XOR U11682 ( .A(n22643), .B(n22642), .Z(n22697) );
  NANDN U11683 ( .A(n10179), .B(n10178), .Z(n10183) );
  NAND U11684 ( .A(n10181), .B(n10180), .Z(n10182) );
  AND U11685 ( .A(n10183), .B(n10182), .Z(n22695) );
  AND U11686 ( .A(a[48]), .B(b[53]), .Z(n22694) );
  XOR U11687 ( .A(n22697), .B(n22696), .Z(n22637) );
  NANDN U11688 ( .A(n10185), .B(n10184), .Z(n10189) );
  NAND U11689 ( .A(n10187), .B(n10186), .Z(n10188) );
  AND U11690 ( .A(n10189), .B(n10188), .Z(n22634) );
  NAND U11691 ( .A(a[49]), .B(b[52]), .Z(n22635) );
  XOR U11692 ( .A(n22637), .B(n22636), .Z(n22631) );
  NANDN U11693 ( .A(n10191), .B(n10190), .Z(n10195) );
  NAND U11694 ( .A(n10193), .B(n10192), .Z(n10194) );
  AND U11695 ( .A(n10195), .B(n10194), .Z(n22629) );
  AND U11696 ( .A(a[50]), .B(b[51]), .Z(n22628) );
  XOR U11697 ( .A(n22631), .B(n22630), .Z(n22624) );
  XOR U11698 ( .A(n22625), .B(n22624), .Z(n22619) );
  NANDN U11699 ( .A(n10197), .B(n10196), .Z(n10201) );
  NAND U11700 ( .A(n10199), .B(n10198), .Z(n10200) );
  AND U11701 ( .A(n10201), .B(n10200), .Z(n22617) );
  AND U11702 ( .A(a[52]), .B(b[49]), .Z(n22616) );
  XOR U11703 ( .A(n22619), .B(n22618), .Z(n22613) );
  NANDN U11704 ( .A(n10203), .B(n10202), .Z(n10207) );
  NAND U11705 ( .A(n10205), .B(n10204), .Z(n10206) );
  AND U11706 ( .A(n10207), .B(n10206), .Z(n22610) );
  NAND U11707 ( .A(a[53]), .B(b[48]), .Z(n22611) );
  XOR U11708 ( .A(n22613), .B(n22612), .Z(n22607) );
  NANDN U11709 ( .A(n10209), .B(n10208), .Z(n10213) );
  NAND U11710 ( .A(n10211), .B(n10210), .Z(n10212) );
  AND U11711 ( .A(n10213), .B(n10212), .Z(n22605) );
  AND U11712 ( .A(a[54]), .B(b[47]), .Z(n22604) );
  XOR U11713 ( .A(n22607), .B(n22606), .Z(n22600) );
  XOR U11714 ( .A(n22601), .B(n22600), .Z(n22595) );
  NANDN U11715 ( .A(n10215), .B(n10214), .Z(n10219) );
  NAND U11716 ( .A(n10217), .B(n10216), .Z(n10218) );
  AND U11717 ( .A(n10219), .B(n10218), .Z(n22593) );
  AND U11718 ( .A(a[56]), .B(b[45]), .Z(n22592) );
  XOR U11719 ( .A(n22595), .B(n22594), .Z(n22589) );
  NAND U11720 ( .A(n10221), .B(n10220), .Z(n10225) );
  NANDN U11721 ( .A(n10223), .B(n10222), .Z(n10224) );
  AND U11722 ( .A(n10225), .B(n10224), .Z(n22587) );
  AND U11723 ( .A(a[57]), .B(b[44]), .Z(n22586) );
  XOR U11724 ( .A(n22587), .B(n22586), .Z(n22588) );
  XOR U11725 ( .A(n22589), .B(n22588), .Z(n22583) );
  NAND U11726 ( .A(n10227), .B(n10226), .Z(n10231) );
  NANDN U11727 ( .A(n10229), .B(n10228), .Z(n10230) );
  NAND U11728 ( .A(n10231), .B(n10230), .Z(n22581) );
  NAND U11729 ( .A(a[58]), .B(b[43]), .Z(n22580) );
  XOR U11730 ( .A(n22581), .B(n22580), .Z(n22582) );
  NANDN U11731 ( .A(n10233), .B(n10232), .Z(n10237) );
  NANDN U11732 ( .A(n10235), .B(n10234), .Z(n10236) );
  AND U11733 ( .A(n10237), .B(n10236), .Z(n22569) );
  AND U11734 ( .A(a[60]), .B(b[41]), .Z(n22568) );
  XOR U11735 ( .A(n22571), .B(n22570), .Z(n22565) );
  AND U11736 ( .A(a[61]), .B(b[40]), .Z(n22562) );
  NANDN U11737 ( .A(n10239), .B(n10238), .Z(n10243) );
  NAND U11738 ( .A(n10241), .B(n10240), .Z(n10242) );
  NAND U11739 ( .A(n10243), .B(n10242), .Z(n22563) );
  XOR U11740 ( .A(n22565), .B(n22564), .Z(n22559) );
  NANDN U11741 ( .A(n10245), .B(n10244), .Z(n10249) );
  NAND U11742 ( .A(n10247), .B(n10246), .Z(n10248) );
  AND U11743 ( .A(n10249), .B(n10248), .Z(n22557) );
  AND U11744 ( .A(a[62]), .B(b[39]), .Z(n22556) );
  XOR U11745 ( .A(n22559), .B(n22558), .Z(n22703) );
  NAND U11746 ( .A(n10251), .B(n10250), .Z(n10255) );
  NANDN U11747 ( .A(n10253), .B(n10252), .Z(n10254) );
  NAND U11748 ( .A(n10255), .B(n10254), .Z(n22701) );
  NAND U11749 ( .A(a[63]), .B(b[38]), .Z(n22700) );
  XOR U11750 ( .A(n22701), .B(n22700), .Z(n22702) );
  NANDN U11751 ( .A(n10257), .B(n10256), .Z(n10261) );
  NAND U11752 ( .A(n10259), .B(n10258), .Z(n10260) );
  NAND U11753 ( .A(n10261), .B(n10260), .Z(n22555) );
  XNOR U11754 ( .A(n22554), .B(n22555), .Z(n24794) );
  NAND U11755 ( .A(a[61]), .B(b[35]), .Z(n10627) );
  AND U11756 ( .A(a[60]), .B(b[35]), .Z(n10620) );
  NAND U11757 ( .A(a[59]), .B(b[35]), .Z(n10615) );
  AND U11758 ( .A(a[58]), .B(b[35]), .Z(n10608) );
  NAND U11759 ( .A(a[57]), .B(b[35]), .Z(n10603) );
  AND U11760 ( .A(a[56]), .B(b[35]), .Z(n10596) );
  NAND U11761 ( .A(a[53]), .B(b[35]), .Z(n10577) );
  AND U11762 ( .A(a[52]), .B(b[35]), .Z(n10572) );
  AND U11763 ( .A(a[51]), .B(b[35]), .Z(n10566) );
  AND U11764 ( .A(a[50]), .B(b[35]), .Z(n10560) );
  AND U11765 ( .A(a[49]), .B(b[35]), .Z(n10554) );
  NAND U11766 ( .A(a[47]), .B(b[35]), .Z(n10543) );
  AND U11767 ( .A(a[46]), .B(b[35]), .Z(n10536) );
  AND U11768 ( .A(a[45]), .B(b[35]), .Z(n10530) );
  AND U11769 ( .A(a[44]), .B(b[35]), .Z(n10524) );
  AND U11770 ( .A(a[43]), .B(b[35]), .Z(n10518) );
  NAND U11771 ( .A(a[42]), .B(b[35]), .Z(n10513) );
  AND U11772 ( .A(a[41]), .B(b[35]), .Z(n10506) );
  NAND U11773 ( .A(a[40]), .B(b[35]), .Z(n10501) );
  AND U11774 ( .A(a[39]), .B(b[35]), .Z(n10494) );
  AND U11775 ( .A(a[38]), .B(b[35]), .Z(n10488) );
  NAND U11776 ( .A(a[36]), .B(b[35]), .Z(n10477) );
  AND U11777 ( .A(a[35]), .B(b[35]), .Z(n10470) );
  AND U11778 ( .A(a[34]), .B(b[35]), .Z(n10464) );
  AND U11779 ( .A(a[33]), .B(b[35]), .Z(n10458) );
  AND U11780 ( .A(a[28]), .B(b[35]), .Z(n10429) );
  NAND U11781 ( .A(n10429), .B(n10430), .Z(n10432) );
  NAND U11782 ( .A(a[27]), .B(b[35]), .Z(n10425) );
  AND U11783 ( .A(a[26]), .B(b[35]), .Z(n10418) );
  XNOR U11784 ( .A(n10267), .B(n10266), .Z(n10419) );
  NANDN U11785 ( .A(n10418), .B(n10419), .Z(n10421) );
  AND U11786 ( .A(a[24]), .B(b[35]), .Z(n10271) );
  NAND U11787 ( .A(n10271), .B(n10270), .Z(n10409) );
  XOR U11788 ( .A(n10271), .B(n10270), .Z(n10708) );
  AND U11789 ( .A(a[22]), .B(b[35]), .Z(n10397) );
  XOR U11790 ( .A(n10273), .B(n10272), .Z(n10396) );
  NAND U11791 ( .A(n10397), .B(n10396), .Z(n10399) );
  AND U11792 ( .A(a[0]), .B(b[35]), .Z(n10999) );
  AND U11793 ( .A(a[1]), .B(b[36]), .Z(n10275) );
  AND U11794 ( .A(n10999), .B(n10275), .Z(n10274) );
  NAND U11795 ( .A(a[2]), .B(n10274), .Z(n10281) );
  NAND U11796 ( .A(n10275), .B(a[0]), .Z(n10276) );
  XNOR U11797 ( .A(a[2]), .B(n10276), .Z(n10277) );
  NAND U11798 ( .A(b[35]), .B(n10277), .Z(n10731) );
  NAND U11799 ( .A(b[36]), .B(a[1]), .Z(n10278) );
  XNOR U11800 ( .A(n10279), .B(n10278), .Z(n10732) );
  NANDN U11801 ( .A(n10731), .B(n10732), .Z(n10280) );
  AND U11802 ( .A(n10281), .B(n10280), .Z(n10282) );
  AND U11803 ( .A(a[3]), .B(b[35]), .Z(n10283) );
  NANDN U11804 ( .A(n10282), .B(n10283), .Z(n10287) );
  NAND U11805 ( .A(n10738), .B(n10737), .Z(n10286) );
  AND U11806 ( .A(n10287), .B(n10286), .Z(n10290) );
  NANDN U11807 ( .A(n10290), .B(n10291), .Z(n10293) );
  AND U11808 ( .A(a[4]), .B(b[35]), .Z(n10722) );
  NAND U11809 ( .A(n10722), .B(n10721), .Z(n10292) );
  AND U11810 ( .A(n10293), .B(n10292), .Z(n10296) );
  XOR U11811 ( .A(n10295), .B(n10294), .Z(n10297) );
  NANDN U11812 ( .A(n10296), .B(n10297), .Z(n10299) );
  NAND U11813 ( .A(a[5]), .B(b[35]), .Z(n10747) );
  NANDN U11814 ( .A(n10747), .B(n10748), .Z(n10298) );
  AND U11815 ( .A(n10299), .B(n10298), .Z(n10302) );
  NANDN U11816 ( .A(n10302), .B(n10303), .Z(n10305) );
  NAND U11817 ( .A(a[6]), .B(b[35]), .Z(n10753) );
  NANDN U11818 ( .A(n10753), .B(n10754), .Z(n10304) );
  AND U11819 ( .A(n10305), .B(n10304), .Z(n10308) );
  XOR U11820 ( .A(n10307), .B(n10306), .Z(n10309) );
  NANDN U11821 ( .A(n10308), .B(n10309), .Z(n10311) );
  NAND U11822 ( .A(a[7]), .B(b[35]), .Z(n10756) );
  NANDN U11823 ( .A(n10756), .B(n10757), .Z(n10310) );
  AND U11824 ( .A(n10311), .B(n10310), .Z(n10314) );
  AND U11825 ( .A(a[8]), .B(b[35]), .Z(n10315) );
  NANDN U11826 ( .A(n10314), .B(n10315), .Z(n10317) );
  XOR U11827 ( .A(n10313), .B(n10312), .Z(n10720) );
  NAND U11828 ( .A(n10720), .B(n10719), .Z(n10316) );
  AND U11829 ( .A(n10317), .B(n10316), .Z(n10320) );
  NANDN U11830 ( .A(n10320), .B(n10321), .Z(n10323) );
  NAND U11831 ( .A(a[9]), .B(b[35]), .Z(n10764) );
  NANDN U11832 ( .A(n10764), .B(n10765), .Z(n10322) );
  AND U11833 ( .A(n10323), .B(n10322), .Z(n10326) );
  NANDN U11834 ( .A(n10326), .B(n10327), .Z(n10329) );
  AND U11835 ( .A(a[10]), .B(b[35]), .Z(n10717) );
  NAND U11836 ( .A(n10718), .B(n10717), .Z(n10328) );
  AND U11837 ( .A(n10329), .B(n10328), .Z(n10330) );
  AND U11838 ( .A(a[11]), .B(b[35]), .Z(n10331) );
  NANDN U11839 ( .A(n10330), .B(n10331), .Z(n10335) );
  NAND U11840 ( .A(n10771), .B(n10770), .Z(n10334) );
  AND U11841 ( .A(n10335), .B(n10334), .Z(n10338) );
  AND U11842 ( .A(a[12]), .B(b[35]), .Z(n10339) );
  NANDN U11843 ( .A(n10338), .B(n10339), .Z(n10341) );
  XOR U11844 ( .A(n10337), .B(n10336), .Z(n10774) );
  NANDN U11845 ( .A(n10774), .B(n10775), .Z(n10340) );
  AND U11846 ( .A(n10341), .B(n10340), .Z(n10344) );
  AND U11847 ( .A(a[13]), .B(b[35]), .Z(n10345) );
  NANDN U11848 ( .A(n10344), .B(n10345), .Z(n10347) );
  XOR U11849 ( .A(n10343), .B(n10342), .Z(n10777) );
  NAND U11850 ( .A(n10777), .B(n10776), .Z(n10346) );
  AND U11851 ( .A(n10347), .B(n10346), .Z(n10350) );
  AND U11852 ( .A(a[14]), .B(b[35]), .Z(n10351) );
  NANDN U11853 ( .A(n10350), .B(n10351), .Z(n10353) );
  XOR U11854 ( .A(n10349), .B(n10348), .Z(n10716) );
  NAND U11855 ( .A(n10716), .B(n10715), .Z(n10352) );
  AND U11856 ( .A(n10353), .B(n10352), .Z(n10356) );
  XOR U11857 ( .A(n10355), .B(n10354), .Z(n10357) );
  NANDN U11858 ( .A(n10356), .B(n10357), .Z(n10359) );
  NAND U11859 ( .A(a[15]), .B(b[35]), .Z(n10784) );
  NANDN U11860 ( .A(n10784), .B(n10785), .Z(n10358) );
  AND U11861 ( .A(n10359), .B(n10358), .Z(n10362) );
  XOR U11862 ( .A(n10361), .B(n10360), .Z(n10363) );
  NANDN U11863 ( .A(n10362), .B(n10363), .Z(n10365) );
  NAND U11864 ( .A(a[16]), .B(b[35]), .Z(n10788) );
  NANDN U11865 ( .A(n10788), .B(n10789), .Z(n10364) );
  AND U11866 ( .A(n10365), .B(n10364), .Z(n10368) );
  XOR U11867 ( .A(n10367), .B(n10366), .Z(n10369) );
  NANDN U11868 ( .A(n10368), .B(n10369), .Z(n10371) );
  AND U11869 ( .A(a[17]), .B(b[35]), .Z(n10795) );
  NAND U11870 ( .A(n10795), .B(n10794), .Z(n10370) );
  AND U11871 ( .A(n10371), .B(n10370), .Z(n10372) );
  AND U11872 ( .A(a[18]), .B(b[35]), .Z(n10373) );
  NANDN U11873 ( .A(n10372), .B(n10373), .Z(n10377) );
  NAND U11874 ( .A(n10713), .B(n10714), .Z(n10376) );
  AND U11875 ( .A(n10377), .B(n10376), .Z(n10380) );
  NANDN U11876 ( .A(n10380), .B(n10381), .Z(n10383) );
  AND U11877 ( .A(a[19]), .B(b[35]), .Z(n10801) );
  NAND U11878 ( .A(n10801), .B(n10800), .Z(n10382) );
  AND U11879 ( .A(n10383), .B(n10382), .Z(n10386) );
  AND U11880 ( .A(a[20]), .B(b[35]), .Z(n10387) );
  NANDN U11881 ( .A(n10386), .B(n10387), .Z(n10389) );
  XOR U11882 ( .A(n10385), .B(n10384), .Z(n10712) );
  NAND U11883 ( .A(n10712), .B(n10711), .Z(n10388) );
  AND U11884 ( .A(n10389), .B(n10388), .Z(n10392) );
  AND U11885 ( .A(a[21]), .B(b[35]), .Z(n10393) );
  NANDN U11886 ( .A(n10392), .B(n10393), .Z(n10395) );
  XOR U11887 ( .A(n10391), .B(n10390), .Z(n10809) );
  NAND U11888 ( .A(n10809), .B(n10808), .Z(n10394) );
  AND U11889 ( .A(n10395), .B(n10394), .Z(n10709) );
  XOR U11890 ( .A(n10397), .B(n10396), .Z(n10710) );
  NANDN U11891 ( .A(n10709), .B(n10710), .Z(n10398) );
  AND U11892 ( .A(n10399), .B(n10398), .Z(n10404) );
  AND U11893 ( .A(a[23]), .B(b[35]), .Z(n10405) );
  NANDN U11894 ( .A(n10404), .B(n10405), .Z(n10407) );
  XOR U11895 ( .A(n10401), .B(n10400), .Z(n10402) );
  XNOR U11896 ( .A(n10403), .B(n10402), .Z(n10815) );
  NAND U11897 ( .A(n10815), .B(n10814), .Z(n10406) );
  NAND U11898 ( .A(n10407), .B(n10406), .Z(n10707) );
  NAND U11899 ( .A(n10708), .B(n10707), .Z(n10408) );
  AND U11900 ( .A(n10409), .B(n10408), .Z(n10414) );
  AND U11901 ( .A(a[25]), .B(b[35]), .Z(n10415) );
  NANDN U11902 ( .A(n10414), .B(n10415), .Z(n10417) );
  XOR U11903 ( .A(n10411), .B(n10410), .Z(n10412) );
  XNOR U11904 ( .A(n10413), .B(n10412), .Z(n10821) );
  NAND U11905 ( .A(n10821), .B(n10820), .Z(n10416) );
  AND U11906 ( .A(n10417), .B(n10416), .Z(n10706) );
  NAND U11907 ( .A(n10706), .B(n10705), .Z(n10420) );
  AND U11908 ( .A(n10421), .B(n10420), .Z(n10426) );
  NANDN U11909 ( .A(n10425), .B(n10426), .Z(n10428) );
  NAND U11910 ( .A(n10827), .B(n10826), .Z(n10427) );
  AND U11911 ( .A(n10428), .B(n10427), .Z(n10830) );
  XOR U11912 ( .A(n10430), .B(n10429), .Z(n10831) );
  NANDN U11913 ( .A(n10830), .B(n10831), .Z(n10431) );
  AND U11914 ( .A(n10432), .B(n10431), .Z(n10435) );
  XOR U11915 ( .A(n10434), .B(n10433), .Z(n10436) );
  NANDN U11916 ( .A(n10435), .B(n10436), .Z(n10438) );
  AND U11917 ( .A(a[29]), .B(b[35]), .Z(n10837) );
  NAND U11918 ( .A(n10837), .B(n10836), .Z(n10437) );
  AND U11919 ( .A(n10438), .B(n10437), .Z(n10442) );
  XNOR U11920 ( .A(n10440), .B(n10439), .Z(n10441) );
  NANDN U11921 ( .A(n10442), .B(n10441), .Z(n10444) );
  NAND U11922 ( .A(a[30]), .B(b[35]), .Z(n10842) );
  XNOR U11923 ( .A(n10442), .B(n10441), .Z(n10843) );
  NANDN U11924 ( .A(n10842), .B(n10843), .Z(n10443) );
  AND U11925 ( .A(n10444), .B(n10443), .Z(n10448) );
  AND U11926 ( .A(a[31]), .B(b[35]), .Z(n10447) );
  NANDN U11927 ( .A(n10448), .B(n10447), .Z(n10450) );
  XOR U11928 ( .A(n10446), .B(n10445), .Z(n10703) );
  XNOR U11929 ( .A(n10448), .B(n10447), .Z(n10704) );
  NANDN U11930 ( .A(n10703), .B(n10704), .Z(n10449) );
  AND U11931 ( .A(n10450), .B(n10449), .Z(n10454) );
  AND U11932 ( .A(a[32]), .B(b[35]), .Z(n10453) );
  NANDN U11933 ( .A(n10454), .B(n10453), .Z(n10456) );
  XOR U11934 ( .A(n10452), .B(n10451), .Z(n10701) );
  XNOR U11935 ( .A(n10454), .B(n10453), .Z(n10702) );
  NANDN U11936 ( .A(n10701), .B(n10702), .Z(n10455) );
  AND U11937 ( .A(n10456), .B(n10455), .Z(n10457) );
  NANDN U11938 ( .A(n10458), .B(n10457), .Z(n10462) );
  XOR U11939 ( .A(n10458), .B(n10457), .Z(n10858) );
  XOR U11940 ( .A(n10460), .B(n10459), .Z(n10859) );
  OR U11941 ( .A(n10858), .B(n10859), .Z(n10461) );
  NAND U11942 ( .A(n10462), .B(n10461), .Z(n10463) );
  NANDN U11943 ( .A(n10464), .B(n10463), .Z(n10468) );
  XOR U11944 ( .A(n10464), .B(n10463), .Z(n10699) );
  XOR U11945 ( .A(n10466), .B(n10465), .Z(n10700) );
  OR U11946 ( .A(n10699), .B(n10700), .Z(n10467) );
  NAND U11947 ( .A(n10468), .B(n10467), .Z(n10469) );
  NANDN U11948 ( .A(n10470), .B(n10469), .Z(n10474) );
  XOR U11949 ( .A(n10470), .B(n10469), .Z(n10695) );
  XOR U11950 ( .A(n10472), .B(n10471), .Z(n10696) );
  OR U11951 ( .A(n10695), .B(n10696), .Z(n10473) );
  AND U11952 ( .A(n10474), .B(n10473), .Z(n10478) );
  NANDN U11953 ( .A(n10477), .B(n10478), .Z(n10480) );
  XOR U11954 ( .A(n10476), .B(n10475), .Z(n10864) );
  XNOR U11955 ( .A(n10478), .B(n10477), .Z(n10865) );
  NANDN U11956 ( .A(n10864), .B(n10865), .Z(n10479) );
  AND U11957 ( .A(n10480), .B(n10479), .Z(n10484) );
  AND U11958 ( .A(a[37]), .B(b[35]), .Z(n10483) );
  NANDN U11959 ( .A(n10484), .B(n10483), .Z(n10486) );
  XOR U11960 ( .A(n10482), .B(n10481), .Z(n10693) );
  XNOR U11961 ( .A(n10484), .B(n10483), .Z(n10694) );
  NANDN U11962 ( .A(n10693), .B(n10694), .Z(n10485) );
  AND U11963 ( .A(n10486), .B(n10485), .Z(n10487) );
  NANDN U11964 ( .A(n10488), .B(n10487), .Z(n10492) );
  XOR U11965 ( .A(n10488), .B(n10487), .Z(n10689) );
  XOR U11966 ( .A(n10490), .B(n10489), .Z(n10690) );
  OR U11967 ( .A(n10689), .B(n10690), .Z(n10491) );
  NAND U11968 ( .A(n10492), .B(n10491), .Z(n10493) );
  NANDN U11969 ( .A(n10494), .B(n10493), .Z(n10498) );
  XOR U11970 ( .A(n10494), .B(n10493), .Z(n10878) );
  XOR U11971 ( .A(n10496), .B(n10495), .Z(n10879) );
  OR U11972 ( .A(n10878), .B(n10879), .Z(n10497) );
  AND U11973 ( .A(n10498), .B(n10497), .Z(n10502) );
  NANDN U11974 ( .A(n10501), .B(n10502), .Z(n10504) );
  XOR U11975 ( .A(n10500), .B(n10499), .Z(n10882) );
  XNOR U11976 ( .A(n10502), .B(n10501), .Z(n10883) );
  NANDN U11977 ( .A(n10882), .B(n10883), .Z(n10503) );
  AND U11978 ( .A(n10504), .B(n10503), .Z(n10505) );
  NANDN U11979 ( .A(n10506), .B(n10505), .Z(n10510) );
  XOR U11980 ( .A(n10506), .B(n10505), .Z(n10685) );
  XOR U11981 ( .A(n10508), .B(n10507), .Z(n10686) );
  OR U11982 ( .A(n10685), .B(n10686), .Z(n10509) );
  AND U11983 ( .A(n10510), .B(n10509), .Z(n10514) );
  NANDN U11984 ( .A(n10513), .B(n10514), .Z(n10516) );
  XOR U11985 ( .A(n10512), .B(n10511), .Z(n10892) );
  XNOR U11986 ( .A(n10514), .B(n10513), .Z(n10893) );
  NANDN U11987 ( .A(n10892), .B(n10893), .Z(n10515) );
  AND U11988 ( .A(n10516), .B(n10515), .Z(n10517) );
  NANDN U11989 ( .A(n10518), .B(n10517), .Z(n10522) );
  XOR U11990 ( .A(n10518), .B(n10517), .Z(n10681) );
  XOR U11991 ( .A(n10520), .B(n10519), .Z(n10682) );
  OR U11992 ( .A(n10681), .B(n10682), .Z(n10521) );
  NAND U11993 ( .A(n10522), .B(n10521), .Z(n10523) );
  NANDN U11994 ( .A(n10524), .B(n10523), .Z(n10528) );
  XOR U11995 ( .A(n10524), .B(n10523), .Z(n10898) );
  XOR U11996 ( .A(n10526), .B(n10525), .Z(n10899) );
  OR U11997 ( .A(n10898), .B(n10899), .Z(n10527) );
  NAND U11998 ( .A(n10528), .B(n10527), .Z(n10529) );
  NANDN U11999 ( .A(n10530), .B(n10529), .Z(n10534) );
  XOR U12000 ( .A(n10530), .B(n10529), .Z(n10677) );
  XOR U12001 ( .A(n10532), .B(n10531), .Z(n10678) );
  OR U12002 ( .A(n10677), .B(n10678), .Z(n10533) );
  NAND U12003 ( .A(n10534), .B(n10533), .Z(n10535) );
  NANDN U12004 ( .A(n10536), .B(n10535), .Z(n10540) );
  XOR U12005 ( .A(n10536), .B(n10535), .Z(n10906) );
  XOR U12006 ( .A(n10538), .B(n10537), .Z(n10907) );
  OR U12007 ( .A(n10906), .B(n10907), .Z(n10539) );
  AND U12008 ( .A(n10540), .B(n10539), .Z(n10544) );
  NANDN U12009 ( .A(n10543), .B(n10544), .Z(n10546) );
  XOR U12010 ( .A(n10542), .B(n10541), .Z(n10673) );
  XNOR U12011 ( .A(n10544), .B(n10543), .Z(n10674) );
  NANDN U12012 ( .A(n10673), .B(n10674), .Z(n10545) );
  AND U12013 ( .A(n10546), .B(n10545), .Z(n10550) );
  AND U12014 ( .A(a[48]), .B(b[35]), .Z(n10549) );
  NANDN U12015 ( .A(n10550), .B(n10549), .Z(n10552) );
  XOR U12016 ( .A(n10548), .B(n10547), .Z(n10916) );
  XNOR U12017 ( .A(n10550), .B(n10549), .Z(n10917) );
  NANDN U12018 ( .A(n10916), .B(n10917), .Z(n10551) );
  AND U12019 ( .A(n10552), .B(n10551), .Z(n10553) );
  NANDN U12020 ( .A(n10554), .B(n10553), .Z(n10558) );
  XOR U12021 ( .A(n10554), .B(n10553), .Z(n10669) );
  XOR U12022 ( .A(n10556), .B(n10555), .Z(n10670) );
  OR U12023 ( .A(n10669), .B(n10670), .Z(n10557) );
  NAND U12024 ( .A(n10558), .B(n10557), .Z(n10559) );
  NANDN U12025 ( .A(n10560), .B(n10559), .Z(n10564) );
  XOR U12026 ( .A(n10560), .B(n10559), .Z(n10665) );
  XOR U12027 ( .A(n10562), .B(n10561), .Z(n10666) );
  OR U12028 ( .A(n10665), .B(n10666), .Z(n10563) );
  NAND U12029 ( .A(n10564), .B(n10563), .Z(n10565) );
  NANDN U12030 ( .A(n10566), .B(n10565), .Z(n10570) );
  XOR U12031 ( .A(n10566), .B(n10565), .Z(n10926) );
  XOR U12032 ( .A(n10568), .B(n10567), .Z(n10927) );
  OR U12033 ( .A(n10926), .B(n10927), .Z(n10569) );
  NAND U12034 ( .A(n10570), .B(n10569), .Z(n10571) );
  NANDN U12035 ( .A(n10572), .B(n10571), .Z(n10576) );
  XOR U12036 ( .A(n10572), .B(n10571), .Z(n10661) );
  XOR U12037 ( .A(n10574), .B(n10573), .Z(n10662) );
  OR U12038 ( .A(n10661), .B(n10662), .Z(n10575) );
  AND U12039 ( .A(n10576), .B(n10575), .Z(n10578) );
  NANDN U12040 ( .A(n10577), .B(n10578), .Z(n10582) );
  XNOR U12041 ( .A(n10578), .B(n10577), .Z(n10660) );
  XNOR U12042 ( .A(n10580), .B(n10579), .Z(n10659) );
  NAND U12043 ( .A(n10660), .B(n10659), .Z(n10581) );
  AND U12044 ( .A(n10582), .B(n10581), .Z(n10586) );
  AND U12045 ( .A(a[54]), .B(b[35]), .Z(n10585) );
  NANDN U12046 ( .A(n10586), .B(n10585), .Z(n10588) );
  XOR U12047 ( .A(n10584), .B(n10583), .Z(n10657) );
  XNOR U12048 ( .A(n10586), .B(n10585), .Z(n10658) );
  NANDN U12049 ( .A(n10657), .B(n10658), .Z(n10587) );
  AND U12050 ( .A(n10588), .B(n10587), .Z(n10592) );
  AND U12051 ( .A(a[55]), .B(b[35]), .Z(n10591) );
  NANDN U12052 ( .A(n10592), .B(n10591), .Z(n10594) );
  XOR U12053 ( .A(n10590), .B(n10589), .Z(n10942) );
  XNOR U12054 ( .A(n10592), .B(n10591), .Z(n10943) );
  NANDN U12055 ( .A(n10942), .B(n10943), .Z(n10593) );
  AND U12056 ( .A(n10594), .B(n10593), .Z(n10595) );
  NANDN U12057 ( .A(n10596), .B(n10595), .Z(n10600) );
  XOR U12058 ( .A(n10596), .B(n10595), .Z(n10653) );
  XOR U12059 ( .A(n10598), .B(n10597), .Z(n10654) );
  OR U12060 ( .A(n10653), .B(n10654), .Z(n10599) );
  AND U12061 ( .A(n10600), .B(n10599), .Z(n10604) );
  NANDN U12062 ( .A(n10603), .B(n10604), .Z(n10606) );
  XOR U12063 ( .A(n10602), .B(n10601), .Z(n10948) );
  XNOR U12064 ( .A(n10604), .B(n10603), .Z(n10949) );
  NANDN U12065 ( .A(n10948), .B(n10949), .Z(n10605) );
  AND U12066 ( .A(n10606), .B(n10605), .Z(n10607) );
  NANDN U12067 ( .A(n10608), .B(n10607), .Z(n10612) );
  XOR U12068 ( .A(n10608), .B(n10607), .Z(n10651) );
  XOR U12069 ( .A(n10610), .B(n10609), .Z(n10652) );
  OR U12070 ( .A(n10651), .B(n10652), .Z(n10611) );
  AND U12071 ( .A(n10612), .B(n10611), .Z(n10616) );
  NANDN U12072 ( .A(n10615), .B(n10616), .Z(n10618) );
  XOR U12073 ( .A(n10614), .B(n10613), .Z(n10960) );
  XNOR U12074 ( .A(n10616), .B(n10615), .Z(n10961) );
  NANDN U12075 ( .A(n10960), .B(n10961), .Z(n10617) );
  AND U12076 ( .A(n10618), .B(n10617), .Z(n10619) );
  NANDN U12077 ( .A(n10620), .B(n10619), .Z(n10624) );
  XOR U12078 ( .A(n10620), .B(n10619), .Z(n10647) );
  XOR U12079 ( .A(n10622), .B(n10621), .Z(n10648) );
  OR U12080 ( .A(n10647), .B(n10648), .Z(n10623) );
  AND U12081 ( .A(n10624), .B(n10623), .Z(n10628) );
  NANDN U12082 ( .A(n10627), .B(n10628), .Z(n10630) );
  XOR U12083 ( .A(n10626), .B(n10625), .Z(n10966) );
  XNOR U12084 ( .A(n10628), .B(n10627), .Z(n10967) );
  NANDN U12085 ( .A(n10966), .B(n10967), .Z(n10629) );
  AND U12086 ( .A(n10630), .B(n10629), .Z(n10634) );
  AND U12087 ( .A(a[62]), .B(b[35]), .Z(n10633) );
  NANDN U12088 ( .A(n10634), .B(n10633), .Z(n10636) );
  XNOR U12089 ( .A(n10632), .B(n10631), .Z(n10975) );
  XNOR U12090 ( .A(n10634), .B(n10633), .Z(n10974) );
  NAND U12091 ( .A(n10975), .B(n10974), .Z(n10635) );
  AND U12092 ( .A(n10636), .B(n10635), .Z(n10640) );
  AND U12093 ( .A(a[63]), .B(b[35]), .Z(n10639) );
  NANDN U12094 ( .A(n10640), .B(n10639), .Z(n10642) );
  XOR U12095 ( .A(n10638), .B(n10637), .Z(n10645) );
  XNOR U12096 ( .A(n10640), .B(n10639), .Z(n10646) );
  NANDN U12097 ( .A(n10645), .B(n10646), .Z(n10641) );
  AND U12098 ( .A(n10642), .B(n10641), .Z(n10979) );
  ANDN U12099 ( .B(n10978), .A(n10979), .Z(n22551) );
  XOR U12100 ( .A(n10644), .B(n10643), .Z(n22550) );
  NANDN U12101 ( .A(n22551), .B(n22550), .Z(n22553) );
  XNOR U12102 ( .A(n10646), .B(n10645), .Z(n11348) );
  AND U12103 ( .A(a[63]), .B(b[34]), .Z(n10973) );
  XOR U12104 ( .A(n10648), .B(n10647), .Z(n10650) );
  AND U12105 ( .A(a[61]), .B(b[34]), .Z(n10649) );
  NANDN U12106 ( .A(n10650), .B(n10649), .Z(n10965) );
  XOR U12107 ( .A(n10650), .B(n10649), .Z(n11335) );
  XOR U12108 ( .A(n10652), .B(n10651), .Z(n10955) );
  AND U12109 ( .A(a[59]), .B(b[34]), .Z(n10954) );
  NANDN U12110 ( .A(n10955), .B(n10954), .Z(n10957) );
  XOR U12111 ( .A(n10654), .B(n10653), .Z(n10656) );
  AND U12112 ( .A(a[57]), .B(b[34]), .Z(n10655) );
  NANDN U12113 ( .A(n10656), .B(n10655), .Z(n10947) );
  XOR U12114 ( .A(n10656), .B(n10655), .Z(n11311) );
  NAND U12115 ( .A(a[55]), .B(b[34]), .Z(n10936) );
  XNOR U12116 ( .A(n10658), .B(n10657), .Z(n10937) );
  NANDN U12117 ( .A(n10936), .B(n10937), .Z(n10939) );
  XOR U12118 ( .A(n10660), .B(n10659), .Z(n10933) );
  XOR U12119 ( .A(n10662), .B(n10661), .Z(n10664) );
  AND U12120 ( .A(a[53]), .B(b[34]), .Z(n10663) );
  NANDN U12121 ( .A(n10664), .B(n10663), .Z(n10931) );
  XOR U12122 ( .A(n10664), .B(n10663), .Z(n11287) );
  XOR U12123 ( .A(n10666), .B(n10665), .Z(n10668) );
  AND U12124 ( .A(a[51]), .B(b[34]), .Z(n10667) );
  NANDN U12125 ( .A(n10668), .B(n10667), .Z(n10923) );
  XOR U12126 ( .A(n10668), .B(n10667), .Z(n11275) );
  XOR U12127 ( .A(n10670), .B(n10669), .Z(n10672) );
  AND U12128 ( .A(a[50]), .B(b[34]), .Z(n10671) );
  NANDN U12129 ( .A(n10672), .B(n10671), .Z(n10921) );
  XOR U12130 ( .A(n10672), .B(n10671), .Z(n11269) );
  NAND U12131 ( .A(a[48]), .B(b[34]), .Z(n10675) );
  XNOR U12132 ( .A(n10674), .B(n10673), .Z(n10676) );
  NANDN U12133 ( .A(n10675), .B(n10676), .Z(n10913) );
  XOR U12134 ( .A(n10676), .B(n10675), .Z(n11257) );
  XOR U12135 ( .A(n10678), .B(n10677), .Z(n10680) );
  AND U12136 ( .A(a[46]), .B(b[34]), .Z(n10679) );
  NANDN U12137 ( .A(n10680), .B(n10679), .Z(n10905) );
  XOR U12138 ( .A(n10680), .B(n10679), .Z(n11245) );
  XOR U12139 ( .A(n10682), .B(n10681), .Z(n10684) );
  AND U12140 ( .A(a[44]), .B(b[34]), .Z(n10683) );
  NANDN U12141 ( .A(n10684), .B(n10683), .Z(n10897) );
  XOR U12142 ( .A(n10684), .B(n10683), .Z(n11233) );
  XOR U12143 ( .A(n10686), .B(n10685), .Z(n10688) );
  AND U12144 ( .A(a[42]), .B(b[34]), .Z(n10687) );
  NANDN U12145 ( .A(n10688), .B(n10687), .Z(n10889) );
  XOR U12146 ( .A(n10688), .B(n10687), .Z(n11221) );
  XOR U12147 ( .A(n10690), .B(n10689), .Z(n10692) );
  AND U12148 ( .A(a[39]), .B(b[34]), .Z(n10691) );
  NANDN U12149 ( .A(n10692), .B(n10691), .Z(n10875) );
  XOR U12150 ( .A(n10692), .B(n10691), .Z(n11203) );
  NAND U12151 ( .A(a[38]), .B(b[34]), .Z(n10870) );
  XNOR U12152 ( .A(n10694), .B(n10693), .Z(n10871) );
  NANDN U12153 ( .A(n10870), .B(n10871), .Z(n10873) );
  XOR U12154 ( .A(n10696), .B(n10695), .Z(n10698) );
  AND U12155 ( .A(a[36]), .B(b[34]), .Z(n10697) );
  NANDN U12156 ( .A(n10698), .B(n10697), .Z(n10863) );
  XOR U12157 ( .A(n10698), .B(n10697), .Z(n11183) );
  XOR U12158 ( .A(n10700), .B(n10699), .Z(n11179) );
  NAND U12159 ( .A(a[35]), .B(b[34]), .Z(n11180) );
  NAND U12160 ( .A(a[33]), .B(b[34]), .Z(n10852) );
  XNOR U12161 ( .A(n10702), .B(n10701), .Z(n10853) );
  NANDN U12162 ( .A(n10852), .B(n10853), .Z(n10855) );
  NAND U12163 ( .A(a[32]), .B(b[34]), .Z(n10848) );
  XNOR U12164 ( .A(n10704), .B(n10703), .Z(n10849) );
  NANDN U12165 ( .A(n10848), .B(n10849), .Z(n10851) );
  NAND U12166 ( .A(a[30]), .B(b[34]), .Z(n10838) );
  XOR U12167 ( .A(n10706), .B(n10705), .Z(n11137) );
  XNOR U12168 ( .A(n10708), .B(n10707), .Z(n11126) );
  XNOR U12169 ( .A(n10712), .B(n10711), .Z(n11109) );
  XNOR U12170 ( .A(n10714), .B(n10713), .Z(n11100) );
  XNOR U12171 ( .A(n10716), .B(n10715), .Z(n11080) );
  NAND U12172 ( .A(a[14]), .B(b[34]), .Z(n10778) );
  XNOR U12173 ( .A(n10718), .B(n10717), .Z(n11053) );
  XNOR U12174 ( .A(n10720), .B(n10719), .Z(n11041) );
  NAND U12175 ( .A(a[8]), .B(b[34]), .Z(n10758) );
  XOR U12176 ( .A(n10722), .B(n10721), .Z(n10743) );
  AND U12177 ( .A(a[0]), .B(b[34]), .Z(n11429) );
  AND U12178 ( .A(a[1]), .B(b[35]), .Z(n10726) );
  AND U12179 ( .A(n11429), .B(n10726), .Z(n10723) );
  NAND U12180 ( .A(a[2]), .B(n10723), .Z(n10730) );
  NAND U12181 ( .A(b[35]), .B(a[1]), .Z(n10724) );
  XOR U12182 ( .A(n10725), .B(n10724), .Z(n11002) );
  NAND U12183 ( .A(n10726), .B(a[0]), .Z(n10727) );
  XNOR U12184 ( .A(a[2]), .B(n10727), .Z(n10728) );
  AND U12185 ( .A(b[34]), .B(n10728), .Z(n11003) );
  NANDN U12186 ( .A(n11002), .B(n11003), .Z(n10729) );
  AND U12187 ( .A(n10730), .B(n10729), .Z(n10733) );
  NANDN U12188 ( .A(n10733), .B(n10734), .Z(n10736) );
  AND U12189 ( .A(a[3]), .B(b[34]), .Z(n11009) );
  NAND U12190 ( .A(n11009), .B(n11008), .Z(n10735) );
  AND U12191 ( .A(n10736), .B(n10735), .Z(n10739) );
  AND U12192 ( .A(a[4]), .B(b[34]), .Z(n10740) );
  NANDN U12193 ( .A(n10739), .B(n10740), .Z(n10742) );
  XOR U12194 ( .A(n10738), .B(n10737), .Z(n11015) );
  NAND U12195 ( .A(n11015), .B(n11014), .Z(n10741) );
  AND U12196 ( .A(n10742), .B(n10741), .Z(n10744) );
  NANDN U12197 ( .A(n10743), .B(n10744), .Z(n10746) );
  AND U12198 ( .A(a[5]), .B(b[34]), .Z(n11022) );
  NANDN U12199 ( .A(n11022), .B(n11023), .Z(n10745) );
  NAND U12200 ( .A(n10746), .B(n10745), .Z(n10749) );
  AND U12201 ( .A(a[6]), .B(b[34]), .Z(n10750) );
  NANDN U12202 ( .A(n10749), .B(n10750), .Z(n10752) );
  NAND U12203 ( .A(n10993), .B(n10992), .Z(n10751) );
  AND U12204 ( .A(n10752), .B(n10751), .Z(n11029) );
  IV U12205 ( .A(n10755), .Z(n11030) );
  NAND U12206 ( .A(a[7]), .B(b[34]), .Z(n11028) );
  NANDN U12207 ( .A(n10758), .B(n10759), .Z(n10761) );
  NAND U12208 ( .A(n11034), .B(n11033), .Z(n10760) );
  NAND U12209 ( .A(n10761), .B(n10760), .Z(n11042) );
  NAND U12210 ( .A(a[9]), .B(b[34]), .Z(n11044) );
  AND U12211 ( .A(a[10]), .B(b[34]), .Z(n10763) );
  NANDN U12212 ( .A(n10762), .B(n10763), .Z(n10767) );
  XNOR U12213 ( .A(n10763), .B(n10762), .Z(n11048) );
  NAND U12214 ( .A(n11048), .B(n11047), .Z(n10766) );
  NAND U12215 ( .A(n10767), .B(n10766), .Z(n11054) );
  NAND U12216 ( .A(a[11]), .B(b[34]), .Z(n11056) );
  AND U12217 ( .A(a[12]), .B(b[34]), .Z(n10769) );
  NANDN U12218 ( .A(n10768), .B(n10769), .Z(n10773) );
  XOR U12219 ( .A(n10769), .B(n10768), .Z(n11061) );
  XOR U12220 ( .A(n10771), .B(n10770), .Z(n11062) );
  NANDN U12221 ( .A(n11061), .B(n11062), .Z(n10772) );
  NAND U12222 ( .A(n10773), .B(n10772), .Z(n11070) );
  NAND U12223 ( .A(a[13]), .B(b[34]), .Z(n11069) );
  NANDN U12224 ( .A(n10778), .B(n10779), .Z(n10781) );
  XOR U12225 ( .A(n10777), .B(n10776), .Z(n11075) );
  NAND U12226 ( .A(n11075), .B(n11074), .Z(n10780) );
  NAND U12227 ( .A(n10781), .B(n10780), .Z(n11081) );
  NAND U12228 ( .A(a[15]), .B(b[34]), .Z(n11083) );
  AND U12229 ( .A(a[16]), .B(b[34]), .Z(n10783) );
  NANDN U12230 ( .A(n10782), .B(n10783), .Z(n10787) );
  XOR U12231 ( .A(n10783), .B(n10782), .Z(n11088) );
  NANDN U12232 ( .A(n11088), .B(n11089), .Z(n10786) );
  AND U12233 ( .A(n10787), .B(n10786), .Z(n10790) );
  NANDN U12234 ( .A(n10790), .B(n10791), .Z(n10793) );
  AND U12235 ( .A(a[17]), .B(b[34]), .Z(n11097) );
  NAND U12236 ( .A(n11097), .B(n11096), .Z(n10792) );
  AND U12237 ( .A(n10793), .B(n10792), .Z(n10796) );
  AND U12238 ( .A(a[18]), .B(b[34]), .Z(n10797) );
  NANDN U12239 ( .A(n10796), .B(n10797), .Z(n10799) );
  XOR U12240 ( .A(n10795), .B(n10794), .Z(n10991) );
  NAND U12241 ( .A(n10991), .B(n10990), .Z(n10798) );
  NAND U12242 ( .A(n10799), .B(n10798), .Z(n11101) );
  NAND U12243 ( .A(a[19]), .B(b[34]), .Z(n11102) );
  AND U12244 ( .A(a[20]), .B(b[34]), .Z(n10803) );
  NANDN U12245 ( .A(n10802), .B(n10803), .Z(n10805) );
  XOR U12246 ( .A(n10801), .B(n10800), .Z(n10989) );
  XNOR U12247 ( .A(n10803), .B(n10802), .Z(n10988) );
  NAND U12248 ( .A(n10989), .B(n10988), .Z(n10804) );
  NAND U12249 ( .A(n10805), .B(n10804), .Z(n11110) );
  NAND U12250 ( .A(a[21]), .B(b[34]), .Z(n11112) );
  AND U12251 ( .A(a[22]), .B(b[34]), .Z(n10807) );
  NANDN U12252 ( .A(n10806), .B(n10807), .Z(n10811) );
  XNOR U12253 ( .A(n10807), .B(n10806), .Z(n10987) );
  XOR U12254 ( .A(n10809), .B(n10808), .Z(n10986) );
  NAND U12255 ( .A(n10987), .B(n10986), .Z(n10810) );
  NAND U12256 ( .A(n10811), .B(n10810), .Z(n11116) );
  NAND U12257 ( .A(a[23]), .B(b[34]), .Z(n11118) );
  AND U12258 ( .A(a[24]), .B(b[34]), .Z(n10813) );
  NANDN U12259 ( .A(n10812), .B(n10813), .Z(n10817) );
  XNOR U12260 ( .A(n10813), .B(n10812), .Z(n10985) );
  XOR U12261 ( .A(n10815), .B(n10814), .Z(n10984) );
  NAND U12262 ( .A(n10985), .B(n10984), .Z(n10816) );
  NAND U12263 ( .A(n10817), .B(n10816), .Z(n11127) );
  AND U12264 ( .A(a[25]), .B(b[34]), .Z(n11125) );
  AND U12265 ( .A(a[26]), .B(b[34]), .Z(n10819) );
  NANDN U12266 ( .A(n10818), .B(n10819), .Z(n10823) );
  XNOR U12267 ( .A(n10819), .B(n10818), .Z(n11131) );
  XOR U12268 ( .A(n10821), .B(n10820), .Z(n11130) );
  NAND U12269 ( .A(n11131), .B(n11130), .Z(n10822) );
  NAND U12270 ( .A(n10823), .B(n10822), .Z(n11138) );
  AND U12271 ( .A(a[27]), .B(b[34]), .Z(n11136) );
  AND U12272 ( .A(a[28]), .B(b[34]), .Z(n10825) );
  NANDN U12273 ( .A(n10824), .B(n10825), .Z(n10829) );
  XNOR U12274 ( .A(n10825), .B(n10824), .Z(n11144) );
  XOR U12275 ( .A(n10827), .B(n10826), .Z(n11143) );
  NAND U12276 ( .A(n11144), .B(n11143), .Z(n10828) );
  AND U12277 ( .A(n10829), .B(n10828), .Z(n10833) );
  NAND U12278 ( .A(n10833), .B(n10832), .Z(n10835) );
  AND U12279 ( .A(a[29]), .B(b[34]), .Z(n11152) );
  XOR U12280 ( .A(n10833), .B(n10832), .Z(n11151) );
  NANDN U12281 ( .A(n11152), .B(n11151), .Z(n10834) );
  AND U12282 ( .A(n10835), .B(n10834), .Z(n10839) );
  NANDN U12283 ( .A(n10838), .B(n10839), .Z(n10841) );
  XOR U12284 ( .A(n10837), .B(n10836), .Z(n11156) );
  NAND U12285 ( .A(n11156), .B(n11155), .Z(n10840) );
  AND U12286 ( .A(n10841), .B(n10840), .Z(n10845) );
  AND U12287 ( .A(a[31]), .B(b[34]), .Z(n10844) );
  NANDN U12288 ( .A(n10845), .B(n10844), .Z(n10847) );
  XNOR U12289 ( .A(n10843), .B(n10842), .Z(n10983) );
  XNOR U12290 ( .A(n10845), .B(n10844), .Z(n10982) );
  NAND U12291 ( .A(n10983), .B(n10982), .Z(n10846) );
  AND U12292 ( .A(n10847), .B(n10846), .Z(n11162) );
  XNOR U12293 ( .A(n10849), .B(n10848), .Z(n11161) );
  NANDN U12294 ( .A(n11162), .B(n11161), .Z(n10850) );
  AND U12295 ( .A(n10851), .B(n10850), .Z(n11168) );
  XNOR U12296 ( .A(n10853), .B(n10852), .Z(n11167) );
  NANDN U12297 ( .A(n11168), .B(n11167), .Z(n10854) );
  AND U12298 ( .A(n10855), .B(n10854), .Z(n10857) );
  AND U12299 ( .A(a[34]), .B(b[34]), .Z(n10856) );
  NANDN U12300 ( .A(n10857), .B(n10856), .Z(n10861) );
  XOR U12301 ( .A(n10857), .B(n10856), .Z(n11175) );
  XOR U12302 ( .A(n10859), .B(n10858), .Z(n11176) );
  OR U12303 ( .A(n11175), .B(n11176), .Z(n10860) );
  NAND U12304 ( .A(n10861), .B(n10860), .Z(n11182) );
  NANDN U12305 ( .A(n11183), .B(n11184), .Z(n10862) );
  AND U12306 ( .A(n10863), .B(n10862), .Z(n10867) );
  AND U12307 ( .A(a[37]), .B(b[34]), .Z(n10866) );
  NANDN U12308 ( .A(n10867), .B(n10866), .Z(n10869) );
  XNOR U12309 ( .A(n10865), .B(n10864), .Z(n11192) );
  XNOR U12310 ( .A(n10867), .B(n10866), .Z(n11191) );
  NAND U12311 ( .A(n11192), .B(n11191), .Z(n10868) );
  AND U12312 ( .A(n10869), .B(n10868), .Z(n11196) );
  XNOR U12313 ( .A(n10871), .B(n10870), .Z(n11195) );
  NANDN U12314 ( .A(n11196), .B(n11195), .Z(n10872) );
  AND U12315 ( .A(n10873), .B(n10872), .Z(n11204) );
  OR U12316 ( .A(n11203), .B(n11204), .Z(n10874) );
  AND U12317 ( .A(n10875), .B(n10874), .Z(n10877) );
  AND U12318 ( .A(a[40]), .B(b[34]), .Z(n10876) );
  NANDN U12319 ( .A(n10877), .B(n10876), .Z(n10881) );
  XOR U12320 ( .A(n10877), .B(n10876), .Z(n11209) );
  XOR U12321 ( .A(n10879), .B(n10878), .Z(n11210) );
  OR U12322 ( .A(n11209), .B(n11210), .Z(n10880) );
  AND U12323 ( .A(n10881), .B(n10880), .Z(n10885) );
  XNOR U12324 ( .A(n10883), .B(n10882), .Z(n10884) );
  NANDN U12325 ( .A(n10885), .B(n10884), .Z(n10887) );
  NAND U12326 ( .A(a[41]), .B(b[34]), .Z(n11213) );
  XNOR U12327 ( .A(n10885), .B(n10884), .Z(n11214) );
  NANDN U12328 ( .A(n11213), .B(n11214), .Z(n10886) );
  AND U12329 ( .A(n10887), .B(n10886), .Z(n11222) );
  OR U12330 ( .A(n11221), .B(n11222), .Z(n10888) );
  AND U12331 ( .A(n10889), .B(n10888), .Z(n10891) );
  AND U12332 ( .A(a[43]), .B(b[34]), .Z(n10890) );
  NANDN U12333 ( .A(n10891), .B(n10890), .Z(n10895) );
  XOR U12334 ( .A(n10891), .B(n10890), .Z(n11225) );
  XNOR U12335 ( .A(n10893), .B(n10892), .Z(n11226) );
  NANDN U12336 ( .A(n11225), .B(n11226), .Z(n10894) );
  AND U12337 ( .A(n10895), .B(n10894), .Z(n11234) );
  OR U12338 ( .A(n11233), .B(n11234), .Z(n10896) );
  AND U12339 ( .A(n10897), .B(n10896), .Z(n10901) );
  AND U12340 ( .A(a[45]), .B(b[34]), .Z(n10900) );
  NANDN U12341 ( .A(n10901), .B(n10900), .Z(n10903) );
  XOR U12342 ( .A(n10899), .B(n10898), .Z(n11238) );
  XNOR U12343 ( .A(n10901), .B(n10900), .Z(n11237) );
  NANDN U12344 ( .A(n11238), .B(n11237), .Z(n10902) );
  AND U12345 ( .A(n10903), .B(n10902), .Z(n11246) );
  OR U12346 ( .A(n11245), .B(n11246), .Z(n10904) );
  AND U12347 ( .A(n10905), .B(n10904), .Z(n10909) );
  AND U12348 ( .A(a[47]), .B(b[34]), .Z(n10908) );
  NANDN U12349 ( .A(n10909), .B(n10908), .Z(n10911) );
  XOR U12350 ( .A(n10907), .B(n10906), .Z(n11250) );
  XNOR U12351 ( .A(n10909), .B(n10908), .Z(n11249) );
  NANDN U12352 ( .A(n11250), .B(n11249), .Z(n10910) );
  AND U12353 ( .A(n10911), .B(n10910), .Z(n11258) );
  OR U12354 ( .A(n11257), .B(n11258), .Z(n10912) );
  AND U12355 ( .A(n10913), .B(n10912), .Z(n10915) );
  AND U12356 ( .A(a[49]), .B(b[34]), .Z(n10914) );
  NANDN U12357 ( .A(n10915), .B(n10914), .Z(n10919) );
  XOR U12358 ( .A(n10915), .B(n10914), .Z(n11261) );
  XNOR U12359 ( .A(n10917), .B(n10916), .Z(n11262) );
  NANDN U12360 ( .A(n11261), .B(n11262), .Z(n10918) );
  AND U12361 ( .A(n10919), .B(n10918), .Z(n11270) );
  OR U12362 ( .A(n11269), .B(n11270), .Z(n10920) );
  AND U12363 ( .A(n10921), .B(n10920), .Z(n11276) );
  OR U12364 ( .A(n11275), .B(n11276), .Z(n10922) );
  AND U12365 ( .A(n10923), .B(n10922), .Z(n10925) );
  AND U12366 ( .A(a[52]), .B(b[34]), .Z(n10924) );
  NANDN U12367 ( .A(n10925), .B(n10924), .Z(n10929) );
  XOR U12368 ( .A(n10925), .B(n10924), .Z(n11281) );
  XOR U12369 ( .A(n10927), .B(n10926), .Z(n11282) );
  OR U12370 ( .A(n11281), .B(n11282), .Z(n10928) );
  AND U12371 ( .A(n10929), .B(n10928), .Z(n11288) );
  OR U12372 ( .A(n11287), .B(n11288), .Z(n10930) );
  AND U12373 ( .A(n10931), .B(n10930), .Z(n10932) );
  NANDN U12374 ( .A(n10933), .B(n10932), .Z(n10935) );
  AND U12375 ( .A(a[54]), .B(b[34]), .Z(n11294) );
  XNOR U12376 ( .A(n10933), .B(n10932), .Z(n11293) );
  NANDN U12377 ( .A(n11294), .B(n11293), .Z(n10934) );
  NAND U12378 ( .A(n10935), .B(n10934), .Z(n11297) );
  XNOR U12379 ( .A(n10937), .B(n10936), .Z(n11298) );
  NANDN U12380 ( .A(n11297), .B(n11298), .Z(n10938) );
  AND U12381 ( .A(n10939), .B(n10938), .Z(n10941) );
  AND U12382 ( .A(a[56]), .B(b[34]), .Z(n10940) );
  NANDN U12383 ( .A(n10941), .B(n10940), .Z(n10945) );
  XOR U12384 ( .A(n10941), .B(n10940), .Z(n11303) );
  XNOR U12385 ( .A(n10943), .B(n10942), .Z(n11304) );
  NANDN U12386 ( .A(n11303), .B(n11304), .Z(n10944) );
  AND U12387 ( .A(n10945), .B(n10944), .Z(n11312) );
  OR U12388 ( .A(n11311), .B(n11312), .Z(n10946) );
  AND U12389 ( .A(n10947), .B(n10946), .Z(n10951) );
  AND U12390 ( .A(a[58]), .B(b[34]), .Z(n10950) );
  NANDN U12391 ( .A(n10951), .B(n10950), .Z(n10953) );
  XOR U12392 ( .A(n10949), .B(n10948), .Z(n11317) );
  XNOR U12393 ( .A(n10951), .B(n10950), .Z(n11318) );
  NANDN U12394 ( .A(n11317), .B(n11318), .Z(n10952) );
  AND U12395 ( .A(n10953), .B(n10952), .Z(n11322) );
  XNOR U12396 ( .A(n10955), .B(n10954), .Z(n11321) );
  NANDN U12397 ( .A(n11322), .B(n11321), .Z(n10956) );
  AND U12398 ( .A(n10957), .B(n10956), .Z(n10959) );
  AND U12399 ( .A(a[60]), .B(b[34]), .Z(n10958) );
  NANDN U12400 ( .A(n10959), .B(n10958), .Z(n10963) );
  XOR U12401 ( .A(n10959), .B(n10958), .Z(n11327) );
  XNOR U12402 ( .A(n10961), .B(n10960), .Z(n11328) );
  NANDN U12403 ( .A(n11327), .B(n11328), .Z(n10962) );
  AND U12404 ( .A(n10963), .B(n10962), .Z(n11336) );
  OR U12405 ( .A(n11335), .B(n11336), .Z(n10964) );
  AND U12406 ( .A(n10965), .B(n10964), .Z(n10969) );
  XNOR U12407 ( .A(n10967), .B(n10966), .Z(n10968) );
  NANDN U12408 ( .A(n10969), .B(n10968), .Z(n10971) );
  NAND U12409 ( .A(a[62]), .B(b[34]), .Z(n11339) );
  XNOR U12410 ( .A(n10969), .B(n10968), .Z(n11340) );
  NANDN U12411 ( .A(n11339), .B(n11340), .Z(n10970) );
  AND U12412 ( .A(n10971), .B(n10970), .Z(n10972) );
  NANDN U12413 ( .A(n10973), .B(n10972), .Z(n10977) );
  XOR U12414 ( .A(n10973), .B(n10972), .Z(n11345) );
  XOR U12415 ( .A(n10975), .B(n10974), .Z(n11346) );
  OR U12416 ( .A(n11345), .B(n11346), .Z(n10976) );
  NAND U12417 ( .A(n10977), .B(n10976), .Z(n11347) );
  ANDN U12418 ( .B(n11348), .A(n11347), .Z(n10980) );
  XNOR U12419 ( .A(n10979), .B(n10978), .Z(n10981) );
  XOR U12420 ( .A(n10981), .B(n10980), .Z(n24790) );
  NAND U12421 ( .A(a[63]), .B(b[33]), .Z(n11341) );
  AND U12422 ( .A(a[62]), .B(b[33]), .Z(n11334) );
  NAND U12423 ( .A(a[59]), .B(b[33]), .Z(n11315) );
  AND U12424 ( .A(a[58]), .B(b[33]), .Z(n11310) );
  NAND U12425 ( .A(a[56]), .B(b[33]), .Z(n11299) );
  AND U12426 ( .A(a[55]), .B(b[33]), .Z(n11292) );
  AND U12427 ( .A(a[54]), .B(b[33]), .Z(n11286) );
  AND U12428 ( .A(a[53]), .B(b[33]), .Z(n11280) );
  AND U12429 ( .A(a[52]), .B(b[33]), .Z(n11274) );
  AND U12430 ( .A(a[51]), .B(b[33]), .Z(n11268) );
  NAND U12431 ( .A(a[50]), .B(b[33]), .Z(n11263) );
  AND U12432 ( .A(a[49]), .B(b[33]), .Z(n11256) );
  NAND U12433 ( .A(a[48]), .B(b[33]), .Z(n11251) );
  AND U12434 ( .A(a[47]), .B(b[33]), .Z(n11244) );
  NAND U12435 ( .A(a[46]), .B(b[33]), .Z(n11239) );
  AND U12436 ( .A(a[45]), .B(b[33]), .Z(n11232) );
  NAND U12437 ( .A(a[44]), .B(b[33]), .Z(n11227) );
  AND U12438 ( .A(a[43]), .B(b[33]), .Z(n11220) );
  NAND U12439 ( .A(a[42]), .B(b[33]), .Z(n11215) );
  AND U12440 ( .A(a[41]), .B(b[33]), .Z(n11208) );
  AND U12441 ( .A(a[40]), .B(b[33]), .Z(n11202) );
  NAND U12442 ( .A(a[39]), .B(b[33]), .Z(n11197) );
  AND U12443 ( .A(a[38]), .B(b[33]), .Z(n11190) );
  AND U12444 ( .A(a[35]), .B(b[33]), .Z(n11174) );
  XNOR U12445 ( .A(n10983), .B(n10982), .Z(n11563) );
  AND U12446 ( .A(a[32]), .B(b[33]), .Z(n11562) );
  AND U12447 ( .A(a[31]), .B(b[33]), .Z(n11157) );
  NAND U12448 ( .A(a[28]), .B(b[33]), .Z(n11139) );
  AND U12449 ( .A(a[26]), .B(b[33]), .Z(n11123) );
  XNOR U12450 ( .A(n10985), .B(n10984), .Z(n11534) );
  XNOR U12451 ( .A(n10987), .B(n10986), .Z(n11526) );
  XNOR U12452 ( .A(n10989), .B(n10988), .Z(n11518) );
  XNOR U12453 ( .A(n10991), .B(n10990), .Z(n11512) );
  XNOR U12454 ( .A(n10993), .B(n10992), .Z(n11463) );
  AND U12455 ( .A(a[4]), .B(b[33]), .Z(n11010) );
  AND U12456 ( .A(a[0]), .B(b[33]), .Z(n11710) );
  AND U12457 ( .A(a[1]), .B(b[34]), .Z(n10995) );
  AND U12458 ( .A(n11710), .B(n10995), .Z(n10994) );
  NAND U12459 ( .A(a[2]), .B(n10994), .Z(n11001) );
  NAND U12460 ( .A(n10995), .B(a[0]), .Z(n10996) );
  XNOR U12461 ( .A(a[2]), .B(n10996), .Z(n10997) );
  NAND U12462 ( .A(b[33]), .B(n10997), .Z(n11435) );
  NAND U12463 ( .A(b[34]), .B(a[1]), .Z(n10998) );
  XNOR U12464 ( .A(n10999), .B(n10998), .Z(n11436) );
  NANDN U12465 ( .A(n11435), .B(n11436), .Z(n11000) );
  AND U12466 ( .A(n11001), .B(n11000), .Z(n11004) );
  NANDN U12467 ( .A(n11004), .B(n11005), .Z(n11007) );
  NAND U12468 ( .A(a[3]), .B(b[33]), .Z(n11443) );
  NANDN U12469 ( .A(n11443), .B(n11444), .Z(n11006) );
  AND U12470 ( .A(n11007), .B(n11006), .Z(n11011) );
  NANDN U12471 ( .A(n11010), .B(n11011), .Z(n11013) );
  XOR U12472 ( .A(n11009), .B(n11008), .Z(n11425) );
  NANDN U12473 ( .A(n11425), .B(n11426), .Z(n11012) );
  AND U12474 ( .A(n11013), .B(n11012), .Z(n11017) );
  XOR U12475 ( .A(n11015), .B(n11014), .Z(n11016) );
  NAND U12476 ( .A(n11017), .B(n11016), .Z(n11019) );
  AND U12477 ( .A(a[5]), .B(b[33]), .Z(n11452) );
  XOR U12478 ( .A(n11017), .B(n11016), .Z(n11451) );
  NAND U12479 ( .A(n11452), .B(n11451), .Z(n11018) );
  AND U12480 ( .A(n11019), .B(n11018), .Z(n11020) );
  AND U12481 ( .A(a[6]), .B(b[33]), .Z(n11021) );
  NANDN U12482 ( .A(n11020), .B(n11021), .Z(n11025) );
  NAND U12483 ( .A(n11457), .B(n11458), .Z(n11024) );
  NAND U12484 ( .A(n11025), .B(n11024), .Z(n11464) );
  NAND U12485 ( .A(a[7]), .B(b[33]), .Z(n11466) );
  AND U12486 ( .A(a[8]), .B(b[33]), .Z(n11026) );
  NANDN U12487 ( .A(n11027), .B(n11026), .Z(n11032) );
  XOR U12488 ( .A(n11027), .B(n11026), .Z(n11471) );
  NANDN U12489 ( .A(n11471), .B(n11472), .Z(n11031) );
  AND U12490 ( .A(n11032), .B(n11031), .Z(n11035) );
  XOR U12491 ( .A(n11034), .B(n11033), .Z(n11036) );
  NANDN U12492 ( .A(n11035), .B(n11036), .Z(n11038) );
  NAND U12493 ( .A(a[9]), .B(b[33]), .Z(n11479) );
  NANDN U12494 ( .A(n11479), .B(n11480), .Z(n11037) );
  AND U12495 ( .A(n11038), .B(n11037), .Z(n11039) );
  AND U12496 ( .A(a[10]), .B(b[33]), .Z(n11040) );
  NANDN U12497 ( .A(n11039), .B(n11040), .Z(n11046) );
  XNOR U12498 ( .A(n11042), .B(n11041), .Z(n11043) );
  XNOR U12499 ( .A(n11044), .B(n11043), .Z(n11423) );
  NAND U12500 ( .A(n11424), .B(n11423), .Z(n11045) );
  AND U12501 ( .A(n11046), .B(n11045), .Z(n11049) );
  XOR U12502 ( .A(n11048), .B(n11047), .Z(n11050) );
  NANDN U12503 ( .A(n11049), .B(n11050), .Z(n11052) );
  NAND U12504 ( .A(a[11]), .B(b[33]), .Z(n11485) );
  NANDN U12505 ( .A(n11485), .B(n11486), .Z(n11051) );
  AND U12506 ( .A(n11052), .B(n11051), .Z(n11057) );
  AND U12507 ( .A(a[12]), .B(b[33]), .Z(n11058) );
  NANDN U12508 ( .A(n11057), .B(n11058), .Z(n11060) );
  XNOR U12509 ( .A(n11054), .B(n11053), .Z(n11055) );
  XNOR U12510 ( .A(n11056), .B(n11055), .Z(n11490) );
  NAND U12511 ( .A(n11490), .B(n11489), .Z(n11059) );
  AND U12512 ( .A(n11060), .B(n11059), .Z(n11063) );
  NANDN U12513 ( .A(n11063), .B(n11064), .Z(n11066) );
  NAND U12514 ( .A(a[13]), .B(b[33]), .Z(n11492) );
  NANDN U12515 ( .A(n11492), .B(n11493), .Z(n11065) );
  AND U12516 ( .A(n11066), .B(n11065), .Z(n11067) );
  AND U12517 ( .A(a[14]), .B(b[33]), .Z(n11068) );
  NANDN U12518 ( .A(n11067), .B(n11068), .Z(n11073) );
  NAND U12519 ( .A(n11422), .B(n11421), .Z(n11072) );
  AND U12520 ( .A(n11073), .B(n11072), .Z(n11076) );
  XOR U12521 ( .A(n11075), .B(n11074), .Z(n11077) );
  NANDN U12522 ( .A(n11076), .B(n11077), .Z(n11079) );
  NAND U12523 ( .A(a[15]), .B(b[33]), .Z(n11500) );
  NANDN U12524 ( .A(n11500), .B(n11501), .Z(n11078) );
  AND U12525 ( .A(n11079), .B(n11078), .Z(n11084) );
  AND U12526 ( .A(a[16]), .B(b[33]), .Z(n11085) );
  NANDN U12527 ( .A(n11084), .B(n11085), .Z(n11087) );
  XNOR U12528 ( .A(n11081), .B(n11080), .Z(n11082) );
  XNOR U12529 ( .A(n11083), .B(n11082), .Z(n11420) );
  NAND U12530 ( .A(n11420), .B(n11419), .Z(n11086) );
  AND U12531 ( .A(n11087), .B(n11086), .Z(n11090) );
  NANDN U12532 ( .A(n11090), .B(n11091), .Z(n11093) );
  NAND U12533 ( .A(a[17]), .B(b[33]), .Z(n11504) );
  NANDN U12534 ( .A(n11504), .B(n11505), .Z(n11092) );
  AND U12535 ( .A(n11093), .B(n11092), .Z(n11094) );
  AND U12536 ( .A(a[18]), .B(b[33]), .Z(n11095) );
  NANDN U12537 ( .A(n11094), .B(n11095), .Z(n11099) );
  XOR U12538 ( .A(n11097), .B(n11096), .Z(n11417) );
  NAND U12539 ( .A(n11418), .B(n11417), .Z(n11098) );
  NAND U12540 ( .A(n11099), .B(n11098), .Z(n11513) );
  NAND U12541 ( .A(a[19]), .B(b[33]), .Z(n11515) );
  AND U12542 ( .A(a[20]), .B(b[33]), .Z(n11103) );
  NANDN U12543 ( .A(n11104), .B(n11103), .Z(n11106) );
  XNOR U12544 ( .A(n11104), .B(n11103), .Z(n11415) );
  NAND U12545 ( .A(n11416), .B(n11415), .Z(n11105) );
  NAND U12546 ( .A(n11106), .B(n11105), .Z(n11519) );
  NAND U12547 ( .A(a[21]), .B(b[33]), .Z(n11521) );
  AND U12548 ( .A(a[22]), .B(b[33]), .Z(n11107) );
  NANDN U12549 ( .A(n11108), .B(n11107), .Z(n11114) );
  XNOR U12550 ( .A(n11108), .B(n11107), .Z(n11414) );
  XNOR U12551 ( .A(n11110), .B(n11109), .Z(n11111) );
  XNOR U12552 ( .A(n11112), .B(n11111), .Z(n11413) );
  NAND U12553 ( .A(n11414), .B(n11413), .Z(n11113) );
  NAND U12554 ( .A(n11114), .B(n11113), .Z(n11527) );
  NAND U12555 ( .A(a[23]), .B(b[33]), .Z(n11529) );
  AND U12556 ( .A(a[24]), .B(b[33]), .Z(n11119) );
  NANDN U12557 ( .A(n11120), .B(n11119), .Z(n11122) );
  XNOR U12558 ( .A(n11116), .B(n11115), .Z(n11117) );
  XNOR U12559 ( .A(n11118), .B(n11117), .Z(n11412) );
  XNOR U12560 ( .A(n11120), .B(n11119), .Z(n11411) );
  NAND U12561 ( .A(n11412), .B(n11411), .Z(n11121) );
  NAND U12562 ( .A(n11122), .B(n11121), .Z(n11535) );
  NAND U12563 ( .A(a[25]), .B(b[33]), .Z(n11537) );
  NANDN U12564 ( .A(n11123), .B(n11124), .Z(n11129) );
  NAND U12565 ( .A(n11409), .B(n11410), .Z(n11128) );
  AND U12566 ( .A(n11129), .B(n11128), .Z(n11132) );
  XNOR U12567 ( .A(n11131), .B(n11130), .Z(n11133) );
  NANDN U12568 ( .A(n11132), .B(n11133), .Z(n11135) );
  AND U12569 ( .A(a[27]), .B(b[33]), .Z(n11544) );
  NANDN U12570 ( .A(n11544), .B(n11545), .Z(n11134) );
  AND U12571 ( .A(n11135), .B(n11134), .Z(n11140) );
  NANDN U12572 ( .A(n11139), .B(n11140), .Z(n11142) );
  NAND U12573 ( .A(n11408), .B(n11407), .Z(n11141) );
  AND U12574 ( .A(n11142), .B(n11141), .Z(n11145) );
  XOR U12575 ( .A(n11144), .B(n11143), .Z(n11146) );
  NANDN U12576 ( .A(n11145), .B(n11146), .Z(n11148) );
  NAND U12577 ( .A(a[29]), .B(b[33]), .Z(n11550) );
  NANDN U12578 ( .A(n11550), .B(n11551), .Z(n11147) );
  AND U12579 ( .A(n11148), .B(n11147), .Z(n11149) );
  AND U12580 ( .A(a[30]), .B(b[33]), .Z(n11150) );
  NANDN U12581 ( .A(n11149), .B(n11150), .Z(n11154) );
  XOR U12582 ( .A(n11152), .B(n11151), .Z(n11405) );
  NAND U12583 ( .A(n11406), .B(n11405), .Z(n11153) );
  AND U12584 ( .A(n11154), .B(n11153), .Z(n11158) );
  NANDN U12585 ( .A(n11157), .B(n11158), .Z(n11160) );
  XOR U12586 ( .A(n11156), .B(n11155), .Z(n11556) );
  NANDN U12587 ( .A(n11556), .B(n11557), .Z(n11159) );
  NAND U12588 ( .A(n11160), .B(n11159), .Z(n11565) );
  AND U12589 ( .A(a[33]), .B(b[33]), .Z(n11163) );
  NANDN U12590 ( .A(n11164), .B(n11163), .Z(n11166) );
  XOR U12591 ( .A(n11162), .B(n11161), .Z(n11403) );
  XNOR U12592 ( .A(n11164), .B(n11163), .Z(n11404) );
  NANDN U12593 ( .A(n11403), .B(n11404), .Z(n11165) );
  AND U12594 ( .A(n11166), .B(n11165), .Z(n11170) );
  AND U12595 ( .A(a[34]), .B(b[33]), .Z(n11169) );
  NANDN U12596 ( .A(n11170), .B(n11169), .Z(n11172) );
  XOR U12597 ( .A(n11168), .B(n11167), .Z(n11572) );
  XNOR U12598 ( .A(n11170), .B(n11169), .Z(n11573) );
  NANDN U12599 ( .A(n11572), .B(n11573), .Z(n11171) );
  AND U12600 ( .A(n11172), .B(n11171), .Z(n11173) );
  NANDN U12601 ( .A(n11174), .B(n11173), .Z(n11178) );
  XOR U12602 ( .A(n11174), .B(n11173), .Z(n11399) );
  XOR U12603 ( .A(n11176), .B(n11175), .Z(n11400) );
  OR U12604 ( .A(n11399), .B(n11400), .Z(n11177) );
  NAND U12605 ( .A(n11178), .B(n11177), .Z(n11581) );
  AND U12606 ( .A(a[36]), .B(b[33]), .Z(n11580) );
  XOR U12607 ( .A(n11180), .B(n11179), .Z(n11181) );
  XNOR U12608 ( .A(n11182), .B(n11181), .Z(n11583) );
  AND U12609 ( .A(a[37]), .B(b[33]), .Z(n11185) );
  NANDN U12610 ( .A(n11186), .B(n11185), .Z(n11188) );
  XOR U12611 ( .A(n11184), .B(n11183), .Z(n11395) );
  XNOR U12612 ( .A(n11186), .B(n11185), .Z(n11396) );
  NANDN U12613 ( .A(n11395), .B(n11396), .Z(n11187) );
  AND U12614 ( .A(n11188), .B(n11187), .Z(n11189) );
  NANDN U12615 ( .A(n11190), .B(n11189), .Z(n11194) );
  XOR U12616 ( .A(n11190), .B(n11189), .Z(n11393) );
  XOR U12617 ( .A(n11192), .B(n11191), .Z(n11394) );
  OR U12618 ( .A(n11393), .B(n11394), .Z(n11193) );
  AND U12619 ( .A(n11194), .B(n11193), .Z(n11198) );
  NANDN U12620 ( .A(n11197), .B(n11198), .Z(n11200) );
  XOR U12621 ( .A(n11196), .B(n11195), .Z(n11391) );
  XNOR U12622 ( .A(n11198), .B(n11197), .Z(n11392) );
  NANDN U12623 ( .A(n11391), .B(n11392), .Z(n11199) );
  AND U12624 ( .A(n11200), .B(n11199), .Z(n11201) );
  NANDN U12625 ( .A(n11202), .B(n11201), .Z(n11206) );
  XOR U12626 ( .A(n11202), .B(n11201), .Z(n11389) );
  XOR U12627 ( .A(n11204), .B(n11203), .Z(n11390) );
  OR U12628 ( .A(n11389), .B(n11390), .Z(n11205) );
  NAND U12629 ( .A(n11206), .B(n11205), .Z(n11207) );
  NANDN U12630 ( .A(n11208), .B(n11207), .Z(n11212) );
  XOR U12631 ( .A(n11208), .B(n11207), .Z(n11387) );
  XOR U12632 ( .A(n11210), .B(n11209), .Z(n11388) );
  OR U12633 ( .A(n11387), .B(n11388), .Z(n11211) );
  AND U12634 ( .A(n11212), .B(n11211), .Z(n11216) );
  NANDN U12635 ( .A(n11215), .B(n11216), .Z(n11218) );
  XOR U12636 ( .A(n11214), .B(n11213), .Z(n11606) );
  XNOR U12637 ( .A(n11216), .B(n11215), .Z(n11607) );
  NANDN U12638 ( .A(n11606), .B(n11607), .Z(n11217) );
  AND U12639 ( .A(n11218), .B(n11217), .Z(n11219) );
  NANDN U12640 ( .A(n11220), .B(n11219), .Z(n11224) );
  XOR U12641 ( .A(n11220), .B(n11219), .Z(n11383) );
  XOR U12642 ( .A(n11222), .B(n11221), .Z(n11384) );
  OR U12643 ( .A(n11383), .B(n11384), .Z(n11223) );
  AND U12644 ( .A(n11224), .B(n11223), .Z(n11228) );
  NANDN U12645 ( .A(n11227), .B(n11228), .Z(n11230) );
  XOR U12646 ( .A(n11226), .B(n11225), .Z(n11614) );
  XNOR U12647 ( .A(n11228), .B(n11227), .Z(n11615) );
  NANDN U12648 ( .A(n11614), .B(n11615), .Z(n11229) );
  AND U12649 ( .A(n11230), .B(n11229), .Z(n11231) );
  NANDN U12650 ( .A(n11232), .B(n11231), .Z(n11236) );
  XOR U12651 ( .A(n11232), .B(n11231), .Z(n11381) );
  XOR U12652 ( .A(n11234), .B(n11233), .Z(n11382) );
  OR U12653 ( .A(n11381), .B(n11382), .Z(n11235) );
  AND U12654 ( .A(n11236), .B(n11235), .Z(n11240) );
  NANDN U12655 ( .A(n11239), .B(n11240), .Z(n11242) );
  XOR U12656 ( .A(n11238), .B(n11237), .Z(n11624) );
  XNOR U12657 ( .A(n11240), .B(n11239), .Z(n11625) );
  NANDN U12658 ( .A(n11624), .B(n11625), .Z(n11241) );
  AND U12659 ( .A(n11242), .B(n11241), .Z(n11243) );
  NANDN U12660 ( .A(n11244), .B(n11243), .Z(n11248) );
  XOR U12661 ( .A(n11244), .B(n11243), .Z(n11377) );
  XOR U12662 ( .A(n11246), .B(n11245), .Z(n11378) );
  OR U12663 ( .A(n11377), .B(n11378), .Z(n11247) );
  AND U12664 ( .A(n11248), .B(n11247), .Z(n11252) );
  NANDN U12665 ( .A(n11251), .B(n11252), .Z(n11254) );
  XOR U12666 ( .A(n11250), .B(n11249), .Z(n11632) );
  XNOR U12667 ( .A(n11252), .B(n11251), .Z(n11633) );
  NANDN U12668 ( .A(n11632), .B(n11633), .Z(n11253) );
  AND U12669 ( .A(n11254), .B(n11253), .Z(n11255) );
  NANDN U12670 ( .A(n11256), .B(n11255), .Z(n11260) );
  XOR U12671 ( .A(n11256), .B(n11255), .Z(n11373) );
  XOR U12672 ( .A(n11258), .B(n11257), .Z(n11374) );
  OR U12673 ( .A(n11373), .B(n11374), .Z(n11259) );
  AND U12674 ( .A(n11260), .B(n11259), .Z(n11264) );
  NANDN U12675 ( .A(n11263), .B(n11264), .Z(n11266) );
  XOR U12676 ( .A(n11262), .B(n11261), .Z(n11640) );
  XNOR U12677 ( .A(n11264), .B(n11263), .Z(n11641) );
  NANDN U12678 ( .A(n11640), .B(n11641), .Z(n11265) );
  AND U12679 ( .A(n11266), .B(n11265), .Z(n11267) );
  NANDN U12680 ( .A(n11268), .B(n11267), .Z(n11272) );
  XOR U12681 ( .A(n11268), .B(n11267), .Z(n11369) );
  XOR U12682 ( .A(n11270), .B(n11269), .Z(n11370) );
  OR U12683 ( .A(n11369), .B(n11370), .Z(n11271) );
  NAND U12684 ( .A(n11272), .B(n11271), .Z(n11273) );
  NANDN U12685 ( .A(n11274), .B(n11273), .Z(n11278) );
  XOR U12686 ( .A(n11274), .B(n11273), .Z(n11367) );
  XOR U12687 ( .A(n11276), .B(n11275), .Z(n11368) );
  OR U12688 ( .A(n11367), .B(n11368), .Z(n11277) );
  NAND U12689 ( .A(n11278), .B(n11277), .Z(n11279) );
  NANDN U12690 ( .A(n11280), .B(n11279), .Z(n11284) );
  XOR U12691 ( .A(n11280), .B(n11279), .Z(n11363) );
  XOR U12692 ( .A(n11282), .B(n11281), .Z(n11364) );
  OR U12693 ( .A(n11363), .B(n11364), .Z(n11283) );
  NAND U12694 ( .A(n11284), .B(n11283), .Z(n11285) );
  NANDN U12695 ( .A(n11286), .B(n11285), .Z(n11290) );
  XOR U12696 ( .A(n11286), .B(n11285), .Z(n11361) );
  XOR U12697 ( .A(n11288), .B(n11287), .Z(n11362) );
  OR U12698 ( .A(n11361), .B(n11362), .Z(n11289) );
  NAND U12699 ( .A(n11290), .B(n11289), .Z(n11291) );
  NANDN U12700 ( .A(n11292), .B(n11291), .Z(n11296) );
  XNOR U12701 ( .A(n11292), .B(n11291), .Z(n11360) );
  XNOR U12702 ( .A(n11294), .B(n11293), .Z(n11359) );
  NAND U12703 ( .A(n11360), .B(n11359), .Z(n11295) );
  AND U12704 ( .A(n11296), .B(n11295), .Z(n11300) );
  NANDN U12705 ( .A(n11299), .B(n11300), .Z(n11302) );
  XOR U12706 ( .A(n11298), .B(n11297), .Z(n11662) );
  XNOR U12707 ( .A(n11300), .B(n11299), .Z(n11663) );
  NANDN U12708 ( .A(n11662), .B(n11663), .Z(n11301) );
  AND U12709 ( .A(n11302), .B(n11301), .Z(n11306) );
  AND U12710 ( .A(a[57]), .B(b[33]), .Z(n11305) );
  NANDN U12711 ( .A(n11306), .B(n11305), .Z(n11308) );
  XOR U12712 ( .A(n11304), .B(n11303), .Z(n11357) );
  XNOR U12713 ( .A(n11306), .B(n11305), .Z(n11358) );
  NANDN U12714 ( .A(n11357), .B(n11358), .Z(n11307) );
  AND U12715 ( .A(n11308), .B(n11307), .Z(n11309) );
  NANDN U12716 ( .A(n11310), .B(n11309), .Z(n11314) );
  XOR U12717 ( .A(n11310), .B(n11309), .Z(n11672) );
  XOR U12718 ( .A(n11312), .B(n11311), .Z(n11673) );
  OR U12719 ( .A(n11672), .B(n11673), .Z(n11313) );
  AND U12720 ( .A(n11314), .B(n11313), .Z(n11316) );
  NANDN U12721 ( .A(n11315), .B(n11316), .Z(n11320) );
  XOR U12722 ( .A(n11316), .B(n11315), .Z(n11355) );
  XNOR U12723 ( .A(n11318), .B(n11317), .Z(n11356) );
  NANDN U12724 ( .A(n11355), .B(n11356), .Z(n11319) );
  AND U12725 ( .A(n11320), .B(n11319), .Z(n11324) );
  AND U12726 ( .A(a[60]), .B(b[33]), .Z(n11323) );
  NANDN U12727 ( .A(n11324), .B(n11323), .Z(n11326) );
  XOR U12728 ( .A(n11322), .B(n11321), .Z(n11682) );
  XNOR U12729 ( .A(n11324), .B(n11323), .Z(n11683) );
  NANDN U12730 ( .A(n11682), .B(n11683), .Z(n11325) );
  AND U12731 ( .A(n11326), .B(n11325), .Z(n11330) );
  AND U12732 ( .A(a[61]), .B(b[33]), .Z(n11329) );
  NANDN U12733 ( .A(n11330), .B(n11329), .Z(n11332) );
  XOR U12734 ( .A(n11328), .B(n11327), .Z(n11353) );
  XNOR U12735 ( .A(n11330), .B(n11329), .Z(n11354) );
  NANDN U12736 ( .A(n11353), .B(n11354), .Z(n11331) );
  AND U12737 ( .A(n11332), .B(n11331), .Z(n11333) );
  NANDN U12738 ( .A(n11334), .B(n11333), .Z(n11338) );
  XOR U12739 ( .A(n11334), .B(n11333), .Z(n11351) );
  XOR U12740 ( .A(n11336), .B(n11335), .Z(n11352) );
  OR U12741 ( .A(n11351), .B(n11352), .Z(n11337) );
  AND U12742 ( .A(n11338), .B(n11337), .Z(n11342) );
  NANDN U12743 ( .A(n11341), .B(n11342), .Z(n11344) );
  XOR U12744 ( .A(n11340), .B(n11339), .Z(n11349) );
  XNOR U12745 ( .A(n11342), .B(n11341), .Z(n11350) );
  NANDN U12746 ( .A(n11349), .B(n11350), .Z(n11343) );
  NAND U12747 ( .A(n11344), .B(n11343), .Z(n22546) );
  XOR U12748 ( .A(n11346), .B(n11345), .Z(n22547) );
  ANDN U12749 ( .B(n22546), .A(n22547), .Z(n22548) );
  XNOR U12750 ( .A(n11348), .B(n11347), .Z(n22549) );
  XOR U12751 ( .A(n11350), .B(n11349), .Z(n12050) );
  XOR U12752 ( .A(n11352), .B(n11351), .Z(n11693) );
  NAND U12753 ( .A(a[62]), .B(b[32]), .Z(n11688) );
  XNOR U12754 ( .A(n11354), .B(n11353), .Z(n11689) );
  NANDN U12755 ( .A(n11688), .B(n11689), .Z(n11691) );
  NAND U12756 ( .A(a[60]), .B(b[32]), .Z(n11678) );
  XNOR U12757 ( .A(n11356), .B(n11355), .Z(n11679) );
  NANDN U12758 ( .A(n11678), .B(n11679), .Z(n11681) );
  NAND U12759 ( .A(a[58]), .B(b[32]), .Z(n11668) );
  XNOR U12760 ( .A(n11358), .B(n11357), .Z(n11669) );
  NANDN U12761 ( .A(n11668), .B(n11669), .Z(n11671) );
  XOR U12762 ( .A(n11360), .B(n11359), .Z(n11659) );
  AND U12763 ( .A(a[56]), .B(b[32]), .Z(n11658) );
  NANDN U12764 ( .A(n11659), .B(n11658), .Z(n11661) );
  XOR U12765 ( .A(n11362), .B(n11361), .Z(n11655) );
  XOR U12766 ( .A(n11364), .B(n11363), .Z(n11366) );
  AND U12767 ( .A(a[54]), .B(b[32]), .Z(n11365) );
  NANDN U12768 ( .A(n11366), .B(n11365), .Z(n11653) );
  XOR U12769 ( .A(n11366), .B(n11365), .Z(n11998) );
  XOR U12770 ( .A(n11368), .B(n11367), .Z(n11649) );
  XOR U12771 ( .A(n11370), .B(n11369), .Z(n11372) );
  AND U12772 ( .A(a[52]), .B(b[32]), .Z(n11371) );
  NANDN U12773 ( .A(n11372), .B(n11371), .Z(n11647) );
  XOR U12774 ( .A(n11372), .B(n11371), .Z(n11986) );
  XOR U12775 ( .A(n11374), .B(n11373), .Z(n11376) );
  AND U12776 ( .A(a[50]), .B(b[32]), .Z(n11375) );
  NANDN U12777 ( .A(n11376), .B(n11375), .Z(n11639) );
  XOR U12778 ( .A(n11376), .B(n11375), .Z(n11974) );
  XOR U12779 ( .A(n11378), .B(n11377), .Z(n11380) );
  AND U12780 ( .A(a[48]), .B(b[32]), .Z(n11379) );
  NANDN U12781 ( .A(n11380), .B(n11379), .Z(n11631) );
  XOR U12782 ( .A(n11380), .B(n11379), .Z(n11962) );
  XOR U12783 ( .A(n11382), .B(n11381), .Z(n11621) );
  AND U12784 ( .A(a[46]), .B(b[32]), .Z(n11620) );
  NANDN U12785 ( .A(n11621), .B(n11620), .Z(n11623) );
  XOR U12786 ( .A(n11384), .B(n11383), .Z(n11386) );
  AND U12787 ( .A(a[44]), .B(b[32]), .Z(n11385) );
  NANDN U12788 ( .A(n11386), .B(n11385), .Z(n11613) );
  XOR U12789 ( .A(n11386), .B(n11385), .Z(n11938) );
  XOR U12790 ( .A(n11388), .B(n11387), .Z(n11603) );
  AND U12791 ( .A(a[42]), .B(b[32]), .Z(n11602) );
  NANDN U12792 ( .A(n11603), .B(n11602), .Z(n11605) );
  XOR U12793 ( .A(n11390), .B(n11389), .Z(n11599) );
  NAND U12794 ( .A(a[40]), .B(b[32]), .Z(n11594) );
  XNOR U12795 ( .A(n11392), .B(n11391), .Z(n11595) );
  NANDN U12796 ( .A(n11594), .B(n11595), .Z(n11597) );
  XOR U12797 ( .A(n11394), .B(n11393), .Z(n11591) );
  NAND U12798 ( .A(a[38]), .B(b[32]), .Z(n11397) );
  XNOR U12799 ( .A(n11396), .B(n11395), .Z(n11398) );
  NANDN U12800 ( .A(n11397), .B(n11398), .Z(n11589) );
  XOR U12801 ( .A(n11398), .B(n11397), .Z(n11900) );
  XOR U12802 ( .A(n11400), .B(n11399), .Z(n11402) );
  AND U12803 ( .A(a[36]), .B(b[32]), .Z(n11401) );
  NANDN U12804 ( .A(n11402), .B(n11401), .Z(n11579) );
  XOR U12805 ( .A(n11402), .B(n11401), .Z(n11890) );
  NAND U12806 ( .A(a[34]), .B(b[32]), .Z(n11568) );
  XNOR U12807 ( .A(n11404), .B(n11403), .Z(n11569) );
  NANDN U12808 ( .A(n11568), .B(n11569), .Z(n11571) );
  AND U12809 ( .A(a[33]), .B(b[32]), .Z(n11561) );
  XNOR U12810 ( .A(n11406), .B(n11405), .Z(n11862) );
  XNOR U12811 ( .A(n11408), .B(n11407), .Z(n11854) );
  NAND U12812 ( .A(a[28]), .B(b[32]), .Z(n11542) );
  AND U12813 ( .A(a[27]), .B(b[32]), .Z(n11847) );
  XOR U12814 ( .A(n11410), .B(n11409), .Z(n11845) );
  XNOR U12815 ( .A(n11412), .B(n11411), .Z(n11839) );
  XNOR U12816 ( .A(n11414), .B(n11413), .Z(n11828) );
  XNOR U12817 ( .A(n11416), .B(n11415), .Z(n11820) );
  XNOR U12818 ( .A(n11418), .B(n11417), .Z(n11814) );
  XNOR U12819 ( .A(n11420), .B(n11419), .Z(n11803) );
  XNOR U12820 ( .A(n11422), .B(n11421), .Z(n11794) );
  NAND U12821 ( .A(a[14]), .B(b[32]), .Z(n11494) );
  XNOR U12822 ( .A(n11424), .B(n11423), .Z(n11771) );
  AND U12823 ( .A(a[0]), .B(b[32]), .Z(n12130) );
  AND U12824 ( .A(a[1]), .B(b[33]), .Z(n11430) );
  AND U12825 ( .A(n12130), .B(n11430), .Z(n11427) );
  NAND U12826 ( .A(a[2]), .B(n11427), .Z(n11434) );
  NAND U12827 ( .A(b[33]), .B(a[1]), .Z(n11428) );
  XOR U12828 ( .A(n11429), .B(n11428), .Z(n11716) );
  NAND U12829 ( .A(n11430), .B(a[0]), .Z(n11431) );
  XNOR U12830 ( .A(a[2]), .B(n11431), .Z(n11432) );
  AND U12831 ( .A(b[32]), .B(n11432), .Z(n11717) );
  NANDN U12832 ( .A(n11716), .B(n11717), .Z(n11433) );
  AND U12833 ( .A(n11434), .B(n11433), .Z(n11437) );
  NANDN U12834 ( .A(n11437), .B(n11438), .Z(n11440) );
  AND U12835 ( .A(a[3]), .B(b[32]), .Z(n11722) );
  NAND U12836 ( .A(n11723), .B(n11722), .Z(n11439) );
  AND U12837 ( .A(n11440), .B(n11439), .Z(n11441) );
  AND U12838 ( .A(a[4]), .B(b[32]), .Z(n11442) );
  NANDN U12839 ( .A(n11441), .B(n11442), .Z(n11446) );
  NAND U12840 ( .A(n11729), .B(n11728), .Z(n11445) );
  NAND U12841 ( .A(n11446), .B(n11445), .Z(n11447) );
  NAND U12842 ( .A(n11448), .B(n11447), .Z(n11450) );
  NAND U12843 ( .A(a[5]), .B(b[32]), .Z(n11734) );
  XOR U12844 ( .A(n11448), .B(n11447), .Z(n11735) );
  NANDN U12845 ( .A(n11734), .B(n11735), .Z(n11449) );
  AND U12846 ( .A(n11450), .B(n11449), .Z(n11453) );
  XOR U12847 ( .A(n11452), .B(n11451), .Z(n11454) );
  NANDN U12848 ( .A(n11453), .B(n11454), .Z(n11456) );
  AND U12849 ( .A(a[6]), .B(b[32]), .Z(n11741) );
  NAND U12850 ( .A(n11741), .B(n11740), .Z(n11455) );
  AND U12851 ( .A(n11456), .B(n11455), .Z(n11460) );
  XNOR U12852 ( .A(n11458), .B(n11457), .Z(n11459) );
  NAND U12853 ( .A(n11460), .B(n11459), .Z(n11462) );
  AND U12854 ( .A(a[7]), .B(b[32]), .Z(n11748) );
  XOR U12855 ( .A(n11460), .B(n11459), .Z(n11749) );
  NANDN U12856 ( .A(n11748), .B(n11749), .Z(n11461) );
  NAND U12857 ( .A(n11462), .B(n11461), .Z(n11467) );
  AND U12858 ( .A(a[8]), .B(b[32]), .Z(n11468) );
  NANDN U12859 ( .A(n11467), .B(n11468), .Z(n11470) );
  XNOR U12860 ( .A(n11464), .B(n11463), .Z(n11465) );
  XOR U12861 ( .A(n11466), .B(n11465), .Z(n11752) );
  NANDN U12862 ( .A(n11752), .B(n11753), .Z(n11469) );
  AND U12863 ( .A(n11470), .B(n11469), .Z(n11473) );
  NANDN U12864 ( .A(n11473), .B(n11474), .Z(n11476) );
  AND U12865 ( .A(a[9]), .B(b[32]), .Z(n11759) );
  NAND U12866 ( .A(n11759), .B(n11758), .Z(n11475) );
  AND U12867 ( .A(n11476), .B(n11475), .Z(n11477) );
  AND U12868 ( .A(a[10]), .B(b[32]), .Z(n11478) );
  NANDN U12869 ( .A(n11477), .B(n11478), .Z(n11482) );
  NAND U12870 ( .A(n11765), .B(n11764), .Z(n11481) );
  NAND U12871 ( .A(n11482), .B(n11481), .Z(n11772) );
  AND U12872 ( .A(a[11]), .B(b[32]), .Z(n11770) );
  AND U12873 ( .A(a[12]), .B(b[32]), .Z(n11484) );
  NANDN U12874 ( .A(n11483), .B(n11484), .Z(n11488) );
  XOR U12875 ( .A(n11484), .B(n11483), .Z(n11773) );
  NANDN U12876 ( .A(n11773), .B(n11774), .Z(n11487) );
  AND U12877 ( .A(n11488), .B(n11487), .Z(n11780) );
  XOR U12878 ( .A(n11490), .B(n11489), .Z(n11491) );
  IV U12879 ( .A(n11491), .Z(n11781) );
  NAND U12880 ( .A(a[13]), .B(b[32]), .Z(n11779) );
  NANDN U12881 ( .A(n11494), .B(n11495), .Z(n11497) );
  NAND U12882 ( .A(n11787), .B(n11786), .Z(n11496) );
  NAND U12883 ( .A(n11497), .B(n11496), .Z(n11795) );
  NAND U12884 ( .A(a[15]), .B(b[32]), .Z(n11797) );
  AND U12885 ( .A(a[16]), .B(b[32]), .Z(n11499) );
  NANDN U12886 ( .A(n11498), .B(n11499), .Z(n11503) );
  XNOR U12887 ( .A(n11499), .B(n11498), .Z(n11801) );
  NAND U12888 ( .A(n11801), .B(n11800), .Z(n11502) );
  NAND U12889 ( .A(n11503), .B(n11502), .Z(n11804) );
  NAND U12890 ( .A(a[17]), .B(b[32]), .Z(n11806) );
  AND U12891 ( .A(a[18]), .B(b[32]), .Z(n11507) );
  NANDN U12892 ( .A(n11506), .B(n11507), .Z(n11509) );
  XNOR U12893 ( .A(n11507), .B(n11506), .Z(n11706) );
  NAND U12894 ( .A(n11707), .B(n11706), .Z(n11508) );
  NAND U12895 ( .A(n11509), .B(n11508), .Z(n11815) );
  AND U12896 ( .A(a[19]), .B(b[32]), .Z(n11813) );
  AND U12897 ( .A(a[20]), .B(b[32]), .Z(n11511) );
  NANDN U12898 ( .A(n11510), .B(n11511), .Z(n11517) );
  XNOR U12899 ( .A(n11511), .B(n11510), .Z(n11819) );
  XNOR U12900 ( .A(n11513), .B(n11512), .Z(n11514) );
  XNOR U12901 ( .A(n11515), .B(n11514), .Z(n11818) );
  NAND U12902 ( .A(n11819), .B(n11818), .Z(n11516) );
  NAND U12903 ( .A(n11517), .B(n11516), .Z(n11821) );
  NAND U12904 ( .A(a[21]), .B(b[32]), .Z(n11823) );
  AND U12905 ( .A(a[22]), .B(b[32]), .Z(n11523) );
  NANDN U12906 ( .A(n11522), .B(n11523), .Z(n11525) );
  XNOR U12907 ( .A(n11519), .B(n11518), .Z(n11520) );
  XNOR U12908 ( .A(n11521), .B(n11520), .Z(n11705) );
  XNOR U12909 ( .A(n11523), .B(n11522), .Z(n11704) );
  NAND U12910 ( .A(n11705), .B(n11704), .Z(n11524) );
  NAND U12911 ( .A(n11525), .B(n11524), .Z(n11829) );
  NAND U12912 ( .A(a[23]), .B(b[32]), .Z(n11831) );
  AND U12913 ( .A(a[24]), .B(b[32]), .Z(n11531) );
  NANDN U12914 ( .A(n11530), .B(n11531), .Z(n11533) );
  XNOR U12915 ( .A(n11527), .B(n11526), .Z(n11528) );
  XNOR U12916 ( .A(n11529), .B(n11528), .Z(n11703) );
  XNOR U12917 ( .A(n11531), .B(n11530), .Z(n11702) );
  NAND U12918 ( .A(n11703), .B(n11702), .Z(n11532) );
  NAND U12919 ( .A(n11533), .B(n11532), .Z(n11840) );
  AND U12920 ( .A(a[25]), .B(b[32]), .Z(n11838) );
  AND U12921 ( .A(a[26]), .B(b[32]), .Z(n11539) );
  NANDN U12922 ( .A(n11538), .B(n11539), .Z(n11541) );
  XNOR U12923 ( .A(n11535), .B(n11534), .Z(n11536) );
  XNOR U12924 ( .A(n11537), .B(n11536), .Z(n11844) );
  XNOR U12925 ( .A(n11539), .B(n11538), .Z(n11843) );
  NAND U12926 ( .A(n11844), .B(n11843), .Z(n11540) );
  NAND U12927 ( .A(n11541), .B(n11540), .Z(n11846) );
  NANDN U12928 ( .A(n11542), .B(n11543), .Z(n11547) );
  NAND U12929 ( .A(n11853), .B(n11852), .Z(n11546) );
  NAND U12930 ( .A(n11547), .B(n11546), .Z(n11855) );
  NAND U12931 ( .A(a[29]), .B(b[32]), .Z(n11857) );
  AND U12932 ( .A(a[30]), .B(b[32]), .Z(n11549) );
  NANDN U12933 ( .A(n11548), .B(n11549), .Z(n11553) );
  XNOR U12934 ( .A(n11549), .B(n11548), .Z(n11701) );
  NAND U12935 ( .A(n11701), .B(n11700), .Z(n11552) );
  NAND U12936 ( .A(n11553), .B(n11552), .Z(n11863) );
  NAND U12937 ( .A(a[31]), .B(b[32]), .Z(n11865) );
  AND U12938 ( .A(a[32]), .B(b[32]), .Z(n11554) );
  NANDN U12939 ( .A(n11555), .B(n11554), .Z(n11559) );
  XOR U12940 ( .A(n11555), .B(n11554), .Z(n11870) );
  NANDN U12941 ( .A(n11870), .B(n11871), .Z(n11558) );
  AND U12942 ( .A(n11559), .B(n11558), .Z(n11560) );
  NANDN U12943 ( .A(n11561), .B(n11560), .Z(n11567) );
  XOR U12944 ( .A(n11561), .B(n11560), .Z(n11698) );
  XOR U12945 ( .A(n11563), .B(n11562), .Z(n11564) );
  XOR U12946 ( .A(n11565), .B(n11564), .Z(n11699) );
  OR U12947 ( .A(n11698), .B(n11699), .Z(n11566) );
  NAND U12948 ( .A(n11567), .B(n11566), .Z(n11876) );
  XNOR U12949 ( .A(n11569), .B(n11568), .Z(n11877) );
  NANDN U12950 ( .A(n11876), .B(n11877), .Z(n11570) );
  AND U12951 ( .A(n11571), .B(n11570), .Z(n11575) );
  XNOR U12952 ( .A(n11573), .B(n11572), .Z(n11574) );
  NANDN U12953 ( .A(n11575), .B(n11574), .Z(n11577) );
  NAND U12954 ( .A(a[35]), .B(b[32]), .Z(n11884) );
  XNOR U12955 ( .A(n11575), .B(n11574), .Z(n11885) );
  NANDN U12956 ( .A(n11884), .B(n11885), .Z(n11576) );
  AND U12957 ( .A(n11577), .B(n11576), .Z(n11891) );
  OR U12958 ( .A(n11890), .B(n11891), .Z(n11578) );
  NAND U12959 ( .A(n11579), .B(n11578), .Z(n11584) );
  XOR U12960 ( .A(n11581), .B(n11580), .Z(n11582) );
  XNOR U12961 ( .A(n11583), .B(n11582), .Z(n11585) );
  NANDN U12962 ( .A(n11584), .B(n11585), .Z(n11587) );
  XOR U12963 ( .A(n11585), .B(n11584), .Z(n11894) );
  AND U12964 ( .A(a[37]), .B(b[32]), .Z(n11895) );
  OR U12965 ( .A(n11894), .B(n11895), .Z(n11586) );
  AND U12966 ( .A(n11587), .B(n11586), .Z(n11901) );
  NANDN U12967 ( .A(n11900), .B(n11901), .Z(n11588) );
  NAND U12968 ( .A(n11589), .B(n11588), .Z(n11590) );
  NANDN U12969 ( .A(n11591), .B(n11590), .Z(n11593) );
  NAND U12970 ( .A(a[39]), .B(b[32]), .Z(n11908) );
  XNOR U12971 ( .A(n11591), .B(n11590), .Z(n11909) );
  NANDN U12972 ( .A(n11908), .B(n11909), .Z(n11592) );
  AND U12973 ( .A(n11593), .B(n11592), .Z(n11913) );
  XNOR U12974 ( .A(n11595), .B(n11594), .Z(n11912) );
  NANDN U12975 ( .A(n11913), .B(n11912), .Z(n11596) );
  NAND U12976 ( .A(n11597), .B(n11596), .Z(n11598) );
  NANDN U12977 ( .A(n11599), .B(n11598), .Z(n11601) );
  NAND U12978 ( .A(a[41]), .B(b[32]), .Z(n11920) );
  XNOR U12979 ( .A(n11599), .B(n11598), .Z(n11921) );
  NANDN U12980 ( .A(n11920), .B(n11921), .Z(n11600) );
  AND U12981 ( .A(n11601), .B(n11600), .Z(n11925) );
  XNOR U12982 ( .A(n11603), .B(n11602), .Z(n11924) );
  NANDN U12983 ( .A(n11925), .B(n11924), .Z(n11604) );
  AND U12984 ( .A(n11605), .B(n11604), .Z(n11609) );
  XNOR U12985 ( .A(n11607), .B(n11606), .Z(n11608) );
  NANDN U12986 ( .A(n11609), .B(n11608), .Z(n11611) );
  NAND U12987 ( .A(a[43]), .B(b[32]), .Z(n11932) );
  XNOR U12988 ( .A(n11609), .B(n11608), .Z(n11933) );
  NANDN U12989 ( .A(n11932), .B(n11933), .Z(n11610) );
  AND U12990 ( .A(n11611), .B(n11610), .Z(n11939) );
  OR U12991 ( .A(n11938), .B(n11939), .Z(n11612) );
  AND U12992 ( .A(n11613), .B(n11612), .Z(n11617) );
  XNOR U12993 ( .A(n11615), .B(n11614), .Z(n11616) );
  NANDN U12994 ( .A(n11617), .B(n11616), .Z(n11619) );
  NAND U12995 ( .A(a[45]), .B(b[32]), .Z(n11944) );
  XNOR U12996 ( .A(n11617), .B(n11616), .Z(n11945) );
  NANDN U12997 ( .A(n11944), .B(n11945), .Z(n11618) );
  AND U12998 ( .A(n11619), .B(n11618), .Z(n11949) );
  XNOR U12999 ( .A(n11621), .B(n11620), .Z(n11948) );
  NANDN U13000 ( .A(n11949), .B(n11948), .Z(n11622) );
  AND U13001 ( .A(n11623), .B(n11622), .Z(n11627) );
  XNOR U13002 ( .A(n11625), .B(n11624), .Z(n11626) );
  NANDN U13003 ( .A(n11627), .B(n11626), .Z(n11629) );
  NAND U13004 ( .A(a[47]), .B(b[32]), .Z(n11956) );
  XNOR U13005 ( .A(n11627), .B(n11626), .Z(n11957) );
  NANDN U13006 ( .A(n11956), .B(n11957), .Z(n11628) );
  AND U13007 ( .A(n11629), .B(n11628), .Z(n11963) );
  OR U13008 ( .A(n11962), .B(n11963), .Z(n11630) );
  AND U13009 ( .A(n11631), .B(n11630), .Z(n11635) );
  XNOR U13010 ( .A(n11633), .B(n11632), .Z(n11634) );
  NANDN U13011 ( .A(n11635), .B(n11634), .Z(n11637) );
  NAND U13012 ( .A(a[49]), .B(b[32]), .Z(n11968) );
  XNOR U13013 ( .A(n11635), .B(n11634), .Z(n11969) );
  NANDN U13014 ( .A(n11968), .B(n11969), .Z(n11636) );
  AND U13015 ( .A(n11637), .B(n11636), .Z(n11975) );
  OR U13016 ( .A(n11974), .B(n11975), .Z(n11638) );
  AND U13017 ( .A(n11639), .B(n11638), .Z(n11643) );
  XNOR U13018 ( .A(n11641), .B(n11640), .Z(n11642) );
  NANDN U13019 ( .A(n11643), .B(n11642), .Z(n11645) );
  NAND U13020 ( .A(a[51]), .B(b[32]), .Z(n11980) );
  XNOR U13021 ( .A(n11643), .B(n11642), .Z(n11981) );
  NANDN U13022 ( .A(n11980), .B(n11981), .Z(n11644) );
  AND U13023 ( .A(n11645), .B(n11644), .Z(n11987) );
  OR U13024 ( .A(n11986), .B(n11987), .Z(n11646) );
  NAND U13025 ( .A(n11647), .B(n11646), .Z(n11648) );
  NANDN U13026 ( .A(n11649), .B(n11648), .Z(n11651) );
  NAND U13027 ( .A(a[53]), .B(b[32]), .Z(n11992) );
  XNOR U13028 ( .A(n11649), .B(n11648), .Z(n11993) );
  NANDN U13029 ( .A(n11992), .B(n11993), .Z(n11650) );
  AND U13030 ( .A(n11651), .B(n11650), .Z(n11999) );
  OR U13031 ( .A(n11998), .B(n11999), .Z(n11652) );
  NAND U13032 ( .A(n11653), .B(n11652), .Z(n11654) );
  NANDN U13033 ( .A(n11655), .B(n11654), .Z(n11657) );
  NAND U13034 ( .A(a[55]), .B(b[32]), .Z(n12004) );
  XNOR U13035 ( .A(n11655), .B(n11654), .Z(n12005) );
  NANDN U13036 ( .A(n12004), .B(n12005), .Z(n11656) );
  AND U13037 ( .A(n11657), .B(n11656), .Z(n12011) );
  XNOR U13038 ( .A(n11659), .B(n11658), .Z(n12010) );
  NANDN U13039 ( .A(n12011), .B(n12010), .Z(n11660) );
  AND U13040 ( .A(n11661), .B(n11660), .Z(n11665) );
  XNOR U13041 ( .A(n11663), .B(n11662), .Z(n11664) );
  NANDN U13042 ( .A(n11665), .B(n11664), .Z(n11667) );
  NAND U13043 ( .A(a[57]), .B(b[32]), .Z(n12016) );
  XNOR U13044 ( .A(n11665), .B(n11664), .Z(n12017) );
  NANDN U13045 ( .A(n12016), .B(n12017), .Z(n11666) );
  AND U13046 ( .A(n11667), .B(n11666), .Z(n12021) );
  XNOR U13047 ( .A(n11669), .B(n11668), .Z(n12020) );
  NANDN U13048 ( .A(n12021), .B(n12020), .Z(n11670) );
  AND U13049 ( .A(n11671), .B(n11670), .Z(n11675) );
  XNOR U13050 ( .A(n11673), .B(n11672), .Z(n11674) );
  NANDN U13051 ( .A(n11675), .B(n11674), .Z(n11677) );
  NAND U13052 ( .A(a[59]), .B(b[32]), .Z(n12028) );
  XNOR U13053 ( .A(n11675), .B(n11674), .Z(n12029) );
  NANDN U13054 ( .A(n12028), .B(n12029), .Z(n11676) );
  AND U13055 ( .A(n11677), .B(n11676), .Z(n12033) );
  XNOR U13056 ( .A(n11679), .B(n11678), .Z(n12032) );
  NANDN U13057 ( .A(n12033), .B(n12032), .Z(n11680) );
  AND U13058 ( .A(n11681), .B(n11680), .Z(n11685) );
  XNOR U13059 ( .A(n11683), .B(n11682), .Z(n11684) );
  NANDN U13060 ( .A(n11685), .B(n11684), .Z(n11687) );
  NAND U13061 ( .A(a[61]), .B(b[32]), .Z(n12040) );
  XNOR U13062 ( .A(n11685), .B(n11684), .Z(n12041) );
  NANDN U13063 ( .A(n12040), .B(n12041), .Z(n11686) );
  AND U13064 ( .A(n11687), .B(n11686), .Z(n12045) );
  XNOR U13065 ( .A(n11689), .B(n11688), .Z(n12044) );
  NANDN U13066 ( .A(n12045), .B(n12044), .Z(n11690) );
  NAND U13067 ( .A(n11691), .B(n11690), .Z(n11692) );
  NANDN U13068 ( .A(n11693), .B(n11692), .Z(n11695) );
  NAND U13069 ( .A(a[63]), .B(b[32]), .Z(n11696) );
  XNOR U13070 ( .A(n11693), .B(n11692), .Z(n11697) );
  NANDN U13071 ( .A(n11696), .B(n11697), .Z(n11694) );
  AND U13072 ( .A(n11695), .B(n11694), .Z(n12051) );
  NOR U13073 ( .A(n12050), .B(n12051), .Z(n24784) );
  XOR U13074 ( .A(n11697), .B(n11696), .Z(n12407) );
  NAND U13075 ( .A(a[56]), .B(b[31]), .Z(n12002) );
  AND U13076 ( .A(a[55]), .B(b[31]), .Z(n11997) );
  NAND U13077 ( .A(a[54]), .B(b[31]), .Z(n11990) );
  AND U13078 ( .A(a[53]), .B(b[31]), .Z(n11985) );
  NAND U13079 ( .A(a[52]), .B(b[31]), .Z(n11978) );
  AND U13080 ( .A(a[51]), .B(b[31]), .Z(n11973) );
  NAND U13081 ( .A(a[50]), .B(b[31]), .Z(n11966) );
  AND U13082 ( .A(a[49]), .B(b[31]), .Z(n11961) );
  NAND U13083 ( .A(a[46]), .B(b[31]), .Z(n11942) );
  AND U13084 ( .A(a[45]), .B(b[31]), .Z(n11937) );
  NAND U13085 ( .A(a[38]), .B(b[31]), .Z(n11896) );
  AND U13086 ( .A(a[37]), .B(b[31]), .Z(n11889) );
  NAND U13087 ( .A(a[35]), .B(b[31]), .Z(n11878) );
  XOR U13088 ( .A(n11699), .B(n11698), .Z(n12287) );
  NAND U13089 ( .A(a[34]), .B(b[31]), .Z(n12288) );
  XNOR U13090 ( .A(n11701), .B(n11700), .Z(n12271) );
  AND U13091 ( .A(a[26]), .B(b[31]), .Z(n11836) );
  XNOR U13092 ( .A(n11703), .B(n11702), .Z(n12247) );
  XNOR U13093 ( .A(n11705), .B(n11704), .Z(n12238) );
  AND U13094 ( .A(a[20]), .B(b[31]), .Z(n11811) );
  XNOR U13095 ( .A(n11707), .B(n11706), .Z(n12219) );
  NAND U13096 ( .A(a[18]), .B(b[31]), .Z(n11807) );
  NAND U13097 ( .A(a[12]), .B(b[31]), .Z(n12122) );
  AND U13098 ( .A(a[4]), .B(b[31]), .Z(n11724) );
  AND U13099 ( .A(a[0]), .B(b[31]), .Z(n12433) );
  AND U13100 ( .A(a[1]), .B(b[32]), .Z(n11711) );
  AND U13101 ( .A(n12433), .B(n11711), .Z(n11708) );
  NAND U13102 ( .A(a[2]), .B(n11708), .Z(n11715) );
  NAND U13103 ( .A(b[32]), .B(a[1]), .Z(n11709) );
  XOR U13104 ( .A(n11710), .B(n11709), .Z(n12136) );
  NAND U13105 ( .A(n11711), .B(a[0]), .Z(n11712) );
  XNOR U13106 ( .A(a[2]), .B(n11712), .Z(n11713) );
  AND U13107 ( .A(b[31]), .B(n11713), .Z(n12137) );
  NANDN U13108 ( .A(n12136), .B(n12137), .Z(n11714) );
  AND U13109 ( .A(n11715), .B(n11714), .Z(n11718) );
  NANDN U13110 ( .A(n11718), .B(n11719), .Z(n11721) );
  NAND U13111 ( .A(a[3]), .B(b[31]), .Z(n12144) );
  NANDN U13112 ( .A(n12144), .B(n12145), .Z(n11720) );
  AND U13113 ( .A(n11721), .B(n11720), .Z(n11725) );
  NANDN U13114 ( .A(n11724), .B(n11725), .Z(n11727) );
  XOR U13115 ( .A(n11723), .B(n11722), .Z(n12126) );
  NANDN U13116 ( .A(n12126), .B(n12127), .Z(n11726) );
  AND U13117 ( .A(n11727), .B(n11726), .Z(n11731) );
  XOR U13118 ( .A(n11729), .B(n11728), .Z(n11730) );
  NAND U13119 ( .A(n11731), .B(n11730), .Z(n11733) );
  AND U13120 ( .A(a[5]), .B(b[31]), .Z(n12153) );
  XOR U13121 ( .A(n11731), .B(n11730), .Z(n12152) );
  NAND U13122 ( .A(n12153), .B(n12152), .Z(n11732) );
  AND U13123 ( .A(n11733), .B(n11732), .Z(n11736) );
  NANDN U13124 ( .A(n11736), .B(n11737), .Z(n11739) );
  NAND U13125 ( .A(a[6]), .B(b[31]), .Z(n12158) );
  NANDN U13126 ( .A(n12158), .B(n12159), .Z(n11738) );
  AND U13127 ( .A(n11739), .B(n11738), .Z(n11742) );
  XOR U13128 ( .A(n11741), .B(n11740), .Z(n11743) );
  NANDN U13129 ( .A(n11742), .B(n11743), .Z(n11745) );
  AND U13130 ( .A(a[7]), .B(b[31]), .Z(n12164) );
  NAND U13131 ( .A(n12165), .B(n12164), .Z(n11744) );
  AND U13132 ( .A(n11745), .B(n11744), .Z(n11746) );
  AND U13133 ( .A(a[8]), .B(b[31]), .Z(n11747) );
  NANDN U13134 ( .A(n11746), .B(n11747), .Z(n11751) );
  NAND U13135 ( .A(n12170), .B(n12171), .Z(n11750) );
  AND U13136 ( .A(n11751), .B(n11750), .Z(n11754) );
  NANDN U13137 ( .A(n11754), .B(n11755), .Z(n11757) );
  AND U13138 ( .A(a[9]), .B(b[31]), .Z(n12177) );
  NAND U13139 ( .A(n12177), .B(n12176), .Z(n11756) );
  AND U13140 ( .A(n11757), .B(n11756), .Z(n11760) );
  AND U13141 ( .A(a[10]), .B(b[31]), .Z(n11761) );
  NANDN U13142 ( .A(n11760), .B(n11761), .Z(n11763) );
  XOR U13143 ( .A(n11759), .B(n11758), .Z(n12183) );
  NAND U13144 ( .A(n12183), .B(n12182), .Z(n11762) );
  AND U13145 ( .A(n11763), .B(n11762), .Z(n11766) );
  XOR U13146 ( .A(n11765), .B(n11764), .Z(n11767) );
  NANDN U13147 ( .A(n11766), .B(n11767), .Z(n11769) );
  NAND U13148 ( .A(a[11]), .B(b[31]), .Z(n12188) );
  NANDN U13149 ( .A(n12188), .B(n12189), .Z(n11768) );
  NAND U13150 ( .A(n11769), .B(n11768), .Z(n12123) );
  NANDN U13151 ( .A(n11776), .B(n11775), .Z(n11778) );
  NAND U13152 ( .A(a[13]), .B(b[31]), .Z(n12194) );
  XNOR U13153 ( .A(n11776), .B(n11775), .Z(n12195) );
  NANDN U13154 ( .A(n12194), .B(n12195), .Z(n11777) );
  AND U13155 ( .A(n11778), .B(n11777), .Z(n11782) );
  AND U13156 ( .A(a[14]), .B(b[31]), .Z(n11783) );
  NANDN U13157 ( .A(n11782), .B(n11783), .Z(n11785) );
  NAND U13158 ( .A(n12201), .B(n12200), .Z(n11784) );
  AND U13159 ( .A(n11785), .B(n11784), .Z(n11788) );
  XOR U13160 ( .A(n11787), .B(n11786), .Z(n11789) );
  NANDN U13161 ( .A(n11788), .B(n11789), .Z(n11791) );
  NAND U13162 ( .A(a[15]), .B(b[31]), .Z(n12208) );
  NANDN U13163 ( .A(n12208), .B(n12209), .Z(n11790) );
  AND U13164 ( .A(n11791), .B(n11790), .Z(n11792) );
  AND U13165 ( .A(a[16]), .B(b[31]), .Z(n11793) );
  NANDN U13166 ( .A(n11792), .B(n11793), .Z(n11799) );
  XNOR U13167 ( .A(n11795), .B(n11794), .Z(n11796) );
  XNOR U13168 ( .A(n11797), .B(n11796), .Z(n12120) );
  NAND U13169 ( .A(n12121), .B(n12120), .Z(n11798) );
  AND U13170 ( .A(n11799), .B(n11798), .Z(n12215) );
  XOR U13171 ( .A(n11801), .B(n11800), .Z(n11802) );
  IV U13172 ( .A(n11802), .Z(n12216) );
  NAND U13173 ( .A(a[17]), .B(b[31]), .Z(n12214) );
  NANDN U13174 ( .A(n11807), .B(n11808), .Z(n11810) );
  XNOR U13175 ( .A(n11804), .B(n11803), .Z(n11805) );
  XNOR U13176 ( .A(n11806), .B(n11805), .Z(n12119) );
  NAND U13177 ( .A(n12119), .B(n12118), .Z(n11809) );
  NAND U13178 ( .A(n11810), .B(n11809), .Z(n12220) );
  NAND U13179 ( .A(a[19]), .B(b[31]), .Z(n12222) );
  NANDN U13180 ( .A(n11811), .B(n11812), .Z(n11817) );
  NAND U13181 ( .A(n12227), .B(n12228), .Z(n11816) );
  NAND U13182 ( .A(n11817), .B(n11816), .Z(n12233) );
  XOR U13183 ( .A(n11819), .B(n11818), .Z(n12232) );
  AND U13184 ( .A(a[21]), .B(b[31]), .Z(n12231) );
  AND U13185 ( .A(a[22]), .B(b[31]), .Z(n11824) );
  NANDN U13186 ( .A(n11825), .B(n11824), .Z(n11827) );
  XNOR U13187 ( .A(n11821), .B(n11820), .Z(n11822) );
  XNOR U13188 ( .A(n11823), .B(n11822), .Z(n12117) );
  XNOR U13189 ( .A(n11825), .B(n11824), .Z(n12116) );
  NAND U13190 ( .A(n12117), .B(n12116), .Z(n11826) );
  NAND U13191 ( .A(n11827), .B(n11826), .Z(n12239) );
  NAND U13192 ( .A(a[23]), .B(b[31]), .Z(n12241) );
  AND U13193 ( .A(a[24]), .B(b[31]), .Z(n11832) );
  NANDN U13194 ( .A(n11833), .B(n11832), .Z(n11835) );
  XNOR U13195 ( .A(n11829), .B(n11828), .Z(n11830) );
  XNOR U13196 ( .A(n11831), .B(n11830), .Z(n12115) );
  XNOR U13197 ( .A(n11833), .B(n11832), .Z(n12114) );
  NAND U13198 ( .A(n12115), .B(n12114), .Z(n11834) );
  NAND U13199 ( .A(n11835), .B(n11834), .Z(n12248) );
  AND U13200 ( .A(a[25]), .B(b[31]), .Z(n12246) );
  NANDN U13201 ( .A(n11836), .B(n11837), .Z(n11842) );
  NAND U13202 ( .A(n12251), .B(n12252), .Z(n11841) );
  NAND U13203 ( .A(n11842), .B(n11841), .Z(n12256) );
  XOR U13204 ( .A(n11844), .B(n11843), .Z(n12255) );
  AND U13205 ( .A(a[27]), .B(b[31]), .Z(n12254) );
  AND U13206 ( .A(a[28]), .B(b[31]), .Z(n11848) );
  NANDN U13207 ( .A(n11849), .B(n11848), .Z(n11851) );
  XNOR U13208 ( .A(n11849), .B(n11848), .Z(n12112) );
  NAND U13209 ( .A(n12113), .B(n12112), .Z(n11850) );
  AND U13210 ( .A(n11851), .B(n11850), .Z(n12261) );
  XOR U13211 ( .A(n11853), .B(n11852), .Z(n12262) );
  NAND U13212 ( .A(a[29]), .B(b[31]), .Z(n12263) );
  AND U13213 ( .A(a[30]), .B(b[31]), .Z(n11858) );
  NANDN U13214 ( .A(n11859), .B(n11858), .Z(n11861) );
  XNOR U13215 ( .A(n11855), .B(n11854), .Z(n11856) );
  XOR U13216 ( .A(n11857), .B(n11856), .Z(n12268) );
  XNOR U13217 ( .A(n11859), .B(n11858), .Z(n12269) );
  NANDN U13218 ( .A(n12268), .B(n12269), .Z(n11860) );
  NAND U13219 ( .A(n11861), .B(n11860), .Z(n12272) );
  NAND U13220 ( .A(a[31]), .B(b[31]), .Z(n12274) );
  AND U13221 ( .A(a[32]), .B(b[31]), .Z(n11866) );
  NANDN U13222 ( .A(n11867), .B(n11866), .Z(n11869) );
  XNOR U13223 ( .A(n11863), .B(n11862), .Z(n11864) );
  XNOR U13224 ( .A(n11865), .B(n11864), .Z(n12111) );
  XNOR U13225 ( .A(n11867), .B(n11866), .Z(n12110) );
  NAND U13226 ( .A(n12111), .B(n12110), .Z(n11868) );
  AND U13227 ( .A(n11869), .B(n11868), .Z(n11873) );
  NAND U13228 ( .A(n11873), .B(n11872), .Z(n11875) );
  XOR U13229 ( .A(n11873), .B(n11872), .Z(n12282) );
  NAND U13230 ( .A(a[33]), .B(b[31]), .Z(n12281) );
  NAND U13231 ( .A(n12282), .B(n12281), .Z(n11874) );
  NAND U13232 ( .A(n11875), .B(n11874), .Z(n12290) );
  NANDN U13233 ( .A(n11878), .B(n11879), .Z(n11881) );
  XOR U13234 ( .A(n11877), .B(n11876), .Z(n12108) );
  XNOR U13235 ( .A(n11879), .B(n11878), .Z(n12109) );
  NANDN U13236 ( .A(n12108), .B(n12109), .Z(n11880) );
  AND U13237 ( .A(n11881), .B(n11880), .Z(n11883) );
  AND U13238 ( .A(a[36]), .B(b[31]), .Z(n11882) );
  NANDN U13239 ( .A(n11883), .B(n11882), .Z(n11887) );
  XOR U13240 ( .A(n11883), .B(n11882), .Z(n12297) );
  XNOR U13241 ( .A(n11885), .B(n11884), .Z(n12298) );
  NANDN U13242 ( .A(n12297), .B(n12298), .Z(n11886) );
  AND U13243 ( .A(n11887), .B(n11886), .Z(n11888) );
  NANDN U13244 ( .A(n11889), .B(n11888), .Z(n11893) );
  XOR U13245 ( .A(n11889), .B(n11888), .Z(n12104) );
  XOR U13246 ( .A(n11891), .B(n11890), .Z(n12105) );
  OR U13247 ( .A(n12104), .B(n12105), .Z(n11892) );
  AND U13248 ( .A(n11893), .B(n11892), .Z(n11897) );
  NANDN U13249 ( .A(n11896), .B(n11897), .Z(n11899) );
  XOR U13250 ( .A(n11895), .B(n11894), .Z(n12306) );
  XNOR U13251 ( .A(n11897), .B(n11896), .Z(n12305) );
  NANDN U13252 ( .A(n12306), .B(n12305), .Z(n11898) );
  AND U13253 ( .A(n11899), .B(n11898), .Z(n11903) );
  AND U13254 ( .A(a[39]), .B(b[31]), .Z(n11902) );
  NANDN U13255 ( .A(n11903), .B(n11902), .Z(n11905) );
  XOR U13256 ( .A(n11901), .B(n11900), .Z(n12100) );
  XNOR U13257 ( .A(n11903), .B(n11902), .Z(n12101) );
  NANDN U13258 ( .A(n12100), .B(n12101), .Z(n11904) );
  AND U13259 ( .A(n11905), .B(n11904), .Z(n11907) );
  AND U13260 ( .A(a[40]), .B(b[31]), .Z(n11906) );
  NANDN U13261 ( .A(n11907), .B(n11906), .Z(n11911) );
  XOR U13262 ( .A(n11907), .B(n11906), .Z(n12313) );
  XNOR U13263 ( .A(n11909), .B(n11908), .Z(n12314) );
  NANDN U13264 ( .A(n12313), .B(n12314), .Z(n11910) );
  AND U13265 ( .A(n11911), .B(n11910), .Z(n11915) );
  AND U13266 ( .A(a[41]), .B(b[31]), .Z(n11914) );
  NANDN U13267 ( .A(n11915), .B(n11914), .Z(n11917) );
  XOR U13268 ( .A(n11913), .B(n11912), .Z(n12096) );
  XNOR U13269 ( .A(n11915), .B(n11914), .Z(n12097) );
  NANDN U13270 ( .A(n12096), .B(n12097), .Z(n11916) );
  AND U13271 ( .A(n11917), .B(n11916), .Z(n11919) );
  AND U13272 ( .A(a[42]), .B(b[31]), .Z(n11918) );
  NANDN U13273 ( .A(n11919), .B(n11918), .Z(n11923) );
  XOR U13274 ( .A(n11919), .B(n11918), .Z(n12321) );
  XNOR U13275 ( .A(n11921), .B(n11920), .Z(n12322) );
  NANDN U13276 ( .A(n12321), .B(n12322), .Z(n11922) );
  AND U13277 ( .A(n11923), .B(n11922), .Z(n11927) );
  AND U13278 ( .A(a[43]), .B(b[31]), .Z(n11926) );
  NANDN U13279 ( .A(n11927), .B(n11926), .Z(n11929) );
  XOR U13280 ( .A(n11925), .B(n11924), .Z(n12092) );
  XNOR U13281 ( .A(n11927), .B(n11926), .Z(n12093) );
  NANDN U13282 ( .A(n12092), .B(n12093), .Z(n11928) );
  AND U13283 ( .A(n11929), .B(n11928), .Z(n11931) );
  AND U13284 ( .A(a[44]), .B(b[31]), .Z(n11930) );
  NANDN U13285 ( .A(n11931), .B(n11930), .Z(n11935) );
  XOR U13286 ( .A(n11931), .B(n11930), .Z(n12329) );
  XNOR U13287 ( .A(n11933), .B(n11932), .Z(n12330) );
  NANDN U13288 ( .A(n12329), .B(n12330), .Z(n11934) );
  AND U13289 ( .A(n11935), .B(n11934), .Z(n11936) );
  NANDN U13290 ( .A(n11937), .B(n11936), .Z(n11941) );
  XOR U13291 ( .A(n11937), .B(n11936), .Z(n12088) );
  XOR U13292 ( .A(n11939), .B(n11938), .Z(n12089) );
  OR U13293 ( .A(n12088), .B(n12089), .Z(n11940) );
  AND U13294 ( .A(n11941), .B(n11940), .Z(n11943) );
  NANDN U13295 ( .A(n11942), .B(n11943), .Z(n11947) );
  XOR U13296 ( .A(n11943), .B(n11942), .Z(n12337) );
  XNOR U13297 ( .A(n11945), .B(n11944), .Z(n12338) );
  NANDN U13298 ( .A(n12337), .B(n12338), .Z(n11946) );
  AND U13299 ( .A(n11947), .B(n11946), .Z(n11951) );
  AND U13300 ( .A(a[47]), .B(b[31]), .Z(n11950) );
  NANDN U13301 ( .A(n11951), .B(n11950), .Z(n11953) );
  XOR U13302 ( .A(n11949), .B(n11948), .Z(n12084) );
  XNOR U13303 ( .A(n11951), .B(n11950), .Z(n12085) );
  NANDN U13304 ( .A(n12084), .B(n12085), .Z(n11952) );
  AND U13305 ( .A(n11953), .B(n11952), .Z(n11955) );
  AND U13306 ( .A(a[48]), .B(b[31]), .Z(n11954) );
  NANDN U13307 ( .A(n11955), .B(n11954), .Z(n11959) );
  XOR U13308 ( .A(n11955), .B(n11954), .Z(n12345) );
  XNOR U13309 ( .A(n11957), .B(n11956), .Z(n12346) );
  NANDN U13310 ( .A(n12345), .B(n12346), .Z(n11958) );
  AND U13311 ( .A(n11959), .B(n11958), .Z(n11960) );
  NANDN U13312 ( .A(n11961), .B(n11960), .Z(n11965) );
  XOR U13313 ( .A(n11961), .B(n11960), .Z(n12080) );
  XOR U13314 ( .A(n11963), .B(n11962), .Z(n12081) );
  OR U13315 ( .A(n12080), .B(n12081), .Z(n11964) );
  AND U13316 ( .A(n11965), .B(n11964), .Z(n11967) );
  NANDN U13317 ( .A(n11966), .B(n11967), .Z(n11971) );
  XOR U13318 ( .A(n11967), .B(n11966), .Z(n12353) );
  XNOR U13319 ( .A(n11969), .B(n11968), .Z(n12354) );
  NANDN U13320 ( .A(n12353), .B(n12354), .Z(n11970) );
  AND U13321 ( .A(n11971), .B(n11970), .Z(n11972) );
  NANDN U13322 ( .A(n11973), .B(n11972), .Z(n11977) );
  XOR U13323 ( .A(n11973), .B(n11972), .Z(n12076) );
  XOR U13324 ( .A(n11975), .B(n11974), .Z(n12077) );
  OR U13325 ( .A(n12076), .B(n12077), .Z(n11976) );
  AND U13326 ( .A(n11977), .B(n11976), .Z(n11979) );
  NANDN U13327 ( .A(n11978), .B(n11979), .Z(n11983) );
  XOR U13328 ( .A(n11979), .B(n11978), .Z(n12361) );
  XNOR U13329 ( .A(n11981), .B(n11980), .Z(n12362) );
  NANDN U13330 ( .A(n12361), .B(n12362), .Z(n11982) );
  AND U13331 ( .A(n11983), .B(n11982), .Z(n11984) );
  NANDN U13332 ( .A(n11985), .B(n11984), .Z(n11989) );
  XOR U13333 ( .A(n11985), .B(n11984), .Z(n12072) );
  XOR U13334 ( .A(n11987), .B(n11986), .Z(n12073) );
  OR U13335 ( .A(n12072), .B(n12073), .Z(n11988) );
  AND U13336 ( .A(n11989), .B(n11988), .Z(n11991) );
  NANDN U13337 ( .A(n11990), .B(n11991), .Z(n11995) );
  XOR U13338 ( .A(n11991), .B(n11990), .Z(n12369) );
  XNOR U13339 ( .A(n11993), .B(n11992), .Z(n12370) );
  NANDN U13340 ( .A(n12369), .B(n12370), .Z(n11994) );
  AND U13341 ( .A(n11995), .B(n11994), .Z(n11996) );
  NANDN U13342 ( .A(n11997), .B(n11996), .Z(n12001) );
  XOR U13343 ( .A(n11997), .B(n11996), .Z(n12068) );
  XOR U13344 ( .A(n11999), .B(n11998), .Z(n12069) );
  OR U13345 ( .A(n12068), .B(n12069), .Z(n12000) );
  AND U13346 ( .A(n12001), .B(n12000), .Z(n12003) );
  NANDN U13347 ( .A(n12002), .B(n12003), .Z(n12007) );
  XOR U13348 ( .A(n12003), .B(n12002), .Z(n12377) );
  XNOR U13349 ( .A(n12005), .B(n12004), .Z(n12378) );
  NANDN U13350 ( .A(n12377), .B(n12378), .Z(n12006) );
  AND U13351 ( .A(n12007), .B(n12006), .Z(n12009) );
  AND U13352 ( .A(a[57]), .B(b[31]), .Z(n12008) );
  NANDN U13353 ( .A(n12009), .B(n12008), .Z(n12013) );
  XOR U13354 ( .A(n12009), .B(n12008), .Z(n12064) );
  XNOR U13355 ( .A(n12011), .B(n12010), .Z(n12065) );
  NANDN U13356 ( .A(n12064), .B(n12065), .Z(n12012) );
  AND U13357 ( .A(n12013), .B(n12012), .Z(n12015) );
  AND U13358 ( .A(a[58]), .B(b[31]), .Z(n12014) );
  NANDN U13359 ( .A(n12015), .B(n12014), .Z(n12019) );
  XOR U13360 ( .A(n12015), .B(n12014), .Z(n12385) );
  XNOR U13361 ( .A(n12017), .B(n12016), .Z(n12386) );
  NANDN U13362 ( .A(n12385), .B(n12386), .Z(n12018) );
  AND U13363 ( .A(n12019), .B(n12018), .Z(n12023) );
  AND U13364 ( .A(a[59]), .B(b[31]), .Z(n12022) );
  NANDN U13365 ( .A(n12023), .B(n12022), .Z(n12025) );
  XOR U13366 ( .A(n12021), .B(n12020), .Z(n12060) );
  XNOR U13367 ( .A(n12023), .B(n12022), .Z(n12061) );
  NANDN U13368 ( .A(n12060), .B(n12061), .Z(n12024) );
  AND U13369 ( .A(n12025), .B(n12024), .Z(n12027) );
  AND U13370 ( .A(a[60]), .B(b[31]), .Z(n12026) );
  NANDN U13371 ( .A(n12027), .B(n12026), .Z(n12031) );
  XOR U13372 ( .A(n12027), .B(n12026), .Z(n12393) );
  XNOR U13373 ( .A(n12029), .B(n12028), .Z(n12394) );
  NANDN U13374 ( .A(n12393), .B(n12394), .Z(n12030) );
  AND U13375 ( .A(n12031), .B(n12030), .Z(n12035) );
  AND U13376 ( .A(a[61]), .B(b[31]), .Z(n12034) );
  NANDN U13377 ( .A(n12035), .B(n12034), .Z(n12037) );
  XOR U13378 ( .A(n12033), .B(n12032), .Z(n12056) );
  XNOR U13379 ( .A(n12035), .B(n12034), .Z(n12057) );
  NANDN U13380 ( .A(n12056), .B(n12057), .Z(n12036) );
  AND U13381 ( .A(n12037), .B(n12036), .Z(n12039) );
  AND U13382 ( .A(a[62]), .B(b[31]), .Z(n12038) );
  NANDN U13383 ( .A(n12039), .B(n12038), .Z(n12043) );
  XOR U13384 ( .A(n12039), .B(n12038), .Z(n12401) );
  XNOR U13385 ( .A(n12041), .B(n12040), .Z(n12402) );
  NANDN U13386 ( .A(n12401), .B(n12402), .Z(n12042) );
  AND U13387 ( .A(n12043), .B(n12042), .Z(n12047) );
  AND U13388 ( .A(a[63]), .B(b[31]), .Z(n12046) );
  NANDN U13389 ( .A(n12047), .B(n12046), .Z(n12049) );
  XOR U13390 ( .A(n12045), .B(n12044), .Z(n12054) );
  XNOR U13391 ( .A(n12047), .B(n12046), .Z(n12055) );
  NANDN U13392 ( .A(n12054), .B(n12055), .Z(n12048) );
  AND U13393 ( .A(n12049), .B(n12048), .Z(n12408) );
  NOR U13394 ( .A(n12407), .B(n12408), .Z(n12053) );
  XNOR U13395 ( .A(n12051), .B(n12050), .Z(n12052) );
  NANDN U13396 ( .A(n12053), .B(n12052), .Z(n22545) );
  XNOR U13397 ( .A(n12053), .B(n12052), .Z(n24782) );
  XOR U13398 ( .A(n12055), .B(n12054), .Z(n12756) );
  NAND U13399 ( .A(a[62]), .B(b[30]), .Z(n12058) );
  XNOR U13400 ( .A(n12057), .B(n12056), .Z(n12059) );
  NANDN U13401 ( .A(n12058), .B(n12059), .Z(n12400) );
  XOR U13402 ( .A(n12059), .B(n12058), .Z(n12750) );
  NAND U13403 ( .A(a[60]), .B(b[30]), .Z(n12062) );
  XNOR U13404 ( .A(n12061), .B(n12060), .Z(n12063) );
  NANDN U13405 ( .A(n12062), .B(n12063), .Z(n12392) );
  XOR U13406 ( .A(n12063), .B(n12062), .Z(n12738) );
  NAND U13407 ( .A(a[58]), .B(b[30]), .Z(n12066) );
  XNOR U13408 ( .A(n12065), .B(n12064), .Z(n12067) );
  NANDN U13409 ( .A(n12066), .B(n12067), .Z(n12384) );
  XOR U13410 ( .A(n12067), .B(n12066), .Z(n12726) );
  XOR U13411 ( .A(n12069), .B(n12068), .Z(n12071) );
  AND U13412 ( .A(a[56]), .B(b[30]), .Z(n12070) );
  NANDN U13413 ( .A(n12071), .B(n12070), .Z(n12376) );
  XOR U13414 ( .A(n12071), .B(n12070), .Z(n12714) );
  XOR U13415 ( .A(n12073), .B(n12072), .Z(n12075) );
  AND U13416 ( .A(a[54]), .B(b[30]), .Z(n12074) );
  NANDN U13417 ( .A(n12075), .B(n12074), .Z(n12368) );
  XOR U13418 ( .A(n12075), .B(n12074), .Z(n12702) );
  XOR U13419 ( .A(n12077), .B(n12076), .Z(n12079) );
  AND U13420 ( .A(a[52]), .B(b[30]), .Z(n12078) );
  NANDN U13421 ( .A(n12079), .B(n12078), .Z(n12360) );
  XOR U13422 ( .A(n12079), .B(n12078), .Z(n12690) );
  XOR U13423 ( .A(n12081), .B(n12080), .Z(n12083) );
  AND U13424 ( .A(a[50]), .B(b[30]), .Z(n12082) );
  NANDN U13425 ( .A(n12083), .B(n12082), .Z(n12352) );
  XOR U13426 ( .A(n12083), .B(n12082), .Z(n12678) );
  NAND U13427 ( .A(a[48]), .B(b[30]), .Z(n12086) );
  XNOR U13428 ( .A(n12085), .B(n12084), .Z(n12087) );
  NANDN U13429 ( .A(n12086), .B(n12087), .Z(n12344) );
  XOR U13430 ( .A(n12087), .B(n12086), .Z(n12666) );
  XOR U13431 ( .A(n12089), .B(n12088), .Z(n12091) );
  AND U13432 ( .A(a[46]), .B(b[30]), .Z(n12090) );
  NANDN U13433 ( .A(n12091), .B(n12090), .Z(n12336) );
  XOR U13434 ( .A(n12091), .B(n12090), .Z(n12654) );
  NAND U13435 ( .A(a[44]), .B(b[30]), .Z(n12094) );
  XNOR U13436 ( .A(n12093), .B(n12092), .Z(n12095) );
  NANDN U13437 ( .A(n12094), .B(n12095), .Z(n12328) );
  XOR U13438 ( .A(n12095), .B(n12094), .Z(n12642) );
  NAND U13439 ( .A(a[42]), .B(b[30]), .Z(n12098) );
  XNOR U13440 ( .A(n12097), .B(n12096), .Z(n12099) );
  NANDN U13441 ( .A(n12098), .B(n12099), .Z(n12320) );
  XOR U13442 ( .A(n12099), .B(n12098), .Z(n12630) );
  NAND U13443 ( .A(a[40]), .B(b[30]), .Z(n12102) );
  XNOR U13444 ( .A(n12101), .B(n12100), .Z(n12103) );
  NANDN U13445 ( .A(n12102), .B(n12103), .Z(n12312) );
  XOR U13446 ( .A(n12103), .B(n12102), .Z(n12618) );
  XOR U13447 ( .A(n12105), .B(n12104), .Z(n12107) );
  AND U13448 ( .A(a[38]), .B(b[30]), .Z(n12106) );
  NANDN U13449 ( .A(n12107), .B(n12106), .Z(n12304) );
  XOR U13450 ( .A(n12107), .B(n12106), .Z(n12606) );
  NAND U13451 ( .A(a[36]), .B(b[30]), .Z(n12293) );
  XNOR U13452 ( .A(n12109), .B(n12108), .Z(n12294) );
  NANDN U13453 ( .A(n12293), .B(n12294), .Z(n12296) );
  XNOR U13454 ( .A(n12111), .B(n12110), .Z(n12582) );
  NAND U13455 ( .A(a[32]), .B(b[30]), .Z(n12275) );
  XNOR U13456 ( .A(n12113), .B(n12112), .Z(n12565) );
  AND U13457 ( .A(a[26]), .B(b[30]), .Z(n12244) );
  XNOR U13458 ( .A(n12115), .B(n12114), .Z(n12547) );
  XNOR U13459 ( .A(n12117), .B(n12116), .Z(n12541) );
  XNOR U13460 ( .A(n12119), .B(n12118), .Z(n12522) );
  XNOR U13461 ( .A(n12121), .B(n12120), .Z(n12518) );
  XNOR U13462 ( .A(n12123), .B(n12122), .Z(n12124) );
  XOR U13463 ( .A(n12125), .B(n12124), .Z(n12500) );
  AND U13464 ( .A(a[8]), .B(b[30]), .Z(n12166) );
  AND U13465 ( .A(b[30]), .B(a[0]), .Z(n12828) );
  AND U13466 ( .A(a[1]), .B(b[31]), .Z(n12131) );
  AND U13467 ( .A(n12828), .B(n12131), .Z(n12128) );
  NAND U13468 ( .A(a[2]), .B(n12128), .Z(n12135) );
  NAND U13469 ( .A(b[31]), .B(a[1]), .Z(n12129) );
  XOR U13470 ( .A(n12130), .B(n12129), .Z(n12439) );
  NAND U13471 ( .A(n12131), .B(a[0]), .Z(n12132) );
  XNOR U13472 ( .A(a[2]), .B(n12132), .Z(n12133) );
  AND U13473 ( .A(b[30]), .B(n12133), .Z(n12440) );
  NANDN U13474 ( .A(n12439), .B(n12440), .Z(n12134) );
  AND U13475 ( .A(n12135), .B(n12134), .Z(n12138) );
  NANDN U13476 ( .A(n12138), .B(n12139), .Z(n12141) );
  AND U13477 ( .A(a[3]), .B(b[30]), .Z(n12445) );
  NAND U13478 ( .A(n12446), .B(n12445), .Z(n12140) );
  AND U13479 ( .A(n12141), .B(n12140), .Z(n12142) );
  AND U13480 ( .A(a[4]), .B(b[30]), .Z(n12143) );
  NANDN U13481 ( .A(n12142), .B(n12143), .Z(n12147) );
  NAND U13482 ( .A(n12452), .B(n12451), .Z(n12146) );
  NAND U13483 ( .A(n12147), .B(n12146), .Z(n12148) );
  NAND U13484 ( .A(n12149), .B(n12148), .Z(n12151) );
  NAND U13485 ( .A(a[5]), .B(b[30]), .Z(n12457) );
  XOR U13486 ( .A(n12149), .B(n12148), .Z(n12458) );
  NANDN U13487 ( .A(n12457), .B(n12458), .Z(n12150) );
  AND U13488 ( .A(n12151), .B(n12150), .Z(n12154) );
  XOR U13489 ( .A(n12153), .B(n12152), .Z(n12155) );
  NANDN U13490 ( .A(n12154), .B(n12155), .Z(n12157) );
  NAND U13491 ( .A(a[6]), .B(b[30]), .Z(n12463) );
  NANDN U13492 ( .A(n12463), .B(n12464), .Z(n12156) );
  AND U13493 ( .A(n12157), .B(n12156), .Z(n12160) );
  NANDN U13494 ( .A(n12160), .B(n12161), .Z(n12163) );
  NAND U13495 ( .A(a[7]), .B(b[30]), .Z(n12471) );
  NANDN U13496 ( .A(n12471), .B(n12472), .Z(n12162) );
  AND U13497 ( .A(n12163), .B(n12162), .Z(n12167) );
  NANDN U13498 ( .A(n12166), .B(n12167), .Z(n12169) );
  XOR U13499 ( .A(n12165), .B(n12164), .Z(n12429) );
  NANDN U13500 ( .A(n12429), .B(n12430), .Z(n12168) );
  AND U13501 ( .A(n12169), .B(n12168), .Z(n12173) );
  XOR U13502 ( .A(n12171), .B(n12170), .Z(n12172) );
  NAND U13503 ( .A(n12173), .B(n12172), .Z(n12175) );
  AND U13504 ( .A(a[9]), .B(b[30]), .Z(n12480) );
  XOR U13505 ( .A(n12173), .B(n12172), .Z(n12479) );
  NAND U13506 ( .A(n12480), .B(n12479), .Z(n12174) );
  AND U13507 ( .A(n12175), .B(n12174), .Z(n12178) );
  AND U13508 ( .A(a[10]), .B(b[30]), .Z(n12179) );
  NANDN U13509 ( .A(n12178), .B(n12179), .Z(n12181) );
  XOR U13510 ( .A(n12177), .B(n12176), .Z(n12486) );
  NAND U13511 ( .A(n12486), .B(n12485), .Z(n12180) );
  AND U13512 ( .A(n12181), .B(n12180), .Z(n12184) );
  XOR U13513 ( .A(n12183), .B(n12182), .Z(n12185) );
  NANDN U13514 ( .A(n12184), .B(n12185), .Z(n12187) );
  AND U13515 ( .A(a[11]), .B(b[30]), .Z(n12492) );
  NAND U13516 ( .A(n12492), .B(n12491), .Z(n12186) );
  AND U13517 ( .A(n12187), .B(n12186), .Z(n12190) );
  AND U13518 ( .A(a[12]), .B(b[30]), .Z(n12191) );
  NANDN U13519 ( .A(n12190), .B(n12191), .Z(n12193) );
  NAND U13520 ( .A(n12428), .B(n12427), .Z(n12192) );
  NAND U13521 ( .A(n12193), .B(n12192), .Z(n12501) );
  AND U13522 ( .A(a[13]), .B(b[30]), .Z(n12499) );
  AND U13523 ( .A(a[14]), .B(b[30]), .Z(n12197) );
  NANDN U13524 ( .A(n12196), .B(n12197), .Z(n12199) );
  XNOR U13525 ( .A(n12197), .B(n12196), .Z(n12504) );
  NAND U13526 ( .A(n12505), .B(n12504), .Z(n12198) );
  AND U13527 ( .A(n12199), .B(n12198), .Z(n12202) );
  XOR U13528 ( .A(n12201), .B(n12200), .Z(n12203) );
  NANDN U13529 ( .A(n12202), .B(n12203), .Z(n12205) );
  AND U13530 ( .A(a[15]), .B(b[30]), .Z(n12507) );
  NAND U13531 ( .A(n12507), .B(n12506), .Z(n12204) );
  AND U13532 ( .A(n12205), .B(n12204), .Z(n12206) );
  AND U13533 ( .A(a[16]), .B(b[30]), .Z(n12207) );
  NANDN U13534 ( .A(n12206), .B(n12207), .Z(n12211) );
  NAND U13535 ( .A(n12513), .B(n12512), .Z(n12210) );
  NAND U13536 ( .A(n12211), .B(n12210), .Z(n12519) );
  AND U13537 ( .A(a[17]), .B(b[30]), .Z(n12517) );
  AND U13538 ( .A(a[18]), .B(b[30]), .Z(n12213) );
  NANDN U13539 ( .A(n12212), .B(n12213), .Z(n12218) );
  XNOR U13540 ( .A(n12213), .B(n12212), .Z(n12426) );
  NAND U13541 ( .A(n12426), .B(n12425), .Z(n12217) );
  NAND U13542 ( .A(n12218), .B(n12217), .Z(n12523) );
  NAND U13543 ( .A(a[19]), .B(b[30]), .Z(n12525) );
  AND U13544 ( .A(a[20]), .B(b[30]), .Z(n12224) );
  NANDN U13545 ( .A(n12223), .B(n12224), .Z(n12226) );
  XNOR U13546 ( .A(n12220), .B(n12219), .Z(n12221) );
  XOR U13547 ( .A(n12222), .B(n12221), .Z(n12530) );
  XNOR U13548 ( .A(n12224), .B(n12223), .Z(n12531) );
  NANDN U13549 ( .A(n12530), .B(n12531), .Z(n12225) );
  AND U13550 ( .A(n12226), .B(n12225), .Z(n12536) );
  XOR U13551 ( .A(n12228), .B(n12227), .Z(n12535) );
  AND U13552 ( .A(a[21]), .B(b[30]), .Z(n12534) );
  AND U13553 ( .A(a[22]), .B(b[30]), .Z(n12230) );
  NANDN U13554 ( .A(n12229), .B(n12230), .Z(n12235) );
  XNOR U13555 ( .A(n12230), .B(n12229), .Z(n12424) );
  NAND U13556 ( .A(n12424), .B(n12423), .Z(n12234) );
  NAND U13557 ( .A(n12235), .B(n12234), .Z(n12542) );
  NAND U13558 ( .A(a[23]), .B(b[30]), .Z(n12544) );
  AND U13559 ( .A(a[24]), .B(b[30]), .Z(n12237) );
  NANDN U13560 ( .A(n12236), .B(n12237), .Z(n12243) );
  XOR U13561 ( .A(n12237), .B(n12236), .Z(n12421) );
  XNOR U13562 ( .A(n12239), .B(n12238), .Z(n12240) );
  XNOR U13563 ( .A(n12241), .B(n12240), .Z(n12422) );
  NANDN U13564 ( .A(n12421), .B(n12422), .Z(n12242) );
  NAND U13565 ( .A(n12243), .B(n12242), .Z(n12548) );
  NAND U13566 ( .A(a[25]), .B(b[30]), .Z(n12550) );
  NANDN U13567 ( .A(n12244), .B(n12245), .Z(n12250) );
  NAND U13568 ( .A(n12555), .B(n12556), .Z(n12249) );
  AND U13569 ( .A(n12250), .B(n12249), .Z(n12557) );
  XOR U13570 ( .A(n12252), .B(n12251), .Z(n12253) );
  IV U13571 ( .A(n12253), .Z(n12558) );
  NAND U13572 ( .A(a[27]), .B(b[30]), .Z(n12560) );
  AND U13573 ( .A(a[28]), .B(b[30]), .Z(n12258) );
  NANDN U13574 ( .A(n12257), .B(n12258), .Z(n12260) );
  XNOR U13575 ( .A(n12258), .B(n12257), .Z(n12419) );
  NAND U13576 ( .A(n12420), .B(n12419), .Z(n12259) );
  NAND U13577 ( .A(n12260), .B(n12259), .Z(n12566) );
  NAND U13578 ( .A(a[29]), .B(b[30]), .Z(n12568) );
  AND U13579 ( .A(a[30]), .B(b[30]), .Z(n12265) );
  NANDN U13580 ( .A(n12264), .B(n12265), .Z(n12267) );
  XNOR U13581 ( .A(n12265), .B(n12264), .Z(n12418) );
  NANDN U13582 ( .A(n12417), .B(n12418), .Z(n12266) );
  AND U13583 ( .A(n12267), .B(n12266), .Z(n12574) );
  IV U13584 ( .A(n12270), .Z(n12575) );
  NAND U13585 ( .A(a[31]), .B(b[30]), .Z(n12573) );
  NANDN U13586 ( .A(n12275), .B(n12276), .Z(n12278) );
  XNOR U13587 ( .A(n12272), .B(n12271), .Z(n12273) );
  XNOR U13588 ( .A(n12274), .B(n12273), .Z(n12416) );
  NAND U13589 ( .A(n12416), .B(n12415), .Z(n12277) );
  NAND U13590 ( .A(n12278), .B(n12277), .Z(n12583) );
  NAND U13591 ( .A(a[33]), .B(b[30]), .Z(n12585) );
  AND U13592 ( .A(a[34]), .B(b[30]), .Z(n12279) );
  NANDN U13593 ( .A(n12280), .B(n12279), .Z(n12284) );
  XOR U13594 ( .A(n12280), .B(n12279), .Z(n12588) );
  XNOR U13595 ( .A(n12282), .B(n12281), .Z(n12589) );
  NANDN U13596 ( .A(n12588), .B(n12589), .Z(n12283) );
  AND U13597 ( .A(n12284), .B(n12283), .Z(n12286) );
  AND U13598 ( .A(a[35]), .B(b[30]), .Z(n12285) );
  NANDN U13599 ( .A(n12286), .B(n12285), .Z(n12292) );
  XOR U13600 ( .A(n12286), .B(n12285), .Z(n12413) );
  XOR U13601 ( .A(n12288), .B(n12287), .Z(n12289) );
  XNOR U13602 ( .A(n12290), .B(n12289), .Z(n12414) );
  NANDN U13603 ( .A(n12413), .B(n12414), .Z(n12291) );
  AND U13604 ( .A(n12292), .B(n12291), .Z(n12595) );
  XNOR U13605 ( .A(n12294), .B(n12293), .Z(n12594) );
  NANDN U13606 ( .A(n12595), .B(n12594), .Z(n12295) );
  AND U13607 ( .A(n12296), .B(n12295), .Z(n12300) );
  XNOR U13608 ( .A(n12298), .B(n12297), .Z(n12299) );
  NANDN U13609 ( .A(n12300), .B(n12299), .Z(n12302) );
  NAND U13610 ( .A(a[37]), .B(b[30]), .Z(n12600) );
  XNOR U13611 ( .A(n12300), .B(n12299), .Z(n12601) );
  NANDN U13612 ( .A(n12600), .B(n12601), .Z(n12301) );
  AND U13613 ( .A(n12302), .B(n12301), .Z(n12607) );
  OR U13614 ( .A(n12606), .B(n12607), .Z(n12303) );
  AND U13615 ( .A(n12304), .B(n12303), .Z(n12308) );
  XNOR U13616 ( .A(n12306), .B(n12305), .Z(n12307) );
  NANDN U13617 ( .A(n12308), .B(n12307), .Z(n12310) );
  NAND U13618 ( .A(a[39]), .B(b[30]), .Z(n12612) );
  XNOR U13619 ( .A(n12308), .B(n12307), .Z(n12613) );
  NANDN U13620 ( .A(n12612), .B(n12613), .Z(n12309) );
  AND U13621 ( .A(n12310), .B(n12309), .Z(n12619) );
  OR U13622 ( .A(n12618), .B(n12619), .Z(n12311) );
  AND U13623 ( .A(n12312), .B(n12311), .Z(n12316) );
  XNOR U13624 ( .A(n12314), .B(n12313), .Z(n12315) );
  NANDN U13625 ( .A(n12316), .B(n12315), .Z(n12318) );
  NAND U13626 ( .A(a[41]), .B(b[30]), .Z(n12624) );
  XNOR U13627 ( .A(n12316), .B(n12315), .Z(n12625) );
  NANDN U13628 ( .A(n12624), .B(n12625), .Z(n12317) );
  AND U13629 ( .A(n12318), .B(n12317), .Z(n12631) );
  OR U13630 ( .A(n12630), .B(n12631), .Z(n12319) );
  AND U13631 ( .A(n12320), .B(n12319), .Z(n12324) );
  XNOR U13632 ( .A(n12322), .B(n12321), .Z(n12323) );
  NANDN U13633 ( .A(n12324), .B(n12323), .Z(n12326) );
  NAND U13634 ( .A(a[43]), .B(b[30]), .Z(n12636) );
  XNOR U13635 ( .A(n12324), .B(n12323), .Z(n12637) );
  NANDN U13636 ( .A(n12636), .B(n12637), .Z(n12325) );
  AND U13637 ( .A(n12326), .B(n12325), .Z(n12643) );
  OR U13638 ( .A(n12642), .B(n12643), .Z(n12327) );
  AND U13639 ( .A(n12328), .B(n12327), .Z(n12332) );
  XNOR U13640 ( .A(n12330), .B(n12329), .Z(n12331) );
  NANDN U13641 ( .A(n12332), .B(n12331), .Z(n12334) );
  NAND U13642 ( .A(a[45]), .B(b[30]), .Z(n12648) );
  XNOR U13643 ( .A(n12332), .B(n12331), .Z(n12649) );
  NANDN U13644 ( .A(n12648), .B(n12649), .Z(n12333) );
  AND U13645 ( .A(n12334), .B(n12333), .Z(n12655) );
  OR U13646 ( .A(n12654), .B(n12655), .Z(n12335) );
  AND U13647 ( .A(n12336), .B(n12335), .Z(n12340) );
  XNOR U13648 ( .A(n12338), .B(n12337), .Z(n12339) );
  NANDN U13649 ( .A(n12340), .B(n12339), .Z(n12342) );
  NAND U13650 ( .A(a[47]), .B(b[30]), .Z(n12660) );
  XNOR U13651 ( .A(n12340), .B(n12339), .Z(n12661) );
  NANDN U13652 ( .A(n12660), .B(n12661), .Z(n12341) );
  AND U13653 ( .A(n12342), .B(n12341), .Z(n12667) );
  OR U13654 ( .A(n12666), .B(n12667), .Z(n12343) );
  AND U13655 ( .A(n12344), .B(n12343), .Z(n12348) );
  XNOR U13656 ( .A(n12346), .B(n12345), .Z(n12347) );
  NANDN U13657 ( .A(n12348), .B(n12347), .Z(n12350) );
  NAND U13658 ( .A(a[49]), .B(b[30]), .Z(n12672) );
  XNOR U13659 ( .A(n12348), .B(n12347), .Z(n12673) );
  NANDN U13660 ( .A(n12672), .B(n12673), .Z(n12349) );
  AND U13661 ( .A(n12350), .B(n12349), .Z(n12679) );
  OR U13662 ( .A(n12678), .B(n12679), .Z(n12351) );
  AND U13663 ( .A(n12352), .B(n12351), .Z(n12356) );
  XNOR U13664 ( .A(n12354), .B(n12353), .Z(n12355) );
  NANDN U13665 ( .A(n12356), .B(n12355), .Z(n12358) );
  NAND U13666 ( .A(a[51]), .B(b[30]), .Z(n12684) );
  XNOR U13667 ( .A(n12356), .B(n12355), .Z(n12685) );
  NANDN U13668 ( .A(n12684), .B(n12685), .Z(n12357) );
  AND U13669 ( .A(n12358), .B(n12357), .Z(n12691) );
  OR U13670 ( .A(n12690), .B(n12691), .Z(n12359) );
  AND U13671 ( .A(n12360), .B(n12359), .Z(n12364) );
  XNOR U13672 ( .A(n12362), .B(n12361), .Z(n12363) );
  NANDN U13673 ( .A(n12364), .B(n12363), .Z(n12366) );
  NAND U13674 ( .A(a[53]), .B(b[30]), .Z(n12696) );
  XNOR U13675 ( .A(n12364), .B(n12363), .Z(n12697) );
  NANDN U13676 ( .A(n12696), .B(n12697), .Z(n12365) );
  AND U13677 ( .A(n12366), .B(n12365), .Z(n12703) );
  OR U13678 ( .A(n12702), .B(n12703), .Z(n12367) );
  AND U13679 ( .A(n12368), .B(n12367), .Z(n12372) );
  XNOR U13680 ( .A(n12370), .B(n12369), .Z(n12371) );
  NANDN U13681 ( .A(n12372), .B(n12371), .Z(n12374) );
  NAND U13682 ( .A(a[55]), .B(b[30]), .Z(n12708) );
  XNOR U13683 ( .A(n12372), .B(n12371), .Z(n12709) );
  NANDN U13684 ( .A(n12708), .B(n12709), .Z(n12373) );
  AND U13685 ( .A(n12374), .B(n12373), .Z(n12715) );
  OR U13686 ( .A(n12714), .B(n12715), .Z(n12375) );
  AND U13687 ( .A(n12376), .B(n12375), .Z(n12380) );
  XNOR U13688 ( .A(n12378), .B(n12377), .Z(n12379) );
  NANDN U13689 ( .A(n12380), .B(n12379), .Z(n12382) );
  NAND U13690 ( .A(a[57]), .B(b[30]), .Z(n12720) );
  XNOR U13691 ( .A(n12380), .B(n12379), .Z(n12721) );
  NANDN U13692 ( .A(n12720), .B(n12721), .Z(n12381) );
  AND U13693 ( .A(n12382), .B(n12381), .Z(n12727) );
  OR U13694 ( .A(n12726), .B(n12727), .Z(n12383) );
  AND U13695 ( .A(n12384), .B(n12383), .Z(n12388) );
  XNOR U13696 ( .A(n12386), .B(n12385), .Z(n12387) );
  NANDN U13697 ( .A(n12388), .B(n12387), .Z(n12390) );
  NAND U13698 ( .A(a[59]), .B(b[30]), .Z(n12734) );
  XNOR U13699 ( .A(n12388), .B(n12387), .Z(n12735) );
  NANDN U13700 ( .A(n12734), .B(n12735), .Z(n12389) );
  AND U13701 ( .A(n12390), .B(n12389), .Z(n12739) );
  OR U13702 ( .A(n12738), .B(n12739), .Z(n12391) );
  AND U13703 ( .A(n12392), .B(n12391), .Z(n12396) );
  XNOR U13704 ( .A(n12394), .B(n12393), .Z(n12395) );
  NANDN U13705 ( .A(n12396), .B(n12395), .Z(n12398) );
  NAND U13706 ( .A(a[61]), .B(b[30]), .Z(n12744) );
  XNOR U13707 ( .A(n12396), .B(n12395), .Z(n12745) );
  NANDN U13708 ( .A(n12744), .B(n12745), .Z(n12397) );
  AND U13709 ( .A(n12398), .B(n12397), .Z(n12751) );
  OR U13710 ( .A(n12750), .B(n12751), .Z(n12399) );
  AND U13711 ( .A(n12400), .B(n12399), .Z(n12404) );
  XNOR U13712 ( .A(n12402), .B(n12401), .Z(n12403) );
  NANDN U13713 ( .A(n12404), .B(n12403), .Z(n12406) );
  NAND U13714 ( .A(a[63]), .B(b[30]), .Z(n12411) );
  XNOR U13715 ( .A(n12404), .B(n12403), .Z(n12412) );
  NANDN U13716 ( .A(n12411), .B(n12412), .Z(n12405) );
  AND U13717 ( .A(n12406), .B(n12405), .Z(n12757) );
  NOR U13718 ( .A(n12756), .B(n12757), .Z(n12410) );
  XNOR U13719 ( .A(n12408), .B(n12407), .Z(n12409) );
  NANDN U13720 ( .A(n12410), .B(n12409), .Z(n22543) );
  XNOR U13721 ( .A(n12410), .B(n12409), .Z(n24780) );
  XNOR U13722 ( .A(n12412), .B(n12411), .Z(n12759) );
  AND U13723 ( .A(a[63]), .B(b[29]), .Z(n12753) );
  NAND U13724 ( .A(a[62]), .B(b[29]), .Z(n12746) );
  AND U13725 ( .A(a[61]), .B(b[29]), .Z(n12741) );
  NAND U13726 ( .A(a[60]), .B(b[29]), .Z(n12732) );
  AND U13727 ( .A(a[59]), .B(b[29]), .Z(n12729) );
  NAND U13728 ( .A(a[58]), .B(b[29]), .Z(n12722) );
  AND U13729 ( .A(a[57]), .B(b[29]), .Z(n12717) );
  NAND U13730 ( .A(a[56]), .B(b[29]), .Z(n12710) );
  AND U13731 ( .A(a[55]), .B(b[29]), .Z(n12705) );
  NAND U13732 ( .A(a[54]), .B(b[29]), .Z(n12698) );
  AND U13733 ( .A(a[53]), .B(b[29]), .Z(n12693) );
  NAND U13734 ( .A(a[52]), .B(b[29]), .Z(n12686) );
  AND U13735 ( .A(a[51]), .B(b[29]), .Z(n12681) );
  NAND U13736 ( .A(a[50]), .B(b[29]), .Z(n12674) );
  AND U13737 ( .A(a[49]), .B(b[29]), .Z(n12669) );
  NAND U13738 ( .A(a[48]), .B(b[29]), .Z(n12662) );
  AND U13739 ( .A(a[47]), .B(b[29]), .Z(n12657) );
  NAND U13740 ( .A(a[46]), .B(b[29]), .Z(n12650) );
  AND U13741 ( .A(a[45]), .B(b[29]), .Z(n12645) );
  NAND U13742 ( .A(a[44]), .B(b[29]), .Z(n12638) );
  AND U13743 ( .A(a[43]), .B(b[29]), .Z(n12633) );
  NAND U13744 ( .A(a[42]), .B(b[29]), .Z(n12626) );
  AND U13745 ( .A(a[41]), .B(b[29]), .Z(n12621) );
  NAND U13746 ( .A(a[40]), .B(b[29]), .Z(n12614) );
  AND U13747 ( .A(a[39]), .B(b[29]), .Z(n12609) );
  NAND U13748 ( .A(a[37]), .B(b[29]), .Z(n12596) );
  AND U13749 ( .A(a[36]), .B(b[29]), .Z(n12983) );
  XOR U13750 ( .A(n12414), .B(n12413), .Z(n12982) );
  XNOR U13751 ( .A(n12416), .B(n12415), .Z(n12968) );
  XNOR U13752 ( .A(n12420), .B(n12419), .Z(n12953) );
  NAND U13753 ( .A(a[28]), .B(b[29]), .Z(n12561) );
  XNOR U13754 ( .A(n12424), .B(n12423), .Z(n12931) );
  XNOR U13755 ( .A(n12426), .B(n12425), .Z(n12918) );
  AND U13756 ( .A(a[14]), .B(b[29]), .Z(n12497) );
  XNOR U13757 ( .A(n12428), .B(n12427), .Z(n12894) );
  AND U13758 ( .A(a[4]), .B(b[29]), .Z(n12447) );
  AND U13759 ( .A(b[29]), .B(a[0]), .Z(n13060) );
  AND U13760 ( .A(a[1]), .B(b[30]), .Z(n12434) );
  AND U13761 ( .A(n13060), .B(n12434), .Z(n12431) );
  NAND U13762 ( .A(a[2]), .B(n12431), .Z(n12438) );
  NAND U13763 ( .A(b[30]), .B(a[1]), .Z(n12432) );
  XOR U13764 ( .A(n12433), .B(n12432), .Z(n12834) );
  NAND U13765 ( .A(n12434), .B(a[0]), .Z(n12435) );
  XNOR U13766 ( .A(a[2]), .B(n12435), .Z(n12436) );
  AND U13767 ( .A(b[29]), .B(n12436), .Z(n12835) );
  NANDN U13768 ( .A(n12834), .B(n12835), .Z(n12437) );
  AND U13769 ( .A(n12438), .B(n12437), .Z(n12441) );
  NANDN U13770 ( .A(n12441), .B(n12442), .Z(n12444) );
  NAND U13771 ( .A(a[3]), .B(b[29]), .Z(n12842) );
  NANDN U13772 ( .A(n12842), .B(n12843), .Z(n12443) );
  AND U13773 ( .A(n12444), .B(n12443), .Z(n12448) );
  NANDN U13774 ( .A(n12447), .B(n12448), .Z(n12450) );
  XOR U13775 ( .A(n12446), .B(n12445), .Z(n12824) );
  NANDN U13776 ( .A(n12824), .B(n12825), .Z(n12449) );
  AND U13777 ( .A(n12450), .B(n12449), .Z(n12454) );
  XOR U13778 ( .A(n12452), .B(n12451), .Z(n12453) );
  NAND U13779 ( .A(n12454), .B(n12453), .Z(n12456) );
  NAND U13780 ( .A(a[5]), .B(b[29]), .Z(n12850) );
  XOR U13781 ( .A(n12454), .B(n12453), .Z(n12851) );
  NANDN U13782 ( .A(n12850), .B(n12851), .Z(n12455) );
  AND U13783 ( .A(n12456), .B(n12455), .Z(n12459) );
  NANDN U13784 ( .A(n12459), .B(n12460), .Z(n12462) );
  NAND U13785 ( .A(a[6]), .B(b[29]), .Z(n12856) );
  NANDN U13786 ( .A(n12856), .B(n12857), .Z(n12461) );
  AND U13787 ( .A(n12462), .B(n12461), .Z(n12465) );
  NANDN U13788 ( .A(n12465), .B(n12466), .Z(n12468) );
  AND U13789 ( .A(a[7]), .B(b[29]), .Z(n12862) );
  NAND U13790 ( .A(n12863), .B(n12862), .Z(n12467) );
  AND U13791 ( .A(n12468), .B(n12467), .Z(n12469) );
  AND U13792 ( .A(a[8]), .B(b[29]), .Z(n12470) );
  NANDN U13793 ( .A(n12469), .B(n12470), .Z(n12474) );
  NAND U13794 ( .A(n12869), .B(n12868), .Z(n12473) );
  NAND U13795 ( .A(n12474), .B(n12473), .Z(n12475) );
  NAND U13796 ( .A(n12476), .B(n12475), .Z(n12478) );
  AND U13797 ( .A(a[9]), .B(b[29]), .Z(n12877) );
  XOR U13798 ( .A(n12476), .B(n12475), .Z(n12876) );
  NAND U13799 ( .A(n12877), .B(n12876), .Z(n12477) );
  AND U13800 ( .A(n12478), .B(n12477), .Z(n12481) );
  AND U13801 ( .A(a[10]), .B(b[29]), .Z(n12482) );
  NANDN U13802 ( .A(n12481), .B(n12482), .Z(n12484) );
  XOR U13803 ( .A(n12480), .B(n12479), .Z(n12881) );
  NAND U13804 ( .A(n12881), .B(n12880), .Z(n12483) );
  AND U13805 ( .A(n12484), .B(n12483), .Z(n12487) );
  XOR U13806 ( .A(n12486), .B(n12485), .Z(n12488) );
  NANDN U13807 ( .A(n12487), .B(n12488), .Z(n12490) );
  AND U13808 ( .A(a[11]), .B(b[29]), .Z(n12887) );
  NAND U13809 ( .A(n12887), .B(n12886), .Z(n12489) );
  AND U13810 ( .A(n12490), .B(n12489), .Z(n12493) );
  AND U13811 ( .A(a[12]), .B(b[29]), .Z(n12494) );
  NANDN U13812 ( .A(n12493), .B(n12494), .Z(n12496) );
  XOR U13813 ( .A(n12492), .B(n12491), .Z(n12823) );
  NAND U13814 ( .A(n12823), .B(n12822), .Z(n12495) );
  NAND U13815 ( .A(n12496), .B(n12495), .Z(n12895) );
  NAND U13816 ( .A(a[13]), .B(b[29]), .Z(n12897) );
  NANDN U13817 ( .A(n12497), .B(n12498), .Z(n12503) );
  NAND U13818 ( .A(n12820), .B(n12821), .Z(n12502) );
  NAND U13819 ( .A(n12503), .B(n12502), .Z(n12902) );
  XOR U13820 ( .A(n12505), .B(n12504), .Z(n12901) );
  AND U13821 ( .A(a[15]), .B(b[29]), .Z(n12900) );
  AND U13822 ( .A(a[16]), .B(b[29]), .Z(n12508) );
  NANDN U13823 ( .A(n12509), .B(n12508), .Z(n12511) );
  XOR U13824 ( .A(n12507), .B(n12506), .Z(n12819) );
  XNOR U13825 ( .A(n12509), .B(n12508), .Z(n12818) );
  NAND U13826 ( .A(n12819), .B(n12818), .Z(n12510) );
  AND U13827 ( .A(n12511), .B(n12510), .Z(n12908) );
  XOR U13828 ( .A(n12513), .B(n12512), .Z(n12514) );
  IV U13829 ( .A(n12514), .Z(n12909) );
  NAND U13830 ( .A(a[17]), .B(b[29]), .Z(n12907) );
  NAND U13831 ( .A(a[18]), .B(b[29]), .Z(n12515) );
  NANDN U13832 ( .A(n12516), .B(n12515), .Z(n12521) );
  XNOR U13833 ( .A(n12516), .B(n12515), .Z(n12816) );
  NAND U13834 ( .A(n12816), .B(n12817), .Z(n12520) );
  AND U13835 ( .A(n12521), .B(n12520), .Z(n12917) );
  AND U13836 ( .A(a[19]), .B(b[29]), .Z(n12916) );
  AND U13837 ( .A(a[20]), .B(b[29]), .Z(n12526) );
  NANDN U13838 ( .A(n12527), .B(n12526), .Z(n12529) );
  XNOR U13839 ( .A(n12523), .B(n12522), .Z(n12524) );
  XNOR U13840 ( .A(n12525), .B(n12524), .Z(n12815) );
  XNOR U13841 ( .A(n12527), .B(n12526), .Z(n12814) );
  NAND U13842 ( .A(n12815), .B(n12814), .Z(n12528) );
  AND U13843 ( .A(n12529), .B(n12528), .Z(n12921) );
  NAND U13844 ( .A(a[21]), .B(b[29]), .Z(n12923) );
  AND U13845 ( .A(a[22]), .B(b[29]), .Z(n12532) );
  NANDN U13846 ( .A(n12533), .B(n12532), .Z(n12538) );
  XNOR U13847 ( .A(n12533), .B(n12532), .Z(n12813) );
  NAND U13848 ( .A(n12813), .B(n12812), .Z(n12537) );
  NAND U13849 ( .A(n12538), .B(n12537), .Z(n12932) );
  AND U13850 ( .A(a[23]), .B(b[29]), .Z(n12930) );
  AND U13851 ( .A(a[24]), .B(b[29]), .Z(n12539) );
  NANDN U13852 ( .A(n12540), .B(n12539), .Z(n12546) );
  XOR U13853 ( .A(n12540), .B(n12539), .Z(n12935) );
  XNOR U13854 ( .A(n12542), .B(n12541), .Z(n12543) );
  XNOR U13855 ( .A(n12544), .B(n12543), .Z(n12936) );
  NANDN U13856 ( .A(n12935), .B(n12936), .Z(n12545) );
  NAND U13857 ( .A(n12546), .B(n12545), .Z(n12941) );
  NAND U13858 ( .A(a[25]), .B(b[29]), .Z(n12939) );
  AND U13859 ( .A(a[26]), .B(b[29]), .Z(n12552) );
  NANDN U13860 ( .A(n12551), .B(n12552), .Z(n12554) );
  XNOR U13861 ( .A(n12548), .B(n12547), .Z(n12549) );
  XNOR U13862 ( .A(n12550), .B(n12549), .Z(n12811) );
  NAND U13863 ( .A(n12811), .B(n12810), .Z(n12553) );
  NAND U13864 ( .A(n12554), .B(n12553), .Z(n12948) );
  XOR U13865 ( .A(n12556), .B(n12555), .Z(n12947) );
  AND U13866 ( .A(a[27]), .B(b[29]), .Z(n12946) );
  NANDN U13867 ( .A(n12561), .B(n12562), .Z(n12564) );
  XOR U13868 ( .A(n12558), .B(n12557), .Z(n12559) );
  XNOR U13869 ( .A(n12560), .B(n12559), .Z(n12809) );
  NAND U13870 ( .A(n12809), .B(n12808), .Z(n12563) );
  NAND U13871 ( .A(n12564), .B(n12563), .Z(n12954) );
  NAND U13872 ( .A(a[29]), .B(b[29]), .Z(n12956) );
  AND U13873 ( .A(a[30]), .B(b[29]), .Z(n12569) );
  NANDN U13874 ( .A(n12570), .B(n12569), .Z(n12572) );
  XNOR U13875 ( .A(n12566), .B(n12565), .Z(n12567) );
  XNOR U13876 ( .A(n12568), .B(n12567), .Z(n12807) );
  XNOR U13877 ( .A(n12570), .B(n12569), .Z(n12806) );
  NAND U13878 ( .A(n12807), .B(n12806), .Z(n12571) );
  NAND U13879 ( .A(n12572), .B(n12571), .Z(n12963) );
  NAND U13880 ( .A(a[31]), .B(b[29]), .Z(n12961) );
  AND U13881 ( .A(a[32]), .B(b[29]), .Z(n12577) );
  NANDN U13882 ( .A(n12576), .B(n12577), .Z(n12579) );
  NAND U13883 ( .A(n12805), .B(n12804), .Z(n12578) );
  NAND U13884 ( .A(n12579), .B(n12578), .Z(n12969) );
  NAND U13885 ( .A(a[33]), .B(b[29]), .Z(n12971) );
  AND U13886 ( .A(a[34]), .B(b[29]), .Z(n12580) );
  NANDN U13887 ( .A(n12581), .B(n12580), .Z(n12587) );
  XNOR U13888 ( .A(n12581), .B(n12580), .Z(n12803) );
  XNOR U13889 ( .A(n12583), .B(n12582), .Z(n12584) );
  XNOR U13890 ( .A(n12585), .B(n12584), .Z(n12802) );
  NAND U13891 ( .A(n12803), .B(n12802), .Z(n12586) );
  AND U13892 ( .A(n12587), .B(n12586), .Z(n12591) );
  NAND U13893 ( .A(n12591), .B(n12590), .Z(n12593) );
  XOR U13894 ( .A(n12591), .B(n12590), .Z(n12977) );
  NAND U13895 ( .A(a[35]), .B(b[29]), .Z(n12976) );
  NAND U13896 ( .A(n12977), .B(n12976), .Z(n12592) );
  AND U13897 ( .A(n12593), .B(n12592), .Z(n12985) );
  NANDN U13898 ( .A(n12596), .B(n12597), .Z(n12599) );
  XOR U13899 ( .A(n12595), .B(n12594), .Z(n12800) );
  XNOR U13900 ( .A(n12597), .B(n12596), .Z(n12801) );
  NANDN U13901 ( .A(n12800), .B(n12801), .Z(n12598) );
  AND U13902 ( .A(n12599), .B(n12598), .Z(n12603) );
  AND U13903 ( .A(a[38]), .B(b[29]), .Z(n12602) );
  NANDN U13904 ( .A(n12603), .B(n12602), .Z(n12605) );
  XOR U13905 ( .A(n12601), .B(n12600), .Z(n12988) );
  XNOR U13906 ( .A(n12603), .B(n12602), .Z(n12989) );
  NANDN U13907 ( .A(n12988), .B(n12989), .Z(n12604) );
  AND U13908 ( .A(n12605), .B(n12604), .Z(n12608) );
  NANDN U13909 ( .A(n12609), .B(n12608), .Z(n12611) );
  XOR U13910 ( .A(n12607), .B(n12606), .Z(n12797) );
  XNOR U13911 ( .A(n12609), .B(n12608), .Z(n12796) );
  NANDN U13912 ( .A(n12797), .B(n12796), .Z(n12610) );
  AND U13913 ( .A(n12611), .B(n12610), .Z(n12615) );
  NANDN U13914 ( .A(n12614), .B(n12615), .Z(n12617) );
  XOR U13915 ( .A(n12613), .B(n12612), .Z(n12992) );
  XNOR U13916 ( .A(n12615), .B(n12614), .Z(n12993) );
  NANDN U13917 ( .A(n12992), .B(n12993), .Z(n12616) );
  AND U13918 ( .A(n12617), .B(n12616), .Z(n12620) );
  NANDN U13919 ( .A(n12621), .B(n12620), .Z(n12623) );
  XOR U13920 ( .A(n12619), .B(n12618), .Z(n12793) );
  XNOR U13921 ( .A(n12621), .B(n12620), .Z(n12792) );
  NANDN U13922 ( .A(n12793), .B(n12792), .Z(n12622) );
  AND U13923 ( .A(n12623), .B(n12622), .Z(n12627) );
  NANDN U13924 ( .A(n12626), .B(n12627), .Z(n12629) );
  XOR U13925 ( .A(n12625), .B(n12624), .Z(n12996) );
  XNOR U13926 ( .A(n12627), .B(n12626), .Z(n12997) );
  NANDN U13927 ( .A(n12996), .B(n12997), .Z(n12628) );
  AND U13928 ( .A(n12629), .B(n12628), .Z(n12632) );
  NANDN U13929 ( .A(n12633), .B(n12632), .Z(n12635) );
  XOR U13930 ( .A(n12631), .B(n12630), .Z(n12789) );
  XNOR U13931 ( .A(n12633), .B(n12632), .Z(n12788) );
  NANDN U13932 ( .A(n12789), .B(n12788), .Z(n12634) );
  AND U13933 ( .A(n12635), .B(n12634), .Z(n12639) );
  NANDN U13934 ( .A(n12638), .B(n12639), .Z(n12641) );
  XOR U13935 ( .A(n12637), .B(n12636), .Z(n13000) );
  XNOR U13936 ( .A(n12639), .B(n12638), .Z(n13001) );
  NANDN U13937 ( .A(n13000), .B(n13001), .Z(n12640) );
  AND U13938 ( .A(n12641), .B(n12640), .Z(n12644) );
  NANDN U13939 ( .A(n12645), .B(n12644), .Z(n12647) );
  XOR U13940 ( .A(n12643), .B(n12642), .Z(n12785) );
  XNOR U13941 ( .A(n12645), .B(n12644), .Z(n12784) );
  NANDN U13942 ( .A(n12785), .B(n12784), .Z(n12646) );
  AND U13943 ( .A(n12647), .B(n12646), .Z(n12651) );
  NANDN U13944 ( .A(n12650), .B(n12651), .Z(n12653) );
  XOR U13945 ( .A(n12649), .B(n12648), .Z(n13004) );
  XNOR U13946 ( .A(n12651), .B(n12650), .Z(n13005) );
  NANDN U13947 ( .A(n13004), .B(n13005), .Z(n12652) );
  AND U13948 ( .A(n12653), .B(n12652), .Z(n12656) );
  NANDN U13949 ( .A(n12657), .B(n12656), .Z(n12659) );
  XOR U13950 ( .A(n12655), .B(n12654), .Z(n12781) );
  XNOR U13951 ( .A(n12657), .B(n12656), .Z(n12780) );
  NANDN U13952 ( .A(n12781), .B(n12780), .Z(n12658) );
  AND U13953 ( .A(n12659), .B(n12658), .Z(n12663) );
  NANDN U13954 ( .A(n12662), .B(n12663), .Z(n12665) );
  XOR U13955 ( .A(n12661), .B(n12660), .Z(n13008) );
  XNOR U13956 ( .A(n12663), .B(n12662), .Z(n13009) );
  NANDN U13957 ( .A(n13008), .B(n13009), .Z(n12664) );
  AND U13958 ( .A(n12665), .B(n12664), .Z(n12668) );
  NANDN U13959 ( .A(n12669), .B(n12668), .Z(n12671) );
  XOR U13960 ( .A(n12667), .B(n12666), .Z(n12777) );
  XNOR U13961 ( .A(n12669), .B(n12668), .Z(n12776) );
  NANDN U13962 ( .A(n12777), .B(n12776), .Z(n12670) );
  AND U13963 ( .A(n12671), .B(n12670), .Z(n12675) );
  NANDN U13964 ( .A(n12674), .B(n12675), .Z(n12677) );
  XOR U13965 ( .A(n12673), .B(n12672), .Z(n13012) );
  XNOR U13966 ( .A(n12675), .B(n12674), .Z(n13013) );
  NANDN U13967 ( .A(n13012), .B(n13013), .Z(n12676) );
  AND U13968 ( .A(n12677), .B(n12676), .Z(n12680) );
  NANDN U13969 ( .A(n12681), .B(n12680), .Z(n12683) );
  XOR U13970 ( .A(n12679), .B(n12678), .Z(n12773) );
  XNOR U13971 ( .A(n12681), .B(n12680), .Z(n12772) );
  NANDN U13972 ( .A(n12773), .B(n12772), .Z(n12682) );
  AND U13973 ( .A(n12683), .B(n12682), .Z(n12687) );
  NANDN U13974 ( .A(n12686), .B(n12687), .Z(n12689) );
  XOR U13975 ( .A(n12685), .B(n12684), .Z(n13016) );
  XNOR U13976 ( .A(n12687), .B(n12686), .Z(n13017) );
  NANDN U13977 ( .A(n13016), .B(n13017), .Z(n12688) );
  AND U13978 ( .A(n12689), .B(n12688), .Z(n12692) );
  NANDN U13979 ( .A(n12693), .B(n12692), .Z(n12695) );
  XOR U13980 ( .A(n12691), .B(n12690), .Z(n12769) );
  XNOR U13981 ( .A(n12693), .B(n12692), .Z(n12768) );
  NANDN U13982 ( .A(n12769), .B(n12768), .Z(n12694) );
  AND U13983 ( .A(n12695), .B(n12694), .Z(n12699) );
  NANDN U13984 ( .A(n12698), .B(n12699), .Z(n12701) );
  XOR U13985 ( .A(n12697), .B(n12696), .Z(n13020) );
  XNOR U13986 ( .A(n12699), .B(n12698), .Z(n13021) );
  NANDN U13987 ( .A(n13020), .B(n13021), .Z(n12700) );
  AND U13988 ( .A(n12701), .B(n12700), .Z(n12704) );
  NANDN U13989 ( .A(n12705), .B(n12704), .Z(n12707) );
  XOR U13990 ( .A(n12703), .B(n12702), .Z(n12765) );
  XNOR U13991 ( .A(n12705), .B(n12704), .Z(n12764) );
  NANDN U13992 ( .A(n12765), .B(n12764), .Z(n12706) );
  AND U13993 ( .A(n12707), .B(n12706), .Z(n12711) );
  NANDN U13994 ( .A(n12710), .B(n12711), .Z(n12713) );
  XOR U13995 ( .A(n12709), .B(n12708), .Z(n13024) );
  XNOR U13996 ( .A(n12711), .B(n12710), .Z(n13025) );
  NANDN U13997 ( .A(n13024), .B(n13025), .Z(n12712) );
  AND U13998 ( .A(n12713), .B(n12712), .Z(n12716) );
  NANDN U13999 ( .A(n12717), .B(n12716), .Z(n12719) );
  XOR U14000 ( .A(n12715), .B(n12714), .Z(n12761) );
  XNOR U14001 ( .A(n12717), .B(n12716), .Z(n12760) );
  NANDN U14002 ( .A(n12761), .B(n12760), .Z(n12718) );
  AND U14003 ( .A(n12719), .B(n12718), .Z(n12723) );
  NANDN U14004 ( .A(n12722), .B(n12723), .Z(n12725) );
  XOR U14005 ( .A(n12721), .B(n12720), .Z(n13028) );
  XNOR U14006 ( .A(n12723), .B(n12722), .Z(n13029) );
  NANDN U14007 ( .A(n13028), .B(n13029), .Z(n12724) );
  AND U14008 ( .A(n12725), .B(n12724), .Z(n12728) );
  NANDN U14009 ( .A(n12729), .B(n12728), .Z(n12731) );
  XOR U14010 ( .A(n12727), .B(n12726), .Z(n13033) );
  XNOR U14011 ( .A(n12729), .B(n12728), .Z(n13032) );
  NANDN U14012 ( .A(n13033), .B(n13032), .Z(n12730) );
  AND U14013 ( .A(n12731), .B(n12730), .Z(n12733) );
  NANDN U14014 ( .A(n12732), .B(n12733), .Z(n12737) );
  XOR U14015 ( .A(n12733), .B(n12732), .Z(n13667) );
  XNOR U14016 ( .A(n12735), .B(n12734), .Z(n13668) );
  NANDN U14017 ( .A(n13667), .B(n13668), .Z(n12736) );
  AND U14018 ( .A(n12737), .B(n12736), .Z(n12740) );
  NANDN U14019 ( .A(n12741), .B(n12740), .Z(n12743) );
  XOR U14020 ( .A(n12739), .B(n12738), .Z(n13680) );
  XNOR U14021 ( .A(n12741), .B(n12740), .Z(n13679) );
  NANDN U14022 ( .A(n13680), .B(n13679), .Z(n12742) );
  AND U14023 ( .A(n12743), .B(n12742), .Z(n12747) );
  NANDN U14024 ( .A(n12746), .B(n12747), .Z(n12749) );
  XOR U14025 ( .A(n12745), .B(n12744), .Z(n13699) );
  XNOR U14026 ( .A(n12747), .B(n12746), .Z(n13700) );
  NANDN U14027 ( .A(n13699), .B(n13700), .Z(n12748) );
  AND U14028 ( .A(n12749), .B(n12748), .Z(n12752) );
  NANDN U14029 ( .A(n12753), .B(n12752), .Z(n12755) );
  XOR U14030 ( .A(n12751), .B(n12750), .Z(n22523) );
  XNOR U14031 ( .A(n12753), .B(n12752), .Z(n22522) );
  NANDN U14032 ( .A(n22523), .B(n22522), .Z(n12754) );
  AND U14033 ( .A(n12755), .B(n12754), .Z(n12758) );
  AND U14034 ( .A(n12759), .B(n12758), .Z(n22539) );
  XNOR U14035 ( .A(n12757), .B(n12756), .Z(n22538) );
  NANDN U14036 ( .A(n22539), .B(n22538), .Z(n22541) );
  XNOR U14037 ( .A(n12759), .B(n12758), .Z(n24776) );
  AND U14038 ( .A(a[58]), .B(b[28]), .Z(n12762) );
  XOR U14039 ( .A(n12761), .B(n12760), .Z(n12763) );
  XNOR U14040 ( .A(n12763), .B(n12762), .Z(n13325) );
  AND U14041 ( .A(a[56]), .B(b[28]), .Z(n12766) );
  XOR U14042 ( .A(n12765), .B(n12764), .Z(n12767) );
  XNOR U14043 ( .A(n12767), .B(n12766), .Z(n13315) );
  AND U14044 ( .A(a[54]), .B(b[28]), .Z(n12770) );
  XOR U14045 ( .A(n12769), .B(n12768), .Z(n12771) );
  XNOR U14046 ( .A(n12771), .B(n12770), .Z(n13305) );
  AND U14047 ( .A(a[52]), .B(b[28]), .Z(n12774) );
  XOR U14048 ( .A(n12773), .B(n12772), .Z(n12775) );
  XNOR U14049 ( .A(n12775), .B(n12774), .Z(n13295) );
  AND U14050 ( .A(a[50]), .B(b[28]), .Z(n12778) );
  XOR U14051 ( .A(n12777), .B(n12776), .Z(n12779) );
  XNOR U14052 ( .A(n12779), .B(n12778), .Z(n13285) );
  AND U14053 ( .A(a[48]), .B(b[28]), .Z(n12782) );
  XOR U14054 ( .A(n12781), .B(n12780), .Z(n12783) );
  XNOR U14055 ( .A(n12783), .B(n12782), .Z(n13275) );
  AND U14056 ( .A(a[46]), .B(b[28]), .Z(n12786) );
  XOR U14057 ( .A(n12785), .B(n12784), .Z(n12787) );
  XNOR U14058 ( .A(n12787), .B(n12786), .Z(n13265) );
  AND U14059 ( .A(a[44]), .B(b[28]), .Z(n12790) );
  XOR U14060 ( .A(n12789), .B(n12788), .Z(n12791) );
  XNOR U14061 ( .A(n12791), .B(n12790), .Z(n13255) );
  AND U14062 ( .A(a[42]), .B(b[28]), .Z(n12794) );
  XOR U14063 ( .A(n12793), .B(n12792), .Z(n12795) );
  XNOR U14064 ( .A(n12795), .B(n12794), .Z(n13245) );
  AND U14065 ( .A(a[40]), .B(b[28]), .Z(n12798) );
  XOR U14066 ( .A(n12797), .B(n12796), .Z(n12799) );
  XNOR U14067 ( .A(n12799), .B(n12798), .Z(n13235) );
  AND U14068 ( .A(a[38]), .B(b[28]), .Z(n12986) );
  XNOR U14069 ( .A(n12801), .B(n12800), .Z(n12987) );
  AND U14070 ( .A(a[37]), .B(b[28]), .Z(n12980) );
  XNOR U14071 ( .A(n12803), .B(n12802), .Z(n13211) );
  XNOR U14072 ( .A(n12805), .B(n12804), .Z(n13205) );
  XNOR U14073 ( .A(n12807), .B(n12806), .Z(n13195) );
  XNOR U14074 ( .A(n12809), .B(n12808), .Z(n13184) );
  XNOR U14075 ( .A(n12811), .B(n12810), .Z(n13178) );
  AND U14076 ( .A(a[24]), .B(b[28]), .Z(n12928) );
  XNOR U14077 ( .A(n12813), .B(n12812), .Z(n13159) );
  XNOR U14078 ( .A(n12815), .B(n12814), .Z(n13151) );
  XOR U14079 ( .A(n12817), .B(n12816), .Z(n13142) );
  XNOR U14080 ( .A(n12819), .B(n12818), .Z(n13135) );
  XOR U14081 ( .A(n12821), .B(n12820), .Z(n13127) );
  XNOR U14082 ( .A(n12823), .B(n12822), .Z(n13118) );
  AND U14083 ( .A(a[8]), .B(b[28]), .Z(n12864) );
  AND U14084 ( .A(b[28]), .B(a[0]), .Z(n13377) );
  AND U14085 ( .A(a[1]), .B(b[29]), .Z(n12829) );
  AND U14086 ( .A(n13377), .B(n12829), .Z(n12826) );
  NAND U14087 ( .A(a[2]), .B(n12826), .Z(n12833) );
  NAND U14088 ( .A(b[29]), .B(a[1]), .Z(n12827) );
  XOR U14089 ( .A(n12828), .B(n12827), .Z(n13066) );
  NAND U14090 ( .A(n12829), .B(a[0]), .Z(n12830) );
  XNOR U14091 ( .A(a[2]), .B(n12830), .Z(n12831) );
  AND U14092 ( .A(b[28]), .B(n12831), .Z(n13067) );
  NANDN U14093 ( .A(n13066), .B(n13067), .Z(n12832) );
  AND U14094 ( .A(n12833), .B(n12832), .Z(n12836) );
  NANDN U14095 ( .A(n12836), .B(n12837), .Z(n12839) );
  AND U14096 ( .A(a[3]), .B(b[28]), .Z(n13072) );
  NAND U14097 ( .A(n13073), .B(n13072), .Z(n12838) );
  AND U14098 ( .A(n12839), .B(n12838), .Z(n12840) );
  AND U14099 ( .A(a[4]), .B(b[28]), .Z(n12841) );
  NANDN U14100 ( .A(n12840), .B(n12841), .Z(n12845) );
  NAND U14101 ( .A(n13079), .B(n13078), .Z(n12844) );
  NAND U14102 ( .A(n12845), .B(n12844), .Z(n12846) );
  NAND U14103 ( .A(n12847), .B(n12846), .Z(n12849) );
  NAND U14104 ( .A(a[5]), .B(b[28]), .Z(n13084) );
  XOR U14105 ( .A(n12847), .B(n12846), .Z(n13085) );
  NANDN U14106 ( .A(n13084), .B(n13085), .Z(n12848) );
  AND U14107 ( .A(n12849), .B(n12848), .Z(n12852) );
  NANDN U14108 ( .A(n12852), .B(n12853), .Z(n12855) );
  NAND U14109 ( .A(a[6]), .B(b[28]), .Z(n13090) );
  NANDN U14110 ( .A(n13090), .B(n13091), .Z(n12854) );
  AND U14111 ( .A(n12855), .B(n12854), .Z(n12858) );
  NANDN U14112 ( .A(n12858), .B(n12859), .Z(n12861) );
  NAND U14113 ( .A(a[7]), .B(b[28]), .Z(n13098) );
  NANDN U14114 ( .A(n13098), .B(n13099), .Z(n12860) );
  AND U14115 ( .A(n12861), .B(n12860), .Z(n12865) );
  NANDN U14116 ( .A(n12864), .B(n12865), .Z(n12867) );
  XOR U14117 ( .A(n12863), .B(n12862), .Z(n13056) );
  NANDN U14118 ( .A(n13056), .B(n13057), .Z(n12866) );
  AND U14119 ( .A(n12867), .B(n12866), .Z(n12871) );
  XOR U14120 ( .A(n12869), .B(n12868), .Z(n12870) );
  NAND U14121 ( .A(n12871), .B(n12870), .Z(n12873) );
  AND U14122 ( .A(a[9]), .B(b[28]), .Z(n13107) );
  XOR U14123 ( .A(n12871), .B(n12870), .Z(n13106) );
  NAND U14124 ( .A(n13107), .B(n13106), .Z(n12872) );
  AND U14125 ( .A(n12873), .B(n12872), .Z(n12874) );
  AND U14126 ( .A(a[10]), .B(b[28]), .Z(n12875) );
  NANDN U14127 ( .A(n12874), .B(n12875), .Z(n12879) );
  XOR U14128 ( .A(n12877), .B(n12876), .Z(n13054) );
  NAND U14129 ( .A(n13055), .B(n13054), .Z(n12878) );
  AND U14130 ( .A(n12879), .B(n12878), .Z(n12882) );
  XOR U14131 ( .A(n12881), .B(n12880), .Z(n12883) );
  NANDN U14132 ( .A(n12882), .B(n12883), .Z(n12885) );
  AND U14133 ( .A(a[11]), .B(b[28]), .Z(n13115) );
  NAND U14134 ( .A(n13115), .B(n13114), .Z(n12884) );
  AND U14135 ( .A(n12885), .B(n12884), .Z(n12888) );
  AND U14136 ( .A(a[12]), .B(b[28]), .Z(n12889) );
  NANDN U14137 ( .A(n12888), .B(n12889), .Z(n12891) );
  XOR U14138 ( .A(n12887), .B(n12886), .Z(n13053) );
  NAND U14139 ( .A(n13053), .B(n13052), .Z(n12890) );
  NAND U14140 ( .A(n12891), .B(n12890), .Z(n13119) );
  NAND U14141 ( .A(a[13]), .B(b[28]), .Z(n13121) );
  AND U14142 ( .A(a[14]), .B(b[28]), .Z(n12893) );
  NANDN U14143 ( .A(n12892), .B(n12893), .Z(n12899) );
  XNOR U14144 ( .A(n12893), .B(n12892), .Z(n13051) );
  XNOR U14145 ( .A(n12895), .B(n12894), .Z(n12896) );
  XNOR U14146 ( .A(n12897), .B(n12896), .Z(n13050) );
  NAND U14147 ( .A(n13051), .B(n13050), .Z(n12898) );
  NAND U14148 ( .A(n12899), .B(n12898), .Z(n13128) );
  AND U14149 ( .A(a[15]), .B(b[28]), .Z(n13126) );
  AND U14150 ( .A(a[16]), .B(b[28]), .Z(n12904) );
  NANDN U14151 ( .A(n12903), .B(n12904), .Z(n12906) );
  XNOR U14152 ( .A(n12904), .B(n12903), .Z(n13048) );
  NAND U14153 ( .A(n13049), .B(n13048), .Z(n12905) );
  NAND U14154 ( .A(n12906), .B(n12905), .Z(n13136) );
  NAND U14155 ( .A(a[17]), .B(b[28]), .Z(n13138) );
  AND U14156 ( .A(a[18]), .B(b[28]), .Z(n12911) );
  NANDN U14157 ( .A(n12910), .B(n12911), .Z(n12913) );
  XNOR U14158 ( .A(n12911), .B(n12910), .Z(n13046) );
  NAND U14159 ( .A(n13047), .B(n13046), .Z(n12912) );
  NAND U14160 ( .A(n12913), .B(n12912), .Z(n13143) );
  AND U14161 ( .A(a[19]), .B(b[28]), .Z(n13141) );
  AND U14162 ( .A(a[20]), .B(b[28]), .Z(n12915) );
  NANDN U14163 ( .A(n12914), .B(n12915), .Z(n12920) );
  XOR U14164 ( .A(n12915), .B(n12914), .Z(n13148) );
  NANDN U14165 ( .A(n13148), .B(n13149), .Z(n12919) );
  NAND U14166 ( .A(n12920), .B(n12919), .Z(n13152) );
  NAND U14167 ( .A(a[21]), .B(b[28]), .Z(n13154) );
  AND U14168 ( .A(a[22]), .B(b[28]), .Z(n12925) );
  NANDN U14169 ( .A(n12924), .B(n12925), .Z(n12927) );
  XNOR U14170 ( .A(n12925), .B(n12924), .Z(n13044) );
  NAND U14171 ( .A(n13045), .B(n13044), .Z(n12926) );
  NAND U14172 ( .A(n12927), .B(n12926), .Z(n13160) );
  NAND U14173 ( .A(a[23]), .B(b[28]), .Z(n13162) );
  NANDN U14174 ( .A(n12928), .B(n12929), .Z(n12934) );
  NAND U14175 ( .A(n13167), .B(n13168), .Z(n12933) );
  NAND U14176 ( .A(n12934), .B(n12933), .Z(n13173) );
  NAND U14177 ( .A(a[25]), .B(b[28]), .Z(n13171) );
  AND U14178 ( .A(a[26]), .B(b[28]), .Z(n12938) );
  NANDN U14179 ( .A(n12937), .B(n12938), .Z(n12943) );
  NAND U14180 ( .A(n13043), .B(n13042), .Z(n12942) );
  NAND U14181 ( .A(n12943), .B(n12942), .Z(n13179) );
  NAND U14182 ( .A(a[27]), .B(b[28]), .Z(n13181) );
  AND U14183 ( .A(a[28]), .B(b[28]), .Z(n12945) );
  NANDN U14184 ( .A(n12944), .B(n12945), .Z(n12950) );
  XNOR U14185 ( .A(n12945), .B(n12944), .Z(n13040) );
  NAND U14186 ( .A(n13040), .B(n13041), .Z(n12949) );
  NAND U14187 ( .A(n12950), .B(n12949), .Z(n13185) );
  NAND U14188 ( .A(a[29]), .B(b[28]), .Z(n13187) );
  AND U14189 ( .A(a[30]), .B(b[28]), .Z(n12952) );
  NANDN U14190 ( .A(n12951), .B(n12952), .Z(n12958) );
  XOR U14191 ( .A(n12952), .B(n12951), .Z(n13192) );
  XNOR U14192 ( .A(n12954), .B(n12953), .Z(n12955) );
  XNOR U14193 ( .A(n12956), .B(n12955), .Z(n13193) );
  NANDN U14194 ( .A(n13192), .B(n13193), .Z(n12957) );
  NAND U14195 ( .A(n12958), .B(n12957), .Z(n13196) );
  NAND U14196 ( .A(a[31]), .B(b[28]), .Z(n13198) );
  AND U14197 ( .A(a[32]), .B(b[28]), .Z(n12960) );
  NANDN U14198 ( .A(n12959), .B(n12960), .Z(n12965) );
  XNOR U14199 ( .A(n12960), .B(n12959), .Z(n13039) );
  NAND U14200 ( .A(n13039), .B(n13038), .Z(n12964) );
  NAND U14201 ( .A(n12965), .B(n12964), .Z(n13206) );
  NAND U14202 ( .A(a[33]), .B(b[28]), .Z(n13208) );
  AND U14203 ( .A(a[34]), .B(b[28]), .Z(n12967) );
  NANDN U14204 ( .A(n12966), .B(n12967), .Z(n12973) );
  XNOR U14205 ( .A(n12967), .B(n12966), .Z(n13037) );
  XNOR U14206 ( .A(n12969), .B(n12968), .Z(n12970) );
  XNOR U14207 ( .A(n12971), .B(n12970), .Z(n13036) );
  NAND U14208 ( .A(n13037), .B(n13036), .Z(n12972) );
  NAND U14209 ( .A(n12973), .B(n12972), .Z(n13212) );
  NAND U14210 ( .A(a[35]), .B(b[28]), .Z(n13214) );
  AND U14211 ( .A(a[36]), .B(b[28]), .Z(n12974) );
  NANDN U14212 ( .A(n12975), .B(n12974), .Z(n12979) );
  XOR U14213 ( .A(n12975), .B(n12974), .Z(n13219) );
  XNOR U14214 ( .A(n12977), .B(n12976), .Z(n13220) );
  NANDN U14215 ( .A(n13219), .B(n13220), .Z(n12978) );
  NAND U14216 ( .A(n12979), .B(n12978), .Z(n12981) );
  XNOR U14217 ( .A(n12981), .B(n12980), .Z(n13034) );
  XOR U14218 ( .A(n12983), .B(n12982), .Z(n12984) );
  XNOR U14219 ( .A(n12985), .B(n12984), .Z(n13035) );
  XOR U14220 ( .A(n12987), .B(n12986), .Z(n13225) );
  XNOR U14221 ( .A(n12989), .B(n12988), .Z(n12990) );
  AND U14222 ( .A(a[39]), .B(b[28]), .Z(n13229) );
  XOR U14223 ( .A(n12991), .B(n12990), .Z(n13230) );
  XNOR U14224 ( .A(n12993), .B(n12992), .Z(n12994) );
  AND U14225 ( .A(a[41]), .B(b[28]), .Z(n13239) );
  XOR U14226 ( .A(n12995), .B(n12994), .Z(n13240) );
  XNOR U14227 ( .A(n12997), .B(n12996), .Z(n12998) );
  AND U14228 ( .A(a[43]), .B(b[28]), .Z(n13249) );
  XOR U14229 ( .A(n12999), .B(n12998), .Z(n13250) );
  XNOR U14230 ( .A(n13001), .B(n13000), .Z(n13002) );
  AND U14231 ( .A(a[45]), .B(b[28]), .Z(n13259) );
  XOR U14232 ( .A(n13003), .B(n13002), .Z(n13260) );
  XNOR U14233 ( .A(n13005), .B(n13004), .Z(n13006) );
  AND U14234 ( .A(a[47]), .B(b[28]), .Z(n13269) );
  XOR U14235 ( .A(n13007), .B(n13006), .Z(n13270) );
  XNOR U14236 ( .A(n13009), .B(n13008), .Z(n13010) );
  AND U14237 ( .A(a[49]), .B(b[28]), .Z(n13279) );
  XOR U14238 ( .A(n13011), .B(n13010), .Z(n13280) );
  XNOR U14239 ( .A(n13013), .B(n13012), .Z(n13014) );
  AND U14240 ( .A(a[51]), .B(b[28]), .Z(n13289) );
  XOR U14241 ( .A(n13015), .B(n13014), .Z(n13290) );
  XNOR U14242 ( .A(n13017), .B(n13016), .Z(n13018) );
  AND U14243 ( .A(a[53]), .B(b[28]), .Z(n13299) );
  XOR U14244 ( .A(n13019), .B(n13018), .Z(n13300) );
  XNOR U14245 ( .A(n13021), .B(n13020), .Z(n13022) );
  AND U14246 ( .A(a[55]), .B(b[28]), .Z(n13309) );
  XOR U14247 ( .A(n13023), .B(n13022), .Z(n13310) );
  XNOR U14248 ( .A(n13025), .B(n13024), .Z(n13026) );
  AND U14249 ( .A(a[57]), .B(b[28]), .Z(n13319) );
  XOR U14250 ( .A(n13027), .B(n13026), .Z(n13320) );
  XNOR U14251 ( .A(n13029), .B(n13028), .Z(n13030) );
  AND U14252 ( .A(a[59]), .B(b[28]), .Z(n13329) );
  XOR U14253 ( .A(n13031), .B(n13030), .Z(n13330) );
  XOR U14254 ( .A(n13033), .B(n13032), .Z(n13661) );
  AND U14255 ( .A(a[60]), .B(b[28]), .Z(n13662) );
  XNOR U14256 ( .A(n13661), .B(n13662), .Z(n13664) );
  XOR U14257 ( .A(n13663), .B(n13664), .Z(n13657) );
  AND U14258 ( .A(a[61]), .B(b[27]), .Z(n13656) );
  NAND U14259 ( .A(a[60]), .B(b[27]), .Z(n13331) );
  AND U14260 ( .A(a[59]), .B(b[27]), .Z(n13324) );
  NAND U14261 ( .A(a[58]), .B(b[27]), .Z(n13321) );
  AND U14262 ( .A(a[57]), .B(b[27]), .Z(n13314) );
  NAND U14263 ( .A(a[56]), .B(b[27]), .Z(n13311) );
  AND U14264 ( .A(a[55]), .B(b[27]), .Z(n13304) );
  NAND U14265 ( .A(a[54]), .B(b[27]), .Z(n13301) );
  AND U14266 ( .A(a[53]), .B(b[27]), .Z(n13294) );
  NAND U14267 ( .A(a[52]), .B(b[27]), .Z(n13291) );
  AND U14268 ( .A(a[51]), .B(b[27]), .Z(n13284) );
  NAND U14269 ( .A(a[50]), .B(b[27]), .Z(n13281) );
  AND U14270 ( .A(a[49]), .B(b[27]), .Z(n13274) );
  NAND U14271 ( .A(a[48]), .B(b[27]), .Z(n13271) );
  AND U14272 ( .A(a[47]), .B(b[27]), .Z(n13264) );
  NAND U14273 ( .A(a[46]), .B(b[27]), .Z(n13261) );
  AND U14274 ( .A(a[45]), .B(b[27]), .Z(n13254) );
  NAND U14275 ( .A(a[44]), .B(b[27]), .Z(n13251) );
  AND U14276 ( .A(a[43]), .B(b[27]), .Z(n13244) );
  NAND U14277 ( .A(a[42]), .B(b[27]), .Z(n13241) );
  AND U14278 ( .A(a[41]), .B(b[27]), .Z(n13234) );
  NAND U14279 ( .A(a[39]), .B(b[27]), .Z(n13227) );
  AND U14280 ( .A(a[38]), .B(b[27]), .Z(n13558) );
  XOR U14281 ( .A(n13035), .B(n13034), .Z(n13557) );
  XNOR U14282 ( .A(n13037), .B(n13036), .Z(n13541) );
  XNOR U14283 ( .A(n13039), .B(n13038), .Z(n13533) );
  NAND U14284 ( .A(a[32]), .B(b[27]), .Z(n13199) );
  XNOR U14285 ( .A(n13041), .B(n13040), .Z(n13519) );
  XNOR U14286 ( .A(n13043), .B(n13042), .Z(n13509) );
  AND U14287 ( .A(a[26]), .B(b[27]), .Z(n13169) );
  XNOR U14288 ( .A(n13045), .B(n13044), .Z(n13490) );
  NAND U14289 ( .A(a[22]), .B(b[27]), .Z(n13155) );
  XNOR U14290 ( .A(n13047), .B(n13046), .Z(n13474) );
  XNOR U14291 ( .A(n13049), .B(n13048), .Z(n13464) );
  XNOR U14292 ( .A(n13051), .B(n13050), .Z(n13458) );
  XNOR U14293 ( .A(n13053), .B(n13052), .Z(n13448) );
  XNOR U14294 ( .A(n13055), .B(n13054), .Z(n13437) );
  AND U14295 ( .A(a[4]), .B(b[27]), .Z(n13074) );
  AND U14296 ( .A(b[27]), .B(a[0]), .Z(n13729) );
  AND U14297 ( .A(a[1]), .B(b[28]), .Z(n13061) );
  AND U14298 ( .A(n13729), .B(n13061), .Z(n13058) );
  NAND U14299 ( .A(a[2]), .B(n13058), .Z(n13065) );
  NAND U14300 ( .A(b[28]), .B(a[1]), .Z(n13059) );
  XOR U14301 ( .A(n13060), .B(n13059), .Z(n13383) );
  NAND U14302 ( .A(n13061), .B(a[0]), .Z(n13062) );
  XNOR U14303 ( .A(a[2]), .B(n13062), .Z(n13063) );
  AND U14304 ( .A(b[27]), .B(n13063), .Z(n13384) );
  NANDN U14305 ( .A(n13383), .B(n13384), .Z(n13064) );
  AND U14306 ( .A(n13065), .B(n13064), .Z(n13068) );
  NANDN U14307 ( .A(n13068), .B(n13069), .Z(n13071) );
  NAND U14308 ( .A(a[3]), .B(b[27]), .Z(n13391) );
  NANDN U14309 ( .A(n13391), .B(n13392), .Z(n13070) );
  AND U14310 ( .A(n13071), .B(n13070), .Z(n13075) );
  NANDN U14311 ( .A(n13074), .B(n13075), .Z(n13077) );
  XOR U14312 ( .A(n13073), .B(n13072), .Z(n13373) );
  NANDN U14313 ( .A(n13373), .B(n13374), .Z(n13076) );
  AND U14314 ( .A(n13077), .B(n13076), .Z(n13081) );
  XOR U14315 ( .A(n13079), .B(n13078), .Z(n13080) );
  NAND U14316 ( .A(n13081), .B(n13080), .Z(n13083) );
  NAND U14317 ( .A(a[5]), .B(b[27]), .Z(n13399) );
  XOR U14318 ( .A(n13081), .B(n13080), .Z(n13400) );
  NANDN U14319 ( .A(n13399), .B(n13400), .Z(n13082) );
  AND U14320 ( .A(n13083), .B(n13082), .Z(n13086) );
  NANDN U14321 ( .A(n13086), .B(n13087), .Z(n13089) );
  NAND U14322 ( .A(a[6]), .B(b[27]), .Z(n13405) );
  NANDN U14323 ( .A(n13405), .B(n13406), .Z(n13088) );
  AND U14324 ( .A(n13089), .B(n13088), .Z(n13092) );
  NANDN U14325 ( .A(n13092), .B(n13093), .Z(n13095) );
  AND U14326 ( .A(a[7]), .B(b[27]), .Z(n13411) );
  NAND U14327 ( .A(n13412), .B(n13411), .Z(n13094) );
  AND U14328 ( .A(n13095), .B(n13094), .Z(n13096) );
  AND U14329 ( .A(a[8]), .B(b[27]), .Z(n13097) );
  NANDN U14330 ( .A(n13096), .B(n13097), .Z(n13101) );
  NAND U14331 ( .A(n13418), .B(n13417), .Z(n13100) );
  NAND U14332 ( .A(n13101), .B(n13100), .Z(n13102) );
  NAND U14333 ( .A(n13103), .B(n13102), .Z(n13105) );
  NAND U14334 ( .A(a[9]), .B(b[27]), .Z(n13423) );
  XOR U14335 ( .A(n13103), .B(n13102), .Z(n13424) );
  NANDN U14336 ( .A(n13423), .B(n13424), .Z(n13104) );
  AND U14337 ( .A(n13105), .B(n13104), .Z(n13108) );
  AND U14338 ( .A(a[10]), .B(b[27]), .Z(n13109) );
  NANDN U14339 ( .A(n13108), .B(n13109), .Z(n13111) );
  XOR U14340 ( .A(n13107), .B(n13106), .Z(n13430) );
  NAND U14341 ( .A(n13430), .B(n13429), .Z(n13110) );
  NAND U14342 ( .A(n13111), .B(n13110), .Z(n13438) );
  AND U14343 ( .A(a[11]), .B(b[27]), .Z(n13436) );
  AND U14344 ( .A(a[12]), .B(b[27]), .Z(n13112) );
  NANDN U14345 ( .A(n13113), .B(n13112), .Z(n13117) );
  XNOR U14346 ( .A(n13113), .B(n13112), .Z(n13443) );
  XOR U14347 ( .A(n13115), .B(n13114), .Z(n13442) );
  NAND U14348 ( .A(n13443), .B(n13442), .Z(n13116) );
  NAND U14349 ( .A(n13117), .B(n13116), .Z(n13449) );
  NAND U14350 ( .A(a[13]), .B(b[27]), .Z(n13451) );
  AND U14351 ( .A(a[14]), .B(b[27]), .Z(n13122) );
  NANDN U14352 ( .A(n13123), .B(n13122), .Z(n13125) );
  XNOR U14353 ( .A(n13119), .B(n13118), .Z(n13120) );
  XNOR U14354 ( .A(n13121), .B(n13120), .Z(n13372) );
  XNOR U14355 ( .A(n13123), .B(n13122), .Z(n13371) );
  NAND U14356 ( .A(n13372), .B(n13371), .Z(n13124) );
  NAND U14357 ( .A(n13125), .B(n13124), .Z(n13459) );
  NAND U14358 ( .A(a[15]), .B(b[27]), .Z(n13461) );
  AND U14359 ( .A(a[16]), .B(b[27]), .Z(n13129) );
  NANDN U14360 ( .A(n13130), .B(n13129), .Z(n13132) );
  XNOR U14361 ( .A(n13130), .B(n13129), .Z(n13369) );
  NAND U14362 ( .A(n13370), .B(n13369), .Z(n13131) );
  NAND U14363 ( .A(n13132), .B(n13131), .Z(n13465) );
  NAND U14364 ( .A(a[17]), .B(b[27]), .Z(n13467) );
  AND U14365 ( .A(a[18]), .B(b[27]), .Z(n13133) );
  NANDN U14366 ( .A(n13134), .B(n13133), .Z(n13140) );
  XNOR U14367 ( .A(n13134), .B(n13133), .Z(n13368) );
  XNOR U14368 ( .A(n13136), .B(n13135), .Z(n13137) );
  XNOR U14369 ( .A(n13138), .B(n13137), .Z(n13367) );
  NAND U14370 ( .A(n13368), .B(n13367), .Z(n13139) );
  NAND U14371 ( .A(n13140), .B(n13139), .Z(n13475) );
  NAND U14372 ( .A(a[19]), .B(b[27]), .Z(n13477) );
  AND U14373 ( .A(a[20]), .B(b[27]), .Z(n13144) );
  NANDN U14374 ( .A(n13145), .B(n13144), .Z(n13147) );
  XNOR U14375 ( .A(n13145), .B(n13144), .Z(n13365) );
  NAND U14376 ( .A(n13366), .B(n13365), .Z(n13146) );
  AND U14377 ( .A(n13147), .B(n13146), .Z(n13483) );
  IV U14378 ( .A(n13150), .Z(n13484) );
  NAND U14379 ( .A(a[21]), .B(b[27]), .Z(n13482) );
  NANDN U14380 ( .A(n13155), .B(n13156), .Z(n13158) );
  XNOR U14381 ( .A(n13152), .B(n13151), .Z(n13153) );
  XNOR U14382 ( .A(n13154), .B(n13153), .Z(n13488) );
  NAND U14383 ( .A(n13488), .B(n13487), .Z(n13157) );
  NAND U14384 ( .A(n13158), .B(n13157), .Z(n13491) );
  NAND U14385 ( .A(a[23]), .B(b[27]), .Z(n13493) );
  AND U14386 ( .A(a[24]), .B(b[27]), .Z(n13163) );
  NANDN U14387 ( .A(n13164), .B(n13163), .Z(n13166) );
  XNOR U14388 ( .A(n13160), .B(n13159), .Z(n13161) );
  XNOR U14389 ( .A(n13162), .B(n13161), .Z(n13364) );
  XNOR U14390 ( .A(n13164), .B(n13163), .Z(n13363) );
  NAND U14391 ( .A(n13364), .B(n13363), .Z(n13165) );
  AND U14392 ( .A(n13166), .B(n13165), .Z(n13501) );
  XNOR U14393 ( .A(n13168), .B(n13167), .Z(n13502) );
  NAND U14394 ( .A(a[25]), .B(b[27]), .Z(n13500) );
  NANDN U14395 ( .A(n13169), .B(n13170), .Z(n13175) );
  NAND U14396 ( .A(n13505), .B(n13506), .Z(n13174) );
  AND U14397 ( .A(n13175), .B(n13174), .Z(n13508) );
  NAND U14398 ( .A(a[27]), .B(b[27]), .Z(n13511) );
  AND U14399 ( .A(a[28]), .B(b[27]), .Z(n13176) );
  NANDN U14400 ( .A(n13177), .B(n13176), .Z(n13183) );
  XOR U14401 ( .A(n13177), .B(n13176), .Z(n13361) );
  XNOR U14402 ( .A(n13179), .B(n13178), .Z(n13180) );
  XNOR U14403 ( .A(n13181), .B(n13180), .Z(n13362) );
  NANDN U14404 ( .A(n13361), .B(n13362), .Z(n13182) );
  NAND U14405 ( .A(n13183), .B(n13182), .Z(n13520) );
  NAND U14406 ( .A(a[29]), .B(b[27]), .Z(n13518) );
  AND U14407 ( .A(a[30]), .B(b[27]), .Z(n13189) );
  NANDN U14408 ( .A(n13188), .B(n13189), .Z(n13191) );
  XNOR U14409 ( .A(n13185), .B(n13184), .Z(n13186) );
  XNOR U14410 ( .A(n13187), .B(n13186), .Z(n13360) );
  NAND U14411 ( .A(n13360), .B(n13359), .Z(n13190) );
  AND U14412 ( .A(n13191), .B(n13190), .Z(n13523) );
  IV U14413 ( .A(n13194), .Z(n13524) );
  AND U14414 ( .A(a[31]), .B(b[27]), .Z(n13526) );
  NANDN U14415 ( .A(n13199), .B(n13200), .Z(n13202) );
  XNOR U14416 ( .A(n13196), .B(n13195), .Z(n13197) );
  XNOR U14417 ( .A(n13198), .B(n13197), .Z(n13532) );
  NAND U14418 ( .A(n13532), .B(n13531), .Z(n13201) );
  NAND U14419 ( .A(n13202), .B(n13201), .Z(n13534) );
  NAND U14420 ( .A(a[33]), .B(b[27]), .Z(n13536) );
  AND U14421 ( .A(a[34]), .B(b[27]), .Z(n13203) );
  NANDN U14422 ( .A(n13204), .B(n13203), .Z(n13210) );
  XNOR U14423 ( .A(n13204), .B(n13203), .Z(n13358) );
  XNOR U14424 ( .A(n13206), .B(n13205), .Z(n13207) );
  XNOR U14425 ( .A(n13208), .B(n13207), .Z(n13357) );
  NAND U14426 ( .A(n13358), .B(n13357), .Z(n13209) );
  NAND U14427 ( .A(n13210), .B(n13209), .Z(n13542) );
  NAND U14428 ( .A(a[35]), .B(b[27]), .Z(n13544) );
  AND U14429 ( .A(a[36]), .B(b[27]), .Z(n13215) );
  NANDN U14430 ( .A(n13216), .B(n13215), .Z(n13218) );
  XNOR U14431 ( .A(n13212), .B(n13211), .Z(n13213) );
  XNOR U14432 ( .A(n13214), .B(n13213), .Z(n13356) );
  XNOR U14433 ( .A(n13216), .B(n13215), .Z(n13355) );
  NAND U14434 ( .A(n13356), .B(n13355), .Z(n13217) );
  AND U14435 ( .A(n13218), .B(n13217), .Z(n13222) );
  NAND U14436 ( .A(n13222), .B(n13221), .Z(n13224) );
  XOR U14437 ( .A(n13222), .B(n13221), .Z(n13552) );
  NAND U14438 ( .A(a[37]), .B(b[27]), .Z(n13551) );
  NAND U14439 ( .A(n13552), .B(n13551), .Z(n13223) );
  AND U14440 ( .A(n13224), .B(n13223), .Z(n13560) );
  XOR U14441 ( .A(n13226), .B(n13225), .Z(n13353) );
  XNOR U14442 ( .A(n13228), .B(n13227), .Z(n13354) );
  AND U14443 ( .A(a[40]), .B(b[27]), .Z(n13231) );
  XOR U14444 ( .A(n13230), .B(n13229), .Z(n13567) );
  XNOR U14445 ( .A(n13232), .B(n13231), .Z(n13568) );
  NANDN U14446 ( .A(n13234), .B(n13233), .Z(n13238) );
  XOR U14447 ( .A(n13234), .B(n13233), .Z(n13351) );
  XOR U14448 ( .A(n13236), .B(n13235), .Z(n13352) );
  NANDN U14449 ( .A(n13351), .B(n13352), .Z(n13237) );
  AND U14450 ( .A(n13238), .B(n13237), .Z(n13242) );
  XOR U14451 ( .A(n13240), .B(n13239), .Z(n13575) );
  XNOR U14452 ( .A(n13242), .B(n13241), .Z(n13576) );
  NANDN U14453 ( .A(n13244), .B(n13243), .Z(n13248) );
  XOR U14454 ( .A(n13244), .B(n13243), .Z(n13349) );
  XOR U14455 ( .A(n13246), .B(n13245), .Z(n13350) );
  NANDN U14456 ( .A(n13349), .B(n13350), .Z(n13247) );
  AND U14457 ( .A(n13248), .B(n13247), .Z(n13252) );
  XOR U14458 ( .A(n13250), .B(n13249), .Z(n13583) );
  XNOR U14459 ( .A(n13252), .B(n13251), .Z(n13584) );
  NANDN U14460 ( .A(n13254), .B(n13253), .Z(n13258) );
  XOR U14461 ( .A(n13254), .B(n13253), .Z(n13347) );
  XOR U14462 ( .A(n13256), .B(n13255), .Z(n13348) );
  NANDN U14463 ( .A(n13347), .B(n13348), .Z(n13257) );
  AND U14464 ( .A(n13258), .B(n13257), .Z(n13262) );
  XOR U14465 ( .A(n13260), .B(n13259), .Z(n13591) );
  XNOR U14466 ( .A(n13262), .B(n13261), .Z(n13592) );
  NANDN U14467 ( .A(n13264), .B(n13263), .Z(n13268) );
  XOR U14468 ( .A(n13264), .B(n13263), .Z(n13345) );
  XOR U14469 ( .A(n13266), .B(n13265), .Z(n13346) );
  NANDN U14470 ( .A(n13345), .B(n13346), .Z(n13267) );
  AND U14471 ( .A(n13268), .B(n13267), .Z(n13272) );
  XOR U14472 ( .A(n13270), .B(n13269), .Z(n13599) );
  XNOR U14473 ( .A(n13272), .B(n13271), .Z(n13600) );
  NANDN U14474 ( .A(n13274), .B(n13273), .Z(n13278) );
  XOR U14475 ( .A(n13274), .B(n13273), .Z(n13343) );
  XOR U14476 ( .A(n13276), .B(n13275), .Z(n13344) );
  NANDN U14477 ( .A(n13343), .B(n13344), .Z(n13277) );
  AND U14478 ( .A(n13278), .B(n13277), .Z(n13282) );
  XOR U14479 ( .A(n13280), .B(n13279), .Z(n13607) );
  XNOR U14480 ( .A(n13282), .B(n13281), .Z(n13608) );
  NANDN U14481 ( .A(n13284), .B(n13283), .Z(n13288) );
  XOR U14482 ( .A(n13284), .B(n13283), .Z(n13341) );
  XOR U14483 ( .A(n13286), .B(n13285), .Z(n13342) );
  NANDN U14484 ( .A(n13341), .B(n13342), .Z(n13287) );
  AND U14485 ( .A(n13288), .B(n13287), .Z(n13292) );
  XOR U14486 ( .A(n13290), .B(n13289), .Z(n13615) );
  XNOR U14487 ( .A(n13292), .B(n13291), .Z(n13616) );
  NANDN U14488 ( .A(n13294), .B(n13293), .Z(n13298) );
  XOR U14489 ( .A(n13294), .B(n13293), .Z(n13339) );
  XOR U14490 ( .A(n13296), .B(n13295), .Z(n13340) );
  NANDN U14491 ( .A(n13339), .B(n13340), .Z(n13297) );
  AND U14492 ( .A(n13298), .B(n13297), .Z(n13302) );
  XOR U14493 ( .A(n13300), .B(n13299), .Z(n13623) );
  XNOR U14494 ( .A(n13302), .B(n13301), .Z(n13624) );
  NANDN U14495 ( .A(n13304), .B(n13303), .Z(n13308) );
  XOR U14496 ( .A(n13304), .B(n13303), .Z(n13337) );
  XOR U14497 ( .A(n13306), .B(n13305), .Z(n13338) );
  NANDN U14498 ( .A(n13337), .B(n13338), .Z(n13307) );
  AND U14499 ( .A(n13308), .B(n13307), .Z(n13312) );
  XOR U14500 ( .A(n13310), .B(n13309), .Z(n13631) );
  XNOR U14501 ( .A(n13312), .B(n13311), .Z(n13632) );
  NANDN U14502 ( .A(n13314), .B(n13313), .Z(n13318) );
  XOR U14503 ( .A(n13314), .B(n13313), .Z(n13335) );
  XOR U14504 ( .A(n13316), .B(n13315), .Z(n13336) );
  NANDN U14505 ( .A(n13335), .B(n13336), .Z(n13317) );
  AND U14506 ( .A(n13318), .B(n13317), .Z(n13322) );
  XOR U14507 ( .A(n13320), .B(n13319), .Z(n13639) );
  XNOR U14508 ( .A(n13322), .B(n13321), .Z(n13640) );
  NANDN U14509 ( .A(n13324), .B(n13323), .Z(n13328) );
  XOR U14510 ( .A(n13324), .B(n13323), .Z(n13333) );
  XOR U14511 ( .A(n13326), .B(n13325), .Z(n13334) );
  NANDN U14512 ( .A(n13333), .B(n13334), .Z(n13327) );
  AND U14513 ( .A(n13328), .B(n13327), .Z(n13332) );
  XOR U14514 ( .A(n13330), .B(n13329), .Z(n13647) );
  XNOR U14515 ( .A(n13332), .B(n13331), .Z(n13648) );
  XOR U14516 ( .A(n13656), .B(n13655), .Z(n13658) );
  XOR U14517 ( .A(n13657), .B(n13658), .Z(n13654) );
  AND U14518 ( .A(a[62]), .B(b[26]), .Z(n13653) );
  XOR U14519 ( .A(n13334), .B(n13333), .Z(n13646) );
  AND U14520 ( .A(a[60]), .B(b[26]), .Z(n13645) );
  XOR U14521 ( .A(n13336), .B(n13335), .Z(n13638) );
  AND U14522 ( .A(a[58]), .B(b[26]), .Z(n13637) );
  XOR U14523 ( .A(n13338), .B(n13337), .Z(n13630) );
  AND U14524 ( .A(a[56]), .B(b[26]), .Z(n13629) );
  XOR U14525 ( .A(n13340), .B(n13339), .Z(n13622) );
  AND U14526 ( .A(a[54]), .B(b[26]), .Z(n13621) );
  XOR U14527 ( .A(n13342), .B(n13341), .Z(n13614) );
  AND U14528 ( .A(a[52]), .B(b[26]), .Z(n13613) );
  XOR U14529 ( .A(n13344), .B(n13343), .Z(n13606) );
  AND U14530 ( .A(a[50]), .B(b[26]), .Z(n13605) );
  XOR U14531 ( .A(n13346), .B(n13345), .Z(n13598) );
  AND U14532 ( .A(a[48]), .B(b[26]), .Z(n13597) );
  XOR U14533 ( .A(n13348), .B(n13347), .Z(n13590) );
  AND U14534 ( .A(a[46]), .B(b[26]), .Z(n13589) );
  XOR U14535 ( .A(n13350), .B(n13349), .Z(n13582) );
  AND U14536 ( .A(a[44]), .B(b[26]), .Z(n13581) );
  XOR U14537 ( .A(n13352), .B(n13351), .Z(n13574) );
  AND U14538 ( .A(a[42]), .B(b[26]), .Z(n13573) );
  NAND U14539 ( .A(a[40]), .B(b[26]), .Z(n13563) );
  XOR U14540 ( .A(n13354), .B(n13353), .Z(n13564) );
  NANDN U14541 ( .A(n13563), .B(n13564), .Z(n13566) );
  XNOR U14542 ( .A(n13356), .B(n13355), .Z(n13904) );
  XNOR U14543 ( .A(n13358), .B(n13357), .Z(n13893) );
  AND U14544 ( .A(a[32]), .B(b[26]), .Z(n13527) );
  XNOR U14545 ( .A(n13360), .B(n13359), .Z(n13878) );
  NAND U14546 ( .A(a[30]), .B(b[26]), .Z(n13516) );
  AND U14547 ( .A(a[28]), .B(b[26]), .Z(n13512) );
  AND U14548 ( .A(a[26]), .B(b[26]), .Z(n13498) );
  XNOR U14549 ( .A(n13364), .B(n13363), .Z(n13848) );
  NAND U14550 ( .A(a[24]), .B(b[26]), .Z(n13494) );
  XNOR U14551 ( .A(n13366), .B(n13365), .Z(n13833) );
  XNOR U14552 ( .A(n13368), .B(n13367), .Z(n13819) );
  XNOR U14553 ( .A(n13370), .B(n13369), .Z(n13811) );
  XNOR U14554 ( .A(n13372), .B(n13371), .Z(n13805) );
  AND U14555 ( .A(a[8]), .B(b[26]), .Z(n13413) );
  AND U14556 ( .A(b[26]), .B(a[0]), .Z(n14096) );
  AND U14557 ( .A(a[1]), .B(b[27]), .Z(n13378) );
  AND U14558 ( .A(n14096), .B(n13378), .Z(n13375) );
  NAND U14559 ( .A(a[2]), .B(n13375), .Z(n13382) );
  NAND U14560 ( .A(b[27]), .B(a[1]), .Z(n13376) );
  XOR U14561 ( .A(n13377), .B(n13376), .Z(n13735) );
  NAND U14562 ( .A(n13378), .B(a[0]), .Z(n13379) );
  XNOR U14563 ( .A(a[2]), .B(n13379), .Z(n13380) );
  AND U14564 ( .A(b[26]), .B(n13380), .Z(n13736) );
  NANDN U14565 ( .A(n13735), .B(n13736), .Z(n13381) );
  AND U14566 ( .A(n13382), .B(n13381), .Z(n13385) );
  NANDN U14567 ( .A(n13385), .B(n13386), .Z(n13388) );
  AND U14568 ( .A(a[3]), .B(b[26]), .Z(n13741) );
  NAND U14569 ( .A(n13742), .B(n13741), .Z(n13387) );
  AND U14570 ( .A(n13388), .B(n13387), .Z(n13389) );
  AND U14571 ( .A(a[4]), .B(b[26]), .Z(n13390) );
  NANDN U14572 ( .A(n13389), .B(n13390), .Z(n13394) );
  NAND U14573 ( .A(n13748), .B(n13747), .Z(n13393) );
  NAND U14574 ( .A(n13394), .B(n13393), .Z(n13395) );
  NAND U14575 ( .A(n13396), .B(n13395), .Z(n13398) );
  NAND U14576 ( .A(a[5]), .B(b[26]), .Z(n13753) );
  XOR U14577 ( .A(n13396), .B(n13395), .Z(n13754) );
  NANDN U14578 ( .A(n13753), .B(n13754), .Z(n13397) );
  AND U14579 ( .A(n13398), .B(n13397), .Z(n13401) );
  NANDN U14580 ( .A(n13401), .B(n13402), .Z(n13404) );
  NAND U14581 ( .A(a[6]), .B(b[26]), .Z(n13759) );
  NANDN U14582 ( .A(n13759), .B(n13760), .Z(n13403) );
  AND U14583 ( .A(n13404), .B(n13403), .Z(n13407) );
  NANDN U14584 ( .A(n13407), .B(n13408), .Z(n13410) );
  NAND U14585 ( .A(a[7]), .B(b[26]), .Z(n13767) );
  NANDN U14586 ( .A(n13767), .B(n13768), .Z(n13409) );
  AND U14587 ( .A(n13410), .B(n13409), .Z(n13414) );
  NANDN U14588 ( .A(n13413), .B(n13414), .Z(n13416) );
  XOR U14589 ( .A(n13412), .B(n13411), .Z(n13725) );
  NANDN U14590 ( .A(n13725), .B(n13726), .Z(n13415) );
  AND U14591 ( .A(n13416), .B(n13415), .Z(n13420) );
  XOR U14592 ( .A(n13418), .B(n13417), .Z(n13419) );
  NAND U14593 ( .A(n13420), .B(n13419), .Z(n13422) );
  NAND U14594 ( .A(a[9]), .B(b[26]), .Z(n13775) );
  XOR U14595 ( .A(n13420), .B(n13419), .Z(n13776) );
  NANDN U14596 ( .A(n13775), .B(n13776), .Z(n13421) );
  AND U14597 ( .A(n13422), .B(n13421), .Z(n13425) );
  AND U14598 ( .A(a[10]), .B(b[26]), .Z(n13426) );
  NANDN U14599 ( .A(n13425), .B(n13426), .Z(n13428) );
  NAND U14600 ( .A(n13782), .B(n13781), .Z(n13427) );
  AND U14601 ( .A(n13428), .B(n13427), .Z(n13431) );
  XOR U14602 ( .A(n13430), .B(n13429), .Z(n13432) );
  NANDN U14603 ( .A(n13431), .B(n13432), .Z(n13434) );
  AND U14604 ( .A(a[11]), .B(b[26]), .Z(n13788) );
  NAND U14605 ( .A(n13788), .B(n13787), .Z(n13433) );
  AND U14606 ( .A(n13434), .B(n13433), .Z(n13721) );
  AND U14607 ( .A(a[12]), .B(b[26]), .Z(n13435) );
  IV U14608 ( .A(n13435), .Z(n13722) );
  OR U14609 ( .A(n13721), .B(n13722), .Z(n13441) );
  ANDN U14610 ( .B(n13721), .A(n13435), .Z(n13439) );
  OR U14611 ( .A(n13439), .B(n13724), .Z(n13440) );
  AND U14612 ( .A(n13441), .B(n13440), .Z(n13794) );
  XOR U14613 ( .A(n13443), .B(n13442), .Z(n13444) );
  IV U14614 ( .A(n13444), .Z(n13793) );
  OR U14615 ( .A(n13794), .B(n13793), .Z(n13447) );
  ANDN U14616 ( .B(n13794), .A(n13444), .Z(n13445) );
  NAND U14617 ( .A(a[13]), .B(b[26]), .Z(n13796) );
  OR U14618 ( .A(n13445), .B(n13796), .Z(n13446) );
  AND U14619 ( .A(n13447), .B(n13446), .Z(n13452) );
  AND U14620 ( .A(a[14]), .B(b[26]), .Z(n13453) );
  NANDN U14621 ( .A(n13452), .B(n13453), .Z(n13455) );
  XNOR U14622 ( .A(n13449), .B(n13448), .Z(n13450) );
  XOR U14623 ( .A(n13451), .B(n13450), .Z(n13797) );
  XNOR U14624 ( .A(n13453), .B(n13452), .Z(n13798) );
  NANDN U14625 ( .A(n13797), .B(n13798), .Z(n13454) );
  NAND U14626 ( .A(n13455), .B(n13454), .Z(n13806) );
  NAND U14627 ( .A(a[15]), .B(b[26]), .Z(n13808) );
  AND U14628 ( .A(a[16]), .B(b[26]), .Z(n13457) );
  NANDN U14629 ( .A(n13456), .B(n13457), .Z(n13463) );
  XNOR U14630 ( .A(n13457), .B(n13456), .Z(n13720) );
  XNOR U14631 ( .A(n13459), .B(n13458), .Z(n13460) );
  XNOR U14632 ( .A(n13461), .B(n13460), .Z(n13719) );
  NAND U14633 ( .A(n13720), .B(n13719), .Z(n13462) );
  NAND U14634 ( .A(n13463), .B(n13462), .Z(n13812) );
  NAND U14635 ( .A(a[17]), .B(b[26]), .Z(n13814) );
  AND U14636 ( .A(a[18]), .B(b[26]), .Z(n13469) );
  NANDN U14637 ( .A(n13468), .B(n13469), .Z(n13471) );
  XNOR U14638 ( .A(n13465), .B(n13464), .Z(n13466) );
  XNOR U14639 ( .A(n13467), .B(n13466), .Z(n13718) );
  XNOR U14640 ( .A(n13469), .B(n13468), .Z(n13717) );
  NAND U14641 ( .A(n13718), .B(n13717), .Z(n13470) );
  NAND U14642 ( .A(n13471), .B(n13470), .Z(n13820) );
  NAND U14643 ( .A(a[19]), .B(b[26]), .Z(n13822) );
  AND U14644 ( .A(a[20]), .B(b[26]), .Z(n13473) );
  NANDN U14645 ( .A(n13472), .B(n13473), .Z(n13479) );
  XNOR U14646 ( .A(n13473), .B(n13472), .Z(n13828) );
  XNOR U14647 ( .A(n13475), .B(n13474), .Z(n13476) );
  XNOR U14648 ( .A(n13477), .B(n13476), .Z(n13827) );
  NAND U14649 ( .A(n13828), .B(n13827), .Z(n13478) );
  NAND U14650 ( .A(n13479), .B(n13478), .Z(n13834) );
  NAND U14651 ( .A(a[21]), .B(b[26]), .Z(n13836) );
  AND U14652 ( .A(a[22]), .B(b[26]), .Z(n13481) );
  NANDN U14653 ( .A(n13480), .B(n13481), .Z(n13486) );
  XNOR U14654 ( .A(n13481), .B(n13480), .Z(n13716) );
  NAND U14655 ( .A(n13716), .B(n13715), .Z(n13485) );
  AND U14656 ( .A(n13486), .B(n13485), .Z(n13844) );
  XOR U14657 ( .A(n13488), .B(n13487), .Z(n13489) );
  IV U14658 ( .A(n13489), .Z(n13845) );
  NAND U14659 ( .A(a[23]), .B(b[26]), .Z(n13843) );
  NANDN U14660 ( .A(n13494), .B(n13495), .Z(n13497) );
  XNOR U14661 ( .A(n13491), .B(n13490), .Z(n13492) );
  XNOR U14662 ( .A(n13493), .B(n13492), .Z(n13714) );
  NAND U14663 ( .A(n13714), .B(n13713), .Z(n13496) );
  NAND U14664 ( .A(n13497), .B(n13496), .Z(n13849) );
  NAND U14665 ( .A(a[25]), .B(b[26]), .Z(n13851) );
  NANDN U14666 ( .A(n13498), .B(n13499), .Z(n13504) );
  NAND U14667 ( .A(n13711), .B(n13712), .Z(n13503) );
  AND U14668 ( .A(n13504), .B(n13503), .Z(n13856) );
  XOR U14669 ( .A(n13506), .B(n13505), .Z(n13507) );
  IV U14670 ( .A(n13507), .Z(n13857) );
  NAND U14671 ( .A(a[27]), .B(b[26]), .Z(n13859) );
  NANDN U14672 ( .A(n13512), .B(n13513), .Z(n13515) );
  XOR U14673 ( .A(n13509), .B(n13508), .Z(n13510) );
  XOR U14674 ( .A(n13511), .B(n13510), .Z(n13709) );
  NANDN U14675 ( .A(n13709), .B(n13710), .Z(n13514) );
  NAND U14676 ( .A(n13515), .B(n13514), .Z(n13868) );
  NAND U14677 ( .A(a[29]), .B(b[26]), .Z(n13866) );
  NANDN U14678 ( .A(n13516), .B(n13517), .Z(n13522) );
  NAND U14679 ( .A(n13872), .B(n13871), .Z(n13521) );
  NAND U14680 ( .A(n13522), .B(n13521), .Z(n13879) );
  NAND U14681 ( .A(a[31]), .B(b[26]), .Z(n13881) );
  NANDN U14682 ( .A(n13527), .B(n13528), .Z(n13530) );
  XOR U14683 ( .A(n13524), .B(n13523), .Z(n13525) );
  XNOR U14684 ( .A(n13526), .B(n13525), .Z(n13885) );
  NAND U14685 ( .A(n13885), .B(n13884), .Z(n13529) );
  NAND U14686 ( .A(n13530), .B(n13529), .Z(n13888) );
  XOR U14687 ( .A(n13532), .B(n13531), .Z(n13887) );
  AND U14688 ( .A(a[33]), .B(b[26]), .Z(n13886) );
  AND U14689 ( .A(a[34]), .B(b[26]), .Z(n13538) );
  NANDN U14690 ( .A(n13537), .B(n13538), .Z(n13540) );
  XNOR U14691 ( .A(n13534), .B(n13533), .Z(n13535) );
  XNOR U14692 ( .A(n13536), .B(n13535), .Z(n13708) );
  XNOR U14693 ( .A(n13538), .B(n13537), .Z(n13707) );
  NAND U14694 ( .A(n13708), .B(n13707), .Z(n13539) );
  NAND U14695 ( .A(n13540), .B(n13539), .Z(n13894) );
  NAND U14696 ( .A(a[35]), .B(b[26]), .Z(n13896) );
  AND U14697 ( .A(a[36]), .B(b[26]), .Z(n13546) );
  NANDN U14698 ( .A(n13545), .B(n13546), .Z(n13548) );
  XNOR U14699 ( .A(n13542), .B(n13541), .Z(n13543) );
  XNOR U14700 ( .A(n13544), .B(n13543), .Z(n13706) );
  XNOR U14701 ( .A(n13546), .B(n13545), .Z(n13705) );
  NAND U14702 ( .A(n13706), .B(n13705), .Z(n13547) );
  NAND U14703 ( .A(n13548), .B(n13547), .Z(n13905) );
  AND U14704 ( .A(a[37]), .B(b[26]), .Z(n13903) );
  AND U14705 ( .A(a[38]), .B(b[26]), .Z(n13549) );
  NANDN U14706 ( .A(n13550), .B(n13549), .Z(n13554) );
  XOR U14707 ( .A(n13550), .B(n13549), .Z(n13908) );
  XNOR U14708 ( .A(n13552), .B(n13551), .Z(n13909) );
  NANDN U14709 ( .A(n13908), .B(n13909), .Z(n13553) );
  AND U14710 ( .A(n13554), .B(n13553), .Z(n13556) );
  AND U14711 ( .A(a[39]), .B(b[26]), .Z(n13555) );
  NANDN U14712 ( .A(n13556), .B(n13555), .Z(n13562) );
  XOR U14713 ( .A(n13556), .B(n13555), .Z(n13703) );
  XOR U14714 ( .A(n13558), .B(n13557), .Z(n13559) );
  XNOR U14715 ( .A(n13560), .B(n13559), .Z(n13704) );
  NANDN U14716 ( .A(n13703), .B(n13704), .Z(n13561) );
  AND U14717 ( .A(n13562), .B(n13561), .Z(n13915) );
  XNOR U14718 ( .A(n13564), .B(n13563), .Z(n13914) );
  NANDN U14719 ( .A(n13915), .B(n13914), .Z(n13565) );
  AND U14720 ( .A(n13566), .B(n13565), .Z(n13570) );
  XOR U14721 ( .A(n13568), .B(n13567), .Z(n13569) );
  NANDN U14722 ( .A(n13570), .B(n13569), .Z(n13572) );
  NAND U14723 ( .A(a[41]), .B(b[26]), .Z(n13920) );
  XNOR U14724 ( .A(n13570), .B(n13569), .Z(n13921) );
  NANDN U14725 ( .A(n13920), .B(n13921), .Z(n13571) );
  AND U14726 ( .A(n13572), .B(n13571), .Z(n13929) );
  XOR U14727 ( .A(n13574), .B(n13573), .Z(n13928) );
  XOR U14728 ( .A(n13576), .B(n13575), .Z(n13577) );
  NANDN U14729 ( .A(n13578), .B(n13577), .Z(n13580) );
  NAND U14730 ( .A(a[43]), .B(b[26]), .Z(n13932) );
  XNOR U14731 ( .A(n13578), .B(n13577), .Z(n13933) );
  NANDN U14732 ( .A(n13932), .B(n13933), .Z(n13579) );
  AND U14733 ( .A(n13580), .B(n13579), .Z(n13941) );
  XOR U14734 ( .A(n13582), .B(n13581), .Z(n13940) );
  XOR U14735 ( .A(n13584), .B(n13583), .Z(n13585) );
  NANDN U14736 ( .A(n13586), .B(n13585), .Z(n13588) );
  NAND U14737 ( .A(a[45]), .B(b[26]), .Z(n13944) );
  XNOR U14738 ( .A(n13586), .B(n13585), .Z(n13945) );
  NANDN U14739 ( .A(n13944), .B(n13945), .Z(n13587) );
  AND U14740 ( .A(n13588), .B(n13587), .Z(n13953) );
  XOR U14741 ( .A(n13590), .B(n13589), .Z(n13952) );
  XOR U14742 ( .A(n13592), .B(n13591), .Z(n13593) );
  NANDN U14743 ( .A(n13594), .B(n13593), .Z(n13596) );
  NAND U14744 ( .A(a[47]), .B(b[26]), .Z(n13956) );
  XNOR U14745 ( .A(n13594), .B(n13593), .Z(n13957) );
  NANDN U14746 ( .A(n13956), .B(n13957), .Z(n13595) );
  AND U14747 ( .A(n13596), .B(n13595), .Z(n13965) );
  XOR U14748 ( .A(n13598), .B(n13597), .Z(n13964) );
  XOR U14749 ( .A(n13600), .B(n13599), .Z(n13601) );
  NANDN U14750 ( .A(n13602), .B(n13601), .Z(n13604) );
  NAND U14751 ( .A(a[49]), .B(b[26]), .Z(n13968) );
  XNOR U14752 ( .A(n13602), .B(n13601), .Z(n13969) );
  NANDN U14753 ( .A(n13968), .B(n13969), .Z(n13603) );
  AND U14754 ( .A(n13604), .B(n13603), .Z(n13977) );
  XOR U14755 ( .A(n13606), .B(n13605), .Z(n13976) );
  XOR U14756 ( .A(n13608), .B(n13607), .Z(n13609) );
  NANDN U14757 ( .A(n13610), .B(n13609), .Z(n13612) );
  NAND U14758 ( .A(a[51]), .B(b[26]), .Z(n13980) );
  XNOR U14759 ( .A(n13610), .B(n13609), .Z(n13981) );
  NANDN U14760 ( .A(n13980), .B(n13981), .Z(n13611) );
  AND U14761 ( .A(n13612), .B(n13611), .Z(n13989) );
  XOR U14762 ( .A(n13614), .B(n13613), .Z(n13988) );
  XOR U14763 ( .A(n13616), .B(n13615), .Z(n13617) );
  NANDN U14764 ( .A(n13618), .B(n13617), .Z(n13620) );
  NAND U14765 ( .A(a[53]), .B(b[26]), .Z(n13992) );
  XNOR U14766 ( .A(n13618), .B(n13617), .Z(n13993) );
  NANDN U14767 ( .A(n13992), .B(n13993), .Z(n13619) );
  AND U14768 ( .A(n13620), .B(n13619), .Z(n14001) );
  XOR U14769 ( .A(n13622), .B(n13621), .Z(n14000) );
  XOR U14770 ( .A(n13624), .B(n13623), .Z(n13625) );
  NANDN U14771 ( .A(n13626), .B(n13625), .Z(n13628) );
  NAND U14772 ( .A(a[55]), .B(b[26]), .Z(n14004) );
  XNOR U14773 ( .A(n13626), .B(n13625), .Z(n14005) );
  NANDN U14774 ( .A(n14004), .B(n14005), .Z(n13627) );
  AND U14775 ( .A(n13628), .B(n13627), .Z(n14013) );
  XOR U14776 ( .A(n13630), .B(n13629), .Z(n14012) );
  XOR U14777 ( .A(n13632), .B(n13631), .Z(n13633) );
  NANDN U14778 ( .A(n13634), .B(n13633), .Z(n13636) );
  NAND U14779 ( .A(a[57]), .B(b[26]), .Z(n14016) );
  XNOR U14780 ( .A(n13634), .B(n13633), .Z(n14017) );
  NANDN U14781 ( .A(n14016), .B(n14017), .Z(n13635) );
  AND U14782 ( .A(n13636), .B(n13635), .Z(n14025) );
  XOR U14783 ( .A(n13638), .B(n13637), .Z(n14024) );
  XOR U14784 ( .A(n13640), .B(n13639), .Z(n13641) );
  NANDN U14785 ( .A(n13642), .B(n13641), .Z(n13644) );
  NAND U14786 ( .A(a[59]), .B(b[26]), .Z(n14028) );
  XNOR U14787 ( .A(n13642), .B(n13641), .Z(n14029) );
  NANDN U14788 ( .A(n14028), .B(n14029), .Z(n13643) );
  AND U14789 ( .A(n13644), .B(n13643), .Z(n14035) );
  XOR U14790 ( .A(n13646), .B(n13645), .Z(n14034) );
  XOR U14791 ( .A(n13648), .B(n13647), .Z(n13649) );
  NANDN U14792 ( .A(n13650), .B(n13649), .Z(n13652) );
  NAND U14793 ( .A(a[61]), .B(b[26]), .Z(n14040) );
  XNOR U14794 ( .A(n13650), .B(n13649), .Z(n14041) );
  NANDN U14795 ( .A(n14040), .B(n14041), .Z(n13651) );
  AND U14796 ( .A(n13652), .B(n13651), .Z(n14045) );
  XOR U14797 ( .A(n13654), .B(n13653), .Z(n14044) );
  NANDN U14798 ( .A(n13656), .B(n13655), .Z(n13660) );
  NANDN U14799 ( .A(n13658), .B(n13657), .Z(n13659) );
  AND U14800 ( .A(n13660), .B(n13659), .Z(n13681) );
  NAND U14801 ( .A(a[62]), .B(b[27]), .Z(n13682) );
  XNOR U14802 ( .A(n13681), .B(n13682), .Z(n13683) );
  NAND U14803 ( .A(n13662), .B(n13661), .Z(n13666) );
  NANDN U14804 ( .A(n13664), .B(n13663), .Z(n13665) );
  NAND U14805 ( .A(n13666), .B(n13665), .Z(n13674) );
  XNOR U14806 ( .A(n13668), .B(n13667), .Z(n13673) );
  XOR U14807 ( .A(n13674), .B(n13673), .Z(n13675) );
  AND U14808 ( .A(a[61]), .B(b[28]), .Z(n13676) );
  XOR U14809 ( .A(n13675), .B(n13676), .Z(n13684) );
  XOR U14810 ( .A(n13683), .B(n13684), .Z(n13669) );
  NANDN U14811 ( .A(n13670), .B(n13669), .Z(n13672) );
  NAND U14812 ( .A(a[63]), .B(b[26]), .Z(n14048) );
  XNOR U14813 ( .A(n13670), .B(n13669), .Z(n14049) );
  NANDN U14814 ( .A(n14048), .B(n14049), .Z(n13671) );
  NAND U14815 ( .A(n13672), .B(n13671), .Z(n13701) );
  NAND U14816 ( .A(n13674), .B(n13673), .Z(n13678) );
  NAND U14817 ( .A(n13676), .B(n13675), .Z(n13677) );
  NAND U14818 ( .A(n13678), .B(n13677), .Z(n13695) );
  XOR U14819 ( .A(n13680), .B(n13679), .Z(n13693) );
  AND U14820 ( .A(a[62]), .B(b[28]), .Z(n13694) );
  XNOR U14821 ( .A(n13693), .B(n13694), .Z(n13696) );
  AND U14822 ( .A(a[63]), .B(b[27]), .Z(n13688) );
  NANDN U14823 ( .A(n13682), .B(n13681), .Z(n13686) );
  NAND U14824 ( .A(n13684), .B(n13683), .Z(n13685) );
  AND U14825 ( .A(n13686), .B(n13685), .Z(n13687) );
  XOR U14826 ( .A(n13689), .B(n13690), .Z(n13702) );
  NANDN U14827 ( .A(n13688), .B(n13687), .Z(n13692) );
  NAND U14828 ( .A(n13690), .B(n13689), .Z(n13691) );
  AND U14829 ( .A(n13692), .B(n13691), .Z(n22521) );
  NAND U14830 ( .A(n13694), .B(n13693), .Z(n13698) );
  NANDN U14831 ( .A(n13696), .B(n13695), .Z(n13697) );
  NAND U14832 ( .A(n13698), .B(n13697), .Z(n22524) );
  XNOR U14833 ( .A(n13700), .B(n13699), .Z(n22525) );
  XOR U14834 ( .A(n22524), .B(n22525), .Z(n22527) );
  AND U14835 ( .A(a[63]), .B(b[28]), .Z(n22526) );
  XOR U14836 ( .A(n22527), .B(n22526), .Z(n22520) );
  XOR U14837 ( .A(n22521), .B(n22520), .Z(n24766) );
  XOR U14838 ( .A(n13702), .B(n13701), .Z(n24760) );
  AND U14839 ( .A(a[63]), .B(b[25]), .Z(n14047) );
  NAND U14840 ( .A(a[62]), .B(b[25]), .Z(n14038) );
  AND U14841 ( .A(a[61]), .B(b[25]), .Z(n14037) );
  NAND U14842 ( .A(a[60]), .B(b[25]), .Z(n14030) );
  AND U14843 ( .A(a[59]), .B(b[25]), .Z(n14023) );
  NAND U14844 ( .A(a[58]), .B(b[25]), .Z(n14018) );
  AND U14845 ( .A(a[57]), .B(b[25]), .Z(n14011) );
  NAND U14846 ( .A(a[56]), .B(b[25]), .Z(n14006) );
  AND U14847 ( .A(a[55]), .B(b[25]), .Z(n13999) );
  NAND U14848 ( .A(a[54]), .B(b[25]), .Z(n13994) );
  AND U14849 ( .A(a[53]), .B(b[25]), .Z(n13987) );
  NAND U14850 ( .A(a[52]), .B(b[25]), .Z(n13982) );
  AND U14851 ( .A(a[51]), .B(b[25]), .Z(n13975) );
  NAND U14852 ( .A(a[50]), .B(b[25]), .Z(n13970) );
  AND U14853 ( .A(a[49]), .B(b[25]), .Z(n13963) );
  NAND U14854 ( .A(a[48]), .B(b[25]), .Z(n13958) );
  AND U14855 ( .A(a[47]), .B(b[25]), .Z(n13951) );
  NAND U14856 ( .A(a[46]), .B(b[25]), .Z(n13946) );
  AND U14857 ( .A(a[45]), .B(b[25]), .Z(n13939) );
  NAND U14858 ( .A(a[44]), .B(b[25]), .Z(n13934) );
  AND U14859 ( .A(a[43]), .B(b[25]), .Z(n13927) );
  NAND U14860 ( .A(a[41]), .B(b[25]), .Z(n13916) );
  AND U14861 ( .A(a[40]), .B(b[25]), .Z(n14285) );
  XOR U14862 ( .A(n13704), .B(n13703), .Z(n14284) );
  AND U14863 ( .A(a[38]), .B(b[25]), .Z(n13901) );
  XNOR U14864 ( .A(n13706), .B(n13705), .Z(n14270) );
  XNOR U14865 ( .A(n13708), .B(n13707), .Z(n14262) );
  NAND U14866 ( .A(a[34]), .B(b[25]), .Z(n13889) );
  AND U14867 ( .A(a[30]), .B(b[25]), .Z(n13864) );
  XOR U14868 ( .A(n13712), .B(n13711), .Z(n14229) );
  XNOR U14869 ( .A(n13714), .B(n13713), .Z(n14218) );
  XNOR U14870 ( .A(n13716), .B(n13715), .Z(n14210) );
  XNOR U14871 ( .A(n13718), .B(n13717), .Z(n14196) );
  XNOR U14872 ( .A(n13720), .B(n13719), .Z(n14186) );
  NAND U14873 ( .A(a[14]), .B(b[25]), .Z(n14174) );
  XOR U14874 ( .A(n13722), .B(n13721), .Z(n13723) );
  XOR U14875 ( .A(n13724), .B(n13723), .Z(n14168) );
  AND U14876 ( .A(a[4]), .B(b[25]), .Z(n13743) );
  AND U14877 ( .A(b[25]), .B(a[0]), .Z(n14414) );
  AND U14878 ( .A(a[1]), .B(b[26]), .Z(n13730) );
  AND U14879 ( .A(n14414), .B(n13730), .Z(n13727) );
  NAND U14880 ( .A(a[2]), .B(n13727), .Z(n13734) );
  NAND U14881 ( .A(b[26]), .B(a[1]), .Z(n13728) );
  XOR U14882 ( .A(n13729), .B(n13728), .Z(n14102) );
  NAND U14883 ( .A(n13730), .B(a[0]), .Z(n13731) );
  XNOR U14884 ( .A(a[2]), .B(n13731), .Z(n13732) );
  AND U14885 ( .A(b[25]), .B(n13732), .Z(n14103) );
  NANDN U14886 ( .A(n14102), .B(n14103), .Z(n13733) );
  AND U14887 ( .A(n13734), .B(n13733), .Z(n13737) );
  NANDN U14888 ( .A(n13737), .B(n13738), .Z(n13740) );
  NAND U14889 ( .A(a[3]), .B(b[25]), .Z(n14110) );
  NANDN U14890 ( .A(n14110), .B(n14111), .Z(n13739) );
  AND U14891 ( .A(n13740), .B(n13739), .Z(n13744) );
  NANDN U14892 ( .A(n13743), .B(n13744), .Z(n13746) );
  XOR U14893 ( .A(n13742), .B(n13741), .Z(n14092) );
  NANDN U14894 ( .A(n14092), .B(n14093), .Z(n13745) );
  AND U14895 ( .A(n13746), .B(n13745), .Z(n13750) );
  XOR U14896 ( .A(n13748), .B(n13747), .Z(n13749) );
  NAND U14897 ( .A(n13750), .B(n13749), .Z(n13752) );
  NAND U14898 ( .A(a[5]), .B(b[25]), .Z(n14118) );
  XOR U14899 ( .A(n13750), .B(n13749), .Z(n14119) );
  NANDN U14900 ( .A(n14118), .B(n14119), .Z(n13751) );
  AND U14901 ( .A(n13752), .B(n13751), .Z(n13755) );
  NANDN U14902 ( .A(n13755), .B(n13756), .Z(n13758) );
  NAND U14903 ( .A(a[6]), .B(b[25]), .Z(n14124) );
  NANDN U14904 ( .A(n14124), .B(n14125), .Z(n13757) );
  AND U14905 ( .A(n13758), .B(n13757), .Z(n13761) );
  NANDN U14906 ( .A(n13761), .B(n13762), .Z(n13764) );
  AND U14907 ( .A(a[7]), .B(b[25]), .Z(n14130) );
  NAND U14908 ( .A(n14131), .B(n14130), .Z(n13763) );
  AND U14909 ( .A(n13764), .B(n13763), .Z(n13765) );
  AND U14910 ( .A(a[8]), .B(b[25]), .Z(n13766) );
  NANDN U14911 ( .A(n13765), .B(n13766), .Z(n13770) );
  NAND U14912 ( .A(n14137), .B(n14136), .Z(n13769) );
  NAND U14913 ( .A(n13770), .B(n13769), .Z(n13771) );
  NAND U14914 ( .A(n13772), .B(n13771), .Z(n13774) );
  NAND U14915 ( .A(a[9]), .B(b[25]), .Z(n14144) );
  XOR U14916 ( .A(n13772), .B(n13771), .Z(n14145) );
  NANDN U14917 ( .A(n14144), .B(n14145), .Z(n13773) );
  AND U14918 ( .A(n13774), .B(n13773), .Z(n13777) );
  AND U14919 ( .A(a[10]), .B(b[25]), .Z(n13778) );
  NANDN U14920 ( .A(n13777), .B(n13778), .Z(n13780) );
  NAND U14921 ( .A(n14149), .B(n14148), .Z(n13779) );
  AND U14922 ( .A(n13780), .B(n13779), .Z(n13783) );
  XOR U14923 ( .A(n13782), .B(n13781), .Z(n13784) );
  NANDN U14924 ( .A(n13783), .B(n13784), .Z(n13786) );
  NAND U14925 ( .A(a[11]), .B(b[25]), .Z(n14156) );
  NANDN U14926 ( .A(n14156), .B(n14157), .Z(n13785) );
  AND U14927 ( .A(n13786), .B(n13785), .Z(n13789) );
  AND U14928 ( .A(a[12]), .B(b[25]), .Z(n13790) );
  NANDN U14929 ( .A(n13789), .B(n13790), .Z(n13792) );
  XOR U14930 ( .A(n13788), .B(n13787), .Z(n14161) );
  NAND U14931 ( .A(n14161), .B(n14160), .Z(n13791) );
  NAND U14932 ( .A(n13792), .B(n13791), .Z(n14169) );
  AND U14933 ( .A(a[13]), .B(b[25]), .Z(n14167) );
  XOR U14934 ( .A(n13794), .B(n13793), .Z(n13795) );
  XOR U14935 ( .A(n13796), .B(n13795), .Z(n14173) );
  NAND U14936 ( .A(n13800), .B(n13799), .Z(n13802) );
  AND U14937 ( .A(a[15]), .B(b[25]), .Z(n14181) );
  XOR U14938 ( .A(n13800), .B(n13799), .Z(n14180) );
  NAND U14939 ( .A(n14181), .B(n14180), .Z(n13801) );
  AND U14940 ( .A(n13802), .B(n13801), .Z(n13803) );
  AND U14941 ( .A(a[16]), .B(b[25]), .Z(n13804) );
  NANDN U14942 ( .A(n13803), .B(n13804), .Z(n13810) );
  XNOR U14943 ( .A(n13806), .B(n13805), .Z(n13807) );
  XNOR U14944 ( .A(n13808), .B(n13807), .Z(n14090) );
  NAND U14945 ( .A(n14091), .B(n14090), .Z(n13809) );
  NAND U14946 ( .A(n13810), .B(n13809), .Z(n14187) );
  NAND U14947 ( .A(a[17]), .B(b[25]), .Z(n14189) );
  AND U14948 ( .A(a[18]), .B(b[25]), .Z(n13815) );
  NANDN U14949 ( .A(n13816), .B(n13815), .Z(n13818) );
  XNOR U14950 ( .A(n13812), .B(n13811), .Z(n13813) );
  XNOR U14951 ( .A(n13814), .B(n13813), .Z(n14089) );
  XNOR U14952 ( .A(n13816), .B(n13815), .Z(n14088) );
  NAND U14953 ( .A(n14089), .B(n14088), .Z(n13817) );
  NAND U14954 ( .A(n13818), .B(n13817), .Z(n14197) );
  NAND U14955 ( .A(a[19]), .B(b[25]), .Z(n14199) );
  AND U14956 ( .A(a[20]), .B(b[25]), .Z(n13823) );
  NANDN U14957 ( .A(n13824), .B(n13823), .Z(n13826) );
  XNOR U14958 ( .A(n13820), .B(n13819), .Z(n13821) );
  XNOR U14959 ( .A(n13822), .B(n13821), .Z(n14087) );
  XNOR U14960 ( .A(n13824), .B(n13823), .Z(n14086) );
  NAND U14961 ( .A(n14087), .B(n14086), .Z(n13825) );
  AND U14962 ( .A(n13826), .B(n13825), .Z(n14202) );
  XOR U14963 ( .A(n13828), .B(n13827), .Z(n13829) );
  IV U14964 ( .A(n13829), .Z(n14203) );
  OR U14965 ( .A(n14202), .B(n14203), .Z(n13832) );
  ANDN U14966 ( .B(n14202), .A(n13829), .Z(n13830) );
  NAND U14967 ( .A(a[21]), .B(b[25]), .Z(n14205) );
  OR U14968 ( .A(n13830), .B(n14205), .Z(n13831) );
  AND U14969 ( .A(n13832), .B(n13831), .Z(n13838) );
  AND U14970 ( .A(a[22]), .B(b[25]), .Z(n13837) );
  NANDN U14971 ( .A(n13838), .B(n13837), .Z(n13840) );
  XNOR U14972 ( .A(n13834), .B(n13833), .Z(n13835) );
  XOR U14973 ( .A(n13836), .B(n13835), .Z(n14084) );
  XNOR U14974 ( .A(n13838), .B(n13837), .Z(n14085) );
  NANDN U14975 ( .A(n14084), .B(n14085), .Z(n13839) );
  NAND U14976 ( .A(n13840), .B(n13839), .Z(n14211) );
  NAND U14977 ( .A(a[23]), .B(b[25]), .Z(n14213) );
  AND U14978 ( .A(a[24]), .B(b[25]), .Z(n13841) );
  NANDN U14979 ( .A(n13842), .B(n13841), .Z(n13847) );
  XOR U14980 ( .A(n13842), .B(n13841), .Z(n14082) );
  NANDN U14981 ( .A(n14082), .B(n14083), .Z(n13846) );
  NAND U14982 ( .A(n13847), .B(n13846), .Z(n14219) );
  NAND U14983 ( .A(a[25]), .B(b[25]), .Z(n14221) );
  AND U14984 ( .A(a[26]), .B(b[25]), .Z(n13852) );
  NANDN U14985 ( .A(n13853), .B(n13852), .Z(n13855) );
  XNOR U14986 ( .A(n13849), .B(n13848), .Z(n13850) );
  XNOR U14987 ( .A(n13851), .B(n13850), .Z(n14081) );
  XNOR U14988 ( .A(n13853), .B(n13852), .Z(n14080) );
  NAND U14989 ( .A(n14081), .B(n14080), .Z(n13854) );
  NAND U14990 ( .A(n13855), .B(n13854), .Z(n14230) );
  AND U14991 ( .A(a[27]), .B(b[25]), .Z(n14228) );
  AND U14992 ( .A(a[28]), .B(b[25]), .Z(n13860) );
  NANDN U14993 ( .A(n13861), .B(n13860), .Z(n13863) );
  XOR U14994 ( .A(n13857), .B(n13856), .Z(n13858) );
  XNOR U14995 ( .A(n13859), .B(n13858), .Z(n14079) );
  XNOR U14996 ( .A(n13861), .B(n13860), .Z(n14078) );
  NAND U14997 ( .A(n14079), .B(n14078), .Z(n13862) );
  NAND U14998 ( .A(n13863), .B(n13862), .Z(n14234) );
  NAND U14999 ( .A(a[29]), .B(b[25]), .Z(n14236) );
  NANDN U15000 ( .A(n13864), .B(n13865), .Z(n13870) );
  NAND U15001 ( .A(n14076), .B(n14077), .Z(n13869) );
  NAND U15002 ( .A(n13870), .B(n13869), .Z(n14245) );
  XOR U15003 ( .A(n13872), .B(n13871), .Z(n14244) );
  NANDN U15004 ( .A(n14245), .B(n14244), .Z(n13875) );
  ANDN U15005 ( .B(n14245), .A(n14244), .Z(n13873) );
  AND U15006 ( .A(a[31]), .B(b[25]), .Z(n14243) );
  NANDN U15007 ( .A(n13873), .B(n14243), .Z(n13874) );
  AND U15008 ( .A(n13875), .B(n13874), .Z(n13877) );
  AND U15009 ( .A(a[32]), .B(b[25]), .Z(n13876) );
  NANDN U15010 ( .A(n13877), .B(n13876), .Z(n13883) );
  XOR U15011 ( .A(n13877), .B(n13876), .Z(n14248) );
  XNOR U15012 ( .A(n13879), .B(n13878), .Z(n13880) );
  XNOR U15013 ( .A(n13881), .B(n13880), .Z(n14249) );
  NANDN U15014 ( .A(n14248), .B(n14249), .Z(n13882) );
  NAND U15015 ( .A(n13883), .B(n13882), .Z(n14254) );
  XOR U15016 ( .A(n13885), .B(n13884), .Z(n14253) );
  AND U15017 ( .A(a[33]), .B(b[25]), .Z(n14256) );
  NANDN U15018 ( .A(n13889), .B(n13890), .Z(n13892) );
  NAND U15019 ( .A(n14075), .B(n14074), .Z(n13891) );
  NAND U15020 ( .A(n13892), .B(n13891), .Z(n14263) );
  AND U15021 ( .A(a[35]), .B(b[25]), .Z(n14261) );
  AND U15022 ( .A(a[36]), .B(b[25]), .Z(n13897) );
  NANDN U15023 ( .A(n13898), .B(n13897), .Z(n13900) );
  XNOR U15024 ( .A(n13894), .B(n13893), .Z(n13895) );
  XNOR U15025 ( .A(n13896), .B(n13895), .Z(n14267) );
  XNOR U15026 ( .A(n13898), .B(n13897), .Z(n14266) );
  NAND U15027 ( .A(n14267), .B(n14266), .Z(n13899) );
  NAND U15028 ( .A(n13900), .B(n13899), .Z(n14271) );
  NAND U15029 ( .A(a[37]), .B(b[25]), .Z(n14273) );
  NANDN U15030 ( .A(n13901), .B(n13902), .Z(n13907) );
  NAND U15031 ( .A(n14072), .B(n14073), .Z(n13906) );
  AND U15032 ( .A(n13907), .B(n13906), .Z(n13910) );
  XOR U15033 ( .A(n13909), .B(n13908), .Z(n13911) );
  NANDN U15034 ( .A(n13910), .B(n13911), .Z(n13913) );
  NAND U15035 ( .A(a[39]), .B(b[25]), .Z(n14278) );
  NAND U15036 ( .A(n14279), .B(n14278), .Z(n13912) );
  AND U15037 ( .A(n13913), .B(n13912), .Z(n14287) );
  NANDN U15038 ( .A(n13916), .B(n13917), .Z(n13919) );
  XOR U15039 ( .A(n13915), .B(n13914), .Z(n14070) );
  XNOR U15040 ( .A(n13917), .B(n13916), .Z(n14071) );
  NANDN U15041 ( .A(n14070), .B(n14071), .Z(n13918) );
  AND U15042 ( .A(n13919), .B(n13918), .Z(n13923) );
  AND U15043 ( .A(a[42]), .B(b[25]), .Z(n13922) );
  NANDN U15044 ( .A(n13923), .B(n13922), .Z(n13925) );
  XOR U15045 ( .A(n13921), .B(n13920), .Z(n14294) );
  XNOR U15046 ( .A(n13923), .B(n13922), .Z(n14295) );
  NANDN U15047 ( .A(n14294), .B(n14295), .Z(n13924) );
  AND U15048 ( .A(n13925), .B(n13924), .Z(n13926) );
  NANDN U15049 ( .A(n13927), .B(n13926), .Z(n13931) );
  XOR U15050 ( .A(n13927), .B(n13926), .Z(n14068) );
  XOR U15051 ( .A(n13929), .B(n13928), .Z(n14069) );
  NANDN U15052 ( .A(n14068), .B(n14069), .Z(n13930) );
  AND U15053 ( .A(n13931), .B(n13930), .Z(n13935) );
  NANDN U15054 ( .A(n13934), .B(n13935), .Z(n13937) );
  XOR U15055 ( .A(n13933), .B(n13932), .Z(n14302) );
  XNOR U15056 ( .A(n13935), .B(n13934), .Z(n14303) );
  NANDN U15057 ( .A(n14302), .B(n14303), .Z(n13936) );
  AND U15058 ( .A(n13937), .B(n13936), .Z(n13938) );
  NANDN U15059 ( .A(n13939), .B(n13938), .Z(n13943) );
  XOR U15060 ( .A(n13939), .B(n13938), .Z(n14066) );
  XOR U15061 ( .A(n13941), .B(n13940), .Z(n14067) );
  NANDN U15062 ( .A(n14066), .B(n14067), .Z(n13942) );
  AND U15063 ( .A(n13943), .B(n13942), .Z(n13947) );
  NANDN U15064 ( .A(n13946), .B(n13947), .Z(n13949) );
  XOR U15065 ( .A(n13945), .B(n13944), .Z(n14310) );
  XNOR U15066 ( .A(n13947), .B(n13946), .Z(n14311) );
  NANDN U15067 ( .A(n14310), .B(n14311), .Z(n13948) );
  AND U15068 ( .A(n13949), .B(n13948), .Z(n13950) );
  NANDN U15069 ( .A(n13951), .B(n13950), .Z(n13955) );
  XOR U15070 ( .A(n13951), .B(n13950), .Z(n14064) );
  XOR U15071 ( .A(n13953), .B(n13952), .Z(n14065) );
  NANDN U15072 ( .A(n14064), .B(n14065), .Z(n13954) );
  AND U15073 ( .A(n13955), .B(n13954), .Z(n13959) );
  NANDN U15074 ( .A(n13958), .B(n13959), .Z(n13961) );
  XOR U15075 ( .A(n13957), .B(n13956), .Z(n14318) );
  XNOR U15076 ( .A(n13959), .B(n13958), .Z(n14319) );
  NANDN U15077 ( .A(n14318), .B(n14319), .Z(n13960) );
  AND U15078 ( .A(n13961), .B(n13960), .Z(n13962) );
  NANDN U15079 ( .A(n13963), .B(n13962), .Z(n13967) );
  XOR U15080 ( .A(n13963), .B(n13962), .Z(n14062) );
  XOR U15081 ( .A(n13965), .B(n13964), .Z(n14063) );
  NANDN U15082 ( .A(n14062), .B(n14063), .Z(n13966) );
  AND U15083 ( .A(n13967), .B(n13966), .Z(n13971) );
  NANDN U15084 ( .A(n13970), .B(n13971), .Z(n13973) );
  XOR U15085 ( .A(n13969), .B(n13968), .Z(n14326) );
  XNOR U15086 ( .A(n13971), .B(n13970), .Z(n14327) );
  NANDN U15087 ( .A(n14326), .B(n14327), .Z(n13972) );
  AND U15088 ( .A(n13973), .B(n13972), .Z(n13974) );
  NANDN U15089 ( .A(n13975), .B(n13974), .Z(n13979) );
  XOR U15090 ( .A(n13975), .B(n13974), .Z(n14060) );
  XOR U15091 ( .A(n13977), .B(n13976), .Z(n14061) );
  NANDN U15092 ( .A(n14060), .B(n14061), .Z(n13978) );
  AND U15093 ( .A(n13979), .B(n13978), .Z(n13983) );
  NANDN U15094 ( .A(n13982), .B(n13983), .Z(n13985) );
  XOR U15095 ( .A(n13981), .B(n13980), .Z(n14334) );
  XNOR U15096 ( .A(n13983), .B(n13982), .Z(n14335) );
  NANDN U15097 ( .A(n14334), .B(n14335), .Z(n13984) );
  AND U15098 ( .A(n13985), .B(n13984), .Z(n13986) );
  NANDN U15099 ( .A(n13987), .B(n13986), .Z(n13991) );
  XOR U15100 ( .A(n13987), .B(n13986), .Z(n14058) );
  XOR U15101 ( .A(n13989), .B(n13988), .Z(n14059) );
  NANDN U15102 ( .A(n14058), .B(n14059), .Z(n13990) );
  AND U15103 ( .A(n13991), .B(n13990), .Z(n13995) );
  NANDN U15104 ( .A(n13994), .B(n13995), .Z(n13997) );
  XOR U15105 ( .A(n13993), .B(n13992), .Z(n14342) );
  XNOR U15106 ( .A(n13995), .B(n13994), .Z(n14343) );
  NANDN U15107 ( .A(n14342), .B(n14343), .Z(n13996) );
  AND U15108 ( .A(n13997), .B(n13996), .Z(n13998) );
  NANDN U15109 ( .A(n13999), .B(n13998), .Z(n14003) );
  XOR U15110 ( .A(n13999), .B(n13998), .Z(n14056) );
  XOR U15111 ( .A(n14001), .B(n14000), .Z(n14057) );
  NANDN U15112 ( .A(n14056), .B(n14057), .Z(n14002) );
  AND U15113 ( .A(n14003), .B(n14002), .Z(n14007) );
  NANDN U15114 ( .A(n14006), .B(n14007), .Z(n14009) );
  XOR U15115 ( .A(n14005), .B(n14004), .Z(n14350) );
  XNOR U15116 ( .A(n14007), .B(n14006), .Z(n14351) );
  NANDN U15117 ( .A(n14350), .B(n14351), .Z(n14008) );
  AND U15118 ( .A(n14009), .B(n14008), .Z(n14010) );
  NANDN U15119 ( .A(n14011), .B(n14010), .Z(n14015) );
  XOR U15120 ( .A(n14011), .B(n14010), .Z(n14054) );
  XOR U15121 ( .A(n14013), .B(n14012), .Z(n14055) );
  NANDN U15122 ( .A(n14054), .B(n14055), .Z(n14014) );
  AND U15123 ( .A(n14015), .B(n14014), .Z(n14019) );
  NANDN U15124 ( .A(n14018), .B(n14019), .Z(n14021) );
  XOR U15125 ( .A(n14017), .B(n14016), .Z(n14358) );
  XNOR U15126 ( .A(n14019), .B(n14018), .Z(n14359) );
  NANDN U15127 ( .A(n14358), .B(n14359), .Z(n14020) );
  AND U15128 ( .A(n14021), .B(n14020), .Z(n14022) );
  NANDN U15129 ( .A(n14023), .B(n14022), .Z(n14027) );
  XOR U15130 ( .A(n14023), .B(n14022), .Z(n14052) );
  XOR U15131 ( .A(n14025), .B(n14024), .Z(n14053) );
  NANDN U15132 ( .A(n14052), .B(n14053), .Z(n14026) );
  AND U15133 ( .A(n14027), .B(n14026), .Z(n14031) );
  NANDN U15134 ( .A(n14030), .B(n14031), .Z(n14033) );
  XOR U15135 ( .A(n14029), .B(n14028), .Z(n14366) );
  XNOR U15136 ( .A(n14031), .B(n14030), .Z(n14367) );
  NANDN U15137 ( .A(n14366), .B(n14367), .Z(n14032) );
  AND U15138 ( .A(n14033), .B(n14032), .Z(n14036) );
  XOR U15139 ( .A(n14035), .B(n14034), .Z(n14051) );
  XNOR U15140 ( .A(n14037), .B(n14036), .Z(n14050) );
  NANDN U15141 ( .A(n14038), .B(n14039), .Z(n14043) );
  XNOR U15142 ( .A(n14039), .B(n14038), .Z(n14375) );
  XNOR U15143 ( .A(n14041), .B(n14040), .Z(n14374) );
  NAND U15144 ( .A(n14375), .B(n14374), .Z(n14042) );
  AND U15145 ( .A(n14043), .B(n14042), .Z(n14046) );
  XOR U15146 ( .A(n14045), .B(n14044), .Z(n14379) );
  XNOR U15147 ( .A(n14047), .B(n14046), .Z(n14378) );
  XNOR U15148 ( .A(n14049), .B(n14048), .Z(n14380) );
  AND U15149 ( .A(n14381), .B(n14380), .Z(n24762) );
  XOR U15150 ( .A(n14051), .B(n14050), .Z(n14373) );
  XOR U15151 ( .A(n14053), .B(n14052), .Z(n14365) );
  XOR U15152 ( .A(n14055), .B(n14054), .Z(n14357) );
  AND U15153 ( .A(a[58]), .B(b[24]), .Z(n14356) );
  XOR U15154 ( .A(n14057), .B(n14056), .Z(n14349) );
  AND U15155 ( .A(a[56]), .B(b[24]), .Z(n14348) );
  XOR U15156 ( .A(n14059), .B(n14058), .Z(n14341) );
  AND U15157 ( .A(a[54]), .B(b[24]), .Z(n14340) );
  XOR U15158 ( .A(n14061), .B(n14060), .Z(n14333) );
  AND U15159 ( .A(a[52]), .B(b[24]), .Z(n14332) );
  XOR U15160 ( .A(n14063), .B(n14062), .Z(n14325) );
  AND U15161 ( .A(a[50]), .B(b[24]), .Z(n14324) );
  XOR U15162 ( .A(n14065), .B(n14064), .Z(n14317) );
  AND U15163 ( .A(a[48]), .B(b[24]), .Z(n14316) );
  XOR U15164 ( .A(n14067), .B(n14066), .Z(n14309) );
  AND U15165 ( .A(a[46]), .B(b[24]), .Z(n14308) );
  XOR U15166 ( .A(n14069), .B(n14068), .Z(n14301) );
  AND U15167 ( .A(a[44]), .B(b[24]), .Z(n14300) );
  NAND U15168 ( .A(a[42]), .B(b[24]), .Z(n14290) );
  XNOR U15169 ( .A(n14071), .B(n14070), .Z(n14291) );
  NANDN U15170 ( .A(n14290), .B(n14291), .Z(n14293) );
  XOR U15171 ( .A(n14073), .B(n14072), .Z(n14587) );
  AND U15172 ( .A(a[36]), .B(b[24]), .Z(n14259) );
  XNOR U15173 ( .A(n14075), .B(n14074), .Z(n14571) );
  NAND U15174 ( .A(a[34]), .B(b[24]), .Z(n14251) );
  NAND U15175 ( .A(a[32]), .B(b[24]), .Z(n14241) );
  XNOR U15176 ( .A(n14077), .B(n14076), .Z(n14558) );
  AND U15177 ( .A(a[30]), .B(b[24]), .Z(n14237) );
  XNOR U15178 ( .A(n14079), .B(n14078), .Z(n14551) );
  XNOR U15179 ( .A(n14081), .B(n14080), .Z(n14541) );
  XNOR U15180 ( .A(n14087), .B(n14086), .Z(n14519) );
  XNOR U15181 ( .A(n14089), .B(n14088), .Z(n14511) );
  XOR U15182 ( .A(n14091), .B(n14090), .Z(n14182) );
  IV U15183 ( .A(n14182), .Z(n14505) );
  AND U15184 ( .A(a[8]), .B(b[24]), .Z(n14132) );
  AND U15185 ( .A(b[24]), .B(a[0]), .Z(n14784) );
  AND U15186 ( .A(a[1]), .B(b[25]), .Z(n14097) );
  AND U15187 ( .A(n14784), .B(n14097), .Z(n14094) );
  NAND U15188 ( .A(a[2]), .B(n14094), .Z(n14101) );
  NAND U15189 ( .A(b[25]), .B(a[1]), .Z(n14095) );
  XOR U15190 ( .A(n14096), .B(n14095), .Z(n14420) );
  NAND U15191 ( .A(n14097), .B(a[0]), .Z(n14098) );
  XNOR U15192 ( .A(a[2]), .B(n14098), .Z(n14099) );
  AND U15193 ( .A(b[24]), .B(n14099), .Z(n14421) );
  NANDN U15194 ( .A(n14420), .B(n14421), .Z(n14100) );
  AND U15195 ( .A(n14101), .B(n14100), .Z(n14104) );
  NANDN U15196 ( .A(n14104), .B(n14105), .Z(n14107) );
  AND U15197 ( .A(a[3]), .B(b[24]), .Z(n14426) );
  NAND U15198 ( .A(n14427), .B(n14426), .Z(n14106) );
  AND U15199 ( .A(n14107), .B(n14106), .Z(n14108) );
  AND U15200 ( .A(a[4]), .B(b[24]), .Z(n14109) );
  NANDN U15201 ( .A(n14108), .B(n14109), .Z(n14113) );
  NAND U15202 ( .A(n14433), .B(n14432), .Z(n14112) );
  NAND U15203 ( .A(n14113), .B(n14112), .Z(n14114) );
  NAND U15204 ( .A(n14115), .B(n14114), .Z(n14117) );
  NAND U15205 ( .A(a[5]), .B(b[24]), .Z(n14438) );
  XOR U15206 ( .A(n14115), .B(n14114), .Z(n14439) );
  NANDN U15207 ( .A(n14438), .B(n14439), .Z(n14116) );
  AND U15208 ( .A(n14117), .B(n14116), .Z(n14120) );
  NANDN U15209 ( .A(n14120), .B(n14121), .Z(n14123) );
  NAND U15210 ( .A(a[6]), .B(b[24]), .Z(n14444) );
  NANDN U15211 ( .A(n14444), .B(n14445), .Z(n14122) );
  AND U15212 ( .A(n14123), .B(n14122), .Z(n14126) );
  NANDN U15213 ( .A(n14126), .B(n14127), .Z(n14129) );
  NAND U15214 ( .A(a[7]), .B(b[24]), .Z(n14452) );
  NANDN U15215 ( .A(n14452), .B(n14453), .Z(n14128) );
  AND U15216 ( .A(n14129), .B(n14128), .Z(n14133) );
  NANDN U15217 ( .A(n14132), .B(n14133), .Z(n14135) );
  XOR U15218 ( .A(n14131), .B(n14130), .Z(n14410) );
  NANDN U15219 ( .A(n14410), .B(n14411), .Z(n14134) );
  AND U15220 ( .A(n14135), .B(n14134), .Z(n14139) );
  XOR U15221 ( .A(n14137), .B(n14136), .Z(n14138) );
  NAND U15222 ( .A(n14139), .B(n14138), .Z(n14141) );
  NAND U15223 ( .A(a[9]), .B(b[24]), .Z(n14460) );
  XOR U15224 ( .A(n14139), .B(n14138), .Z(n14461) );
  NANDN U15225 ( .A(n14460), .B(n14461), .Z(n14140) );
  AND U15226 ( .A(n14141), .B(n14140), .Z(n14142) );
  AND U15227 ( .A(a[10]), .B(b[24]), .Z(n14143) );
  NANDN U15228 ( .A(n14142), .B(n14143), .Z(n14147) );
  NAND U15229 ( .A(n14467), .B(n14466), .Z(n14146) );
  AND U15230 ( .A(n14147), .B(n14146), .Z(n14150) );
  XOR U15231 ( .A(n14149), .B(n14148), .Z(n14151) );
  NANDN U15232 ( .A(n14150), .B(n14151), .Z(n14153) );
  NAND U15233 ( .A(a[11]), .B(b[24]), .Z(n14472) );
  NANDN U15234 ( .A(n14472), .B(n14473), .Z(n14152) );
  AND U15235 ( .A(n14153), .B(n14152), .Z(n14154) );
  AND U15236 ( .A(a[12]), .B(b[24]), .Z(n14155) );
  NANDN U15237 ( .A(n14154), .B(n14155), .Z(n14159) );
  NAND U15238 ( .A(n14479), .B(n14478), .Z(n14158) );
  AND U15239 ( .A(n14159), .B(n14158), .Z(n14162) );
  XOR U15240 ( .A(n14161), .B(n14160), .Z(n14163) );
  NANDN U15241 ( .A(n14162), .B(n14163), .Z(n14165) );
  NAND U15242 ( .A(a[13]), .B(b[24]), .Z(n14484) );
  NANDN U15243 ( .A(n14484), .B(n14485), .Z(n14164) );
  AND U15244 ( .A(n14165), .B(n14164), .Z(n14490) );
  AND U15245 ( .A(a[14]), .B(b[24]), .Z(n14166) );
  IV U15246 ( .A(n14166), .Z(n14491) );
  OR U15247 ( .A(n14490), .B(n14491), .Z(n14172) );
  ANDN U15248 ( .B(n14490), .A(n14166), .Z(n14170) );
  OR U15249 ( .A(n14170), .B(n14493), .Z(n14171) );
  AND U15250 ( .A(n14172), .B(n14171), .Z(n14177) );
  NANDN U15251 ( .A(n14177), .B(n14176), .Z(n14179) );
  XOR U15252 ( .A(n14177), .B(n14176), .Z(n14498) );
  AND U15253 ( .A(a[15]), .B(b[24]), .Z(n14499) );
  NANDN U15254 ( .A(n14498), .B(n14499), .Z(n14178) );
  NAND U15255 ( .A(n14179), .B(n14178), .Z(n14406) );
  NAND U15256 ( .A(a[16]), .B(b[24]), .Z(n14407) );
  XOR U15257 ( .A(n14181), .B(n14180), .Z(n14409) );
  NANDN U15258 ( .A(n14505), .B(n14506), .Z(n14185) );
  NOR U15259 ( .A(n14182), .B(n14506), .Z(n14183) );
  AND U15260 ( .A(a[17]), .B(b[24]), .Z(n14504) );
  NANDN U15261 ( .A(n14183), .B(n14504), .Z(n14184) );
  AND U15262 ( .A(n14185), .B(n14184), .Z(n14190) );
  AND U15263 ( .A(a[18]), .B(b[24]), .Z(n14191) );
  NANDN U15264 ( .A(n14190), .B(n14191), .Z(n14193) );
  XNOR U15265 ( .A(n14187), .B(n14186), .Z(n14188) );
  XNOR U15266 ( .A(n14189), .B(n14188), .Z(n14405) );
  XNOR U15267 ( .A(n14191), .B(n14190), .Z(n14404) );
  NAND U15268 ( .A(n14405), .B(n14404), .Z(n14192) );
  NAND U15269 ( .A(n14193), .B(n14192), .Z(n14512) );
  NAND U15270 ( .A(a[19]), .B(b[24]), .Z(n14514) );
  AND U15271 ( .A(a[20]), .B(b[24]), .Z(n14195) );
  NANDN U15272 ( .A(n14194), .B(n14195), .Z(n14201) );
  XNOR U15273 ( .A(n14195), .B(n14194), .Z(n14403) );
  XNOR U15274 ( .A(n14197), .B(n14196), .Z(n14198) );
  XNOR U15275 ( .A(n14199), .B(n14198), .Z(n14402) );
  NAND U15276 ( .A(n14403), .B(n14402), .Z(n14200) );
  NAND U15277 ( .A(n14201), .B(n14200), .Z(n14520) );
  NAND U15278 ( .A(a[21]), .B(b[24]), .Z(n14522) );
  AND U15279 ( .A(a[22]), .B(b[24]), .Z(n14207) );
  NANDN U15280 ( .A(n14206), .B(n14207), .Z(n14209) );
  XOR U15281 ( .A(n14203), .B(n14202), .Z(n14204) );
  XNOR U15282 ( .A(n14205), .B(n14204), .Z(n14401) );
  XNOR U15283 ( .A(n14207), .B(n14206), .Z(n14400) );
  NAND U15284 ( .A(n14401), .B(n14400), .Z(n14208) );
  NAND U15285 ( .A(n14209), .B(n14208), .Z(n14529) );
  NAND U15286 ( .A(a[23]), .B(b[24]), .Z(n14527) );
  AND U15287 ( .A(a[24]), .B(b[24]), .Z(n14215) );
  NANDN U15288 ( .A(n14214), .B(n14215), .Z(n14217) );
  XNOR U15289 ( .A(n14211), .B(n14210), .Z(n14212) );
  XNOR U15290 ( .A(n14213), .B(n14212), .Z(n14399) );
  NAND U15291 ( .A(n14399), .B(n14398), .Z(n14216) );
  NAND U15292 ( .A(n14217), .B(n14216), .Z(n14536) );
  NAND U15293 ( .A(a[25]), .B(b[24]), .Z(n14534) );
  AND U15294 ( .A(a[26]), .B(b[24]), .Z(n14223) );
  NANDN U15295 ( .A(n14222), .B(n14223), .Z(n14225) );
  XNOR U15296 ( .A(n14219), .B(n14218), .Z(n14220) );
  XNOR U15297 ( .A(n14221), .B(n14220), .Z(n14397) );
  NAND U15298 ( .A(n14397), .B(n14396), .Z(n14224) );
  NAND U15299 ( .A(n14225), .B(n14224), .Z(n14542) );
  NAND U15300 ( .A(a[27]), .B(b[24]), .Z(n14544) );
  AND U15301 ( .A(a[28]), .B(b[24]), .Z(n14227) );
  NANDN U15302 ( .A(n14226), .B(n14227), .Z(n14232) );
  XNOR U15303 ( .A(n14227), .B(n14226), .Z(n14395) );
  NAND U15304 ( .A(n14395), .B(n14394), .Z(n14231) );
  NAND U15305 ( .A(n14232), .B(n14231), .Z(n14552) );
  NAND U15306 ( .A(a[29]), .B(b[24]), .Z(n14554) );
  NANDN U15307 ( .A(n14237), .B(n14238), .Z(n14240) );
  XOR U15308 ( .A(n14234), .B(n14233), .Z(n14235) );
  XOR U15309 ( .A(n14236), .B(n14235), .Z(n14392) );
  NANDN U15310 ( .A(n14392), .B(n14393), .Z(n14239) );
  NAND U15311 ( .A(n14240), .B(n14239), .Z(n14559) );
  NAND U15312 ( .A(a[31]), .B(b[24]), .Z(n14557) );
  NANDN U15313 ( .A(n14241), .B(n14242), .Z(n14247) );
  NAND U15314 ( .A(n14391), .B(n14390), .Z(n14246) );
  AND U15315 ( .A(n14247), .B(n14246), .Z(n14565) );
  IV U15316 ( .A(n14250), .Z(n14566) );
  NAND U15317 ( .A(a[33]), .B(b[24]), .Z(n14564) );
  NANDN U15318 ( .A(n14251), .B(n14252), .Z(n14258) );
  XOR U15319 ( .A(n14254), .B(n14253), .Z(n14255) );
  XNOR U15320 ( .A(n14256), .B(n14255), .Z(n14388) );
  NAND U15321 ( .A(n14389), .B(n14388), .Z(n14257) );
  NAND U15322 ( .A(n14258), .B(n14257), .Z(n14572) );
  NAND U15323 ( .A(a[35]), .B(b[24]), .Z(n14574) );
  NANDN U15324 ( .A(n14259), .B(n14260), .Z(n14265) );
  NAND U15325 ( .A(n14386), .B(n14387), .Z(n14264) );
  NAND U15326 ( .A(n14265), .B(n14264), .Z(n14581) );
  XOR U15327 ( .A(n14267), .B(n14266), .Z(n14580) );
  AND U15328 ( .A(a[37]), .B(b[24]), .Z(n14579) );
  AND U15329 ( .A(a[38]), .B(b[24]), .Z(n14269) );
  NANDN U15330 ( .A(n14268), .B(n14269), .Z(n14275) );
  XNOR U15331 ( .A(n14269), .B(n14268), .Z(n14385) );
  XNOR U15332 ( .A(n14271), .B(n14270), .Z(n14272) );
  XNOR U15333 ( .A(n14273), .B(n14272), .Z(n14384) );
  NAND U15334 ( .A(n14385), .B(n14384), .Z(n14274) );
  NAND U15335 ( .A(n14275), .B(n14274), .Z(n14588) );
  AND U15336 ( .A(a[39]), .B(b[24]), .Z(n14586) );
  AND U15337 ( .A(a[40]), .B(b[24]), .Z(n14276) );
  NANDN U15338 ( .A(n14277), .B(n14276), .Z(n14281) );
  XOR U15339 ( .A(n14277), .B(n14276), .Z(n14593) );
  XNOR U15340 ( .A(n14279), .B(n14278), .Z(n14594) );
  NANDN U15341 ( .A(n14593), .B(n14594), .Z(n14280) );
  AND U15342 ( .A(n14281), .B(n14280), .Z(n14283) );
  AND U15343 ( .A(a[41]), .B(b[24]), .Z(n14282) );
  NANDN U15344 ( .A(n14283), .B(n14282), .Z(n14289) );
  XOR U15345 ( .A(n14283), .B(n14282), .Z(n14382) );
  XOR U15346 ( .A(n14285), .B(n14284), .Z(n14286) );
  XNOR U15347 ( .A(n14287), .B(n14286), .Z(n14383) );
  NANDN U15348 ( .A(n14382), .B(n14383), .Z(n14288) );
  AND U15349 ( .A(n14289), .B(n14288), .Z(n14600) );
  XNOR U15350 ( .A(n14291), .B(n14290), .Z(n14599) );
  NANDN U15351 ( .A(n14600), .B(n14599), .Z(n14292) );
  AND U15352 ( .A(n14293), .B(n14292), .Z(n14297) );
  XNOR U15353 ( .A(n14295), .B(n14294), .Z(n14296) );
  NANDN U15354 ( .A(n14297), .B(n14296), .Z(n14299) );
  NAND U15355 ( .A(a[43]), .B(b[24]), .Z(n14605) );
  XNOR U15356 ( .A(n14297), .B(n14296), .Z(n14606) );
  NANDN U15357 ( .A(n14605), .B(n14606), .Z(n14298) );
  AND U15358 ( .A(n14299), .B(n14298), .Z(n14614) );
  XOR U15359 ( .A(n14301), .B(n14300), .Z(n14613) );
  XNOR U15360 ( .A(n14303), .B(n14302), .Z(n14304) );
  NANDN U15361 ( .A(n14305), .B(n14304), .Z(n14307) );
  NAND U15362 ( .A(a[45]), .B(b[24]), .Z(n14617) );
  XNOR U15363 ( .A(n14305), .B(n14304), .Z(n14618) );
  NANDN U15364 ( .A(n14617), .B(n14618), .Z(n14306) );
  AND U15365 ( .A(n14307), .B(n14306), .Z(n14626) );
  XOR U15366 ( .A(n14309), .B(n14308), .Z(n14625) );
  XNOR U15367 ( .A(n14311), .B(n14310), .Z(n14312) );
  NANDN U15368 ( .A(n14313), .B(n14312), .Z(n14315) );
  NAND U15369 ( .A(a[47]), .B(b[24]), .Z(n14629) );
  XNOR U15370 ( .A(n14313), .B(n14312), .Z(n14630) );
  NANDN U15371 ( .A(n14629), .B(n14630), .Z(n14314) );
  AND U15372 ( .A(n14315), .B(n14314), .Z(n14638) );
  XOR U15373 ( .A(n14317), .B(n14316), .Z(n14637) );
  XNOR U15374 ( .A(n14319), .B(n14318), .Z(n14320) );
  NANDN U15375 ( .A(n14321), .B(n14320), .Z(n14323) );
  NAND U15376 ( .A(a[49]), .B(b[24]), .Z(n14641) );
  XNOR U15377 ( .A(n14321), .B(n14320), .Z(n14642) );
  NANDN U15378 ( .A(n14641), .B(n14642), .Z(n14322) );
  AND U15379 ( .A(n14323), .B(n14322), .Z(n14650) );
  XOR U15380 ( .A(n14325), .B(n14324), .Z(n14649) );
  XNOR U15381 ( .A(n14327), .B(n14326), .Z(n14328) );
  NANDN U15382 ( .A(n14329), .B(n14328), .Z(n14331) );
  NAND U15383 ( .A(a[51]), .B(b[24]), .Z(n14653) );
  XNOR U15384 ( .A(n14329), .B(n14328), .Z(n14654) );
  NANDN U15385 ( .A(n14653), .B(n14654), .Z(n14330) );
  AND U15386 ( .A(n14331), .B(n14330), .Z(n14662) );
  XOR U15387 ( .A(n14333), .B(n14332), .Z(n14661) );
  XNOR U15388 ( .A(n14335), .B(n14334), .Z(n14336) );
  NANDN U15389 ( .A(n14337), .B(n14336), .Z(n14339) );
  NAND U15390 ( .A(a[53]), .B(b[24]), .Z(n14665) );
  XNOR U15391 ( .A(n14337), .B(n14336), .Z(n14666) );
  NANDN U15392 ( .A(n14665), .B(n14666), .Z(n14338) );
  AND U15393 ( .A(n14339), .B(n14338), .Z(n14674) );
  XOR U15394 ( .A(n14341), .B(n14340), .Z(n14673) );
  XNOR U15395 ( .A(n14343), .B(n14342), .Z(n14344) );
  NANDN U15396 ( .A(n14345), .B(n14344), .Z(n14347) );
  NAND U15397 ( .A(a[55]), .B(b[24]), .Z(n14677) );
  XNOR U15398 ( .A(n14345), .B(n14344), .Z(n14678) );
  NANDN U15399 ( .A(n14677), .B(n14678), .Z(n14346) );
  AND U15400 ( .A(n14347), .B(n14346), .Z(n14686) );
  XOR U15401 ( .A(n14349), .B(n14348), .Z(n14685) );
  XNOR U15402 ( .A(n14351), .B(n14350), .Z(n14352) );
  NANDN U15403 ( .A(n14353), .B(n14352), .Z(n14355) );
  NAND U15404 ( .A(a[57]), .B(b[24]), .Z(n14689) );
  XNOR U15405 ( .A(n14353), .B(n14352), .Z(n14690) );
  NANDN U15406 ( .A(n14689), .B(n14690), .Z(n14354) );
  AND U15407 ( .A(n14355), .B(n14354), .Z(n14698) );
  XOR U15408 ( .A(n14357), .B(n14356), .Z(n14697) );
  XNOR U15409 ( .A(n14359), .B(n14358), .Z(n14360) );
  NANDN U15410 ( .A(n14361), .B(n14360), .Z(n14363) );
  NAND U15411 ( .A(a[59]), .B(b[24]), .Z(n14701) );
  XNOR U15412 ( .A(n14361), .B(n14360), .Z(n14702) );
  NANDN U15413 ( .A(n14701), .B(n14702), .Z(n14362) );
  NAND U15414 ( .A(n14363), .B(n14362), .Z(n14364) );
  XOR U15415 ( .A(n14365), .B(n14364), .Z(n14710) );
  AND U15416 ( .A(a[60]), .B(b[24]), .Z(n14709) );
  AND U15417 ( .A(a[61]), .B(b[24]), .Z(n14368) );
  NANDN U15418 ( .A(n14369), .B(n14368), .Z(n14371) );
  XOR U15419 ( .A(n14367), .B(n14366), .Z(n14715) );
  XNOR U15420 ( .A(n14369), .B(n14368), .Z(n14716) );
  NANDN U15421 ( .A(n14715), .B(n14716), .Z(n14370) );
  NAND U15422 ( .A(n14371), .B(n14370), .Z(n14372) );
  AND U15423 ( .A(a[62]), .B(b[24]), .Z(n14721) );
  XNOR U15424 ( .A(n14373), .B(n14372), .Z(n14722) );
  AND U15425 ( .A(a[63]), .B(b[24]), .Z(n14376) );
  XOR U15426 ( .A(n14375), .B(n14374), .Z(n14723) );
  XOR U15427 ( .A(n14377), .B(n14376), .Z(n14724) );
  XOR U15428 ( .A(n14379), .B(n14378), .Z(n14726) );
  ANDN U15429 ( .B(n14725), .A(n14726), .Z(n24755) );
  XOR U15430 ( .A(n14381), .B(n14380), .Z(n24756) );
  NAND U15431 ( .A(a[62]), .B(b[23]), .Z(n14713) );
  AND U15432 ( .A(a[61]), .B(b[23]), .Z(n14708) );
  NAND U15433 ( .A(a[60]), .B(b[23]), .Z(n14703) );
  AND U15434 ( .A(a[59]), .B(b[23]), .Z(n14696) );
  NAND U15435 ( .A(a[58]), .B(b[23]), .Z(n14691) );
  AND U15436 ( .A(a[57]), .B(b[23]), .Z(n14684) );
  NAND U15437 ( .A(a[56]), .B(b[23]), .Z(n14679) );
  AND U15438 ( .A(a[55]), .B(b[23]), .Z(n14672) );
  NAND U15439 ( .A(a[54]), .B(b[23]), .Z(n14667) );
  AND U15440 ( .A(a[53]), .B(b[23]), .Z(n14660) );
  NAND U15441 ( .A(a[52]), .B(b[23]), .Z(n14655) );
  AND U15442 ( .A(a[51]), .B(b[23]), .Z(n14648) );
  NAND U15443 ( .A(a[50]), .B(b[23]), .Z(n14643) );
  AND U15444 ( .A(a[49]), .B(b[23]), .Z(n14636) );
  NAND U15445 ( .A(a[48]), .B(b[23]), .Z(n14631) );
  AND U15446 ( .A(a[47]), .B(b[23]), .Z(n14624) );
  NAND U15447 ( .A(a[46]), .B(b[23]), .Z(n14619) );
  AND U15448 ( .A(a[45]), .B(b[23]), .Z(n14612) );
  NAND U15449 ( .A(a[43]), .B(b[23]), .Z(n14601) );
  AND U15450 ( .A(a[42]), .B(b[23]), .Z(n14984) );
  XOR U15451 ( .A(n14383), .B(n14382), .Z(n14983) );
  XNOR U15452 ( .A(n14385), .B(n14384), .Z(n14969) );
  XOR U15453 ( .A(n14387), .B(n14386), .Z(n14965) );
  XNOR U15454 ( .A(n14389), .B(n14388), .Z(n14954) );
  XNOR U15455 ( .A(n14391), .B(n14390), .Z(n14940) );
  XNOR U15456 ( .A(n14395), .B(n14394), .Z(n14927) );
  XNOR U15457 ( .A(n14397), .B(n14396), .Z(n14919) );
  XNOR U15458 ( .A(n14399), .B(n14398), .Z(n14909) );
  XNOR U15459 ( .A(n14401), .B(n14400), .Z(n14903) );
  XNOR U15460 ( .A(n14403), .B(n14402), .Z(n14895) );
  XOR U15461 ( .A(n14405), .B(n14404), .Z(n14507) );
  IV U15462 ( .A(n14507), .Z(n14880) );
  NAND U15463 ( .A(a[18]), .B(b[23]), .Z(n14772) );
  XNOR U15464 ( .A(n14407), .B(n14406), .Z(n14408) );
  XOR U15465 ( .A(n14409), .B(n14408), .Z(n14500) );
  IV U15466 ( .A(n14500), .Z(n14874) );
  AND U15467 ( .A(a[16]), .B(b[23]), .Z(n14777) );
  AND U15468 ( .A(a[4]), .B(b[23]), .Z(n14429) );
  AND U15469 ( .A(b[23]), .B(a[0]), .Z(n15107) );
  AND U15470 ( .A(a[1]), .B(b[24]), .Z(n14415) );
  AND U15471 ( .A(n15107), .B(n14415), .Z(n14412) );
  NAND U15472 ( .A(a[2]), .B(n14412), .Z(n14419) );
  NAND U15473 ( .A(b[24]), .B(a[1]), .Z(n14413) );
  XOR U15474 ( .A(n14414), .B(n14413), .Z(n14790) );
  NAND U15475 ( .A(n14415), .B(a[0]), .Z(n14416) );
  XNOR U15476 ( .A(a[2]), .B(n14416), .Z(n14417) );
  AND U15477 ( .A(b[23]), .B(n14417), .Z(n14791) );
  NANDN U15478 ( .A(n14790), .B(n14791), .Z(n14418) );
  AND U15479 ( .A(n14419), .B(n14418), .Z(n14423) );
  NANDN U15480 ( .A(n14423), .B(n14422), .Z(n14425) );
  NAND U15481 ( .A(a[3]), .B(b[23]), .Z(n14798) );
  XNOR U15482 ( .A(n14423), .B(n14422), .Z(n14799) );
  NANDN U15483 ( .A(n14798), .B(n14799), .Z(n14424) );
  AND U15484 ( .A(n14425), .B(n14424), .Z(n14428) );
  NANDN U15485 ( .A(n14429), .B(n14428), .Z(n14431) );
  XOR U15486 ( .A(n14427), .B(n14426), .Z(n14781) );
  XNOR U15487 ( .A(n14429), .B(n14428), .Z(n14780) );
  NANDN U15488 ( .A(n14781), .B(n14780), .Z(n14430) );
  AND U15489 ( .A(n14431), .B(n14430), .Z(n14435) );
  XOR U15490 ( .A(n14433), .B(n14432), .Z(n14434) );
  NAND U15491 ( .A(n14435), .B(n14434), .Z(n14437) );
  NAND U15492 ( .A(a[5]), .B(b[23]), .Z(n14806) );
  XOR U15493 ( .A(n14435), .B(n14434), .Z(n14807) );
  NANDN U15494 ( .A(n14806), .B(n14807), .Z(n14436) );
  AND U15495 ( .A(n14437), .B(n14436), .Z(n14441) );
  NANDN U15496 ( .A(n14441), .B(n14440), .Z(n14443) );
  NAND U15497 ( .A(a[6]), .B(b[23]), .Z(n14812) );
  XNOR U15498 ( .A(n14441), .B(n14440), .Z(n14813) );
  NANDN U15499 ( .A(n14812), .B(n14813), .Z(n14442) );
  AND U15500 ( .A(n14443), .B(n14442), .Z(n14446) );
  NANDN U15501 ( .A(n14446), .B(n14447), .Z(n14449) );
  AND U15502 ( .A(a[7]), .B(b[23]), .Z(n14818) );
  NAND U15503 ( .A(n14819), .B(n14818), .Z(n14448) );
  AND U15504 ( .A(n14449), .B(n14448), .Z(n14450) );
  AND U15505 ( .A(a[8]), .B(b[23]), .Z(n14451) );
  NANDN U15506 ( .A(n14450), .B(n14451), .Z(n14455) );
  NAND U15507 ( .A(n14825), .B(n14824), .Z(n14454) );
  NAND U15508 ( .A(n14455), .B(n14454), .Z(n14456) );
  NAND U15509 ( .A(n14457), .B(n14456), .Z(n14459) );
  NAND U15510 ( .A(a[9]), .B(b[23]), .Z(n14832) );
  XOR U15511 ( .A(n14457), .B(n14456), .Z(n14833) );
  NANDN U15512 ( .A(n14832), .B(n14833), .Z(n14458) );
  AND U15513 ( .A(n14459), .B(n14458), .Z(n14462) );
  AND U15514 ( .A(a[10]), .B(b[23]), .Z(n14463) );
  NANDN U15515 ( .A(n14462), .B(n14463), .Z(n14465) );
  NAND U15516 ( .A(n14837), .B(n14836), .Z(n14464) );
  AND U15517 ( .A(n14465), .B(n14464), .Z(n14468) );
  XOR U15518 ( .A(n14467), .B(n14466), .Z(n14469) );
  NANDN U15519 ( .A(n14468), .B(n14469), .Z(n14471) );
  NAND U15520 ( .A(a[11]), .B(b[23]), .Z(n14844) );
  NANDN U15521 ( .A(n14844), .B(n14845), .Z(n14470) );
  AND U15522 ( .A(n14471), .B(n14470), .Z(n14474) );
  AND U15523 ( .A(a[12]), .B(b[23]), .Z(n14475) );
  NANDN U15524 ( .A(n14474), .B(n14475), .Z(n14477) );
  NAND U15525 ( .A(n14849), .B(n14848), .Z(n14476) );
  AND U15526 ( .A(n14477), .B(n14476), .Z(n14480) );
  XOR U15527 ( .A(n14479), .B(n14478), .Z(n14481) );
  NANDN U15528 ( .A(n14480), .B(n14481), .Z(n14483) );
  NAND U15529 ( .A(a[13]), .B(b[23]), .Z(n14854) );
  NANDN U15530 ( .A(n14854), .B(n14855), .Z(n14482) );
  AND U15531 ( .A(n14483), .B(n14482), .Z(n14486) );
  AND U15532 ( .A(a[14]), .B(b[23]), .Z(n14487) );
  NANDN U15533 ( .A(n14486), .B(n14487), .Z(n14489) );
  NAND U15534 ( .A(n14861), .B(n14860), .Z(n14488) );
  AND U15535 ( .A(n14489), .B(n14488), .Z(n14495) );
  XOR U15536 ( .A(n14491), .B(n14490), .Z(n14492) );
  XOR U15537 ( .A(n14493), .B(n14492), .Z(n14494) );
  NAND U15538 ( .A(n14495), .B(n14494), .Z(n14497) );
  XOR U15539 ( .A(n14495), .B(n14494), .Z(n14869) );
  NAND U15540 ( .A(a[15]), .B(b[23]), .Z(n14868) );
  NAND U15541 ( .A(n14869), .B(n14868), .Z(n14496) );
  AND U15542 ( .A(n14497), .B(n14496), .Z(n14776) );
  NANDN U15543 ( .A(n14874), .B(n14873), .Z(n14503) );
  NOR U15544 ( .A(n14500), .B(n14873), .Z(n14501) );
  AND U15545 ( .A(a[17]), .B(b[23]), .Z(n14872) );
  NANDN U15546 ( .A(n14501), .B(n14872), .Z(n14502) );
  AND U15547 ( .A(n14503), .B(n14502), .Z(n14773) );
  NANDN U15548 ( .A(n14880), .B(n14881), .Z(n14510) );
  NOR U15549 ( .A(n14507), .B(n14881), .Z(n14508) );
  NAND U15550 ( .A(a[19]), .B(b[23]), .Z(n14883) );
  OR U15551 ( .A(n14508), .B(n14883), .Z(n14509) );
  AND U15552 ( .A(n14510), .B(n14509), .Z(n14516) );
  AND U15553 ( .A(a[20]), .B(b[23]), .Z(n14515) );
  NANDN U15554 ( .A(n14516), .B(n14515), .Z(n14518) );
  XNOR U15555 ( .A(n14512), .B(n14511), .Z(n14513) );
  XNOR U15556 ( .A(n14514), .B(n14513), .Z(n14888) );
  XNOR U15557 ( .A(n14516), .B(n14515), .Z(n14887) );
  NAND U15558 ( .A(n14888), .B(n14887), .Z(n14517) );
  NAND U15559 ( .A(n14518), .B(n14517), .Z(n14896) );
  NAND U15560 ( .A(a[21]), .B(b[23]), .Z(n14898) );
  AND U15561 ( .A(a[22]), .B(b[23]), .Z(n14523) );
  NANDN U15562 ( .A(n14524), .B(n14523), .Z(n14526) );
  XNOR U15563 ( .A(n14520), .B(n14519), .Z(n14521) );
  XNOR U15564 ( .A(n14522), .B(n14521), .Z(n14771) );
  XNOR U15565 ( .A(n14524), .B(n14523), .Z(n14770) );
  NAND U15566 ( .A(n14771), .B(n14770), .Z(n14525) );
  NAND U15567 ( .A(n14526), .B(n14525), .Z(n14904) );
  NAND U15568 ( .A(a[23]), .B(b[23]), .Z(n14906) );
  AND U15569 ( .A(a[24]), .B(b[23]), .Z(n14530) );
  NANDN U15570 ( .A(n14531), .B(n14530), .Z(n14533) );
  XNOR U15571 ( .A(n14531), .B(n14530), .Z(n14768) );
  NAND U15572 ( .A(n14769), .B(n14768), .Z(n14532) );
  NAND U15573 ( .A(n14533), .B(n14532), .Z(n14910) );
  NAND U15574 ( .A(a[25]), .B(b[23]), .Z(n14912) );
  AND U15575 ( .A(a[26]), .B(b[23]), .Z(n14537) );
  NANDN U15576 ( .A(n14538), .B(n14537), .Z(n14540) );
  XNOR U15577 ( .A(n14538), .B(n14537), .Z(n14766) );
  NAND U15578 ( .A(n14767), .B(n14766), .Z(n14539) );
  NAND U15579 ( .A(n14540), .B(n14539), .Z(n14920) );
  NAND U15580 ( .A(a[27]), .B(b[23]), .Z(n14922) );
  AND U15581 ( .A(a[28]), .B(b[23]), .Z(n14545) );
  NANDN U15582 ( .A(n14546), .B(n14545), .Z(n14548) );
  XNOR U15583 ( .A(n14542), .B(n14541), .Z(n14543) );
  XNOR U15584 ( .A(n14544), .B(n14543), .Z(n14765) );
  XNOR U15585 ( .A(n14546), .B(n14545), .Z(n14764) );
  NAND U15586 ( .A(n14765), .B(n14764), .Z(n14547) );
  NAND U15587 ( .A(n14548), .B(n14547), .Z(n14928) );
  NAND U15588 ( .A(a[29]), .B(b[23]), .Z(n14930) );
  AND U15589 ( .A(a[30]), .B(b[23]), .Z(n14549) );
  NANDN U15590 ( .A(n14550), .B(n14549), .Z(n14556) );
  XNOR U15591 ( .A(n14550), .B(n14549), .Z(n14763) );
  XNOR U15592 ( .A(n14552), .B(n14551), .Z(n14553) );
  XNOR U15593 ( .A(n14554), .B(n14553), .Z(n14762) );
  NAND U15594 ( .A(n14763), .B(n14762), .Z(n14555) );
  NAND U15595 ( .A(n14556), .B(n14555), .Z(n14935) );
  AND U15596 ( .A(a[31]), .B(b[23]), .Z(n14933) );
  AND U15597 ( .A(a[32]), .B(b[23]), .Z(n14560) );
  NANDN U15598 ( .A(n14561), .B(n14560), .Z(n14563) );
  XNOR U15599 ( .A(n14561), .B(n14560), .Z(n14760) );
  NAND U15600 ( .A(n14761), .B(n14760), .Z(n14562) );
  NAND U15601 ( .A(n14563), .B(n14562), .Z(n14941) );
  NAND U15602 ( .A(a[33]), .B(b[23]), .Z(n14943) );
  AND U15603 ( .A(a[34]), .B(b[23]), .Z(n14567) );
  NANDN U15604 ( .A(n14568), .B(n14567), .Z(n14570) );
  XNOR U15605 ( .A(n14568), .B(n14567), .Z(n14948) );
  NAND U15606 ( .A(n14949), .B(n14948), .Z(n14569) );
  NAND U15607 ( .A(n14570), .B(n14569), .Z(n14955) );
  NAND U15608 ( .A(a[35]), .B(b[23]), .Z(n14957) );
  AND U15609 ( .A(a[36]), .B(b[23]), .Z(n14575) );
  NANDN U15610 ( .A(n14576), .B(n14575), .Z(n14578) );
  XNOR U15611 ( .A(n14572), .B(n14571), .Z(n14573) );
  XNOR U15612 ( .A(n14574), .B(n14573), .Z(n14759) );
  XNOR U15613 ( .A(n14576), .B(n14575), .Z(n14758) );
  NAND U15614 ( .A(n14759), .B(n14758), .Z(n14577) );
  NAND U15615 ( .A(n14578), .B(n14577), .Z(n14966) );
  AND U15616 ( .A(a[37]), .B(b[23]), .Z(n14964) );
  AND U15617 ( .A(a[38]), .B(b[23]), .Z(n14582) );
  NANDN U15618 ( .A(n14583), .B(n14582), .Z(n14585) );
  XNOR U15619 ( .A(n14583), .B(n14582), .Z(n14756) );
  NAND U15620 ( .A(n14757), .B(n14756), .Z(n14584) );
  NAND U15621 ( .A(n14585), .B(n14584), .Z(n14970) );
  NAND U15622 ( .A(a[39]), .B(b[23]), .Z(n14972) );
  AND U15623 ( .A(a[40]), .B(b[23]), .Z(n14589) );
  NANDN U15624 ( .A(n14590), .B(n14589), .Z(n14592) );
  XNOR U15625 ( .A(n14590), .B(n14589), .Z(n14754) );
  NAND U15626 ( .A(n14755), .B(n14754), .Z(n14591) );
  AND U15627 ( .A(n14592), .B(n14591), .Z(n14596) );
  NAND U15628 ( .A(n14596), .B(n14595), .Z(n14598) );
  XOR U15629 ( .A(n14596), .B(n14595), .Z(n14978) );
  NAND U15630 ( .A(a[41]), .B(b[23]), .Z(n14977) );
  NAND U15631 ( .A(n14978), .B(n14977), .Z(n14597) );
  AND U15632 ( .A(n14598), .B(n14597), .Z(n14986) );
  NANDN U15633 ( .A(n14601), .B(n14602), .Z(n14604) );
  XOR U15634 ( .A(n14600), .B(n14599), .Z(n14752) );
  XNOR U15635 ( .A(n14602), .B(n14601), .Z(n14753) );
  NANDN U15636 ( .A(n14752), .B(n14753), .Z(n14603) );
  AND U15637 ( .A(n14604), .B(n14603), .Z(n14608) );
  AND U15638 ( .A(a[44]), .B(b[23]), .Z(n14607) );
  NANDN U15639 ( .A(n14608), .B(n14607), .Z(n14610) );
  XOR U15640 ( .A(n14606), .B(n14605), .Z(n14995) );
  XNOR U15641 ( .A(n14608), .B(n14607), .Z(n14996) );
  NANDN U15642 ( .A(n14995), .B(n14996), .Z(n14609) );
  AND U15643 ( .A(n14610), .B(n14609), .Z(n14611) );
  NANDN U15644 ( .A(n14612), .B(n14611), .Z(n14616) );
  XOR U15645 ( .A(n14612), .B(n14611), .Z(n14750) );
  XOR U15646 ( .A(n14614), .B(n14613), .Z(n14751) );
  NANDN U15647 ( .A(n14750), .B(n14751), .Z(n14615) );
  AND U15648 ( .A(n14616), .B(n14615), .Z(n14620) );
  NANDN U15649 ( .A(n14619), .B(n14620), .Z(n14622) );
  XOR U15650 ( .A(n14618), .B(n14617), .Z(n15003) );
  XNOR U15651 ( .A(n14620), .B(n14619), .Z(n15004) );
  NANDN U15652 ( .A(n15003), .B(n15004), .Z(n14621) );
  AND U15653 ( .A(n14622), .B(n14621), .Z(n14623) );
  NANDN U15654 ( .A(n14624), .B(n14623), .Z(n14628) );
  XOR U15655 ( .A(n14624), .B(n14623), .Z(n14748) );
  XOR U15656 ( .A(n14626), .B(n14625), .Z(n14749) );
  NANDN U15657 ( .A(n14748), .B(n14749), .Z(n14627) );
  AND U15658 ( .A(n14628), .B(n14627), .Z(n14632) );
  NANDN U15659 ( .A(n14631), .B(n14632), .Z(n14634) );
  XOR U15660 ( .A(n14630), .B(n14629), .Z(n15011) );
  XNOR U15661 ( .A(n14632), .B(n14631), .Z(n15012) );
  NANDN U15662 ( .A(n15011), .B(n15012), .Z(n14633) );
  AND U15663 ( .A(n14634), .B(n14633), .Z(n14635) );
  NANDN U15664 ( .A(n14636), .B(n14635), .Z(n14640) );
  XOR U15665 ( .A(n14636), .B(n14635), .Z(n14746) );
  XOR U15666 ( .A(n14638), .B(n14637), .Z(n14747) );
  NANDN U15667 ( .A(n14746), .B(n14747), .Z(n14639) );
  AND U15668 ( .A(n14640), .B(n14639), .Z(n14644) );
  NANDN U15669 ( .A(n14643), .B(n14644), .Z(n14646) );
  XOR U15670 ( .A(n14642), .B(n14641), .Z(n15019) );
  XNOR U15671 ( .A(n14644), .B(n14643), .Z(n15020) );
  NANDN U15672 ( .A(n15019), .B(n15020), .Z(n14645) );
  AND U15673 ( .A(n14646), .B(n14645), .Z(n14647) );
  NANDN U15674 ( .A(n14648), .B(n14647), .Z(n14652) );
  XOR U15675 ( .A(n14648), .B(n14647), .Z(n14744) );
  XOR U15676 ( .A(n14650), .B(n14649), .Z(n14745) );
  NANDN U15677 ( .A(n14744), .B(n14745), .Z(n14651) );
  AND U15678 ( .A(n14652), .B(n14651), .Z(n14656) );
  NANDN U15679 ( .A(n14655), .B(n14656), .Z(n14658) );
  XOR U15680 ( .A(n14654), .B(n14653), .Z(n15027) );
  XNOR U15681 ( .A(n14656), .B(n14655), .Z(n15028) );
  NANDN U15682 ( .A(n15027), .B(n15028), .Z(n14657) );
  AND U15683 ( .A(n14658), .B(n14657), .Z(n14659) );
  NANDN U15684 ( .A(n14660), .B(n14659), .Z(n14664) );
  XOR U15685 ( .A(n14660), .B(n14659), .Z(n14742) );
  XOR U15686 ( .A(n14662), .B(n14661), .Z(n14743) );
  NANDN U15687 ( .A(n14742), .B(n14743), .Z(n14663) );
  AND U15688 ( .A(n14664), .B(n14663), .Z(n14668) );
  NANDN U15689 ( .A(n14667), .B(n14668), .Z(n14670) );
  XOR U15690 ( .A(n14666), .B(n14665), .Z(n15035) );
  XNOR U15691 ( .A(n14668), .B(n14667), .Z(n15036) );
  NANDN U15692 ( .A(n15035), .B(n15036), .Z(n14669) );
  AND U15693 ( .A(n14670), .B(n14669), .Z(n14671) );
  NANDN U15694 ( .A(n14672), .B(n14671), .Z(n14676) );
  XOR U15695 ( .A(n14672), .B(n14671), .Z(n14740) );
  XOR U15696 ( .A(n14674), .B(n14673), .Z(n14741) );
  NANDN U15697 ( .A(n14740), .B(n14741), .Z(n14675) );
  AND U15698 ( .A(n14676), .B(n14675), .Z(n14680) );
  NANDN U15699 ( .A(n14679), .B(n14680), .Z(n14682) );
  XOR U15700 ( .A(n14678), .B(n14677), .Z(n15043) );
  XNOR U15701 ( .A(n14680), .B(n14679), .Z(n15044) );
  NANDN U15702 ( .A(n15043), .B(n15044), .Z(n14681) );
  AND U15703 ( .A(n14682), .B(n14681), .Z(n14683) );
  NANDN U15704 ( .A(n14684), .B(n14683), .Z(n14688) );
  XOR U15705 ( .A(n14684), .B(n14683), .Z(n14738) );
  XOR U15706 ( .A(n14686), .B(n14685), .Z(n14739) );
  NANDN U15707 ( .A(n14738), .B(n14739), .Z(n14687) );
  AND U15708 ( .A(n14688), .B(n14687), .Z(n14692) );
  NANDN U15709 ( .A(n14691), .B(n14692), .Z(n14694) );
  XOR U15710 ( .A(n14690), .B(n14689), .Z(n15051) );
  XNOR U15711 ( .A(n14692), .B(n14691), .Z(n15052) );
  NANDN U15712 ( .A(n15051), .B(n15052), .Z(n14693) );
  AND U15713 ( .A(n14694), .B(n14693), .Z(n14695) );
  NANDN U15714 ( .A(n14696), .B(n14695), .Z(n14700) );
  XOR U15715 ( .A(n14696), .B(n14695), .Z(n14736) );
  XOR U15716 ( .A(n14698), .B(n14697), .Z(n14737) );
  NANDN U15717 ( .A(n14736), .B(n14737), .Z(n14699) );
  AND U15718 ( .A(n14700), .B(n14699), .Z(n14704) );
  NANDN U15719 ( .A(n14703), .B(n14704), .Z(n14706) );
  XOR U15720 ( .A(n14702), .B(n14701), .Z(n15059) );
  XNOR U15721 ( .A(n14704), .B(n14703), .Z(n15060) );
  NANDN U15722 ( .A(n15059), .B(n15060), .Z(n14705) );
  AND U15723 ( .A(n14706), .B(n14705), .Z(n14707) );
  NANDN U15724 ( .A(n14708), .B(n14707), .Z(n14712) );
  XOR U15725 ( .A(n14708), .B(n14707), .Z(n14732) );
  XOR U15726 ( .A(n14710), .B(n14709), .Z(n14733) );
  OR U15727 ( .A(n14732), .B(n14733), .Z(n14711) );
  AND U15728 ( .A(n14712), .B(n14711), .Z(n14714) );
  NANDN U15729 ( .A(n14713), .B(n14714), .Z(n14718) );
  XOR U15730 ( .A(n14714), .B(n14713), .Z(n15067) );
  XNOR U15731 ( .A(n14716), .B(n14715), .Z(n15068) );
  NANDN U15732 ( .A(n15067), .B(n15068), .Z(n14717) );
  AND U15733 ( .A(n14718), .B(n14717), .Z(n14719) );
  NAND U15734 ( .A(a[63]), .B(b[23]), .Z(n14720) );
  XNOR U15735 ( .A(n14720), .B(n14719), .Z(n14730) );
  XOR U15736 ( .A(n14722), .B(n14721), .Z(n14731) );
  XOR U15737 ( .A(n14724), .B(n14723), .Z(n14728) );
  NAND U15738 ( .A(n14729), .B(n14728), .Z(n24746) );
  IV U15739 ( .A(n24746), .Z(n14727) );
  XOR U15740 ( .A(n14726), .B(n14725), .Z(n24745) );
  NANDN U15741 ( .A(n14727), .B(n24745), .Z(n24753) );
  XOR U15742 ( .A(n14729), .B(n14728), .Z(n24739) );
  XOR U15743 ( .A(n14731), .B(n14730), .Z(n15074) );
  XOR U15744 ( .A(n14733), .B(n14732), .Z(n14735) );
  AND U15745 ( .A(a[62]), .B(b[22]), .Z(n14734) );
  NANDN U15746 ( .A(n14735), .B(n14734), .Z(n15066) );
  XOR U15747 ( .A(n14735), .B(n14734), .Z(n15419) );
  XOR U15748 ( .A(n14737), .B(n14736), .Z(n15058) );
  AND U15749 ( .A(a[60]), .B(b[22]), .Z(n15057) );
  XOR U15750 ( .A(n14739), .B(n14738), .Z(n15050) );
  AND U15751 ( .A(a[58]), .B(b[22]), .Z(n15049) );
  XOR U15752 ( .A(n14741), .B(n14740), .Z(n15042) );
  AND U15753 ( .A(a[56]), .B(b[22]), .Z(n15041) );
  XOR U15754 ( .A(n14743), .B(n14742), .Z(n15034) );
  AND U15755 ( .A(a[54]), .B(b[22]), .Z(n15033) );
  XOR U15756 ( .A(n14745), .B(n14744), .Z(n15026) );
  AND U15757 ( .A(a[52]), .B(b[22]), .Z(n15025) );
  XOR U15758 ( .A(n14747), .B(n14746), .Z(n15018) );
  AND U15759 ( .A(a[50]), .B(b[22]), .Z(n15017) );
  XOR U15760 ( .A(n14749), .B(n14748), .Z(n15010) );
  AND U15761 ( .A(a[48]), .B(b[22]), .Z(n15009) );
  XOR U15762 ( .A(n14751), .B(n14750), .Z(n15002) );
  AND U15763 ( .A(a[46]), .B(b[22]), .Z(n15001) );
  NAND U15764 ( .A(a[44]), .B(b[22]), .Z(n14991) );
  XNOR U15765 ( .A(n14753), .B(n14752), .Z(n14992) );
  NANDN U15766 ( .A(n14991), .B(n14992), .Z(n14994) );
  XNOR U15767 ( .A(n14755), .B(n14754), .Z(n15299) );
  XNOR U15768 ( .A(n14757), .B(n14756), .Z(n15290) );
  XNOR U15769 ( .A(n14759), .B(n14758), .Z(n15282) );
  XNOR U15770 ( .A(n14761), .B(n14760), .Z(n15264) );
  XNOR U15771 ( .A(n14763), .B(n14762), .Z(n15256) );
  XNOR U15772 ( .A(n14765), .B(n14764), .Z(n15248) );
  XNOR U15773 ( .A(n14767), .B(n14766), .Z(n15242) );
  XNOR U15774 ( .A(n14769), .B(n14768), .Z(n15232) );
  XNOR U15775 ( .A(n14771), .B(n14770), .Z(n15224) );
  XOR U15776 ( .A(n14773), .B(n14772), .Z(n14774) );
  XOR U15777 ( .A(n14775), .B(n14774), .Z(n14875) );
  IV U15778 ( .A(n14875), .Z(n15205) );
  NAND U15779 ( .A(a[18]), .B(b[22]), .Z(n15098) );
  XNOR U15780 ( .A(n14777), .B(n14776), .Z(n14778) );
  XOR U15781 ( .A(n14779), .B(n14778), .Z(n15196) );
  AND U15782 ( .A(a[8]), .B(b[22]), .Z(n14820) );
  XOR U15783 ( .A(n14781), .B(n14780), .Z(n14803) );
  AND U15784 ( .A(b[22]), .B(a[0]), .Z(n15474) );
  AND U15785 ( .A(a[1]), .B(b[23]), .Z(n14785) );
  AND U15786 ( .A(n15474), .B(n14785), .Z(n14782) );
  NAND U15787 ( .A(a[2]), .B(n14782), .Z(n14789) );
  NAND U15788 ( .A(b[23]), .B(a[1]), .Z(n14783) );
  XOR U15789 ( .A(n14784), .B(n14783), .Z(n15113) );
  NAND U15790 ( .A(n14785), .B(a[0]), .Z(n14786) );
  XNOR U15791 ( .A(a[2]), .B(n14786), .Z(n14787) );
  AND U15792 ( .A(b[22]), .B(n14787), .Z(n15114) );
  NANDN U15793 ( .A(n15113), .B(n15114), .Z(n14788) );
  AND U15794 ( .A(n14789), .B(n14788), .Z(n14793) );
  XNOR U15795 ( .A(n14791), .B(n14790), .Z(n14792) );
  NANDN U15796 ( .A(n14793), .B(n14792), .Z(n14795) );
  XNOR U15797 ( .A(n14793), .B(n14792), .Z(n15120) );
  AND U15798 ( .A(a[3]), .B(b[22]), .Z(n15119) );
  NAND U15799 ( .A(n15120), .B(n15119), .Z(n14794) );
  AND U15800 ( .A(n14795), .B(n14794), .Z(n14797) );
  AND U15801 ( .A(a[4]), .B(b[22]), .Z(n14796) );
  NANDN U15802 ( .A(n14797), .B(n14796), .Z(n14801) );
  XNOR U15803 ( .A(n14797), .B(n14796), .Z(n15126) );
  XNOR U15804 ( .A(n14799), .B(n14798), .Z(n15125) );
  NAND U15805 ( .A(n15126), .B(n15125), .Z(n14800) );
  NAND U15806 ( .A(n14801), .B(n14800), .Z(n14802) );
  NAND U15807 ( .A(n14803), .B(n14802), .Z(n14805) );
  NAND U15808 ( .A(a[5]), .B(b[22]), .Z(n15131) );
  XOR U15809 ( .A(n14803), .B(n14802), .Z(n15132) );
  NANDN U15810 ( .A(n15131), .B(n15132), .Z(n14804) );
  AND U15811 ( .A(n14805), .B(n14804), .Z(n14809) );
  XNOR U15812 ( .A(n14807), .B(n14806), .Z(n14808) );
  NANDN U15813 ( .A(n14809), .B(n14808), .Z(n14811) );
  NAND U15814 ( .A(a[6]), .B(b[22]), .Z(n15137) );
  XNOR U15815 ( .A(n14809), .B(n14808), .Z(n15138) );
  NANDN U15816 ( .A(n15137), .B(n15138), .Z(n14810) );
  AND U15817 ( .A(n14811), .B(n14810), .Z(n14815) );
  XNOR U15818 ( .A(n14813), .B(n14812), .Z(n14814) );
  NANDN U15819 ( .A(n14815), .B(n14814), .Z(n14817) );
  NAND U15820 ( .A(a[7]), .B(b[22]), .Z(n15145) );
  XNOR U15821 ( .A(n14815), .B(n14814), .Z(n15146) );
  NANDN U15822 ( .A(n15145), .B(n15146), .Z(n14816) );
  AND U15823 ( .A(n14817), .B(n14816), .Z(n14821) );
  NANDN U15824 ( .A(n14820), .B(n14821), .Z(n14823) );
  XOR U15825 ( .A(n14819), .B(n14818), .Z(n15103) );
  NANDN U15826 ( .A(n15103), .B(n15104), .Z(n14822) );
  AND U15827 ( .A(n14823), .B(n14822), .Z(n14827) );
  XOR U15828 ( .A(n14825), .B(n14824), .Z(n14826) );
  NAND U15829 ( .A(n14827), .B(n14826), .Z(n14829) );
  NAND U15830 ( .A(a[9]), .B(b[22]), .Z(n15153) );
  XOR U15831 ( .A(n14827), .B(n14826), .Z(n15154) );
  NANDN U15832 ( .A(n15153), .B(n15154), .Z(n14828) );
  AND U15833 ( .A(n14829), .B(n14828), .Z(n14830) );
  AND U15834 ( .A(a[10]), .B(b[22]), .Z(n14831) );
  NANDN U15835 ( .A(n14830), .B(n14831), .Z(n14835) );
  NAND U15836 ( .A(n15160), .B(n15159), .Z(n14834) );
  AND U15837 ( .A(n14835), .B(n14834), .Z(n14838) );
  XOR U15838 ( .A(n14837), .B(n14836), .Z(n14839) );
  NANDN U15839 ( .A(n14838), .B(n14839), .Z(n14841) );
  NAND U15840 ( .A(a[11]), .B(b[22]), .Z(n15165) );
  NANDN U15841 ( .A(n15165), .B(n15166), .Z(n14840) );
  AND U15842 ( .A(n14841), .B(n14840), .Z(n14842) );
  AND U15843 ( .A(a[12]), .B(b[22]), .Z(n14843) );
  NANDN U15844 ( .A(n14842), .B(n14843), .Z(n14847) );
  NAND U15845 ( .A(n15172), .B(n15171), .Z(n14846) );
  AND U15846 ( .A(n14847), .B(n14846), .Z(n14850) );
  XOR U15847 ( .A(n14849), .B(n14848), .Z(n14851) );
  NANDN U15848 ( .A(n14850), .B(n14851), .Z(n14853) );
  NAND U15849 ( .A(a[13]), .B(b[22]), .Z(n15177) );
  NANDN U15850 ( .A(n15177), .B(n15178), .Z(n14852) );
  AND U15851 ( .A(n14853), .B(n14852), .Z(n14856) );
  AND U15852 ( .A(a[14]), .B(b[22]), .Z(n14857) );
  NANDN U15853 ( .A(n14856), .B(n14857), .Z(n14859) );
  NAND U15854 ( .A(n15184), .B(n15183), .Z(n14858) );
  AND U15855 ( .A(n14859), .B(n14858), .Z(n14862) );
  XOR U15856 ( .A(n14861), .B(n14860), .Z(n14863) );
  NANDN U15857 ( .A(n14862), .B(n14863), .Z(n14865) );
  AND U15858 ( .A(a[15]), .B(b[22]), .Z(n15190) );
  NAND U15859 ( .A(n15190), .B(n15189), .Z(n14864) );
  AND U15860 ( .A(n14865), .B(n14864), .Z(n14866) );
  AND U15861 ( .A(a[16]), .B(b[22]), .Z(n14867) );
  NANDN U15862 ( .A(n14866), .B(n14867), .Z(n14871) );
  XNOR U15863 ( .A(n14869), .B(n14868), .Z(n15101) );
  NAND U15864 ( .A(n15102), .B(n15101), .Z(n14870) );
  NAND U15865 ( .A(n14871), .B(n14870), .Z(n15195) );
  NAND U15866 ( .A(a[17]), .B(b[22]), .Z(n15197) );
  NANDN U15867 ( .A(n15205), .B(n15204), .Z(n14878) );
  NOR U15868 ( .A(n14875), .B(n15204), .Z(n14876) );
  AND U15869 ( .A(a[19]), .B(b[22]), .Z(n15203) );
  NANDN U15870 ( .A(n14876), .B(n15203), .Z(n14877) );
  AND U15871 ( .A(n14878), .B(n14877), .Z(n15209) );
  AND U15872 ( .A(a[20]), .B(b[22]), .Z(n14879) );
  IV U15873 ( .A(n14879), .Z(n15210) );
  OR U15874 ( .A(n15209), .B(n15210), .Z(n14886) );
  ANDN U15875 ( .B(n15209), .A(n14879), .Z(n14884) );
  XOR U15876 ( .A(n14881), .B(n14880), .Z(n14882) );
  XNOR U15877 ( .A(n14883), .B(n14882), .Z(n15212) );
  OR U15878 ( .A(n14884), .B(n15212), .Z(n14885) );
  AND U15879 ( .A(n14886), .B(n14885), .Z(n15216) );
  XOR U15880 ( .A(n14888), .B(n14887), .Z(n14889) );
  IV U15881 ( .A(n14889), .Z(n15215) );
  OR U15882 ( .A(n15216), .B(n15215), .Z(n14892) );
  ANDN U15883 ( .B(n15216), .A(n14889), .Z(n14890) );
  AND U15884 ( .A(a[21]), .B(b[22]), .Z(n15214) );
  NANDN U15885 ( .A(n14890), .B(n15214), .Z(n14891) );
  AND U15886 ( .A(n14892), .B(n14891), .Z(n14894) );
  AND U15887 ( .A(a[22]), .B(b[22]), .Z(n14893) );
  NANDN U15888 ( .A(n14894), .B(n14893), .Z(n14900) );
  XOR U15889 ( .A(n14894), .B(n14893), .Z(n15095) );
  XNOR U15890 ( .A(n14896), .B(n14895), .Z(n14897) );
  XNOR U15891 ( .A(n14898), .B(n14897), .Z(n15096) );
  NANDN U15892 ( .A(n15095), .B(n15096), .Z(n14899) );
  NAND U15893 ( .A(n14900), .B(n14899), .Z(n15225) );
  NAND U15894 ( .A(a[23]), .B(b[22]), .Z(n15227) );
  AND U15895 ( .A(a[24]), .B(b[22]), .Z(n14902) );
  NANDN U15896 ( .A(n14901), .B(n14902), .Z(n14908) );
  XNOR U15897 ( .A(n14902), .B(n14901), .Z(n15094) );
  XNOR U15898 ( .A(n14904), .B(n14903), .Z(n14905) );
  XNOR U15899 ( .A(n14906), .B(n14905), .Z(n15093) );
  NAND U15900 ( .A(n15094), .B(n15093), .Z(n14907) );
  NAND U15901 ( .A(n14908), .B(n14907), .Z(n15233) );
  NAND U15902 ( .A(a[25]), .B(b[22]), .Z(n15235) );
  AND U15903 ( .A(a[26]), .B(b[22]), .Z(n14914) );
  NANDN U15904 ( .A(n14913), .B(n14914), .Z(n14916) );
  XNOR U15905 ( .A(n14910), .B(n14909), .Z(n14911) );
  XNOR U15906 ( .A(n14912), .B(n14911), .Z(n15092) );
  XNOR U15907 ( .A(n14914), .B(n14913), .Z(n15091) );
  NAND U15908 ( .A(n15092), .B(n15091), .Z(n14915) );
  NAND U15909 ( .A(n14916), .B(n14915), .Z(n15243) );
  NAND U15910 ( .A(a[27]), .B(b[22]), .Z(n15245) );
  AND U15911 ( .A(a[28]), .B(b[22]), .Z(n14918) );
  NANDN U15912 ( .A(n14917), .B(n14918), .Z(n14924) );
  XNOR U15913 ( .A(n14918), .B(n14917), .Z(n15090) );
  XNOR U15914 ( .A(n14920), .B(n14919), .Z(n14921) );
  XNOR U15915 ( .A(n14922), .B(n14921), .Z(n15089) );
  NAND U15916 ( .A(n15090), .B(n15089), .Z(n14923) );
  NAND U15917 ( .A(n14924), .B(n14923), .Z(n15249) );
  NAND U15918 ( .A(a[29]), .B(b[22]), .Z(n15251) );
  AND U15919 ( .A(a[30]), .B(b[22]), .Z(n14926) );
  NANDN U15920 ( .A(n14925), .B(n14926), .Z(n14932) );
  XNOR U15921 ( .A(n14926), .B(n14925), .Z(n15088) );
  XNOR U15922 ( .A(n14928), .B(n14927), .Z(n14929) );
  XNOR U15923 ( .A(n14930), .B(n14929), .Z(n15087) );
  NAND U15924 ( .A(n15088), .B(n15087), .Z(n14931) );
  NAND U15925 ( .A(n14932), .B(n14931), .Z(n15257) );
  NAND U15926 ( .A(a[31]), .B(b[22]), .Z(n15259) );
  AND U15927 ( .A(a[32]), .B(b[22]), .Z(n14937) );
  NANDN U15928 ( .A(n14936), .B(n14937), .Z(n14939) );
  XNOR U15929 ( .A(n14937), .B(n14936), .Z(n15085) );
  NAND U15930 ( .A(n15086), .B(n15085), .Z(n14938) );
  NAND U15931 ( .A(n14939), .B(n14938), .Z(n15265) );
  NAND U15932 ( .A(a[33]), .B(b[22]), .Z(n15267) );
  AND U15933 ( .A(a[34]), .B(b[22]), .Z(n14945) );
  NANDN U15934 ( .A(n14944), .B(n14945), .Z(n14947) );
  XNOR U15935 ( .A(n14941), .B(n14940), .Z(n14942) );
  XNOR U15936 ( .A(n14943), .B(n14942), .Z(n15084) );
  XNOR U15937 ( .A(n14945), .B(n14944), .Z(n15083) );
  NAND U15938 ( .A(n15084), .B(n15083), .Z(n14946) );
  AND U15939 ( .A(n14947), .B(n14946), .Z(n15274) );
  XOR U15940 ( .A(n14949), .B(n14948), .Z(n14950) );
  IV U15941 ( .A(n14950), .Z(n15275) );
  OR U15942 ( .A(n15274), .B(n15275), .Z(n14953) );
  ANDN U15943 ( .B(n15274), .A(n14950), .Z(n14951) );
  NAND U15944 ( .A(a[35]), .B(b[22]), .Z(n15277) );
  OR U15945 ( .A(n14951), .B(n15277), .Z(n14952) );
  AND U15946 ( .A(n14953), .B(n14952), .Z(n14958) );
  AND U15947 ( .A(a[36]), .B(b[22]), .Z(n14959) );
  NANDN U15948 ( .A(n14958), .B(n14959), .Z(n14961) );
  XNOR U15949 ( .A(n14955), .B(n14954), .Z(n14956) );
  XNOR U15950 ( .A(n14957), .B(n14956), .Z(n15082) );
  XNOR U15951 ( .A(n14959), .B(n14958), .Z(n15081) );
  NAND U15952 ( .A(n15082), .B(n15081), .Z(n14960) );
  NAND U15953 ( .A(n14961), .B(n14960), .Z(n15283) );
  NAND U15954 ( .A(a[37]), .B(b[22]), .Z(n15285) );
  AND U15955 ( .A(a[38]), .B(b[22]), .Z(n14963) );
  NANDN U15956 ( .A(n14962), .B(n14963), .Z(n14968) );
  XNOR U15957 ( .A(n14963), .B(n14962), .Z(n15080) );
  NAND U15958 ( .A(n15080), .B(n15079), .Z(n14967) );
  NAND U15959 ( .A(n14968), .B(n14967), .Z(n15291) );
  NAND U15960 ( .A(a[39]), .B(b[22]), .Z(n15293) );
  AND U15961 ( .A(a[40]), .B(b[22]), .Z(n14974) );
  NANDN U15962 ( .A(n14973), .B(n14974), .Z(n14976) );
  XNOR U15963 ( .A(n14970), .B(n14969), .Z(n14971) );
  XOR U15964 ( .A(n14972), .B(n14971), .Z(n15296) );
  XNOR U15965 ( .A(n14974), .B(n14973), .Z(n15297) );
  NANDN U15966 ( .A(n15296), .B(n15297), .Z(n14975) );
  NAND U15967 ( .A(n14976), .B(n14975), .Z(n15300) );
  NAND U15968 ( .A(a[41]), .B(b[22]), .Z(n15302) );
  AND U15969 ( .A(a[42]), .B(b[22]), .Z(n14979) );
  NANDN U15970 ( .A(n14980), .B(n14979), .Z(n14982) );
  XOR U15971 ( .A(n14978), .B(n14977), .Z(n15307) );
  XNOR U15972 ( .A(n14980), .B(n14979), .Z(n15308) );
  NANDN U15973 ( .A(n15307), .B(n15308), .Z(n14981) );
  AND U15974 ( .A(n14982), .B(n14981), .Z(n14988) );
  AND U15975 ( .A(a[43]), .B(b[22]), .Z(n14987) );
  NANDN U15976 ( .A(n14988), .B(n14987), .Z(n14990) );
  XOR U15977 ( .A(n14984), .B(n14983), .Z(n14985) );
  XNOR U15978 ( .A(n14986), .B(n14985), .Z(n15078) );
  XNOR U15979 ( .A(n14988), .B(n14987), .Z(n15077) );
  NAND U15980 ( .A(n15078), .B(n15077), .Z(n14989) );
  AND U15981 ( .A(n14990), .B(n14989), .Z(n15314) );
  XNOR U15982 ( .A(n14992), .B(n14991), .Z(n15313) );
  NANDN U15983 ( .A(n15314), .B(n15313), .Z(n14993) );
  AND U15984 ( .A(n14994), .B(n14993), .Z(n14998) );
  XNOR U15985 ( .A(n14996), .B(n14995), .Z(n14997) );
  NANDN U15986 ( .A(n14998), .B(n14997), .Z(n15000) );
  NAND U15987 ( .A(a[45]), .B(b[22]), .Z(n15315) );
  XNOR U15988 ( .A(n14998), .B(n14997), .Z(n15316) );
  NANDN U15989 ( .A(n15315), .B(n15316), .Z(n14999) );
  AND U15990 ( .A(n15000), .B(n14999), .Z(n15324) );
  XOR U15991 ( .A(n15002), .B(n15001), .Z(n15323) );
  XNOR U15992 ( .A(n15004), .B(n15003), .Z(n15005) );
  NANDN U15993 ( .A(n15006), .B(n15005), .Z(n15008) );
  NAND U15994 ( .A(a[47]), .B(b[22]), .Z(n15327) );
  XNOR U15995 ( .A(n15006), .B(n15005), .Z(n15328) );
  NANDN U15996 ( .A(n15327), .B(n15328), .Z(n15007) );
  AND U15997 ( .A(n15008), .B(n15007), .Z(n15336) );
  XOR U15998 ( .A(n15010), .B(n15009), .Z(n15335) );
  XNOR U15999 ( .A(n15012), .B(n15011), .Z(n15013) );
  NANDN U16000 ( .A(n15014), .B(n15013), .Z(n15016) );
  NAND U16001 ( .A(a[49]), .B(b[22]), .Z(n15339) );
  XNOR U16002 ( .A(n15014), .B(n15013), .Z(n15340) );
  NANDN U16003 ( .A(n15339), .B(n15340), .Z(n15015) );
  AND U16004 ( .A(n15016), .B(n15015), .Z(n15348) );
  XOR U16005 ( .A(n15018), .B(n15017), .Z(n15347) );
  XNOR U16006 ( .A(n15020), .B(n15019), .Z(n15021) );
  NANDN U16007 ( .A(n15022), .B(n15021), .Z(n15024) );
  NAND U16008 ( .A(a[51]), .B(b[22]), .Z(n15351) );
  XNOR U16009 ( .A(n15022), .B(n15021), .Z(n15352) );
  NANDN U16010 ( .A(n15351), .B(n15352), .Z(n15023) );
  AND U16011 ( .A(n15024), .B(n15023), .Z(n15360) );
  XOR U16012 ( .A(n15026), .B(n15025), .Z(n15359) );
  XNOR U16013 ( .A(n15028), .B(n15027), .Z(n15029) );
  NANDN U16014 ( .A(n15030), .B(n15029), .Z(n15032) );
  NAND U16015 ( .A(a[53]), .B(b[22]), .Z(n15363) );
  XNOR U16016 ( .A(n15030), .B(n15029), .Z(n15364) );
  NANDN U16017 ( .A(n15363), .B(n15364), .Z(n15031) );
  AND U16018 ( .A(n15032), .B(n15031), .Z(n15372) );
  XOR U16019 ( .A(n15034), .B(n15033), .Z(n15371) );
  XNOR U16020 ( .A(n15036), .B(n15035), .Z(n15037) );
  NANDN U16021 ( .A(n15038), .B(n15037), .Z(n15040) );
  NAND U16022 ( .A(a[55]), .B(b[22]), .Z(n15375) );
  XNOR U16023 ( .A(n15038), .B(n15037), .Z(n15376) );
  NANDN U16024 ( .A(n15375), .B(n15376), .Z(n15039) );
  AND U16025 ( .A(n15040), .B(n15039), .Z(n15384) );
  XOR U16026 ( .A(n15042), .B(n15041), .Z(n15383) );
  XNOR U16027 ( .A(n15044), .B(n15043), .Z(n15045) );
  NANDN U16028 ( .A(n15046), .B(n15045), .Z(n15048) );
  NAND U16029 ( .A(a[57]), .B(b[22]), .Z(n15387) );
  XNOR U16030 ( .A(n15046), .B(n15045), .Z(n15388) );
  NANDN U16031 ( .A(n15387), .B(n15388), .Z(n15047) );
  AND U16032 ( .A(n15048), .B(n15047), .Z(n15396) );
  XOR U16033 ( .A(n15050), .B(n15049), .Z(n15395) );
  XNOR U16034 ( .A(n15052), .B(n15051), .Z(n15053) );
  NANDN U16035 ( .A(n15054), .B(n15053), .Z(n15056) );
  NAND U16036 ( .A(a[59]), .B(b[22]), .Z(n15399) );
  XNOR U16037 ( .A(n15054), .B(n15053), .Z(n15400) );
  NANDN U16038 ( .A(n15399), .B(n15400), .Z(n15055) );
  AND U16039 ( .A(n15056), .B(n15055), .Z(n15408) );
  XOR U16040 ( .A(n15058), .B(n15057), .Z(n15407) );
  XNOR U16041 ( .A(n15060), .B(n15059), .Z(n15061) );
  NANDN U16042 ( .A(n15062), .B(n15061), .Z(n15064) );
  NAND U16043 ( .A(a[61]), .B(b[22]), .Z(n15411) );
  XNOR U16044 ( .A(n15062), .B(n15061), .Z(n15412) );
  NANDN U16045 ( .A(n15411), .B(n15412), .Z(n15063) );
  AND U16046 ( .A(n15064), .B(n15063), .Z(n15420) );
  OR U16047 ( .A(n15419), .B(n15420), .Z(n15065) );
  AND U16048 ( .A(n15066), .B(n15065), .Z(n15070) );
  XNOR U16049 ( .A(n15068), .B(n15067), .Z(n15069) );
  NANDN U16050 ( .A(n15070), .B(n15069), .Z(n15072) );
  NAND U16051 ( .A(a[63]), .B(b[22]), .Z(n15075) );
  XNOR U16052 ( .A(n15070), .B(n15069), .Z(n15076) );
  NANDN U16053 ( .A(n15075), .B(n15076), .Z(n15071) );
  AND U16054 ( .A(n15072), .B(n15071), .Z(n15073) );
  NOR U16055 ( .A(n15074), .B(n15073), .Z(n24740) );
  NOR U16056 ( .A(n24739), .B(n24740), .Z(n24750) );
  XNOR U16057 ( .A(n15074), .B(n15073), .Z(n24737) );
  XNOR U16058 ( .A(n15076), .B(n15075), .Z(n15764) );
  AND U16059 ( .A(a[63]), .B(b[21]), .Z(n15418) );
  NAND U16060 ( .A(a[62]), .B(b[21]), .Z(n15413) );
  AND U16061 ( .A(a[61]), .B(b[21]), .Z(n15406) );
  NAND U16062 ( .A(a[60]), .B(b[21]), .Z(n15401) );
  AND U16063 ( .A(a[59]), .B(b[21]), .Z(n15394) );
  NAND U16064 ( .A(a[58]), .B(b[21]), .Z(n15389) );
  AND U16065 ( .A(a[57]), .B(b[21]), .Z(n15382) );
  NAND U16066 ( .A(a[56]), .B(b[21]), .Z(n15377) );
  AND U16067 ( .A(a[55]), .B(b[21]), .Z(n15370) );
  NAND U16068 ( .A(a[54]), .B(b[21]), .Z(n15365) );
  AND U16069 ( .A(a[53]), .B(b[21]), .Z(n15358) );
  NAND U16070 ( .A(a[52]), .B(b[21]), .Z(n15353) );
  AND U16071 ( .A(a[51]), .B(b[21]), .Z(n15346) );
  NAND U16072 ( .A(a[50]), .B(b[21]), .Z(n15341) );
  AND U16073 ( .A(a[49]), .B(b[21]), .Z(n15334) );
  NAND U16074 ( .A(a[48]), .B(b[21]), .Z(n15329) );
  AND U16075 ( .A(a[47]), .B(b[21]), .Z(n15322) );
  NAND U16076 ( .A(a[46]), .B(b[21]), .Z(n15317) );
  NAND U16077 ( .A(a[45]), .B(b[21]), .Z(n15443) );
  XNOR U16078 ( .A(n15078), .B(n15077), .Z(n15682) );
  AND U16079 ( .A(a[44]), .B(b[21]), .Z(n15681) );
  NAND U16080 ( .A(a[42]), .B(b[21]), .Z(n15303) );
  XNOR U16081 ( .A(n15080), .B(n15079), .Z(n15659) );
  XNOR U16082 ( .A(n15082), .B(n15081), .Z(n15651) );
  XNOR U16083 ( .A(n15084), .B(n15083), .Z(n15640) );
  XNOR U16084 ( .A(n15086), .B(n15085), .Z(n15630) );
  XNOR U16085 ( .A(n15088), .B(n15087), .Z(n15624) );
  XNOR U16086 ( .A(n15090), .B(n15089), .Z(n15614) );
  XNOR U16087 ( .A(n15092), .B(n15091), .Z(n15603) );
  XNOR U16088 ( .A(n15094), .B(n15093), .Z(n15595) );
  NAND U16089 ( .A(a[24]), .B(b[21]), .Z(n15228) );
  AND U16090 ( .A(a[22]), .B(b[21]), .Z(n15213) );
  IV U16091 ( .A(n15213), .Z(n15458) );
  NAND U16092 ( .A(a[20]), .B(b[21]), .Z(n15462) );
  IV U16093 ( .A(n15462), .Z(n15202) );
  XOR U16094 ( .A(n15098), .B(n15097), .Z(n15099) );
  XNOR U16095 ( .A(n15100), .B(n15099), .Z(n15572) );
  XNOR U16096 ( .A(n15102), .B(n15101), .Z(n15562) );
  AND U16097 ( .A(a[4]), .B(b[21]), .Z(n15122) );
  AND U16098 ( .A(b[21]), .B(a[0]), .Z(n15801) );
  AND U16099 ( .A(a[1]), .B(b[22]), .Z(n15108) );
  AND U16100 ( .A(n15801), .B(n15108), .Z(n15105) );
  NAND U16101 ( .A(a[2]), .B(n15105), .Z(n15112) );
  NAND U16102 ( .A(b[22]), .B(a[1]), .Z(n15106) );
  XOR U16103 ( .A(n15107), .B(n15106), .Z(n15480) );
  NAND U16104 ( .A(n15108), .B(a[0]), .Z(n15109) );
  XNOR U16105 ( .A(a[2]), .B(n15109), .Z(n15110) );
  AND U16106 ( .A(b[21]), .B(n15110), .Z(n15481) );
  NANDN U16107 ( .A(n15480), .B(n15481), .Z(n15111) );
  AND U16108 ( .A(n15112), .B(n15111), .Z(n15116) );
  XNOR U16109 ( .A(n15114), .B(n15113), .Z(n15115) );
  NANDN U16110 ( .A(n15116), .B(n15115), .Z(n15118) );
  NAND U16111 ( .A(a[3]), .B(b[21]), .Z(n15488) );
  XNOR U16112 ( .A(n15116), .B(n15115), .Z(n15489) );
  NANDN U16113 ( .A(n15488), .B(n15489), .Z(n15117) );
  AND U16114 ( .A(n15118), .B(n15117), .Z(n15121) );
  NANDN U16115 ( .A(n15122), .B(n15121), .Z(n15124) );
  XOR U16116 ( .A(n15120), .B(n15119), .Z(n15471) );
  XNOR U16117 ( .A(n15122), .B(n15121), .Z(n15470) );
  NANDN U16118 ( .A(n15471), .B(n15470), .Z(n15123) );
  AND U16119 ( .A(n15124), .B(n15123), .Z(n15128) );
  XOR U16120 ( .A(n15126), .B(n15125), .Z(n15127) );
  NAND U16121 ( .A(n15128), .B(n15127), .Z(n15130) );
  NAND U16122 ( .A(a[5]), .B(b[21]), .Z(n15496) );
  XOR U16123 ( .A(n15128), .B(n15127), .Z(n15497) );
  NANDN U16124 ( .A(n15496), .B(n15497), .Z(n15129) );
  AND U16125 ( .A(n15130), .B(n15129), .Z(n15134) );
  XNOR U16126 ( .A(n15132), .B(n15131), .Z(n15133) );
  NANDN U16127 ( .A(n15134), .B(n15133), .Z(n15136) );
  NAND U16128 ( .A(a[6]), .B(b[21]), .Z(n15502) );
  XNOR U16129 ( .A(n15134), .B(n15133), .Z(n15503) );
  NANDN U16130 ( .A(n15502), .B(n15503), .Z(n15135) );
  AND U16131 ( .A(n15136), .B(n15135), .Z(n15140) );
  XNOR U16132 ( .A(n15138), .B(n15137), .Z(n15139) );
  NANDN U16133 ( .A(n15140), .B(n15139), .Z(n15142) );
  XNOR U16134 ( .A(n15140), .B(n15139), .Z(n15509) );
  AND U16135 ( .A(a[7]), .B(b[21]), .Z(n15508) );
  NAND U16136 ( .A(n15509), .B(n15508), .Z(n15141) );
  AND U16137 ( .A(n15142), .B(n15141), .Z(n15144) );
  AND U16138 ( .A(a[8]), .B(b[21]), .Z(n15143) );
  NANDN U16139 ( .A(n15144), .B(n15143), .Z(n15148) );
  XNOR U16140 ( .A(n15144), .B(n15143), .Z(n15515) );
  XNOR U16141 ( .A(n15146), .B(n15145), .Z(n15514) );
  NAND U16142 ( .A(n15515), .B(n15514), .Z(n15147) );
  NAND U16143 ( .A(n15148), .B(n15147), .Z(n15149) );
  NAND U16144 ( .A(n15150), .B(n15149), .Z(n15152) );
  NAND U16145 ( .A(a[9]), .B(b[21]), .Z(n15522) );
  XOR U16146 ( .A(n15150), .B(n15149), .Z(n15523) );
  NANDN U16147 ( .A(n15522), .B(n15523), .Z(n15151) );
  AND U16148 ( .A(n15152), .B(n15151), .Z(n15156) );
  AND U16149 ( .A(a[10]), .B(b[21]), .Z(n15155) );
  NANDN U16150 ( .A(n15156), .B(n15155), .Z(n15158) );
  XNOR U16151 ( .A(n15156), .B(n15155), .Z(n15526) );
  NAND U16152 ( .A(n15527), .B(n15526), .Z(n15157) );
  AND U16153 ( .A(n15158), .B(n15157), .Z(n15162) );
  XOR U16154 ( .A(n15160), .B(n15159), .Z(n15161) );
  NANDN U16155 ( .A(n15162), .B(n15161), .Z(n15164) );
  NAND U16156 ( .A(a[11]), .B(b[21]), .Z(n15534) );
  XNOR U16157 ( .A(n15162), .B(n15161), .Z(n15535) );
  NANDN U16158 ( .A(n15534), .B(n15535), .Z(n15163) );
  AND U16159 ( .A(n15164), .B(n15163), .Z(n15168) );
  AND U16160 ( .A(a[12]), .B(b[21]), .Z(n15167) );
  NANDN U16161 ( .A(n15168), .B(n15167), .Z(n15170) );
  XNOR U16162 ( .A(n15168), .B(n15167), .Z(n15538) );
  NAND U16163 ( .A(n15539), .B(n15538), .Z(n15169) );
  AND U16164 ( .A(n15170), .B(n15169), .Z(n15174) );
  XOR U16165 ( .A(n15172), .B(n15171), .Z(n15173) );
  NANDN U16166 ( .A(n15174), .B(n15173), .Z(n15176) );
  NAND U16167 ( .A(a[13]), .B(b[21]), .Z(n15546) );
  XNOR U16168 ( .A(n15174), .B(n15173), .Z(n15547) );
  NANDN U16169 ( .A(n15546), .B(n15547), .Z(n15175) );
  AND U16170 ( .A(n15176), .B(n15175), .Z(n15180) );
  AND U16171 ( .A(a[14]), .B(b[21]), .Z(n15179) );
  NANDN U16172 ( .A(n15180), .B(n15179), .Z(n15182) );
  XNOR U16173 ( .A(n15180), .B(n15179), .Z(n15550) );
  NAND U16174 ( .A(n15551), .B(n15550), .Z(n15181) );
  AND U16175 ( .A(n15182), .B(n15181), .Z(n15186) );
  XOR U16176 ( .A(n15184), .B(n15183), .Z(n15185) );
  NANDN U16177 ( .A(n15186), .B(n15185), .Z(n15188) );
  NAND U16178 ( .A(a[15]), .B(b[21]), .Z(n15558) );
  XNOR U16179 ( .A(n15186), .B(n15185), .Z(n15559) );
  NANDN U16180 ( .A(n15558), .B(n15559), .Z(n15187) );
  AND U16181 ( .A(n15188), .B(n15187), .Z(n15192) );
  AND U16182 ( .A(a[16]), .B(b[21]), .Z(n15191) );
  NANDN U16183 ( .A(n15192), .B(n15191), .Z(n15194) );
  XOR U16184 ( .A(n15190), .B(n15189), .Z(n15469) );
  XNOR U16185 ( .A(n15192), .B(n15191), .Z(n15468) );
  NAND U16186 ( .A(n15469), .B(n15468), .Z(n15193) );
  NAND U16187 ( .A(n15194), .B(n15193), .Z(n15563) );
  NAND U16188 ( .A(a[17]), .B(b[21]), .Z(n15565) );
  AND U16189 ( .A(a[18]), .B(b[21]), .Z(n15198) );
  NANDN U16190 ( .A(n15199), .B(n15198), .Z(n15201) );
  XNOR U16191 ( .A(n15199), .B(n15198), .Z(n15466) );
  NAND U16192 ( .A(n15467), .B(n15466), .Z(n15200) );
  NAND U16193 ( .A(n15201), .B(n15200), .Z(n15573) );
  NAND U16194 ( .A(a[19]), .B(b[21]), .Z(n15575) );
  NANDN U16195 ( .A(n15202), .B(n15463), .Z(n15208) );
  NOR U16196 ( .A(n15462), .B(n15463), .Z(n15206) );
  OR U16197 ( .A(n15206), .B(n15465), .Z(n15207) );
  AND U16198 ( .A(n15208), .B(n15207), .Z(n15578) );
  XOR U16199 ( .A(n15210), .B(n15209), .Z(n15211) );
  XOR U16200 ( .A(n15212), .B(n15211), .Z(n15579) );
  AND U16201 ( .A(a[21]), .B(b[21]), .Z(n15581) );
  NANDN U16202 ( .A(n15458), .B(n15459), .Z(n15219) );
  NOR U16203 ( .A(n15213), .B(n15459), .Z(n15217) );
  OR U16204 ( .A(n15217), .B(n15461), .Z(n15218) );
  AND U16205 ( .A(n15219), .B(n15218), .Z(n15587) );
  NANDN U16206 ( .A(n15220), .B(n15587), .Z(n15223) );
  IV U16207 ( .A(n15220), .Z(n15588) );
  NOR U16208 ( .A(n15588), .B(n15587), .Z(n15221) );
  NAND U16209 ( .A(a[23]), .B(b[21]), .Z(n15586) );
  NANDN U16210 ( .A(n15221), .B(n15586), .Z(n15222) );
  AND U16211 ( .A(n15223), .B(n15222), .Z(n15229) );
  NANDN U16212 ( .A(n15228), .B(n15229), .Z(n15231) );
  XNOR U16213 ( .A(n15225), .B(n15224), .Z(n15226) );
  XNOR U16214 ( .A(n15227), .B(n15226), .Z(n15590) );
  NAND U16215 ( .A(n15590), .B(n15589), .Z(n15230) );
  NAND U16216 ( .A(n15231), .B(n15230), .Z(n15596) );
  NAND U16217 ( .A(a[25]), .B(b[21]), .Z(n15598) );
  AND U16218 ( .A(a[26]), .B(b[21]), .Z(n15236) );
  NANDN U16219 ( .A(n15237), .B(n15236), .Z(n15239) );
  XNOR U16220 ( .A(n15233), .B(n15232), .Z(n15234) );
  XNOR U16221 ( .A(n15235), .B(n15234), .Z(n15457) );
  XNOR U16222 ( .A(n15237), .B(n15236), .Z(n15456) );
  NAND U16223 ( .A(n15457), .B(n15456), .Z(n15238) );
  NAND U16224 ( .A(n15239), .B(n15238), .Z(n15604) );
  NAND U16225 ( .A(a[27]), .B(b[21]), .Z(n15606) );
  AND U16226 ( .A(a[28]), .B(b[21]), .Z(n15240) );
  NANDN U16227 ( .A(n15241), .B(n15240), .Z(n15247) );
  XOR U16228 ( .A(n15241), .B(n15240), .Z(n15611) );
  XNOR U16229 ( .A(n15243), .B(n15242), .Z(n15244) );
  XNOR U16230 ( .A(n15245), .B(n15244), .Z(n15612) );
  NANDN U16231 ( .A(n15611), .B(n15612), .Z(n15246) );
  NAND U16232 ( .A(n15247), .B(n15246), .Z(n15615) );
  NAND U16233 ( .A(a[29]), .B(b[21]), .Z(n15617) );
  AND U16234 ( .A(a[30]), .B(b[21]), .Z(n15252) );
  NANDN U16235 ( .A(n15253), .B(n15252), .Z(n15255) );
  XNOR U16236 ( .A(n15249), .B(n15248), .Z(n15250) );
  XNOR U16237 ( .A(n15251), .B(n15250), .Z(n15455) );
  XNOR U16238 ( .A(n15253), .B(n15252), .Z(n15454) );
  NAND U16239 ( .A(n15455), .B(n15454), .Z(n15254) );
  NAND U16240 ( .A(n15255), .B(n15254), .Z(n15625) );
  NAND U16241 ( .A(a[31]), .B(b[21]), .Z(n15627) );
  AND U16242 ( .A(a[32]), .B(b[21]), .Z(n15260) );
  NANDN U16243 ( .A(n15261), .B(n15260), .Z(n15263) );
  XNOR U16244 ( .A(n15257), .B(n15256), .Z(n15258) );
  XNOR U16245 ( .A(n15259), .B(n15258), .Z(n15453) );
  XNOR U16246 ( .A(n15261), .B(n15260), .Z(n15452) );
  NAND U16247 ( .A(n15453), .B(n15452), .Z(n15262) );
  NAND U16248 ( .A(n15263), .B(n15262), .Z(n15631) );
  NAND U16249 ( .A(a[33]), .B(b[21]), .Z(n15633) );
  AND U16250 ( .A(a[34]), .B(b[21]), .Z(n15268) );
  NANDN U16251 ( .A(n15269), .B(n15268), .Z(n15271) );
  XNOR U16252 ( .A(n15265), .B(n15264), .Z(n15266) );
  XNOR U16253 ( .A(n15267), .B(n15266), .Z(n15451) );
  XNOR U16254 ( .A(n15269), .B(n15268), .Z(n15450) );
  NAND U16255 ( .A(n15451), .B(n15450), .Z(n15270) );
  NAND U16256 ( .A(n15271), .B(n15270), .Z(n15641) );
  NAND U16257 ( .A(a[35]), .B(b[21]), .Z(n15643) );
  AND U16258 ( .A(a[36]), .B(b[21]), .Z(n15272) );
  NANDN U16259 ( .A(n15273), .B(n15272), .Z(n15279) );
  XOR U16260 ( .A(n15273), .B(n15272), .Z(n15646) );
  XOR U16261 ( .A(n15275), .B(n15274), .Z(n15276) );
  XNOR U16262 ( .A(n15277), .B(n15276), .Z(n15647) );
  NANDN U16263 ( .A(n15646), .B(n15647), .Z(n15278) );
  NAND U16264 ( .A(n15279), .B(n15278), .Z(n15652) );
  NAND U16265 ( .A(a[37]), .B(b[21]), .Z(n15654) );
  AND U16266 ( .A(a[38]), .B(b[21]), .Z(n15280) );
  NANDN U16267 ( .A(n15281), .B(n15280), .Z(n15287) );
  XNOR U16268 ( .A(n15281), .B(n15280), .Z(n15449) );
  XNOR U16269 ( .A(n15283), .B(n15282), .Z(n15284) );
  XNOR U16270 ( .A(n15285), .B(n15284), .Z(n15448) );
  NAND U16271 ( .A(n15449), .B(n15448), .Z(n15286) );
  NAND U16272 ( .A(n15287), .B(n15286), .Z(n15660) );
  NAND U16273 ( .A(a[39]), .B(b[21]), .Z(n15662) );
  AND U16274 ( .A(a[40]), .B(b[21]), .Z(n15288) );
  NANDN U16275 ( .A(n15289), .B(n15288), .Z(n15295) );
  XOR U16276 ( .A(n15289), .B(n15288), .Z(n15665) );
  XNOR U16277 ( .A(n15291), .B(n15290), .Z(n15292) );
  XNOR U16278 ( .A(n15293), .B(n15292), .Z(n15666) );
  NANDN U16279 ( .A(n15665), .B(n15666), .Z(n15294) );
  AND U16280 ( .A(n15295), .B(n15294), .Z(n15671) );
  IV U16281 ( .A(n15298), .Z(n15672) );
  NAND U16282 ( .A(a[41]), .B(b[21]), .Z(n15670) );
  NANDN U16283 ( .A(n15303), .B(n15304), .Z(n15306) );
  XNOR U16284 ( .A(n15300), .B(n15299), .Z(n15301) );
  XNOR U16285 ( .A(n15302), .B(n15301), .Z(n15447) );
  NAND U16286 ( .A(n15447), .B(n15446), .Z(n15305) );
  AND U16287 ( .A(n15306), .B(n15305), .Z(n15309) );
  NANDN U16288 ( .A(n15309), .B(n15310), .Z(n15312) );
  AND U16289 ( .A(a[43]), .B(b[21]), .Z(n15676) );
  NAND U16290 ( .A(n15676), .B(n15675), .Z(n15311) );
  NAND U16291 ( .A(n15312), .B(n15311), .Z(n15684) );
  XOR U16292 ( .A(n15314), .B(n15313), .Z(n15445) );
  NANDN U16293 ( .A(n15317), .B(n15318), .Z(n15320) );
  XOR U16294 ( .A(n15316), .B(n15315), .Z(n15693) );
  XNOR U16295 ( .A(n15318), .B(n15317), .Z(n15694) );
  NANDN U16296 ( .A(n15693), .B(n15694), .Z(n15319) );
  AND U16297 ( .A(n15320), .B(n15319), .Z(n15321) );
  NANDN U16298 ( .A(n15322), .B(n15321), .Z(n15326) );
  XOR U16299 ( .A(n15322), .B(n15321), .Z(n15440) );
  XOR U16300 ( .A(n15324), .B(n15323), .Z(n15441) );
  NANDN U16301 ( .A(n15440), .B(n15441), .Z(n15325) );
  AND U16302 ( .A(n15326), .B(n15325), .Z(n15330) );
  NANDN U16303 ( .A(n15329), .B(n15330), .Z(n15332) );
  XOR U16304 ( .A(n15328), .B(n15327), .Z(n15701) );
  XNOR U16305 ( .A(n15330), .B(n15329), .Z(n15702) );
  NANDN U16306 ( .A(n15701), .B(n15702), .Z(n15331) );
  AND U16307 ( .A(n15332), .B(n15331), .Z(n15333) );
  NANDN U16308 ( .A(n15334), .B(n15333), .Z(n15338) );
  XOR U16309 ( .A(n15334), .B(n15333), .Z(n15438) );
  XOR U16310 ( .A(n15336), .B(n15335), .Z(n15439) );
  NANDN U16311 ( .A(n15438), .B(n15439), .Z(n15337) );
  AND U16312 ( .A(n15338), .B(n15337), .Z(n15342) );
  NANDN U16313 ( .A(n15341), .B(n15342), .Z(n15344) );
  XOR U16314 ( .A(n15340), .B(n15339), .Z(n15709) );
  XNOR U16315 ( .A(n15342), .B(n15341), .Z(n15710) );
  NANDN U16316 ( .A(n15709), .B(n15710), .Z(n15343) );
  AND U16317 ( .A(n15344), .B(n15343), .Z(n15345) );
  NANDN U16318 ( .A(n15346), .B(n15345), .Z(n15350) );
  XOR U16319 ( .A(n15346), .B(n15345), .Z(n15436) );
  XOR U16320 ( .A(n15348), .B(n15347), .Z(n15437) );
  NANDN U16321 ( .A(n15436), .B(n15437), .Z(n15349) );
  AND U16322 ( .A(n15350), .B(n15349), .Z(n15354) );
  NANDN U16323 ( .A(n15353), .B(n15354), .Z(n15356) );
  XOR U16324 ( .A(n15352), .B(n15351), .Z(n15717) );
  XNOR U16325 ( .A(n15354), .B(n15353), .Z(n15718) );
  NANDN U16326 ( .A(n15717), .B(n15718), .Z(n15355) );
  AND U16327 ( .A(n15356), .B(n15355), .Z(n15357) );
  NANDN U16328 ( .A(n15358), .B(n15357), .Z(n15362) );
  XOR U16329 ( .A(n15358), .B(n15357), .Z(n15434) );
  XOR U16330 ( .A(n15360), .B(n15359), .Z(n15435) );
  NANDN U16331 ( .A(n15434), .B(n15435), .Z(n15361) );
  AND U16332 ( .A(n15362), .B(n15361), .Z(n15366) );
  NANDN U16333 ( .A(n15365), .B(n15366), .Z(n15368) );
  XOR U16334 ( .A(n15364), .B(n15363), .Z(n15725) );
  XNOR U16335 ( .A(n15366), .B(n15365), .Z(n15726) );
  NANDN U16336 ( .A(n15725), .B(n15726), .Z(n15367) );
  AND U16337 ( .A(n15368), .B(n15367), .Z(n15369) );
  NANDN U16338 ( .A(n15370), .B(n15369), .Z(n15374) );
  XOR U16339 ( .A(n15370), .B(n15369), .Z(n15432) );
  XOR U16340 ( .A(n15372), .B(n15371), .Z(n15433) );
  NANDN U16341 ( .A(n15432), .B(n15433), .Z(n15373) );
  AND U16342 ( .A(n15374), .B(n15373), .Z(n15378) );
  NANDN U16343 ( .A(n15377), .B(n15378), .Z(n15380) );
  XOR U16344 ( .A(n15376), .B(n15375), .Z(n15733) );
  XNOR U16345 ( .A(n15378), .B(n15377), .Z(n15734) );
  NANDN U16346 ( .A(n15733), .B(n15734), .Z(n15379) );
  AND U16347 ( .A(n15380), .B(n15379), .Z(n15381) );
  NANDN U16348 ( .A(n15382), .B(n15381), .Z(n15386) );
  XOR U16349 ( .A(n15382), .B(n15381), .Z(n15430) );
  XOR U16350 ( .A(n15384), .B(n15383), .Z(n15431) );
  NANDN U16351 ( .A(n15430), .B(n15431), .Z(n15385) );
  AND U16352 ( .A(n15386), .B(n15385), .Z(n15390) );
  NANDN U16353 ( .A(n15389), .B(n15390), .Z(n15392) );
  XOR U16354 ( .A(n15388), .B(n15387), .Z(n15741) );
  XNOR U16355 ( .A(n15390), .B(n15389), .Z(n15742) );
  NANDN U16356 ( .A(n15741), .B(n15742), .Z(n15391) );
  AND U16357 ( .A(n15392), .B(n15391), .Z(n15393) );
  NANDN U16358 ( .A(n15394), .B(n15393), .Z(n15398) );
  XOR U16359 ( .A(n15394), .B(n15393), .Z(n15428) );
  XOR U16360 ( .A(n15396), .B(n15395), .Z(n15429) );
  NANDN U16361 ( .A(n15428), .B(n15429), .Z(n15397) );
  AND U16362 ( .A(n15398), .B(n15397), .Z(n15402) );
  NANDN U16363 ( .A(n15401), .B(n15402), .Z(n15404) );
  XOR U16364 ( .A(n15400), .B(n15399), .Z(n15749) );
  XNOR U16365 ( .A(n15402), .B(n15401), .Z(n15750) );
  NANDN U16366 ( .A(n15749), .B(n15750), .Z(n15403) );
  AND U16367 ( .A(n15404), .B(n15403), .Z(n15405) );
  NANDN U16368 ( .A(n15406), .B(n15405), .Z(n15410) );
  XOR U16369 ( .A(n15406), .B(n15405), .Z(n15426) );
  XOR U16370 ( .A(n15408), .B(n15407), .Z(n15427) );
  NANDN U16371 ( .A(n15426), .B(n15427), .Z(n15409) );
  AND U16372 ( .A(n15410), .B(n15409), .Z(n15414) );
  NANDN U16373 ( .A(n15413), .B(n15414), .Z(n15416) );
  XOR U16374 ( .A(n15412), .B(n15411), .Z(n15757) );
  XNOR U16375 ( .A(n15414), .B(n15413), .Z(n15758) );
  NANDN U16376 ( .A(n15757), .B(n15758), .Z(n15415) );
  AND U16377 ( .A(n15416), .B(n15415), .Z(n15417) );
  NANDN U16378 ( .A(n15418), .B(n15417), .Z(n15422) );
  XOR U16379 ( .A(n15418), .B(n15417), .Z(n15424) );
  XOR U16380 ( .A(n15420), .B(n15419), .Z(n15425) );
  OR U16381 ( .A(n15424), .B(n15425), .Z(n15421) );
  AND U16382 ( .A(n15422), .B(n15421), .Z(n15763) );
  AND U16383 ( .A(n15764), .B(n15763), .Z(n15423) );
  IV U16384 ( .A(n15423), .Z(n24738) );
  NANDN U16385 ( .A(n15423), .B(n24737), .Z(n24744) );
  XOR U16386 ( .A(n15425), .B(n15424), .Z(n16114) );
  XOR U16387 ( .A(n15427), .B(n15426), .Z(n15756) );
  AND U16388 ( .A(a[62]), .B(b[20]), .Z(n15755) );
  XOR U16389 ( .A(n15429), .B(n15428), .Z(n15748) );
  AND U16390 ( .A(a[60]), .B(b[20]), .Z(n15747) );
  XOR U16391 ( .A(n15431), .B(n15430), .Z(n15740) );
  AND U16392 ( .A(a[58]), .B(b[20]), .Z(n15739) );
  XOR U16393 ( .A(n15433), .B(n15432), .Z(n15732) );
  AND U16394 ( .A(a[56]), .B(b[20]), .Z(n15731) );
  XOR U16395 ( .A(n15435), .B(n15434), .Z(n15724) );
  AND U16396 ( .A(a[54]), .B(b[20]), .Z(n15723) );
  XOR U16397 ( .A(n15437), .B(n15436), .Z(n15716) );
  AND U16398 ( .A(a[52]), .B(b[20]), .Z(n15715) );
  XOR U16399 ( .A(n15439), .B(n15438), .Z(n15708) );
  AND U16400 ( .A(a[50]), .B(b[20]), .Z(n15707) );
  XOR U16401 ( .A(n15441), .B(n15440), .Z(n15700) );
  AND U16402 ( .A(a[48]), .B(b[20]), .Z(n15699) );
  NAND U16403 ( .A(a[46]), .B(b[20]), .Z(n15689) );
  XOR U16404 ( .A(n15443), .B(n15442), .Z(n15444) );
  XNOR U16405 ( .A(n15445), .B(n15444), .Z(n15690) );
  NANDN U16406 ( .A(n15689), .B(n15690), .Z(n15692) );
  XNOR U16407 ( .A(n15447), .B(n15446), .Z(n16001) );
  NAND U16408 ( .A(a[42]), .B(b[20]), .Z(n15668) );
  XNOR U16409 ( .A(n15449), .B(n15448), .Z(n15985) );
  NAND U16410 ( .A(a[38]), .B(b[20]), .Z(n15649) );
  XNOR U16411 ( .A(n15451), .B(n15450), .Z(n15968) );
  XNOR U16412 ( .A(n15453), .B(n15452), .Z(n15962) );
  XNOR U16413 ( .A(n15455), .B(n15454), .Z(n15952) );
  NAND U16414 ( .A(a[30]), .B(b[20]), .Z(n15618) );
  XNOR U16415 ( .A(n15457), .B(n15456), .Z(n15937) );
  NAND U16416 ( .A(a[26]), .B(b[20]), .Z(n15599) );
  NAND U16417 ( .A(a[24]), .B(b[20]), .Z(n15922) );
  XOR U16418 ( .A(n15459), .B(n15458), .Z(n15460) );
  XOR U16419 ( .A(n15461), .B(n15460), .Z(n15582) );
  IV U16420 ( .A(n15582), .Z(n15915) );
  NAND U16421 ( .A(a[22]), .B(b[20]), .Z(n15788) );
  XOR U16422 ( .A(n15463), .B(n15462), .Z(n15464) );
  XNOR U16423 ( .A(n15465), .B(n15464), .Z(n15905) );
  XNOR U16424 ( .A(n15467), .B(n15466), .Z(n15897) );
  XNOR U16425 ( .A(n15469), .B(n15468), .Z(n15891) );
  AND U16426 ( .A(a[8]), .B(b[20]), .Z(n15511) );
  XOR U16427 ( .A(n15471), .B(n15470), .Z(n15493) );
  AND U16428 ( .A(b[20]), .B(a[0]), .Z(n16166) );
  AND U16429 ( .A(a[1]), .B(b[21]), .Z(n15475) );
  AND U16430 ( .A(n16166), .B(n15475), .Z(n15472) );
  NAND U16431 ( .A(a[2]), .B(n15472), .Z(n15479) );
  NAND U16432 ( .A(b[21]), .B(a[1]), .Z(n15473) );
  XOR U16433 ( .A(n15474), .B(n15473), .Z(n15807) );
  NAND U16434 ( .A(n15475), .B(a[0]), .Z(n15476) );
  XNOR U16435 ( .A(a[2]), .B(n15476), .Z(n15477) );
  AND U16436 ( .A(b[20]), .B(n15477), .Z(n15808) );
  NANDN U16437 ( .A(n15807), .B(n15808), .Z(n15478) );
  AND U16438 ( .A(n15479), .B(n15478), .Z(n15483) );
  XNOR U16439 ( .A(n15481), .B(n15480), .Z(n15482) );
  NANDN U16440 ( .A(n15483), .B(n15482), .Z(n15485) );
  XNOR U16441 ( .A(n15483), .B(n15482), .Z(n15814) );
  AND U16442 ( .A(a[3]), .B(b[20]), .Z(n15813) );
  NAND U16443 ( .A(n15814), .B(n15813), .Z(n15484) );
  AND U16444 ( .A(n15485), .B(n15484), .Z(n15487) );
  AND U16445 ( .A(a[4]), .B(b[20]), .Z(n15486) );
  NANDN U16446 ( .A(n15487), .B(n15486), .Z(n15491) );
  XNOR U16447 ( .A(n15487), .B(n15486), .Z(n15820) );
  XNOR U16448 ( .A(n15489), .B(n15488), .Z(n15819) );
  NAND U16449 ( .A(n15820), .B(n15819), .Z(n15490) );
  NAND U16450 ( .A(n15491), .B(n15490), .Z(n15492) );
  NAND U16451 ( .A(n15493), .B(n15492), .Z(n15495) );
  NAND U16452 ( .A(a[5]), .B(b[20]), .Z(n15825) );
  XOR U16453 ( .A(n15493), .B(n15492), .Z(n15826) );
  NANDN U16454 ( .A(n15825), .B(n15826), .Z(n15494) );
  AND U16455 ( .A(n15495), .B(n15494), .Z(n15499) );
  XNOR U16456 ( .A(n15497), .B(n15496), .Z(n15498) );
  NANDN U16457 ( .A(n15499), .B(n15498), .Z(n15501) );
  NAND U16458 ( .A(a[6]), .B(b[20]), .Z(n15831) );
  XNOR U16459 ( .A(n15499), .B(n15498), .Z(n15832) );
  NANDN U16460 ( .A(n15831), .B(n15832), .Z(n15500) );
  AND U16461 ( .A(n15501), .B(n15500), .Z(n15505) );
  XNOR U16462 ( .A(n15503), .B(n15502), .Z(n15504) );
  NANDN U16463 ( .A(n15505), .B(n15504), .Z(n15507) );
  NAND U16464 ( .A(a[7]), .B(b[20]), .Z(n15839) );
  XNOR U16465 ( .A(n15505), .B(n15504), .Z(n15840) );
  NANDN U16466 ( .A(n15839), .B(n15840), .Z(n15506) );
  AND U16467 ( .A(n15507), .B(n15506), .Z(n15510) );
  NANDN U16468 ( .A(n15511), .B(n15510), .Z(n15513) );
  XOR U16469 ( .A(n15509), .B(n15508), .Z(n15798) );
  XNOR U16470 ( .A(n15511), .B(n15510), .Z(n15797) );
  NANDN U16471 ( .A(n15798), .B(n15797), .Z(n15512) );
  AND U16472 ( .A(n15513), .B(n15512), .Z(n15517) );
  XOR U16473 ( .A(n15515), .B(n15514), .Z(n15516) );
  NAND U16474 ( .A(n15517), .B(n15516), .Z(n15519) );
  NAND U16475 ( .A(a[9]), .B(b[20]), .Z(n15847) );
  XOR U16476 ( .A(n15517), .B(n15516), .Z(n15848) );
  NANDN U16477 ( .A(n15847), .B(n15848), .Z(n15518) );
  AND U16478 ( .A(n15519), .B(n15518), .Z(n15521) );
  AND U16479 ( .A(a[10]), .B(b[20]), .Z(n15520) );
  NANDN U16480 ( .A(n15521), .B(n15520), .Z(n15525) );
  XNOR U16481 ( .A(n15521), .B(n15520), .Z(n15854) );
  XNOR U16482 ( .A(n15523), .B(n15522), .Z(n15853) );
  NAND U16483 ( .A(n15854), .B(n15853), .Z(n15524) );
  AND U16484 ( .A(n15525), .B(n15524), .Z(n15529) );
  XOR U16485 ( .A(n15527), .B(n15526), .Z(n15528) );
  NANDN U16486 ( .A(n15529), .B(n15528), .Z(n15531) );
  NAND U16487 ( .A(a[11]), .B(b[20]), .Z(n15859) );
  XNOR U16488 ( .A(n15529), .B(n15528), .Z(n15860) );
  NANDN U16489 ( .A(n15859), .B(n15860), .Z(n15530) );
  AND U16490 ( .A(n15531), .B(n15530), .Z(n15533) );
  AND U16491 ( .A(a[12]), .B(b[20]), .Z(n15532) );
  NANDN U16492 ( .A(n15533), .B(n15532), .Z(n15537) );
  XNOR U16493 ( .A(n15533), .B(n15532), .Z(n15866) );
  XNOR U16494 ( .A(n15535), .B(n15534), .Z(n15865) );
  NAND U16495 ( .A(n15866), .B(n15865), .Z(n15536) );
  AND U16496 ( .A(n15537), .B(n15536), .Z(n15541) );
  XOR U16497 ( .A(n15539), .B(n15538), .Z(n15540) );
  NANDN U16498 ( .A(n15541), .B(n15540), .Z(n15543) );
  NAND U16499 ( .A(a[13]), .B(b[20]), .Z(n15871) );
  XNOR U16500 ( .A(n15541), .B(n15540), .Z(n15872) );
  NANDN U16501 ( .A(n15871), .B(n15872), .Z(n15542) );
  AND U16502 ( .A(n15543), .B(n15542), .Z(n15545) );
  AND U16503 ( .A(a[14]), .B(b[20]), .Z(n15544) );
  NANDN U16504 ( .A(n15545), .B(n15544), .Z(n15549) );
  XNOR U16505 ( .A(n15545), .B(n15544), .Z(n15878) );
  XNOR U16506 ( .A(n15547), .B(n15546), .Z(n15877) );
  NAND U16507 ( .A(n15878), .B(n15877), .Z(n15548) );
  AND U16508 ( .A(n15549), .B(n15548), .Z(n15553) );
  XOR U16509 ( .A(n15551), .B(n15550), .Z(n15552) );
  NANDN U16510 ( .A(n15553), .B(n15552), .Z(n15555) );
  NAND U16511 ( .A(a[15]), .B(b[20]), .Z(n15883) );
  XNOR U16512 ( .A(n15553), .B(n15552), .Z(n15884) );
  NANDN U16513 ( .A(n15883), .B(n15884), .Z(n15554) );
  AND U16514 ( .A(n15555), .B(n15554), .Z(n15557) );
  AND U16515 ( .A(a[16]), .B(b[20]), .Z(n15556) );
  NANDN U16516 ( .A(n15557), .B(n15556), .Z(n15561) );
  XNOR U16517 ( .A(n15557), .B(n15556), .Z(n15796) );
  XNOR U16518 ( .A(n15559), .B(n15558), .Z(n15795) );
  NAND U16519 ( .A(n15796), .B(n15795), .Z(n15560) );
  NAND U16520 ( .A(n15561), .B(n15560), .Z(n15892) );
  NAND U16521 ( .A(a[17]), .B(b[20]), .Z(n15894) );
  AND U16522 ( .A(a[18]), .B(b[20]), .Z(n15567) );
  NANDN U16523 ( .A(n15566), .B(n15567), .Z(n15569) );
  XNOR U16524 ( .A(n15563), .B(n15562), .Z(n15564) );
  XNOR U16525 ( .A(n15565), .B(n15564), .Z(n15794) );
  XNOR U16526 ( .A(n15567), .B(n15566), .Z(n15793) );
  NAND U16527 ( .A(n15794), .B(n15793), .Z(n15568) );
  NAND U16528 ( .A(n15569), .B(n15568), .Z(n15898) );
  NAND U16529 ( .A(a[19]), .B(b[20]), .Z(n15900) );
  AND U16530 ( .A(a[20]), .B(b[20]), .Z(n15571) );
  NANDN U16531 ( .A(n15570), .B(n15571), .Z(n15577) );
  XOR U16532 ( .A(n15571), .B(n15570), .Z(n15791) );
  XNOR U16533 ( .A(n15573), .B(n15572), .Z(n15574) );
  XNOR U16534 ( .A(n15575), .B(n15574), .Z(n15792) );
  NANDN U16535 ( .A(n15791), .B(n15792), .Z(n15576) );
  NAND U16536 ( .A(n15577), .B(n15576), .Z(n15906) );
  NAND U16537 ( .A(a[21]), .B(b[20]), .Z(n15908) );
  XOR U16538 ( .A(n15579), .B(n15578), .Z(n15580) );
  XNOR U16539 ( .A(n15581), .B(n15580), .Z(n15790) );
  NANDN U16540 ( .A(n15915), .B(n15914), .Z(n15585) );
  NOR U16541 ( .A(n15582), .B(n15914), .Z(n15583) );
  NAND U16542 ( .A(a[23]), .B(b[20]), .Z(n15917) );
  OR U16543 ( .A(n15583), .B(n15917), .Z(n15584) );
  AND U16544 ( .A(n15585), .B(n15584), .Z(n15921) );
  XOR U16545 ( .A(n15590), .B(n15589), .Z(n15591) );
  OR U16546 ( .A(n15929), .B(n15591), .Z(n15594) );
  AND U16547 ( .A(a[25]), .B(b[20]), .Z(n15932) );
  IV U16548 ( .A(n15591), .Z(n15930) );
  ANDN U16549 ( .B(n15929), .A(n15930), .Z(n15592) );
  OR U16550 ( .A(n15932), .B(n15592), .Z(n15593) );
  AND U16551 ( .A(n15594), .B(n15593), .Z(n15600) );
  NANDN U16552 ( .A(n15599), .B(n15600), .Z(n15602) );
  XNOR U16553 ( .A(n15596), .B(n15595), .Z(n15597) );
  XNOR U16554 ( .A(n15598), .B(n15597), .Z(n15786) );
  NAND U16555 ( .A(n15786), .B(n15785), .Z(n15601) );
  NAND U16556 ( .A(n15602), .B(n15601), .Z(n15938) );
  NAND U16557 ( .A(a[27]), .B(b[20]), .Z(n15940) );
  AND U16558 ( .A(a[28]), .B(b[20]), .Z(n15608) );
  NANDN U16559 ( .A(n15607), .B(n15608), .Z(n15610) );
  XNOR U16560 ( .A(n15604), .B(n15603), .Z(n15605) );
  XNOR U16561 ( .A(n15606), .B(n15605), .Z(n15784) );
  XNOR U16562 ( .A(n15608), .B(n15607), .Z(n15783) );
  NAND U16563 ( .A(n15784), .B(n15783), .Z(n15609) );
  AND U16564 ( .A(n15610), .B(n15609), .Z(n15948) );
  IV U16565 ( .A(n15613), .Z(n15949) );
  NAND U16566 ( .A(a[29]), .B(b[20]), .Z(n15947) );
  NANDN U16567 ( .A(n15618), .B(n15619), .Z(n15621) );
  XNOR U16568 ( .A(n15615), .B(n15614), .Z(n15616) );
  XNOR U16569 ( .A(n15617), .B(n15616), .Z(n15782) );
  NAND U16570 ( .A(n15782), .B(n15781), .Z(n15620) );
  NAND U16571 ( .A(n15621), .B(n15620), .Z(n15953) );
  NAND U16572 ( .A(a[31]), .B(b[20]), .Z(n15955) );
  AND U16573 ( .A(a[32]), .B(b[20]), .Z(n15623) );
  NANDN U16574 ( .A(n15622), .B(n15623), .Z(n15629) );
  XNOR U16575 ( .A(n15623), .B(n15622), .Z(n15780) );
  XNOR U16576 ( .A(n15625), .B(n15624), .Z(n15626) );
  XNOR U16577 ( .A(n15627), .B(n15626), .Z(n15779) );
  NAND U16578 ( .A(n15780), .B(n15779), .Z(n15628) );
  NAND U16579 ( .A(n15629), .B(n15628), .Z(n15963) );
  NAND U16580 ( .A(a[33]), .B(b[20]), .Z(n15965) );
  AND U16581 ( .A(a[34]), .B(b[20]), .Z(n15635) );
  NANDN U16582 ( .A(n15634), .B(n15635), .Z(n15637) );
  XNOR U16583 ( .A(n15631), .B(n15630), .Z(n15632) );
  XNOR U16584 ( .A(n15633), .B(n15632), .Z(n15778) );
  XNOR U16585 ( .A(n15635), .B(n15634), .Z(n15777) );
  NAND U16586 ( .A(n15778), .B(n15777), .Z(n15636) );
  NAND U16587 ( .A(n15637), .B(n15636), .Z(n15969) );
  NAND U16588 ( .A(a[35]), .B(b[20]), .Z(n15971) );
  AND U16589 ( .A(a[36]), .B(b[20]), .Z(n15639) );
  NANDN U16590 ( .A(n15638), .B(n15639), .Z(n15645) );
  XNOR U16591 ( .A(n15639), .B(n15638), .Z(n15776) );
  XNOR U16592 ( .A(n15641), .B(n15640), .Z(n15642) );
  XNOR U16593 ( .A(n15643), .B(n15642), .Z(n15775) );
  NAND U16594 ( .A(n15776), .B(n15775), .Z(n15644) );
  AND U16595 ( .A(n15645), .B(n15644), .Z(n15979) );
  IV U16596 ( .A(n15648), .Z(n15980) );
  NAND U16597 ( .A(a[37]), .B(b[20]), .Z(n15978) );
  NANDN U16598 ( .A(n15649), .B(n15650), .Z(n15656) );
  XNOR U16599 ( .A(n15652), .B(n15651), .Z(n15653) );
  XNOR U16600 ( .A(n15654), .B(n15653), .Z(n15983) );
  NAND U16601 ( .A(n15984), .B(n15983), .Z(n15655) );
  NAND U16602 ( .A(n15656), .B(n15655), .Z(n15986) );
  NAND U16603 ( .A(a[39]), .B(b[20]), .Z(n15988) );
  AND U16604 ( .A(a[40]), .B(b[20]), .Z(n15658) );
  NANDN U16605 ( .A(n15657), .B(n15658), .Z(n15664) );
  XOR U16606 ( .A(n15658), .B(n15657), .Z(n15773) );
  XNOR U16607 ( .A(n15660), .B(n15659), .Z(n15661) );
  XNOR U16608 ( .A(n15662), .B(n15661), .Z(n15774) );
  NANDN U16609 ( .A(n15773), .B(n15774), .Z(n15663) );
  AND U16610 ( .A(n15664), .B(n15663), .Z(n15993) );
  IV U16611 ( .A(n15667), .Z(n15994) );
  AND U16612 ( .A(a[41]), .B(b[20]), .Z(n15996) );
  NANDN U16613 ( .A(n15668), .B(n15669), .Z(n15674) );
  NAND U16614 ( .A(n15772), .B(n15771), .Z(n15673) );
  NAND U16615 ( .A(n15674), .B(n15673), .Z(n16002) );
  NAND U16616 ( .A(a[43]), .B(b[20]), .Z(n16004) );
  AND U16617 ( .A(a[44]), .B(b[20]), .Z(n15677) );
  NANDN U16618 ( .A(n15678), .B(n15677), .Z(n15680) );
  XOR U16619 ( .A(n15676), .B(n15675), .Z(n15770) );
  XNOR U16620 ( .A(n15678), .B(n15677), .Z(n15769) );
  NAND U16621 ( .A(n15770), .B(n15769), .Z(n15679) );
  AND U16622 ( .A(n15680), .B(n15679), .Z(n15686) );
  AND U16623 ( .A(a[45]), .B(b[20]), .Z(n15685) );
  NANDN U16624 ( .A(n15686), .B(n15685), .Z(n15688) );
  XOR U16625 ( .A(n15682), .B(n15681), .Z(n15683) );
  XOR U16626 ( .A(n15684), .B(n15683), .Z(n15768) );
  XNOR U16627 ( .A(n15686), .B(n15685), .Z(n15767) );
  NANDN U16628 ( .A(n15768), .B(n15767), .Z(n15687) );
  AND U16629 ( .A(n15688), .B(n15687), .Z(n16014) );
  XNOR U16630 ( .A(n15690), .B(n15689), .Z(n16013) );
  NANDN U16631 ( .A(n16014), .B(n16013), .Z(n15691) );
  AND U16632 ( .A(n15692), .B(n15691), .Z(n15696) );
  XNOR U16633 ( .A(n15694), .B(n15693), .Z(n15695) );
  NANDN U16634 ( .A(n15696), .B(n15695), .Z(n15698) );
  NAND U16635 ( .A(a[47]), .B(b[20]), .Z(n16019) );
  XNOR U16636 ( .A(n15696), .B(n15695), .Z(n16020) );
  NANDN U16637 ( .A(n16019), .B(n16020), .Z(n15697) );
  AND U16638 ( .A(n15698), .B(n15697), .Z(n16026) );
  XOR U16639 ( .A(n15700), .B(n15699), .Z(n16025) );
  XNOR U16640 ( .A(n15702), .B(n15701), .Z(n15703) );
  NANDN U16641 ( .A(n15704), .B(n15703), .Z(n15706) );
  NAND U16642 ( .A(a[49]), .B(b[20]), .Z(n16027) );
  XNOR U16643 ( .A(n15704), .B(n15703), .Z(n16028) );
  NANDN U16644 ( .A(n16027), .B(n16028), .Z(n15705) );
  AND U16645 ( .A(n15706), .B(n15705), .Z(n16036) );
  XOR U16646 ( .A(n15708), .B(n15707), .Z(n16035) );
  XNOR U16647 ( .A(n15710), .B(n15709), .Z(n15711) );
  NANDN U16648 ( .A(n15712), .B(n15711), .Z(n15714) );
  NAND U16649 ( .A(a[51]), .B(b[20]), .Z(n16039) );
  XNOR U16650 ( .A(n15712), .B(n15711), .Z(n16040) );
  NANDN U16651 ( .A(n16039), .B(n16040), .Z(n15713) );
  AND U16652 ( .A(n15714), .B(n15713), .Z(n16048) );
  XOR U16653 ( .A(n15716), .B(n15715), .Z(n16047) );
  XNOR U16654 ( .A(n15718), .B(n15717), .Z(n15719) );
  NANDN U16655 ( .A(n15720), .B(n15719), .Z(n15722) );
  NAND U16656 ( .A(a[53]), .B(b[20]), .Z(n16051) );
  XNOR U16657 ( .A(n15720), .B(n15719), .Z(n16052) );
  NANDN U16658 ( .A(n16051), .B(n16052), .Z(n15721) );
  AND U16659 ( .A(n15722), .B(n15721), .Z(n16060) );
  XOR U16660 ( .A(n15724), .B(n15723), .Z(n16059) );
  XNOR U16661 ( .A(n15726), .B(n15725), .Z(n15727) );
  NANDN U16662 ( .A(n15728), .B(n15727), .Z(n15730) );
  NAND U16663 ( .A(a[55]), .B(b[20]), .Z(n16063) );
  XNOR U16664 ( .A(n15728), .B(n15727), .Z(n16064) );
  NANDN U16665 ( .A(n16063), .B(n16064), .Z(n15729) );
  AND U16666 ( .A(n15730), .B(n15729), .Z(n16072) );
  XOR U16667 ( .A(n15732), .B(n15731), .Z(n16071) );
  XNOR U16668 ( .A(n15734), .B(n15733), .Z(n15735) );
  NANDN U16669 ( .A(n15736), .B(n15735), .Z(n15738) );
  NAND U16670 ( .A(a[57]), .B(b[20]), .Z(n16075) );
  XNOR U16671 ( .A(n15736), .B(n15735), .Z(n16076) );
  NANDN U16672 ( .A(n16075), .B(n16076), .Z(n15737) );
  AND U16673 ( .A(n15738), .B(n15737), .Z(n16084) );
  XOR U16674 ( .A(n15740), .B(n15739), .Z(n16083) );
  XNOR U16675 ( .A(n15742), .B(n15741), .Z(n15743) );
  NANDN U16676 ( .A(n15744), .B(n15743), .Z(n15746) );
  NAND U16677 ( .A(a[59]), .B(b[20]), .Z(n16087) );
  XNOR U16678 ( .A(n15744), .B(n15743), .Z(n16088) );
  NANDN U16679 ( .A(n16087), .B(n16088), .Z(n15745) );
  AND U16680 ( .A(n15746), .B(n15745), .Z(n16096) );
  XOR U16681 ( .A(n15748), .B(n15747), .Z(n16095) );
  XNOR U16682 ( .A(n15750), .B(n15749), .Z(n15751) );
  NANDN U16683 ( .A(n15752), .B(n15751), .Z(n15754) );
  NAND U16684 ( .A(a[61]), .B(b[20]), .Z(n16099) );
  XNOR U16685 ( .A(n15752), .B(n15751), .Z(n16100) );
  NANDN U16686 ( .A(n16099), .B(n16100), .Z(n15753) );
  AND U16687 ( .A(n15754), .B(n15753), .Z(n16108) );
  XOR U16688 ( .A(n15756), .B(n15755), .Z(n16107) );
  XNOR U16689 ( .A(n15758), .B(n15757), .Z(n15759) );
  NANDN U16690 ( .A(n15760), .B(n15759), .Z(n15762) );
  NAND U16691 ( .A(a[63]), .B(b[20]), .Z(n16111) );
  XNOR U16692 ( .A(n15760), .B(n15759), .Z(n16112) );
  NANDN U16693 ( .A(n16111), .B(n16112), .Z(n15761) );
  AND U16694 ( .A(n15762), .B(n15761), .Z(n16113) );
  NOR U16695 ( .A(n16114), .B(n16113), .Z(n15766) );
  XNOR U16696 ( .A(n15764), .B(n15763), .Z(n15765) );
  NANDN U16697 ( .A(n15766), .B(n15765), .Z(n22519) );
  XNOR U16698 ( .A(n15766), .B(n15765), .Z(n24736) );
  AND U16699 ( .A(a[63]), .B(b[19]), .Z(n16106) );
  NAND U16700 ( .A(a[62]), .B(b[19]), .Z(n16101) );
  AND U16701 ( .A(a[61]), .B(b[19]), .Z(n16094) );
  NAND U16702 ( .A(a[60]), .B(b[19]), .Z(n16089) );
  AND U16703 ( .A(a[59]), .B(b[19]), .Z(n16082) );
  NAND U16704 ( .A(a[58]), .B(b[19]), .Z(n16077) );
  AND U16705 ( .A(a[57]), .B(b[19]), .Z(n16070) );
  NAND U16706 ( .A(a[56]), .B(b[19]), .Z(n16065) );
  AND U16707 ( .A(a[55]), .B(b[19]), .Z(n16058) );
  NAND U16708 ( .A(a[54]), .B(b[19]), .Z(n16053) );
  AND U16709 ( .A(a[53]), .B(b[19]), .Z(n16046) );
  NAND U16710 ( .A(a[52]), .B(b[19]), .Z(n16041) );
  AND U16711 ( .A(a[51]), .B(b[19]), .Z(n16034) );
  NAND U16712 ( .A(a[47]), .B(b[19]), .Z(n16015) );
  AND U16713 ( .A(a[46]), .B(b[19]), .Z(n16386) );
  XOR U16714 ( .A(n15768), .B(n15767), .Z(n16385) );
  XOR U16715 ( .A(n15770), .B(n15769), .Z(n16009) );
  XNOR U16716 ( .A(n15772), .B(n15771), .Z(n16374) );
  AND U16717 ( .A(a[42]), .B(b[19]), .Z(n15997) );
  NAND U16718 ( .A(a[40]), .B(b[19]), .Z(n15989) );
  XNOR U16719 ( .A(n15776), .B(n15775), .Z(n16340) );
  XNOR U16720 ( .A(n15778), .B(n15777), .Z(n16330) );
  XNOR U16721 ( .A(n15780), .B(n15779), .Z(n16322) );
  XNOR U16722 ( .A(n15782), .B(n15781), .Z(n16314) );
  XNOR U16723 ( .A(n15784), .B(n15783), .Z(n16310) );
  XOR U16724 ( .A(n15786), .B(n15785), .Z(n15933) );
  IV U16725 ( .A(n15933), .Z(n16301) );
  NAND U16726 ( .A(a[26]), .B(b[19]), .Z(n16293) );
  XOR U16727 ( .A(n15788), .B(n15787), .Z(n15789) );
  XNOR U16728 ( .A(n15790), .B(n15789), .Z(n16281) );
  NAND U16729 ( .A(a[22]), .B(b[19]), .Z(n15909) );
  XNOR U16730 ( .A(n15794), .B(n15793), .Z(n16262) );
  XNOR U16731 ( .A(n15796), .B(n15795), .Z(n16256) );
  XOR U16732 ( .A(n15798), .B(n15797), .Z(n15844) );
  AND U16733 ( .A(a[4]), .B(b[19]), .Z(n15816) );
  AND U16734 ( .A(b[19]), .B(a[0]), .Z(n16503) );
  AND U16735 ( .A(a[1]), .B(b[20]), .Z(n15802) );
  AND U16736 ( .A(n16503), .B(n15802), .Z(n15799) );
  NAND U16737 ( .A(a[2]), .B(n15799), .Z(n15806) );
  NAND U16738 ( .A(b[20]), .B(a[1]), .Z(n15800) );
  XOR U16739 ( .A(n15801), .B(n15800), .Z(n16172) );
  NAND U16740 ( .A(n15802), .B(a[0]), .Z(n15803) );
  XNOR U16741 ( .A(a[2]), .B(n15803), .Z(n15804) );
  AND U16742 ( .A(b[19]), .B(n15804), .Z(n16173) );
  NANDN U16743 ( .A(n16172), .B(n16173), .Z(n15805) );
  AND U16744 ( .A(n15806), .B(n15805), .Z(n15810) );
  XNOR U16745 ( .A(n15808), .B(n15807), .Z(n15809) );
  NANDN U16746 ( .A(n15810), .B(n15809), .Z(n15812) );
  NAND U16747 ( .A(a[3]), .B(b[19]), .Z(n16180) );
  XNOR U16748 ( .A(n15810), .B(n15809), .Z(n16181) );
  NANDN U16749 ( .A(n16180), .B(n16181), .Z(n15811) );
  AND U16750 ( .A(n15812), .B(n15811), .Z(n15815) );
  NANDN U16751 ( .A(n15816), .B(n15815), .Z(n15818) );
  XOR U16752 ( .A(n15814), .B(n15813), .Z(n16163) );
  XNOR U16753 ( .A(n15816), .B(n15815), .Z(n16162) );
  NANDN U16754 ( .A(n16163), .B(n16162), .Z(n15817) );
  AND U16755 ( .A(n15818), .B(n15817), .Z(n15822) );
  XOR U16756 ( .A(n15820), .B(n15819), .Z(n15821) );
  NAND U16757 ( .A(n15822), .B(n15821), .Z(n15824) );
  NAND U16758 ( .A(a[5]), .B(b[19]), .Z(n16188) );
  XOR U16759 ( .A(n15822), .B(n15821), .Z(n16189) );
  NANDN U16760 ( .A(n16188), .B(n16189), .Z(n15823) );
  AND U16761 ( .A(n15824), .B(n15823), .Z(n15828) );
  XNOR U16762 ( .A(n15826), .B(n15825), .Z(n15827) );
  NANDN U16763 ( .A(n15828), .B(n15827), .Z(n15830) );
  NAND U16764 ( .A(a[6]), .B(b[19]), .Z(n16194) );
  XNOR U16765 ( .A(n15828), .B(n15827), .Z(n16195) );
  NANDN U16766 ( .A(n16194), .B(n16195), .Z(n15829) );
  AND U16767 ( .A(n15830), .B(n15829), .Z(n15834) );
  XNOR U16768 ( .A(n15832), .B(n15831), .Z(n15833) );
  NANDN U16769 ( .A(n15834), .B(n15833), .Z(n15836) );
  XNOR U16770 ( .A(n15834), .B(n15833), .Z(n16201) );
  AND U16771 ( .A(a[7]), .B(b[19]), .Z(n16200) );
  NAND U16772 ( .A(n16201), .B(n16200), .Z(n15835) );
  AND U16773 ( .A(n15836), .B(n15835), .Z(n15838) );
  AND U16774 ( .A(a[8]), .B(b[19]), .Z(n15837) );
  NANDN U16775 ( .A(n15838), .B(n15837), .Z(n15842) );
  XNOR U16776 ( .A(n15838), .B(n15837), .Z(n16207) );
  XNOR U16777 ( .A(n15840), .B(n15839), .Z(n16206) );
  NAND U16778 ( .A(n16207), .B(n16206), .Z(n15841) );
  NAND U16779 ( .A(n15842), .B(n15841), .Z(n15843) );
  NAND U16780 ( .A(n15844), .B(n15843), .Z(n15846) );
  NAND U16781 ( .A(a[9]), .B(b[19]), .Z(n16214) );
  XOR U16782 ( .A(n15844), .B(n15843), .Z(n16215) );
  NANDN U16783 ( .A(n16214), .B(n16215), .Z(n15845) );
  AND U16784 ( .A(n15846), .B(n15845), .Z(n15850) );
  AND U16785 ( .A(a[10]), .B(b[19]), .Z(n15849) );
  NANDN U16786 ( .A(n15850), .B(n15849), .Z(n15852) );
  XNOR U16787 ( .A(n15848), .B(n15847), .Z(n16219) );
  XNOR U16788 ( .A(n15850), .B(n15849), .Z(n16218) );
  NAND U16789 ( .A(n16219), .B(n16218), .Z(n15851) );
  AND U16790 ( .A(n15852), .B(n15851), .Z(n15856) );
  XOR U16791 ( .A(n15854), .B(n15853), .Z(n15855) );
  NANDN U16792 ( .A(n15856), .B(n15855), .Z(n15858) );
  NAND U16793 ( .A(a[11]), .B(b[19]), .Z(n16226) );
  XNOR U16794 ( .A(n15856), .B(n15855), .Z(n16227) );
  NANDN U16795 ( .A(n16226), .B(n16227), .Z(n15857) );
  AND U16796 ( .A(n15858), .B(n15857), .Z(n15862) );
  AND U16797 ( .A(a[12]), .B(b[19]), .Z(n15861) );
  NANDN U16798 ( .A(n15862), .B(n15861), .Z(n15864) );
  XNOR U16799 ( .A(n15860), .B(n15859), .Z(n16231) );
  XNOR U16800 ( .A(n15862), .B(n15861), .Z(n16230) );
  NAND U16801 ( .A(n16231), .B(n16230), .Z(n15863) );
  AND U16802 ( .A(n15864), .B(n15863), .Z(n15868) );
  XOR U16803 ( .A(n15866), .B(n15865), .Z(n15867) );
  NANDN U16804 ( .A(n15868), .B(n15867), .Z(n15870) );
  NAND U16805 ( .A(a[13]), .B(b[19]), .Z(n16238) );
  XNOR U16806 ( .A(n15868), .B(n15867), .Z(n16239) );
  NANDN U16807 ( .A(n16238), .B(n16239), .Z(n15869) );
  AND U16808 ( .A(n15870), .B(n15869), .Z(n15874) );
  AND U16809 ( .A(a[14]), .B(b[19]), .Z(n15873) );
  NANDN U16810 ( .A(n15874), .B(n15873), .Z(n15876) );
  XNOR U16811 ( .A(n15872), .B(n15871), .Z(n16243) );
  XNOR U16812 ( .A(n15874), .B(n15873), .Z(n16242) );
  NAND U16813 ( .A(n16243), .B(n16242), .Z(n15875) );
  AND U16814 ( .A(n15876), .B(n15875), .Z(n15880) );
  XOR U16815 ( .A(n15878), .B(n15877), .Z(n15879) );
  NANDN U16816 ( .A(n15880), .B(n15879), .Z(n15882) );
  NAND U16817 ( .A(a[15]), .B(b[19]), .Z(n16250) );
  XNOR U16818 ( .A(n15880), .B(n15879), .Z(n16251) );
  NANDN U16819 ( .A(n16250), .B(n16251), .Z(n15881) );
  AND U16820 ( .A(n15882), .B(n15881), .Z(n15886) );
  AND U16821 ( .A(a[16]), .B(b[19]), .Z(n15885) );
  NANDN U16822 ( .A(n15886), .B(n15885), .Z(n15888) );
  XNOR U16823 ( .A(n15884), .B(n15883), .Z(n16161) );
  XNOR U16824 ( .A(n15886), .B(n15885), .Z(n16160) );
  NAND U16825 ( .A(n16161), .B(n16160), .Z(n15887) );
  NAND U16826 ( .A(n15888), .B(n15887), .Z(n16257) );
  NAND U16827 ( .A(a[17]), .B(b[19]), .Z(n16259) );
  AND U16828 ( .A(a[18]), .B(b[19]), .Z(n15889) );
  NANDN U16829 ( .A(n15890), .B(n15889), .Z(n15896) );
  XOR U16830 ( .A(n15890), .B(n15889), .Z(n16158) );
  XNOR U16831 ( .A(n15892), .B(n15891), .Z(n15893) );
  XNOR U16832 ( .A(n15894), .B(n15893), .Z(n16159) );
  NANDN U16833 ( .A(n16158), .B(n16159), .Z(n15895) );
  NAND U16834 ( .A(n15896), .B(n15895), .Z(n16263) );
  NAND U16835 ( .A(a[19]), .B(b[19]), .Z(n16265) );
  AND U16836 ( .A(a[20]), .B(b[19]), .Z(n15901) );
  NANDN U16837 ( .A(n15902), .B(n15901), .Z(n15904) );
  XNOR U16838 ( .A(n15898), .B(n15897), .Z(n15899) );
  XNOR U16839 ( .A(n15900), .B(n15899), .Z(n16157) );
  XNOR U16840 ( .A(n15902), .B(n15901), .Z(n16156) );
  NAND U16841 ( .A(n16157), .B(n16156), .Z(n15903) );
  AND U16842 ( .A(n15904), .B(n15903), .Z(n16272) );
  NAND U16843 ( .A(a[21]), .B(b[19]), .Z(n16275) );
  NANDN U16844 ( .A(n15909), .B(n15910), .Z(n15912) );
  XNOR U16845 ( .A(n15906), .B(n15905), .Z(n15907) );
  XNOR U16846 ( .A(n15908), .B(n15907), .Z(n16155) );
  XNOR U16847 ( .A(n15910), .B(n15909), .Z(n16154) );
  NAND U16848 ( .A(n16155), .B(n16154), .Z(n15911) );
  NAND U16849 ( .A(n15912), .B(n15911), .Z(n16282) );
  AND U16850 ( .A(a[23]), .B(b[19]), .Z(n16280) );
  AND U16851 ( .A(a[24]), .B(b[19]), .Z(n15913) );
  IV U16852 ( .A(n15913), .Z(n16153) );
  OR U16853 ( .A(n16152), .B(n16153), .Z(n15920) );
  ANDN U16854 ( .B(n16152), .A(n15913), .Z(n15918) );
  XOR U16855 ( .A(n15915), .B(n15914), .Z(n15916) );
  XOR U16856 ( .A(n15917), .B(n15916), .Z(n16151) );
  NANDN U16857 ( .A(n15918), .B(n16151), .Z(n15919) );
  AND U16858 ( .A(n15920), .B(n15919), .Z(n16288) );
  XOR U16859 ( .A(n15922), .B(n15921), .Z(n15923) );
  XOR U16860 ( .A(n15924), .B(n15923), .Z(n15925) );
  IV U16861 ( .A(n15925), .Z(n16287) );
  OR U16862 ( .A(n16288), .B(n16287), .Z(n15928) );
  ANDN U16863 ( .B(n16288), .A(n15925), .Z(n15926) );
  AND U16864 ( .A(a[25]), .B(b[19]), .Z(n16286) );
  NANDN U16865 ( .A(n15926), .B(n16286), .Z(n15927) );
  AND U16866 ( .A(n15928), .B(n15927), .Z(n16292) );
  XOR U16867 ( .A(n15930), .B(n15929), .Z(n15931) );
  XNOR U16868 ( .A(n15932), .B(n15931), .Z(n16295) );
  NANDN U16869 ( .A(n16301), .B(n16302), .Z(n15936) );
  NOR U16870 ( .A(n15933), .B(n16302), .Z(n15934) );
  AND U16871 ( .A(a[27]), .B(b[19]), .Z(n16300) );
  NANDN U16872 ( .A(n15934), .B(n16300), .Z(n15935) );
  AND U16873 ( .A(n15936), .B(n15935), .Z(n15942) );
  AND U16874 ( .A(a[28]), .B(b[19]), .Z(n15941) );
  NANDN U16875 ( .A(n15942), .B(n15941), .Z(n15944) );
  XNOR U16876 ( .A(n15938), .B(n15937), .Z(n15939) );
  XNOR U16877 ( .A(n15940), .B(n15939), .Z(n16150) );
  XNOR U16878 ( .A(n15942), .B(n15941), .Z(n16149) );
  NAND U16879 ( .A(n16150), .B(n16149), .Z(n15943) );
  NAND U16880 ( .A(n15944), .B(n15943), .Z(n16311) );
  AND U16881 ( .A(a[29]), .B(b[19]), .Z(n16309) );
  AND U16882 ( .A(a[30]), .B(b[19]), .Z(n15945) );
  NANDN U16883 ( .A(n15946), .B(n15945), .Z(n15951) );
  XOR U16884 ( .A(n15946), .B(n15945), .Z(n16147) );
  NANDN U16885 ( .A(n16147), .B(n16148), .Z(n15950) );
  NAND U16886 ( .A(n15951), .B(n15950), .Z(n16315) );
  NAND U16887 ( .A(a[31]), .B(b[19]), .Z(n16317) );
  AND U16888 ( .A(a[32]), .B(b[19]), .Z(n15956) );
  NANDN U16889 ( .A(n15957), .B(n15956), .Z(n15959) );
  XNOR U16890 ( .A(n15953), .B(n15952), .Z(n15954) );
  XNOR U16891 ( .A(n15955), .B(n15954), .Z(n16146) );
  XNOR U16892 ( .A(n15957), .B(n15956), .Z(n16145) );
  NAND U16893 ( .A(n16146), .B(n16145), .Z(n15958) );
  NAND U16894 ( .A(n15959), .B(n15958), .Z(n16323) );
  NAND U16895 ( .A(a[33]), .B(b[19]), .Z(n16325) );
  AND U16896 ( .A(a[34]), .B(b[19]), .Z(n15960) );
  NANDN U16897 ( .A(n15961), .B(n15960), .Z(n15967) );
  XNOR U16898 ( .A(n15961), .B(n15960), .Z(n16144) );
  XNOR U16899 ( .A(n15963), .B(n15962), .Z(n15964) );
  XNOR U16900 ( .A(n15965), .B(n15964), .Z(n16143) );
  NAND U16901 ( .A(n16144), .B(n16143), .Z(n15966) );
  NAND U16902 ( .A(n15967), .B(n15966), .Z(n16331) );
  NAND U16903 ( .A(a[35]), .B(b[19]), .Z(n16333) );
  AND U16904 ( .A(a[36]), .B(b[19]), .Z(n15972) );
  NANDN U16905 ( .A(n15973), .B(n15972), .Z(n15975) );
  XNOR U16906 ( .A(n15969), .B(n15968), .Z(n15970) );
  XNOR U16907 ( .A(n15971), .B(n15970), .Z(n16142) );
  XNOR U16908 ( .A(n15973), .B(n15972), .Z(n16141) );
  NAND U16909 ( .A(n16142), .B(n16141), .Z(n15974) );
  NAND U16910 ( .A(n15975), .B(n15974), .Z(n16341) );
  NAND U16911 ( .A(a[37]), .B(b[19]), .Z(n16343) );
  AND U16912 ( .A(a[38]), .B(b[19]), .Z(n15976) );
  NANDN U16913 ( .A(n15977), .B(n15976), .Z(n15982) );
  XNOR U16914 ( .A(n15977), .B(n15976), .Z(n16140) );
  NAND U16915 ( .A(n16140), .B(n16139), .Z(n15981) );
  NAND U16916 ( .A(n15982), .B(n15981), .Z(n16346) );
  XNOR U16917 ( .A(n15984), .B(n15983), .Z(n16347) );
  NAND U16918 ( .A(a[39]), .B(b[19]), .Z(n16348) );
  NANDN U16919 ( .A(n15989), .B(n15990), .Z(n15992) );
  XNOR U16920 ( .A(n15986), .B(n15985), .Z(n15987) );
  XNOR U16921 ( .A(n15988), .B(n15987), .Z(n16354) );
  NAND U16922 ( .A(n16354), .B(n16353), .Z(n15991) );
  NAND U16923 ( .A(n15992), .B(n15991), .Z(n16360) );
  AND U16924 ( .A(a[41]), .B(b[19]), .Z(n16362) );
  NANDN U16925 ( .A(n15997), .B(n15998), .Z(n16000) );
  XOR U16926 ( .A(n15994), .B(n15993), .Z(n15995) );
  XOR U16927 ( .A(n15996), .B(n15995), .Z(n16367) );
  NANDN U16928 ( .A(n16367), .B(n16368), .Z(n15999) );
  AND U16929 ( .A(n16000), .B(n15999), .Z(n16373) );
  AND U16930 ( .A(a[43]), .B(b[19]), .Z(n16372) );
  AND U16931 ( .A(a[44]), .B(b[19]), .Z(n16005) );
  NANDN U16932 ( .A(n16006), .B(n16005), .Z(n16008) );
  XNOR U16933 ( .A(n16002), .B(n16001), .Z(n16003) );
  XNOR U16934 ( .A(n16004), .B(n16003), .Z(n16138) );
  XNOR U16935 ( .A(n16006), .B(n16005), .Z(n16137) );
  NAND U16936 ( .A(n16138), .B(n16137), .Z(n16007) );
  AND U16937 ( .A(n16008), .B(n16007), .Z(n16010) );
  NANDN U16938 ( .A(n16009), .B(n16010), .Z(n16012) );
  NAND U16939 ( .A(a[45]), .B(b[19]), .Z(n16379) );
  NAND U16940 ( .A(n16380), .B(n16379), .Z(n16011) );
  AND U16941 ( .A(n16012), .B(n16011), .Z(n16388) );
  NANDN U16942 ( .A(n16015), .B(n16016), .Z(n16018) );
  XOR U16943 ( .A(n16014), .B(n16013), .Z(n16135) );
  XNOR U16944 ( .A(n16016), .B(n16015), .Z(n16136) );
  NANDN U16945 ( .A(n16135), .B(n16136), .Z(n16017) );
  AND U16946 ( .A(n16018), .B(n16017), .Z(n16022) );
  AND U16947 ( .A(a[48]), .B(b[19]), .Z(n16021) );
  NANDN U16948 ( .A(n16022), .B(n16021), .Z(n16024) );
  XOR U16949 ( .A(n16020), .B(n16019), .Z(n16395) );
  XNOR U16950 ( .A(n16022), .B(n16021), .Z(n16396) );
  NANDN U16951 ( .A(n16395), .B(n16396), .Z(n16023) );
  AND U16952 ( .A(n16024), .B(n16023), .Z(n16132) );
  NAND U16953 ( .A(a[49]), .B(b[19]), .Z(n16131) );
  XOR U16954 ( .A(n16026), .B(n16025), .Z(n16134) );
  AND U16955 ( .A(a[50]), .B(b[19]), .Z(n16029) );
  NANDN U16956 ( .A(n16030), .B(n16029), .Z(n16032) );
  XOR U16957 ( .A(n16028), .B(n16027), .Z(n16405) );
  XNOR U16958 ( .A(n16030), .B(n16029), .Z(n16406) );
  NANDN U16959 ( .A(n16405), .B(n16406), .Z(n16031) );
  AND U16960 ( .A(n16032), .B(n16031), .Z(n16033) );
  NANDN U16961 ( .A(n16034), .B(n16033), .Z(n16038) );
  XOR U16962 ( .A(n16034), .B(n16033), .Z(n16129) );
  XOR U16963 ( .A(n16036), .B(n16035), .Z(n16130) );
  NANDN U16964 ( .A(n16129), .B(n16130), .Z(n16037) );
  AND U16965 ( .A(n16038), .B(n16037), .Z(n16042) );
  NANDN U16966 ( .A(n16041), .B(n16042), .Z(n16044) );
  XOR U16967 ( .A(n16040), .B(n16039), .Z(n16413) );
  XNOR U16968 ( .A(n16042), .B(n16041), .Z(n16414) );
  NANDN U16969 ( .A(n16413), .B(n16414), .Z(n16043) );
  AND U16970 ( .A(n16044), .B(n16043), .Z(n16045) );
  NANDN U16971 ( .A(n16046), .B(n16045), .Z(n16050) );
  XOR U16972 ( .A(n16046), .B(n16045), .Z(n16127) );
  XOR U16973 ( .A(n16048), .B(n16047), .Z(n16128) );
  NANDN U16974 ( .A(n16127), .B(n16128), .Z(n16049) );
  AND U16975 ( .A(n16050), .B(n16049), .Z(n16054) );
  NANDN U16976 ( .A(n16053), .B(n16054), .Z(n16056) );
  XOR U16977 ( .A(n16052), .B(n16051), .Z(n16421) );
  XNOR U16978 ( .A(n16054), .B(n16053), .Z(n16422) );
  NANDN U16979 ( .A(n16421), .B(n16422), .Z(n16055) );
  AND U16980 ( .A(n16056), .B(n16055), .Z(n16057) );
  NANDN U16981 ( .A(n16058), .B(n16057), .Z(n16062) );
  XOR U16982 ( .A(n16058), .B(n16057), .Z(n16125) );
  XOR U16983 ( .A(n16060), .B(n16059), .Z(n16126) );
  NANDN U16984 ( .A(n16125), .B(n16126), .Z(n16061) );
  AND U16985 ( .A(n16062), .B(n16061), .Z(n16066) );
  NANDN U16986 ( .A(n16065), .B(n16066), .Z(n16068) );
  XOR U16987 ( .A(n16064), .B(n16063), .Z(n16429) );
  XNOR U16988 ( .A(n16066), .B(n16065), .Z(n16430) );
  NANDN U16989 ( .A(n16429), .B(n16430), .Z(n16067) );
  AND U16990 ( .A(n16068), .B(n16067), .Z(n16069) );
  NANDN U16991 ( .A(n16070), .B(n16069), .Z(n16074) );
  XOR U16992 ( .A(n16070), .B(n16069), .Z(n16123) );
  XOR U16993 ( .A(n16072), .B(n16071), .Z(n16124) );
  NANDN U16994 ( .A(n16123), .B(n16124), .Z(n16073) );
  AND U16995 ( .A(n16074), .B(n16073), .Z(n16078) );
  NANDN U16996 ( .A(n16077), .B(n16078), .Z(n16080) );
  XOR U16997 ( .A(n16076), .B(n16075), .Z(n16437) );
  XNOR U16998 ( .A(n16078), .B(n16077), .Z(n16438) );
  NANDN U16999 ( .A(n16437), .B(n16438), .Z(n16079) );
  AND U17000 ( .A(n16080), .B(n16079), .Z(n16081) );
  NANDN U17001 ( .A(n16082), .B(n16081), .Z(n16086) );
  XOR U17002 ( .A(n16082), .B(n16081), .Z(n16121) );
  XOR U17003 ( .A(n16084), .B(n16083), .Z(n16122) );
  NANDN U17004 ( .A(n16121), .B(n16122), .Z(n16085) );
  AND U17005 ( .A(n16086), .B(n16085), .Z(n16090) );
  NANDN U17006 ( .A(n16089), .B(n16090), .Z(n16092) );
  XOR U17007 ( .A(n16088), .B(n16087), .Z(n16445) );
  XNOR U17008 ( .A(n16090), .B(n16089), .Z(n16446) );
  NANDN U17009 ( .A(n16445), .B(n16446), .Z(n16091) );
  AND U17010 ( .A(n16092), .B(n16091), .Z(n16093) );
  NANDN U17011 ( .A(n16094), .B(n16093), .Z(n16098) );
  XOR U17012 ( .A(n16094), .B(n16093), .Z(n16119) );
  XOR U17013 ( .A(n16096), .B(n16095), .Z(n16120) );
  NANDN U17014 ( .A(n16119), .B(n16120), .Z(n16097) );
  AND U17015 ( .A(n16098), .B(n16097), .Z(n16102) );
  NANDN U17016 ( .A(n16101), .B(n16102), .Z(n16104) );
  XOR U17017 ( .A(n16100), .B(n16099), .Z(n16453) );
  XNOR U17018 ( .A(n16102), .B(n16101), .Z(n16454) );
  NANDN U17019 ( .A(n16453), .B(n16454), .Z(n16103) );
  AND U17020 ( .A(n16104), .B(n16103), .Z(n16105) );
  NANDN U17021 ( .A(n16106), .B(n16105), .Z(n16110) );
  XOR U17022 ( .A(n16106), .B(n16105), .Z(n16117) );
  XOR U17023 ( .A(n16108), .B(n16107), .Z(n16118) );
  NANDN U17024 ( .A(n16117), .B(n16118), .Z(n16109) );
  AND U17025 ( .A(n16110), .B(n16109), .Z(n16460) );
  XNOR U17026 ( .A(n16112), .B(n16111), .Z(n16459) );
  AND U17027 ( .A(n16460), .B(n16459), .Z(n16116) );
  XNOR U17028 ( .A(n16114), .B(n16113), .Z(n16115) );
  NANDN U17029 ( .A(n16116), .B(n16115), .Z(n22517) );
  XNOR U17030 ( .A(n16116), .B(n16115), .Z(n24734) );
  XOR U17031 ( .A(n16118), .B(n16117), .Z(n16804) );
  XOR U17032 ( .A(n16120), .B(n16119), .Z(n16452) );
  XOR U17033 ( .A(n16122), .B(n16121), .Z(n16444) );
  AND U17034 ( .A(a[60]), .B(b[18]), .Z(n16443) );
  XOR U17035 ( .A(n16124), .B(n16123), .Z(n16436) );
  AND U17036 ( .A(a[58]), .B(b[18]), .Z(n16435) );
  XOR U17037 ( .A(n16126), .B(n16125), .Z(n16428) );
  AND U17038 ( .A(a[56]), .B(b[18]), .Z(n16427) );
  XOR U17039 ( .A(n16128), .B(n16127), .Z(n16420) );
  AND U17040 ( .A(a[54]), .B(b[18]), .Z(n16419) );
  XOR U17041 ( .A(n16130), .B(n16129), .Z(n16412) );
  AND U17042 ( .A(a[52]), .B(b[18]), .Z(n16411) );
  NAND U17043 ( .A(a[50]), .B(b[18]), .Z(n16401) );
  XOR U17044 ( .A(n16132), .B(n16131), .Z(n16133) );
  XNOR U17045 ( .A(n16134), .B(n16133), .Z(n16402) );
  NANDN U17046 ( .A(n16401), .B(n16402), .Z(n16404) );
  NAND U17047 ( .A(a[48]), .B(b[18]), .Z(n16391) );
  XNOR U17048 ( .A(n16136), .B(n16135), .Z(n16392) );
  NANDN U17049 ( .A(n16391), .B(n16392), .Z(n16394) );
  XNOR U17050 ( .A(n16138), .B(n16137), .Z(n16703) );
  AND U17051 ( .A(a[42]), .B(b[18]), .Z(n16363) );
  XNOR U17052 ( .A(n16140), .B(n16139), .Z(n16676) );
  XNOR U17053 ( .A(n16142), .B(n16141), .Z(n16668) );
  XNOR U17054 ( .A(n16144), .B(n16143), .Z(n16660) );
  XNOR U17055 ( .A(n16146), .B(n16145), .Z(n16652) );
  NAND U17056 ( .A(a[32]), .B(b[18]), .Z(n16318) );
  AND U17057 ( .A(a[30]), .B(b[18]), .Z(n16307) );
  XOR U17058 ( .A(n16150), .B(n16149), .Z(n16303) );
  IV U17059 ( .A(n16303), .Z(n16640) );
  NAND U17060 ( .A(a[28]), .B(b[18]), .Z(n16482) );
  AND U17061 ( .A(a[24]), .B(b[18]), .Z(n16278) );
  XNOR U17062 ( .A(n16155), .B(n16154), .Z(n16615) );
  XNOR U17063 ( .A(n16157), .B(n16156), .Z(n16607) );
  NAND U17064 ( .A(a[20]), .B(b[18]), .Z(n16266) );
  XNOR U17065 ( .A(n16159), .B(n16158), .Z(n16600) );
  XNOR U17066 ( .A(n16161), .B(n16160), .Z(n16593) );
  AND U17067 ( .A(a[8]), .B(b[18]), .Z(n16203) );
  XOR U17068 ( .A(n16163), .B(n16162), .Z(n16185) );
  AND U17069 ( .A(b[18]), .B(a[0]), .Z(n16853) );
  AND U17070 ( .A(a[1]), .B(b[19]), .Z(n16167) );
  AND U17071 ( .A(n16853), .B(n16167), .Z(n16164) );
  NAND U17072 ( .A(a[2]), .B(n16164), .Z(n16171) );
  NAND U17073 ( .A(b[19]), .B(a[1]), .Z(n16165) );
  XOR U17074 ( .A(n16166), .B(n16165), .Z(n16509) );
  NAND U17075 ( .A(n16167), .B(a[0]), .Z(n16168) );
  XNOR U17076 ( .A(a[2]), .B(n16168), .Z(n16169) );
  AND U17077 ( .A(b[18]), .B(n16169), .Z(n16510) );
  NANDN U17078 ( .A(n16509), .B(n16510), .Z(n16170) );
  AND U17079 ( .A(n16171), .B(n16170), .Z(n16175) );
  XNOR U17080 ( .A(n16173), .B(n16172), .Z(n16174) );
  NANDN U17081 ( .A(n16175), .B(n16174), .Z(n16177) );
  XNOR U17082 ( .A(n16175), .B(n16174), .Z(n16516) );
  AND U17083 ( .A(a[3]), .B(b[18]), .Z(n16515) );
  NAND U17084 ( .A(n16516), .B(n16515), .Z(n16176) );
  AND U17085 ( .A(n16177), .B(n16176), .Z(n16179) );
  AND U17086 ( .A(a[4]), .B(b[18]), .Z(n16178) );
  NANDN U17087 ( .A(n16179), .B(n16178), .Z(n16183) );
  XNOR U17088 ( .A(n16179), .B(n16178), .Z(n16522) );
  XNOR U17089 ( .A(n16181), .B(n16180), .Z(n16521) );
  NAND U17090 ( .A(n16522), .B(n16521), .Z(n16182) );
  NAND U17091 ( .A(n16183), .B(n16182), .Z(n16184) );
  NAND U17092 ( .A(n16185), .B(n16184), .Z(n16187) );
  NAND U17093 ( .A(a[5]), .B(b[18]), .Z(n16527) );
  XOR U17094 ( .A(n16185), .B(n16184), .Z(n16528) );
  NANDN U17095 ( .A(n16527), .B(n16528), .Z(n16186) );
  AND U17096 ( .A(n16187), .B(n16186), .Z(n16191) );
  XNOR U17097 ( .A(n16189), .B(n16188), .Z(n16190) );
  NANDN U17098 ( .A(n16191), .B(n16190), .Z(n16193) );
  NAND U17099 ( .A(a[6]), .B(b[18]), .Z(n16533) );
  XNOR U17100 ( .A(n16191), .B(n16190), .Z(n16534) );
  NANDN U17101 ( .A(n16533), .B(n16534), .Z(n16192) );
  AND U17102 ( .A(n16193), .B(n16192), .Z(n16197) );
  XNOR U17103 ( .A(n16195), .B(n16194), .Z(n16196) );
  NANDN U17104 ( .A(n16197), .B(n16196), .Z(n16199) );
  NAND U17105 ( .A(a[7]), .B(b[18]), .Z(n16541) );
  XNOR U17106 ( .A(n16197), .B(n16196), .Z(n16542) );
  NANDN U17107 ( .A(n16541), .B(n16542), .Z(n16198) );
  AND U17108 ( .A(n16199), .B(n16198), .Z(n16202) );
  NANDN U17109 ( .A(n16203), .B(n16202), .Z(n16205) );
  XOR U17110 ( .A(n16201), .B(n16200), .Z(n16500) );
  XNOR U17111 ( .A(n16203), .B(n16202), .Z(n16499) );
  NANDN U17112 ( .A(n16500), .B(n16499), .Z(n16204) );
  AND U17113 ( .A(n16205), .B(n16204), .Z(n16209) );
  XOR U17114 ( .A(n16207), .B(n16206), .Z(n16208) );
  NAND U17115 ( .A(n16209), .B(n16208), .Z(n16211) );
  NAND U17116 ( .A(a[9]), .B(b[18]), .Z(n16549) );
  XOR U17117 ( .A(n16209), .B(n16208), .Z(n16550) );
  NANDN U17118 ( .A(n16549), .B(n16550), .Z(n16210) );
  AND U17119 ( .A(n16211), .B(n16210), .Z(n16213) );
  AND U17120 ( .A(a[10]), .B(b[18]), .Z(n16212) );
  NANDN U17121 ( .A(n16213), .B(n16212), .Z(n16217) );
  XNOR U17122 ( .A(n16213), .B(n16212), .Z(n16556) );
  XNOR U17123 ( .A(n16215), .B(n16214), .Z(n16555) );
  NAND U17124 ( .A(n16556), .B(n16555), .Z(n16216) );
  AND U17125 ( .A(n16217), .B(n16216), .Z(n16221) );
  XOR U17126 ( .A(n16219), .B(n16218), .Z(n16220) );
  NANDN U17127 ( .A(n16221), .B(n16220), .Z(n16223) );
  NAND U17128 ( .A(a[11]), .B(b[18]), .Z(n16561) );
  XNOR U17129 ( .A(n16221), .B(n16220), .Z(n16562) );
  NANDN U17130 ( .A(n16561), .B(n16562), .Z(n16222) );
  AND U17131 ( .A(n16223), .B(n16222), .Z(n16225) );
  AND U17132 ( .A(a[12]), .B(b[18]), .Z(n16224) );
  NANDN U17133 ( .A(n16225), .B(n16224), .Z(n16229) );
  XNOR U17134 ( .A(n16225), .B(n16224), .Z(n16568) );
  XNOR U17135 ( .A(n16227), .B(n16226), .Z(n16567) );
  NAND U17136 ( .A(n16568), .B(n16567), .Z(n16228) );
  AND U17137 ( .A(n16229), .B(n16228), .Z(n16233) );
  XOR U17138 ( .A(n16231), .B(n16230), .Z(n16232) );
  NANDN U17139 ( .A(n16233), .B(n16232), .Z(n16235) );
  NAND U17140 ( .A(a[13]), .B(b[18]), .Z(n16573) );
  XNOR U17141 ( .A(n16233), .B(n16232), .Z(n16574) );
  NANDN U17142 ( .A(n16573), .B(n16574), .Z(n16234) );
  AND U17143 ( .A(n16235), .B(n16234), .Z(n16237) );
  AND U17144 ( .A(a[14]), .B(b[18]), .Z(n16236) );
  NANDN U17145 ( .A(n16237), .B(n16236), .Z(n16241) );
  XNOR U17146 ( .A(n16237), .B(n16236), .Z(n16580) );
  XNOR U17147 ( .A(n16239), .B(n16238), .Z(n16579) );
  NAND U17148 ( .A(n16580), .B(n16579), .Z(n16240) );
  AND U17149 ( .A(n16241), .B(n16240), .Z(n16245) );
  XOR U17150 ( .A(n16243), .B(n16242), .Z(n16244) );
  NANDN U17151 ( .A(n16245), .B(n16244), .Z(n16247) );
  NAND U17152 ( .A(a[15]), .B(b[18]), .Z(n16585) );
  XNOR U17153 ( .A(n16245), .B(n16244), .Z(n16586) );
  NANDN U17154 ( .A(n16585), .B(n16586), .Z(n16246) );
  AND U17155 ( .A(n16247), .B(n16246), .Z(n16249) );
  AND U17156 ( .A(a[16]), .B(b[18]), .Z(n16248) );
  NANDN U17157 ( .A(n16249), .B(n16248), .Z(n16253) );
  XNOR U17158 ( .A(n16249), .B(n16248), .Z(n16498) );
  XNOR U17159 ( .A(n16251), .B(n16250), .Z(n16497) );
  NAND U17160 ( .A(n16498), .B(n16497), .Z(n16252) );
  NAND U17161 ( .A(n16253), .B(n16252), .Z(n16594) );
  NAND U17162 ( .A(a[17]), .B(b[18]), .Z(n16596) );
  AND U17163 ( .A(a[18]), .B(b[18]), .Z(n16254) );
  NANDN U17164 ( .A(n16255), .B(n16254), .Z(n16261) );
  XOR U17165 ( .A(n16255), .B(n16254), .Z(n16495) );
  XNOR U17166 ( .A(n16257), .B(n16256), .Z(n16258) );
  XNOR U17167 ( .A(n16259), .B(n16258), .Z(n16496) );
  NANDN U17168 ( .A(n16495), .B(n16496), .Z(n16260) );
  AND U17169 ( .A(n16261), .B(n16260), .Z(n16599) );
  NAND U17170 ( .A(a[19]), .B(b[18]), .Z(n16602) );
  NANDN U17171 ( .A(n16266), .B(n16267), .Z(n16269) );
  XNOR U17172 ( .A(n16263), .B(n16262), .Z(n16264) );
  XNOR U17173 ( .A(n16265), .B(n16264), .Z(n16494) );
  XNOR U17174 ( .A(n16267), .B(n16266), .Z(n16493) );
  NAND U17175 ( .A(n16494), .B(n16493), .Z(n16268) );
  NAND U17176 ( .A(n16269), .B(n16268), .Z(n16608) );
  NAND U17177 ( .A(a[21]), .B(b[18]), .Z(n16610) );
  AND U17178 ( .A(a[22]), .B(b[18]), .Z(n16270) );
  NANDN U17179 ( .A(n16271), .B(n16270), .Z(n16277) );
  XOR U17180 ( .A(n16271), .B(n16270), .Z(n16491) );
  XNOR U17181 ( .A(n16273), .B(n16272), .Z(n16274) );
  XNOR U17182 ( .A(n16275), .B(n16274), .Z(n16492) );
  NANDN U17183 ( .A(n16491), .B(n16492), .Z(n16276) );
  NAND U17184 ( .A(n16277), .B(n16276), .Z(n16616) );
  NAND U17185 ( .A(a[23]), .B(b[18]), .Z(n16618) );
  NANDN U17186 ( .A(n16278), .B(n16279), .Z(n16284) );
  NAND U17187 ( .A(n16489), .B(n16490), .Z(n16283) );
  AND U17188 ( .A(n16284), .B(n16283), .Z(n16626) );
  AND U17189 ( .A(a[25]), .B(b[18]), .Z(n16625) );
  AND U17190 ( .A(a[26]), .B(b[18]), .Z(n16285) );
  IV U17191 ( .A(n16285), .Z(n16486) );
  OR U17192 ( .A(n16485), .B(n16486), .Z(n16291) );
  ANDN U17193 ( .B(n16485), .A(n16285), .Z(n16289) );
  OR U17194 ( .A(n16289), .B(n16488), .Z(n16290) );
  AND U17195 ( .A(n16291), .B(n16290), .Z(n16631) );
  XOR U17196 ( .A(n16293), .B(n16292), .Z(n16294) );
  XOR U17197 ( .A(n16295), .B(n16294), .Z(n16296) );
  IV U17198 ( .A(n16296), .Z(n16630) );
  OR U17199 ( .A(n16631), .B(n16630), .Z(n16299) );
  ANDN U17200 ( .B(n16631), .A(n16296), .Z(n16297) );
  NAND U17201 ( .A(a[27]), .B(b[18]), .Z(n16633) );
  OR U17202 ( .A(n16297), .B(n16633), .Z(n16298) );
  AND U17203 ( .A(n16299), .B(n16298), .Z(n16481) );
  NANDN U17204 ( .A(n16640), .B(n16639), .Z(n16306) );
  NOR U17205 ( .A(n16303), .B(n16639), .Z(n16304) );
  AND U17206 ( .A(a[29]), .B(b[18]), .Z(n16638) );
  NANDN U17207 ( .A(n16304), .B(n16638), .Z(n16305) );
  AND U17208 ( .A(n16306), .B(n16305), .Z(n16308) );
  NANDN U17209 ( .A(n16307), .B(n16308), .Z(n16313) );
  NAND U17210 ( .A(n16479), .B(n16480), .Z(n16312) );
  NAND U17211 ( .A(n16313), .B(n16312), .Z(n16648) );
  AND U17212 ( .A(a[31]), .B(b[18]), .Z(n16649) );
  NANDN U17213 ( .A(n16318), .B(n16319), .Z(n16321) );
  XNOR U17214 ( .A(n16315), .B(n16314), .Z(n16316) );
  XNOR U17215 ( .A(n16317), .B(n16316), .Z(n16478) );
  NAND U17216 ( .A(n16478), .B(n16477), .Z(n16320) );
  NAND U17217 ( .A(n16321), .B(n16320), .Z(n16653) );
  NAND U17218 ( .A(a[33]), .B(b[18]), .Z(n16655) );
  AND U17219 ( .A(a[34]), .B(b[18]), .Z(n16327) );
  NANDN U17220 ( .A(n16326), .B(n16327), .Z(n16329) );
  XNOR U17221 ( .A(n16323), .B(n16322), .Z(n16324) );
  XNOR U17222 ( .A(n16325), .B(n16324), .Z(n16476) );
  XNOR U17223 ( .A(n16327), .B(n16326), .Z(n16475) );
  NAND U17224 ( .A(n16476), .B(n16475), .Z(n16328) );
  NAND U17225 ( .A(n16329), .B(n16328), .Z(n16661) );
  NAND U17226 ( .A(a[35]), .B(b[18]), .Z(n16663) );
  AND U17227 ( .A(a[36]), .B(b[18]), .Z(n16335) );
  NANDN U17228 ( .A(n16334), .B(n16335), .Z(n16337) );
  XNOR U17229 ( .A(n16331), .B(n16330), .Z(n16332) );
  XNOR U17230 ( .A(n16333), .B(n16332), .Z(n16474) );
  XNOR U17231 ( .A(n16335), .B(n16334), .Z(n16473) );
  NAND U17232 ( .A(n16474), .B(n16473), .Z(n16336) );
  NAND U17233 ( .A(n16337), .B(n16336), .Z(n16669) );
  NAND U17234 ( .A(a[37]), .B(b[18]), .Z(n16671) );
  AND U17235 ( .A(a[38]), .B(b[18]), .Z(n16339) );
  NANDN U17236 ( .A(n16338), .B(n16339), .Z(n16345) );
  XNOR U17237 ( .A(n16339), .B(n16338), .Z(n16472) );
  XNOR U17238 ( .A(n16341), .B(n16340), .Z(n16342) );
  XNOR U17239 ( .A(n16343), .B(n16342), .Z(n16471) );
  NAND U17240 ( .A(n16472), .B(n16471), .Z(n16344) );
  NAND U17241 ( .A(n16345), .B(n16344), .Z(n16677) );
  NAND U17242 ( .A(a[39]), .B(b[18]), .Z(n16679) );
  AND U17243 ( .A(a[40]), .B(b[18]), .Z(n16350) );
  NANDN U17244 ( .A(n16349), .B(n16350), .Z(n16352) );
  XNOR U17245 ( .A(n16350), .B(n16349), .Z(n16685) );
  NANDN U17246 ( .A(n16684), .B(n16685), .Z(n16351) );
  AND U17247 ( .A(n16352), .B(n16351), .Z(n16687) );
  XOR U17248 ( .A(n16354), .B(n16353), .Z(n16355) );
  IV U17249 ( .A(n16355), .Z(n16688) );
  OR U17250 ( .A(n16687), .B(n16688), .Z(n16358) );
  ANDN U17251 ( .B(n16687), .A(n16355), .Z(n16356) );
  NAND U17252 ( .A(a[41]), .B(b[18]), .Z(n16690) );
  OR U17253 ( .A(n16356), .B(n16690), .Z(n16357) );
  AND U17254 ( .A(n16358), .B(n16357), .Z(n16364) );
  NANDN U17255 ( .A(n16363), .B(n16364), .Z(n16366) );
  XNOR U17256 ( .A(n16360), .B(n16359), .Z(n16361) );
  XOR U17257 ( .A(n16362), .B(n16361), .Z(n16469) );
  NANDN U17258 ( .A(n16469), .B(n16470), .Z(n16365) );
  AND U17259 ( .A(n16366), .B(n16365), .Z(n16697) );
  IV U17260 ( .A(n16369), .Z(n16698) );
  NAND U17261 ( .A(a[43]), .B(b[18]), .Z(n16700) );
  AND U17262 ( .A(a[44]), .B(b[18]), .Z(n16371) );
  NANDN U17263 ( .A(n16370), .B(n16371), .Z(n16376) );
  XNOR U17264 ( .A(n16371), .B(n16370), .Z(n16468) );
  NAND U17265 ( .A(n16468), .B(n16467), .Z(n16375) );
  NAND U17266 ( .A(n16376), .B(n16375), .Z(n16704) );
  NAND U17267 ( .A(a[45]), .B(b[18]), .Z(n16706) );
  AND U17268 ( .A(a[46]), .B(b[18]), .Z(n16377) );
  NANDN U17269 ( .A(n16378), .B(n16377), .Z(n16382) );
  XOR U17270 ( .A(n16378), .B(n16377), .Z(n16711) );
  XNOR U17271 ( .A(n16380), .B(n16379), .Z(n16712) );
  NANDN U17272 ( .A(n16711), .B(n16712), .Z(n16381) );
  AND U17273 ( .A(n16382), .B(n16381), .Z(n16384) );
  AND U17274 ( .A(a[47]), .B(b[18]), .Z(n16383) );
  NANDN U17275 ( .A(n16384), .B(n16383), .Z(n16390) );
  XOR U17276 ( .A(n16384), .B(n16383), .Z(n16465) );
  XOR U17277 ( .A(n16386), .B(n16385), .Z(n16387) );
  XNOR U17278 ( .A(n16388), .B(n16387), .Z(n16466) );
  NANDN U17279 ( .A(n16465), .B(n16466), .Z(n16389) );
  AND U17280 ( .A(n16390), .B(n16389), .Z(n16718) );
  XNOR U17281 ( .A(n16392), .B(n16391), .Z(n16717) );
  NANDN U17282 ( .A(n16718), .B(n16717), .Z(n16393) );
  AND U17283 ( .A(n16394), .B(n16393), .Z(n16398) );
  XNOR U17284 ( .A(n16396), .B(n16395), .Z(n16397) );
  NANDN U17285 ( .A(n16398), .B(n16397), .Z(n16400) );
  NAND U17286 ( .A(a[49]), .B(b[18]), .Z(n16723) );
  XNOR U17287 ( .A(n16398), .B(n16397), .Z(n16724) );
  NANDN U17288 ( .A(n16723), .B(n16724), .Z(n16399) );
  AND U17289 ( .A(n16400), .B(n16399), .Z(n16730) );
  XNOR U17290 ( .A(n16402), .B(n16401), .Z(n16729) );
  NANDN U17291 ( .A(n16730), .B(n16729), .Z(n16403) );
  AND U17292 ( .A(n16404), .B(n16403), .Z(n16408) );
  XNOR U17293 ( .A(n16406), .B(n16405), .Z(n16407) );
  NANDN U17294 ( .A(n16408), .B(n16407), .Z(n16410) );
  NAND U17295 ( .A(a[51]), .B(b[18]), .Z(n16735) );
  XNOR U17296 ( .A(n16408), .B(n16407), .Z(n16736) );
  NANDN U17297 ( .A(n16735), .B(n16736), .Z(n16409) );
  AND U17298 ( .A(n16410), .B(n16409), .Z(n16742) );
  XOR U17299 ( .A(n16412), .B(n16411), .Z(n16741) );
  XNOR U17300 ( .A(n16414), .B(n16413), .Z(n16415) );
  NANDN U17301 ( .A(n16416), .B(n16415), .Z(n16418) );
  NAND U17302 ( .A(a[53]), .B(b[18]), .Z(n16743) );
  XNOR U17303 ( .A(n16416), .B(n16415), .Z(n16744) );
  NANDN U17304 ( .A(n16743), .B(n16744), .Z(n16417) );
  AND U17305 ( .A(n16418), .B(n16417), .Z(n16752) );
  XOR U17306 ( .A(n16420), .B(n16419), .Z(n16751) );
  XNOR U17307 ( .A(n16422), .B(n16421), .Z(n16423) );
  NANDN U17308 ( .A(n16424), .B(n16423), .Z(n16426) );
  NAND U17309 ( .A(a[55]), .B(b[18]), .Z(n16755) );
  XNOR U17310 ( .A(n16424), .B(n16423), .Z(n16756) );
  NANDN U17311 ( .A(n16755), .B(n16756), .Z(n16425) );
  AND U17312 ( .A(n16426), .B(n16425), .Z(n16764) );
  XOR U17313 ( .A(n16428), .B(n16427), .Z(n16763) );
  XNOR U17314 ( .A(n16430), .B(n16429), .Z(n16431) );
  NANDN U17315 ( .A(n16432), .B(n16431), .Z(n16434) );
  NAND U17316 ( .A(a[57]), .B(b[18]), .Z(n16767) );
  XNOR U17317 ( .A(n16432), .B(n16431), .Z(n16768) );
  NANDN U17318 ( .A(n16767), .B(n16768), .Z(n16433) );
  AND U17319 ( .A(n16434), .B(n16433), .Z(n16776) );
  XOR U17320 ( .A(n16436), .B(n16435), .Z(n16775) );
  XNOR U17321 ( .A(n16438), .B(n16437), .Z(n16439) );
  NANDN U17322 ( .A(n16440), .B(n16439), .Z(n16442) );
  NAND U17323 ( .A(a[59]), .B(b[18]), .Z(n16779) );
  XNOR U17324 ( .A(n16440), .B(n16439), .Z(n16780) );
  NANDN U17325 ( .A(n16779), .B(n16780), .Z(n16441) );
  AND U17326 ( .A(n16442), .B(n16441), .Z(n16788) );
  XOR U17327 ( .A(n16444), .B(n16443), .Z(n16787) );
  XNOR U17328 ( .A(n16446), .B(n16445), .Z(n16447) );
  NANDN U17329 ( .A(n16448), .B(n16447), .Z(n16450) );
  NAND U17330 ( .A(a[61]), .B(b[18]), .Z(n16791) );
  XNOR U17331 ( .A(n16448), .B(n16447), .Z(n16792) );
  NANDN U17332 ( .A(n16791), .B(n16792), .Z(n16449) );
  NAND U17333 ( .A(n16450), .B(n16449), .Z(n16451) );
  XOR U17334 ( .A(n16452), .B(n16451), .Z(n16800) );
  AND U17335 ( .A(a[62]), .B(b[18]), .Z(n16799) );
  XNOR U17336 ( .A(n16454), .B(n16453), .Z(n16455) );
  NANDN U17337 ( .A(n16456), .B(n16455), .Z(n16458) );
  NAND U17338 ( .A(a[63]), .B(b[18]), .Z(n16463) );
  XNOR U17339 ( .A(n16456), .B(n16455), .Z(n16464) );
  NANDN U17340 ( .A(n16463), .B(n16464), .Z(n16457) );
  AND U17341 ( .A(n16458), .B(n16457), .Z(n16803) );
  XNOR U17342 ( .A(n16460), .B(n16459), .Z(n16461) );
  NANDN U17343 ( .A(n16462), .B(n16461), .Z(n22515) );
  XNOR U17344 ( .A(n16462), .B(n16461), .Z(n24732) );
  XNOR U17345 ( .A(n16464), .B(n16463), .Z(n17150) );
  AND U17346 ( .A(a[63]), .B(b[17]), .Z(n16798) );
  NAND U17347 ( .A(a[62]), .B(b[17]), .Z(n16793) );
  AND U17348 ( .A(a[61]), .B(b[17]), .Z(n16786) );
  NAND U17349 ( .A(a[60]), .B(b[17]), .Z(n16781) );
  AND U17350 ( .A(a[59]), .B(b[17]), .Z(n16774) );
  NAND U17351 ( .A(a[58]), .B(b[17]), .Z(n16769) );
  AND U17352 ( .A(a[57]), .B(b[17]), .Z(n16762) );
  NAND U17353 ( .A(a[56]), .B(b[17]), .Z(n16757) );
  AND U17354 ( .A(a[55]), .B(b[17]), .Z(n16750) );
  NAND U17355 ( .A(a[54]), .B(b[17]), .Z(n16745) );
  AND U17356 ( .A(a[53]), .B(b[17]), .Z(n16814) );
  NAND U17357 ( .A(a[49]), .B(b[17]), .Z(n16719) );
  AND U17358 ( .A(a[48]), .B(b[17]), .Z(n17082) );
  XOR U17359 ( .A(n16466), .B(n16465), .Z(n17081) );
  XNOR U17360 ( .A(n16468), .B(n16467), .Z(n17067) );
  NAND U17361 ( .A(a[42]), .B(b[17]), .Z(n16691) );
  XNOR U17362 ( .A(n16472), .B(n16471), .Z(n17045) );
  XNOR U17363 ( .A(n16474), .B(n16473), .Z(n17034) );
  XNOR U17364 ( .A(n16476), .B(n16475), .Z(n17024) );
  XNOR U17365 ( .A(n16478), .B(n16477), .Z(n17016) );
  XOR U17366 ( .A(n16480), .B(n16479), .Z(n16641) );
  NAND U17367 ( .A(a[30]), .B(b[17]), .Z(n17000) );
  XOR U17368 ( .A(n16482), .B(n16481), .Z(n16483) );
  XOR U17369 ( .A(n16484), .B(n16483), .Z(n16634) );
  IV U17370 ( .A(n16634), .Z(n16994) );
  NAND U17371 ( .A(a[28]), .B(b[17]), .Z(n16989) );
  XOR U17372 ( .A(n16486), .B(n16485), .Z(n16487) );
  XOR U17373 ( .A(n16488), .B(n16487), .Z(n16981) );
  XOR U17374 ( .A(n16490), .B(n16489), .Z(n16975) );
  NAND U17375 ( .A(a[24]), .B(b[17]), .Z(n16619) );
  XNOR U17376 ( .A(n16492), .B(n16491), .Z(n16966) );
  XNOR U17377 ( .A(n16494), .B(n16493), .Z(n16959) );
  NAND U17378 ( .A(a[20]), .B(b[17]), .Z(n16603) );
  XNOR U17379 ( .A(n16496), .B(n16495), .Z(n16950) );
  XNOR U17380 ( .A(n16498), .B(n16497), .Z(n16941) );
  XOR U17381 ( .A(n16500), .B(n16499), .Z(n16546) );
  AND U17382 ( .A(a[4]), .B(b[17]), .Z(n16518) );
  AND U17383 ( .A(b[17]), .B(a[0]), .Z(n17187) );
  AND U17384 ( .A(a[1]), .B(b[18]), .Z(n16504) );
  AND U17385 ( .A(n17187), .B(n16504), .Z(n16501) );
  NAND U17386 ( .A(a[2]), .B(n16501), .Z(n16508) );
  NAND U17387 ( .A(b[18]), .B(a[1]), .Z(n16502) );
  XOR U17388 ( .A(n16503), .B(n16502), .Z(n16859) );
  NAND U17389 ( .A(n16504), .B(a[0]), .Z(n16505) );
  XNOR U17390 ( .A(a[2]), .B(n16505), .Z(n16506) );
  AND U17391 ( .A(b[17]), .B(n16506), .Z(n16860) );
  NANDN U17392 ( .A(n16859), .B(n16860), .Z(n16507) );
  AND U17393 ( .A(n16508), .B(n16507), .Z(n16512) );
  XNOR U17394 ( .A(n16510), .B(n16509), .Z(n16511) );
  NANDN U17395 ( .A(n16512), .B(n16511), .Z(n16514) );
  NAND U17396 ( .A(a[3]), .B(b[17]), .Z(n16867) );
  XNOR U17397 ( .A(n16512), .B(n16511), .Z(n16868) );
  NANDN U17398 ( .A(n16867), .B(n16868), .Z(n16513) );
  AND U17399 ( .A(n16514), .B(n16513), .Z(n16517) );
  NANDN U17400 ( .A(n16518), .B(n16517), .Z(n16520) );
  XOR U17401 ( .A(n16516), .B(n16515), .Z(n16850) );
  XNOR U17402 ( .A(n16518), .B(n16517), .Z(n16849) );
  NANDN U17403 ( .A(n16850), .B(n16849), .Z(n16519) );
  AND U17404 ( .A(n16520), .B(n16519), .Z(n16524) );
  XOR U17405 ( .A(n16522), .B(n16521), .Z(n16523) );
  NAND U17406 ( .A(n16524), .B(n16523), .Z(n16526) );
  NAND U17407 ( .A(a[5]), .B(b[17]), .Z(n16875) );
  XOR U17408 ( .A(n16524), .B(n16523), .Z(n16876) );
  NANDN U17409 ( .A(n16875), .B(n16876), .Z(n16525) );
  AND U17410 ( .A(n16526), .B(n16525), .Z(n16530) );
  XNOR U17411 ( .A(n16528), .B(n16527), .Z(n16529) );
  NANDN U17412 ( .A(n16530), .B(n16529), .Z(n16532) );
  NAND U17413 ( .A(a[6]), .B(b[17]), .Z(n16881) );
  XNOR U17414 ( .A(n16530), .B(n16529), .Z(n16882) );
  NANDN U17415 ( .A(n16881), .B(n16882), .Z(n16531) );
  AND U17416 ( .A(n16532), .B(n16531), .Z(n16536) );
  XNOR U17417 ( .A(n16534), .B(n16533), .Z(n16535) );
  NANDN U17418 ( .A(n16536), .B(n16535), .Z(n16538) );
  XNOR U17419 ( .A(n16536), .B(n16535), .Z(n16888) );
  AND U17420 ( .A(a[7]), .B(b[17]), .Z(n16887) );
  NAND U17421 ( .A(n16888), .B(n16887), .Z(n16537) );
  AND U17422 ( .A(n16538), .B(n16537), .Z(n16540) );
  AND U17423 ( .A(a[8]), .B(b[17]), .Z(n16539) );
  NANDN U17424 ( .A(n16540), .B(n16539), .Z(n16544) );
  XNOR U17425 ( .A(n16540), .B(n16539), .Z(n16894) );
  XNOR U17426 ( .A(n16542), .B(n16541), .Z(n16893) );
  NAND U17427 ( .A(n16894), .B(n16893), .Z(n16543) );
  NAND U17428 ( .A(n16544), .B(n16543), .Z(n16545) );
  NAND U17429 ( .A(n16546), .B(n16545), .Z(n16548) );
  NAND U17430 ( .A(a[9]), .B(b[17]), .Z(n16901) );
  XOR U17431 ( .A(n16546), .B(n16545), .Z(n16902) );
  NANDN U17432 ( .A(n16901), .B(n16902), .Z(n16547) );
  AND U17433 ( .A(n16548), .B(n16547), .Z(n16552) );
  AND U17434 ( .A(a[10]), .B(b[17]), .Z(n16551) );
  NANDN U17435 ( .A(n16552), .B(n16551), .Z(n16554) );
  XNOR U17436 ( .A(n16550), .B(n16549), .Z(n16906) );
  XNOR U17437 ( .A(n16552), .B(n16551), .Z(n16905) );
  NAND U17438 ( .A(n16906), .B(n16905), .Z(n16553) );
  AND U17439 ( .A(n16554), .B(n16553), .Z(n16558) );
  XOR U17440 ( .A(n16556), .B(n16555), .Z(n16557) );
  NANDN U17441 ( .A(n16558), .B(n16557), .Z(n16560) );
  NAND U17442 ( .A(a[11]), .B(b[17]), .Z(n16913) );
  XNOR U17443 ( .A(n16558), .B(n16557), .Z(n16914) );
  NANDN U17444 ( .A(n16913), .B(n16914), .Z(n16559) );
  AND U17445 ( .A(n16560), .B(n16559), .Z(n16564) );
  AND U17446 ( .A(a[12]), .B(b[17]), .Z(n16563) );
  NANDN U17447 ( .A(n16564), .B(n16563), .Z(n16566) );
  XNOR U17448 ( .A(n16562), .B(n16561), .Z(n16918) );
  XNOR U17449 ( .A(n16564), .B(n16563), .Z(n16917) );
  NAND U17450 ( .A(n16918), .B(n16917), .Z(n16565) );
  AND U17451 ( .A(n16566), .B(n16565), .Z(n16570) );
  XOR U17452 ( .A(n16568), .B(n16567), .Z(n16569) );
  NANDN U17453 ( .A(n16570), .B(n16569), .Z(n16572) );
  NAND U17454 ( .A(a[13]), .B(b[17]), .Z(n16925) );
  XNOR U17455 ( .A(n16570), .B(n16569), .Z(n16926) );
  NANDN U17456 ( .A(n16925), .B(n16926), .Z(n16571) );
  AND U17457 ( .A(n16572), .B(n16571), .Z(n16576) );
  AND U17458 ( .A(a[14]), .B(b[17]), .Z(n16575) );
  NANDN U17459 ( .A(n16576), .B(n16575), .Z(n16578) );
  XNOR U17460 ( .A(n16574), .B(n16573), .Z(n16930) );
  XNOR U17461 ( .A(n16576), .B(n16575), .Z(n16929) );
  NAND U17462 ( .A(n16930), .B(n16929), .Z(n16577) );
  AND U17463 ( .A(n16578), .B(n16577), .Z(n16582) );
  XOR U17464 ( .A(n16580), .B(n16579), .Z(n16581) );
  NANDN U17465 ( .A(n16582), .B(n16581), .Z(n16584) );
  NAND U17466 ( .A(a[15]), .B(b[17]), .Z(n16937) );
  XNOR U17467 ( .A(n16582), .B(n16581), .Z(n16938) );
  NANDN U17468 ( .A(n16937), .B(n16938), .Z(n16583) );
  AND U17469 ( .A(n16584), .B(n16583), .Z(n16588) );
  AND U17470 ( .A(a[16]), .B(b[17]), .Z(n16587) );
  NANDN U17471 ( .A(n16588), .B(n16587), .Z(n16590) );
  XNOR U17472 ( .A(n16586), .B(n16585), .Z(n16848) );
  XNOR U17473 ( .A(n16588), .B(n16587), .Z(n16847) );
  NAND U17474 ( .A(n16848), .B(n16847), .Z(n16589) );
  NAND U17475 ( .A(n16590), .B(n16589), .Z(n16942) );
  NAND U17476 ( .A(a[17]), .B(b[17]), .Z(n16944) );
  AND U17477 ( .A(a[18]), .B(b[17]), .Z(n16591) );
  NANDN U17478 ( .A(n16592), .B(n16591), .Z(n16598) );
  XOR U17479 ( .A(n16592), .B(n16591), .Z(n16845) );
  XNOR U17480 ( .A(n16594), .B(n16593), .Z(n16595) );
  XNOR U17481 ( .A(n16596), .B(n16595), .Z(n16846) );
  NANDN U17482 ( .A(n16845), .B(n16846), .Z(n16597) );
  AND U17483 ( .A(n16598), .B(n16597), .Z(n16949) );
  NAND U17484 ( .A(a[19]), .B(b[17]), .Z(n16952) );
  NANDN U17485 ( .A(n16603), .B(n16604), .Z(n16606) );
  XNOR U17486 ( .A(n16600), .B(n16599), .Z(n16601) );
  XNOR U17487 ( .A(n16602), .B(n16601), .Z(n16844) );
  XNOR U17488 ( .A(n16604), .B(n16603), .Z(n16843) );
  NAND U17489 ( .A(n16844), .B(n16843), .Z(n16605) );
  NAND U17490 ( .A(n16606), .B(n16605), .Z(n16960) );
  NAND U17491 ( .A(a[21]), .B(b[17]), .Z(n16962) );
  AND U17492 ( .A(a[22]), .B(b[17]), .Z(n16611) );
  NANDN U17493 ( .A(n16612), .B(n16611), .Z(n16614) );
  XNOR U17494 ( .A(n16608), .B(n16607), .Z(n16609) );
  XNOR U17495 ( .A(n16610), .B(n16609), .Z(n16842) );
  XNOR U17496 ( .A(n16612), .B(n16611), .Z(n16841) );
  NAND U17497 ( .A(n16842), .B(n16841), .Z(n16613) );
  AND U17498 ( .A(n16614), .B(n16613), .Z(n16965) );
  NAND U17499 ( .A(a[23]), .B(b[17]), .Z(n16968) );
  NANDN U17500 ( .A(n16619), .B(n16620), .Z(n16622) );
  XNOR U17501 ( .A(n16616), .B(n16615), .Z(n16617) );
  XNOR U17502 ( .A(n16618), .B(n16617), .Z(n16840) );
  XNOR U17503 ( .A(n16620), .B(n16619), .Z(n16839) );
  NAND U17504 ( .A(n16840), .B(n16839), .Z(n16621) );
  NAND U17505 ( .A(n16622), .B(n16621), .Z(n16976) );
  AND U17506 ( .A(a[25]), .B(b[17]), .Z(n16978) );
  AND U17507 ( .A(a[26]), .B(b[17]), .Z(n16623) );
  NANDN U17508 ( .A(n16624), .B(n16623), .Z(n16629) );
  XNOR U17509 ( .A(n16624), .B(n16623), .Z(n16838) );
  NAND U17510 ( .A(n16838), .B(n16837), .Z(n16628) );
  NAND U17511 ( .A(n16629), .B(n16628), .Z(n16982) );
  NAND U17512 ( .A(a[27]), .B(b[17]), .Z(n16983) );
  XOR U17513 ( .A(n16631), .B(n16630), .Z(n16632) );
  XOR U17514 ( .A(n16633), .B(n16632), .Z(n16988) );
  NANDN U17515 ( .A(n16994), .B(n16993), .Z(n16637) );
  NOR U17516 ( .A(n16634), .B(n16993), .Z(n16635) );
  NAND U17517 ( .A(a[29]), .B(b[17]), .Z(n16996) );
  OR U17518 ( .A(n16635), .B(n16996), .Z(n16636) );
  AND U17519 ( .A(n16637), .B(n16636), .Z(n17001) );
  NANDN U17520 ( .A(n16641), .B(n17008), .Z(n16644) );
  IV U17521 ( .A(n16641), .Z(n17009) );
  NOR U17522 ( .A(n17009), .B(n17008), .Z(n16642) );
  NAND U17523 ( .A(a[31]), .B(b[17]), .Z(n17011) );
  OR U17524 ( .A(n16642), .B(n17011), .Z(n16643) );
  AND U17525 ( .A(n16644), .B(n16643), .Z(n16646) );
  AND U17526 ( .A(a[32]), .B(b[17]), .Z(n16645) );
  NANDN U17527 ( .A(n16646), .B(n16645), .Z(n16651) );
  XNOR U17528 ( .A(n16646), .B(n16645), .Z(n16836) );
  NAND U17529 ( .A(n16836), .B(n16835), .Z(n16650) );
  NAND U17530 ( .A(n16651), .B(n16650), .Z(n17017) );
  NAND U17531 ( .A(a[33]), .B(b[17]), .Z(n17019) );
  AND U17532 ( .A(a[34]), .B(b[17]), .Z(n16656) );
  NANDN U17533 ( .A(n16657), .B(n16656), .Z(n16659) );
  XNOR U17534 ( .A(n16653), .B(n16652), .Z(n16654) );
  XNOR U17535 ( .A(n16655), .B(n16654), .Z(n16834) );
  XNOR U17536 ( .A(n16657), .B(n16656), .Z(n16833) );
  NAND U17537 ( .A(n16834), .B(n16833), .Z(n16658) );
  NAND U17538 ( .A(n16659), .B(n16658), .Z(n17025) );
  NAND U17539 ( .A(a[35]), .B(b[17]), .Z(n17027) );
  AND U17540 ( .A(a[36]), .B(b[17]), .Z(n16664) );
  NANDN U17541 ( .A(n16665), .B(n16664), .Z(n16667) );
  XNOR U17542 ( .A(n16661), .B(n16660), .Z(n16662) );
  XNOR U17543 ( .A(n16663), .B(n16662), .Z(n16832) );
  XNOR U17544 ( .A(n16665), .B(n16664), .Z(n16831) );
  NAND U17545 ( .A(n16832), .B(n16831), .Z(n16666) );
  NAND U17546 ( .A(n16667), .B(n16666), .Z(n17035) );
  NAND U17547 ( .A(a[37]), .B(b[17]), .Z(n17037) );
  AND U17548 ( .A(a[38]), .B(b[17]), .Z(n16672) );
  NANDN U17549 ( .A(n16673), .B(n16672), .Z(n16675) );
  XNOR U17550 ( .A(n16669), .B(n16668), .Z(n16670) );
  XOR U17551 ( .A(n16671), .B(n16670), .Z(n17040) );
  XNOR U17552 ( .A(n16673), .B(n16672), .Z(n17041) );
  NANDN U17553 ( .A(n17040), .B(n17041), .Z(n16674) );
  NAND U17554 ( .A(n16675), .B(n16674), .Z(n17046) );
  NAND U17555 ( .A(a[39]), .B(b[17]), .Z(n17048) );
  AND U17556 ( .A(a[40]), .B(b[17]), .Z(n16680) );
  NANDN U17557 ( .A(n16681), .B(n16680), .Z(n16683) );
  XNOR U17558 ( .A(n16677), .B(n16676), .Z(n16678) );
  XNOR U17559 ( .A(n16679), .B(n16678), .Z(n16830) );
  XNOR U17560 ( .A(n16681), .B(n16680), .Z(n16829) );
  NAND U17561 ( .A(n16830), .B(n16829), .Z(n16682) );
  AND U17562 ( .A(n16683), .B(n16682), .Z(n17052) );
  IV U17563 ( .A(n16686), .Z(n17053) );
  NAND U17564 ( .A(a[41]), .B(b[17]), .Z(n17051) );
  NANDN U17565 ( .A(n16691), .B(n16692), .Z(n16694) );
  XOR U17566 ( .A(n16688), .B(n16687), .Z(n16689) );
  XNOR U17567 ( .A(n16690), .B(n16689), .Z(n16828) );
  NAND U17568 ( .A(n16828), .B(n16827), .Z(n16693) );
  NAND U17569 ( .A(n16694), .B(n16693), .Z(n17059) );
  NAND U17570 ( .A(a[43]), .B(b[17]), .Z(n17060) );
  AND U17571 ( .A(a[44]), .B(b[17]), .Z(n16695) );
  NANDN U17572 ( .A(n16696), .B(n16695), .Z(n16702) );
  XOR U17573 ( .A(n16696), .B(n16695), .Z(n16825) );
  XOR U17574 ( .A(n16698), .B(n16697), .Z(n16699) );
  XNOR U17575 ( .A(n16700), .B(n16699), .Z(n16826) );
  NANDN U17576 ( .A(n16825), .B(n16826), .Z(n16701) );
  NAND U17577 ( .A(n16702), .B(n16701), .Z(n17068) );
  NAND U17578 ( .A(a[45]), .B(b[17]), .Z(n17070) );
  AND U17579 ( .A(a[46]), .B(b[17]), .Z(n16707) );
  NANDN U17580 ( .A(n16708), .B(n16707), .Z(n16710) );
  XNOR U17581 ( .A(n16704), .B(n16703), .Z(n16705) );
  XNOR U17582 ( .A(n16706), .B(n16705), .Z(n16824) );
  XNOR U17583 ( .A(n16708), .B(n16707), .Z(n16823) );
  NAND U17584 ( .A(n16824), .B(n16823), .Z(n16709) );
  AND U17585 ( .A(n16710), .B(n16709), .Z(n16714) );
  NAND U17586 ( .A(n16714), .B(n16713), .Z(n16716) );
  XOR U17587 ( .A(n16714), .B(n16713), .Z(n17076) );
  NAND U17588 ( .A(a[47]), .B(b[17]), .Z(n17075) );
  NAND U17589 ( .A(n17076), .B(n17075), .Z(n16715) );
  AND U17590 ( .A(n16716), .B(n16715), .Z(n17084) );
  NANDN U17591 ( .A(n16719), .B(n16720), .Z(n16722) );
  XOR U17592 ( .A(n16718), .B(n16717), .Z(n16821) );
  XNOR U17593 ( .A(n16720), .B(n16719), .Z(n16822) );
  NANDN U17594 ( .A(n16821), .B(n16822), .Z(n16721) );
  AND U17595 ( .A(n16722), .B(n16721), .Z(n16726) );
  AND U17596 ( .A(a[50]), .B(b[17]), .Z(n16725) );
  NANDN U17597 ( .A(n16726), .B(n16725), .Z(n16728) );
  XOR U17598 ( .A(n16724), .B(n16723), .Z(n17091) );
  XNOR U17599 ( .A(n16726), .B(n16725), .Z(n17092) );
  NANDN U17600 ( .A(n17091), .B(n17092), .Z(n16727) );
  AND U17601 ( .A(n16728), .B(n16727), .Z(n16732) );
  AND U17602 ( .A(a[51]), .B(b[17]), .Z(n16731) );
  NANDN U17603 ( .A(n16732), .B(n16731), .Z(n16734) );
  XOR U17604 ( .A(n16730), .B(n16729), .Z(n16817) );
  XNOR U17605 ( .A(n16732), .B(n16731), .Z(n16818) );
  NANDN U17606 ( .A(n16817), .B(n16818), .Z(n16733) );
  AND U17607 ( .A(n16734), .B(n16733), .Z(n16738) );
  AND U17608 ( .A(a[52]), .B(b[17]), .Z(n16737) );
  NANDN U17609 ( .A(n16738), .B(n16737), .Z(n16740) );
  XOR U17610 ( .A(n16736), .B(n16735), .Z(n17099) );
  XNOR U17611 ( .A(n16738), .B(n16737), .Z(n17100) );
  NANDN U17612 ( .A(n17099), .B(n17100), .Z(n16739) );
  NAND U17613 ( .A(n16740), .B(n16739), .Z(n16813) );
  XOR U17614 ( .A(n16742), .B(n16741), .Z(n16816) );
  NANDN U17615 ( .A(n16745), .B(n16746), .Z(n16748) );
  XOR U17616 ( .A(n16744), .B(n16743), .Z(n17109) );
  XNOR U17617 ( .A(n16746), .B(n16745), .Z(n17110) );
  NANDN U17618 ( .A(n17109), .B(n17110), .Z(n16747) );
  AND U17619 ( .A(n16748), .B(n16747), .Z(n16749) );
  NANDN U17620 ( .A(n16750), .B(n16749), .Z(n16754) );
  XOR U17621 ( .A(n16750), .B(n16749), .Z(n16811) );
  XOR U17622 ( .A(n16752), .B(n16751), .Z(n16812) );
  NANDN U17623 ( .A(n16811), .B(n16812), .Z(n16753) );
  AND U17624 ( .A(n16754), .B(n16753), .Z(n16758) );
  NANDN U17625 ( .A(n16757), .B(n16758), .Z(n16760) );
  XOR U17626 ( .A(n16756), .B(n16755), .Z(n17117) );
  XNOR U17627 ( .A(n16758), .B(n16757), .Z(n17118) );
  NANDN U17628 ( .A(n17117), .B(n17118), .Z(n16759) );
  AND U17629 ( .A(n16760), .B(n16759), .Z(n16761) );
  NANDN U17630 ( .A(n16762), .B(n16761), .Z(n16766) );
  XOR U17631 ( .A(n16762), .B(n16761), .Z(n16809) );
  XOR U17632 ( .A(n16764), .B(n16763), .Z(n16810) );
  NANDN U17633 ( .A(n16809), .B(n16810), .Z(n16765) );
  AND U17634 ( .A(n16766), .B(n16765), .Z(n16770) );
  NANDN U17635 ( .A(n16769), .B(n16770), .Z(n16772) );
  XOR U17636 ( .A(n16768), .B(n16767), .Z(n17125) );
  XNOR U17637 ( .A(n16770), .B(n16769), .Z(n17126) );
  NANDN U17638 ( .A(n17125), .B(n17126), .Z(n16771) );
  AND U17639 ( .A(n16772), .B(n16771), .Z(n16773) );
  NANDN U17640 ( .A(n16774), .B(n16773), .Z(n16778) );
  XOR U17641 ( .A(n16774), .B(n16773), .Z(n16807) );
  XOR U17642 ( .A(n16776), .B(n16775), .Z(n16808) );
  NANDN U17643 ( .A(n16807), .B(n16808), .Z(n16777) );
  AND U17644 ( .A(n16778), .B(n16777), .Z(n16782) );
  NANDN U17645 ( .A(n16781), .B(n16782), .Z(n16784) );
  XOR U17646 ( .A(n16780), .B(n16779), .Z(n17133) );
  XNOR U17647 ( .A(n16782), .B(n16781), .Z(n17134) );
  NANDN U17648 ( .A(n17133), .B(n17134), .Z(n16783) );
  AND U17649 ( .A(n16784), .B(n16783), .Z(n16785) );
  NANDN U17650 ( .A(n16786), .B(n16785), .Z(n16790) );
  XOR U17651 ( .A(n16786), .B(n16785), .Z(n16805) );
  XOR U17652 ( .A(n16788), .B(n16787), .Z(n16806) );
  NANDN U17653 ( .A(n16805), .B(n16806), .Z(n16789) );
  AND U17654 ( .A(n16790), .B(n16789), .Z(n16794) );
  NANDN U17655 ( .A(n16793), .B(n16794), .Z(n16796) );
  XOR U17656 ( .A(n16792), .B(n16791), .Z(n17141) );
  XNOR U17657 ( .A(n16794), .B(n16793), .Z(n17142) );
  NANDN U17658 ( .A(n17141), .B(n17142), .Z(n16795) );
  AND U17659 ( .A(n16796), .B(n16795), .Z(n16797) );
  NANDN U17660 ( .A(n16798), .B(n16797), .Z(n16802) );
  XOR U17661 ( .A(n16798), .B(n16797), .Z(n17147) );
  XOR U17662 ( .A(n16800), .B(n16799), .Z(n17148) );
  OR U17663 ( .A(n17147), .B(n17148), .Z(n16801) );
  NAND U17664 ( .A(n16802), .B(n16801), .Z(n17149) );
  ANDN U17665 ( .B(n17150), .A(n17149), .Z(n22511) );
  XOR U17666 ( .A(n16804), .B(n16803), .Z(n22510) );
  NANDN U17667 ( .A(n22511), .B(n22510), .Z(n22513) );
  XOR U17668 ( .A(n16806), .B(n16805), .Z(n17140) );
  AND U17669 ( .A(a[62]), .B(b[16]), .Z(n17139) );
  XOR U17670 ( .A(n16808), .B(n16807), .Z(n17132) );
  AND U17671 ( .A(a[60]), .B(b[16]), .Z(n17131) );
  XOR U17672 ( .A(n16810), .B(n16809), .Z(n17124) );
  AND U17673 ( .A(a[58]), .B(b[16]), .Z(n17123) );
  XOR U17674 ( .A(n16812), .B(n16811), .Z(n17116) );
  AND U17675 ( .A(a[56]), .B(b[16]), .Z(n17115) );
  XOR U17676 ( .A(n16814), .B(n16813), .Z(n16815) );
  XOR U17677 ( .A(n16816), .B(n16815), .Z(n17106) );
  AND U17678 ( .A(a[54]), .B(b[16]), .Z(n17105) );
  NANDN U17679 ( .A(n17106), .B(n17105), .Z(n17108) );
  NAND U17680 ( .A(a[52]), .B(b[16]), .Z(n16819) );
  XNOR U17681 ( .A(n16818), .B(n16817), .Z(n16820) );
  NANDN U17682 ( .A(n16819), .B(n16820), .Z(n17098) );
  XOR U17683 ( .A(n16820), .B(n16819), .Z(n17435) );
  NAND U17684 ( .A(a[50]), .B(b[16]), .Z(n17087) );
  XNOR U17685 ( .A(n16822), .B(n16821), .Z(n17088) );
  NANDN U17686 ( .A(n17087), .B(n17088), .Z(n17090) );
  XNOR U17687 ( .A(n16824), .B(n16823), .Z(n17407) );
  NAND U17688 ( .A(a[46]), .B(b[16]), .Z(n17065) );
  AND U17689 ( .A(a[44]), .B(b[16]), .Z(n17061) );
  XNOR U17690 ( .A(n16828), .B(n16827), .Z(n17392) );
  XNOR U17691 ( .A(n16830), .B(n16829), .Z(n17386) );
  NAND U17692 ( .A(a[40]), .B(b[16]), .Z(n17043) );
  XNOR U17693 ( .A(n16832), .B(n16831), .Z(n17371) );
  XNOR U17694 ( .A(n16834), .B(n16833), .Z(n17363) );
  XOR U17695 ( .A(n16836), .B(n16835), .Z(n17012) );
  IV U17696 ( .A(n17012), .Z(n17348) );
  NAND U17697 ( .A(a[32]), .B(b[16]), .Z(n17340) );
  AND U17698 ( .A(a[30]), .B(b[16]), .Z(n16992) );
  IV U17699 ( .A(n16992), .Z(n17168) );
  XNOR U17700 ( .A(n16838), .B(n16837), .Z(n17317) );
  XNOR U17701 ( .A(n16840), .B(n16839), .Z(n17309) );
  XNOR U17702 ( .A(n16842), .B(n16841), .Z(n17301) );
  XNOR U17703 ( .A(n16844), .B(n16843), .Z(n17291) );
  NAND U17704 ( .A(a[20]), .B(b[16]), .Z(n16953) );
  XNOR U17705 ( .A(n16846), .B(n16845), .Z(n17284) );
  XNOR U17706 ( .A(n16848), .B(n16847), .Z(n17275) );
  AND U17707 ( .A(a[8]), .B(b[16]), .Z(n16890) );
  XOR U17708 ( .A(n16850), .B(n16849), .Z(n16872) );
  AND U17709 ( .A(b[16]), .B(a[0]), .Z(n17557) );
  AND U17710 ( .A(a[1]), .B(b[17]), .Z(n16854) );
  AND U17711 ( .A(n17557), .B(n16854), .Z(n16851) );
  NAND U17712 ( .A(a[2]), .B(n16851), .Z(n16858) );
  NAND U17713 ( .A(b[17]), .B(a[1]), .Z(n16852) );
  XOR U17714 ( .A(n16853), .B(n16852), .Z(n17193) );
  NAND U17715 ( .A(n16854), .B(a[0]), .Z(n16855) );
  XNOR U17716 ( .A(a[2]), .B(n16855), .Z(n16856) );
  AND U17717 ( .A(b[16]), .B(n16856), .Z(n17194) );
  NANDN U17718 ( .A(n17193), .B(n17194), .Z(n16857) );
  AND U17719 ( .A(n16858), .B(n16857), .Z(n16862) );
  XNOR U17720 ( .A(n16860), .B(n16859), .Z(n16861) );
  NANDN U17721 ( .A(n16862), .B(n16861), .Z(n16864) );
  XNOR U17722 ( .A(n16862), .B(n16861), .Z(n17200) );
  AND U17723 ( .A(a[3]), .B(b[16]), .Z(n17199) );
  NAND U17724 ( .A(n17200), .B(n17199), .Z(n16863) );
  AND U17725 ( .A(n16864), .B(n16863), .Z(n16866) );
  AND U17726 ( .A(a[4]), .B(b[16]), .Z(n16865) );
  NANDN U17727 ( .A(n16866), .B(n16865), .Z(n16870) );
  XNOR U17728 ( .A(n16866), .B(n16865), .Z(n17206) );
  XNOR U17729 ( .A(n16868), .B(n16867), .Z(n17205) );
  NAND U17730 ( .A(n17206), .B(n17205), .Z(n16869) );
  NAND U17731 ( .A(n16870), .B(n16869), .Z(n16871) );
  NAND U17732 ( .A(n16872), .B(n16871), .Z(n16874) );
  NAND U17733 ( .A(a[5]), .B(b[16]), .Z(n17211) );
  XOR U17734 ( .A(n16872), .B(n16871), .Z(n17212) );
  NANDN U17735 ( .A(n17211), .B(n17212), .Z(n16873) );
  AND U17736 ( .A(n16874), .B(n16873), .Z(n16878) );
  XNOR U17737 ( .A(n16876), .B(n16875), .Z(n16877) );
  NANDN U17738 ( .A(n16878), .B(n16877), .Z(n16880) );
  NAND U17739 ( .A(a[6]), .B(b[16]), .Z(n17217) );
  XNOR U17740 ( .A(n16878), .B(n16877), .Z(n17218) );
  NANDN U17741 ( .A(n17217), .B(n17218), .Z(n16879) );
  AND U17742 ( .A(n16880), .B(n16879), .Z(n16884) );
  XNOR U17743 ( .A(n16882), .B(n16881), .Z(n16883) );
  NANDN U17744 ( .A(n16884), .B(n16883), .Z(n16886) );
  NAND U17745 ( .A(a[7]), .B(b[16]), .Z(n17225) );
  XNOR U17746 ( .A(n16884), .B(n16883), .Z(n17226) );
  NANDN U17747 ( .A(n17225), .B(n17226), .Z(n16885) );
  AND U17748 ( .A(n16886), .B(n16885), .Z(n16889) );
  NANDN U17749 ( .A(n16890), .B(n16889), .Z(n16892) );
  XOR U17750 ( .A(n16888), .B(n16887), .Z(n17184) );
  XNOR U17751 ( .A(n16890), .B(n16889), .Z(n17183) );
  NANDN U17752 ( .A(n17184), .B(n17183), .Z(n16891) );
  AND U17753 ( .A(n16892), .B(n16891), .Z(n16896) );
  XOR U17754 ( .A(n16894), .B(n16893), .Z(n16895) );
  NAND U17755 ( .A(n16896), .B(n16895), .Z(n16898) );
  NAND U17756 ( .A(a[9]), .B(b[16]), .Z(n17233) );
  XOR U17757 ( .A(n16896), .B(n16895), .Z(n17234) );
  NANDN U17758 ( .A(n17233), .B(n17234), .Z(n16897) );
  AND U17759 ( .A(n16898), .B(n16897), .Z(n16900) );
  AND U17760 ( .A(a[10]), .B(b[16]), .Z(n16899) );
  NANDN U17761 ( .A(n16900), .B(n16899), .Z(n16904) );
  XNOR U17762 ( .A(n16900), .B(n16899), .Z(n17240) );
  XNOR U17763 ( .A(n16902), .B(n16901), .Z(n17239) );
  NAND U17764 ( .A(n17240), .B(n17239), .Z(n16903) );
  AND U17765 ( .A(n16904), .B(n16903), .Z(n16908) );
  XOR U17766 ( .A(n16906), .B(n16905), .Z(n16907) );
  NANDN U17767 ( .A(n16908), .B(n16907), .Z(n16910) );
  NAND U17768 ( .A(a[11]), .B(b[16]), .Z(n17245) );
  XNOR U17769 ( .A(n16908), .B(n16907), .Z(n17246) );
  NANDN U17770 ( .A(n17245), .B(n17246), .Z(n16909) );
  AND U17771 ( .A(n16910), .B(n16909), .Z(n16912) );
  AND U17772 ( .A(a[12]), .B(b[16]), .Z(n16911) );
  NANDN U17773 ( .A(n16912), .B(n16911), .Z(n16916) );
  XNOR U17774 ( .A(n16912), .B(n16911), .Z(n17252) );
  XNOR U17775 ( .A(n16914), .B(n16913), .Z(n17251) );
  NAND U17776 ( .A(n17252), .B(n17251), .Z(n16915) );
  AND U17777 ( .A(n16916), .B(n16915), .Z(n16920) );
  XOR U17778 ( .A(n16918), .B(n16917), .Z(n16919) );
  NANDN U17779 ( .A(n16920), .B(n16919), .Z(n16922) );
  NAND U17780 ( .A(a[13]), .B(b[16]), .Z(n17257) );
  XNOR U17781 ( .A(n16920), .B(n16919), .Z(n17258) );
  NANDN U17782 ( .A(n17257), .B(n17258), .Z(n16921) );
  AND U17783 ( .A(n16922), .B(n16921), .Z(n16924) );
  AND U17784 ( .A(a[14]), .B(b[16]), .Z(n16923) );
  NANDN U17785 ( .A(n16924), .B(n16923), .Z(n16928) );
  XNOR U17786 ( .A(n16924), .B(n16923), .Z(n17264) );
  XNOR U17787 ( .A(n16926), .B(n16925), .Z(n17263) );
  NAND U17788 ( .A(n17264), .B(n17263), .Z(n16927) );
  AND U17789 ( .A(n16928), .B(n16927), .Z(n16932) );
  XOR U17790 ( .A(n16930), .B(n16929), .Z(n16931) );
  NANDN U17791 ( .A(n16932), .B(n16931), .Z(n16934) );
  NAND U17792 ( .A(a[15]), .B(b[16]), .Z(n17269) );
  XNOR U17793 ( .A(n16932), .B(n16931), .Z(n17270) );
  NANDN U17794 ( .A(n17269), .B(n17270), .Z(n16933) );
  AND U17795 ( .A(n16934), .B(n16933), .Z(n16936) );
  AND U17796 ( .A(a[16]), .B(b[16]), .Z(n16935) );
  NANDN U17797 ( .A(n16936), .B(n16935), .Z(n16940) );
  XNOR U17798 ( .A(n16936), .B(n16935), .Z(n17182) );
  XNOR U17799 ( .A(n16938), .B(n16937), .Z(n17181) );
  NAND U17800 ( .A(n17182), .B(n17181), .Z(n16939) );
  NAND U17801 ( .A(n16940), .B(n16939), .Z(n17276) );
  NAND U17802 ( .A(a[17]), .B(b[16]), .Z(n17278) );
  AND U17803 ( .A(a[18]), .B(b[16]), .Z(n16945) );
  NANDN U17804 ( .A(n16946), .B(n16945), .Z(n16948) );
  XNOR U17805 ( .A(n16942), .B(n16941), .Z(n16943) );
  XNOR U17806 ( .A(n16944), .B(n16943), .Z(n17180) );
  XNOR U17807 ( .A(n16946), .B(n16945), .Z(n17179) );
  NAND U17808 ( .A(n17180), .B(n17179), .Z(n16947) );
  AND U17809 ( .A(n16948), .B(n16947), .Z(n17283) );
  NAND U17810 ( .A(a[19]), .B(b[16]), .Z(n17286) );
  NANDN U17811 ( .A(n16953), .B(n16954), .Z(n16956) );
  XNOR U17812 ( .A(n16950), .B(n16949), .Z(n16951) );
  XNOR U17813 ( .A(n16952), .B(n16951), .Z(n17178) );
  XNOR U17814 ( .A(n16954), .B(n16953), .Z(n17177) );
  NAND U17815 ( .A(n17178), .B(n17177), .Z(n16955) );
  NAND U17816 ( .A(n16956), .B(n16955), .Z(n17292) );
  NAND U17817 ( .A(a[21]), .B(b[16]), .Z(n17294) );
  AND U17818 ( .A(a[22]), .B(b[16]), .Z(n16957) );
  NANDN U17819 ( .A(n16958), .B(n16957), .Z(n16964) );
  XOR U17820 ( .A(n16958), .B(n16957), .Z(n17299) );
  XNOR U17821 ( .A(n16960), .B(n16959), .Z(n16961) );
  XNOR U17822 ( .A(n16962), .B(n16961), .Z(n17300) );
  NANDN U17823 ( .A(n17299), .B(n17300), .Z(n16963) );
  NAND U17824 ( .A(n16964), .B(n16963), .Z(n17302) );
  NAND U17825 ( .A(a[23]), .B(b[16]), .Z(n17304) );
  AND U17826 ( .A(a[24]), .B(b[16]), .Z(n16969) );
  NANDN U17827 ( .A(n16970), .B(n16969), .Z(n16972) );
  XNOR U17828 ( .A(n16966), .B(n16965), .Z(n16967) );
  XNOR U17829 ( .A(n16968), .B(n16967), .Z(n17176) );
  XNOR U17830 ( .A(n16970), .B(n16969), .Z(n17175) );
  NAND U17831 ( .A(n17176), .B(n17175), .Z(n16971) );
  NAND U17832 ( .A(n16972), .B(n16971), .Z(n17310) );
  NAND U17833 ( .A(a[25]), .B(b[16]), .Z(n17312) );
  AND U17834 ( .A(a[26]), .B(b[16]), .Z(n16973) );
  NANDN U17835 ( .A(n16974), .B(n16973), .Z(n16980) );
  XOR U17836 ( .A(n16974), .B(n16973), .Z(n17173) );
  XOR U17837 ( .A(n16976), .B(n16975), .Z(n16977) );
  XNOR U17838 ( .A(n16978), .B(n16977), .Z(n17174) );
  NANDN U17839 ( .A(n17173), .B(n17174), .Z(n16979) );
  NAND U17840 ( .A(n16980), .B(n16979), .Z(n17318) );
  NAND U17841 ( .A(a[27]), .B(b[16]), .Z(n17320) );
  AND U17842 ( .A(a[28]), .B(b[16]), .Z(n16985) );
  NANDN U17843 ( .A(n16984), .B(n16985), .Z(n16987) );
  XNOR U17844 ( .A(n16985), .B(n16984), .Z(n17171) );
  NAND U17845 ( .A(n17172), .B(n17171), .Z(n16986) );
  AND U17846 ( .A(n16987), .B(n16986), .Z(n17326) );
  IV U17847 ( .A(n16991), .Z(n17327) );
  NAND U17848 ( .A(a[29]), .B(b[16]), .Z(n17325) );
  NANDN U17849 ( .A(n17168), .B(n17167), .Z(n16999) );
  NOR U17850 ( .A(n16992), .B(n17167), .Z(n16997) );
  XOR U17851 ( .A(n16994), .B(n16993), .Z(n16995) );
  XNOR U17852 ( .A(n16996), .B(n16995), .Z(n17170) );
  OR U17853 ( .A(n16997), .B(n17170), .Z(n16998) );
  AND U17854 ( .A(n16999), .B(n16998), .Z(n17335) );
  XOR U17855 ( .A(n17001), .B(n17000), .Z(n17002) );
  XOR U17856 ( .A(n17003), .B(n17002), .Z(n17004) );
  IV U17857 ( .A(n17004), .Z(n17334) );
  OR U17858 ( .A(n17335), .B(n17334), .Z(n17007) );
  ANDN U17859 ( .B(n17335), .A(n17004), .Z(n17005) );
  AND U17860 ( .A(a[31]), .B(b[16]), .Z(n17333) );
  NANDN U17861 ( .A(n17005), .B(n17333), .Z(n17006) );
  AND U17862 ( .A(n17007), .B(n17006), .Z(n17339) );
  XOR U17863 ( .A(n17009), .B(n17008), .Z(n17010) );
  XNOR U17864 ( .A(n17011), .B(n17010), .Z(n17342) );
  NANDN U17865 ( .A(n17348), .B(n17349), .Z(n17015) );
  NOR U17866 ( .A(n17012), .B(n17349), .Z(n17013) );
  NAND U17867 ( .A(a[33]), .B(b[16]), .Z(n17351) );
  OR U17868 ( .A(n17013), .B(n17351), .Z(n17014) );
  AND U17869 ( .A(n17015), .B(n17014), .Z(n17021) );
  AND U17870 ( .A(a[34]), .B(b[16]), .Z(n17020) );
  NANDN U17871 ( .A(n17021), .B(n17020), .Z(n17023) );
  XNOR U17872 ( .A(n17017), .B(n17016), .Z(n17018) );
  XNOR U17873 ( .A(n17019), .B(n17018), .Z(n17356) );
  XNOR U17874 ( .A(n17021), .B(n17020), .Z(n17355) );
  NAND U17875 ( .A(n17356), .B(n17355), .Z(n17022) );
  NAND U17876 ( .A(n17023), .B(n17022), .Z(n17364) );
  NAND U17877 ( .A(a[35]), .B(b[16]), .Z(n17366) );
  AND U17878 ( .A(a[36]), .B(b[16]), .Z(n17029) );
  NANDN U17879 ( .A(n17028), .B(n17029), .Z(n17031) );
  XNOR U17880 ( .A(n17025), .B(n17024), .Z(n17026) );
  XNOR U17881 ( .A(n17027), .B(n17026), .Z(n17166) );
  XNOR U17882 ( .A(n17029), .B(n17028), .Z(n17165) );
  NAND U17883 ( .A(n17166), .B(n17165), .Z(n17030) );
  NAND U17884 ( .A(n17031), .B(n17030), .Z(n17372) );
  NAND U17885 ( .A(a[37]), .B(b[16]), .Z(n17374) );
  AND U17886 ( .A(a[38]), .B(b[16]), .Z(n17033) );
  NANDN U17887 ( .A(n17032), .B(n17033), .Z(n17039) );
  XNOR U17888 ( .A(n17033), .B(n17032), .Z(n17164) );
  XNOR U17889 ( .A(n17035), .B(n17034), .Z(n17036) );
  XNOR U17890 ( .A(n17037), .B(n17036), .Z(n17163) );
  NAND U17891 ( .A(n17164), .B(n17163), .Z(n17038) );
  AND U17892 ( .A(n17039), .B(n17038), .Z(n17378) );
  IV U17893 ( .A(n17042), .Z(n17379) );
  NAND U17894 ( .A(a[39]), .B(b[16]), .Z(n17377) );
  NANDN U17895 ( .A(n17043), .B(n17044), .Z(n17050) );
  XNOR U17896 ( .A(n17046), .B(n17045), .Z(n17047) );
  XNOR U17897 ( .A(n17048), .B(n17047), .Z(n17161) );
  NAND U17898 ( .A(n17162), .B(n17161), .Z(n17049) );
  NAND U17899 ( .A(n17050), .B(n17049), .Z(n17387) );
  NAND U17900 ( .A(a[41]), .B(b[16]), .Z(n17389) );
  AND U17901 ( .A(a[42]), .B(b[16]), .Z(n17055) );
  NANDN U17902 ( .A(n17054), .B(n17055), .Z(n17057) );
  XNOR U17903 ( .A(n17055), .B(n17054), .Z(n17159) );
  NAND U17904 ( .A(n17160), .B(n17159), .Z(n17056) );
  NAND U17905 ( .A(n17057), .B(n17056), .Z(n17393) );
  NAND U17906 ( .A(a[43]), .B(b[16]), .Z(n17395) );
  NANDN U17907 ( .A(n17061), .B(n17062), .Z(n17064) );
  NANDN U17908 ( .A(n17157), .B(n17158), .Z(n17063) );
  NAND U17909 ( .A(n17064), .B(n17063), .Z(n17401) );
  AND U17910 ( .A(a[45]), .B(b[16]), .Z(n17402) );
  NANDN U17911 ( .A(n17065), .B(n17066), .Z(n17072) );
  XNOR U17912 ( .A(n17068), .B(n17067), .Z(n17069) );
  XNOR U17913 ( .A(n17070), .B(n17069), .Z(n17155) );
  NAND U17914 ( .A(n17156), .B(n17155), .Z(n17071) );
  NAND U17915 ( .A(n17072), .B(n17071), .Z(n17408) );
  NAND U17916 ( .A(a[47]), .B(b[16]), .Z(n17410) );
  AND U17917 ( .A(a[48]), .B(b[16]), .Z(n17073) );
  NANDN U17918 ( .A(n17074), .B(n17073), .Z(n17078) );
  XOR U17919 ( .A(n17074), .B(n17073), .Z(n17415) );
  XNOR U17920 ( .A(n17076), .B(n17075), .Z(n17416) );
  NANDN U17921 ( .A(n17415), .B(n17416), .Z(n17077) );
  AND U17922 ( .A(n17078), .B(n17077), .Z(n17080) );
  AND U17923 ( .A(a[49]), .B(b[16]), .Z(n17079) );
  NANDN U17924 ( .A(n17080), .B(n17079), .Z(n17086) );
  XOR U17925 ( .A(n17080), .B(n17079), .Z(n17153) );
  XOR U17926 ( .A(n17082), .B(n17081), .Z(n17083) );
  XNOR U17927 ( .A(n17084), .B(n17083), .Z(n17154) );
  NANDN U17928 ( .A(n17153), .B(n17154), .Z(n17085) );
  AND U17929 ( .A(n17086), .B(n17085), .Z(n17422) );
  XNOR U17930 ( .A(n17088), .B(n17087), .Z(n17421) );
  NANDN U17931 ( .A(n17422), .B(n17421), .Z(n17089) );
  AND U17932 ( .A(n17090), .B(n17089), .Z(n17094) );
  XNOR U17933 ( .A(n17092), .B(n17091), .Z(n17093) );
  NANDN U17934 ( .A(n17094), .B(n17093), .Z(n17096) );
  NAND U17935 ( .A(a[51]), .B(b[16]), .Z(n17427) );
  XNOR U17936 ( .A(n17094), .B(n17093), .Z(n17428) );
  NANDN U17937 ( .A(n17427), .B(n17428), .Z(n17095) );
  AND U17938 ( .A(n17096), .B(n17095), .Z(n17436) );
  OR U17939 ( .A(n17435), .B(n17436), .Z(n17097) );
  AND U17940 ( .A(n17098), .B(n17097), .Z(n17102) );
  XNOR U17941 ( .A(n17100), .B(n17099), .Z(n17101) );
  NANDN U17942 ( .A(n17102), .B(n17101), .Z(n17104) );
  NAND U17943 ( .A(a[53]), .B(b[16]), .Z(n17439) );
  XNOR U17944 ( .A(n17102), .B(n17101), .Z(n17440) );
  NANDN U17945 ( .A(n17439), .B(n17440), .Z(n17103) );
  AND U17946 ( .A(n17104), .B(n17103), .Z(n17446) );
  XNOR U17947 ( .A(n17106), .B(n17105), .Z(n17445) );
  NANDN U17948 ( .A(n17446), .B(n17445), .Z(n17107) );
  AND U17949 ( .A(n17108), .B(n17107), .Z(n17112) );
  XNOR U17950 ( .A(n17110), .B(n17109), .Z(n17111) );
  NANDN U17951 ( .A(n17112), .B(n17111), .Z(n17114) );
  NAND U17952 ( .A(a[55]), .B(b[16]), .Z(n17451) );
  XNOR U17953 ( .A(n17112), .B(n17111), .Z(n17452) );
  NANDN U17954 ( .A(n17451), .B(n17452), .Z(n17113) );
  AND U17955 ( .A(n17114), .B(n17113), .Z(n17458) );
  XOR U17956 ( .A(n17116), .B(n17115), .Z(n17457) );
  XNOR U17957 ( .A(n17118), .B(n17117), .Z(n17119) );
  NANDN U17958 ( .A(n17120), .B(n17119), .Z(n17122) );
  NAND U17959 ( .A(a[57]), .B(b[16]), .Z(n17459) );
  XNOR U17960 ( .A(n17120), .B(n17119), .Z(n17460) );
  NANDN U17961 ( .A(n17459), .B(n17460), .Z(n17121) );
  AND U17962 ( .A(n17122), .B(n17121), .Z(n17468) );
  XOR U17963 ( .A(n17124), .B(n17123), .Z(n17467) );
  XNOR U17964 ( .A(n17126), .B(n17125), .Z(n17127) );
  NANDN U17965 ( .A(n17128), .B(n17127), .Z(n17130) );
  NAND U17966 ( .A(a[59]), .B(b[16]), .Z(n17471) );
  XNOR U17967 ( .A(n17128), .B(n17127), .Z(n17472) );
  NANDN U17968 ( .A(n17471), .B(n17472), .Z(n17129) );
  AND U17969 ( .A(n17130), .B(n17129), .Z(n17480) );
  XOR U17970 ( .A(n17132), .B(n17131), .Z(n17479) );
  XNOR U17971 ( .A(n17134), .B(n17133), .Z(n17135) );
  NANDN U17972 ( .A(n17136), .B(n17135), .Z(n17138) );
  NAND U17973 ( .A(a[61]), .B(b[16]), .Z(n17483) );
  XNOR U17974 ( .A(n17136), .B(n17135), .Z(n17484) );
  NANDN U17975 ( .A(n17483), .B(n17484), .Z(n17137) );
  AND U17976 ( .A(n17138), .B(n17137), .Z(n17492) );
  XOR U17977 ( .A(n17140), .B(n17139), .Z(n17491) );
  XNOR U17978 ( .A(n17142), .B(n17141), .Z(n17143) );
  NANDN U17979 ( .A(n17144), .B(n17143), .Z(n17146) );
  NAND U17980 ( .A(a[63]), .B(b[16]), .Z(n17495) );
  XNOR U17981 ( .A(n17144), .B(n17143), .Z(n17496) );
  NANDN U17982 ( .A(n17495), .B(n17496), .Z(n17145) );
  NAND U17983 ( .A(n17146), .B(n17145), .Z(n17497) );
  XOR U17984 ( .A(n17148), .B(n17147), .Z(n17498) );
  ANDN U17985 ( .B(n17497), .A(n17498), .Z(n17151) );
  XNOR U17986 ( .A(n17150), .B(n17149), .Z(n17152) );
  XOR U17987 ( .A(n17152), .B(n17151), .Z(n24728) );
  AND U17988 ( .A(a[63]), .B(b[15]), .Z(n17490) );
  NAND U17989 ( .A(a[62]), .B(b[15]), .Z(n17485) );
  AND U17990 ( .A(a[61]), .B(b[15]), .Z(n17478) );
  NAND U17991 ( .A(a[60]), .B(b[15]), .Z(n17473) );
  AND U17992 ( .A(a[59]), .B(b[15]), .Z(n17466) );
  NAND U17993 ( .A(a[58]), .B(b[15]), .Z(n17461) );
  NAND U17994 ( .A(a[54]), .B(b[15]), .Z(n17441) );
  AND U17995 ( .A(a[53]), .B(b[15]), .Z(n17434) );
  NAND U17996 ( .A(a[51]), .B(b[15]), .Z(n17423) );
  AND U17997 ( .A(a[50]), .B(b[15]), .Z(n17779) );
  XOR U17998 ( .A(n17154), .B(n17153), .Z(n17778) );
  XNOR U17999 ( .A(n17156), .B(n17155), .Z(n17764) );
  XNOR U18000 ( .A(n17160), .B(n17159), .Z(n17751) );
  XNOR U18001 ( .A(n17162), .B(n17161), .Z(n17745) );
  XNOR U18002 ( .A(n17164), .B(n17163), .Z(n17736) );
  XNOR U18003 ( .A(n17166), .B(n17165), .Z(n17730) );
  XOR U18004 ( .A(n17168), .B(n17167), .Z(n17169) );
  XNOR U18005 ( .A(n17170), .B(n17169), .Z(n17701) );
  XNOR U18006 ( .A(n17172), .B(n17171), .Z(n17693) );
  NAND U18007 ( .A(a[28]), .B(b[15]), .Z(n17321) );
  XNOR U18008 ( .A(n17174), .B(n17173), .Z(n17686) );
  XNOR U18009 ( .A(n17176), .B(n17175), .Z(n17679) );
  XNOR U18010 ( .A(n17178), .B(n17177), .Z(n17661) );
  XNOR U18011 ( .A(n17180), .B(n17179), .Z(n17655) );
  XNOR U18012 ( .A(n17182), .B(n17181), .Z(n17645) );
  XOR U18013 ( .A(n17184), .B(n17183), .Z(n17230) );
  AND U18014 ( .A(a[4]), .B(b[15]), .Z(n17202) );
  AND U18015 ( .A(b[15]), .B(a[0]), .Z(n17880) );
  AND U18016 ( .A(a[1]), .B(b[16]), .Z(n17188) );
  AND U18017 ( .A(n17880), .B(n17188), .Z(n17185) );
  NAND U18018 ( .A(a[2]), .B(n17185), .Z(n17192) );
  NAND U18019 ( .A(b[16]), .B(a[1]), .Z(n17186) );
  XOR U18020 ( .A(n17187), .B(n17186), .Z(n17563) );
  NAND U18021 ( .A(n17188), .B(a[0]), .Z(n17189) );
  XNOR U18022 ( .A(a[2]), .B(n17189), .Z(n17190) );
  AND U18023 ( .A(b[15]), .B(n17190), .Z(n17564) );
  NANDN U18024 ( .A(n17563), .B(n17564), .Z(n17191) );
  AND U18025 ( .A(n17192), .B(n17191), .Z(n17196) );
  XNOR U18026 ( .A(n17194), .B(n17193), .Z(n17195) );
  NANDN U18027 ( .A(n17196), .B(n17195), .Z(n17198) );
  NAND U18028 ( .A(a[3]), .B(b[15]), .Z(n17571) );
  XNOR U18029 ( .A(n17196), .B(n17195), .Z(n17572) );
  NANDN U18030 ( .A(n17571), .B(n17572), .Z(n17197) );
  AND U18031 ( .A(n17198), .B(n17197), .Z(n17201) );
  NANDN U18032 ( .A(n17202), .B(n17201), .Z(n17204) );
  XOR U18033 ( .A(n17200), .B(n17199), .Z(n17554) );
  XNOR U18034 ( .A(n17202), .B(n17201), .Z(n17553) );
  NANDN U18035 ( .A(n17554), .B(n17553), .Z(n17203) );
  AND U18036 ( .A(n17204), .B(n17203), .Z(n17208) );
  XOR U18037 ( .A(n17206), .B(n17205), .Z(n17207) );
  NAND U18038 ( .A(n17208), .B(n17207), .Z(n17210) );
  NAND U18039 ( .A(a[5]), .B(b[15]), .Z(n17579) );
  XOR U18040 ( .A(n17208), .B(n17207), .Z(n17580) );
  NANDN U18041 ( .A(n17579), .B(n17580), .Z(n17209) );
  AND U18042 ( .A(n17210), .B(n17209), .Z(n17214) );
  XNOR U18043 ( .A(n17212), .B(n17211), .Z(n17213) );
  NANDN U18044 ( .A(n17214), .B(n17213), .Z(n17216) );
  NAND U18045 ( .A(a[6]), .B(b[15]), .Z(n17585) );
  XNOR U18046 ( .A(n17214), .B(n17213), .Z(n17586) );
  NANDN U18047 ( .A(n17585), .B(n17586), .Z(n17215) );
  AND U18048 ( .A(n17216), .B(n17215), .Z(n17220) );
  XNOR U18049 ( .A(n17218), .B(n17217), .Z(n17219) );
  NANDN U18050 ( .A(n17220), .B(n17219), .Z(n17222) );
  XNOR U18051 ( .A(n17220), .B(n17219), .Z(n17592) );
  AND U18052 ( .A(a[7]), .B(b[15]), .Z(n17591) );
  NAND U18053 ( .A(n17592), .B(n17591), .Z(n17221) );
  AND U18054 ( .A(n17222), .B(n17221), .Z(n17224) );
  AND U18055 ( .A(a[8]), .B(b[15]), .Z(n17223) );
  NANDN U18056 ( .A(n17224), .B(n17223), .Z(n17228) );
  XNOR U18057 ( .A(n17224), .B(n17223), .Z(n17598) );
  XNOR U18058 ( .A(n17226), .B(n17225), .Z(n17597) );
  NAND U18059 ( .A(n17598), .B(n17597), .Z(n17227) );
  NAND U18060 ( .A(n17228), .B(n17227), .Z(n17229) );
  NAND U18061 ( .A(n17230), .B(n17229), .Z(n17232) );
  NAND U18062 ( .A(a[9]), .B(b[15]), .Z(n17605) );
  XOR U18063 ( .A(n17230), .B(n17229), .Z(n17606) );
  NANDN U18064 ( .A(n17605), .B(n17606), .Z(n17231) );
  AND U18065 ( .A(n17232), .B(n17231), .Z(n17236) );
  AND U18066 ( .A(a[10]), .B(b[15]), .Z(n17235) );
  NANDN U18067 ( .A(n17236), .B(n17235), .Z(n17238) );
  XNOR U18068 ( .A(n17234), .B(n17233), .Z(n17610) );
  XNOR U18069 ( .A(n17236), .B(n17235), .Z(n17609) );
  NAND U18070 ( .A(n17610), .B(n17609), .Z(n17237) );
  AND U18071 ( .A(n17238), .B(n17237), .Z(n17242) );
  XOR U18072 ( .A(n17240), .B(n17239), .Z(n17241) );
  NANDN U18073 ( .A(n17242), .B(n17241), .Z(n17244) );
  NAND U18074 ( .A(a[11]), .B(b[15]), .Z(n17617) );
  XNOR U18075 ( .A(n17242), .B(n17241), .Z(n17618) );
  NANDN U18076 ( .A(n17617), .B(n17618), .Z(n17243) );
  AND U18077 ( .A(n17244), .B(n17243), .Z(n17248) );
  AND U18078 ( .A(a[12]), .B(b[15]), .Z(n17247) );
  NANDN U18079 ( .A(n17248), .B(n17247), .Z(n17250) );
  XNOR U18080 ( .A(n17246), .B(n17245), .Z(n17622) );
  XNOR U18081 ( .A(n17248), .B(n17247), .Z(n17621) );
  NAND U18082 ( .A(n17622), .B(n17621), .Z(n17249) );
  AND U18083 ( .A(n17250), .B(n17249), .Z(n17254) );
  XOR U18084 ( .A(n17252), .B(n17251), .Z(n17253) );
  NANDN U18085 ( .A(n17254), .B(n17253), .Z(n17256) );
  NAND U18086 ( .A(a[13]), .B(b[15]), .Z(n17629) );
  XNOR U18087 ( .A(n17254), .B(n17253), .Z(n17630) );
  NANDN U18088 ( .A(n17629), .B(n17630), .Z(n17255) );
  AND U18089 ( .A(n17256), .B(n17255), .Z(n17260) );
  AND U18090 ( .A(a[14]), .B(b[15]), .Z(n17259) );
  NANDN U18091 ( .A(n17260), .B(n17259), .Z(n17262) );
  XNOR U18092 ( .A(n17258), .B(n17257), .Z(n17634) );
  XNOR U18093 ( .A(n17260), .B(n17259), .Z(n17633) );
  NAND U18094 ( .A(n17634), .B(n17633), .Z(n17261) );
  AND U18095 ( .A(n17262), .B(n17261), .Z(n17266) );
  XOR U18096 ( .A(n17264), .B(n17263), .Z(n17265) );
  NANDN U18097 ( .A(n17266), .B(n17265), .Z(n17268) );
  NAND U18098 ( .A(a[15]), .B(b[15]), .Z(n17641) );
  XNOR U18099 ( .A(n17266), .B(n17265), .Z(n17642) );
  NANDN U18100 ( .A(n17641), .B(n17642), .Z(n17267) );
  AND U18101 ( .A(n17268), .B(n17267), .Z(n17272) );
  AND U18102 ( .A(a[16]), .B(b[15]), .Z(n17271) );
  NANDN U18103 ( .A(n17272), .B(n17271), .Z(n17274) );
  XNOR U18104 ( .A(n17270), .B(n17269), .Z(n17552) );
  XNOR U18105 ( .A(n17272), .B(n17271), .Z(n17551) );
  NAND U18106 ( .A(n17552), .B(n17551), .Z(n17273) );
  NAND U18107 ( .A(n17274), .B(n17273), .Z(n17646) );
  NAND U18108 ( .A(a[17]), .B(b[15]), .Z(n17648) );
  AND U18109 ( .A(a[18]), .B(b[15]), .Z(n17279) );
  NANDN U18110 ( .A(n17280), .B(n17279), .Z(n17282) );
  XNOR U18111 ( .A(n17276), .B(n17275), .Z(n17277) );
  XNOR U18112 ( .A(n17278), .B(n17277), .Z(n17550) );
  XNOR U18113 ( .A(n17280), .B(n17279), .Z(n17549) );
  NAND U18114 ( .A(n17550), .B(n17549), .Z(n17281) );
  NAND U18115 ( .A(n17282), .B(n17281), .Z(n17656) );
  NAND U18116 ( .A(a[19]), .B(b[15]), .Z(n17658) );
  AND U18117 ( .A(a[20]), .B(b[15]), .Z(n17287) );
  NANDN U18118 ( .A(n17288), .B(n17287), .Z(n17290) );
  XNOR U18119 ( .A(n17284), .B(n17283), .Z(n17285) );
  XNOR U18120 ( .A(n17286), .B(n17285), .Z(n17548) );
  XNOR U18121 ( .A(n17288), .B(n17287), .Z(n17547) );
  NAND U18122 ( .A(n17548), .B(n17547), .Z(n17289) );
  NAND U18123 ( .A(n17290), .B(n17289), .Z(n17662) );
  NAND U18124 ( .A(a[21]), .B(b[15]), .Z(n17664) );
  AND U18125 ( .A(a[22]), .B(b[15]), .Z(n17295) );
  NANDN U18126 ( .A(n17296), .B(n17295), .Z(n17298) );
  XNOR U18127 ( .A(n17292), .B(n17291), .Z(n17293) );
  XNOR U18128 ( .A(n17294), .B(n17293), .Z(n17546) );
  XNOR U18129 ( .A(n17296), .B(n17295), .Z(n17545) );
  NAND U18130 ( .A(n17546), .B(n17545), .Z(n17297) );
  AND U18131 ( .A(n17298), .B(n17297), .Z(n17670) );
  XNOR U18132 ( .A(n17300), .B(n17299), .Z(n17669) );
  NAND U18133 ( .A(a[23]), .B(b[15]), .Z(n17672) );
  AND U18134 ( .A(a[24]), .B(b[15]), .Z(n17305) );
  NANDN U18135 ( .A(n17306), .B(n17305), .Z(n17308) );
  XNOR U18136 ( .A(n17302), .B(n17301), .Z(n17303) );
  XNOR U18137 ( .A(n17304), .B(n17303), .Z(n17544) );
  XNOR U18138 ( .A(n17306), .B(n17305), .Z(n17543) );
  NAND U18139 ( .A(n17544), .B(n17543), .Z(n17307) );
  NAND U18140 ( .A(n17308), .B(n17307), .Z(n17680) );
  NAND U18141 ( .A(a[25]), .B(b[15]), .Z(n17682) );
  AND U18142 ( .A(a[26]), .B(b[15]), .Z(n17313) );
  NANDN U18143 ( .A(n17314), .B(n17313), .Z(n17316) );
  XNOR U18144 ( .A(n17310), .B(n17309), .Z(n17311) );
  XNOR U18145 ( .A(n17312), .B(n17311), .Z(n17542) );
  XNOR U18146 ( .A(n17314), .B(n17313), .Z(n17541) );
  NAND U18147 ( .A(n17542), .B(n17541), .Z(n17315) );
  AND U18148 ( .A(n17316), .B(n17315), .Z(n17685) );
  NAND U18149 ( .A(a[27]), .B(b[15]), .Z(n17688) );
  NANDN U18150 ( .A(n17321), .B(n17322), .Z(n17324) );
  XNOR U18151 ( .A(n17318), .B(n17317), .Z(n17319) );
  XNOR U18152 ( .A(n17320), .B(n17319), .Z(n17540) );
  XNOR U18153 ( .A(n17322), .B(n17321), .Z(n17539) );
  NAND U18154 ( .A(n17540), .B(n17539), .Z(n17323) );
  NAND U18155 ( .A(n17324), .B(n17323), .Z(n17694) );
  NAND U18156 ( .A(a[29]), .B(b[15]), .Z(n17696) );
  AND U18157 ( .A(a[30]), .B(b[15]), .Z(n17328) );
  NANDN U18158 ( .A(n17329), .B(n17328), .Z(n17331) );
  XNOR U18159 ( .A(n17329), .B(n17328), .Z(n17537) );
  NAND U18160 ( .A(n17538), .B(n17537), .Z(n17330) );
  NAND U18161 ( .A(n17331), .B(n17330), .Z(n17702) );
  NAND U18162 ( .A(a[31]), .B(b[15]), .Z(n17704) );
  AND U18163 ( .A(a[32]), .B(b[15]), .Z(n17332) );
  IV U18164 ( .A(n17332), .Z(n17533) );
  OR U18165 ( .A(n17534), .B(n17533), .Z(n17338) );
  ANDN U18166 ( .B(n17534), .A(n17332), .Z(n17336) );
  OR U18167 ( .A(n17336), .B(n17536), .Z(n17337) );
  AND U18168 ( .A(n17338), .B(n17337), .Z(n17712) );
  XOR U18169 ( .A(n17340), .B(n17339), .Z(n17341) );
  XOR U18170 ( .A(n17342), .B(n17341), .Z(n17343) );
  IV U18171 ( .A(n17343), .Z(n17711) );
  OR U18172 ( .A(n17712), .B(n17711), .Z(n17346) );
  ANDN U18173 ( .B(n17712), .A(n17343), .Z(n17344) );
  AND U18174 ( .A(a[33]), .B(b[15]), .Z(n17710) );
  NANDN U18175 ( .A(n17344), .B(n17710), .Z(n17345) );
  AND U18176 ( .A(n17346), .B(n17345), .Z(n17718) );
  AND U18177 ( .A(a[34]), .B(b[15]), .Z(n17347) );
  IV U18178 ( .A(n17347), .Z(n17717) );
  OR U18179 ( .A(n17718), .B(n17717), .Z(n17354) );
  ANDN U18180 ( .B(n17718), .A(n17347), .Z(n17352) );
  XOR U18181 ( .A(n17349), .B(n17348), .Z(n17350) );
  XOR U18182 ( .A(n17351), .B(n17350), .Z(n17716) );
  NANDN U18183 ( .A(n17352), .B(n17716), .Z(n17353) );
  AND U18184 ( .A(n17354), .B(n17353), .Z(n17720) );
  XOR U18185 ( .A(n17356), .B(n17355), .Z(n17357) );
  IV U18186 ( .A(n17357), .Z(n17719) );
  OR U18187 ( .A(n17720), .B(n17719), .Z(n17360) );
  ANDN U18188 ( .B(n17720), .A(n17357), .Z(n17358) );
  NAND U18189 ( .A(a[35]), .B(b[15]), .Z(n17722) );
  OR U18190 ( .A(n17358), .B(n17722), .Z(n17359) );
  AND U18191 ( .A(n17360), .B(n17359), .Z(n17362) );
  AND U18192 ( .A(a[36]), .B(b[15]), .Z(n17361) );
  NANDN U18193 ( .A(n17362), .B(n17361), .Z(n17368) );
  XNOR U18194 ( .A(n17362), .B(n17361), .Z(n17532) );
  XNOR U18195 ( .A(n17364), .B(n17363), .Z(n17365) );
  XNOR U18196 ( .A(n17366), .B(n17365), .Z(n17531) );
  NAND U18197 ( .A(n17532), .B(n17531), .Z(n17367) );
  NAND U18198 ( .A(n17368), .B(n17367), .Z(n17731) );
  AND U18199 ( .A(a[37]), .B(b[15]), .Z(n17729) );
  AND U18200 ( .A(a[38]), .B(b[15]), .Z(n17369) );
  NANDN U18201 ( .A(n17370), .B(n17369), .Z(n17376) );
  XOR U18202 ( .A(n17370), .B(n17369), .Z(n17529) );
  XNOR U18203 ( .A(n17372), .B(n17371), .Z(n17373) );
  XNOR U18204 ( .A(n17374), .B(n17373), .Z(n17530) );
  NANDN U18205 ( .A(n17529), .B(n17530), .Z(n17375) );
  NAND U18206 ( .A(n17376), .B(n17375), .Z(n17737) );
  NAND U18207 ( .A(a[39]), .B(b[15]), .Z(n17739) );
  AND U18208 ( .A(a[40]), .B(b[15]), .Z(n17380) );
  NANDN U18209 ( .A(n17381), .B(n17380), .Z(n17383) );
  XNOR U18210 ( .A(n17381), .B(n17380), .Z(n17527) );
  NAND U18211 ( .A(n17528), .B(n17527), .Z(n17382) );
  NAND U18212 ( .A(n17383), .B(n17382), .Z(n17746) );
  AND U18213 ( .A(a[41]), .B(b[15]), .Z(n17744) );
  AND U18214 ( .A(a[42]), .B(b[15]), .Z(n17384) );
  NANDN U18215 ( .A(n17385), .B(n17384), .Z(n17391) );
  XNOR U18216 ( .A(n17385), .B(n17384), .Z(n17526) );
  XNOR U18217 ( .A(n17387), .B(n17386), .Z(n17388) );
  XNOR U18218 ( .A(n17389), .B(n17388), .Z(n17525) );
  NAND U18219 ( .A(n17526), .B(n17525), .Z(n17390) );
  NAND U18220 ( .A(n17391), .B(n17390), .Z(n17752) );
  NAND U18221 ( .A(a[43]), .B(b[15]), .Z(n17754) );
  AND U18222 ( .A(a[44]), .B(b[15]), .Z(n17396) );
  NANDN U18223 ( .A(n17397), .B(n17396), .Z(n17399) );
  XNOR U18224 ( .A(n17393), .B(n17392), .Z(n17394) );
  XNOR U18225 ( .A(n17395), .B(n17394), .Z(n17524) );
  XNOR U18226 ( .A(n17397), .B(n17396), .Z(n17523) );
  NAND U18227 ( .A(n17524), .B(n17523), .Z(n17398) );
  NAND U18228 ( .A(n17399), .B(n17398), .Z(n17759) );
  AND U18229 ( .A(a[45]), .B(b[15]), .Z(n17757) );
  AND U18230 ( .A(a[46]), .B(b[15]), .Z(n17403) );
  NANDN U18231 ( .A(n17404), .B(n17403), .Z(n17406) );
  XNOR U18232 ( .A(n17404), .B(n17403), .Z(n17521) );
  NAND U18233 ( .A(n17522), .B(n17521), .Z(n17405) );
  NAND U18234 ( .A(n17406), .B(n17405), .Z(n17765) );
  NAND U18235 ( .A(a[47]), .B(b[15]), .Z(n17767) );
  AND U18236 ( .A(a[48]), .B(b[15]), .Z(n17411) );
  NANDN U18237 ( .A(n17412), .B(n17411), .Z(n17414) );
  XNOR U18238 ( .A(n17408), .B(n17407), .Z(n17409) );
  XNOR U18239 ( .A(n17410), .B(n17409), .Z(n17520) );
  XNOR U18240 ( .A(n17412), .B(n17411), .Z(n17519) );
  NAND U18241 ( .A(n17520), .B(n17519), .Z(n17413) );
  AND U18242 ( .A(n17414), .B(n17413), .Z(n17418) );
  NAND U18243 ( .A(n17418), .B(n17417), .Z(n17420) );
  XOR U18244 ( .A(n17418), .B(n17417), .Z(n17775) );
  NAND U18245 ( .A(a[49]), .B(b[15]), .Z(n17774) );
  NAND U18246 ( .A(n17775), .B(n17774), .Z(n17419) );
  AND U18247 ( .A(n17420), .B(n17419), .Z(n17781) );
  NANDN U18248 ( .A(n17423), .B(n17424), .Z(n17426) );
  XOR U18249 ( .A(n17422), .B(n17421), .Z(n17517) );
  XNOR U18250 ( .A(n17424), .B(n17423), .Z(n17518) );
  NANDN U18251 ( .A(n17517), .B(n17518), .Z(n17425) );
  AND U18252 ( .A(n17426), .B(n17425), .Z(n17430) );
  AND U18253 ( .A(a[52]), .B(b[15]), .Z(n17429) );
  NANDN U18254 ( .A(n17430), .B(n17429), .Z(n17432) );
  XOR U18255 ( .A(n17428), .B(n17427), .Z(n17790) );
  XNOR U18256 ( .A(n17430), .B(n17429), .Z(n17791) );
  NANDN U18257 ( .A(n17790), .B(n17791), .Z(n17431) );
  AND U18258 ( .A(n17432), .B(n17431), .Z(n17433) );
  NANDN U18259 ( .A(n17434), .B(n17433), .Z(n17438) );
  XOR U18260 ( .A(n17434), .B(n17433), .Z(n17513) );
  XOR U18261 ( .A(n17436), .B(n17435), .Z(n17514) );
  OR U18262 ( .A(n17513), .B(n17514), .Z(n17437) );
  AND U18263 ( .A(n17438), .B(n17437), .Z(n17442) );
  NANDN U18264 ( .A(n17441), .B(n17442), .Z(n17444) );
  XOR U18265 ( .A(n17440), .B(n17439), .Z(n17798) );
  XNOR U18266 ( .A(n17442), .B(n17441), .Z(n17799) );
  NANDN U18267 ( .A(n17798), .B(n17799), .Z(n17443) );
  AND U18268 ( .A(n17444), .B(n17443), .Z(n17448) );
  AND U18269 ( .A(a[55]), .B(b[15]), .Z(n17447) );
  NANDN U18270 ( .A(n17448), .B(n17447), .Z(n17450) );
  XOR U18271 ( .A(n17446), .B(n17445), .Z(n17509) );
  XNOR U18272 ( .A(n17448), .B(n17447), .Z(n17510) );
  NANDN U18273 ( .A(n17509), .B(n17510), .Z(n17449) );
  AND U18274 ( .A(n17450), .B(n17449), .Z(n17454) );
  AND U18275 ( .A(a[56]), .B(b[15]), .Z(n17453) );
  NANDN U18276 ( .A(n17454), .B(n17453), .Z(n17456) );
  XOR U18277 ( .A(n17452), .B(n17451), .Z(n17806) );
  XNOR U18278 ( .A(n17454), .B(n17453), .Z(n17807) );
  NANDN U18279 ( .A(n17806), .B(n17807), .Z(n17455) );
  AND U18280 ( .A(n17456), .B(n17455), .Z(n17505) );
  NAND U18281 ( .A(a[57]), .B(b[15]), .Z(n17506) );
  XOR U18282 ( .A(n17458), .B(n17457), .Z(n17508) );
  NANDN U18283 ( .A(n17461), .B(n17462), .Z(n17464) );
  XOR U18284 ( .A(n17460), .B(n17459), .Z(n17816) );
  XNOR U18285 ( .A(n17462), .B(n17461), .Z(n17817) );
  NANDN U18286 ( .A(n17816), .B(n17817), .Z(n17463) );
  AND U18287 ( .A(n17464), .B(n17463), .Z(n17465) );
  NANDN U18288 ( .A(n17466), .B(n17465), .Z(n17470) );
  XOR U18289 ( .A(n17466), .B(n17465), .Z(n17503) );
  XOR U18290 ( .A(n17468), .B(n17467), .Z(n17504) );
  NANDN U18291 ( .A(n17503), .B(n17504), .Z(n17469) );
  AND U18292 ( .A(n17470), .B(n17469), .Z(n17474) );
  NANDN U18293 ( .A(n17473), .B(n17474), .Z(n17476) );
  XOR U18294 ( .A(n17472), .B(n17471), .Z(n17824) );
  XNOR U18295 ( .A(n17474), .B(n17473), .Z(n17825) );
  NANDN U18296 ( .A(n17824), .B(n17825), .Z(n17475) );
  AND U18297 ( .A(n17476), .B(n17475), .Z(n17477) );
  NANDN U18298 ( .A(n17478), .B(n17477), .Z(n17482) );
  XOR U18299 ( .A(n17478), .B(n17477), .Z(n17501) );
  XOR U18300 ( .A(n17480), .B(n17479), .Z(n17502) );
  NANDN U18301 ( .A(n17501), .B(n17502), .Z(n17481) );
  AND U18302 ( .A(n17482), .B(n17481), .Z(n17486) );
  NANDN U18303 ( .A(n17485), .B(n17486), .Z(n17488) );
  XOR U18304 ( .A(n17484), .B(n17483), .Z(n17832) );
  XNOR U18305 ( .A(n17486), .B(n17485), .Z(n17833) );
  NANDN U18306 ( .A(n17832), .B(n17833), .Z(n17487) );
  AND U18307 ( .A(n17488), .B(n17487), .Z(n17489) );
  NANDN U18308 ( .A(n17490), .B(n17489), .Z(n17494) );
  XOR U18309 ( .A(n17490), .B(n17489), .Z(n17499) );
  XOR U18310 ( .A(n17492), .B(n17491), .Z(n17500) );
  NANDN U18311 ( .A(n17499), .B(n17500), .Z(n17493) );
  AND U18312 ( .A(n17494), .B(n17493), .Z(n22507) );
  XOR U18313 ( .A(n17496), .B(n17495), .Z(n22506) );
  ANDN U18314 ( .B(n22507), .A(n22506), .Z(n22508) );
  XNOR U18315 ( .A(n17498), .B(n17497), .Z(n22509) );
  XOR U18316 ( .A(n17500), .B(n17499), .Z(n18163) );
  XOR U18317 ( .A(n17502), .B(n17501), .Z(n17831) );
  AND U18318 ( .A(a[62]), .B(b[14]), .Z(n17830) );
  XOR U18319 ( .A(n17504), .B(n17503), .Z(n17823) );
  AND U18320 ( .A(a[60]), .B(b[14]), .Z(n17822) );
  NAND U18321 ( .A(a[58]), .B(b[14]), .Z(n17812) );
  XOR U18322 ( .A(n17506), .B(n17505), .Z(n17507) );
  XNOR U18323 ( .A(n17508), .B(n17507), .Z(n17813) );
  NANDN U18324 ( .A(n17812), .B(n17813), .Z(n17815) );
  NAND U18325 ( .A(a[56]), .B(b[14]), .Z(n17511) );
  XNOR U18326 ( .A(n17510), .B(n17509), .Z(n17512) );
  NANDN U18327 ( .A(n17511), .B(n17512), .Z(n17805) );
  XOR U18328 ( .A(n17512), .B(n17511), .Z(n18124) );
  XOR U18329 ( .A(n17514), .B(n17513), .Z(n17516) );
  AND U18330 ( .A(a[54]), .B(b[14]), .Z(n17515) );
  NANDN U18331 ( .A(n17516), .B(n17515), .Z(n17797) );
  XOR U18332 ( .A(n17516), .B(n17515), .Z(n18112) );
  NAND U18333 ( .A(a[52]), .B(b[14]), .Z(n17786) );
  XNOR U18334 ( .A(n17518), .B(n17517), .Z(n17787) );
  NANDN U18335 ( .A(n17786), .B(n17787), .Z(n17789) );
  XNOR U18336 ( .A(n17520), .B(n17519), .Z(n18092) );
  XNOR U18337 ( .A(n17522), .B(n17521), .Z(n18082) );
  XNOR U18338 ( .A(n17524), .B(n17523), .Z(n18074) );
  XNOR U18339 ( .A(n17526), .B(n17525), .Z(n18069) );
  AND U18340 ( .A(a[42]), .B(b[14]), .Z(n17742) );
  XNOR U18341 ( .A(n17528), .B(n17527), .Z(n18059) );
  NAND U18342 ( .A(a[40]), .B(b[14]), .Z(n17734) );
  AND U18343 ( .A(a[38]), .B(b[14]), .Z(n17727) );
  XOR U18344 ( .A(n17532), .B(n17531), .Z(n17723) );
  IV U18345 ( .A(n17723), .Z(n18048) );
  NAND U18346 ( .A(a[36]), .B(b[14]), .Z(n17851) );
  XOR U18347 ( .A(n17534), .B(n17533), .Z(n17535) );
  XOR U18348 ( .A(n17536), .B(n17535), .Z(n18034) );
  XNOR U18349 ( .A(n17538), .B(n17537), .Z(n18024) );
  XNOR U18350 ( .A(n17540), .B(n17539), .Z(n18016) );
  XNOR U18351 ( .A(n17542), .B(n17541), .Z(n18008) );
  XNOR U18352 ( .A(n17544), .B(n17543), .Z(n18000) );
  XNOR U18353 ( .A(n17546), .B(n17545), .Z(n17992) );
  XNOR U18354 ( .A(n17548), .B(n17547), .Z(n17984) );
  XNOR U18355 ( .A(n17550), .B(n17549), .Z(n17976) );
  XNOR U18356 ( .A(n17552), .B(n17551), .Z(n17968) );
  AND U18357 ( .A(a[8]), .B(b[14]), .Z(n17594) );
  XOR U18358 ( .A(n17554), .B(n17553), .Z(n17576) );
  AND U18359 ( .A(b[14]), .B(a[0]), .Z(n18224) );
  AND U18360 ( .A(a[1]), .B(b[15]), .Z(n17558) );
  AND U18361 ( .A(n18224), .B(n17558), .Z(n17555) );
  NAND U18362 ( .A(a[2]), .B(n17555), .Z(n17562) );
  NAND U18363 ( .A(b[15]), .B(a[1]), .Z(n17556) );
  XOR U18364 ( .A(n17557), .B(n17556), .Z(n17886) );
  NAND U18365 ( .A(n17558), .B(a[0]), .Z(n17559) );
  XNOR U18366 ( .A(a[2]), .B(n17559), .Z(n17560) );
  AND U18367 ( .A(b[14]), .B(n17560), .Z(n17887) );
  NANDN U18368 ( .A(n17886), .B(n17887), .Z(n17561) );
  AND U18369 ( .A(n17562), .B(n17561), .Z(n17566) );
  XNOR U18370 ( .A(n17564), .B(n17563), .Z(n17565) );
  NANDN U18371 ( .A(n17566), .B(n17565), .Z(n17568) );
  XNOR U18372 ( .A(n17566), .B(n17565), .Z(n17893) );
  AND U18373 ( .A(a[3]), .B(b[14]), .Z(n17892) );
  NAND U18374 ( .A(n17893), .B(n17892), .Z(n17567) );
  AND U18375 ( .A(n17568), .B(n17567), .Z(n17570) );
  AND U18376 ( .A(a[4]), .B(b[14]), .Z(n17569) );
  NANDN U18377 ( .A(n17570), .B(n17569), .Z(n17574) );
  XNOR U18378 ( .A(n17570), .B(n17569), .Z(n17899) );
  XNOR U18379 ( .A(n17572), .B(n17571), .Z(n17898) );
  NAND U18380 ( .A(n17899), .B(n17898), .Z(n17573) );
  NAND U18381 ( .A(n17574), .B(n17573), .Z(n17575) );
  NAND U18382 ( .A(n17576), .B(n17575), .Z(n17578) );
  NAND U18383 ( .A(a[5]), .B(b[14]), .Z(n17904) );
  XOR U18384 ( .A(n17576), .B(n17575), .Z(n17905) );
  NANDN U18385 ( .A(n17904), .B(n17905), .Z(n17577) );
  AND U18386 ( .A(n17578), .B(n17577), .Z(n17582) );
  XNOR U18387 ( .A(n17580), .B(n17579), .Z(n17581) );
  NANDN U18388 ( .A(n17582), .B(n17581), .Z(n17584) );
  NAND U18389 ( .A(a[6]), .B(b[14]), .Z(n17910) );
  XNOR U18390 ( .A(n17582), .B(n17581), .Z(n17911) );
  NANDN U18391 ( .A(n17910), .B(n17911), .Z(n17583) );
  AND U18392 ( .A(n17584), .B(n17583), .Z(n17588) );
  XNOR U18393 ( .A(n17586), .B(n17585), .Z(n17587) );
  NANDN U18394 ( .A(n17588), .B(n17587), .Z(n17590) );
  NAND U18395 ( .A(a[7]), .B(b[14]), .Z(n17918) );
  XNOR U18396 ( .A(n17588), .B(n17587), .Z(n17919) );
  NANDN U18397 ( .A(n17918), .B(n17919), .Z(n17589) );
  AND U18398 ( .A(n17590), .B(n17589), .Z(n17593) );
  NANDN U18399 ( .A(n17594), .B(n17593), .Z(n17596) );
  XOR U18400 ( .A(n17592), .B(n17591), .Z(n17877) );
  XNOR U18401 ( .A(n17594), .B(n17593), .Z(n17876) );
  NANDN U18402 ( .A(n17877), .B(n17876), .Z(n17595) );
  AND U18403 ( .A(n17596), .B(n17595), .Z(n17600) );
  XOR U18404 ( .A(n17598), .B(n17597), .Z(n17599) );
  NAND U18405 ( .A(n17600), .B(n17599), .Z(n17602) );
  NAND U18406 ( .A(a[9]), .B(b[14]), .Z(n17926) );
  XOR U18407 ( .A(n17600), .B(n17599), .Z(n17927) );
  NANDN U18408 ( .A(n17926), .B(n17927), .Z(n17601) );
  AND U18409 ( .A(n17602), .B(n17601), .Z(n17604) );
  AND U18410 ( .A(a[10]), .B(b[14]), .Z(n17603) );
  NANDN U18411 ( .A(n17604), .B(n17603), .Z(n17608) );
  XNOR U18412 ( .A(n17604), .B(n17603), .Z(n17933) );
  XNOR U18413 ( .A(n17606), .B(n17605), .Z(n17932) );
  NAND U18414 ( .A(n17933), .B(n17932), .Z(n17607) );
  AND U18415 ( .A(n17608), .B(n17607), .Z(n17612) );
  XOR U18416 ( .A(n17610), .B(n17609), .Z(n17611) );
  NANDN U18417 ( .A(n17612), .B(n17611), .Z(n17614) );
  NAND U18418 ( .A(a[11]), .B(b[14]), .Z(n17938) );
  XNOR U18419 ( .A(n17612), .B(n17611), .Z(n17939) );
  NANDN U18420 ( .A(n17938), .B(n17939), .Z(n17613) );
  AND U18421 ( .A(n17614), .B(n17613), .Z(n17616) );
  AND U18422 ( .A(a[12]), .B(b[14]), .Z(n17615) );
  NANDN U18423 ( .A(n17616), .B(n17615), .Z(n17620) );
  XNOR U18424 ( .A(n17616), .B(n17615), .Z(n17945) );
  XNOR U18425 ( .A(n17618), .B(n17617), .Z(n17944) );
  NAND U18426 ( .A(n17945), .B(n17944), .Z(n17619) );
  AND U18427 ( .A(n17620), .B(n17619), .Z(n17624) );
  XOR U18428 ( .A(n17622), .B(n17621), .Z(n17623) );
  NANDN U18429 ( .A(n17624), .B(n17623), .Z(n17626) );
  NAND U18430 ( .A(a[13]), .B(b[14]), .Z(n17950) );
  XNOR U18431 ( .A(n17624), .B(n17623), .Z(n17951) );
  NANDN U18432 ( .A(n17950), .B(n17951), .Z(n17625) );
  AND U18433 ( .A(n17626), .B(n17625), .Z(n17628) );
  AND U18434 ( .A(a[14]), .B(b[14]), .Z(n17627) );
  NANDN U18435 ( .A(n17628), .B(n17627), .Z(n17632) );
  XNOR U18436 ( .A(n17628), .B(n17627), .Z(n17957) );
  XNOR U18437 ( .A(n17630), .B(n17629), .Z(n17956) );
  NAND U18438 ( .A(n17957), .B(n17956), .Z(n17631) );
  AND U18439 ( .A(n17632), .B(n17631), .Z(n17636) );
  XOR U18440 ( .A(n17634), .B(n17633), .Z(n17635) );
  NANDN U18441 ( .A(n17636), .B(n17635), .Z(n17638) );
  NAND U18442 ( .A(a[15]), .B(b[14]), .Z(n17962) );
  XNOR U18443 ( .A(n17636), .B(n17635), .Z(n17963) );
  NANDN U18444 ( .A(n17962), .B(n17963), .Z(n17637) );
  AND U18445 ( .A(n17638), .B(n17637), .Z(n17640) );
  AND U18446 ( .A(a[16]), .B(b[14]), .Z(n17639) );
  NANDN U18447 ( .A(n17640), .B(n17639), .Z(n17644) );
  XNOR U18448 ( .A(n17640), .B(n17639), .Z(n17875) );
  XNOR U18449 ( .A(n17642), .B(n17641), .Z(n17874) );
  NAND U18450 ( .A(n17875), .B(n17874), .Z(n17643) );
  NAND U18451 ( .A(n17644), .B(n17643), .Z(n17969) );
  NAND U18452 ( .A(a[17]), .B(b[14]), .Z(n17971) );
  AND U18453 ( .A(a[18]), .B(b[14]), .Z(n17649) );
  NANDN U18454 ( .A(n17650), .B(n17649), .Z(n17652) );
  XNOR U18455 ( .A(n17646), .B(n17645), .Z(n17647) );
  XNOR U18456 ( .A(n17648), .B(n17647), .Z(n17873) );
  XNOR U18457 ( .A(n17650), .B(n17649), .Z(n17872) );
  NAND U18458 ( .A(n17873), .B(n17872), .Z(n17651) );
  NAND U18459 ( .A(n17652), .B(n17651), .Z(n17977) );
  NAND U18460 ( .A(a[19]), .B(b[14]), .Z(n17979) );
  AND U18461 ( .A(a[20]), .B(b[14]), .Z(n17653) );
  NANDN U18462 ( .A(n17654), .B(n17653), .Z(n17660) );
  XOR U18463 ( .A(n17654), .B(n17653), .Z(n17870) );
  XNOR U18464 ( .A(n17656), .B(n17655), .Z(n17657) );
  XNOR U18465 ( .A(n17658), .B(n17657), .Z(n17871) );
  NANDN U18466 ( .A(n17870), .B(n17871), .Z(n17659) );
  NAND U18467 ( .A(n17660), .B(n17659), .Z(n17985) );
  NAND U18468 ( .A(a[21]), .B(b[14]), .Z(n17987) );
  AND U18469 ( .A(a[22]), .B(b[14]), .Z(n17665) );
  NANDN U18470 ( .A(n17666), .B(n17665), .Z(n17668) );
  XNOR U18471 ( .A(n17662), .B(n17661), .Z(n17663) );
  XNOR U18472 ( .A(n17664), .B(n17663), .Z(n17869) );
  XNOR U18473 ( .A(n17666), .B(n17665), .Z(n17868) );
  NAND U18474 ( .A(n17869), .B(n17868), .Z(n17667) );
  NAND U18475 ( .A(n17668), .B(n17667), .Z(n17993) );
  NAND U18476 ( .A(a[23]), .B(b[14]), .Z(n17995) );
  AND U18477 ( .A(a[24]), .B(b[14]), .Z(n17673) );
  NANDN U18478 ( .A(n17674), .B(n17673), .Z(n17676) );
  XNOR U18479 ( .A(n17670), .B(n17669), .Z(n17671) );
  XNOR U18480 ( .A(n17672), .B(n17671), .Z(n17867) );
  XNOR U18481 ( .A(n17674), .B(n17673), .Z(n17866) );
  NAND U18482 ( .A(n17867), .B(n17866), .Z(n17675) );
  NAND U18483 ( .A(n17676), .B(n17675), .Z(n18001) );
  NAND U18484 ( .A(a[25]), .B(b[14]), .Z(n18003) );
  AND U18485 ( .A(a[26]), .B(b[14]), .Z(n17677) );
  NANDN U18486 ( .A(n17678), .B(n17677), .Z(n17684) );
  XOR U18487 ( .A(n17678), .B(n17677), .Z(n17864) );
  XNOR U18488 ( .A(n17680), .B(n17679), .Z(n17681) );
  XNOR U18489 ( .A(n17682), .B(n17681), .Z(n17865) );
  NANDN U18490 ( .A(n17864), .B(n17865), .Z(n17683) );
  NAND U18491 ( .A(n17684), .B(n17683), .Z(n18009) );
  NAND U18492 ( .A(a[27]), .B(b[14]), .Z(n18011) );
  AND U18493 ( .A(a[28]), .B(b[14]), .Z(n17689) );
  NANDN U18494 ( .A(n17690), .B(n17689), .Z(n17692) );
  XNOR U18495 ( .A(n17686), .B(n17685), .Z(n17687) );
  XNOR U18496 ( .A(n17688), .B(n17687), .Z(n17863) );
  XNOR U18497 ( .A(n17690), .B(n17689), .Z(n17862) );
  NAND U18498 ( .A(n17863), .B(n17862), .Z(n17691) );
  NAND U18499 ( .A(n17692), .B(n17691), .Z(n18017) );
  NAND U18500 ( .A(a[29]), .B(b[14]), .Z(n18019) );
  AND U18501 ( .A(a[30]), .B(b[14]), .Z(n17697) );
  NANDN U18502 ( .A(n17698), .B(n17697), .Z(n17700) );
  XNOR U18503 ( .A(n17694), .B(n17693), .Z(n17695) );
  XNOR U18504 ( .A(n17696), .B(n17695), .Z(n17861) );
  XNOR U18505 ( .A(n17698), .B(n17697), .Z(n17860) );
  NAND U18506 ( .A(n17861), .B(n17860), .Z(n17699) );
  NAND U18507 ( .A(n17700), .B(n17699), .Z(n18025) );
  NAND U18508 ( .A(a[31]), .B(b[14]), .Z(n18027) );
  AND U18509 ( .A(a[32]), .B(b[14]), .Z(n17705) );
  NANDN U18510 ( .A(n17706), .B(n17705), .Z(n17708) );
  XNOR U18511 ( .A(n17702), .B(n17701), .Z(n17703) );
  XNOR U18512 ( .A(n17704), .B(n17703), .Z(n17859) );
  XNOR U18513 ( .A(n17706), .B(n17705), .Z(n17858) );
  NAND U18514 ( .A(n17859), .B(n17858), .Z(n17707) );
  NAND U18515 ( .A(n17708), .B(n17707), .Z(n18035) );
  NAND U18516 ( .A(a[33]), .B(b[14]), .Z(n18036) );
  AND U18517 ( .A(a[34]), .B(b[14]), .Z(n17709) );
  IV U18518 ( .A(n17709), .Z(n17855) );
  OR U18519 ( .A(n17854), .B(n17855), .Z(n17715) );
  ANDN U18520 ( .B(n17854), .A(n17709), .Z(n17713) );
  OR U18521 ( .A(n17713), .B(n17857), .Z(n17714) );
  AND U18522 ( .A(n17715), .B(n17714), .Z(n18040) );
  NAND U18523 ( .A(a[35]), .B(b[14]), .Z(n18042) );
  XOR U18524 ( .A(n17720), .B(n17719), .Z(n17721) );
  XNOR U18525 ( .A(n17722), .B(n17721), .Z(n17853) );
  NANDN U18526 ( .A(n18048), .B(n18049), .Z(n17726) );
  NOR U18527 ( .A(n17723), .B(n18049), .Z(n17724) );
  AND U18528 ( .A(a[37]), .B(b[14]), .Z(n18047) );
  NANDN U18529 ( .A(n17724), .B(n18047), .Z(n17725) );
  AND U18530 ( .A(n17726), .B(n17725), .Z(n17728) );
  NANDN U18531 ( .A(n17727), .B(n17728), .Z(n17733) );
  NAND U18532 ( .A(n18050), .B(n18051), .Z(n17732) );
  NAND U18533 ( .A(n17733), .B(n17732), .Z(n18053) );
  AND U18534 ( .A(a[39]), .B(b[14]), .Z(n18054) );
  NANDN U18535 ( .A(n17734), .B(n17735), .Z(n17741) );
  XNOR U18536 ( .A(n17737), .B(n17736), .Z(n17738) );
  XNOR U18537 ( .A(n17739), .B(n17738), .Z(n17848) );
  NAND U18538 ( .A(n17849), .B(n17848), .Z(n17740) );
  NAND U18539 ( .A(n17741), .B(n17740), .Z(n18060) );
  NAND U18540 ( .A(a[41]), .B(b[14]), .Z(n18062) );
  NANDN U18541 ( .A(n17742), .B(n17743), .Z(n17748) );
  NAND U18542 ( .A(n17846), .B(n17847), .Z(n17747) );
  AND U18543 ( .A(n17748), .B(n17747), .Z(n18068) );
  AND U18544 ( .A(a[43]), .B(b[14]), .Z(n18067) );
  AND U18545 ( .A(a[44]), .B(b[14]), .Z(n17750) );
  NANDN U18546 ( .A(n17749), .B(n17750), .Z(n17756) );
  XNOR U18547 ( .A(n17750), .B(n17749), .Z(n17845) );
  XNOR U18548 ( .A(n17752), .B(n17751), .Z(n17753) );
  XNOR U18549 ( .A(n17754), .B(n17753), .Z(n17844) );
  NAND U18550 ( .A(n17845), .B(n17844), .Z(n17755) );
  NAND U18551 ( .A(n17756), .B(n17755), .Z(n18075) );
  NAND U18552 ( .A(a[45]), .B(b[14]), .Z(n18077) );
  AND U18553 ( .A(a[46]), .B(b[14]), .Z(n17761) );
  NANDN U18554 ( .A(n17760), .B(n17761), .Z(n17763) );
  XNOR U18555 ( .A(n17761), .B(n17760), .Z(n17842) );
  NAND U18556 ( .A(n17843), .B(n17842), .Z(n17762) );
  NAND U18557 ( .A(n17763), .B(n17762), .Z(n18083) );
  NAND U18558 ( .A(a[47]), .B(b[14]), .Z(n18085) );
  AND U18559 ( .A(a[48]), .B(b[14]), .Z(n17769) );
  NANDN U18560 ( .A(n17768), .B(n17769), .Z(n17771) );
  XNOR U18561 ( .A(n17765), .B(n17764), .Z(n17766) );
  XNOR U18562 ( .A(n17767), .B(n17766), .Z(n17841) );
  XNOR U18563 ( .A(n17769), .B(n17768), .Z(n17840) );
  NAND U18564 ( .A(n17841), .B(n17840), .Z(n17770) );
  NAND U18565 ( .A(n17771), .B(n17770), .Z(n18093) );
  NAND U18566 ( .A(a[49]), .B(b[14]), .Z(n18095) );
  AND U18567 ( .A(a[50]), .B(b[14]), .Z(n17772) );
  NANDN U18568 ( .A(n17773), .B(n17772), .Z(n17777) );
  XOR U18569 ( .A(n17773), .B(n17772), .Z(n18098) );
  XNOR U18570 ( .A(n17775), .B(n17774), .Z(n18099) );
  NANDN U18571 ( .A(n18098), .B(n18099), .Z(n17776) );
  AND U18572 ( .A(n17777), .B(n17776), .Z(n17783) );
  AND U18573 ( .A(a[51]), .B(b[14]), .Z(n17782) );
  NANDN U18574 ( .A(n17783), .B(n17782), .Z(n17785) );
  XOR U18575 ( .A(n17779), .B(n17778), .Z(n17780) );
  XNOR U18576 ( .A(n17781), .B(n17780), .Z(n17839) );
  XNOR U18577 ( .A(n17783), .B(n17782), .Z(n17838) );
  NAND U18578 ( .A(n17839), .B(n17838), .Z(n17784) );
  AND U18579 ( .A(n17785), .B(n17784), .Z(n18105) );
  XNOR U18580 ( .A(n17787), .B(n17786), .Z(n18104) );
  NANDN U18581 ( .A(n18105), .B(n18104), .Z(n17788) );
  AND U18582 ( .A(n17789), .B(n17788), .Z(n17793) );
  XNOR U18583 ( .A(n17791), .B(n17790), .Z(n17792) );
  NANDN U18584 ( .A(n17793), .B(n17792), .Z(n17795) );
  NAND U18585 ( .A(a[53]), .B(b[14]), .Z(n18106) );
  XNOR U18586 ( .A(n17793), .B(n17792), .Z(n18107) );
  NANDN U18587 ( .A(n18106), .B(n18107), .Z(n17794) );
  AND U18588 ( .A(n17795), .B(n17794), .Z(n18113) );
  OR U18589 ( .A(n18112), .B(n18113), .Z(n17796) );
  AND U18590 ( .A(n17797), .B(n17796), .Z(n17801) );
  XNOR U18591 ( .A(n17799), .B(n17798), .Z(n17800) );
  NANDN U18592 ( .A(n17801), .B(n17800), .Z(n17803) );
  NAND U18593 ( .A(a[55]), .B(b[14]), .Z(n18118) );
  XNOR U18594 ( .A(n17801), .B(n17800), .Z(n18119) );
  NANDN U18595 ( .A(n18118), .B(n18119), .Z(n17802) );
  AND U18596 ( .A(n17803), .B(n17802), .Z(n18125) );
  OR U18597 ( .A(n18124), .B(n18125), .Z(n17804) );
  AND U18598 ( .A(n17805), .B(n17804), .Z(n17809) );
  XNOR U18599 ( .A(n17807), .B(n17806), .Z(n17808) );
  NANDN U18600 ( .A(n17809), .B(n17808), .Z(n17811) );
  NAND U18601 ( .A(a[57]), .B(b[14]), .Z(n18130) );
  XNOR U18602 ( .A(n17809), .B(n17808), .Z(n18131) );
  NANDN U18603 ( .A(n18130), .B(n18131), .Z(n17810) );
  AND U18604 ( .A(n17811), .B(n17810), .Z(n18137) );
  XNOR U18605 ( .A(n17813), .B(n17812), .Z(n18136) );
  NANDN U18606 ( .A(n18137), .B(n18136), .Z(n17814) );
  AND U18607 ( .A(n17815), .B(n17814), .Z(n17819) );
  XNOR U18608 ( .A(n17817), .B(n17816), .Z(n17818) );
  NANDN U18609 ( .A(n17819), .B(n17818), .Z(n17821) );
  NAND U18610 ( .A(a[59]), .B(b[14]), .Z(n18142) );
  XNOR U18611 ( .A(n17819), .B(n17818), .Z(n18143) );
  NANDN U18612 ( .A(n18142), .B(n18143), .Z(n17820) );
  AND U18613 ( .A(n17821), .B(n17820), .Z(n18149) );
  XOR U18614 ( .A(n17823), .B(n17822), .Z(n18148) );
  XNOR U18615 ( .A(n17825), .B(n17824), .Z(n17826) );
  NANDN U18616 ( .A(n17827), .B(n17826), .Z(n17829) );
  NAND U18617 ( .A(a[61]), .B(b[14]), .Z(n18152) );
  XNOR U18618 ( .A(n17827), .B(n17826), .Z(n18153) );
  NANDN U18619 ( .A(n18152), .B(n18153), .Z(n17828) );
  AND U18620 ( .A(n17829), .B(n17828), .Z(n18157) );
  XOR U18621 ( .A(n17831), .B(n17830), .Z(n18156) );
  XNOR U18622 ( .A(n17833), .B(n17832), .Z(n17834) );
  NANDN U18623 ( .A(n17835), .B(n17834), .Z(n17837) );
  NAND U18624 ( .A(a[63]), .B(b[14]), .Z(n18160) );
  XNOR U18625 ( .A(n17835), .B(n17834), .Z(n18161) );
  NANDN U18626 ( .A(n18160), .B(n18161), .Z(n17836) );
  AND U18627 ( .A(n17837), .B(n17836), .Z(n18162) );
  AND U18628 ( .A(a[63]), .B(b[13]), .Z(n18159) );
  NAND U18629 ( .A(a[62]), .B(b[13]), .Z(n18150) );
  NAND U18630 ( .A(a[58]), .B(b[13]), .Z(n18132) );
  AND U18631 ( .A(a[57]), .B(b[13]), .Z(n18127) );
  NAND U18632 ( .A(a[56]), .B(b[13]), .Z(n18120) );
  AND U18633 ( .A(a[55]), .B(b[13]), .Z(n18115) );
  NAND U18634 ( .A(a[54]), .B(b[13]), .Z(n18108) );
  NAND U18635 ( .A(a[53]), .B(b[13]), .Z(n18179) );
  XNOR U18636 ( .A(n17839), .B(n17838), .Z(n18458) );
  AND U18637 ( .A(a[52]), .B(b[13]), .Z(n18457) );
  XNOR U18638 ( .A(n17841), .B(n17840), .Z(n18442) );
  XNOR U18639 ( .A(n17843), .B(n17842), .Z(n18432) );
  XNOR U18640 ( .A(n17845), .B(n17844), .Z(n18425) );
  XOR U18641 ( .A(n17847), .B(n17846), .Z(n18415) );
  XNOR U18642 ( .A(n17849), .B(n17848), .Z(n18409) );
  NAND U18643 ( .A(a[40]), .B(b[13]), .Z(n18055) );
  NAND U18644 ( .A(a[38]), .B(b[13]), .Z(n18194) );
  XOR U18645 ( .A(n17851), .B(n17850), .Z(n17852) );
  XOR U18646 ( .A(n17853), .B(n17852), .Z(n18043) );
  IV U18647 ( .A(n18043), .Z(n18395) );
  NAND U18648 ( .A(a[36]), .B(b[13]), .Z(n18198) );
  XOR U18649 ( .A(n17855), .B(n17854), .Z(n17856) );
  XOR U18650 ( .A(n17857), .B(n17856), .Z(n18386) );
  XNOR U18651 ( .A(n17859), .B(n17858), .Z(n18378) );
  XNOR U18652 ( .A(n17861), .B(n17860), .Z(n18370) );
  XNOR U18653 ( .A(n17863), .B(n17862), .Z(n18362) );
  NAND U18654 ( .A(a[28]), .B(b[13]), .Z(n18012) );
  XNOR U18655 ( .A(n17865), .B(n17864), .Z(n18355) );
  XNOR U18656 ( .A(n17867), .B(n17866), .Z(n18346) );
  XNOR U18657 ( .A(n17869), .B(n17868), .Z(n18340) );
  NAND U18658 ( .A(a[22]), .B(b[13]), .Z(n17988) );
  XNOR U18659 ( .A(n17871), .B(n17870), .Z(n18331) );
  XNOR U18660 ( .A(n17873), .B(n17872), .Z(n18322) );
  XNOR U18661 ( .A(n17875), .B(n17874), .Z(n18312) );
  XOR U18662 ( .A(n17877), .B(n17876), .Z(n17923) );
  AND U18663 ( .A(a[4]), .B(b[13]), .Z(n17895) );
  AND U18664 ( .A(b[13]), .B(a[0]), .Z(n18533) );
  AND U18665 ( .A(a[1]), .B(b[14]), .Z(n17881) );
  AND U18666 ( .A(n18533), .B(n17881), .Z(n17878) );
  NAND U18667 ( .A(a[2]), .B(n17878), .Z(n17885) );
  NAND U18668 ( .A(b[14]), .B(a[1]), .Z(n17879) );
  XOR U18669 ( .A(n17880), .B(n17879), .Z(n18230) );
  NAND U18670 ( .A(n17881), .B(a[0]), .Z(n17882) );
  XNOR U18671 ( .A(a[2]), .B(n17882), .Z(n17883) );
  AND U18672 ( .A(b[13]), .B(n17883), .Z(n18231) );
  NANDN U18673 ( .A(n18230), .B(n18231), .Z(n17884) );
  AND U18674 ( .A(n17885), .B(n17884), .Z(n17889) );
  XNOR U18675 ( .A(n17887), .B(n17886), .Z(n17888) );
  NANDN U18676 ( .A(n17889), .B(n17888), .Z(n17891) );
  NAND U18677 ( .A(a[3]), .B(b[13]), .Z(n18238) );
  XNOR U18678 ( .A(n17889), .B(n17888), .Z(n18239) );
  NANDN U18679 ( .A(n18238), .B(n18239), .Z(n17890) );
  AND U18680 ( .A(n17891), .B(n17890), .Z(n17894) );
  NANDN U18681 ( .A(n17895), .B(n17894), .Z(n17897) );
  XOR U18682 ( .A(n17893), .B(n17892), .Z(n18221) );
  XNOR U18683 ( .A(n17895), .B(n17894), .Z(n18220) );
  NANDN U18684 ( .A(n18221), .B(n18220), .Z(n17896) );
  AND U18685 ( .A(n17897), .B(n17896), .Z(n17901) );
  XOR U18686 ( .A(n17899), .B(n17898), .Z(n17900) );
  NAND U18687 ( .A(n17901), .B(n17900), .Z(n17903) );
  NAND U18688 ( .A(a[5]), .B(b[13]), .Z(n18246) );
  XOR U18689 ( .A(n17901), .B(n17900), .Z(n18247) );
  NANDN U18690 ( .A(n18246), .B(n18247), .Z(n17902) );
  AND U18691 ( .A(n17903), .B(n17902), .Z(n17907) );
  XNOR U18692 ( .A(n17905), .B(n17904), .Z(n17906) );
  NANDN U18693 ( .A(n17907), .B(n17906), .Z(n17909) );
  NAND U18694 ( .A(a[6]), .B(b[13]), .Z(n18252) );
  XNOR U18695 ( .A(n17907), .B(n17906), .Z(n18253) );
  NANDN U18696 ( .A(n18252), .B(n18253), .Z(n17908) );
  AND U18697 ( .A(n17909), .B(n17908), .Z(n17913) );
  XNOR U18698 ( .A(n17911), .B(n17910), .Z(n17912) );
  NANDN U18699 ( .A(n17913), .B(n17912), .Z(n17915) );
  XNOR U18700 ( .A(n17913), .B(n17912), .Z(n18259) );
  AND U18701 ( .A(a[7]), .B(b[13]), .Z(n18258) );
  NAND U18702 ( .A(n18259), .B(n18258), .Z(n17914) );
  AND U18703 ( .A(n17915), .B(n17914), .Z(n17917) );
  AND U18704 ( .A(a[8]), .B(b[13]), .Z(n17916) );
  NANDN U18705 ( .A(n17917), .B(n17916), .Z(n17921) );
  XNOR U18706 ( .A(n17917), .B(n17916), .Z(n18265) );
  XNOR U18707 ( .A(n17919), .B(n17918), .Z(n18264) );
  NAND U18708 ( .A(n18265), .B(n18264), .Z(n17920) );
  NAND U18709 ( .A(n17921), .B(n17920), .Z(n17922) );
  NAND U18710 ( .A(n17923), .B(n17922), .Z(n17925) );
  NAND U18711 ( .A(a[9]), .B(b[13]), .Z(n18272) );
  XOR U18712 ( .A(n17923), .B(n17922), .Z(n18273) );
  NANDN U18713 ( .A(n18272), .B(n18273), .Z(n17924) );
  AND U18714 ( .A(n17925), .B(n17924), .Z(n17929) );
  AND U18715 ( .A(a[10]), .B(b[13]), .Z(n17928) );
  NANDN U18716 ( .A(n17929), .B(n17928), .Z(n17931) );
  XNOR U18717 ( .A(n17927), .B(n17926), .Z(n18277) );
  XNOR U18718 ( .A(n17929), .B(n17928), .Z(n18276) );
  NAND U18719 ( .A(n18277), .B(n18276), .Z(n17930) );
  AND U18720 ( .A(n17931), .B(n17930), .Z(n17935) );
  XOR U18721 ( .A(n17933), .B(n17932), .Z(n17934) );
  NANDN U18722 ( .A(n17935), .B(n17934), .Z(n17937) );
  NAND U18723 ( .A(a[11]), .B(b[13]), .Z(n18284) );
  XNOR U18724 ( .A(n17935), .B(n17934), .Z(n18285) );
  NANDN U18725 ( .A(n18284), .B(n18285), .Z(n17936) );
  AND U18726 ( .A(n17937), .B(n17936), .Z(n17941) );
  AND U18727 ( .A(a[12]), .B(b[13]), .Z(n17940) );
  NANDN U18728 ( .A(n17941), .B(n17940), .Z(n17943) );
  XNOR U18729 ( .A(n17939), .B(n17938), .Z(n18289) );
  XNOR U18730 ( .A(n17941), .B(n17940), .Z(n18288) );
  NAND U18731 ( .A(n18289), .B(n18288), .Z(n17942) );
  AND U18732 ( .A(n17943), .B(n17942), .Z(n17947) );
  XOR U18733 ( .A(n17945), .B(n17944), .Z(n17946) );
  NANDN U18734 ( .A(n17947), .B(n17946), .Z(n17949) );
  NAND U18735 ( .A(a[13]), .B(b[13]), .Z(n18296) );
  XNOR U18736 ( .A(n17947), .B(n17946), .Z(n18297) );
  NANDN U18737 ( .A(n18296), .B(n18297), .Z(n17948) );
  AND U18738 ( .A(n17949), .B(n17948), .Z(n17953) );
  AND U18739 ( .A(a[14]), .B(b[13]), .Z(n17952) );
  NANDN U18740 ( .A(n17953), .B(n17952), .Z(n17955) );
  XNOR U18741 ( .A(n17951), .B(n17950), .Z(n18301) );
  XNOR U18742 ( .A(n17953), .B(n17952), .Z(n18300) );
  NAND U18743 ( .A(n18301), .B(n18300), .Z(n17954) );
  AND U18744 ( .A(n17955), .B(n17954), .Z(n17959) );
  XOR U18745 ( .A(n17957), .B(n17956), .Z(n17958) );
  NANDN U18746 ( .A(n17959), .B(n17958), .Z(n17961) );
  NAND U18747 ( .A(a[15]), .B(b[13]), .Z(n18308) );
  XNOR U18748 ( .A(n17959), .B(n17958), .Z(n18309) );
  NANDN U18749 ( .A(n18308), .B(n18309), .Z(n17960) );
  AND U18750 ( .A(n17961), .B(n17960), .Z(n17965) );
  AND U18751 ( .A(a[16]), .B(b[13]), .Z(n17964) );
  NANDN U18752 ( .A(n17965), .B(n17964), .Z(n17967) );
  XNOR U18753 ( .A(n17963), .B(n17962), .Z(n18219) );
  XNOR U18754 ( .A(n17965), .B(n17964), .Z(n18218) );
  NAND U18755 ( .A(n18219), .B(n18218), .Z(n17966) );
  NAND U18756 ( .A(n17967), .B(n17966), .Z(n18313) );
  NAND U18757 ( .A(a[17]), .B(b[13]), .Z(n18315) );
  AND U18758 ( .A(a[18]), .B(b[13]), .Z(n17972) );
  NANDN U18759 ( .A(n17973), .B(n17972), .Z(n17975) );
  XNOR U18760 ( .A(n17969), .B(n17968), .Z(n17970) );
  XNOR U18761 ( .A(n17971), .B(n17970), .Z(n18217) );
  XNOR U18762 ( .A(n17973), .B(n17972), .Z(n18216) );
  NAND U18763 ( .A(n18217), .B(n18216), .Z(n17974) );
  NAND U18764 ( .A(n17975), .B(n17974), .Z(n18323) );
  AND U18765 ( .A(a[19]), .B(b[13]), .Z(n18325) );
  AND U18766 ( .A(a[20]), .B(b[13]), .Z(n17980) );
  NANDN U18767 ( .A(n17981), .B(n17980), .Z(n17983) );
  XNOR U18768 ( .A(n17977), .B(n17976), .Z(n17978) );
  XNOR U18769 ( .A(n17979), .B(n17978), .Z(n18329) );
  XNOR U18770 ( .A(n17981), .B(n17980), .Z(n18328) );
  NAND U18771 ( .A(n18329), .B(n18328), .Z(n17982) );
  AND U18772 ( .A(n17983), .B(n17982), .Z(n18330) );
  NAND U18773 ( .A(a[21]), .B(b[13]), .Z(n18333) );
  NANDN U18774 ( .A(n17988), .B(n17989), .Z(n17991) );
  XNOR U18775 ( .A(n17985), .B(n17984), .Z(n17986) );
  XNOR U18776 ( .A(n17987), .B(n17986), .Z(n18215) );
  XNOR U18777 ( .A(n17989), .B(n17988), .Z(n18214) );
  NAND U18778 ( .A(n18215), .B(n18214), .Z(n17990) );
  NAND U18779 ( .A(n17991), .B(n17990), .Z(n18341) );
  NAND U18780 ( .A(a[23]), .B(b[13]), .Z(n18343) );
  AND U18781 ( .A(a[24]), .B(b[13]), .Z(n17996) );
  NANDN U18782 ( .A(n17997), .B(n17996), .Z(n17999) );
  XNOR U18783 ( .A(n17993), .B(n17992), .Z(n17994) );
  XNOR U18784 ( .A(n17995), .B(n17994), .Z(n18213) );
  XNOR U18785 ( .A(n17997), .B(n17996), .Z(n18212) );
  NAND U18786 ( .A(n18213), .B(n18212), .Z(n17998) );
  NAND U18787 ( .A(n17999), .B(n17998), .Z(n18347) );
  NAND U18788 ( .A(a[25]), .B(b[13]), .Z(n18349) );
  AND U18789 ( .A(a[26]), .B(b[13]), .Z(n18004) );
  NANDN U18790 ( .A(n18005), .B(n18004), .Z(n18007) );
  XNOR U18791 ( .A(n18001), .B(n18000), .Z(n18002) );
  XNOR U18792 ( .A(n18003), .B(n18002), .Z(n18211) );
  XNOR U18793 ( .A(n18005), .B(n18004), .Z(n18210) );
  NAND U18794 ( .A(n18211), .B(n18210), .Z(n18006) );
  AND U18795 ( .A(n18007), .B(n18006), .Z(n18354) );
  NAND U18796 ( .A(a[27]), .B(b[13]), .Z(n18357) );
  NANDN U18797 ( .A(n18012), .B(n18013), .Z(n18015) );
  XNOR U18798 ( .A(n18009), .B(n18008), .Z(n18010) );
  XNOR U18799 ( .A(n18011), .B(n18010), .Z(n18209) );
  XNOR U18800 ( .A(n18013), .B(n18012), .Z(n18208) );
  NAND U18801 ( .A(n18209), .B(n18208), .Z(n18014) );
  NAND U18802 ( .A(n18015), .B(n18014), .Z(n18363) );
  NAND U18803 ( .A(a[29]), .B(b[13]), .Z(n18365) );
  AND U18804 ( .A(a[30]), .B(b[13]), .Z(n18020) );
  NANDN U18805 ( .A(n18021), .B(n18020), .Z(n18023) );
  XNOR U18806 ( .A(n18017), .B(n18016), .Z(n18018) );
  XNOR U18807 ( .A(n18019), .B(n18018), .Z(n18207) );
  XNOR U18808 ( .A(n18021), .B(n18020), .Z(n18206) );
  NAND U18809 ( .A(n18207), .B(n18206), .Z(n18022) );
  NAND U18810 ( .A(n18023), .B(n18022), .Z(n18371) );
  NAND U18811 ( .A(a[31]), .B(b[13]), .Z(n18373) );
  AND U18812 ( .A(a[32]), .B(b[13]), .Z(n18028) );
  NANDN U18813 ( .A(n18029), .B(n18028), .Z(n18031) );
  XNOR U18814 ( .A(n18025), .B(n18024), .Z(n18026) );
  XNOR U18815 ( .A(n18027), .B(n18026), .Z(n18205) );
  XNOR U18816 ( .A(n18029), .B(n18028), .Z(n18204) );
  NAND U18817 ( .A(n18205), .B(n18204), .Z(n18030) );
  NAND U18818 ( .A(n18031), .B(n18030), .Z(n18379) );
  NAND U18819 ( .A(a[33]), .B(b[13]), .Z(n18381) );
  AND U18820 ( .A(a[34]), .B(b[13]), .Z(n18032) );
  NANDN U18821 ( .A(n18033), .B(n18032), .Z(n18038) );
  XNOR U18822 ( .A(n18033), .B(n18032), .Z(n18203) );
  NAND U18823 ( .A(n18203), .B(n18202), .Z(n18037) );
  NAND U18824 ( .A(n18038), .B(n18037), .Z(n18387) );
  NAND U18825 ( .A(a[35]), .B(b[13]), .Z(n18388) );
  XOR U18826 ( .A(n18040), .B(n18039), .Z(n18041) );
  XNOR U18827 ( .A(n18042), .B(n18041), .Z(n18201) );
  NANDN U18828 ( .A(n18395), .B(n18394), .Z(n18046) );
  NOR U18829 ( .A(n18043), .B(n18394), .Z(n18044) );
  AND U18830 ( .A(a[37]), .B(b[13]), .Z(n18393) );
  NANDN U18831 ( .A(n18044), .B(n18393), .Z(n18045) );
  AND U18832 ( .A(n18046), .B(n18045), .Z(n18195) );
  XNOR U18833 ( .A(n18051), .B(n18050), .Z(n18401) );
  NAND U18834 ( .A(a[39]), .B(b[13]), .Z(n18400) );
  NANDN U18835 ( .A(n18055), .B(n18056), .Z(n18058) );
  NAND U18836 ( .A(n18193), .B(n18192), .Z(n18057) );
  NAND U18837 ( .A(n18058), .B(n18057), .Z(n18410) );
  NAND U18838 ( .A(a[41]), .B(b[13]), .Z(n18412) );
  AND U18839 ( .A(a[42]), .B(b[13]), .Z(n18063) );
  NANDN U18840 ( .A(n18064), .B(n18063), .Z(n18066) );
  XNOR U18841 ( .A(n18060), .B(n18059), .Z(n18061) );
  XNOR U18842 ( .A(n18062), .B(n18061), .Z(n18191) );
  XNOR U18843 ( .A(n18064), .B(n18063), .Z(n18190) );
  NAND U18844 ( .A(n18191), .B(n18190), .Z(n18065) );
  NAND U18845 ( .A(n18066), .B(n18065), .Z(n18416) );
  NAND U18846 ( .A(a[43]), .B(b[13]), .Z(n18418) );
  AND U18847 ( .A(a[44]), .B(b[13]), .Z(n18070) );
  NANDN U18848 ( .A(n18071), .B(n18070), .Z(n18073) );
  XNOR U18849 ( .A(n18071), .B(n18070), .Z(n18188) );
  NAND U18850 ( .A(n18189), .B(n18188), .Z(n18072) );
  NAND U18851 ( .A(n18073), .B(n18072), .Z(n18426) );
  NAND U18852 ( .A(a[45]), .B(b[13]), .Z(n18428) );
  AND U18853 ( .A(a[46]), .B(b[13]), .Z(n18078) );
  NANDN U18854 ( .A(n18079), .B(n18078), .Z(n18081) );
  XNOR U18855 ( .A(n18075), .B(n18074), .Z(n18076) );
  XNOR U18856 ( .A(n18077), .B(n18076), .Z(n18187) );
  XNOR U18857 ( .A(n18079), .B(n18078), .Z(n18186) );
  NAND U18858 ( .A(n18187), .B(n18186), .Z(n18080) );
  NAND U18859 ( .A(n18081), .B(n18080), .Z(n18433) );
  NAND U18860 ( .A(a[47]), .B(b[13]), .Z(n18435) );
  AND U18861 ( .A(a[48]), .B(b[13]), .Z(n18086) );
  NANDN U18862 ( .A(n18087), .B(n18086), .Z(n18089) );
  XNOR U18863 ( .A(n18083), .B(n18082), .Z(n18084) );
  XNOR U18864 ( .A(n18085), .B(n18084), .Z(n18185) );
  XNOR U18865 ( .A(n18087), .B(n18086), .Z(n18184) );
  NAND U18866 ( .A(n18185), .B(n18184), .Z(n18088) );
  NAND U18867 ( .A(n18089), .B(n18088), .Z(n18443) );
  AND U18868 ( .A(a[49]), .B(b[13]), .Z(n18441) );
  AND U18869 ( .A(a[50]), .B(b[13]), .Z(n18090) );
  NANDN U18870 ( .A(n18091), .B(n18090), .Z(n18097) );
  XNOR U18871 ( .A(n18091), .B(n18090), .Z(n18183) );
  XNOR U18872 ( .A(n18093), .B(n18092), .Z(n18094) );
  XNOR U18873 ( .A(n18095), .B(n18094), .Z(n18182) );
  NAND U18874 ( .A(n18183), .B(n18182), .Z(n18096) );
  AND U18875 ( .A(n18097), .B(n18096), .Z(n18101) );
  NAND U18876 ( .A(n18101), .B(n18100), .Z(n18103) );
  AND U18877 ( .A(a[51]), .B(b[13]), .Z(n18449) );
  XOR U18878 ( .A(n18101), .B(n18100), .Z(n18450) );
  NANDN U18879 ( .A(n18449), .B(n18450), .Z(n18102) );
  AND U18880 ( .A(n18103), .B(n18102), .Z(n18460) );
  XOR U18881 ( .A(n18105), .B(n18104), .Z(n18181) );
  NANDN U18882 ( .A(n18108), .B(n18109), .Z(n18111) );
  XOR U18883 ( .A(n18107), .B(n18106), .Z(n18463) );
  XNOR U18884 ( .A(n18109), .B(n18108), .Z(n18464) );
  NANDN U18885 ( .A(n18463), .B(n18464), .Z(n18110) );
  AND U18886 ( .A(n18111), .B(n18110), .Z(n18114) );
  NANDN U18887 ( .A(n18115), .B(n18114), .Z(n18117) );
  XOR U18888 ( .A(n18113), .B(n18112), .Z(n18177) );
  XNOR U18889 ( .A(n18115), .B(n18114), .Z(n18176) );
  NANDN U18890 ( .A(n18177), .B(n18176), .Z(n18116) );
  AND U18891 ( .A(n18117), .B(n18116), .Z(n18121) );
  NANDN U18892 ( .A(n18120), .B(n18121), .Z(n18123) );
  XOR U18893 ( .A(n18119), .B(n18118), .Z(n18469) );
  XNOR U18894 ( .A(n18121), .B(n18120), .Z(n18470) );
  NANDN U18895 ( .A(n18469), .B(n18470), .Z(n18122) );
  AND U18896 ( .A(n18123), .B(n18122), .Z(n18126) );
  NANDN U18897 ( .A(n18127), .B(n18126), .Z(n18129) );
  XOR U18898 ( .A(n18125), .B(n18124), .Z(n18175) );
  XNOR U18899 ( .A(n18127), .B(n18126), .Z(n18174) );
  NANDN U18900 ( .A(n18175), .B(n18174), .Z(n18128) );
  AND U18901 ( .A(n18129), .B(n18128), .Z(n18133) );
  NANDN U18902 ( .A(n18132), .B(n18133), .Z(n18135) );
  XOR U18903 ( .A(n18131), .B(n18130), .Z(n18475) );
  XNOR U18904 ( .A(n18133), .B(n18132), .Z(n18476) );
  NANDN U18905 ( .A(n18475), .B(n18476), .Z(n18134) );
  AND U18906 ( .A(n18135), .B(n18134), .Z(n18139) );
  AND U18907 ( .A(a[59]), .B(b[13]), .Z(n18138) );
  NANDN U18908 ( .A(n18139), .B(n18138), .Z(n18141) );
  XOR U18909 ( .A(n18137), .B(n18136), .Z(n18172) );
  XNOR U18910 ( .A(n18139), .B(n18138), .Z(n18173) );
  NANDN U18911 ( .A(n18172), .B(n18173), .Z(n18140) );
  AND U18912 ( .A(n18141), .B(n18140), .Z(n18145) );
  AND U18913 ( .A(a[60]), .B(b[13]), .Z(n18144) );
  NANDN U18914 ( .A(n18145), .B(n18144), .Z(n18147) );
  XOR U18915 ( .A(n18143), .B(n18142), .Z(n18481) );
  XNOR U18916 ( .A(n18145), .B(n18144), .Z(n18482) );
  NANDN U18917 ( .A(n18481), .B(n18482), .Z(n18146) );
  AND U18918 ( .A(n18147), .B(n18146), .Z(n18168) );
  NAND U18919 ( .A(a[61]), .B(b[13]), .Z(n18169) );
  XOR U18920 ( .A(n18149), .B(n18148), .Z(n18171) );
  NANDN U18921 ( .A(n18150), .B(n18151), .Z(n18155) );
  XNOR U18922 ( .A(n18151), .B(n18150), .Z(n18167) );
  XNOR U18923 ( .A(n18153), .B(n18152), .Z(n18166) );
  NAND U18924 ( .A(n18167), .B(n18166), .Z(n18154) );
  AND U18925 ( .A(n18155), .B(n18154), .Z(n18158) );
  XOR U18926 ( .A(n18157), .B(n18156), .Z(n18488) );
  XNOR U18927 ( .A(n18159), .B(n18158), .Z(n18487) );
  XNOR U18928 ( .A(n18161), .B(n18160), .Z(n18489) );
  AND U18929 ( .A(n18490), .B(n18489), .Z(n18165) );
  XOR U18930 ( .A(n18163), .B(n18162), .Z(n18164) );
  NANDN U18931 ( .A(n18165), .B(n18164), .Z(n22505) );
  XNOR U18932 ( .A(n18165), .B(n18164), .Z(n24720) );
  XOR U18933 ( .A(n18167), .B(n18166), .Z(n18485) );
  AND U18934 ( .A(a[62]), .B(b[12]), .Z(n18810) );
  XOR U18935 ( .A(n18169), .B(n18168), .Z(n18170) );
  XOR U18936 ( .A(n18171), .B(n18170), .Z(n18813) );
  AND U18937 ( .A(a[60]), .B(b[12]), .Z(n18479) );
  XNOR U18938 ( .A(n18173), .B(n18172), .Z(n18480) );
  XOR U18939 ( .A(n18175), .B(n18174), .Z(n18474) );
  AND U18940 ( .A(a[58]), .B(b[12]), .Z(n18473) );
  XOR U18941 ( .A(n18177), .B(n18176), .Z(n18468) );
  AND U18942 ( .A(a[56]), .B(b[12]), .Z(n18467) );
  AND U18943 ( .A(a[54]), .B(b[12]), .Z(n18461) );
  XOR U18944 ( .A(n18179), .B(n18178), .Z(n18180) );
  XNOR U18945 ( .A(n18181), .B(n18180), .Z(n18462) );
  AND U18946 ( .A(a[53]), .B(b[12]), .Z(n18455) );
  XOR U18947 ( .A(n18183), .B(n18182), .Z(n18773) );
  XOR U18948 ( .A(n18185), .B(n18184), .Z(n18765) );
  XOR U18949 ( .A(n18187), .B(n18186), .Z(n18755) );
  XNOR U18950 ( .A(n18189), .B(n18188), .Z(n18744) );
  AND U18951 ( .A(a[44]), .B(b[12]), .Z(n18419) );
  XNOR U18952 ( .A(n18191), .B(n18190), .Z(n18734) );
  XOR U18953 ( .A(n18193), .B(n18192), .Z(n18403) );
  IV U18954 ( .A(n18403), .Z(n18726) );
  NAND U18955 ( .A(a[40]), .B(b[12]), .Z(n18718) );
  XOR U18956 ( .A(n18195), .B(n18194), .Z(n18196) );
  XOR U18957 ( .A(n18197), .B(n18196), .Z(n18396) );
  IV U18958 ( .A(n18396), .Z(n18711) );
  NAND U18959 ( .A(a[38]), .B(b[12]), .Z(n18504) );
  XOR U18960 ( .A(n18199), .B(n18198), .Z(n18200) );
  XNOR U18961 ( .A(n18201), .B(n18200), .Z(n18703) );
  XNOR U18962 ( .A(n18203), .B(n18202), .Z(n18693) );
  XNOR U18963 ( .A(n18205), .B(n18204), .Z(n18685) );
  XNOR U18964 ( .A(n18207), .B(n18206), .Z(n18677) );
  XNOR U18965 ( .A(n18209), .B(n18208), .Z(n18669) );
  XNOR U18966 ( .A(n18211), .B(n18210), .Z(n18661) );
  XNOR U18967 ( .A(n18213), .B(n18212), .Z(n18653) );
  XNOR U18968 ( .A(n18215), .B(n18214), .Z(n18645) );
  AND U18969 ( .A(a[20]), .B(b[12]), .Z(n18321) );
  XNOR U18970 ( .A(n18217), .B(n18216), .Z(n18629) );
  NAND U18971 ( .A(a[18]), .B(b[12]), .Z(n18316) );
  XOR U18972 ( .A(n18219), .B(n18218), .Z(n18622) );
  AND U18973 ( .A(a[8]), .B(b[12]), .Z(n18261) );
  XOR U18974 ( .A(n18221), .B(n18220), .Z(n18243) );
  AND U18975 ( .A(a[1]), .B(b[13]), .Z(n18225) );
  AND U18976 ( .A(b[12]), .B(a[0]), .Z(n18866) );
  AND U18977 ( .A(n18225), .B(n18866), .Z(n18222) );
  NAND U18978 ( .A(a[2]), .B(n18222), .Z(n18229) );
  NAND U18979 ( .A(b[13]), .B(a[1]), .Z(n18223) );
  XOR U18980 ( .A(n18224), .B(n18223), .Z(n18539) );
  NAND U18981 ( .A(n18225), .B(a[0]), .Z(n18226) );
  XNOR U18982 ( .A(a[2]), .B(n18226), .Z(n18227) );
  AND U18983 ( .A(b[12]), .B(n18227), .Z(n18540) );
  NANDN U18984 ( .A(n18539), .B(n18540), .Z(n18228) );
  AND U18985 ( .A(n18229), .B(n18228), .Z(n18233) );
  XNOR U18986 ( .A(n18231), .B(n18230), .Z(n18232) );
  NANDN U18987 ( .A(n18233), .B(n18232), .Z(n18235) );
  XNOR U18988 ( .A(n18233), .B(n18232), .Z(n18546) );
  AND U18989 ( .A(a[3]), .B(b[12]), .Z(n18545) );
  NAND U18990 ( .A(n18546), .B(n18545), .Z(n18234) );
  AND U18991 ( .A(n18235), .B(n18234), .Z(n18237) );
  AND U18992 ( .A(a[4]), .B(b[12]), .Z(n18236) );
  NANDN U18993 ( .A(n18237), .B(n18236), .Z(n18241) );
  XNOR U18994 ( .A(n18237), .B(n18236), .Z(n18552) );
  XNOR U18995 ( .A(n18239), .B(n18238), .Z(n18551) );
  NAND U18996 ( .A(n18552), .B(n18551), .Z(n18240) );
  NAND U18997 ( .A(n18241), .B(n18240), .Z(n18242) );
  NAND U18998 ( .A(n18243), .B(n18242), .Z(n18245) );
  NAND U18999 ( .A(a[5]), .B(b[12]), .Z(n18557) );
  XOR U19000 ( .A(n18243), .B(n18242), .Z(n18558) );
  NANDN U19001 ( .A(n18557), .B(n18558), .Z(n18244) );
  AND U19002 ( .A(n18245), .B(n18244), .Z(n18249) );
  XNOR U19003 ( .A(n18247), .B(n18246), .Z(n18248) );
  NANDN U19004 ( .A(n18249), .B(n18248), .Z(n18251) );
  NAND U19005 ( .A(a[6]), .B(b[12]), .Z(n18563) );
  XNOR U19006 ( .A(n18249), .B(n18248), .Z(n18564) );
  NANDN U19007 ( .A(n18563), .B(n18564), .Z(n18250) );
  AND U19008 ( .A(n18251), .B(n18250), .Z(n18255) );
  XNOR U19009 ( .A(n18253), .B(n18252), .Z(n18254) );
  NANDN U19010 ( .A(n18255), .B(n18254), .Z(n18257) );
  NAND U19011 ( .A(a[7]), .B(b[12]), .Z(n18571) );
  XNOR U19012 ( .A(n18255), .B(n18254), .Z(n18572) );
  NANDN U19013 ( .A(n18571), .B(n18572), .Z(n18256) );
  AND U19014 ( .A(n18257), .B(n18256), .Z(n18260) );
  NANDN U19015 ( .A(n18261), .B(n18260), .Z(n18263) );
  XOR U19016 ( .A(n18259), .B(n18258), .Z(n18530) );
  XNOR U19017 ( .A(n18261), .B(n18260), .Z(n18529) );
  NANDN U19018 ( .A(n18530), .B(n18529), .Z(n18262) );
  AND U19019 ( .A(n18263), .B(n18262), .Z(n18267) );
  XOR U19020 ( .A(n18265), .B(n18264), .Z(n18266) );
  NAND U19021 ( .A(n18267), .B(n18266), .Z(n18269) );
  NAND U19022 ( .A(a[9]), .B(b[12]), .Z(n18579) );
  XOR U19023 ( .A(n18267), .B(n18266), .Z(n18580) );
  NANDN U19024 ( .A(n18579), .B(n18580), .Z(n18268) );
  AND U19025 ( .A(n18269), .B(n18268), .Z(n18271) );
  AND U19026 ( .A(a[10]), .B(b[12]), .Z(n18270) );
  NANDN U19027 ( .A(n18271), .B(n18270), .Z(n18275) );
  XNOR U19028 ( .A(n18271), .B(n18270), .Z(n18586) );
  XNOR U19029 ( .A(n18273), .B(n18272), .Z(n18585) );
  NAND U19030 ( .A(n18586), .B(n18585), .Z(n18274) );
  AND U19031 ( .A(n18275), .B(n18274), .Z(n18279) );
  XOR U19032 ( .A(n18277), .B(n18276), .Z(n18278) );
  NANDN U19033 ( .A(n18279), .B(n18278), .Z(n18281) );
  NAND U19034 ( .A(a[11]), .B(b[12]), .Z(n18591) );
  XNOR U19035 ( .A(n18279), .B(n18278), .Z(n18592) );
  NANDN U19036 ( .A(n18591), .B(n18592), .Z(n18280) );
  AND U19037 ( .A(n18281), .B(n18280), .Z(n18283) );
  AND U19038 ( .A(a[12]), .B(b[12]), .Z(n18282) );
  NANDN U19039 ( .A(n18283), .B(n18282), .Z(n18287) );
  XNOR U19040 ( .A(n18283), .B(n18282), .Z(n18598) );
  XNOR U19041 ( .A(n18285), .B(n18284), .Z(n18597) );
  NAND U19042 ( .A(n18598), .B(n18597), .Z(n18286) );
  AND U19043 ( .A(n18287), .B(n18286), .Z(n18291) );
  XOR U19044 ( .A(n18289), .B(n18288), .Z(n18290) );
  NANDN U19045 ( .A(n18291), .B(n18290), .Z(n18293) );
  NAND U19046 ( .A(a[13]), .B(b[12]), .Z(n18603) );
  XNOR U19047 ( .A(n18291), .B(n18290), .Z(n18604) );
  NANDN U19048 ( .A(n18603), .B(n18604), .Z(n18292) );
  AND U19049 ( .A(n18293), .B(n18292), .Z(n18295) );
  AND U19050 ( .A(a[14]), .B(b[12]), .Z(n18294) );
  NANDN U19051 ( .A(n18295), .B(n18294), .Z(n18299) );
  XNOR U19052 ( .A(n18295), .B(n18294), .Z(n18610) );
  XNOR U19053 ( .A(n18297), .B(n18296), .Z(n18609) );
  NAND U19054 ( .A(n18610), .B(n18609), .Z(n18298) );
  AND U19055 ( .A(n18299), .B(n18298), .Z(n18303) );
  XOR U19056 ( .A(n18301), .B(n18300), .Z(n18302) );
  NANDN U19057 ( .A(n18303), .B(n18302), .Z(n18305) );
  NAND U19058 ( .A(a[15]), .B(b[12]), .Z(n18615) );
  XNOR U19059 ( .A(n18303), .B(n18302), .Z(n18616) );
  NANDN U19060 ( .A(n18615), .B(n18616), .Z(n18304) );
  AND U19061 ( .A(n18305), .B(n18304), .Z(n18307) );
  AND U19062 ( .A(a[16]), .B(b[12]), .Z(n18306) );
  NANDN U19063 ( .A(n18307), .B(n18306), .Z(n18311) );
  XNOR U19064 ( .A(n18307), .B(n18306), .Z(n18528) );
  XNOR U19065 ( .A(n18309), .B(n18308), .Z(n18527) );
  NAND U19066 ( .A(n18528), .B(n18527), .Z(n18310) );
  AND U19067 ( .A(n18311), .B(n18310), .Z(n18621) );
  NAND U19068 ( .A(a[17]), .B(b[12]), .Z(n18624) );
  NANDN U19069 ( .A(n18316), .B(n18317), .Z(n18319) );
  XNOR U19070 ( .A(n18313), .B(n18312), .Z(n18314) );
  XNOR U19071 ( .A(n18315), .B(n18314), .Z(n18526) );
  XNOR U19072 ( .A(n18317), .B(n18316), .Z(n18525) );
  NAND U19073 ( .A(n18526), .B(n18525), .Z(n18318) );
  NAND U19074 ( .A(n18319), .B(n18318), .Z(n18630) );
  NAND U19075 ( .A(a[19]), .B(b[12]), .Z(n18632) );
  NANDN U19076 ( .A(n18321), .B(n18320), .Z(n18327) );
  XNOR U19077 ( .A(n18321), .B(n18320), .Z(n18523) );
  XNOR U19078 ( .A(n18323), .B(n18322), .Z(n18324) );
  XNOR U19079 ( .A(n18325), .B(n18324), .Z(n18524) );
  NAND U19080 ( .A(n18523), .B(n18524), .Z(n18326) );
  NAND U19081 ( .A(n18327), .B(n18326), .Z(n18638) );
  XOR U19082 ( .A(n18329), .B(n18328), .Z(n18637) );
  AND U19083 ( .A(a[21]), .B(b[12]), .Z(n18640) );
  AND U19084 ( .A(a[22]), .B(b[12]), .Z(n18334) );
  NANDN U19085 ( .A(n18335), .B(n18334), .Z(n18337) );
  XNOR U19086 ( .A(n18331), .B(n18330), .Z(n18332) );
  XNOR U19087 ( .A(n18333), .B(n18332), .Z(n18522) );
  XNOR U19088 ( .A(n18335), .B(n18334), .Z(n18521) );
  NAND U19089 ( .A(n18522), .B(n18521), .Z(n18336) );
  NAND U19090 ( .A(n18337), .B(n18336), .Z(n18646) );
  NAND U19091 ( .A(a[23]), .B(b[12]), .Z(n18648) );
  AND U19092 ( .A(a[24]), .B(b[12]), .Z(n18338) );
  NANDN U19093 ( .A(n18339), .B(n18338), .Z(n18345) );
  XOR U19094 ( .A(n18339), .B(n18338), .Z(n18519) );
  XNOR U19095 ( .A(n18341), .B(n18340), .Z(n18342) );
  XNOR U19096 ( .A(n18343), .B(n18342), .Z(n18520) );
  NANDN U19097 ( .A(n18519), .B(n18520), .Z(n18344) );
  NAND U19098 ( .A(n18345), .B(n18344), .Z(n18654) );
  NAND U19099 ( .A(a[25]), .B(b[12]), .Z(n18656) );
  AND U19100 ( .A(a[26]), .B(b[12]), .Z(n18350) );
  NANDN U19101 ( .A(n18351), .B(n18350), .Z(n18353) );
  XNOR U19102 ( .A(n18347), .B(n18346), .Z(n18348) );
  XNOR U19103 ( .A(n18349), .B(n18348), .Z(n18518) );
  XNOR U19104 ( .A(n18351), .B(n18350), .Z(n18517) );
  NAND U19105 ( .A(n18518), .B(n18517), .Z(n18352) );
  NAND U19106 ( .A(n18353), .B(n18352), .Z(n18662) );
  NAND U19107 ( .A(a[27]), .B(b[12]), .Z(n18664) );
  AND U19108 ( .A(a[28]), .B(b[12]), .Z(n18358) );
  NANDN U19109 ( .A(n18359), .B(n18358), .Z(n18361) );
  XNOR U19110 ( .A(n18355), .B(n18354), .Z(n18356) );
  XNOR U19111 ( .A(n18357), .B(n18356), .Z(n18516) );
  XNOR U19112 ( .A(n18359), .B(n18358), .Z(n18515) );
  NAND U19113 ( .A(n18516), .B(n18515), .Z(n18360) );
  NAND U19114 ( .A(n18361), .B(n18360), .Z(n18670) );
  NAND U19115 ( .A(a[29]), .B(b[12]), .Z(n18672) );
  AND U19116 ( .A(a[30]), .B(b[12]), .Z(n18366) );
  NANDN U19117 ( .A(n18367), .B(n18366), .Z(n18369) );
  XNOR U19118 ( .A(n18363), .B(n18362), .Z(n18364) );
  XNOR U19119 ( .A(n18365), .B(n18364), .Z(n18514) );
  XNOR U19120 ( .A(n18367), .B(n18366), .Z(n18513) );
  NAND U19121 ( .A(n18514), .B(n18513), .Z(n18368) );
  NAND U19122 ( .A(n18369), .B(n18368), .Z(n18678) );
  NAND U19123 ( .A(a[31]), .B(b[12]), .Z(n18680) );
  AND U19124 ( .A(a[32]), .B(b[12]), .Z(n18374) );
  NANDN U19125 ( .A(n18375), .B(n18374), .Z(n18377) );
  XNOR U19126 ( .A(n18371), .B(n18370), .Z(n18372) );
  XNOR U19127 ( .A(n18373), .B(n18372), .Z(n18512) );
  XNOR U19128 ( .A(n18375), .B(n18374), .Z(n18511) );
  NAND U19129 ( .A(n18512), .B(n18511), .Z(n18376) );
  NAND U19130 ( .A(n18377), .B(n18376), .Z(n18686) );
  NAND U19131 ( .A(a[33]), .B(b[12]), .Z(n18688) );
  AND U19132 ( .A(a[34]), .B(b[12]), .Z(n18382) );
  NANDN U19133 ( .A(n18383), .B(n18382), .Z(n18385) );
  XNOR U19134 ( .A(n18379), .B(n18378), .Z(n18380) );
  XNOR U19135 ( .A(n18381), .B(n18380), .Z(n18510) );
  XNOR U19136 ( .A(n18383), .B(n18382), .Z(n18509) );
  NAND U19137 ( .A(n18510), .B(n18509), .Z(n18384) );
  NAND U19138 ( .A(n18385), .B(n18384), .Z(n18694) );
  NAND U19139 ( .A(a[35]), .B(b[12]), .Z(n18696) );
  AND U19140 ( .A(a[36]), .B(b[12]), .Z(n18389) );
  NANDN U19141 ( .A(n18390), .B(n18389), .Z(n18392) );
  XNOR U19142 ( .A(n18390), .B(n18389), .Z(n18507) );
  NAND U19143 ( .A(n18508), .B(n18507), .Z(n18391) );
  NAND U19144 ( .A(n18392), .B(n18391), .Z(n18704) );
  NAND U19145 ( .A(a[37]), .B(b[12]), .Z(n18706) );
  NANDN U19146 ( .A(n18711), .B(n18710), .Z(n18399) );
  NOR U19147 ( .A(n18396), .B(n18710), .Z(n18397) );
  NAND U19148 ( .A(a[39]), .B(b[12]), .Z(n18713) );
  OR U19149 ( .A(n18397), .B(n18713), .Z(n18398) );
  AND U19150 ( .A(n18399), .B(n18398), .Z(n18717) );
  NANDN U19151 ( .A(n18726), .B(n18727), .Z(n18406) );
  NOR U19152 ( .A(n18403), .B(n18727), .Z(n18404) );
  AND U19153 ( .A(a[41]), .B(b[12]), .Z(n18725) );
  NANDN U19154 ( .A(n18404), .B(n18725), .Z(n18405) );
  AND U19155 ( .A(n18406), .B(n18405), .Z(n18407) );
  AND U19156 ( .A(a[42]), .B(b[12]), .Z(n18408) );
  NANDN U19157 ( .A(n18407), .B(n18408), .Z(n18414) );
  XNOR U19158 ( .A(n18408), .B(n18407), .Z(n18502) );
  XNOR U19159 ( .A(n18410), .B(n18409), .Z(n18411) );
  XNOR U19160 ( .A(n18412), .B(n18411), .Z(n18501) );
  NAND U19161 ( .A(n18502), .B(n18501), .Z(n18413) );
  NAND U19162 ( .A(n18414), .B(n18413), .Z(n18735) );
  NAND U19163 ( .A(a[43]), .B(b[12]), .Z(n18737) );
  NANDN U19164 ( .A(n18419), .B(n18420), .Z(n18422) );
  XOR U19165 ( .A(n18416), .B(n18415), .Z(n18417) );
  XNOR U19166 ( .A(n18418), .B(n18417), .Z(n18741) );
  NAND U19167 ( .A(n18741), .B(n18740), .Z(n18421) );
  AND U19168 ( .A(n18422), .B(n18421), .Z(n18743) );
  AND U19169 ( .A(a[45]), .B(b[12]), .Z(n18742) );
  AND U19170 ( .A(a[46]), .B(b[12]), .Z(n18423) );
  NANDN U19171 ( .A(n18424), .B(n18423), .Z(n18430) );
  XOR U19172 ( .A(n18424), .B(n18423), .Z(n18749) );
  XNOR U19173 ( .A(n18426), .B(n18425), .Z(n18427) );
  XNOR U19174 ( .A(n18428), .B(n18427), .Z(n18750) );
  NANDN U19175 ( .A(n18749), .B(n18750), .Z(n18429) );
  NAND U19176 ( .A(n18430), .B(n18429), .Z(n18431) );
  IV U19177 ( .A(n18431), .Z(n18752) );
  NAND U19178 ( .A(a[47]), .B(b[12]), .Z(n18753) );
  AND U19179 ( .A(a[48]), .B(b[12]), .Z(n18437) );
  NANDN U19180 ( .A(n18436), .B(n18437), .Z(n18439) );
  XNOR U19181 ( .A(n18433), .B(n18432), .Z(n18434) );
  XNOR U19182 ( .A(n18435), .B(n18434), .Z(n18500) );
  XNOR U19183 ( .A(n18437), .B(n18436), .Z(n18499) );
  NAND U19184 ( .A(n18500), .B(n18499), .Z(n18438) );
  NAND U19185 ( .A(n18439), .B(n18438), .Z(n18440) );
  IV U19186 ( .A(n18440), .Z(n18762) );
  NAND U19187 ( .A(a[49]), .B(b[12]), .Z(n18763) );
  AND U19188 ( .A(a[50]), .B(b[12]), .Z(n18445) );
  NANDN U19189 ( .A(n18444), .B(n18445), .Z(n18447) );
  XNOR U19190 ( .A(n18445), .B(n18444), .Z(n18498) );
  NANDN U19191 ( .A(n18497), .B(n18498), .Z(n18446) );
  NAND U19192 ( .A(n18447), .B(n18446), .Z(n18448) );
  IV U19193 ( .A(n18448), .Z(n18770) );
  NAND U19194 ( .A(a[51]), .B(b[12]), .Z(n18771) );
  AND U19195 ( .A(a[52]), .B(b[12]), .Z(n18451) );
  NANDN U19196 ( .A(n18452), .B(n18451), .Z(n18454) );
  XNOR U19197 ( .A(n18452), .B(n18451), .Z(n18496) );
  NANDN U19198 ( .A(n18495), .B(n18496), .Z(n18453) );
  NAND U19199 ( .A(n18454), .B(n18453), .Z(n18456) );
  XNOR U19200 ( .A(n18456), .B(n18455), .Z(n18493) );
  XOR U19201 ( .A(n18458), .B(n18457), .Z(n18459) );
  XNOR U19202 ( .A(n18460), .B(n18459), .Z(n18494) );
  XOR U19203 ( .A(n18462), .B(n18461), .Z(n18780) );
  XNOR U19204 ( .A(n18464), .B(n18463), .Z(n18465) );
  XOR U19205 ( .A(n18466), .B(n18465), .Z(n18783) );
  AND U19206 ( .A(a[55]), .B(b[12]), .Z(n18782) );
  XOR U19207 ( .A(n18468), .B(n18467), .Z(n18786) );
  XNOR U19208 ( .A(n18470), .B(n18469), .Z(n18471) );
  XOR U19209 ( .A(n18472), .B(n18471), .Z(n18789) );
  AND U19210 ( .A(a[57]), .B(b[12]), .Z(n18788) );
  XOR U19211 ( .A(n18474), .B(n18473), .Z(n18792) );
  XNOR U19212 ( .A(n18476), .B(n18475), .Z(n18477) );
  XOR U19213 ( .A(n18478), .B(n18477), .Z(n18797) );
  AND U19214 ( .A(a[59]), .B(b[12]), .Z(n18796) );
  XOR U19215 ( .A(n18480), .B(n18479), .Z(n18800) );
  XNOR U19216 ( .A(n18482), .B(n18481), .Z(n18483) );
  XOR U19217 ( .A(n18484), .B(n18483), .Z(n18805) );
  AND U19218 ( .A(a[61]), .B(b[12]), .Z(n18804) );
  AND U19219 ( .A(a[63]), .B(b[12]), .Z(n18814) );
  XOR U19220 ( .A(n18486), .B(n18485), .Z(n18815) );
  XOR U19221 ( .A(n18488), .B(n18487), .Z(n18492) );
  XOR U19222 ( .A(n18490), .B(n18489), .Z(n24716) );
  XOR U19223 ( .A(n18492), .B(n18491), .Z(n24705) );
  AND U19224 ( .A(a[62]), .B(b[11]), .Z(n18806) );
  NAND U19225 ( .A(a[61]), .B(b[11]), .Z(n18803) );
  AND U19226 ( .A(a[60]), .B(b[11]), .Z(n18798) );
  NAND U19227 ( .A(a[59]), .B(b[11]), .Z(n18795) );
  AND U19228 ( .A(a[58]), .B(b[11]), .Z(n18790) );
  AND U19229 ( .A(a[56]), .B(b[11]), .Z(n18784) );
  NAND U19230 ( .A(a[54]), .B(b[11]), .Z(n19132) );
  XOR U19231 ( .A(n18494), .B(n18493), .Z(n19135) );
  XNOR U19232 ( .A(n18500), .B(n18499), .Z(n19108) );
  NAND U19233 ( .A(a[48]), .B(b[11]), .Z(n18756) );
  NAND U19234 ( .A(a[46]), .B(b[11]), .Z(n18745) );
  XOR U19235 ( .A(n18502), .B(n18501), .Z(n18728) );
  IV U19236 ( .A(n18728), .Z(n19071) );
  NAND U19237 ( .A(a[42]), .B(b[11]), .Z(n18838) );
  AND U19238 ( .A(a[40]), .B(b[11]), .Z(n18709) );
  IV U19239 ( .A(n18709), .Z(n19054) );
  XOR U19240 ( .A(n18504), .B(n18503), .Z(n18505) );
  XOR U19241 ( .A(n18506), .B(n18505), .Z(n19047) );
  XNOR U19242 ( .A(n18508), .B(n18507), .Z(n19040) );
  XNOR U19243 ( .A(n18510), .B(n18509), .Z(n19030) );
  XNOR U19244 ( .A(n18512), .B(n18511), .Z(n19022) );
  XNOR U19245 ( .A(n18514), .B(n18513), .Z(n19014) );
  XNOR U19246 ( .A(n18516), .B(n18515), .Z(n19004) );
  XNOR U19247 ( .A(n18518), .B(n18517), .Z(n18996) );
  NAND U19248 ( .A(a[26]), .B(b[11]), .Z(n18657) );
  XNOR U19249 ( .A(n18520), .B(n18519), .Z(n18989) );
  XNOR U19250 ( .A(n18522), .B(n18521), .Z(n18980) );
  NAND U19251 ( .A(a[22]), .B(b[11]), .Z(n18641) );
  XNOR U19252 ( .A(n18524), .B(n18523), .Z(n18971) );
  XNOR U19253 ( .A(n18526), .B(n18525), .Z(n18962) );
  XNOR U19254 ( .A(n18528), .B(n18527), .Z(n18954) );
  XOR U19255 ( .A(n18530), .B(n18529), .Z(n18576) );
  AND U19256 ( .A(a[4]), .B(b[11]), .Z(n18548) );
  AND U19257 ( .A(a[0]), .B(b[11]), .Z(n19208) );
  AND U19258 ( .A(a[1]), .B(b[12]), .Z(n18534) );
  AND U19259 ( .A(n19208), .B(n18534), .Z(n18531) );
  NAND U19260 ( .A(a[2]), .B(n18531), .Z(n18538) );
  NAND U19261 ( .A(b[12]), .B(a[1]), .Z(n18532) );
  XOR U19262 ( .A(n18533), .B(n18532), .Z(n18872) );
  NAND U19263 ( .A(n18534), .B(a[0]), .Z(n18535) );
  XNOR U19264 ( .A(a[2]), .B(n18535), .Z(n18536) );
  AND U19265 ( .A(b[11]), .B(n18536), .Z(n18873) );
  NANDN U19266 ( .A(n18872), .B(n18873), .Z(n18537) );
  AND U19267 ( .A(n18538), .B(n18537), .Z(n18542) );
  XNOR U19268 ( .A(n18540), .B(n18539), .Z(n18541) );
  NANDN U19269 ( .A(n18542), .B(n18541), .Z(n18544) );
  NAND U19270 ( .A(a[3]), .B(b[11]), .Z(n18880) );
  XNOR U19271 ( .A(n18542), .B(n18541), .Z(n18881) );
  NANDN U19272 ( .A(n18880), .B(n18881), .Z(n18543) );
  AND U19273 ( .A(n18544), .B(n18543), .Z(n18547) );
  NANDN U19274 ( .A(n18548), .B(n18547), .Z(n18550) );
  XOR U19275 ( .A(n18546), .B(n18545), .Z(n18863) );
  XNOR U19276 ( .A(n18548), .B(n18547), .Z(n18862) );
  NANDN U19277 ( .A(n18863), .B(n18862), .Z(n18549) );
  AND U19278 ( .A(n18550), .B(n18549), .Z(n18554) );
  XOR U19279 ( .A(n18552), .B(n18551), .Z(n18553) );
  NAND U19280 ( .A(n18554), .B(n18553), .Z(n18556) );
  NAND U19281 ( .A(a[5]), .B(b[11]), .Z(n18888) );
  XOR U19282 ( .A(n18554), .B(n18553), .Z(n18889) );
  NANDN U19283 ( .A(n18888), .B(n18889), .Z(n18555) );
  AND U19284 ( .A(n18556), .B(n18555), .Z(n18560) );
  XNOR U19285 ( .A(n18558), .B(n18557), .Z(n18559) );
  NANDN U19286 ( .A(n18560), .B(n18559), .Z(n18562) );
  NAND U19287 ( .A(a[6]), .B(b[11]), .Z(n18894) );
  XNOR U19288 ( .A(n18560), .B(n18559), .Z(n18895) );
  NANDN U19289 ( .A(n18894), .B(n18895), .Z(n18561) );
  AND U19290 ( .A(n18562), .B(n18561), .Z(n18566) );
  XNOR U19291 ( .A(n18564), .B(n18563), .Z(n18565) );
  NANDN U19292 ( .A(n18566), .B(n18565), .Z(n18568) );
  XNOR U19293 ( .A(n18566), .B(n18565), .Z(n18901) );
  AND U19294 ( .A(a[7]), .B(b[11]), .Z(n18900) );
  NAND U19295 ( .A(n18901), .B(n18900), .Z(n18567) );
  AND U19296 ( .A(n18568), .B(n18567), .Z(n18570) );
  AND U19297 ( .A(a[8]), .B(b[11]), .Z(n18569) );
  NANDN U19298 ( .A(n18570), .B(n18569), .Z(n18574) );
  XNOR U19299 ( .A(n18570), .B(n18569), .Z(n18907) );
  XNOR U19300 ( .A(n18572), .B(n18571), .Z(n18906) );
  NAND U19301 ( .A(n18907), .B(n18906), .Z(n18573) );
  NAND U19302 ( .A(n18574), .B(n18573), .Z(n18575) );
  NAND U19303 ( .A(n18576), .B(n18575), .Z(n18578) );
  NAND U19304 ( .A(a[9]), .B(b[11]), .Z(n18914) );
  XOR U19305 ( .A(n18576), .B(n18575), .Z(n18915) );
  NANDN U19306 ( .A(n18914), .B(n18915), .Z(n18577) );
  AND U19307 ( .A(n18578), .B(n18577), .Z(n18582) );
  AND U19308 ( .A(a[10]), .B(b[11]), .Z(n18581) );
  NANDN U19309 ( .A(n18582), .B(n18581), .Z(n18584) );
  XNOR U19310 ( .A(n18580), .B(n18579), .Z(n18919) );
  XNOR U19311 ( .A(n18582), .B(n18581), .Z(n18918) );
  NAND U19312 ( .A(n18919), .B(n18918), .Z(n18583) );
  AND U19313 ( .A(n18584), .B(n18583), .Z(n18588) );
  XOR U19314 ( .A(n18586), .B(n18585), .Z(n18587) );
  NANDN U19315 ( .A(n18588), .B(n18587), .Z(n18590) );
  NAND U19316 ( .A(a[11]), .B(b[11]), .Z(n18926) );
  XNOR U19317 ( .A(n18588), .B(n18587), .Z(n18927) );
  NANDN U19318 ( .A(n18926), .B(n18927), .Z(n18589) );
  AND U19319 ( .A(n18590), .B(n18589), .Z(n18594) );
  AND U19320 ( .A(a[12]), .B(b[11]), .Z(n18593) );
  NANDN U19321 ( .A(n18594), .B(n18593), .Z(n18596) );
  XNOR U19322 ( .A(n18592), .B(n18591), .Z(n18931) );
  XNOR U19323 ( .A(n18594), .B(n18593), .Z(n18930) );
  NAND U19324 ( .A(n18931), .B(n18930), .Z(n18595) );
  AND U19325 ( .A(n18596), .B(n18595), .Z(n18600) );
  XOR U19326 ( .A(n18598), .B(n18597), .Z(n18599) );
  NANDN U19327 ( .A(n18600), .B(n18599), .Z(n18602) );
  NAND U19328 ( .A(a[13]), .B(b[11]), .Z(n18938) );
  XNOR U19329 ( .A(n18600), .B(n18599), .Z(n18939) );
  NANDN U19330 ( .A(n18938), .B(n18939), .Z(n18601) );
  AND U19331 ( .A(n18602), .B(n18601), .Z(n18606) );
  AND U19332 ( .A(a[14]), .B(b[11]), .Z(n18605) );
  NANDN U19333 ( .A(n18606), .B(n18605), .Z(n18608) );
  XNOR U19334 ( .A(n18604), .B(n18603), .Z(n18943) );
  XNOR U19335 ( .A(n18606), .B(n18605), .Z(n18942) );
  NAND U19336 ( .A(n18943), .B(n18942), .Z(n18607) );
  AND U19337 ( .A(n18608), .B(n18607), .Z(n18612) );
  XOR U19338 ( .A(n18610), .B(n18609), .Z(n18611) );
  NANDN U19339 ( .A(n18612), .B(n18611), .Z(n18614) );
  NAND U19340 ( .A(a[15]), .B(b[11]), .Z(n18950) );
  XNOR U19341 ( .A(n18612), .B(n18611), .Z(n18951) );
  NANDN U19342 ( .A(n18950), .B(n18951), .Z(n18613) );
  AND U19343 ( .A(n18614), .B(n18613), .Z(n18618) );
  AND U19344 ( .A(a[16]), .B(b[11]), .Z(n18617) );
  NANDN U19345 ( .A(n18618), .B(n18617), .Z(n18620) );
  XNOR U19346 ( .A(n18616), .B(n18615), .Z(n18861) );
  XNOR U19347 ( .A(n18618), .B(n18617), .Z(n18860) );
  NAND U19348 ( .A(n18861), .B(n18860), .Z(n18619) );
  NAND U19349 ( .A(n18620), .B(n18619), .Z(n18955) );
  NAND U19350 ( .A(a[17]), .B(b[11]), .Z(n18957) );
  AND U19351 ( .A(a[18]), .B(b[11]), .Z(n18625) );
  NANDN U19352 ( .A(n18626), .B(n18625), .Z(n18628) );
  XNOR U19353 ( .A(n18622), .B(n18621), .Z(n18623) );
  XNOR U19354 ( .A(n18624), .B(n18623), .Z(n18859) );
  XNOR U19355 ( .A(n18626), .B(n18625), .Z(n18858) );
  NAND U19356 ( .A(n18859), .B(n18858), .Z(n18627) );
  NAND U19357 ( .A(n18628), .B(n18627), .Z(n18963) );
  NAND U19358 ( .A(a[19]), .B(b[11]), .Z(n18965) );
  AND U19359 ( .A(a[20]), .B(b[11]), .Z(n18633) );
  NANDN U19360 ( .A(n18634), .B(n18633), .Z(n18636) );
  XNOR U19361 ( .A(n18630), .B(n18629), .Z(n18631) );
  XNOR U19362 ( .A(n18632), .B(n18631), .Z(n18857) );
  XNOR U19363 ( .A(n18634), .B(n18633), .Z(n18856) );
  NAND U19364 ( .A(n18857), .B(n18856), .Z(n18635) );
  AND U19365 ( .A(n18636), .B(n18635), .Z(n18970) );
  AND U19366 ( .A(a[21]), .B(b[11]), .Z(n18973) );
  NANDN U19367 ( .A(n18641), .B(n18642), .Z(n18644) );
  XOR U19368 ( .A(n18638), .B(n18637), .Z(n18639) );
  XNOR U19369 ( .A(n18640), .B(n18639), .Z(n18855) );
  XNOR U19370 ( .A(n18642), .B(n18641), .Z(n18854) );
  NAND U19371 ( .A(n18855), .B(n18854), .Z(n18643) );
  NAND U19372 ( .A(n18644), .B(n18643), .Z(n18981) );
  AND U19373 ( .A(a[23]), .B(b[11]), .Z(n18983) );
  AND U19374 ( .A(a[24]), .B(b[11]), .Z(n18649) );
  NANDN U19375 ( .A(n18650), .B(n18649), .Z(n18652) );
  XNOR U19376 ( .A(n18646), .B(n18645), .Z(n18647) );
  XNOR U19377 ( .A(n18648), .B(n18647), .Z(n18987) );
  XNOR U19378 ( .A(n18650), .B(n18649), .Z(n18986) );
  NAND U19379 ( .A(n18987), .B(n18986), .Z(n18651) );
  AND U19380 ( .A(n18652), .B(n18651), .Z(n18988) );
  AND U19381 ( .A(a[25]), .B(b[11]), .Z(n18991) );
  NANDN U19382 ( .A(n18657), .B(n18658), .Z(n18660) );
  XNOR U19383 ( .A(n18654), .B(n18653), .Z(n18655) );
  XNOR U19384 ( .A(n18656), .B(n18655), .Z(n18853) );
  XNOR U19385 ( .A(n18658), .B(n18657), .Z(n18852) );
  NAND U19386 ( .A(n18853), .B(n18852), .Z(n18659) );
  NAND U19387 ( .A(n18660), .B(n18659), .Z(n18997) );
  NAND U19388 ( .A(a[27]), .B(b[11]), .Z(n18999) );
  AND U19389 ( .A(a[28]), .B(b[11]), .Z(n18665) );
  NANDN U19390 ( .A(n18666), .B(n18665), .Z(n18668) );
  XNOR U19391 ( .A(n18662), .B(n18661), .Z(n18663) );
  XNOR U19392 ( .A(n18664), .B(n18663), .Z(n18851) );
  XNOR U19393 ( .A(n18666), .B(n18665), .Z(n18850) );
  NAND U19394 ( .A(n18851), .B(n18850), .Z(n18667) );
  NAND U19395 ( .A(n18668), .B(n18667), .Z(n19005) );
  NAND U19396 ( .A(a[29]), .B(b[11]), .Z(n19007) );
  AND U19397 ( .A(a[30]), .B(b[11]), .Z(n18673) );
  NANDN U19398 ( .A(n18674), .B(n18673), .Z(n18676) );
  XNOR U19399 ( .A(n18670), .B(n18669), .Z(n18671) );
  XNOR U19400 ( .A(n18672), .B(n18671), .Z(n18849) );
  XNOR U19401 ( .A(n18674), .B(n18673), .Z(n18848) );
  NAND U19402 ( .A(n18849), .B(n18848), .Z(n18675) );
  NAND U19403 ( .A(n18676), .B(n18675), .Z(n19015) );
  AND U19404 ( .A(a[31]), .B(b[11]), .Z(n19017) );
  AND U19405 ( .A(a[32]), .B(b[11]), .Z(n18681) );
  NANDN U19406 ( .A(n18682), .B(n18681), .Z(n18684) );
  XNOR U19407 ( .A(n18678), .B(n18677), .Z(n18679) );
  XNOR U19408 ( .A(n18680), .B(n18679), .Z(n19021) );
  XNOR U19409 ( .A(n18682), .B(n18681), .Z(n19020) );
  NAND U19410 ( .A(n19021), .B(n19020), .Z(n18683) );
  NAND U19411 ( .A(n18684), .B(n18683), .Z(n19023) );
  NAND U19412 ( .A(a[33]), .B(b[11]), .Z(n19025) );
  AND U19413 ( .A(a[34]), .B(b[11]), .Z(n18689) );
  NANDN U19414 ( .A(n18690), .B(n18689), .Z(n18692) );
  XNOR U19415 ( .A(n18686), .B(n18685), .Z(n18687) );
  XNOR U19416 ( .A(n18688), .B(n18687), .Z(n18847) );
  XNOR U19417 ( .A(n18690), .B(n18689), .Z(n18846) );
  NAND U19418 ( .A(n18847), .B(n18846), .Z(n18691) );
  NAND U19419 ( .A(n18692), .B(n18691), .Z(n19031) );
  NAND U19420 ( .A(a[35]), .B(b[11]), .Z(n19033) );
  AND U19421 ( .A(a[36]), .B(b[11]), .Z(n18697) );
  NANDN U19422 ( .A(n18698), .B(n18697), .Z(n18700) );
  XNOR U19423 ( .A(n18694), .B(n18693), .Z(n18695) );
  XNOR U19424 ( .A(n18696), .B(n18695), .Z(n18845) );
  XNOR U19425 ( .A(n18698), .B(n18697), .Z(n18844) );
  NAND U19426 ( .A(n18845), .B(n18844), .Z(n18699) );
  NAND U19427 ( .A(n18700), .B(n18699), .Z(n19041) );
  NAND U19428 ( .A(a[37]), .B(b[11]), .Z(n19043) );
  AND U19429 ( .A(a[38]), .B(b[11]), .Z(n18701) );
  NANDN U19430 ( .A(n18702), .B(n18701), .Z(n18708) );
  XNOR U19431 ( .A(n18702), .B(n18701), .Z(n18843) );
  XNOR U19432 ( .A(n18704), .B(n18703), .Z(n18705) );
  XNOR U19433 ( .A(n18706), .B(n18705), .Z(n18842) );
  NAND U19434 ( .A(n18843), .B(n18842), .Z(n18707) );
  AND U19435 ( .A(n18708), .B(n18707), .Z(n19046) );
  NAND U19436 ( .A(a[39]), .B(b[11]), .Z(n19049) );
  NANDN U19437 ( .A(n19054), .B(n19055), .Z(n18716) );
  NOR U19438 ( .A(n18709), .B(n19055), .Z(n18714) );
  XOR U19439 ( .A(n18711), .B(n18710), .Z(n18712) );
  XNOR U19440 ( .A(n18713), .B(n18712), .Z(n19057) );
  OR U19441 ( .A(n18714), .B(n19057), .Z(n18715) );
  AND U19442 ( .A(n18716), .B(n18715), .Z(n19063) );
  XOR U19443 ( .A(n18718), .B(n18717), .Z(n18719) );
  XOR U19444 ( .A(n18720), .B(n18719), .Z(n18721) );
  IV U19445 ( .A(n18721), .Z(n19062) );
  OR U19446 ( .A(n19063), .B(n19062), .Z(n18724) );
  ANDN U19447 ( .B(n19063), .A(n18721), .Z(n18722) );
  NAND U19448 ( .A(a[41]), .B(b[11]), .Z(n19065) );
  OR U19449 ( .A(n18722), .B(n19065), .Z(n18723) );
  AND U19450 ( .A(n18724), .B(n18723), .Z(n18839) );
  NANDN U19451 ( .A(n19071), .B(n19072), .Z(n18731) );
  NOR U19452 ( .A(n18728), .B(n19072), .Z(n18729) );
  NAND U19453 ( .A(a[43]), .B(b[11]), .Z(n19074) );
  OR U19454 ( .A(n18729), .B(n19074), .Z(n18730) );
  AND U19455 ( .A(n18731), .B(n18730), .Z(n18733) );
  AND U19456 ( .A(a[44]), .B(b[11]), .Z(n18732) );
  NANDN U19457 ( .A(n18733), .B(n18732), .Z(n18739) );
  XOR U19458 ( .A(n18733), .B(n18732), .Z(n18836) );
  XNOR U19459 ( .A(n18735), .B(n18734), .Z(n18736) );
  XNOR U19460 ( .A(n18737), .B(n18736), .Z(n18837) );
  NANDN U19461 ( .A(n18836), .B(n18837), .Z(n18738) );
  NAND U19462 ( .A(n18739), .B(n18738), .Z(n19085) );
  XOR U19463 ( .A(n18741), .B(n18740), .Z(n19084) );
  AND U19464 ( .A(a[45]), .B(b[11]), .Z(n19087) );
  NANDN U19465 ( .A(n18745), .B(n18746), .Z(n18748) );
  NAND U19466 ( .A(n19091), .B(n19090), .Z(n18747) );
  AND U19467 ( .A(n18748), .B(n18747), .Z(n19099) );
  IV U19468 ( .A(n18751), .Z(n19100) );
  NAND U19469 ( .A(a[47]), .B(b[11]), .Z(n19098) );
  NANDN U19470 ( .A(n18756), .B(n18757), .Z(n18759) );
  XOR U19471 ( .A(n18753), .B(n18752), .Z(n18754) );
  XOR U19472 ( .A(n18755), .B(n18754), .Z(n19104) );
  NAND U19473 ( .A(n19104), .B(n19103), .Z(n18758) );
  NAND U19474 ( .A(n18759), .B(n18758), .Z(n19109) );
  NAND U19475 ( .A(a[49]), .B(b[11]), .Z(n19111) );
  AND U19476 ( .A(a[50]), .B(b[11]), .Z(n18760) );
  NANDN U19477 ( .A(n18761), .B(n18760), .Z(n18767) );
  XNOR U19478 ( .A(n18761), .B(n18760), .Z(n18835) );
  XOR U19479 ( .A(n18763), .B(n18762), .Z(n18764) );
  XOR U19480 ( .A(n18765), .B(n18764), .Z(n18834) );
  NAND U19481 ( .A(n18835), .B(n18834), .Z(n18766) );
  NAND U19482 ( .A(n18767), .B(n18766), .Z(n19117) );
  NAND U19483 ( .A(a[51]), .B(b[11]), .Z(n19119) );
  AND U19484 ( .A(a[52]), .B(b[11]), .Z(n18768) );
  NANDN U19485 ( .A(n18769), .B(n18768), .Z(n18775) );
  XOR U19486 ( .A(n18769), .B(n18768), .Z(n19122) );
  XOR U19487 ( .A(n18771), .B(n18770), .Z(n18772) );
  XOR U19488 ( .A(n18773), .B(n18772), .Z(n19123) );
  NANDN U19489 ( .A(n19122), .B(n19123), .Z(n18774) );
  AND U19490 ( .A(n18775), .B(n18774), .Z(n18777) );
  NANDN U19491 ( .A(n18776), .B(n18777), .Z(n18779) );
  NAND U19492 ( .A(a[53]), .B(b[11]), .Z(n19124) );
  NAND U19493 ( .A(n19125), .B(n19124), .Z(n18778) );
  AND U19494 ( .A(n18779), .B(n18778), .Z(n19133) );
  NAND U19495 ( .A(a[55]), .B(b[11]), .Z(n18828) );
  XOR U19496 ( .A(n18781), .B(n18780), .Z(n18829) );
  XOR U19497 ( .A(n18783), .B(n18782), .Z(n19136) );
  XOR U19498 ( .A(n18785), .B(n18784), .Z(n19137) );
  NAND U19499 ( .A(a[57]), .B(b[11]), .Z(n18824) );
  XOR U19500 ( .A(n18787), .B(n18786), .Z(n18825) );
  XOR U19501 ( .A(n18789), .B(n18788), .Z(n19142) );
  XOR U19502 ( .A(n18791), .B(n18790), .Z(n19143) );
  XOR U19503 ( .A(n18793), .B(n18792), .Z(n18821) );
  XOR U19504 ( .A(n18795), .B(n18794), .Z(n18820) );
  XOR U19505 ( .A(n18797), .B(n18796), .Z(n19146) );
  XOR U19506 ( .A(n18799), .B(n18798), .Z(n19147) );
  XOR U19507 ( .A(n18801), .B(n18800), .Z(n18819) );
  XOR U19508 ( .A(n18803), .B(n18802), .Z(n18818) );
  XOR U19509 ( .A(n18805), .B(n18804), .Z(n19152) );
  XOR U19510 ( .A(n18807), .B(n18806), .Z(n19153) );
  NAND U19511 ( .A(a[63]), .B(b[11]), .Z(n18809) );
  XNOR U19512 ( .A(n18809), .B(n18808), .Z(n18816) );
  XOR U19513 ( .A(n18811), .B(n18810), .Z(n18812) );
  XOR U19514 ( .A(n18813), .B(n18812), .Z(n18817) );
  XOR U19515 ( .A(n18815), .B(n18814), .Z(n19156) );
  AND U19516 ( .A(n19157), .B(n19156), .Z(n24706) );
  NANDN U19517 ( .A(n24706), .B(n24705), .Z(n24713) );
  XOR U19518 ( .A(n18817), .B(n18816), .Z(n19480) );
  XOR U19519 ( .A(n18819), .B(n18818), .Z(n19151) );
  AND U19520 ( .A(a[62]), .B(b[10]), .Z(n19150) );
  AND U19521 ( .A(a[60]), .B(b[10]), .Z(n18822) );
  XOR U19522 ( .A(n18821), .B(n18820), .Z(n18823) );
  XNOR U19523 ( .A(n18823), .B(n18822), .Z(n19467) );
  AND U19524 ( .A(a[58]), .B(b[10]), .Z(n19140) );
  XOR U19525 ( .A(n18825), .B(n18824), .Z(n18826) );
  XOR U19526 ( .A(n18827), .B(n18826), .Z(n19141) );
  XOR U19527 ( .A(n18829), .B(n18828), .Z(n18830) );
  XNOR U19528 ( .A(n18831), .B(n18830), .Z(n18833) );
  AND U19529 ( .A(a[56]), .B(b[10]), .Z(n18832) );
  XOR U19530 ( .A(n18833), .B(n18832), .Z(n19451) );
  AND U19531 ( .A(a[55]), .B(b[10]), .Z(n19130) );
  XNOR U19532 ( .A(n18835), .B(n18834), .Z(n19431) );
  NAND U19533 ( .A(a[50]), .B(b[10]), .Z(n19106) );
  NAND U19534 ( .A(a[46]), .B(b[10]), .Z(n19082) );
  XOR U19535 ( .A(n18839), .B(n18838), .Z(n18840) );
  XOR U19536 ( .A(n18841), .B(n18840), .Z(n19066) );
  IV U19537 ( .A(n19066), .Z(n19403) );
  NAND U19538 ( .A(a[42]), .B(b[10]), .Z(n19176) );
  XNOR U19539 ( .A(n18843), .B(n18842), .Z(n19385) );
  XNOR U19540 ( .A(n18845), .B(n18844), .Z(n19375) );
  XNOR U19541 ( .A(n18847), .B(n18846), .Z(n19367) );
  AND U19542 ( .A(a[32]), .B(b[10]), .Z(n19013) );
  XNOR U19543 ( .A(n18849), .B(n18848), .Z(n19351) );
  XNOR U19544 ( .A(n18851), .B(n18850), .Z(n19343) );
  NAND U19545 ( .A(a[28]), .B(b[10]), .Z(n19000) );
  XOR U19546 ( .A(n18853), .B(n18852), .Z(n19336) );
  AND U19547 ( .A(a[26]), .B(b[10]), .Z(n18993) );
  AND U19548 ( .A(a[24]), .B(b[10]), .Z(n18979) );
  XNOR U19549 ( .A(n18855), .B(n18854), .Z(n19317) );
  XNOR U19550 ( .A(n18857), .B(n18856), .Z(n19309) );
  XNOR U19551 ( .A(n18859), .B(n18858), .Z(n19301) );
  XNOR U19552 ( .A(n18861), .B(n18860), .Z(n19293) );
  AND U19553 ( .A(a[8]), .B(b[10]), .Z(n18903) );
  XOR U19554 ( .A(n18863), .B(n18862), .Z(n18885) );
  AND U19555 ( .A(a[0]), .B(b[10]), .Z(n19542) );
  AND U19556 ( .A(a[1]), .B(b[11]), .Z(n18867) );
  AND U19557 ( .A(n19542), .B(n18867), .Z(n18864) );
  NAND U19558 ( .A(a[2]), .B(n18864), .Z(n18871) );
  NAND U19559 ( .A(b[11]), .B(a[1]), .Z(n18865) );
  XOR U19560 ( .A(n18866), .B(n18865), .Z(n19211) );
  NAND U19561 ( .A(n18867), .B(a[0]), .Z(n18868) );
  XNOR U19562 ( .A(a[2]), .B(n18868), .Z(n18869) );
  AND U19563 ( .A(b[10]), .B(n18869), .Z(n19212) );
  NANDN U19564 ( .A(n19211), .B(n19212), .Z(n18870) );
  AND U19565 ( .A(n18871), .B(n18870), .Z(n18875) );
  XNOR U19566 ( .A(n18873), .B(n18872), .Z(n18874) );
  NANDN U19567 ( .A(n18875), .B(n18874), .Z(n18877) );
  XNOR U19568 ( .A(n18875), .B(n18874), .Z(n19218) );
  AND U19569 ( .A(a[3]), .B(b[10]), .Z(n19217) );
  NAND U19570 ( .A(n19218), .B(n19217), .Z(n18876) );
  AND U19571 ( .A(n18877), .B(n18876), .Z(n18879) );
  AND U19572 ( .A(a[4]), .B(b[10]), .Z(n18878) );
  NANDN U19573 ( .A(n18879), .B(n18878), .Z(n18883) );
  XNOR U19574 ( .A(n18879), .B(n18878), .Z(n19224) );
  XNOR U19575 ( .A(n18881), .B(n18880), .Z(n19223) );
  NAND U19576 ( .A(n19224), .B(n19223), .Z(n18882) );
  NAND U19577 ( .A(n18883), .B(n18882), .Z(n18884) );
  NAND U19578 ( .A(n18885), .B(n18884), .Z(n18887) );
  NAND U19579 ( .A(a[5]), .B(b[10]), .Z(n19229) );
  XOR U19580 ( .A(n18885), .B(n18884), .Z(n19230) );
  NANDN U19581 ( .A(n19229), .B(n19230), .Z(n18886) );
  AND U19582 ( .A(n18887), .B(n18886), .Z(n18891) );
  XNOR U19583 ( .A(n18889), .B(n18888), .Z(n18890) );
  NANDN U19584 ( .A(n18891), .B(n18890), .Z(n18893) );
  NAND U19585 ( .A(a[6]), .B(b[10]), .Z(n19235) );
  XNOR U19586 ( .A(n18891), .B(n18890), .Z(n19236) );
  NANDN U19587 ( .A(n19235), .B(n19236), .Z(n18892) );
  AND U19588 ( .A(n18893), .B(n18892), .Z(n18897) );
  XNOR U19589 ( .A(n18895), .B(n18894), .Z(n18896) );
  NANDN U19590 ( .A(n18897), .B(n18896), .Z(n18899) );
  NAND U19591 ( .A(a[7]), .B(b[10]), .Z(n19243) );
  XNOR U19592 ( .A(n18897), .B(n18896), .Z(n19244) );
  NANDN U19593 ( .A(n19243), .B(n19244), .Z(n18898) );
  AND U19594 ( .A(n18899), .B(n18898), .Z(n18902) );
  NANDN U19595 ( .A(n18903), .B(n18902), .Z(n18905) );
  XOR U19596 ( .A(n18901), .B(n18900), .Z(n19202) );
  XNOR U19597 ( .A(n18903), .B(n18902), .Z(n19201) );
  NANDN U19598 ( .A(n19202), .B(n19201), .Z(n18904) );
  AND U19599 ( .A(n18905), .B(n18904), .Z(n18909) );
  XOR U19600 ( .A(n18907), .B(n18906), .Z(n18908) );
  NAND U19601 ( .A(n18909), .B(n18908), .Z(n18911) );
  NAND U19602 ( .A(a[9]), .B(b[10]), .Z(n19251) );
  XOR U19603 ( .A(n18909), .B(n18908), .Z(n19252) );
  NANDN U19604 ( .A(n19251), .B(n19252), .Z(n18910) );
  AND U19605 ( .A(n18911), .B(n18910), .Z(n18913) );
  AND U19606 ( .A(a[10]), .B(b[10]), .Z(n18912) );
  NANDN U19607 ( .A(n18913), .B(n18912), .Z(n18917) );
  XNOR U19608 ( .A(n18913), .B(n18912), .Z(n19258) );
  XNOR U19609 ( .A(n18915), .B(n18914), .Z(n19257) );
  NAND U19610 ( .A(n19258), .B(n19257), .Z(n18916) );
  AND U19611 ( .A(n18917), .B(n18916), .Z(n18921) );
  XOR U19612 ( .A(n18919), .B(n18918), .Z(n18920) );
  NANDN U19613 ( .A(n18921), .B(n18920), .Z(n18923) );
  NAND U19614 ( .A(a[11]), .B(b[10]), .Z(n19263) );
  XNOR U19615 ( .A(n18921), .B(n18920), .Z(n19264) );
  NANDN U19616 ( .A(n19263), .B(n19264), .Z(n18922) );
  AND U19617 ( .A(n18923), .B(n18922), .Z(n18925) );
  AND U19618 ( .A(a[12]), .B(b[10]), .Z(n18924) );
  NANDN U19619 ( .A(n18925), .B(n18924), .Z(n18929) );
  XNOR U19620 ( .A(n18925), .B(n18924), .Z(n19270) );
  XNOR U19621 ( .A(n18927), .B(n18926), .Z(n19269) );
  NAND U19622 ( .A(n19270), .B(n19269), .Z(n18928) );
  AND U19623 ( .A(n18929), .B(n18928), .Z(n18933) );
  XOR U19624 ( .A(n18931), .B(n18930), .Z(n18932) );
  NANDN U19625 ( .A(n18933), .B(n18932), .Z(n18935) );
  NAND U19626 ( .A(a[13]), .B(b[10]), .Z(n19275) );
  XNOR U19627 ( .A(n18933), .B(n18932), .Z(n19276) );
  NANDN U19628 ( .A(n19275), .B(n19276), .Z(n18934) );
  AND U19629 ( .A(n18935), .B(n18934), .Z(n18937) );
  AND U19630 ( .A(a[14]), .B(b[10]), .Z(n18936) );
  NANDN U19631 ( .A(n18937), .B(n18936), .Z(n18941) );
  XNOR U19632 ( .A(n18937), .B(n18936), .Z(n19282) );
  XNOR U19633 ( .A(n18939), .B(n18938), .Z(n19281) );
  NAND U19634 ( .A(n19282), .B(n19281), .Z(n18940) );
  AND U19635 ( .A(n18941), .B(n18940), .Z(n18945) );
  XOR U19636 ( .A(n18943), .B(n18942), .Z(n18944) );
  NANDN U19637 ( .A(n18945), .B(n18944), .Z(n18947) );
  NAND U19638 ( .A(a[15]), .B(b[10]), .Z(n19287) );
  XNOR U19639 ( .A(n18945), .B(n18944), .Z(n19288) );
  NANDN U19640 ( .A(n19287), .B(n19288), .Z(n18946) );
  AND U19641 ( .A(n18947), .B(n18946), .Z(n18949) );
  AND U19642 ( .A(a[16]), .B(b[10]), .Z(n18948) );
  NANDN U19643 ( .A(n18949), .B(n18948), .Z(n18953) );
  XNOR U19644 ( .A(n18949), .B(n18948), .Z(n19200) );
  XNOR U19645 ( .A(n18951), .B(n18950), .Z(n19199) );
  NAND U19646 ( .A(n19200), .B(n19199), .Z(n18952) );
  NAND U19647 ( .A(n18953), .B(n18952), .Z(n19294) );
  NAND U19648 ( .A(a[17]), .B(b[10]), .Z(n19296) );
  AND U19649 ( .A(a[18]), .B(b[10]), .Z(n18958) );
  NANDN U19650 ( .A(n18959), .B(n18958), .Z(n18961) );
  XNOR U19651 ( .A(n18955), .B(n18954), .Z(n18956) );
  XNOR U19652 ( .A(n18957), .B(n18956), .Z(n19198) );
  XNOR U19653 ( .A(n18959), .B(n18958), .Z(n19197) );
  NAND U19654 ( .A(n19198), .B(n19197), .Z(n18960) );
  NAND U19655 ( .A(n18961), .B(n18960), .Z(n19302) );
  NAND U19656 ( .A(a[19]), .B(b[10]), .Z(n19304) );
  AND U19657 ( .A(a[20]), .B(b[10]), .Z(n18966) );
  NANDN U19658 ( .A(n18967), .B(n18966), .Z(n18969) );
  XNOR U19659 ( .A(n18963), .B(n18962), .Z(n18964) );
  XNOR U19660 ( .A(n18965), .B(n18964), .Z(n19196) );
  XNOR U19661 ( .A(n18967), .B(n18966), .Z(n19195) );
  NAND U19662 ( .A(n19196), .B(n19195), .Z(n18968) );
  NAND U19663 ( .A(n18969), .B(n18968), .Z(n19310) );
  NAND U19664 ( .A(a[21]), .B(b[10]), .Z(n19312) );
  AND U19665 ( .A(a[22]), .B(b[10]), .Z(n18974) );
  NANDN U19666 ( .A(n18975), .B(n18974), .Z(n18977) );
  XOR U19667 ( .A(n18971), .B(n18970), .Z(n18972) );
  XNOR U19668 ( .A(n18973), .B(n18972), .Z(n19194) );
  XNOR U19669 ( .A(n18975), .B(n18974), .Z(n19193) );
  NAND U19670 ( .A(n19194), .B(n19193), .Z(n18976) );
  NAND U19671 ( .A(n18977), .B(n18976), .Z(n19318) );
  NAND U19672 ( .A(a[23]), .B(b[10]), .Z(n19320) );
  NANDN U19673 ( .A(n18979), .B(n18978), .Z(n18985) );
  XNOR U19674 ( .A(n18979), .B(n18978), .Z(n19191) );
  XNOR U19675 ( .A(n18981), .B(n18980), .Z(n18982) );
  XNOR U19676 ( .A(n18983), .B(n18982), .Z(n19192) );
  NAND U19677 ( .A(n19191), .B(n19192), .Z(n18984) );
  NAND U19678 ( .A(n18985), .B(n18984), .Z(n19328) );
  XOR U19679 ( .A(n18987), .B(n18986), .Z(n19327) );
  AND U19680 ( .A(a[25]), .B(b[10]), .Z(n19330) );
  NANDN U19681 ( .A(n18993), .B(n18992), .Z(n18995) );
  XNOR U19682 ( .A(n18989), .B(n18988), .Z(n18990) );
  XNOR U19683 ( .A(n18991), .B(n18990), .Z(n19334) );
  XNOR U19684 ( .A(n18993), .B(n18992), .Z(n19333) );
  NAND U19685 ( .A(n19334), .B(n19333), .Z(n18994) );
  NAND U19686 ( .A(n18995), .B(n18994), .Z(n19335) );
  AND U19687 ( .A(a[27]), .B(b[10]), .Z(n19338) );
  NANDN U19688 ( .A(n19000), .B(n19001), .Z(n19003) );
  XNOR U19689 ( .A(n18997), .B(n18996), .Z(n18998) );
  XNOR U19690 ( .A(n18999), .B(n18998), .Z(n19190) );
  XNOR U19691 ( .A(n19001), .B(n19000), .Z(n19189) );
  NAND U19692 ( .A(n19190), .B(n19189), .Z(n19002) );
  NAND U19693 ( .A(n19003), .B(n19002), .Z(n19344) );
  NAND U19694 ( .A(a[29]), .B(b[10]), .Z(n19346) );
  AND U19695 ( .A(a[30]), .B(b[10]), .Z(n19008) );
  NANDN U19696 ( .A(n19009), .B(n19008), .Z(n19011) );
  XNOR U19697 ( .A(n19005), .B(n19004), .Z(n19006) );
  XNOR U19698 ( .A(n19007), .B(n19006), .Z(n19188) );
  XNOR U19699 ( .A(n19009), .B(n19008), .Z(n19187) );
  NAND U19700 ( .A(n19188), .B(n19187), .Z(n19010) );
  NAND U19701 ( .A(n19011), .B(n19010), .Z(n19352) );
  NAND U19702 ( .A(a[31]), .B(b[10]), .Z(n19354) );
  NANDN U19703 ( .A(n19013), .B(n19012), .Z(n19019) );
  XNOR U19704 ( .A(n19013), .B(n19012), .Z(n19185) );
  XNOR U19705 ( .A(n19015), .B(n19014), .Z(n19016) );
  XNOR U19706 ( .A(n19017), .B(n19016), .Z(n19186) );
  NAND U19707 ( .A(n19185), .B(n19186), .Z(n19018) );
  NAND U19708 ( .A(n19019), .B(n19018), .Z(n19360) );
  XOR U19709 ( .A(n19021), .B(n19020), .Z(n19359) );
  AND U19710 ( .A(a[33]), .B(b[10]), .Z(n19362) );
  AND U19711 ( .A(a[34]), .B(b[10]), .Z(n19026) );
  NANDN U19712 ( .A(n19027), .B(n19026), .Z(n19029) );
  XNOR U19713 ( .A(n19023), .B(n19022), .Z(n19024) );
  XNOR U19714 ( .A(n19025), .B(n19024), .Z(n19184) );
  XNOR U19715 ( .A(n19027), .B(n19026), .Z(n19183) );
  NAND U19716 ( .A(n19184), .B(n19183), .Z(n19028) );
  NAND U19717 ( .A(n19029), .B(n19028), .Z(n19368) );
  NAND U19718 ( .A(a[35]), .B(b[10]), .Z(n19370) );
  AND U19719 ( .A(a[36]), .B(b[10]), .Z(n19034) );
  NANDN U19720 ( .A(n19035), .B(n19034), .Z(n19037) );
  XNOR U19721 ( .A(n19031), .B(n19030), .Z(n19032) );
  XNOR U19722 ( .A(n19033), .B(n19032), .Z(n19182) );
  XNOR U19723 ( .A(n19035), .B(n19034), .Z(n19181) );
  NAND U19724 ( .A(n19182), .B(n19181), .Z(n19036) );
  NAND U19725 ( .A(n19037), .B(n19036), .Z(n19376) );
  NAND U19726 ( .A(a[37]), .B(b[10]), .Z(n19378) );
  AND U19727 ( .A(a[38]), .B(b[10]), .Z(n19038) );
  NANDN U19728 ( .A(n19039), .B(n19038), .Z(n19045) );
  XOR U19729 ( .A(n19039), .B(n19038), .Z(n19383) );
  XNOR U19730 ( .A(n19041), .B(n19040), .Z(n19042) );
  XNOR U19731 ( .A(n19043), .B(n19042), .Z(n19384) );
  NANDN U19732 ( .A(n19383), .B(n19384), .Z(n19044) );
  NAND U19733 ( .A(n19045), .B(n19044), .Z(n19386) );
  NAND U19734 ( .A(a[39]), .B(b[10]), .Z(n19388) );
  AND U19735 ( .A(a[40]), .B(b[10]), .Z(n19050) );
  NANDN U19736 ( .A(n19051), .B(n19050), .Z(n19053) );
  XNOR U19737 ( .A(n19047), .B(n19046), .Z(n19048) );
  XNOR U19738 ( .A(n19049), .B(n19048), .Z(n19180) );
  XNOR U19739 ( .A(n19051), .B(n19050), .Z(n19179) );
  NAND U19740 ( .A(n19180), .B(n19179), .Z(n19052) );
  AND U19741 ( .A(n19053), .B(n19052), .Z(n19395) );
  XOR U19742 ( .A(n19055), .B(n19054), .Z(n19056) );
  XOR U19743 ( .A(n19057), .B(n19056), .Z(n19058) );
  IV U19744 ( .A(n19058), .Z(n19396) );
  OR U19745 ( .A(n19395), .B(n19396), .Z(n19061) );
  ANDN U19746 ( .B(n19395), .A(n19058), .Z(n19059) );
  NAND U19747 ( .A(a[41]), .B(b[10]), .Z(n19398) );
  OR U19748 ( .A(n19059), .B(n19398), .Z(n19060) );
  AND U19749 ( .A(n19061), .B(n19060), .Z(n19175) );
  XOR U19750 ( .A(n19063), .B(n19062), .Z(n19064) );
  XOR U19751 ( .A(n19065), .B(n19064), .Z(n19178) );
  NANDN U19752 ( .A(n19403), .B(n19402), .Z(n19069) );
  NOR U19753 ( .A(n19066), .B(n19402), .Z(n19067) );
  AND U19754 ( .A(a[43]), .B(b[10]), .Z(n19405) );
  NANDN U19755 ( .A(n19067), .B(n19405), .Z(n19068) );
  AND U19756 ( .A(n19069), .B(n19068), .Z(n19173) );
  AND U19757 ( .A(a[44]), .B(b[10]), .Z(n19070) );
  IV U19758 ( .A(n19070), .Z(n19174) );
  OR U19759 ( .A(n19173), .B(n19174), .Z(n19077) );
  ANDN U19760 ( .B(n19173), .A(n19070), .Z(n19075) );
  XOR U19761 ( .A(n19072), .B(n19071), .Z(n19073) );
  XOR U19762 ( .A(n19074), .B(n19073), .Z(n19172) );
  NANDN U19763 ( .A(n19075), .B(n19172), .Z(n19076) );
  AND U19764 ( .A(n19077), .B(n19076), .Z(n19410) );
  NANDN U19765 ( .A(n19078), .B(n19410), .Z(n19081) );
  IV U19766 ( .A(n19078), .Z(n19411) );
  NOR U19767 ( .A(n19411), .B(n19410), .Z(n19079) );
  NAND U19768 ( .A(a[45]), .B(b[10]), .Z(n19409) );
  NANDN U19769 ( .A(n19079), .B(n19409), .Z(n19080) );
  AND U19770 ( .A(n19081), .B(n19080), .Z(n19083) );
  NANDN U19771 ( .A(n19082), .B(n19083), .Z(n19089) );
  XOR U19772 ( .A(n19085), .B(n19084), .Z(n19086) );
  XNOR U19773 ( .A(n19087), .B(n19086), .Z(n19170) );
  NAND U19774 ( .A(n19171), .B(n19170), .Z(n19088) );
  AND U19775 ( .A(n19089), .B(n19088), .Z(n19416) );
  XOR U19776 ( .A(n19091), .B(n19090), .Z(n19092) );
  IV U19777 ( .A(n19092), .Z(n19417) );
  OR U19778 ( .A(n19416), .B(n19417), .Z(n19095) );
  ANDN U19779 ( .B(n19416), .A(n19092), .Z(n19093) );
  NAND U19780 ( .A(a[47]), .B(b[10]), .Z(n19419) );
  OR U19781 ( .A(n19093), .B(n19419), .Z(n19094) );
  AND U19782 ( .A(n19095), .B(n19094), .Z(n19096) );
  AND U19783 ( .A(a[48]), .B(b[10]), .Z(n19097) );
  NANDN U19784 ( .A(n19096), .B(n19097), .Z(n19102) );
  XNOR U19785 ( .A(n19097), .B(n19096), .Z(n19169) );
  NAND U19786 ( .A(n19169), .B(n19168), .Z(n19101) );
  AND U19787 ( .A(n19102), .B(n19101), .Z(n19425) );
  XOR U19788 ( .A(n19104), .B(n19103), .Z(n19105) );
  IV U19789 ( .A(n19105), .Z(n19426) );
  NAND U19790 ( .A(a[49]), .B(b[10]), .Z(n19424) );
  NANDN U19791 ( .A(n19106), .B(n19107), .Z(n19113) );
  XNOR U19792 ( .A(n19109), .B(n19108), .Z(n19110) );
  XNOR U19793 ( .A(n19111), .B(n19110), .Z(n19166) );
  NAND U19794 ( .A(n19167), .B(n19166), .Z(n19112) );
  NAND U19795 ( .A(n19113), .B(n19112), .Z(n19432) );
  NAND U19796 ( .A(a[51]), .B(b[10]), .Z(n19434) );
  NAND U19797 ( .A(a[52]), .B(b[10]), .Z(n19115) );
  NAND U19798 ( .A(n19114), .B(n19115), .Z(n19121) );
  XOR U19799 ( .A(n19115), .B(n19114), .Z(n19164) );
  XNOR U19800 ( .A(n19117), .B(n19116), .Z(n19118) );
  XOR U19801 ( .A(n19119), .B(n19118), .Z(n19165) );
  NAND U19802 ( .A(n19164), .B(n19165), .Z(n19120) );
  NAND U19803 ( .A(n19121), .B(n19120), .Z(n19442) );
  NAND U19804 ( .A(a[53]), .B(b[10]), .Z(n19444) );
  AND U19805 ( .A(a[54]), .B(b[10]), .Z(n19126) );
  NANDN U19806 ( .A(n19127), .B(n19126), .Z(n19129) );
  XOR U19807 ( .A(n19125), .B(n19124), .Z(n19162) );
  XNOR U19808 ( .A(n19127), .B(n19126), .Z(n19163) );
  NANDN U19809 ( .A(n19162), .B(n19163), .Z(n19128) );
  NAND U19810 ( .A(n19129), .B(n19128), .Z(n19131) );
  XNOR U19811 ( .A(n19131), .B(n19130), .Z(n19160) );
  XOR U19812 ( .A(n19133), .B(n19132), .Z(n19134) );
  XOR U19813 ( .A(n19135), .B(n19134), .Z(n19161) );
  XOR U19814 ( .A(n19137), .B(n19136), .Z(n19138) );
  XOR U19815 ( .A(n19139), .B(n19138), .Z(n19456) );
  AND U19816 ( .A(a[57]), .B(b[10]), .Z(n19455) );
  XOR U19817 ( .A(n19141), .B(n19140), .Z(n19459) );
  XOR U19818 ( .A(n19143), .B(n19142), .Z(n19144) );
  XOR U19819 ( .A(n19145), .B(n19144), .Z(n19464) );
  AND U19820 ( .A(a[59]), .B(b[10]), .Z(n19463) );
  XOR U19821 ( .A(n19147), .B(n19146), .Z(n19148) );
  XOR U19822 ( .A(n19149), .B(n19148), .Z(n19472) );
  AND U19823 ( .A(a[61]), .B(b[10]), .Z(n19471) );
  XOR U19824 ( .A(n19151), .B(n19150), .Z(n19475) );
  XOR U19825 ( .A(n19153), .B(n19152), .Z(n19154) );
  XOR U19826 ( .A(n19155), .B(n19154), .Z(n19159) );
  AND U19827 ( .A(a[63]), .B(b[10]), .Z(n19158) );
  XOR U19828 ( .A(n19157), .B(n19156), .Z(n24701) );
  IV U19829 ( .A(n24701), .Z(n19481) );
  NANDN U19830 ( .A(n24702), .B(n19481), .Z(n24710) );
  XOR U19831 ( .A(n19159), .B(n19158), .Z(n20149) );
  NAND U19832 ( .A(a[63]), .B(b[9]), .Z(n19478) );
  AND U19833 ( .A(a[60]), .B(b[9]), .Z(n19465) );
  NAND U19834 ( .A(a[59]), .B(b[9]), .Z(n19462) );
  AND U19835 ( .A(a[57]), .B(b[9]), .Z(n19453) );
  AND U19836 ( .A(a[56]), .B(b[9]), .Z(n19802) );
  XOR U19837 ( .A(n19161), .B(n19160), .Z(n19801) );
  XNOR U19838 ( .A(n19165), .B(n19164), .Z(n19786) );
  XNOR U19839 ( .A(n19167), .B(n19166), .Z(n19775) );
  XNOR U19840 ( .A(n19169), .B(n19168), .Z(n19767) );
  XOR U19841 ( .A(n19171), .B(n19170), .Z(n19412) );
  IV U19842 ( .A(n19412), .Z(n19761) );
  NAND U19843 ( .A(a[46]), .B(b[9]), .Z(n19752) );
  AND U19844 ( .A(a[44]), .B(b[9]), .Z(n19508) );
  XOR U19845 ( .A(n19176), .B(n19175), .Z(n19177) );
  XOR U19846 ( .A(n19178), .B(n19177), .Z(n19736) );
  XNOR U19847 ( .A(n19180), .B(n19179), .Z(n19730) );
  XNOR U19848 ( .A(n19182), .B(n19181), .Z(n19712) );
  XNOR U19849 ( .A(n19184), .B(n19183), .Z(n19704) );
  XOR U19850 ( .A(n19186), .B(n19185), .Z(n19697) );
  XNOR U19851 ( .A(n19188), .B(n19187), .Z(n19688) );
  XNOR U19852 ( .A(n19190), .B(n19189), .Z(n19680) );
  NAND U19853 ( .A(a[28]), .B(b[9]), .Z(n19339) );
  XOR U19854 ( .A(n19192), .B(n19191), .Z(n19662) );
  XNOR U19855 ( .A(n19194), .B(n19193), .Z(n19654) );
  XNOR U19856 ( .A(n19196), .B(n19195), .Z(n19648) );
  XNOR U19857 ( .A(n19198), .B(n19197), .Z(n19638) );
  XNOR U19858 ( .A(n19200), .B(n19199), .Z(n19632) );
  XOR U19859 ( .A(n19202), .B(n19201), .Z(n19248) );
  AND U19860 ( .A(a[4]), .B(b[9]), .Z(n19220) );
  AND U19861 ( .A(a[0]), .B(b[9]), .Z(n19875) );
  AND U19862 ( .A(a[1]), .B(b[10]), .Z(n19204) );
  AND U19863 ( .A(n19875), .B(n19204), .Z(n19203) );
  NAND U19864 ( .A(a[2]), .B(n19203), .Z(n19210) );
  NAND U19865 ( .A(n19204), .B(a[0]), .Z(n19205) );
  XNOR U19866 ( .A(a[2]), .B(n19205), .Z(n19206) );
  NAND U19867 ( .A(b[9]), .B(n19206), .Z(n19548) );
  NAND U19868 ( .A(b[10]), .B(a[1]), .Z(n19207) );
  XNOR U19869 ( .A(n19208), .B(n19207), .Z(n19549) );
  NANDN U19870 ( .A(n19548), .B(n19549), .Z(n19209) );
  AND U19871 ( .A(n19210), .B(n19209), .Z(n19214) );
  XNOR U19872 ( .A(n19212), .B(n19211), .Z(n19213) );
  NANDN U19873 ( .A(n19214), .B(n19213), .Z(n19216) );
  NAND U19874 ( .A(a[3]), .B(b[9]), .Z(n19556) );
  XNOR U19875 ( .A(n19214), .B(n19213), .Z(n19557) );
  NANDN U19876 ( .A(n19556), .B(n19557), .Z(n19215) );
  AND U19877 ( .A(n19216), .B(n19215), .Z(n19219) );
  NANDN U19878 ( .A(n19220), .B(n19219), .Z(n19222) );
  XOR U19879 ( .A(n19218), .B(n19217), .Z(n19539) );
  XNOR U19880 ( .A(n19220), .B(n19219), .Z(n19538) );
  NANDN U19881 ( .A(n19539), .B(n19538), .Z(n19221) );
  AND U19882 ( .A(n19222), .B(n19221), .Z(n19226) );
  XOR U19883 ( .A(n19224), .B(n19223), .Z(n19225) );
  NAND U19884 ( .A(n19226), .B(n19225), .Z(n19228) );
  NAND U19885 ( .A(a[5]), .B(b[9]), .Z(n19564) );
  XOR U19886 ( .A(n19226), .B(n19225), .Z(n19565) );
  NANDN U19887 ( .A(n19564), .B(n19565), .Z(n19227) );
  AND U19888 ( .A(n19228), .B(n19227), .Z(n19232) );
  XNOR U19889 ( .A(n19230), .B(n19229), .Z(n19231) );
  NANDN U19890 ( .A(n19232), .B(n19231), .Z(n19234) );
  NAND U19891 ( .A(a[6]), .B(b[9]), .Z(n19570) );
  XNOR U19892 ( .A(n19232), .B(n19231), .Z(n19571) );
  NANDN U19893 ( .A(n19570), .B(n19571), .Z(n19233) );
  AND U19894 ( .A(n19234), .B(n19233), .Z(n19238) );
  XNOR U19895 ( .A(n19236), .B(n19235), .Z(n19237) );
  NANDN U19896 ( .A(n19238), .B(n19237), .Z(n19240) );
  XNOR U19897 ( .A(n19238), .B(n19237), .Z(n19577) );
  AND U19898 ( .A(a[7]), .B(b[9]), .Z(n19576) );
  NAND U19899 ( .A(n19577), .B(n19576), .Z(n19239) );
  AND U19900 ( .A(n19240), .B(n19239), .Z(n19242) );
  AND U19901 ( .A(a[8]), .B(b[9]), .Z(n19241) );
  NANDN U19902 ( .A(n19242), .B(n19241), .Z(n19246) );
  XNOR U19903 ( .A(n19242), .B(n19241), .Z(n19583) );
  XNOR U19904 ( .A(n19244), .B(n19243), .Z(n19582) );
  NAND U19905 ( .A(n19583), .B(n19582), .Z(n19245) );
  NAND U19906 ( .A(n19246), .B(n19245), .Z(n19247) );
  NAND U19907 ( .A(n19248), .B(n19247), .Z(n19250) );
  NAND U19908 ( .A(a[9]), .B(b[9]), .Z(n19590) );
  XOR U19909 ( .A(n19248), .B(n19247), .Z(n19591) );
  NANDN U19910 ( .A(n19590), .B(n19591), .Z(n19249) );
  AND U19911 ( .A(n19250), .B(n19249), .Z(n19254) );
  AND U19912 ( .A(a[10]), .B(b[9]), .Z(n19253) );
  NANDN U19913 ( .A(n19254), .B(n19253), .Z(n19256) );
  XNOR U19914 ( .A(n19252), .B(n19251), .Z(n19595) );
  XNOR U19915 ( .A(n19254), .B(n19253), .Z(n19594) );
  NAND U19916 ( .A(n19595), .B(n19594), .Z(n19255) );
  AND U19917 ( .A(n19256), .B(n19255), .Z(n19260) );
  XOR U19918 ( .A(n19258), .B(n19257), .Z(n19259) );
  NANDN U19919 ( .A(n19260), .B(n19259), .Z(n19262) );
  NAND U19920 ( .A(a[11]), .B(b[9]), .Z(n19602) );
  XNOR U19921 ( .A(n19260), .B(n19259), .Z(n19603) );
  NANDN U19922 ( .A(n19602), .B(n19603), .Z(n19261) );
  AND U19923 ( .A(n19262), .B(n19261), .Z(n19266) );
  AND U19924 ( .A(a[12]), .B(b[9]), .Z(n19265) );
  NANDN U19925 ( .A(n19266), .B(n19265), .Z(n19268) );
  XNOR U19926 ( .A(n19264), .B(n19263), .Z(n19607) );
  XNOR U19927 ( .A(n19266), .B(n19265), .Z(n19606) );
  NAND U19928 ( .A(n19607), .B(n19606), .Z(n19267) );
  AND U19929 ( .A(n19268), .B(n19267), .Z(n19272) );
  XOR U19930 ( .A(n19270), .B(n19269), .Z(n19271) );
  NANDN U19931 ( .A(n19272), .B(n19271), .Z(n19274) );
  NAND U19932 ( .A(a[13]), .B(b[9]), .Z(n19614) );
  XNOR U19933 ( .A(n19272), .B(n19271), .Z(n19615) );
  NANDN U19934 ( .A(n19614), .B(n19615), .Z(n19273) );
  AND U19935 ( .A(n19274), .B(n19273), .Z(n19278) );
  AND U19936 ( .A(a[14]), .B(b[9]), .Z(n19277) );
  NANDN U19937 ( .A(n19278), .B(n19277), .Z(n19280) );
  XNOR U19938 ( .A(n19276), .B(n19275), .Z(n19619) );
  XNOR U19939 ( .A(n19278), .B(n19277), .Z(n19618) );
  NAND U19940 ( .A(n19619), .B(n19618), .Z(n19279) );
  AND U19941 ( .A(n19280), .B(n19279), .Z(n19284) );
  XOR U19942 ( .A(n19282), .B(n19281), .Z(n19283) );
  NANDN U19943 ( .A(n19284), .B(n19283), .Z(n19286) );
  NAND U19944 ( .A(a[15]), .B(b[9]), .Z(n19626) );
  XNOR U19945 ( .A(n19284), .B(n19283), .Z(n19627) );
  NANDN U19946 ( .A(n19626), .B(n19627), .Z(n19285) );
  AND U19947 ( .A(n19286), .B(n19285), .Z(n19290) );
  AND U19948 ( .A(a[16]), .B(b[9]), .Z(n19289) );
  NANDN U19949 ( .A(n19290), .B(n19289), .Z(n19292) );
  XNOR U19950 ( .A(n19288), .B(n19287), .Z(n19537) );
  XNOR U19951 ( .A(n19290), .B(n19289), .Z(n19536) );
  NAND U19952 ( .A(n19537), .B(n19536), .Z(n19291) );
  NAND U19953 ( .A(n19292), .B(n19291), .Z(n19633) );
  NAND U19954 ( .A(a[17]), .B(b[9]), .Z(n19635) );
  AND U19955 ( .A(a[18]), .B(b[9]), .Z(n19297) );
  NANDN U19956 ( .A(n19298), .B(n19297), .Z(n19300) );
  XNOR U19957 ( .A(n19294), .B(n19293), .Z(n19295) );
  XNOR U19958 ( .A(n19296), .B(n19295), .Z(n19535) );
  XNOR U19959 ( .A(n19298), .B(n19297), .Z(n19534) );
  NAND U19960 ( .A(n19535), .B(n19534), .Z(n19299) );
  NAND U19961 ( .A(n19300), .B(n19299), .Z(n19639) );
  NAND U19962 ( .A(a[19]), .B(b[9]), .Z(n19641) );
  AND U19963 ( .A(a[20]), .B(b[9]), .Z(n19305) );
  NANDN U19964 ( .A(n19306), .B(n19305), .Z(n19308) );
  XNOR U19965 ( .A(n19302), .B(n19301), .Z(n19303) );
  XNOR U19966 ( .A(n19304), .B(n19303), .Z(n19533) );
  XNOR U19967 ( .A(n19306), .B(n19305), .Z(n19532) );
  NAND U19968 ( .A(n19533), .B(n19532), .Z(n19307) );
  NAND U19969 ( .A(n19308), .B(n19307), .Z(n19649) );
  NAND U19970 ( .A(a[21]), .B(b[9]), .Z(n19651) );
  AND U19971 ( .A(a[22]), .B(b[9]), .Z(n19313) );
  NANDN U19972 ( .A(n19314), .B(n19313), .Z(n19316) );
  XNOR U19973 ( .A(n19310), .B(n19309), .Z(n19311) );
  XNOR U19974 ( .A(n19312), .B(n19311), .Z(n19531) );
  XNOR U19975 ( .A(n19314), .B(n19313), .Z(n19530) );
  NAND U19976 ( .A(n19531), .B(n19530), .Z(n19315) );
  NAND U19977 ( .A(n19316), .B(n19315), .Z(n19655) );
  NAND U19978 ( .A(a[23]), .B(b[9]), .Z(n19657) );
  AND U19979 ( .A(a[24]), .B(b[9]), .Z(n19321) );
  NANDN U19980 ( .A(n19322), .B(n19321), .Z(n19324) );
  XNOR U19981 ( .A(n19318), .B(n19317), .Z(n19319) );
  XNOR U19982 ( .A(n19320), .B(n19319), .Z(n19529) );
  XNOR U19983 ( .A(n19322), .B(n19321), .Z(n19528) );
  NAND U19984 ( .A(n19529), .B(n19528), .Z(n19323) );
  NAND U19985 ( .A(n19324), .B(n19323), .Z(n19663) );
  NAND U19986 ( .A(a[25]), .B(b[9]), .Z(n19665) );
  AND U19987 ( .A(a[26]), .B(b[9]), .Z(n19325) );
  NANDN U19988 ( .A(n19326), .B(n19325), .Z(n19332) );
  XOR U19989 ( .A(n19326), .B(n19325), .Z(n19526) );
  XOR U19990 ( .A(n19328), .B(n19327), .Z(n19329) );
  XNOR U19991 ( .A(n19330), .B(n19329), .Z(n19527) );
  NANDN U19992 ( .A(n19526), .B(n19527), .Z(n19331) );
  NAND U19993 ( .A(n19332), .B(n19331), .Z(n19671) );
  XOR U19994 ( .A(n19334), .B(n19333), .Z(n19670) );
  AND U19995 ( .A(a[27]), .B(b[9]), .Z(n19673) );
  NANDN U19996 ( .A(n19339), .B(n19340), .Z(n19342) );
  XOR U19997 ( .A(n19336), .B(n19335), .Z(n19337) );
  XNOR U19998 ( .A(n19338), .B(n19337), .Z(n19525) );
  XNOR U19999 ( .A(n19340), .B(n19339), .Z(n19524) );
  NAND U20000 ( .A(n19525), .B(n19524), .Z(n19341) );
  NAND U20001 ( .A(n19342), .B(n19341), .Z(n19681) );
  AND U20002 ( .A(a[29]), .B(b[9]), .Z(n19683) );
  AND U20003 ( .A(a[30]), .B(b[9]), .Z(n19347) );
  NANDN U20004 ( .A(n19348), .B(n19347), .Z(n19350) );
  XNOR U20005 ( .A(n19344), .B(n19343), .Z(n19345) );
  XNOR U20006 ( .A(n19346), .B(n19345), .Z(n19687) );
  XNOR U20007 ( .A(n19348), .B(n19347), .Z(n19686) );
  NAND U20008 ( .A(n19687), .B(n19686), .Z(n19349) );
  NAND U20009 ( .A(n19350), .B(n19349), .Z(n19689) );
  NAND U20010 ( .A(a[31]), .B(b[9]), .Z(n19691) );
  AND U20011 ( .A(a[32]), .B(b[9]), .Z(n19355) );
  NANDN U20012 ( .A(n19356), .B(n19355), .Z(n19358) );
  XNOR U20013 ( .A(n19352), .B(n19351), .Z(n19353) );
  XNOR U20014 ( .A(n19354), .B(n19353), .Z(n19523) );
  XNOR U20015 ( .A(n19356), .B(n19355), .Z(n19522) );
  NAND U20016 ( .A(n19523), .B(n19522), .Z(n19357) );
  NAND U20017 ( .A(n19358), .B(n19357), .Z(n19696) );
  AND U20018 ( .A(a[33]), .B(b[9]), .Z(n19699) );
  AND U20019 ( .A(a[34]), .B(b[9]), .Z(n19363) );
  NANDN U20020 ( .A(n19364), .B(n19363), .Z(n19366) );
  XOR U20021 ( .A(n19360), .B(n19359), .Z(n19361) );
  XNOR U20022 ( .A(n19362), .B(n19361), .Z(n19521) );
  XNOR U20023 ( .A(n19364), .B(n19363), .Z(n19520) );
  NAND U20024 ( .A(n19521), .B(n19520), .Z(n19365) );
  NAND U20025 ( .A(n19366), .B(n19365), .Z(n19705) );
  NAND U20026 ( .A(a[35]), .B(b[9]), .Z(n19707) );
  AND U20027 ( .A(a[36]), .B(b[9]), .Z(n19371) );
  NANDN U20028 ( .A(n19372), .B(n19371), .Z(n19374) );
  XNOR U20029 ( .A(n19368), .B(n19367), .Z(n19369) );
  XNOR U20030 ( .A(n19370), .B(n19369), .Z(n19519) );
  XNOR U20031 ( .A(n19372), .B(n19371), .Z(n19518) );
  NAND U20032 ( .A(n19519), .B(n19518), .Z(n19373) );
  NAND U20033 ( .A(n19374), .B(n19373), .Z(n19713) );
  NAND U20034 ( .A(a[37]), .B(b[9]), .Z(n19715) );
  AND U20035 ( .A(a[38]), .B(b[9]), .Z(n19379) );
  NANDN U20036 ( .A(n19380), .B(n19379), .Z(n19382) );
  XNOR U20037 ( .A(n19376), .B(n19375), .Z(n19377) );
  XNOR U20038 ( .A(n19378), .B(n19377), .Z(n19517) );
  XNOR U20039 ( .A(n19380), .B(n19379), .Z(n19516) );
  NAND U20040 ( .A(n19517), .B(n19516), .Z(n19381) );
  AND U20041 ( .A(n19382), .B(n19381), .Z(n19721) );
  XNOR U20042 ( .A(n19384), .B(n19383), .Z(n19720) );
  NAND U20043 ( .A(a[39]), .B(b[9]), .Z(n19723) );
  AND U20044 ( .A(a[40]), .B(b[9]), .Z(n19389) );
  NANDN U20045 ( .A(n19390), .B(n19389), .Z(n19392) );
  XNOR U20046 ( .A(n19386), .B(n19385), .Z(n19387) );
  XNOR U20047 ( .A(n19388), .B(n19387), .Z(n19515) );
  XNOR U20048 ( .A(n19390), .B(n19389), .Z(n19514) );
  NAND U20049 ( .A(n19515), .B(n19514), .Z(n19391) );
  NAND U20050 ( .A(n19392), .B(n19391), .Z(n19731) );
  NAND U20051 ( .A(a[41]), .B(b[9]), .Z(n19733) );
  AND U20052 ( .A(a[42]), .B(b[9]), .Z(n19393) );
  NANDN U20053 ( .A(n19394), .B(n19393), .Z(n19400) );
  XNOR U20054 ( .A(n19394), .B(n19393), .Z(n19513) );
  XOR U20055 ( .A(n19396), .B(n19395), .Z(n19397) );
  XNOR U20056 ( .A(n19398), .B(n19397), .Z(n19512) );
  NAND U20057 ( .A(n19513), .B(n19512), .Z(n19399) );
  NAND U20058 ( .A(n19400), .B(n19399), .Z(n19737) );
  NAND U20059 ( .A(a[43]), .B(b[9]), .Z(n19739) );
  IV U20060 ( .A(n19401), .Z(n19509) );
  OR U20061 ( .A(n19508), .B(n19509), .Z(n19408) );
  ANDN U20062 ( .B(n19508), .A(n19401), .Z(n19406) );
  XOR U20063 ( .A(n19403), .B(n19402), .Z(n19404) );
  XNOR U20064 ( .A(n19405), .B(n19404), .Z(n19511) );
  OR U20065 ( .A(n19406), .B(n19511), .Z(n19407) );
  AND U20066 ( .A(n19408), .B(n19407), .Z(n19745) );
  NAND U20067 ( .A(a[45]), .B(b[9]), .Z(n19748) );
  NANDN U20068 ( .A(n19761), .B(n19762), .Z(n19415) );
  NOR U20069 ( .A(n19412), .B(n19762), .Z(n19413) );
  AND U20070 ( .A(a[47]), .B(b[9]), .Z(n19760) );
  NANDN U20071 ( .A(n19413), .B(n19760), .Z(n19414) );
  AND U20072 ( .A(n19415), .B(n19414), .Z(n19421) );
  AND U20073 ( .A(a[48]), .B(b[9]), .Z(n19420) );
  NANDN U20074 ( .A(n19421), .B(n19420), .Z(n19423) );
  XOR U20075 ( .A(n19417), .B(n19416), .Z(n19418) );
  XNOR U20076 ( .A(n19419), .B(n19418), .Z(n19507) );
  XNOR U20077 ( .A(n19421), .B(n19420), .Z(n19506) );
  NAND U20078 ( .A(n19507), .B(n19506), .Z(n19422) );
  NAND U20079 ( .A(n19423), .B(n19422), .Z(n19768) );
  NAND U20080 ( .A(a[49]), .B(b[9]), .Z(n19770) );
  AND U20081 ( .A(a[50]), .B(b[9]), .Z(n19427) );
  NANDN U20082 ( .A(n19428), .B(n19427), .Z(n19430) );
  XNOR U20083 ( .A(n19428), .B(n19427), .Z(n19504) );
  NAND U20084 ( .A(n19505), .B(n19504), .Z(n19429) );
  NAND U20085 ( .A(n19430), .B(n19429), .Z(n19776) );
  NAND U20086 ( .A(a[51]), .B(b[9]), .Z(n19778) );
  AND U20087 ( .A(a[52]), .B(b[9]), .Z(n19435) );
  NANDN U20088 ( .A(n19436), .B(n19435), .Z(n19438) );
  XNOR U20089 ( .A(n19432), .B(n19431), .Z(n19433) );
  XNOR U20090 ( .A(n19434), .B(n19433), .Z(n19503) );
  XNOR U20091 ( .A(n19436), .B(n19435), .Z(n19502) );
  NAND U20092 ( .A(n19503), .B(n19502), .Z(n19437) );
  AND U20093 ( .A(n19438), .B(n19437), .Z(n19785) );
  AND U20094 ( .A(a[53]), .B(b[9]), .Z(n19788) );
  AND U20095 ( .A(a[54]), .B(b[9]), .Z(n19439) );
  NAND U20096 ( .A(n19440), .B(n19439), .Z(n19446) );
  XOR U20097 ( .A(n19440), .B(n19439), .Z(n19792) );
  XOR U20098 ( .A(n19442), .B(n19441), .Z(n19443) );
  XOR U20099 ( .A(n19444), .B(n19443), .Z(n19791) );
  NAND U20100 ( .A(n19792), .B(n19791), .Z(n19445) );
  AND U20101 ( .A(n19446), .B(n19445), .Z(n19448) );
  NANDN U20102 ( .A(n19447), .B(n19448), .Z(n19450) );
  NAND U20103 ( .A(a[55]), .B(b[9]), .Z(n19795) );
  NAND U20104 ( .A(n19796), .B(n19795), .Z(n19449) );
  AND U20105 ( .A(n19450), .B(n19449), .Z(n19804) );
  XNOR U20106 ( .A(n19452), .B(n19451), .Z(n19498) );
  XOR U20107 ( .A(n19454), .B(n19453), .Z(n19499) );
  AND U20108 ( .A(a[58]), .B(b[9]), .Z(n19457) );
  XOR U20109 ( .A(n19456), .B(n19455), .Z(n19496) );
  XOR U20110 ( .A(n19458), .B(n19457), .Z(n19497) );
  XOR U20111 ( .A(n19460), .B(n19459), .Z(n19493) );
  XOR U20112 ( .A(n19462), .B(n19461), .Z(n19492) );
  XOR U20113 ( .A(n19464), .B(n19463), .Z(n19490) );
  XOR U20114 ( .A(n19466), .B(n19465), .Z(n19491) );
  AND U20115 ( .A(a[61]), .B(b[9]), .Z(n19469) );
  XOR U20116 ( .A(n19468), .B(n19467), .Z(n19486) );
  XOR U20117 ( .A(n19470), .B(n19469), .Z(n19487) );
  AND U20118 ( .A(a[62]), .B(b[9]), .Z(n19473) );
  XOR U20119 ( .A(n19472), .B(n19471), .Z(n19484) );
  XOR U20120 ( .A(n19474), .B(n19473), .Z(n19485) );
  XOR U20121 ( .A(n19476), .B(n19475), .Z(n19483) );
  XOR U20122 ( .A(n19478), .B(n19477), .Z(n19482) );
  XOR U20123 ( .A(n19480), .B(n19479), .Z(n24697) );
  NANDN U20124 ( .A(n24698), .B(n24697), .Z(n24703) );
  XOR U20125 ( .A(n19483), .B(n19482), .Z(n20148) );
  XOR U20126 ( .A(n19485), .B(n19484), .Z(n19821) );
  XNOR U20127 ( .A(n19487), .B(n19486), .Z(n19489) );
  AND U20128 ( .A(a[62]), .B(b[8]), .Z(n19488) );
  NAND U20129 ( .A(n19489), .B(n19488), .Z(n19820) );
  XOR U20130 ( .A(n19489), .B(n19488), .Z(n20141) );
  XOR U20131 ( .A(n19491), .B(n19490), .Z(n19815) );
  AND U20132 ( .A(a[60]), .B(b[8]), .Z(n19494) );
  XOR U20133 ( .A(n19493), .B(n19492), .Z(n19495) );
  NAND U20134 ( .A(n19494), .B(n19495), .Z(n19814) );
  XOR U20135 ( .A(n19495), .B(n19494), .Z(n20133) );
  XOR U20136 ( .A(n19497), .B(n19496), .Z(n19809) );
  XNOR U20137 ( .A(n19499), .B(n19498), .Z(n19501) );
  AND U20138 ( .A(a[58]), .B(b[8]), .Z(n19500) );
  NAND U20139 ( .A(n19501), .B(n19500), .Z(n19808) );
  XOR U20140 ( .A(n19501), .B(n19500), .Z(n20127) );
  AND U20141 ( .A(a[57]), .B(b[8]), .Z(n19799) );
  XNOR U20142 ( .A(n19503), .B(n19502), .Z(n20106) );
  XNOR U20143 ( .A(n19505), .B(n19504), .Z(n20100) );
  XOR U20144 ( .A(n19507), .B(n19506), .Z(n19763) );
  IV U20145 ( .A(n19763), .Z(n20092) );
  NAND U20146 ( .A(a[48]), .B(b[8]), .Z(n19834) );
  XOR U20147 ( .A(n19509), .B(n19508), .Z(n19510) );
  XNOR U20148 ( .A(n19511), .B(n19510), .Z(n20075) );
  XNOR U20149 ( .A(n19513), .B(n19512), .Z(n20067) );
  XNOR U20150 ( .A(n19515), .B(n19514), .Z(n20059) );
  XNOR U20151 ( .A(n19517), .B(n19516), .Z(n20051) );
  XNOR U20152 ( .A(n19519), .B(n19518), .Z(n20043) );
  XNOR U20153 ( .A(n19521), .B(n19520), .Z(n20035) );
  XNOR U20154 ( .A(n19523), .B(n19522), .Z(n20027) );
  AND U20155 ( .A(a[30]), .B(b[8]), .Z(n19679) );
  XNOR U20156 ( .A(n19525), .B(n19524), .Z(n20011) );
  NAND U20157 ( .A(a[28]), .B(b[8]), .Z(n19674) );
  XNOR U20158 ( .A(n19527), .B(n19526), .Z(n20004) );
  AND U20159 ( .A(a[26]), .B(b[8]), .Z(n19667) );
  XNOR U20160 ( .A(n19529), .B(n19528), .Z(n19995) );
  XNOR U20161 ( .A(n19531), .B(n19530), .Z(n19987) );
  XNOR U20162 ( .A(n19533), .B(n19532), .Z(n19981) );
  XNOR U20163 ( .A(n19535), .B(n19534), .Z(n19971) );
  XNOR U20164 ( .A(n19537), .B(n19536), .Z(n19963) );
  AND U20165 ( .A(a[8]), .B(b[8]), .Z(n19579) );
  XOR U20166 ( .A(n19539), .B(n19538), .Z(n19561) );
  AND U20167 ( .A(a[0]), .B(b[8]), .Z(n20210) );
  AND U20168 ( .A(a[1]), .B(b[9]), .Z(n19543) );
  AND U20169 ( .A(n20210), .B(n19543), .Z(n19540) );
  NAND U20170 ( .A(a[2]), .B(n19540), .Z(n19547) );
  NAND U20171 ( .A(b[9]), .B(a[1]), .Z(n19541) );
  XOR U20172 ( .A(n19542), .B(n19541), .Z(n19881) );
  NAND U20173 ( .A(n19543), .B(a[0]), .Z(n19544) );
  XNOR U20174 ( .A(a[2]), .B(n19544), .Z(n19545) );
  AND U20175 ( .A(b[8]), .B(n19545), .Z(n19882) );
  NANDN U20176 ( .A(n19881), .B(n19882), .Z(n19546) );
  AND U20177 ( .A(n19547), .B(n19546), .Z(n19550) );
  NANDN U20178 ( .A(n19550), .B(n19551), .Z(n19553) );
  NAND U20179 ( .A(a[3]), .B(b[8]), .Z(n19889) );
  NANDN U20180 ( .A(n19889), .B(n19890), .Z(n19552) );
  AND U20181 ( .A(n19553), .B(n19552), .Z(n19555) );
  AND U20182 ( .A(a[4]), .B(b[8]), .Z(n19554) );
  NANDN U20183 ( .A(n19555), .B(n19554), .Z(n19559) );
  XNOR U20184 ( .A(n19555), .B(n19554), .Z(n19894) );
  XNOR U20185 ( .A(n19557), .B(n19556), .Z(n19893) );
  NAND U20186 ( .A(n19894), .B(n19893), .Z(n19558) );
  NAND U20187 ( .A(n19559), .B(n19558), .Z(n19560) );
  NAND U20188 ( .A(n19561), .B(n19560), .Z(n19563) );
  NAND U20189 ( .A(a[5]), .B(b[8]), .Z(n19899) );
  XOR U20190 ( .A(n19561), .B(n19560), .Z(n19900) );
  NANDN U20191 ( .A(n19899), .B(n19900), .Z(n19562) );
  AND U20192 ( .A(n19563), .B(n19562), .Z(n19567) );
  XNOR U20193 ( .A(n19565), .B(n19564), .Z(n19566) );
  NANDN U20194 ( .A(n19567), .B(n19566), .Z(n19569) );
  NAND U20195 ( .A(a[6]), .B(b[8]), .Z(n19905) );
  XNOR U20196 ( .A(n19567), .B(n19566), .Z(n19906) );
  NANDN U20197 ( .A(n19905), .B(n19906), .Z(n19568) );
  AND U20198 ( .A(n19569), .B(n19568), .Z(n19573) );
  XNOR U20199 ( .A(n19571), .B(n19570), .Z(n19572) );
  NANDN U20200 ( .A(n19573), .B(n19572), .Z(n19575) );
  NAND U20201 ( .A(a[7]), .B(b[8]), .Z(n19913) );
  XNOR U20202 ( .A(n19573), .B(n19572), .Z(n19914) );
  NANDN U20203 ( .A(n19913), .B(n19914), .Z(n19574) );
  AND U20204 ( .A(n19575), .B(n19574), .Z(n19578) );
  NANDN U20205 ( .A(n19579), .B(n19578), .Z(n19581) );
  XOR U20206 ( .A(n19577), .B(n19576), .Z(n19872) );
  XNOR U20207 ( .A(n19579), .B(n19578), .Z(n19871) );
  NANDN U20208 ( .A(n19872), .B(n19871), .Z(n19580) );
  AND U20209 ( .A(n19581), .B(n19580), .Z(n19585) );
  XOR U20210 ( .A(n19583), .B(n19582), .Z(n19584) );
  NAND U20211 ( .A(n19585), .B(n19584), .Z(n19587) );
  NAND U20212 ( .A(a[9]), .B(b[8]), .Z(n19921) );
  XOR U20213 ( .A(n19585), .B(n19584), .Z(n19922) );
  NANDN U20214 ( .A(n19921), .B(n19922), .Z(n19586) );
  AND U20215 ( .A(n19587), .B(n19586), .Z(n19589) );
  AND U20216 ( .A(a[10]), .B(b[8]), .Z(n19588) );
  NANDN U20217 ( .A(n19589), .B(n19588), .Z(n19593) );
  XNOR U20218 ( .A(n19589), .B(n19588), .Z(n19928) );
  XNOR U20219 ( .A(n19591), .B(n19590), .Z(n19927) );
  NAND U20220 ( .A(n19928), .B(n19927), .Z(n19592) );
  AND U20221 ( .A(n19593), .B(n19592), .Z(n19597) );
  XOR U20222 ( .A(n19595), .B(n19594), .Z(n19596) );
  NANDN U20223 ( .A(n19597), .B(n19596), .Z(n19599) );
  NAND U20224 ( .A(a[11]), .B(b[8]), .Z(n19933) );
  XNOR U20225 ( .A(n19597), .B(n19596), .Z(n19934) );
  NANDN U20226 ( .A(n19933), .B(n19934), .Z(n19598) );
  AND U20227 ( .A(n19599), .B(n19598), .Z(n19601) );
  AND U20228 ( .A(a[12]), .B(b[8]), .Z(n19600) );
  NANDN U20229 ( .A(n19601), .B(n19600), .Z(n19605) );
  XNOR U20230 ( .A(n19601), .B(n19600), .Z(n19940) );
  XNOR U20231 ( .A(n19603), .B(n19602), .Z(n19939) );
  NAND U20232 ( .A(n19940), .B(n19939), .Z(n19604) );
  AND U20233 ( .A(n19605), .B(n19604), .Z(n19609) );
  XOR U20234 ( .A(n19607), .B(n19606), .Z(n19608) );
  NANDN U20235 ( .A(n19609), .B(n19608), .Z(n19611) );
  NAND U20236 ( .A(a[13]), .B(b[8]), .Z(n19945) );
  XNOR U20237 ( .A(n19609), .B(n19608), .Z(n19946) );
  NANDN U20238 ( .A(n19945), .B(n19946), .Z(n19610) );
  AND U20239 ( .A(n19611), .B(n19610), .Z(n19613) );
  AND U20240 ( .A(a[14]), .B(b[8]), .Z(n19612) );
  NANDN U20241 ( .A(n19613), .B(n19612), .Z(n19617) );
  XNOR U20242 ( .A(n19613), .B(n19612), .Z(n19952) );
  XNOR U20243 ( .A(n19615), .B(n19614), .Z(n19951) );
  NAND U20244 ( .A(n19952), .B(n19951), .Z(n19616) );
  AND U20245 ( .A(n19617), .B(n19616), .Z(n19621) );
  XOR U20246 ( .A(n19619), .B(n19618), .Z(n19620) );
  NANDN U20247 ( .A(n19621), .B(n19620), .Z(n19623) );
  NAND U20248 ( .A(a[15]), .B(b[8]), .Z(n19957) );
  XNOR U20249 ( .A(n19621), .B(n19620), .Z(n19958) );
  NANDN U20250 ( .A(n19957), .B(n19958), .Z(n19622) );
  AND U20251 ( .A(n19623), .B(n19622), .Z(n19625) );
  AND U20252 ( .A(a[16]), .B(b[8]), .Z(n19624) );
  NANDN U20253 ( .A(n19625), .B(n19624), .Z(n19629) );
  XNOR U20254 ( .A(n19625), .B(n19624), .Z(n19870) );
  XNOR U20255 ( .A(n19627), .B(n19626), .Z(n19869) );
  NAND U20256 ( .A(n19870), .B(n19869), .Z(n19628) );
  NAND U20257 ( .A(n19629), .B(n19628), .Z(n19964) );
  NAND U20258 ( .A(a[17]), .B(b[8]), .Z(n19966) );
  AND U20259 ( .A(a[18]), .B(b[8]), .Z(n19630) );
  NANDN U20260 ( .A(n19631), .B(n19630), .Z(n19637) );
  XOR U20261 ( .A(n19631), .B(n19630), .Z(n19867) );
  XNOR U20262 ( .A(n19633), .B(n19632), .Z(n19634) );
  XNOR U20263 ( .A(n19635), .B(n19634), .Z(n19868) );
  NANDN U20264 ( .A(n19867), .B(n19868), .Z(n19636) );
  NAND U20265 ( .A(n19637), .B(n19636), .Z(n19972) );
  NAND U20266 ( .A(a[19]), .B(b[8]), .Z(n19974) );
  AND U20267 ( .A(a[20]), .B(b[8]), .Z(n19642) );
  NANDN U20268 ( .A(n19643), .B(n19642), .Z(n19645) );
  XNOR U20269 ( .A(n19639), .B(n19638), .Z(n19640) );
  XNOR U20270 ( .A(n19641), .B(n19640), .Z(n19866) );
  XNOR U20271 ( .A(n19643), .B(n19642), .Z(n19865) );
  NAND U20272 ( .A(n19866), .B(n19865), .Z(n19644) );
  NAND U20273 ( .A(n19645), .B(n19644), .Z(n19982) );
  NAND U20274 ( .A(a[21]), .B(b[8]), .Z(n19984) );
  AND U20275 ( .A(a[22]), .B(b[8]), .Z(n19646) );
  NANDN U20276 ( .A(n19647), .B(n19646), .Z(n19653) );
  XOR U20277 ( .A(n19647), .B(n19646), .Z(n19863) );
  XNOR U20278 ( .A(n19649), .B(n19648), .Z(n19650) );
  XNOR U20279 ( .A(n19651), .B(n19650), .Z(n19864) );
  NANDN U20280 ( .A(n19863), .B(n19864), .Z(n19652) );
  NAND U20281 ( .A(n19653), .B(n19652), .Z(n19988) );
  NAND U20282 ( .A(a[23]), .B(b[8]), .Z(n19990) );
  AND U20283 ( .A(a[24]), .B(b[8]), .Z(n19658) );
  NANDN U20284 ( .A(n19659), .B(n19658), .Z(n19661) );
  XNOR U20285 ( .A(n19655), .B(n19654), .Z(n19656) );
  XNOR U20286 ( .A(n19657), .B(n19656), .Z(n19862) );
  XNOR U20287 ( .A(n19659), .B(n19658), .Z(n19861) );
  NAND U20288 ( .A(n19862), .B(n19861), .Z(n19660) );
  NAND U20289 ( .A(n19661), .B(n19660), .Z(n19996) );
  NAND U20290 ( .A(a[25]), .B(b[8]), .Z(n19998) );
  NANDN U20291 ( .A(n19667), .B(n19666), .Z(n19669) );
  XOR U20292 ( .A(n19663), .B(n19662), .Z(n19664) );
  XOR U20293 ( .A(n19665), .B(n19664), .Z(n19860) );
  XNOR U20294 ( .A(n19667), .B(n19666), .Z(n19859) );
  NANDN U20295 ( .A(n19860), .B(n19859), .Z(n19668) );
  NAND U20296 ( .A(n19669), .B(n19668), .Z(n20003) );
  AND U20297 ( .A(a[27]), .B(b[8]), .Z(n20006) );
  NANDN U20298 ( .A(n19674), .B(n19675), .Z(n19677) );
  XOR U20299 ( .A(n19671), .B(n19670), .Z(n19672) );
  XNOR U20300 ( .A(n19673), .B(n19672), .Z(n19858) );
  XNOR U20301 ( .A(n19675), .B(n19674), .Z(n19857) );
  NAND U20302 ( .A(n19858), .B(n19857), .Z(n19676) );
  NAND U20303 ( .A(n19677), .B(n19676), .Z(n20012) );
  NAND U20304 ( .A(a[29]), .B(b[8]), .Z(n20014) );
  NANDN U20305 ( .A(n19679), .B(n19678), .Z(n19685) );
  XNOR U20306 ( .A(n19679), .B(n19678), .Z(n19855) );
  XNOR U20307 ( .A(n19681), .B(n19680), .Z(n19682) );
  XNOR U20308 ( .A(n19683), .B(n19682), .Z(n19856) );
  NAND U20309 ( .A(n19855), .B(n19856), .Z(n19684) );
  NAND U20310 ( .A(n19685), .B(n19684), .Z(n20020) );
  XOR U20311 ( .A(n19687), .B(n19686), .Z(n20019) );
  AND U20312 ( .A(a[31]), .B(b[8]), .Z(n20022) );
  AND U20313 ( .A(a[32]), .B(b[8]), .Z(n19692) );
  NANDN U20314 ( .A(n19693), .B(n19692), .Z(n19695) );
  XNOR U20315 ( .A(n19689), .B(n19688), .Z(n19690) );
  XNOR U20316 ( .A(n19691), .B(n19690), .Z(n19854) );
  XNOR U20317 ( .A(n19693), .B(n19692), .Z(n19853) );
  NAND U20318 ( .A(n19854), .B(n19853), .Z(n19694) );
  NAND U20319 ( .A(n19695), .B(n19694), .Z(n20028) );
  NAND U20320 ( .A(a[33]), .B(b[8]), .Z(n20030) );
  AND U20321 ( .A(a[34]), .B(b[8]), .Z(n19700) );
  NANDN U20322 ( .A(n19701), .B(n19700), .Z(n19703) );
  XOR U20323 ( .A(n19697), .B(n19696), .Z(n19698) );
  XNOR U20324 ( .A(n19699), .B(n19698), .Z(n19852) );
  XNOR U20325 ( .A(n19701), .B(n19700), .Z(n19851) );
  NAND U20326 ( .A(n19852), .B(n19851), .Z(n19702) );
  NAND U20327 ( .A(n19703), .B(n19702), .Z(n20036) );
  NAND U20328 ( .A(a[35]), .B(b[8]), .Z(n20038) );
  AND U20329 ( .A(a[36]), .B(b[8]), .Z(n19708) );
  NANDN U20330 ( .A(n19709), .B(n19708), .Z(n19711) );
  XNOR U20331 ( .A(n19705), .B(n19704), .Z(n19706) );
  XNOR U20332 ( .A(n19707), .B(n19706), .Z(n19850) );
  XNOR U20333 ( .A(n19709), .B(n19708), .Z(n19849) );
  NAND U20334 ( .A(n19850), .B(n19849), .Z(n19710) );
  NAND U20335 ( .A(n19711), .B(n19710), .Z(n20044) );
  NAND U20336 ( .A(a[37]), .B(b[8]), .Z(n20046) );
  AND U20337 ( .A(a[38]), .B(b[8]), .Z(n19716) );
  NANDN U20338 ( .A(n19717), .B(n19716), .Z(n19719) );
  XNOR U20339 ( .A(n19713), .B(n19712), .Z(n19714) );
  XNOR U20340 ( .A(n19715), .B(n19714), .Z(n19848) );
  XNOR U20341 ( .A(n19717), .B(n19716), .Z(n19847) );
  NAND U20342 ( .A(n19848), .B(n19847), .Z(n19718) );
  NAND U20343 ( .A(n19719), .B(n19718), .Z(n20052) );
  NAND U20344 ( .A(a[39]), .B(b[8]), .Z(n20054) );
  AND U20345 ( .A(a[40]), .B(b[8]), .Z(n19724) );
  NANDN U20346 ( .A(n19725), .B(n19724), .Z(n19727) );
  XNOR U20347 ( .A(n19721), .B(n19720), .Z(n19722) );
  XNOR U20348 ( .A(n19723), .B(n19722), .Z(n19846) );
  XNOR U20349 ( .A(n19725), .B(n19724), .Z(n19845) );
  NAND U20350 ( .A(n19846), .B(n19845), .Z(n19726) );
  NAND U20351 ( .A(n19727), .B(n19726), .Z(n20060) );
  NAND U20352 ( .A(a[41]), .B(b[8]), .Z(n20062) );
  AND U20353 ( .A(a[42]), .B(b[8]), .Z(n19728) );
  NANDN U20354 ( .A(n19729), .B(n19728), .Z(n19735) );
  XOR U20355 ( .A(n19729), .B(n19728), .Z(n19843) );
  XNOR U20356 ( .A(n19731), .B(n19730), .Z(n19732) );
  XNOR U20357 ( .A(n19733), .B(n19732), .Z(n19844) );
  NANDN U20358 ( .A(n19843), .B(n19844), .Z(n19734) );
  NAND U20359 ( .A(n19735), .B(n19734), .Z(n20068) );
  NAND U20360 ( .A(a[43]), .B(b[8]), .Z(n20070) );
  AND U20361 ( .A(a[44]), .B(b[8]), .Z(n19741) );
  NANDN U20362 ( .A(n19740), .B(n19741), .Z(n19743) );
  XNOR U20363 ( .A(n19737), .B(n19736), .Z(n19738) );
  XNOR U20364 ( .A(n19739), .B(n19738), .Z(n19842) );
  XNOR U20365 ( .A(n19741), .B(n19740), .Z(n19841) );
  NAND U20366 ( .A(n19842), .B(n19841), .Z(n19742) );
  NAND U20367 ( .A(n19743), .B(n19742), .Z(n20076) );
  NAND U20368 ( .A(a[45]), .B(b[8]), .Z(n20078) );
  AND U20369 ( .A(a[46]), .B(b[8]), .Z(n19744) );
  IV U20370 ( .A(n19744), .Z(n19837) );
  OR U20371 ( .A(n19838), .B(n19837), .Z(n19751) );
  ANDN U20372 ( .B(n19838), .A(n19744), .Z(n19749) );
  XOR U20373 ( .A(n19746), .B(n19745), .Z(n19747) );
  XOR U20374 ( .A(n19748), .B(n19747), .Z(n19840) );
  NANDN U20375 ( .A(n19749), .B(n19840), .Z(n19750) );
  AND U20376 ( .A(n19751), .B(n19750), .Z(n20084) );
  XOR U20377 ( .A(n19753), .B(n19752), .Z(n19754) );
  XOR U20378 ( .A(n19755), .B(n19754), .Z(n19756) );
  IV U20379 ( .A(n19756), .Z(n20083) );
  OR U20380 ( .A(n20084), .B(n20083), .Z(n19759) );
  ANDN U20381 ( .B(n20084), .A(n19756), .Z(n19757) );
  NAND U20382 ( .A(a[47]), .B(b[8]), .Z(n20086) );
  OR U20383 ( .A(n19757), .B(n20086), .Z(n19758) );
  AND U20384 ( .A(n19759), .B(n19758), .Z(n19833) );
  NANDN U20385 ( .A(n20092), .B(n20093), .Z(n19766) );
  NOR U20386 ( .A(n19763), .B(n20093), .Z(n19764) );
  AND U20387 ( .A(a[49]), .B(b[8]), .Z(n20091) );
  NANDN U20388 ( .A(n19764), .B(n20091), .Z(n19765) );
  AND U20389 ( .A(n19766), .B(n19765), .Z(n19771) );
  AND U20390 ( .A(a[50]), .B(b[8]), .Z(n19772) );
  NANDN U20391 ( .A(n19771), .B(n19772), .Z(n19774) );
  XNOR U20392 ( .A(n19768), .B(n19767), .Z(n19769) );
  XNOR U20393 ( .A(n19770), .B(n19769), .Z(n19832) );
  XNOR U20394 ( .A(n19772), .B(n19771), .Z(n19831) );
  NAND U20395 ( .A(n19832), .B(n19831), .Z(n19773) );
  NAND U20396 ( .A(n19774), .B(n19773), .Z(n20101) );
  NAND U20397 ( .A(a[51]), .B(b[8]), .Z(n20103) );
  AND U20398 ( .A(a[52]), .B(b[8]), .Z(n19780) );
  NANDN U20399 ( .A(n19779), .B(n19780), .Z(n19782) );
  XNOR U20400 ( .A(n19776), .B(n19775), .Z(n19777) );
  XNOR U20401 ( .A(n19778), .B(n19777), .Z(n19830) );
  XNOR U20402 ( .A(n19780), .B(n19779), .Z(n19829) );
  NAND U20403 ( .A(n19830), .B(n19829), .Z(n19781) );
  NAND U20404 ( .A(n19782), .B(n19781), .Z(n20107) );
  NAND U20405 ( .A(a[53]), .B(b[8]), .Z(n20109) );
  NAND U20406 ( .A(a[54]), .B(b[8]), .Z(n19783) );
  NAND U20407 ( .A(n19784), .B(n19783), .Z(n19790) );
  XOR U20408 ( .A(n19784), .B(n19783), .Z(n19827) );
  XOR U20409 ( .A(n19786), .B(n19785), .Z(n19787) );
  XOR U20410 ( .A(n19788), .B(n19787), .Z(n19828) );
  NAND U20411 ( .A(n19827), .B(n19828), .Z(n19789) );
  NAND U20412 ( .A(n19790), .B(n19789), .Z(n20115) );
  XOR U20413 ( .A(n19792), .B(n19791), .Z(n20114) );
  NAND U20414 ( .A(a[55]), .B(b[8]), .Z(n20116) );
  AND U20415 ( .A(a[56]), .B(b[8]), .Z(n19793) );
  NANDN U20416 ( .A(n19794), .B(n19793), .Z(n19798) );
  XOR U20417 ( .A(n19794), .B(n19793), .Z(n20121) );
  XNOR U20418 ( .A(n19796), .B(n19795), .Z(n20122) );
  NANDN U20419 ( .A(n20121), .B(n20122), .Z(n19797) );
  NAND U20420 ( .A(n19798), .B(n19797), .Z(n19800) );
  NAND U20421 ( .A(n19799), .B(n19800), .Z(n19806) );
  XNOR U20422 ( .A(n19800), .B(n19799), .Z(n19825) );
  XOR U20423 ( .A(n19802), .B(n19801), .Z(n19803) );
  XNOR U20424 ( .A(n19804), .B(n19803), .Z(n19826) );
  NANDN U20425 ( .A(n19825), .B(n19826), .Z(n19805) );
  NAND U20426 ( .A(n19806), .B(n19805), .Z(n20128) );
  NAND U20427 ( .A(n20127), .B(n20128), .Z(n19807) );
  NAND U20428 ( .A(n19808), .B(n19807), .Z(n19810) );
  NAND U20429 ( .A(n19809), .B(n19810), .Z(n19812) );
  XOR U20430 ( .A(n19810), .B(n19809), .Z(n20130) );
  AND U20431 ( .A(a[59]), .B(b[8]), .Z(n20129) );
  NAND U20432 ( .A(n20130), .B(n20129), .Z(n19811) );
  NAND U20433 ( .A(n19812), .B(n19811), .Z(n20134) );
  NAND U20434 ( .A(n20133), .B(n20134), .Z(n19813) );
  NAND U20435 ( .A(n19814), .B(n19813), .Z(n19816) );
  NAND U20436 ( .A(n19815), .B(n19816), .Z(n19818) );
  XOR U20437 ( .A(n19816), .B(n19815), .Z(n20138) );
  AND U20438 ( .A(a[61]), .B(b[8]), .Z(n20137) );
  NAND U20439 ( .A(n20138), .B(n20137), .Z(n19817) );
  NAND U20440 ( .A(n19818), .B(n19817), .Z(n20142) );
  NAND U20441 ( .A(n20141), .B(n20142), .Z(n19819) );
  NAND U20442 ( .A(n19820), .B(n19819), .Z(n19822) );
  NAND U20443 ( .A(n19821), .B(n19822), .Z(n19824) );
  XOR U20444 ( .A(n19822), .B(n19821), .Z(n20146) );
  AND U20445 ( .A(a[63]), .B(b[8]), .Z(n20145) );
  NAND U20446 ( .A(n20146), .B(n20145), .Z(n19823) );
  NAND U20447 ( .A(n19824), .B(n19823), .Z(n20147) );
  XNOR U20448 ( .A(n20148), .B(n20147), .Z(n24683) );
  NAND U20449 ( .A(a[63]), .B(b[7]), .Z(n20144) );
  AND U20450 ( .A(a[62]), .B(b[7]), .Z(n20139) );
  NAND U20451 ( .A(a[61]), .B(b[7]), .Z(n20136) );
  AND U20452 ( .A(a[60]), .B(b[7]), .Z(n20131) );
  AND U20453 ( .A(a[59]), .B(b[7]), .Z(n20159) );
  XNOR U20454 ( .A(n19826), .B(n19825), .Z(n20462) );
  NAND U20455 ( .A(a[58]), .B(b[7]), .Z(n20465) );
  NAND U20456 ( .A(a[56]), .B(b[7]), .Z(n20117) );
  XNOR U20457 ( .A(n19828), .B(n19827), .Z(n20447) );
  XNOR U20458 ( .A(n19830), .B(n19829), .Z(n20440) );
  XOR U20459 ( .A(n19832), .B(n19831), .Z(n20094) );
  IV U20460 ( .A(n20094), .Z(n20432) );
  NAND U20461 ( .A(a[50]), .B(b[7]), .Z(n20168) );
  XOR U20462 ( .A(n19834), .B(n19833), .Z(n19835) );
  XOR U20463 ( .A(n19836), .B(n19835), .Z(n20087) );
  IV U20464 ( .A(n20087), .Z(n20426) );
  NAND U20465 ( .A(a[48]), .B(b[7]), .Z(n20172) );
  XOR U20466 ( .A(n19838), .B(n19837), .Z(n19839) );
  XNOR U20467 ( .A(n19840), .B(n19839), .Z(n20416) );
  XNOR U20468 ( .A(n19842), .B(n19841), .Z(n20408) );
  NAND U20469 ( .A(a[44]), .B(b[7]), .Z(n20071) );
  XNOR U20470 ( .A(n19844), .B(n19843), .Z(n20399) );
  XNOR U20471 ( .A(n19846), .B(n19845), .Z(n20390) );
  XNOR U20472 ( .A(n19848), .B(n19847), .Z(n20382) );
  XNOR U20473 ( .A(n19850), .B(n19849), .Z(n20374) );
  XNOR U20474 ( .A(n19852), .B(n19851), .Z(n20366) );
  XNOR U20475 ( .A(n19854), .B(n19853), .Z(n20360) );
  XOR U20476 ( .A(n19856), .B(n19855), .Z(n20349) );
  XNOR U20477 ( .A(n19858), .B(n19857), .Z(n20340) );
  XNOR U20478 ( .A(n19860), .B(n19859), .Z(n20330) );
  XNOR U20479 ( .A(n19862), .B(n19861), .Z(n20322) );
  NAND U20480 ( .A(a[24]), .B(b[7]), .Z(n19991) );
  XNOR U20481 ( .A(n19864), .B(n19863), .Z(n20315) );
  XNOR U20482 ( .A(n19866), .B(n19865), .Z(n20308) );
  NAND U20483 ( .A(a[20]), .B(b[7]), .Z(n19975) );
  XNOR U20484 ( .A(n19868), .B(n19867), .Z(n20299) );
  XNOR U20485 ( .A(n19870), .B(n19869), .Z(n20290) );
  XOR U20486 ( .A(n19872), .B(n19871), .Z(n19918) );
  AND U20487 ( .A(a[0]), .B(b[7]), .Z(n20531) );
  AND U20488 ( .A(a[1]), .B(b[8]), .Z(n19876) );
  AND U20489 ( .A(n20531), .B(n19876), .Z(n19873) );
  NAND U20490 ( .A(a[2]), .B(n19873), .Z(n19880) );
  NAND U20491 ( .A(b[8]), .B(a[1]), .Z(n19874) );
  XOR U20492 ( .A(n19875), .B(n19874), .Z(n20216) );
  NAND U20493 ( .A(n19876), .B(a[0]), .Z(n19877) );
  XNOR U20494 ( .A(a[2]), .B(n19877), .Z(n19878) );
  AND U20495 ( .A(b[7]), .B(n19878), .Z(n20217) );
  NANDN U20496 ( .A(n20216), .B(n20217), .Z(n19879) );
  AND U20497 ( .A(n19880), .B(n19879), .Z(n19883) );
  NANDN U20498 ( .A(n19883), .B(n19884), .Z(n19886) );
  NAND U20499 ( .A(a[3]), .B(b[7]), .Z(n20222) );
  NANDN U20500 ( .A(n20222), .B(n20223), .Z(n19885) );
  AND U20501 ( .A(n19886), .B(n19885), .Z(n19887) );
  AND U20502 ( .A(a[4]), .B(b[7]), .Z(n19888) );
  NANDN U20503 ( .A(n19887), .B(n19888), .Z(n19892) );
  NAND U20504 ( .A(n20207), .B(n20206), .Z(n19891) );
  AND U20505 ( .A(n19892), .B(n19891), .Z(n19896) );
  XOR U20506 ( .A(n19894), .B(n19893), .Z(n19895) );
  NANDN U20507 ( .A(n19896), .B(n19895), .Z(n19898) );
  XNOR U20508 ( .A(n19896), .B(n19895), .Z(n20205) );
  AND U20509 ( .A(a[5]), .B(b[7]), .Z(n20204) );
  NAND U20510 ( .A(n20205), .B(n20204), .Z(n19897) );
  AND U20511 ( .A(n19898), .B(n19897), .Z(n19902) );
  XNOR U20512 ( .A(n19900), .B(n19899), .Z(n19901) );
  NANDN U20513 ( .A(n19902), .B(n19901), .Z(n19904) );
  NAND U20514 ( .A(a[6]), .B(b[7]), .Z(n20202) );
  XNOR U20515 ( .A(n19902), .B(n19901), .Z(n20203) );
  NANDN U20516 ( .A(n20202), .B(n20203), .Z(n19903) );
  AND U20517 ( .A(n19904), .B(n19903), .Z(n19908) );
  XNOR U20518 ( .A(n19906), .B(n19905), .Z(n19907) );
  NANDN U20519 ( .A(n19908), .B(n19907), .Z(n19910) );
  NAND U20520 ( .A(a[7]), .B(b[7]), .Z(n20238) );
  XNOR U20521 ( .A(n19908), .B(n19907), .Z(n20239) );
  NANDN U20522 ( .A(n20238), .B(n20239), .Z(n19909) );
  AND U20523 ( .A(n19910), .B(n19909), .Z(n19912) );
  AND U20524 ( .A(a[8]), .B(b[7]), .Z(n19911) );
  NANDN U20525 ( .A(n19912), .B(n19911), .Z(n19916) );
  XNOR U20526 ( .A(n19912), .B(n19911), .Z(n20243) );
  XNOR U20527 ( .A(n19914), .B(n19913), .Z(n20242) );
  NAND U20528 ( .A(n20243), .B(n20242), .Z(n19915) );
  NAND U20529 ( .A(n19916), .B(n19915), .Z(n19917) );
  NAND U20530 ( .A(n19918), .B(n19917), .Z(n19920) );
  XOR U20531 ( .A(n19918), .B(n19917), .Z(n20249) );
  AND U20532 ( .A(a[9]), .B(b[7]), .Z(n20248) );
  NAND U20533 ( .A(n20249), .B(n20248), .Z(n19919) );
  AND U20534 ( .A(n19920), .B(n19919), .Z(n19924) );
  AND U20535 ( .A(a[10]), .B(b[7]), .Z(n19923) );
  NANDN U20536 ( .A(n19924), .B(n19923), .Z(n19926) );
  XNOR U20537 ( .A(n19922), .B(n19921), .Z(n20255) );
  XNOR U20538 ( .A(n19924), .B(n19923), .Z(n20254) );
  NAND U20539 ( .A(n20255), .B(n20254), .Z(n19925) );
  AND U20540 ( .A(n19926), .B(n19925), .Z(n19930) );
  XOR U20541 ( .A(n19928), .B(n19927), .Z(n19929) );
  NANDN U20542 ( .A(n19930), .B(n19929), .Z(n19932) );
  NAND U20543 ( .A(a[11]), .B(b[7]), .Z(n20262) );
  XNOR U20544 ( .A(n19930), .B(n19929), .Z(n20263) );
  NANDN U20545 ( .A(n20262), .B(n20263), .Z(n19931) );
  AND U20546 ( .A(n19932), .B(n19931), .Z(n19936) );
  AND U20547 ( .A(a[12]), .B(b[7]), .Z(n19935) );
  NANDN U20548 ( .A(n19936), .B(n19935), .Z(n19938) );
  XNOR U20549 ( .A(n19934), .B(n19933), .Z(n20267) );
  XNOR U20550 ( .A(n19936), .B(n19935), .Z(n20266) );
  NAND U20551 ( .A(n20267), .B(n20266), .Z(n19937) );
  AND U20552 ( .A(n19938), .B(n19937), .Z(n19942) );
  XOR U20553 ( .A(n19940), .B(n19939), .Z(n19941) );
  NANDN U20554 ( .A(n19942), .B(n19941), .Z(n19944) );
  NAND U20555 ( .A(a[13]), .B(b[7]), .Z(n20274) );
  XNOR U20556 ( .A(n19942), .B(n19941), .Z(n20275) );
  NANDN U20557 ( .A(n20274), .B(n20275), .Z(n19943) );
  AND U20558 ( .A(n19944), .B(n19943), .Z(n19948) );
  AND U20559 ( .A(a[14]), .B(b[7]), .Z(n19947) );
  NANDN U20560 ( .A(n19948), .B(n19947), .Z(n19950) );
  XNOR U20561 ( .A(n19946), .B(n19945), .Z(n20279) );
  XNOR U20562 ( .A(n19948), .B(n19947), .Z(n20278) );
  NAND U20563 ( .A(n20279), .B(n20278), .Z(n19949) );
  AND U20564 ( .A(n19950), .B(n19949), .Z(n19954) );
  XOR U20565 ( .A(n19952), .B(n19951), .Z(n19953) );
  NANDN U20566 ( .A(n19954), .B(n19953), .Z(n19956) );
  NAND U20567 ( .A(a[15]), .B(b[7]), .Z(n20286) );
  XNOR U20568 ( .A(n19954), .B(n19953), .Z(n20287) );
  NANDN U20569 ( .A(n20286), .B(n20287), .Z(n19955) );
  AND U20570 ( .A(n19956), .B(n19955), .Z(n19960) );
  AND U20571 ( .A(a[16]), .B(b[7]), .Z(n19959) );
  NANDN U20572 ( .A(n19960), .B(n19959), .Z(n19962) );
  XNOR U20573 ( .A(n19958), .B(n19957), .Z(n20201) );
  XNOR U20574 ( .A(n19960), .B(n19959), .Z(n20200) );
  NAND U20575 ( .A(n20201), .B(n20200), .Z(n19961) );
  NAND U20576 ( .A(n19962), .B(n19961), .Z(n20291) );
  NAND U20577 ( .A(a[17]), .B(b[7]), .Z(n20293) );
  AND U20578 ( .A(a[18]), .B(b[7]), .Z(n19967) );
  NANDN U20579 ( .A(n19968), .B(n19967), .Z(n19970) );
  XNOR U20580 ( .A(n19964), .B(n19963), .Z(n19965) );
  XNOR U20581 ( .A(n19966), .B(n19965), .Z(n20199) );
  XNOR U20582 ( .A(n19968), .B(n19967), .Z(n20198) );
  NAND U20583 ( .A(n20199), .B(n20198), .Z(n19969) );
  AND U20584 ( .A(n19970), .B(n19969), .Z(n20298) );
  NAND U20585 ( .A(a[19]), .B(b[7]), .Z(n20301) );
  NANDN U20586 ( .A(n19975), .B(n19976), .Z(n19978) );
  XNOR U20587 ( .A(n19972), .B(n19971), .Z(n19973) );
  XNOR U20588 ( .A(n19974), .B(n19973), .Z(n20197) );
  XNOR U20589 ( .A(n19976), .B(n19975), .Z(n20196) );
  NAND U20590 ( .A(n20197), .B(n20196), .Z(n19977) );
  NAND U20591 ( .A(n19978), .B(n19977), .Z(n20309) );
  AND U20592 ( .A(a[21]), .B(b[7]), .Z(n20311) );
  AND U20593 ( .A(a[22]), .B(b[7]), .Z(n19979) );
  NANDN U20594 ( .A(n19980), .B(n19979), .Z(n19986) );
  XOR U20595 ( .A(n19980), .B(n19979), .Z(n20194) );
  XNOR U20596 ( .A(n19982), .B(n19981), .Z(n19983) );
  XNOR U20597 ( .A(n19984), .B(n19983), .Z(n20195) );
  NANDN U20598 ( .A(n20194), .B(n20195), .Z(n19985) );
  AND U20599 ( .A(n19986), .B(n19985), .Z(n20314) );
  NAND U20600 ( .A(a[23]), .B(b[7]), .Z(n20317) );
  NANDN U20601 ( .A(n19991), .B(n19992), .Z(n19994) );
  XNOR U20602 ( .A(n19988), .B(n19987), .Z(n19989) );
  XNOR U20603 ( .A(n19990), .B(n19989), .Z(n20193) );
  XNOR U20604 ( .A(n19992), .B(n19991), .Z(n20192) );
  NAND U20605 ( .A(n20193), .B(n20192), .Z(n19993) );
  NAND U20606 ( .A(n19994), .B(n19993), .Z(n20323) );
  NAND U20607 ( .A(a[25]), .B(b[7]), .Z(n20325) );
  AND U20608 ( .A(a[26]), .B(b[7]), .Z(n19999) );
  NANDN U20609 ( .A(n20000), .B(n19999), .Z(n20002) );
  XNOR U20610 ( .A(n19996), .B(n19995), .Z(n19997) );
  XNOR U20611 ( .A(n19998), .B(n19997), .Z(n20191) );
  XNOR U20612 ( .A(n20000), .B(n19999), .Z(n20190) );
  NAND U20613 ( .A(n20191), .B(n20190), .Z(n20001) );
  NAND U20614 ( .A(n20002), .B(n20001), .Z(n20331) );
  NAND U20615 ( .A(a[27]), .B(b[7]), .Z(n20333) );
  AND U20616 ( .A(a[28]), .B(b[7]), .Z(n20007) );
  NANDN U20617 ( .A(n20008), .B(n20007), .Z(n20010) );
  XOR U20618 ( .A(n20004), .B(n20003), .Z(n20005) );
  XNOR U20619 ( .A(n20006), .B(n20005), .Z(n20339) );
  XNOR U20620 ( .A(n20008), .B(n20007), .Z(n20338) );
  NAND U20621 ( .A(n20339), .B(n20338), .Z(n20009) );
  NAND U20622 ( .A(n20010), .B(n20009), .Z(n20341) );
  NAND U20623 ( .A(a[29]), .B(b[7]), .Z(n20343) );
  AND U20624 ( .A(a[30]), .B(b[7]), .Z(n20015) );
  NANDN U20625 ( .A(n20016), .B(n20015), .Z(n20018) );
  XNOR U20626 ( .A(n20012), .B(n20011), .Z(n20013) );
  XNOR U20627 ( .A(n20014), .B(n20013), .Z(n20189) );
  XNOR U20628 ( .A(n20016), .B(n20015), .Z(n20188) );
  NAND U20629 ( .A(n20189), .B(n20188), .Z(n20017) );
  NAND U20630 ( .A(n20018), .B(n20017), .Z(n20348) );
  NAND U20631 ( .A(a[31]), .B(b[7]), .Z(n20351) );
  AND U20632 ( .A(a[32]), .B(b[7]), .Z(n20023) );
  NANDN U20633 ( .A(n20024), .B(n20023), .Z(n20026) );
  XOR U20634 ( .A(n20020), .B(n20019), .Z(n20021) );
  XNOR U20635 ( .A(n20022), .B(n20021), .Z(n20357) );
  XNOR U20636 ( .A(n20024), .B(n20023), .Z(n20356) );
  NAND U20637 ( .A(n20357), .B(n20356), .Z(n20025) );
  NAND U20638 ( .A(n20026), .B(n20025), .Z(n20361) );
  NAND U20639 ( .A(a[33]), .B(b[7]), .Z(n20363) );
  AND U20640 ( .A(a[34]), .B(b[7]), .Z(n20031) );
  NANDN U20641 ( .A(n20032), .B(n20031), .Z(n20034) );
  XNOR U20642 ( .A(n20028), .B(n20027), .Z(n20029) );
  XNOR U20643 ( .A(n20030), .B(n20029), .Z(n20187) );
  XNOR U20644 ( .A(n20032), .B(n20031), .Z(n20186) );
  NAND U20645 ( .A(n20187), .B(n20186), .Z(n20033) );
  NAND U20646 ( .A(n20034), .B(n20033), .Z(n20367) );
  NAND U20647 ( .A(a[35]), .B(b[7]), .Z(n20369) );
  AND U20648 ( .A(a[36]), .B(b[7]), .Z(n20039) );
  NANDN U20649 ( .A(n20040), .B(n20039), .Z(n20042) );
  XNOR U20650 ( .A(n20036), .B(n20035), .Z(n20037) );
  XNOR U20651 ( .A(n20038), .B(n20037), .Z(n20185) );
  XNOR U20652 ( .A(n20040), .B(n20039), .Z(n20184) );
  NAND U20653 ( .A(n20185), .B(n20184), .Z(n20041) );
  NAND U20654 ( .A(n20042), .B(n20041), .Z(n20375) );
  NAND U20655 ( .A(a[37]), .B(b[7]), .Z(n20377) );
  AND U20656 ( .A(a[38]), .B(b[7]), .Z(n20047) );
  NANDN U20657 ( .A(n20048), .B(n20047), .Z(n20050) );
  XNOR U20658 ( .A(n20044), .B(n20043), .Z(n20045) );
  XNOR U20659 ( .A(n20046), .B(n20045), .Z(n20183) );
  XNOR U20660 ( .A(n20048), .B(n20047), .Z(n20182) );
  NAND U20661 ( .A(n20183), .B(n20182), .Z(n20049) );
  NAND U20662 ( .A(n20050), .B(n20049), .Z(n20383) );
  NAND U20663 ( .A(a[39]), .B(b[7]), .Z(n20385) );
  AND U20664 ( .A(a[40]), .B(b[7]), .Z(n20055) );
  NANDN U20665 ( .A(n20056), .B(n20055), .Z(n20058) );
  XNOR U20666 ( .A(n20052), .B(n20051), .Z(n20053) );
  XNOR U20667 ( .A(n20054), .B(n20053), .Z(n20181) );
  XNOR U20668 ( .A(n20056), .B(n20055), .Z(n20180) );
  NAND U20669 ( .A(n20181), .B(n20180), .Z(n20057) );
  NAND U20670 ( .A(n20058), .B(n20057), .Z(n20391) );
  NAND U20671 ( .A(a[41]), .B(b[7]), .Z(n20393) );
  AND U20672 ( .A(a[42]), .B(b[7]), .Z(n20063) );
  NANDN U20673 ( .A(n20064), .B(n20063), .Z(n20066) );
  XNOR U20674 ( .A(n20060), .B(n20059), .Z(n20061) );
  XNOR U20675 ( .A(n20062), .B(n20061), .Z(n20179) );
  XNOR U20676 ( .A(n20064), .B(n20063), .Z(n20178) );
  NAND U20677 ( .A(n20179), .B(n20178), .Z(n20065) );
  AND U20678 ( .A(n20066), .B(n20065), .Z(n20398) );
  NAND U20679 ( .A(a[43]), .B(b[7]), .Z(n20401) );
  NANDN U20680 ( .A(n20071), .B(n20072), .Z(n20074) );
  XNOR U20681 ( .A(n20068), .B(n20067), .Z(n20069) );
  XNOR U20682 ( .A(n20070), .B(n20069), .Z(n20407) );
  XNOR U20683 ( .A(n20072), .B(n20071), .Z(n20406) );
  NAND U20684 ( .A(n20407), .B(n20406), .Z(n20073) );
  NAND U20685 ( .A(n20074), .B(n20073), .Z(n20409) );
  NAND U20686 ( .A(a[45]), .B(b[7]), .Z(n20411) );
  AND U20687 ( .A(a[46]), .B(b[7]), .Z(n20079) );
  NANDN U20688 ( .A(n20080), .B(n20079), .Z(n20082) );
  XNOR U20689 ( .A(n20076), .B(n20075), .Z(n20077) );
  XNOR U20690 ( .A(n20078), .B(n20077), .Z(n20177) );
  XNOR U20691 ( .A(n20080), .B(n20079), .Z(n20176) );
  NAND U20692 ( .A(n20177), .B(n20176), .Z(n20081) );
  NAND U20693 ( .A(n20082), .B(n20081), .Z(n20417) );
  NAND U20694 ( .A(a[47]), .B(b[7]), .Z(n20419) );
  XOR U20695 ( .A(n20084), .B(n20083), .Z(n20085) );
  XNOR U20696 ( .A(n20086), .B(n20085), .Z(n20175) );
  NANDN U20697 ( .A(n20426), .B(n20425), .Z(n20090) );
  NOR U20698 ( .A(n20087), .B(n20425), .Z(n20088) );
  AND U20699 ( .A(a[49]), .B(b[7]), .Z(n20424) );
  NANDN U20700 ( .A(n20088), .B(n20424), .Z(n20089) );
  AND U20701 ( .A(n20090), .B(n20089), .Z(n20169) );
  NANDN U20702 ( .A(n20432), .B(n20433), .Z(n20097) );
  NOR U20703 ( .A(n20094), .B(n20433), .Z(n20095) );
  AND U20704 ( .A(a[51]), .B(b[7]), .Z(n20431) );
  NANDN U20705 ( .A(n20095), .B(n20431), .Z(n20096) );
  AND U20706 ( .A(n20097), .B(n20096), .Z(n20099) );
  AND U20707 ( .A(a[52]), .B(b[7]), .Z(n20098) );
  NANDN U20708 ( .A(n20099), .B(n20098), .Z(n20105) );
  XNOR U20709 ( .A(n20099), .B(n20098), .Z(n20167) );
  XNOR U20710 ( .A(n20101), .B(n20100), .Z(n20102) );
  XNOR U20711 ( .A(n20103), .B(n20102), .Z(n20166) );
  NAND U20712 ( .A(n20167), .B(n20166), .Z(n20104) );
  NAND U20713 ( .A(n20105), .B(n20104), .Z(n20441) );
  NAND U20714 ( .A(a[53]), .B(b[7]), .Z(n20443) );
  AND U20715 ( .A(a[54]), .B(b[7]), .Z(n20110) );
  NANDN U20716 ( .A(n20111), .B(n20110), .Z(n20113) );
  XNOR U20717 ( .A(n20107), .B(n20106), .Z(n20108) );
  XNOR U20718 ( .A(n20109), .B(n20108), .Z(n20165) );
  XNOR U20719 ( .A(n20111), .B(n20110), .Z(n20164) );
  NAND U20720 ( .A(n20165), .B(n20164), .Z(n20112) );
  AND U20721 ( .A(n20113), .B(n20112), .Z(n20446) );
  AND U20722 ( .A(a[55]), .B(b[7]), .Z(n20449) );
  NANDN U20723 ( .A(n20117), .B(n20118), .Z(n20120) );
  NAND U20724 ( .A(n20163), .B(n20162), .Z(n20119) );
  AND U20725 ( .A(n20120), .B(n20119), .Z(n20124) );
  NAND U20726 ( .A(n20124), .B(n20123), .Z(n20126) );
  XOR U20727 ( .A(n20124), .B(n20123), .Z(n20455) );
  NAND U20728 ( .A(a[57]), .B(b[7]), .Z(n20454) );
  NAND U20729 ( .A(n20455), .B(n20454), .Z(n20125) );
  NAND U20730 ( .A(n20126), .B(n20125), .Z(n20463) );
  XOR U20731 ( .A(n20128), .B(n20127), .Z(n20157) );
  XOR U20732 ( .A(n20130), .B(n20129), .Z(n20468) );
  XOR U20733 ( .A(n20132), .B(n20131), .Z(n20469) );
  XOR U20734 ( .A(n20134), .B(n20133), .Z(n20153) );
  XOR U20735 ( .A(n20136), .B(n20135), .Z(n20152) );
  XOR U20736 ( .A(n20138), .B(n20137), .Z(n20472) );
  XOR U20737 ( .A(n20140), .B(n20139), .Z(n20473) );
  XOR U20738 ( .A(n20142), .B(n20141), .Z(n20477) );
  XOR U20739 ( .A(n20144), .B(n20143), .Z(n20476) );
  XOR U20740 ( .A(n20146), .B(n20145), .Z(n20478) );
  NANDN U20741 ( .A(n24683), .B(n24684), .Z(n24692) );
  NAND U20742 ( .A(n20148), .B(n20147), .Z(n24694) );
  XOR U20743 ( .A(n20150), .B(n20149), .Z(n24693) );
  NANDN U20744 ( .A(n24694), .B(n24693), .Z(n20151) );
  NAND U20745 ( .A(n24692), .B(n20151), .Z(n22500) );
  NANDN U20746 ( .A(n24684), .B(n24683), .Z(n20481) );
  AND U20747 ( .A(a[62]), .B(b[6]), .Z(n20154) );
  XOR U20748 ( .A(n20153), .B(n20152), .Z(n20155) );
  XNOR U20749 ( .A(n20155), .B(n20154), .Z(n20810) );
  XNOR U20750 ( .A(n20157), .B(n20156), .Z(n20158) );
  XOR U20751 ( .A(n20159), .B(n20158), .Z(n20161) );
  AND U20752 ( .A(a[60]), .B(b[6]), .Z(n20160) );
  NAND U20753 ( .A(n20161), .B(n20160), .Z(n20467) );
  XNOR U20754 ( .A(n20161), .B(n20160), .Z(n20799) );
  AND U20755 ( .A(a[59]), .B(b[6]), .Z(n20460) );
  XNOR U20756 ( .A(n20163), .B(n20162), .Z(n20784) );
  XNOR U20757 ( .A(n20165), .B(n20164), .Z(n20778) );
  XOR U20758 ( .A(n20167), .B(n20166), .Z(n20434) );
  IV U20759 ( .A(n20434), .Z(n20763) );
  NAND U20760 ( .A(a[52]), .B(b[6]), .Z(n20759) );
  XOR U20761 ( .A(n20169), .B(n20168), .Z(n20170) );
  XOR U20762 ( .A(n20171), .B(n20170), .Z(n20427) );
  IV U20763 ( .A(n20427), .Z(n20757) );
  NAND U20764 ( .A(a[50]), .B(b[6]), .Z(n20490) );
  XOR U20765 ( .A(n20173), .B(n20172), .Z(n20174) );
  XNOR U20766 ( .A(n20175), .B(n20174), .Z(n20749) );
  XNOR U20767 ( .A(n20177), .B(n20176), .Z(n20739) );
  XNOR U20768 ( .A(n20179), .B(n20178), .Z(n20723) );
  XNOR U20769 ( .A(n20181), .B(n20180), .Z(n20715) );
  XNOR U20770 ( .A(n20183), .B(n20182), .Z(n20707) );
  XNOR U20771 ( .A(n20185), .B(n20184), .Z(n20699) );
  XNOR U20772 ( .A(n20187), .B(n20186), .Z(n20691) );
  AND U20773 ( .A(a[32]), .B(b[6]), .Z(n20353) );
  XNOR U20774 ( .A(n20189), .B(n20188), .Z(n20675) );
  AND U20775 ( .A(a[28]), .B(b[6]), .Z(n20335) );
  XNOR U20776 ( .A(n20191), .B(n20190), .Z(n20659) );
  XNOR U20777 ( .A(n20193), .B(n20192), .Z(n20651) );
  NAND U20778 ( .A(a[24]), .B(b[6]), .Z(n20318) );
  XNOR U20779 ( .A(n20195), .B(n20194), .Z(n20644) );
  AND U20780 ( .A(a[22]), .B(b[6]), .Z(n20307) );
  XNOR U20781 ( .A(n20197), .B(n20196), .Z(n20635) );
  XNOR U20782 ( .A(n20199), .B(n20198), .Z(n20627) );
  XNOR U20783 ( .A(n20201), .B(n20200), .Z(n20619) );
  AND U20784 ( .A(a[10]), .B(b[6]), .Z(n20251) );
  XNOR U20785 ( .A(n20203), .B(n20202), .Z(n20236) );
  XOR U20786 ( .A(n20205), .B(n20204), .Z(n20233) );
  NAND U20787 ( .A(a[5]), .B(b[6]), .Z(n20228) );
  XOR U20788 ( .A(n20207), .B(n20206), .Z(n20229) );
  NANDN U20789 ( .A(n20228), .B(n20229), .Z(n20231) );
  AND U20790 ( .A(a[0]), .B(b[6]), .Z(n20868) );
  AND U20791 ( .A(a[1]), .B(b[7]), .Z(n20211) );
  AND U20792 ( .A(n20868), .B(n20211), .Z(n20208) );
  NAND U20793 ( .A(a[2]), .B(n20208), .Z(n20215) );
  NAND U20794 ( .A(b[7]), .B(a[1]), .Z(n20209) );
  XOR U20795 ( .A(n20210), .B(n20209), .Z(n20537) );
  NAND U20796 ( .A(n20211), .B(a[0]), .Z(n20212) );
  XNOR U20797 ( .A(a[2]), .B(n20212), .Z(n20213) );
  AND U20798 ( .A(b[6]), .B(n20213), .Z(n20538) );
  NANDN U20799 ( .A(n20537), .B(n20538), .Z(n20214) );
  AND U20800 ( .A(n20215), .B(n20214), .Z(n20218) );
  NANDN U20801 ( .A(n20218), .B(n20219), .Z(n20221) );
  AND U20802 ( .A(a[3]), .B(b[6]), .Z(n20543) );
  NAND U20803 ( .A(n20544), .B(n20543), .Z(n20220) );
  AND U20804 ( .A(n20221), .B(n20220), .Z(n20224) );
  AND U20805 ( .A(a[4]), .B(b[6]), .Z(n20225) );
  NANDN U20806 ( .A(n20224), .B(n20225), .Z(n20227) );
  NAND U20807 ( .A(n20550), .B(n20549), .Z(n20226) );
  AND U20808 ( .A(n20227), .B(n20226), .Z(n20555) );
  NANDN U20809 ( .A(n20555), .B(n20556), .Z(n20230) );
  AND U20810 ( .A(n20231), .B(n20230), .Z(n20232) );
  NANDN U20811 ( .A(n20233), .B(n20232), .Z(n20235) );
  XOR U20812 ( .A(n20233), .B(n20232), .Z(n20527) );
  AND U20813 ( .A(a[6]), .B(b[6]), .Z(n20528) );
  OR U20814 ( .A(n20527), .B(n20528), .Z(n20234) );
  AND U20815 ( .A(n20235), .B(n20234), .Z(n20237) );
  NAND U20816 ( .A(a[7]), .B(b[6]), .Z(n20567) );
  XOR U20817 ( .A(n20237), .B(n20236), .Z(n20568) );
  AND U20818 ( .A(a[8]), .B(b[6]), .Z(n20240) );
  XNOR U20819 ( .A(n20239), .B(n20238), .Z(n20571) );
  XNOR U20820 ( .A(n20241), .B(n20240), .Z(n20572) );
  XOR U20821 ( .A(n20243), .B(n20242), .Z(n20244) );
  NANDN U20822 ( .A(n20245), .B(n20244), .Z(n20247) );
  NAND U20823 ( .A(a[9]), .B(b[6]), .Z(n20577) );
  XNOR U20824 ( .A(n20245), .B(n20244), .Z(n20578) );
  NANDN U20825 ( .A(n20577), .B(n20578), .Z(n20246) );
  AND U20826 ( .A(n20247), .B(n20246), .Z(n20250) );
  NANDN U20827 ( .A(n20251), .B(n20250), .Z(n20253) );
  XOR U20828 ( .A(n20249), .B(n20248), .Z(n20584) );
  XNOR U20829 ( .A(n20251), .B(n20250), .Z(n20583) );
  NANDN U20830 ( .A(n20584), .B(n20583), .Z(n20252) );
  AND U20831 ( .A(n20253), .B(n20252), .Z(n20257) );
  XOR U20832 ( .A(n20255), .B(n20254), .Z(n20256) );
  NAND U20833 ( .A(n20257), .B(n20256), .Z(n20259) );
  NAND U20834 ( .A(a[11]), .B(b[6]), .Z(n20589) );
  XOR U20835 ( .A(n20257), .B(n20256), .Z(n20590) );
  NANDN U20836 ( .A(n20589), .B(n20590), .Z(n20258) );
  AND U20837 ( .A(n20259), .B(n20258), .Z(n20261) );
  AND U20838 ( .A(a[12]), .B(b[6]), .Z(n20260) );
  NANDN U20839 ( .A(n20261), .B(n20260), .Z(n20265) );
  XNOR U20840 ( .A(n20261), .B(n20260), .Z(n20596) );
  XNOR U20841 ( .A(n20263), .B(n20262), .Z(n20595) );
  NAND U20842 ( .A(n20596), .B(n20595), .Z(n20264) );
  AND U20843 ( .A(n20265), .B(n20264), .Z(n20269) );
  XOR U20844 ( .A(n20267), .B(n20266), .Z(n20268) );
  NANDN U20845 ( .A(n20269), .B(n20268), .Z(n20271) );
  NAND U20846 ( .A(a[13]), .B(b[6]), .Z(n20601) );
  XNOR U20847 ( .A(n20269), .B(n20268), .Z(n20602) );
  NANDN U20848 ( .A(n20601), .B(n20602), .Z(n20270) );
  AND U20849 ( .A(n20271), .B(n20270), .Z(n20273) );
  AND U20850 ( .A(a[14]), .B(b[6]), .Z(n20272) );
  NANDN U20851 ( .A(n20273), .B(n20272), .Z(n20277) );
  XNOR U20852 ( .A(n20273), .B(n20272), .Z(n20608) );
  XNOR U20853 ( .A(n20275), .B(n20274), .Z(n20607) );
  NAND U20854 ( .A(n20608), .B(n20607), .Z(n20276) );
  AND U20855 ( .A(n20277), .B(n20276), .Z(n20281) );
  XOR U20856 ( .A(n20279), .B(n20278), .Z(n20280) );
  NANDN U20857 ( .A(n20281), .B(n20280), .Z(n20283) );
  NAND U20858 ( .A(a[15]), .B(b[6]), .Z(n20613) );
  XNOR U20859 ( .A(n20281), .B(n20280), .Z(n20614) );
  NANDN U20860 ( .A(n20613), .B(n20614), .Z(n20282) );
  AND U20861 ( .A(n20283), .B(n20282), .Z(n20285) );
  AND U20862 ( .A(a[16]), .B(b[6]), .Z(n20284) );
  NANDN U20863 ( .A(n20285), .B(n20284), .Z(n20289) );
  XNOR U20864 ( .A(n20285), .B(n20284), .Z(n20526) );
  XNOR U20865 ( .A(n20287), .B(n20286), .Z(n20525) );
  NAND U20866 ( .A(n20526), .B(n20525), .Z(n20288) );
  NAND U20867 ( .A(n20289), .B(n20288), .Z(n20620) );
  NAND U20868 ( .A(a[17]), .B(b[6]), .Z(n20622) );
  AND U20869 ( .A(a[18]), .B(b[6]), .Z(n20294) );
  NANDN U20870 ( .A(n20295), .B(n20294), .Z(n20297) );
  XNOR U20871 ( .A(n20291), .B(n20290), .Z(n20292) );
  XNOR U20872 ( .A(n20293), .B(n20292), .Z(n20524) );
  XNOR U20873 ( .A(n20295), .B(n20294), .Z(n20523) );
  NAND U20874 ( .A(n20524), .B(n20523), .Z(n20296) );
  NAND U20875 ( .A(n20297), .B(n20296), .Z(n20628) );
  NAND U20876 ( .A(a[19]), .B(b[6]), .Z(n20630) );
  AND U20877 ( .A(a[20]), .B(b[6]), .Z(n20302) );
  NANDN U20878 ( .A(n20303), .B(n20302), .Z(n20305) );
  XNOR U20879 ( .A(n20299), .B(n20298), .Z(n20300) );
  XNOR U20880 ( .A(n20301), .B(n20300), .Z(n20522) );
  XNOR U20881 ( .A(n20303), .B(n20302), .Z(n20521) );
  NAND U20882 ( .A(n20522), .B(n20521), .Z(n20304) );
  NAND U20883 ( .A(n20305), .B(n20304), .Z(n20636) );
  NAND U20884 ( .A(a[21]), .B(b[6]), .Z(n20638) );
  NANDN U20885 ( .A(n20307), .B(n20306), .Z(n20313) );
  XNOR U20886 ( .A(n20307), .B(n20306), .Z(n20519) );
  XNOR U20887 ( .A(n20309), .B(n20308), .Z(n20310) );
  XNOR U20888 ( .A(n20311), .B(n20310), .Z(n20520) );
  NAND U20889 ( .A(n20519), .B(n20520), .Z(n20312) );
  NAND U20890 ( .A(n20313), .B(n20312), .Z(n20643) );
  AND U20891 ( .A(a[23]), .B(b[6]), .Z(n20646) );
  NANDN U20892 ( .A(n20318), .B(n20319), .Z(n20321) );
  XNOR U20893 ( .A(n20315), .B(n20314), .Z(n20316) );
  XNOR U20894 ( .A(n20317), .B(n20316), .Z(n20518) );
  XNOR U20895 ( .A(n20319), .B(n20318), .Z(n20517) );
  NAND U20896 ( .A(n20518), .B(n20517), .Z(n20320) );
  NAND U20897 ( .A(n20321), .B(n20320), .Z(n20652) );
  NAND U20898 ( .A(a[25]), .B(b[6]), .Z(n20654) );
  AND U20899 ( .A(a[26]), .B(b[6]), .Z(n20326) );
  NANDN U20900 ( .A(n20327), .B(n20326), .Z(n20329) );
  XNOR U20901 ( .A(n20323), .B(n20322), .Z(n20324) );
  XNOR U20902 ( .A(n20325), .B(n20324), .Z(n20516) );
  XNOR U20903 ( .A(n20327), .B(n20326), .Z(n20515) );
  NAND U20904 ( .A(n20516), .B(n20515), .Z(n20328) );
  NAND U20905 ( .A(n20329), .B(n20328), .Z(n20660) );
  NAND U20906 ( .A(a[27]), .B(b[6]), .Z(n20662) );
  NANDN U20907 ( .A(n20335), .B(n20334), .Z(n20337) );
  XOR U20908 ( .A(n20331), .B(n20330), .Z(n20332) );
  XOR U20909 ( .A(n20333), .B(n20332), .Z(n20514) );
  XNOR U20910 ( .A(n20335), .B(n20334), .Z(n20513) );
  NANDN U20911 ( .A(n20514), .B(n20513), .Z(n20336) );
  NAND U20912 ( .A(n20337), .B(n20336), .Z(n20668) );
  XOR U20913 ( .A(n20339), .B(n20338), .Z(n20667) );
  AND U20914 ( .A(a[29]), .B(b[6]), .Z(n20670) );
  AND U20915 ( .A(a[30]), .B(b[6]), .Z(n20344) );
  NANDN U20916 ( .A(n20345), .B(n20344), .Z(n20347) );
  XNOR U20917 ( .A(n20341), .B(n20340), .Z(n20342) );
  XNOR U20918 ( .A(n20343), .B(n20342), .Z(n20512) );
  XNOR U20919 ( .A(n20345), .B(n20344), .Z(n20511) );
  NAND U20920 ( .A(n20512), .B(n20511), .Z(n20346) );
  NAND U20921 ( .A(n20347), .B(n20346), .Z(n20676) );
  NAND U20922 ( .A(a[31]), .B(b[6]), .Z(n20678) );
  NANDN U20923 ( .A(n20353), .B(n20352), .Z(n20355) );
  XOR U20924 ( .A(n20349), .B(n20348), .Z(n20350) );
  XOR U20925 ( .A(n20351), .B(n20350), .Z(n20510) );
  XNOR U20926 ( .A(n20353), .B(n20352), .Z(n20509) );
  NANDN U20927 ( .A(n20510), .B(n20509), .Z(n20354) );
  NAND U20928 ( .A(n20355), .B(n20354), .Z(n20686) );
  XOR U20929 ( .A(n20357), .B(n20356), .Z(n20685) );
  AND U20930 ( .A(a[33]), .B(b[6]), .Z(n20688) );
  AND U20931 ( .A(a[34]), .B(b[6]), .Z(n20358) );
  NANDN U20932 ( .A(n20359), .B(n20358), .Z(n20365) );
  XOR U20933 ( .A(n20359), .B(n20358), .Z(n20507) );
  XNOR U20934 ( .A(n20361), .B(n20360), .Z(n20362) );
  XNOR U20935 ( .A(n20363), .B(n20362), .Z(n20508) );
  NANDN U20936 ( .A(n20507), .B(n20508), .Z(n20364) );
  NAND U20937 ( .A(n20365), .B(n20364), .Z(n20692) );
  NAND U20938 ( .A(a[35]), .B(b[6]), .Z(n20694) );
  AND U20939 ( .A(a[36]), .B(b[6]), .Z(n20370) );
  NANDN U20940 ( .A(n20371), .B(n20370), .Z(n20373) );
  XNOR U20941 ( .A(n20367), .B(n20366), .Z(n20368) );
  XNOR U20942 ( .A(n20369), .B(n20368), .Z(n20506) );
  XNOR U20943 ( .A(n20371), .B(n20370), .Z(n20505) );
  NAND U20944 ( .A(n20506), .B(n20505), .Z(n20372) );
  NAND U20945 ( .A(n20373), .B(n20372), .Z(n20700) );
  NAND U20946 ( .A(a[37]), .B(b[6]), .Z(n20702) );
  AND U20947 ( .A(a[38]), .B(b[6]), .Z(n20378) );
  NANDN U20948 ( .A(n20379), .B(n20378), .Z(n20381) );
  XNOR U20949 ( .A(n20375), .B(n20374), .Z(n20376) );
  XNOR U20950 ( .A(n20377), .B(n20376), .Z(n20504) );
  XNOR U20951 ( .A(n20379), .B(n20378), .Z(n20503) );
  NAND U20952 ( .A(n20504), .B(n20503), .Z(n20380) );
  NAND U20953 ( .A(n20381), .B(n20380), .Z(n20708) );
  NAND U20954 ( .A(a[39]), .B(b[6]), .Z(n20710) );
  AND U20955 ( .A(a[40]), .B(b[6]), .Z(n20386) );
  NANDN U20956 ( .A(n20387), .B(n20386), .Z(n20389) );
  XNOR U20957 ( .A(n20383), .B(n20382), .Z(n20384) );
  XNOR U20958 ( .A(n20385), .B(n20384), .Z(n20502) );
  XNOR U20959 ( .A(n20387), .B(n20386), .Z(n20501) );
  NAND U20960 ( .A(n20502), .B(n20501), .Z(n20388) );
  NAND U20961 ( .A(n20389), .B(n20388), .Z(n20716) );
  NAND U20962 ( .A(a[41]), .B(b[6]), .Z(n20718) );
  AND U20963 ( .A(a[42]), .B(b[6]), .Z(n20394) );
  NANDN U20964 ( .A(n20395), .B(n20394), .Z(n20397) );
  XNOR U20965 ( .A(n20391), .B(n20390), .Z(n20392) );
  XNOR U20966 ( .A(n20393), .B(n20392), .Z(n20500) );
  XNOR U20967 ( .A(n20395), .B(n20394), .Z(n20499) );
  NAND U20968 ( .A(n20500), .B(n20499), .Z(n20396) );
  NAND U20969 ( .A(n20397), .B(n20396), .Z(n20724) );
  NAND U20970 ( .A(a[43]), .B(b[6]), .Z(n20726) );
  AND U20971 ( .A(a[44]), .B(b[6]), .Z(n20402) );
  NANDN U20972 ( .A(n20403), .B(n20402), .Z(n20405) );
  XNOR U20973 ( .A(n20399), .B(n20398), .Z(n20400) );
  XNOR U20974 ( .A(n20401), .B(n20400), .Z(n20498) );
  XNOR U20975 ( .A(n20403), .B(n20402), .Z(n20497) );
  NAND U20976 ( .A(n20498), .B(n20497), .Z(n20404) );
  AND U20977 ( .A(n20405), .B(n20404), .Z(n20732) );
  XOR U20978 ( .A(n20407), .B(n20406), .Z(n20731) );
  NAND U20979 ( .A(a[45]), .B(b[6]), .Z(n20734) );
  AND U20980 ( .A(a[46]), .B(b[6]), .Z(n20412) );
  NANDN U20981 ( .A(n20413), .B(n20412), .Z(n20415) );
  XNOR U20982 ( .A(n20409), .B(n20408), .Z(n20410) );
  XNOR U20983 ( .A(n20411), .B(n20410), .Z(n20496) );
  XNOR U20984 ( .A(n20413), .B(n20412), .Z(n20495) );
  NAND U20985 ( .A(n20496), .B(n20495), .Z(n20414) );
  NAND U20986 ( .A(n20415), .B(n20414), .Z(n20740) );
  NAND U20987 ( .A(a[47]), .B(b[6]), .Z(n20742) );
  AND U20988 ( .A(a[48]), .B(b[6]), .Z(n20420) );
  NANDN U20989 ( .A(n20421), .B(n20420), .Z(n20423) );
  XNOR U20990 ( .A(n20417), .B(n20416), .Z(n20418) );
  XNOR U20991 ( .A(n20419), .B(n20418), .Z(n20494) );
  XNOR U20992 ( .A(n20421), .B(n20420), .Z(n20493) );
  NAND U20993 ( .A(n20494), .B(n20493), .Z(n20422) );
  NAND U20994 ( .A(n20423), .B(n20422), .Z(n20750) );
  NAND U20995 ( .A(a[49]), .B(b[6]), .Z(n20752) );
  NANDN U20996 ( .A(n20757), .B(n20756), .Z(n20430) );
  NOR U20997 ( .A(n20427), .B(n20756), .Z(n20428) );
  AND U20998 ( .A(a[51]), .B(b[6]), .Z(n20755) );
  NANDN U20999 ( .A(n20428), .B(n20755), .Z(n20429) );
  AND U21000 ( .A(n20430), .B(n20429), .Z(n20758) );
  NANDN U21001 ( .A(n20763), .B(n20764), .Z(n20437) );
  NOR U21002 ( .A(n20434), .B(n20764), .Z(n20435) );
  NAND U21003 ( .A(a[53]), .B(b[6]), .Z(n20766) );
  OR U21004 ( .A(n20435), .B(n20766), .Z(n20436) );
  AND U21005 ( .A(n20437), .B(n20436), .Z(n20438) );
  AND U21006 ( .A(a[54]), .B(b[6]), .Z(n20439) );
  NANDN U21007 ( .A(n20438), .B(n20439), .Z(n20445) );
  XNOR U21008 ( .A(n20439), .B(n20438), .Z(n20771) );
  XNOR U21009 ( .A(n20441), .B(n20440), .Z(n20442) );
  XNOR U21010 ( .A(n20443), .B(n20442), .Z(n20770) );
  NAND U21011 ( .A(n20771), .B(n20770), .Z(n20444) );
  NAND U21012 ( .A(n20445), .B(n20444), .Z(n20779) );
  NAND U21013 ( .A(a[55]), .B(b[6]), .Z(n20781) );
  AND U21014 ( .A(a[56]), .B(b[6]), .Z(n20451) );
  NANDN U21015 ( .A(n20450), .B(n20451), .Z(n20453) );
  XOR U21016 ( .A(n20447), .B(n20446), .Z(n20448) );
  XNOR U21017 ( .A(n20449), .B(n20448), .Z(n20488) );
  XNOR U21018 ( .A(n20451), .B(n20450), .Z(n20487) );
  NAND U21019 ( .A(n20488), .B(n20487), .Z(n20452) );
  NAND U21020 ( .A(n20453), .B(n20452), .Z(n20785) );
  NAND U21021 ( .A(a[57]), .B(b[6]), .Z(n20787) );
  AND U21022 ( .A(a[58]), .B(b[6]), .Z(n20456) );
  NANDN U21023 ( .A(n20457), .B(n20456), .Z(n20459) );
  XOR U21024 ( .A(n20455), .B(n20454), .Z(n20792) );
  XNOR U21025 ( .A(n20457), .B(n20456), .Z(n20793) );
  NANDN U21026 ( .A(n20792), .B(n20793), .Z(n20458) );
  NAND U21027 ( .A(n20459), .B(n20458), .Z(n20461) );
  XNOR U21028 ( .A(n20461), .B(n20460), .Z(n20485) );
  XOR U21029 ( .A(n20463), .B(n20462), .Z(n20464) );
  XOR U21030 ( .A(n20465), .B(n20464), .Z(n20486) );
  NANDN U21031 ( .A(n20799), .B(n20800), .Z(n20466) );
  NAND U21032 ( .A(n20467), .B(n20466), .Z(n20471) );
  XOR U21033 ( .A(n20469), .B(n20468), .Z(n20470) );
  AND U21034 ( .A(a[61]), .B(b[6]), .Z(n20804) );
  XOR U21035 ( .A(n20471), .B(n20470), .Z(n20805) );
  XOR U21036 ( .A(n20473), .B(n20472), .Z(n20474) );
  AND U21037 ( .A(a[63]), .B(b[6]), .Z(n20814) );
  XOR U21038 ( .A(n20475), .B(n20474), .Z(n20815) );
  XOR U21039 ( .A(n20477), .B(n20476), .Z(n20484) );
  XOR U21040 ( .A(n20479), .B(n20478), .Z(n24681) );
  IV U21041 ( .A(n24681), .Z(n20482) );
  NANDN U21042 ( .A(n24682), .B(n20482), .Z(n20480) );
  AND U21043 ( .A(n20481), .B(n20480), .Z(n22498) );
  ANDN U21044 ( .B(n24682), .A(n20482), .Z(n24688) );
  XNOR U21045 ( .A(n20484), .B(n20483), .Z(n24677) );
  AND U21046 ( .A(a[63]), .B(b[5]), .Z(n20809) );
  AND U21047 ( .A(a[61]), .B(b[5]), .Z(n20798) );
  IV U21048 ( .A(n20798), .Z(n20818) );
  AND U21049 ( .A(a[60]), .B(b[5]), .Z(n21139) );
  XOR U21050 ( .A(n20486), .B(n20485), .Z(n21138) );
  XNOR U21051 ( .A(n20488), .B(n20487), .Z(n21126) );
  AND U21052 ( .A(a[54]), .B(b[5]), .Z(n20762) );
  IV U21053 ( .A(n20762), .Z(n21108) );
  NAND U21054 ( .A(a[52]), .B(b[5]), .Z(n20826) );
  XOR U21055 ( .A(n20490), .B(n20489), .Z(n20491) );
  XNOR U21056 ( .A(n20492), .B(n20491), .Z(n21092) );
  XNOR U21057 ( .A(n20494), .B(n20493), .Z(n21084) );
  XNOR U21058 ( .A(n20496), .B(n20495), .Z(n21076) );
  XNOR U21059 ( .A(n20498), .B(n20497), .Z(n21070) );
  XNOR U21060 ( .A(n20500), .B(n20499), .Z(n21060) );
  XNOR U21061 ( .A(n20502), .B(n20501), .Z(n21052) );
  XNOR U21062 ( .A(n20504), .B(n20503), .Z(n21044) );
  XNOR U21063 ( .A(n20506), .B(n20505), .Z(n21036) );
  NAND U21064 ( .A(a[36]), .B(b[5]), .Z(n20695) );
  XNOR U21065 ( .A(n20508), .B(n20507), .Z(n21029) );
  XNOR U21066 ( .A(n20510), .B(n20509), .Z(n21020) );
  XNOR U21067 ( .A(n20512), .B(n20511), .Z(n21012) );
  NAND U21068 ( .A(a[30]), .B(b[5]), .Z(n20671) );
  XOR U21069 ( .A(n20514), .B(n20513), .Z(n21003) );
  XNOR U21070 ( .A(n20516), .B(n20515), .Z(n20994) );
  XNOR U21071 ( .A(n20518), .B(n20517), .Z(n20986) );
  XOR U21072 ( .A(n20520), .B(n20519), .Z(n20977) );
  XNOR U21073 ( .A(n20522), .B(n20521), .Z(n20968) );
  XNOR U21074 ( .A(n20524), .B(n20523), .Z(n20960) );
  XNOR U21075 ( .A(n20526), .B(n20525), .Z(n20952) );
  XOR U21076 ( .A(n20528), .B(n20527), .Z(n20562) );
  AND U21077 ( .A(a[4]), .B(b[5]), .Z(n20545) );
  AND U21078 ( .A(a[0]), .B(b[5]), .Z(n21200) );
  AND U21079 ( .A(a[1]), .B(b[6]), .Z(n20532) );
  AND U21080 ( .A(n21200), .B(n20532), .Z(n20529) );
  NAND U21081 ( .A(a[2]), .B(n20529), .Z(n20536) );
  NAND U21082 ( .A(b[6]), .B(a[1]), .Z(n20530) );
  XOR U21083 ( .A(n20531), .B(n20530), .Z(n20874) );
  NAND U21084 ( .A(n20532), .B(a[0]), .Z(n20533) );
  XNOR U21085 ( .A(a[2]), .B(n20533), .Z(n20534) );
  AND U21086 ( .A(b[5]), .B(n20534), .Z(n20875) );
  NANDN U21087 ( .A(n20874), .B(n20875), .Z(n20535) );
  AND U21088 ( .A(n20536), .B(n20535), .Z(n20539) );
  NANDN U21089 ( .A(n20539), .B(n20540), .Z(n20542) );
  NAND U21090 ( .A(a[3]), .B(b[5]), .Z(n20882) );
  NANDN U21091 ( .A(n20882), .B(n20883), .Z(n20541) );
  AND U21092 ( .A(n20542), .B(n20541), .Z(n20546) );
  NANDN U21093 ( .A(n20545), .B(n20546), .Z(n20548) );
  XOR U21094 ( .A(n20544), .B(n20543), .Z(n20864) );
  NANDN U21095 ( .A(n20864), .B(n20865), .Z(n20547) );
  AND U21096 ( .A(n20548), .B(n20547), .Z(n20552) );
  XOR U21097 ( .A(n20550), .B(n20549), .Z(n20551) );
  NAND U21098 ( .A(n20552), .B(n20551), .Z(n20554) );
  NAND U21099 ( .A(a[5]), .B(b[5]), .Z(n20890) );
  XOR U21100 ( .A(n20552), .B(n20551), .Z(n20891) );
  NANDN U21101 ( .A(n20890), .B(n20891), .Z(n20553) );
  AND U21102 ( .A(n20554), .B(n20553), .Z(n20557) );
  NANDN U21103 ( .A(n20557), .B(n20558), .Z(n20560) );
  AND U21104 ( .A(a[6]), .B(b[5]), .Z(n20897) );
  NAND U21105 ( .A(n20897), .B(n20896), .Z(n20559) );
  NAND U21106 ( .A(n20560), .B(n20559), .Z(n20561) );
  NANDN U21107 ( .A(n20562), .B(n20561), .Z(n20564) );
  XNOR U21108 ( .A(n20562), .B(n20561), .Z(n20905) );
  AND U21109 ( .A(a[7]), .B(b[5]), .Z(n20904) );
  NAND U21110 ( .A(n20905), .B(n20904), .Z(n20563) );
  AND U21111 ( .A(n20564), .B(n20563), .Z(n20566) );
  AND U21112 ( .A(a[8]), .B(b[5]), .Z(n20565) );
  NANDN U21113 ( .A(n20566), .B(n20565), .Z(n20570) );
  XOR U21114 ( .A(n20566), .B(n20565), .Z(n20862) );
  XNOR U21115 ( .A(n20568), .B(n20567), .Z(n20863) );
  NANDN U21116 ( .A(n20862), .B(n20863), .Z(n20569) );
  AND U21117 ( .A(n20570), .B(n20569), .Z(n20574) );
  XOR U21118 ( .A(n20572), .B(n20571), .Z(n20573) );
  NANDN U21119 ( .A(n20574), .B(n20573), .Z(n20576) );
  NAND U21120 ( .A(a[9]), .B(b[5]), .Z(n20912) );
  XNOR U21121 ( .A(n20574), .B(n20573), .Z(n20913) );
  NANDN U21122 ( .A(n20912), .B(n20913), .Z(n20575) );
  AND U21123 ( .A(n20576), .B(n20575), .Z(n20580) );
  AND U21124 ( .A(a[10]), .B(b[5]), .Z(n20579) );
  NANDN U21125 ( .A(n20580), .B(n20579), .Z(n20582) );
  XNOR U21126 ( .A(n20578), .B(n20577), .Z(n20919) );
  XNOR U21127 ( .A(n20580), .B(n20579), .Z(n20918) );
  NAND U21128 ( .A(n20919), .B(n20918), .Z(n20581) );
  AND U21129 ( .A(n20582), .B(n20581), .Z(n20586) );
  XOR U21130 ( .A(n20584), .B(n20583), .Z(n20585) );
  NANDN U21131 ( .A(n20586), .B(n20585), .Z(n20588) );
  NAND U21132 ( .A(a[11]), .B(b[5]), .Z(n20924) );
  XNOR U21133 ( .A(n20586), .B(n20585), .Z(n20925) );
  NANDN U21134 ( .A(n20924), .B(n20925), .Z(n20587) );
  AND U21135 ( .A(n20588), .B(n20587), .Z(n20592) );
  AND U21136 ( .A(a[12]), .B(b[5]), .Z(n20591) );
  NANDN U21137 ( .A(n20592), .B(n20591), .Z(n20594) );
  XNOR U21138 ( .A(n20590), .B(n20589), .Z(n20929) );
  XNOR U21139 ( .A(n20592), .B(n20591), .Z(n20928) );
  NAND U21140 ( .A(n20929), .B(n20928), .Z(n20593) );
  AND U21141 ( .A(n20594), .B(n20593), .Z(n20598) );
  XOR U21142 ( .A(n20596), .B(n20595), .Z(n20597) );
  NANDN U21143 ( .A(n20598), .B(n20597), .Z(n20600) );
  NAND U21144 ( .A(a[13]), .B(b[5]), .Z(n20936) );
  XNOR U21145 ( .A(n20598), .B(n20597), .Z(n20937) );
  NANDN U21146 ( .A(n20936), .B(n20937), .Z(n20599) );
  AND U21147 ( .A(n20600), .B(n20599), .Z(n20604) );
  AND U21148 ( .A(a[14]), .B(b[5]), .Z(n20603) );
  NANDN U21149 ( .A(n20604), .B(n20603), .Z(n20606) );
  XNOR U21150 ( .A(n20602), .B(n20601), .Z(n20941) );
  XNOR U21151 ( .A(n20604), .B(n20603), .Z(n20940) );
  NAND U21152 ( .A(n20941), .B(n20940), .Z(n20605) );
  AND U21153 ( .A(n20606), .B(n20605), .Z(n20610) );
  XOR U21154 ( .A(n20608), .B(n20607), .Z(n20609) );
  NANDN U21155 ( .A(n20610), .B(n20609), .Z(n20612) );
  NAND U21156 ( .A(a[15]), .B(b[5]), .Z(n20948) );
  XNOR U21157 ( .A(n20610), .B(n20609), .Z(n20949) );
  NANDN U21158 ( .A(n20948), .B(n20949), .Z(n20611) );
  AND U21159 ( .A(n20612), .B(n20611), .Z(n20616) );
  AND U21160 ( .A(a[16]), .B(b[5]), .Z(n20615) );
  NANDN U21161 ( .A(n20616), .B(n20615), .Z(n20618) );
  XNOR U21162 ( .A(n20614), .B(n20613), .Z(n20861) );
  XNOR U21163 ( .A(n20616), .B(n20615), .Z(n20860) );
  NAND U21164 ( .A(n20861), .B(n20860), .Z(n20617) );
  NAND U21165 ( .A(n20618), .B(n20617), .Z(n20953) );
  NAND U21166 ( .A(a[17]), .B(b[5]), .Z(n20955) );
  AND U21167 ( .A(a[18]), .B(b[5]), .Z(n20623) );
  NANDN U21168 ( .A(n20624), .B(n20623), .Z(n20626) );
  XNOR U21169 ( .A(n20620), .B(n20619), .Z(n20621) );
  XNOR U21170 ( .A(n20622), .B(n20621), .Z(n20859) );
  XNOR U21171 ( .A(n20624), .B(n20623), .Z(n20858) );
  NAND U21172 ( .A(n20859), .B(n20858), .Z(n20625) );
  NAND U21173 ( .A(n20626), .B(n20625), .Z(n20961) );
  NAND U21174 ( .A(a[19]), .B(b[5]), .Z(n20963) );
  AND U21175 ( .A(a[20]), .B(b[5]), .Z(n20631) );
  NANDN U21176 ( .A(n20632), .B(n20631), .Z(n20634) );
  XNOR U21177 ( .A(n20628), .B(n20627), .Z(n20629) );
  XNOR U21178 ( .A(n20630), .B(n20629), .Z(n20857) );
  XNOR U21179 ( .A(n20632), .B(n20631), .Z(n20856) );
  NAND U21180 ( .A(n20857), .B(n20856), .Z(n20633) );
  NAND U21181 ( .A(n20634), .B(n20633), .Z(n20969) );
  NAND U21182 ( .A(a[21]), .B(b[5]), .Z(n20971) );
  AND U21183 ( .A(a[22]), .B(b[5]), .Z(n20639) );
  NANDN U21184 ( .A(n20640), .B(n20639), .Z(n20642) );
  XNOR U21185 ( .A(n20636), .B(n20635), .Z(n20637) );
  XNOR U21186 ( .A(n20638), .B(n20637), .Z(n20855) );
  XNOR U21187 ( .A(n20640), .B(n20639), .Z(n20854) );
  NAND U21188 ( .A(n20855), .B(n20854), .Z(n20641) );
  NAND U21189 ( .A(n20642), .B(n20641), .Z(n20976) );
  NAND U21190 ( .A(a[23]), .B(b[5]), .Z(n20979) );
  AND U21191 ( .A(a[24]), .B(b[5]), .Z(n20647) );
  NANDN U21192 ( .A(n20648), .B(n20647), .Z(n20650) );
  XOR U21193 ( .A(n20644), .B(n20643), .Z(n20645) );
  XNOR U21194 ( .A(n20646), .B(n20645), .Z(n20985) );
  XNOR U21195 ( .A(n20648), .B(n20647), .Z(n20984) );
  NAND U21196 ( .A(n20985), .B(n20984), .Z(n20649) );
  NAND U21197 ( .A(n20650), .B(n20649), .Z(n20987) );
  NAND U21198 ( .A(a[25]), .B(b[5]), .Z(n20989) );
  AND U21199 ( .A(a[26]), .B(b[5]), .Z(n20655) );
  NANDN U21200 ( .A(n20656), .B(n20655), .Z(n20658) );
  XNOR U21201 ( .A(n20652), .B(n20651), .Z(n20653) );
  XNOR U21202 ( .A(n20654), .B(n20653), .Z(n20853) );
  XNOR U21203 ( .A(n20656), .B(n20655), .Z(n20852) );
  NAND U21204 ( .A(n20853), .B(n20852), .Z(n20657) );
  NAND U21205 ( .A(n20658), .B(n20657), .Z(n20995) );
  NAND U21206 ( .A(a[27]), .B(b[5]), .Z(n20997) );
  AND U21207 ( .A(a[28]), .B(b[5]), .Z(n20663) );
  NANDN U21208 ( .A(n20664), .B(n20663), .Z(n20666) );
  XNOR U21209 ( .A(n20660), .B(n20659), .Z(n20661) );
  XNOR U21210 ( .A(n20662), .B(n20661), .Z(n20851) );
  XNOR U21211 ( .A(n20664), .B(n20663), .Z(n20850) );
  NAND U21212 ( .A(n20851), .B(n20850), .Z(n20665) );
  AND U21213 ( .A(n20666), .B(n20665), .Z(n21002) );
  AND U21214 ( .A(a[29]), .B(b[5]), .Z(n21005) );
  NANDN U21215 ( .A(n20671), .B(n20672), .Z(n20674) );
  XOR U21216 ( .A(n20668), .B(n20667), .Z(n20669) );
  XNOR U21217 ( .A(n20670), .B(n20669), .Z(n20849) );
  XNOR U21218 ( .A(n20672), .B(n20671), .Z(n20848) );
  NAND U21219 ( .A(n20849), .B(n20848), .Z(n20673) );
  NAND U21220 ( .A(n20674), .B(n20673), .Z(n21013) );
  AND U21221 ( .A(a[31]), .B(b[5]), .Z(n21015) );
  AND U21222 ( .A(a[32]), .B(b[5]), .Z(n20679) );
  NANDN U21223 ( .A(n20680), .B(n20679), .Z(n20682) );
  XNOR U21224 ( .A(n20676), .B(n20675), .Z(n20677) );
  XNOR U21225 ( .A(n20678), .B(n20677), .Z(n21019) );
  XNOR U21226 ( .A(n20680), .B(n20679), .Z(n21018) );
  NAND U21227 ( .A(n21019), .B(n21018), .Z(n20681) );
  NAND U21228 ( .A(n20682), .B(n20681), .Z(n21021) );
  AND U21229 ( .A(a[33]), .B(b[5]), .Z(n21023) );
  AND U21230 ( .A(a[34]), .B(b[5]), .Z(n20683) );
  NANDN U21231 ( .A(n20684), .B(n20683), .Z(n20690) );
  XOR U21232 ( .A(n20684), .B(n20683), .Z(n20846) );
  XOR U21233 ( .A(n20686), .B(n20685), .Z(n20687) );
  XNOR U21234 ( .A(n20688), .B(n20687), .Z(n20847) );
  NANDN U21235 ( .A(n20846), .B(n20847), .Z(n20689) );
  AND U21236 ( .A(n20690), .B(n20689), .Z(n21028) );
  NAND U21237 ( .A(a[35]), .B(b[5]), .Z(n21031) );
  NANDN U21238 ( .A(n20695), .B(n20696), .Z(n20698) );
  XNOR U21239 ( .A(n20692), .B(n20691), .Z(n20693) );
  XNOR U21240 ( .A(n20694), .B(n20693), .Z(n20845) );
  XNOR U21241 ( .A(n20696), .B(n20695), .Z(n20844) );
  NAND U21242 ( .A(n20845), .B(n20844), .Z(n20697) );
  NAND U21243 ( .A(n20698), .B(n20697), .Z(n21037) );
  NAND U21244 ( .A(a[37]), .B(b[5]), .Z(n21039) );
  AND U21245 ( .A(a[38]), .B(b[5]), .Z(n20703) );
  NANDN U21246 ( .A(n20704), .B(n20703), .Z(n20706) );
  XNOR U21247 ( .A(n20700), .B(n20699), .Z(n20701) );
  XNOR U21248 ( .A(n20702), .B(n20701), .Z(n20843) );
  XNOR U21249 ( .A(n20704), .B(n20703), .Z(n20842) );
  NAND U21250 ( .A(n20843), .B(n20842), .Z(n20705) );
  NAND U21251 ( .A(n20706), .B(n20705), .Z(n21045) );
  NAND U21252 ( .A(a[39]), .B(b[5]), .Z(n21047) );
  AND U21253 ( .A(a[40]), .B(b[5]), .Z(n20711) );
  NANDN U21254 ( .A(n20712), .B(n20711), .Z(n20714) );
  XNOR U21255 ( .A(n20708), .B(n20707), .Z(n20709) );
  XNOR U21256 ( .A(n20710), .B(n20709), .Z(n20841) );
  XNOR U21257 ( .A(n20712), .B(n20711), .Z(n20840) );
  NAND U21258 ( .A(n20841), .B(n20840), .Z(n20713) );
  NAND U21259 ( .A(n20714), .B(n20713), .Z(n21053) );
  NAND U21260 ( .A(a[41]), .B(b[5]), .Z(n21055) );
  AND U21261 ( .A(a[42]), .B(b[5]), .Z(n20719) );
  NANDN U21262 ( .A(n20720), .B(n20719), .Z(n20722) );
  XNOR U21263 ( .A(n20716), .B(n20715), .Z(n20717) );
  XNOR U21264 ( .A(n20718), .B(n20717), .Z(n20839) );
  XNOR U21265 ( .A(n20720), .B(n20719), .Z(n20838) );
  NAND U21266 ( .A(n20839), .B(n20838), .Z(n20721) );
  NAND U21267 ( .A(n20722), .B(n20721), .Z(n21061) );
  NAND U21268 ( .A(a[43]), .B(b[5]), .Z(n21063) );
  AND U21269 ( .A(a[44]), .B(b[5]), .Z(n20727) );
  NANDN U21270 ( .A(n20728), .B(n20727), .Z(n20730) );
  XNOR U21271 ( .A(n20724), .B(n20723), .Z(n20725) );
  XNOR U21272 ( .A(n20726), .B(n20725), .Z(n20837) );
  XNOR U21273 ( .A(n20728), .B(n20727), .Z(n20836) );
  NAND U21274 ( .A(n20837), .B(n20836), .Z(n20729) );
  NAND U21275 ( .A(n20730), .B(n20729), .Z(n21071) );
  NAND U21276 ( .A(a[45]), .B(b[5]), .Z(n21073) );
  AND U21277 ( .A(a[46]), .B(b[5]), .Z(n20735) );
  NANDN U21278 ( .A(n20736), .B(n20735), .Z(n20738) );
  XNOR U21279 ( .A(n20732), .B(n20731), .Z(n20733) );
  XNOR U21280 ( .A(n20734), .B(n20733), .Z(n20835) );
  XNOR U21281 ( .A(n20736), .B(n20735), .Z(n20834) );
  NAND U21282 ( .A(n20835), .B(n20834), .Z(n20737) );
  NAND U21283 ( .A(n20738), .B(n20737), .Z(n21077) );
  NAND U21284 ( .A(a[47]), .B(b[5]), .Z(n21079) );
  AND U21285 ( .A(a[48]), .B(b[5]), .Z(n20743) );
  NANDN U21286 ( .A(n20744), .B(n20743), .Z(n20746) );
  XNOR U21287 ( .A(n20740), .B(n20739), .Z(n20741) );
  XNOR U21288 ( .A(n20742), .B(n20741), .Z(n20833) );
  XNOR U21289 ( .A(n20744), .B(n20743), .Z(n20832) );
  NAND U21290 ( .A(n20833), .B(n20832), .Z(n20745) );
  NAND U21291 ( .A(n20746), .B(n20745), .Z(n21085) );
  NAND U21292 ( .A(a[49]), .B(b[5]), .Z(n21087) );
  AND U21293 ( .A(a[50]), .B(b[5]), .Z(n20747) );
  NANDN U21294 ( .A(n20748), .B(n20747), .Z(n20754) );
  XNOR U21295 ( .A(n20748), .B(n20747), .Z(n20831) );
  XNOR U21296 ( .A(n20750), .B(n20749), .Z(n20751) );
  XNOR U21297 ( .A(n20752), .B(n20751), .Z(n20830) );
  NAND U21298 ( .A(n20831), .B(n20830), .Z(n20753) );
  NAND U21299 ( .A(n20754), .B(n20753), .Z(n21093) );
  NAND U21300 ( .A(a[51]), .B(b[5]), .Z(n21095) );
  XOR U21301 ( .A(n20759), .B(n20758), .Z(n20760) );
  XOR U21302 ( .A(n20761), .B(n20760), .Z(n21102) );
  NAND U21303 ( .A(a[53]), .B(b[5]), .Z(n21104) );
  NANDN U21304 ( .A(n21108), .B(n21109), .Z(n20769) );
  NOR U21305 ( .A(n20762), .B(n21109), .Z(n20767) );
  XOR U21306 ( .A(n20764), .B(n20763), .Z(n20765) );
  XNOR U21307 ( .A(n20766), .B(n20765), .Z(n21111) );
  OR U21308 ( .A(n20767), .B(n21111), .Z(n20768) );
  AND U21309 ( .A(n20769), .B(n20768), .Z(n21117) );
  XOR U21310 ( .A(n20771), .B(n20770), .Z(n20772) );
  IV U21311 ( .A(n20772), .Z(n21116) );
  OR U21312 ( .A(n21117), .B(n21116), .Z(n20775) );
  ANDN U21313 ( .B(n21117), .A(n20772), .Z(n20773) );
  NAND U21314 ( .A(a[55]), .B(b[5]), .Z(n21119) );
  OR U21315 ( .A(n20773), .B(n21119), .Z(n20774) );
  AND U21316 ( .A(n20775), .B(n20774), .Z(n20777) );
  AND U21317 ( .A(a[56]), .B(b[5]), .Z(n20776) );
  NANDN U21318 ( .A(n20777), .B(n20776), .Z(n20783) );
  XNOR U21319 ( .A(n20777), .B(n20776), .Z(n20825) );
  XNOR U21320 ( .A(n20779), .B(n20778), .Z(n20780) );
  XNOR U21321 ( .A(n20781), .B(n20780), .Z(n20824) );
  NAND U21322 ( .A(n20825), .B(n20824), .Z(n20782) );
  NAND U21323 ( .A(n20783), .B(n20782), .Z(n21127) );
  NAND U21324 ( .A(a[57]), .B(b[5]), .Z(n21129) );
  AND U21325 ( .A(a[58]), .B(b[5]), .Z(n20788) );
  NANDN U21326 ( .A(n20789), .B(n20788), .Z(n20791) );
  XNOR U21327 ( .A(n20785), .B(n20784), .Z(n20786) );
  XNOR U21328 ( .A(n20787), .B(n20786), .Z(n20823) );
  XNOR U21329 ( .A(n20789), .B(n20788), .Z(n20822) );
  NAND U21330 ( .A(n20823), .B(n20822), .Z(n20790) );
  AND U21331 ( .A(n20791), .B(n20790), .Z(n20794) );
  NANDN U21332 ( .A(n20794), .B(n20795), .Z(n20797) );
  AND U21333 ( .A(a[59]), .B(b[5]), .Z(n21135) );
  NAND U21334 ( .A(n21135), .B(n21134), .Z(n20796) );
  NAND U21335 ( .A(n20797), .B(n20796), .Z(n21141) );
  NANDN U21336 ( .A(n20818), .B(n20819), .Z(n20803) );
  NOR U21337 ( .A(n20798), .B(n20819), .Z(n20801) );
  XOR U21338 ( .A(n20800), .B(n20799), .Z(n20821) );
  OR U21339 ( .A(n20801), .B(n20821), .Z(n20802) );
  AND U21340 ( .A(n20803), .B(n20802), .Z(n20807) );
  AND U21341 ( .A(a[62]), .B(b[5]), .Z(n20806) );
  XOR U21342 ( .A(n20805), .B(n20804), .Z(n21146) );
  XNOR U21343 ( .A(n20807), .B(n20806), .Z(n21147) );
  NANDN U21344 ( .A(n20809), .B(n20808), .Z(n20813) );
  XOR U21345 ( .A(n20809), .B(n20808), .Z(n20816) );
  XOR U21346 ( .A(n20811), .B(n20810), .Z(n20817) );
  NANDN U21347 ( .A(n20816), .B(n20817), .Z(n20812) );
  AND U21348 ( .A(n20813), .B(n20812), .Z(n21153) );
  XOR U21349 ( .A(n20815), .B(n20814), .Z(n21152) );
  AND U21350 ( .A(n21153), .B(n21152), .Z(n24678) );
  XOR U21351 ( .A(n20817), .B(n20816), .Z(n22496) );
  XOR U21352 ( .A(n20819), .B(n20818), .Z(n20820) );
  XNOR U21353 ( .A(n20821), .B(n20820), .Z(n21481) );
  AND U21354 ( .A(a[62]), .B(b[4]), .Z(n21480) );
  XNOR U21355 ( .A(n20823), .B(n20822), .Z(n21468) );
  XOR U21356 ( .A(n20825), .B(n20824), .Z(n21120) );
  IV U21357 ( .A(n21120), .Z(n21456) );
  NAND U21358 ( .A(a[56]), .B(b[4]), .Z(n21448) );
  AND U21359 ( .A(a[54]), .B(b[4]), .Z(n21100) );
  IV U21360 ( .A(n21100), .Z(n21156) );
  XOR U21361 ( .A(n20827), .B(n20826), .Z(n20828) );
  XOR U21362 ( .A(n20829), .B(n20828), .Z(n21433) );
  XNOR U21363 ( .A(n20831), .B(n20830), .Z(n21424) );
  XNOR U21364 ( .A(n20833), .B(n20832), .Z(n21416) );
  XNOR U21365 ( .A(n20835), .B(n20834), .Z(n21408) );
  XNOR U21366 ( .A(n20837), .B(n20836), .Z(n21400) );
  XNOR U21367 ( .A(n20839), .B(n20838), .Z(n21392) );
  XNOR U21368 ( .A(n20841), .B(n20840), .Z(n21384) );
  XNOR U21369 ( .A(n20843), .B(n20842), .Z(n21376) );
  XNOR U21370 ( .A(n20845), .B(n20844), .Z(n21368) );
  NAND U21371 ( .A(a[36]), .B(b[4]), .Z(n21032) );
  XNOR U21372 ( .A(n20847), .B(n20846), .Z(n21363) );
  AND U21373 ( .A(a[32]), .B(b[4]), .Z(n21011) );
  XNOR U21374 ( .A(n20849), .B(n20848), .Z(n21344) );
  XNOR U21375 ( .A(n20851), .B(n20850), .Z(n21336) );
  XNOR U21376 ( .A(n20853), .B(n20852), .Z(n21328) );
  AND U21377 ( .A(a[24]), .B(b[4]), .Z(n20981) );
  XNOR U21378 ( .A(n20855), .B(n20854), .Z(n21312) );
  XNOR U21379 ( .A(n20857), .B(n20856), .Z(n21304) );
  XNOR U21380 ( .A(n20859), .B(n20858), .Z(n21296) );
  XNOR U21381 ( .A(n20861), .B(n20860), .Z(n21288) );
  XOR U21382 ( .A(n20863), .B(n20862), .Z(n20908) );
  AND U21383 ( .A(a[8]), .B(b[4]), .Z(n20903) );
  AND U21384 ( .A(a[1]), .B(b[5]), .Z(n20869) );
  AND U21385 ( .A(b[4]), .B(a[0]), .Z(n21530) );
  AND U21386 ( .A(n20869), .B(n21530), .Z(n20866) );
  NAND U21387 ( .A(a[2]), .B(n20866), .Z(n20873) );
  NAND U21388 ( .A(b[5]), .B(a[1]), .Z(n20867) );
  XOR U21389 ( .A(n20868), .B(n20867), .Z(n21206) );
  NAND U21390 ( .A(n20869), .B(a[0]), .Z(n20870) );
  XNOR U21391 ( .A(a[2]), .B(n20870), .Z(n20871) );
  AND U21392 ( .A(b[4]), .B(n20871), .Z(n21207) );
  NANDN U21393 ( .A(n21206), .B(n21207), .Z(n20872) );
  AND U21394 ( .A(n20873), .B(n20872), .Z(n20876) );
  NANDN U21395 ( .A(n20876), .B(n20877), .Z(n20879) );
  NAND U21396 ( .A(a[3]), .B(b[4]), .Z(n21212) );
  NANDN U21397 ( .A(n21212), .B(n21213), .Z(n20878) );
  AND U21398 ( .A(n20879), .B(n20878), .Z(n20880) );
  AND U21399 ( .A(a[4]), .B(b[4]), .Z(n20881) );
  NANDN U21400 ( .A(n20880), .B(n20881), .Z(n20885) );
  NAND U21401 ( .A(n21217), .B(n21216), .Z(n20884) );
  NAND U21402 ( .A(n20885), .B(n20884), .Z(n20886) );
  NAND U21403 ( .A(n20887), .B(n20886), .Z(n20889) );
  NAND U21404 ( .A(a[5]), .B(b[4]), .Z(n21222) );
  XOR U21405 ( .A(n20887), .B(n20886), .Z(n21223) );
  NANDN U21406 ( .A(n21222), .B(n21223), .Z(n20888) );
  AND U21407 ( .A(n20889), .B(n20888), .Z(n20892) );
  NANDN U21408 ( .A(n20892), .B(n20893), .Z(n20895) );
  NAND U21409 ( .A(a[6]), .B(b[4]), .Z(n21228) );
  NANDN U21410 ( .A(n21228), .B(n21229), .Z(n20894) );
  AND U21411 ( .A(n20895), .B(n20894), .Z(n20898) );
  XOR U21412 ( .A(n20897), .B(n20896), .Z(n20899) );
  NANDN U21413 ( .A(n20898), .B(n20899), .Z(n20901) );
  NAND U21414 ( .A(a[7]), .B(b[4]), .Z(n21236) );
  NANDN U21415 ( .A(n21236), .B(n21237), .Z(n20900) );
  AND U21416 ( .A(n20901), .B(n20900), .Z(n20902) );
  NANDN U21417 ( .A(n20903), .B(n20902), .Z(n20907) );
  XOR U21418 ( .A(n20903), .B(n20902), .Z(n21240) );
  XOR U21419 ( .A(n20905), .B(n20904), .Z(n21241) );
  OR U21420 ( .A(n21240), .B(n21241), .Z(n20906) );
  AND U21421 ( .A(n20907), .B(n20906), .Z(n20909) );
  NANDN U21422 ( .A(n20908), .B(n20909), .Z(n20911) );
  NAND U21423 ( .A(a[9]), .B(b[4]), .Z(n21248) );
  XNOR U21424 ( .A(n20909), .B(n20908), .Z(n21249) );
  NANDN U21425 ( .A(n21248), .B(n21249), .Z(n20910) );
  AND U21426 ( .A(n20911), .B(n20910), .Z(n20915) );
  AND U21427 ( .A(a[10]), .B(b[4]), .Z(n20914) );
  NANDN U21428 ( .A(n20915), .B(n20914), .Z(n20917) );
  XOR U21429 ( .A(n20913), .B(n20912), .Z(n21252) );
  XNOR U21430 ( .A(n20915), .B(n20914), .Z(n21253) );
  NANDN U21431 ( .A(n21252), .B(n21253), .Z(n20916) );
  AND U21432 ( .A(n20917), .B(n20916), .Z(n20921) );
  XOR U21433 ( .A(n20919), .B(n20918), .Z(n20920) );
  NANDN U21434 ( .A(n20921), .B(n20920), .Z(n20923) );
  NAND U21435 ( .A(a[11]), .B(b[4]), .Z(n21260) );
  XNOR U21436 ( .A(n20921), .B(n20920), .Z(n21261) );
  NANDN U21437 ( .A(n21260), .B(n21261), .Z(n20922) );
  AND U21438 ( .A(n20923), .B(n20922), .Z(n20927) );
  AND U21439 ( .A(a[12]), .B(b[4]), .Z(n20926) );
  XNOR U21440 ( .A(n20925), .B(n20924), .Z(n21264) );
  XNOR U21441 ( .A(n20927), .B(n20926), .Z(n21265) );
  XOR U21442 ( .A(n20929), .B(n20928), .Z(n20930) );
  NANDN U21443 ( .A(n20931), .B(n20930), .Z(n20933) );
  NAND U21444 ( .A(a[13]), .B(b[4]), .Z(n21270) );
  XNOR U21445 ( .A(n20931), .B(n20930), .Z(n21271) );
  NANDN U21446 ( .A(n21270), .B(n21271), .Z(n20932) );
  AND U21447 ( .A(n20933), .B(n20932), .Z(n20935) );
  AND U21448 ( .A(a[14]), .B(b[4]), .Z(n20934) );
  NANDN U21449 ( .A(n20935), .B(n20934), .Z(n20939) );
  XNOR U21450 ( .A(n20935), .B(n20934), .Z(n21277) );
  XNOR U21451 ( .A(n20937), .B(n20936), .Z(n21276) );
  NAND U21452 ( .A(n21277), .B(n21276), .Z(n20938) );
  AND U21453 ( .A(n20939), .B(n20938), .Z(n20943) );
  XOR U21454 ( .A(n20941), .B(n20940), .Z(n20942) );
  NANDN U21455 ( .A(n20943), .B(n20942), .Z(n20945) );
  NAND U21456 ( .A(a[15]), .B(b[4]), .Z(n21282) );
  XNOR U21457 ( .A(n20943), .B(n20942), .Z(n21283) );
  NANDN U21458 ( .A(n21282), .B(n21283), .Z(n20944) );
  AND U21459 ( .A(n20945), .B(n20944), .Z(n20947) );
  AND U21460 ( .A(a[16]), .B(b[4]), .Z(n20946) );
  NANDN U21461 ( .A(n20947), .B(n20946), .Z(n20951) );
  XNOR U21462 ( .A(n20947), .B(n20946), .Z(n21197) );
  XNOR U21463 ( .A(n20949), .B(n20948), .Z(n21196) );
  NAND U21464 ( .A(n21197), .B(n21196), .Z(n20950) );
  NAND U21465 ( .A(n20951), .B(n20950), .Z(n21289) );
  NAND U21466 ( .A(a[17]), .B(b[4]), .Z(n21291) );
  AND U21467 ( .A(a[18]), .B(b[4]), .Z(n20956) );
  NANDN U21468 ( .A(n20957), .B(n20956), .Z(n20959) );
  XNOR U21469 ( .A(n20953), .B(n20952), .Z(n20954) );
  XNOR U21470 ( .A(n20955), .B(n20954), .Z(n21195) );
  XNOR U21471 ( .A(n20957), .B(n20956), .Z(n21194) );
  NAND U21472 ( .A(n21195), .B(n21194), .Z(n20958) );
  NAND U21473 ( .A(n20959), .B(n20958), .Z(n21297) );
  NAND U21474 ( .A(a[19]), .B(b[4]), .Z(n21299) );
  AND U21475 ( .A(a[20]), .B(b[4]), .Z(n20964) );
  NANDN U21476 ( .A(n20965), .B(n20964), .Z(n20967) );
  XNOR U21477 ( .A(n20961), .B(n20960), .Z(n20962) );
  XNOR U21478 ( .A(n20963), .B(n20962), .Z(n21193) );
  XNOR U21479 ( .A(n20965), .B(n20964), .Z(n21192) );
  NAND U21480 ( .A(n21193), .B(n21192), .Z(n20966) );
  NAND U21481 ( .A(n20967), .B(n20966), .Z(n21305) );
  NAND U21482 ( .A(a[21]), .B(b[4]), .Z(n21307) );
  AND U21483 ( .A(a[22]), .B(b[4]), .Z(n20972) );
  NANDN U21484 ( .A(n20973), .B(n20972), .Z(n20975) );
  XNOR U21485 ( .A(n20969), .B(n20968), .Z(n20970) );
  XNOR U21486 ( .A(n20971), .B(n20970), .Z(n21191) );
  XNOR U21487 ( .A(n20973), .B(n20972), .Z(n21190) );
  NAND U21488 ( .A(n21191), .B(n21190), .Z(n20974) );
  NAND U21489 ( .A(n20975), .B(n20974), .Z(n21313) );
  NAND U21490 ( .A(a[23]), .B(b[4]), .Z(n21315) );
  NANDN U21491 ( .A(n20981), .B(n20980), .Z(n20983) );
  XOR U21492 ( .A(n20977), .B(n20976), .Z(n20978) );
  XOR U21493 ( .A(n20979), .B(n20978), .Z(n21189) );
  XNOR U21494 ( .A(n20981), .B(n20980), .Z(n21188) );
  NANDN U21495 ( .A(n21189), .B(n21188), .Z(n20982) );
  NAND U21496 ( .A(n20983), .B(n20982), .Z(n21321) );
  XOR U21497 ( .A(n20985), .B(n20984), .Z(n21320) );
  AND U21498 ( .A(a[25]), .B(b[4]), .Z(n21323) );
  AND U21499 ( .A(a[26]), .B(b[4]), .Z(n20990) );
  NANDN U21500 ( .A(n20991), .B(n20990), .Z(n20993) );
  XNOR U21501 ( .A(n20987), .B(n20986), .Z(n20988) );
  XNOR U21502 ( .A(n20989), .B(n20988), .Z(n21187) );
  XNOR U21503 ( .A(n20991), .B(n20990), .Z(n21186) );
  NAND U21504 ( .A(n21187), .B(n21186), .Z(n20992) );
  NAND U21505 ( .A(n20993), .B(n20992), .Z(n21329) );
  NAND U21506 ( .A(a[27]), .B(b[4]), .Z(n21331) );
  AND U21507 ( .A(a[28]), .B(b[4]), .Z(n20998) );
  NANDN U21508 ( .A(n20999), .B(n20998), .Z(n21001) );
  XNOR U21509 ( .A(n20995), .B(n20994), .Z(n20996) );
  XNOR U21510 ( .A(n20997), .B(n20996), .Z(n21185) );
  XNOR U21511 ( .A(n20999), .B(n20998), .Z(n21184) );
  NAND U21512 ( .A(n21185), .B(n21184), .Z(n21000) );
  NAND U21513 ( .A(n21001), .B(n21000), .Z(n21337) );
  NAND U21514 ( .A(a[29]), .B(b[4]), .Z(n21339) );
  AND U21515 ( .A(a[30]), .B(b[4]), .Z(n21006) );
  NANDN U21516 ( .A(n21007), .B(n21006), .Z(n21009) );
  XOR U21517 ( .A(n21003), .B(n21002), .Z(n21004) );
  XNOR U21518 ( .A(n21005), .B(n21004), .Z(n21183) );
  XNOR U21519 ( .A(n21007), .B(n21006), .Z(n21182) );
  NAND U21520 ( .A(n21183), .B(n21182), .Z(n21008) );
  NAND U21521 ( .A(n21009), .B(n21008), .Z(n21345) );
  NAND U21522 ( .A(a[31]), .B(b[4]), .Z(n21347) );
  NANDN U21523 ( .A(n21011), .B(n21010), .Z(n21017) );
  XNOR U21524 ( .A(n21011), .B(n21010), .Z(n21180) );
  XNOR U21525 ( .A(n21013), .B(n21012), .Z(n21014) );
  XNOR U21526 ( .A(n21015), .B(n21014), .Z(n21181) );
  NAND U21527 ( .A(n21180), .B(n21181), .Z(n21016) );
  NAND U21528 ( .A(n21017), .B(n21016), .Z(n21353) );
  XOR U21529 ( .A(n21019), .B(n21018), .Z(n21352) );
  AND U21530 ( .A(a[33]), .B(b[4]), .Z(n21355) );
  AND U21531 ( .A(a[34]), .B(b[4]), .Z(n21024) );
  NANDN U21532 ( .A(n21025), .B(n21024), .Z(n21027) );
  XOR U21533 ( .A(n21021), .B(n21020), .Z(n21022) );
  XNOR U21534 ( .A(n21023), .B(n21022), .Z(n21179) );
  XNOR U21535 ( .A(n21025), .B(n21024), .Z(n21178) );
  NAND U21536 ( .A(n21179), .B(n21178), .Z(n21026) );
  AND U21537 ( .A(n21027), .B(n21026), .Z(n21362) );
  NAND U21538 ( .A(a[35]), .B(b[4]), .Z(n21365) );
  NANDN U21539 ( .A(n21032), .B(n21033), .Z(n21035) );
  XNOR U21540 ( .A(n21029), .B(n21028), .Z(n21030) );
  XNOR U21541 ( .A(n21031), .B(n21030), .Z(n21177) );
  XNOR U21542 ( .A(n21033), .B(n21032), .Z(n21176) );
  NAND U21543 ( .A(n21177), .B(n21176), .Z(n21034) );
  NAND U21544 ( .A(n21035), .B(n21034), .Z(n21369) );
  NAND U21545 ( .A(a[37]), .B(b[4]), .Z(n21371) );
  AND U21546 ( .A(a[38]), .B(b[4]), .Z(n21040) );
  NANDN U21547 ( .A(n21041), .B(n21040), .Z(n21043) );
  XNOR U21548 ( .A(n21037), .B(n21036), .Z(n21038) );
  XNOR U21549 ( .A(n21039), .B(n21038), .Z(n21175) );
  XNOR U21550 ( .A(n21041), .B(n21040), .Z(n21174) );
  NAND U21551 ( .A(n21175), .B(n21174), .Z(n21042) );
  NAND U21552 ( .A(n21043), .B(n21042), .Z(n21377) );
  NAND U21553 ( .A(a[39]), .B(b[4]), .Z(n21379) );
  AND U21554 ( .A(a[40]), .B(b[4]), .Z(n21048) );
  NANDN U21555 ( .A(n21049), .B(n21048), .Z(n21051) );
  XNOR U21556 ( .A(n21045), .B(n21044), .Z(n21046) );
  XNOR U21557 ( .A(n21047), .B(n21046), .Z(n21173) );
  XNOR U21558 ( .A(n21049), .B(n21048), .Z(n21172) );
  NAND U21559 ( .A(n21173), .B(n21172), .Z(n21050) );
  NAND U21560 ( .A(n21051), .B(n21050), .Z(n21385) );
  NAND U21561 ( .A(a[41]), .B(b[4]), .Z(n21387) );
  AND U21562 ( .A(a[42]), .B(b[4]), .Z(n21056) );
  NANDN U21563 ( .A(n21057), .B(n21056), .Z(n21059) );
  XNOR U21564 ( .A(n21053), .B(n21052), .Z(n21054) );
  XNOR U21565 ( .A(n21055), .B(n21054), .Z(n21171) );
  XNOR U21566 ( .A(n21057), .B(n21056), .Z(n21170) );
  NAND U21567 ( .A(n21171), .B(n21170), .Z(n21058) );
  NAND U21568 ( .A(n21059), .B(n21058), .Z(n21393) );
  NAND U21569 ( .A(a[43]), .B(b[4]), .Z(n21395) );
  AND U21570 ( .A(a[44]), .B(b[4]), .Z(n21064) );
  NANDN U21571 ( .A(n21065), .B(n21064), .Z(n21067) );
  XNOR U21572 ( .A(n21061), .B(n21060), .Z(n21062) );
  XNOR U21573 ( .A(n21063), .B(n21062), .Z(n21169) );
  XNOR U21574 ( .A(n21065), .B(n21064), .Z(n21168) );
  NAND U21575 ( .A(n21169), .B(n21168), .Z(n21066) );
  NAND U21576 ( .A(n21067), .B(n21066), .Z(n21401) );
  NAND U21577 ( .A(a[45]), .B(b[4]), .Z(n21403) );
  AND U21578 ( .A(a[46]), .B(b[4]), .Z(n21068) );
  NANDN U21579 ( .A(n21069), .B(n21068), .Z(n21075) );
  XOR U21580 ( .A(n21069), .B(n21068), .Z(n21166) );
  XNOR U21581 ( .A(n21071), .B(n21070), .Z(n21072) );
  XNOR U21582 ( .A(n21073), .B(n21072), .Z(n21167) );
  NANDN U21583 ( .A(n21166), .B(n21167), .Z(n21074) );
  NAND U21584 ( .A(n21075), .B(n21074), .Z(n21409) );
  NAND U21585 ( .A(a[47]), .B(b[4]), .Z(n21411) );
  AND U21586 ( .A(a[48]), .B(b[4]), .Z(n21080) );
  NANDN U21587 ( .A(n21081), .B(n21080), .Z(n21083) );
  XNOR U21588 ( .A(n21077), .B(n21076), .Z(n21078) );
  XNOR U21589 ( .A(n21079), .B(n21078), .Z(n21165) );
  XNOR U21590 ( .A(n21081), .B(n21080), .Z(n21164) );
  NAND U21591 ( .A(n21165), .B(n21164), .Z(n21082) );
  NAND U21592 ( .A(n21083), .B(n21082), .Z(n21417) );
  NAND U21593 ( .A(a[49]), .B(b[4]), .Z(n21419) );
  AND U21594 ( .A(a[50]), .B(b[4]), .Z(n21088) );
  NANDN U21595 ( .A(n21089), .B(n21088), .Z(n21091) );
  XNOR U21596 ( .A(n21085), .B(n21084), .Z(n21086) );
  XNOR U21597 ( .A(n21087), .B(n21086), .Z(n21163) );
  XNOR U21598 ( .A(n21089), .B(n21088), .Z(n21162) );
  NAND U21599 ( .A(n21163), .B(n21162), .Z(n21090) );
  NAND U21600 ( .A(n21091), .B(n21090), .Z(n21425) );
  NAND U21601 ( .A(a[51]), .B(b[4]), .Z(n21427) );
  AND U21602 ( .A(a[52]), .B(b[4]), .Z(n21096) );
  NANDN U21603 ( .A(n21097), .B(n21096), .Z(n21099) );
  XNOR U21604 ( .A(n21093), .B(n21092), .Z(n21094) );
  XNOR U21605 ( .A(n21095), .B(n21094), .Z(n21161) );
  XNOR U21606 ( .A(n21097), .B(n21096), .Z(n21160) );
  NAND U21607 ( .A(n21161), .B(n21160), .Z(n21098) );
  AND U21608 ( .A(n21099), .B(n21098), .Z(n21432) );
  NAND U21609 ( .A(a[53]), .B(b[4]), .Z(n21435) );
  NANDN U21610 ( .A(n21156), .B(n21157), .Z(n21107) );
  NOR U21611 ( .A(n21100), .B(n21157), .Z(n21105) );
  XNOR U21612 ( .A(n21102), .B(n21101), .Z(n21103) );
  XNOR U21613 ( .A(n21104), .B(n21103), .Z(n21159) );
  OR U21614 ( .A(n21105), .B(n21159), .Z(n21106) );
  AND U21615 ( .A(n21107), .B(n21106), .Z(n21442) );
  XOR U21616 ( .A(n21109), .B(n21108), .Z(n21110) );
  XOR U21617 ( .A(n21111), .B(n21110), .Z(n21112) );
  IV U21618 ( .A(n21112), .Z(n21441) );
  OR U21619 ( .A(n21442), .B(n21441), .Z(n21115) );
  ANDN U21620 ( .B(n21442), .A(n21112), .Z(n21113) );
  AND U21621 ( .A(a[55]), .B(b[4]), .Z(n21444) );
  NANDN U21622 ( .A(n21113), .B(n21444), .Z(n21114) );
  AND U21623 ( .A(n21115), .B(n21114), .Z(n21449) );
  XOR U21624 ( .A(n21117), .B(n21116), .Z(n21118) );
  XNOR U21625 ( .A(n21119), .B(n21118), .Z(n21451) );
  NANDN U21626 ( .A(n21456), .B(n21457), .Z(n21123) );
  NOR U21627 ( .A(n21120), .B(n21457), .Z(n21121) );
  AND U21628 ( .A(a[57]), .B(b[4]), .Z(n21459) );
  NANDN U21629 ( .A(n21121), .B(n21459), .Z(n21122) );
  AND U21630 ( .A(n21123), .B(n21122), .Z(n21124) );
  AND U21631 ( .A(a[58]), .B(b[4]), .Z(n21125) );
  NANDN U21632 ( .A(n21124), .B(n21125), .Z(n21131) );
  XOR U21633 ( .A(n21125), .B(n21124), .Z(n21460) );
  XNOR U21634 ( .A(n21127), .B(n21126), .Z(n21128) );
  XNOR U21635 ( .A(n21129), .B(n21128), .Z(n21461) );
  NANDN U21636 ( .A(n21460), .B(n21461), .Z(n21130) );
  NAND U21637 ( .A(n21131), .B(n21130), .Z(n21469) );
  NAND U21638 ( .A(a[59]), .B(b[4]), .Z(n21471) );
  AND U21639 ( .A(a[60]), .B(b[4]), .Z(n21132) );
  NANDN U21640 ( .A(n21133), .B(n21132), .Z(n21137) );
  XOR U21641 ( .A(n21133), .B(n21132), .Z(n21474) );
  XOR U21642 ( .A(n21135), .B(n21134), .Z(n21475) );
  NANDN U21643 ( .A(n21474), .B(n21475), .Z(n21136) );
  AND U21644 ( .A(n21137), .B(n21136), .Z(n21143) );
  AND U21645 ( .A(a[61]), .B(b[4]), .Z(n21142) );
  NANDN U21646 ( .A(n21143), .B(n21142), .Z(n21145) );
  XOR U21647 ( .A(n21139), .B(n21138), .Z(n21140) );
  XOR U21648 ( .A(n21141), .B(n21140), .Z(n21154) );
  XNOR U21649 ( .A(n21143), .B(n21142), .Z(n21155) );
  NANDN U21650 ( .A(n21154), .B(n21155), .Z(n21144) );
  NAND U21651 ( .A(n21145), .B(n21144), .Z(n21483) );
  XOR U21652 ( .A(n21147), .B(n21146), .Z(n21148) );
  NANDN U21653 ( .A(n21149), .B(n21148), .Z(n21151) );
  NAND U21654 ( .A(a[63]), .B(b[4]), .Z(n21488) );
  XNOR U21655 ( .A(n21149), .B(n21148), .Z(n21489) );
  NANDN U21656 ( .A(n21488), .B(n21489), .Z(n21150) );
  AND U21657 ( .A(n21151), .B(n21150), .Z(n22495) );
  XOR U21658 ( .A(n21153), .B(n21152), .Z(n24673) );
  NAND U21659 ( .A(a[63]), .B(b[3]), .Z(n21484) );
  AND U21660 ( .A(a[62]), .B(b[3]), .Z(n21823) );
  XOR U21661 ( .A(n21155), .B(n21154), .Z(n21822) );
  NAND U21662 ( .A(a[60]), .B(b[3]), .Z(n21466) );
  NAND U21663 ( .A(a[58]), .B(b[3]), .Z(n21795) );
  XOR U21664 ( .A(n21157), .B(n21156), .Z(n21158) );
  XNOR U21665 ( .A(n21159), .B(n21158), .Z(n21778) );
  XNOR U21666 ( .A(n21161), .B(n21160), .Z(n21770) );
  XNOR U21667 ( .A(n21163), .B(n21162), .Z(n21760) );
  XNOR U21668 ( .A(n21165), .B(n21164), .Z(n21752) );
  NAND U21669 ( .A(a[48]), .B(b[3]), .Z(n21412) );
  XNOR U21670 ( .A(n21167), .B(n21166), .Z(n21745) );
  XNOR U21671 ( .A(n21169), .B(n21168), .Z(n21736) );
  XNOR U21672 ( .A(n21171), .B(n21170), .Z(n21728) );
  XNOR U21673 ( .A(n21173), .B(n21172), .Z(n21720) );
  XNOR U21674 ( .A(n21175), .B(n21174), .Z(n21712) );
  XNOR U21675 ( .A(n21177), .B(n21176), .Z(n21702) );
  XNOR U21676 ( .A(n21179), .B(n21178), .Z(n21696) );
  NAND U21677 ( .A(a[34]), .B(b[3]), .Z(n21356) );
  XNOR U21678 ( .A(n21181), .B(n21180), .Z(n21687) );
  XNOR U21679 ( .A(n21183), .B(n21182), .Z(n21678) );
  XNOR U21680 ( .A(n21185), .B(n21184), .Z(n21670) );
  XNOR U21681 ( .A(n21187), .B(n21186), .Z(n21660) );
  XNOR U21682 ( .A(n21189), .B(n21188), .Z(n21652) );
  XNOR U21683 ( .A(n21191), .B(n21190), .Z(n21644) );
  XNOR U21684 ( .A(n21193), .B(n21192), .Z(n21636) );
  XNOR U21685 ( .A(n21195), .B(n21194), .Z(n21628) );
  XNOR U21686 ( .A(n21197), .B(n21196), .Z(n21620) );
  AND U21687 ( .A(b[3]), .B(a[0]), .Z(n21853) );
  AND U21688 ( .A(a[1]), .B(b[4]), .Z(n21201) );
  AND U21689 ( .A(n21853), .B(n21201), .Z(n21198) );
  NAND U21690 ( .A(a[2]), .B(n21198), .Z(n21205) );
  NAND U21691 ( .A(b[4]), .B(a[1]), .Z(n21199) );
  XOR U21692 ( .A(n21200), .B(n21199), .Z(n21536) );
  NAND U21693 ( .A(n21201), .B(a[0]), .Z(n21202) );
  XNOR U21694 ( .A(a[2]), .B(n21202), .Z(n21203) );
  AND U21695 ( .A(b[3]), .B(n21203), .Z(n21537) );
  NANDN U21696 ( .A(n21536), .B(n21537), .Z(n21204) );
  AND U21697 ( .A(n21205), .B(n21204), .Z(n21209) );
  NANDN U21698 ( .A(n21209), .B(n21208), .Z(n21211) );
  XNOR U21699 ( .A(n21209), .B(n21208), .Z(n21545) );
  AND U21700 ( .A(a[3]), .B(b[3]), .Z(n21544) );
  NAND U21701 ( .A(n21545), .B(n21544), .Z(n21210) );
  AND U21702 ( .A(n21211), .B(n21210), .Z(n21215) );
  AND U21703 ( .A(a[4]), .B(b[3]), .Z(n21214) );
  XNOR U21704 ( .A(n21215), .B(n21214), .Z(n21549) );
  XOR U21705 ( .A(n21217), .B(n21216), .Z(n21219) );
  NANDN U21706 ( .A(n21218), .B(n21219), .Z(n21221) );
  AND U21707 ( .A(a[5]), .B(b[3]), .Z(n21526) );
  NAND U21708 ( .A(n21527), .B(n21526), .Z(n21220) );
  AND U21709 ( .A(n21221), .B(n21220), .Z(n21224) );
  NANDN U21710 ( .A(n21224), .B(n21225), .Z(n21227) );
  NAND U21711 ( .A(a[6]), .B(b[3]), .Z(n21558) );
  NANDN U21712 ( .A(n21558), .B(n21559), .Z(n21226) );
  AND U21713 ( .A(n21227), .B(n21226), .Z(n21230) );
  NANDN U21714 ( .A(n21230), .B(n21231), .Z(n21233) );
  NAND U21715 ( .A(a[7]), .B(b[3]), .Z(n21566) );
  NANDN U21716 ( .A(n21566), .B(n21567), .Z(n21232) );
  AND U21717 ( .A(n21233), .B(n21232), .Z(n21234) );
  AND U21718 ( .A(a[8]), .B(b[3]), .Z(n21235) );
  NANDN U21719 ( .A(n21234), .B(n21235), .Z(n21239) );
  NAND U21720 ( .A(n21571), .B(n21570), .Z(n21238) );
  AND U21721 ( .A(n21239), .B(n21238), .Z(n21243) );
  XNOR U21722 ( .A(n21241), .B(n21240), .Z(n21242) );
  NANDN U21723 ( .A(n21243), .B(n21242), .Z(n21245) );
  NAND U21724 ( .A(a[9]), .B(b[3]), .Z(n21576) );
  XNOR U21725 ( .A(n21243), .B(n21242), .Z(n21577) );
  NANDN U21726 ( .A(n21576), .B(n21577), .Z(n21244) );
  AND U21727 ( .A(n21245), .B(n21244), .Z(n21247) );
  AND U21728 ( .A(a[10]), .B(b[3]), .Z(n21246) );
  NANDN U21729 ( .A(n21247), .B(n21246), .Z(n21251) );
  XOR U21730 ( .A(n21247), .B(n21246), .Z(n21582) );
  XNOR U21731 ( .A(n21249), .B(n21248), .Z(n21583) );
  NANDN U21732 ( .A(n21582), .B(n21583), .Z(n21250) );
  AND U21733 ( .A(n21251), .B(n21250), .Z(n21255) );
  XNOR U21734 ( .A(n21253), .B(n21252), .Z(n21254) );
  NANDN U21735 ( .A(n21255), .B(n21254), .Z(n21257) );
  NAND U21736 ( .A(a[11]), .B(b[3]), .Z(n21588) );
  XNOR U21737 ( .A(n21255), .B(n21254), .Z(n21589) );
  NANDN U21738 ( .A(n21588), .B(n21589), .Z(n21256) );
  AND U21739 ( .A(n21257), .B(n21256), .Z(n21259) );
  AND U21740 ( .A(a[12]), .B(b[3]), .Z(n21258) );
  NANDN U21741 ( .A(n21259), .B(n21258), .Z(n21263) );
  XOR U21742 ( .A(n21259), .B(n21258), .Z(n21594) );
  XNOR U21743 ( .A(n21261), .B(n21260), .Z(n21595) );
  NANDN U21744 ( .A(n21594), .B(n21595), .Z(n21262) );
  AND U21745 ( .A(n21263), .B(n21262), .Z(n21267) );
  XOR U21746 ( .A(n21265), .B(n21264), .Z(n21266) );
  NANDN U21747 ( .A(n21267), .B(n21266), .Z(n21269) );
  NAND U21748 ( .A(a[13]), .B(b[3]), .Z(n21600) );
  XNOR U21749 ( .A(n21267), .B(n21266), .Z(n21601) );
  NANDN U21750 ( .A(n21600), .B(n21601), .Z(n21268) );
  AND U21751 ( .A(n21269), .B(n21268), .Z(n21273) );
  AND U21752 ( .A(a[14]), .B(b[3]), .Z(n21272) );
  NANDN U21753 ( .A(n21273), .B(n21272), .Z(n21275) );
  XNOR U21754 ( .A(n21271), .B(n21270), .Z(n21607) );
  XNOR U21755 ( .A(n21273), .B(n21272), .Z(n21606) );
  NAND U21756 ( .A(n21607), .B(n21606), .Z(n21274) );
  AND U21757 ( .A(n21275), .B(n21274), .Z(n21279) );
  XOR U21758 ( .A(n21277), .B(n21276), .Z(n21278) );
  NANDN U21759 ( .A(n21279), .B(n21278), .Z(n21281) );
  NAND U21760 ( .A(a[15]), .B(b[3]), .Z(n21614) );
  XNOR U21761 ( .A(n21279), .B(n21278), .Z(n21615) );
  NANDN U21762 ( .A(n21614), .B(n21615), .Z(n21280) );
  AND U21763 ( .A(n21281), .B(n21280), .Z(n21285) );
  AND U21764 ( .A(a[16]), .B(b[3]), .Z(n21284) );
  NANDN U21765 ( .A(n21285), .B(n21284), .Z(n21287) );
  XNOR U21766 ( .A(n21283), .B(n21282), .Z(n21525) );
  XNOR U21767 ( .A(n21285), .B(n21284), .Z(n21524) );
  NAND U21768 ( .A(n21525), .B(n21524), .Z(n21286) );
  NAND U21769 ( .A(n21287), .B(n21286), .Z(n21621) );
  NAND U21770 ( .A(a[17]), .B(b[3]), .Z(n21623) );
  AND U21771 ( .A(a[18]), .B(b[3]), .Z(n21292) );
  NANDN U21772 ( .A(n21293), .B(n21292), .Z(n21295) );
  XNOR U21773 ( .A(n21289), .B(n21288), .Z(n21290) );
  XNOR U21774 ( .A(n21291), .B(n21290), .Z(n21523) );
  XNOR U21775 ( .A(n21293), .B(n21292), .Z(n21522) );
  NAND U21776 ( .A(n21523), .B(n21522), .Z(n21294) );
  NAND U21777 ( .A(n21295), .B(n21294), .Z(n21629) );
  NAND U21778 ( .A(a[19]), .B(b[3]), .Z(n21631) );
  AND U21779 ( .A(a[20]), .B(b[3]), .Z(n21300) );
  NANDN U21780 ( .A(n21301), .B(n21300), .Z(n21303) );
  XNOR U21781 ( .A(n21297), .B(n21296), .Z(n21298) );
  XNOR U21782 ( .A(n21299), .B(n21298), .Z(n21521) );
  XNOR U21783 ( .A(n21301), .B(n21300), .Z(n21520) );
  NAND U21784 ( .A(n21521), .B(n21520), .Z(n21302) );
  NAND U21785 ( .A(n21303), .B(n21302), .Z(n21637) );
  NAND U21786 ( .A(a[21]), .B(b[3]), .Z(n21639) );
  AND U21787 ( .A(a[22]), .B(b[3]), .Z(n21308) );
  NANDN U21788 ( .A(n21309), .B(n21308), .Z(n21311) );
  XNOR U21789 ( .A(n21305), .B(n21304), .Z(n21306) );
  XNOR U21790 ( .A(n21307), .B(n21306), .Z(n21519) );
  XNOR U21791 ( .A(n21309), .B(n21308), .Z(n21518) );
  NAND U21792 ( .A(n21519), .B(n21518), .Z(n21310) );
  NAND U21793 ( .A(n21311), .B(n21310), .Z(n21645) );
  NAND U21794 ( .A(a[23]), .B(b[3]), .Z(n21647) );
  AND U21795 ( .A(a[24]), .B(b[3]), .Z(n21316) );
  NANDN U21796 ( .A(n21317), .B(n21316), .Z(n21319) );
  XNOR U21797 ( .A(n21313), .B(n21312), .Z(n21314) );
  XNOR U21798 ( .A(n21315), .B(n21314), .Z(n21517) );
  XNOR U21799 ( .A(n21317), .B(n21316), .Z(n21516) );
  NAND U21800 ( .A(n21517), .B(n21516), .Z(n21318) );
  NAND U21801 ( .A(n21319), .B(n21318), .Z(n21653) );
  AND U21802 ( .A(a[25]), .B(b[3]), .Z(n21655) );
  AND U21803 ( .A(a[26]), .B(b[3]), .Z(n21324) );
  NANDN U21804 ( .A(n21325), .B(n21324), .Z(n21327) );
  XOR U21805 ( .A(n21321), .B(n21320), .Z(n21322) );
  XNOR U21806 ( .A(n21323), .B(n21322), .Z(n21515) );
  XNOR U21807 ( .A(n21325), .B(n21324), .Z(n21514) );
  NAND U21808 ( .A(n21515), .B(n21514), .Z(n21326) );
  NAND U21809 ( .A(n21327), .B(n21326), .Z(n21661) );
  AND U21810 ( .A(a[27]), .B(b[3]), .Z(n21663) );
  AND U21811 ( .A(a[28]), .B(b[3]), .Z(n21332) );
  NANDN U21812 ( .A(n21333), .B(n21332), .Z(n21335) );
  XNOR U21813 ( .A(n21329), .B(n21328), .Z(n21330) );
  XNOR U21814 ( .A(n21331), .B(n21330), .Z(n21667) );
  XNOR U21815 ( .A(n21333), .B(n21332), .Z(n21666) );
  NAND U21816 ( .A(n21667), .B(n21666), .Z(n21334) );
  NAND U21817 ( .A(n21335), .B(n21334), .Z(n21671) );
  NAND U21818 ( .A(a[29]), .B(b[3]), .Z(n21673) );
  AND U21819 ( .A(a[30]), .B(b[3]), .Z(n21340) );
  NANDN U21820 ( .A(n21341), .B(n21340), .Z(n21343) );
  XNOR U21821 ( .A(n21337), .B(n21336), .Z(n21338) );
  XNOR U21822 ( .A(n21339), .B(n21338), .Z(n21513) );
  XNOR U21823 ( .A(n21341), .B(n21340), .Z(n21512) );
  NAND U21824 ( .A(n21513), .B(n21512), .Z(n21342) );
  NAND U21825 ( .A(n21343), .B(n21342), .Z(n21679) );
  NAND U21826 ( .A(a[31]), .B(b[3]), .Z(n21681) );
  AND U21827 ( .A(a[32]), .B(b[3]), .Z(n21348) );
  NANDN U21828 ( .A(n21349), .B(n21348), .Z(n21351) );
  XNOR U21829 ( .A(n21345), .B(n21344), .Z(n21346) );
  XNOR U21830 ( .A(n21347), .B(n21346), .Z(n21511) );
  XNOR U21831 ( .A(n21349), .B(n21348), .Z(n21510) );
  NAND U21832 ( .A(n21511), .B(n21510), .Z(n21350) );
  AND U21833 ( .A(n21351), .B(n21350), .Z(n21686) );
  NAND U21834 ( .A(a[33]), .B(b[3]), .Z(n21689) );
  NANDN U21835 ( .A(n21356), .B(n21357), .Z(n21359) );
  XOR U21836 ( .A(n21353), .B(n21352), .Z(n21354) );
  XNOR U21837 ( .A(n21355), .B(n21354), .Z(n21693) );
  XNOR U21838 ( .A(n21357), .B(n21356), .Z(n21692) );
  NAND U21839 ( .A(n21693), .B(n21692), .Z(n21358) );
  NAND U21840 ( .A(n21359), .B(n21358), .Z(n21697) );
  NAND U21841 ( .A(a[35]), .B(b[3]), .Z(n21699) );
  AND U21842 ( .A(a[36]), .B(b[3]), .Z(n21360) );
  NANDN U21843 ( .A(n21361), .B(n21360), .Z(n21367) );
  XOR U21844 ( .A(n21361), .B(n21360), .Z(n21508) );
  XNOR U21845 ( .A(n21363), .B(n21362), .Z(n21364) );
  XNOR U21846 ( .A(n21365), .B(n21364), .Z(n21509) );
  NANDN U21847 ( .A(n21508), .B(n21509), .Z(n21366) );
  NAND U21848 ( .A(n21367), .B(n21366), .Z(n21703) );
  NAND U21849 ( .A(a[37]), .B(b[3]), .Z(n21705) );
  AND U21850 ( .A(a[38]), .B(b[3]), .Z(n21372) );
  NANDN U21851 ( .A(n21373), .B(n21372), .Z(n21375) );
  XNOR U21852 ( .A(n21369), .B(n21368), .Z(n21370) );
  XNOR U21853 ( .A(n21371), .B(n21370), .Z(n21507) );
  XNOR U21854 ( .A(n21373), .B(n21372), .Z(n21506) );
  NAND U21855 ( .A(n21507), .B(n21506), .Z(n21374) );
  NAND U21856 ( .A(n21375), .B(n21374), .Z(n21713) );
  NAND U21857 ( .A(a[39]), .B(b[3]), .Z(n21715) );
  AND U21858 ( .A(a[40]), .B(b[3]), .Z(n21380) );
  NANDN U21859 ( .A(n21381), .B(n21380), .Z(n21383) );
  XNOR U21860 ( .A(n21377), .B(n21376), .Z(n21378) );
  XNOR U21861 ( .A(n21379), .B(n21378), .Z(n21505) );
  XNOR U21862 ( .A(n21381), .B(n21380), .Z(n21504) );
  NAND U21863 ( .A(n21505), .B(n21504), .Z(n21382) );
  NAND U21864 ( .A(n21383), .B(n21382), .Z(n21721) );
  NAND U21865 ( .A(a[41]), .B(b[3]), .Z(n21723) );
  AND U21866 ( .A(a[42]), .B(b[3]), .Z(n21388) );
  NANDN U21867 ( .A(n21389), .B(n21388), .Z(n21391) );
  XNOR U21868 ( .A(n21385), .B(n21384), .Z(n21386) );
  XNOR U21869 ( .A(n21387), .B(n21386), .Z(n21503) );
  XNOR U21870 ( .A(n21389), .B(n21388), .Z(n21502) );
  NAND U21871 ( .A(n21503), .B(n21502), .Z(n21390) );
  NAND U21872 ( .A(n21391), .B(n21390), .Z(n21729) );
  NAND U21873 ( .A(a[43]), .B(b[3]), .Z(n21731) );
  AND U21874 ( .A(a[44]), .B(b[3]), .Z(n21396) );
  NANDN U21875 ( .A(n21397), .B(n21396), .Z(n21399) );
  XNOR U21876 ( .A(n21393), .B(n21392), .Z(n21394) );
  XNOR U21877 ( .A(n21395), .B(n21394), .Z(n21501) );
  XNOR U21878 ( .A(n21397), .B(n21396), .Z(n21500) );
  NAND U21879 ( .A(n21501), .B(n21500), .Z(n21398) );
  NAND U21880 ( .A(n21399), .B(n21398), .Z(n21737) );
  NAND U21881 ( .A(a[45]), .B(b[3]), .Z(n21739) );
  AND U21882 ( .A(a[46]), .B(b[3]), .Z(n21404) );
  NANDN U21883 ( .A(n21405), .B(n21404), .Z(n21407) );
  XNOR U21884 ( .A(n21401), .B(n21400), .Z(n21402) );
  XNOR U21885 ( .A(n21403), .B(n21402), .Z(n21499) );
  XNOR U21886 ( .A(n21405), .B(n21404), .Z(n21498) );
  NAND U21887 ( .A(n21499), .B(n21498), .Z(n21406) );
  AND U21888 ( .A(n21407), .B(n21406), .Z(n21744) );
  NAND U21889 ( .A(a[47]), .B(b[3]), .Z(n21747) );
  NANDN U21890 ( .A(n21412), .B(n21413), .Z(n21415) );
  XNOR U21891 ( .A(n21409), .B(n21408), .Z(n21410) );
  XNOR U21892 ( .A(n21411), .B(n21410), .Z(n21497) );
  XNOR U21893 ( .A(n21413), .B(n21412), .Z(n21496) );
  NAND U21894 ( .A(n21497), .B(n21496), .Z(n21414) );
  NAND U21895 ( .A(n21415), .B(n21414), .Z(n21753) );
  NAND U21896 ( .A(a[49]), .B(b[3]), .Z(n21755) );
  AND U21897 ( .A(a[50]), .B(b[3]), .Z(n21420) );
  NANDN U21898 ( .A(n21421), .B(n21420), .Z(n21423) );
  XNOR U21899 ( .A(n21417), .B(n21416), .Z(n21418) );
  XNOR U21900 ( .A(n21419), .B(n21418), .Z(n21495) );
  XNOR U21901 ( .A(n21421), .B(n21420), .Z(n21494) );
  NAND U21902 ( .A(n21495), .B(n21494), .Z(n21422) );
  NAND U21903 ( .A(n21423), .B(n21422), .Z(n21761) );
  AND U21904 ( .A(a[51]), .B(b[3]), .Z(n21763) );
  AND U21905 ( .A(a[52]), .B(b[3]), .Z(n21428) );
  NANDN U21906 ( .A(n21429), .B(n21428), .Z(n21431) );
  XNOR U21907 ( .A(n21425), .B(n21424), .Z(n21426) );
  XNOR U21908 ( .A(n21427), .B(n21426), .Z(n21767) );
  XNOR U21909 ( .A(n21429), .B(n21428), .Z(n21766) );
  NAND U21910 ( .A(n21767), .B(n21766), .Z(n21430) );
  NAND U21911 ( .A(n21431), .B(n21430), .Z(n21771) );
  NAND U21912 ( .A(a[53]), .B(b[3]), .Z(n21773) );
  AND U21913 ( .A(a[54]), .B(b[3]), .Z(n21436) );
  NANDN U21914 ( .A(n21437), .B(n21436), .Z(n21439) );
  XNOR U21915 ( .A(n21433), .B(n21432), .Z(n21434) );
  XNOR U21916 ( .A(n21435), .B(n21434), .Z(n21493) );
  XNOR U21917 ( .A(n21437), .B(n21436), .Z(n21492) );
  NAND U21918 ( .A(n21493), .B(n21492), .Z(n21438) );
  NAND U21919 ( .A(n21439), .B(n21438), .Z(n21779) );
  NAND U21920 ( .A(a[55]), .B(b[3]), .Z(n21781) );
  AND U21921 ( .A(a[56]), .B(b[3]), .Z(n21440) );
  IV U21922 ( .A(n21440), .Z(n21785) );
  OR U21923 ( .A(n21784), .B(n21785), .Z(n21447) );
  ANDN U21924 ( .B(n21784), .A(n21440), .Z(n21445) );
  XOR U21925 ( .A(n21442), .B(n21441), .Z(n21443) );
  XNOR U21926 ( .A(n21444), .B(n21443), .Z(n21787) );
  OR U21927 ( .A(n21445), .B(n21787), .Z(n21446) );
  AND U21928 ( .A(n21447), .B(n21446), .Z(n21792) );
  XOR U21929 ( .A(n21449), .B(n21448), .Z(n21450) );
  XOR U21930 ( .A(n21451), .B(n21450), .Z(n21452) );
  IV U21931 ( .A(n21452), .Z(n21791) );
  OR U21932 ( .A(n21792), .B(n21791), .Z(n21455) );
  ANDN U21933 ( .B(n21792), .A(n21452), .Z(n21453) );
  AND U21934 ( .A(a[57]), .B(b[3]), .Z(n21794) );
  NANDN U21935 ( .A(n21453), .B(n21794), .Z(n21454) );
  AND U21936 ( .A(n21455), .B(n21454), .Z(n21796) );
  XOR U21937 ( .A(n21457), .B(n21456), .Z(n21458) );
  XNOR U21938 ( .A(n21459), .B(n21458), .Z(n21798) );
  OR U21939 ( .A(n21805), .B(n21462), .Z(n21465) );
  IV U21940 ( .A(n21462), .Z(n21806) );
  ANDN U21941 ( .B(n21805), .A(n21806), .Z(n21463) );
  NAND U21942 ( .A(a[59]), .B(b[3]), .Z(n21804) );
  NANDN U21943 ( .A(n21463), .B(n21804), .Z(n21464) );
  AND U21944 ( .A(n21465), .B(n21464), .Z(n21467) );
  NANDN U21945 ( .A(n21466), .B(n21467), .Z(n21473) );
  XNOR U21946 ( .A(n21469), .B(n21468), .Z(n21470) );
  XNOR U21947 ( .A(n21471), .B(n21470), .Z(n21810) );
  NAND U21948 ( .A(n21811), .B(n21810), .Z(n21472) );
  AND U21949 ( .A(n21473), .B(n21472), .Z(n21476) );
  NANDN U21950 ( .A(n21476), .B(n21477), .Z(n21479) );
  NAND U21951 ( .A(a[61]), .B(b[3]), .Z(n21816) );
  NANDN U21952 ( .A(n21816), .B(n21817), .Z(n21478) );
  NAND U21953 ( .A(n21479), .B(n21478), .Z(n21825) );
  NANDN U21954 ( .A(n21484), .B(n21485), .Z(n21487) );
  XOR U21955 ( .A(n21481), .B(n21480), .Z(n21482) );
  XOR U21956 ( .A(n21483), .B(n21482), .Z(n21491) );
  XNOR U21957 ( .A(n21485), .B(n21484), .Z(n21490) );
  NANDN U21958 ( .A(n21491), .B(n21490), .Z(n21486) );
  AND U21959 ( .A(n21487), .B(n21486), .Z(n22493) );
  XNOR U21960 ( .A(n21489), .B(n21488), .Z(n22494) );
  XNOR U21961 ( .A(n21491), .B(n21490), .Z(n21830) );
  XNOR U21962 ( .A(n21493), .B(n21492), .Z(n22124) );
  AND U21963 ( .A(a[52]), .B(b[2]), .Z(n21759) );
  XNOR U21964 ( .A(n21495), .B(n21494), .Z(n22104) );
  XNOR U21965 ( .A(n21497), .B(n21496), .Z(n22094) );
  XNOR U21966 ( .A(n21499), .B(n21498), .Z(n22084) );
  XNOR U21967 ( .A(n21501), .B(n21500), .Z(n22074) );
  XNOR U21968 ( .A(n21503), .B(n21502), .Z(n22064) );
  XNOR U21969 ( .A(n21505), .B(n21504), .Z(n22054) );
  XNOR U21970 ( .A(n21507), .B(n21506), .Z(n22044) );
  NAND U21971 ( .A(a[38]), .B(b[2]), .Z(n21706) );
  XNOR U21972 ( .A(n21509), .B(n21508), .Z(n22039) );
  AND U21973 ( .A(a[34]), .B(b[2]), .Z(n21685) );
  XNOR U21974 ( .A(n21511), .B(n21510), .Z(n22018) );
  XNOR U21975 ( .A(n21513), .B(n21512), .Z(n22008) );
  AND U21976 ( .A(a[28]), .B(b[2]), .Z(n21659) );
  XNOR U21977 ( .A(n21515), .B(n21514), .Z(n21988) );
  XNOR U21978 ( .A(n21517), .B(n21516), .Z(n21978) );
  XNOR U21979 ( .A(n21519), .B(n21518), .Z(n21968) );
  XNOR U21980 ( .A(n21521), .B(n21520), .Z(n21962) );
  XNOR U21981 ( .A(n21523), .B(n21522), .Z(n21952) );
  XNOR U21982 ( .A(n21525), .B(n21524), .Z(n21942) );
  XOR U21983 ( .A(n21527), .B(n21526), .Z(n21554) );
  AND U21984 ( .A(a[4]), .B(b[2]), .Z(n21543) );
  AND U21985 ( .A(a[0]), .B(b[2]), .Z(n22172) );
  AND U21986 ( .A(a[1]), .B(b[3]), .Z(n21531) );
  AND U21987 ( .A(n22172), .B(n21531), .Z(n21528) );
  NAND U21988 ( .A(a[2]), .B(n21528), .Z(n21535) );
  NAND U21989 ( .A(b[3]), .B(a[1]), .Z(n21529) );
  XOR U21990 ( .A(n21530), .B(n21529), .Z(n21856) );
  NAND U21991 ( .A(n21531), .B(a[0]), .Z(n21532) );
  XNOR U21992 ( .A(a[2]), .B(n21532), .Z(n21533) );
  AND U21993 ( .A(b[2]), .B(n21533), .Z(n21857) );
  NANDN U21994 ( .A(n21856), .B(n21857), .Z(n21534) );
  AND U21995 ( .A(n21535), .B(n21534), .Z(n21539) );
  XNOR U21996 ( .A(n21537), .B(n21536), .Z(n21538) );
  NANDN U21997 ( .A(n21539), .B(n21538), .Z(n21541) );
  NAND U21998 ( .A(a[3]), .B(b[2]), .Z(n21864) );
  XNOR U21999 ( .A(n21539), .B(n21538), .Z(n21865) );
  NANDN U22000 ( .A(n21864), .B(n21865), .Z(n21540) );
  AND U22001 ( .A(n21541), .B(n21540), .Z(n21542) );
  NANDN U22002 ( .A(n21543), .B(n21542), .Z(n21547) );
  XOR U22003 ( .A(n21543), .B(n21542), .Z(n21846) );
  XOR U22004 ( .A(n21545), .B(n21544), .Z(n21847) );
  OR U22005 ( .A(n21846), .B(n21847), .Z(n21546) );
  NAND U22006 ( .A(n21547), .B(n21546), .Z(n21550) );
  XOR U22007 ( .A(n21549), .B(n21548), .Z(n21551) );
  NANDN U22008 ( .A(n21550), .B(n21551), .Z(n21553) );
  NAND U22009 ( .A(a[5]), .B(b[2]), .Z(n21872) );
  XNOR U22010 ( .A(n21551), .B(n21550), .Z(n21873) );
  NANDN U22011 ( .A(n21872), .B(n21873), .Z(n21552) );
  AND U22012 ( .A(n21553), .B(n21552), .Z(n21555) );
  NANDN U22013 ( .A(n21554), .B(n21555), .Z(n21557) );
  AND U22014 ( .A(a[6]), .B(b[2]), .Z(n21844) );
  NANDN U22015 ( .A(n21844), .B(n21845), .Z(n21556) );
  AND U22016 ( .A(n21557), .B(n21556), .Z(n21561) );
  NAND U22017 ( .A(n21561), .B(n21560), .Z(n21563) );
  NAND U22018 ( .A(a[7]), .B(b[2]), .Z(n21884) );
  XOR U22019 ( .A(n21561), .B(n21560), .Z(n21885) );
  NANDN U22020 ( .A(n21884), .B(n21885), .Z(n21562) );
  AND U22021 ( .A(n21563), .B(n21562), .Z(n21564) );
  AND U22022 ( .A(a[8]), .B(b[2]), .Z(n21565) );
  NANDN U22023 ( .A(n21564), .B(n21565), .Z(n21569) );
  NAND U22024 ( .A(n21889), .B(n21888), .Z(n21568) );
  AND U22025 ( .A(n21569), .B(n21568), .Z(n21572) );
  XOR U22026 ( .A(n21571), .B(n21570), .Z(n21573) );
  NANDN U22027 ( .A(n21572), .B(n21573), .Z(n21575) );
  NAND U22028 ( .A(a[9]), .B(b[2]), .Z(n21894) );
  NANDN U22029 ( .A(n21894), .B(n21895), .Z(n21574) );
  AND U22030 ( .A(n21575), .B(n21574), .Z(n21579) );
  AND U22031 ( .A(a[10]), .B(b[2]), .Z(n21578) );
  NANDN U22032 ( .A(n21579), .B(n21578), .Z(n21581) );
  XOR U22033 ( .A(n21577), .B(n21576), .Z(n21900) );
  XNOR U22034 ( .A(n21579), .B(n21578), .Z(n21901) );
  NANDN U22035 ( .A(n21900), .B(n21901), .Z(n21580) );
  AND U22036 ( .A(n21581), .B(n21580), .Z(n21585) );
  XNOR U22037 ( .A(n21583), .B(n21582), .Z(n21584) );
  NANDN U22038 ( .A(n21585), .B(n21584), .Z(n21587) );
  NAND U22039 ( .A(a[11]), .B(b[2]), .Z(n21906) );
  XNOR U22040 ( .A(n21585), .B(n21584), .Z(n21907) );
  NANDN U22041 ( .A(n21906), .B(n21907), .Z(n21586) );
  AND U22042 ( .A(n21587), .B(n21586), .Z(n21591) );
  AND U22043 ( .A(a[12]), .B(b[2]), .Z(n21590) );
  NANDN U22044 ( .A(n21591), .B(n21590), .Z(n21593) );
  XOR U22045 ( .A(n21589), .B(n21588), .Z(n21912) );
  XNOR U22046 ( .A(n21591), .B(n21590), .Z(n21913) );
  NANDN U22047 ( .A(n21912), .B(n21913), .Z(n21592) );
  AND U22048 ( .A(n21593), .B(n21592), .Z(n21597) );
  XNOR U22049 ( .A(n21595), .B(n21594), .Z(n21596) );
  NANDN U22050 ( .A(n21597), .B(n21596), .Z(n21599) );
  NAND U22051 ( .A(a[13]), .B(b[2]), .Z(n21918) );
  XNOR U22052 ( .A(n21597), .B(n21596), .Z(n21919) );
  NANDN U22053 ( .A(n21918), .B(n21919), .Z(n21598) );
  AND U22054 ( .A(n21599), .B(n21598), .Z(n21603) );
  AND U22055 ( .A(a[14]), .B(b[2]), .Z(n21602) );
  NANDN U22056 ( .A(n21603), .B(n21602), .Z(n21605) );
  XOR U22057 ( .A(n21601), .B(n21600), .Z(n21924) );
  XNOR U22058 ( .A(n21603), .B(n21602), .Z(n21925) );
  NANDN U22059 ( .A(n21924), .B(n21925), .Z(n21604) );
  AND U22060 ( .A(n21605), .B(n21604), .Z(n21609) );
  XOR U22061 ( .A(n21607), .B(n21606), .Z(n21608) );
  NANDN U22062 ( .A(n21609), .B(n21608), .Z(n21611) );
  NAND U22063 ( .A(a[15]), .B(b[2]), .Z(n21930) );
  XNOR U22064 ( .A(n21609), .B(n21608), .Z(n21931) );
  NANDN U22065 ( .A(n21930), .B(n21931), .Z(n21610) );
  AND U22066 ( .A(n21611), .B(n21610), .Z(n21613) );
  AND U22067 ( .A(a[16]), .B(b[2]), .Z(n21612) );
  NANDN U22068 ( .A(n21613), .B(n21612), .Z(n21617) );
  XNOR U22069 ( .A(n21613), .B(n21612), .Z(n21937) );
  XNOR U22070 ( .A(n21615), .B(n21614), .Z(n21936) );
  NAND U22071 ( .A(n21937), .B(n21936), .Z(n21616) );
  NAND U22072 ( .A(n21617), .B(n21616), .Z(n21943) );
  AND U22073 ( .A(a[17]), .B(b[2]), .Z(n21945) );
  AND U22074 ( .A(a[18]), .B(b[2]), .Z(n21618) );
  NANDN U22075 ( .A(n21619), .B(n21618), .Z(n21625) );
  XOR U22076 ( .A(n21619), .B(n21618), .Z(n21946) );
  XNOR U22077 ( .A(n21621), .B(n21620), .Z(n21622) );
  XNOR U22078 ( .A(n21623), .B(n21622), .Z(n21947) );
  NANDN U22079 ( .A(n21946), .B(n21947), .Z(n21624) );
  NAND U22080 ( .A(n21625), .B(n21624), .Z(n21953) );
  AND U22081 ( .A(a[19]), .B(b[2]), .Z(n21955) );
  AND U22082 ( .A(a[20]), .B(b[2]), .Z(n21626) );
  NANDN U22083 ( .A(n21627), .B(n21626), .Z(n21633) );
  XOR U22084 ( .A(n21627), .B(n21626), .Z(n21956) );
  XNOR U22085 ( .A(n21629), .B(n21628), .Z(n21630) );
  XNOR U22086 ( .A(n21631), .B(n21630), .Z(n21957) );
  NANDN U22087 ( .A(n21956), .B(n21957), .Z(n21632) );
  NAND U22088 ( .A(n21633), .B(n21632), .Z(n21963) );
  NAND U22089 ( .A(a[21]), .B(b[2]), .Z(n21965) );
  AND U22090 ( .A(a[22]), .B(b[2]), .Z(n21634) );
  NANDN U22091 ( .A(n21635), .B(n21634), .Z(n21641) );
  XOR U22092 ( .A(n21635), .B(n21634), .Z(n21842) );
  XNOR U22093 ( .A(n21637), .B(n21636), .Z(n21638) );
  XNOR U22094 ( .A(n21639), .B(n21638), .Z(n21843) );
  NANDN U22095 ( .A(n21842), .B(n21843), .Z(n21640) );
  NAND U22096 ( .A(n21641), .B(n21640), .Z(n21969) );
  AND U22097 ( .A(a[23]), .B(b[2]), .Z(n21971) );
  AND U22098 ( .A(a[24]), .B(b[2]), .Z(n21642) );
  NANDN U22099 ( .A(n21643), .B(n21642), .Z(n21649) );
  XOR U22100 ( .A(n21643), .B(n21642), .Z(n21972) );
  XNOR U22101 ( .A(n21645), .B(n21644), .Z(n21646) );
  XNOR U22102 ( .A(n21647), .B(n21646), .Z(n21973) );
  NANDN U22103 ( .A(n21972), .B(n21973), .Z(n21648) );
  NAND U22104 ( .A(n21649), .B(n21648), .Z(n21979) );
  AND U22105 ( .A(a[25]), .B(b[2]), .Z(n21981) );
  AND U22106 ( .A(a[26]), .B(b[2]), .Z(n21650) );
  NANDN U22107 ( .A(n21651), .B(n21650), .Z(n21657) );
  XOR U22108 ( .A(n21651), .B(n21650), .Z(n21982) );
  XOR U22109 ( .A(n21653), .B(n21652), .Z(n21654) );
  XNOR U22110 ( .A(n21655), .B(n21654), .Z(n21983) );
  NANDN U22111 ( .A(n21982), .B(n21983), .Z(n21656) );
  NAND U22112 ( .A(n21657), .B(n21656), .Z(n21989) );
  AND U22113 ( .A(a[27]), .B(b[2]), .Z(n21991) );
  NANDN U22114 ( .A(n21659), .B(n21658), .Z(n21665) );
  XNOR U22115 ( .A(n21659), .B(n21658), .Z(n21992) );
  XNOR U22116 ( .A(n21661), .B(n21660), .Z(n21662) );
  XNOR U22117 ( .A(n21663), .B(n21662), .Z(n21993) );
  NAND U22118 ( .A(n21992), .B(n21993), .Z(n21664) );
  NAND U22119 ( .A(n21665), .B(n21664), .Z(n21999) );
  XOR U22120 ( .A(n21667), .B(n21666), .Z(n21998) );
  NAND U22121 ( .A(a[29]), .B(b[2]), .Z(n22001) );
  AND U22122 ( .A(a[30]), .B(b[2]), .Z(n21668) );
  NANDN U22123 ( .A(n21669), .B(n21668), .Z(n21675) );
  XOR U22124 ( .A(n21669), .B(n21668), .Z(n22002) );
  XNOR U22125 ( .A(n21671), .B(n21670), .Z(n21672) );
  XNOR U22126 ( .A(n21673), .B(n21672), .Z(n22003) );
  NANDN U22127 ( .A(n22002), .B(n22003), .Z(n21674) );
  NAND U22128 ( .A(n21675), .B(n21674), .Z(n22009) );
  AND U22129 ( .A(a[31]), .B(b[2]), .Z(n22011) );
  AND U22130 ( .A(a[32]), .B(b[2]), .Z(n21676) );
  NANDN U22131 ( .A(n21677), .B(n21676), .Z(n21683) );
  XOR U22132 ( .A(n21677), .B(n21676), .Z(n22012) );
  XNOR U22133 ( .A(n21679), .B(n21678), .Z(n21680) );
  XNOR U22134 ( .A(n21681), .B(n21680), .Z(n22013) );
  NANDN U22135 ( .A(n22012), .B(n22013), .Z(n21682) );
  NAND U22136 ( .A(n21683), .B(n21682), .Z(n22019) );
  AND U22137 ( .A(a[33]), .B(b[2]), .Z(n22021) );
  NANDN U22138 ( .A(n21685), .B(n21684), .Z(n21691) );
  XNOR U22139 ( .A(n21685), .B(n21684), .Z(n22022) );
  XOR U22140 ( .A(n21687), .B(n21686), .Z(n21688) );
  XNOR U22141 ( .A(n21689), .B(n21688), .Z(n22023) );
  NAND U22142 ( .A(n22022), .B(n22023), .Z(n21690) );
  NAND U22143 ( .A(n21691), .B(n21690), .Z(n22029) );
  XOR U22144 ( .A(n21693), .B(n21692), .Z(n22028) );
  NAND U22145 ( .A(a[35]), .B(b[2]), .Z(n22031) );
  AND U22146 ( .A(a[36]), .B(b[2]), .Z(n21694) );
  NANDN U22147 ( .A(n21695), .B(n21694), .Z(n21701) );
  XOR U22148 ( .A(n21695), .B(n21694), .Z(n22032) );
  XNOR U22149 ( .A(n21697), .B(n21696), .Z(n21698) );
  XNOR U22150 ( .A(n21699), .B(n21698), .Z(n22033) );
  NANDN U22151 ( .A(n22032), .B(n22033), .Z(n21700) );
  AND U22152 ( .A(n21701), .B(n21700), .Z(n22038) );
  NAND U22153 ( .A(a[37]), .B(b[2]), .Z(n22041) );
  NANDN U22154 ( .A(n21706), .B(n21707), .Z(n21709) );
  XNOR U22155 ( .A(n21703), .B(n21702), .Z(n21704) );
  XNOR U22156 ( .A(n21705), .B(n21704), .Z(n21841) );
  XNOR U22157 ( .A(n21707), .B(n21706), .Z(n21840) );
  NAND U22158 ( .A(n21841), .B(n21840), .Z(n21708) );
  NAND U22159 ( .A(n21709), .B(n21708), .Z(n22045) );
  AND U22160 ( .A(a[39]), .B(b[2]), .Z(n22047) );
  AND U22161 ( .A(a[40]), .B(b[2]), .Z(n21710) );
  NANDN U22162 ( .A(n21711), .B(n21710), .Z(n21717) );
  XOR U22163 ( .A(n21711), .B(n21710), .Z(n22048) );
  XNOR U22164 ( .A(n21713), .B(n21712), .Z(n21714) );
  XNOR U22165 ( .A(n21715), .B(n21714), .Z(n22049) );
  NANDN U22166 ( .A(n22048), .B(n22049), .Z(n21716) );
  NAND U22167 ( .A(n21717), .B(n21716), .Z(n22055) );
  AND U22168 ( .A(a[41]), .B(b[2]), .Z(n22057) );
  AND U22169 ( .A(a[42]), .B(b[2]), .Z(n21718) );
  NANDN U22170 ( .A(n21719), .B(n21718), .Z(n21725) );
  XOR U22171 ( .A(n21719), .B(n21718), .Z(n22058) );
  XNOR U22172 ( .A(n21721), .B(n21720), .Z(n21722) );
  XNOR U22173 ( .A(n21723), .B(n21722), .Z(n22059) );
  NANDN U22174 ( .A(n22058), .B(n22059), .Z(n21724) );
  NAND U22175 ( .A(n21725), .B(n21724), .Z(n22065) );
  AND U22176 ( .A(a[43]), .B(b[2]), .Z(n22067) );
  AND U22177 ( .A(a[44]), .B(b[2]), .Z(n21726) );
  NANDN U22178 ( .A(n21727), .B(n21726), .Z(n21733) );
  XOR U22179 ( .A(n21727), .B(n21726), .Z(n22068) );
  XNOR U22180 ( .A(n21729), .B(n21728), .Z(n21730) );
  XNOR U22181 ( .A(n21731), .B(n21730), .Z(n22069) );
  NANDN U22182 ( .A(n22068), .B(n22069), .Z(n21732) );
  NAND U22183 ( .A(n21733), .B(n21732), .Z(n22075) );
  AND U22184 ( .A(a[45]), .B(b[2]), .Z(n22077) );
  AND U22185 ( .A(a[46]), .B(b[2]), .Z(n21734) );
  NANDN U22186 ( .A(n21735), .B(n21734), .Z(n21741) );
  XOR U22187 ( .A(n21735), .B(n21734), .Z(n22078) );
  XNOR U22188 ( .A(n21737), .B(n21736), .Z(n21738) );
  XNOR U22189 ( .A(n21739), .B(n21738), .Z(n22079) );
  NANDN U22190 ( .A(n22078), .B(n22079), .Z(n21740) );
  NAND U22191 ( .A(n21741), .B(n21740), .Z(n22085) );
  AND U22192 ( .A(a[47]), .B(b[2]), .Z(n22087) );
  AND U22193 ( .A(a[48]), .B(b[2]), .Z(n21742) );
  NANDN U22194 ( .A(n21743), .B(n21742), .Z(n21749) );
  XOR U22195 ( .A(n21743), .B(n21742), .Z(n22088) );
  XNOR U22196 ( .A(n21745), .B(n21744), .Z(n21746) );
  XNOR U22197 ( .A(n21747), .B(n21746), .Z(n22089) );
  NANDN U22198 ( .A(n22088), .B(n22089), .Z(n21748) );
  NAND U22199 ( .A(n21749), .B(n21748), .Z(n22095) );
  AND U22200 ( .A(a[49]), .B(b[2]), .Z(n22097) );
  AND U22201 ( .A(a[50]), .B(b[2]), .Z(n21750) );
  NANDN U22202 ( .A(n21751), .B(n21750), .Z(n21757) );
  XOR U22203 ( .A(n21751), .B(n21750), .Z(n22098) );
  XNOR U22204 ( .A(n21753), .B(n21752), .Z(n21754) );
  XNOR U22205 ( .A(n21755), .B(n21754), .Z(n22099) );
  NANDN U22206 ( .A(n22098), .B(n22099), .Z(n21756) );
  NAND U22207 ( .A(n21757), .B(n21756), .Z(n22105) );
  AND U22208 ( .A(a[51]), .B(b[2]), .Z(n22107) );
  NANDN U22209 ( .A(n21759), .B(n21758), .Z(n21765) );
  XNOR U22210 ( .A(n21759), .B(n21758), .Z(n22108) );
  XNOR U22211 ( .A(n21761), .B(n21760), .Z(n21762) );
  XNOR U22212 ( .A(n21763), .B(n21762), .Z(n22109) );
  NAND U22213 ( .A(n22108), .B(n22109), .Z(n21764) );
  NAND U22214 ( .A(n21765), .B(n21764), .Z(n22115) );
  XOR U22215 ( .A(n21767), .B(n21766), .Z(n22114) );
  NAND U22216 ( .A(a[53]), .B(b[2]), .Z(n22117) );
  AND U22217 ( .A(a[54]), .B(b[2]), .Z(n21768) );
  NANDN U22218 ( .A(n21769), .B(n21768), .Z(n21775) );
  XOR U22219 ( .A(n21769), .B(n21768), .Z(n22118) );
  XNOR U22220 ( .A(n21771), .B(n21770), .Z(n21772) );
  XNOR U22221 ( .A(n21773), .B(n21772), .Z(n22119) );
  NANDN U22222 ( .A(n22118), .B(n22119), .Z(n21774) );
  NAND U22223 ( .A(n21775), .B(n21774), .Z(n22125) );
  AND U22224 ( .A(a[55]), .B(b[2]), .Z(n22127) );
  AND U22225 ( .A(a[56]), .B(b[2]), .Z(n21776) );
  NANDN U22226 ( .A(n21777), .B(n21776), .Z(n21783) );
  XOR U22227 ( .A(n21777), .B(n21776), .Z(n22128) );
  XNOR U22228 ( .A(n21779), .B(n21778), .Z(n21780) );
  XNOR U22229 ( .A(n21781), .B(n21780), .Z(n22129) );
  NANDN U22230 ( .A(n22128), .B(n22129), .Z(n21782) );
  NAND U22231 ( .A(n21783), .B(n21782), .Z(n21788) );
  XOR U22232 ( .A(n21785), .B(n21784), .Z(n21786) );
  XOR U22233 ( .A(n21787), .B(n21786), .Z(n21789) );
  NANDN U22234 ( .A(n21788), .B(n21789), .Z(n22134) );
  NAND U22235 ( .A(a[57]), .B(b[2]), .Z(n22137) );
  NANDN U22236 ( .A(n21789), .B(n21788), .Z(n22135) );
  NAND U22237 ( .A(n22137), .B(n22135), .Z(n21790) );
  NAND U22238 ( .A(n22134), .B(n21790), .Z(n21837) );
  AND U22239 ( .A(a[58]), .B(b[2]), .Z(n21836) );
  XOR U22240 ( .A(n21792), .B(n21791), .Z(n21793) );
  XNOR U22241 ( .A(n21794), .B(n21793), .Z(n21839) );
  XOR U22242 ( .A(n21796), .B(n21795), .Z(n21797) );
  XOR U22243 ( .A(n21798), .B(n21797), .Z(n21799) );
  IV U22244 ( .A(n21799), .Z(n22139) );
  OR U22245 ( .A(n22140), .B(n22139), .Z(n21802) );
  ANDN U22246 ( .B(n22140), .A(n21799), .Z(n21800) );
  AND U22247 ( .A(a[59]), .B(b[2]), .Z(n22142) );
  NANDN U22248 ( .A(n21800), .B(n22142), .Z(n21801) );
  AND U22249 ( .A(n21802), .B(n21801), .Z(n21833) );
  AND U22250 ( .A(a[60]), .B(b[2]), .Z(n21803) );
  IV U22251 ( .A(n21803), .Z(n21832) );
  OR U22252 ( .A(n21833), .B(n21832), .Z(n21809) );
  ANDN U22253 ( .B(n21833), .A(n21803), .Z(n21807) );
  OR U22254 ( .A(n21807), .B(n21835), .Z(n21808) );
  AND U22255 ( .A(n21809), .B(n21808), .Z(n22150) );
  XOR U22256 ( .A(n21811), .B(n21810), .Z(n21812) );
  IV U22257 ( .A(n21812), .Z(n22149) );
  OR U22258 ( .A(n22150), .B(n22149), .Z(n21815) );
  ANDN U22259 ( .B(n22150), .A(n21812), .Z(n21813) );
  AND U22260 ( .A(a[61]), .B(b[2]), .Z(n22148) );
  NANDN U22261 ( .A(n21813), .B(n22148), .Z(n21814) );
  AND U22262 ( .A(n21815), .B(n21814), .Z(n21819) );
  AND U22263 ( .A(a[62]), .B(b[2]), .Z(n21818) );
  NANDN U22264 ( .A(n21819), .B(n21818), .Z(n21821) );
  XNOR U22265 ( .A(n21819), .B(n21818), .Z(n22151) );
  NAND U22266 ( .A(n22152), .B(n22151), .Z(n21820) );
  AND U22267 ( .A(n21821), .B(n21820), .Z(n21827) );
  AND U22268 ( .A(a[63]), .B(b[2]), .Z(n21826) );
  NANDN U22269 ( .A(n21827), .B(n21826), .Z(n21829) );
  XOR U22270 ( .A(n21823), .B(n21822), .Z(n21824) );
  XOR U22271 ( .A(n21825), .B(n21824), .Z(n22158) );
  XNOR U22272 ( .A(n21827), .B(n21826), .Z(n22157) );
  NANDN U22273 ( .A(n22158), .B(n22157), .Z(n21828) );
  AND U22274 ( .A(n21829), .B(n21828), .Z(n21831) );
  ANDN U22275 ( .B(n21830), .A(n21831), .Z(n24663) );
  XNOR U22276 ( .A(n21831), .B(n21830), .Z(n24662) );
  XOR U22277 ( .A(n21833), .B(n21832), .Z(n21834) );
  XOR U22278 ( .A(n21835), .B(n21834), .Z(n22147) );
  AND U22279 ( .A(a[60]), .B(b[1]), .Z(n22138) );
  IV U22280 ( .A(n22138), .Z(n22475) );
  XOR U22281 ( .A(n21837), .B(n21836), .Z(n21838) );
  XOR U22282 ( .A(n21839), .B(n21838), .Z(n22470) );
  AND U22283 ( .A(a[58]), .B(b[1]), .Z(n22461) );
  AND U22284 ( .A(a[56]), .B(b[1]), .Z(n22453) );
  AND U22285 ( .A(a[54]), .B(b[1]), .Z(n22443) );
  AND U22286 ( .A(a[52]), .B(b[1]), .Z(n22433) );
  AND U22287 ( .A(a[50]), .B(b[1]), .Z(n22423) );
  AND U22288 ( .A(a[48]), .B(b[1]), .Z(n22413) );
  AND U22289 ( .A(a[46]), .B(b[1]), .Z(n22403) );
  AND U22290 ( .A(a[44]), .B(b[1]), .Z(n22393) );
  AND U22291 ( .A(a[42]), .B(b[1]), .Z(n22383) );
  AND U22292 ( .A(a[40]), .B(b[1]), .Z(n22373) );
  XOR U22293 ( .A(n21841), .B(n21840), .Z(n22042) );
  AND U22294 ( .A(a[36]), .B(b[1]), .Z(n22353) );
  AND U22295 ( .A(a[34]), .B(b[1]), .Z(n22343) );
  AND U22296 ( .A(a[32]), .B(b[1]), .Z(n22333) );
  AND U22297 ( .A(a[30]), .B(b[1]), .Z(n22323) );
  AND U22298 ( .A(a[28]), .B(b[1]), .Z(n22313) );
  AND U22299 ( .A(a[26]), .B(b[1]), .Z(n22303) );
  AND U22300 ( .A(a[24]), .B(b[1]), .Z(n22293) );
  XNOR U22301 ( .A(n21843), .B(n21842), .Z(n21966) );
  AND U22302 ( .A(a[20]), .B(b[1]), .Z(n22273) );
  AND U22303 ( .A(a[18]), .B(b[1]), .Z(n22263) );
  XOR U22304 ( .A(n21847), .B(n21846), .Z(n21869) );
  AND U22305 ( .A(a[0]), .B(b[1]), .Z(n24972) );
  AND U22306 ( .A(a[1]), .B(b[2]), .Z(n21849) );
  AND U22307 ( .A(n24972), .B(n21849), .Z(n21848) );
  NAND U22308 ( .A(a[2]), .B(n21848), .Z(n21855) );
  NAND U22309 ( .A(n21849), .B(a[0]), .Z(n21850) );
  XNOR U22310 ( .A(a[2]), .B(n21850), .Z(n21851) );
  AND U22311 ( .A(b[1]), .B(n21851), .Z(n22178) );
  NAND U22312 ( .A(b[2]), .B(a[1]), .Z(n21852) );
  XNOR U22313 ( .A(n21853), .B(n21852), .Z(n22177) );
  NAND U22314 ( .A(n22178), .B(n22177), .Z(n21854) );
  AND U22315 ( .A(n21855), .B(n21854), .Z(n21859) );
  XNOR U22316 ( .A(n21857), .B(n21856), .Z(n21858) );
  NANDN U22317 ( .A(n21859), .B(n21858), .Z(n21861) );
  NAND U22318 ( .A(a[3]), .B(b[1]), .Z(n22181) );
  XNOR U22319 ( .A(n21859), .B(n21858), .Z(n22182) );
  NANDN U22320 ( .A(n22181), .B(n22182), .Z(n21860) );
  AND U22321 ( .A(n21861), .B(n21860), .Z(n21863) );
  AND U22322 ( .A(a[4]), .B(b[1]), .Z(n21862) );
  NANDN U22323 ( .A(n21863), .B(n21862), .Z(n21867) );
  XNOR U22324 ( .A(n21863), .B(n21862), .Z(n22190) );
  XNOR U22325 ( .A(n21865), .B(n21864), .Z(n22189) );
  NAND U22326 ( .A(n22190), .B(n22189), .Z(n21866) );
  NAND U22327 ( .A(n21867), .B(n21866), .Z(n21868) );
  NANDN U22328 ( .A(n21869), .B(n21868), .Z(n21871) );
  XNOR U22329 ( .A(n21869), .B(n21868), .Z(n22196) );
  AND U22330 ( .A(a[5]), .B(b[1]), .Z(n22195) );
  NAND U22331 ( .A(n22196), .B(n22195), .Z(n21870) );
  AND U22332 ( .A(n21871), .B(n21870), .Z(n21875) );
  XNOR U22333 ( .A(n21873), .B(n21872), .Z(n21874) );
  NANDN U22334 ( .A(n21875), .B(n21874), .Z(n21877) );
  XNOR U22335 ( .A(n21875), .B(n21874), .Z(n22202) );
  AND U22336 ( .A(a[6]), .B(b[1]), .Z(n22201) );
  NAND U22337 ( .A(n22202), .B(n22201), .Z(n21876) );
  NAND U22338 ( .A(n21877), .B(n21876), .Z(n21878) );
  NAND U22339 ( .A(n21879), .B(n21878), .Z(n21881) );
  NAND U22340 ( .A(a[7]), .B(b[1]), .Z(n22205) );
  XOR U22341 ( .A(n21879), .B(n21878), .Z(n22206) );
  NANDN U22342 ( .A(n22205), .B(n22206), .Z(n21880) );
  AND U22343 ( .A(n21881), .B(n21880), .Z(n21883) );
  AND U22344 ( .A(a[8]), .B(b[1]), .Z(n21882) );
  NANDN U22345 ( .A(n21883), .B(n21882), .Z(n21887) );
  XNOR U22346 ( .A(n21883), .B(n21882), .Z(n22214) );
  NAND U22347 ( .A(n22214), .B(n22213), .Z(n21886) );
  AND U22348 ( .A(n21887), .B(n21886), .Z(n21890) );
  XOR U22349 ( .A(n21889), .B(n21888), .Z(n21891) );
  NANDN U22350 ( .A(n21890), .B(n21891), .Z(n21893) );
  AND U22351 ( .A(a[9]), .B(b[1]), .Z(n22165) );
  NAND U22352 ( .A(n22166), .B(n22165), .Z(n21892) );
  AND U22353 ( .A(n21893), .B(n21892), .Z(n21896) );
  AND U22354 ( .A(a[10]), .B(b[1]), .Z(n21897) );
  NANDN U22355 ( .A(n21896), .B(n21897), .Z(n21899) );
  NAND U22356 ( .A(n22220), .B(n22219), .Z(n21898) );
  AND U22357 ( .A(n21899), .B(n21898), .Z(n21903) );
  XNOR U22358 ( .A(n21901), .B(n21900), .Z(n21902) );
  NANDN U22359 ( .A(n21903), .B(n21902), .Z(n21905) );
  NAND U22360 ( .A(a[11]), .B(b[1]), .Z(n22225) );
  XNOR U22361 ( .A(n21903), .B(n21902), .Z(n22226) );
  NANDN U22362 ( .A(n22225), .B(n22226), .Z(n21904) );
  AND U22363 ( .A(n21905), .B(n21904), .Z(n21909) );
  AND U22364 ( .A(a[12]), .B(b[1]), .Z(n21908) );
  NANDN U22365 ( .A(n21909), .B(n21908), .Z(n21911) );
  XNOR U22366 ( .A(n21907), .B(n21906), .Z(n22232) );
  XNOR U22367 ( .A(n21909), .B(n21908), .Z(n22231) );
  NAND U22368 ( .A(n22232), .B(n22231), .Z(n21910) );
  AND U22369 ( .A(n21911), .B(n21910), .Z(n21915) );
  XNOR U22370 ( .A(n21913), .B(n21912), .Z(n21914) );
  NANDN U22371 ( .A(n21915), .B(n21914), .Z(n21917) );
  NAND U22372 ( .A(a[13]), .B(b[1]), .Z(n22237) );
  XNOR U22373 ( .A(n21915), .B(n21914), .Z(n22238) );
  NANDN U22374 ( .A(n22237), .B(n22238), .Z(n21916) );
  AND U22375 ( .A(n21917), .B(n21916), .Z(n21921) );
  AND U22376 ( .A(a[14]), .B(b[1]), .Z(n21920) );
  NANDN U22377 ( .A(n21921), .B(n21920), .Z(n21923) );
  XNOR U22378 ( .A(n21919), .B(n21918), .Z(n22244) );
  XNOR U22379 ( .A(n21921), .B(n21920), .Z(n22243) );
  NAND U22380 ( .A(n22244), .B(n22243), .Z(n21922) );
  AND U22381 ( .A(n21923), .B(n21922), .Z(n21927) );
  XNOR U22382 ( .A(n21925), .B(n21924), .Z(n21926) );
  NANDN U22383 ( .A(n21927), .B(n21926), .Z(n21929) );
  NAND U22384 ( .A(a[15]), .B(b[1]), .Z(n22249) );
  XNOR U22385 ( .A(n21927), .B(n21926), .Z(n22250) );
  NANDN U22386 ( .A(n22249), .B(n22250), .Z(n21928) );
  AND U22387 ( .A(n21929), .B(n21928), .Z(n21933) );
  AND U22388 ( .A(a[16]), .B(b[1]), .Z(n21932) );
  NANDN U22389 ( .A(n21933), .B(n21932), .Z(n21935) );
  XNOR U22390 ( .A(n21931), .B(n21930), .Z(n22256) );
  XNOR U22391 ( .A(n21933), .B(n21932), .Z(n22255) );
  NAND U22392 ( .A(n22256), .B(n22255), .Z(n21934) );
  AND U22393 ( .A(n21935), .B(n21934), .Z(n21939) );
  XOR U22394 ( .A(n21937), .B(n21936), .Z(n21938) );
  NANDN U22395 ( .A(n21939), .B(n21938), .Z(n21941) );
  NAND U22396 ( .A(a[17]), .B(b[1]), .Z(n22259) );
  XNOR U22397 ( .A(n21939), .B(n21938), .Z(n22260) );
  NANDN U22398 ( .A(n22259), .B(n22260), .Z(n21940) );
  NAND U22399 ( .A(n21941), .B(n21940), .Z(n22264) );
  XNOR U22400 ( .A(n21943), .B(n21942), .Z(n21944) );
  XNOR U22401 ( .A(n21945), .B(n21944), .Z(n22266) );
  XNOR U22402 ( .A(n21947), .B(n21946), .Z(n21948) );
  NANDN U22403 ( .A(n21949), .B(n21948), .Z(n21951) );
  NAND U22404 ( .A(a[19]), .B(b[1]), .Z(n22269) );
  XNOR U22405 ( .A(n21949), .B(n21948), .Z(n22270) );
  NANDN U22406 ( .A(n22269), .B(n22270), .Z(n21950) );
  NAND U22407 ( .A(n21951), .B(n21950), .Z(n22274) );
  XNOR U22408 ( .A(n21953), .B(n21952), .Z(n21954) );
  XNOR U22409 ( .A(n21955), .B(n21954), .Z(n22276) );
  XNOR U22410 ( .A(n21957), .B(n21956), .Z(n21958) );
  NANDN U22411 ( .A(n21959), .B(n21958), .Z(n21961) );
  NAND U22412 ( .A(a[21]), .B(b[1]), .Z(n22279) );
  XNOR U22413 ( .A(n21959), .B(n21958), .Z(n22280) );
  NANDN U22414 ( .A(n22279), .B(n22280), .Z(n21960) );
  AND U22415 ( .A(n21961), .B(n21960), .Z(n22283) );
  NAND U22416 ( .A(a[22]), .B(b[1]), .Z(n22284) );
  XNOR U22417 ( .A(n21963), .B(n21962), .Z(n21964) );
  XNOR U22418 ( .A(n21965), .B(n21964), .Z(n22286) );
  NAND U22419 ( .A(a[23]), .B(b[1]), .Z(n22289) );
  XOR U22420 ( .A(n21967), .B(n21966), .Z(n22290) );
  XNOR U22421 ( .A(n21969), .B(n21968), .Z(n21970) );
  XNOR U22422 ( .A(n21971), .B(n21970), .Z(n22296) );
  XNOR U22423 ( .A(n21973), .B(n21972), .Z(n21974) );
  NANDN U22424 ( .A(n21975), .B(n21974), .Z(n21977) );
  XNOR U22425 ( .A(n21975), .B(n21974), .Z(n22300) );
  AND U22426 ( .A(a[25]), .B(b[1]), .Z(n22299) );
  NAND U22427 ( .A(n22300), .B(n22299), .Z(n21976) );
  NAND U22428 ( .A(n21977), .B(n21976), .Z(n22304) );
  XNOR U22429 ( .A(n21979), .B(n21978), .Z(n21980) );
  XNOR U22430 ( .A(n21981), .B(n21980), .Z(n22306) );
  XNOR U22431 ( .A(n21983), .B(n21982), .Z(n21984) );
  NANDN U22432 ( .A(n21985), .B(n21984), .Z(n21987) );
  NAND U22433 ( .A(a[27]), .B(b[1]), .Z(n22309) );
  XNOR U22434 ( .A(n21985), .B(n21984), .Z(n22310) );
  NANDN U22435 ( .A(n22309), .B(n22310), .Z(n21986) );
  NAND U22436 ( .A(n21987), .B(n21986), .Z(n22314) );
  XNOR U22437 ( .A(n21989), .B(n21988), .Z(n21990) );
  XNOR U22438 ( .A(n21991), .B(n21990), .Z(n22316) );
  XNOR U22439 ( .A(n21993), .B(n21992), .Z(n21994) );
  NANDN U22440 ( .A(n21995), .B(n21994), .Z(n21997) );
  NAND U22441 ( .A(a[29]), .B(b[1]), .Z(n22319) );
  XNOR U22442 ( .A(n21995), .B(n21994), .Z(n22320) );
  NANDN U22443 ( .A(n22319), .B(n22320), .Z(n21996) );
  NAND U22444 ( .A(n21997), .B(n21996), .Z(n22324) );
  XOR U22445 ( .A(n21999), .B(n21998), .Z(n22000) );
  XOR U22446 ( .A(n22001), .B(n22000), .Z(n22326) );
  XNOR U22447 ( .A(n22003), .B(n22002), .Z(n22004) );
  NANDN U22448 ( .A(n22005), .B(n22004), .Z(n22007) );
  XNOR U22449 ( .A(n22005), .B(n22004), .Z(n22330) );
  AND U22450 ( .A(a[31]), .B(b[1]), .Z(n22329) );
  NAND U22451 ( .A(n22330), .B(n22329), .Z(n22006) );
  NAND U22452 ( .A(n22007), .B(n22006), .Z(n22334) );
  XNOR U22453 ( .A(n22009), .B(n22008), .Z(n22010) );
  XNOR U22454 ( .A(n22011), .B(n22010), .Z(n22336) );
  XNOR U22455 ( .A(n22013), .B(n22012), .Z(n22014) );
  NANDN U22456 ( .A(n22015), .B(n22014), .Z(n22017) );
  NAND U22457 ( .A(a[33]), .B(b[1]), .Z(n22339) );
  XNOR U22458 ( .A(n22015), .B(n22014), .Z(n22340) );
  NANDN U22459 ( .A(n22339), .B(n22340), .Z(n22016) );
  NAND U22460 ( .A(n22017), .B(n22016), .Z(n22344) );
  XNOR U22461 ( .A(n22019), .B(n22018), .Z(n22020) );
  XNOR U22462 ( .A(n22021), .B(n22020), .Z(n22346) );
  XNOR U22463 ( .A(n22023), .B(n22022), .Z(n22024) );
  NANDN U22464 ( .A(n22025), .B(n22024), .Z(n22027) );
  NAND U22465 ( .A(a[35]), .B(b[1]), .Z(n22349) );
  XNOR U22466 ( .A(n22025), .B(n22024), .Z(n22350) );
  NANDN U22467 ( .A(n22349), .B(n22350), .Z(n22026) );
  NAND U22468 ( .A(n22027), .B(n22026), .Z(n22354) );
  XOR U22469 ( .A(n22029), .B(n22028), .Z(n22030) );
  XOR U22470 ( .A(n22031), .B(n22030), .Z(n22356) );
  XNOR U22471 ( .A(n22033), .B(n22032), .Z(n22034) );
  NANDN U22472 ( .A(n22035), .B(n22034), .Z(n22037) );
  NAND U22473 ( .A(a[37]), .B(b[1]), .Z(n22359) );
  XNOR U22474 ( .A(n22035), .B(n22034), .Z(n22360) );
  NANDN U22475 ( .A(n22359), .B(n22360), .Z(n22036) );
  AND U22476 ( .A(n22037), .B(n22036), .Z(n22363) );
  NAND U22477 ( .A(a[38]), .B(b[1]), .Z(n22364) );
  XNOR U22478 ( .A(n22039), .B(n22038), .Z(n22040) );
  XNOR U22479 ( .A(n22041), .B(n22040), .Z(n22366) );
  NAND U22480 ( .A(a[39]), .B(b[1]), .Z(n22369) );
  XOR U22481 ( .A(n22043), .B(n22042), .Z(n22370) );
  XNOR U22482 ( .A(n22045), .B(n22044), .Z(n22046) );
  XNOR U22483 ( .A(n22047), .B(n22046), .Z(n22376) );
  XNOR U22484 ( .A(n22049), .B(n22048), .Z(n22050) );
  NANDN U22485 ( .A(n22051), .B(n22050), .Z(n22053) );
  NAND U22486 ( .A(a[41]), .B(b[1]), .Z(n22379) );
  XNOR U22487 ( .A(n22051), .B(n22050), .Z(n22380) );
  NANDN U22488 ( .A(n22379), .B(n22380), .Z(n22052) );
  NAND U22489 ( .A(n22053), .B(n22052), .Z(n22384) );
  XNOR U22490 ( .A(n22055), .B(n22054), .Z(n22056) );
  XNOR U22491 ( .A(n22057), .B(n22056), .Z(n22386) );
  XNOR U22492 ( .A(n22059), .B(n22058), .Z(n22060) );
  NANDN U22493 ( .A(n22061), .B(n22060), .Z(n22063) );
  XNOR U22494 ( .A(n22061), .B(n22060), .Z(n22390) );
  AND U22495 ( .A(a[43]), .B(b[1]), .Z(n22389) );
  NAND U22496 ( .A(n22390), .B(n22389), .Z(n22062) );
  NAND U22497 ( .A(n22063), .B(n22062), .Z(n22394) );
  XNOR U22498 ( .A(n22065), .B(n22064), .Z(n22066) );
  XNOR U22499 ( .A(n22067), .B(n22066), .Z(n22396) );
  XNOR U22500 ( .A(n22069), .B(n22068), .Z(n22070) );
  NANDN U22501 ( .A(n22071), .B(n22070), .Z(n22073) );
  NAND U22502 ( .A(a[45]), .B(b[1]), .Z(n22399) );
  XNOR U22503 ( .A(n22071), .B(n22070), .Z(n22400) );
  NANDN U22504 ( .A(n22399), .B(n22400), .Z(n22072) );
  NAND U22505 ( .A(n22073), .B(n22072), .Z(n22404) );
  XNOR U22506 ( .A(n22075), .B(n22074), .Z(n22076) );
  XNOR U22507 ( .A(n22077), .B(n22076), .Z(n22406) );
  XNOR U22508 ( .A(n22079), .B(n22078), .Z(n22080) );
  NANDN U22509 ( .A(n22081), .B(n22080), .Z(n22083) );
  NAND U22510 ( .A(a[47]), .B(b[1]), .Z(n22409) );
  XNOR U22511 ( .A(n22081), .B(n22080), .Z(n22410) );
  NANDN U22512 ( .A(n22409), .B(n22410), .Z(n22082) );
  NAND U22513 ( .A(n22083), .B(n22082), .Z(n22414) );
  XNOR U22514 ( .A(n22085), .B(n22084), .Z(n22086) );
  XNOR U22515 ( .A(n22087), .B(n22086), .Z(n22416) );
  XNOR U22516 ( .A(n22089), .B(n22088), .Z(n22090) );
  NANDN U22517 ( .A(n22091), .B(n22090), .Z(n22093) );
  NAND U22518 ( .A(a[49]), .B(b[1]), .Z(n22419) );
  XNOR U22519 ( .A(n22091), .B(n22090), .Z(n22420) );
  NANDN U22520 ( .A(n22419), .B(n22420), .Z(n22092) );
  NAND U22521 ( .A(n22093), .B(n22092), .Z(n22424) );
  XNOR U22522 ( .A(n22095), .B(n22094), .Z(n22096) );
  XNOR U22523 ( .A(n22097), .B(n22096), .Z(n22426) );
  XNOR U22524 ( .A(n22099), .B(n22098), .Z(n22100) );
  NANDN U22525 ( .A(n22101), .B(n22100), .Z(n22103) );
  XNOR U22526 ( .A(n22101), .B(n22100), .Z(n22430) );
  AND U22527 ( .A(a[51]), .B(b[1]), .Z(n22429) );
  NAND U22528 ( .A(n22430), .B(n22429), .Z(n22102) );
  NAND U22529 ( .A(n22103), .B(n22102), .Z(n22434) );
  XNOR U22530 ( .A(n22105), .B(n22104), .Z(n22106) );
  XNOR U22531 ( .A(n22107), .B(n22106), .Z(n22436) );
  XNOR U22532 ( .A(n22109), .B(n22108), .Z(n22110) );
  NANDN U22533 ( .A(n22111), .B(n22110), .Z(n22113) );
  NAND U22534 ( .A(a[53]), .B(b[1]), .Z(n22439) );
  XNOR U22535 ( .A(n22111), .B(n22110), .Z(n22440) );
  NANDN U22536 ( .A(n22439), .B(n22440), .Z(n22112) );
  NAND U22537 ( .A(n22113), .B(n22112), .Z(n22444) );
  XOR U22538 ( .A(n22115), .B(n22114), .Z(n22116) );
  XOR U22539 ( .A(n22117), .B(n22116), .Z(n22446) );
  XNOR U22540 ( .A(n22119), .B(n22118), .Z(n22120) );
  NANDN U22541 ( .A(n22121), .B(n22120), .Z(n22123) );
  XNOR U22542 ( .A(n22121), .B(n22120), .Z(n22450) );
  AND U22543 ( .A(a[55]), .B(b[1]), .Z(n22449) );
  NAND U22544 ( .A(n22450), .B(n22449), .Z(n22122) );
  NAND U22545 ( .A(n22123), .B(n22122), .Z(n22454) );
  XNOR U22546 ( .A(n22125), .B(n22124), .Z(n22126) );
  XNOR U22547 ( .A(n22127), .B(n22126), .Z(n22456) );
  XNOR U22548 ( .A(n22129), .B(n22128), .Z(n22130) );
  NANDN U22549 ( .A(n22131), .B(n22130), .Z(n22133) );
  NAND U22550 ( .A(a[57]), .B(b[1]), .Z(n22459) );
  XNOR U22551 ( .A(n22131), .B(n22130), .Z(n22460) );
  NANDN U22552 ( .A(n22459), .B(n22460), .Z(n22132) );
  NAND U22553 ( .A(n22133), .B(n22132), .Z(n22462) );
  NAND U22554 ( .A(n22135), .B(n22134), .Z(n22136) );
  XOR U22555 ( .A(n22137), .B(n22136), .Z(n22464) );
  NAND U22556 ( .A(a[59]), .B(b[1]), .Z(n22472) );
  NANDN U22557 ( .A(n22475), .B(n22476), .Z(n22145) );
  NOR U22558 ( .A(n22138), .B(n22476), .Z(n22143) );
  XOR U22559 ( .A(n22140), .B(n22139), .Z(n22141) );
  XNOR U22560 ( .A(n22142), .B(n22141), .Z(n22478) );
  OR U22561 ( .A(n22143), .B(n22478), .Z(n22144) );
  AND U22562 ( .A(n22145), .B(n22144), .Z(n22146) );
  AND U22563 ( .A(a[61]), .B(b[1]), .Z(n22164) );
  XOR U22564 ( .A(n22147), .B(n22146), .Z(n22163) );
  AND U22565 ( .A(a[62]), .B(b[1]), .Z(n22483) );
  XOR U22566 ( .A(n22152), .B(n22151), .Z(n22153) );
  IV U22567 ( .A(n22153), .Z(n22159) );
  OR U22568 ( .A(n22160), .B(n22159), .Z(n22156) );
  ANDN U22569 ( .B(n22160), .A(n22153), .Z(n22154) );
  NAND U22570 ( .A(a[63]), .B(b[1]), .Z(n22162) );
  OR U22571 ( .A(n22154), .B(n22162), .Z(n22155) );
  AND U22572 ( .A(n22156), .B(n22155), .Z(n22490) );
  XNOR U22573 ( .A(n22158), .B(n22157), .Z(n22489) );
  NANDN U22574 ( .A(n22490), .B(n22489), .Z(n22492) );
  XOR U22575 ( .A(n22160), .B(n22159), .Z(n22161) );
  XNOR U22576 ( .A(n22162), .B(n22161), .Z(n24960) );
  XOR U22577 ( .A(n22164), .B(n22163), .Z(n24956) );
  AND U22578 ( .A(a[59]), .B(b[0]), .Z(n22466) );
  NAND U22579 ( .A(a[58]), .B(b[0]), .Z(n24940) );
  AND U22580 ( .A(a[57]), .B(b[0]), .Z(n22452) );
  AND U22581 ( .A(a[56]), .B(b[0]), .Z(n24934) );
  AND U22582 ( .A(a[53]), .B(b[0]), .Z(n22432) );
  AND U22583 ( .A(a[52]), .B(b[0]), .Z(n24922) );
  AND U22584 ( .A(a[45]), .B(b[0]), .Z(n22392) );
  AND U22585 ( .A(a[44]), .B(b[0]), .Z(n24896) );
  AND U22586 ( .A(a[33]), .B(b[0]), .Z(n22332) );
  AND U22587 ( .A(a[32]), .B(b[0]), .Z(n24858) );
  AND U22588 ( .A(a[29]), .B(b[0]), .Z(n22312) );
  NAND U22589 ( .A(a[28]), .B(b[0]), .Z(n24844) );
  AND U22590 ( .A(a[27]), .B(b[0]), .Z(n22302) );
  AND U22591 ( .A(a[26]), .B(b[0]), .Z(n24838) );
  AND U22592 ( .A(a[25]), .B(b[0]), .Z(n22292) );
  NAND U22593 ( .A(a[24]), .B(b[0]), .Z(n24832) );
  AND U22594 ( .A(a[19]), .B(b[0]), .Z(n22262) );
  NAND U22595 ( .A(a[18]), .B(b[0]), .Z(n24812) );
  AND U22596 ( .A(a[17]), .B(b[0]), .Z(n22254) );
  AND U22597 ( .A(a[15]), .B(b[0]), .Z(n22242) );
  AND U22598 ( .A(a[13]), .B(b[0]), .Z(n22230) );
  AND U22599 ( .A(a[11]), .B(b[0]), .Z(n22217) );
  XOR U22600 ( .A(n22166), .B(n22165), .Z(n24966) );
  AND U22601 ( .A(a[10]), .B(b[0]), .Z(n24965) );
  AND U22602 ( .A(a[9]), .B(b[0]), .Z(n22212) );
  AND U22603 ( .A(a[7]), .B(b[0]), .Z(n22200) );
  AND U22604 ( .A(a[5]), .B(b[0]), .Z(n22188) );
  AND U22605 ( .A(a[3]), .B(b[0]), .Z(n22176) );
  AND U22606 ( .A(b[1]), .B(a[1]), .Z(n22171) );
  AND U22607 ( .A(a[0]), .B(b[0]), .Z(c[0]) );
  NAND U22608 ( .A(n22171), .B(c[0]), .Z(n22168) );
  NAND U22609 ( .A(a[2]), .B(b[0]), .Z(n22167) );
  AND U22610 ( .A(n22168), .B(n22167), .Z(n22174) );
  XNOR U22611 ( .A(a[2]), .B(n22168), .Z(n22170) );
  NANDN U22612 ( .A(b[0]), .B(a[2]), .Z(n22169) );
  NAND U22613 ( .A(n22170), .B(n22169), .Z(n24797) );
  XNOR U22614 ( .A(n22172), .B(n22171), .Z(n24798) );
  NANDN U22615 ( .A(n24797), .B(n24798), .Z(n22173) );
  NANDN U22616 ( .A(n22174), .B(n22173), .Z(n22175) );
  NANDN U22617 ( .A(n22176), .B(n22175), .Z(n22180) );
  XNOR U22618 ( .A(n22176), .B(n22175), .Z(n24824) );
  XNOR U22619 ( .A(n22178), .B(n22177), .Z(n24823) );
  NAND U22620 ( .A(n24824), .B(n24823), .Z(n22179) );
  NAND U22621 ( .A(n22180), .B(n22179), .Z(n22183) );
  XNOR U22622 ( .A(n22182), .B(n22181), .Z(n22184) );
  NANDN U22623 ( .A(n22183), .B(n22184), .Z(n22186) );
  XNOR U22624 ( .A(n22184), .B(n22183), .Z(n24856) );
  AND U22625 ( .A(a[4]), .B(b[0]), .Z(n24855) );
  NAND U22626 ( .A(n24856), .B(n24855), .Z(n22185) );
  AND U22627 ( .A(n22186), .B(n22185), .Z(n22187) );
  NANDN U22628 ( .A(n22188), .B(n22187), .Z(n22192) );
  XNOR U22629 ( .A(n22188), .B(n22187), .Z(n24888) );
  XNOR U22630 ( .A(n22190), .B(n22189), .Z(n24887) );
  NAND U22631 ( .A(n24888), .B(n24887), .Z(n22191) );
  AND U22632 ( .A(n22192), .B(n22191), .Z(n22194) );
  NAND U22633 ( .A(a[6]), .B(b[0]), .Z(n22193) );
  NANDN U22634 ( .A(n22194), .B(n22193), .Z(n22198) );
  XNOR U22635 ( .A(n22194), .B(n22193), .Z(n24920) );
  XNOR U22636 ( .A(n22196), .B(n22195), .Z(n24919) );
  NAND U22637 ( .A(n24920), .B(n24919), .Z(n22197) );
  NAND U22638 ( .A(n22198), .B(n22197), .Z(n22199) );
  NANDN U22639 ( .A(n22200), .B(n22199), .Z(n22204) );
  XNOR U22640 ( .A(n22200), .B(n22199), .Z(n24952) );
  XNOR U22641 ( .A(n22202), .B(n22201), .Z(n24951) );
  NAND U22642 ( .A(n24952), .B(n24951), .Z(n22203) );
  NAND U22643 ( .A(n22204), .B(n22203), .Z(n22207) );
  AND U22644 ( .A(a[8]), .B(b[0]), .Z(n22208) );
  NANDN U22645 ( .A(n22207), .B(n22208), .Z(n22210) );
  XNOR U22646 ( .A(n22206), .B(n22205), .Z(n24962) );
  XNOR U22647 ( .A(n22208), .B(n22207), .Z(n24961) );
  NAND U22648 ( .A(n24962), .B(n24961), .Z(n22209) );
  AND U22649 ( .A(n22210), .B(n22209), .Z(n22211) );
  NANDN U22650 ( .A(n22212), .B(n22211), .Z(n22216) );
  XNOR U22651 ( .A(n22212), .B(n22211), .Z(n24964) );
  XNOR U22652 ( .A(n22214), .B(n22213), .Z(n24963) );
  NAND U22653 ( .A(n24964), .B(n24963), .Z(n22215) );
  NAND U22654 ( .A(n22216), .B(n22215), .Z(n24968) );
  NANDN U22655 ( .A(n22217), .B(n22218), .Z(n22222) );
  XNOR U22656 ( .A(n22220), .B(n22219), .Z(n24969) );
  NAND U22657 ( .A(n24970), .B(n24969), .Z(n22221) );
  NAND U22658 ( .A(n22222), .B(n22221), .Z(n22223) );
  AND U22659 ( .A(a[12]), .B(b[0]), .Z(n22224) );
  NANDN U22660 ( .A(n22223), .B(n22224), .Z(n22228) );
  XNOR U22661 ( .A(n22224), .B(n22223), .Z(n24800) );
  XNOR U22662 ( .A(n22226), .B(n22225), .Z(n24799) );
  NAND U22663 ( .A(n24800), .B(n24799), .Z(n22227) );
  AND U22664 ( .A(n22228), .B(n22227), .Z(n22229) );
  NANDN U22665 ( .A(n22230), .B(n22229), .Z(n22234) );
  XNOR U22666 ( .A(n22230), .B(n22229), .Z(n24802) );
  XNOR U22667 ( .A(n22232), .B(n22231), .Z(n24801) );
  NAND U22668 ( .A(n24802), .B(n24801), .Z(n22233) );
  NAND U22669 ( .A(n22234), .B(n22233), .Z(n22235) );
  AND U22670 ( .A(a[14]), .B(b[0]), .Z(n22236) );
  NANDN U22671 ( .A(n22235), .B(n22236), .Z(n22240) );
  XNOR U22672 ( .A(n22236), .B(n22235), .Z(n24804) );
  XNOR U22673 ( .A(n22238), .B(n22237), .Z(n24803) );
  NAND U22674 ( .A(n24804), .B(n24803), .Z(n22239) );
  AND U22675 ( .A(n22240), .B(n22239), .Z(n22241) );
  NANDN U22676 ( .A(n22242), .B(n22241), .Z(n22246) );
  XNOR U22677 ( .A(n22242), .B(n22241), .Z(n24806) );
  XNOR U22678 ( .A(n22244), .B(n22243), .Z(n24805) );
  NAND U22679 ( .A(n24806), .B(n24805), .Z(n22245) );
  NAND U22680 ( .A(n22246), .B(n22245), .Z(n22247) );
  AND U22681 ( .A(a[16]), .B(b[0]), .Z(n22248) );
  NANDN U22682 ( .A(n22247), .B(n22248), .Z(n22252) );
  XNOR U22683 ( .A(n22248), .B(n22247), .Z(n24808) );
  XNOR U22684 ( .A(n22250), .B(n22249), .Z(n24807) );
  NAND U22685 ( .A(n24808), .B(n24807), .Z(n22251) );
  AND U22686 ( .A(n22252), .B(n22251), .Z(n22253) );
  NANDN U22687 ( .A(n22254), .B(n22253), .Z(n22258) );
  XNOR U22688 ( .A(n22254), .B(n22253), .Z(n24810) );
  XNOR U22689 ( .A(n22256), .B(n22255), .Z(n24809) );
  NAND U22690 ( .A(n24810), .B(n24809), .Z(n22257) );
  AND U22691 ( .A(n22258), .B(n22257), .Z(n24811) );
  XNOR U22692 ( .A(n22260), .B(n22259), .Z(n24814) );
  NANDN U22693 ( .A(n22262), .B(n22261), .Z(n22268) );
  XNOR U22694 ( .A(n22262), .B(n22261), .Z(n24816) );
  XOR U22695 ( .A(n22264), .B(n22263), .Z(n22265) );
  XOR U22696 ( .A(n22266), .B(n22265), .Z(n24815) );
  NAND U22697 ( .A(n24816), .B(n24815), .Z(n22267) );
  AND U22698 ( .A(n22268), .B(n22267), .Z(n24818) );
  NAND U22699 ( .A(a[20]), .B(b[0]), .Z(n24817) );
  XNOR U22700 ( .A(n22270), .B(n22269), .Z(n24820) );
  NAND U22701 ( .A(a[21]), .B(b[0]), .Z(n22271) );
  NANDN U22702 ( .A(n22272), .B(n22271), .Z(n22278) );
  XNOR U22703 ( .A(n22272), .B(n22271), .Z(n24822) );
  XOR U22704 ( .A(n22274), .B(n22273), .Z(n22275) );
  XOR U22705 ( .A(n22276), .B(n22275), .Z(n24821) );
  NAND U22706 ( .A(n24822), .B(n24821), .Z(n22277) );
  AND U22707 ( .A(n22278), .B(n22277), .Z(n24826) );
  NAND U22708 ( .A(a[22]), .B(b[0]), .Z(n24825) );
  XNOR U22709 ( .A(n22280), .B(n22279), .Z(n24828) );
  NAND U22710 ( .A(a[23]), .B(b[0]), .Z(n22281) );
  NANDN U22711 ( .A(n22282), .B(n22281), .Z(n22288) );
  XNOR U22712 ( .A(n22282), .B(n22281), .Z(n24830) );
  XOR U22713 ( .A(n22284), .B(n22283), .Z(n22285) );
  XNOR U22714 ( .A(n22286), .B(n22285), .Z(n24829) );
  NAND U22715 ( .A(n24830), .B(n24829), .Z(n22287) );
  AND U22716 ( .A(n22288), .B(n22287), .Z(n24831) );
  XNOR U22717 ( .A(n22290), .B(n22289), .Z(n24834) );
  NANDN U22718 ( .A(n22292), .B(n22291), .Z(n22298) );
  XNOR U22719 ( .A(n22292), .B(n22291), .Z(n24836) );
  XOR U22720 ( .A(n22294), .B(n22293), .Z(n22295) );
  XOR U22721 ( .A(n22296), .B(n22295), .Z(n24835) );
  NAND U22722 ( .A(n24836), .B(n24835), .Z(n22297) );
  AND U22723 ( .A(n22298), .B(n22297), .Z(n24837) );
  XNOR U22724 ( .A(n22300), .B(n22299), .Z(n24840) );
  NANDN U22725 ( .A(n22302), .B(n22301), .Z(n22308) );
  XNOR U22726 ( .A(n22302), .B(n22301), .Z(n24842) );
  XOR U22727 ( .A(n22304), .B(n22303), .Z(n22305) );
  XOR U22728 ( .A(n22306), .B(n22305), .Z(n24841) );
  NAND U22729 ( .A(n24842), .B(n24841), .Z(n22307) );
  AND U22730 ( .A(n22308), .B(n22307), .Z(n24843) );
  XNOR U22731 ( .A(n22310), .B(n22309), .Z(n24846) );
  NANDN U22732 ( .A(n22312), .B(n22311), .Z(n22318) );
  XNOR U22733 ( .A(n22312), .B(n22311), .Z(n24848) );
  XOR U22734 ( .A(n22314), .B(n22313), .Z(n22315) );
  XOR U22735 ( .A(n22316), .B(n22315), .Z(n24847) );
  NAND U22736 ( .A(n24848), .B(n24847), .Z(n22317) );
  AND U22737 ( .A(n22318), .B(n22317), .Z(n24850) );
  NAND U22738 ( .A(a[30]), .B(b[0]), .Z(n24849) );
  XNOR U22739 ( .A(n22320), .B(n22319), .Z(n24852) );
  NAND U22740 ( .A(a[31]), .B(b[0]), .Z(n22321) );
  NANDN U22741 ( .A(n22322), .B(n22321), .Z(n22328) );
  XNOR U22742 ( .A(n22322), .B(n22321), .Z(n24854) );
  XOR U22743 ( .A(n22324), .B(n22323), .Z(n22325) );
  XNOR U22744 ( .A(n22326), .B(n22325), .Z(n24853) );
  NAND U22745 ( .A(n24854), .B(n24853), .Z(n22327) );
  AND U22746 ( .A(n22328), .B(n22327), .Z(n24857) );
  XNOR U22747 ( .A(n22330), .B(n22329), .Z(n24860) );
  NANDN U22748 ( .A(n22332), .B(n22331), .Z(n22338) );
  XNOR U22749 ( .A(n22332), .B(n22331), .Z(n24862) );
  XOR U22750 ( .A(n22334), .B(n22333), .Z(n22335) );
  XOR U22751 ( .A(n22336), .B(n22335), .Z(n24861) );
  NAND U22752 ( .A(n24862), .B(n24861), .Z(n22337) );
  AND U22753 ( .A(n22338), .B(n22337), .Z(n24864) );
  NAND U22754 ( .A(a[34]), .B(b[0]), .Z(n24863) );
  XNOR U22755 ( .A(n22340), .B(n22339), .Z(n24866) );
  NAND U22756 ( .A(a[35]), .B(b[0]), .Z(n22341) );
  NANDN U22757 ( .A(n22342), .B(n22341), .Z(n22348) );
  XNOR U22758 ( .A(n22342), .B(n22341), .Z(n24868) );
  XOR U22759 ( .A(n22344), .B(n22343), .Z(n22345) );
  XOR U22760 ( .A(n22346), .B(n22345), .Z(n24867) );
  NAND U22761 ( .A(n24868), .B(n24867), .Z(n22347) );
  AND U22762 ( .A(n22348), .B(n22347), .Z(n24870) );
  NAND U22763 ( .A(a[36]), .B(b[0]), .Z(n24869) );
  XNOR U22764 ( .A(n22350), .B(n22349), .Z(n24872) );
  NAND U22765 ( .A(a[37]), .B(b[0]), .Z(n22351) );
  NANDN U22766 ( .A(n22352), .B(n22351), .Z(n22358) );
  XNOR U22767 ( .A(n22352), .B(n22351), .Z(n24874) );
  XOR U22768 ( .A(n22354), .B(n22353), .Z(n22355) );
  XNOR U22769 ( .A(n22356), .B(n22355), .Z(n24873) );
  NAND U22770 ( .A(n24874), .B(n24873), .Z(n22357) );
  AND U22771 ( .A(n22358), .B(n22357), .Z(n24876) );
  NAND U22772 ( .A(a[38]), .B(b[0]), .Z(n24875) );
  XNOR U22773 ( .A(n22360), .B(n22359), .Z(n24878) );
  NAND U22774 ( .A(a[39]), .B(b[0]), .Z(n22361) );
  NANDN U22775 ( .A(n22362), .B(n22361), .Z(n22368) );
  XNOR U22776 ( .A(n22362), .B(n22361), .Z(n24880) );
  XOR U22777 ( .A(n22364), .B(n22363), .Z(n22365) );
  XNOR U22778 ( .A(n22366), .B(n22365), .Z(n24879) );
  NAND U22779 ( .A(n24880), .B(n24879), .Z(n22367) );
  AND U22780 ( .A(n22368), .B(n22367), .Z(n24882) );
  NAND U22781 ( .A(a[40]), .B(b[0]), .Z(n24881) );
  XNOR U22782 ( .A(n22370), .B(n22369), .Z(n24884) );
  NAND U22783 ( .A(a[41]), .B(b[0]), .Z(n22371) );
  NANDN U22784 ( .A(n22372), .B(n22371), .Z(n22378) );
  XNOR U22785 ( .A(n22372), .B(n22371), .Z(n24886) );
  XOR U22786 ( .A(n22374), .B(n22373), .Z(n22375) );
  XOR U22787 ( .A(n22376), .B(n22375), .Z(n24885) );
  NAND U22788 ( .A(n24886), .B(n24885), .Z(n22377) );
  AND U22789 ( .A(n22378), .B(n22377), .Z(n24890) );
  NAND U22790 ( .A(a[42]), .B(b[0]), .Z(n24889) );
  XNOR U22791 ( .A(n22380), .B(n22379), .Z(n24892) );
  NAND U22792 ( .A(a[43]), .B(b[0]), .Z(n22381) );
  NANDN U22793 ( .A(n22382), .B(n22381), .Z(n22388) );
  XNOR U22794 ( .A(n22382), .B(n22381), .Z(n24894) );
  XOR U22795 ( .A(n22384), .B(n22383), .Z(n22385) );
  XOR U22796 ( .A(n22386), .B(n22385), .Z(n24893) );
  NAND U22797 ( .A(n24894), .B(n24893), .Z(n22387) );
  AND U22798 ( .A(n22388), .B(n22387), .Z(n24895) );
  XNOR U22799 ( .A(n22390), .B(n22389), .Z(n24898) );
  NANDN U22800 ( .A(n22392), .B(n22391), .Z(n22398) );
  XNOR U22801 ( .A(n22392), .B(n22391), .Z(n24900) );
  XOR U22802 ( .A(n22394), .B(n22393), .Z(n22395) );
  XOR U22803 ( .A(n22396), .B(n22395), .Z(n24899) );
  NAND U22804 ( .A(n24900), .B(n24899), .Z(n22397) );
  AND U22805 ( .A(n22398), .B(n22397), .Z(n24902) );
  NAND U22806 ( .A(a[46]), .B(b[0]), .Z(n24901) );
  XNOR U22807 ( .A(n22400), .B(n22399), .Z(n24904) );
  NAND U22808 ( .A(a[47]), .B(b[0]), .Z(n22401) );
  NANDN U22809 ( .A(n22402), .B(n22401), .Z(n22408) );
  XNOR U22810 ( .A(n22402), .B(n22401), .Z(n24906) );
  XOR U22811 ( .A(n22404), .B(n22403), .Z(n22405) );
  XOR U22812 ( .A(n22406), .B(n22405), .Z(n24905) );
  NAND U22813 ( .A(n24906), .B(n24905), .Z(n22407) );
  AND U22814 ( .A(n22408), .B(n22407), .Z(n24908) );
  NAND U22815 ( .A(a[48]), .B(b[0]), .Z(n24907) );
  XNOR U22816 ( .A(n22410), .B(n22409), .Z(n24910) );
  NAND U22817 ( .A(a[49]), .B(b[0]), .Z(n22411) );
  NANDN U22818 ( .A(n22412), .B(n22411), .Z(n22418) );
  XNOR U22819 ( .A(n22412), .B(n22411), .Z(n24912) );
  XOR U22820 ( .A(n22414), .B(n22413), .Z(n22415) );
  XOR U22821 ( .A(n22416), .B(n22415), .Z(n24911) );
  NAND U22822 ( .A(n24912), .B(n24911), .Z(n22417) );
  AND U22823 ( .A(n22418), .B(n22417), .Z(n24914) );
  NAND U22824 ( .A(a[50]), .B(b[0]), .Z(n24913) );
  XNOR U22825 ( .A(n22420), .B(n22419), .Z(n24916) );
  NAND U22826 ( .A(a[51]), .B(b[0]), .Z(n22421) );
  NANDN U22827 ( .A(n22422), .B(n22421), .Z(n22428) );
  XNOR U22828 ( .A(n22422), .B(n22421), .Z(n24918) );
  XOR U22829 ( .A(n22424), .B(n22423), .Z(n22425) );
  XOR U22830 ( .A(n22426), .B(n22425), .Z(n24917) );
  NAND U22831 ( .A(n24918), .B(n24917), .Z(n22427) );
  AND U22832 ( .A(n22428), .B(n22427), .Z(n24921) );
  XNOR U22833 ( .A(n22430), .B(n22429), .Z(n24924) );
  NANDN U22834 ( .A(n22432), .B(n22431), .Z(n22438) );
  XNOR U22835 ( .A(n22432), .B(n22431), .Z(n24926) );
  XOR U22836 ( .A(n22434), .B(n22433), .Z(n22435) );
  XOR U22837 ( .A(n22436), .B(n22435), .Z(n24925) );
  NAND U22838 ( .A(n24926), .B(n24925), .Z(n22437) );
  AND U22839 ( .A(n22438), .B(n22437), .Z(n24928) );
  NAND U22840 ( .A(a[54]), .B(b[0]), .Z(n24927) );
  XNOR U22841 ( .A(n22440), .B(n22439), .Z(n24930) );
  NAND U22842 ( .A(a[55]), .B(b[0]), .Z(n22441) );
  NANDN U22843 ( .A(n22442), .B(n22441), .Z(n22448) );
  XNOR U22844 ( .A(n22442), .B(n22441), .Z(n24932) );
  XOR U22845 ( .A(n22444), .B(n22443), .Z(n22445) );
  XNOR U22846 ( .A(n22446), .B(n22445), .Z(n24931) );
  NAND U22847 ( .A(n24932), .B(n24931), .Z(n22447) );
  AND U22848 ( .A(n22448), .B(n22447), .Z(n24933) );
  XNOR U22849 ( .A(n22450), .B(n22449), .Z(n24936) );
  NANDN U22850 ( .A(n22452), .B(n22451), .Z(n22458) );
  XNOR U22851 ( .A(n22452), .B(n22451), .Z(n24938) );
  XOR U22852 ( .A(n22454), .B(n22453), .Z(n22455) );
  XOR U22853 ( .A(n22456), .B(n22455), .Z(n24937) );
  NAND U22854 ( .A(n24938), .B(n24937), .Z(n22457) );
  AND U22855 ( .A(n22458), .B(n22457), .Z(n24939) );
  XNOR U22856 ( .A(n22460), .B(n22459), .Z(n24942) );
  NANDN U22857 ( .A(n22466), .B(n22465), .Z(n22468) );
  XOR U22858 ( .A(n22462), .B(n22461), .Z(n22463) );
  XNOR U22859 ( .A(n22464), .B(n22463), .Z(n24944) );
  XNOR U22860 ( .A(n22466), .B(n22465), .Z(n24943) );
  NAND U22861 ( .A(n24944), .B(n24943), .Z(n22467) );
  AND U22862 ( .A(n22468), .B(n22467), .Z(n24946) );
  NAND U22863 ( .A(a[60]), .B(b[0]), .Z(n24945) );
  XNOR U22864 ( .A(n22470), .B(n22469), .Z(n22471) );
  XNOR U22865 ( .A(n22472), .B(n22471), .Z(n24948) );
  NAND U22866 ( .A(a[61]), .B(b[0]), .Z(n22473) );
  NANDN U22867 ( .A(n22474), .B(n22473), .Z(n22480) );
  XNOR U22868 ( .A(n22474), .B(n22473), .Z(n24950) );
  XOR U22869 ( .A(n22476), .B(n22475), .Z(n22477) );
  XNOR U22870 ( .A(n22478), .B(n22477), .Z(n24949) );
  NAND U22871 ( .A(n24950), .B(n24949), .Z(n22479) );
  NAND U22872 ( .A(n22480), .B(n22479), .Z(n24954) );
  AND U22873 ( .A(a[62]), .B(b[0]), .Z(n24953) );
  NAND U22874 ( .A(a[63]), .B(b[0]), .Z(n22481) );
  NANDN U22875 ( .A(n22482), .B(n22481), .Z(n22488) );
  XNOR U22876 ( .A(n22482), .B(n22481), .Z(n24958) );
  XOR U22877 ( .A(n22484), .B(n22483), .Z(n22485) );
  XNOR U22878 ( .A(n22486), .B(n22485), .Z(n24957) );
  NAND U22879 ( .A(n24958), .B(n24957), .Z(n22487) );
  AND U22880 ( .A(n22488), .B(n22487), .Z(n24959) );
  AND U22881 ( .A(n24960), .B(n24959), .Z(n24660) );
  XNOR U22882 ( .A(n22490), .B(n22489), .Z(n24659) );
  NAND U22883 ( .A(n24660), .B(n24659), .Z(n22491) );
  NAND U22884 ( .A(n22492), .B(n22491), .Z(n24661) );
  AND U22885 ( .A(n24662), .B(n24661), .Z(n24666) );
  ANDN U22886 ( .B(n22494), .A(n22493), .Z(n24668) );
  XOR U22887 ( .A(n22496), .B(n22495), .Z(n24667) );
  ANDN U22888 ( .B(n24668), .A(n24667), .Z(n24672) );
  NANDN U22889 ( .A(n24688), .B(n24686), .Z(n22497) );
  NAND U22890 ( .A(n22498), .B(n22497), .Z(n22499) );
  NANDN U22891 ( .A(n22500), .B(n22499), .Z(n22502) );
  NANDN U22892 ( .A(n24693), .B(n24694), .Z(n22501) );
  AND U22893 ( .A(n22502), .B(n22501), .Z(n24700) );
  NANDN U22894 ( .A(n24697), .B(n24698), .Z(n22503) );
  NAND U22895 ( .A(n24700), .B(n22503), .Z(n24704) );
  NAND U22896 ( .A(n24720), .B(n24719), .Z(n22504) );
  NAND U22897 ( .A(n22505), .B(n22504), .Z(n24721) );
  XNOR U22898 ( .A(n22507), .B(n22506), .Z(n24724) );
  XOR U22899 ( .A(n22509), .B(n22508), .Z(n24725) );
  XNOR U22900 ( .A(n22511), .B(n22510), .Z(n24729) );
  NAND U22901 ( .A(n24730), .B(n24729), .Z(n22512) );
  NAND U22902 ( .A(n22513), .B(n22512), .Z(n24731) );
  NAND U22903 ( .A(n24732), .B(n24731), .Z(n22514) );
  NAND U22904 ( .A(n22515), .B(n22514), .Z(n24733) );
  NAND U22905 ( .A(n24734), .B(n24733), .Z(n22516) );
  NAND U22906 ( .A(n22517), .B(n22516), .Z(n24735) );
  NAND U22907 ( .A(n24736), .B(n24735), .Z(n22518) );
  NAND U22908 ( .A(n22519), .B(n22518), .Z(n24741) );
  NAND U22909 ( .A(n22521), .B(n22520), .Z(n24768) );
  XOR U22910 ( .A(n22523), .B(n22522), .Z(n22531) );
  NAND U22911 ( .A(n22525), .B(n22524), .Z(n22529) );
  NAND U22912 ( .A(n22527), .B(n22526), .Z(n22528) );
  NAND U22913 ( .A(n22529), .B(n22528), .Z(n22530) );
  XNOR U22914 ( .A(n22531), .B(n22530), .Z(n24767) );
  NAND U22915 ( .A(n24770), .B(n24772), .Z(n22533) );
  NAND U22916 ( .A(n22531), .B(n22530), .Z(n24773) );
  OR U22917 ( .A(n22533), .B(n24773), .Z(n22532) );
  NAND U22918 ( .A(n24776), .B(n22532), .Z(n22537) );
  AND U22919 ( .A(n22533), .B(n24773), .Z(n22535) );
  OR U22920 ( .A(n24767), .B(n24768), .Z(n22534) );
  NAND U22921 ( .A(n22535), .B(n22534), .Z(n22536) );
  NAND U22922 ( .A(n22537), .B(n22536), .Z(n24778) );
  XNOR U22923 ( .A(n22539), .B(n22538), .Z(n24777) );
  NAND U22924 ( .A(n24778), .B(n24777), .Z(n22540) );
  NAND U22925 ( .A(n22541), .B(n22540), .Z(n24779) );
  NAND U22926 ( .A(n24780), .B(n24779), .Z(n22542) );
  NAND U22927 ( .A(n22543), .B(n22542), .Z(n24781) );
  NAND U22928 ( .A(n24782), .B(n24781), .Z(n22544) );
  NAND U22929 ( .A(n22545), .B(n22544), .Z(n24783) );
  XNOR U22930 ( .A(n22547), .B(n22546), .Z(n24786) );
  XOR U22931 ( .A(n22549), .B(n22548), .Z(n24787) );
  XNOR U22932 ( .A(n22551), .B(n22550), .Z(n24791) );
  NAND U22933 ( .A(n24792), .B(n24791), .Z(n22552) );
  AND U22934 ( .A(n22553), .B(n22552), .Z(n24796) );
  NAND U22935 ( .A(n22555), .B(n22554), .Z(n22846) );
  NANDN U22936 ( .A(n22557), .B(n22556), .Z(n22561) );
  NAND U22937 ( .A(n22559), .B(n22558), .Z(n22560) );
  AND U22938 ( .A(n22561), .B(n22560), .Z(n22710) );
  AND U22939 ( .A(a[63]), .B(b[39]), .Z(n22709) );
  XNOR U22940 ( .A(n22710), .B(n22709), .Z(n22711) );
  NANDN U22941 ( .A(n22563), .B(n22562), .Z(n22567) );
  NAND U22942 ( .A(n22565), .B(n22564), .Z(n22566) );
  AND U22943 ( .A(n22567), .B(n22566), .Z(n22718) );
  NANDN U22944 ( .A(n22569), .B(n22568), .Z(n22573) );
  NAND U22945 ( .A(n22571), .B(n22570), .Z(n22572) );
  NAND U22946 ( .A(n22573), .B(n22572), .Z(n22841) );
  AND U22947 ( .A(a[61]), .B(b[41]), .Z(n22842) );
  XOR U22948 ( .A(n22841), .B(n22842), .Z(n22843) );
  NAND U22949 ( .A(n22575), .B(n22574), .Z(n22579) );
  NANDN U22950 ( .A(n22577), .B(n22576), .Z(n22578) );
  NAND U22951 ( .A(n22579), .B(n22578), .Z(n22724) );
  NAND U22952 ( .A(n22581), .B(n22580), .Z(n22585) );
  NANDN U22953 ( .A(n22583), .B(n22582), .Z(n22584) );
  AND U22954 ( .A(n22585), .B(n22584), .Z(n22838) );
  AND U22955 ( .A(a[59]), .B(b[43]), .Z(n22837) );
  XOR U22956 ( .A(n22838), .B(n22837), .Z(n22839) );
  NAND U22957 ( .A(n22587), .B(n22586), .Z(n22591) );
  NAND U22958 ( .A(n22589), .B(n22588), .Z(n22590) );
  NAND U22959 ( .A(n22591), .B(n22590), .Z(n22728) );
  NANDN U22960 ( .A(n22593), .B(n22592), .Z(n22597) );
  NAND U22961 ( .A(n22595), .B(n22594), .Z(n22596) );
  AND U22962 ( .A(n22597), .B(n22596), .Z(n22832) );
  AND U22963 ( .A(a[57]), .B(b[45]), .Z(n22831) );
  XNOR U22964 ( .A(n22832), .B(n22831), .Z(n22833) );
  NANDN U22965 ( .A(n22599), .B(n22598), .Z(n22603) );
  NAND U22966 ( .A(n22601), .B(n22600), .Z(n22602) );
  AND U22967 ( .A(n22603), .B(n22602), .Z(n22732) );
  NANDN U22968 ( .A(n22605), .B(n22604), .Z(n22609) );
  NAND U22969 ( .A(n22607), .B(n22606), .Z(n22608) );
  AND U22970 ( .A(n22609), .B(n22608), .Z(n22826) );
  AND U22971 ( .A(a[55]), .B(b[47]), .Z(n22825) );
  XNOR U22972 ( .A(n22826), .B(n22825), .Z(n22827) );
  NANDN U22973 ( .A(n22611), .B(n22610), .Z(n22615) );
  NAND U22974 ( .A(n22613), .B(n22612), .Z(n22614) );
  AND U22975 ( .A(n22615), .B(n22614), .Z(n22738) );
  NANDN U22976 ( .A(n22617), .B(n22616), .Z(n22621) );
  NAND U22977 ( .A(n22619), .B(n22618), .Z(n22620) );
  AND U22978 ( .A(n22621), .B(n22620), .Z(n22820) );
  AND U22979 ( .A(a[53]), .B(b[49]), .Z(n22819) );
  XNOR U22980 ( .A(n22820), .B(n22819), .Z(n22821) );
  NANDN U22981 ( .A(n22623), .B(n22622), .Z(n22627) );
  NAND U22982 ( .A(n22625), .B(n22624), .Z(n22626) );
  AND U22983 ( .A(n22627), .B(n22626), .Z(n22744) );
  NANDN U22984 ( .A(n22629), .B(n22628), .Z(n22633) );
  NAND U22985 ( .A(n22631), .B(n22630), .Z(n22632) );
  AND U22986 ( .A(n22633), .B(n22632), .Z(n22814) );
  AND U22987 ( .A(a[51]), .B(b[51]), .Z(n22813) );
  XNOR U22988 ( .A(n22814), .B(n22813), .Z(n22815) );
  NANDN U22989 ( .A(n22635), .B(n22634), .Z(n22639) );
  NAND U22990 ( .A(n22637), .B(n22636), .Z(n22638) );
  AND U22991 ( .A(n22639), .B(n22638), .Z(n22750) );
  NANDN U22992 ( .A(n22641), .B(n22640), .Z(n22645) );
  NAND U22993 ( .A(n22643), .B(n22642), .Z(n22644) );
  AND U22994 ( .A(n22645), .B(n22644), .Z(n22755) );
  NANDN U22995 ( .A(n22647), .B(n22646), .Z(n22651) );
  NAND U22996 ( .A(n22649), .B(n22648), .Z(n22650) );
  AND U22997 ( .A(n22651), .B(n22650), .Z(n22802) );
  AND U22998 ( .A(a[47]), .B(b[55]), .Z(n22801) );
  XNOR U22999 ( .A(n22802), .B(n22801), .Z(n22803) );
  NANDN U23000 ( .A(n22653), .B(n22652), .Z(n22657) );
  NAND U23001 ( .A(n22655), .B(n22654), .Z(n22656) );
  AND U23002 ( .A(n22657), .B(n22656), .Z(n22762) );
  NANDN U23003 ( .A(n22659), .B(n22658), .Z(n22663) );
  NAND U23004 ( .A(n22661), .B(n22660), .Z(n22662) );
  AND U23005 ( .A(n22663), .B(n22662), .Z(n22796) );
  AND U23006 ( .A(a[45]), .B(b[57]), .Z(n22795) );
  XNOR U23007 ( .A(n22796), .B(n22795), .Z(n22797) );
  NANDN U23008 ( .A(n22665), .B(n22664), .Z(n22669) );
  NANDN U23009 ( .A(n22667), .B(n22666), .Z(n22668) );
  AND U23010 ( .A(n22669), .B(n22668), .Z(n22768) );
  NANDN U23011 ( .A(n22671), .B(n22670), .Z(n22675) );
  NAND U23012 ( .A(n22673), .B(n22672), .Z(n22674) );
  AND U23013 ( .A(n22675), .B(n22674), .Z(n22771) );
  NAND U23014 ( .A(a[43]), .B(b[59]), .Z(n22772) );
  XNOR U23015 ( .A(n22771), .B(n22772), .Z(n22773) );
  NANDN U23016 ( .A(n22677), .B(n22676), .Z(n22681) );
  NANDN U23017 ( .A(n22679), .B(n22678), .Z(n22680) );
  AND U23018 ( .A(n22681), .B(n22680), .Z(n22777) );
  NAND U23019 ( .A(a[42]), .B(b[60]), .Z(n22778) );
  XNOR U23020 ( .A(n22777), .B(n22778), .Z(n22779) );
  NANDN U23021 ( .A(n22683), .B(n22682), .Z(n22687) );
  NAND U23022 ( .A(n22685), .B(n22684), .Z(n22686) );
  AND U23023 ( .A(n22687), .B(n22686), .Z(n22790) );
  NANDN U23024 ( .A(n22689), .B(n22688), .Z(n22693) );
  NAND U23025 ( .A(n22691), .B(n22690), .Z(n22692) );
  AND U23026 ( .A(n22693), .B(n22692), .Z(n22786) );
  AND U23027 ( .A(b[63]), .B(a[39]), .Z(n22783) );
  NAND U23028 ( .A(b[62]), .B(a[40]), .Z(n22784) );
  XNOR U23029 ( .A(n22783), .B(n22784), .Z(n22785) );
  XNOR U23030 ( .A(n22786), .B(n22785), .Z(n22789) );
  XNOR U23031 ( .A(n22790), .B(n22789), .Z(n22791) );
  NAND U23032 ( .A(a[41]), .B(b[61]), .Z(n22792) );
  XOR U23033 ( .A(n22791), .B(n22792), .Z(n22780) );
  XOR U23034 ( .A(n22779), .B(n22780), .Z(n22774) );
  XNOR U23035 ( .A(n22773), .B(n22774), .Z(n22765) );
  NAND U23036 ( .A(a[44]), .B(b[58]), .Z(n22766) );
  XNOR U23037 ( .A(n22765), .B(n22766), .Z(n22767) );
  XOR U23038 ( .A(n22768), .B(n22767), .Z(n22798) );
  XNOR U23039 ( .A(n22797), .B(n22798), .Z(n22759) );
  NAND U23040 ( .A(a[46]), .B(b[56]), .Z(n22760) );
  XNOR U23041 ( .A(n22759), .B(n22760), .Z(n22761) );
  XOR U23042 ( .A(n22762), .B(n22761), .Z(n22804) );
  XNOR U23043 ( .A(n22803), .B(n22804), .Z(n22753) );
  NAND U23044 ( .A(a[48]), .B(b[54]), .Z(n22754) );
  XOR U23045 ( .A(n22753), .B(n22754), .Z(n22756) );
  XOR U23046 ( .A(n22755), .B(n22756), .Z(n22809) );
  AND U23047 ( .A(a[49]), .B(b[53]), .Z(n22808) );
  NANDN U23048 ( .A(n22695), .B(n22694), .Z(n22699) );
  NAND U23049 ( .A(n22697), .B(n22696), .Z(n22698) );
  AND U23050 ( .A(n22699), .B(n22698), .Z(n22807) );
  XOR U23051 ( .A(n22808), .B(n22807), .Z(n22810) );
  XOR U23052 ( .A(n22809), .B(n22810), .Z(n22748) );
  AND U23053 ( .A(a[50]), .B(b[52]), .Z(n22747) );
  XNOR U23054 ( .A(n22748), .B(n22747), .Z(n22749) );
  XOR U23055 ( .A(n22750), .B(n22749), .Z(n22816) );
  XNOR U23056 ( .A(n22815), .B(n22816), .Z(n22741) );
  NAND U23057 ( .A(a[52]), .B(b[50]), .Z(n22742) );
  XNOR U23058 ( .A(n22741), .B(n22742), .Z(n22743) );
  XOR U23059 ( .A(n22744), .B(n22743), .Z(n22822) );
  XNOR U23060 ( .A(n22821), .B(n22822), .Z(n22735) );
  NAND U23061 ( .A(a[54]), .B(b[48]), .Z(n22736) );
  XNOR U23062 ( .A(n22735), .B(n22736), .Z(n22737) );
  XOR U23063 ( .A(n22738), .B(n22737), .Z(n22828) );
  XNOR U23064 ( .A(n22827), .B(n22828), .Z(n22729) );
  NAND U23065 ( .A(a[56]), .B(b[46]), .Z(n22730) );
  XNOR U23066 ( .A(n22729), .B(n22730), .Z(n22731) );
  XOR U23067 ( .A(n22732), .B(n22731), .Z(n22834) );
  XNOR U23068 ( .A(n22833), .B(n22834), .Z(n22726) );
  AND U23069 ( .A(a[58]), .B(b[44]), .Z(n22725) );
  XOR U23070 ( .A(n22726), .B(n22725), .Z(n22727) );
  XNOR U23071 ( .A(n22728), .B(n22727), .Z(n22840) );
  XNOR U23072 ( .A(n22839), .B(n22840), .Z(n22722) );
  AND U23073 ( .A(a[60]), .B(b[42]), .Z(n22721) );
  XOR U23074 ( .A(n22722), .B(n22721), .Z(n22723) );
  XNOR U23075 ( .A(n22724), .B(n22723), .Z(n22844) );
  XNOR U23076 ( .A(n22843), .B(n22844), .Z(n22715) );
  NAND U23077 ( .A(a[62]), .B(b[40]), .Z(n22716) );
  XNOR U23078 ( .A(n22715), .B(n22716), .Z(n22717) );
  XOR U23079 ( .A(n22718), .B(n22717), .Z(n22712) );
  XNOR U23080 ( .A(n22711), .B(n22712), .Z(n22708) );
  NAND U23081 ( .A(n22701), .B(n22700), .Z(n22705) );
  NANDN U23082 ( .A(n22703), .B(n22702), .Z(n22704) );
  AND U23083 ( .A(n22705), .B(n22704), .Z(n22707) );
  XOR U23084 ( .A(n22708), .B(n22707), .Z(n22845) );
  XOR U23085 ( .A(n22846), .B(n22845), .Z(n22706) );
  XNOR U23086 ( .A(n22847), .B(n22706), .Z(c[102]) );
  NAND U23087 ( .A(n22708), .B(n22707), .Z(n22851) );
  NANDN U23088 ( .A(n22710), .B(n22709), .Z(n22714) );
  NANDN U23089 ( .A(n22712), .B(n22711), .Z(n22713) );
  AND U23090 ( .A(n22714), .B(n22713), .Z(n22983) );
  NANDN U23091 ( .A(n22716), .B(n22715), .Z(n22720) );
  NANDN U23092 ( .A(n22718), .B(n22717), .Z(n22719) );
  AND U23093 ( .A(n22720), .B(n22719), .Z(n22853) );
  AND U23094 ( .A(a[63]), .B(b[40]), .Z(n22852) );
  XNOR U23095 ( .A(n22853), .B(n22852), .Z(n22854) );
  AND U23096 ( .A(a[61]), .B(b[42]), .Z(n22863) );
  XOR U23097 ( .A(n22862), .B(n22863), .Z(n22865) );
  AND U23098 ( .A(a[59]), .B(b[44]), .Z(n22871) );
  XOR U23099 ( .A(n22870), .B(n22871), .Z(n22873) );
  NANDN U23100 ( .A(n22730), .B(n22729), .Z(n22734) );
  NANDN U23101 ( .A(n22732), .B(n22731), .Z(n22733) );
  AND U23102 ( .A(n22734), .B(n22733), .Z(n22881) );
  AND U23103 ( .A(a[57]), .B(b[46]), .Z(n22880) );
  XNOR U23104 ( .A(n22881), .B(n22880), .Z(n22882) );
  NANDN U23105 ( .A(n22736), .B(n22735), .Z(n22740) );
  NANDN U23106 ( .A(n22738), .B(n22737), .Z(n22739) );
  AND U23107 ( .A(n22740), .B(n22739), .Z(n22893) );
  AND U23108 ( .A(a[55]), .B(b[48]), .Z(n22892) );
  XNOR U23109 ( .A(n22893), .B(n22892), .Z(n22894) );
  NANDN U23110 ( .A(n22742), .B(n22741), .Z(n22746) );
  NANDN U23111 ( .A(n22744), .B(n22743), .Z(n22745) );
  AND U23112 ( .A(n22746), .B(n22745), .Z(n22905) );
  AND U23113 ( .A(a[53]), .B(b[50]), .Z(n22904) );
  XNOR U23114 ( .A(n22905), .B(n22904), .Z(n22906) );
  NANDN U23115 ( .A(n22748), .B(n22747), .Z(n22752) );
  NANDN U23116 ( .A(n22750), .B(n22749), .Z(n22751) );
  AND U23117 ( .A(n22752), .B(n22751), .Z(n22917) );
  AND U23118 ( .A(a[51]), .B(b[52]), .Z(n22916) );
  XNOR U23119 ( .A(n22917), .B(n22916), .Z(n22918) );
  NANDN U23120 ( .A(n22754), .B(n22753), .Z(n22758) );
  OR U23121 ( .A(n22756), .B(n22755), .Z(n22757) );
  AND U23122 ( .A(n22758), .B(n22757), .Z(n22929) );
  AND U23123 ( .A(a[49]), .B(b[54]), .Z(n22928) );
  XNOR U23124 ( .A(n22929), .B(n22928), .Z(n22930) );
  AND U23125 ( .A(a[47]), .B(b[56]), .Z(n22941) );
  NANDN U23126 ( .A(n22760), .B(n22759), .Z(n22764) );
  NANDN U23127 ( .A(n22762), .B(n22761), .Z(n22763) );
  AND U23128 ( .A(n22764), .B(n22763), .Z(n22940) );
  XNOR U23129 ( .A(n22941), .B(n22940), .Z(n22943) );
  AND U23130 ( .A(a[46]), .B(b[57]), .Z(n22949) );
  NANDN U23131 ( .A(n22766), .B(n22765), .Z(n22770) );
  NANDN U23132 ( .A(n22768), .B(n22767), .Z(n22769) );
  AND U23133 ( .A(n22770), .B(n22769), .Z(n22954) );
  NANDN U23134 ( .A(n22772), .B(n22771), .Z(n22776) );
  NANDN U23135 ( .A(n22774), .B(n22773), .Z(n22775) );
  AND U23136 ( .A(n22776), .B(n22775), .Z(n22977) );
  AND U23137 ( .A(a[44]), .B(b[59]), .Z(n22976) );
  XNOR U23138 ( .A(n22977), .B(n22976), .Z(n22978) );
  NANDN U23139 ( .A(n22778), .B(n22777), .Z(n22782) );
  NANDN U23140 ( .A(n22780), .B(n22779), .Z(n22781) );
  AND U23141 ( .A(n22782), .B(n22781), .Z(n22961) );
  NANDN U23142 ( .A(n22784), .B(n22783), .Z(n22788) );
  NANDN U23143 ( .A(n22786), .B(n22785), .Z(n22787) );
  AND U23144 ( .A(n22788), .B(n22787), .Z(n22966) );
  AND U23145 ( .A(b[62]), .B(a[41]), .Z(n22964) );
  NAND U23146 ( .A(b[63]), .B(a[40]), .Z(n22965) );
  XOR U23147 ( .A(n22964), .B(n22965), .Z(n22967) );
  XOR U23148 ( .A(n22966), .B(n22967), .Z(n22972) );
  AND U23149 ( .A(a[42]), .B(b[61]), .Z(n22971) );
  NANDN U23150 ( .A(n22790), .B(n22789), .Z(n22794) );
  NANDN U23151 ( .A(n22792), .B(n22791), .Z(n22793) );
  AND U23152 ( .A(n22794), .B(n22793), .Z(n22970) );
  XOR U23153 ( .A(n22971), .B(n22970), .Z(n22973) );
  XOR U23154 ( .A(n22972), .B(n22973), .Z(n22959) );
  AND U23155 ( .A(a[43]), .B(b[60]), .Z(n22958) );
  XNOR U23156 ( .A(n22959), .B(n22958), .Z(n22960) );
  XOR U23157 ( .A(n22961), .B(n22960), .Z(n22979) );
  XNOR U23158 ( .A(n22978), .B(n22979), .Z(n22952) );
  NAND U23159 ( .A(a[45]), .B(b[58]), .Z(n22953) );
  XOR U23160 ( .A(n22952), .B(n22953), .Z(n22955) );
  XOR U23161 ( .A(n22954), .B(n22955), .Z(n22947) );
  NANDN U23162 ( .A(n22796), .B(n22795), .Z(n22800) );
  NANDN U23163 ( .A(n22798), .B(n22797), .Z(n22799) );
  AND U23164 ( .A(n22800), .B(n22799), .Z(n22946) );
  XNOR U23165 ( .A(n22947), .B(n22946), .Z(n22948) );
  XNOR U23166 ( .A(n22949), .B(n22948), .Z(n22942) );
  XOR U23167 ( .A(n22943), .B(n22942), .Z(n22937) );
  NANDN U23168 ( .A(n22802), .B(n22801), .Z(n22806) );
  NANDN U23169 ( .A(n22804), .B(n22803), .Z(n22805) );
  AND U23170 ( .A(n22806), .B(n22805), .Z(n22935) );
  AND U23171 ( .A(a[48]), .B(b[55]), .Z(n22934) );
  XNOR U23172 ( .A(n22935), .B(n22934), .Z(n22936) );
  XOR U23173 ( .A(n22937), .B(n22936), .Z(n22931) );
  XNOR U23174 ( .A(n22930), .B(n22931), .Z(n22924) );
  NANDN U23175 ( .A(n22808), .B(n22807), .Z(n22812) );
  OR U23176 ( .A(n22810), .B(n22809), .Z(n22811) );
  AND U23177 ( .A(n22812), .B(n22811), .Z(n22922) );
  NAND U23178 ( .A(a[50]), .B(b[53]), .Z(n22923) );
  XOR U23179 ( .A(n22922), .B(n22923), .Z(n22925) );
  XOR U23180 ( .A(n22924), .B(n22925), .Z(n22919) );
  XNOR U23181 ( .A(n22918), .B(n22919), .Z(n22912) );
  NANDN U23182 ( .A(n22814), .B(n22813), .Z(n22818) );
  NANDN U23183 ( .A(n22816), .B(n22815), .Z(n22817) );
  AND U23184 ( .A(n22818), .B(n22817), .Z(n22911) );
  AND U23185 ( .A(a[52]), .B(b[51]), .Z(n22910) );
  XOR U23186 ( .A(n22911), .B(n22910), .Z(n22913) );
  XOR U23187 ( .A(n22912), .B(n22913), .Z(n22907) );
  XNOR U23188 ( .A(n22906), .B(n22907), .Z(n22900) );
  NANDN U23189 ( .A(n22820), .B(n22819), .Z(n22824) );
  NANDN U23190 ( .A(n22822), .B(n22821), .Z(n22823) );
  AND U23191 ( .A(n22824), .B(n22823), .Z(n22899) );
  AND U23192 ( .A(a[54]), .B(b[49]), .Z(n22898) );
  XOR U23193 ( .A(n22899), .B(n22898), .Z(n22901) );
  XOR U23194 ( .A(n22900), .B(n22901), .Z(n22895) );
  XNOR U23195 ( .A(n22894), .B(n22895), .Z(n22888) );
  NANDN U23196 ( .A(n22826), .B(n22825), .Z(n22830) );
  NANDN U23197 ( .A(n22828), .B(n22827), .Z(n22829) );
  AND U23198 ( .A(n22830), .B(n22829), .Z(n22887) );
  AND U23199 ( .A(a[56]), .B(b[47]), .Z(n22886) );
  XOR U23200 ( .A(n22887), .B(n22886), .Z(n22889) );
  XOR U23201 ( .A(n22888), .B(n22889), .Z(n22883) );
  XNOR U23202 ( .A(n22882), .B(n22883), .Z(n22877) );
  NANDN U23203 ( .A(n22832), .B(n22831), .Z(n22836) );
  NANDN U23204 ( .A(n22834), .B(n22833), .Z(n22835) );
  AND U23205 ( .A(n22836), .B(n22835), .Z(n22875) );
  AND U23206 ( .A(a[58]), .B(b[45]), .Z(n22874) );
  XNOR U23207 ( .A(n22875), .B(n22874), .Z(n22876) );
  XOR U23208 ( .A(n22877), .B(n22876), .Z(n22872) );
  XOR U23209 ( .A(n22873), .B(n22872), .Z(n22869) );
  AND U23210 ( .A(a[60]), .B(b[43]), .Z(n22867) );
  XOR U23211 ( .A(n22866), .B(n22867), .Z(n22868) );
  XOR U23212 ( .A(n22869), .B(n22868), .Z(n22864) );
  XOR U23213 ( .A(n22865), .B(n22864), .Z(n22860) );
  AND U23214 ( .A(a[62]), .B(b[41]), .Z(n22858) );
  XNOR U23215 ( .A(n22859), .B(n22858), .Z(n22861) );
  XOR U23216 ( .A(n22860), .B(n22861), .Z(n22855) );
  XNOR U23217 ( .A(n22854), .B(n22855), .Z(n22982) );
  XOR U23218 ( .A(n22983), .B(n22982), .Z(n22849) );
  XOR U23219 ( .A(n22849), .B(n22850), .Z(n22848) );
  XNOR U23220 ( .A(n22851), .B(n22848), .Z(c[103]) );
  NANDN U23221 ( .A(n22853), .B(n22852), .Z(n22857) );
  NANDN U23222 ( .A(n22855), .B(n22854), .Z(n22856) );
  NAND U23223 ( .A(n22857), .B(n22856), .Z(n22990) );
  AND U23224 ( .A(a[63]), .B(b[41]), .Z(n22993) );
  XOR U23225 ( .A(n22992), .B(n22993), .Z(n22994) );
  AND U23226 ( .A(a[61]), .B(b[43]), .Z(n23109) );
  XOR U23227 ( .A(n23108), .B(n23109), .Z(n23110) );
  NANDN U23228 ( .A(n22875), .B(n22874), .Z(n22879) );
  NAND U23229 ( .A(n22877), .B(n22876), .Z(n22878) );
  AND U23230 ( .A(n22879), .B(n22878), .Z(n23103) );
  AND U23231 ( .A(a[59]), .B(b[45]), .Z(n23102) );
  XNOR U23232 ( .A(n23103), .B(n23102), .Z(n23104) );
  NANDN U23233 ( .A(n22881), .B(n22880), .Z(n22885) );
  NANDN U23234 ( .A(n22883), .B(n22882), .Z(n22884) );
  AND U23235 ( .A(n22885), .B(n22884), .Z(n23003) );
  NANDN U23236 ( .A(n22887), .B(n22886), .Z(n22891) );
  NANDN U23237 ( .A(n22889), .B(n22888), .Z(n22890) );
  AND U23238 ( .A(n22891), .B(n22890), .Z(n23097) );
  AND U23239 ( .A(a[57]), .B(b[47]), .Z(n23096) );
  XNOR U23240 ( .A(n23097), .B(n23096), .Z(n23098) );
  NANDN U23241 ( .A(n22893), .B(n22892), .Z(n22897) );
  NANDN U23242 ( .A(n22895), .B(n22894), .Z(n22896) );
  AND U23243 ( .A(n22897), .B(n22896), .Z(n23009) );
  NANDN U23244 ( .A(n22899), .B(n22898), .Z(n22903) );
  NANDN U23245 ( .A(n22901), .B(n22900), .Z(n22902) );
  AND U23246 ( .A(n22903), .B(n22902), .Z(n23091) );
  AND U23247 ( .A(a[55]), .B(b[49]), .Z(n23090) );
  XNOR U23248 ( .A(n23091), .B(n23090), .Z(n23092) );
  NANDN U23249 ( .A(n22905), .B(n22904), .Z(n22909) );
  NANDN U23250 ( .A(n22907), .B(n22906), .Z(n22908) );
  AND U23251 ( .A(n22909), .B(n22908), .Z(n23015) );
  NANDN U23252 ( .A(n22911), .B(n22910), .Z(n22915) );
  NANDN U23253 ( .A(n22913), .B(n22912), .Z(n22914) );
  AND U23254 ( .A(n22915), .B(n22914), .Z(n23085) );
  AND U23255 ( .A(a[53]), .B(b[51]), .Z(n23084) );
  XNOR U23256 ( .A(n23085), .B(n23084), .Z(n23086) );
  NANDN U23257 ( .A(n22917), .B(n22916), .Z(n22921) );
  NANDN U23258 ( .A(n22919), .B(n22918), .Z(n22920) );
  AND U23259 ( .A(n22921), .B(n22920), .Z(n23021) );
  NANDN U23260 ( .A(n22923), .B(n22922), .Z(n22927) );
  NANDN U23261 ( .A(n22925), .B(n22924), .Z(n22926) );
  AND U23262 ( .A(n22927), .B(n22926), .Z(n23079) );
  AND U23263 ( .A(a[51]), .B(b[53]), .Z(n23078) );
  XNOR U23264 ( .A(n23079), .B(n23078), .Z(n23080) );
  NANDN U23265 ( .A(n22929), .B(n22928), .Z(n22933) );
  NANDN U23266 ( .A(n22931), .B(n22930), .Z(n22932) );
  AND U23267 ( .A(n22933), .B(n22932), .Z(n23027) );
  NANDN U23268 ( .A(n22935), .B(n22934), .Z(n22939) );
  NANDN U23269 ( .A(n22937), .B(n22936), .Z(n22938) );
  AND U23270 ( .A(n22939), .B(n22938), .Z(n23073) );
  AND U23271 ( .A(a[49]), .B(b[55]), .Z(n23072) );
  XNOR U23272 ( .A(n23073), .B(n23072), .Z(n23074) );
  NANDN U23273 ( .A(n22941), .B(n22940), .Z(n22945) );
  NAND U23274 ( .A(n22943), .B(n22942), .Z(n22944) );
  AND U23275 ( .A(n22945), .B(n22944), .Z(n23032) );
  AND U23276 ( .A(a[47]), .B(b[57]), .Z(n23068) );
  NANDN U23277 ( .A(n22947), .B(n22946), .Z(n22951) );
  NANDN U23278 ( .A(n22949), .B(n22948), .Z(n22950) );
  AND U23279 ( .A(n22951), .B(n22950), .Z(n23067) );
  NANDN U23280 ( .A(n22953), .B(n22952), .Z(n22957) );
  OR U23281 ( .A(n22955), .B(n22954), .Z(n22956) );
  AND U23282 ( .A(n22957), .B(n22956), .Z(n23037) );
  AND U23283 ( .A(a[46]), .B(b[58]), .Z(n23036) );
  XNOR U23284 ( .A(n23037), .B(n23036), .Z(n23039) );
  NANDN U23285 ( .A(n22959), .B(n22958), .Z(n22963) );
  NANDN U23286 ( .A(n22961), .B(n22960), .Z(n22962) );
  AND U23287 ( .A(n22963), .B(n22962), .Z(n23049) );
  AND U23288 ( .A(a[44]), .B(b[60]), .Z(n23048) );
  XNOR U23289 ( .A(n23049), .B(n23048), .Z(n23050) );
  NANDN U23290 ( .A(n22965), .B(n22964), .Z(n22969) );
  OR U23291 ( .A(n22967), .B(n22966), .Z(n22968) );
  AND U23292 ( .A(n22969), .B(n22968), .Z(n23061) );
  AND U23293 ( .A(b[62]), .B(a[42]), .Z(n23060) );
  XNOR U23294 ( .A(n23061), .B(n23060), .Z(n23062) );
  NAND U23295 ( .A(b[63]), .B(a[41]), .Z(n23063) );
  XNOR U23296 ( .A(n23062), .B(n23063), .Z(n23056) );
  NANDN U23297 ( .A(n22971), .B(n22970), .Z(n22975) );
  OR U23298 ( .A(n22973), .B(n22972), .Z(n22974) );
  AND U23299 ( .A(n22975), .B(n22974), .Z(n23054) );
  NAND U23300 ( .A(a[43]), .B(b[61]), .Z(n23055) );
  XOR U23301 ( .A(n23054), .B(n23055), .Z(n23057) );
  XOR U23302 ( .A(n23056), .B(n23057), .Z(n23051) );
  XNOR U23303 ( .A(n23050), .B(n23051), .Z(n23044) );
  NANDN U23304 ( .A(n22977), .B(n22976), .Z(n22981) );
  NANDN U23305 ( .A(n22979), .B(n22978), .Z(n22980) );
  AND U23306 ( .A(n22981), .B(n22980), .Z(n23043) );
  AND U23307 ( .A(a[45]), .B(b[59]), .Z(n23042) );
  XOR U23308 ( .A(n23043), .B(n23042), .Z(n23045) );
  XNOR U23309 ( .A(n23044), .B(n23045), .Z(n23038) );
  XNOR U23310 ( .A(n23039), .B(n23038), .Z(n23066) );
  XOR U23311 ( .A(n23067), .B(n23066), .Z(n23069) );
  XOR U23312 ( .A(n23068), .B(n23069), .Z(n23031) );
  AND U23313 ( .A(a[48]), .B(b[56]), .Z(n23030) );
  XOR U23314 ( .A(n23031), .B(n23030), .Z(n23033) );
  XOR U23315 ( .A(n23032), .B(n23033), .Z(n23075) );
  XNOR U23316 ( .A(n23074), .B(n23075), .Z(n23024) );
  NAND U23317 ( .A(a[50]), .B(b[54]), .Z(n23025) );
  XNOR U23318 ( .A(n23024), .B(n23025), .Z(n23026) );
  XOR U23319 ( .A(n23027), .B(n23026), .Z(n23081) );
  XNOR U23320 ( .A(n23080), .B(n23081), .Z(n23018) );
  NAND U23321 ( .A(a[52]), .B(b[52]), .Z(n23019) );
  XNOR U23322 ( .A(n23018), .B(n23019), .Z(n23020) );
  XOR U23323 ( .A(n23021), .B(n23020), .Z(n23087) );
  XNOR U23324 ( .A(n23086), .B(n23087), .Z(n23012) );
  NAND U23325 ( .A(a[54]), .B(b[50]), .Z(n23013) );
  XNOR U23326 ( .A(n23012), .B(n23013), .Z(n23014) );
  XOR U23327 ( .A(n23015), .B(n23014), .Z(n23093) );
  XNOR U23328 ( .A(n23092), .B(n23093), .Z(n23006) );
  NAND U23329 ( .A(a[56]), .B(b[48]), .Z(n23007) );
  XNOR U23330 ( .A(n23006), .B(n23007), .Z(n23008) );
  XOR U23331 ( .A(n23009), .B(n23008), .Z(n23099) );
  XNOR U23332 ( .A(n23098), .B(n23099), .Z(n23000) );
  NAND U23333 ( .A(a[58]), .B(b[46]), .Z(n23001) );
  XNOR U23334 ( .A(n23000), .B(n23001), .Z(n23002) );
  XOR U23335 ( .A(n23003), .B(n23002), .Z(n23105) );
  XNOR U23336 ( .A(n23104), .B(n23105), .Z(n22997) );
  AND U23337 ( .A(a[60]), .B(b[44]), .Z(n22996) );
  XOR U23338 ( .A(n22997), .B(n22996), .Z(n22998) );
  XNOR U23339 ( .A(n22999), .B(n22998), .Z(n23111) );
  XNOR U23340 ( .A(n23110), .B(n23111), .Z(n23113) );
  AND U23341 ( .A(a[62]), .B(b[42]), .Z(n23112) );
  XOR U23342 ( .A(n23113), .B(n23112), .Z(n23114) );
  XNOR U23343 ( .A(n23115), .B(n23114), .Z(n22995) );
  XNOR U23344 ( .A(n22994), .B(n22995), .Z(n22991) );
  XOR U23345 ( .A(n22990), .B(n22991), .Z(n22986) );
  NANDN U23346 ( .A(n22983), .B(n22982), .Z(n22985) );
  XOR U23347 ( .A(n22986), .B(n22985), .Z(n22984) );
  XNOR U23348 ( .A(n22988), .B(n22984), .Z(c[104]) );
  ANDN U23349 ( .B(n22986), .A(n22985), .Z(n22989) );
  NANDN U23350 ( .A(n22986), .B(n22985), .Z(n22987) );
  AND U23351 ( .A(n22988), .B(n22987), .Z(n23241) );
  OR U23352 ( .A(n22989), .B(n23241), .Z(n23239) );
  AND U23353 ( .A(n22991), .B(n22990), .Z(n23243) );
  AND U23354 ( .A(a[61]), .B(b[44]), .Z(n23128) );
  XOR U23355 ( .A(n23127), .B(n23128), .Z(n23130) );
  NANDN U23356 ( .A(n23001), .B(n23000), .Z(n23005) );
  NANDN U23357 ( .A(n23003), .B(n23002), .Z(n23004) );
  AND U23358 ( .A(n23005), .B(n23004), .Z(n23132) );
  AND U23359 ( .A(a[59]), .B(b[46]), .Z(n23131) );
  XNOR U23360 ( .A(n23132), .B(n23131), .Z(n23133) );
  NANDN U23361 ( .A(n23007), .B(n23006), .Z(n23011) );
  NANDN U23362 ( .A(n23009), .B(n23008), .Z(n23010) );
  AND U23363 ( .A(n23011), .B(n23010), .Z(n23144) );
  AND U23364 ( .A(a[57]), .B(b[48]), .Z(n23143) );
  XNOR U23365 ( .A(n23144), .B(n23143), .Z(n23145) );
  NANDN U23366 ( .A(n23013), .B(n23012), .Z(n23017) );
  NANDN U23367 ( .A(n23015), .B(n23014), .Z(n23016) );
  AND U23368 ( .A(n23017), .B(n23016), .Z(n23156) );
  AND U23369 ( .A(a[55]), .B(b[50]), .Z(n23155) );
  XNOR U23370 ( .A(n23156), .B(n23155), .Z(n23157) );
  NANDN U23371 ( .A(n23019), .B(n23018), .Z(n23023) );
  NANDN U23372 ( .A(n23021), .B(n23020), .Z(n23022) );
  AND U23373 ( .A(n23023), .B(n23022), .Z(n23168) );
  AND U23374 ( .A(a[53]), .B(b[52]), .Z(n23167) );
  XNOR U23375 ( .A(n23168), .B(n23167), .Z(n23169) );
  NANDN U23376 ( .A(n23025), .B(n23024), .Z(n23029) );
  NANDN U23377 ( .A(n23027), .B(n23026), .Z(n23028) );
  AND U23378 ( .A(n23029), .B(n23028), .Z(n23180) );
  AND U23379 ( .A(a[51]), .B(b[54]), .Z(n23179) );
  XNOR U23380 ( .A(n23180), .B(n23179), .Z(n23181) );
  AND U23381 ( .A(a[49]), .B(b[56]), .Z(n23192) );
  NANDN U23382 ( .A(n23031), .B(n23030), .Z(n23035) );
  NANDN U23383 ( .A(n23033), .B(n23032), .Z(n23034) );
  AND U23384 ( .A(n23035), .B(n23034), .Z(n23191) );
  XNOR U23385 ( .A(n23192), .B(n23191), .Z(n23194) );
  AND U23386 ( .A(a[48]), .B(b[57]), .Z(n23230) );
  NANDN U23387 ( .A(n23037), .B(n23036), .Z(n23041) );
  NAND U23388 ( .A(n23039), .B(n23038), .Z(n23040) );
  AND U23389 ( .A(n23041), .B(n23040), .Z(n23199) );
  NANDN U23390 ( .A(n23043), .B(n23042), .Z(n23047) );
  NANDN U23391 ( .A(n23045), .B(n23044), .Z(n23046) );
  AND U23392 ( .A(n23047), .B(n23046), .Z(n23222) );
  AND U23393 ( .A(a[46]), .B(b[59]), .Z(n23221) );
  XNOR U23394 ( .A(n23222), .B(n23221), .Z(n23223) );
  NANDN U23395 ( .A(n23049), .B(n23048), .Z(n23053) );
  NANDN U23396 ( .A(n23051), .B(n23050), .Z(n23052) );
  AND U23397 ( .A(n23053), .B(n23052), .Z(n23206) );
  NANDN U23398 ( .A(n23055), .B(n23054), .Z(n23059) );
  NANDN U23399 ( .A(n23057), .B(n23056), .Z(n23058) );
  AND U23400 ( .A(n23059), .B(n23058), .Z(n23216) );
  AND U23401 ( .A(a[44]), .B(b[61]), .Z(n23215) );
  XNOR U23402 ( .A(n23216), .B(n23215), .Z(n23217) );
  NANDN U23403 ( .A(n23061), .B(n23060), .Z(n23065) );
  NANDN U23404 ( .A(n23063), .B(n23062), .Z(n23064) );
  AND U23405 ( .A(n23065), .B(n23064), .Z(n23210) );
  AND U23406 ( .A(b[62]), .B(a[43]), .Z(n23209) );
  XNOR U23407 ( .A(n23210), .B(n23209), .Z(n23211) );
  NAND U23408 ( .A(b[63]), .B(a[42]), .Z(n23212) );
  XOR U23409 ( .A(n23211), .B(n23212), .Z(n23218) );
  XNOR U23410 ( .A(n23217), .B(n23218), .Z(n23203) );
  NAND U23411 ( .A(a[45]), .B(b[60]), .Z(n23204) );
  XNOR U23412 ( .A(n23203), .B(n23204), .Z(n23205) );
  XOR U23413 ( .A(n23206), .B(n23205), .Z(n23224) );
  XNOR U23414 ( .A(n23223), .B(n23224), .Z(n23197) );
  NAND U23415 ( .A(a[47]), .B(b[58]), .Z(n23198) );
  XOR U23416 ( .A(n23197), .B(n23198), .Z(n23200) );
  XOR U23417 ( .A(n23199), .B(n23200), .Z(n23228) );
  NANDN U23418 ( .A(n23067), .B(n23066), .Z(n23071) );
  OR U23419 ( .A(n23069), .B(n23068), .Z(n23070) );
  NAND U23420 ( .A(n23071), .B(n23070), .Z(n23227) );
  XNOR U23421 ( .A(n23228), .B(n23227), .Z(n23229) );
  XNOR U23422 ( .A(n23230), .B(n23229), .Z(n23193) );
  XOR U23423 ( .A(n23194), .B(n23193), .Z(n23188) );
  NANDN U23424 ( .A(n23073), .B(n23072), .Z(n23077) );
  NANDN U23425 ( .A(n23075), .B(n23074), .Z(n23076) );
  AND U23426 ( .A(n23077), .B(n23076), .Z(n23186) );
  AND U23427 ( .A(a[50]), .B(b[55]), .Z(n23185) );
  XNOR U23428 ( .A(n23186), .B(n23185), .Z(n23187) );
  XOR U23429 ( .A(n23188), .B(n23187), .Z(n23182) );
  XNOR U23430 ( .A(n23181), .B(n23182), .Z(n23175) );
  NANDN U23431 ( .A(n23079), .B(n23078), .Z(n23083) );
  NANDN U23432 ( .A(n23081), .B(n23080), .Z(n23082) );
  AND U23433 ( .A(n23083), .B(n23082), .Z(n23174) );
  AND U23434 ( .A(a[52]), .B(b[53]), .Z(n23173) );
  XOR U23435 ( .A(n23174), .B(n23173), .Z(n23176) );
  XOR U23436 ( .A(n23175), .B(n23176), .Z(n23170) );
  XNOR U23437 ( .A(n23169), .B(n23170), .Z(n23163) );
  NANDN U23438 ( .A(n23085), .B(n23084), .Z(n23089) );
  NANDN U23439 ( .A(n23087), .B(n23086), .Z(n23088) );
  AND U23440 ( .A(n23089), .B(n23088), .Z(n23162) );
  AND U23441 ( .A(a[54]), .B(b[51]), .Z(n23161) );
  XOR U23442 ( .A(n23162), .B(n23161), .Z(n23164) );
  XOR U23443 ( .A(n23163), .B(n23164), .Z(n23158) );
  XNOR U23444 ( .A(n23157), .B(n23158), .Z(n23151) );
  NANDN U23445 ( .A(n23091), .B(n23090), .Z(n23095) );
  NANDN U23446 ( .A(n23093), .B(n23092), .Z(n23094) );
  AND U23447 ( .A(n23095), .B(n23094), .Z(n23150) );
  AND U23448 ( .A(a[56]), .B(b[49]), .Z(n23149) );
  XOR U23449 ( .A(n23150), .B(n23149), .Z(n23152) );
  XOR U23450 ( .A(n23151), .B(n23152), .Z(n23146) );
  XNOR U23451 ( .A(n23145), .B(n23146), .Z(n23139) );
  NANDN U23452 ( .A(n23097), .B(n23096), .Z(n23101) );
  NANDN U23453 ( .A(n23099), .B(n23098), .Z(n23100) );
  AND U23454 ( .A(n23101), .B(n23100), .Z(n23138) );
  AND U23455 ( .A(a[58]), .B(b[47]), .Z(n23137) );
  XOR U23456 ( .A(n23138), .B(n23137), .Z(n23140) );
  XOR U23457 ( .A(n23139), .B(n23140), .Z(n23134) );
  XNOR U23458 ( .A(n23133), .B(n23134), .Z(n23236) );
  NANDN U23459 ( .A(n23103), .B(n23102), .Z(n23107) );
  NANDN U23460 ( .A(n23105), .B(n23104), .Z(n23106) );
  AND U23461 ( .A(n23107), .B(n23106), .Z(n23234) );
  AND U23462 ( .A(a[60]), .B(b[45]), .Z(n23233) );
  XNOR U23463 ( .A(n23234), .B(n23233), .Z(n23235) );
  XOR U23464 ( .A(n23236), .B(n23235), .Z(n23129) );
  XOR U23465 ( .A(n23130), .B(n23129), .Z(n23125) );
  AND U23466 ( .A(a[62]), .B(b[43]), .Z(n23123) );
  XNOR U23467 ( .A(n23124), .B(n23123), .Z(n23126) );
  XNOR U23468 ( .A(n23125), .B(n23126), .Z(n23121) );
  AND U23469 ( .A(a[63]), .B(b[42]), .Z(n23119) );
  XNOR U23470 ( .A(n23120), .B(n23119), .Z(n23122) );
  XNOR U23471 ( .A(n23121), .B(n23122), .Z(n23118) );
  XOR U23472 ( .A(n23117), .B(n23118), .Z(n23240) );
  XNOR U23473 ( .A(n23243), .B(n23240), .Z(n23116) );
  XNOR U23474 ( .A(n23239), .B(n23116), .Z(c[105]) );
  IV U23475 ( .A(n23715), .Z(n23246) );
  AND U23476 ( .A(a[63]), .B(b[43]), .Z(n23364) );
  XOR U23477 ( .A(n23363), .B(n23364), .Z(n23365) );
  NANDN U23478 ( .A(n23132), .B(n23131), .Z(n23136) );
  NANDN U23479 ( .A(n23134), .B(n23133), .Z(n23135) );
  AND U23480 ( .A(n23136), .B(n23135), .Z(n23253) );
  NANDN U23481 ( .A(n23138), .B(n23137), .Z(n23142) );
  NANDN U23482 ( .A(n23140), .B(n23139), .Z(n23141) );
  AND U23483 ( .A(n23142), .B(n23141), .Z(n23348) );
  AND U23484 ( .A(a[59]), .B(b[47]), .Z(n23347) );
  XNOR U23485 ( .A(n23348), .B(n23347), .Z(n23349) );
  NANDN U23486 ( .A(n23144), .B(n23143), .Z(n23148) );
  NANDN U23487 ( .A(n23146), .B(n23145), .Z(n23147) );
  AND U23488 ( .A(n23148), .B(n23147), .Z(n23260) );
  NANDN U23489 ( .A(n23150), .B(n23149), .Z(n23154) );
  NANDN U23490 ( .A(n23152), .B(n23151), .Z(n23153) );
  AND U23491 ( .A(n23154), .B(n23153), .Z(n23342) );
  AND U23492 ( .A(a[57]), .B(b[49]), .Z(n23341) );
  XNOR U23493 ( .A(n23342), .B(n23341), .Z(n23343) );
  NANDN U23494 ( .A(n23156), .B(n23155), .Z(n23160) );
  NANDN U23495 ( .A(n23158), .B(n23157), .Z(n23159) );
  AND U23496 ( .A(n23160), .B(n23159), .Z(n23266) );
  NANDN U23497 ( .A(n23162), .B(n23161), .Z(n23166) );
  NANDN U23498 ( .A(n23164), .B(n23163), .Z(n23165) );
  AND U23499 ( .A(n23166), .B(n23165), .Z(n23336) );
  AND U23500 ( .A(a[55]), .B(b[51]), .Z(n23335) );
  XNOR U23501 ( .A(n23336), .B(n23335), .Z(n23337) );
  NANDN U23502 ( .A(n23168), .B(n23167), .Z(n23172) );
  NANDN U23503 ( .A(n23170), .B(n23169), .Z(n23171) );
  AND U23504 ( .A(n23172), .B(n23171), .Z(n23272) );
  NANDN U23505 ( .A(n23174), .B(n23173), .Z(n23178) );
  NANDN U23506 ( .A(n23176), .B(n23175), .Z(n23177) );
  AND U23507 ( .A(n23178), .B(n23177), .Z(n23330) );
  AND U23508 ( .A(a[53]), .B(b[53]), .Z(n23329) );
  XNOR U23509 ( .A(n23330), .B(n23329), .Z(n23331) );
  NANDN U23510 ( .A(n23180), .B(n23179), .Z(n23184) );
  NANDN U23511 ( .A(n23182), .B(n23181), .Z(n23183) );
  AND U23512 ( .A(n23184), .B(n23183), .Z(n23278) );
  NANDN U23513 ( .A(n23186), .B(n23185), .Z(n23190) );
  NANDN U23514 ( .A(n23188), .B(n23187), .Z(n23189) );
  AND U23515 ( .A(n23190), .B(n23189), .Z(n23324) );
  AND U23516 ( .A(a[51]), .B(b[55]), .Z(n23323) );
  XNOR U23517 ( .A(n23324), .B(n23323), .Z(n23325) );
  NANDN U23518 ( .A(n23192), .B(n23191), .Z(n23196) );
  NAND U23519 ( .A(n23194), .B(n23193), .Z(n23195) );
  AND U23520 ( .A(n23196), .B(n23195), .Z(n23283) );
  NANDN U23521 ( .A(n23198), .B(n23197), .Z(n23202) );
  OR U23522 ( .A(n23200), .B(n23199), .Z(n23201) );
  AND U23523 ( .A(n23202), .B(n23201), .Z(n23288) );
  AND U23524 ( .A(a[48]), .B(b[58]), .Z(n23287) );
  XNOR U23525 ( .A(n23288), .B(n23287), .Z(n23289) );
  NANDN U23526 ( .A(n23204), .B(n23203), .Z(n23208) );
  NANDN U23527 ( .A(n23206), .B(n23205), .Z(n23207) );
  AND U23528 ( .A(n23208), .B(n23207), .Z(n23300) );
  AND U23529 ( .A(a[46]), .B(b[60]), .Z(n23299) );
  XNOR U23530 ( .A(n23300), .B(n23299), .Z(n23301) );
  NANDN U23531 ( .A(n23210), .B(n23209), .Z(n23214) );
  NANDN U23532 ( .A(n23212), .B(n23211), .Z(n23213) );
  AND U23533 ( .A(n23214), .B(n23213), .Z(n23312) );
  AND U23534 ( .A(b[62]), .B(a[44]), .Z(n23311) );
  XNOR U23535 ( .A(n23312), .B(n23311), .Z(n23313) );
  NAND U23536 ( .A(b[63]), .B(a[43]), .Z(n23314) );
  XNOR U23537 ( .A(n23313), .B(n23314), .Z(n23307) );
  NANDN U23538 ( .A(n23216), .B(n23215), .Z(n23220) );
  NANDN U23539 ( .A(n23218), .B(n23217), .Z(n23219) );
  AND U23540 ( .A(n23220), .B(n23219), .Z(n23306) );
  AND U23541 ( .A(a[45]), .B(b[61]), .Z(n23305) );
  XOR U23542 ( .A(n23306), .B(n23305), .Z(n23308) );
  XOR U23543 ( .A(n23307), .B(n23308), .Z(n23302) );
  XNOR U23544 ( .A(n23301), .B(n23302), .Z(n23295) );
  NANDN U23545 ( .A(n23222), .B(n23221), .Z(n23226) );
  NANDN U23546 ( .A(n23224), .B(n23223), .Z(n23225) );
  AND U23547 ( .A(n23226), .B(n23225), .Z(n23294) );
  AND U23548 ( .A(a[47]), .B(b[59]), .Z(n23293) );
  XOR U23549 ( .A(n23294), .B(n23293), .Z(n23296) );
  XOR U23550 ( .A(n23295), .B(n23296), .Z(n23290) );
  XNOR U23551 ( .A(n23289), .B(n23290), .Z(n23317) );
  NANDN U23552 ( .A(n23228), .B(n23227), .Z(n23232) );
  NANDN U23553 ( .A(n23230), .B(n23229), .Z(n23231) );
  NAND U23554 ( .A(n23232), .B(n23231), .Z(n23318) );
  XNOR U23555 ( .A(n23317), .B(n23318), .Z(n23319) );
  NAND U23556 ( .A(a[49]), .B(b[57]), .Z(n23320) );
  XNOR U23557 ( .A(n23319), .B(n23320), .Z(n23281) );
  NAND U23558 ( .A(a[50]), .B(b[56]), .Z(n23282) );
  XOR U23559 ( .A(n23281), .B(n23282), .Z(n23284) );
  XOR U23560 ( .A(n23283), .B(n23284), .Z(n23326) );
  XNOR U23561 ( .A(n23325), .B(n23326), .Z(n23275) );
  NAND U23562 ( .A(a[52]), .B(b[54]), .Z(n23276) );
  XNOR U23563 ( .A(n23275), .B(n23276), .Z(n23277) );
  XOR U23564 ( .A(n23278), .B(n23277), .Z(n23332) );
  XNOR U23565 ( .A(n23331), .B(n23332), .Z(n23269) );
  NAND U23566 ( .A(a[54]), .B(b[52]), .Z(n23270) );
  XNOR U23567 ( .A(n23269), .B(n23270), .Z(n23271) );
  XOR U23568 ( .A(n23272), .B(n23271), .Z(n23338) );
  XNOR U23569 ( .A(n23337), .B(n23338), .Z(n23263) );
  NAND U23570 ( .A(a[56]), .B(b[50]), .Z(n23264) );
  XNOR U23571 ( .A(n23263), .B(n23264), .Z(n23265) );
  XOR U23572 ( .A(n23266), .B(n23265), .Z(n23344) );
  XNOR U23573 ( .A(n23343), .B(n23344), .Z(n23257) );
  NAND U23574 ( .A(a[58]), .B(b[48]), .Z(n23258) );
  XNOR U23575 ( .A(n23257), .B(n23258), .Z(n23259) );
  XOR U23576 ( .A(n23260), .B(n23259), .Z(n23350) );
  XNOR U23577 ( .A(n23349), .B(n23350), .Z(n23251) );
  NAND U23578 ( .A(a[60]), .B(b[46]), .Z(n23252) );
  XOR U23579 ( .A(n23251), .B(n23252), .Z(n23254) );
  XOR U23580 ( .A(n23253), .B(n23254), .Z(n23356) );
  AND U23581 ( .A(a[61]), .B(b[45]), .Z(n23354) );
  NANDN U23582 ( .A(n23234), .B(n23233), .Z(n23238) );
  NAND U23583 ( .A(n23236), .B(n23235), .Z(n23237) );
  AND U23584 ( .A(n23238), .B(n23237), .Z(n23353) );
  XNOR U23585 ( .A(n23354), .B(n23353), .Z(n23355) );
  XOR U23586 ( .A(n23356), .B(n23355), .Z(n23360) );
  AND U23587 ( .A(a[62]), .B(b[44]), .Z(n23359) );
  XNOR U23588 ( .A(n23360), .B(n23359), .Z(n23362) );
  XOR U23589 ( .A(n23361), .B(n23362), .Z(n23366) );
  XOR U23590 ( .A(n23365), .B(n23366), .Z(n23250) );
  XNOR U23591 ( .A(n23249), .B(n23250), .Z(n23714) );
  XOR U23592 ( .A(n23246), .B(n23714), .Z(n23247) );
  NAND U23593 ( .A(n23240), .B(n23239), .Z(n23245) );
  OR U23594 ( .A(n23241), .B(n23240), .Z(n23242) );
  NAND U23595 ( .A(n23243), .B(n23242), .Z(n23244) );
  NAND U23596 ( .A(n23245), .B(n23244), .Z(n23716) );
  XOR U23597 ( .A(n23247), .B(n23716), .Z(c[106]) );
  OR U23598 ( .A(n23714), .B(n23246), .Z(n23711) );
  NAND U23599 ( .A(n23247), .B(n23716), .Z(n23248) );
  AND U23600 ( .A(n23711), .B(n23248), .Z(n23482) );
  NOR U23601 ( .A(n23250), .B(n23249), .Z(n23709) );
  NANDN U23602 ( .A(n23252), .B(n23251), .Z(n23256) );
  OR U23603 ( .A(n23254), .B(n23253), .Z(n23255) );
  AND U23604 ( .A(n23256), .B(n23255), .Z(n23376) );
  AND U23605 ( .A(a[61]), .B(b[46]), .Z(n23375) );
  XNOR U23606 ( .A(n23376), .B(n23375), .Z(n23377) );
  NANDN U23607 ( .A(n23258), .B(n23257), .Z(n23262) );
  NANDN U23608 ( .A(n23260), .B(n23259), .Z(n23261) );
  AND U23609 ( .A(n23262), .B(n23261), .Z(n23388) );
  AND U23610 ( .A(a[59]), .B(b[48]), .Z(n23387) );
  XNOR U23611 ( .A(n23388), .B(n23387), .Z(n23389) );
  NANDN U23612 ( .A(n23264), .B(n23263), .Z(n23268) );
  NANDN U23613 ( .A(n23266), .B(n23265), .Z(n23267) );
  AND U23614 ( .A(n23268), .B(n23267), .Z(n23394) );
  AND U23615 ( .A(a[57]), .B(b[50]), .Z(n23393) );
  XNOR U23616 ( .A(n23394), .B(n23393), .Z(n23395) );
  NANDN U23617 ( .A(n23270), .B(n23269), .Z(n23274) );
  NANDN U23618 ( .A(n23272), .B(n23271), .Z(n23273) );
  AND U23619 ( .A(n23274), .B(n23273), .Z(n23400) );
  AND U23620 ( .A(a[55]), .B(b[52]), .Z(n23399) );
  XNOR U23621 ( .A(n23400), .B(n23399), .Z(n23401) );
  NANDN U23622 ( .A(n23276), .B(n23275), .Z(n23280) );
  NANDN U23623 ( .A(n23278), .B(n23277), .Z(n23279) );
  AND U23624 ( .A(n23280), .B(n23279), .Z(n23412) );
  AND U23625 ( .A(a[53]), .B(b[54]), .Z(n23411) );
  XNOR U23626 ( .A(n23412), .B(n23411), .Z(n23413) );
  AND U23627 ( .A(a[51]), .B(b[56]), .Z(n23424) );
  NANDN U23628 ( .A(n23282), .B(n23281), .Z(n23286) );
  NANDN U23629 ( .A(n23284), .B(n23283), .Z(n23285) );
  AND U23630 ( .A(n23286), .B(n23285), .Z(n23423) );
  XNOR U23631 ( .A(n23424), .B(n23423), .Z(n23426) );
  AND U23632 ( .A(a[50]), .B(b[57]), .Z(n23462) );
  NANDN U23633 ( .A(n23288), .B(n23287), .Z(n23292) );
  NANDN U23634 ( .A(n23290), .B(n23289), .Z(n23291) );
  AND U23635 ( .A(n23292), .B(n23291), .Z(n23431) );
  NANDN U23636 ( .A(n23294), .B(n23293), .Z(n23298) );
  NANDN U23637 ( .A(n23296), .B(n23295), .Z(n23297) );
  AND U23638 ( .A(n23298), .B(n23297), .Z(n23454) );
  AND U23639 ( .A(a[48]), .B(b[59]), .Z(n23453) );
  XNOR U23640 ( .A(n23454), .B(n23453), .Z(n23455) );
  NANDN U23641 ( .A(n23300), .B(n23299), .Z(n23304) );
  NANDN U23642 ( .A(n23302), .B(n23301), .Z(n23303) );
  AND U23643 ( .A(n23304), .B(n23303), .Z(n23450) );
  NANDN U23644 ( .A(n23306), .B(n23305), .Z(n23310) );
  NANDN U23645 ( .A(n23308), .B(n23307), .Z(n23309) );
  AND U23646 ( .A(n23310), .B(n23309), .Z(n23442) );
  AND U23647 ( .A(a[46]), .B(b[61]), .Z(n23441) );
  XNOR U23648 ( .A(n23442), .B(n23441), .Z(n23443) );
  NANDN U23649 ( .A(n23312), .B(n23311), .Z(n23316) );
  NANDN U23650 ( .A(n23314), .B(n23313), .Z(n23315) );
  AND U23651 ( .A(n23316), .B(n23315), .Z(n23438) );
  AND U23652 ( .A(b[62]), .B(a[45]), .Z(n23435) );
  NAND U23653 ( .A(b[63]), .B(a[44]), .Z(n23436) );
  XNOR U23654 ( .A(n23435), .B(n23436), .Z(n23437) );
  XOR U23655 ( .A(n23438), .B(n23437), .Z(n23444) );
  XNOR U23656 ( .A(n23443), .B(n23444), .Z(n23447) );
  NAND U23657 ( .A(a[47]), .B(b[60]), .Z(n23448) );
  XNOR U23658 ( .A(n23447), .B(n23448), .Z(n23449) );
  XOR U23659 ( .A(n23450), .B(n23449), .Z(n23456) );
  XNOR U23660 ( .A(n23455), .B(n23456), .Z(n23429) );
  NAND U23661 ( .A(a[49]), .B(b[58]), .Z(n23430) );
  XOR U23662 ( .A(n23429), .B(n23430), .Z(n23432) );
  XOR U23663 ( .A(n23431), .B(n23432), .Z(n23460) );
  NANDN U23664 ( .A(n23318), .B(n23317), .Z(n23322) );
  NANDN U23665 ( .A(n23320), .B(n23319), .Z(n23321) );
  AND U23666 ( .A(n23322), .B(n23321), .Z(n23459) );
  XNOR U23667 ( .A(n23460), .B(n23459), .Z(n23461) );
  XNOR U23668 ( .A(n23462), .B(n23461), .Z(n23425) );
  XOR U23669 ( .A(n23426), .B(n23425), .Z(n23420) );
  NANDN U23670 ( .A(n23324), .B(n23323), .Z(n23328) );
  NANDN U23671 ( .A(n23326), .B(n23325), .Z(n23327) );
  AND U23672 ( .A(n23328), .B(n23327), .Z(n23418) );
  AND U23673 ( .A(a[52]), .B(b[55]), .Z(n23417) );
  XNOR U23674 ( .A(n23418), .B(n23417), .Z(n23419) );
  XOR U23675 ( .A(n23420), .B(n23419), .Z(n23414) );
  XNOR U23676 ( .A(n23413), .B(n23414), .Z(n23407) );
  NANDN U23677 ( .A(n23330), .B(n23329), .Z(n23334) );
  NANDN U23678 ( .A(n23332), .B(n23331), .Z(n23333) );
  AND U23679 ( .A(n23334), .B(n23333), .Z(n23406) );
  AND U23680 ( .A(a[54]), .B(b[53]), .Z(n23405) );
  XOR U23681 ( .A(n23406), .B(n23405), .Z(n23408) );
  XOR U23682 ( .A(n23407), .B(n23408), .Z(n23402) );
  XNOR U23683 ( .A(n23401), .B(n23402), .Z(n23467) );
  NANDN U23684 ( .A(n23336), .B(n23335), .Z(n23340) );
  NANDN U23685 ( .A(n23338), .B(n23337), .Z(n23339) );
  AND U23686 ( .A(n23340), .B(n23339), .Z(n23466) );
  AND U23687 ( .A(a[56]), .B(b[51]), .Z(n23465) );
  XOR U23688 ( .A(n23466), .B(n23465), .Z(n23468) );
  XOR U23689 ( .A(n23467), .B(n23468), .Z(n23396) );
  XNOR U23690 ( .A(n23395), .B(n23396), .Z(n23473) );
  NANDN U23691 ( .A(n23342), .B(n23341), .Z(n23346) );
  NANDN U23692 ( .A(n23344), .B(n23343), .Z(n23345) );
  AND U23693 ( .A(n23346), .B(n23345), .Z(n23472) );
  AND U23694 ( .A(a[58]), .B(b[49]), .Z(n23471) );
  XOR U23695 ( .A(n23472), .B(n23471), .Z(n23474) );
  XOR U23696 ( .A(n23473), .B(n23474), .Z(n23390) );
  XNOR U23697 ( .A(n23389), .B(n23390), .Z(n23383) );
  NANDN U23698 ( .A(n23348), .B(n23347), .Z(n23352) );
  NANDN U23699 ( .A(n23350), .B(n23349), .Z(n23351) );
  AND U23700 ( .A(n23352), .B(n23351), .Z(n23382) );
  AND U23701 ( .A(a[60]), .B(b[47]), .Z(n23381) );
  XOR U23702 ( .A(n23382), .B(n23381), .Z(n23384) );
  XOR U23703 ( .A(n23383), .B(n23384), .Z(n23378) );
  XNOR U23704 ( .A(n23377), .B(n23378), .Z(n23371) );
  NANDN U23705 ( .A(n23354), .B(n23353), .Z(n23358) );
  NANDN U23706 ( .A(n23356), .B(n23355), .Z(n23357) );
  AND U23707 ( .A(n23358), .B(n23357), .Z(n23369) );
  NAND U23708 ( .A(a[62]), .B(b[45]), .Z(n23370) );
  XOR U23709 ( .A(n23369), .B(n23370), .Z(n23372) );
  XOR U23710 ( .A(n23371), .B(n23372), .Z(n23479) );
  NAND U23711 ( .A(a[63]), .B(b[44]), .Z(n23477) );
  XOR U23712 ( .A(n23477), .B(n23478), .Z(n23480) );
  XOR U23713 ( .A(n23479), .B(n23480), .Z(n23368) );
  XOR U23714 ( .A(n23368), .B(n23367), .Z(n23710) );
  XNOR U23715 ( .A(n23709), .B(n23710), .Z(n23481) );
  XNOR U23716 ( .A(n23482), .B(n23481), .Z(c[107]) );
  IV U23717 ( .A(n23486), .Z(n23705) );
  NANDN U23718 ( .A(n23370), .B(n23369), .Z(n23374) );
  NANDN U23719 ( .A(n23372), .B(n23371), .Z(n23373) );
  AND U23720 ( .A(n23374), .B(n23373), .Z(n23489) );
  AND U23721 ( .A(a[63]), .B(b[45]), .Z(n23488) );
  XNOR U23722 ( .A(n23489), .B(n23488), .Z(n23490) );
  NANDN U23723 ( .A(n23376), .B(n23375), .Z(n23380) );
  NANDN U23724 ( .A(n23378), .B(n23377), .Z(n23379) );
  AND U23725 ( .A(n23380), .B(n23379), .Z(n23497) );
  NANDN U23726 ( .A(n23382), .B(n23381), .Z(n23386) );
  NANDN U23727 ( .A(n23384), .B(n23383), .Z(n23385) );
  AND U23728 ( .A(n23386), .B(n23385), .Z(n23591) );
  AND U23729 ( .A(a[61]), .B(b[47]), .Z(n23590) );
  XNOR U23730 ( .A(n23591), .B(n23590), .Z(n23592) );
  NANDN U23731 ( .A(n23388), .B(n23387), .Z(n23392) );
  NANDN U23732 ( .A(n23390), .B(n23389), .Z(n23391) );
  AND U23733 ( .A(n23392), .B(n23391), .Z(n23503) );
  NANDN U23734 ( .A(n23394), .B(n23393), .Z(n23398) );
  NANDN U23735 ( .A(n23396), .B(n23395), .Z(n23397) );
  AND U23736 ( .A(n23398), .B(n23397), .Z(n23580) );
  NANDN U23737 ( .A(n23400), .B(n23399), .Z(n23404) );
  NANDN U23738 ( .A(n23402), .B(n23401), .Z(n23403) );
  AND U23739 ( .A(n23404), .B(n23403), .Z(n23508) );
  NANDN U23740 ( .A(n23406), .B(n23405), .Z(n23410) );
  NANDN U23741 ( .A(n23408), .B(n23407), .Z(n23409) );
  AND U23742 ( .A(n23410), .B(n23409), .Z(n23567) );
  AND U23743 ( .A(a[55]), .B(b[53]), .Z(n23566) );
  XNOR U23744 ( .A(n23567), .B(n23566), .Z(n23568) );
  NANDN U23745 ( .A(n23412), .B(n23411), .Z(n23416) );
  NANDN U23746 ( .A(n23414), .B(n23413), .Z(n23415) );
  AND U23747 ( .A(n23416), .B(n23415), .Z(n23563) );
  NANDN U23748 ( .A(n23418), .B(n23417), .Z(n23422) );
  NANDN U23749 ( .A(n23420), .B(n23419), .Z(n23421) );
  AND U23750 ( .A(n23422), .B(n23421), .Z(n23555) );
  AND U23751 ( .A(a[53]), .B(b[55]), .Z(n23554) );
  XNOR U23752 ( .A(n23555), .B(n23554), .Z(n23556) );
  NANDN U23753 ( .A(n23424), .B(n23423), .Z(n23428) );
  NAND U23754 ( .A(n23426), .B(n23425), .Z(n23427) );
  AND U23755 ( .A(n23428), .B(n23427), .Z(n23514) );
  NANDN U23756 ( .A(n23430), .B(n23429), .Z(n23434) );
  OR U23757 ( .A(n23432), .B(n23431), .Z(n23433) );
  AND U23758 ( .A(n23434), .B(n23433), .Z(n23519) );
  AND U23759 ( .A(a[50]), .B(b[58]), .Z(n23518) );
  XNOR U23760 ( .A(n23519), .B(n23518), .Z(n23520) );
  NANDN U23761 ( .A(n23436), .B(n23435), .Z(n23440) );
  NANDN U23762 ( .A(n23438), .B(n23437), .Z(n23439) );
  AND U23763 ( .A(n23440), .B(n23439), .Z(n23543) );
  AND U23764 ( .A(b[62]), .B(a[46]), .Z(n23542) );
  XNOR U23765 ( .A(n23543), .B(n23542), .Z(n23544) );
  NAND U23766 ( .A(b[63]), .B(a[45]), .Z(n23545) );
  XNOR U23767 ( .A(n23544), .B(n23545), .Z(n23539) );
  NANDN U23768 ( .A(n23442), .B(n23441), .Z(n23446) );
  NANDN U23769 ( .A(n23444), .B(n23443), .Z(n23445) );
  AND U23770 ( .A(n23446), .B(n23445), .Z(n23537) );
  AND U23771 ( .A(a[47]), .B(b[61]), .Z(n23536) );
  XNOR U23772 ( .A(n23537), .B(n23536), .Z(n23538) );
  XOR U23773 ( .A(n23539), .B(n23538), .Z(n23532) );
  AND U23774 ( .A(a[48]), .B(b[60]), .Z(n23531) );
  NANDN U23775 ( .A(n23448), .B(n23447), .Z(n23452) );
  NANDN U23776 ( .A(n23450), .B(n23449), .Z(n23451) );
  AND U23777 ( .A(n23452), .B(n23451), .Z(n23530) );
  XOR U23778 ( .A(n23531), .B(n23530), .Z(n23533) );
  XOR U23779 ( .A(n23532), .B(n23533), .Z(n23527) );
  NANDN U23780 ( .A(n23454), .B(n23453), .Z(n23458) );
  NANDN U23781 ( .A(n23456), .B(n23455), .Z(n23457) );
  AND U23782 ( .A(n23458), .B(n23457), .Z(n23525) );
  AND U23783 ( .A(a[49]), .B(b[59]), .Z(n23524) );
  XNOR U23784 ( .A(n23525), .B(n23524), .Z(n23526) );
  XOR U23785 ( .A(n23527), .B(n23526), .Z(n23521) );
  XNOR U23786 ( .A(n23520), .B(n23521), .Z(n23548) );
  NANDN U23787 ( .A(n23460), .B(n23459), .Z(n23464) );
  NANDN U23788 ( .A(n23462), .B(n23461), .Z(n23463) );
  NAND U23789 ( .A(n23464), .B(n23463), .Z(n23549) );
  XNOR U23790 ( .A(n23548), .B(n23549), .Z(n23550) );
  NAND U23791 ( .A(a[51]), .B(b[57]), .Z(n23551) );
  XNOR U23792 ( .A(n23550), .B(n23551), .Z(n23512) );
  NAND U23793 ( .A(a[52]), .B(b[56]), .Z(n23513) );
  XOR U23794 ( .A(n23512), .B(n23513), .Z(n23515) );
  XOR U23795 ( .A(n23514), .B(n23515), .Z(n23557) );
  XNOR U23796 ( .A(n23556), .B(n23557), .Z(n23560) );
  NAND U23797 ( .A(a[54]), .B(b[54]), .Z(n23561) );
  XNOR U23798 ( .A(n23560), .B(n23561), .Z(n23562) );
  XOR U23799 ( .A(n23563), .B(n23562), .Z(n23569) );
  XNOR U23800 ( .A(n23568), .B(n23569), .Z(n23506) );
  NAND U23801 ( .A(a[56]), .B(b[52]), .Z(n23507) );
  XOR U23802 ( .A(n23506), .B(n23507), .Z(n23509) );
  XOR U23803 ( .A(n23508), .B(n23509), .Z(n23574) );
  AND U23804 ( .A(a[57]), .B(b[51]), .Z(n23573) );
  NANDN U23805 ( .A(n23466), .B(n23465), .Z(n23470) );
  NANDN U23806 ( .A(n23468), .B(n23467), .Z(n23469) );
  AND U23807 ( .A(n23470), .B(n23469), .Z(n23572) );
  XOR U23808 ( .A(n23573), .B(n23572), .Z(n23575) );
  XOR U23809 ( .A(n23574), .B(n23575), .Z(n23579) );
  AND U23810 ( .A(a[58]), .B(b[50]), .Z(n23578) );
  XOR U23811 ( .A(n23579), .B(n23578), .Z(n23581) );
  XOR U23812 ( .A(n23580), .B(n23581), .Z(n23586) );
  AND U23813 ( .A(a[59]), .B(b[49]), .Z(n23585) );
  NANDN U23814 ( .A(n23472), .B(n23471), .Z(n23476) );
  NANDN U23815 ( .A(n23474), .B(n23473), .Z(n23475) );
  AND U23816 ( .A(n23476), .B(n23475), .Z(n23584) );
  XOR U23817 ( .A(n23585), .B(n23584), .Z(n23587) );
  XOR U23818 ( .A(n23586), .B(n23587), .Z(n23501) );
  AND U23819 ( .A(a[60]), .B(b[48]), .Z(n23500) );
  XNOR U23820 ( .A(n23501), .B(n23500), .Z(n23502) );
  XOR U23821 ( .A(n23503), .B(n23502), .Z(n23593) );
  XNOR U23822 ( .A(n23592), .B(n23593), .Z(n23494) );
  NAND U23823 ( .A(a[62]), .B(b[46]), .Z(n23495) );
  XNOR U23824 ( .A(n23494), .B(n23495), .Z(n23496) );
  XOR U23825 ( .A(n23497), .B(n23496), .Z(n23491) );
  XNOR U23826 ( .A(n23490), .B(n23491), .Z(n23597) );
  XNOR U23827 ( .A(n23597), .B(n23596), .Z(n23706) );
  XOR U23828 ( .A(n23705), .B(n23706), .Z(n23485) );
  NANDN U23829 ( .A(n23709), .B(n23710), .Z(n23708) );
  NAND U23830 ( .A(n23482), .B(n23481), .Z(n23483) );
  NAND U23831 ( .A(n23708), .B(n23483), .Z(n23484) );
  XNOR U23832 ( .A(n23485), .B(n23484), .Z(c[108]) );
  NAND U23833 ( .A(n23485), .B(n23484), .Z(n23487) );
  NANDN U23834 ( .A(n23486), .B(n23706), .Z(n23707) );
  AND U23835 ( .A(n23487), .B(n23707), .Z(n23599) );
  NANDN U23836 ( .A(n23489), .B(n23488), .Z(n23493) );
  NANDN U23837 ( .A(n23491), .B(n23490), .Z(n23492) );
  AND U23838 ( .A(n23493), .B(n23492), .Z(n23702) );
  NANDN U23839 ( .A(n23495), .B(n23494), .Z(n23499) );
  NANDN U23840 ( .A(n23497), .B(n23496), .Z(n23498) );
  AND U23841 ( .A(n23499), .B(n23498), .Z(n23601) );
  AND U23842 ( .A(a[63]), .B(b[46]), .Z(n23600) );
  XNOR U23843 ( .A(n23601), .B(n23600), .Z(n23602) );
  NANDN U23844 ( .A(n23501), .B(n23500), .Z(n23505) );
  NANDN U23845 ( .A(n23503), .B(n23502), .Z(n23504) );
  AND U23846 ( .A(n23505), .B(n23504), .Z(n23613) );
  AND U23847 ( .A(a[61]), .B(b[48]), .Z(n23612) );
  XNOR U23848 ( .A(n23613), .B(n23612), .Z(n23614) );
  NANDN U23849 ( .A(n23507), .B(n23506), .Z(n23511) );
  OR U23850 ( .A(n23509), .B(n23508), .Z(n23510) );
  AND U23851 ( .A(n23511), .B(n23510), .Z(n23637) );
  AND U23852 ( .A(a[57]), .B(b[52]), .Z(n23636) );
  XNOR U23853 ( .A(n23637), .B(n23636), .Z(n23638) );
  AND U23854 ( .A(a[53]), .B(b[56]), .Z(n23661) );
  NANDN U23855 ( .A(n23513), .B(n23512), .Z(n23517) );
  NANDN U23856 ( .A(n23515), .B(n23514), .Z(n23516) );
  AND U23857 ( .A(n23517), .B(n23516), .Z(n23660) );
  XNOR U23858 ( .A(n23661), .B(n23660), .Z(n23663) );
  AND U23859 ( .A(a[52]), .B(b[57]), .Z(n23699) );
  NANDN U23860 ( .A(n23519), .B(n23518), .Z(n23523) );
  NANDN U23861 ( .A(n23521), .B(n23520), .Z(n23522) );
  AND U23862 ( .A(n23523), .B(n23522), .Z(n23668) );
  NANDN U23863 ( .A(n23525), .B(n23524), .Z(n23529) );
  NANDN U23864 ( .A(n23527), .B(n23526), .Z(n23528) );
  AND U23865 ( .A(n23529), .B(n23528), .Z(n23691) );
  AND U23866 ( .A(a[50]), .B(b[59]), .Z(n23690) );
  XNOR U23867 ( .A(n23691), .B(n23690), .Z(n23692) );
  NANDN U23868 ( .A(n23531), .B(n23530), .Z(n23535) );
  OR U23869 ( .A(n23533), .B(n23532), .Z(n23534) );
  AND U23870 ( .A(n23535), .B(n23534), .Z(n23674) );
  NANDN U23871 ( .A(n23537), .B(n23536), .Z(n23541) );
  NAND U23872 ( .A(n23539), .B(n23538), .Z(n23540) );
  AND U23873 ( .A(n23541), .B(n23540), .Z(n23685) );
  AND U23874 ( .A(a[48]), .B(b[61]), .Z(n23684) );
  XNOR U23875 ( .A(n23685), .B(n23684), .Z(n23686) );
  NANDN U23876 ( .A(n23543), .B(n23542), .Z(n23547) );
  NANDN U23877 ( .A(n23545), .B(n23544), .Z(n23546) );
  AND U23878 ( .A(n23547), .B(n23546), .Z(n23681) );
  AND U23879 ( .A(b[62]), .B(a[47]), .Z(n23678) );
  NAND U23880 ( .A(b[63]), .B(a[46]), .Z(n23679) );
  XNOR U23881 ( .A(n23678), .B(n23679), .Z(n23680) );
  XOR U23882 ( .A(n23681), .B(n23680), .Z(n23687) );
  XNOR U23883 ( .A(n23686), .B(n23687), .Z(n23672) );
  NAND U23884 ( .A(a[49]), .B(b[60]), .Z(n23673) );
  XOR U23885 ( .A(n23672), .B(n23673), .Z(n23675) );
  XOR U23886 ( .A(n23674), .B(n23675), .Z(n23693) );
  XNOR U23887 ( .A(n23692), .B(n23693), .Z(n23666) );
  NAND U23888 ( .A(a[51]), .B(b[58]), .Z(n23667) );
  XOR U23889 ( .A(n23666), .B(n23667), .Z(n23669) );
  XOR U23890 ( .A(n23668), .B(n23669), .Z(n23697) );
  NANDN U23891 ( .A(n23549), .B(n23548), .Z(n23553) );
  NANDN U23892 ( .A(n23551), .B(n23550), .Z(n23552) );
  AND U23893 ( .A(n23553), .B(n23552), .Z(n23696) );
  XNOR U23894 ( .A(n23697), .B(n23696), .Z(n23698) );
  XNOR U23895 ( .A(n23699), .B(n23698), .Z(n23662) );
  XOR U23896 ( .A(n23663), .B(n23662), .Z(n23656) );
  NANDN U23897 ( .A(n23555), .B(n23554), .Z(n23559) );
  NANDN U23898 ( .A(n23557), .B(n23556), .Z(n23558) );
  AND U23899 ( .A(n23559), .B(n23558), .Z(n23655) );
  AND U23900 ( .A(a[54]), .B(b[55]), .Z(n23654) );
  XOR U23901 ( .A(n23655), .B(n23654), .Z(n23657) );
  XOR U23902 ( .A(n23656), .B(n23657), .Z(n23650) );
  AND U23903 ( .A(a[55]), .B(b[54]), .Z(n23649) );
  NANDN U23904 ( .A(n23561), .B(n23560), .Z(n23565) );
  NANDN U23905 ( .A(n23563), .B(n23562), .Z(n23564) );
  AND U23906 ( .A(n23565), .B(n23564), .Z(n23648) );
  XOR U23907 ( .A(n23649), .B(n23648), .Z(n23651) );
  XOR U23908 ( .A(n23650), .B(n23651), .Z(n23645) );
  NANDN U23909 ( .A(n23567), .B(n23566), .Z(n23571) );
  NANDN U23910 ( .A(n23569), .B(n23568), .Z(n23570) );
  AND U23911 ( .A(n23571), .B(n23570), .Z(n23643) );
  AND U23912 ( .A(a[56]), .B(b[53]), .Z(n23642) );
  XNOR U23913 ( .A(n23643), .B(n23642), .Z(n23644) );
  XOR U23914 ( .A(n23645), .B(n23644), .Z(n23639) );
  XNOR U23915 ( .A(n23638), .B(n23639), .Z(n23633) );
  NANDN U23916 ( .A(n23573), .B(n23572), .Z(n23577) );
  OR U23917 ( .A(n23575), .B(n23574), .Z(n23576) );
  AND U23918 ( .A(n23577), .B(n23576), .Z(n23630) );
  NAND U23919 ( .A(a[58]), .B(b[51]), .Z(n23631) );
  XNOR U23920 ( .A(n23630), .B(n23631), .Z(n23632) );
  XOR U23921 ( .A(n23633), .B(n23632), .Z(n23626) );
  AND U23922 ( .A(a[59]), .B(b[50]), .Z(n23625) );
  NANDN U23923 ( .A(n23579), .B(n23578), .Z(n23583) );
  OR U23924 ( .A(n23581), .B(n23580), .Z(n23582) );
  AND U23925 ( .A(n23583), .B(n23582), .Z(n23624) );
  XOR U23926 ( .A(n23625), .B(n23624), .Z(n23627) );
  XOR U23927 ( .A(n23626), .B(n23627), .Z(n23621) );
  NANDN U23928 ( .A(n23585), .B(n23584), .Z(n23589) );
  OR U23929 ( .A(n23587), .B(n23586), .Z(n23588) );
  AND U23930 ( .A(n23589), .B(n23588), .Z(n23618) );
  NAND U23931 ( .A(a[60]), .B(b[49]), .Z(n23619) );
  XNOR U23932 ( .A(n23618), .B(n23619), .Z(n23620) );
  XOR U23933 ( .A(n23621), .B(n23620), .Z(n23615) );
  XNOR U23934 ( .A(n23614), .B(n23615), .Z(n23608) );
  NANDN U23935 ( .A(n23591), .B(n23590), .Z(n23595) );
  NANDN U23936 ( .A(n23593), .B(n23592), .Z(n23594) );
  AND U23937 ( .A(n23595), .B(n23594), .Z(n23607) );
  AND U23938 ( .A(a[62]), .B(b[47]), .Z(n23606) );
  XOR U23939 ( .A(n23607), .B(n23606), .Z(n23609) );
  XOR U23940 ( .A(n23608), .B(n23609), .Z(n23603) );
  XNOR U23941 ( .A(n23602), .B(n23603), .Z(n23703) );
  XOR U23942 ( .A(n23702), .B(n23703), .Z(n23712) );
  NAND U23943 ( .A(n23597), .B(n23596), .Z(n23713) );
  IV U23944 ( .A(n23713), .Z(n23704) );
  XOR U23945 ( .A(n23712), .B(n23704), .Z(n23598) );
  XNOR U23946 ( .A(n23599), .B(n23598), .Z(c[109]) );
  NANDN U23947 ( .A(n23601), .B(n23600), .Z(n23605) );
  NANDN U23948 ( .A(n23603), .B(n23602), .Z(n23604) );
  AND U23949 ( .A(n23605), .B(n23604), .Z(n23813) );
  NANDN U23950 ( .A(n23607), .B(n23606), .Z(n23611) );
  NANDN U23951 ( .A(n23609), .B(n23608), .Z(n23610) );
  AND U23952 ( .A(n23611), .B(n23610), .Z(n23718) );
  AND U23953 ( .A(a[63]), .B(b[47]), .Z(n23717) );
  XNOR U23954 ( .A(n23718), .B(n23717), .Z(n23719) );
  NANDN U23955 ( .A(n23613), .B(n23612), .Z(n23617) );
  NANDN U23956 ( .A(n23615), .B(n23614), .Z(n23616) );
  AND U23957 ( .A(n23617), .B(n23616), .Z(n23726) );
  NANDN U23958 ( .A(n23619), .B(n23618), .Z(n23623) );
  NANDN U23959 ( .A(n23621), .B(n23620), .Z(n23622) );
  AND U23960 ( .A(n23623), .B(n23622), .Z(n23808) );
  AND U23961 ( .A(a[61]), .B(b[49]), .Z(n23807) );
  XNOR U23962 ( .A(n23808), .B(n23807), .Z(n23809) );
  NANDN U23963 ( .A(n23625), .B(n23624), .Z(n23629) );
  OR U23964 ( .A(n23627), .B(n23626), .Z(n23628) );
  AND U23965 ( .A(n23629), .B(n23628), .Z(n23731) );
  NANDN U23966 ( .A(n23631), .B(n23630), .Z(n23635) );
  NAND U23967 ( .A(n23633), .B(n23632), .Z(n23634) );
  AND U23968 ( .A(n23635), .B(n23634), .Z(n23802) );
  AND U23969 ( .A(a[59]), .B(b[51]), .Z(n23801) );
  XNOR U23970 ( .A(n23802), .B(n23801), .Z(n23803) );
  NANDN U23971 ( .A(n23637), .B(n23636), .Z(n23641) );
  NANDN U23972 ( .A(n23639), .B(n23638), .Z(n23640) );
  AND U23973 ( .A(n23641), .B(n23640), .Z(n23738) );
  NANDN U23974 ( .A(n23643), .B(n23642), .Z(n23647) );
  NANDN U23975 ( .A(n23645), .B(n23644), .Z(n23646) );
  AND U23976 ( .A(n23647), .B(n23646), .Z(n23796) );
  AND U23977 ( .A(a[57]), .B(b[53]), .Z(n23795) );
  XNOR U23978 ( .A(n23796), .B(n23795), .Z(n23797) );
  NANDN U23979 ( .A(n23649), .B(n23648), .Z(n23653) );
  OR U23980 ( .A(n23651), .B(n23650), .Z(n23652) );
  AND U23981 ( .A(n23653), .B(n23652), .Z(n23743) );
  NANDN U23982 ( .A(n23655), .B(n23654), .Z(n23659) );
  OR U23983 ( .A(n23657), .B(n23656), .Z(n23658) );
  AND U23984 ( .A(n23659), .B(n23658), .Z(n23790) );
  AND U23985 ( .A(a[55]), .B(b[55]), .Z(n23789) );
  XNOR U23986 ( .A(n23790), .B(n23789), .Z(n23791) );
  NANDN U23987 ( .A(n23661), .B(n23660), .Z(n23665) );
  NAND U23988 ( .A(n23663), .B(n23662), .Z(n23664) );
  AND U23989 ( .A(n23665), .B(n23664), .Z(n23749) );
  NANDN U23990 ( .A(n23667), .B(n23666), .Z(n23671) );
  OR U23991 ( .A(n23669), .B(n23668), .Z(n23670) );
  AND U23992 ( .A(n23671), .B(n23670), .Z(n23754) );
  AND U23993 ( .A(a[52]), .B(b[58]), .Z(n23753) );
  XNOR U23994 ( .A(n23754), .B(n23753), .Z(n23755) );
  NANDN U23995 ( .A(n23673), .B(n23672), .Z(n23677) );
  NANDN U23996 ( .A(n23675), .B(n23674), .Z(n23676) );
  AND U23997 ( .A(n23677), .B(n23676), .Z(n23766) );
  AND U23998 ( .A(a[50]), .B(b[60]), .Z(n23765) );
  XNOR U23999 ( .A(n23766), .B(n23765), .Z(n23767) );
  NANDN U24000 ( .A(n23679), .B(n23678), .Z(n23683) );
  NANDN U24001 ( .A(n23681), .B(n23680), .Z(n23682) );
  AND U24002 ( .A(n23683), .B(n23682), .Z(n23778) );
  AND U24003 ( .A(b[62]), .B(a[48]), .Z(n23777) );
  XNOR U24004 ( .A(n23778), .B(n23777), .Z(n23779) );
  NAND U24005 ( .A(b[63]), .B(a[47]), .Z(n23780) );
  XNOR U24006 ( .A(n23779), .B(n23780), .Z(n23773) );
  NANDN U24007 ( .A(n23685), .B(n23684), .Z(n23689) );
  NANDN U24008 ( .A(n23687), .B(n23686), .Z(n23688) );
  AND U24009 ( .A(n23689), .B(n23688), .Z(n23772) );
  AND U24010 ( .A(a[49]), .B(b[61]), .Z(n23771) );
  XOR U24011 ( .A(n23772), .B(n23771), .Z(n23774) );
  XOR U24012 ( .A(n23773), .B(n23774), .Z(n23768) );
  XNOR U24013 ( .A(n23767), .B(n23768), .Z(n23761) );
  NANDN U24014 ( .A(n23691), .B(n23690), .Z(n23695) );
  NANDN U24015 ( .A(n23693), .B(n23692), .Z(n23694) );
  AND U24016 ( .A(n23695), .B(n23694), .Z(n23760) );
  AND U24017 ( .A(a[51]), .B(b[59]), .Z(n23759) );
  XOR U24018 ( .A(n23760), .B(n23759), .Z(n23762) );
  XOR U24019 ( .A(n23761), .B(n23762), .Z(n23756) );
  XNOR U24020 ( .A(n23755), .B(n23756), .Z(n23783) );
  NANDN U24021 ( .A(n23697), .B(n23696), .Z(n23701) );
  NANDN U24022 ( .A(n23699), .B(n23698), .Z(n23700) );
  NAND U24023 ( .A(n23701), .B(n23700), .Z(n23784) );
  XNOR U24024 ( .A(n23783), .B(n23784), .Z(n23785) );
  NAND U24025 ( .A(a[53]), .B(b[57]), .Z(n23786) );
  XNOR U24026 ( .A(n23785), .B(n23786), .Z(n23747) );
  NAND U24027 ( .A(a[54]), .B(b[56]), .Z(n23748) );
  XOR U24028 ( .A(n23747), .B(n23748), .Z(n23750) );
  XOR U24029 ( .A(n23749), .B(n23750), .Z(n23792) );
  XNOR U24030 ( .A(n23791), .B(n23792), .Z(n23741) );
  NAND U24031 ( .A(a[56]), .B(b[54]), .Z(n23742) );
  XOR U24032 ( .A(n23741), .B(n23742), .Z(n23744) );
  XOR U24033 ( .A(n23743), .B(n23744), .Z(n23798) );
  XNOR U24034 ( .A(n23797), .B(n23798), .Z(n23735) );
  NAND U24035 ( .A(a[58]), .B(b[52]), .Z(n23736) );
  XNOR U24036 ( .A(n23735), .B(n23736), .Z(n23737) );
  XOR U24037 ( .A(n23738), .B(n23737), .Z(n23804) );
  XNOR U24038 ( .A(n23803), .B(n23804), .Z(n23729) );
  NAND U24039 ( .A(a[60]), .B(b[50]), .Z(n23730) );
  XOR U24040 ( .A(n23729), .B(n23730), .Z(n23732) );
  XOR U24041 ( .A(n23731), .B(n23732), .Z(n23810) );
  XNOR U24042 ( .A(n23809), .B(n23810), .Z(n23723) );
  NAND U24043 ( .A(a[62]), .B(b[48]), .Z(n23724) );
  XNOR U24044 ( .A(n23723), .B(n23724), .Z(n23725) );
  XOR U24045 ( .A(n23726), .B(n23725), .Z(n23720) );
  XNOR U24046 ( .A(n23719), .B(n23720), .Z(n23814) );
  XNOR U24047 ( .A(n23813), .B(n23814), .Z(n23816) );
  ANDN U24048 ( .B(n23703), .A(n23702), .Z(n23815) );
  XOR U24049 ( .A(n23816), .B(n23815), .Z(n23818) );
  XOR U24050 ( .A(n23818), .B(n23817), .Z(c[110]) );
  NANDN U24051 ( .A(n23718), .B(n23717), .Z(n23722) );
  NANDN U24052 ( .A(n23720), .B(n23719), .Z(n23721) );
  AND U24053 ( .A(n23722), .B(n23721), .Z(n23909) );
  NANDN U24054 ( .A(n23724), .B(n23723), .Z(n23728) );
  NANDN U24055 ( .A(n23726), .B(n23725), .Z(n23727) );
  AND U24056 ( .A(n23728), .B(n23727), .Z(n23820) );
  AND U24057 ( .A(a[63]), .B(b[48]), .Z(n23819) );
  XNOR U24058 ( .A(n23820), .B(n23819), .Z(n23821) );
  NANDN U24059 ( .A(n23730), .B(n23729), .Z(n23734) );
  NANDN U24060 ( .A(n23732), .B(n23731), .Z(n23733) );
  AND U24061 ( .A(n23734), .B(n23733), .Z(n23832) );
  AND U24062 ( .A(a[61]), .B(b[50]), .Z(n23831) );
  XNOR U24063 ( .A(n23832), .B(n23831), .Z(n23833) );
  NANDN U24064 ( .A(n23736), .B(n23735), .Z(n23740) );
  NANDN U24065 ( .A(n23738), .B(n23737), .Z(n23739) );
  AND U24066 ( .A(n23740), .B(n23739), .Z(n23844) );
  AND U24067 ( .A(a[59]), .B(b[52]), .Z(n23843) );
  XNOR U24068 ( .A(n23844), .B(n23843), .Z(n23845) );
  NANDN U24069 ( .A(n23742), .B(n23741), .Z(n23746) );
  NANDN U24070 ( .A(n23744), .B(n23743), .Z(n23745) );
  AND U24071 ( .A(n23746), .B(n23745), .Z(n23856) );
  AND U24072 ( .A(a[57]), .B(b[54]), .Z(n23855) );
  XNOR U24073 ( .A(n23856), .B(n23855), .Z(n23857) );
  AND U24074 ( .A(a[55]), .B(b[56]), .Z(n23868) );
  NANDN U24075 ( .A(n23748), .B(n23747), .Z(n23752) );
  NANDN U24076 ( .A(n23750), .B(n23749), .Z(n23751) );
  AND U24077 ( .A(n23752), .B(n23751), .Z(n23867) );
  XNOR U24078 ( .A(n23868), .B(n23867), .Z(n23870) );
  AND U24079 ( .A(a[54]), .B(b[57]), .Z(n23906) );
  NANDN U24080 ( .A(n23754), .B(n23753), .Z(n23758) );
  NANDN U24081 ( .A(n23756), .B(n23755), .Z(n23757) );
  AND U24082 ( .A(n23758), .B(n23757), .Z(n23875) );
  NANDN U24083 ( .A(n23760), .B(n23759), .Z(n23764) );
  NANDN U24084 ( .A(n23762), .B(n23761), .Z(n23763) );
  AND U24085 ( .A(n23764), .B(n23763), .Z(n23898) );
  AND U24086 ( .A(a[52]), .B(b[59]), .Z(n23897) );
  XNOR U24087 ( .A(n23898), .B(n23897), .Z(n23899) );
  NANDN U24088 ( .A(n23766), .B(n23765), .Z(n23770) );
  NANDN U24089 ( .A(n23768), .B(n23767), .Z(n23769) );
  AND U24090 ( .A(n23770), .B(n23769), .Z(n23882) );
  NANDN U24091 ( .A(n23772), .B(n23771), .Z(n23776) );
  NANDN U24092 ( .A(n23774), .B(n23773), .Z(n23775) );
  AND U24093 ( .A(n23776), .B(n23775), .Z(n23892) );
  AND U24094 ( .A(a[50]), .B(b[61]), .Z(n23891) );
  XNOR U24095 ( .A(n23892), .B(n23891), .Z(n23893) );
  NANDN U24096 ( .A(n23778), .B(n23777), .Z(n23782) );
  NANDN U24097 ( .A(n23780), .B(n23779), .Z(n23781) );
  AND U24098 ( .A(n23782), .B(n23781), .Z(n23886) );
  AND U24099 ( .A(b[62]), .B(a[49]), .Z(n23885) );
  XNOR U24100 ( .A(n23886), .B(n23885), .Z(n23887) );
  NAND U24101 ( .A(b[63]), .B(a[48]), .Z(n23888) );
  XOR U24102 ( .A(n23887), .B(n23888), .Z(n23894) );
  XNOR U24103 ( .A(n23893), .B(n23894), .Z(n23879) );
  NAND U24104 ( .A(a[51]), .B(b[60]), .Z(n23880) );
  XNOR U24105 ( .A(n23879), .B(n23880), .Z(n23881) );
  XOR U24106 ( .A(n23882), .B(n23881), .Z(n23900) );
  XNOR U24107 ( .A(n23899), .B(n23900), .Z(n23873) );
  NAND U24108 ( .A(a[53]), .B(b[58]), .Z(n23874) );
  XOR U24109 ( .A(n23873), .B(n23874), .Z(n23876) );
  XOR U24110 ( .A(n23875), .B(n23876), .Z(n23904) );
  NANDN U24111 ( .A(n23784), .B(n23783), .Z(n23788) );
  NANDN U24112 ( .A(n23786), .B(n23785), .Z(n23787) );
  AND U24113 ( .A(n23788), .B(n23787), .Z(n23903) );
  XNOR U24114 ( .A(n23904), .B(n23903), .Z(n23905) );
  XNOR U24115 ( .A(n23906), .B(n23905), .Z(n23869) );
  XOR U24116 ( .A(n23870), .B(n23869), .Z(n23864) );
  NANDN U24117 ( .A(n23790), .B(n23789), .Z(n23794) );
  NANDN U24118 ( .A(n23792), .B(n23791), .Z(n23793) );
  AND U24119 ( .A(n23794), .B(n23793), .Z(n23862) );
  AND U24120 ( .A(a[56]), .B(b[55]), .Z(n23861) );
  XNOR U24121 ( .A(n23862), .B(n23861), .Z(n23863) );
  XOR U24122 ( .A(n23864), .B(n23863), .Z(n23858) );
  XNOR U24123 ( .A(n23857), .B(n23858), .Z(n23851) );
  NANDN U24124 ( .A(n23796), .B(n23795), .Z(n23800) );
  NANDN U24125 ( .A(n23798), .B(n23797), .Z(n23799) );
  AND U24126 ( .A(n23800), .B(n23799), .Z(n23850) );
  AND U24127 ( .A(a[58]), .B(b[53]), .Z(n23849) );
  XOR U24128 ( .A(n23850), .B(n23849), .Z(n23852) );
  XOR U24129 ( .A(n23851), .B(n23852), .Z(n23846) );
  XNOR U24130 ( .A(n23845), .B(n23846), .Z(n23839) );
  NANDN U24131 ( .A(n23802), .B(n23801), .Z(n23806) );
  NANDN U24132 ( .A(n23804), .B(n23803), .Z(n23805) );
  AND U24133 ( .A(n23806), .B(n23805), .Z(n23838) );
  AND U24134 ( .A(a[60]), .B(b[51]), .Z(n23837) );
  XOR U24135 ( .A(n23838), .B(n23837), .Z(n23840) );
  XOR U24136 ( .A(n23839), .B(n23840), .Z(n23834) );
  XNOR U24137 ( .A(n23833), .B(n23834), .Z(n23827) );
  NANDN U24138 ( .A(n23808), .B(n23807), .Z(n23812) );
  NANDN U24139 ( .A(n23810), .B(n23809), .Z(n23811) );
  AND U24140 ( .A(n23812), .B(n23811), .Z(n23826) );
  AND U24141 ( .A(a[62]), .B(b[49]), .Z(n23825) );
  XOR U24142 ( .A(n23826), .B(n23825), .Z(n23828) );
  XOR U24143 ( .A(n23827), .B(n23828), .Z(n23822) );
  XNOR U24144 ( .A(n23821), .B(n23822), .Z(n23910) );
  XNOR U24145 ( .A(n23909), .B(n23910), .Z(n23912) );
  ANDN U24146 ( .B(n23814), .A(n23813), .Z(n23911) );
  XOR U24147 ( .A(n23912), .B(n23911), .Z(n23914) );
  XOR U24148 ( .A(n23914), .B(n23913), .Z(c[111]) );
  NANDN U24149 ( .A(n23820), .B(n23819), .Z(n23824) );
  NANDN U24150 ( .A(n23822), .B(n23821), .Z(n23823) );
  AND U24151 ( .A(n23824), .B(n23823), .Z(n23919) );
  NANDN U24152 ( .A(n23826), .B(n23825), .Z(n23830) );
  NANDN U24153 ( .A(n23828), .B(n23827), .Z(n23829) );
  AND U24154 ( .A(n23830), .B(n23829), .Z(n24000) );
  AND U24155 ( .A(a[63]), .B(b[49]), .Z(n23999) );
  XNOR U24156 ( .A(n24000), .B(n23999), .Z(n24001) );
  NANDN U24157 ( .A(n23832), .B(n23831), .Z(n23836) );
  NANDN U24158 ( .A(n23834), .B(n23833), .Z(n23835) );
  AND U24159 ( .A(n23836), .B(n23835), .Z(n23996) );
  NANDN U24160 ( .A(n23838), .B(n23837), .Z(n23842) );
  NANDN U24161 ( .A(n23840), .B(n23839), .Z(n23841) );
  AND U24162 ( .A(n23842), .B(n23841), .Z(n23988) );
  AND U24163 ( .A(a[61]), .B(b[51]), .Z(n23987) );
  XNOR U24164 ( .A(n23988), .B(n23987), .Z(n23989) );
  NANDN U24165 ( .A(n23844), .B(n23843), .Z(n23848) );
  NANDN U24166 ( .A(n23846), .B(n23845), .Z(n23847) );
  AND U24167 ( .A(n23848), .B(n23847), .Z(n23924) );
  NANDN U24168 ( .A(n23850), .B(n23849), .Z(n23854) );
  NANDN U24169 ( .A(n23852), .B(n23851), .Z(n23853) );
  AND U24170 ( .A(n23854), .B(n23853), .Z(n23982) );
  AND U24171 ( .A(a[59]), .B(b[53]), .Z(n23981) );
  XNOR U24172 ( .A(n23982), .B(n23981), .Z(n23983) );
  NANDN U24173 ( .A(n23856), .B(n23855), .Z(n23860) );
  NANDN U24174 ( .A(n23858), .B(n23857), .Z(n23859) );
  AND U24175 ( .A(n23860), .B(n23859), .Z(n23978) );
  NANDN U24176 ( .A(n23862), .B(n23861), .Z(n23866) );
  NANDN U24177 ( .A(n23864), .B(n23863), .Z(n23865) );
  AND U24178 ( .A(n23866), .B(n23865), .Z(n23970) );
  AND U24179 ( .A(a[57]), .B(b[55]), .Z(n23969) );
  XNOR U24180 ( .A(n23970), .B(n23969), .Z(n23971) );
  NANDN U24181 ( .A(n23868), .B(n23867), .Z(n23872) );
  NAND U24182 ( .A(n23870), .B(n23869), .Z(n23871) );
  AND U24183 ( .A(n23872), .B(n23871), .Z(n23929) );
  NANDN U24184 ( .A(n23874), .B(n23873), .Z(n23878) );
  OR U24185 ( .A(n23876), .B(n23875), .Z(n23877) );
  AND U24186 ( .A(n23878), .B(n23877), .Z(n23934) );
  AND U24187 ( .A(a[54]), .B(b[58]), .Z(n23933) );
  XNOR U24188 ( .A(n23934), .B(n23933), .Z(n23935) );
  NANDN U24189 ( .A(n23880), .B(n23879), .Z(n23884) );
  NANDN U24190 ( .A(n23882), .B(n23881), .Z(n23883) );
  AND U24191 ( .A(n23884), .B(n23883), .Z(n23946) );
  AND U24192 ( .A(a[52]), .B(b[60]), .Z(n23945) );
  XNOR U24193 ( .A(n23946), .B(n23945), .Z(n23947) );
  NANDN U24194 ( .A(n23886), .B(n23885), .Z(n23890) );
  NANDN U24195 ( .A(n23888), .B(n23887), .Z(n23889) );
  AND U24196 ( .A(n23890), .B(n23889), .Z(n23952) );
  AND U24197 ( .A(b[62]), .B(a[50]), .Z(n23951) );
  XNOR U24198 ( .A(n23952), .B(n23951), .Z(n23953) );
  NAND U24199 ( .A(b[63]), .B(a[49]), .Z(n23954) );
  XNOR U24200 ( .A(n23953), .B(n23954), .Z(n23959) );
  NANDN U24201 ( .A(n23892), .B(n23891), .Z(n23896) );
  NANDN U24202 ( .A(n23894), .B(n23893), .Z(n23895) );
  AND U24203 ( .A(n23896), .B(n23895), .Z(n23958) );
  AND U24204 ( .A(a[51]), .B(b[61]), .Z(n23957) );
  XOR U24205 ( .A(n23958), .B(n23957), .Z(n23960) );
  XOR U24206 ( .A(n23959), .B(n23960), .Z(n23948) );
  XNOR U24207 ( .A(n23947), .B(n23948), .Z(n23941) );
  NANDN U24208 ( .A(n23898), .B(n23897), .Z(n23902) );
  NANDN U24209 ( .A(n23900), .B(n23899), .Z(n23901) );
  AND U24210 ( .A(n23902), .B(n23901), .Z(n23940) );
  AND U24211 ( .A(a[53]), .B(b[59]), .Z(n23939) );
  XOR U24212 ( .A(n23940), .B(n23939), .Z(n23942) );
  XOR U24213 ( .A(n23941), .B(n23942), .Z(n23936) );
  XNOR U24214 ( .A(n23935), .B(n23936), .Z(n23963) );
  NANDN U24215 ( .A(n23904), .B(n23903), .Z(n23908) );
  NANDN U24216 ( .A(n23906), .B(n23905), .Z(n23907) );
  NAND U24217 ( .A(n23908), .B(n23907), .Z(n23964) );
  XNOR U24218 ( .A(n23963), .B(n23964), .Z(n23965) );
  NAND U24219 ( .A(a[55]), .B(b[57]), .Z(n23966) );
  XNOR U24220 ( .A(n23965), .B(n23966), .Z(n23927) );
  NAND U24221 ( .A(a[56]), .B(b[56]), .Z(n23928) );
  XOR U24222 ( .A(n23927), .B(n23928), .Z(n23930) );
  XOR U24223 ( .A(n23929), .B(n23930), .Z(n23972) );
  XNOR U24224 ( .A(n23971), .B(n23972), .Z(n23975) );
  NAND U24225 ( .A(a[58]), .B(b[54]), .Z(n23976) );
  XNOR U24226 ( .A(n23975), .B(n23976), .Z(n23977) );
  XOR U24227 ( .A(n23978), .B(n23977), .Z(n23984) );
  XNOR U24228 ( .A(n23983), .B(n23984), .Z(n23921) );
  NAND U24229 ( .A(a[60]), .B(b[52]), .Z(n23922) );
  XNOR U24230 ( .A(n23921), .B(n23922), .Z(n23923) );
  XOR U24231 ( .A(n23924), .B(n23923), .Z(n23990) );
  XNOR U24232 ( .A(n23989), .B(n23990), .Z(n23993) );
  NAND U24233 ( .A(a[62]), .B(b[50]), .Z(n23994) );
  XNOR U24234 ( .A(n23993), .B(n23994), .Z(n23995) );
  XOR U24235 ( .A(n23996), .B(n23995), .Z(n24002) );
  XNOR U24236 ( .A(n24001), .B(n24002), .Z(n23920) );
  XNOR U24237 ( .A(n23919), .B(n23920), .Z(n23916) );
  ANDN U24238 ( .B(n23910), .A(n23909), .Z(n23915) );
  XOR U24239 ( .A(n23916), .B(n23915), .Z(n23918) );
  XOR U24240 ( .A(n23918), .B(n23917), .Z(c[112]) );
  ANDN U24241 ( .B(n23920), .A(n23919), .Z(n24086) );
  NANDN U24242 ( .A(n23922), .B(n23921), .Z(n23926) );
  NANDN U24243 ( .A(n23924), .B(n23923), .Z(n23925) );
  AND U24244 ( .A(n23926), .B(n23925), .Z(n24014) );
  AND U24245 ( .A(a[61]), .B(b[52]), .Z(n24013) );
  XNOR U24246 ( .A(n24014), .B(n24013), .Z(n24015) );
  AND U24247 ( .A(a[57]), .B(b[56]), .Z(n24038) );
  NANDN U24248 ( .A(n23928), .B(n23927), .Z(n23932) );
  NANDN U24249 ( .A(n23930), .B(n23929), .Z(n23931) );
  AND U24250 ( .A(n23932), .B(n23931), .Z(n24037) );
  XNOR U24251 ( .A(n24038), .B(n24037), .Z(n24040) );
  AND U24252 ( .A(a[56]), .B(b[57]), .Z(n24076) );
  NANDN U24253 ( .A(n23934), .B(n23933), .Z(n23938) );
  NANDN U24254 ( .A(n23936), .B(n23935), .Z(n23937) );
  AND U24255 ( .A(n23938), .B(n23937), .Z(n24045) );
  NANDN U24256 ( .A(n23940), .B(n23939), .Z(n23944) );
  NANDN U24257 ( .A(n23942), .B(n23941), .Z(n23943) );
  AND U24258 ( .A(n23944), .B(n23943), .Z(n24068) );
  AND U24259 ( .A(a[54]), .B(b[59]), .Z(n24067) );
  XNOR U24260 ( .A(n24068), .B(n24067), .Z(n24069) );
  NANDN U24261 ( .A(n23946), .B(n23945), .Z(n23950) );
  NANDN U24262 ( .A(n23948), .B(n23947), .Z(n23949) );
  AND U24263 ( .A(n23950), .B(n23949), .Z(n24052) );
  NANDN U24264 ( .A(n23952), .B(n23951), .Z(n23956) );
  NANDN U24265 ( .A(n23954), .B(n23953), .Z(n23955) );
  AND U24266 ( .A(n23956), .B(n23955), .Z(n24058) );
  AND U24267 ( .A(b[62]), .B(a[51]), .Z(n24055) );
  NAND U24268 ( .A(b[63]), .B(a[50]), .Z(n24056) );
  XNOR U24269 ( .A(n24055), .B(n24056), .Z(n24057) );
  XNOR U24270 ( .A(n24058), .B(n24057), .Z(n24063) );
  NANDN U24271 ( .A(n23958), .B(n23957), .Z(n23962) );
  NANDN U24272 ( .A(n23960), .B(n23959), .Z(n23961) );
  AND U24273 ( .A(n23962), .B(n23961), .Z(n24062) );
  AND U24274 ( .A(a[52]), .B(b[61]), .Z(n24061) );
  XOR U24275 ( .A(n24062), .B(n24061), .Z(n24064) );
  XNOR U24276 ( .A(n24063), .B(n24064), .Z(n24049) );
  NAND U24277 ( .A(a[53]), .B(b[60]), .Z(n24050) );
  XNOR U24278 ( .A(n24049), .B(n24050), .Z(n24051) );
  XOR U24279 ( .A(n24052), .B(n24051), .Z(n24070) );
  XNOR U24280 ( .A(n24069), .B(n24070), .Z(n24043) );
  NAND U24281 ( .A(a[55]), .B(b[58]), .Z(n24044) );
  XOR U24282 ( .A(n24043), .B(n24044), .Z(n24046) );
  XOR U24283 ( .A(n24045), .B(n24046), .Z(n24074) );
  NANDN U24284 ( .A(n23964), .B(n23963), .Z(n23968) );
  NANDN U24285 ( .A(n23966), .B(n23965), .Z(n23967) );
  AND U24286 ( .A(n23968), .B(n23967), .Z(n24073) );
  XNOR U24287 ( .A(n24074), .B(n24073), .Z(n24075) );
  XNOR U24288 ( .A(n24076), .B(n24075), .Z(n24039) );
  XOR U24289 ( .A(n24040), .B(n24039), .Z(n24033) );
  NANDN U24290 ( .A(n23970), .B(n23969), .Z(n23974) );
  NANDN U24291 ( .A(n23972), .B(n23971), .Z(n23973) );
  AND U24292 ( .A(n23974), .B(n23973), .Z(n24032) );
  AND U24293 ( .A(a[58]), .B(b[55]), .Z(n24031) );
  XOR U24294 ( .A(n24032), .B(n24031), .Z(n24034) );
  XOR U24295 ( .A(n24033), .B(n24034), .Z(n24027) );
  AND U24296 ( .A(a[59]), .B(b[54]), .Z(n24026) );
  NANDN U24297 ( .A(n23976), .B(n23975), .Z(n23980) );
  NANDN U24298 ( .A(n23978), .B(n23977), .Z(n23979) );
  AND U24299 ( .A(n23980), .B(n23979), .Z(n24025) );
  XOR U24300 ( .A(n24026), .B(n24025), .Z(n24028) );
  XOR U24301 ( .A(n24027), .B(n24028), .Z(n24022) );
  NANDN U24302 ( .A(n23982), .B(n23981), .Z(n23986) );
  NANDN U24303 ( .A(n23984), .B(n23983), .Z(n23985) );
  AND U24304 ( .A(n23986), .B(n23985), .Z(n24020) );
  AND U24305 ( .A(a[60]), .B(b[53]), .Z(n24019) );
  XNOR U24306 ( .A(n24020), .B(n24019), .Z(n24021) );
  XOR U24307 ( .A(n24022), .B(n24021), .Z(n24016) );
  XNOR U24308 ( .A(n24015), .B(n24016), .Z(n24010) );
  NANDN U24309 ( .A(n23988), .B(n23987), .Z(n23992) );
  NANDN U24310 ( .A(n23990), .B(n23989), .Z(n23991) );
  AND U24311 ( .A(n23992), .B(n23991), .Z(n24008) );
  AND U24312 ( .A(a[62]), .B(b[51]), .Z(n24007) );
  XNOR U24313 ( .A(n24008), .B(n24007), .Z(n24009) );
  XOR U24314 ( .A(n24010), .B(n24009), .Z(n24081) );
  AND U24315 ( .A(a[63]), .B(b[50]), .Z(n24080) );
  NANDN U24316 ( .A(n23994), .B(n23993), .Z(n23998) );
  NANDN U24317 ( .A(n23996), .B(n23995), .Z(n23997) );
  AND U24318 ( .A(n23998), .B(n23997), .Z(n24079) );
  XOR U24319 ( .A(n24080), .B(n24079), .Z(n24082) );
  XOR U24320 ( .A(n24081), .B(n24082), .Z(n24006) );
  NANDN U24321 ( .A(n24000), .B(n23999), .Z(n24004) );
  NANDN U24322 ( .A(n24002), .B(n24001), .Z(n24003) );
  AND U24323 ( .A(n24004), .B(n24003), .Z(n24005) );
  XNOR U24324 ( .A(n24006), .B(n24005), .Z(n24085) );
  XNOR U24325 ( .A(n24086), .B(n24085), .Z(n24087) );
  XNOR U24326 ( .A(n24088), .B(n24087), .Z(c[113]) );
  NOR U24327 ( .A(n24006), .B(n24005), .Z(n24166) );
  NANDN U24328 ( .A(n24008), .B(n24007), .Z(n24012) );
  NAND U24329 ( .A(n24010), .B(n24009), .Z(n24011) );
  AND U24330 ( .A(n24012), .B(n24011), .Z(n24092) );
  AND U24331 ( .A(a[63]), .B(b[51]), .Z(n24091) );
  XNOR U24332 ( .A(n24092), .B(n24091), .Z(n24093) );
  NANDN U24333 ( .A(n24014), .B(n24013), .Z(n24018) );
  NANDN U24334 ( .A(n24016), .B(n24015), .Z(n24017) );
  AND U24335 ( .A(n24018), .B(n24017), .Z(n24100) );
  NANDN U24336 ( .A(n24020), .B(n24019), .Z(n24024) );
  NANDN U24337 ( .A(n24022), .B(n24021), .Z(n24023) );
  AND U24338 ( .A(n24024), .B(n24023), .Z(n24158) );
  AND U24339 ( .A(a[61]), .B(b[53]), .Z(n24157) );
  XNOR U24340 ( .A(n24158), .B(n24157), .Z(n24159) );
  NANDN U24341 ( .A(n24026), .B(n24025), .Z(n24030) );
  OR U24342 ( .A(n24028), .B(n24027), .Z(n24029) );
  AND U24343 ( .A(n24030), .B(n24029), .Z(n24105) );
  NANDN U24344 ( .A(n24032), .B(n24031), .Z(n24036) );
  OR U24345 ( .A(n24034), .B(n24033), .Z(n24035) );
  AND U24346 ( .A(n24036), .B(n24035), .Z(n24152) );
  AND U24347 ( .A(a[59]), .B(b[55]), .Z(n24151) );
  XNOR U24348 ( .A(n24152), .B(n24151), .Z(n24153) );
  NANDN U24349 ( .A(n24038), .B(n24037), .Z(n24042) );
  NAND U24350 ( .A(n24040), .B(n24039), .Z(n24041) );
  AND U24351 ( .A(n24042), .B(n24041), .Z(n24111) );
  NANDN U24352 ( .A(n24044), .B(n24043), .Z(n24048) );
  OR U24353 ( .A(n24046), .B(n24045), .Z(n24047) );
  AND U24354 ( .A(n24048), .B(n24047), .Z(n24116) );
  AND U24355 ( .A(a[56]), .B(b[58]), .Z(n24115) );
  XNOR U24356 ( .A(n24116), .B(n24115), .Z(n24117) );
  NANDN U24357 ( .A(n24050), .B(n24049), .Z(n24054) );
  NANDN U24358 ( .A(n24052), .B(n24051), .Z(n24053) );
  AND U24359 ( .A(n24054), .B(n24053), .Z(n24128) );
  AND U24360 ( .A(a[54]), .B(b[60]), .Z(n24127) );
  XNOR U24361 ( .A(n24128), .B(n24127), .Z(n24129) );
  NANDN U24362 ( .A(n24056), .B(n24055), .Z(n24060) );
  NANDN U24363 ( .A(n24058), .B(n24057), .Z(n24059) );
  AND U24364 ( .A(n24060), .B(n24059), .Z(n24134) );
  AND U24365 ( .A(b[62]), .B(a[52]), .Z(n24133) );
  XNOR U24366 ( .A(n24134), .B(n24133), .Z(n24135) );
  NAND U24367 ( .A(b[63]), .B(a[51]), .Z(n24136) );
  XNOR U24368 ( .A(n24135), .B(n24136), .Z(n24141) );
  NANDN U24369 ( .A(n24062), .B(n24061), .Z(n24066) );
  NANDN U24370 ( .A(n24064), .B(n24063), .Z(n24065) );
  AND U24371 ( .A(n24066), .B(n24065), .Z(n24140) );
  AND U24372 ( .A(a[53]), .B(b[61]), .Z(n24139) );
  XOR U24373 ( .A(n24140), .B(n24139), .Z(n24142) );
  XOR U24374 ( .A(n24141), .B(n24142), .Z(n24130) );
  XNOR U24375 ( .A(n24129), .B(n24130), .Z(n24123) );
  NANDN U24376 ( .A(n24068), .B(n24067), .Z(n24072) );
  NANDN U24377 ( .A(n24070), .B(n24069), .Z(n24071) );
  AND U24378 ( .A(n24072), .B(n24071), .Z(n24122) );
  AND U24379 ( .A(a[55]), .B(b[59]), .Z(n24121) );
  XOR U24380 ( .A(n24122), .B(n24121), .Z(n24124) );
  XOR U24381 ( .A(n24123), .B(n24124), .Z(n24118) );
  XNOR U24382 ( .A(n24117), .B(n24118), .Z(n24145) );
  NANDN U24383 ( .A(n24074), .B(n24073), .Z(n24078) );
  NANDN U24384 ( .A(n24076), .B(n24075), .Z(n24077) );
  NAND U24385 ( .A(n24078), .B(n24077), .Z(n24146) );
  XNOR U24386 ( .A(n24145), .B(n24146), .Z(n24147) );
  NAND U24387 ( .A(a[57]), .B(b[57]), .Z(n24148) );
  XNOR U24388 ( .A(n24147), .B(n24148), .Z(n24109) );
  NAND U24389 ( .A(a[58]), .B(b[56]), .Z(n24110) );
  XOR U24390 ( .A(n24109), .B(n24110), .Z(n24112) );
  XOR U24391 ( .A(n24111), .B(n24112), .Z(n24154) );
  XNOR U24392 ( .A(n24153), .B(n24154), .Z(n24103) );
  NAND U24393 ( .A(a[60]), .B(b[54]), .Z(n24104) );
  XOR U24394 ( .A(n24103), .B(n24104), .Z(n24106) );
  XOR U24395 ( .A(n24105), .B(n24106), .Z(n24160) );
  XNOR U24396 ( .A(n24159), .B(n24160), .Z(n24097) );
  NAND U24397 ( .A(a[62]), .B(b[52]), .Z(n24098) );
  XNOR U24398 ( .A(n24097), .B(n24098), .Z(n24099) );
  XOR U24399 ( .A(n24100), .B(n24099), .Z(n24094) );
  XNOR U24400 ( .A(n24093), .B(n24094), .Z(n24164) );
  NANDN U24401 ( .A(n24080), .B(n24079), .Z(n24084) );
  OR U24402 ( .A(n24082), .B(n24081), .Z(n24083) );
  AND U24403 ( .A(n24084), .B(n24083), .Z(n24163) );
  XNOR U24404 ( .A(n24164), .B(n24163), .Z(n24165) );
  XNOR U24405 ( .A(n24166), .B(n24165), .Z(n24168) );
  NANDN U24406 ( .A(n24086), .B(n24085), .Z(n24090) );
  NAND U24407 ( .A(n24088), .B(n24087), .Z(n24089) );
  NAND U24408 ( .A(n24090), .B(n24089), .Z(n24167) );
  XNOR U24409 ( .A(n24168), .B(n24167), .Z(c[114]) );
  NANDN U24410 ( .A(n24092), .B(n24091), .Z(n24096) );
  NANDN U24411 ( .A(n24094), .B(n24093), .Z(n24095) );
  AND U24412 ( .A(n24096), .B(n24095), .Z(n24177) );
  NANDN U24413 ( .A(n24098), .B(n24097), .Z(n24102) );
  NANDN U24414 ( .A(n24100), .B(n24099), .Z(n24101) );
  AND U24415 ( .A(n24102), .B(n24101), .Z(n24180) );
  AND U24416 ( .A(a[63]), .B(b[52]), .Z(n24179) );
  XNOR U24417 ( .A(n24180), .B(n24179), .Z(n24181) );
  NANDN U24418 ( .A(n24104), .B(n24103), .Z(n24108) );
  NANDN U24419 ( .A(n24106), .B(n24105), .Z(n24107) );
  AND U24420 ( .A(n24108), .B(n24107), .Z(n24192) );
  AND U24421 ( .A(a[61]), .B(b[54]), .Z(n24191) );
  XNOR U24422 ( .A(n24192), .B(n24191), .Z(n24193) );
  AND U24423 ( .A(a[59]), .B(b[56]), .Z(n24204) );
  NANDN U24424 ( .A(n24110), .B(n24109), .Z(n24114) );
  NANDN U24425 ( .A(n24112), .B(n24111), .Z(n24113) );
  AND U24426 ( .A(n24114), .B(n24113), .Z(n24203) );
  XNOR U24427 ( .A(n24204), .B(n24203), .Z(n24206) );
  AND U24428 ( .A(a[58]), .B(b[57]), .Z(n24242) );
  NANDN U24429 ( .A(n24116), .B(n24115), .Z(n24120) );
  NANDN U24430 ( .A(n24118), .B(n24117), .Z(n24119) );
  AND U24431 ( .A(n24120), .B(n24119), .Z(n24211) );
  NANDN U24432 ( .A(n24122), .B(n24121), .Z(n24126) );
  NANDN U24433 ( .A(n24124), .B(n24123), .Z(n24125) );
  AND U24434 ( .A(n24126), .B(n24125), .Z(n24234) );
  AND U24435 ( .A(a[56]), .B(b[59]), .Z(n24233) );
  XNOR U24436 ( .A(n24234), .B(n24233), .Z(n24235) );
  NANDN U24437 ( .A(n24128), .B(n24127), .Z(n24132) );
  NANDN U24438 ( .A(n24130), .B(n24129), .Z(n24131) );
  AND U24439 ( .A(n24132), .B(n24131), .Z(n24218) );
  NANDN U24440 ( .A(n24134), .B(n24133), .Z(n24138) );
  NANDN U24441 ( .A(n24136), .B(n24135), .Z(n24137) );
  AND U24442 ( .A(n24138), .B(n24137), .Z(n24222) );
  AND U24443 ( .A(b[62]), .B(a[53]), .Z(n24221) );
  XNOR U24444 ( .A(n24222), .B(n24221), .Z(n24223) );
  NAND U24445 ( .A(b[63]), .B(a[52]), .Z(n24224) );
  XNOR U24446 ( .A(n24223), .B(n24224), .Z(n24229) );
  NANDN U24447 ( .A(n24140), .B(n24139), .Z(n24144) );
  NANDN U24448 ( .A(n24142), .B(n24141), .Z(n24143) );
  AND U24449 ( .A(n24144), .B(n24143), .Z(n24228) );
  AND U24450 ( .A(a[54]), .B(b[61]), .Z(n24227) );
  XOR U24451 ( .A(n24228), .B(n24227), .Z(n24230) );
  XNOR U24452 ( .A(n24229), .B(n24230), .Z(n24215) );
  NAND U24453 ( .A(a[55]), .B(b[60]), .Z(n24216) );
  XNOR U24454 ( .A(n24215), .B(n24216), .Z(n24217) );
  XOR U24455 ( .A(n24218), .B(n24217), .Z(n24236) );
  XNOR U24456 ( .A(n24235), .B(n24236), .Z(n24209) );
  NAND U24457 ( .A(a[57]), .B(b[58]), .Z(n24210) );
  XOR U24458 ( .A(n24209), .B(n24210), .Z(n24212) );
  XOR U24459 ( .A(n24211), .B(n24212), .Z(n24240) );
  NANDN U24460 ( .A(n24146), .B(n24145), .Z(n24150) );
  NANDN U24461 ( .A(n24148), .B(n24147), .Z(n24149) );
  AND U24462 ( .A(n24150), .B(n24149), .Z(n24239) );
  XNOR U24463 ( .A(n24240), .B(n24239), .Z(n24241) );
  XNOR U24464 ( .A(n24242), .B(n24241), .Z(n24205) );
  XOR U24465 ( .A(n24206), .B(n24205), .Z(n24200) );
  NANDN U24466 ( .A(n24152), .B(n24151), .Z(n24156) );
  NANDN U24467 ( .A(n24154), .B(n24153), .Z(n24155) );
  AND U24468 ( .A(n24156), .B(n24155), .Z(n24198) );
  AND U24469 ( .A(a[60]), .B(b[55]), .Z(n24197) );
  XNOR U24470 ( .A(n24198), .B(n24197), .Z(n24199) );
  XOR U24471 ( .A(n24200), .B(n24199), .Z(n24194) );
  XNOR U24472 ( .A(n24193), .B(n24194), .Z(n24187) );
  NANDN U24473 ( .A(n24158), .B(n24157), .Z(n24162) );
  NANDN U24474 ( .A(n24160), .B(n24159), .Z(n24161) );
  AND U24475 ( .A(n24162), .B(n24161), .Z(n24186) );
  AND U24476 ( .A(a[62]), .B(b[53]), .Z(n24185) );
  XOR U24477 ( .A(n24186), .B(n24185), .Z(n24188) );
  XOR U24478 ( .A(n24187), .B(n24188), .Z(n24182) );
  XNOR U24479 ( .A(n24181), .B(n24182), .Z(n24178) );
  XNOR U24480 ( .A(n24177), .B(n24178), .Z(n24171) );
  NAND U24481 ( .A(n24164), .B(n24163), .Z(n24172) );
  XNOR U24482 ( .A(n24171), .B(n24172), .Z(n24174) );
  NANDN U24483 ( .A(n24166), .B(n24165), .Z(n24170) );
  NAND U24484 ( .A(n24168), .B(n24167), .Z(n24169) );
  AND U24485 ( .A(n24170), .B(n24169), .Z(n24173) );
  XOR U24486 ( .A(n24174), .B(n24173), .Z(c[115]) );
  NANDN U24487 ( .A(n24172), .B(n24171), .Z(n24176) );
  NAND U24488 ( .A(n24174), .B(n24173), .Z(n24175) );
  AND U24489 ( .A(n24176), .B(n24175), .Z(n24310) );
  ANDN U24490 ( .B(n24178), .A(n24177), .Z(n24308) );
  NANDN U24491 ( .A(n24180), .B(n24179), .Z(n24184) );
  NANDN U24492 ( .A(n24182), .B(n24181), .Z(n24183) );
  AND U24493 ( .A(n24184), .B(n24183), .Z(n24245) );
  NANDN U24494 ( .A(n24186), .B(n24185), .Z(n24190) );
  NANDN U24495 ( .A(n24188), .B(n24187), .Z(n24189) );
  AND U24496 ( .A(n24190), .B(n24189), .Z(n24248) );
  AND U24497 ( .A(a[63]), .B(b[53]), .Z(n24247) );
  XNOR U24498 ( .A(n24248), .B(n24247), .Z(n24249) );
  NANDN U24499 ( .A(n24192), .B(n24191), .Z(n24196) );
  NANDN U24500 ( .A(n24194), .B(n24193), .Z(n24195) );
  AND U24501 ( .A(n24196), .B(n24195), .Z(n24256) );
  NANDN U24502 ( .A(n24198), .B(n24197), .Z(n24202) );
  NANDN U24503 ( .A(n24200), .B(n24199), .Z(n24201) );
  AND U24504 ( .A(n24202), .B(n24201), .Z(n24302) );
  AND U24505 ( .A(a[61]), .B(b[55]), .Z(n24301) );
  XNOR U24506 ( .A(n24302), .B(n24301), .Z(n24303) );
  NANDN U24507 ( .A(n24204), .B(n24203), .Z(n24208) );
  NAND U24508 ( .A(n24206), .B(n24205), .Z(n24207) );
  AND U24509 ( .A(n24208), .B(n24207), .Z(n24261) );
  NANDN U24510 ( .A(n24210), .B(n24209), .Z(n24214) );
  OR U24511 ( .A(n24212), .B(n24211), .Z(n24213) );
  AND U24512 ( .A(n24214), .B(n24213), .Z(n24266) );
  AND U24513 ( .A(a[58]), .B(b[58]), .Z(n24265) );
  XNOR U24514 ( .A(n24266), .B(n24265), .Z(n24267) );
  NANDN U24515 ( .A(n24216), .B(n24215), .Z(n24220) );
  NANDN U24516 ( .A(n24218), .B(n24217), .Z(n24219) );
  AND U24517 ( .A(n24220), .B(n24219), .Z(n24278) );
  AND U24518 ( .A(a[56]), .B(b[60]), .Z(n24277) );
  XNOR U24519 ( .A(n24278), .B(n24277), .Z(n24279) );
  NANDN U24520 ( .A(n24222), .B(n24221), .Z(n24226) );
  NANDN U24521 ( .A(n24224), .B(n24223), .Z(n24225) );
  AND U24522 ( .A(n24226), .B(n24225), .Z(n24290) );
  AND U24523 ( .A(b[62]), .B(a[54]), .Z(n24289) );
  XNOR U24524 ( .A(n24290), .B(n24289), .Z(n24291) );
  NAND U24525 ( .A(b[63]), .B(a[53]), .Z(n24292) );
  XNOR U24526 ( .A(n24291), .B(n24292), .Z(n24285) );
  NANDN U24527 ( .A(n24228), .B(n24227), .Z(n24232) );
  NANDN U24528 ( .A(n24230), .B(n24229), .Z(n24231) );
  AND U24529 ( .A(n24232), .B(n24231), .Z(n24284) );
  AND U24530 ( .A(a[55]), .B(b[61]), .Z(n24283) );
  XOR U24531 ( .A(n24284), .B(n24283), .Z(n24286) );
  XOR U24532 ( .A(n24285), .B(n24286), .Z(n24280) );
  XNOR U24533 ( .A(n24279), .B(n24280), .Z(n24273) );
  NANDN U24534 ( .A(n24234), .B(n24233), .Z(n24238) );
  NANDN U24535 ( .A(n24236), .B(n24235), .Z(n24237) );
  AND U24536 ( .A(n24238), .B(n24237), .Z(n24272) );
  AND U24537 ( .A(a[57]), .B(b[59]), .Z(n24271) );
  XOR U24538 ( .A(n24272), .B(n24271), .Z(n24274) );
  XOR U24539 ( .A(n24273), .B(n24274), .Z(n24268) );
  XNOR U24540 ( .A(n24267), .B(n24268), .Z(n24295) );
  NANDN U24541 ( .A(n24240), .B(n24239), .Z(n24244) );
  NANDN U24542 ( .A(n24242), .B(n24241), .Z(n24243) );
  NAND U24543 ( .A(n24244), .B(n24243), .Z(n24296) );
  XNOR U24544 ( .A(n24295), .B(n24296), .Z(n24297) );
  NAND U24545 ( .A(a[59]), .B(b[57]), .Z(n24298) );
  XNOR U24546 ( .A(n24297), .B(n24298), .Z(n24259) );
  NAND U24547 ( .A(a[60]), .B(b[56]), .Z(n24260) );
  XOR U24548 ( .A(n24259), .B(n24260), .Z(n24262) );
  XOR U24549 ( .A(n24261), .B(n24262), .Z(n24304) );
  XNOR U24550 ( .A(n24303), .B(n24304), .Z(n24253) );
  NAND U24551 ( .A(a[62]), .B(b[54]), .Z(n24254) );
  XNOR U24552 ( .A(n24253), .B(n24254), .Z(n24255) );
  XOR U24553 ( .A(n24256), .B(n24255), .Z(n24250) );
  XOR U24554 ( .A(n24249), .B(n24250), .Z(n24246) );
  XNOR U24555 ( .A(n24245), .B(n24246), .Z(n24307) );
  XNOR U24556 ( .A(n24308), .B(n24307), .Z(n24309) );
  XNOR U24557 ( .A(n24310), .B(n24309), .Z(c[116]) );
  NOR U24558 ( .A(n24246), .B(n24245), .Z(n24370) );
  NANDN U24559 ( .A(n24248), .B(n24247), .Z(n24252) );
  NANDN U24560 ( .A(n24250), .B(n24249), .Z(n24251) );
  AND U24561 ( .A(n24252), .B(n24251), .Z(n24313) );
  NANDN U24562 ( .A(n24254), .B(n24253), .Z(n24258) );
  NANDN U24563 ( .A(n24256), .B(n24255), .Z(n24257) );
  AND U24564 ( .A(n24258), .B(n24257), .Z(n24316) );
  AND U24565 ( .A(a[63]), .B(b[54]), .Z(n24315) );
  XNOR U24566 ( .A(n24316), .B(n24315), .Z(n24317) );
  AND U24567 ( .A(a[61]), .B(b[56]), .Z(n24328) );
  NANDN U24568 ( .A(n24260), .B(n24259), .Z(n24264) );
  NANDN U24569 ( .A(n24262), .B(n24261), .Z(n24263) );
  AND U24570 ( .A(n24264), .B(n24263), .Z(n24327) );
  XNOR U24571 ( .A(n24328), .B(n24327), .Z(n24330) );
  AND U24572 ( .A(a[60]), .B(b[57]), .Z(n24366) );
  NANDN U24573 ( .A(n24266), .B(n24265), .Z(n24270) );
  NANDN U24574 ( .A(n24268), .B(n24267), .Z(n24269) );
  AND U24575 ( .A(n24270), .B(n24269), .Z(n24335) );
  NANDN U24576 ( .A(n24272), .B(n24271), .Z(n24276) );
  NANDN U24577 ( .A(n24274), .B(n24273), .Z(n24275) );
  AND U24578 ( .A(n24276), .B(n24275), .Z(n24358) );
  AND U24579 ( .A(a[58]), .B(b[59]), .Z(n24357) );
  XNOR U24580 ( .A(n24358), .B(n24357), .Z(n24359) );
  NANDN U24581 ( .A(n24278), .B(n24277), .Z(n24282) );
  NANDN U24582 ( .A(n24280), .B(n24279), .Z(n24281) );
  AND U24583 ( .A(n24282), .B(n24281), .Z(n24342) );
  NANDN U24584 ( .A(n24284), .B(n24283), .Z(n24288) );
  NANDN U24585 ( .A(n24286), .B(n24285), .Z(n24287) );
  AND U24586 ( .A(n24288), .B(n24287), .Z(n24352) );
  AND U24587 ( .A(a[56]), .B(b[61]), .Z(n24351) );
  XNOR U24588 ( .A(n24352), .B(n24351), .Z(n24353) );
  NANDN U24589 ( .A(n24290), .B(n24289), .Z(n24294) );
  NANDN U24590 ( .A(n24292), .B(n24291), .Z(n24293) );
  AND U24591 ( .A(n24294), .B(n24293), .Z(n24346) );
  AND U24592 ( .A(b[62]), .B(a[55]), .Z(n24345) );
  XNOR U24593 ( .A(n24346), .B(n24345), .Z(n24347) );
  NAND U24594 ( .A(b[63]), .B(a[54]), .Z(n24348) );
  XOR U24595 ( .A(n24347), .B(n24348), .Z(n24354) );
  XNOR U24596 ( .A(n24353), .B(n24354), .Z(n24339) );
  NAND U24597 ( .A(a[57]), .B(b[60]), .Z(n24340) );
  XNOR U24598 ( .A(n24339), .B(n24340), .Z(n24341) );
  XOR U24599 ( .A(n24342), .B(n24341), .Z(n24360) );
  XNOR U24600 ( .A(n24359), .B(n24360), .Z(n24333) );
  NAND U24601 ( .A(a[59]), .B(b[58]), .Z(n24334) );
  XOR U24602 ( .A(n24333), .B(n24334), .Z(n24336) );
  XOR U24603 ( .A(n24335), .B(n24336), .Z(n24364) );
  NANDN U24604 ( .A(n24296), .B(n24295), .Z(n24300) );
  NANDN U24605 ( .A(n24298), .B(n24297), .Z(n24299) );
  AND U24606 ( .A(n24300), .B(n24299), .Z(n24363) );
  XNOR U24607 ( .A(n24364), .B(n24363), .Z(n24365) );
  XNOR U24608 ( .A(n24366), .B(n24365), .Z(n24329) );
  XOR U24609 ( .A(n24330), .B(n24329), .Z(n24324) );
  NANDN U24610 ( .A(n24302), .B(n24301), .Z(n24306) );
  NANDN U24611 ( .A(n24304), .B(n24303), .Z(n24305) );
  AND U24612 ( .A(n24306), .B(n24305), .Z(n24322) );
  AND U24613 ( .A(a[62]), .B(b[55]), .Z(n24321) );
  XNOR U24614 ( .A(n24322), .B(n24321), .Z(n24323) );
  XOR U24615 ( .A(n24324), .B(n24323), .Z(n24318) );
  XOR U24616 ( .A(n24317), .B(n24318), .Z(n24314) );
  XNOR U24617 ( .A(n24313), .B(n24314), .Z(n24369) );
  XNOR U24618 ( .A(n24370), .B(n24369), .Z(n24372) );
  NANDN U24619 ( .A(n24308), .B(n24307), .Z(n24312) );
  NAND U24620 ( .A(n24310), .B(n24309), .Z(n24311) );
  NAND U24621 ( .A(n24312), .B(n24311), .Z(n24371) );
  XNOR U24622 ( .A(n24372), .B(n24371), .Z(c[117]) );
  NOR U24623 ( .A(n24314), .B(n24313), .Z(n24426) );
  NANDN U24624 ( .A(n24316), .B(n24315), .Z(n24320) );
  NANDN U24625 ( .A(n24318), .B(n24317), .Z(n24319) );
  AND U24626 ( .A(n24320), .B(n24319), .Z(n24375) );
  NANDN U24627 ( .A(n24322), .B(n24321), .Z(n24326) );
  NANDN U24628 ( .A(n24324), .B(n24323), .Z(n24325) );
  AND U24629 ( .A(n24326), .B(n24325), .Z(n24420) );
  AND U24630 ( .A(a[63]), .B(b[55]), .Z(n24419) );
  XNOR U24631 ( .A(n24420), .B(n24419), .Z(n24421) );
  NANDN U24632 ( .A(n24328), .B(n24327), .Z(n24332) );
  NAND U24633 ( .A(n24330), .B(n24329), .Z(n24331) );
  AND U24634 ( .A(n24332), .B(n24331), .Z(n24379) );
  NANDN U24635 ( .A(n24334), .B(n24333), .Z(n24338) );
  OR U24636 ( .A(n24336), .B(n24335), .Z(n24337) );
  AND U24637 ( .A(n24338), .B(n24337), .Z(n24384) );
  AND U24638 ( .A(a[60]), .B(b[58]), .Z(n24383) );
  XNOR U24639 ( .A(n24384), .B(n24383), .Z(n24385) );
  NANDN U24640 ( .A(n24340), .B(n24339), .Z(n24344) );
  NANDN U24641 ( .A(n24342), .B(n24341), .Z(n24343) );
  AND U24642 ( .A(n24344), .B(n24343), .Z(n24390) );
  AND U24643 ( .A(a[58]), .B(b[60]), .Z(n24389) );
  XNOR U24644 ( .A(n24390), .B(n24389), .Z(n24391) );
  NANDN U24645 ( .A(n24346), .B(n24345), .Z(n24350) );
  NANDN U24646 ( .A(n24348), .B(n24347), .Z(n24349) );
  AND U24647 ( .A(n24350), .B(n24349), .Z(n24402) );
  AND U24648 ( .A(b[62]), .B(a[56]), .Z(n24401) );
  XNOR U24649 ( .A(n24402), .B(n24401), .Z(n24403) );
  NAND U24650 ( .A(b[63]), .B(a[55]), .Z(n24404) );
  XNOR U24651 ( .A(n24403), .B(n24404), .Z(n24397) );
  NANDN U24652 ( .A(n24352), .B(n24351), .Z(n24356) );
  NANDN U24653 ( .A(n24354), .B(n24353), .Z(n24355) );
  AND U24654 ( .A(n24356), .B(n24355), .Z(n24396) );
  AND U24655 ( .A(a[57]), .B(b[61]), .Z(n24395) );
  XOR U24656 ( .A(n24396), .B(n24395), .Z(n24398) );
  XOR U24657 ( .A(n24397), .B(n24398), .Z(n24392) );
  XNOR U24658 ( .A(n24391), .B(n24392), .Z(n24409) );
  NANDN U24659 ( .A(n24358), .B(n24357), .Z(n24362) );
  NANDN U24660 ( .A(n24360), .B(n24359), .Z(n24361) );
  AND U24661 ( .A(n24362), .B(n24361), .Z(n24408) );
  AND U24662 ( .A(a[59]), .B(b[59]), .Z(n24407) );
  XOR U24663 ( .A(n24408), .B(n24407), .Z(n24410) );
  XOR U24664 ( .A(n24409), .B(n24410), .Z(n24386) );
  XNOR U24665 ( .A(n24385), .B(n24386), .Z(n24413) );
  NANDN U24666 ( .A(n24364), .B(n24363), .Z(n24368) );
  NANDN U24667 ( .A(n24366), .B(n24365), .Z(n24367) );
  NAND U24668 ( .A(n24368), .B(n24367), .Z(n24414) );
  XNOR U24669 ( .A(n24413), .B(n24414), .Z(n24415) );
  NAND U24670 ( .A(a[61]), .B(b[57]), .Z(n24416) );
  XNOR U24671 ( .A(n24415), .B(n24416), .Z(n24377) );
  NAND U24672 ( .A(a[62]), .B(b[56]), .Z(n24378) );
  XOR U24673 ( .A(n24377), .B(n24378), .Z(n24380) );
  XOR U24674 ( .A(n24379), .B(n24380), .Z(n24422) );
  XOR U24675 ( .A(n24421), .B(n24422), .Z(n24376) );
  XNOR U24676 ( .A(n24375), .B(n24376), .Z(n24425) );
  XNOR U24677 ( .A(n24426), .B(n24425), .Z(n24428) );
  NANDN U24678 ( .A(n24370), .B(n24369), .Z(n24374) );
  NAND U24679 ( .A(n24372), .B(n24371), .Z(n24373) );
  NAND U24680 ( .A(n24374), .B(n24373), .Z(n24427) );
  XNOR U24681 ( .A(n24428), .B(n24427), .Z(c[118]) );
  NOR U24682 ( .A(n24376), .B(n24375), .Z(n24476) );
  AND U24683 ( .A(a[63]), .B(b[56]), .Z(n24470) );
  NANDN U24684 ( .A(n24378), .B(n24377), .Z(n24382) );
  NANDN U24685 ( .A(n24380), .B(n24379), .Z(n24381) );
  AND U24686 ( .A(n24382), .B(n24381), .Z(n24469) );
  XNOR U24687 ( .A(n24470), .B(n24469), .Z(n24472) );
  AND U24688 ( .A(a[62]), .B(b[57]), .Z(n24466) );
  NANDN U24689 ( .A(n24384), .B(n24383), .Z(n24388) );
  NANDN U24690 ( .A(n24386), .B(n24385), .Z(n24387) );
  AND U24691 ( .A(n24388), .B(n24387), .Z(n24459) );
  NANDN U24692 ( .A(n24390), .B(n24389), .Z(n24394) );
  NANDN U24693 ( .A(n24392), .B(n24391), .Z(n24393) );
  AND U24694 ( .A(n24394), .B(n24393), .Z(n24435) );
  NANDN U24695 ( .A(n24396), .B(n24395), .Z(n24400) );
  NANDN U24696 ( .A(n24398), .B(n24397), .Z(n24399) );
  AND U24697 ( .A(n24400), .B(n24399), .Z(n24446) );
  AND U24698 ( .A(a[58]), .B(b[61]), .Z(n24445) );
  XNOR U24699 ( .A(n24446), .B(n24445), .Z(n24447) );
  NANDN U24700 ( .A(n24402), .B(n24401), .Z(n24406) );
  NANDN U24701 ( .A(n24404), .B(n24403), .Z(n24405) );
  AND U24702 ( .A(n24406), .B(n24405), .Z(n24442) );
  AND U24703 ( .A(b[62]), .B(a[57]), .Z(n24439) );
  NAND U24704 ( .A(b[63]), .B(a[56]), .Z(n24440) );
  XNOR U24705 ( .A(n24439), .B(n24440), .Z(n24441) );
  XOR U24706 ( .A(n24442), .B(n24441), .Z(n24448) );
  XNOR U24707 ( .A(n24447), .B(n24448), .Z(n24433) );
  NAND U24708 ( .A(a[59]), .B(b[60]), .Z(n24434) );
  XOR U24709 ( .A(n24433), .B(n24434), .Z(n24436) );
  XOR U24710 ( .A(n24435), .B(n24436), .Z(n24453) );
  AND U24711 ( .A(a[60]), .B(b[59]), .Z(n24452) );
  NANDN U24712 ( .A(n24408), .B(n24407), .Z(n24412) );
  NANDN U24713 ( .A(n24410), .B(n24409), .Z(n24411) );
  AND U24714 ( .A(n24412), .B(n24411), .Z(n24451) );
  XOR U24715 ( .A(n24452), .B(n24451), .Z(n24454) );
  XOR U24716 ( .A(n24453), .B(n24454), .Z(n24458) );
  AND U24717 ( .A(a[61]), .B(b[58]), .Z(n24457) );
  XOR U24718 ( .A(n24458), .B(n24457), .Z(n24460) );
  XOR U24719 ( .A(n24459), .B(n24460), .Z(n24464) );
  NANDN U24720 ( .A(n24414), .B(n24413), .Z(n24418) );
  NANDN U24721 ( .A(n24416), .B(n24415), .Z(n24417) );
  AND U24722 ( .A(n24418), .B(n24417), .Z(n24463) );
  XNOR U24723 ( .A(n24464), .B(n24463), .Z(n24465) );
  XNOR U24724 ( .A(n24466), .B(n24465), .Z(n24471) );
  XOR U24725 ( .A(n24472), .B(n24471), .Z(n24432) );
  NANDN U24726 ( .A(n24420), .B(n24419), .Z(n24424) );
  NANDN U24727 ( .A(n24422), .B(n24421), .Z(n24423) );
  AND U24728 ( .A(n24424), .B(n24423), .Z(n24431) );
  XNOR U24729 ( .A(n24432), .B(n24431), .Z(n24475) );
  XNOR U24730 ( .A(n24476), .B(n24475), .Z(n24478) );
  NANDN U24731 ( .A(n24426), .B(n24425), .Z(n24430) );
  NAND U24732 ( .A(n24428), .B(n24427), .Z(n24429) );
  NAND U24733 ( .A(n24430), .B(n24429), .Z(n24477) );
  XNOR U24734 ( .A(n24478), .B(n24477), .Z(c[119]) );
  NOR U24735 ( .A(n24432), .B(n24431), .Z(n24520) );
  NANDN U24736 ( .A(n24434), .B(n24433), .Z(n24438) );
  OR U24737 ( .A(n24436), .B(n24435), .Z(n24437) );
  AND U24738 ( .A(n24438), .B(n24437), .Z(n24496) );
  AND U24739 ( .A(a[60]), .B(b[60]), .Z(n24495) );
  XNOR U24740 ( .A(n24496), .B(n24495), .Z(n24497) );
  NANDN U24741 ( .A(n24440), .B(n24439), .Z(n24444) );
  NANDN U24742 ( .A(n24442), .B(n24441), .Z(n24443) );
  AND U24743 ( .A(n24444), .B(n24443), .Z(n24502) );
  AND U24744 ( .A(b[62]), .B(a[58]), .Z(n24501) );
  XNOR U24745 ( .A(n24502), .B(n24501), .Z(n24503) );
  NAND U24746 ( .A(b[63]), .B(a[57]), .Z(n24504) );
  XNOR U24747 ( .A(n24503), .B(n24504), .Z(n24509) );
  NANDN U24748 ( .A(n24446), .B(n24445), .Z(n24450) );
  NANDN U24749 ( .A(n24448), .B(n24447), .Z(n24449) );
  AND U24750 ( .A(n24450), .B(n24449), .Z(n24508) );
  AND U24751 ( .A(a[59]), .B(b[61]), .Z(n24507) );
  XOR U24752 ( .A(n24508), .B(n24507), .Z(n24510) );
  XOR U24753 ( .A(n24509), .B(n24510), .Z(n24498) );
  XNOR U24754 ( .A(n24497), .B(n24498), .Z(n24516) );
  NANDN U24755 ( .A(n24452), .B(n24451), .Z(n24456) );
  OR U24756 ( .A(n24454), .B(n24453), .Z(n24455) );
  AND U24757 ( .A(n24456), .B(n24455), .Z(n24513) );
  NAND U24758 ( .A(a[61]), .B(b[59]), .Z(n24514) );
  XNOR U24759 ( .A(n24513), .B(n24514), .Z(n24515) );
  XOR U24760 ( .A(n24516), .B(n24515), .Z(n24491) );
  AND U24761 ( .A(a[62]), .B(b[58]), .Z(n24490) );
  NANDN U24762 ( .A(n24458), .B(n24457), .Z(n24462) );
  OR U24763 ( .A(n24460), .B(n24459), .Z(n24461) );
  AND U24764 ( .A(n24462), .B(n24461), .Z(n24489) );
  XOR U24765 ( .A(n24490), .B(n24489), .Z(n24492) );
  XOR U24766 ( .A(n24491), .B(n24492), .Z(n24484) );
  NANDN U24767 ( .A(n24464), .B(n24463), .Z(n24468) );
  NANDN U24768 ( .A(n24466), .B(n24465), .Z(n24467) );
  AND U24769 ( .A(n24468), .B(n24467), .Z(n24483) );
  XNOR U24770 ( .A(n24484), .B(n24483), .Z(n24485) );
  NAND U24771 ( .A(a[63]), .B(b[57]), .Z(n24486) );
  XNOR U24772 ( .A(n24485), .B(n24486), .Z(n24482) );
  NANDN U24773 ( .A(n24470), .B(n24469), .Z(n24474) );
  NAND U24774 ( .A(n24472), .B(n24471), .Z(n24473) );
  AND U24775 ( .A(n24474), .B(n24473), .Z(n24481) );
  XNOR U24776 ( .A(n24482), .B(n24481), .Z(n24519) );
  XNOR U24777 ( .A(n24520), .B(n24519), .Z(n24522) );
  NANDN U24778 ( .A(n24476), .B(n24475), .Z(n24480) );
  NAND U24779 ( .A(n24478), .B(n24477), .Z(n24479) );
  NAND U24780 ( .A(n24480), .B(n24479), .Z(n24521) );
  XNOR U24781 ( .A(n24522), .B(n24521), .Z(c[120]) );
  AND U24782 ( .A(n24482), .B(n24481), .Z(n24558) );
  NANDN U24783 ( .A(n24484), .B(n24483), .Z(n24488) );
  NANDN U24784 ( .A(n24486), .B(n24485), .Z(n24487) );
  AND U24785 ( .A(n24488), .B(n24487), .Z(n24525) );
  NANDN U24786 ( .A(n24490), .B(n24489), .Z(n24494) );
  OR U24787 ( .A(n24492), .B(n24491), .Z(n24493) );
  AND U24788 ( .A(n24494), .B(n24493), .Z(n24527) );
  NAND U24789 ( .A(a[63]), .B(b[58]), .Z(n24528) );
  XNOR U24790 ( .A(n24527), .B(n24528), .Z(n24529) );
  NANDN U24791 ( .A(n24496), .B(n24495), .Z(n24500) );
  NANDN U24792 ( .A(n24498), .B(n24497), .Z(n24499) );
  AND U24793 ( .A(n24500), .B(n24499), .Z(n24540) );
  AND U24794 ( .A(a[61]), .B(b[60]), .Z(n24539) );
  XNOR U24795 ( .A(n24540), .B(n24539), .Z(n24541) );
  NANDN U24796 ( .A(n24502), .B(n24501), .Z(n24506) );
  NANDN U24797 ( .A(n24504), .B(n24503), .Z(n24505) );
  AND U24798 ( .A(n24506), .B(n24505), .Z(n24552) );
  AND U24799 ( .A(b[62]), .B(a[59]), .Z(n24551) );
  XNOR U24800 ( .A(n24552), .B(n24551), .Z(n24553) );
  NAND U24801 ( .A(b[63]), .B(a[58]), .Z(n24554) );
  XNOR U24802 ( .A(n24553), .B(n24554), .Z(n24547) );
  NANDN U24803 ( .A(n24508), .B(n24507), .Z(n24512) );
  NANDN U24804 ( .A(n24510), .B(n24509), .Z(n24511) );
  AND U24805 ( .A(n24512), .B(n24511), .Z(n24546) );
  AND U24806 ( .A(a[60]), .B(b[61]), .Z(n24545) );
  XOR U24807 ( .A(n24546), .B(n24545), .Z(n24548) );
  XOR U24808 ( .A(n24547), .B(n24548), .Z(n24542) );
  XNOR U24809 ( .A(n24541), .B(n24542), .Z(n24535) );
  NANDN U24810 ( .A(n24514), .B(n24513), .Z(n24518) );
  NAND U24811 ( .A(n24516), .B(n24515), .Z(n24517) );
  AND U24812 ( .A(n24518), .B(n24517), .Z(n24534) );
  AND U24813 ( .A(a[62]), .B(b[59]), .Z(n24533) );
  XOR U24814 ( .A(n24534), .B(n24533), .Z(n24536) );
  XOR U24815 ( .A(n24535), .B(n24536), .Z(n24530) );
  XOR U24816 ( .A(n24529), .B(n24530), .Z(n24526) );
  XNOR U24817 ( .A(n24525), .B(n24526), .Z(n24557) );
  XNOR U24818 ( .A(n24558), .B(n24557), .Z(n24560) );
  NANDN U24819 ( .A(n24520), .B(n24519), .Z(n24524) );
  NAND U24820 ( .A(n24522), .B(n24521), .Z(n24523) );
  NAND U24821 ( .A(n24524), .B(n24523), .Z(n24559) );
  XNOR U24822 ( .A(n24560), .B(n24559), .Z(c[121]) );
  NOR U24823 ( .A(n24526), .B(n24525), .Z(n24590) );
  NANDN U24824 ( .A(n24528), .B(n24527), .Z(n24532) );
  NANDN U24825 ( .A(n24530), .B(n24529), .Z(n24531) );
  AND U24826 ( .A(n24532), .B(n24531), .Z(n24563) );
  NANDN U24827 ( .A(n24534), .B(n24533), .Z(n24538) );
  NANDN U24828 ( .A(n24536), .B(n24535), .Z(n24537) );
  AND U24829 ( .A(n24538), .B(n24537), .Z(n24566) );
  AND U24830 ( .A(a[63]), .B(b[59]), .Z(n24565) );
  XNOR U24831 ( .A(n24566), .B(n24565), .Z(n24567) );
  NANDN U24832 ( .A(n24540), .B(n24539), .Z(n24544) );
  NANDN U24833 ( .A(n24542), .B(n24541), .Z(n24543) );
  AND U24834 ( .A(n24544), .B(n24543), .Z(n24574) );
  NANDN U24835 ( .A(n24546), .B(n24545), .Z(n24550) );
  NANDN U24836 ( .A(n24548), .B(n24547), .Z(n24549) );
  AND U24837 ( .A(n24550), .B(n24549), .Z(n24584) );
  AND U24838 ( .A(a[61]), .B(b[61]), .Z(n24583) );
  XNOR U24839 ( .A(n24584), .B(n24583), .Z(n24585) );
  NANDN U24840 ( .A(n24552), .B(n24551), .Z(n24556) );
  NANDN U24841 ( .A(n24554), .B(n24553), .Z(n24555) );
  AND U24842 ( .A(n24556), .B(n24555), .Z(n24580) );
  AND U24843 ( .A(b[62]), .B(a[60]), .Z(n24577) );
  NAND U24844 ( .A(b[63]), .B(a[59]), .Z(n24578) );
  XNOR U24845 ( .A(n24577), .B(n24578), .Z(n24579) );
  XOR U24846 ( .A(n24580), .B(n24579), .Z(n24586) );
  XNOR U24847 ( .A(n24585), .B(n24586), .Z(n24571) );
  NAND U24848 ( .A(a[62]), .B(b[60]), .Z(n24572) );
  XNOR U24849 ( .A(n24571), .B(n24572), .Z(n24573) );
  XOR U24850 ( .A(n24574), .B(n24573), .Z(n24568) );
  XOR U24851 ( .A(n24567), .B(n24568), .Z(n24564) );
  XNOR U24852 ( .A(n24563), .B(n24564), .Z(n24589) );
  XNOR U24853 ( .A(n24590), .B(n24589), .Z(n24592) );
  NANDN U24854 ( .A(n24558), .B(n24557), .Z(n24562) );
  NAND U24855 ( .A(n24560), .B(n24559), .Z(n24561) );
  NAND U24856 ( .A(n24562), .B(n24561), .Z(n24591) );
  XNOR U24857 ( .A(n24592), .B(n24591), .Z(c[122]) );
  NOR U24858 ( .A(n24564), .B(n24563), .Z(n24616) );
  NANDN U24859 ( .A(n24566), .B(n24565), .Z(n24570) );
  NANDN U24860 ( .A(n24568), .B(n24567), .Z(n24569) );
  AND U24861 ( .A(n24570), .B(n24569), .Z(n24595) );
  NANDN U24862 ( .A(n24572), .B(n24571), .Z(n24576) );
  NANDN U24863 ( .A(n24574), .B(n24573), .Z(n24575) );
  AND U24864 ( .A(n24576), .B(n24575), .Z(n24598) );
  AND U24865 ( .A(a[63]), .B(b[60]), .Z(n24597) );
  XNOR U24866 ( .A(n24598), .B(n24597), .Z(n24599) );
  NANDN U24867 ( .A(n24578), .B(n24577), .Z(n24582) );
  NANDN U24868 ( .A(n24580), .B(n24579), .Z(n24581) );
  AND U24869 ( .A(n24582), .B(n24581), .Z(n24604) );
  AND U24870 ( .A(b[62]), .B(a[61]), .Z(n24603) );
  XNOR U24871 ( .A(n24604), .B(n24603), .Z(n24605) );
  NAND U24872 ( .A(b[63]), .B(a[60]), .Z(n24606) );
  XNOR U24873 ( .A(n24605), .B(n24606), .Z(n24611) );
  NANDN U24874 ( .A(n24584), .B(n24583), .Z(n24588) );
  NANDN U24875 ( .A(n24586), .B(n24585), .Z(n24587) );
  AND U24876 ( .A(n24588), .B(n24587), .Z(n24610) );
  AND U24877 ( .A(a[62]), .B(b[61]), .Z(n24609) );
  XOR U24878 ( .A(n24610), .B(n24609), .Z(n24612) );
  XOR U24879 ( .A(n24611), .B(n24612), .Z(n24600) );
  XOR U24880 ( .A(n24599), .B(n24600), .Z(n24596) );
  XNOR U24881 ( .A(n24595), .B(n24596), .Z(n24615) );
  XNOR U24882 ( .A(n24616), .B(n24615), .Z(n24618) );
  NANDN U24883 ( .A(n24590), .B(n24589), .Z(n24594) );
  NAND U24884 ( .A(n24592), .B(n24591), .Z(n24593) );
  NAND U24885 ( .A(n24594), .B(n24593), .Z(n24617) );
  XNOR U24886 ( .A(n24618), .B(n24617), .Z(c[123]) );
  NOR U24887 ( .A(n24596), .B(n24595), .Z(n24636) );
  NANDN U24888 ( .A(n24598), .B(n24597), .Z(n24602) );
  NANDN U24889 ( .A(n24600), .B(n24599), .Z(n24601) );
  AND U24890 ( .A(n24602), .B(n24601), .Z(n24621) );
  NANDN U24891 ( .A(n24604), .B(n24603), .Z(n24608) );
  NANDN U24892 ( .A(n24606), .B(n24605), .Z(n24607) );
  AND U24893 ( .A(n24608), .B(n24607), .Z(n24626) );
  AND U24894 ( .A(b[62]), .B(a[62]), .Z(n24623) );
  NAND U24895 ( .A(a[61]), .B(b[63]), .Z(n24624) );
  XNOR U24896 ( .A(n24623), .B(n24624), .Z(n24625) );
  XNOR U24897 ( .A(n24626), .B(n24625), .Z(n24631) );
  NANDN U24898 ( .A(n24610), .B(n24609), .Z(n24614) );
  NANDN U24899 ( .A(n24612), .B(n24611), .Z(n24613) );
  AND U24900 ( .A(n24614), .B(n24613), .Z(n24630) );
  AND U24901 ( .A(a[63]), .B(b[61]), .Z(n24629) );
  XOR U24902 ( .A(n24630), .B(n24629), .Z(n24632) );
  XOR U24903 ( .A(n24631), .B(n24632), .Z(n24622) );
  XNOR U24904 ( .A(n24621), .B(n24622), .Z(n24635) );
  XNOR U24905 ( .A(n24636), .B(n24635), .Z(n24638) );
  NANDN U24906 ( .A(n24616), .B(n24615), .Z(n24620) );
  NAND U24907 ( .A(n24618), .B(n24617), .Z(n24619) );
  NAND U24908 ( .A(n24620), .B(n24619), .Z(n24637) );
  XNOR U24909 ( .A(n24638), .B(n24637), .Z(c[124]) );
  NOR U24910 ( .A(n24622), .B(n24621), .Z(n24649) );
  NAND U24911 ( .A(a[62]), .B(b[63]), .Z(n24645) );
  NAND U24912 ( .A(a[63]), .B(b[62]), .Z(n24644) );
  NANDN U24913 ( .A(n24624), .B(n24623), .Z(n24628) );
  NANDN U24914 ( .A(n24626), .B(n24625), .Z(n24627) );
  AND U24915 ( .A(n24628), .B(n24627), .Z(n24643) );
  XNOR U24916 ( .A(n24644), .B(n24643), .Z(n24646) );
  XOR U24917 ( .A(n24645), .B(n24646), .Z(n24641) );
  NANDN U24918 ( .A(n24630), .B(n24629), .Z(n24634) );
  NANDN U24919 ( .A(n24632), .B(n24631), .Z(n24633) );
  AND U24920 ( .A(n24634), .B(n24633), .Z(n24642) );
  XOR U24921 ( .A(n24641), .B(n24642), .Z(n24648) );
  XNOR U24922 ( .A(n24649), .B(n24648), .Z(n24651) );
  NANDN U24923 ( .A(n24636), .B(n24635), .Z(n24640) );
  NAND U24924 ( .A(n24638), .B(n24637), .Z(n24639) );
  NAND U24925 ( .A(n24640), .B(n24639), .Z(n24650) );
  XNOR U24926 ( .A(n24651), .B(n24650), .Z(c[125]) );
  NAND U24927 ( .A(b[63]), .B(a[63]), .Z(n24647) );
  XOR U24928 ( .A(n24654), .B(n24647), .Z(n24657) );
  XNOR U24929 ( .A(n24658), .B(n24657), .Z(n24656) );
  NANDN U24930 ( .A(n24649), .B(n24648), .Z(n24653) );
  NAND U24931 ( .A(n24651), .B(n24650), .Z(n24652) );
  NAND U24932 ( .A(n24653), .B(n24652), .Z(n24655) );
  XNOR U24933 ( .A(n24656), .B(n24655), .Z(c[126]) );
  XOR U24934 ( .A(n24660), .B(n24659), .Z(c[65]) );
  XOR U24935 ( .A(n24662), .B(n24661), .Z(c[66]) );
  XNOR U24936 ( .A(n24664), .B(n24663), .Z(n24665) );
  XNOR U24937 ( .A(n24666), .B(n24665), .Z(c[67]) );
  XNOR U24938 ( .A(n24668), .B(n24667), .Z(n24669) );
  XOR U24939 ( .A(n24670), .B(n24669), .Z(c[68]) );
  NAND U24940 ( .A(n24670), .B(n24669), .Z(n24671) );
  NANDN U24941 ( .A(n24672), .B(n24671), .Z(n24676) );
  XNOR U24942 ( .A(n24674), .B(n24673), .Z(n24675) );
  XNOR U24943 ( .A(n24676), .B(n24675), .Z(c[69]) );
  XNOR U24944 ( .A(n24678), .B(n24677), .Z(n24679) );
  XNOR U24945 ( .A(n24680), .B(n24679), .Z(c[70]) );
  XOR U24946 ( .A(n24682), .B(n24681), .Z(n24685) );
  XNOR U24947 ( .A(n24686), .B(n24685), .Z(c[71]) );
  XNOR U24948 ( .A(n24684), .B(n24683), .Z(n24690) );
  NANDN U24949 ( .A(n24686), .B(n24685), .Z(n24687) );
  NANDN U24950 ( .A(n24688), .B(n24687), .Z(n24689) );
  XOR U24951 ( .A(n24690), .B(n24689), .Z(c[72]) );
  NAND U24952 ( .A(n24690), .B(n24689), .Z(n24691) );
  NAND U24953 ( .A(n24692), .B(n24691), .Z(n24696) );
  XOR U24954 ( .A(n24694), .B(n24693), .Z(n24695) );
  XNOR U24955 ( .A(n24696), .B(n24695), .Z(c[73]) );
  XOR U24956 ( .A(n24698), .B(n24697), .Z(n24699) );
  XNOR U24957 ( .A(n24700), .B(n24699), .Z(c[74]) );
  XOR U24958 ( .A(n24702), .B(n24701), .Z(n24708) );
  AND U24959 ( .A(n24704), .B(n24703), .Z(n24707) );
  XNOR U24960 ( .A(n24708), .B(n24707), .Z(c[75]) );
  XNOR U24961 ( .A(n24706), .B(n24705), .Z(n24712) );
  NAND U24962 ( .A(n24708), .B(n24707), .Z(n24709) );
  NAND U24963 ( .A(n24710), .B(n24709), .Z(n24711) );
  XNOR U24964 ( .A(n24712), .B(n24711), .Z(c[76]) );
  NAND U24965 ( .A(n24712), .B(n24711), .Z(n24714) );
  AND U24966 ( .A(n24714), .B(n24713), .Z(n24718) );
  XNOR U24967 ( .A(n24716), .B(n24715), .Z(n24717) );
  XNOR U24968 ( .A(n24718), .B(n24717), .Z(c[77]) );
  XNOR U24969 ( .A(n24720), .B(n24719), .Z(c[78]) );
  XOR U24970 ( .A(n24722), .B(n24721), .Z(n24723) );
  XNOR U24971 ( .A(n24724), .B(n24723), .Z(c[79]) );
  XOR U24972 ( .A(n24726), .B(n24725), .Z(c[80]) );
  XOR U24973 ( .A(n24728), .B(n24727), .Z(c[81]) );
  XNOR U24974 ( .A(n24730), .B(n24729), .Z(c[82]) );
  XNOR U24975 ( .A(n24732), .B(n24731), .Z(c[83]) );
  XNOR U24976 ( .A(n24734), .B(n24733), .Z(c[84]) );
  XNOR U24977 ( .A(n24736), .B(n24735), .Z(c[85]) );
  XOR U24978 ( .A(n24738), .B(n24737), .Z(n24742) );
  XNOR U24979 ( .A(n24742), .B(n24741), .Z(c[86]) );
  XOR U24980 ( .A(n24740), .B(n24739), .Z(n24748) );
  NAND U24981 ( .A(n24742), .B(n24741), .Z(n24743) );
  NAND U24982 ( .A(n24744), .B(n24743), .Z(n24747) );
  XNOR U24983 ( .A(n24748), .B(n24747), .Z(c[87]) );
  XOR U24984 ( .A(n24746), .B(n24745), .Z(n24752) );
  NAND U24985 ( .A(n24748), .B(n24747), .Z(n24749) );
  NANDN U24986 ( .A(n24750), .B(n24749), .Z(n24751) );
  XNOR U24987 ( .A(n24752), .B(n24751), .Z(c[88]) );
  NAND U24988 ( .A(n24752), .B(n24751), .Z(n24754) );
  AND U24989 ( .A(n24754), .B(n24753), .Z(n24758) );
  XNOR U24990 ( .A(n24756), .B(n24755), .Z(n24757) );
  XNOR U24991 ( .A(n24758), .B(n24757), .Z(c[89]) );
  XOR U24992 ( .A(n24760), .B(n24759), .Z(n24761) );
  XOR U24993 ( .A(n24762), .B(n24761), .Z(c[90]) );
  XNOR U24994 ( .A(n24764), .B(n24763), .Z(n24765) );
  XOR U24995 ( .A(n24766), .B(n24765), .Z(c[91]) );
  XOR U24996 ( .A(n24768), .B(n24767), .Z(n24769) );
  XOR U24997 ( .A(n24770), .B(n24769), .Z(c[92]) );
  NANDN U24998 ( .A(n24770), .B(n24769), .Z(n24771) );
  AND U24999 ( .A(n24772), .B(n24771), .Z(n24774) );
  XNOR U25000 ( .A(n24774), .B(n24773), .Z(n24775) );
  XNOR U25001 ( .A(n24776), .B(n24775), .Z(c[93]) );
  XNOR U25002 ( .A(n24778), .B(n24777), .Z(c[94]) );
  XNOR U25003 ( .A(n24780), .B(n24779), .Z(c[95]) );
  XNOR U25004 ( .A(n24782), .B(n24781), .Z(c[96]) );
  XOR U25005 ( .A(n24784), .B(n24783), .Z(n24785) );
  XNOR U25006 ( .A(n24786), .B(n24785), .Z(c[97]) );
  XOR U25007 ( .A(n24788), .B(n24787), .Z(c[98]) );
  XOR U25008 ( .A(n24790), .B(n24789), .Z(c[99]) );
  XNOR U25009 ( .A(n24792), .B(n24791), .Z(c[100]) );
  XOR U25010 ( .A(n24794), .B(n24793), .Z(n24795) );
  XNOR U25011 ( .A(n24796), .B(n24795), .Z(c[101]) );
  XOR U25012 ( .A(n24798), .B(n24797), .Z(c[2]) );
  XOR U25013 ( .A(n24800), .B(n24799), .Z(c[12]) );
  XNOR U25014 ( .A(n24802), .B(n24801), .Z(c[13]) );
  XOR U25015 ( .A(n24804), .B(n24803), .Z(c[14]) );
  XNOR U25016 ( .A(n24806), .B(n24805), .Z(c[15]) );
  XOR U25017 ( .A(n24808), .B(n24807), .Z(c[16]) );
  XNOR U25018 ( .A(n24810), .B(n24809), .Z(c[17]) );
  XOR U25019 ( .A(n24812), .B(n24811), .Z(n24813) );
  XNOR U25020 ( .A(n24814), .B(n24813), .Z(c[18]) );
  XNOR U25021 ( .A(n24816), .B(n24815), .Z(c[19]) );
  XOR U25022 ( .A(n24818), .B(n24817), .Z(n24819) );
  XNOR U25023 ( .A(n24820), .B(n24819), .Z(c[20]) );
  XNOR U25024 ( .A(n24822), .B(n24821), .Z(c[21]) );
  XNOR U25025 ( .A(n24824), .B(n24823), .Z(c[3]) );
  XOR U25026 ( .A(n24826), .B(n24825), .Z(n24827) );
  XNOR U25027 ( .A(n24828), .B(n24827), .Z(c[22]) );
  XNOR U25028 ( .A(n24830), .B(n24829), .Z(c[23]) );
  XOR U25029 ( .A(n24832), .B(n24831), .Z(n24833) );
  XNOR U25030 ( .A(n24834), .B(n24833), .Z(c[24]) );
  XNOR U25031 ( .A(n24836), .B(n24835), .Z(c[25]) );
  XOR U25032 ( .A(n24838), .B(n24837), .Z(n24839) );
  XNOR U25033 ( .A(n24840), .B(n24839), .Z(c[26]) );
  XNOR U25034 ( .A(n24842), .B(n24841), .Z(c[27]) );
  XOR U25035 ( .A(n24844), .B(n24843), .Z(n24845) );
  XNOR U25036 ( .A(n24846), .B(n24845), .Z(c[28]) );
  XNOR U25037 ( .A(n24848), .B(n24847), .Z(c[29]) );
  XOR U25038 ( .A(n24850), .B(n24849), .Z(n24851) );
  XNOR U25039 ( .A(n24852), .B(n24851), .Z(c[30]) );
  XNOR U25040 ( .A(n24854), .B(n24853), .Z(c[31]) );
  XOR U25041 ( .A(n24856), .B(n24855), .Z(c[4]) );
  XOR U25042 ( .A(n24858), .B(n24857), .Z(n24859) );
  XNOR U25043 ( .A(n24860), .B(n24859), .Z(c[32]) );
  XNOR U25044 ( .A(n24862), .B(n24861), .Z(c[33]) );
  XOR U25045 ( .A(n24864), .B(n24863), .Z(n24865) );
  XNOR U25046 ( .A(n24866), .B(n24865), .Z(c[34]) );
  XNOR U25047 ( .A(n24868), .B(n24867), .Z(c[35]) );
  XOR U25048 ( .A(n24870), .B(n24869), .Z(n24871) );
  XNOR U25049 ( .A(n24872), .B(n24871), .Z(c[36]) );
  XNOR U25050 ( .A(n24874), .B(n24873), .Z(c[37]) );
  XOR U25051 ( .A(n24876), .B(n24875), .Z(n24877) );
  XNOR U25052 ( .A(n24878), .B(n24877), .Z(c[38]) );
  XNOR U25053 ( .A(n24880), .B(n24879), .Z(c[39]) );
  XOR U25054 ( .A(n24882), .B(n24881), .Z(n24883) );
  XNOR U25055 ( .A(n24884), .B(n24883), .Z(c[40]) );
  XNOR U25056 ( .A(n24886), .B(n24885), .Z(c[41]) );
  XNOR U25057 ( .A(n24888), .B(n24887), .Z(c[5]) );
  XOR U25058 ( .A(n24890), .B(n24889), .Z(n24891) );
  XNOR U25059 ( .A(n24892), .B(n24891), .Z(c[42]) );
  XNOR U25060 ( .A(n24894), .B(n24893), .Z(c[43]) );
  XOR U25061 ( .A(n24896), .B(n24895), .Z(n24897) );
  XNOR U25062 ( .A(n24898), .B(n24897), .Z(c[44]) );
  XNOR U25063 ( .A(n24900), .B(n24899), .Z(c[45]) );
  XOR U25064 ( .A(n24902), .B(n24901), .Z(n24903) );
  XNOR U25065 ( .A(n24904), .B(n24903), .Z(c[46]) );
  XNOR U25066 ( .A(n24906), .B(n24905), .Z(c[47]) );
  XOR U25067 ( .A(n24908), .B(n24907), .Z(n24909) );
  XNOR U25068 ( .A(n24910), .B(n24909), .Z(c[48]) );
  XNOR U25069 ( .A(n24912), .B(n24911), .Z(c[49]) );
  XOR U25070 ( .A(n24914), .B(n24913), .Z(n24915) );
  XNOR U25071 ( .A(n24916), .B(n24915), .Z(c[50]) );
  XNOR U25072 ( .A(n24918), .B(n24917), .Z(c[51]) );
  XNOR U25073 ( .A(n24920), .B(n24919), .Z(c[6]) );
  XOR U25074 ( .A(n24922), .B(n24921), .Z(n24923) );
  XNOR U25075 ( .A(n24924), .B(n24923), .Z(c[52]) );
  XNOR U25076 ( .A(n24926), .B(n24925), .Z(c[53]) );
  XOR U25077 ( .A(n24928), .B(n24927), .Z(n24929) );
  XNOR U25078 ( .A(n24930), .B(n24929), .Z(c[54]) );
  XNOR U25079 ( .A(n24932), .B(n24931), .Z(c[55]) );
  XOR U25080 ( .A(n24934), .B(n24933), .Z(n24935) );
  XNOR U25081 ( .A(n24936), .B(n24935), .Z(c[56]) );
  XNOR U25082 ( .A(n24938), .B(n24937), .Z(c[57]) );
  XOR U25083 ( .A(n24940), .B(n24939), .Z(n24941) );
  XNOR U25084 ( .A(n24942), .B(n24941), .Z(c[58]) );
  XNOR U25085 ( .A(n24944), .B(n24943), .Z(c[59]) );
  XOR U25086 ( .A(n24946), .B(n24945), .Z(n24947) );
  XNOR U25087 ( .A(n24948), .B(n24947), .Z(c[60]) );
  XNOR U25088 ( .A(n24950), .B(n24949), .Z(c[61]) );
  XNOR U25089 ( .A(n24952), .B(n24951), .Z(c[7]) );
  XOR U25090 ( .A(n24954), .B(n24953), .Z(n24955) );
  XNOR U25091 ( .A(n24956), .B(n24955), .Z(c[62]) );
  XNOR U25092 ( .A(n24958), .B(n24957), .Z(c[63]) );
  XOR U25093 ( .A(n24960), .B(n24959), .Z(c[64]) );
  XOR U25094 ( .A(n24962), .B(n24961), .Z(c[8]) );
  XNOR U25095 ( .A(n24964), .B(n24963), .Z(c[9]) );
  XOR U25096 ( .A(n24966), .B(n24965), .Z(n24967) );
  XNOR U25097 ( .A(n24968), .B(n24967), .Z(c[10]) );
  XNOR U25098 ( .A(n24970), .B(n24969), .Z(c[11]) );
  NAND U25099 ( .A(b[0]), .B(a[1]), .Z(n24971) );
  XNOR U25100 ( .A(n24972), .B(n24971), .Z(c[1]) );
endmodule

