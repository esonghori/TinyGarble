
module mult_N128_CC64 ( clk, rst, a, b, c );
  input [127:0] a;
  input [1:0] b;
  output [127:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991;
  wire   [127:2] swire;
  wire   [255:128] sreg;

  DFF \sreg_reg[128]  ( .D(swire[2]), .CLK(clk), .RST(rst), .Q(sreg[128]) );
  DFF \sreg_reg[129]  ( .D(swire[3]), .CLK(clk), .RST(rst), .Q(sreg[129]) );
  DFF \sreg_reg[130]  ( .D(swire[4]), .CLK(clk), .RST(rst), .Q(sreg[130]) );
  DFF \sreg_reg[131]  ( .D(swire[5]), .CLK(clk), .RST(rst), .Q(sreg[131]) );
  DFF \sreg_reg[132]  ( .D(swire[6]), .CLK(clk), .RST(rst), .Q(sreg[132]) );
  DFF \sreg_reg[133]  ( .D(swire[7]), .CLK(clk), .RST(rst), .Q(sreg[133]) );
  DFF \sreg_reg[134]  ( .D(swire[8]), .CLK(clk), .RST(rst), .Q(sreg[134]) );
  DFF \sreg_reg[135]  ( .D(swire[9]), .CLK(clk), .RST(rst), .Q(sreg[135]) );
  DFF \sreg_reg[136]  ( .D(swire[10]), .CLK(clk), .RST(rst), .Q(sreg[136]) );
  DFF \sreg_reg[137]  ( .D(swire[11]), .CLK(clk), .RST(rst), .Q(sreg[137]) );
  DFF \sreg_reg[138]  ( .D(swire[12]), .CLK(clk), .RST(rst), .Q(sreg[138]) );
  DFF \sreg_reg[139]  ( .D(swire[13]), .CLK(clk), .RST(rst), .Q(sreg[139]) );
  DFF \sreg_reg[140]  ( .D(swire[14]), .CLK(clk), .RST(rst), .Q(sreg[140]) );
  DFF \sreg_reg[141]  ( .D(swire[15]), .CLK(clk), .RST(rst), .Q(sreg[141]) );
  DFF \sreg_reg[142]  ( .D(swire[16]), .CLK(clk), .RST(rst), .Q(sreg[142]) );
  DFF \sreg_reg[143]  ( .D(swire[17]), .CLK(clk), .RST(rst), .Q(sreg[143]) );
  DFF \sreg_reg[144]  ( .D(swire[18]), .CLK(clk), .RST(rst), .Q(sreg[144]) );
  DFF \sreg_reg[145]  ( .D(swire[19]), .CLK(clk), .RST(rst), .Q(sreg[145]) );
  DFF \sreg_reg[146]  ( .D(swire[20]), .CLK(clk), .RST(rst), .Q(sreg[146]) );
  DFF \sreg_reg[147]  ( .D(swire[21]), .CLK(clk), .RST(rst), .Q(sreg[147]) );
  DFF \sreg_reg[148]  ( .D(swire[22]), .CLK(clk), .RST(rst), .Q(sreg[148]) );
  DFF \sreg_reg[149]  ( .D(swire[23]), .CLK(clk), .RST(rst), .Q(sreg[149]) );
  DFF \sreg_reg[150]  ( .D(swire[24]), .CLK(clk), .RST(rst), .Q(sreg[150]) );
  DFF \sreg_reg[151]  ( .D(swire[25]), .CLK(clk), .RST(rst), .Q(sreg[151]) );
  DFF \sreg_reg[152]  ( .D(swire[26]), .CLK(clk), .RST(rst), .Q(sreg[152]) );
  DFF \sreg_reg[153]  ( .D(swire[27]), .CLK(clk), .RST(rst), .Q(sreg[153]) );
  DFF \sreg_reg[154]  ( .D(swire[28]), .CLK(clk), .RST(rst), .Q(sreg[154]) );
  DFF \sreg_reg[155]  ( .D(swire[29]), .CLK(clk), .RST(rst), .Q(sreg[155]) );
  DFF \sreg_reg[156]  ( .D(swire[30]), .CLK(clk), .RST(rst), .Q(sreg[156]) );
  DFF \sreg_reg[157]  ( .D(swire[31]), .CLK(clk), .RST(rst), .Q(sreg[157]) );
  DFF \sreg_reg[158]  ( .D(swire[32]), .CLK(clk), .RST(rst), .Q(sreg[158]) );
  DFF \sreg_reg[159]  ( .D(swire[33]), .CLK(clk), .RST(rst), .Q(sreg[159]) );
  DFF \sreg_reg[160]  ( .D(swire[34]), .CLK(clk), .RST(rst), .Q(sreg[160]) );
  DFF \sreg_reg[161]  ( .D(swire[35]), .CLK(clk), .RST(rst), .Q(sreg[161]) );
  DFF \sreg_reg[162]  ( .D(swire[36]), .CLK(clk), .RST(rst), .Q(sreg[162]) );
  DFF \sreg_reg[163]  ( .D(swire[37]), .CLK(clk), .RST(rst), .Q(sreg[163]) );
  DFF \sreg_reg[164]  ( .D(swire[38]), .CLK(clk), .RST(rst), .Q(sreg[164]) );
  DFF \sreg_reg[165]  ( .D(swire[39]), .CLK(clk), .RST(rst), .Q(sreg[165]) );
  DFF \sreg_reg[166]  ( .D(swire[40]), .CLK(clk), .RST(rst), .Q(sreg[166]) );
  DFF \sreg_reg[167]  ( .D(swire[41]), .CLK(clk), .RST(rst), .Q(sreg[167]) );
  DFF \sreg_reg[168]  ( .D(swire[42]), .CLK(clk), .RST(rst), .Q(sreg[168]) );
  DFF \sreg_reg[169]  ( .D(swire[43]), .CLK(clk), .RST(rst), .Q(sreg[169]) );
  DFF \sreg_reg[170]  ( .D(swire[44]), .CLK(clk), .RST(rst), .Q(sreg[170]) );
  DFF \sreg_reg[171]  ( .D(swire[45]), .CLK(clk), .RST(rst), .Q(sreg[171]) );
  DFF \sreg_reg[172]  ( .D(swire[46]), .CLK(clk), .RST(rst), .Q(sreg[172]) );
  DFF \sreg_reg[173]  ( .D(swire[47]), .CLK(clk), .RST(rst), .Q(sreg[173]) );
  DFF \sreg_reg[174]  ( .D(swire[48]), .CLK(clk), .RST(rst), .Q(sreg[174]) );
  DFF \sreg_reg[175]  ( .D(swire[49]), .CLK(clk), .RST(rst), .Q(sreg[175]) );
  DFF \sreg_reg[176]  ( .D(swire[50]), .CLK(clk), .RST(rst), .Q(sreg[176]) );
  DFF \sreg_reg[177]  ( .D(swire[51]), .CLK(clk), .RST(rst), .Q(sreg[177]) );
  DFF \sreg_reg[178]  ( .D(swire[52]), .CLK(clk), .RST(rst), .Q(sreg[178]) );
  DFF \sreg_reg[179]  ( .D(swire[53]), .CLK(clk), .RST(rst), .Q(sreg[179]) );
  DFF \sreg_reg[180]  ( .D(swire[54]), .CLK(clk), .RST(rst), .Q(sreg[180]) );
  DFF \sreg_reg[181]  ( .D(swire[55]), .CLK(clk), .RST(rst), .Q(sreg[181]) );
  DFF \sreg_reg[182]  ( .D(swire[56]), .CLK(clk), .RST(rst), .Q(sreg[182]) );
  DFF \sreg_reg[183]  ( .D(swire[57]), .CLK(clk), .RST(rst), .Q(sreg[183]) );
  DFF \sreg_reg[184]  ( .D(swire[58]), .CLK(clk), .RST(rst), .Q(sreg[184]) );
  DFF \sreg_reg[185]  ( .D(swire[59]), .CLK(clk), .RST(rst), .Q(sreg[185]) );
  DFF \sreg_reg[186]  ( .D(swire[60]), .CLK(clk), .RST(rst), .Q(sreg[186]) );
  DFF \sreg_reg[187]  ( .D(swire[61]), .CLK(clk), .RST(rst), .Q(sreg[187]) );
  DFF \sreg_reg[188]  ( .D(swire[62]), .CLK(clk), .RST(rst), .Q(sreg[188]) );
  DFF \sreg_reg[189]  ( .D(swire[63]), .CLK(clk), .RST(rst), .Q(sreg[189]) );
  DFF \sreg_reg[190]  ( .D(swire[64]), .CLK(clk), .RST(rst), .Q(sreg[190]) );
  DFF \sreg_reg[191]  ( .D(swire[65]), .CLK(clk), .RST(rst), .Q(sreg[191]) );
  DFF \sreg_reg[192]  ( .D(swire[66]), .CLK(clk), .RST(rst), .Q(sreg[192]) );
  DFF \sreg_reg[193]  ( .D(swire[67]), .CLK(clk), .RST(rst), .Q(sreg[193]) );
  DFF \sreg_reg[194]  ( .D(swire[68]), .CLK(clk), .RST(rst), .Q(sreg[194]) );
  DFF \sreg_reg[195]  ( .D(swire[69]), .CLK(clk), .RST(rst), .Q(sreg[195]) );
  DFF \sreg_reg[196]  ( .D(swire[70]), .CLK(clk), .RST(rst), .Q(sreg[196]) );
  DFF \sreg_reg[197]  ( .D(swire[71]), .CLK(clk), .RST(rst), .Q(sreg[197]) );
  DFF \sreg_reg[198]  ( .D(swire[72]), .CLK(clk), .RST(rst), .Q(sreg[198]) );
  DFF \sreg_reg[199]  ( .D(swire[73]), .CLK(clk), .RST(rst), .Q(sreg[199]) );
  DFF \sreg_reg[200]  ( .D(swire[74]), .CLK(clk), .RST(rst), .Q(sreg[200]) );
  DFF \sreg_reg[201]  ( .D(swire[75]), .CLK(clk), .RST(rst), .Q(sreg[201]) );
  DFF \sreg_reg[202]  ( .D(swire[76]), .CLK(clk), .RST(rst), .Q(sreg[202]) );
  DFF \sreg_reg[203]  ( .D(swire[77]), .CLK(clk), .RST(rst), .Q(sreg[203]) );
  DFF \sreg_reg[204]  ( .D(swire[78]), .CLK(clk), .RST(rst), .Q(sreg[204]) );
  DFF \sreg_reg[205]  ( .D(swire[79]), .CLK(clk), .RST(rst), .Q(sreg[205]) );
  DFF \sreg_reg[206]  ( .D(swire[80]), .CLK(clk), .RST(rst), .Q(sreg[206]) );
  DFF \sreg_reg[207]  ( .D(swire[81]), .CLK(clk), .RST(rst), .Q(sreg[207]) );
  DFF \sreg_reg[208]  ( .D(swire[82]), .CLK(clk), .RST(rst), .Q(sreg[208]) );
  DFF \sreg_reg[209]  ( .D(swire[83]), .CLK(clk), .RST(rst), .Q(sreg[209]) );
  DFF \sreg_reg[210]  ( .D(swire[84]), .CLK(clk), .RST(rst), .Q(sreg[210]) );
  DFF \sreg_reg[211]  ( .D(swire[85]), .CLK(clk), .RST(rst), .Q(sreg[211]) );
  DFF \sreg_reg[212]  ( .D(swire[86]), .CLK(clk), .RST(rst), .Q(sreg[212]) );
  DFF \sreg_reg[213]  ( .D(swire[87]), .CLK(clk), .RST(rst), .Q(sreg[213]) );
  DFF \sreg_reg[214]  ( .D(swire[88]), .CLK(clk), .RST(rst), .Q(sreg[214]) );
  DFF \sreg_reg[215]  ( .D(swire[89]), .CLK(clk), .RST(rst), .Q(sreg[215]) );
  DFF \sreg_reg[216]  ( .D(swire[90]), .CLK(clk), .RST(rst), .Q(sreg[216]) );
  DFF \sreg_reg[217]  ( .D(swire[91]), .CLK(clk), .RST(rst), .Q(sreg[217]) );
  DFF \sreg_reg[218]  ( .D(swire[92]), .CLK(clk), .RST(rst), .Q(sreg[218]) );
  DFF \sreg_reg[219]  ( .D(swire[93]), .CLK(clk), .RST(rst), .Q(sreg[219]) );
  DFF \sreg_reg[220]  ( .D(swire[94]), .CLK(clk), .RST(rst), .Q(sreg[220]) );
  DFF \sreg_reg[221]  ( .D(swire[95]), .CLK(clk), .RST(rst), .Q(sreg[221]) );
  DFF \sreg_reg[222]  ( .D(swire[96]), .CLK(clk), .RST(rst), .Q(sreg[222]) );
  DFF \sreg_reg[223]  ( .D(swire[97]), .CLK(clk), .RST(rst), .Q(sreg[223]) );
  DFF \sreg_reg[224]  ( .D(swire[98]), .CLK(clk), .RST(rst), .Q(sreg[224]) );
  DFF \sreg_reg[225]  ( .D(swire[99]), .CLK(clk), .RST(rst), .Q(sreg[225]) );
  DFF \sreg_reg[226]  ( .D(swire[100]), .CLK(clk), .RST(rst), .Q(sreg[226]) );
  DFF \sreg_reg[227]  ( .D(swire[101]), .CLK(clk), .RST(rst), .Q(sreg[227]) );
  DFF \sreg_reg[228]  ( .D(swire[102]), .CLK(clk), .RST(rst), .Q(sreg[228]) );
  DFF \sreg_reg[229]  ( .D(swire[103]), .CLK(clk), .RST(rst), .Q(sreg[229]) );
  DFF \sreg_reg[230]  ( .D(swire[104]), .CLK(clk), .RST(rst), .Q(sreg[230]) );
  DFF \sreg_reg[231]  ( .D(swire[105]), .CLK(clk), .RST(rst), .Q(sreg[231]) );
  DFF \sreg_reg[232]  ( .D(swire[106]), .CLK(clk), .RST(rst), .Q(sreg[232]) );
  DFF \sreg_reg[233]  ( .D(swire[107]), .CLK(clk), .RST(rst), .Q(sreg[233]) );
  DFF \sreg_reg[234]  ( .D(swire[108]), .CLK(clk), .RST(rst), .Q(sreg[234]) );
  DFF \sreg_reg[235]  ( .D(swire[109]), .CLK(clk), .RST(rst), .Q(sreg[235]) );
  DFF \sreg_reg[236]  ( .D(swire[110]), .CLK(clk), .RST(rst), .Q(sreg[236]) );
  DFF \sreg_reg[237]  ( .D(swire[111]), .CLK(clk), .RST(rst), .Q(sreg[237]) );
  DFF \sreg_reg[238]  ( .D(swire[112]), .CLK(clk), .RST(rst), .Q(sreg[238]) );
  DFF \sreg_reg[239]  ( .D(swire[113]), .CLK(clk), .RST(rst), .Q(sreg[239]) );
  DFF \sreg_reg[240]  ( .D(swire[114]), .CLK(clk), .RST(rst), .Q(sreg[240]) );
  DFF \sreg_reg[241]  ( .D(swire[115]), .CLK(clk), .RST(rst), .Q(sreg[241]) );
  DFF \sreg_reg[242]  ( .D(swire[116]), .CLK(clk), .RST(rst), .Q(sreg[242]) );
  DFF \sreg_reg[243]  ( .D(swire[117]), .CLK(clk), .RST(rst), .Q(sreg[243]) );
  DFF \sreg_reg[244]  ( .D(swire[118]), .CLK(clk), .RST(rst), .Q(sreg[244]) );
  DFF \sreg_reg[245]  ( .D(swire[119]), .CLK(clk), .RST(rst), .Q(sreg[245]) );
  DFF \sreg_reg[246]  ( .D(swire[120]), .CLK(clk), .RST(rst), .Q(sreg[246]) );
  DFF \sreg_reg[247]  ( .D(swire[121]), .CLK(clk), .RST(rst), .Q(sreg[247]) );
  DFF \sreg_reg[248]  ( .D(swire[122]), .CLK(clk), .RST(rst), .Q(sreg[248]) );
  DFF \sreg_reg[249]  ( .D(swire[123]), .CLK(clk), .RST(rst), .Q(sreg[249]) );
  DFF \sreg_reg[250]  ( .D(swire[124]), .CLK(clk), .RST(rst), .Q(sreg[250]) );
  DFF \sreg_reg[251]  ( .D(swire[125]), .CLK(clk), .RST(rst), .Q(sreg[251]) );
  DFF \sreg_reg[252]  ( .D(swire[126]), .CLK(clk), .RST(rst), .Q(sreg[252]) );
  DFF \sreg_reg[253]  ( .D(swire[127]), .CLK(clk), .RST(rst), .Q(sreg[253]) );
  DFF \sreg_reg[127]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[125]) );
  DFF \sreg_reg[126]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[124]) );
  DFF \sreg_reg[125]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[123]) );
  DFF \sreg_reg[124]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[122]) );
  DFF \sreg_reg[123]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[121]) );
  DFF \sreg_reg[122]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[120]) );
  DFF \sreg_reg[121]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[120]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[119]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[118]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[117]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[116]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[115]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[114]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[113]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[112]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[111]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[110]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[109]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[108]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[107]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[106]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[105]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[104]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[103]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[102]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[101]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[100]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[99]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[98]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[97]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[96]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[95]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[94]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[93]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[92]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[91]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[90]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[89]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[88]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[87]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[86]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[85]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[84]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[83]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[82]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[81]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[80]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[79]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[78]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[77]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[76]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[75]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[74]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[73]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[72]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[71]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[70]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[69]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[68]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[67]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[66]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[65]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[64]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[63]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[62]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[61]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[60]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[59]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[58]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[57]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[56]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[55]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[54]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[53]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[52]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[51]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[50]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[49]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[48]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[47]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[46]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[45]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[44]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[43]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[42]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[41]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[40]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[39]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[38]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[37]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[36]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[35]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[34]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[33]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[32]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[31]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[30]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[29]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[28]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[27]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[26]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[25]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[24]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[23]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[22]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[21]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[20]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[19]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[18]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[17]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[16]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[15]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[14]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[13]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[12]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[11]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[10]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[9]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[8]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[7]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[6]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[5]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[4]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[3]  ( .D(c[3]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[2]  ( .D(c[2]), .CLK(clk), .RST(rst), .Q(c[0]) );
  XNOR U5 ( .A(n1), .B(n2), .Z(swire[9]) );
  XNOR U6 ( .A(n3), .B(n4), .Z(swire[99]) );
  XNOR U7 ( .A(n5), .B(n6), .Z(swire[98]) );
  XNOR U8 ( .A(n7), .B(n8), .Z(swire[97]) );
  XNOR U9 ( .A(n9), .B(n10), .Z(swire[96]) );
  XNOR U10 ( .A(n11), .B(n12), .Z(swire[95]) );
  XNOR U11 ( .A(n13), .B(n14), .Z(swire[94]) );
  XNOR U12 ( .A(n15), .B(n16), .Z(swire[93]) );
  XNOR U13 ( .A(n17), .B(n18), .Z(swire[92]) );
  XNOR U14 ( .A(n19), .B(n20), .Z(swire[91]) );
  XNOR U15 ( .A(n21), .B(n22), .Z(swire[90]) );
  XNOR U16 ( .A(n23), .B(n24), .Z(swire[8]) );
  XNOR U17 ( .A(n25), .B(n26), .Z(swire[89]) );
  XNOR U18 ( .A(n27), .B(n28), .Z(swire[88]) );
  XNOR U19 ( .A(n29), .B(n30), .Z(swire[87]) );
  XNOR U20 ( .A(n31), .B(n32), .Z(swire[86]) );
  XNOR U21 ( .A(n33), .B(n34), .Z(swire[85]) );
  XNOR U22 ( .A(n35), .B(n36), .Z(swire[84]) );
  XNOR U23 ( .A(n37), .B(n38), .Z(swire[83]) );
  XNOR U24 ( .A(n39), .B(n40), .Z(swire[82]) );
  XNOR U25 ( .A(n41), .B(n42), .Z(swire[81]) );
  XNOR U26 ( .A(n43), .B(n44), .Z(swire[80]) );
  XNOR U27 ( .A(n45), .B(n46), .Z(swire[7]) );
  XNOR U28 ( .A(n47), .B(n48), .Z(swire[79]) );
  XNOR U29 ( .A(n49), .B(n50), .Z(swire[78]) );
  XNOR U30 ( .A(n51), .B(n52), .Z(swire[77]) );
  XNOR U31 ( .A(n53), .B(n54), .Z(swire[76]) );
  XNOR U32 ( .A(n55), .B(n56), .Z(swire[75]) );
  XNOR U33 ( .A(n57), .B(n58), .Z(swire[74]) );
  XNOR U34 ( .A(n59), .B(n60), .Z(swire[73]) );
  XNOR U35 ( .A(n61), .B(n62), .Z(swire[72]) );
  XNOR U36 ( .A(n63), .B(n64), .Z(swire[71]) );
  XNOR U37 ( .A(n65), .B(n66), .Z(swire[70]) );
  XNOR U38 ( .A(n67), .B(n68), .Z(swire[6]) );
  XNOR U39 ( .A(n69), .B(n70), .Z(swire[69]) );
  XNOR U40 ( .A(n71), .B(n72), .Z(swire[68]) );
  XNOR U41 ( .A(n73), .B(n74), .Z(swire[67]) );
  XNOR U42 ( .A(n75), .B(n76), .Z(swire[66]) );
  XNOR U43 ( .A(n77), .B(n78), .Z(swire[65]) );
  XNOR U44 ( .A(n79), .B(n80), .Z(swire[64]) );
  XNOR U45 ( .A(n81), .B(n82), .Z(swire[63]) );
  XNOR U46 ( .A(n83), .B(n84), .Z(swire[62]) );
  XNOR U47 ( .A(n85), .B(n86), .Z(swire[61]) );
  XNOR U48 ( .A(n87), .B(n88), .Z(swire[60]) );
  XNOR U49 ( .A(n89), .B(n90), .Z(swire[5]) );
  XNOR U50 ( .A(n91), .B(n92), .Z(swire[59]) );
  XNOR U51 ( .A(n93), .B(n94), .Z(swire[58]) );
  XNOR U52 ( .A(n95), .B(n96), .Z(swire[57]) );
  XNOR U53 ( .A(n97), .B(n98), .Z(swire[56]) );
  XNOR U54 ( .A(n99), .B(n100), .Z(swire[55]) );
  XNOR U55 ( .A(n101), .B(n102), .Z(swire[54]) );
  XNOR U56 ( .A(n103), .B(n104), .Z(swire[53]) );
  XNOR U57 ( .A(n105), .B(n106), .Z(swire[52]) );
  XNOR U58 ( .A(n107), .B(n108), .Z(swire[51]) );
  XNOR U59 ( .A(n109), .B(n110), .Z(swire[50]) );
  XNOR U60 ( .A(n111), .B(n112), .Z(swire[4]) );
  XNOR U61 ( .A(n113), .B(n114), .Z(swire[49]) );
  XNOR U62 ( .A(n115), .B(n116), .Z(swire[48]) );
  XNOR U63 ( .A(n117), .B(n118), .Z(swire[47]) );
  XNOR U64 ( .A(n119), .B(n120), .Z(swire[46]) );
  XNOR U65 ( .A(n121), .B(n122), .Z(swire[45]) );
  XNOR U66 ( .A(n123), .B(n124), .Z(swire[44]) );
  XNOR U67 ( .A(n125), .B(n126), .Z(swire[43]) );
  XNOR U68 ( .A(n127), .B(n128), .Z(swire[42]) );
  XNOR U69 ( .A(n129), .B(n130), .Z(swire[41]) );
  XNOR U70 ( .A(n131), .B(n132), .Z(swire[40]) );
  XNOR U71 ( .A(n133), .B(n134), .Z(swire[3]) );
  XNOR U72 ( .A(n135), .B(n136), .Z(swire[39]) );
  XNOR U73 ( .A(n137), .B(n138), .Z(swire[38]) );
  XNOR U74 ( .A(n139), .B(n140), .Z(swire[37]) );
  XNOR U75 ( .A(n141), .B(n142), .Z(swire[36]) );
  XNOR U76 ( .A(n143), .B(n144), .Z(swire[35]) );
  XNOR U77 ( .A(n145), .B(n146), .Z(swire[34]) );
  XNOR U78 ( .A(n147), .B(n148), .Z(swire[33]) );
  XNOR U79 ( .A(n149), .B(n150), .Z(swire[32]) );
  XNOR U80 ( .A(n151), .B(n152), .Z(swire[31]) );
  XNOR U81 ( .A(n153), .B(n154), .Z(swire[30]) );
  XNOR U82 ( .A(n155), .B(n156), .Z(swire[2]) );
  XNOR U83 ( .A(n157), .B(n158), .Z(swire[29]) );
  XNOR U84 ( .A(n159), .B(n160), .Z(swire[28]) );
  XNOR U85 ( .A(n161), .B(n162), .Z(swire[27]) );
  XNOR U86 ( .A(n163), .B(n164), .Z(swire[26]) );
  XNOR U87 ( .A(n165), .B(n166), .Z(swire[25]) );
  XNOR U88 ( .A(n167), .B(n168), .Z(swire[24]) );
  XNOR U89 ( .A(n169), .B(n170), .Z(swire[23]) );
  XNOR U90 ( .A(n171), .B(n172), .Z(swire[22]) );
  XNOR U91 ( .A(n173), .B(n174), .Z(swire[21]) );
  XNOR U92 ( .A(n175), .B(n176), .Z(swire[20]) );
  XNOR U93 ( .A(n177), .B(n178), .Z(swire[19]) );
  XNOR U94 ( .A(n179), .B(n180), .Z(swire[18]) );
  XNOR U95 ( .A(n181), .B(n182), .Z(swire[17]) );
  XNOR U96 ( .A(n183), .B(n184), .Z(swire[16]) );
  XNOR U97 ( .A(n185), .B(n186), .Z(swire[15]) );
  XNOR U98 ( .A(n187), .B(n188), .Z(swire[14]) );
  XNOR U99 ( .A(n189), .B(n190), .Z(swire[13]) );
  XNOR U100 ( .A(n191), .B(n192), .Z(swire[12]) );
  XOR U101 ( .A(n193), .B(n194), .Z(swire[127]) );
  AND U102 ( .A(a[127]), .B(b[0]), .Z(n194) );
  AND U103 ( .A(b[1]), .B(a[126]), .Z(n193) );
  XOR U104 ( .A(n195), .B(n196), .Z(swire[126]) );
  AND U105 ( .A(a[126]), .B(b[0]), .Z(n196) );
  AND U106 ( .A(b[1]), .B(a[125]), .Z(n195) );
  XOR U107 ( .A(n197), .B(n198), .Z(swire[125]) );
  XOR U108 ( .A(sreg[253]), .B(n199), .Z(n198) );
  AND U109 ( .A(b[1]), .B(a[124]), .Z(n199) );
  AND U110 ( .A(a[125]), .B(b[0]), .Z(n197) );
  XOR U111 ( .A(n200), .B(n201), .Z(swire[124]) );
  XOR U112 ( .A(sreg[252]), .B(n202), .Z(n201) );
  AND U113 ( .A(b[1]), .B(a[123]), .Z(n202) );
  AND U114 ( .A(a[124]), .B(b[0]), .Z(n200) );
  XOR U115 ( .A(n203), .B(n204), .Z(swire[123]) );
  XOR U116 ( .A(sreg[251]), .B(n205), .Z(n204) );
  XOR U117 ( .A(n205), .B(n206), .Z(n203) );
  XOR U118 ( .A(n207), .B(n208), .Z(n206) );
  AND U119 ( .A(a[123]), .B(b[0]), .Z(n208) );
  AND U120 ( .A(b[1]), .B(a[122]), .Z(n207) );
  XOR U121 ( .A(n209), .B(n210), .Z(n205) );
  ANDN U122 ( .B(n211), .A(n212), .Z(n209) );
  XNOR U123 ( .A(n211), .B(n212), .Z(swire[122]) );
  XOR U124 ( .A(sreg[250]), .B(n213), .Z(n212) );
  XOR U125 ( .A(n213), .B(n214), .Z(n211) );
  XOR U126 ( .A(n215), .B(n216), .Z(n214) );
  NAND U127 ( .A(b[0]), .B(a[122]), .Z(n216) );
  AND U128 ( .A(b[1]), .B(a[121]), .Z(n215) );
  IV U129 ( .A(n210), .Z(n213) );
  XOR U130 ( .A(n217), .B(n218), .Z(n210) );
  ANDN U131 ( .B(n219), .A(n220), .Z(n217) );
  XNOR U132 ( .A(n219), .B(n220), .Z(swire[121]) );
  XOR U133 ( .A(sreg[249]), .B(n221), .Z(n220) );
  XOR U134 ( .A(n221), .B(n222), .Z(n219) );
  XOR U135 ( .A(n223), .B(n224), .Z(n222) );
  NAND U136 ( .A(b[0]), .B(a[121]), .Z(n224) );
  AND U137 ( .A(b[1]), .B(a[120]), .Z(n223) );
  IV U138 ( .A(n218), .Z(n221) );
  XOR U139 ( .A(n225), .B(n226), .Z(n218) );
  ANDN U140 ( .B(n227), .A(n228), .Z(n225) );
  XNOR U141 ( .A(n227), .B(n228), .Z(swire[120]) );
  XOR U142 ( .A(sreg[248]), .B(n229), .Z(n228) );
  XOR U143 ( .A(n229), .B(n230), .Z(n227) );
  XOR U144 ( .A(n231), .B(n232), .Z(n230) );
  NAND U145 ( .A(b[0]), .B(a[120]), .Z(n232) );
  AND U146 ( .A(b[1]), .B(a[119]), .Z(n231) );
  IV U147 ( .A(n226), .Z(n229) );
  XOR U148 ( .A(n233), .B(n234), .Z(n226) );
  ANDN U149 ( .B(n235), .A(n236), .Z(n233) );
  XNOR U150 ( .A(n237), .B(n238), .Z(swire[11]) );
  XNOR U151 ( .A(n235), .B(n236), .Z(swire[119]) );
  XOR U152 ( .A(sreg[247]), .B(n239), .Z(n236) );
  XOR U153 ( .A(n239), .B(n240), .Z(n235) );
  XOR U154 ( .A(n241), .B(n242), .Z(n240) );
  NAND U155 ( .A(b[0]), .B(a[119]), .Z(n242) );
  AND U156 ( .A(b[1]), .B(a[118]), .Z(n241) );
  IV U157 ( .A(n234), .Z(n239) );
  XOR U158 ( .A(n243), .B(n244), .Z(n234) );
  ANDN U159 ( .B(n245), .A(n246), .Z(n243) );
  XNOR U160 ( .A(n245), .B(n246), .Z(swire[118]) );
  XOR U161 ( .A(sreg[246]), .B(n247), .Z(n246) );
  XOR U162 ( .A(n247), .B(n248), .Z(n245) );
  XOR U163 ( .A(n249), .B(n250), .Z(n248) );
  NAND U164 ( .A(b[0]), .B(a[118]), .Z(n250) );
  AND U165 ( .A(b[1]), .B(a[117]), .Z(n249) );
  IV U166 ( .A(n244), .Z(n247) );
  XOR U167 ( .A(n251), .B(n252), .Z(n244) );
  ANDN U168 ( .B(n253), .A(n254), .Z(n251) );
  XNOR U169 ( .A(n253), .B(n254), .Z(swire[117]) );
  XOR U170 ( .A(sreg[245]), .B(n255), .Z(n254) );
  XOR U171 ( .A(n255), .B(n256), .Z(n253) );
  XOR U172 ( .A(n257), .B(n258), .Z(n256) );
  NAND U173 ( .A(b[0]), .B(a[117]), .Z(n258) );
  AND U174 ( .A(b[1]), .B(a[116]), .Z(n257) );
  IV U175 ( .A(n252), .Z(n255) );
  XOR U176 ( .A(n259), .B(n260), .Z(n252) );
  ANDN U177 ( .B(n261), .A(n262), .Z(n259) );
  XNOR U178 ( .A(n261), .B(n262), .Z(swire[116]) );
  XOR U179 ( .A(sreg[244]), .B(n263), .Z(n262) );
  XOR U180 ( .A(n263), .B(n264), .Z(n261) );
  XOR U181 ( .A(n265), .B(n266), .Z(n264) );
  NAND U182 ( .A(b[0]), .B(a[116]), .Z(n266) );
  AND U183 ( .A(b[1]), .B(a[115]), .Z(n265) );
  IV U184 ( .A(n260), .Z(n263) );
  XOR U185 ( .A(n267), .B(n268), .Z(n260) );
  ANDN U186 ( .B(n269), .A(n270), .Z(n267) );
  XNOR U187 ( .A(n269), .B(n270), .Z(swire[115]) );
  XOR U188 ( .A(sreg[243]), .B(n271), .Z(n270) );
  XOR U189 ( .A(n271), .B(n272), .Z(n269) );
  XOR U190 ( .A(n273), .B(n274), .Z(n272) );
  NAND U191 ( .A(b[0]), .B(a[115]), .Z(n274) );
  AND U192 ( .A(b[1]), .B(a[114]), .Z(n273) );
  IV U193 ( .A(n268), .Z(n271) );
  XOR U194 ( .A(n275), .B(n276), .Z(n268) );
  ANDN U195 ( .B(n277), .A(n278), .Z(n275) );
  XNOR U196 ( .A(n277), .B(n278), .Z(swire[114]) );
  XOR U197 ( .A(sreg[242]), .B(n279), .Z(n278) );
  XOR U198 ( .A(n279), .B(n280), .Z(n277) );
  XOR U199 ( .A(n281), .B(n282), .Z(n280) );
  NAND U200 ( .A(b[0]), .B(a[114]), .Z(n282) );
  AND U201 ( .A(b[1]), .B(a[113]), .Z(n281) );
  IV U202 ( .A(n276), .Z(n279) );
  XOR U203 ( .A(n283), .B(n284), .Z(n276) );
  ANDN U204 ( .B(n285), .A(n286), .Z(n283) );
  XNOR U205 ( .A(n285), .B(n286), .Z(swire[113]) );
  XOR U206 ( .A(sreg[241]), .B(n287), .Z(n286) );
  XOR U207 ( .A(n287), .B(n288), .Z(n285) );
  XOR U208 ( .A(n289), .B(n290), .Z(n288) );
  NAND U209 ( .A(b[0]), .B(a[113]), .Z(n290) );
  AND U210 ( .A(b[1]), .B(a[112]), .Z(n289) );
  IV U211 ( .A(n284), .Z(n287) );
  XOR U212 ( .A(n291), .B(n292), .Z(n284) );
  ANDN U213 ( .B(n293), .A(n294), .Z(n291) );
  XNOR U214 ( .A(n293), .B(n294), .Z(swire[112]) );
  XOR U215 ( .A(sreg[240]), .B(n295), .Z(n294) );
  XOR U216 ( .A(n295), .B(n296), .Z(n293) );
  XOR U217 ( .A(n297), .B(n298), .Z(n296) );
  NAND U218 ( .A(b[0]), .B(a[112]), .Z(n298) );
  AND U219 ( .A(b[1]), .B(a[111]), .Z(n297) );
  IV U220 ( .A(n292), .Z(n295) );
  XOR U221 ( .A(n299), .B(n300), .Z(n292) );
  ANDN U222 ( .B(n301), .A(n302), .Z(n299) );
  XNOR U223 ( .A(n301), .B(n302), .Z(swire[111]) );
  XOR U224 ( .A(sreg[239]), .B(n303), .Z(n302) );
  XOR U225 ( .A(n303), .B(n304), .Z(n301) );
  XOR U226 ( .A(n305), .B(n306), .Z(n304) );
  NAND U227 ( .A(b[0]), .B(a[111]), .Z(n306) );
  AND U228 ( .A(b[1]), .B(a[110]), .Z(n305) );
  IV U229 ( .A(n300), .Z(n303) );
  XOR U230 ( .A(n307), .B(n308), .Z(n300) );
  ANDN U231 ( .B(n309), .A(n310), .Z(n307) );
  XNOR U232 ( .A(n309), .B(n310), .Z(swire[110]) );
  XOR U233 ( .A(sreg[238]), .B(n311), .Z(n310) );
  XOR U234 ( .A(n311), .B(n312), .Z(n309) );
  XOR U235 ( .A(n313), .B(n314), .Z(n312) );
  NAND U236 ( .A(b[0]), .B(a[110]), .Z(n314) );
  AND U237 ( .A(b[1]), .B(a[109]), .Z(n313) );
  IV U238 ( .A(n308), .Z(n311) );
  XOR U239 ( .A(n315), .B(n316), .Z(n308) );
  ANDN U240 ( .B(n317), .A(n318), .Z(n315) );
  XNOR U241 ( .A(n319), .B(n320), .Z(swire[10]) );
  XNOR U242 ( .A(n317), .B(n318), .Z(swire[109]) );
  XOR U243 ( .A(sreg[237]), .B(n321), .Z(n318) );
  XOR U244 ( .A(n321), .B(n322), .Z(n317) );
  XOR U245 ( .A(n323), .B(n324), .Z(n322) );
  NAND U246 ( .A(b[0]), .B(a[109]), .Z(n324) );
  AND U247 ( .A(b[1]), .B(a[108]), .Z(n323) );
  IV U248 ( .A(n316), .Z(n321) );
  XOR U249 ( .A(n325), .B(n326), .Z(n316) );
  ANDN U250 ( .B(n327), .A(n328), .Z(n325) );
  XNOR U251 ( .A(n327), .B(n328), .Z(swire[108]) );
  XOR U252 ( .A(sreg[236]), .B(n329), .Z(n328) );
  XOR U253 ( .A(n329), .B(n330), .Z(n327) );
  XOR U254 ( .A(n331), .B(n332), .Z(n330) );
  NAND U255 ( .A(b[0]), .B(a[108]), .Z(n332) );
  AND U256 ( .A(b[1]), .B(a[107]), .Z(n331) );
  IV U257 ( .A(n326), .Z(n329) );
  XOR U258 ( .A(n333), .B(n334), .Z(n326) );
  ANDN U259 ( .B(n335), .A(n336), .Z(n333) );
  XNOR U260 ( .A(n335), .B(n336), .Z(swire[107]) );
  XOR U261 ( .A(sreg[235]), .B(n337), .Z(n336) );
  XOR U262 ( .A(n337), .B(n338), .Z(n335) );
  XOR U263 ( .A(n339), .B(n340), .Z(n338) );
  NAND U264 ( .A(b[0]), .B(a[107]), .Z(n340) );
  AND U265 ( .A(b[1]), .B(a[106]), .Z(n339) );
  IV U266 ( .A(n334), .Z(n337) );
  XOR U267 ( .A(n341), .B(n342), .Z(n334) );
  ANDN U268 ( .B(n343), .A(n344), .Z(n341) );
  XNOR U269 ( .A(n343), .B(n344), .Z(swire[106]) );
  XOR U270 ( .A(sreg[234]), .B(n345), .Z(n344) );
  XOR U271 ( .A(n345), .B(n346), .Z(n343) );
  XOR U272 ( .A(n347), .B(n348), .Z(n346) );
  NAND U273 ( .A(b[0]), .B(a[106]), .Z(n348) );
  AND U274 ( .A(b[1]), .B(a[105]), .Z(n347) );
  IV U275 ( .A(n342), .Z(n345) );
  XOR U276 ( .A(n349), .B(n350), .Z(n342) );
  ANDN U277 ( .B(n351), .A(n352), .Z(n349) );
  XNOR U278 ( .A(n351), .B(n352), .Z(swire[105]) );
  XOR U279 ( .A(sreg[233]), .B(n353), .Z(n352) );
  XOR U280 ( .A(n353), .B(n354), .Z(n351) );
  XOR U281 ( .A(n355), .B(n356), .Z(n354) );
  NAND U282 ( .A(b[0]), .B(a[105]), .Z(n356) );
  AND U283 ( .A(b[1]), .B(a[104]), .Z(n355) );
  IV U284 ( .A(n350), .Z(n353) );
  XOR U285 ( .A(n357), .B(n358), .Z(n350) );
  ANDN U286 ( .B(n359), .A(n360), .Z(n357) );
  XNOR U287 ( .A(n359), .B(n360), .Z(swire[104]) );
  XOR U288 ( .A(sreg[232]), .B(n361), .Z(n360) );
  XOR U289 ( .A(n361), .B(n362), .Z(n359) );
  XOR U290 ( .A(n363), .B(n364), .Z(n362) );
  NAND U291 ( .A(b[0]), .B(a[104]), .Z(n364) );
  AND U292 ( .A(b[1]), .B(a[103]), .Z(n363) );
  IV U293 ( .A(n358), .Z(n361) );
  XOR U294 ( .A(n365), .B(n366), .Z(n358) );
  ANDN U295 ( .B(n367), .A(n368), .Z(n365) );
  XNOR U296 ( .A(n367), .B(n368), .Z(swire[103]) );
  XOR U297 ( .A(sreg[231]), .B(n369), .Z(n368) );
  XOR U298 ( .A(n369), .B(n370), .Z(n367) );
  XOR U299 ( .A(n371), .B(n372), .Z(n370) );
  NAND U300 ( .A(b[0]), .B(a[103]), .Z(n372) );
  AND U301 ( .A(b[1]), .B(a[102]), .Z(n371) );
  IV U302 ( .A(n366), .Z(n369) );
  XOR U303 ( .A(n373), .B(n374), .Z(n366) );
  ANDN U304 ( .B(n375), .A(n376), .Z(n373) );
  XNOR U305 ( .A(n375), .B(n376), .Z(swire[102]) );
  XOR U306 ( .A(sreg[230]), .B(n377), .Z(n376) );
  XOR U307 ( .A(n377), .B(n378), .Z(n375) );
  XOR U308 ( .A(n379), .B(n380), .Z(n378) );
  NAND U309 ( .A(b[0]), .B(a[102]), .Z(n380) );
  AND U310 ( .A(b[1]), .B(a[101]), .Z(n379) );
  IV U311 ( .A(n374), .Z(n377) );
  XOR U312 ( .A(n381), .B(n382), .Z(n374) );
  ANDN U313 ( .B(n383), .A(n384), .Z(n381) );
  XNOR U314 ( .A(n383), .B(n384), .Z(swire[101]) );
  XOR U315 ( .A(sreg[229]), .B(n385), .Z(n384) );
  XOR U316 ( .A(n385), .B(n386), .Z(n383) );
  XOR U317 ( .A(n387), .B(n388), .Z(n386) );
  NAND U318 ( .A(b[0]), .B(a[101]), .Z(n388) );
  AND U319 ( .A(b[1]), .B(a[100]), .Z(n387) );
  IV U320 ( .A(n382), .Z(n385) );
  XOR U321 ( .A(n389), .B(n390), .Z(n382) );
  ANDN U322 ( .B(n391), .A(n392), .Z(n389) );
  XNOR U323 ( .A(n391), .B(n392), .Z(swire[100]) );
  XOR U324 ( .A(sreg[228]), .B(n393), .Z(n392) );
  XOR U325 ( .A(n393), .B(n394), .Z(n391) );
  XOR U326 ( .A(n395), .B(n396), .Z(n394) );
  NAND U327 ( .A(b[0]), .B(a[100]), .Z(n396) );
  AND U328 ( .A(a[99]), .B(b[1]), .Z(n395) );
  IV U329 ( .A(n390), .Z(n393) );
  XOR U330 ( .A(n397), .B(n398), .Z(n390) );
  ANDN U331 ( .B(n4), .A(n3), .Z(n397) );
  XOR U332 ( .A(sreg[227]), .B(n399), .Z(n3) );
  XOR U333 ( .A(n399), .B(n400), .Z(n4) );
  XOR U334 ( .A(n401), .B(n402), .Z(n400) );
  NAND U335 ( .A(b[1]), .B(a[98]), .Z(n402) );
  AND U336 ( .A(b[0]), .B(a[99]), .Z(n401) );
  IV U337 ( .A(n398), .Z(n399) );
  XOR U338 ( .A(n403), .B(n404), .Z(n398) );
  ANDN U339 ( .B(n5), .A(n6), .Z(n403) );
  XOR U340 ( .A(sreg[226]), .B(n405), .Z(n6) );
  XOR U341 ( .A(n405), .B(n406), .Z(n5) );
  XOR U342 ( .A(n407), .B(n408), .Z(n406) );
  NAND U343 ( .A(b[1]), .B(a[97]), .Z(n408) );
  AND U344 ( .A(b[0]), .B(a[98]), .Z(n407) );
  IV U345 ( .A(n404), .Z(n405) );
  XOR U346 ( .A(n409), .B(n410), .Z(n404) );
  ANDN U347 ( .B(n7), .A(n8), .Z(n409) );
  XOR U348 ( .A(sreg[225]), .B(n411), .Z(n8) );
  XOR U349 ( .A(n411), .B(n412), .Z(n7) );
  XOR U350 ( .A(n413), .B(n414), .Z(n412) );
  NAND U351 ( .A(b[1]), .B(a[96]), .Z(n414) );
  AND U352 ( .A(b[0]), .B(a[97]), .Z(n413) );
  IV U353 ( .A(n410), .Z(n411) );
  XOR U354 ( .A(n415), .B(n416), .Z(n410) );
  ANDN U355 ( .B(n9), .A(n10), .Z(n415) );
  XOR U356 ( .A(sreg[224]), .B(n417), .Z(n10) );
  XOR U357 ( .A(n417), .B(n418), .Z(n9) );
  XOR U358 ( .A(n419), .B(n420), .Z(n418) );
  NAND U359 ( .A(b[1]), .B(a[95]), .Z(n420) );
  AND U360 ( .A(b[0]), .B(a[96]), .Z(n419) );
  IV U361 ( .A(n416), .Z(n417) );
  XOR U362 ( .A(n421), .B(n422), .Z(n416) );
  ANDN U363 ( .B(n11), .A(n12), .Z(n421) );
  XOR U364 ( .A(sreg[223]), .B(n423), .Z(n12) );
  XOR U365 ( .A(n423), .B(n424), .Z(n11) );
  XOR U366 ( .A(n425), .B(n426), .Z(n424) );
  NAND U367 ( .A(b[1]), .B(a[94]), .Z(n426) );
  AND U368 ( .A(b[0]), .B(a[95]), .Z(n425) );
  IV U369 ( .A(n422), .Z(n423) );
  XOR U370 ( .A(n427), .B(n428), .Z(n422) );
  ANDN U371 ( .B(n13), .A(n14), .Z(n427) );
  XOR U372 ( .A(sreg[222]), .B(n429), .Z(n14) );
  XOR U373 ( .A(n429), .B(n430), .Z(n13) );
  XOR U374 ( .A(n431), .B(n432), .Z(n430) );
  NAND U375 ( .A(b[1]), .B(a[93]), .Z(n432) );
  AND U376 ( .A(b[0]), .B(a[94]), .Z(n431) );
  IV U377 ( .A(n428), .Z(n429) );
  XOR U378 ( .A(n433), .B(n434), .Z(n428) );
  ANDN U379 ( .B(n15), .A(n16), .Z(n433) );
  XOR U380 ( .A(sreg[221]), .B(n435), .Z(n16) );
  XOR U381 ( .A(n435), .B(n436), .Z(n15) );
  XOR U382 ( .A(n437), .B(n438), .Z(n436) );
  NAND U383 ( .A(b[1]), .B(a[92]), .Z(n438) );
  AND U384 ( .A(b[0]), .B(a[93]), .Z(n437) );
  IV U385 ( .A(n434), .Z(n435) );
  XOR U386 ( .A(n439), .B(n440), .Z(n434) );
  ANDN U387 ( .B(n17), .A(n18), .Z(n439) );
  XOR U388 ( .A(sreg[220]), .B(n441), .Z(n18) );
  XOR U389 ( .A(n441), .B(n442), .Z(n17) );
  XOR U390 ( .A(n443), .B(n444), .Z(n442) );
  NAND U391 ( .A(b[1]), .B(a[91]), .Z(n444) );
  AND U392 ( .A(b[0]), .B(a[92]), .Z(n443) );
  IV U393 ( .A(n440), .Z(n441) );
  XOR U394 ( .A(n445), .B(n446), .Z(n440) );
  ANDN U395 ( .B(n19), .A(n20), .Z(n445) );
  XOR U396 ( .A(sreg[219]), .B(n447), .Z(n20) );
  XOR U397 ( .A(n447), .B(n448), .Z(n19) );
  XOR U398 ( .A(n449), .B(n450), .Z(n448) );
  NAND U399 ( .A(b[1]), .B(a[90]), .Z(n450) );
  AND U400 ( .A(b[0]), .B(a[91]), .Z(n449) );
  IV U401 ( .A(n446), .Z(n447) );
  XOR U402 ( .A(n451), .B(n452), .Z(n446) );
  ANDN U403 ( .B(n21), .A(n22), .Z(n451) );
  XOR U404 ( .A(sreg[218]), .B(n453), .Z(n22) );
  XOR U405 ( .A(n453), .B(n454), .Z(n21) );
  XOR U406 ( .A(n455), .B(n456), .Z(n454) );
  NAND U407 ( .A(b[1]), .B(a[89]), .Z(n456) );
  AND U408 ( .A(b[0]), .B(a[90]), .Z(n455) );
  IV U409 ( .A(n452), .Z(n453) );
  XOR U410 ( .A(n457), .B(n458), .Z(n452) );
  ANDN U411 ( .B(n25), .A(n26), .Z(n457) );
  XOR U412 ( .A(sreg[217]), .B(n459), .Z(n26) );
  XOR U413 ( .A(n459), .B(n460), .Z(n25) );
  XOR U414 ( .A(n461), .B(n462), .Z(n460) );
  NAND U415 ( .A(b[1]), .B(a[88]), .Z(n462) );
  AND U416 ( .A(b[0]), .B(a[89]), .Z(n461) );
  IV U417 ( .A(n458), .Z(n459) );
  XOR U418 ( .A(n463), .B(n464), .Z(n458) );
  ANDN U419 ( .B(n27), .A(n28), .Z(n463) );
  XOR U420 ( .A(sreg[216]), .B(n465), .Z(n28) );
  XOR U421 ( .A(n465), .B(n466), .Z(n27) );
  XOR U422 ( .A(n467), .B(n468), .Z(n466) );
  NAND U423 ( .A(b[1]), .B(a[87]), .Z(n468) );
  AND U424 ( .A(b[0]), .B(a[88]), .Z(n467) );
  IV U425 ( .A(n464), .Z(n465) );
  XOR U426 ( .A(n469), .B(n470), .Z(n464) );
  ANDN U427 ( .B(n29), .A(n30), .Z(n469) );
  XOR U428 ( .A(sreg[215]), .B(n471), .Z(n30) );
  XOR U429 ( .A(n471), .B(n472), .Z(n29) );
  XOR U430 ( .A(n473), .B(n474), .Z(n472) );
  NAND U431 ( .A(b[1]), .B(a[86]), .Z(n474) );
  AND U432 ( .A(b[0]), .B(a[87]), .Z(n473) );
  IV U433 ( .A(n470), .Z(n471) );
  XOR U434 ( .A(n475), .B(n476), .Z(n470) );
  ANDN U435 ( .B(n31), .A(n32), .Z(n475) );
  XOR U436 ( .A(sreg[214]), .B(n477), .Z(n32) );
  XOR U437 ( .A(n477), .B(n478), .Z(n31) );
  XOR U438 ( .A(n479), .B(n480), .Z(n478) );
  NAND U439 ( .A(b[1]), .B(a[85]), .Z(n480) );
  AND U440 ( .A(b[0]), .B(a[86]), .Z(n479) );
  IV U441 ( .A(n476), .Z(n477) );
  XOR U442 ( .A(n481), .B(n482), .Z(n476) );
  ANDN U443 ( .B(n33), .A(n34), .Z(n481) );
  XOR U444 ( .A(sreg[213]), .B(n483), .Z(n34) );
  XOR U445 ( .A(n483), .B(n484), .Z(n33) );
  XOR U446 ( .A(n485), .B(n486), .Z(n484) );
  NAND U447 ( .A(b[1]), .B(a[84]), .Z(n486) );
  AND U448 ( .A(b[0]), .B(a[85]), .Z(n485) );
  IV U449 ( .A(n482), .Z(n483) );
  XOR U450 ( .A(n487), .B(n488), .Z(n482) );
  ANDN U451 ( .B(n35), .A(n36), .Z(n487) );
  XOR U452 ( .A(sreg[212]), .B(n489), .Z(n36) );
  XOR U453 ( .A(n489), .B(n490), .Z(n35) );
  XOR U454 ( .A(n491), .B(n492), .Z(n490) );
  NAND U455 ( .A(b[1]), .B(a[83]), .Z(n492) );
  AND U456 ( .A(b[0]), .B(a[84]), .Z(n491) );
  IV U457 ( .A(n488), .Z(n489) );
  XOR U458 ( .A(n493), .B(n494), .Z(n488) );
  ANDN U459 ( .B(n37), .A(n38), .Z(n493) );
  XOR U460 ( .A(sreg[211]), .B(n495), .Z(n38) );
  XOR U461 ( .A(n495), .B(n496), .Z(n37) );
  XOR U462 ( .A(n497), .B(n498), .Z(n496) );
  NAND U463 ( .A(b[1]), .B(a[82]), .Z(n498) );
  AND U464 ( .A(b[0]), .B(a[83]), .Z(n497) );
  IV U465 ( .A(n494), .Z(n495) );
  XOR U466 ( .A(n499), .B(n500), .Z(n494) );
  ANDN U467 ( .B(n39), .A(n40), .Z(n499) );
  XOR U468 ( .A(sreg[210]), .B(n501), .Z(n40) );
  XOR U469 ( .A(n501), .B(n502), .Z(n39) );
  XOR U470 ( .A(n503), .B(n504), .Z(n502) );
  NAND U471 ( .A(b[1]), .B(a[81]), .Z(n504) );
  AND U472 ( .A(b[0]), .B(a[82]), .Z(n503) );
  IV U473 ( .A(n500), .Z(n501) );
  XOR U474 ( .A(n505), .B(n506), .Z(n500) );
  ANDN U475 ( .B(n41), .A(n42), .Z(n505) );
  XOR U476 ( .A(sreg[209]), .B(n507), .Z(n42) );
  XOR U477 ( .A(n507), .B(n508), .Z(n41) );
  XOR U478 ( .A(n509), .B(n510), .Z(n508) );
  NAND U479 ( .A(b[1]), .B(a[80]), .Z(n510) );
  AND U480 ( .A(b[0]), .B(a[81]), .Z(n509) );
  IV U481 ( .A(n506), .Z(n507) );
  XOR U482 ( .A(n511), .B(n512), .Z(n506) );
  ANDN U483 ( .B(n43), .A(n44), .Z(n511) );
  XOR U484 ( .A(sreg[208]), .B(n513), .Z(n44) );
  XOR U485 ( .A(n513), .B(n514), .Z(n43) );
  XOR U486 ( .A(n515), .B(n516), .Z(n514) );
  NAND U487 ( .A(b[1]), .B(a[79]), .Z(n516) );
  AND U488 ( .A(b[0]), .B(a[80]), .Z(n515) );
  IV U489 ( .A(n512), .Z(n513) );
  XOR U490 ( .A(n517), .B(n518), .Z(n512) );
  ANDN U491 ( .B(n47), .A(n48), .Z(n517) );
  XOR U492 ( .A(sreg[207]), .B(n519), .Z(n48) );
  XOR U493 ( .A(n519), .B(n520), .Z(n47) );
  XOR U494 ( .A(n521), .B(n522), .Z(n520) );
  NAND U495 ( .A(b[1]), .B(a[78]), .Z(n522) );
  AND U496 ( .A(b[0]), .B(a[79]), .Z(n521) );
  IV U497 ( .A(n518), .Z(n519) );
  XOR U498 ( .A(n523), .B(n524), .Z(n518) );
  ANDN U499 ( .B(n49), .A(n50), .Z(n523) );
  XOR U500 ( .A(sreg[206]), .B(n525), .Z(n50) );
  XOR U501 ( .A(n525), .B(n526), .Z(n49) );
  XOR U502 ( .A(n527), .B(n528), .Z(n526) );
  NAND U503 ( .A(b[1]), .B(a[77]), .Z(n528) );
  AND U504 ( .A(b[0]), .B(a[78]), .Z(n527) );
  IV U505 ( .A(n524), .Z(n525) );
  XOR U506 ( .A(n529), .B(n530), .Z(n524) );
  ANDN U507 ( .B(n51), .A(n52), .Z(n529) );
  XOR U508 ( .A(sreg[205]), .B(n531), .Z(n52) );
  XOR U509 ( .A(n531), .B(n532), .Z(n51) );
  XOR U510 ( .A(n533), .B(n534), .Z(n532) );
  NAND U511 ( .A(b[1]), .B(a[76]), .Z(n534) );
  AND U512 ( .A(b[0]), .B(a[77]), .Z(n533) );
  IV U513 ( .A(n530), .Z(n531) );
  XOR U514 ( .A(n535), .B(n536), .Z(n530) );
  ANDN U515 ( .B(n53), .A(n54), .Z(n535) );
  XOR U516 ( .A(sreg[204]), .B(n537), .Z(n54) );
  XOR U517 ( .A(n537), .B(n538), .Z(n53) );
  XOR U518 ( .A(n539), .B(n540), .Z(n538) );
  NAND U519 ( .A(b[1]), .B(a[75]), .Z(n540) );
  AND U520 ( .A(b[0]), .B(a[76]), .Z(n539) );
  IV U521 ( .A(n536), .Z(n537) );
  XOR U522 ( .A(n541), .B(n542), .Z(n536) );
  ANDN U523 ( .B(n55), .A(n56), .Z(n541) );
  XOR U524 ( .A(sreg[203]), .B(n543), .Z(n56) );
  XOR U525 ( .A(n543), .B(n544), .Z(n55) );
  XOR U526 ( .A(n545), .B(n546), .Z(n544) );
  NAND U527 ( .A(b[1]), .B(a[74]), .Z(n546) );
  AND U528 ( .A(b[0]), .B(a[75]), .Z(n545) );
  IV U529 ( .A(n542), .Z(n543) );
  XOR U530 ( .A(n547), .B(n548), .Z(n542) );
  ANDN U531 ( .B(n57), .A(n58), .Z(n547) );
  XOR U532 ( .A(sreg[202]), .B(n549), .Z(n58) );
  XOR U533 ( .A(n549), .B(n550), .Z(n57) );
  XOR U534 ( .A(n551), .B(n552), .Z(n550) );
  NAND U535 ( .A(b[1]), .B(a[73]), .Z(n552) );
  AND U536 ( .A(b[0]), .B(a[74]), .Z(n551) );
  IV U537 ( .A(n548), .Z(n549) );
  XOR U538 ( .A(n553), .B(n554), .Z(n548) );
  ANDN U539 ( .B(n59), .A(n60), .Z(n553) );
  XOR U540 ( .A(sreg[201]), .B(n555), .Z(n60) );
  XOR U541 ( .A(n555), .B(n556), .Z(n59) );
  XOR U542 ( .A(n557), .B(n558), .Z(n556) );
  NAND U543 ( .A(b[1]), .B(a[72]), .Z(n558) );
  AND U544 ( .A(b[0]), .B(a[73]), .Z(n557) );
  IV U545 ( .A(n554), .Z(n555) );
  XOR U546 ( .A(n559), .B(n560), .Z(n554) );
  ANDN U547 ( .B(n61), .A(n62), .Z(n559) );
  XOR U548 ( .A(sreg[200]), .B(n561), .Z(n62) );
  XOR U549 ( .A(n561), .B(n562), .Z(n61) );
  XOR U550 ( .A(n563), .B(n564), .Z(n562) );
  NAND U551 ( .A(b[1]), .B(a[71]), .Z(n564) );
  AND U552 ( .A(b[0]), .B(a[72]), .Z(n563) );
  IV U553 ( .A(n560), .Z(n561) );
  XOR U554 ( .A(n565), .B(n566), .Z(n560) );
  ANDN U555 ( .B(n63), .A(n64), .Z(n565) );
  XOR U556 ( .A(sreg[199]), .B(n567), .Z(n64) );
  XOR U557 ( .A(n567), .B(n568), .Z(n63) );
  XOR U558 ( .A(n569), .B(n570), .Z(n568) );
  NAND U559 ( .A(b[1]), .B(a[70]), .Z(n570) );
  AND U560 ( .A(b[0]), .B(a[71]), .Z(n569) );
  IV U561 ( .A(n566), .Z(n567) );
  XOR U562 ( .A(n571), .B(n572), .Z(n566) );
  ANDN U563 ( .B(n65), .A(n66), .Z(n571) );
  XOR U564 ( .A(sreg[198]), .B(n573), .Z(n66) );
  XOR U565 ( .A(n573), .B(n574), .Z(n65) );
  XOR U566 ( .A(n575), .B(n576), .Z(n574) );
  NAND U567 ( .A(b[1]), .B(a[69]), .Z(n576) );
  AND U568 ( .A(b[0]), .B(a[70]), .Z(n575) );
  IV U569 ( .A(n572), .Z(n573) );
  XOR U570 ( .A(n577), .B(n578), .Z(n572) );
  ANDN U571 ( .B(n69), .A(n70), .Z(n577) );
  XOR U572 ( .A(sreg[197]), .B(n579), .Z(n70) );
  XOR U573 ( .A(n579), .B(n580), .Z(n69) );
  XOR U574 ( .A(n581), .B(n582), .Z(n580) );
  NAND U575 ( .A(b[1]), .B(a[68]), .Z(n582) );
  AND U576 ( .A(b[0]), .B(a[69]), .Z(n581) );
  IV U577 ( .A(n578), .Z(n579) );
  XOR U578 ( .A(n583), .B(n584), .Z(n578) );
  ANDN U579 ( .B(n71), .A(n72), .Z(n583) );
  XOR U580 ( .A(sreg[196]), .B(n585), .Z(n72) );
  XOR U581 ( .A(n585), .B(n586), .Z(n71) );
  XOR U582 ( .A(n587), .B(n588), .Z(n586) );
  NAND U583 ( .A(b[1]), .B(a[67]), .Z(n588) );
  AND U584 ( .A(b[0]), .B(a[68]), .Z(n587) );
  IV U585 ( .A(n584), .Z(n585) );
  XOR U586 ( .A(n589), .B(n590), .Z(n584) );
  ANDN U587 ( .B(n73), .A(n74), .Z(n589) );
  XOR U588 ( .A(sreg[195]), .B(n591), .Z(n74) );
  XOR U589 ( .A(n591), .B(n592), .Z(n73) );
  XOR U590 ( .A(n593), .B(n594), .Z(n592) );
  NAND U591 ( .A(b[1]), .B(a[66]), .Z(n594) );
  AND U592 ( .A(b[0]), .B(a[67]), .Z(n593) );
  IV U593 ( .A(n590), .Z(n591) );
  XOR U594 ( .A(n595), .B(n596), .Z(n590) );
  ANDN U595 ( .B(n75), .A(n76), .Z(n595) );
  XOR U596 ( .A(sreg[194]), .B(n597), .Z(n76) );
  XOR U597 ( .A(n597), .B(n598), .Z(n75) );
  XOR U598 ( .A(n599), .B(n600), .Z(n598) );
  NAND U599 ( .A(b[1]), .B(a[65]), .Z(n600) );
  AND U600 ( .A(b[0]), .B(a[66]), .Z(n599) );
  IV U601 ( .A(n596), .Z(n597) );
  XOR U602 ( .A(n601), .B(n602), .Z(n596) );
  ANDN U603 ( .B(n77), .A(n78), .Z(n601) );
  XOR U604 ( .A(sreg[193]), .B(n603), .Z(n78) );
  XOR U605 ( .A(n603), .B(n604), .Z(n77) );
  XOR U606 ( .A(n605), .B(n606), .Z(n604) );
  NAND U607 ( .A(b[1]), .B(a[64]), .Z(n606) );
  AND U608 ( .A(b[0]), .B(a[65]), .Z(n605) );
  IV U609 ( .A(n602), .Z(n603) );
  XOR U610 ( .A(n607), .B(n608), .Z(n602) );
  ANDN U611 ( .B(n79), .A(n80), .Z(n607) );
  XOR U612 ( .A(sreg[192]), .B(n609), .Z(n80) );
  XOR U613 ( .A(n609), .B(n610), .Z(n79) );
  XOR U614 ( .A(n611), .B(n612), .Z(n610) );
  NAND U615 ( .A(b[1]), .B(a[63]), .Z(n612) );
  AND U616 ( .A(b[0]), .B(a[64]), .Z(n611) );
  IV U617 ( .A(n608), .Z(n609) );
  XOR U618 ( .A(n613), .B(n614), .Z(n608) );
  ANDN U619 ( .B(n81), .A(n82), .Z(n613) );
  XOR U620 ( .A(sreg[191]), .B(n615), .Z(n82) );
  XOR U621 ( .A(n615), .B(n616), .Z(n81) );
  XOR U622 ( .A(n617), .B(n618), .Z(n616) );
  NAND U623 ( .A(b[1]), .B(a[62]), .Z(n618) );
  AND U624 ( .A(b[0]), .B(a[63]), .Z(n617) );
  IV U625 ( .A(n614), .Z(n615) );
  XOR U626 ( .A(n619), .B(n620), .Z(n614) );
  ANDN U627 ( .B(n83), .A(n84), .Z(n619) );
  XOR U628 ( .A(sreg[190]), .B(n621), .Z(n84) );
  XOR U629 ( .A(n621), .B(n622), .Z(n83) );
  XOR U630 ( .A(n623), .B(n624), .Z(n622) );
  NAND U631 ( .A(b[1]), .B(a[61]), .Z(n624) );
  AND U632 ( .A(b[0]), .B(a[62]), .Z(n623) );
  IV U633 ( .A(n620), .Z(n621) );
  XOR U634 ( .A(n625), .B(n626), .Z(n620) );
  ANDN U635 ( .B(n85), .A(n86), .Z(n625) );
  XOR U636 ( .A(sreg[189]), .B(n627), .Z(n86) );
  XOR U637 ( .A(n627), .B(n628), .Z(n85) );
  XOR U638 ( .A(n629), .B(n630), .Z(n628) );
  NAND U639 ( .A(b[1]), .B(a[60]), .Z(n630) );
  AND U640 ( .A(b[0]), .B(a[61]), .Z(n629) );
  IV U641 ( .A(n626), .Z(n627) );
  XOR U642 ( .A(n631), .B(n632), .Z(n626) );
  ANDN U643 ( .B(n87), .A(n88), .Z(n631) );
  XOR U644 ( .A(sreg[188]), .B(n633), .Z(n88) );
  XOR U645 ( .A(n633), .B(n634), .Z(n87) );
  XOR U646 ( .A(n635), .B(n636), .Z(n634) );
  NAND U647 ( .A(b[1]), .B(a[59]), .Z(n636) );
  AND U648 ( .A(b[0]), .B(a[60]), .Z(n635) );
  IV U649 ( .A(n632), .Z(n633) );
  XOR U650 ( .A(n637), .B(n638), .Z(n632) );
  ANDN U651 ( .B(n91), .A(n92), .Z(n637) );
  XOR U652 ( .A(sreg[187]), .B(n639), .Z(n92) );
  XOR U653 ( .A(n639), .B(n640), .Z(n91) );
  XOR U654 ( .A(n641), .B(n642), .Z(n640) );
  NAND U655 ( .A(b[1]), .B(a[58]), .Z(n642) );
  AND U656 ( .A(b[0]), .B(a[59]), .Z(n641) );
  IV U657 ( .A(n638), .Z(n639) );
  XOR U658 ( .A(n643), .B(n644), .Z(n638) );
  ANDN U659 ( .B(n93), .A(n94), .Z(n643) );
  XOR U660 ( .A(sreg[186]), .B(n645), .Z(n94) );
  XOR U661 ( .A(n645), .B(n646), .Z(n93) );
  XOR U662 ( .A(n647), .B(n648), .Z(n646) );
  NAND U663 ( .A(b[1]), .B(a[57]), .Z(n648) );
  AND U664 ( .A(b[0]), .B(a[58]), .Z(n647) );
  IV U665 ( .A(n644), .Z(n645) );
  XOR U666 ( .A(n649), .B(n650), .Z(n644) );
  ANDN U667 ( .B(n95), .A(n96), .Z(n649) );
  XOR U668 ( .A(sreg[185]), .B(n651), .Z(n96) );
  XOR U669 ( .A(n651), .B(n652), .Z(n95) );
  XOR U670 ( .A(n653), .B(n654), .Z(n652) );
  NAND U671 ( .A(b[1]), .B(a[56]), .Z(n654) );
  AND U672 ( .A(b[0]), .B(a[57]), .Z(n653) );
  IV U673 ( .A(n650), .Z(n651) );
  XOR U674 ( .A(n655), .B(n656), .Z(n650) );
  ANDN U675 ( .B(n97), .A(n98), .Z(n655) );
  XOR U676 ( .A(sreg[184]), .B(n657), .Z(n98) );
  XOR U677 ( .A(n657), .B(n658), .Z(n97) );
  XOR U678 ( .A(n659), .B(n660), .Z(n658) );
  NAND U679 ( .A(b[1]), .B(a[55]), .Z(n660) );
  AND U680 ( .A(b[0]), .B(a[56]), .Z(n659) );
  IV U681 ( .A(n656), .Z(n657) );
  XOR U682 ( .A(n661), .B(n662), .Z(n656) );
  ANDN U683 ( .B(n99), .A(n100), .Z(n661) );
  XOR U684 ( .A(sreg[183]), .B(n663), .Z(n100) );
  XOR U685 ( .A(n663), .B(n664), .Z(n99) );
  XOR U686 ( .A(n665), .B(n666), .Z(n664) );
  NAND U687 ( .A(b[1]), .B(a[54]), .Z(n666) );
  AND U688 ( .A(b[0]), .B(a[55]), .Z(n665) );
  IV U689 ( .A(n662), .Z(n663) );
  XOR U690 ( .A(n667), .B(n668), .Z(n662) );
  ANDN U691 ( .B(n101), .A(n102), .Z(n667) );
  XOR U692 ( .A(sreg[182]), .B(n669), .Z(n102) );
  XOR U693 ( .A(n669), .B(n670), .Z(n101) );
  XOR U694 ( .A(n671), .B(n672), .Z(n670) );
  NAND U695 ( .A(b[1]), .B(a[53]), .Z(n672) );
  AND U696 ( .A(b[0]), .B(a[54]), .Z(n671) );
  IV U697 ( .A(n668), .Z(n669) );
  XOR U698 ( .A(n673), .B(n674), .Z(n668) );
  ANDN U699 ( .B(n103), .A(n104), .Z(n673) );
  XOR U700 ( .A(sreg[181]), .B(n675), .Z(n104) );
  XOR U701 ( .A(n675), .B(n676), .Z(n103) );
  XOR U702 ( .A(n677), .B(n678), .Z(n676) );
  NAND U703 ( .A(b[1]), .B(a[52]), .Z(n678) );
  AND U704 ( .A(b[0]), .B(a[53]), .Z(n677) );
  IV U705 ( .A(n674), .Z(n675) );
  XOR U706 ( .A(n679), .B(n680), .Z(n674) );
  ANDN U707 ( .B(n105), .A(n106), .Z(n679) );
  XOR U708 ( .A(sreg[180]), .B(n681), .Z(n106) );
  XOR U709 ( .A(n681), .B(n682), .Z(n105) );
  XOR U710 ( .A(n683), .B(n684), .Z(n682) );
  NAND U711 ( .A(b[1]), .B(a[51]), .Z(n684) );
  AND U712 ( .A(b[0]), .B(a[52]), .Z(n683) );
  IV U713 ( .A(n680), .Z(n681) );
  XOR U714 ( .A(n685), .B(n686), .Z(n680) );
  ANDN U715 ( .B(n107), .A(n108), .Z(n685) );
  XOR U716 ( .A(sreg[179]), .B(n687), .Z(n108) );
  XOR U717 ( .A(n687), .B(n688), .Z(n107) );
  XOR U718 ( .A(n689), .B(n690), .Z(n688) );
  NAND U719 ( .A(b[1]), .B(a[50]), .Z(n690) );
  AND U720 ( .A(b[0]), .B(a[51]), .Z(n689) );
  IV U721 ( .A(n686), .Z(n687) );
  XOR U722 ( .A(n691), .B(n692), .Z(n686) );
  ANDN U723 ( .B(n109), .A(n110), .Z(n691) );
  XOR U724 ( .A(sreg[178]), .B(n693), .Z(n110) );
  XOR U725 ( .A(n693), .B(n694), .Z(n109) );
  XOR U726 ( .A(n695), .B(n696), .Z(n694) );
  NAND U727 ( .A(b[1]), .B(a[49]), .Z(n696) );
  AND U728 ( .A(b[0]), .B(a[50]), .Z(n695) );
  IV U729 ( .A(n692), .Z(n693) );
  XOR U730 ( .A(n697), .B(n698), .Z(n692) );
  ANDN U731 ( .B(n113), .A(n114), .Z(n697) );
  XOR U732 ( .A(sreg[177]), .B(n699), .Z(n114) );
  XOR U733 ( .A(n699), .B(n700), .Z(n113) );
  XOR U734 ( .A(n701), .B(n702), .Z(n700) );
  NAND U735 ( .A(b[1]), .B(a[48]), .Z(n702) );
  AND U736 ( .A(b[0]), .B(a[49]), .Z(n701) );
  IV U737 ( .A(n698), .Z(n699) );
  XOR U738 ( .A(n703), .B(n704), .Z(n698) );
  ANDN U739 ( .B(n115), .A(n116), .Z(n703) );
  XOR U740 ( .A(sreg[176]), .B(n705), .Z(n116) );
  XOR U741 ( .A(n705), .B(n706), .Z(n115) );
  XOR U742 ( .A(n707), .B(n708), .Z(n706) );
  NAND U743 ( .A(b[1]), .B(a[47]), .Z(n708) );
  AND U744 ( .A(b[0]), .B(a[48]), .Z(n707) );
  IV U745 ( .A(n704), .Z(n705) );
  XOR U746 ( .A(n709), .B(n710), .Z(n704) );
  ANDN U747 ( .B(n117), .A(n118), .Z(n709) );
  XOR U748 ( .A(sreg[175]), .B(n711), .Z(n118) );
  XOR U749 ( .A(n711), .B(n712), .Z(n117) );
  XOR U750 ( .A(n713), .B(n714), .Z(n712) );
  NAND U751 ( .A(b[1]), .B(a[46]), .Z(n714) );
  AND U752 ( .A(b[0]), .B(a[47]), .Z(n713) );
  IV U753 ( .A(n710), .Z(n711) );
  XOR U754 ( .A(n715), .B(n716), .Z(n710) );
  ANDN U755 ( .B(n119), .A(n120), .Z(n715) );
  XOR U756 ( .A(sreg[174]), .B(n717), .Z(n120) );
  XOR U757 ( .A(n717), .B(n718), .Z(n119) );
  XOR U758 ( .A(n719), .B(n720), .Z(n718) );
  NAND U759 ( .A(b[1]), .B(a[45]), .Z(n720) );
  AND U760 ( .A(b[0]), .B(a[46]), .Z(n719) );
  IV U761 ( .A(n716), .Z(n717) );
  XOR U762 ( .A(n721), .B(n722), .Z(n716) );
  ANDN U763 ( .B(n121), .A(n122), .Z(n721) );
  XOR U764 ( .A(sreg[173]), .B(n723), .Z(n122) );
  XOR U765 ( .A(n723), .B(n724), .Z(n121) );
  XOR U766 ( .A(n725), .B(n726), .Z(n724) );
  NAND U767 ( .A(b[1]), .B(a[44]), .Z(n726) );
  AND U768 ( .A(b[0]), .B(a[45]), .Z(n725) );
  IV U769 ( .A(n722), .Z(n723) );
  XOR U770 ( .A(n727), .B(n728), .Z(n722) );
  ANDN U771 ( .B(n123), .A(n124), .Z(n727) );
  XOR U772 ( .A(sreg[172]), .B(n729), .Z(n124) );
  XOR U773 ( .A(n729), .B(n730), .Z(n123) );
  XOR U774 ( .A(n731), .B(n732), .Z(n730) );
  NAND U775 ( .A(b[1]), .B(a[43]), .Z(n732) );
  AND U776 ( .A(b[0]), .B(a[44]), .Z(n731) );
  IV U777 ( .A(n728), .Z(n729) );
  XOR U778 ( .A(n733), .B(n734), .Z(n728) );
  ANDN U779 ( .B(n125), .A(n126), .Z(n733) );
  XOR U780 ( .A(sreg[171]), .B(n735), .Z(n126) );
  XOR U781 ( .A(n735), .B(n736), .Z(n125) );
  XOR U782 ( .A(n737), .B(n738), .Z(n736) );
  NAND U783 ( .A(b[1]), .B(a[42]), .Z(n738) );
  AND U784 ( .A(b[0]), .B(a[43]), .Z(n737) );
  IV U785 ( .A(n734), .Z(n735) );
  XOR U786 ( .A(n739), .B(n740), .Z(n734) );
  ANDN U787 ( .B(n127), .A(n128), .Z(n739) );
  XOR U788 ( .A(sreg[170]), .B(n741), .Z(n128) );
  XOR U789 ( .A(n741), .B(n742), .Z(n127) );
  XOR U790 ( .A(n743), .B(n744), .Z(n742) );
  NAND U791 ( .A(b[1]), .B(a[41]), .Z(n744) );
  AND U792 ( .A(b[0]), .B(a[42]), .Z(n743) );
  IV U793 ( .A(n740), .Z(n741) );
  XOR U794 ( .A(n745), .B(n746), .Z(n740) );
  ANDN U795 ( .B(n129), .A(n130), .Z(n745) );
  XOR U796 ( .A(sreg[169]), .B(n747), .Z(n130) );
  XOR U797 ( .A(n747), .B(n748), .Z(n129) );
  XOR U798 ( .A(n749), .B(n750), .Z(n748) );
  NAND U799 ( .A(b[1]), .B(a[40]), .Z(n750) );
  AND U800 ( .A(b[0]), .B(a[41]), .Z(n749) );
  IV U801 ( .A(n746), .Z(n747) );
  XOR U802 ( .A(n751), .B(n752), .Z(n746) );
  ANDN U803 ( .B(n131), .A(n132), .Z(n751) );
  XOR U804 ( .A(sreg[168]), .B(n753), .Z(n132) );
  XOR U805 ( .A(n753), .B(n754), .Z(n131) );
  XOR U806 ( .A(n755), .B(n756), .Z(n754) );
  NAND U807 ( .A(b[1]), .B(a[39]), .Z(n756) );
  AND U808 ( .A(b[0]), .B(a[40]), .Z(n755) );
  IV U809 ( .A(n752), .Z(n753) );
  XOR U810 ( .A(n757), .B(n758), .Z(n752) );
  ANDN U811 ( .B(n135), .A(n136), .Z(n757) );
  XOR U812 ( .A(sreg[167]), .B(n759), .Z(n136) );
  XOR U813 ( .A(n759), .B(n760), .Z(n135) );
  XOR U814 ( .A(n761), .B(n762), .Z(n760) );
  NAND U815 ( .A(b[1]), .B(a[38]), .Z(n762) );
  AND U816 ( .A(b[0]), .B(a[39]), .Z(n761) );
  IV U817 ( .A(n758), .Z(n759) );
  XOR U818 ( .A(n763), .B(n764), .Z(n758) );
  ANDN U819 ( .B(n137), .A(n138), .Z(n763) );
  XOR U820 ( .A(sreg[166]), .B(n765), .Z(n138) );
  XOR U821 ( .A(n765), .B(n766), .Z(n137) );
  XOR U822 ( .A(n767), .B(n768), .Z(n766) );
  NAND U823 ( .A(b[1]), .B(a[37]), .Z(n768) );
  AND U824 ( .A(b[0]), .B(a[38]), .Z(n767) );
  IV U825 ( .A(n764), .Z(n765) );
  XOR U826 ( .A(n769), .B(n770), .Z(n764) );
  ANDN U827 ( .B(n139), .A(n140), .Z(n769) );
  XOR U828 ( .A(sreg[165]), .B(n771), .Z(n140) );
  XOR U829 ( .A(n771), .B(n772), .Z(n139) );
  XOR U830 ( .A(n773), .B(n774), .Z(n772) );
  NAND U831 ( .A(b[1]), .B(a[36]), .Z(n774) );
  AND U832 ( .A(b[0]), .B(a[37]), .Z(n773) );
  IV U833 ( .A(n770), .Z(n771) );
  XOR U834 ( .A(n775), .B(n776), .Z(n770) );
  ANDN U835 ( .B(n141), .A(n142), .Z(n775) );
  XOR U836 ( .A(sreg[164]), .B(n777), .Z(n142) );
  XOR U837 ( .A(n777), .B(n778), .Z(n141) );
  XOR U838 ( .A(n779), .B(n780), .Z(n778) );
  NAND U839 ( .A(b[1]), .B(a[35]), .Z(n780) );
  AND U840 ( .A(b[0]), .B(a[36]), .Z(n779) );
  IV U841 ( .A(n776), .Z(n777) );
  XOR U842 ( .A(n781), .B(n782), .Z(n776) );
  ANDN U843 ( .B(n143), .A(n144), .Z(n781) );
  XOR U844 ( .A(sreg[163]), .B(n783), .Z(n144) );
  XOR U845 ( .A(n783), .B(n784), .Z(n143) );
  XOR U846 ( .A(n785), .B(n786), .Z(n784) );
  NAND U847 ( .A(b[1]), .B(a[34]), .Z(n786) );
  AND U848 ( .A(b[0]), .B(a[35]), .Z(n785) );
  IV U849 ( .A(n782), .Z(n783) );
  XOR U850 ( .A(n787), .B(n788), .Z(n782) );
  ANDN U851 ( .B(n145), .A(n146), .Z(n787) );
  XOR U852 ( .A(sreg[162]), .B(n789), .Z(n146) );
  XOR U853 ( .A(n789), .B(n790), .Z(n145) );
  XOR U854 ( .A(n791), .B(n792), .Z(n790) );
  NAND U855 ( .A(b[1]), .B(a[33]), .Z(n792) );
  AND U856 ( .A(b[0]), .B(a[34]), .Z(n791) );
  IV U857 ( .A(n788), .Z(n789) );
  XOR U858 ( .A(n793), .B(n794), .Z(n788) );
  ANDN U859 ( .B(n147), .A(n148), .Z(n793) );
  XOR U860 ( .A(sreg[161]), .B(n795), .Z(n148) );
  XOR U861 ( .A(n795), .B(n796), .Z(n147) );
  XOR U862 ( .A(n797), .B(n798), .Z(n796) );
  NAND U863 ( .A(b[1]), .B(a[32]), .Z(n798) );
  AND U864 ( .A(b[0]), .B(a[33]), .Z(n797) );
  IV U865 ( .A(n794), .Z(n795) );
  XOR U866 ( .A(n799), .B(n800), .Z(n794) );
  ANDN U867 ( .B(n149), .A(n150), .Z(n799) );
  XOR U868 ( .A(sreg[160]), .B(n801), .Z(n150) );
  XOR U869 ( .A(n801), .B(n802), .Z(n149) );
  XOR U870 ( .A(n803), .B(n804), .Z(n802) );
  NAND U871 ( .A(b[1]), .B(a[31]), .Z(n804) );
  AND U872 ( .A(b[0]), .B(a[32]), .Z(n803) );
  IV U873 ( .A(n800), .Z(n801) );
  XOR U874 ( .A(n805), .B(n806), .Z(n800) );
  ANDN U875 ( .B(n151), .A(n152), .Z(n805) );
  XOR U876 ( .A(sreg[159]), .B(n807), .Z(n152) );
  XOR U877 ( .A(n807), .B(n808), .Z(n151) );
  XOR U878 ( .A(n809), .B(n810), .Z(n808) );
  NAND U879 ( .A(b[1]), .B(a[30]), .Z(n810) );
  AND U880 ( .A(b[0]), .B(a[31]), .Z(n809) );
  IV U881 ( .A(n806), .Z(n807) );
  XOR U882 ( .A(n811), .B(n812), .Z(n806) );
  ANDN U883 ( .B(n153), .A(n154), .Z(n811) );
  XOR U884 ( .A(sreg[158]), .B(n813), .Z(n154) );
  XOR U885 ( .A(n813), .B(n814), .Z(n153) );
  XOR U886 ( .A(n815), .B(n816), .Z(n814) );
  NAND U887 ( .A(b[1]), .B(a[29]), .Z(n816) );
  AND U888 ( .A(b[0]), .B(a[30]), .Z(n815) );
  IV U889 ( .A(n812), .Z(n813) );
  XOR U890 ( .A(n817), .B(n818), .Z(n812) );
  ANDN U891 ( .B(n157), .A(n158), .Z(n817) );
  XOR U892 ( .A(sreg[157]), .B(n819), .Z(n158) );
  XOR U893 ( .A(n819), .B(n820), .Z(n157) );
  XOR U894 ( .A(n821), .B(n822), .Z(n820) );
  NAND U895 ( .A(b[1]), .B(a[28]), .Z(n822) );
  AND U896 ( .A(b[0]), .B(a[29]), .Z(n821) );
  IV U897 ( .A(n818), .Z(n819) );
  XOR U898 ( .A(n823), .B(n824), .Z(n818) );
  ANDN U899 ( .B(n159), .A(n160), .Z(n823) );
  XOR U900 ( .A(sreg[156]), .B(n825), .Z(n160) );
  XOR U901 ( .A(n825), .B(n826), .Z(n159) );
  XOR U902 ( .A(n827), .B(n828), .Z(n826) );
  NAND U903 ( .A(b[1]), .B(a[27]), .Z(n828) );
  AND U904 ( .A(b[0]), .B(a[28]), .Z(n827) );
  IV U905 ( .A(n824), .Z(n825) );
  XOR U906 ( .A(n829), .B(n830), .Z(n824) );
  ANDN U907 ( .B(n161), .A(n162), .Z(n829) );
  XOR U908 ( .A(sreg[155]), .B(n831), .Z(n162) );
  XOR U909 ( .A(n831), .B(n832), .Z(n161) );
  XOR U910 ( .A(n833), .B(n834), .Z(n832) );
  NAND U911 ( .A(b[1]), .B(a[26]), .Z(n834) );
  AND U912 ( .A(b[0]), .B(a[27]), .Z(n833) );
  IV U913 ( .A(n830), .Z(n831) );
  XOR U914 ( .A(n835), .B(n836), .Z(n830) );
  ANDN U915 ( .B(n163), .A(n164), .Z(n835) );
  XOR U916 ( .A(sreg[154]), .B(n837), .Z(n164) );
  XOR U917 ( .A(n837), .B(n838), .Z(n163) );
  XOR U918 ( .A(n839), .B(n840), .Z(n838) );
  NAND U919 ( .A(b[1]), .B(a[25]), .Z(n840) );
  AND U920 ( .A(b[0]), .B(a[26]), .Z(n839) );
  IV U921 ( .A(n836), .Z(n837) );
  XOR U922 ( .A(n841), .B(n842), .Z(n836) );
  ANDN U923 ( .B(n165), .A(n166), .Z(n841) );
  XOR U924 ( .A(sreg[153]), .B(n843), .Z(n166) );
  XOR U925 ( .A(n843), .B(n844), .Z(n165) );
  XOR U926 ( .A(n845), .B(n846), .Z(n844) );
  NAND U927 ( .A(b[1]), .B(a[24]), .Z(n846) );
  AND U928 ( .A(b[0]), .B(a[25]), .Z(n845) );
  IV U929 ( .A(n842), .Z(n843) );
  XOR U930 ( .A(n847), .B(n848), .Z(n842) );
  ANDN U931 ( .B(n167), .A(n168), .Z(n847) );
  XOR U932 ( .A(sreg[152]), .B(n849), .Z(n168) );
  XOR U933 ( .A(n849), .B(n850), .Z(n167) );
  XOR U934 ( .A(n851), .B(n852), .Z(n850) );
  NAND U935 ( .A(b[1]), .B(a[23]), .Z(n852) );
  AND U936 ( .A(b[0]), .B(a[24]), .Z(n851) );
  IV U937 ( .A(n848), .Z(n849) );
  XOR U938 ( .A(n853), .B(n854), .Z(n848) );
  ANDN U939 ( .B(n169), .A(n170), .Z(n853) );
  XOR U940 ( .A(sreg[151]), .B(n855), .Z(n170) );
  XOR U941 ( .A(n855), .B(n856), .Z(n169) );
  XOR U942 ( .A(n857), .B(n858), .Z(n856) );
  NAND U943 ( .A(b[1]), .B(a[22]), .Z(n858) );
  AND U944 ( .A(b[0]), .B(a[23]), .Z(n857) );
  IV U945 ( .A(n854), .Z(n855) );
  XOR U946 ( .A(n859), .B(n860), .Z(n854) );
  ANDN U947 ( .B(n171), .A(n172), .Z(n859) );
  XOR U948 ( .A(sreg[150]), .B(n861), .Z(n172) );
  XOR U949 ( .A(n861), .B(n862), .Z(n171) );
  XOR U950 ( .A(n863), .B(n864), .Z(n862) );
  NAND U951 ( .A(b[1]), .B(a[21]), .Z(n864) );
  AND U952 ( .A(b[0]), .B(a[22]), .Z(n863) );
  IV U953 ( .A(n860), .Z(n861) );
  XOR U954 ( .A(n865), .B(n866), .Z(n860) );
  ANDN U955 ( .B(n173), .A(n174), .Z(n865) );
  XOR U956 ( .A(sreg[149]), .B(n867), .Z(n174) );
  XOR U957 ( .A(n867), .B(n868), .Z(n173) );
  XOR U958 ( .A(n869), .B(n870), .Z(n868) );
  NAND U959 ( .A(b[1]), .B(a[20]), .Z(n870) );
  AND U960 ( .A(b[0]), .B(a[21]), .Z(n869) );
  IV U961 ( .A(n866), .Z(n867) );
  XOR U962 ( .A(n871), .B(n872), .Z(n866) );
  ANDN U963 ( .B(n175), .A(n176), .Z(n871) );
  XOR U964 ( .A(sreg[148]), .B(n873), .Z(n176) );
  XOR U965 ( .A(n873), .B(n874), .Z(n175) );
  XOR U966 ( .A(n875), .B(n876), .Z(n874) );
  NAND U967 ( .A(b[1]), .B(a[19]), .Z(n876) );
  AND U968 ( .A(b[0]), .B(a[20]), .Z(n875) );
  IV U969 ( .A(n872), .Z(n873) );
  XOR U970 ( .A(n877), .B(n878), .Z(n872) );
  ANDN U971 ( .B(n177), .A(n178), .Z(n877) );
  XOR U972 ( .A(sreg[147]), .B(n879), .Z(n178) );
  XOR U973 ( .A(n879), .B(n880), .Z(n177) );
  XOR U974 ( .A(n881), .B(n882), .Z(n880) );
  NAND U975 ( .A(b[1]), .B(a[18]), .Z(n882) );
  AND U976 ( .A(b[0]), .B(a[19]), .Z(n881) );
  IV U977 ( .A(n878), .Z(n879) );
  XOR U978 ( .A(n883), .B(n884), .Z(n878) );
  ANDN U979 ( .B(n179), .A(n180), .Z(n883) );
  XOR U980 ( .A(sreg[146]), .B(n885), .Z(n180) );
  XOR U981 ( .A(n885), .B(n886), .Z(n179) );
  XOR U982 ( .A(n887), .B(n888), .Z(n886) );
  NAND U983 ( .A(b[1]), .B(a[17]), .Z(n888) );
  AND U984 ( .A(b[0]), .B(a[18]), .Z(n887) );
  IV U985 ( .A(n884), .Z(n885) );
  XOR U986 ( .A(n889), .B(n890), .Z(n884) );
  ANDN U987 ( .B(n181), .A(n182), .Z(n889) );
  XOR U988 ( .A(sreg[145]), .B(n891), .Z(n182) );
  XOR U989 ( .A(n891), .B(n892), .Z(n181) );
  XOR U990 ( .A(n893), .B(n894), .Z(n892) );
  NAND U991 ( .A(b[1]), .B(a[16]), .Z(n894) );
  AND U992 ( .A(b[0]), .B(a[17]), .Z(n893) );
  IV U993 ( .A(n890), .Z(n891) );
  XOR U994 ( .A(n895), .B(n896), .Z(n890) );
  ANDN U995 ( .B(n183), .A(n184), .Z(n895) );
  XOR U996 ( .A(sreg[144]), .B(n897), .Z(n184) );
  XOR U997 ( .A(n897), .B(n898), .Z(n183) );
  XOR U998 ( .A(n899), .B(n900), .Z(n898) );
  NAND U999 ( .A(b[1]), .B(a[15]), .Z(n900) );
  AND U1000 ( .A(b[0]), .B(a[16]), .Z(n899) );
  IV U1001 ( .A(n896), .Z(n897) );
  XOR U1002 ( .A(n901), .B(n902), .Z(n896) );
  ANDN U1003 ( .B(n185), .A(n186), .Z(n901) );
  XOR U1004 ( .A(sreg[143]), .B(n903), .Z(n186) );
  XOR U1005 ( .A(n903), .B(n904), .Z(n185) );
  XOR U1006 ( .A(n905), .B(n906), .Z(n904) );
  NAND U1007 ( .A(b[1]), .B(a[14]), .Z(n906) );
  AND U1008 ( .A(b[0]), .B(a[15]), .Z(n905) );
  IV U1009 ( .A(n902), .Z(n903) );
  XOR U1010 ( .A(n907), .B(n908), .Z(n902) );
  ANDN U1011 ( .B(n187), .A(n188), .Z(n907) );
  XOR U1012 ( .A(sreg[142]), .B(n909), .Z(n188) );
  XOR U1013 ( .A(n909), .B(n910), .Z(n187) );
  XOR U1014 ( .A(n911), .B(n912), .Z(n910) );
  NAND U1015 ( .A(b[1]), .B(a[13]), .Z(n912) );
  AND U1016 ( .A(b[0]), .B(a[14]), .Z(n911) );
  IV U1017 ( .A(n908), .Z(n909) );
  XOR U1018 ( .A(n913), .B(n914), .Z(n908) );
  ANDN U1019 ( .B(n189), .A(n190), .Z(n913) );
  XOR U1020 ( .A(sreg[141]), .B(n915), .Z(n190) );
  XOR U1021 ( .A(n915), .B(n916), .Z(n189) );
  XOR U1022 ( .A(n917), .B(n918), .Z(n916) );
  NAND U1023 ( .A(b[1]), .B(a[12]), .Z(n918) );
  AND U1024 ( .A(b[0]), .B(a[13]), .Z(n917) );
  IV U1025 ( .A(n914), .Z(n915) );
  XOR U1026 ( .A(n919), .B(n920), .Z(n914) );
  ANDN U1027 ( .B(n191), .A(n192), .Z(n919) );
  XOR U1028 ( .A(sreg[140]), .B(n921), .Z(n192) );
  XOR U1029 ( .A(n921), .B(n922), .Z(n191) );
  XOR U1030 ( .A(n923), .B(n924), .Z(n922) );
  NAND U1031 ( .A(b[1]), .B(a[11]), .Z(n924) );
  AND U1032 ( .A(b[0]), .B(a[12]), .Z(n923) );
  IV U1033 ( .A(n920), .Z(n921) );
  XOR U1034 ( .A(n925), .B(n926), .Z(n920) );
  ANDN U1035 ( .B(n237), .A(n238), .Z(n925) );
  XOR U1036 ( .A(sreg[139]), .B(n927), .Z(n238) );
  XOR U1037 ( .A(n927), .B(n928), .Z(n237) );
  XOR U1038 ( .A(n929), .B(n930), .Z(n928) );
  NAND U1039 ( .A(b[1]), .B(a[10]), .Z(n930) );
  AND U1040 ( .A(b[0]), .B(a[11]), .Z(n929) );
  IV U1041 ( .A(n926), .Z(n927) );
  XOR U1042 ( .A(n931), .B(n932), .Z(n926) );
  ANDN U1043 ( .B(n319), .A(n320), .Z(n931) );
  XOR U1044 ( .A(sreg[138]), .B(n933), .Z(n320) );
  XOR U1045 ( .A(n933), .B(n934), .Z(n319) );
  XOR U1046 ( .A(n935), .B(n936), .Z(n934) );
  NAND U1047 ( .A(b[1]), .B(a[9]), .Z(n936) );
  AND U1048 ( .A(b[0]), .B(a[10]), .Z(n935) );
  IV U1049 ( .A(n932), .Z(n933) );
  XOR U1050 ( .A(n937), .B(n938), .Z(n932) );
  ANDN U1051 ( .B(n2), .A(n1), .Z(n937) );
  XOR U1052 ( .A(sreg[137]), .B(n939), .Z(n1) );
  XOR U1053 ( .A(n939), .B(n940), .Z(n2) );
  XOR U1054 ( .A(n941), .B(n942), .Z(n940) );
  NAND U1055 ( .A(b[1]), .B(a[8]), .Z(n942) );
  AND U1056 ( .A(b[0]), .B(a[9]), .Z(n941) );
  IV U1057 ( .A(n938), .Z(n939) );
  XOR U1058 ( .A(n943), .B(n944), .Z(n938) );
  ANDN U1059 ( .B(n23), .A(n24), .Z(n943) );
  XOR U1060 ( .A(sreg[136]), .B(n945), .Z(n24) );
  XOR U1061 ( .A(n945), .B(n946), .Z(n23) );
  XOR U1062 ( .A(n947), .B(n948), .Z(n946) );
  NAND U1063 ( .A(a[7]), .B(b[1]), .Z(n948) );
  AND U1064 ( .A(a[8]), .B(b[0]), .Z(n947) );
  IV U1065 ( .A(n944), .Z(n945) );
  XOR U1066 ( .A(n949), .B(n950), .Z(n944) );
  ANDN U1067 ( .B(n45), .A(n46), .Z(n949) );
  XOR U1068 ( .A(sreg[135]), .B(n951), .Z(n46) );
  XOR U1069 ( .A(n951), .B(n952), .Z(n45) );
  XOR U1070 ( .A(n953), .B(n954), .Z(n952) );
  NAND U1071 ( .A(b[1]), .B(a[6]), .Z(n954) );
  AND U1072 ( .A(a[7]), .B(b[0]), .Z(n953) );
  IV U1073 ( .A(n950), .Z(n951) );
  XOR U1074 ( .A(n955), .B(n956), .Z(n950) );
  ANDN U1075 ( .B(n67), .A(n68), .Z(n955) );
  XOR U1076 ( .A(sreg[134]), .B(n957), .Z(n68) );
  XOR U1077 ( .A(n957), .B(n958), .Z(n67) );
  XOR U1078 ( .A(n959), .B(n960), .Z(n958) );
  NAND U1079 ( .A(b[1]), .B(a[5]), .Z(n960) );
  AND U1080 ( .A(b[0]), .B(a[6]), .Z(n959) );
  IV U1081 ( .A(n956), .Z(n957) );
  XOR U1082 ( .A(n961), .B(n962), .Z(n956) );
  ANDN U1083 ( .B(n89), .A(n90), .Z(n961) );
  XOR U1084 ( .A(sreg[133]), .B(n963), .Z(n90) );
  XOR U1085 ( .A(n963), .B(n964), .Z(n89) );
  XOR U1086 ( .A(n965), .B(n966), .Z(n964) );
  NAND U1087 ( .A(b[1]), .B(a[4]), .Z(n966) );
  AND U1088 ( .A(b[0]), .B(a[5]), .Z(n965) );
  IV U1089 ( .A(n962), .Z(n963) );
  XOR U1090 ( .A(n967), .B(n968), .Z(n962) );
  ANDN U1091 ( .B(n111), .A(n112), .Z(n967) );
  XOR U1092 ( .A(sreg[132]), .B(n969), .Z(n112) );
  XOR U1093 ( .A(n969), .B(n970), .Z(n111) );
  XOR U1094 ( .A(n971), .B(n972), .Z(n970) );
  NAND U1095 ( .A(b[1]), .B(a[3]), .Z(n972) );
  AND U1096 ( .A(b[0]), .B(a[4]), .Z(n971) );
  IV U1097 ( .A(n968), .Z(n969) );
  XOR U1098 ( .A(n973), .B(n974), .Z(n968) );
  ANDN U1099 ( .B(n133), .A(n134), .Z(n973) );
  XOR U1100 ( .A(sreg[131]), .B(n975), .Z(n134) );
  XOR U1101 ( .A(n975), .B(n976), .Z(n133) );
  XOR U1102 ( .A(n977), .B(n978), .Z(n976) );
  NAND U1103 ( .A(b[1]), .B(a[2]), .Z(n978) );
  AND U1104 ( .A(b[0]), .B(a[3]), .Z(n977) );
  IV U1105 ( .A(n974), .Z(n975) );
  XNOR U1106 ( .A(n979), .B(n980), .Z(n974) );
  ANDN U1107 ( .B(n155), .A(n156), .Z(n979) );
  XOR U1108 ( .A(sreg[130]), .B(n980), .Z(n156) );
  XOR U1109 ( .A(n980), .B(n981), .Z(n155) );
  XOR U1110 ( .A(n982), .B(n983), .Z(n981) );
  NAND U1111 ( .A(b[1]), .B(a[1]), .Z(n983) );
  AND U1112 ( .A(b[0]), .B(a[2]), .Z(n982) );
  XOR U1113 ( .A(n984), .B(n985), .Z(n980) );
  NAND U1114 ( .A(n986), .B(n987), .Z(n985) );
  XOR U1115 ( .A(n986), .B(n987), .Z(c[127]) );
  XOR U1116 ( .A(sreg[129]), .B(n984), .Z(n987) );
  XNOR U1117 ( .A(n984), .B(n988), .Z(n986) );
  XOR U1118 ( .A(n989), .B(n990), .Z(n988) );
  NAND U1119 ( .A(b[0]), .B(a[1]), .Z(n990) );
  AND U1120 ( .A(b[1]), .B(a[0]), .Z(n989) );
  ANDN U1121 ( .B(sreg[128]), .A(n991), .Z(n984) );
  XNOR U1122 ( .A(sreg[128]), .B(n991), .Z(c[126]) );
  NAND U1123 ( .A(a[0]), .B(b[0]), .Z(n991) );
endmodule

