
module mult_N256_CC32 ( clk, rst, a, b, c );
  input [255:0] a;
  input [7:0] b;
  output [511:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583;
  wire   [511:0] sreg;

  DFF \sreg_reg[503]  ( .D(c[511]), .CLK(clk), .RST(rst), .Q(sreg[503]) );
  DFF \sreg_reg[502]  ( .D(c[510]), .CLK(clk), .RST(rst), .Q(sreg[502]) );
  DFF \sreg_reg[501]  ( .D(c[509]), .CLK(clk), .RST(rst), .Q(sreg[501]) );
  DFF \sreg_reg[500]  ( .D(c[508]), .CLK(clk), .RST(rst), .Q(sreg[500]) );
  DFF \sreg_reg[499]  ( .D(c[507]), .CLK(clk), .RST(rst), .Q(sreg[499]) );
  DFF \sreg_reg[498]  ( .D(c[506]), .CLK(clk), .RST(rst), .Q(sreg[498]) );
  DFF \sreg_reg[497]  ( .D(c[505]), .CLK(clk), .RST(rst), .Q(sreg[497]) );
  DFF \sreg_reg[496]  ( .D(c[504]), .CLK(clk), .RST(rst), .Q(sreg[496]) );
  DFF \sreg_reg[495]  ( .D(c[503]), .CLK(clk), .RST(rst), .Q(sreg[495]) );
  DFF \sreg_reg[494]  ( .D(c[502]), .CLK(clk), .RST(rst), .Q(sreg[494]) );
  DFF \sreg_reg[493]  ( .D(c[501]), .CLK(clk), .RST(rst), .Q(sreg[493]) );
  DFF \sreg_reg[492]  ( .D(c[500]), .CLK(clk), .RST(rst), .Q(sreg[492]) );
  DFF \sreg_reg[491]  ( .D(c[499]), .CLK(clk), .RST(rst), .Q(sreg[491]) );
  DFF \sreg_reg[490]  ( .D(c[498]), .CLK(clk), .RST(rst), .Q(sreg[490]) );
  DFF \sreg_reg[489]  ( .D(c[497]), .CLK(clk), .RST(rst), .Q(sreg[489]) );
  DFF \sreg_reg[488]  ( .D(c[496]), .CLK(clk), .RST(rst), .Q(sreg[488]) );
  DFF \sreg_reg[487]  ( .D(c[495]), .CLK(clk), .RST(rst), .Q(sreg[487]) );
  DFF \sreg_reg[486]  ( .D(c[494]), .CLK(clk), .RST(rst), .Q(sreg[486]) );
  DFF \sreg_reg[485]  ( .D(c[493]), .CLK(clk), .RST(rst), .Q(sreg[485]) );
  DFF \sreg_reg[484]  ( .D(c[492]), .CLK(clk), .RST(rst), .Q(sreg[484]) );
  DFF \sreg_reg[483]  ( .D(c[491]), .CLK(clk), .RST(rst), .Q(sreg[483]) );
  DFF \sreg_reg[482]  ( .D(c[490]), .CLK(clk), .RST(rst), .Q(sreg[482]) );
  DFF \sreg_reg[481]  ( .D(c[489]), .CLK(clk), .RST(rst), .Q(sreg[481]) );
  DFF \sreg_reg[480]  ( .D(c[488]), .CLK(clk), .RST(rst), .Q(sreg[480]) );
  DFF \sreg_reg[479]  ( .D(c[487]), .CLK(clk), .RST(rst), .Q(sreg[479]) );
  DFF \sreg_reg[478]  ( .D(c[486]), .CLK(clk), .RST(rst), .Q(sreg[478]) );
  DFF \sreg_reg[477]  ( .D(c[485]), .CLK(clk), .RST(rst), .Q(sreg[477]) );
  DFF \sreg_reg[476]  ( .D(c[484]), .CLK(clk), .RST(rst), .Q(sreg[476]) );
  DFF \sreg_reg[475]  ( .D(c[483]), .CLK(clk), .RST(rst), .Q(sreg[475]) );
  DFF \sreg_reg[474]  ( .D(c[482]), .CLK(clk), .RST(rst), .Q(sreg[474]) );
  DFF \sreg_reg[473]  ( .D(c[481]), .CLK(clk), .RST(rst), .Q(sreg[473]) );
  DFF \sreg_reg[472]  ( .D(c[480]), .CLK(clk), .RST(rst), .Q(sreg[472]) );
  DFF \sreg_reg[471]  ( .D(c[479]), .CLK(clk), .RST(rst), .Q(sreg[471]) );
  DFF \sreg_reg[470]  ( .D(c[478]), .CLK(clk), .RST(rst), .Q(sreg[470]) );
  DFF \sreg_reg[469]  ( .D(c[477]), .CLK(clk), .RST(rst), .Q(sreg[469]) );
  DFF \sreg_reg[468]  ( .D(c[476]), .CLK(clk), .RST(rst), .Q(sreg[468]) );
  DFF \sreg_reg[467]  ( .D(c[475]), .CLK(clk), .RST(rst), .Q(sreg[467]) );
  DFF \sreg_reg[466]  ( .D(c[474]), .CLK(clk), .RST(rst), .Q(sreg[466]) );
  DFF \sreg_reg[465]  ( .D(c[473]), .CLK(clk), .RST(rst), .Q(sreg[465]) );
  DFF \sreg_reg[464]  ( .D(c[472]), .CLK(clk), .RST(rst), .Q(sreg[464]) );
  DFF \sreg_reg[463]  ( .D(c[471]), .CLK(clk), .RST(rst), .Q(sreg[463]) );
  DFF \sreg_reg[462]  ( .D(c[470]), .CLK(clk), .RST(rst), .Q(sreg[462]) );
  DFF \sreg_reg[461]  ( .D(c[469]), .CLK(clk), .RST(rst), .Q(sreg[461]) );
  DFF \sreg_reg[460]  ( .D(c[468]), .CLK(clk), .RST(rst), .Q(sreg[460]) );
  DFF \sreg_reg[459]  ( .D(c[467]), .CLK(clk), .RST(rst), .Q(sreg[459]) );
  DFF \sreg_reg[458]  ( .D(c[466]), .CLK(clk), .RST(rst), .Q(sreg[458]) );
  DFF \sreg_reg[457]  ( .D(c[465]), .CLK(clk), .RST(rst), .Q(sreg[457]) );
  DFF \sreg_reg[456]  ( .D(c[464]), .CLK(clk), .RST(rst), .Q(sreg[456]) );
  DFF \sreg_reg[455]  ( .D(c[463]), .CLK(clk), .RST(rst), .Q(sreg[455]) );
  DFF \sreg_reg[454]  ( .D(c[462]), .CLK(clk), .RST(rst), .Q(sreg[454]) );
  DFF \sreg_reg[453]  ( .D(c[461]), .CLK(clk), .RST(rst), .Q(sreg[453]) );
  DFF \sreg_reg[452]  ( .D(c[460]), .CLK(clk), .RST(rst), .Q(sreg[452]) );
  DFF \sreg_reg[451]  ( .D(c[459]), .CLK(clk), .RST(rst), .Q(sreg[451]) );
  DFF \sreg_reg[450]  ( .D(c[458]), .CLK(clk), .RST(rst), .Q(sreg[450]) );
  DFF \sreg_reg[449]  ( .D(c[457]), .CLK(clk), .RST(rst), .Q(sreg[449]) );
  DFF \sreg_reg[448]  ( .D(c[456]), .CLK(clk), .RST(rst), .Q(sreg[448]) );
  DFF \sreg_reg[447]  ( .D(c[455]), .CLK(clk), .RST(rst), .Q(sreg[447]) );
  DFF \sreg_reg[446]  ( .D(c[454]), .CLK(clk), .RST(rst), .Q(sreg[446]) );
  DFF \sreg_reg[445]  ( .D(c[453]), .CLK(clk), .RST(rst), .Q(sreg[445]) );
  DFF \sreg_reg[444]  ( .D(c[452]), .CLK(clk), .RST(rst), .Q(sreg[444]) );
  DFF \sreg_reg[443]  ( .D(c[451]), .CLK(clk), .RST(rst), .Q(sreg[443]) );
  DFF \sreg_reg[442]  ( .D(c[450]), .CLK(clk), .RST(rst), .Q(sreg[442]) );
  DFF \sreg_reg[441]  ( .D(c[449]), .CLK(clk), .RST(rst), .Q(sreg[441]) );
  DFF \sreg_reg[440]  ( .D(c[448]), .CLK(clk), .RST(rst), .Q(sreg[440]) );
  DFF \sreg_reg[439]  ( .D(c[447]), .CLK(clk), .RST(rst), .Q(sreg[439]) );
  DFF \sreg_reg[438]  ( .D(c[446]), .CLK(clk), .RST(rst), .Q(sreg[438]) );
  DFF \sreg_reg[437]  ( .D(c[445]), .CLK(clk), .RST(rst), .Q(sreg[437]) );
  DFF \sreg_reg[436]  ( .D(c[444]), .CLK(clk), .RST(rst), .Q(sreg[436]) );
  DFF \sreg_reg[435]  ( .D(c[443]), .CLK(clk), .RST(rst), .Q(sreg[435]) );
  DFF \sreg_reg[434]  ( .D(c[442]), .CLK(clk), .RST(rst), .Q(sreg[434]) );
  DFF \sreg_reg[433]  ( .D(c[441]), .CLK(clk), .RST(rst), .Q(sreg[433]) );
  DFF \sreg_reg[432]  ( .D(c[440]), .CLK(clk), .RST(rst), .Q(sreg[432]) );
  DFF \sreg_reg[431]  ( .D(c[439]), .CLK(clk), .RST(rst), .Q(sreg[431]) );
  DFF \sreg_reg[430]  ( .D(c[438]), .CLK(clk), .RST(rst), .Q(sreg[430]) );
  DFF \sreg_reg[429]  ( .D(c[437]), .CLK(clk), .RST(rst), .Q(sreg[429]) );
  DFF \sreg_reg[428]  ( .D(c[436]), .CLK(clk), .RST(rst), .Q(sreg[428]) );
  DFF \sreg_reg[427]  ( .D(c[435]), .CLK(clk), .RST(rst), .Q(sreg[427]) );
  DFF \sreg_reg[426]  ( .D(c[434]), .CLK(clk), .RST(rst), .Q(sreg[426]) );
  DFF \sreg_reg[425]  ( .D(c[433]), .CLK(clk), .RST(rst), .Q(sreg[425]) );
  DFF \sreg_reg[424]  ( .D(c[432]), .CLK(clk), .RST(rst), .Q(sreg[424]) );
  DFF \sreg_reg[423]  ( .D(c[431]), .CLK(clk), .RST(rst), .Q(sreg[423]) );
  DFF \sreg_reg[422]  ( .D(c[430]), .CLK(clk), .RST(rst), .Q(sreg[422]) );
  DFF \sreg_reg[421]  ( .D(c[429]), .CLK(clk), .RST(rst), .Q(sreg[421]) );
  DFF \sreg_reg[420]  ( .D(c[428]), .CLK(clk), .RST(rst), .Q(sreg[420]) );
  DFF \sreg_reg[419]  ( .D(c[427]), .CLK(clk), .RST(rst), .Q(sreg[419]) );
  DFF \sreg_reg[418]  ( .D(c[426]), .CLK(clk), .RST(rst), .Q(sreg[418]) );
  DFF \sreg_reg[417]  ( .D(c[425]), .CLK(clk), .RST(rst), .Q(sreg[417]) );
  DFF \sreg_reg[416]  ( .D(c[424]), .CLK(clk), .RST(rst), .Q(sreg[416]) );
  DFF \sreg_reg[415]  ( .D(c[423]), .CLK(clk), .RST(rst), .Q(sreg[415]) );
  DFF \sreg_reg[414]  ( .D(c[422]), .CLK(clk), .RST(rst), .Q(sreg[414]) );
  DFF \sreg_reg[413]  ( .D(c[421]), .CLK(clk), .RST(rst), .Q(sreg[413]) );
  DFF \sreg_reg[412]  ( .D(c[420]), .CLK(clk), .RST(rst), .Q(sreg[412]) );
  DFF \sreg_reg[411]  ( .D(c[419]), .CLK(clk), .RST(rst), .Q(sreg[411]) );
  DFF \sreg_reg[410]  ( .D(c[418]), .CLK(clk), .RST(rst), .Q(sreg[410]) );
  DFF \sreg_reg[409]  ( .D(c[417]), .CLK(clk), .RST(rst), .Q(sreg[409]) );
  DFF \sreg_reg[408]  ( .D(c[416]), .CLK(clk), .RST(rst), .Q(sreg[408]) );
  DFF \sreg_reg[407]  ( .D(c[415]), .CLK(clk), .RST(rst), .Q(sreg[407]) );
  DFF \sreg_reg[406]  ( .D(c[414]), .CLK(clk), .RST(rst), .Q(sreg[406]) );
  DFF \sreg_reg[405]  ( .D(c[413]), .CLK(clk), .RST(rst), .Q(sreg[405]) );
  DFF \sreg_reg[404]  ( .D(c[412]), .CLK(clk), .RST(rst), .Q(sreg[404]) );
  DFF \sreg_reg[403]  ( .D(c[411]), .CLK(clk), .RST(rst), .Q(sreg[403]) );
  DFF \sreg_reg[402]  ( .D(c[410]), .CLK(clk), .RST(rst), .Q(sreg[402]) );
  DFF \sreg_reg[401]  ( .D(c[409]), .CLK(clk), .RST(rst), .Q(sreg[401]) );
  DFF \sreg_reg[400]  ( .D(c[408]), .CLK(clk), .RST(rst), .Q(sreg[400]) );
  DFF \sreg_reg[399]  ( .D(c[407]), .CLK(clk), .RST(rst), .Q(sreg[399]) );
  DFF \sreg_reg[398]  ( .D(c[406]), .CLK(clk), .RST(rst), .Q(sreg[398]) );
  DFF \sreg_reg[397]  ( .D(c[405]), .CLK(clk), .RST(rst), .Q(sreg[397]) );
  DFF \sreg_reg[396]  ( .D(c[404]), .CLK(clk), .RST(rst), .Q(sreg[396]) );
  DFF \sreg_reg[395]  ( .D(c[403]), .CLK(clk), .RST(rst), .Q(sreg[395]) );
  DFF \sreg_reg[394]  ( .D(c[402]), .CLK(clk), .RST(rst), .Q(sreg[394]) );
  DFF \sreg_reg[393]  ( .D(c[401]), .CLK(clk), .RST(rst), .Q(sreg[393]) );
  DFF \sreg_reg[392]  ( .D(c[400]), .CLK(clk), .RST(rst), .Q(sreg[392]) );
  DFF \sreg_reg[391]  ( .D(c[399]), .CLK(clk), .RST(rst), .Q(sreg[391]) );
  DFF \sreg_reg[390]  ( .D(c[398]), .CLK(clk), .RST(rst), .Q(sreg[390]) );
  DFF \sreg_reg[389]  ( .D(c[397]), .CLK(clk), .RST(rst), .Q(sreg[389]) );
  DFF \sreg_reg[388]  ( .D(c[396]), .CLK(clk), .RST(rst), .Q(sreg[388]) );
  DFF \sreg_reg[387]  ( .D(c[395]), .CLK(clk), .RST(rst), .Q(sreg[387]) );
  DFF \sreg_reg[386]  ( .D(c[394]), .CLK(clk), .RST(rst), .Q(sreg[386]) );
  DFF \sreg_reg[385]  ( .D(c[393]), .CLK(clk), .RST(rst), .Q(sreg[385]) );
  DFF \sreg_reg[384]  ( .D(c[392]), .CLK(clk), .RST(rst), .Q(sreg[384]) );
  DFF \sreg_reg[383]  ( .D(c[391]), .CLK(clk), .RST(rst), .Q(sreg[383]) );
  DFF \sreg_reg[382]  ( .D(c[390]), .CLK(clk), .RST(rst), .Q(sreg[382]) );
  DFF \sreg_reg[381]  ( .D(c[389]), .CLK(clk), .RST(rst), .Q(sreg[381]) );
  DFF \sreg_reg[380]  ( .D(c[388]), .CLK(clk), .RST(rst), .Q(sreg[380]) );
  DFF \sreg_reg[379]  ( .D(c[387]), .CLK(clk), .RST(rst), .Q(sreg[379]) );
  DFF \sreg_reg[378]  ( .D(c[386]), .CLK(clk), .RST(rst), .Q(sreg[378]) );
  DFF \sreg_reg[377]  ( .D(c[385]), .CLK(clk), .RST(rst), .Q(sreg[377]) );
  DFF \sreg_reg[376]  ( .D(c[384]), .CLK(clk), .RST(rst), .Q(sreg[376]) );
  DFF \sreg_reg[375]  ( .D(c[383]), .CLK(clk), .RST(rst), .Q(sreg[375]) );
  DFF \sreg_reg[374]  ( .D(c[382]), .CLK(clk), .RST(rst), .Q(sreg[374]) );
  DFF \sreg_reg[373]  ( .D(c[381]), .CLK(clk), .RST(rst), .Q(sreg[373]) );
  DFF \sreg_reg[372]  ( .D(c[380]), .CLK(clk), .RST(rst), .Q(sreg[372]) );
  DFF \sreg_reg[371]  ( .D(c[379]), .CLK(clk), .RST(rst), .Q(sreg[371]) );
  DFF \sreg_reg[370]  ( .D(c[378]), .CLK(clk), .RST(rst), .Q(sreg[370]) );
  DFF \sreg_reg[369]  ( .D(c[377]), .CLK(clk), .RST(rst), .Q(sreg[369]) );
  DFF \sreg_reg[368]  ( .D(c[376]), .CLK(clk), .RST(rst), .Q(sreg[368]) );
  DFF \sreg_reg[367]  ( .D(c[375]), .CLK(clk), .RST(rst), .Q(sreg[367]) );
  DFF \sreg_reg[366]  ( .D(c[374]), .CLK(clk), .RST(rst), .Q(sreg[366]) );
  DFF \sreg_reg[365]  ( .D(c[373]), .CLK(clk), .RST(rst), .Q(sreg[365]) );
  DFF \sreg_reg[364]  ( .D(c[372]), .CLK(clk), .RST(rst), .Q(sreg[364]) );
  DFF \sreg_reg[363]  ( .D(c[371]), .CLK(clk), .RST(rst), .Q(sreg[363]) );
  DFF \sreg_reg[362]  ( .D(c[370]), .CLK(clk), .RST(rst), .Q(sreg[362]) );
  DFF \sreg_reg[361]  ( .D(c[369]), .CLK(clk), .RST(rst), .Q(sreg[361]) );
  DFF \sreg_reg[360]  ( .D(c[368]), .CLK(clk), .RST(rst), .Q(sreg[360]) );
  DFF \sreg_reg[359]  ( .D(c[367]), .CLK(clk), .RST(rst), .Q(sreg[359]) );
  DFF \sreg_reg[358]  ( .D(c[366]), .CLK(clk), .RST(rst), .Q(sreg[358]) );
  DFF \sreg_reg[357]  ( .D(c[365]), .CLK(clk), .RST(rst), .Q(sreg[357]) );
  DFF \sreg_reg[356]  ( .D(c[364]), .CLK(clk), .RST(rst), .Q(sreg[356]) );
  DFF \sreg_reg[355]  ( .D(c[363]), .CLK(clk), .RST(rst), .Q(sreg[355]) );
  DFF \sreg_reg[354]  ( .D(c[362]), .CLK(clk), .RST(rst), .Q(sreg[354]) );
  DFF \sreg_reg[353]  ( .D(c[361]), .CLK(clk), .RST(rst), .Q(sreg[353]) );
  DFF \sreg_reg[352]  ( .D(c[360]), .CLK(clk), .RST(rst), .Q(sreg[352]) );
  DFF \sreg_reg[351]  ( .D(c[359]), .CLK(clk), .RST(rst), .Q(sreg[351]) );
  DFF \sreg_reg[350]  ( .D(c[358]), .CLK(clk), .RST(rst), .Q(sreg[350]) );
  DFF \sreg_reg[349]  ( .D(c[357]), .CLK(clk), .RST(rst), .Q(sreg[349]) );
  DFF \sreg_reg[348]  ( .D(c[356]), .CLK(clk), .RST(rst), .Q(sreg[348]) );
  DFF \sreg_reg[347]  ( .D(c[355]), .CLK(clk), .RST(rst), .Q(sreg[347]) );
  DFF \sreg_reg[346]  ( .D(c[354]), .CLK(clk), .RST(rst), .Q(sreg[346]) );
  DFF \sreg_reg[345]  ( .D(c[353]), .CLK(clk), .RST(rst), .Q(sreg[345]) );
  DFF \sreg_reg[344]  ( .D(c[352]), .CLK(clk), .RST(rst), .Q(sreg[344]) );
  DFF \sreg_reg[343]  ( .D(c[351]), .CLK(clk), .RST(rst), .Q(sreg[343]) );
  DFF \sreg_reg[342]  ( .D(c[350]), .CLK(clk), .RST(rst), .Q(sreg[342]) );
  DFF \sreg_reg[341]  ( .D(c[349]), .CLK(clk), .RST(rst), .Q(sreg[341]) );
  DFF \sreg_reg[340]  ( .D(c[348]), .CLK(clk), .RST(rst), .Q(sreg[340]) );
  DFF \sreg_reg[339]  ( .D(c[347]), .CLK(clk), .RST(rst), .Q(sreg[339]) );
  DFF \sreg_reg[338]  ( .D(c[346]), .CLK(clk), .RST(rst), .Q(sreg[338]) );
  DFF \sreg_reg[337]  ( .D(c[345]), .CLK(clk), .RST(rst), .Q(sreg[337]) );
  DFF \sreg_reg[336]  ( .D(c[344]), .CLK(clk), .RST(rst), .Q(sreg[336]) );
  DFF \sreg_reg[335]  ( .D(c[343]), .CLK(clk), .RST(rst), .Q(sreg[335]) );
  DFF \sreg_reg[334]  ( .D(c[342]), .CLK(clk), .RST(rst), .Q(sreg[334]) );
  DFF \sreg_reg[333]  ( .D(c[341]), .CLK(clk), .RST(rst), .Q(sreg[333]) );
  DFF \sreg_reg[332]  ( .D(c[340]), .CLK(clk), .RST(rst), .Q(sreg[332]) );
  DFF \sreg_reg[331]  ( .D(c[339]), .CLK(clk), .RST(rst), .Q(sreg[331]) );
  DFF \sreg_reg[330]  ( .D(c[338]), .CLK(clk), .RST(rst), .Q(sreg[330]) );
  DFF \sreg_reg[329]  ( .D(c[337]), .CLK(clk), .RST(rst), .Q(sreg[329]) );
  DFF \sreg_reg[328]  ( .D(c[336]), .CLK(clk), .RST(rst), .Q(sreg[328]) );
  DFF \sreg_reg[327]  ( .D(c[335]), .CLK(clk), .RST(rst), .Q(sreg[327]) );
  DFF \sreg_reg[326]  ( .D(c[334]), .CLK(clk), .RST(rst), .Q(sreg[326]) );
  DFF \sreg_reg[325]  ( .D(c[333]), .CLK(clk), .RST(rst), .Q(sreg[325]) );
  DFF \sreg_reg[324]  ( .D(c[332]), .CLK(clk), .RST(rst), .Q(sreg[324]) );
  DFF \sreg_reg[323]  ( .D(c[331]), .CLK(clk), .RST(rst), .Q(sreg[323]) );
  DFF \sreg_reg[322]  ( .D(c[330]), .CLK(clk), .RST(rst), .Q(sreg[322]) );
  DFF \sreg_reg[321]  ( .D(c[329]), .CLK(clk), .RST(rst), .Q(sreg[321]) );
  DFF \sreg_reg[320]  ( .D(c[328]), .CLK(clk), .RST(rst), .Q(sreg[320]) );
  DFF \sreg_reg[319]  ( .D(c[327]), .CLK(clk), .RST(rst), .Q(sreg[319]) );
  DFF \sreg_reg[318]  ( .D(c[326]), .CLK(clk), .RST(rst), .Q(sreg[318]) );
  DFF \sreg_reg[317]  ( .D(c[325]), .CLK(clk), .RST(rst), .Q(sreg[317]) );
  DFF \sreg_reg[316]  ( .D(c[324]), .CLK(clk), .RST(rst), .Q(sreg[316]) );
  DFF \sreg_reg[315]  ( .D(c[323]), .CLK(clk), .RST(rst), .Q(sreg[315]) );
  DFF \sreg_reg[314]  ( .D(c[322]), .CLK(clk), .RST(rst), .Q(sreg[314]) );
  DFF \sreg_reg[313]  ( .D(c[321]), .CLK(clk), .RST(rst), .Q(sreg[313]) );
  DFF \sreg_reg[312]  ( .D(c[320]), .CLK(clk), .RST(rst), .Q(sreg[312]) );
  DFF \sreg_reg[311]  ( .D(c[319]), .CLK(clk), .RST(rst), .Q(sreg[311]) );
  DFF \sreg_reg[310]  ( .D(c[318]), .CLK(clk), .RST(rst), .Q(sreg[310]) );
  DFF \sreg_reg[309]  ( .D(c[317]), .CLK(clk), .RST(rst), .Q(sreg[309]) );
  DFF \sreg_reg[308]  ( .D(c[316]), .CLK(clk), .RST(rst), .Q(sreg[308]) );
  DFF \sreg_reg[307]  ( .D(c[315]), .CLK(clk), .RST(rst), .Q(sreg[307]) );
  DFF \sreg_reg[306]  ( .D(c[314]), .CLK(clk), .RST(rst), .Q(sreg[306]) );
  DFF \sreg_reg[305]  ( .D(c[313]), .CLK(clk), .RST(rst), .Q(sreg[305]) );
  DFF \sreg_reg[304]  ( .D(c[312]), .CLK(clk), .RST(rst), .Q(sreg[304]) );
  DFF \sreg_reg[303]  ( .D(c[311]), .CLK(clk), .RST(rst), .Q(sreg[303]) );
  DFF \sreg_reg[302]  ( .D(c[310]), .CLK(clk), .RST(rst), .Q(sreg[302]) );
  DFF \sreg_reg[301]  ( .D(c[309]), .CLK(clk), .RST(rst), .Q(sreg[301]) );
  DFF \sreg_reg[300]  ( .D(c[308]), .CLK(clk), .RST(rst), .Q(sreg[300]) );
  DFF \sreg_reg[299]  ( .D(c[307]), .CLK(clk), .RST(rst), .Q(sreg[299]) );
  DFF \sreg_reg[298]  ( .D(c[306]), .CLK(clk), .RST(rst), .Q(sreg[298]) );
  DFF \sreg_reg[297]  ( .D(c[305]), .CLK(clk), .RST(rst), .Q(sreg[297]) );
  DFF \sreg_reg[296]  ( .D(c[304]), .CLK(clk), .RST(rst), .Q(sreg[296]) );
  DFF \sreg_reg[295]  ( .D(c[303]), .CLK(clk), .RST(rst), .Q(sreg[295]) );
  DFF \sreg_reg[294]  ( .D(c[302]), .CLK(clk), .RST(rst), .Q(sreg[294]) );
  DFF \sreg_reg[293]  ( .D(c[301]), .CLK(clk), .RST(rst), .Q(sreg[293]) );
  DFF \sreg_reg[292]  ( .D(c[300]), .CLK(clk), .RST(rst), .Q(sreg[292]) );
  DFF \sreg_reg[291]  ( .D(c[299]), .CLK(clk), .RST(rst), .Q(sreg[291]) );
  DFF \sreg_reg[290]  ( .D(c[298]), .CLK(clk), .RST(rst), .Q(sreg[290]) );
  DFF \sreg_reg[289]  ( .D(c[297]), .CLK(clk), .RST(rst), .Q(sreg[289]) );
  DFF \sreg_reg[288]  ( .D(c[296]), .CLK(clk), .RST(rst), .Q(sreg[288]) );
  DFF \sreg_reg[287]  ( .D(c[295]), .CLK(clk), .RST(rst), .Q(sreg[287]) );
  DFF \sreg_reg[286]  ( .D(c[294]), .CLK(clk), .RST(rst), .Q(sreg[286]) );
  DFF \sreg_reg[285]  ( .D(c[293]), .CLK(clk), .RST(rst), .Q(sreg[285]) );
  DFF \sreg_reg[284]  ( .D(c[292]), .CLK(clk), .RST(rst), .Q(sreg[284]) );
  DFF \sreg_reg[283]  ( .D(c[291]), .CLK(clk), .RST(rst), .Q(sreg[283]) );
  DFF \sreg_reg[282]  ( .D(c[290]), .CLK(clk), .RST(rst), .Q(sreg[282]) );
  DFF \sreg_reg[281]  ( .D(c[289]), .CLK(clk), .RST(rst), .Q(sreg[281]) );
  DFF \sreg_reg[280]  ( .D(c[288]), .CLK(clk), .RST(rst), .Q(sreg[280]) );
  DFF \sreg_reg[279]  ( .D(c[287]), .CLK(clk), .RST(rst), .Q(sreg[279]) );
  DFF \sreg_reg[278]  ( .D(c[286]), .CLK(clk), .RST(rst), .Q(sreg[278]) );
  DFF \sreg_reg[277]  ( .D(c[285]), .CLK(clk), .RST(rst), .Q(sreg[277]) );
  DFF \sreg_reg[276]  ( .D(c[284]), .CLK(clk), .RST(rst), .Q(sreg[276]) );
  DFF \sreg_reg[275]  ( .D(c[283]), .CLK(clk), .RST(rst), .Q(sreg[275]) );
  DFF \sreg_reg[274]  ( .D(c[282]), .CLK(clk), .RST(rst), .Q(sreg[274]) );
  DFF \sreg_reg[273]  ( .D(c[281]), .CLK(clk), .RST(rst), .Q(sreg[273]) );
  DFF \sreg_reg[272]  ( .D(c[280]), .CLK(clk), .RST(rst), .Q(sreg[272]) );
  DFF \sreg_reg[271]  ( .D(c[279]), .CLK(clk), .RST(rst), .Q(sreg[271]) );
  DFF \sreg_reg[270]  ( .D(c[278]), .CLK(clk), .RST(rst), .Q(sreg[270]) );
  DFF \sreg_reg[269]  ( .D(c[277]), .CLK(clk), .RST(rst), .Q(sreg[269]) );
  DFF \sreg_reg[268]  ( .D(c[276]), .CLK(clk), .RST(rst), .Q(sreg[268]) );
  DFF \sreg_reg[267]  ( .D(c[275]), .CLK(clk), .RST(rst), .Q(sreg[267]) );
  DFF \sreg_reg[266]  ( .D(c[274]), .CLK(clk), .RST(rst), .Q(sreg[266]) );
  DFF \sreg_reg[265]  ( .D(c[273]), .CLK(clk), .RST(rst), .Q(sreg[265]) );
  DFF \sreg_reg[264]  ( .D(c[272]), .CLK(clk), .RST(rst), .Q(sreg[264]) );
  DFF \sreg_reg[263]  ( .D(c[271]), .CLK(clk), .RST(rst), .Q(sreg[263]) );
  DFF \sreg_reg[262]  ( .D(c[270]), .CLK(clk), .RST(rst), .Q(sreg[262]) );
  DFF \sreg_reg[261]  ( .D(c[269]), .CLK(clk), .RST(rst), .Q(sreg[261]) );
  DFF \sreg_reg[260]  ( .D(c[268]), .CLK(clk), .RST(rst), .Q(sreg[260]) );
  DFF \sreg_reg[259]  ( .D(c[267]), .CLK(clk), .RST(rst), .Q(sreg[259]) );
  DFF \sreg_reg[258]  ( .D(c[266]), .CLK(clk), .RST(rst), .Q(sreg[258]) );
  DFF \sreg_reg[257]  ( .D(c[265]), .CLK(clk), .RST(rst), .Q(sreg[257]) );
  DFF \sreg_reg[256]  ( .D(c[264]), .CLK(clk), .RST(rst), .Q(sreg[256]) );
  DFF \sreg_reg[255]  ( .D(c[263]), .CLK(clk), .RST(rst), .Q(sreg[255]) );
  DFF \sreg_reg[254]  ( .D(c[262]), .CLK(clk), .RST(rst), .Q(sreg[254]) );
  DFF \sreg_reg[253]  ( .D(c[261]), .CLK(clk), .RST(rst), .Q(sreg[253]) );
  DFF \sreg_reg[252]  ( .D(c[260]), .CLK(clk), .RST(rst), .Q(sreg[252]) );
  DFF \sreg_reg[251]  ( .D(c[259]), .CLK(clk), .RST(rst), .Q(sreg[251]) );
  DFF \sreg_reg[250]  ( .D(c[258]), .CLK(clk), .RST(rst), .Q(sreg[250]) );
  DFF \sreg_reg[249]  ( .D(c[257]), .CLK(clk), .RST(rst), .Q(sreg[249]) );
  DFF \sreg_reg[248]  ( .D(c[256]), .CLK(clk), .RST(rst), .Q(sreg[248]) );
  DFF \sreg_reg[247]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(c[247]) );
  DFF \sreg_reg[246]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(c[246]) );
  DFF \sreg_reg[245]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(c[245]) );
  DFF \sreg_reg[244]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(c[244]) );
  DFF \sreg_reg[243]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(c[243]) );
  DFF \sreg_reg[242]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(c[242]) );
  DFF \sreg_reg[241]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(c[241]) );
  DFF \sreg_reg[240]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(c[240]) );
  DFF \sreg_reg[239]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(c[239]) );
  DFF \sreg_reg[238]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(c[238]) );
  DFF \sreg_reg[237]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(c[237]) );
  DFF \sreg_reg[236]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(c[236]) );
  DFF \sreg_reg[235]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(c[235]) );
  DFF \sreg_reg[234]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(c[234]) );
  DFF \sreg_reg[233]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(c[233]) );
  DFF \sreg_reg[232]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(c[232]) );
  DFF \sreg_reg[231]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(c[231]) );
  DFF \sreg_reg[230]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(c[230]) );
  DFF \sreg_reg[229]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(c[229]) );
  DFF \sreg_reg[228]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(c[228]) );
  DFF \sreg_reg[227]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(c[227]) );
  DFF \sreg_reg[226]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(c[226]) );
  DFF \sreg_reg[225]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(c[225]) );
  DFF \sreg_reg[224]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(c[224]) );
  DFF \sreg_reg[223]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(c[223]) );
  DFF \sreg_reg[222]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(c[222]) );
  DFF \sreg_reg[221]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(c[221]) );
  DFF \sreg_reg[220]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(c[220]) );
  DFF \sreg_reg[219]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(c[219]) );
  DFF \sreg_reg[218]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(c[218]) );
  DFF \sreg_reg[217]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(c[217]) );
  DFF \sreg_reg[216]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(c[216]) );
  DFF \sreg_reg[215]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(c[215]) );
  DFF \sreg_reg[214]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(c[214]) );
  DFF \sreg_reg[213]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(c[213]) );
  DFF \sreg_reg[212]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(c[212]) );
  DFF \sreg_reg[211]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(c[211]) );
  DFF \sreg_reg[210]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(c[210]) );
  DFF \sreg_reg[209]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(c[209]) );
  DFF \sreg_reg[208]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(c[208]) );
  DFF \sreg_reg[207]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(c[207]) );
  DFF \sreg_reg[206]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(c[206]) );
  DFF \sreg_reg[205]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(c[205]) );
  DFF \sreg_reg[204]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(c[204]) );
  DFF \sreg_reg[203]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(c[203]) );
  DFF \sreg_reg[202]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(c[202]) );
  DFF \sreg_reg[201]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(c[201]) );
  DFF \sreg_reg[200]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(c[200]) );
  DFF \sreg_reg[199]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(c[199]) );
  DFF \sreg_reg[198]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(c[198]) );
  DFF \sreg_reg[197]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(c[197]) );
  DFF \sreg_reg[196]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(c[196]) );
  DFF \sreg_reg[195]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(c[195]) );
  DFF \sreg_reg[194]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(c[194]) );
  DFF \sreg_reg[193]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(c[193]) );
  DFF \sreg_reg[192]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(c[192]) );
  DFF \sreg_reg[191]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(c[191]) );
  DFF \sreg_reg[190]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(c[190]) );
  DFF \sreg_reg[189]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(c[189]) );
  DFF \sreg_reg[188]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(c[188]) );
  DFF \sreg_reg[187]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(c[187]) );
  DFF \sreg_reg[186]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(c[186]) );
  DFF \sreg_reg[185]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(c[185]) );
  DFF \sreg_reg[184]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(c[184]) );
  DFF \sreg_reg[183]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(c[183]) );
  DFF \sreg_reg[182]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(c[182]) );
  DFF \sreg_reg[181]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(c[181]) );
  DFF \sreg_reg[180]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(c[180]) );
  DFF \sreg_reg[179]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(c[179]) );
  DFF \sreg_reg[178]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(c[178]) );
  DFF \sreg_reg[177]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(c[177]) );
  DFF \sreg_reg[176]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(c[176]) );
  DFF \sreg_reg[175]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(c[175]) );
  DFF \sreg_reg[174]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(c[174]) );
  DFF \sreg_reg[173]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(c[173]) );
  DFF \sreg_reg[172]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(c[172]) );
  DFF \sreg_reg[171]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(c[171]) );
  DFF \sreg_reg[170]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(c[170]) );
  DFF \sreg_reg[169]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(c[169]) );
  DFF \sreg_reg[168]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(c[168]) );
  DFF \sreg_reg[167]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(c[167]) );
  DFF \sreg_reg[166]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(c[166]) );
  DFF \sreg_reg[165]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(c[165]) );
  DFF \sreg_reg[164]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(c[164]) );
  DFF \sreg_reg[163]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(c[163]) );
  DFF \sreg_reg[162]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(c[162]) );
  DFF \sreg_reg[161]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(c[161]) );
  DFF \sreg_reg[160]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(c[160]) );
  DFF \sreg_reg[159]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(c[159]) );
  DFF \sreg_reg[158]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(c[158]) );
  DFF \sreg_reg[157]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(c[157]) );
  DFF \sreg_reg[156]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(c[156]) );
  DFF \sreg_reg[155]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(c[155]) );
  DFF \sreg_reg[154]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(c[154]) );
  DFF \sreg_reg[153]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(c[153]) );
  DFF \sreg_reg[152]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(c[152]) );
  DFF \sreg_reg[151]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(c[151]) );
  DFF \sreg_reg[150]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(c[150]) );
  DFF \sreg_reg[149]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(c[149]) );
  DFF \sreg_reg[148]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(c[148]) );
  DFF \sreg_reg[147]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(c[147]) );
  DFF \sreg_reg[146]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(c[146]) );
  DFF \sreg_reg[145]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(c[145]) );
  DFF \sreg_reg[144]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(c[144]) );
  DFF \sreg_reg[143]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(c[143]) );
  DFF \sreg_reg[142]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(c[142]) );
  DFF \sreg_reg[141]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(c[141]) );
  DFF \sreg_reg[140]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(c[140]) );
  DFF \sreg_reg[139]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(c[139]) );
  DFF \sreg_reg[138]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(c[138]) );
  DFF \sreg_reg[137]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(c[137]) );
  DFF \sreg_reg[136]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(c[136]) );
  DFF \sreg_reg[135]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(c[135]) );
  DFF \sreg_reg[134]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(c[134]) );
  DFF \sreg_reg[133]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(c[133]) );
  DFF \sreg_reg[132]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(c[132]) );
  DFF \sreg_reg[131]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(c[131]) );
  DFF \sreg_reg[130]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(c[130]) );
  DFF \sreg_reg[129]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(c[129]) );
  DFF \sreg_reg[128]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(c[128]) );
  DFF \sreg_reg[127]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(c[127]) );
  DFF \sreg_reg[126]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(c[126]) );
  DFF \sreg_reg[125]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(c[125]) );
  DFF \sreg_reg[124]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(c[124]) );
  DFF \sreg_reg[123]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(c[123]) );
  DFF \sreg_reg[122]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(c[122]) );
  DFF \sreg_reg[121]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(c[121]) );
  DFF \sreg_reg[120]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(c[120]) );
  DFF \sreg_reg[119]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[118]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[117]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[116]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[115]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[114]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[113]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[112]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[111]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[110]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[109]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[108]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[107]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[106]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[105]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[104]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[103]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[102]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[101]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[100]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[99]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[98]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[97]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[96]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[95]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[94]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[93]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[92]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[91]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[90]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[89]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[88]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[87]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[86]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[85]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[84]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[83]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[82]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[81]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[80]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[79]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[78]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[77]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[76]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[75]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[74]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[73]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[72]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[71]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[70]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[69]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[68]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[67]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[66]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[65]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[64]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[63]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[62]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[0]) );
  NAND U11 ( .A(n1179), .B(n1178), .Z(n1) );
  NAND U12 ( .A(n1176), .B(n1177), .Z(n2) );
  NAND U13 ( .A(n1), .B(n2), .Z(n1186) );
  NAND U14 ( .A(n1645), .B(n1644), .Z(n3) );
  NAND U15 ( .A(n1642), .B(n1643), .Z(n4) );
  NAND U16 ( .A(n3), .B(n4), .Z(n1652) );
  NAND U17 ( .A(n2462), .B(n2463), .Z(n5) );
  NANDN U18 ( .A(n2461), .B(n2460), .Z(n6) );
  NAND U19 ( .A(n5), .B(n6), .Z(n2470) );
  NAND U20 ( .A(n8738), .B(n8739), .Z(n7) );
  NANDN U21 ( .A(n8737), .B(n8736), .Z(n8) );
  NAND U22 ( .A(n7), .B(n8), .Z(n8746) );
  XOR U23 ( .A(n10533), .B(n10532), .Z(n9) );
  NANDN U24 ( .A(n10531), .B(n9), .Z(n10) );
  NAND U25 ( .A(n10533), .B(n10532), .Z(n11) );
  AND U26 ( .A(n10), .B(n11), .Z(n10564) );
  NAND U27 ( .A(n2773), .B(n2772), .Z(n12) );
  NAND U28 ( .A(n2770), .B(n2771), .Z(n13) );
  NAND U29 ( .A(n12), .B(n13), .Z(n2780) );
  NAND U30 ( .A(n2811), .B(n2812), .Z(n14) );
  NANDN U31 ( .A(n2810), .B(n2809), .Z(n15) );
  NAND U32 ( .A(n14), .B(n15), .Z(n2819) );
  NAND U33 ( .A(n584), .B(n582), .Z(n16) );
  XOR U34 ( .A(n582), .B(n584), .Z(n17) );
  NANDN U35 ( .A(n583), .B(n17), .Z(n18) );
  NAND U36 ( .A(n16), .B(n18), .Z(n612) );
  NAND U37 ( .A(n916), .B(n917), .Z(n19) );
  NANDN U38 ( .A(n915), .B(n914), .Z(n20) );
  NAND U39 ( .A(n19), .B(n20), .Z(n956) );
  NAND U40 ( .A(n1033), .B(n1034), .Z(n21) );
  NANDN U41 ( .A(n1032), .B(n1031), .Z(n22) );
  NAND U42 ( .A(n21), .B(n22), .Z(n1073) );
  NAND U43 ( .A(n1150), .B(n1151), .Z(n23) );
  NANDN U44 ( .A(n1149), .B(n1148), .Z(n24) );
  NAND U45 ( .A(n23), .B(n24), .Z(n1188) );
  NAND U46 ( .A(n1265), .B(n1266), .Z(n25) );
  NANDN U47 ( .A(n1264), .B(n1263), .Z(n26) );
  NAND U48 ( .A(n25), .B(n26), .Z(n1305) );
  NAND U49 ( .A(n1382), .B(n1383), .Z(n27) );
  NANDN U50 ( .A(n1381), .B(n1380), .Z(n28) );
  NAND U51 ( .A(n27), .B(n28), .Z(n1422) );
  NAND U52 ( .A(n1499), .B(n1500), .Z(n29) );
  NANDN U53 ( .A(n1498), .B(n1497), .Z(n30) );
  NAND U54 ( .A(n29), .B(n30), .Z(n1539) );
  NAND U55 ( .A(n1616), .B(n1617), .Z(n31) );
  NANDN U56 ( .A(n1615), .B(n1614), .Z(n32) );
  NAND U57 ( .A(n31), .B(n32), .Z(n1654) );
  NAND U58 ( .A(n1731), .B(n1732), .Z(n33) );
  NANDN U59 ( .A(n1730), .B(n1729), .Z(n34) );
  NAND U60 ( .A(n33), .B(n34), .Z(n1771) );
  NAND U61 ( .A(n1848), .B(n1849), .Z(n35) );
  NANDN U62 ( .A(n1847), .B(n1846), .Z(n36) );
  NAND U63 ( .A(n35), .B(n36), .Z(n1888) );
  NAND U64 ( .A(n1965), .B(n1966), .Z(n37) );
  NANDN U65 ( .A(n1964), .B(n1963), .Z(n38) );
  NAND U66 ( .A(n37), .B(n38), .Z(n2005) );
  NAND U67 ( .A(n2082), .B(n2083), .Z(n39) );
  NANDN U68 ( .A(n2081), .B(n2080), .Z(n40) );
  NAND U69 ( .A(n39), .B(n40), .Z(n2122) );
  NAND U70 ( .A(n2199), .B(n2200), .Z(n41) );
  NANDN U71 ( .A(n2198), .B(n2197), .Z(n42) );
  NAND U72 ( .A(n41), .B(n42), .Z(n2239) );
  NAND U73 ( .A(n2316), .B(n2317), .Z(n43) );
  NANDN U74 ( .A(n2315), .B(n2314), .Z(n44) );
  NAND U75 ( .A(n43), .B(n44), .Z(n2356) );
  NAND U76 ( .A(n2434), .B(n2435), .Z(n45) );
  NANDN U77 ( .A(n2433), .B(n2432), .Z(n46) );
  NAND U78 ( .A(n45), .B(n46), .Z(n2472) );
  NAND U79 ( .A(n2549), .B(n2550), .Z(n47) );
  NANDN U80 ( .A(n2548), .B(n2547), .Z(n48) );
  NAND U81 ( .A(n47), .B(n48), .Z(n2589) );
  NAND U82 ( .A(n2666), .B(n2667), .Z(n49) );
  NANDN U83 ( .A(n2665), .B(n2664), .Z(n50) );
  NAND U84 ( .A(n49), .B(n50), .Z(n2706) );
  NAND U85 ( .A(n2898), .B(n2899), .Z(n51) );
  NANDN U86 ( .A(n2897), .B(n2896), .Z(n52) );
  NAND U87 ( .A(n51), .B(n52), .Z(n2938) );
  NAND U88 ( .A(n3015), .B(n3016), .Z(n53) );
  NANDN U89 ( .A(n3014), .B(n3013), .Z(n54) );
  NAND U90 ( .A(n53), .B(n54), .Z(n3055) );
  NAND U91 ( .A(n3132), .B(n3133), .Z(n55) );
  NANDN U92 ( .A(n3131), .B(n3130), .Z(n56) );
  NAND U93 ( .A(n55), .B(n56), .Z(n3172) );
  NAND U94 ( .A(n3249), .B(n3250), .Z(n57) );
  NANDN U95 ( .A(n3248), .B(n3247), .Z(n58) );
  NAND U96 ( .A(n57), .B(n58), .Z(n3289) );
  NAND U97 ( .A(n3366), .B(n3367), .Z(n59) );
  NANDN U98 ( .A(n3365), .B(n3364), .Z(n60) );
  NAND U99 ( .A(n59), .B(n60), .Z(n3406) );
  NAND U100 ( .A(n3483), .B(n3484), .Z(n61) );
  NANDN U101 ( .A(n3482), .B(n3481), .Z(n62) );
  NAND U102 ( .A(n61), .B(n62), .Z(n3523) );
  NAND U103 ( .A(n3600), .B(n3601), .Z(n63) );
  NANDN U104 ( .A(n3599), .B(n3598), .Z(n64) );
  NAND U105 ( .A(n63), .B(n64), .Z(n3640) );
  NAND U106 ( .A(n3717), .B(n3718), .Z(n65) );
  NANDN U107 ( .A(n3716), .B(n3715), .Z(n66) );
  NAND U108 ( .A(n65), .B(n66), .Z(n3757) );
  NAND U109 ( .A(n3834), .B(n3835), .Z(n67) );
  NANDN U110 ( .A(n3833), .B(n3832), .Z(n68) );
  NAND U111 ( .A(n67), .B(n68), .Z(n3874) );
  NAND U112 ( .A(n3951), .B(n3952), .Z(n69) );
  NANDN U113 ( .A(n3950), .B(n3949), .Z(n70) );
  NAND U114 ( .A(n69), .B(n70), .Z(n3991) );
  NAND U115 ( .A(n4068), .B(n4069), .Z(n71) );
  NANDN U116 ( .A(n4067), .B(n4066), .Z(n72) );
  NAND U117 ( .A(n71), .B(n72), .Z(n4108) );
  NAND U118 ( .A(n4185), .B(n4186), .Z(n73) );
  NANDN U119 ( .A(n4184), .B(n4183), .Z(n74) );
  NAND U120 ( .A(n73), .B(n74), .Z(n4225) );
  NAND U121 ( .A(n4302), .B(n4303), .Z(n75) );
  NANDN U122 ( .A(n4301), .B(n4300), .Z(n76) );
  NAND U123 ( .A(n75), .B(n76), .Z(n4342) );
  NAND U124 ( .A(n4419), .B(n4420), .Z(n77) );
  NANDN U125 ( .A(n4418), .B(n4417), .Z(n78) );
  NAND U126 ( .A(n77), .B(n78), .Z(n4459) );
  NAND U127 ( .A(n4536), .B(n4537), .Z(n79) );
  NANDN U128 ( .A(n4535), .B(n4534), .Z(n80) );
  NAND U129 ( .A(n79), .B(n80), .Z(n4576) );
  NAND U130 ( .A(n4653), .B(n4654), .Z(n81) );
  NANDN U131 ( .A(n4652), .B(n4651), .Z(n82) );
  NAND U132 ( .A(n81), .B(n82), .Z(n4693) );
  NAND U133 ( .A(n4770), .B(n4771), .Z(n83) );
  NANDN U134 ( .A(n4769), .B(n4768), .Z(n84) );
  NAND U135 ( .A(n83), .B(n84), .Z(n4810) );
  NAND U136 ( .A(n4887), .B(n4888), .Z(n85) );
  NANDN U137 ( .A(n4886), .B(n4885), .Z(n86) );
  NAND U138 ( .A(n85), .B(n86), .Z(n4927) );
  NAND U139 ( .A(n5004), .B(n5005), .Z(n87) );
  NANDN U140 ( .A(n5003), .B(n5002), .Z(n88) );
  NAND U141 ( .A(n87), .B(n88), .Z(n5044) );
  NAND U142 ( .A(n5121), .B(n5122), .Z(n89) );
  NANDN U143 ( .A(n5120), .B(n5119), .Z(n90) );
  NAND U144 ( .A(n89), .B(n90), .Z(n5161) );
  NAND U145 ( .A(n5238), .B(n5239), .Z(n91) );
  NANDN U146 ( .A(n5237), .B(n5236), .Z(n92) );
  NAND U147 ( .A(n91), .B(n92), .Z(n5278) );
  NAND U148 ( .A(n5355), .B(n5356), .Z(n93) );
  NANDN U149 ( .A(n5354), .B(n5353), .Z(n94) );
  NAND U150 ( .A(n93), .B(n94), .Z(n5395) );
  NAND U151 ( .A(n5472), .B(n5473), .Z(n95) );
  NANDN U152 ( .A(n5471), .B(n5470), .Z(n96) );
  NAND U153 ( .A(n95), .B(n96), .Z(n5512) );
  NAND U154 ( .A(n5589), .B(n5590), .Z(n97) );
  NANDN U155 ( .A(n5588), .B(n5587), .Z(n98) );
  NAND U156 ( .A(n97), .B(n98), .Z(n5629) );
  NAND U157 ( .A(n5706), .B(n5707), .Z(n99) );
  NANDN U158 ( .A(n5705), .B(n5704), .Z(n100) );
  NAND U159 ( .A(n99), .B(n100), .Z(n5746) );
  NAND U160 ( .A(n5823), .B(n5824), .Z(n101) );
  NANDN U161 ( .A(n5822), .B(n5821), .Z(n102) );
  NAND U162 ( .A(n101), .B(n102), .Z(n5863) );
  NAND U163 ( .A(n5940), .B(n5941), .Z(n103) );
  NANDN U164 ( .A(n5939), .B(n5938), .Z(n104) );
  NAND U165 ( .A(n103), .B(n104), .Z(n5980) );
  NAND U166 ( .A(n6057), .B(n6058), .Z(n105) );
  NANDN U167 ( .A(n6056), .B(n6055), .Z(n106) );
  NAND U168 ( .A(n105), .B(n106), .Z(n6097) );
  NAND U169 ( .A(n6174), .B(n6175), .Z(n107) );
  NANDN U170 ( .A(n6173), .B(n6172), .Z(n108) );
  NAND U171 ( .A(n107), .B(n108), .Z(n6214) );
  NAND U172 ( .A(n6291), .B(n6292), .Z(n109) );
  NANDN U173 ( .A(n6290), .B(n6289), .Z(n110) );
  NAND U174 ( .A(n109), .B(n110), .Z(n6331) );
  NAND U175 ( .A(n6408), .B(n6409), .Z(n111) );
  NANDN U176 ( .A(n6407), .B(n6406), .Z(n112) );
  NAND U177 ( .A(n111), .B(n112), .Z(n6448) );
  NAND U178 ( .A(n6525), .B(n6526), .Z(n113) );
  NANDN U179 ( .A(n6524), .B(n6523), .Z(n114) );
  NAND U180 ( .A(n113), .B(n114), .Z(n6565) );
  NAND U181 ( .A(n6642), .B(n6643), .Z(n115) );
  NANDN U182 ( .A(n6641), .B(n6640), .Z(n116) );
  NAND U183 ( .A(n115), .B(n116), .Z(n6682) );
  NAND U184 ( .A(n6759), .B(n6760), .Z(n117) );
  NANDN U185 ( .A(n6758), .B(n6757), .Z(n118) );
  NAND U186 ( .A(n117), .B(n118), .Z(n6799) );
  NAND U187 ( .A(n6876), .B(n6877), .Z(n119) );
  NANDN U188 ( .A(n6875), .B(n6874), .Z(n120) );
  NAND U189 ( .A(n119), .B(n120), .Z(n6916) );
  NAND U190 ( .A(n6993), .B(n6994), .Z(n121) );
  NANDN U191 ( .A(n6992), .B(n6991), .Z(n122) );
  NAND U192 ( .A(n121), .B(n122), .Z(n7033) );
  NAND U193 ( .A(n7110), .B(n7111), .Z(n123) );
  NANDN U194 ( .A(n7109), .B(n7108), .Z(n124) );
  NAND U195 ( .A(n123), .B(n124), .Z(n7150) );
  NAND U196 ( .A(n7227), .B(n7228), .Z(n125) );
  NANDN U197 ( .A(n7226), .B(n7225), .Z(n126) );
  NAND U198 ( .A(n125), .B(n126), .Z(n7267) );
  NAND U199 ( .A(n7344), .B(n7345), .Z(n127) );
  NANDN U200 ( .A(n7343), .B(n7342), .Z(n128) );
  NAND U201 ( .A(n127), .B(n128), .Z(n7384) );
  NAND U202 ( .A(n7461), .B(n7462), .Z(n129) );
  NANDN U203 ( .A(n7460), .B(n7459), .Z(n130) );
  NAND U204 ( .A(n129), .B(n130), .Z(n7501) );
  NAND U205 ( .A(n7578), .B(n7579), .Z(n131) );
  NANDN U206 ( .A(n7577), .B(n7576), .Z(n132) );
  NAND U207 ( .A(n131), .B(n132), .Z(n7618) );
  NAND U208 ( .A(n7695), .B(n7696), .Z(n133) );
  NANDN U209 ( .A(n7694), .B(n7693), .Z(n134) );
  NAND U210 ( .A(n133), .B(n134), .Z(n7735) );
  NAND U211 ( .A(n7812), .B(n7813), .Z(n135) );
  NANDN U212 ( .A(n7811), .B(n7810), .Z(n136) );
  NAND U213 ( .A(n135), .B(n136), .Z(n7852) );
  NAND U214 ( .A(n7929), .B(n7930), .Z(n137) );
  NANDN U215 ( .A(n7928), .B(n7927), .Z(n138) );
  NAND U216 ( .A(n137), .B(n138), .Z(n7969) );
  NAND U217 ( .A(n8046), .B(n8047), .Z(n139) );
  NANDN U218 ( .A(n8045), .B(n8044), .Z(n140) );
  NAND U219 ( .A(n139), .B(n140), .Z(n8086) );
  NAND U220 ( .A(n8163), .B(n8164), .Z(n141) );
  NANDN U221 ( .A(n8162), .B(n8161), .Z(n142) );
  NAND U222 ( .A(n141), .B(n142), .Z(n8203) );
  NAND U223 ( .A(n8280), .B(n8281), .Z(n143) );
  NANDN U224 ( .A(n8279), .B(n8278), .Z(n144) );
  NAND U225 ( .A(n143), .B(n144), .Z(n8320) );
  NAND U226 ( .A(n8397), .B(n8398), .Z(n145) );
  NANDN U227 ( .A(n8396), .B(n8395), .Z(n146) );
  NAND U228 ( .A(n145), .B(n146), .Z(n8437) );
  NAND U229 ( .A(n8514), .B(n8515), .Z(n147) );
  NANDN U230 ( .A(n8513), .B(n8512), .Z(n148) );
  NAND U231 ( .A(n147), .B(n148), .Z(n8554) );
  NAND U232 ( .A(n8631), .B(n8632), .Z(n149) );
  NANDN U233 ( .A(n8630), .B(n8629), .Z(n150) );
  NAND U234 ( .A(n149), .B(n150), .Z(n8672) );
  NAND U235 ( .A(n8747), .B(n8748), .Z(n151) );
  NANDN U236 ( .A(n8746), .B(n8745), .Z(n152) );
  NAND U237 ( .A(n151), .B(n152), .Z(n8787) );
  NAND U238 ( .A(n8864), .B(n8865), .Z(n153) );
  NANDN U239 ( .A(n8863), .B(n8862), .Z(n154) );
  NAND U240 ( .A(n153), .B(n154), .Z(n8904) );
  NAND U241 ( .A(n8981), .B(n8982), .Z(n155) );
  NANDN U242 ( .A(n8980), .B(n8979), .Z(n156) );
  NAND U243 ( .A(n155), .B(n156), .Z(n9021) );
  NAND U244 ( .A(n9098), .B(n9099), .Z(n157) );
  NANDN U245 ( .A(n9097), .B(n9096), .Z(n158) );
  NAND U246 ( .A(n157), .B(n158), .Z(n9138) );
  NAND U247 ( .A(n9215), .B(n9216), .Z(n159) );
  NANDN U248 ( .A(n9214), .B(n9213), .Z(n160) );
  NAND U249 ( .A(n159), .B(n160), .Z(n9255) );
  NAND U250 ( .A(n9332), .B(n9333), .Z(n161) );
  NANDN U251 ( .A(n9331), .B(n9330), .Z(n162) );
  NAND U252 ( .A(n161), .B(n162), .Z(n9372) );
  NAND U253 ( .A(n9449), .B(n9450), .Z(n163) );
  NANDN U254 ( .A(n9448), .B(n9447), .Z(n164) );
  NAND U255 ( .A(n163), .B(n164), .Z(n9489) );
  NAND U256 ( .A(n9566), .B(n9567), .Z(n165) );
  NANDN U257 ( .A(n9565), .B(n9564), .Z(n166) );
  NAND U258 ( .A(n165), .B(n166), .Z(n9606) );
  NAND U259 ( .A(n9683), .B(n9684), .Z(n167) );
  NANDN U260 ( .A(n9682), .B(n9681), .Z(n168) );
  NAND U261 ( .A(n167), .B(n168), .Z(n9723) );
  NAND U262 ( .A(n9800), .B(n9801), .Z(n169) );
  NANDN U263 ( .A(n9799), .B(n9798), .Z(n170) );
  NAND U264 ( .A(n169), .B(n170), .Z(n9840) );
  NAND U265 ( .A(n9917), .B(n9918), .Z(n171) );
  NANDN U266 ( .A(n9916), .B(n9915), .Z(n172) );
  NAND U267 ( .A(n171), .B(n172), .Z(n9957) );
  NAND U268 ( .A(n10034), .B(n10035), .Z(n173) );
  NANDN U269 ( .A(n10033), .B(n10032), .Z(n174) );
  NAND U270 ( .A(n173), .B(n174), .Z(n10074) );
  NAND U271 ( .A(n10151), .B(n10152), .Z(n175) );
  NANDN U272 ( .A(n10150), .B(n10149), .Z(n176) );
  NAND U273 ( .A(n175), .B(n176), .Z(n10191) );
  NAND U274 ( .A(n10268), .B(n10269), .Z(n177) );
  NANDN U275 ( .A(n10267), .B(n10266), .Z(n178) );
  NAND U276 ( .A(n177), .B(n178), .Z(n10308) );
  XOR U277 ( .A(n10567), .B(n10568), .Z(n10562) );
  NAND U278 ( .A(n838), .B(n839), .Z(n179) );
  NANDN U279 ( .A(n837), .B(n836), .Z(n180) );
  NAND U280 ( .A(n179), .B(n180), .Z(n878) );
  NAND U281 ( .A(n955), .B(n956), .Z(n181) );
  NANDN U282 ( .A(n954), .B(n953), .Z(n182) );
  NAND U283 ( .A(n181), .B(n182), .Z(n995) );
  NAND U284 ( .A(n1072), .B(n1073), .Z(n183) );
  NANDN U285 ( .A(n1071), .B(n1070), .Z(n184) );
  NAND U286 ( .A(n183), .B(n184), .Z(n1112) );
  NAND U287 ( .A(n1187), .B(n1188), .Z(n185) );
  NANDN U288 ( .A(n1186), .B(n1185), .Z(n186) );
  NAND U289 ( .A(n185), .B(n186), .Z(n1227) );
  NAND U290 ( .A(n1304), .B(n1305), .Z(n187) );
  NANDN U291 ( .A(n1303), .B(n1302), .Z(n188) );
  NAND U292 ( .A(n187), .B(n188), .Z(n1344) );
  NAND U293 ( .A(n1421), .B(n1422), .Z(n189) );
  NANDN U294 ( .A(n1420), .B(n1419), .Z(n190) );
  NAND U295 ( .A(n189), .B(n190), .Z(n1461) );
  NAND U296 ( .A(n1538), .B(n1539), .Z(n191) );
  NANDN U297 ( .A(n1537), .B(n1536), .Z(n192) );
  NAND U298 ( .A(n191), .B(n192), .Z(n1578) );
  NAND U299 ( .A(n1653), .B(n1654), .Z(n193) );
  NANDN U300 ( .A(n1652), .B(n1651), .Z(n194) );
  NAND U301 ( .A(n193), .B(n194), .Z(n1693) );
  NAND U302 ( .A(n1770), .B(n1771), .Z(n195) );
  NANDN U303 ( .A(n1769), .B(n1768), .Z(n196) );
  NAND U304 ( .A(n195), .B(n196), .Z(n1810) );
  NAND U305 ( .A(n1887), .B(n1888), .Z(n197) );
  NANDN U306 ( .A(n1886), .B(n1885), .Z(n198) );
  NAND U307 ( .A(n197), .B(n198), .Z(n1927) );
  NAND U308 ( .A(n2004), .B(n2005), .Z(n199) );
  NANDN U309 ( .A(n2003), .B(n2002), .Z(n200) );
  NAND U310 ( .A(n199), .B(n200), .Z(n2044) );
  NAND U311 ( .A(n2121), .B(n2122), .Z(n201) );
  NANDN U312 ( .A(n2120), .B(n2119), .Z(n202) );
  NAND U313 ( .A(n201), .B(n202), .Z(n2161) );
  NAND U314 ( .A(n2238), .B(n2239), .Z(n203) );
  NANDN U315 ( .A(n2237), .B(n2236), .Z(n204) );
  NAND U316 ( .A(n203), .B(n204), .Z(n2278) );
  NAND U317 ( .A(n2355), .B(n2356), .Z(n205) );
  NANDN U318 ( .A(n2354), .B(n2353), .Z(n206) );
  NAND U319 ( .A(n205), .B(n206), .Z(n2396) );
  NAND U320 ( .A(n2471), .B(n2472), .Z(n207) );
  NANDN U321 ( .A(n2470), .B(n2469), .Z(n208) );
  NAND U322 ( .A(n207), .B(n208), .Z(n2511) );
  NAND U323 ( .A(n2588), .B(n2589), .Z(n209) );
  NANDN U324 ( .A(n2587), .B(n2586), .Z(n210) );
  NAND U325 ( .A(n209), .B(n210), .Z(n2628) );
  NAND U326 ( .A(n2705), .B(n2706), .Z(n211) );
  NANDN U327 ( .A(n2704), .B(n2703), .Z(n212) );
  NAND U328 ( .A(n211), .B(n212), .Z(n2745) );
  NAND U329 ( .A(n2820), .B(n2821), .Z(n213) );
  NANDN U330 ( .A(n2819), .B(n2818), .Z(n214) );
  NAND U331 ( .A(n213), .B(n214), .Z(n2860) );
  NAND U332 ( .A(n2937), .B(n2938), .Z(n215) );
  NANDN U333 ( .A(n2936), .B(n2935), .Z(n216) );
  NAND U334 ( .A(n215), .B(n216), .Z(n2977) );
  NAND U335 ( .A(n3054), .B(n3055), .Z(n217) );
  NANDN U336 ( .A(n3053), .B(n3052), .Z(n218) );
  NAND U337 ( .A(n217), .B(n218), .Z(n3094) );
  NAND U338 ( .A(n3171), .B(n3172), .Z(n219) );
  NANDN U339 ( .A(n3170), .B(n3169), .Z(n220) );
  NAND U340 ( .A(n219), .B(n220), .Z(n3211) );
  NAND U341 ( .A(n3288), .B(n3289), .Z(n221) );
  NANDN U342 ( .A(n3287), .B(n3286), .Z(n222) );
  NAND U343 ( .A(n221), .B(n222), .Z(n3328) );
  NAND U344 ( .A(n3405), .B(n3406), .Z(n223) );
  NANDN U345 ( .A(n3404), .B(n3403), .Z(n224) );
  NAND U346 ( .A(n223), .B(n224), .Z(n3445) );
  NAND U347 ( .A(n3522), .B(n3523), .Z(n225) );
  NANDN U348 ( .A(n3521), .B(n3520), .Z(n226) );
  NAND U349 ( .A(n225), .B(n226), .Z(n3562) );
  NAND U350 ( .A(n3639), .B(n3640), .Z(n227) );
  NANDN U351 ( .A(n3638), .B(n3637), .Z(n228) );
  NAND U352 ( .A(n227), .B(n228), .Z(n3679) );
  NAND U353 ( .A(n3756), .B(n3757), .Z(n229) );
  NANDN U354 ( .A(n3755), .B(n3754), .Z(n230) );
  NAND U355 ( .A(n229), .B(n230), .Z(n3796) );
  NAND U356 ( .A(n3873), .B(n3874), .Z(n231) );
  NANDN U357 ( .A(n3872), .B(n3871), .Z(n232) );
  NAND U358 ( .A(n231), .B(n232), .Z(n3913) );
  NAND U359 ( .A(n3990), .B(n3991), .Z(n233) );
  NANDN U360 ( .A(n3989), .B(n3988), .Z(n234) );
  NAND U361 ( .A(n233), .B(n234), .Z(n4030) );
  NAND U362 ( .A(n4107), .B(n4108), .Z(n235) );
  NANDN U363 ( .A(n4106), .B(n4105), .Z(n236) );
  NAND U364 ( .A(n235), .B(n236), .Z(n4147) );
  NAND U365 ( .A(n4224), .B(n4225), .Z(n237) );
  NANDN U366 ( .A(n4223), .B(n4222), .Z(n238) );
  NAND U367 ( .A(n237), .B(n238), .Z(n4264) );
  NAND U368 ( .A(n4341), .B(n4342), .Z(n239) );
  NANDN U369 ( .A(n4340), .B(n4339), .Z(n240) );
  NAND U370 ( .A(n239), .B(n240), .Z(n4381) );
  NAND U371 ( .A(n4458), .B(n4459), .Z(n241) );
  NANDN U372 ( .A(n4457), .B(n4456), .Z(n242) );
  NAND U373 ( .A(n241), .B(n242), .Z(n4498) );
  NAND U374 ( .A(n4575), .B(n4576), .Z(n243) );
  NANDN U375 ( .A(n4574), .B(n4573), .Z(n244) );
  NAND U376 ( .A(n243), .B(n244), .Z(n4615) );
  NAND U377 ( .A(n4692), .B(n4693), .Z(n245) );
  NANDN U378 ( .A(n4691), .B(n4690), .Z(n246) );
  NAND U379 ( .A(n245), .B(n246), .Z(n4732) );
  NAND U380 ( .A(n4809), .B(n4810), .Z(n247) );
  NANDN U381 ( .A(n4808), .B(n4807), .Z(n248) );
  NAND U382 ( .A(n247), .B(n248), .Z(n4849) );
  NAND U383 ( .A(n4926), .B(n4927), .Z(n249) );
  NANDN U384 ( .A(n4925), .B(n4924), .Z(n250) );
  NAND U385 ( .A(n249), .B(n250), .Z(n4966) );
  NAND U386 ( .A(n5043), .B(n5044), .Z(n251) );
  NANDN U387 ( .A(n5042), .B(n5041), .Z(n252) );
  NAND U388 ( .A(n251), .B(n252), .Z(n5083) );
  NAND U389 ( .A(n5160), .B(n5161), .Z(n253) );
  NANDN U390 ( .A(n5159), .B(n5158), .Z(n254) );
  NAND U391 ( .A(n253), .B(n254), .Z(n5200) );
  NAND U392 ( .A(n5277), .B(n5278), .Z(n255) );
  NANDN U393 ( .A(n5276), .B(n5275), .Z(n256) );
  NAND U394 ( .A(n255), .B(n256), .Z(n5317) );
  NAND U395 ( .A(n5394), .B(n5395), .Z(n257) );
  NANDN U396 ( .A(n5393), .B(n5392), .Z(n258) );
  NAND U397 ( .A(n257), .B(n258), .Z(n5434) );
  NAND U398 ( .A(n5511), .B(n5512), .Z(n259) );
  NANDN U399 ( .A(n5510), .B(n5509), .Z(n260) );
  NAND U400 ( .A(n259), .B(n260), .Z(n5551) );
  NAND U401 ( .A(n5628), .B(n5629), .Z(n261) );
  NANDN U402 ( .A(n5627), .B(n5626), .Z(n262) );
  NAND U403 ( .A(n261), .B(n262), .Z(n5668) );
  NAND U404 ( .A(n5745), .B(n5746), .Z(n263) );
  NANDN U405 ( .A(n5744), .B(n5743), .Z(n264) );
  NAND U406 ( .A(n263), .B(n264), .Z(n5785) );
  NAND U407 ( .A(n5862), .B(n5863), .Z(n265) );
  NANDN U408 ( .A(n5861), .B(n5860), .Z(n266) );
  NAND U409 ( .A(n265), .B(n266), .Z(n5902) );
  NAND U410 ( .A(n5979), .B(n5980), .Z(n267) );
  NANDN U411 ( .A(n5978), .B(n5977), .Z(n268) );
  NAND U412 ( .A(n267), .B(n268), .Z(n6019) );
  NAND U413 ( .A(n6096), .B(n6097), .Z(n269) );
  NANDN U414 ( .A(n6095), .B(n6094), .Z(n270) );
  NAND U415 ( .A(n269), .B(n270), .Z(n6136) );
  NAND U416 ( .A(n6213), .B(n6214), .Z(n271) );
  NANDN U417 ( .A(n6212), .B(n6211), .Z(n272) );
  NAND U418 ( .A(n271), .B(n272), .Z(n6253) );
  NAND U419 ( .A(n6330), .B(n6331), .Z(n273) );
  NANDN U420 ( .A(n6329), .B(n6328), .Z(n274) );
  NAND U421 ( .A(n273), .B(n274), .Z(n6370) );
  NAND U422 ( .A(n6447), .B(n6448), .Z(n275) );
  NANDN U423 ( .A(n6446), .B(n6445), .Z(n276) );
  NAND U424 ( .A(n275), .B(n276), .Z(n6487) );
  NAND U425 ( .A(n6564), .B(n6565), .Z(n277) );
  NANDN U426 ( .A(n6563), .B(n6562), .Z(n278) );
  NAND U427 ( .A(n277), .B(n278), .Z(n6604) );
  NAND U428 ( .A(n6681), .B(n6682), .Z(n279) );
  NANDN U429 ( .A(n6680), .B(n6679), .Z(n280) );
  NAND U430 ( .A(n279), .B(n280), .Z(n6721) );
  NAND U431 ( .A(n6798), .B(n6799), .Z(n281) );
  NANDN U432 ( .A(n6797), .B(n6796), .Z(n282) );
  NAND U433 ( .A(n281), .B(n282), .Z(n6838) );
  NAND U434 ( .A(n6915), .B(n6916), .Z(n283) );
  NANDN U435 ( .A(n6914), .B(n6913), .Z(n284) );
  NAND U436 ( .A(n283), .B(n284), .Z(n6955) );
  NAND U437 ( .A(n7032), .B(n7033), .Z(n285) );
  NANDN U438 ( .A(n7031), .B(n7030), .Z(n286) );
  NAND U439 ( .A(n285), .B(n286), .Z(n7072) );
  NAND U440 ( .A(n7149), .B(n7150), .Z(n287) );
  NANDN U441 ( .A(n7148), .B(n7147), .Z(n288) );
  NAND U442 ( .A(n287), .B(n288), .Z(n7189) );
  NAND U443 ( .A(n7266), .B(n7267), .Z(n289) );
  NANDN U444 ( .A(n7265), .B(n7264), .Z(n290) );
  NAND U445 ( .A(n289), .B(n290), .Z(n7306) );
  NAND U446 ( .A(n7383), .B(n7384), .Z(n291) );
  NANDN U447 ( .A(n7382), .B(n7381), .Z(n292) );
  NAND U448 ( .A(n291), .B(n292), .Z(n7423) );
  NAND U449 ( .A(n7500), .B(n7501), .Z(n293) );
  NANDN U450 ( .A(n7499), .B(n7498), .Z(n294) );
  NAND U451 ( .A(n293), .B(n294), .Z(n7540) );
  NAND U452 ( .A(n7617), .B(n7618), .Z(n295) );
  NANDN U453 ( .A(n7616), .B(n7615), .Z(n296) );
  NAND U454 ( .A(n295), .B(n296), .Z(n7657) );
  NAND U455 ( .A(n7734), .B(n7735), .Z(n297) );
  NANDN U456 ( .A(n7733), .B(n7732), .Z(n298) );
  NAND U457 ( .A(n297), .B(n298), .Z(n7774) );
  NAND U458 ( .A(n7851), .B(n7852), .Z(n299) );
  NANDN U459 ( .A(n7850), .B(n7849), .Z(n300) );
  NAND U460 ( .A(n299), .B(n300), .Z(n7891) );
  NAND U461 ( .A(n7968), .B(n7969), .Z(n301) );
  NANDN U462 ( .A(n7967), .B(n7966), .Z(n302) );
  NAND U463 ( .A(n301), .B(n302), .Z(n8008) );
  NAND U464 ( .A(n8085), .B(n8086), .Z(n303) );
  NANDN U465 ( .A(n8084), .B(n8083), .Z(n304) );
  NAND U466 ( .A(n303), .B(n304), .Z(n8125) );
  NAND U467 ( .A(n8202), .B(n8203), .Z(n305) );
  NANDN U468 ( .A(n8201), .B(n8200), .Z(n306) );
  NAND U469 ( .A(n305), .B(n306), .Z(n8242) );
  NAND U470 ( .A(n8319), .B(n8320), .Z(n307) );
  NANDN U471 ( .A(n8318), .B(n8317), .Z(n308) );
  NAND U472 ( .A(n307), .B(n308), .Z(n8359) );
  NAND U473 ( .A(n8436), .B(n8437), .Z(n309) );
  NANDN U474 ( .A(n8435), .B(n8434), .Z(n310) );
  NAND U475 ( .A(n309), .B(n310), .Z(n8476) );
  NAND U476 ( .A(n8553), .B(n8554), .Z(n311) );
  NANDN U477 ( .A(n8552), .B(n8551), .Z(n312) );
  NAND U478 ( .A(n311), .B(n312), .Z(n8593) );
  NAND U479 ( .A(n8671), .B(n8672), .Z(n313) );
  NANDN U480 ( .A(n8670), .B(n8669), .Z(n314) );
  NAND U481 ( .A(n313), .B(n314), .Z(n8711) );
  NAND U482 ( .A(n8786), .B(n8787), .Z(n315) );
  NANDN U483 ( .A(n8785), .B(n8784), .Z(n316) );
  NAND U484 ( .A(n315), .B(n316), .Z(n8826) );
  NAND U485 ( .A(n8903), .B(n8904), .Z(n317) );
  NANDN U486 ( .A(n8902), .B(n8901), .Z(n318) );
  NAND U487 ( .A(n317), .B(n318), .Z(n8943) );
  NAND U488 ( .A(n9020), .B(n9021), .Z(n319) );
  NANDN U489 ( .A(n9019), .B(n9018), .Z(n320) );
  NAND U490 ( .A(n319), .B(n320), .Z(n9060) );
  NAND U491 ( .A(n9137), .B(n9138), .Z(n321) );
  NANDN U492 ( .A(n9136), .B(n9135), .Z(n322) );
  NAND U493 ( .A(n321), .B(n322), .Z(n9177) );
  NAND U494 ( .A(n9254), .B(n9255), .Z(n323) );
  NANDN U495 ( .A(n9253), .B(n9252), .Z(n324) );
  NAND U496 ( .A(n323), .B(n324), .Z(n9294) );
  NAND U497 ( .A(n9371), .B(n9372), .Z(n325) );
  NANDN U498 ( .A(n9370), .B(n9369), .Z(n326) );
  NAND U499 ( .A(n325), .B(n326), .Z(n9411) );
  NAND U500 ( .A(n9488), .B(n9489), .Z(n327) );
  NANDN U501 ( .A(n9487), .B(n9486), .Z(n328) );
  NAND U502 ( .A(n327), .B(n328), .Z(n9528) );
  NAND U503 ( .A(n9605), .B(n9606), .Z(n329) );
  NANDN U504 ( .A(n9604), .B(n9603), .Z(n330) );
  NAND U505 ( .A(n329), .B(n330), .Z(n9645) );
  NAND U506 ( .A(n9722), .B(n9723), .Z(n331) );
  NANDN U507 ( .A(n9721), .B(n9720), .Z(n332) );
  NAND U508 ( .A(n331), .B(n332), .Z(n9762) );
  NAND U509 ( .A(n9839), .B(n9840), .Z(n333) );
  NANDN U510 ( .A(n9838), .B(n9837), .Z(n334) );
  NAND U511 ( .A(n333), .B(n334), .Z(n9879) );
  NAND U512 ( .A(n9956), .B(n9957), .Z(n335) );
  NANDN U513 ( .A(n9955), .B(n9954), .Z(n336) );
  NAND U514 ( .A(n335), .B(n336), .Z(n9996) );
  NAND U515 ( .A(n10073), .B(n10074), .Z(n337) );
  NANDN U516 ( .A(n10072), .B(n10071), .Z(n338) );
  NAND U517 ( .A(n337), .B(n338), .Z(n10113) );
  NAND U518 ( .A(n10190), .B(n10191), .Z(n339) );
  NANDN U519 ( .A(n10189), .B(n10188), .Z(n340) );
  NAND U520 ( .A(n339), .B(n340), .Z(n10230) );
  NAND U521 ( .A(n10307), .B(n10308), .Z(n341) );
  NANDN U522 ( .A(n10306), .B(n10305), .Z(n342) );
  NAND U523 ( .A(n341), .B(n342), .Z(n10349) );
  XOR U524 ( .A(n573), .B(n571), .Z(n343) );
  NAND U525 ( .A(n343), .B(n572), .Z(n344) );
  NAND U526 ( .A(n573), .B(n571), .Z(n345) );
  AND U527 ( .A(n344), .B(n345), .Z(n584) );
  XOR U528 ( .A(n10564), .B(n10562), .Z(n346) );
  NANDN U529 ( .A(n10563), .B(n346), .Z(n347) );
  NAND U530 ( .A(n10564), .B(n10562), .Z(n348) );
  AND U531 ( .A(n347), .B(n348), .Z(n10578) );
  XNOR U532 ( .A(n10411), .B(n10412), .Z(n10404) );
  NAND U533 ( .A(n645), .B(n646), .Z(n349) );
  NANDN U534 ( .A(n644), .B(n643), .Z(n350) );
  NAND U535 ( .A(n349), .B(n350), .Z(n689) );
  XOR U536 ( .A(n10471), .B(n10472), .Z(n10474) );
  NAND U537 ( .A(n877), .B(n878), .Z(n351) );
  NANDN U538 ( .A(n876), .B(n875), .Z(n352) );
  NAND U539 ( .A(n351), .B(n352), .Z(n917) );
  NAND U540 ( .A(n994), .B(n995), .Z(n353) );
  NANDN U541 ( .A(n993), .B(n992), .Z(n354) );
  NAND U542 ( .A(n353), .B(n354), .Z(n1034) );
  NAND U543 ( .A(n1111), .B(n1112), .Z(n355) );
  NANDN U544 ( .A(n1110), .B(n1109), .Z(n356) );
  NAND U545 ( .A(n355), .B(n356), .Z(n1151) );
  NAND U546 ( .A(n1226), .B(n1227), .Z(n357) );
  NANDN U547 ( .A(n1225), .B(n1224), .Z(n358) );
  NAND U548 ( .A(n357), .B(n358), .Z(n1266) );
  NAND U549 ( .A(n1343), .B(n1344), .Z(n359) );
  NANDN U550 ( .A(n1342), .B(n1341), .Z(n360) );
  NAND U551 ( .A(n359), .B(n360), .Z(n1383) );
  NAND U552 ( .A(n1460), .B(n1461), .Z(n361) );
  NANDN U553 ( .A(n1459), .B(n1458), .Z(n362) );
  NAND U554 ( .A(n361), .B(n362), .Z(n1500) );
  NAND U555 ( .A(n1577), .B(n1578), .Z(n363) );
  NANDN U556 ( .A(n1576), .B(n1575), .Z(n364) );
  NAND U557 ( .A(n363), .B(n364), .Z(n1617) );
  NAND U558 ( .A(n1692), .B(n1693), .Z(n365) );
  NANDN U559 ( .A(n1691), .B(n1690), .Z(n366) );
  NAND U560 ( .A(n365), .B(n366), .Z(n1732) );
  NAND U561 ( .A(n1809), .B(n1810), .Z(n367) );
  NANDN U562 ( .A(n1808), .B(n1807), .Z(n368) );
  NAND U563 ( .A(n367), .B(n368), .Z(n1849) );
  NAND U564 ( .A(n1926), .B(n1927), .Z(n369) );
  NANDN U565 ( .A(n1925), .B(n1924), .Z(n370) );
  NAND U566 ( .A(n369), .B(n370), .Z(n1966) );
  NAND U567 ( .A(n2043), .B(n2044), .Z(n371) );
  NANDN U568 ( .A(n2042), .B(n2041), .Z(n372) );
  NAND U569 ( .A(n371), .B(n372), .Z(n2083) );
  NAND U570 ( .A(n2160), .B(n2161), .Z(n373) );
  NANDN U571 ( .A(n2159), .B(n2158), .Z(n374) );
  NAND U572 ( .A(n373), .B(n374), .Z(n2200) );
  NAND U573 ( .A(n2277), .B(n2278), .Z(n375) );
  NANDN U574 ( .A(n2276), .B(n2275), .Z(n376) );
  NAND U575 ( .A(n375), .B(n376), .Z(n2317) );
  NAND U576 ( .A(n2395), .B(n2396), .Z(n377) );
  NANDN U577 ( .A(n2394), .B(n2393), .Z(n378) );
  NAND U578 ( .A(n377), .B(n378), .Z(n2435) );
  NAND U579 ( .A(n2510), .B(n2511), .Z(n379) );
  NANDN U580 ( .A(n2509), .B(n2508), .Z(n380) );
  NAND U581 ( .A(n379), .B(n380), .Z(n2550) );
  NAND U582 ( .A(n2627), .B(n2628), .Z(n381) );
  NANDN U583 ( .A(n2626), .B(n2625), .Z(n382) );
  NAND U584 ( .A(n381), .B(n382), .Z(n2667) );
  NAND U585 ( .A(n2744), .B(n2745), .Z(n383) );
  NANDN U586 ( .A(n2743), .B(n2742), .Z(n384) );
  NAND U587 ( .A(n383), .B(n384), .Z(n2782) );
  NAND U588 ( .A(n2859), .B(n2860), .Z(n385) );
  NANDN U589 ( .A(n2858), .B(n2857), .Z(n386) );
  NAND U590 ( .A(n385), .B(n386), .Z(n2899) );
  NAND U591 ( .A(n2976), .B(n2977), .Z(n387) );
  NANDN U592 ( .A(n2975), .B(n2974), .Z(n388) );
  NAND U593 ( .A(n387), .B(n388), .Z(n3016) );
  NAND U594 ( .A(n3093), .B(n3094), .Z(n389) );
  NANDN U595 ( .A(n3092), .B(n3091), .Z(n390) );
  NAND U596 ( .A(n389), .B(n390), .Z(n3133) );
  NAND U597 ( .A(n3210), .B(n3211), .Z(n391) );
  NANDN U598 ( .A(n3209), .B(n3208), .Z(n392) );
  NAND U599 ( .A(n391), .B(n392), .Z(n3250) );
  NAND U600 ( .A(n3327), .B(n3328), .Z(n393) );
  NANDN U601 ( .A(n3326), .B(n3325), .Z(n394) );
  NAND U602 ( .A(n393), .B(n394), .Z(n3367) );
  NAND U603 ( .A(n3444), .B(n3445), .Z(n395) );
  NANDN U604 ( .A(n3443), .B(n3442), .Z(n396) );
  NAND U605 ( .A(n395), .B(n396), .Z(n3484) );
  NAND U606 ( .A(n3561), .B(n3562), .Z(n397) );
  NANDN U607 ( .A(n3560), .B(n3559), .Z(n398) );
  NAND U608 ( .A(n397), .B(n398), .Z(n3601) );
  NAND U609 ( .A(n3678), .B(n3679), .Z(n399) );
  NANDN U610 ( .A(n3677), .B(n3676), .Z(n400) );
  NAND U611 ( .A(n399), .B(n400), .Z(n3718) );
  NAND U612 ( .A(n3795), .B(n3796), .Z(n401) );
  NANDN U613 ( .A(n3794), .B(n3793), .Z(n402) );
  NAND U614 ( .A(n401), .B(n402), .Z(n3835) );
  NAND U615 ( .A(n3912), .B(n3913), .Z(n403) );
  NANDN U616 ( .A(n3911), .B(n3910), .Z(n404) );
  NAND U617 ( .A(n403), .B(n404), .Z(n3952) );
  NAND U618 ( .A(n4029), .B(n4030), .Z(n405) );
  NANDN U619 ( .A(n4028), .B(n4027), .Z(n406) );
  NAND U620 ( .A(n405), .B(n406), .Z(n4069) );
  NAND U621 ( .A(n4146), .B(n4147), .Z(n407) );
  NANDN U622 ( .A(n4145), .B(n4144), .Z(n408) );
  NAND U623 ( .A(n407), .B(n408), .Z(n4186) );
  NAND U624 ( .A(n4263), .B(n4264), .Z(n409) );
  NANDN U625 ( .A(n4262), .B(n4261), .Z(n410) );
  NAND U626 ( .A(n409), .B(n410), .Z(n4303) );
  NAND U627 ( .A(n4380), .B(n4381), .Z(n411) );
  NANDN U628 ( .A(n4379), .B(n4378), .Z(n412) );
  NAND U629 ( .A(n411), .B(n412), .Z(n4420) );
  NAND U630 ( .A(n4497), .B(n4498), .Z(n413) );
  NANDN U631 ( .A(n4496), .B(n4495), .Z(n414) );
  NAND U632 ( .A(n413), .B(n414), .Z(n4537) );
  NAND U633 ( .A(n4614), .B(n4615), .Z(n415) );
  NANDN U634 ( .A(n4613), .B(n4612), .Z(n416) );
  NAND U635 ( .A(n415), .B(n416), .Z(n4654) );
  NAND U636 ( .A(n4731), .B(n4732), .Z(n417) );
  NANDN U637 ( .A(n4730), .B(n4729), .Z(n418) );
  NAND U638 ( .A(n417), .B(n418), .Z(n4771) );
  NAND U639 ( .A(n4848), .B(n4849), .Z(n419) );
  NANDN U640 ( .A(n4847), .B(n4846), .Z(n420) );
  NAND U641 ( .A(n419), .B(n420), .Z(n4888) );
  NAND U642 ( .A(n4965), .B(n4966), .Z(n421) );
  NANDN U643 ( .A(n4964), .B(n4963), .Z(n422) );
  NAND U644 ( .A(n421), .B(n422), .Z(n5005) );
  NAND U645 ( .A(n5082), .B(n5083), .Z(n423) );
  NANDN U646 ( .A(n5081), .B(n5080), .Z(n424) );
  NAND U647 ( .A(n423), .B(n424), .Z(n5122) );
  NAND U648 ( .A(n5199), .B(n5200), .Z(n425) );
  NANDN U649 ( .A(n5198), .B(n5197), .Z(n426) );
  NAND U650 ( .A(n425), .B(n426), .Z(n5239) );
  NAND U651 ( .A(n5316), .B(n5317), .Z(n427) );
  NANDN U652 ( .A(n5315), .B(n5314), .Z(n428) );
  NAND U653 ( .A(n427), .B(n428), .Z(n5356) );
  NAND U654 ( .A(n5433), .B(n5434), .Z(n429) );
  NANDN U655 ( .A(n5432), .B(n5431), .Z(n430) );
  NAND U656 ( .A(n429), .B(n430), .Z(n5473) );
  NAND U657 ( .A(n5550), .B(n5551), .Z(n431) );
  NANDN U658 ( .A(n5549), .B(n5548), .Z(n432) );
  NAND U659 ( .A(n431), .B(n432), .Z(n5590) );
  NAND U660 ( .A(n5667), .B(n5668), .Z(n433) );
  NANDN U661 ( .A(n5666), .B(n5665), .Z(n434) );
  NAND U662 ( .A(n433), .B(n434), .Z(n5707) );
  NAND U663 ( .A(n5784), .B(n5785), .Z(n435) );
  NANDN U664 ( .A(n5783), .B(n5782), .Z(n436) );
  NAND U665 ( .A(n435), .B(n436), .Z(n5824) );
  NAND U666 ( .A(n5901), .B(n5902), .Z(n437) );
  NANDN U667 ( .A(n5900), .B(n5899), .Z(n438) );
  NAND U668 ( .A(n437), .B(n438), .Z(n5941) );
  NAND U669 ( .A(n6018), .B(n6019), .Z(n439) );
  NANDN U670 ( .A(n6017), .B(n6016), .Z(n440) );
  NAND U671 ( .A(n439), .B(n440), .Z(n6058) );
  NAND U672 ( .A(n6135), .B(n6136), .Z(n441) );
  NANDN U673 ( .A(n6134), .B(n6133), .Z(n442) );
  NAND U674 ( .A(n441), .B(n442), .Z(n6175) );
  NAND U675 ( .A(n6252), .B(n6253), .Z(n443) );
  NANDN U676 ( .A(n6251), .B(n6250), .Z(n444) );
  NAND U677 ( .A(n443), .B(n444), .Z(n6292) );
  NAND U678 ( .A(n6369), .B(n6370), .Z(n445) );
  NANDN U679 ( .A(n6368), .B(n6367), .Z(n446) );
  NAND U680 ( .A(n445), .B(n446), .Z(n6409) );
  NAND U681 ( .A(n6486), .B(n6487), .Z(n447) );
  NANDN U682 ( .A(n6485), .B(n6484), .Z(n448) );
  NAND U683 ( .A(n447), .B(n448), .Z(n6526) );
  NAND U684 ( .A(n6603), .B(n6604), .Z(n449) );
  NANDN U685 ( .A(n6602), .B(n6601), .Z(n450) );
  NAND U686 ( .A(n449), .B(n450), .Z(n6643) );
  NAND U687 ( .A(n6720), .B(n6721), .Z(n451) );
  NANDN U688 ( .A(n6719), .B(n6718), .Z(n452) );
  NAND U689 ( .A(n451), .B(n452), .Z(n6760) );
  NAND U690 ( .A(n6837), .B(n6838), .Z(n453) );
  NANDN U691 ( .A(n6836), .B(n6835), .Z(n454) );
  NAND U692 ( .A(n453), .B(n454), .Z(n6877) );
  NAND U693 ( .A(n6954), .B(n6955), .Z(n455) );
  NANDN U694 ( .A(n6953), .B(n6952), .Z(n456) );
  NAND U695 ( .A(n455), .B(n456), .Z(n6994) );
  NAND U696 ( .A(n7071), .B(n7072), .Z(n457) );
  NANDN U697 ( .A(n7070), .B(n7069), .Z(n458) );
  NAND U698 ( .A(n457), .B(n458), .Z(n7111) );
  NAND U699 ( .A(n7188), .B(n7189), .Z(n459) );
  NANDN U700 ( .A(n7187), .B(n7186), .Z(n460) );
  NAND U701 ( .A(n459), .B(n460), .Z(n7228) );
  NAND U702 ( .A(n7305), .B(n7306), .Z(n461) );
  NANDN U703 ( .A(n7304), .B(n7303), .Z(n462) );
  NAND U704 ( .A(n461), .B(n462), .Z(n7345) );
  NAND U705 ( .A(n7422), .B(n7423), .Z(n463) );
  NANDN U706 ( .A(n7421), .B(n7420), .Z(n464) );
  NAND U707 ( .A(n463), .B(n464), .Z(n7462) );
  NAND U708 ( .A(n7539), .B(n7540), .Z(n465) );
  NANDN U709 ( .A(n7538), .B(n7537), .Z(n466) );
  NAND U710 ( .A(n465), .B(n466), .Z(n7579) );
  NAND U711 ( .A(n7656), .B(n7657), .Z(n467) );
  NANDN U712 ( .A(n7655), .B(n7654), .Z(n468) );
  NAND U713 ( .A(n467), .B(n468), .Z(n7696) );
  NAND U714 ( .A(n7773), .B(n7774), .Z(n469) );
  NANDN U715 ( .A(n7772), .B(n7771), .Z(n470) );
  NAND U716 ( .A(n469), .B(n470), .Z(n7813) );
  NAND U717 ( .A(n7890), .B(n7891), .Z(n471) );
  NANDN U718 ( .A(n7889), .B(n7888), .Z(n472) );
  NAND U719 ( .A(n471), .B(n472), .Z(n7930) );
  NAND U720 ( .A(n8007), .B(n8008), .Z(n473) );
  NANDN U721 ( .A(n8006), .B(n8005), .Z(n474) );
  NAND U722 ( .A(n473), .B(n474), .Z(n8047) );
  NAND U723 ( .A(n8124), .B(n8125), .Z(n475) );
  NANDN U724 ( .A(n8123), .B(n8122), .Z(n476) );
  NAND U725 ( .A(n475), .B(n476), .Z(n8164) );
  NAND U726 ( .A(n8241), .B(n8242), .Z(n477) );
  NANDN U727 ( .A(n8240), .B(n8239), .Z(n478) );
  NAND U728 ( .A(n477), .B(n478), .Z(n8281) );
  NAND U729 ( .A(n8358), .B(n8359), .Z(n479) );
  NANDN U730 ( .A(n8357), .B(n8356), .Z(n480) );
  NAND U731 ( .A(n479), .B(n480), .Z(n8398) );
  NAND U732 ( .A(n8475), .B(n8476), .Z(n481) );
  NANDN U733 ( .A(n8474), .B(n8473), .Z(n482) );
  NAND U734 ( .A(n481), .B(n482), .Z(n8515) );
  NAND U735 ( .A(n8592), .B(n8593), .Z(n483) );
  NANDN U736 ( .A(n8591), .B(n8590), .Z(n484) );
  NAND U737 ( .A(n483), .B(n484), .Z(n8632) );
  NAND U738 ( .A(n8710), .B(n8711), .Z(n485) );
  NANDN U739 ( .A(n8709), .B(n8708), .Z(n486) );
  NAND U740 ( .A(n485), .B(n486), .Z(n8748) );
  NAND U741 ( .A(n8825), .B(n8826), .Z(n487) );
  NANDN U742 ( .A(n8824), .B(n8823), .Z(n488) );
  NAND U743 ( .A(n487), .B(n488), .Z(n8865) );
  NAND U744 ( .A(n8942), .B(n8943), .Z(n489) );
  NANDN U745 ( .A(n8941), .B(n8940), .Z(n490) );
  NAND U746 ( .A(n489), .B(n490), .Z(n8982) );
  NAND U747 ( .A(n9059), .B(n9060), .Z(n491) );
  NANDN U748 ( .A(n9058), .B(n9057), .Z(n492) );
  NAND U749 ( .A(n491), .B(n492), .Z(n9099) );
  NAND U750 ( .A(n9176), .B(n9177), .Z(n493) );
  NANDN U751 ( .A(n9175), .B(n9174), .Z(n494) );
  NAND U752 ( .A(n493), .B(n494), .Z(n9216) );
  NAND U753 ( .A(n9293), .B(n9294), .Z(n495) );
  NANDN U754 ( .A(n9292), .B(n9291), .Z(n496) );
  NAND U755 ( .A(n495), .B(n496), .Z(n9333) );
  NAND U756 ( .A(n9410), .B(n9411), .Z(n497) );
  NANDN U757 ( .A(n9409), .B(n9408), .Z(n498) );
  NAND U758 ( .A(n497), .B(n498), .Z(n9450) );
  NAND U759 ( .A(n9527), .B(n9528), .Z(n499) );
  NANDN U760 ( .A(n9526), .B(n9525), .Z(n500) );
  NAND U761 ( .A(n499), .B(n500), .Z(n9567) );
  NAND U762 ( .A(n9644), .B(n9645), .Z(n501) );
  NANDN U763 ( .A(n9643), .B(n9642), .Z(n502) );
  NAND U764 ( .A(n501), .B(n502), .Z(n9684) );
  NAND U765 ( .A(n9761), .B(n9762), .Z(n503) );
  NANDN U766 ( .A(n9760), .B(n9759), .Z(n504) );
  NAND U767 ( .A(n503), .B(n504), .Z(n9801) );
  NAND U768 ( .A(n9878), .B(n9879), .Z(n505) );
  NANDN U769 ( .A(n9877), .B(n9876), .Z(n506) );
  NAND U770 ( .A(n505), .B(n506), .Z(n9918) );
  NAND U771 ( .A(n9995), .B(n9996), .Z(n507) );
  NANDN U772 ( .A(n9994), .B(n9993), .Z(n508) );
  NAND U773 ( .A(n507), .B(n508), .Z(n10035) );
  NAND U774 ( .A(n10112), .B(n10113), .Z(n509) );
  NANDN U775 ( .A(n10111), .B(n10110), .Z(n510) );
  NAND U776 ( .A(n509), .B(n510), .Z(n10152) );
  NAND U777 ( .A(n10229), .B(n10230), .Z(n511) );
  NANDN U778 ( .A(n10228), .B(n10227), .Z(n512) );
  NAND U779 ( .A(n511), .B(n512), .Z(n10269) );
  XOR U780 ( .A(n10499), .B(n10500), .Z(n10501) );
  XNOR U781 ( .A(n10542), .B(n10541), .Z(n10534) );
  ANDN U782 ( .B(n575), .A(n574), .Z(n583) );
  NAND U783 ( .A(n10348), .B(n10349), .Z(n513) );
  NANDN U784 ( .A(n10347), .B(n10346), .Z(n514) );
  NAND U785 ( .A(n513), .B(n514), .Z(n10389) );
  XNOR U786 ( .A(n10577), .B(n10576), .Z(n515) );
  XOR U787 ( .A(n10575), .B(n10574), .Z(n516) );
  AND U788 ( .A(n515), .B(n516), .Z(n517) );
  NANDN U789 ( .A(n10578), .B(n10579), .Z(n518) );
  XNOR U790 ( .A(n10578), .B(n10579), .Z(n519) );
  NAND U791 ( .A(n519), .B(n10580), .Z(n520) );
  AND U792 ( .A(n518), .B(n520), .Z(n521) );
  XNOR U793 ( .A(n517), .B(n521), .Z(n522) );
  XNOR U794 ( .A(a[255]), .B(n10581), .Z(n523) );
  NANDN U795 ( .A(n529), .B(n523), .Z(n524) );
  XNOR U796 ( .A(n522), .B(n524), .Z(n525) );
  NANDN U797 ( .A(n10583), .B(n10582), .Z(n526) );
  XNOR U798 ( .A(n525), .B(n526), .Z(c[511]) );
  IV U799 ( .A(b[0]), .Z(n527) );
  IV U800 ( .A(b[3]), .Z(n528) );
  IV U801 ( .A(b[7]), .Z(n529) );
  NANDN U802 ( .A(n527), .B(a[0]), .Z(n531) );
  XNOR U803 ( .A(n531), .B(sreg[248]), .Z(c[248]) );
  IV U804 ( .A(b[1]), .Z(n10434) );
  ANDN U805 ( .B(a[0]), .A(n10434), .Z(n530) );
  NANDN U806 ( .A(n527), .B(a[1]), .Z(n536) );
  XNOR U807 ( .A(n530), .B(n536), .Z(n539) );
  XNOR U808 ( .A(sreg[249]), .B(n539), .Z(n541) );
  NANDN U809 ( .A(n531), .B(sreg[248]), .Z(n540) );
  XOR U810 ( .A(n541), .B(n540), .Z(c[249]) );
  NANDN U811 ( .A(n527), .B(a[2]), .Z(n532) );
  XOR U812 ( .A(n10434), .B(n532), .Z(n534) );
  NANDN U813 ( .A(b[0]), .B(a[1]), .Z(n533) );
  NAND U814 ( .A(n534), .B(n533), .Z(n544) );
  IV U815 ( .A(a[0]), .Z(n709) );
  NANDN U816 ( .A(n709), .B(b[2]), .Z(n535) );
  XOR U817 ( .A(n10434), .B(n535), .Z(n538) );
  OR U818 ( .A(n536), .B(a[0]), .Z(n537) );
  AND U819 ( .A(n538), .B(n537), .Z(n545) );
  XOR U820 ( .A(n544), .B(n545), .Z(n562) );
  NAND U821 ( .A(sreg[249]), .B(n539), .Z(n543) );
  OR U822 ( .A(n541), .B(n540), .Z(n542) );
  NAND U823 ( .A(n543), .B(n542), .Z(n560) );
  XNOR U824 ( .A(n560), .B(sreg[250]), .Z(n561) );
  XOR U825 ( .A(n562), .B(n561), .Z(c[250]) );
  ANDN U826 ( .B(n545), .A(n544), .Z(n573) );
  XNOR U827 ( .A(n528), .B(a[0]), .Z(n548) );
  XNOR U828 ( .A(n528), .B(b[1]), .Z(n547) );
  XNOR U829 ( .A(n528), .B(b[2]), .Z(n546) );
  AND U830 ( .A(n547), .B(n546), .Z(n10399) );
  NAND U831 ( .A(n548), .B(n10399), .Z(n550) );
  XNOR U832 ( .A(n528), .B(a[1]), .Z(n568) );
  XNOR U833 ( .A(n10434), .B(b[2]), .Z(n10398) );
  NAND U834 ( .A(n568), .B(n10398), .Z(n549) );
  AND U835 ( .A(n550), .B(n549), .Z(n574) );
  NANDN U836 ( .A(n527), .B(a[3]), .Z(n551) );
  XOR U837 ( .A(n10434), .B(n551), .Z(n553) );
  NANDN U838 ( .A(b[0]), .B(a[2]), .Z(n552) );
  AND U839 ( .A(n553), .B(n552), .Z(n575) );
  XNOR U840 ( .A(n574), .B(n575), .Z(n572) );
  OR U841 ( .A(b[2]), .B(n10434), .Z(n555) );
  NANDN U842 ( .A(n528), .B(b[2]), .Z(n554) );
  AND U843 ( .A(n555), .B(n554), .Z(n557) );
  NANDN U844 ( .A(a[0]), .B(n10398), .Z(n556) );
  NANDN U845 ( .A(n557), .B(n556), .Z(n558) );
  AND U846 ( .A(n558), .B(b[3]), .Z(n571) );
  XOR U847 ( .A(n572), .B(n571), .Z(n559) );
  XOR U848 ( .A(n573), .B(n559), .Z(n577) );
  XNOR U849 ( .A(sreg[251]), .B(n577), .Z(n579) );
  NAND U850 ( .A(n560), .B(sreg[250]), .Z(n564) );
  OR U851 ( .A(n562), .B(n561), .Z(n563) );
  AND U852 ( .A(n564), .B(n563), .Z(n578) );
  XOR U853 ( .A(n579), .B(n578), .Z(c[251]) );
  NANDN U854 ( .A(n527), .B(a[4]), .Z(n565) );
  XOR U855 ( .A(n10434), .B(n565), .Z(n567) );
  NANDN U856 ( .A(b[0]), .B(a[3]), .Z(n566) );
  AND U857 ( .A(n567), .B(n566), .Z(n598) );
  XNOR U858 ( .A(n528), .B(a[2]), .Z(n595) );
  NAND U859 ( .A(n595), .B(n10398), .Z(n570) );
  NAND U860 ( .A(n568), .B(n10399), .Z(n569) );
  AND U861 ( .A(n570), .B(n569), .Z(n599) );
  XOR U862 ( .A(n598), .B(n599), .Z(n601) );
  IV U863 ( .A(b[4]), .Z(n10521) );
  XOR U864 ( .A(n528), .B(n10521), .Z(n10481) );
  NANDN U865 ( .A(n709), .B(n10481), .Z(n600) );
  XNOR U866 ( .A(n601), .B(n600), .Z(n582) );
  XNOR U867 ( .A(n584), .B(n583), .Z(n576) );
  XNOR U868 ( .A(n582), .B(n576), .Z(n605) );
  NAND U869 ( .A(n577), .B(sreg[251]), .Z(n581) );
  OR U870 ( .A(n579), .B(n578), .Z(n580) );
  NAND U871 ( .A(n581), .B(n580), .Z(n604) );
  XNOR U872 ( .A(n604), .B(sreg[252]), .Z(n606) );
  XNOR U873 ( .A(n605), .B(n606), .Z(c[252]) );
  NANDN U874 ( .A(n527), .B(a[5]), .Z(n585) );
  XOR U875 ( .A(n10434), .B(n585), .Z(n587) );
  NANDN U876 ( .A(b[0]), .B(a[4]), .Z(n586) );
  AND U877 ( .A(n587), .B(n586), .Z(n615) );
  XOR U878 ( .A(b[5]), .B(a[1]), .Z(n623) );
  AND U879 ( .A(n10481), .B(n623), .Z(n592) );
  XNOR U880 ( .A(b[5]), .B(n709), .Z(n590) );
  XNOR U881 ( .A(b[5]), .B(n528), .Z(n589) );
  XNOR U882 ( .A(b[5]), .B(n10521), .Z(n588) );
  AND U883 ( .A(n589), .B(n588), .Z(n10482) );
  NAND U884 ( .A(n590), .B(n10482), .Z(n591) );
  NANDN U885 ( .A(n592), .B(n591), .Z(n616) );
  XNOR U886 ( .A(n615), .B(n616), .Z(n629) );
  NANDN U887 ( .A(n528), .B(b[4]), .Z(n10520) );
  AND U888 ( .A(n10520), .B(b[5]), .Z(n10552) );
  XNOR U889 ( .A(n10521), .B(b[3]), .Z(n593) );
  NANDN U890 ( .A(n709), .B(n593), .Z(n594) );
  NAND U891 ( .A(n10552), .B(n594), .Z(n626) );
  XNOR U892 ( .A(b[3]), .B(a[3]), .Z(n617) );
  NANDN U893 ( .A(n617), .B(n10398), .Z(n597) );
  NAND U894 ( .A(n10399), .B(n595), .Z(n596) );
  NAND U895 ( .A(n597), .B(n596), .Z(n627) );
  XNOR U896 ( .A(n626), .B(n627), .Z(n628) );
  XOR U897 ( .A(n629), .B(n628), .Z(n610) );
  NANDN U898 ( .A(n599), .B(n598), .Z(n603) );
  OR U899 ( .A(n601), .B(n600), .Z(n602) );
  AND U900 ( .A(n603), .B(n602), .Z(n609) );
  XOR U901 ( .A(n610), .B(n609), .Z(n611) );
  XNOR U902 ( .A(n612), .B(n611), .Z(n632) );
  XNOR U903 ( .A(sreg[253]), .B(n632), .Z(n634) );
  NAND U904 ( .A(n604), .B(sreg[252]), .Z(n608) );
  NANDN U905 ( .A(n606), .B(n605), .Z(n607) );
  AND U906 ( .A(n608), .B(n607), .Z(n633) );
  XOR U907 ( .A(n634), .B(n633), .Z(c[253]) );
  OR U908 ( .A(n610), .B(n609), .Z(n614) );
  NANDN U909 ( .A(n612), .B(n611), .Z(n613) );
  NAND U910 ( .A(n614), .B(n613), .Z(n640) );
  AND U911 ( .A(n616), .B(n615), .Z(n667) );
  XNOR U912 ( .A(n528), .B(a[4]), .Z(n661) );
  NAND U913 ( .A(n661), .B(n10398), .Z(n619) );
  NANDN U914 ( .A(n617), .B(n10399), .Z(n618) );
  NAND U915 ( .A(n619), .B(n618), .Z(n646) );
  NANDN U916 ( .A(n527), .B(a[6]), .Z(n620) );
  XOR U917 ( .A(n10434), .B(n620), .Z(n622) );
  NANDN U918 ( .A(b[0]), .B(a[5]), .Z(n621) );
  AND U919 ( .A(n622), .B(n621), .Z(n643) );
  XOR U920 ( .A(b[5]), .B(b[6]), .Z(n10545) );
  NANDN U921 ( .A(n709), .B(n10545), .Z(n644) );
  XNOR U922 ( .A(n643), .B(n644), .Z(n645) );
  XNOR U923 ( .A(n646), .B(n645), .Z(n664) );
  XOR U924 ( .A(b[5]), .B(a[2]), .Z(n647) );
  NAND U925 ( .A(n10481), .B(n647), .Z(n625) );
  NAND U926 ( .A(n10482), .B(n623), .Z(n624) );
  NAND U927 ( .A(n625), .B(n624), .Z(n665) );
  XNOR U928 ( .A(n664), .B(n665), .Z(n666) );
  XOR U929 ( .A(n667), .B(n666), .Z(n637) );
  NANDN U930 ( .A(n627), .B(n626), .Z(n631) );
  NAND U931 ( .A(n629), .B(n628), .Z(n630) );
  NAND U932 ( .A(n631), .B(n630), .Z(n638) );
  XNOR U933 ( .A(n637), .B(n638), .Z(n639) );
  XNOR U934 ( .A(n640), .B(n639), .Z(n672) );
  NAND U935 ( .A(sreg[253]), .B(n632), .Z(n636) );
  OR U936 ( .A(n634), .B(n633), .Z(n635) );
  NAND U937 ( .A(n636), .B(n635), .Z(n670) );
  XNOR U938 ( .A(n670), .B(sreg[254]), .Z(n671) );
  XOR U939 ( .A(n672), .B(n671), .Z(c[254]) );
  NANDN U940 ( .A(n638), .B(n637), .Z(n642) );
  NAND U941 ( .A(n640), .B(n639), .Z(n641) );
  NAND U942 ( .A(n642), .B(n641), .Z(n683) );
  XOR U943 ( .A(b[5]), .B(a[3]), .Z(n710) );
  NAND U944 ( .A(n710), .B(n10481), .Z(n649) );
  NAND U945 ( .A(n647), .B(n10482), .Z(n648) );
  NAND U946 ( .A(n649), .B(n648), .Z(n699) );
  XNOR U947 ( .A(n529), .B(a[1]), .Z(n703) );
  AND U948 ( .A(n10545), .B(n703), .Z(n653) );
  XNOR U949 ( .A(n529), .B(a[0]), .Z(n651) );
  XOR U950 ( .A(b[7]), .B(b[5]), .Z(n650) );
  XNOR U951 ( .A(b[5]), .B(b[6]), .Z(n10557) );
  AND U952 ( .A(n650), .B(n10557), .Z(n10546) );
  NAND U953 ( .A(n651), .B(n10546), .Z(n652) );
  NANDN U954 ( .A(n653), .B(n652), .Z(n698) );
  XNOR U955 ( .A(n699), .B(n698), .Z(n695) );
  OR U956 ( .A(b[5]), .B(a[0]), .Z(n654) );
  NAND U957 ( .A(b[6]), .B(n654), .Z(n656) );
  ANDN U958 ( .B(b[5]), .A(n709), .Z(n655) );
  ANDN U959 ( .B(n656), .A(n655), .Z(n657) );
  AND U960 ( .A(n657), .B(b[7]), .Z(n692) );
  NANDN U961 ( .A(n527), .B(a[7]), .Z(n658) );
  XOR U962 ( .A(n10434), .B(n658), .Z(n660) );
  NANDN U963 ( .A(b[0]), .B(a[6]), .Z(n659) );
  AND U964 ( .A(n660), .B(n659), .Z(n693) );
  XOR U965 ( .A(n692), .B(n693), .Z(n694) );
  XOR U966 ( .A(n695), .B(n694), .Z(n686) );
  XOR U967 ( .A(n528), .B(a[5]), .Z(n700) );
  NANDN U968 ( .A(n700), .B(n10398), .Z(n663) );
  NAND U969 ( .A(n10399), .B(n661), .Z(n662) );
  AND U970 ( .A(n663), .B(n662), .Z(n687) );
  XNOR U971 ( .A(n686), .B(n687), .Z(n688) );
  XNOR U972 ( .A(n689), .B(n688), .Z(n680) );
  NANDN U973 ( .A(n665), .B(n664), .Z(n669) );
  NANDN U974 ( .A(n667), .B(n666), .Z(n668) );
  NAND U975 ( .A(n669), .B(n668), .Z(n681) );
  XNOR U976 ( .A(n680), .B(n681), .Z(n682) );
  XOR U977 ( .A(n683), .B(n682), .Z(n675) );
  XNOR U978 ( .A(sreg[255]), .B(n675), .Z(n677) );
  NAND U979 ( .A(n670), .B(sreg[254]), .Z(n674) );
  OR U980 ( .A(n672), .B(n671), .Z(n673) );
  AND U981 ( .A(n674), .B(n673), .Z(n676) );
  XOR U982 ( .A(n677), .B(n676), .Z(c[255]) );
  NAND U983 ( .A(sreg[255]), .B(n675), .Z(n679) );
  OR U984 ( .A(n677), .B(n676), .Z(n678) );
  NAND U985 ( .A(n679), .B(n678), .Z(n749) );
  XNOR U986 ( .A(n749), .B(sreg[256]), .Z(n751) );
  NANDN U987 ( .A(n681), .B(n680), .Z(n685) );
  NAND U988 ( .A(n683), .B(n682), .Z(n684) );
  NAND U989 ( .A(n685), .B(n684), .Z(n746) );
  NAND U990 ( .A(n687), .B(n686), .Z(n691) );
  OR U991 ( .A(n689), .B(n688), .Z(n690) );
  NAND U992 ( .A(n691), .B(n690), .Z(n744) );
  OR U993 ( .A(n693), .B(n692), .Z(n697) );
  NAND U994 ( .A(n695), .B(n694), .Z(n696) );
  NAND U995 ( .A(n697), .B(n696), .Z(n737) );
  NAND U996 ( .A(n699), .B(n698), .Z(n734) );
  XNOR U997 ( .A(b[3]), .B(a[6]), .Z(n716) );
  NANDN U998 ( .A(n716), .B(n10398), .Z(n702) );
  NANDN U999 ( .A(n700), .B(n10399), .Z(n701) );
  NAND U1000 ( .A(n702), .B(n701), .Z(n732) );
  XNOR U1001 ( .A(b[7]), .B(a[2]), .Z(n713) );
  NANDN U1002 ( .A(n713), .B(n10545), .Z(n705) );
  NAND U1003 ( .A(n10546), .B(n703), .Z(n704) );
  AND U1004 ( .A(n705), .B(n704), .Z(n731) );
  XNOR U1005 ( .A(n732), .B(n731), .Z(n733) );
  XNOR U1006 ( .A(n734), .B(n733), .Z(n738) );
  XNOR U1007 ( .A(n737), .B(n738), .Z(n739) );
  NANDN U1008 ( .A(n527), .B(a[8]), .Z(n706) );
  XOR U1009 ( .A(n10434), .B(n706), .Z(n708) );
  NANDN U1010 ( .A(b[0]), .B(a[7]), .Z(n707) );
  AND U1011 ( .A(n708), .B(n707), .Z(n728) );
  ANDN U1012 ( .B(b[7]), .A(n709), .Z(n725) );
  XOR U1013 ( .A(b[5]), .B(a[4]), .Z(n722) );
  NAND U1014 ( .A(n10481), .B(n722), .Z(n712) );
  NAND U1015 ( .A(n10482), .B(n710), .Z(n711) );
  NAND U1016 ( .A(n712), .B(n711), .Z(n726) );
  XOR U1017 ( .A(n725), .B(n726), .Z(n727) );
  XOR U1018 ( .A(n728), .B(n727), .Z(n740) );
  XNOR U1019 ( .A(n739), .B(n740), .Z(n743) );
  XNOR U1020 ( .A(n744), .B(n743), .Z(n745) );
  XOR U1021 ( .A(n746), .B(n745), .Z(n750) );
  XOR U1022 ( .A(n751), .B(n750), .Z(c[256]) );
  XNOR U1023 ( .A(b[7]), .B(a[3]), .Z(n772) );
  NANDN U1024 ( .A(n772), .B(n10545), .Z(n715) );
  NANDN U1025 ( .A(n713), .B(n10546), .Z(n714) );
  NAND U1026 ( .A(n715), .B(n714), .Z(n760) );
  XNOR U1027 ( .A(b[3]), .B(a[7]), .Z(n775) );
  NANDN U1028 ( .A(n775), .B(n10398), .Z(n718) );
  NANDN U1029 ( .A(n716), .B(n10399), .Z(n717) );
  AND U1030 ( .A(n718), .B(n717), .Z(n761) );
  XNOR U1031 ( .A(n760), .B(n761), .Z(n762) );
  NANDN U1032 ( .A(n527), .B(a[9]), .Z(n719) );
  XOR U1033 ( .A(n10434), .B(n719), .Z(n721) );
  NANDN U1034 ( .A(b[0]), .B(a[8]), .Z(n720) );
  AND U1035 ( .A(n721), .B(n720), .Z(n768) );
  XOR U1036 ( .A(b[5]), .B(a[5]), .Z(n781) );
  NAND U1037 ( .A(n781), .B(n10481), .Z(n724) );
  NAND U1038 ( .A(n722), .B(n10482), .Z(n723) );
  NAND U1039 ( .A(n724), .B(n723), .Z(n766) );
  NANDN U1040 ( .A(n529), .B(a[1]), .Z(n767) );
  XNOR U1041 ( .A(n766), .B(n767), .Z(n769) );
  XOR U1042 ( .A(n768), .B(n769), .Z(n763) );
  XOR U1043 ( .A(n762), .B(n763), .Z(n784) );
  OR U1044 ( .A(n726), .B(n725), .Z(n730) );
  NANDN U1045 ( .A(n728), .B(n727), .Z(n729) );
  AND U1046 ( .A(n730), .B(n729), .Z(n785) );
  XNOR U1047 ( .A(n784), .B(n785), .Z(n787) );
  NANDN U1048 ( .A(n732), .B(n731), .Z(n736) );
  NAND U1049 ( .A(n734), .B(n733), .Z(n735) );
  AND U1050 ( .A(n736), .B(n735), .Z(n786) );
  XNOR U1051 ( .A(n787), .B(n786), .Z(n754) );
  NANDN U1052 ( .A(n738), .B(n737), .Z(n742) );
  NANDN U1053 ( .A(n740), .B(n739), .Z(n741) );
  AND U1054 ( .A(n742), .B(n741), .Z(n755) );
  XNOR U1055 ( .A(n754), .B(n755), .Z(n757) );
  NAND U1056 ( .A(n744), .B(n743), .Z(n748) );
  OR U1057 ( .A(n746), .B(n745), .Z(n747) );
  AND U1058 ( .A(n748), .B(n747), .Z(n756) );
  XNOR U1059 ( .A(n757), .B(n756), .Z(n790) );
  XNOR U1060 ( .A(sreg[257]), .B(n790), .Z(n792) );
  NAND U1061 ( .A(n749), .B(sreg[256]), .Z(n753) );
  OR U1062 ( .A(n751), .B(n750), .Z(n752) );
  AND U1063 ( .A(n753), .B(n752), .Z(n791) );
  XOR U1064 ( .A(n792), .B(n791), .Z(c[257]) );
  NAND U1065 ( .A(n755), .B(n754), .Z(n759) );
  NANDN U1066 ( .A(n757), .B(n756), .Z(n758) );
  NAND U1067 ( .A(n759), .B(n758), .Z(n797) );
  NANDN U1068 ( .A(n761), .B(n760), .Z(n765) );
  NAND U1069 ( .A(n763), .B(n762), .Z(n764) );
  NAND U1070 ( .A(n765), .B(n764), .Z(n828) );
  NANDN U1071 ( .A(n767), .B(n766), .Z(n771) );
  NAND U1072 ( .A(n769), .B(n768), .Z(n770) );
  NAND U1073 ( .A(n771), .B(n770), .Z(n826) );
  XNOR U1074 ( .A(b[7]), .B(a[4]), .Z(n813) );
  NANDN U1075 ( .A(n813), .B(n10545), .Z(n774) );
  NANDN U1076 ( .A(n772), .B(n10546), .Z(n773) );
  NAND U1077 ( .A(n774), .B(n773), .Z(n801) );
  XNOR U1078 ( .A(b[3]), .B(a[8]), .Z(n816) );
  NANDN U1079 ( .A(n816), .B(n10398), .Z(n777) );
  NANDN U1080 ( .A(n775), .B(n10399), .Z(n776) );
  AND U1081 ( .A(n777), .B(n776), .Z(n802) );
  XNOR U1082 ( .A(n801), .B(n802), .Z(n803) );
  NANDN U1083 ( .A(n527), .B(a[10]), .Z(n778) );
  XOR U1084 ( .A(n10434), .B(n778), .Z(n780) );
  NANDN U1085 ( .A(b[0]), .B(a[9]), .Z(n779) );
  AND U1086 ( .A(n780), .B(n779), .Z(n809) );
  XOR U1087 ( .A(b[5]), .B(a[6]), .Z(n822) );
  NAND U1088 ( .A(n822), .B(n10481), .Z(n783) );
  NAND U1089 ( .A(n781), .B(n10482), .Z(n782) );
  NAND U1090 ( .A(n783), .B(n782), .Z(n807) );
  NANDN U1091 ( .A(n529), .B(a[2]), .Z(n808) );
  XNOR U1092 ( .A(n807), .B(n808), .Z(n810) );
  XOR U1093 ( .A(n809), .B(n810), .Z(n804) );
  XOR U1094 ( .A(n803), .B(n804), .Z(n825) );
  XOR U1095 ( .A(n826), .B(n825), .Z(n827) );
  XNOR U1096 ( .A(n828), .B(n827), .Z(n795) );
  NAND U1097 ( .A(n785), .B(n784), .Z(n789) );
  NANDN U1098 ( .A(n787), .B(n786), .Z(n788) );
  NAND U1099 ( .A(n789), .B(n788), .Z(n796) );
  XOR U1100 ( .A(n795), .B(n796), .Z(n798) );
  XNOR U1101 ( .A(n797), .B(n798), .Z(n831) );
  XNOR U1102 ( .A(n831), .B(sreg[258]), .Z(n833) );
  NAND U1103 ( .A(sreg[257]), .B(n790), .Z(n794) );
  OR U1104 ( .A(n792), .B(n791), .Z(n793) );
  AND U1105 ( .A(n794), .B(n793), .Z(n832) );
  XOR U1106 ( .A(n833), .B(n832), .Z(c[258]) );
  NANDN U1107 ( .A(n796), .B(n795), .Z(n800) );
  OR U1108 ( .A(n798), .B(n797), .Z(n799) );
  NAND U1109 ( .A(n800), .B(n799), .Z(n839) );
  NANDN U1110 ( .A(n802), .B(n801), .Z(n806) );
  NAND U1111 ( .A(n804), .B(n803), .Z(n805) );
  NAND U1112 ( .A(n806), .B(n805), .Z(n867) );
  NANDN U1113 ( .A(n808), .B(n807), .Z(n812) );
  NAND U1114 ( .A(n810), .B(n809), .Z(n811) );
  NAND U1115 ( .A(n812), .B(n811), .Z(n865) );
  XNOR U1116 ( .A(b[7]), .B(a[5]), .Z(n852) );
  NANDN U1117 ( .A(n852), .B(n10545), .Z(n815) );
  NANDN U1118 ( .A(n813), .B(n10546), .Z(n814) );
  NAND U1119 ( .A(n815), .B(n814), .Z(n840) );
  XNOR U1120 ( .A(b[3]), .B(a[9]), .Z(n855) );
  NANDN U1121 ( .A(n855), .B(n10398), .Z(n818) );
  NANDN U1122 ( .A(n816), .B(n10399), .Z(n817) );
  AND U1123 ( .A(n818), .B(n817), .Z(n841) );
  XNOR U1124 ( .A(n840), .B(n841), .Z(n842) );
  NANDN U1125 ( .A(n527), .B(a[11]), .Z(n819) );
  XOR U1126 ( .A(n10434), .B(n819), .Z(n821) );
  NANDN U1127 ( .A(b[0]), .B(a[10]), .Z(n820) );
  AND U1128 ( .A(n821), .B(n820), .Z(n848) );
  XOR U1129 ( .A(b[5]), .B(a[7]), .Z(n861) );
  NAND U1130 ( .A(n861), .B(n10481), .Z(n824) );
  NAND U1131 ( .A(n822), .B(n10482), .Z(n823) );
  NAND U1132 ( .A(n824), .B(n823), .Z(n846) );
  NANDN U1133 ( .A(n529), .B(a[3]), .Z(n847) );
  XNOR U1134 ( .A(n846), .B(n847), .Z(n849) );
  XOR U1135 ( .A(n848), .B(n849), .Z(n843) );
  XOR U1136 ( .A(n842), .B(n843), .Z(n864) );
  XOR U1137 ( .A(n865), .B(n864), .Z(n866) );
  XNOR U1138 ( .A(n867), .B(n866), .Z(n836) );
  NAND U1139 ( .A(n826), .B(n825), .Z(n830) );
  NAND U1140 ( .A(n828), .B(n827), .Z(n829) );
  NAND U1141 ( .A(n830), .B(n829), .Z(n837) );
  XNOR U1142 ( .A(n836), .B(n837), .Z(n838) );
  XNOR U1143 ( .A(n839), .B(n838), .Z(n870) );
  XNOR U1144 ( .A(n870), .B(sreg[259]), .Z(n872) );
  NAND U1145 ( .A(n831), .B(sreg[258]), .Z(n835) );
  OR U1146 ( .A(n833), .B(n832), .Z(n834) );
  AND U1147 ( .A(n835), .B(n834), .Z(n871) );
  XOR U1148 ( .A(n872), .B(n871), .Z(c[259]) );
  NANDN U1149 ( .A(n841), .B(n840), .Z(n845) );
  NAND U1150 ( .A(n843), .B(n842), .Z(n844) );
  NAND U1151 ( .A(n845), .B(n844), .Z(n906) );
  NANDN U1152 ( .A(n847), .B(n846), .Z(n851) );
  NAND U1153 ( .A(n849), .B(n848), .Z(n850) );
  NAND U1154 ( .A(n851), .B(n850), .Z(n904) );
  XNOR U1155 ( .A(b[7]), .B(a[6]), .Z(n891) );
  NANDN U1156 ( .A(n891), .B(n10545), .Z(n854) );
  NANDN U1157 ( .A(n852), .B(n10546), .Z(n853) );
  NAND U1158 ( .A(n854), .B(n853), .Z(n879) );
  XNOR U1159 ( .A(b[3]), .B(a[10]), .Z(n894) );
  NANDN U1160 ( .A(n894), .B(n10398), .Z(n857) );
  NANDN U1161 ( .A(n855), .B(n10399), .Z(n856) );
  AND U1162 ( .A(n857), .B(n856), .Z(n880) );
  XNOR U1163 ( .A(n879), .B(n880), .Z(n881) );
  NANDN U1164 ( .A(n527), .B(a[12]), .Z(n858) );
  XOR U1165 ( .A(n10434), .B(n858), .Z(n860) );
  NANDN U1166 ( .A(b[0]), .B(a[11]), .Z(n859) );
  AND U1167 ( .A(n860), .B(n859), .Z(n887) );
  XOR U1168 ( .A(b[5]), .B(a[8]), .Z(n900) );
  NAND U1169 ( .A(n900), .B(n10481), .Z(n863) );
  NAND U1170 ( .A(n861), .B(n10482), .Z(n862) );
  NAND U1171 ( .A(n863), .B(n862), .Z(n885) );
  NANDN U1172 ( .A(n529), .B(a[4]), .Z(n886) );
  XNOR U1173 ( .A(n885), .B(n886), .Z(n888) );
  XOR U1174 ( .A(n887), .B(n888), .Z(n882) );
  XOR U1175 ( .A(n881), .B(n882), .Z(n903) );
  XOR U1176 ( .A(n904), .B(n903), .Z(n905) );
  XNOR U1177 ( .A(n906), .B(n905), .Z(n875) );
  NAND U1178 ( .A(n865), .B(n864), .Z(n869) );
  NAND U1179 ( .A(n867), .B(n866), .Z(n868) );
  NAND U1180 ( .A(n869), .B(n868), .Z(n876) );
  XNOR U1181 ( .A(n875), .B(n876), .Z(n877) );
  XNOR U1182 ( .A(n878), .B(n877), .Z(n909) );
  XNOR U1183 ( .A(n909), .B(sreg[260]), .Z(n911) );
  NAND U1184 ( .A(n870), .B(sreg[259]), .Z(n874) );
  OR U1185 ( .A(n872), .B(n871), .Z(n873) );
  AND U1186 ( .A(n874), .B(n873), .Z(n910) );
  XOR U1187 ( .A(n911), .B(n910), .Z(c[260]) );
  NANDN U1188 ( .A(n880), .B(n879), .Z(n884) );
  NAND U1189 ( .A(n882), .B(n881), .Z(n883) );
  NAND U1190 ( .A(n884), .B(n883), .Z(n945) );
  NANDN U1191 ( .A(n886), .B(n885), .Z(n890) );
  NAND U1192 ( .A(n888), .B(n887), .Z(n889) );
  NAND U1193 ( .A(n890), .B(n889), .Z(n943) );
  XNOR U1194 ( .A(b[7]), .B(a[7]), .Z(n930) );
  NANDN U1195 ( .A(n930), .B(n10545), .Z(n893) );
  NANDN U1196 ( .A(n891), .B(n10546), .Z(n892) );
  NAND U1197 ( .A(n893), .B(n892), .Z(n918) );
  XNOR U1198 ( .A(b[3]), .B(a[11]), .Z(n933) );
  NANDN U1199 ( .A(n933), .B(n10398), .Z(n896) );
  NANDN U1200 ( .A(n894), .B(n10399), .Z(n895) );
  AND U1201 ( .A(n896), .B(n895), .Z(n919) );
  XNOR U1202 ( .A(n918), .B(n919), .Z(n920) );
  NANDN U1203 ( .A(n527), .B(a[13]), .Z(n897) );
  XOR U1204 ( .A(n10434), .B(n897), .Z(n899) );
  NANDN U1205 ( .A(b[0]), .B(a[12]), .Z(n898) );
  AND U1206 ( .A(n899), .B(n898), .Z(n926) );
  XOR U1207 ( .A(b[5]), .B(a[9]), .Z(n939) );
  NAND U1208 ( .A(n939), .B(n10481), .Z(n902) );
  NAND U1209 ( .A(n900), .B(n10482), .Z(n901) );
  NAND U1210 ( .A(n902), .B(n901), .Z(n924) );
  NANDN U1211 ( .A(n529), .B(a[5]), .Z(n925) );
  XNOR U1212 ( .A(n924), .B(n925), .Z(n927) );
  XOR U1213 ( .A(n926), .B(n927), .Z(n921) );
  XOR U1214 ( .A(n920), .B(n921), .Z(n942) );
  XOR U1215 ( .A(n943), .B(n942), .Z(n944) );
  XNOR U1216 ( .A(n945), .B(n944), .Z(n914) );
  NAND U1217 ( .A(n904), .B(n903), .Z(n908) );
  NAND U1218 ( .A(n906), .B(n905), .Z(n907) );
  NAND U1219 ( .A(n908), .B(n907), .Z(n915) );
  XNOR U1220 ( .A(n914), .B(n915), .Z(n916) );
  XNOR U1221 ( .A(n917), .B(n916), .Z(n948) );
  XNOR U1222 ( .A(n948), .B(sreg[261]), .Z(n950) );
  NAND U1223 ( .A(n909), .B(sreg[260]), .Z(n913) );
  OR U1224 ( .A(n911), .B(n910), .Z(n912) );
  AND U1225 ( .A(n913), .B(n912), .Z(n949) );
  XOR U1226 ( .A(n950), .B(n949), .Z(c[261]) );
  NANDN U1227 ( .A(n919), .B(n918), .Z(n923) );
  NAND U1228 ( .A(n921), .B(n920), .Z(n922) );
  NAND U1229 ( .A(n923), .B(n922), .Z(n984) );
  NANDN U1230 ( .A(n925), .B(n924), .Z(n929) );
  NAND U1231 ( .A(n927), .B(n926), .Z(n928) );
  NAND U1232 ( .A(n929), .B(n928), .Z(n982) );
  XNOR U1233 ( .A(b[7]), .B(a[8]), .Z(n969) );
  NANDN U1234 ( .A(n969), .B(n10545), .Z(n932) );
  NANDN U1235 ( .A(n930), .B(n10546), .Z(n931) );
  NAND U1236 ( .A(n932), .B(n931), .Z(n957) );
  XNOR U1237 ( .A(b[3]), .B(a[12]), .Z(n972) );
  NANDN U1238 ( .A(n972), .B(n10398), .Z(n935) );
  NANDN U1239 ( .A(n933), .B(n10399), .Z(n934) );
  AND U1240 ( .A(n935), .B(n934), .Z(n958) );
  XNOR U1241 ( .A(n957), .B(n958), .Z(n959) );
  NANDN U1242 ( .A(n527), .B(a[14]), .Z(n936) );
  XOR U1243 ( .A(n10434), .B(n936), .Z(n938) );
  NANDN U1244 ( .A(b[0]), .B(a[13]), .Z(n937) );
  AND U1245 ( .A(n938), .B(n937), .Z(n965) );
  XOR U1246 ( .A(b[5]), .B(a[10]), .Z(n978) );
  NAND U1247 ( .A(n978), .B(n10481), .Z(n941) );
  NAND U1248 ( .A(n939), .B(n10482), .Z(n940) );
  NAND U1249 ( .A(n941), .B(n940), .Z(n963) );
  NANDN U1250 ( .A(n529), .B(a[6]), .Z(n964) );
  XNOR U1251 ( .A(n963), .B(n964), .Z(n966) );
  XOR U1252 ( .A(n965), .B(n966), .Z(n960) );
  XOR U1253 ( .A(n959), .B(n960), .Z(n981) );
  XOR U1254 ( .A(n982), .B(n981), .Z(n983) );
  XNOR U1255 ( .A(n984), .B(n983), .Z(n953) );
  NAND U1256 ( .A(n943), .B(n942), .Z(n947) );
  NAND U1257 ( .A(n945), .B(n944), .Z(n946) );
  NAND U1258 ( .A(n947), .B(n946), .Z(n954) );
  XNOR U1259 ( .A(n953), .B(n954), .Z(n955) );
  XNOR U1260 ( .A(n956), .B(n955), .Z(n987) );
  XNOR U1261 ( .A(n987), .B(sreg[262]), .Z(n989) );
  NAND U1262 ( .A(n948), .B(sreg[261]), .Z(n952) );
  OR U1263 ( .A(n950), .B(n949), .Z(n951) );
  AND U1264 ( .A(n952), .B(n951), .Z(n988) );
  XOR U1265 ( .A(n989), .B(n988), .Z(c[262]) );
  NANDN U1266 ( .A(n958), .B(n957), .Z(n962) );
  NAND U1267 ( .A(n960), .B(n959), .Z(n961) );
  NAND U1268 ( .A(n962), .B(n961), .Z(n1023) );
  NANDN U1269 ( .A(n964), .B(n963), .Z(n968) );
  NAND U1270 ( .A(n966), .B(n965), .Z(n967) );
  NAND U1271 ( .A(n968), .B(n967), .Z(n1021) );
  XNOR U1272 ( .A(b[7]), .B(a[9]), .Z(n1008) );
  NANDN U1273 ( .A(n1008), .B(n10545), .Z(n971) );
  NANDN U1274 ( .A(n969), .B(n10546), .Z(n970) );
  NAND U1275 ( .A(n971), .B(n970), .Z(n996) );
  XNOR U1276 ( .A(b[3]), .B(a[13]), .Z(n1011) );
  NANDN U1277 ( .A(n1011), .B(n10398), .Z(n974) );
  NANDN U1278 ( .A(n972), .B(n10399), .Z(n973) );
  AND U1279 ( .A(n974), .B(n973), .Z(n997) );
  XNOR U1280 ( .A(n996), .B(n997), .Z(n998) );
  NANDN U1281 ( .A(n527), .B(a[15]), .Z(n975) );
  XOR U1282 ( .A(n10434), .B(n975), .Z(n977) );
  NANDN U1283 ( .A(b[0]), .B(a[14]), .Z(n976) );
  AND U1284 ( .A(n977), .B(n976), .Z(n1004) );
  XOR U1285 ( .A(b[5]), .B(a[11]), .Z(n1017) );
  NAND U1286 ( .A(n1017), .B(n10481), .Z(n980) );
  NAND U1287 ( .A(n978), .B(n10482), .Z(n979) );
  NAND U1288 ( .A(n980), .B(n979), .Z(n1002) );
  NANDN U1289 ( .A(n529), .B(a[7]), .Z(n1003) );
  XNOR U1290 ( .A(n1002), .B(n1003), .Z(n1005) );
  XOR U1291 ( .A(n1004), .B(n1005), .Z(n999) );
  XOR U1292 ( .A(n998), .B(n999), .Z(n1020) );
  XOR U1293 ( .A(n1021), .B(n1020), .Z(n1022) );
  XNOR U1294 ( .A(n1023), .B(n1022), .Z(n992) );
  NAND U1295 ( .A(n982), .B(n981), .Z(n986) );
  NAND U1296 ( .A(n984), .B(n983), .Z(n985) );
  NAND U1297 ( .A(n986), .B(n985), .Z(n993) );
  XNOR U1298 ( .A(n992), .B(n993), .Z(n994) );
  XNOR U1299 ( .A(n995), .B(n994), .Z(n1026) );
  XNOR U1300 ( .A(n1026), .B(sreg[263]), .Z(n1028) );
  NAND U1301 ( .A(n987), .B(sreg[262]), .Z(n991) );
  OR U1302 ( .A(n989), .B(n988), .Z(n990) );
  AND U1303 ( .A(n991), .B(n990), .Z(n1027) );
  XOR U1304 ( .A(n1028), .B(n1027), .Z(c[263]) );
  NANDN U1305 ( .A(n997), .B(n996), .Z(n1001) );
  NAND U1306 ( .A(n999), .B(n998), .Z(n1000) );
  NAND U1307 ( .A(n1001), .B(n1000), .Z(n1062) );
  NANDN U1308 ( .A(n1003), .B(n1002), .Z(n1007) );
  NAND U1309 ( .A(n1005), .B(n1004), .Z(n1006) );
  NAND U1310 ( .A(n1007), .B(n1006), .Z(n1060) );
  XNOR U1311 ( .A(b[7]), .B(a[10]), .Z(n1047) );
  NANDN U1312 ( .A(n1047), .B(n10545), .Z(n1010) );
  NANDN U1313 ( .A(n1008), .B(n10546), .Z(n1009) );
  NAND U1314 ( .A(n1010), .B(n1009), .Z(n1035) );
  XNOR U1315 ( .A(b[3]), .B(a[14]), .Z(n1050) );
  NANDN U1316 ( .A(n1050), .B(n10398), .Z(n1013) );
  NANDN U1317 ( .A(n1011), .B(n10399), .Z(n1012) );
  AND U1318 ( .A(n1013), .B(n1012), .Z(n1036) );
  XNOR U1319 ( .A(n1035), .B(n1036), .Z(n1037) );
  NANDN U1320 ( .A(n527), .B(a[16]), .Z(n1014) );
  XOR U1321 ( .A(n10434), .B(n1014), .Z(n1016) );
  NANDN U1322 ( .A(b[0]), .B(a[15]), .Z(n1015) );
  AND U1323 ( .A(n1016), .B(n1015), .Z(n1043) );
  XOR U1324 ( .A(b[5]), .B(a[12]), .Z(n1056) );
  NAND U1325 ( .A(n1056), .B(n10481), .Z(n1019) );
  NAND U1326 ( .A(n1017), .B(n10482), .Z(n1018) );
  NAND U1327 ( .A(n1019), .B(n1018), .Z(n1041) );
  NANDN U1328 ( .A(n529), .B(a[8]), .Z(n1042) );
  XNOR U1329 ( .A(n1041), .B(n1042), .Z(n1044) );
  XOR U1330 ( .A(n1043), .B(n1044), .Z(n1038) );
  XOR U1331 ( .A(n1037), .B(n1038), .Z(n1059) );
  XOR U1332 ( .A(n1060), .B(n1059), .Z(n1061) );
  XNOR U1333 ( .A(n1062), .B(n1061), .Z(n1031) );
  NAND U1334 ( .A(n1021), .B(n1020), .Z(n1025) );
  NAND U1335 ( .A(n1023), .B(n1022), .Z(n1024) );
  NAND U1336 ( .A(n1025), .B(n1024), .Z(n1032) );
  XNOR U1337 ( .A(n1031), .B(n1032), .Z(n1033) );
  XNOR U1338 ( .A(n1034), .B(n1033), .Z(n1065) );
  XNOR U1339 ( .A(n1065), .B(sreg[264]), .Z(n1067) );
  NAND U1340 ( .A(n1026), .B(sreg[263]), .Z(n1030) );
  OR U1341 ( .A(n1028), .B(n1027), .Z(n1029) );
  AND U1342 ( .A(n1030), .B(n1029), .Z(n1066) );
  XOR U1343 ( .A(n1067), .B(n1066), .Z(c[264]) );
  NANDN U1344 ( .A(n1036), .B(n1035), .Z(n1040) );
  NAND U1345 ( .A(n1038), .B(n1037), .Z(n1039) );
  NAND U1346 ( .A(n1040), .B(n1039), .Z(n1101) );
  NANDN U1347 ( .A(n1042), .B(n1041), .Z(n1046) );
  NAND U1348 ( .A(n1044), .B(n1043), .Z(n1045) );
  NAND U1349 ( .A(n1046), .B(n1045), .Z(n1099) );
  XNOR U1350 ( .A(b[7]), .B(a[11]), .Z(n1092) );
  NANDN U1351 ( .A(n1092), .B(n10545), .Z(n1049) );
  NANDN U1352 ( .A(n1047), .B(n10546), .Z(n1048) );
  NAND U1353 ( .A(n1049), .B(n1048), .Z(n1074) );
  XNOR U1354 ( .A(b[3]), .B(a[15]), .Z(n1095) );
  NANDN U1355 ( .A(n1095), .B(n10398), .Z(n1052) );
  NANDN U1356 ( .A(n1050), .B(n10399), .Z(n1051) );
  AND U1357 ( .A(n1052), .B(n1051), .Z(n1075) );
  XNOR U1358 ( .A(n1074), .B(n1075), .Z(n1076) );
  NANDN U1359 ( .A(n527), .B(a[17]), .Z(n1053) );
  XOR U1360 ( .A(n10434), .B(n1053), .Z(n1055) );
  NANDN U1361 ( .A(b[0]), .B(a[16]), .Z(n1054) );
  AND U1362 ( .A(n1055), .B(n1054), .Z(n1082) );
  XOR U1363 ( .A(b[5]), .B(a[13]), .Z(n1089) );
  NAND U1364 ( .A(n1089), .B(n10481), .Z(n1058) );
  NAND U1365 ( .A(n1056), .B(n10482), .Z(n1057) );
  NAND U1366 ( .A(n1058), .B(n1057), .Z(n1080) );
  NANDN U1367 ( .A(n529), .B(a[9]), .Z(n1081) );
  XNOR U1368 ( .A(n1080), .B(n1081), .Z(n1083) );
  XOR U1369 ( .A(n1082), .B(n1083), .Z(n1077) );
  XOR U1370 ( .A(n1076), .B(n1077), .Z(n1098) );
  XOR U1371 ( .A(n1099), .B(n1098), .Z(n1100) );
  XNOR U1372 ( .A(n1101), .B(n1100), .Z(n1070) );
  NAND U1373 ( .A(n1060), .B(n1059), .Z(n1064) );
  NAND U1374 ( .A(n1062), .B(n1061), .Z(n1063) );
  NAND U1375 ( .A(n1064), .B(n1063), .Z(n1071) );
  XNOR U1376 ( .A(n1070), .B(n1071), .Z(n1072) );
  XNOR U1377 ( .A(n1073), .B(n1072), .Z(n1104) );
  XNOR U1378 ( .A(n1104), .B(sreg[265]), .Z(n1106) );
  NAND U1379 ( .A(n1065), .B(sreg[264]), .Z(n1069) );
  OR U1380 ( .A(n1067), .B(n1066), .Z(n1068) );
  AND U1381 ( .A(n1069), .B(n1068), .Z(n1105) );
  XOR U1382 ( .A(n1106), .B(n1105), .Z(c[265]) );
  NANDN U1383 ( .A(n1075), .B(n1074), .Z(n1079) );
  NAND U1384 ( .A(n1077), .B(n1076), .Z(n1078) );
  NAND U1385 ( .A(n1079), .B(n1078), .Z(n1140) );
  NANDN U1386 ( .A(n1081), .B(n1080), .Z(n1085) );
  NAND U1387 ( .A(n1083), .B(n1082), .Z(n1084) );
  NAND U1388 ( .A(n1085), .B(n1084), .Z(n1138) );
  NANDN U1389 ( .A(n527), .B(a[18]), .Z(n1086) );
  XOR U1390 ( .A(n10434), .B(n1086), .Z(n1088) );
  NANDN U1391 ( .A(b[0]), .B(a[17]), .Z(n1087) );
  AND U1392 ( .A(n1088), .B(n1087), .Z(n1121) );
  XOR U1393 ( .A(b[5]), .B(a[14]), .Z(n1125) );
  NAND U1394 ( .A(n1125), .B(n10481), .Z(n1091) );
  NAND U1395 ( .A(n1089), .B(n10482), .Z(n1090) );
  NAND U1396 ( .A(n1091), .B(n1090), .Z(n1119) );
  NANDN U1397 ( .A(n529), .B(a[10]), .Z(n1120) );
  XNOR U1398 ( .A(n1119), .B(n1120), .Z(n1122) );
  XOR U1399 ( .A(n1121), .B(n1122), .Z(n1115) );
  XNOR U1400 ( .A(b[7]), .B(a[12]), .Z(n1131) );
  NANDN U1401 ( .A(n1131), .B(n10545), .Z(n1094) );
  NANDN U1402 ( .A(n1092), .B(n10546), .Z(n1093) );
  NAND U1403 ( .A(n1094), .B(n1093), .Z(n1113) );
  XNOR U1404 ( .A(b[3]), .B(a[16]), .Z(n1134) );
  NANDN U1405 ( .A(n1134), .B(n10398), .Z(n1097) );
  NANDN U1406 ( .A(n1095), .B(n10399), .Z(n1096) );
  AND U1407 ( .A(n1097), .B(n1096), .Z(n1114) );
  XNOR U1408 ( .A(n1113), .B(n1114), .Z(n1116) );
  XOR U1409 ( .A(n1115), .B(n1116), .Z(n1137) );
  XOR U1410 ( .A(n1138), .B(n1137), .Z(n1139) );
  XNOR U1411 ( .A(n1140), .B(n1139), .Z(n1109) );
  NAND U1412 ( .A(n1099), .B(n1098), .Z(n1103) );
  NAND U1413 ( .A(n1101), .B(n1100), .Z(n1102) );
  NAND U1414 ( .A(n1103), .B(n1102), .Z(n1110) );
  XNOR U1415 ( .A(n1109), .B(n1110), .Z(n1111) );
  XNOR U1416 ( .A(n1112), .B(n1111), .Z(n1143) );
  XNOR U1417 ( .A(n1143), .B(sreg[266]), .Z(n1145) );
  NAND U1418 ( .A(n1104), .B(sreg[265]), .Z(n1108) );
  OR U1419 ( .A(n1106), .B(n1105), .Z(n1107) );
  AND U1420 ( .A(n1108), .B(n1107), .Z(n1144) );
  XOR U1421 ( .A(n1145), .B(n1144), .Z(c[266]) );
  NANDN U1422 ( .A(n1114), .B(n1113), .Z(n1118) );
  NAND U1423 ( .A(n1116), .B(n1115), .Z(n1117) );
  NAND U1424 ( .A(n1118), .B(n1117), .Z(n1179) );
  NANDN U1425 ( .A(n1120), .B(n1119), .Z(n1124) );
  NAND U1426 ( .A(n1122), .B(n1121), .Z(n1123) );
  NAND U1427 ( .A(n1124), .B(n1123), .Z(n1177) );
  XOR U1428 ( .A(b[5]), .B(a[15]), .Z(n1161) );
  NAND U1429 ( .A(n10481), .B(n1161), .Z(n1127) );
  NAND U1430 ( .A(n10482), .B(n1125), .Z(n1126) );
  AND U1431 ( .A(n1127), .B(n1126), .Z(n1170) );
  NANDN U1432 ( .A(n529), .B(a[11]), .Z(n1171) );
  XOR U1433 ( .A(n1170), .B(n1171), .Z(n1173) );
  NANDN U1434 ( .A(n527), .B(a[19]), .Z(n1128) );
  XOR U1435 ( .A(n10434), .B(n1128), .Z(n1130) );
  NANDN U1436 ( .A(b[0]), .B(a[18]), .Z(n1129) );
  AND U1437 ( .A(n1130), .B(n1129), .Z(n1172) );
  XNOR U1438 ( .A(n1173), .B(n1172), .Z(n1167) );
  XNOR U1439 ( .A(b[7]), .B(a[13]), .Z(n1152) );
  NANDN U1440 ( .A(n1152), .B(n10545), .Z(n1133) );
  NANDN U1441 ( .A(n1131), .B(n10546), .Z(n1132) );
  NAND U1442 ( .A(n1133), .B(n1132), .Z(n1164) );
  XNOR U1443 ( .A(b[3]), .B(a[17]), .Z(n1155) );
  NANDN U1444 ( .A(n1155), .B(n10398), .Z(n1136) );
  NANDN U1445 ( .A(n1134), .B(n10399), .Z(n1135) );
  AND U1446 ( .A(n1136), .B(n1135), .Z(n1165) );
  XNOR U1447 ( .A(n1164), .B(n1165), .Z(n1166) );
  XNOR U1448 ( .A(n1167), .B(n1166), .Z(n1176) );
  XOR U1449 ( .A(n1177), .B(n1176), .Z(n1178) );
  XNOR U1450 ( .A(n1179), .B(n1178), .Z(n1148) );
  NAND U1451 ( .A(n1138), .B(n1137), .Z(n1142) );
  NAND U1452 ( .A(n1140), .B(n1139), .Z(n1141) );
  NAND U1453 ( .A(n1142), .B(n1141), .Z(n1149) );
  XNOR U1454 ( .A(n1148), .B(n1149), .Z(n1150) );
  XNOR U1455 ( .A(n1151), .B(n1150), .Z(n1180) );
  XNOR U1456 ( .A(n1180), .B(sreg[267]), .Z(n1182) );
  NAND U1457 ( .A(n1143), .B(sreg[266]), .Z(n1147) );
  OR U1458 ( .A(n1145), .B(n1144), .Z(n1146) );
  AND U1459 ( .A(n1147), .B(n1146), .Z(n1181) );
  XOR U1460 ( .A(n1182), .B(n1181), .Z(c[267]) );
  XNOR U1461 ( .A(b[7]), .B(a[14]), .Z(n1201) );
  NANDN U1462 ( .A(n1201), .B(n10545), .Z(n1154) );
  NANDN U1463 ( .A(n1152), .B(n10546), .Z(n1153) );
  NAND U1464 ( .A(n1154), .B(n1153), .Z(n1189) );
  XNOR U1465 ( .A(b[3]), .B(a[18]), .Z(n1204) );
  NANDN U1466 ( .A(n1204), .B(n10398), .Z(n1157) );
  NANDN U1467 ( .A(n1155), .B(n10399), .Z(n1156) );
  AND U1468 ( .A(n1157), .B(n1156), .Z(n1190) );
  XNOR U1469 ( .A(n1189), .B(n1190), .Z(n1191) );
  NANDN U1470 ( .A(n527), .B(a[20]), .Z(n1158) );
  XOR U1471 ( .A(n10434), .B(n1158), .Z(n1160) );
  NANDN U1472 ( .A(b[0]), .B(a[19]), .Z(n1159) );
  AND U1473 ( .A(n1160), .B(n1159), .Z(n1197) );
  XOR U1474 ( .A(b[5]), .B(a[16]), .Z(n1210) );
  NAND U1475 ( .A(n1210), .B(n10481), .Z(n1163) );
  NAND U1476 ( .A(n1161), .B(n10482), .Z(n1162) );
  NAND U1477 ( .A(n1163), .B(n1162), .Z(n1195) );
  NANDN U1478 ( .A(n529), .B(a[12]), .Z(n1196) );
  XNOR U1479 ( .A(n1195), .B(n1196), .Z(n1198) );
  XOR U1480 ( .A(n1197), .B(n1198), .Z(n1192) );
  XOR U1481 ( .A(n1191), .B(n1192), .Z(n1215) );
  NANDN U1482 ( .A(n1165), .B(n1164), .Z(n1169) );
  NANDN U1483 ( .A(n1167), .B(n1166), .Z(n1168) );
  NAND U1484 ( .A(n1169), .B(n1168), .Z(n1213) );
  OR U1485 ( .A(n1171), .B(n1170), .Z(n1175) );
  NAND U1486 ( .A(n1173), .B(n1172), .Z(n1174) );
  AND U1487 ( .A(n1175), .B(n1174), .Z(n1214) );
  XNOR U1488 ( .A(n1213), .B(n1214), .Z(n1216) );
  XNOR U1489 ( .A(n1215), .B(n1216), .Z(n1185) );
  XNOR U1490 ( .A(n1185), .B(n1186), .Z(n1187) );
  XNOR U1491 ( .A(n1188), .B(n1187), .Z(n1219) );
  XNOR U1492 ( .A(n1219), .B(sreg[268]), .Z(n1221) );
  NAND U1493 ( .A(n1180), .B(sreg[267]), .Z(n1184) );
  OR U1494 ( .A(n1182), .B(n1181), .Z(n1183) );
  AND U1495 ( .A(n1184), .B(n1183), .Z(n1220) );
  XOR U1496 ( .A(n1221), .B(n1220), .Z(c[268]) );
  NANDN U1497 ( .A(n1190), .B(n1189), .Z(n1194) );
  NAND U1498 ( .A(n1192), .B(n1191), .Z(n1193) );
  NAND U1499 ( .A(n1194), .B(n1193), .Z(n1255) );
  NANDN U1500 ( .A(n1196), .B(n1195), .Z(n1200) );
  NAND U1501 ( .A(n1198), .B(n1197), .Z(n1199) );
  NAND U1502 ( .A(n1200), .B(n1199), .Z(n1253) );
  XNOR U1503 ( .A(b[7]), .B(a[15]), .Z(n1240) );
  NANDN U1504 ( .A(n1240), .B(n10545), .Z(n1203) );
  NANDN U1505 ( .A(n1201), .B(n10546), .Z(n1202) );
  NAND U1506 ( .A(n1203), .B(n1202), .Z(n1228) );
  XNOR U1507 ( .A(b[3]), .B(a[19]), .Z(n1243) );
  NANDN U1508 ( .A(n1243), .B(n10398), .Z(n1206) );
  NANDN U1509 ( .A(n1204), .B(n10399), .Z(n1205) );
  AND U1510 ( .A(n1206), .B(n1205), .Z(n1229) );
  XNOR U1511 ( .A(n1228), .B(n1229), .Z(n1230) );
  NANDN U1512 ( .A(n527), .B(a[21]), .Z(n1207) );
  XOR U1513 ( .A(n10434), .B(n1207), .Z(n1209) );
  NANDN U1514 ( .A(b[0]), .B(a[20]), .Z(n1208) );
  AND U1515 ( .A(n1209), .B(n1208), .Z(n1236) );
  XOR U1516 ( .A(b[5]), .B(a[17]), .Z(n1249) );
  NAND U1517 ( .A(n1249), .B(n10481), .Z(n1212) );
  NAND U1518 ( .A(n1210), .B(n10482), .Z(n1211) );
  NAND U1519 ( .A(n1212), .B(n1211), .Z(n1234) );
  NANDN U1520 ( .A(n529), .B(a[13]), .Z(n1235) );
  XNOR U1521 ( .A(n1234), .B(n1235), .Z(n1237) );
  XOR U1522 ( .A(n1236), .B(n1237), .Z(n1231) );
  XOR U1523 ( .A(n1230), .B(n1231), .Z(n1252) );
  XOR U1524 ( .A(n1253), .B(n1252), .Z(n1254) );
  XNOR U1525 ( .A(n1255), .B(n1254), .Z(n1224) );
  NANDN U1526 ( .A(n1214), .B(n1213), .Z(n1218) );
  NAND U1527 ( .A(n1216), .B(n1215), .Z(n1217) );
  NAND U1528 ( .A(n1218), .B(n1217), .Z(n1225) );
  XNOR U1529 ( .A(n1224), .B(n1225), .Z(n1226) );
  XNOR U1530 ( .A(n1227), .B(n1226), .Z(n1258) );
  XNOR U1531 ( .A(n1258), .B(sreg[269]), .Z(n1260) );
  NAND U1532 ( .A(n1219), .B(sreg[268]), .Z(n1223) );
  OR U1533 ( .A(n1221), .B(n1220), .Z(n1222) );
  AND U1534 ( .A(n1223), .B(n1222), .Z(n1259) );
  XOR U1535 ( .A(n1260), .B(n1259), .Z(c[269]) );
  NANDN U1536 ( .A(n1229), .B(n1228), .Z(n1233) );
  NAND U1537 ( .A(n1231), .B(n1230), .Z(n1232) );
  NAND U1538 ( .A(n1233), .B(n1232), .Z(n1294) );
  NANDN U1539 ( .A(n1235), .B(n1234), .Z(n1239) );
  NAND U1540 ( .A(n1237), .B(n1236), .Z(n1238) );
  NAND U1541 ( .A(n1239), .B(n1238), .Z(n1292) );
  XNOR U1542 ( .A(b[7]), .B(a[16]), .Z(n1279) );
  NANDN U1543 ( .A(n1279), .B(n10545), .Z(n1242) );
  NANDN U1544 ( .A(n1240), .B(n10546), .Z(n1241) );
  NAND U1545 ( .A(n1242), .B(n1241), .Z(n1267) );
  XNOR U1546 ( .A(b[3]), .B(a[20]), .Z(n1282) );
  NANDN U1547 ( .A(n1282), .B(n10398), .Z(n1245) );
  NANDN U1548 ( .A(n1243), .B(n10399), .Z(n1244) );
  AND U1549 ( .A(n1245), .B(n1244), .Z(n1268) );
  XNOR U1550 ( .A(n1267), .B(n1268), .Z(n1269) );
  NANDN U1551 ( .A(n527), .B(a[22]), .Z(n1246) );
  XOR U1552 ( .A(n10434), .B(n1246), .Z(n1248) );
  NANDN U1553 ( .A(b[0]), .B(a[21]), .Z(n1247) );
  AND U1554 ( .A(n1248), .B(n1247), .Z(n1275) );
  XOR U1555 ( .A(b[5]), .B(a[18]), .Z(n1288) );
  NAND U1556 ( .A(n1288), .B(n10481), .Z(n1251) );
  NAND U1557 ( .A(n1249), .B(n10482), .Z(n1250) );
  NAND U1558 ( .A(n1251), .B(n1250), .Z(n1273) );
  NANDN U1559 ( .A(n529), .B(a[14]), .Z(n1274) );
  XNOR U1560 ( .A(n1273), .B(n1274), .Z(n1276) );
  XOR U1561 ( .A(n1275), .B(n1276), .Z(n1270) );
  XOR U1562 ( .A(n1269), .B(n1270), .Z(n1291) );
  XOR U1563 ( .A(n1292), .B(n1291), .Z(n1293) );
  XNOR U1564 ( .A(n1294), .B(n1293), .Z(n1263) );
  NAND U1565 ( .A(n1253), .B(n1252), .Z(n1257) );
  NAND U1566 ( .A(n1255), .B(n1254), .Z(n1256) );
  NAND U1567 ( .A(n1257), .B(n1256), .Z(n1264) );
  XNOR U1568 ( .A(n1263), .B(n1264), .Z(n1265) );
  XNOR U1569 ( .A(n1266), .B(n1265), .Z(n1297) );
  XNOR U1570 ( .A(n1297), .B(sreg[270]), .Z(n1299) );
  NAND U1571 ( .A(n1258), .B(sreg[269]), .Z(n1262) );
  OR U1572 ( .A(n1260), .B(n1259), .Z(n1261) );
  AND U1573 ( .A(n1262), .B(n1261), .Z(n1298) );
  XOR U1574 ( .A(n1299), .B(n1298), .Z(c[270]) );
  NANDN U1575 ( .A(n1268), .B(n1267), .Z(n1272) );
  NAND U1576 ( .A(n1270), .B(n1269), .Z(n1271) );
  NAND U1577 ( .A(n1272), .B(n1271), .Z(n1333) );
  NANDN U1578 ( .A(n1274), .B(n1273), .Z(n1278) );
  NAND U1579 ( .A(n1276), .B(n1275), .Z(n1277) );
  NAND U1580 ( .A(n1278), .B(n1277), .Z(n1331) );
  XNOR U1581 ( .A(b[7]), .B(a[17]), .Z(n1318) );
  NANDN U1582 ( .A(n1318), .B(n10545), .Z(n1281) );
  NANDN U1583 ( .A(n1279), .B(n10546), .Z(n1280) );
  NAND U1584 ( .A(n1281), .B(n1280), .Z(n1306) );
  XNOR U1585 ( .A(b[3]), .B(a[21]), .Z(n1321) );
  NANDN U1586 ( .A(n1321), .B(n10398), .Z(n1284) );
  NANDN U1587 ( .A(n1282), .B(n10399), .Z(n1283) );
  AND U1588 ( .A(n1284), .B(n1283), .Z(n1307) );
  XNOR U1589 ( .A(n1306), .B(n1307), .Z(n1308) );
  NANDN U1590 ( .A(n527), .B(a[23]), .Z(n1285) );
  XOR U1591 ( .A(n10434), .B(n1285), .Z(n1287) );
  NANDN U1592 ( .A(b[0]), .B(a[22]), .Z(n1286) );
  AND U1593 ( .A(n1287), .B(n1286), .Z(n1314) );
  XOR U1594 ( .A(b[5]), .B(a[19]), .Z(n1327) );
  NAND U1595 ( .A(n1327), .B(n10481), .Z(n1290) );
  NAND U1596 ( .A(n1288), .B(n10482), .Z(n1289) );
  NAND U1597 ( .A(n1290), .B(n1289), .Z(n1312) );
  NANDN U1598 ( .A(n529), .B(a[15]), .Z(n1313) );
  XNOR U1599 ( .A(n1312), .B(n1313), .Z(n1315) );
  XOR U1600 ( .A(n1314), .B(n1315), .Z(n1309) );
  XOR U1601 ( .A(n1308), .B(n1309), .Z(n1330) );
  XOR U1602 ( .A(n1331), .B(n1330), .Z(n1332) );
  XNOR U1603 ( .A(n1333), .B(n1332), .Z(n1302) );
  NAND U1604 ( .A(n1292), .B(n1291), .Z(n1296) );
  NAND U1605 ( .A(n1294), .B(n1293), .Z(n1295) );
  NAND U1606 ( .A(n1296), .B(n1295), .Z(n1303) );
  XNOR U1607 ( .A(n1302), .B(n1303), .Z(n1304) );
  XNOR U1608 ( .A(n1305), .B(n1304), .Z(n1336) );
  XNOR U1609 ( .A(n1336), .B(sreg[271]), .Z(n1338) );
  NAND U1610 ( .A(n1297), .B(sreg[270]), .Z(n1301) );
  OR U1611 ( .A(n1299), .B(n1298), .Z(n1300) );
  AND U1612 ( .A(n1301), .B(n1300), .Z(n1337) );
  XOR U1613 ( .A(n1338), .B(n1337), .Z(c[271]) );
  NANDN U1614 ( .A(n1307), .B(n1306), .Z(n1311) );
  NAND U1615 ( .A(n1309), .B(n1308), .Z(n1310) );
  NAND U1616 ( .A(n1311), .B(n1310), .Z(n1372) );
  NANDN U1617 ( .A(n1313), .B(n1312), .Z(n1317) );
  NAND U1618 ( .A(n1315), .B(n1314), .Z(n1316) );
  NAND U1619 ( .A(n1317), .B(n1316), .Z(n1370) );
  XNOR U1620 ( .A(b[7]), .B(a[18]), .Z(n1357) );
  NANDN U1621 ( .A(n1357), .B(n10545), .Z(n1320) );
  NANDN U1622 ( .A(n1318), .B(n10546), .Z(n1319) );
  NAND U1623 ( .A(n1320), .B(n1319), .Z(n1345) );
  XNOR U1624 ( .A(b[3]), .B(a[22]), .Z(n1360) );
  NANDN U1625 ( .A(n1360), .B(n10398), .Z(n1323) );
  NANDN U1626 ( .A(n1321), .B(n10399), .Z(n1322) );
  AND U1627 ( .A(n1323), .B(n1322), .Z(n1346) );
  XNOR U1628 ( .A(n1345), .B(n1346), .Z(n1347) );
  NANDN U1629 ( .A(n527), .B(a[24]), .Z(n1324) );
  XOR U1630 ( .A(n10434), .B(n1324), .Z(n1326) );
  NANDN U1631 ( .A(b[0]), .B(a[23]), .Z(n1325) );
  AND U1632 ( .A(n1326), .B(n1325), .Z(n1353) );
  XOR U1633 ( .A(b[5]), .B(a[20]), .Z(n1366) );
  NAND U1634 ( .A(n1366), .B(n10481), .Z(n1329) );
  NAND U1635 ( .A(n1327), .B(n10482), .Z(n1328) );
  NAND U1636 ( .A(n1329), .B(n1328), .Z(n1351) );
  NANDN U1637 ( .A(n529), .B(a[16]), .Z(n1352) );
  XNOR U1638 ( .A(n1351), .B(n1352), .Z(n1354) );
  XOR U1639 ( .A(n1353), .B(n1354), .Z(n1348) );
  XOR U1640 ( .A(n1347), .B(n1348), .Z(n1369) );
  XOR U1641 ( .A(n1370), .B(n1369), .Z(n1371) );
  XNOR U1642 ( .A(n1372), .B(n1371), .Z(n1341) );
  NAND U1643 ( .A(n1331), .B(n1330), .Z(n1335) );
  NAND U1644 ( .A(n1333), .B(n1332), .Z(n1334) );
  NAND U1645 ( .A(n1335), .B(n1334), .Z(n1342) );
  XNOR U1646 ( .A(n1341), .B(n1342), .Z(n1343) );
  XNOR U1647 ( .A(n1344), .B(n1343), .Z(n1375) );
  XNOR U1648 ( .A(n1375), .B(sreg[272]), .Z(n1377) );
  NAND U1649 ( .A(n1336), .B(sreg[271]), .Z(n1340) );
  OR U1650 ( .A(n1338), .B(n1337), .Z(n1339) );
  AND U1651 ( .A(n1340), .B(n1339), .Z(n1376) );
  XOR U1652 ( .A(n1377), .B(n1376), .Z(c[272]) );
  NANDN U1653 ( .A(n1346), .B(n1345), .Z(n1350) );
  NAND U1654 ( .A(n1348), .B(n1347), .Z(n1349) );
  NAND U1655 ( .A(n1350), .B(n1349), .Z(n1411) );
  NANDN U1656 ( .A(n1352), .B(n1351), .Z(n1356) );
  NAND U1657 ( .A(n1354), .B(n1353), .Z(n1355) );
  NAND U1658 ( .A(n1356), .B(n1355), .Z(n1409) );
  XNOR U1659 ( .A(b[7]), .B(a[19]), .Z(n1396) );
  NANDN U1660 ( .A(n1396), .B(n10545), .Z(n1359) );
  NANDN U1661 ( .A(n1357), .B(n10546), .Z(n1358) );
  NAND U1662 ( .A(n1359), .B(n1358), .Z(n1384) );
  XNOR U1663 ( .A(b[3]), .B(a[23]), .Z(n1399) );
  NANDN U1664 ( .A(n1399), .B(n10398), .Z(n1362) );
  NANDN U1665 ( .A(n1360), .B(n10399), .Z(n1361) );
  AND U1666 ( .A(n1362), .B(n1361), .Z(n1385) );
  XNOR U1667 ( .A(n1384), .B(n1385), .Z(n1386) );
  NANDN U1668 ( .A(n527), .B(a[25]), .Z(n1363) );
  XOR U1669 ( .A(n10434), .B(n1363), .Z(n1365) );
  NANDN U1670 ( .A(b[0]), .B(a[24]), .Z(n1364) );
  AND U1671 ( .A(n1365), .B(n1364), .Z(n1392) );
  XOR U1672 ( .A(b[5]), .B(a[21]), .Z(n1405) );
  NAND U1673 ( .A(n1405), .B(n10481), .Z(n1368) );
  NAND U1674 ( .A(n1366), .B(n10482), .Z(n1367) );
  NAND U1675 ( .A(n1368), .B(n1367), .Z(n1390) );
  NANDN U1676 ( .A(n529), .B(a[17]), .Z(n1391) );
  XNOR U1677 ( .A(n1390), .B(n1391), .Z(n1393) );
  XOR U1678 ( .A(n1392), .B(n1393), .Z(n1387) );
  XOR U1679 ( .A(n1386), .B(n1387), .Z(n1408) );
  XOR U1680 ( .A(n1409), .B(n1408), .Z(n1410) );
  XNOR U1681 ( .A(n1411), .B(n1410), .Z(n1380) );
  NAND U1682 ( .A(n1370), .B(n1369), .Z(n1374) );
  NAND U1683 ( .A(n1372), .B(n1371), .Z(n1373) );
  NAND U1684 ( .A(n1374), .B(n1373), .Z(n1381) );
  XNOR U1685 ( .A(n1380), .B(n1381), .Z(n1382) );
  XNOR U1686 ( .A(n1383), .B(n1382), .Z(n1414) );
  XNOR U1687 ( .A(n1414), .B(sreg[273]), .Z(n1416) );
  NAND U1688 ( .A(n1375), .B(sreg[272]), .Z(n1379) );
  OR U1689 ( .A(n1377), .B(n1376), .Z(n1378) );
  AND U1690 ( .A(n1379), .B(n1378), .Z(n1415) );
  XOR U1691 ( .A(n1416), .B(n1415), .Z(c[273]) );
  NANDN U1692 ( .A(n1385), .B(n1384), .Z(n1389) );
  NAND U1693 ( .A(n1387), .B(n1386), .Z(n1388) );
  NAND U1694 ( .A(n1389), .B(n1388), .Z(n1450) );
  NANDN U1695 ( .A(n1391), .B(n1390), .Z(n1395) );
  NAND U1696 ( .A(n1393), .B(n1392), .Z(n1394) );
  NAND U1697 ( .A(n1395), .B(n1394), .Z(n1448) );
  XNOR U1698 ( .A(b[7]), .B(a[20]), .Z(n1435) );
  NANDN U1699 ( .A(n1435), .B(n10545), .Z(n1398) );
  NANDN U1700 ( .A(n1396), .B(n10546), .Z(n1397) );
  NAND U1701 ( .A(n1398), .B(n1397), .Z(n1423) );
  XNOR U1702 ( .A(b[3]), .B(a[24]), .Z(n1438) );
  NANDN U1703 ( .A(n1438), .B(n10398), .Z(n1401) );
  NANDN U1704 ( .A(n1399), .B(n10399), .Z(n1400) );
  AND U1705 ( .A(n1401), .B(n1400), .Z(n1424) );
  XNOR U1706 ( .A(n1423), .B(n1424), .Z(n1425) );
  NANDN U1707 ( .A(n527), .B(a[26]), .Z(n1402) );
  XOR U1708 ( .A(n10434), .B(n1402), .Z(n1404) );
  NANDN U1709 ( .A(b[0]), .B(a[25]), .Z(n1403) );
  AND U1710 ( .A(n1404), .B(n1403), .Z(n1431) );
  XOR U1711 ( .A(b[5]), .B(a[22]), .Z(n1444) );
  NAND U1712 ( .A(n1444), .B(n10481), .Z(n1407) );
  NAND U1713 ( .A(n1405), .B(n10482), .Z(n1406) );
  NAND U1714 ( .A(n1407), .B(n1406), .Z(n1429) );
  NANDN U1715 ( .A(n529), .B(a[18]), .Z(n1430) );
  XNOR U1716 ( .A(n1429), .B(n1430), .Z(n1432) );
  XOR U1717 ( .A(n1431), .B(n1432), .Z(n1426) );
  XOR U1718 ( .A(n1425), .B(n1426), .Z(n1447) );
  XOR U1719 ( .A(n1448), .B(n1447), .Z(n1449) );
  XNOR U1720 ( .A(n1450), .B(n1449), .Z(n1419) );
  NAND U1721 ( .A(n1409), .B(n1408), .Z(n1413) );
  NAND U1722 ( .A(n1411), .B(n1410), .Z(n1412) );
  NAND U1723 ( .A(n1413), .B(n1412), .Z(n1420) );
  XNOR U1724 ( .A(n1419), .B(n1420), .Z(n1421) );
  XNOR U1725 ( .A(n1422), .B(n1421), .Z(n1453) );
  XNOR U1726 ( .A(n1453), .B(sreg[274]), .Z(n1455) );
  NAND U1727 ( .A(n1414), .B(sreg[273]), .Z(n1418) );
  OR U1728 ( .A(n1416), .B(n1415), .Z(n1417) );
  AND U1729 ( .A(n1418), .B(n1417), .Z(n1454) );
  XOR U1730 ( .A(n1455), .B(n1454), .Z(c[274]) );
  NANDN U1731 ( .A(n1424), .B(n1423), .Z(n1428) );
  NAND U1732 ( .A(n1426), .B(n1425), .Z(n1427) );
  NAND U1733 ( .A(n1428), .B(n1427), .Z(n1489) );
  NANDN U1734 ( .A(n1430), .B(n1429), .Z(n1434) );
  NAND U1735 ( .A(n1432), .B(n1431), .Z(n1433) );
  NAND U1736 ( .A(n1434), .B(n1433), .Z(n1487) );
  XNOR U1737 ( .A(b[7]), .B(a[21]), .Z(n1474) );
  NANDN U1738 ( .A(n1474), .B(n10545), .Z(n1437) );
  NANDN U1739 ( .A(n1435), .B(n10546), .Z(n1436) );
  NAND U1740 ( .A(n1437), .B(n1436), .Z(n1462) );
  XNOR U1741 ( .A(b[3]), .B(a[25]), .Z(n1477) );
  NANDN U1742 ( .A(n1477), .B(n10398), .Z(n1440) );
  NANDN U1743 ( .A(n1438), .B(n10399), .Z(n1439) );
  AND U1744 ( .A(n1440), .B(n1439), .Z(n1463) );
  XNOR U1745 ( .A(n1462), .B(n1463), .Z(n1464) );
  NANDN U1746 ( .A(n527), .B(a[27]), .Z(n1441) );
  XOR U1747 ( .A(n10434), .B(n1441), .Z(n1443) );
  NANDN U1748 ( .A(b[0]), .B(a[26]), .Z(n1442) );
  AND U1749 ( .A(n1443), .B(n1442), .Z(n1470) );
  XOR U1750 ( .A(b[5]), .B(a[23]), .Z(n1483) );
  NAND U1751 ( .A(n1483), .B(n10481), .Z(n1446) );
  NAND U1752 ( .A(n1444), .B(n10482), .Z(n1445) );
  NAND U1753 ( .A(n1446), .B(n1445), .Z(n1468) );
  NANDN U1754 ( .A(n529), .B(a[19]), .Z(n1469) );
  XNOR U1755 ( .A(n1468), .B(n1469), .Z(n1471) );
  XOR U1756 ( .A(n1470), .B(n1471), .Z(n1465) );
  XOR U1757 ( .A(n1464), .B(n1465), .Z(n1486) );
  XOR U1758 ( .A(n1487), .B(n1486), .Z(n1488) );
  XNOR U1759 ( .A(n1489), .B(n1488), .Z(n1458) );
  NAND U1760 ( .A(n1448), .B(n1447), .Z(n1452) );
  NAND U1761 ( .A(n1450), .B(n1449), .Z(n1451) );
  NAND U1762 ( .A(n1452), .B(n1451), .Z(n1459) );
  XNOR U1763 ( .A(n1458), .B(n1459), .Z(n1460) );
  XNOR U1764 ( .A(n1461), .B(n1460), .Z(n1492) );
  XNOR U1765 ( .A(n1492), .B(sreg[275]), .Z(n1494) );
  NAND U1766 ( .A(n1453), .B(sreg[274]), .Z(n1457) );
  OR U1767 ( .A(n1455), .B(n1454), .Z(n1456) );
  AND U1768 ( .A(n1457), .B(n1456), .Z(n1493) );
  XOR U1769 ( .A(n1494), .B(n1493), .Z(c[275]) );
  NANDN U1770 ( .A(n1463), .B(n1462), .Z(n1467) );
  NAND U1771 ( .A(n1465), .B(n1464), .Z(n1466) );
  NAND U1772 ( .A(n1467), .B(n1466), .Z(n1528) );
  NANDN U1773 ( .A(n1469), .B(n1468), .Z(n1473) );
  NAND U1774 ( .A(n1471), .B(n1470), .Z(n1472) );
  NAND U1775 ( .A(n1473), .B(n1472), .Z(n1526) );
  XNOR U1776 ( .A(b[7]), .B(a[22]), .Z(n1513) );
  NANDN U1777 ( .A(n1513), .B(n10545), .Z(n1476) );
  NANDN U1778 ( .A(n1474), .B(n10546), .Z(n1475) );
  NAND U1779 ( .A(n1476), .B(n1475), .Z(n1501) );
  XNOR U1780 ( .A(b[3]), .B(a[26]), .Z(n1516) );
  NANDN U1781 ( .A(n1516), .B(n10398), .Z(n1479) );
  NANDN U1782 ( .A(n1477), .B(n10399), .Z(n1478) );
  AND U1783 ( .A(n1479), .B(n1478), .Z(n1502) );
  XNOR U1784 ( .A(n1501), .B(n1502), .Z(n1503) );
  NANDN U1785 ( .A(n527), .B(a[28]), .Z(n1480) );
  XOR U1786 ( .A(n10434), .B(n1480), .Z(n1482) );
  NANDN U1787 ( .A(b[0]), .B(a[27]), .Z(n1481) );
  AND U1788 ( .A(n1482), .B(n1481), .Z(n1509) );
  XOR U1789 ( .A(b[5]), .B(a[24]), .Z(n1522) );
  NAND U1790 ( .A(n1522), .B(n10481), .Z(n1485) );
  NAND U1791 ( .A(n1483), .B(n10482), .Z(n1484) );
  NAND U1792 ( .A(n1485), .B(n1484), .Z(n1507) );
  NANDN U1793 ( .A(n529), .B(a[20]), .Z(n1508) );
  XNOR U1794 ( .A(n1507), .B(n1508), .Z(n1510) );
  XOR U1795 ( .A(n1509), .B(n1510), .Z(n1504) );
  XOR U1796 ( .A(n1503), .B(n1504), .Z(n1525) );
  XOR U1797 ( .A(n1526), .B(n1525), .Z(n1527) );
  XNOR U1798 ( .A(n1528), .B(n1527), .Z(n1497) );
  NAND U1799 ( .A(n1487), .B(n1486), .Z(n1491) );
  NAND U1800 ( .A(n1489), .B(n1488), .Z(n1490) );
  NAND U1801 ( .A(n1491), .B(n1490), .Z(n1498) );
  XNOR U1802 ( .A(n1497), .B(n1498), .Z(n1499) );
  XNOR U1803 ( .A(n1500), .B(n1499), .Z(n1531) );
  XNOR U1804 ( .A(n1531), .B(sreg[276]), .Z(n1533) );
  NAND U1805 ( .A(n1492), .B(sreg[275]), .Z(n1496) );
  OR U1806 ( .A(n1494), .B(n1493), .Z(n1495) );
  AND U1807 ( .A(n1496), .B(n1495), .Z(n1532) );
  XOR U1808 ( .A(n1533), .B(n1532), .Z(c[276]) );
  NANDN U1809 ( .A(n1502), .B(n1501), .Z(n1506) );
  NAND U1810 ( .A(n1504), .B(n1503), .Z(n1505) );
  NAND U1811 ( .A(n1506), .B(n1505), .Z(n1567) );
  NANDN U1812 ( .A(n1508), .B(n1507), .Z(n1512) );
  NAND U1813 ( .A(n1510), .B(n1509), .Z(n1511) );
  NAND U1814 ( .A(n1512), .B(n1511), .Z(n1565) );
  XNOR U1815 ( .A(b[7]), .B(a[23]), .Z(n1552) );
  NANDN U1816 ( .A(n1552), .B(n10545), .Z(n1515) );
  NANDN U1817 ( .A(n1513), .B(n10546), .Z(n1514) );
  NAND U1818 ( .A(n1515), .B(n1514), .Z(n1540) );
  XNOR U1819 ( .A(b[3]), .B(a[27]), .Z(n1555) );
  NANDN U1820 ( .A(n1555), .B(n10398), .Z(n1518) );
  NANDN U1821 ( .A(n1516), .B(n10399), .Z(n1517) );
  AND U1822 ( .A(n1518), .B(n1517), .Z(n1541) );
  XNOR U1823 ( .A(n1540), .B(n1541), .Z(n1542) );
  NANDN U1824 ( .A(n527), .B(a[29]), .Z(n1519) );
  XOR U1825 ( .A(n10434), .B(n1519), .Z(n1521) );
  NANDN U1826 ( .A(b[0]), .B(a[28]), .Z(n1520) );
  AND U1827 ( .A(n1521), .B(n1520), .Z(n1548) );
  XOR U1828 ( .A(b[5]), .B(a[25]), .Z(n1561) );
  NAND U1829 ( .A(n1561), .B(n10481), .Z(n1524) );
  NAND U1830 ( .A(n1522), .B(n10482), .Z(n1523) );
  NAND U1831 ( .A(n1524), .B(n1523), .Z(n1546) );
  NANDN U1832 ( .A(n529), .B(a[21]), .Z(n1547) );
  XNOR U1833 ( .A(n1546), .B(n1547), .Z(n1549) );
  XOR U1834 ( .A(n1548), .B(n1549), .Z(n1543) );
  XOR U1835 ( .A(n1542), .B(n1543), .Z(n1564) );
  XOR U1836 ( .A(n1565), .B(n1564), .Z(n1566) );
  XNOR U1837 ( .A(n1567), .B(n1566), .Z(n1536) );
  NAND U1838 ( .A(n1526), .B(n1525), .Z(n1530) );
  NAND U1839 ( .A(n1528), .B(n1527), .Z(n1529) );
  NAND U1840 ( .A(n1530), .B(n1529), .Z(n1537) );
  XNOR U1841 ( .A(n1536), .B(n1537), .Z(n1538) );
  XNOR U1842 ( .A(n1539), .B(n1538), .Z(n1570) );
  XNOR U1843 ( .A(n1570), .B(sreg[277]), .Z(n1572) );
  NAND U1844 ( .A(n1531), .B(sreg[276]), .Z(n1535) );
  OR U1845 ( .A(n1533), .B(n1532), .Z(n1534) );
  AND U1846 ( .A(n1535), .B(n1534), .Z(n1571) );
  XOR U1847 ( .A(n1572), .B(n1571), .Z(c[277]) );
  NANDN U1848 ( .A(n1541), .B(n1540), .Z(n1545) );
  NAND U1849 ( .A(n1543), .B(n1542), .Z(n1544) );
  NAND U1850 ( .A(n1545), .B(n1544), .Z(n1606) );
  NANDN U1851 ( .A(n1547), .B(n1546), .Z(n1551) );
  NAND U1852 ( .A(n1549), .B(n1548), .Z(n1550) );
  NAND U1853 ( .A(n1551), .B(n1550), .Z(n1604) );
  XNOR U1854 ( .A(b[7]), .B(a[24]), .Z(n1591) );
  NANDN U1855 ( .A(n1591), .B(n10545), .Z(n1554) );
  NANDN U1856 ( .A(n1552), .B(n10546), .Z(n1553) );
  NAND U1857 ( .A(n1554), .B(n1553), .Z(n1579) );
  XNOR U1858 ( .A(b[3]), .B(a[28]), .Z(n1594) );
  NANDN U1859 ( .A(n1594), .B(n10398), .Z(n1557) );
  NANDN U1860 ( .A(n1555), .B(n10399), .Z(n1556) );
  AND U1861 ( .A(n1557), .B(n1556), .Z(n1580) );
  XNOR U1862 ( .A(n1579), .B(n1580), .Z(n1581) );
  NANDN U1863 ( .A(n527), .B(a[30]), .Z(n1558) );
  XOR U1864 ( .A(n10434), .B(n1558), .Z(n1560) );
  NANDN U1865 ( .A(b[0]), .B(a[29]), .Z(n1559) );
  AND U1866 ( .A(n1560), .B(n1559), .Z(n1587) );
  XOR U1867 ( .A(b[5]), .B(a[26]), .Z(n1600) );
  NAND U1868 ( .A(n1600), .B(n10481), .Z(n1563) );
  NAND U1869 ( .A(n1561), .B(n10482), .Z(n1562) );
  NAND U1870 ( .A(n1563), .B(n1562), .Z(n1585) );
  NANDN U1871 ( .A(n529), .B(a[22]), .Z(n1586) );
  XNOR U1872 ( .A(n1585), .B(n1586), .Z(n1588) );
  XOR U1873 ( .A(n1587), .B(n1588), .Z(n1582) );
  XOR U1874 ( .A(n1581), .B(n1582), .Z(n1603) );
  XOR U1875 ( .A(n1604), .B(n1603), .Z(n1605) );
  XNOR U1876 ( .A(n1606), .B(n1605), .Z(n1575) );
  NAND U1877 ( .A(n1565), .B(n1564), .Z(n1569) );
  NAND U1878 ( .A(n1567), .B(n1566), .Z(n1568) );
  NAND U1879 ( .A(n1569), .B(n1568), .Z(n1576) );
  XNOR U1880 ( .A(n1575), .B(n1576), .Z(n1577) );
  XNOR U1881 ( .A(n1578), .B(n1577), .Z(n1609) );
  XNOR U1882 ( .A(n1609), .B(sreg[278]), .Z(n1611) );
  NAND U1883 ( .A(n1570), .B(sreg[277]), .Z(n1574) );
  OR U1884 ( .A(n1572), .B(n1571), .Z(n1573) );
  AND U1885 ( .A(n1574), .B(n1573), .Z(n1610) );
  XOR U1886 ( .A(n1611), .B(n1610), .Z(c[278]) );
  NANDN U1887 ( .A(n1580), .B(n1579), .Z(n1584) );
  NAND U1888 ( .A(n1582), .B(n1581), .Z(n1583) );
  NAND U1889 ( .A(n1584), .B(n1583), .Z(n1645) );
  NANDN U1890 ( .A(n1586), .B(n1585), .Z(n1590) );
  NAND U1891 ( .A(n1588), .B(n1587), .Z(n1589) );
  NAND U1892 ( .A(n1590), .B(n1589), .Z(n1643) );
  XNOR U1893 ( .A(b[7]), .B(a[25]), .Z(n1618) );
  NANDN U1894 ( .A(n1618), .B(n10545), .Z(n1593) );
  NANDN U1895 ( .A(n1591), .B(n10546), .Z(n1592) );
  NAND U1896 ( .A(n1593), .B(n1592), .Z(n1630) );
  XNOR U1897 ( .A(b[3]), .B(a[29]), .Z(n1621) );
  NANDN U1898 ( .A(n1621), .B(n10398), .Z(n1596) );
  NANDN U1899 ( .A(n1594), .B(n10399), .Z(n1595) );
  AND U1900 ( .A(n1596), .B(n1595), .Z(n1631) );
  XNOR U1901 ( .A(n1630), .B(n1631), .Z(n1632) );
  NANDN U1902 ( .A(n527), .B(a[31]), .Z(n1597) );
  XOR U1903 ( .A(n10434), .B(n1597), .Z(n1599) );
  NANDN U1904 ( .A(b[0]), .B(a[30]), .Z(n1598) );
  AND U1905 ( .A(n1599), .B(n1598), .Z(n1638) );
  XOR U1906 ( .A(b[5]), .B(a[27]), .Z(n1627) );
  NAND U1907 ( .A(n10481), .B(n1627), .Z(n1602) );
  NAND U1908 ( .A(n10482), .B(n1600), .Z(n1601) );
  AND U1909 ( .A(n1602), .B(n1601), .Z(n1636) );
  NANDN U1910 ( .A(n529), .B(a[23]), .Z(n1637) );
  XOR U1911 ( .A(n1636), .B(n1637), .Z(n1639) );
  XNOR U1912 ( .A(n1638), .B(n1639), .Z(n1633) );
  XNOR U1913 ( .A(n1632), .B(n1633), .Z(n1642) );
  XOR U1914 ( .A(n1643), .B(n1642), .Z(n1644) );
  XNOR U1915 ( .A(n1645), .B(n1644), .Z(n1614) );
  NAND U1916 ( .A(n1604), .B(n1603), .Z(n1608) );
  NAND U1917 ( .A(n1606), .B(n1605), .Z(n1607) );
  NAND U1918 ( .A(n1608), .B(n1607), .Z(n1615) );
  XNOR U1919 ( .A(n1614), .B(n1615), .Z(n1616) );
  XNOR U1920 ( .A(n1617), .B(n1616), .Z(n1646) );
  XNOR U1921 ( .A(n1646), .B(sreg[279]), .Z(n1648) );
  NAND U1922 ( .A(n1609), .B(sreg[278]), .Z(n1613) );
  OR U1923 ( .A(n1611), .B(n1610), .Z(n1612) );
  AND U1924 ( .A(n1613), .B(n1612), .Z(n1647) );
  XOR U1925 ( .A(n1648), .B(n1647), .Z(c[279]) );
  XNOR U1926 ( .A(b[7]), .B(a[26]), .Z(n1673) );
  NANDN U1927 ( .A(n1673), .B(n10545), .Z(n1620) );
  NANDN U1928 ( .A(n1618), .B(n10546), .Z(n1619) );
  NAND U1929 ( .A(n1620), .B(n1619), .Z(n1655) );
  XNOR U1930 ( .A(b[3]), .B(a[30]), .Z(n1676) );
  NANDN U1931 ( .A(n1676), .B(n10398), .Z(n1623) );
  NANDN U1932 ( .A(n1621), .B(n10399), .Z(n1622) );
  AND U1933 ( .A(n1623), .B(n1622), .Z(n1656) );
  XNOR U1934 ( .A(n1655), .B(n1656), .Z(n1657) );
  NANDN U1935 ( .A(n527), .B(a[32]), .Z(n1624) );
  XOR U1936 ( .A(n10434), .B(n1624), .Z(n1626) );
  NANDN U1937 ( .A(b[0]), .B(a[31]), .Z(n1625) );
  AND U1938 ( .A(n1626), .B(n1625), .Z(n1663) );
  XOR U1939 ( .A(b[5]), .B(a[28]), .Z(n1670) );
  NAND U1940 ( .A(n1670), .B(n10481), .Z(n1629) );
  NAND U1941 ( .A(n1627), .B(n10482), .Z(n1628) );
  NAND U1942 ( .A(n1629), .B(n1628), .Z(n1661) );
  NANDN U1943 ( .A(n529), .B(a[24]), .Z(n1662) );
  XNOR U1944 ( .A(n1661), .B(n1662), .Z(n1664) );
  XOR U1945 ( .A(n1663), .B(n1664), .Z(n1658) );
  XOR U1946 ( .A(n1657), .B(n1658), .Z(n1681) );
  NANDN U1947 ( .A(n1631), .B(n1630), .Z(n1635) );
  NANDN U1948 ( .A(n1633), .B(n1632), .Z(n1634) );
  NAND U1949 ( .A(n1635), .B(n1634), .Z(n1679) );
  OR U1950 ( .A(n1637), .B(n1636), .Z(n1641) );
  NAND U1951 ( .A(n1639), .B(n1638), .Z(n1640) );
  AND U1952 ( .A(n1641), .B(n1640), .Z(n1680) );
  XNOR U1953 ( .A(n1679), .B(n1680), .Z(n1682) );
  XNOR U1954 ( .A(n1681), .B(n1682), .Z(n1651) );
  XNOR U1955 ( .A(n1651), .B(n1652), .Z(n1653) );
  XNOR U1956 ( .A(n1654), .B(n1653), .Z(n1685) );
  XNOR U1957 ( .A(n1685), .B(sreg[280]), .Z(n1687) );
  NAND U1958 ( .A(n1646), .B(sreg[279]), .Z(n1650) );
  OR U1959 ( .A(n1648), .B(n1647), .Z(n1649) );
  AND U1960 ( .A(n1650), .B(n1649), .Z(n1686) );
  XOR U1961 ( .A(n1687), .B(n1686), .Z(c[280]) );
  NANDN U1962 ( .A(n1656), .B(n1655), .Z(n1660) );
  NAND U1963 ( .A(n1658), .B(n1657), .Z(n1659) );
  NAND U1964 ( .A(n1660), .B(n1659), .Z(n1721) );
  NANDN U1965 ( .A(n1662), .B(n1661), .Z(n1666) );
  NAND U1966 ( .A(n1664), .B(n1663), .Z(n1665) );
  NAND U1967 ( .A(n1666), .B(n1665), .Z(n1719) );
  NANDN U1968 ( .A(n527), .B(a[33]), .Z(n1667) );
  XOR U1969 ( .A(n10434), .B(n1667), .Z(n1669) );
  NANDN U1970 ( .A(b[0]), .B(a[32]), .Z(n1668) );
  AND U1971 ( .A(n1669), .B(n1668), .Z(n1702) );
  XOR U1972 ( .A(b[5]), .B(a[29]), .Z(n1715) );
  NAND U1973 ( .A(n1715), .B(n10481), .Z(n1672) );
  NAND U1974 ( .A(n1670), .B(n10482), .Z(n1671) );
  NAND U1975 ( .A(n1672), .B(n1671), .Z(n1700) );
  NANDN U1976 ( .A(n529), .B(a[25]), .Z(n1701) );
  XNOR U1977 ( .A(n1700), .B(n1701), .Z(n1703) );
  XOR U1978 ( .A(n1702), .B(n1703), .Z(n1696) );
  XNOR U1979 ( .A(b[7]), .B(a[27]), .Z(n1706) );
  NANDN U1980 ( .A(n1706), .B(n10545), .Z(n1675) );
  NANDN U1981 ( .A(n1673), .B(n10546), .Z(n1674) );
  NAND U1982 ( .A(n1675), .B(n1674), .Z(n1694) );
  XNOR U1983 ( .A(b[3]), .B(a[31]), .Z(n1709) );
  NANDN U1984 ( .A(n1709), .B(n10398), .Z(n1678) );
  NANDN U1985 ( .A(n1676), .B(n10399), .Z(n1677) );
  AND U1986 ( .A(n1678), .B(n1677), .Z(n1695) );
  XNOR U1987 ( .A(n1694), .B(n1695), .Z(n1697) );
  XOR U1988 ( .A(n1696), .B(n1697), .Z(n1718) );
  XOR U1989 ( .A(n1719), .B(n1718), .Z(n1720) );
  XNOR U1990 ( .A(n1721), .B(n1720), .Z(n1690) );
  NANDN U1991 ( .A(n1680), .B(n1679), .Z(n1684) );
  NAND U1992 ( .A(n1682), .B(n1681), .Z(n1683) );
  NAND U1993 ( .A(n1684), .B(n1683), .Z(n1691) );
  XNOR U1994 ( .A(n1690), .B(n1691), .Z(n1692) );
  XNOR U1995 ( .A(n1693), .B(n1692), .Z(n1724) );
  XNOR U1996 ( .A(n1724), .B(sreg[281]), .Z(n1726) );
  NAND U1997 ( .A(n1685), .B(sreg[280]), .Z(n1689) );
  OR U1998 ( .A(n1687), .B(n1686), .Z(n1688) );
  AND U1999 ( .A(n1689), .B(n1688), .Z(n1725) );
  XOR U2000 ( .A(n1726), .B(n1725), .Z(c[281]) );
  NANDN U2001 ( .A(n1695), .B(n1694), .Z(n1699) );
  NAND U2002 ( .A(n1697), .B(n1696), .Z(n1698) );
  NAND U2003 ( .A(n1699), .B(n1698), .Z(n1760) );
  NANDN U2004 ( .A(n1701), .B(n1700), .Z(n1705) );
  NAND U2005 ( .A(n1703), .B(n1702), .Z(n1704) );
  NAND U2006 ( .A(n1705), .B(n1704), .Z(n1758) );
  XNOR U2007 ( .A(b[7]), .B(a[28]), .Z(n1745) );
  NANDN U2008 ( .A(n1745), .B(n10545), .Z(n1708) );
  NANDN U2009 ( .A(n1706), .B(n10546), .Z(n1707) );
  NAND U2010 ( .A(n1708), .B(n1707), .Z(n1733) );
  XNOR U2011 ( .A(b[3]), .B(a[32]), .Z(n1748) );
  NANDN U2012 ( .A(n1748), .B(n10398), .Z(n1711) );
  NANDN U2013 ( .A(n1709), .B(n10399), .Z(n1710) );
  AND U2014 ( .A(n1711), .B(n1710), .Z(n1734) );
  XNOR U2015 ( .A(n1733), .B(n1734), .Z(n1735) );
  NANDN U2016 ( .A(n527), .B(a[34]), .Z(n1712) );
  XOR U2017 ( .A(n10434), .B(n1712), .Z(n1714) );
  NANDN U2018 ( .A(b[0]), .B(a[33]), .Z(n1713) );
  AND U2019 ( .A(n1714), .B(n1713), .Z(n1741) );
  XOR U2020 ( .A(b[5]), .B(a[30]), .Z(n1754) );
  NAND U2021 ( .A(n1754), .B(n10481), .Z(n1717) );
  NAND U2022 ( .A(n1715), .B(n10482), .Z(n1716) );
  NAND U2023 ( .A(n1717), .B(n1716), .Z(n1739) );
  NANDN U2024 ( .A(n529), .B(a[26]), .Z(n1740) );
  XNOR U2025 ( .A(n1739), .B(n1740), .Z(n1742) );
  XOR U2026 ( .A(n1741), .B(n1742), .Z(n1736) );
  XOR U2027 ( .A(n1735), .B(n1736), .Z(n1757) );
  XOR U2028 ( .A(n1758), .B(n1757), .Z(n1759) );
  XNOR U2029 ( .A(n1760), .B(n1759), .Z(n1729) );
  NAND U2030 ( .A(n1719), .B(n1718), .Z(n1723) );
  NAND U2031 ( .A(n1721), .B(n1720), .Z(n1722) );
  NAND U2032 ( .A(n1723), .B(n1722), .Z(n1730) );
  XNOR U2033 ( .A(n1729), .B(n1730), .Z(n1731) );
  XNOR U2034 ( .A(n1732), .B(n1731), .Z(n1763) );
  XNOR U2035 ( .A(n1763), .B(sreg[282]), .Z(n1765) );
  NAND U2036 ( .A(n1724), .B(sreg[281]), .Z(n1728) );
  OR U2037 ( .A(n1726), .B(n1725), .Z(n1727) );
  AND U2038 ( .A(n1728), .B(n1727), .Z(n1764) );
  XOR U2039 ( .A(n1765), .B(n1764), .Z(c[282]) );
  NANDN U2040 ( .A(n1734), .B(n1733), .Z(n1738) );
  NAND U2041 ( .A(n1736), .B(n1735), .Z(n1737) );
  NAND U2042 ( .A(n1738), .B(n1737), .Z(n1799) );
  NANDN U2043 ( .A(n1740), .B(n1739), .Z(n1744) );
  NAND U2044 ( .A(n1742), .B(n1741), .Z(n1743) );
  NAND U2045 ( .A(n1744), .B(n1743), .Z(n1797) );
  XNOR U2046 ( .A(b[7]), .B(a[29]), .Z(n1784) );
  NANDN U2047 ( .A(n1784), .B(n10545), .Z(n1747) );
  NANDN U2048 ( .A(n1745), .B(n10546), .Z(n1746) );
  NAND U2049 ( .A(n1747), .B(n1746), .Z(n1772) );
  XNOR U2050 ( .A(b[3]), .B(a[33]), .Z(n1787) );
  NANDN U2051 ( .A(n1787), .B(n10398), .Z(n1750) );
  NANDN U2052 ( .A(n1748), .B(n10399), .Z(n1749) );
  AND U2053 ( .A(n1750), .B(n1749), .Z(n1773) );
  XNOR U2054 ( .A(n1772), .B(n1773), .Z(n1774) );
  NANDN U2055 ( .A(n527), .B(a[35]), .Z(n1751) );
  XOR U2056 ( .A(n10434), .B(n1751), .Z(n1753) );
  NANDN U2057 ( .A(b[0]), .B(a[34]), .Z(n1752) );
  AND U2058 ( .A(n1753), .B(n1752), .Z(n1780) );
  XOR U2059 ( .A(b[5]), .B(a[31]), .Z(n1793) );
  NAND U2060 ( .A(n1793), .B(n10481), .Z(n1756) );
  NAND U2061 ( .A(n1754), .B(n10482), .Z(n1755) );
  NAND U2062 ( .A(n1756), .B(n1755), .Z(n1778) );
  NANDN U2063 ( .A(n529), .B(a[27]), .Z(n1779) );
  XNOR U2064 ( .A(n1778), .B(n1779), .Z(n1781) );
  XOR U2065 ( .A(n1780), .B(n1781), .Z(n1775) );
  XOR U2066 ( .A(n1774), .B(n1775), .Z(n1796) );
  XOR U2067 ( .A(n1797), .B(n1796), .Z(n1798) );
  XNOR U2068 ( .A(n1799), .B(n1798), .Z(n1768) );
  NAND U2069 ( .A(n1758), .B(n1757), .Z(n1762) );
  NAND U2070 ( .A(n1760), .B(n1759), .Z(n1761) );
  NAND U2071 ( .A(n1762), .B(n1761), .Z(n1769) );
  XNOR U2072 ( .A(n1768), .B(n1769), .Z(n1770) );
  XNOR U2073 ( .A(n1771), .B(n1770), .Z(n1802) );
  XNOR U2074 ( .A(n1802), .B(sreg[283]), .Z(n1804) );
  NAND U2075 ( .A(n1763), .B(sreg[282]), .Z(n1767) );
  OR U2076 ( .A(n1765), .B(n1764), .Z(n1766) );
  AND U2077 ( .A(n1767), .B(n1766), .Z(n1803) );
  XOR U2078 ( .A(n1804), .B(n1803), .Z(c[283]) );
  NANDN U2079 ( .A(n1773), .B(n1772), .Z(n1777) );
  NAND U2080 ( .A(n1775), .B(n1774), .Z(n1776) );
  NAND U2081 ( .A(n1777), .B(n1776), .Z(n1838) );
  NANDN U2082 ( .A(n1779), .B(n1778), .Z(n1783) );
  NAND U2083 ( .A(n1781), .B(n1780), .Z(n1782) );
  NAND U2084 ( .A(n1783), .B(n1782), .Z(n1836) );
  XNOR U2085 ( .A(b[7]), .B(a[30]), .Z(n1823) );
  NANDN U2086 ( .A(n1823), .B(n10545), .Z(n1786) );
  NANDN U2087 ( .A(n1784), .B(n10546), .Z(n1785) );
  NAND U2088 ( .A(n1786), .B(n1785), .Z(n1811) );
  XNOR U2089 ( .A(b[3]), .B(a[34]), .Z(n1826) );
  NANDN U2090 ( .A(n1826), .B(n10398), .Z(n1789) );
  NANDN U2091 ( .A(n1787), .B(n10399), .Z(n1788) );
  AND U2092 ( .A(n1789), .B(n1788), .Z(n1812) );
  XNOR U2093 ( .A(n1811), .B(n1812), .Z(n1813) );
  NANDN U2094 ( .A(n527), .B(a[36]), .Z(n1790) );
  XOR U2095 ( .A(n10434), .B(n1790), .Z(n1792) );
  NANDN U2096 ( .A(b[0]), .B(a[35]), .Z(n1791) );
  AND U2097 ( .A(n1792), .B(n1791), .Z(n1819) );
  XOR U2098 ( .A(b[5]), .B(a[32]), .Z(n1832) );
  NAND U2099 ( .A(n1832), .B(n10481), .Z(n1795) );
  NAND U2100 ( .A(n1793), .B(n10482), .Z(n1794) );
  NAND U2101 ( .A(n1795), .B(n1794), .Z(n1817) );
  NANDN U2102 ( .A(n529), .B(a[28]), .Z(n1818) );
  XNOR U2103 ( .A(n1817), .B(n1818), .Z(n1820) );
  XOR U2104 ( .A(n1819), .B(n1820), .Z(n1814) );
  XOR U2105 ( .A(n1813), .B(n1814), .Z(n1835) );
  XOR U2106 ( .A(n1836), .B(n1835), .Z(n1837) );
  XNOR U2107 ( .A(n1838), .B(n1837), .Z(n1807) );
  NAND U2108 ( .A(n1797), .B(n1796), .Z(n1801) );
  NAND U2109 ( .A(n1799), .B(n1798), .Z(n1800) );
  NAND U2110 ( .A(n1801), .B(n1800), .Z(n1808) );
  XNOR U2111 ( .A(n1807), .B(n1808), .Z(n1809) );
  XNOR U2112 ( .A(n1810), .B(n1809), .Z(n1841) );
  XNOR U2113 ( .A(n1841), .B(sreg[284]), .Z(n1843) );
  NAND U2114 ( .A(n1802), .B(sreg[283]), .Z(n1806) );
  OR U2115 ( .A(n1804), .B(n1803), .Z(n1805) );
  AND U2116 ( .A(n1806), .B(n1805), .Z(n1842) );
  XOR U2117 ( .A(n1843), .B(n1842), .Z(c[284]) );
  NANDN U2118 ( .A(n1812), .B(n1811), .Z(n1816) );
  NAND U2119 ( .A(n1814), .B(n1813), .Z(n1815) );
  NAND U2120 ( .A(n1816), .B(n1815), .Z(n1877) );
  NANDN U2121 ( .A(n1818), .B(n1817), .Z(n1822) );
  NAND U2122 ( .A(n1820), .B(n1819), .Z(n1821) );
  NAND U2123 ( .A(n1822), .B(n1821), .Z(n1875) );
  XNOR U2124 ( .A(b[7]), .B(a[31]), .Z(n1862) );
  NANDN U2125 ( .A(n1862), .B(n10545), .Z(n1825) );
  NANDN U2126 ( .A(n1823), .B(n10546), .Z(n1824) );
  NAND U2127 ( .A(n1825), .B(n1824), .Z(n1850) );
  XNOR U2128 ( .A(b[3]), .B(a[35]), .Z(n1865) );
  NANDN U2129 ( .A(n1865), .B(n10398), .Z(n1828) );
  NANDN U2130 ( .A(n1826), .B(n10399), .Z(n1827) );
  AND U2131 ( .A(n1828), .B(n1827), .Z(n1851) );
  XNOR U2132 ( .A(n1850), .B(n1851), .Z(n1852) );
  NANDN U2133 ( .A(n527), .B(a[37]), .Z(n1829) );
  XOR U2134 ( .A(n10434), .B(n1829), .Z(n1831) );
  NANDN U2135 ( .A(b[0]), .B(a[36]), .Z(n1830) );
  AND U2136 ( .A(n1831), .B(n1830), .Z(n1858) );
  XOR U2137 ( .A(b[5]), .B(a[33]), .Z(n1871) );
  NAND U2138 ( .A(n1871), .B(n10481), .Z(n1834) );
  NAND U2139 ( .A(n1832), .B(n10482), .Z(n1833) );
  NAND U2140 ( .A(n1834), .B(n1833), .Z(n1856) );
  NANDN U2141 ( .A(n529), .B(a[29]), .Z(n1857) );
  XNOR U2142 ( .A(n1856), .B(n1857), .Z(n1859) );
  XOR U2143 ( .A(n1858), .B(n1859), .Z(n1853) );
  XOR U2144 ( .A(n1852), .B(n1853), .Z(n1874) );
  XOR U2145 ( .A(n1875), .B(n1874), .Z(n1876) );
  XNOR U2146 ( .A(n1877), .B(n1876), .Z(n1846) );
  NAND U2147 ( .A(n1836), .B(n1835), .Z(n1840) );
  NAND U2148 ( .A(n1838), .B(n1837), .Z(n1839) );
  NAND U2149 ( .A(n1840), .B(n1839), .Z(n1847) );
  XNOR U2150 ( .A(n1846), .B(n1847), .Z(n1848) );
  XNOR U2151 ( .A(n1849), .B(n1848), .Z(n1880) );
  XNOR U2152 ( .A(n1880), .B(sreg[285]), .Z(n1882) );
  NAND U2153 ( .A(n1841), .B(sreg[284]), .Z(n1845) );
  OR U2154 ( .A(n1843), .B(n1842), .Z(n1844) );
  AND U2155 ( .A(n1845), .B(n1844), .Z(n1881) );
  XOR U2156 ( .A(n1882), .B(n1881), .Z(c[285]) );
  NANDN U2157 ( .A(n1851), .B(n1850), .Z(n1855) );
  NAND U2158 ( .A(n1853), .B(n1852), .Z(n1854) );
  NAND U2159 ( .A(n1855), .B(n1854), .Z(n1916) );
  NANDN U2160 ( .A(n1857), .B(n1856), .Z(n1861) );
  NAND U2161 ( .A(n1859), .B(n1858), .Z(n1860) );
  NAND U2162 ( .A(n1861), .B(n1860), .Z(n1914) );
  XNOR U2163 ( .A(b[7]), .B(a[32]), .Z(n1907) );
  NANDN U2164 ( .A(n1907), .B(n10545), .Z(n1864) );
  NANDN U2165 ( .A(n1862), .B(n10546), .Z(n1863) );
  NAND U2166 ( .A(n1864), .B(n1863), .Z(n1889) );
  XNOR U2167 ( .A(b[3]), .B(a[36]), .Z(n1910) );
  NANDN U2168 ( .A(n1910), .B(n10398), .Z(n1867) );
  NANDN U2169 ( .A(n1865), .B(n10399), .Z(n1866) );
  AND U2170 ( .A(n1867), .B(n1866), .Z(n1890) );
  XNOR U2171 ( .A(n1889), .B(n1890), .Z(n1891) );
  NANDN U2172 ( .A(n527), .B(a[38]), .Z(n1868) );
  XOR U2173 ( .A(n10434), .B(n1868), .Z(n1870) );
  NANDN U2174 ( .A(b[0]), .B(a[37]), .Z(n1869) );
  AND U2175 ( .A(n1870), .B(n1869), .Z(n1897) );
  XOR U2176 ( .A(b[5]), .B(a[34]), .Z(n1904) );
  NAND U2177 ( .A(n1904), .B(n10481), .Z(n1873) );
  NAND U2178 ( .A(n1871), .B(n10482), .Z(n1872) );
  NAND U2179 ( .A(n1873), .B(n1872), .Z(n1895) );
  NANDN U2180 ( .A(n529), .B(a[30]), .Z(n1896) );
  XNOR U2181 ( .A(n1895), .B(n1896), .Z(n1898) );
  XOR U2182 ( .A(n1897), .B(n1898), .Z(n1892) );
  XOR U2183 ( .A(n1891), .B(n1892), .Z(n1913) );
  XOR U2184 ( .A(n1914), .B(n1913), .Z(n1915) );
  XNOR U2185 ( .A(n1916), .B(n1915), .Z(n1885) );
  NAND U2186 ( .A(n1875), .B(n1874), .Z(n1879) );
  NAND U2187 ( .A(n1877), .B(n1876), .Z(n1878) );
  NAND U2188 ( .A(n1879), .B(n1878), .Z(n1886) );
  XNOR U2189 ( .A(n1885), .B(n1886), .Z(n1887) );
  XNOR U2190 ( .A(n1888), .B(n1887), .Z(n1919) );
  XNOR U2191 ( .A(n1919), .B(sreg[286]), .Z(n1921) );
  NAND U2192 ( .A(n1880), .B(sreg[285]), .Z(n1884) );
  OR U2193 ( .A(n1882), .B(n1881), .Z(n1883) );
  AND U2194 ( .A(n1884), .B(n1883), .Z(n1920) );
  XOR U2195 ( .A(n1921), .B(n1920), .Z(c[286]) );
  NANDN U2196 ( .A(n1890), .B(n1889), .Z(n1894) );
  NAND U2197 ( .A(n1892), .B(n1891), .Z(n1893) );
  NAND U2198 ( .A(n1894), .B(n1893), .Z(n1955) );
  NANDN U2199 ( .A(n1896), .B(n1895), .Z(n1900) );
  NAND U2200 ( .A(n1898), .B(n1897), .Z(n1899) );
  NAND U2201 ( .A(n1900), .B(n1899), .Z(n1953) );
  NANDN U2202 ( .A(n527), .B(a[39]), .Z(n1901) );
  XOR U2203 ( .A(n10434), .B(n1901), .Z(n1903) );
  NANDN U2204 ( .A(b[0]), .B(a[38]), .Z(n1902) );
  AND U2205 ( .A(n1903), .B(n1902), .Z(n1936) );
  XOR U2206 ( .A(b[5]), .B(a[35]), .Z(n1949) );
  NAND U2207 ( .A(n1949), .B(n10481), .Z(n1906) );
  NAND U2208 ( .A(n1904), .B(n10482), .Z(n1905) );
  NAND U2209 ( .A(n1906), .B(n1905), .Z(n1934) );
  NANDN U2210 ( .A(n529), .B(a[31]), .Z(n1935) );
  XNOR U2211 ( .A(n1934), .B(n1935), .Z(n1937) );
  XOR U2212 ( .A(n1936), .B(n1937), .Z(n1930) );
  XNOR U2213 ( .A(b[7]), .B(a[33]), .Z(n1940) );
  NANDN U2214 ( .A(n1940), .B(n10545), .Z(n1909) );
  NANDN U2215 ( .A(n1907), .B(n10546), .Z(n1908) );
  NAND U2216 ( .A(n1909), .B(n1908), .Z(n1928) );
  XNOR U2217 ( .A(b[3]), .B(a[37]), .Z(n1943) );
  NANDN U2218 ( .A(n1943), .B(n10398), .Z(n1912) );
  NANDN U2219 ( .A(n1910), .B(n10399), .Z(n1911) );
  AND U2220 ( .A(n1912), .B(n1911), .Z(n1929) );
  XNOR U2221 ( .A(n1928), .B(n1929), .Z(n1931) );
  XOR U2222 ( .A(n1930), .B(n1931), .Z(n1952) );
  XOR U2223 ( .A(n1953), .B(n1952), .Z(n1954) );
  XNOR U2224 ( .A(n1955), .B(n1954), .Z(n1924) );
  NAND U2225 ( .A(n1914), .B(n1913), .Z(n1918) );
  NAND U2226 ( .A(n1916), .B(n1915), .Z(n1917) );
  NAND U2227 ( .A(n1918), .B(n1917), .Z(n1925) );
  XNOR U2228 ( .A(n1924), .B(n1925), .Z(n1926) );
  XNOR U2229 ( .A(n1927), .B(n1926), .Z(n1958) );
  XNOR U2230 ( .A(n1958), .B(sreg[287]), .Z(n1960) );
  NAND U2231 ( .A(n1919), .B(sreg[286]), .Z(n1923) );
  OR U2232 ( .A(n1921), .B(n1920), .Z(n1922) );
  AND U2233 ( .A(n1923), .B(n1922), .Z(n1959) );
  XOR U2234 ( .A(n1960), .B(n1959), .Z(c[287]) );
  NANDN U2235 ( .A(n1929), .B(n1928), .Z(n1933) );
  NAND U2236 ( .A(n1931), .B(n1930), .Z(n1932) );
  NAND U2237 ( .A(n1933), .B(n1932), .Z(n1994) );
  NANDN U2238 ( .A(n1935), .B(n1934), .Z(n1939) );
  NAND U2239 ( .A(n1937), .B(n1936), .Z(n1938) );
  NAND U2240 ( .A(n1939), .B(n1938), .Z(n1992) );
  XNOR U2241 ( .A(b[7]), .B(a[34]), .Z(n1979) );
  NANDN U2242 ( .A(n1979), .B(n10545), .Z(n1942) );
  NANDN U2243 ( .A(n1940), .B(n10546), .Z(n1941) );
  NAND U2244 ( .A(n1942), .B(n1941), .Z(n1967) );
  XNOR U2245 ( .A(b[3]), .B(a[38]), .Z(n1982) );
  NANDN U2246 ( .A(n1982), .B(n10398), .Z(n1945) );
  NANDN U2247 ( .A(n1943), .B(n10399), .Z(n1944) );
  AND U2248 ( .A(n1945), .B(n1944), .Z(n1968) );
  XNOR U2249 ( .A(n1967), .B(n1968), .Z(n1969) );
  NANDN U2250 ( .A(n527), .B(a[40]), .Z(n1946) );
  XOR U2251 ( .A(n10434), .B(n1946), .Z(n1948) );
  NANDN U2252 ( .A(b[0]), .B(a[39]), .Z(n1947) );
  AND U2253 ( .A(n1948), .B(n1947), .Z(n1975) );
  XOR U2254 ( .A(b[5]), .B(a[36]), .Z(n1988) );
  NAND U2255 ( .A(n1988), .B(n10481), .Z(n1951) );
  NAND U2256 ( .A(n1949), .B(n10482), .Z(n1950) );
  NAND U2257 ( .A(n1951), .B(n1950), .Z(n1973) );
  NANDN U2258 ( .A(n529), .B(a[32]), .Z(n1974) );
  XNOR U2259 ( .A(n1973), .B(n1974), .Z(n1976) );
  XOR U2260 ( .A(n1975), .B(n1976), .Z(n1970) );
  XOR U2261 ( .A(n1969), .B(n1970), .Z(n1991) );
  XOR U2262 ( .A(n1992), .B(n1991), .Z(n1993) );
  XNOR U2263 ( .A(n1994), .B(n1993), .Z(n1963) );
  NAND U2264 ( .A(n1953), .B(n1952), .Z(n1957) );
  NAND U2265 ( .A(n1955), .B(n1954), .Z(n1956) );
  NAND U2266 ( .A(n1957), .B(n1956), .Z(n1964) );
  XNOR U2267 ( .A(n1963), .B(n1964), .Z(n1965) );
  XNOR U2268 ( .A(n1966), .B(n1965), .Z(n1997) );
  XNOR U2269 ( .A(n1997), .B(sreg[288]), .Z(n1999) );
  NAND U2270 ( .A(n1958), .B(sreg[287]), .Z(n1962) );
  OR U2271 ( .A(n1960), .B(n1959), .Z(n1961) );
  AND U2272 ( .A(n1962), .B(n1961), .Z(n1998) );
  XOR U2273 ( .A(n1999), .B(n1998), .Z(c[288]) );
  NANDN U2274 ( .A(n1968), .B(n1967), .Z(n1972) );
  NAND U2275 ( .A(n1970), .B(n1969), .Z(n1971) );
  NAND U2276 ( .A(n1972), .B(n1971), .Z(n2033) );
  NANDN U2277 ( .A(n1974), .B(n1973), .Z(n1978) );
  NAND U2278 ( .A(n1976), .B(n1975), .Z(n1977) );
  NAND U2279 ( .A(n1978), .B(n1977), .Z(n2031) );
  XNOR U2280 ( .A(b[7]), .B(a[35]), .Z(n2018) );
  NANDN U2281 ( .A(n2018), .B(n10545), .Z(n1981) );
  NANDN U2282 ( .A(n1979), .B(n10546), .Z(n1980) );
  NAND U2283 ( .A(n1981), .B(n1980), .Z(n2006) );
  XNOR U2284 ( .A(b[3]), .B(a[39]), .Z(n2021) );
  NANDN U2285 ( .A(n2021), .B(n10398), .Z(n1984) );
  NANDN U2286 ( .A(n1982), .B(n10399), .Z(n1983) );
  AND U2287 ( .A(n1984), .B(n1983), .Z(n2007) );
  XNOR U2288 ( .A(n2006), .B(n2007), .Z(n2008) );
  NANDN U2289 ( .A(n527), .B(a[41]), .Z(n1985) );
  XOR U2290 ( .A(n10434), .B(n1985), .Z(n1987) );
  NANDN U2291 ( .A(b[0]), .B(a[40]), .Z(n1986) );
  AND U2292 ( .A(n1987), .B(n1986), .Z(n2014) );
  XOR U2293 ( .A(b[5]), .B(a[37]), .Z(n2027) );
  NAND U2294 ( .A(n2027), .B(n10481), .Z(n1990) );
  NAND U2295 ( .A(n1988), .B(n10482), .Z(n1989) );
  NAND U2296 ( .A(n1990), .B(n1989), .Z(n2012) );
  NANDN U2297 ( .A(n529), .B(a[33]), .Z(n2013) );
  XNOR U2298 ( .A(n2012), .B(n2013), .Z(n2015) );
  XOR U2299 ( .A(n2014), .B(n2015), .Z(n2009) );
  XOR U2300 ( .A(n2008), .B(n2009), .Z(n2030) );
  XOR U2301 ( .A(n2031), .B(n2030), .Z(n2032) );
  XNOR U2302 ( .A(n2033), .B(n2032), .Z(n2002) );
  NAND U2303 ( .A(n1992), .B(n1991), .Z(n1996) );
  NAND U2304 ( .A(n1994), .B(n1993), .Z(n1995) );
  NAND U2305 ( .A(n1996), .B(n1995), .Z(n2003) );
  XNOR U2306 ( .A(n2002), .B(n2003), .Z(n2004) );
  XNOR U2307 ( .A(n2005), .B(n2004), .Z(n2036) );
  XNOR U2308 ( .A(n2036), .B(sreg[289]), .Z(n2038) );
  NAND U2309 ( .A(n1997), .B(sreg[288]), .Z(n2001) );
  OR U2310 ( .A(n1999), .B(n1998), .Z(n2000) );
  AND U2311 ( .A(n2001), .B(n2000), .Z(n2037) );
  XOR U2312 ( .A(n2038), .B(n2037), .Z(c[289]) );
  NANDN U2313 ( .A(n2007), .B(n2006), .Z(n2011) );
  NAND U2314 ( .A(n2009), .B(n2008), .Z(n2010) );
  NAND U2315 ( .A(n2011), .B(n2010), .Z(n2072) );
  NANDN U2316 ( .A(n2013), .B(n2012), .Z(n2017) );
  NAND U2317 ( .A(n2015), .B(n2014), .Z(n2016) );
  NAND U2318 ( .A(n2017), .B(n2016), .Z(n2070) );
  XNOR U2319 ( .A(b[7]), .B(a[36]), .Z(n2057) );
  NANDN U2320 ( .A(n2057), .B(n10545), .Z(n2020) );
  NANDN U2321 ( .A(n2018), .B(n10546), .Z(n2019) );
  NAND U2322 ( .A(n2020), .B(n2019), .Z(n2045) );
  XNOR U2323 ( .A(b[3]), .B(a[40]), .Z(n2060) );
  NANDN U2324 ( .A(n2060), .B(n10398), .Z(n2023) );
  NANDN U2325 ( .A(n2021), .B(n10399), .Z(n2022) );
  AND U2326 ( .A(n2023), .B(n2022), .Z(n2046) );
  XNOR U2327 ( .A(n2045), .B(n2046), .Z(n2047) );
  NANDN U2328 ( .A(n527), .B(a[42]), .Z(n2024) );
  XOR U2329 ( .A(n10434), .B(n2024), .Z(n2026) );
  NANDN U2330 ( .A(b[0]), .B(a[41]), .Z(n2025) );
  AND U2331 ( .A(n2026), .B(n2025), .Z(n2053) );
  XOR U2332 ( .A(b[5]), .B(a[38]), .Z(n2066) );
  NAND U2333 ( .A(n2066), .B(n10481), .Z(n2029) );
  NAND U2334 ( .A(n2027), .B(n10482), .Z(n2028) );
  NAND U2335 ( .A(n2029), .B(n2028), .Z(n2051) );
  NANDN U2336 ( .A(n529), .B(a[34]), .Z(n2052) );
  XNOR U2337 ( .A(n2051), .B(n2052), .Z(n2054) );
  XOR U2338 ( .A(n2053), .B(n2054), .Z(n2048) );
  XOR U2339 ( .A(n2047), .B(n2048), .Z(n2069) );
  XOR U2340 ( .A(n2070), .B(n2069), .Z(n2071) );
  XNOR U2341 ( .A(n2072), .B(n2071), .Z(n2041) );
  NAND U2342 ( .A(n2031), .B(n2030), .Z(n2035) );
  NAND U2343 ( .A(n2033), .B(n2032), .Z(n2034) );
  NAND U2344 ( .A(n2035), .B(n2034), .Z(n2042) );
  XNOR U2345 ( .A(n2041), .B(n2042), .Z(n2043) );
  XNOR U2346 ( .A(n2044), .B(n2043), .Z(n2075) );
  XNOR U2347 ( .A(n2075), .B(sreg[290]), .Z(n2077) );
  NAND U2348 ( .A(n2036), .B(sreg[289]), .Z(n2040) );
  OR U2349 ( .A(n2038), .B(n2037), .Z(n2039) );
  AND U2350 ( .A(n2040), .B(n2039), .Z(n2076) );
  XOR U2351 ( .A(n2077), .B(n2076), .Z(c[290]) );
  NANDN U2352 ( .A(n2046), .B(n2045), .Z(n2050) );
  NAND U2353 ( .A(n2048), .B(n2047), .Z(n2049) );
  NAND U2354 ( .A(n2050), .B(n2049), .Z(n2111) );
  NANDN U2355 ( .A(n2052), .B(n2051), .Z(n2056) );
  NAND U2356 ( .A(n2054), .B(n2053), .Z(n2055) );
  NAND U2357 ( .A(n2056), .B(n2055), .Z(n2109) );
  XNOR U2358 ( .A(b[7]), .B(a[37]), .Z(n2096) );
  NANDN U2359 ( .A(n2096), .B(n10545), .Z(n2059) );
  NANDN U2360 ( .A(n2057), .B(n10546), .Z(n2058) );
  NAND U2361 ( .A(n2059), .B(n2058), .Z(n2084) );
  XNOR U2362 ( .A(b[3]), .B(a[41]), .Z(n2099) );
  NANDN U2363 ( .A(n2099), .B(n10398), .Z(n2062) );
  NANDN U2364 ( .A(n2060), .B(n10399), .Z(n2061) );
  AND U2365 ( .A(n2062), .B(n2061), .Z(n2085) );
  XNOR U2366 ( .A(n2084), .B(n2085), .Z(n2086) );
  NANDN U2367 ( .A(n527), .B(a[43]), .Z(n2063) );
  XOR U2368 ( .A(n10434), .B(n2063), .Z(n2065) );
  NANDN U2369 ( .A(b[0]), .B(a[42]), .Z(n2064) );
  AND U2370 ( .A(n2065), .B(n2064), .Z(n2092) );
  XOR U2371 ( .A(b[5]), .B(a[39]), .Z(n2105) );
  NAND U2372 ( .A(n2105), .B(n10481), .Z(n2068) );
  NAND U2373 ( .A(n2066), .B(n10482), .Z(n2067) );
  NAND U2374 ( .A(n2068), .B(n2067), .Z(n2090) );
  NANDN U2375 ( .A(n529), .B(a[35]), .Z(n2091) );
  XNOR U2376 ( .A(n2090), .B(n2091), .Z(n2093) );
  XOR U2377 ( .A(n2092), .B(n2093), .Z(n2087) );
  XOR U2378 ( .A(n2086), .B(n2087), .Z(n2108) );
  XOR U2379 ( .A(n2109), .B(n2108), .Z(n2110) );
  XNOR U2380 ( .A(n2111), .B(n2110), .Z(n2080) );
  NAND U2381 ( .A(n2070), .B(n2069), .Z(n2074) );
  NAND U2382 ( .A(n2072), .B(n2071), .Z(n2073) );
  NAND U2383 ( .A(n2074), .B(n2073), .Z(n2081) );
  XNOR U2384 ( .A(n2080), .B(n2081), .Z(n2082) );
  XNOR U2385 ( .A(n2083), .B(n2082), .Z(n2114) );
  XNOR U2386 ( .A(n2114), .B(sreg[291]), .Z(n2116) );
  NAND U2387 ( .A(n2075), .B(sreg[290]), .Z(n2079) );
  OR U2388 ( .A(n2077), .B(n2076), .Z(n2078) );
  AND U2389 ( .A(n2079), .B(n2078), .Z(n2115) );
  XOR U2390 ( .A(n2116), .B(n2115), .Z(c[291]) );
  NANDN U2391 ( .A(n2085), .B(n2084), .Z(n2089) );
  NAND U2392 ( .A(n2087), .B(n2086), .Z(n2088) );
  NAND U2393 ( .A(n2089), .B(n2088), .Z(n2150) );
  NANDN U2394 ( .A(n2091), .B(n2090), .Z(n2095) );
  NAND U2395 ( .A(n2093), .B(n2092), .Z(n2094) );
  NAND U2396 ( .A(n2095), .B(n2094), .Z(n2148) );
  XNOR U2397 ( .A(b[7]), .B(a[38]), .Z(n2135) );
  NANDN U2398 ( .A(n2135), .B(n10545), .Z(n2098) );
  NANDN U2399 ( .A(n2096), .B(n10546), .Z(n2097) );
  NAND U2400 ( .A(n2098), .B(n2097), .Z(n2123) );
  XNOR U2401 ( .A(b[3]), .B(a[42]), .Z(n2138) );
  NANDN U2402 ( .A(n2138), .B(n10398), .Z(n2101) );
  NANDN U2403 ( .A(n2099), .B(n10399), .Z(n2100) );
  AND U2404 ( .A(n2101), .B(n2100), .Z(n2124) );
  XNOR U2405 ( .A(n2123), .B(n2124), .Z(n2125) );
  NANDN U2406 ( .A(n527), .B(a[44]), .Z(n2102) );
  XOR U2407 ( .A(n10434), .B(n2102), .Z(n2104) );
  IV U2408 ( .A(a[43]), .Z(n2369) );
  NANDN U2409 ( .A(n2369), .B(n527), .Z(n2103) );
  AND U2410 ( .A(n2104), .B(n2103), .Z(n2131) );
  XOR U2411 ( .A(b[5]), .B(a[40]), .Z(n2144) );
  NAND U2412 ( .A(n2144), .B(n10481), .Z(n2107) );
  NAND U2413 ( .A(n2105), .B(n10482), .Z(n2106) );
  NAND U2414 ( .A(n2107), .B(n2106), .Z(n2129) );
  NANDN U2415 ( .A(n529), .B(a[36]), .Z(n2130) );
  XNOR U2416 ( .A(n2129), .B(n2130), .Z(n2132) );
  XOR U2417 ( .A(n2131), .B(n2132), .Z(n2126) );
  XOR U2418 ( .A(n2125), .B(n2126), .Z(n2147) );
  XOR U2419 ( .A(n2148), .B(n2147), .Z(n2149) );
  XNOR U2420 ( .A(n2150), .B(n2149), .Z(n2119) );
  NAND U2421 ( .A(n2109), .B(n2108), .Z(n2113) );
  NAND U2422 ( .A(n2111), .B(n2110), .Z(n2112) );
  NAND U2423 ( .A(n2113), .B(n2112), .Z(n2120) );
  XNOR U2424 ( .A(n2119), .B(n2120), .Z(n2121) );
  XNOR U2425 ( .A(n2122), .B(n2121), .Z(n2153) );
  XNOR U2426 ( .A(n2153), .B(sreg[292]), .Z(n2155) );
  NAND U2427 ( .A(n2114), .B(sreg[291]), .Z(n2118) );
  OR U2428 ( .A(n2116), .B(n2115), .Z(n2117) );
  AND U2429 ( .A(n2118), .B(n2117), .Z(n2154) );
  XOR U2430 ( .A(n2155), .B(n2154), .Z(c[292]) );
  NANDN U2431 ( .A(n2124), .B(n2123), .Z(n2128) );
  NAND U2432 ( .A(n2126), .B(n2125), .Z(n2127) );
  NAND U2433 ( .A(n2128), .B(n2127), .Z(n2189) );
  NANDN U2434 ( .A(n2130), .B(n2129), .Z(n2134) );
  NAND U2435 ( .A(n2132), .B(n2131), .Z(n2133) );
  NAND U2436 ( .A(n2134), .B(n2133), .Z(n2187) );
  XNOR U2437 ( .A(b[7]), .B(a[39]), .Z(n2174) );
  NANDN U2438 ( .A(n2174), .B(n10545), .Z(n2137) );
  NANDN U2439 ( .A(n2135), .B(n10546), .Z(n2136) );
  NAND U2440 ( .A(n2137), .B(n2136), .Z(n2162) );
  XOR U2441 ( .A(b[3]), .B(n2369), .Z(n2177) );
  NANDN U2442 ( .A(n2177), .B(n10398), .Z(n2140) );
  NANDN U2443 ( .A(n2138), .B(n10399), .Z(n2139) );
  AND U2444 ( .A(n2140), .B(n2139), .Z(n2163) );
  XNOR U2445 ( .A(n2162), .B(n2163), .Z(n2164) );
  NANDN U2446 ( .A(n527), .B(a[45]), .Z(n2141) );
  XOR U2447 ( .A(n10434), .B(n2141), .Z(n2143) );
  NANDN U2448 ( .A(b[0]), .B(a[44]), .Z(n2142) );
  AND U2449 ( .A(n2143), .B(n2142), .Z(n2170) );
  XOR U2450 ( .A(b[5]), .B(a[41]), .Z(n2183) );
  NAND U2451 ( .A(n2183), .B(n10481), .Z(n2146) );
  NAND U2452 ( .A(n2144), .B(n10482), .Z(n2145) );
  NAND U2453 ( .A(n2146), .B(n2145), .Z(n2168) );
  NANDN U2454 ( .A(n529), .B(a[37]), .Z(n2169) );
  XNOR U2455 ( .A(n2168), .B(n2169), .Z(n2171) );
  XOR U2456 ( .A(n2170), .B(n2171), .Z(n2165) );
  XOR U2457 ( .A(n2164), .B(n2165), .Z(n2186) );
  XOR U2458 ( .A(n2187), .B(n2186), .Z(n2188) );
  XNOR U2459 ( .A(n2189), .B(n2188), .Z(n2158) );
  NAND U2460 ( .A(n2148), .B(n2147), .Z(n2152) );
  NAND U2461 ( .A(n2150), .B(n2149), .Z(n2151) );
  NAND U2462 ( .A(n2152), .B(n2151), .Z(n2159) );
  XNOR U2463 ( .A(n2158), .B(n2159), .Z(n2160) );
  XNOR U2464 ( .A(n2161), .B(n2160), .Z(n2192) );
  XNOR U2465 ( .A(n2192), .B(sreg[293]), .Z(n2194) );
  NAND U2466 ( .A(n2153), .B(sreg[292]), .Z(n2157) );
  OR U2467 ( .A(n2155), .B(n2154), .Z(n2156) );
  AND U2468 ( .A(n2157), .B(n2156), .Z(n2193) );
  XOR U2469 ( .A(n2194), .B(n2193), .Z(c[293]) );
  NANDN U2470 ( .A(n2163), .B(n2162), .Z(n2167) );
  NAND U2471 ( .A(n2165), .B(n2164), .Z(n2166) );
  NAND U2472 ( .A(n2167), .B(n2166), .Z(n2228) );
  NANDN U2473 ( .A(n2169), .B(n2168), .Z(n2173) );
  NAND U2474 ( .A(n2171), .B(n2170), .Z(n2172) );
  NAND U2475 ( .A(n2173), .B(n2172), .Z(n2226) );
  XNOR U2476 ( .A(b[7]), .B(a[40]), .Z(n2213) );
  NANDN U2477 ( .A(n2213), .B(n10545), .Z(n2176) );
  NANDN U2478 ( .A(n2174), .B(n10546), .Z(n2175) );
  NAND U2479 ( .A(n2176), .B(n2175), .Z(n2201) );
  XNOR U2480 ( .A(b[3]), .B(a[44]), .Z(n2216) );
  NANDN U2481 ( .A(n2216), .B(n10398), .Z(n2179) );
  NANDN U2482 ( .A(n2177), .B(n10399), .Z(n2178) );
  AND U2483 ( .A(n2179), .B(n2178), .Z(n2202) );
  XNOR U2484 ( .A(n2201), .B(n2202), .Z(n2203) );
  NANDN U2485 ( .A(n527), .B(a[46]), .Z(n2180) );
  XOR U2486 ( .A(n10434), .B(n2180), .Z(n2182) );
  NANDN U2487 ( .A(b[0]), .B(a[45]), .Z(n2181) );
  AND U2488 ( .A(n2182), .B(n2181), .Z(n2209) );
  XOR U2489 ( .A(b[5]), .B(a[42]), .Z(n2222) );
  NAND U2490 ( .A(n2222), .B(n10481), .Z(n2185) );
  NAND U2491 ( .A(n2183), .B(n10482), .Z(n2184) );
  NAND U2492 ( .A(n2185), .B(n2184), .Z(n2207) );
  NANDN U2493 ( .A(n529), .B(a[38]), .Z(n2208) );
  XNOR U2494 ( .A(n2207), .B(n2208), .Z(n2210) );
  XOR U2495 ( .A(n2209), .B(n2210), .Z(n2204) );
  XOR U2496 ( .A(n2203), .B(n2204), .Z(n2225) );
  XOR U2497 ( .A(n2226), .B(n2225), .Z(n2227) );
  XNOR U2498 ( .A(n2228), .B(n2227), .Z(n2197) );
  NAND U2499 ( .A(n2187), .B(n2186), .Z(n2191) );
  NAND U2500 ( .A(n2189), .B(n2188), .Z(n2190) );
  NAND U2501 ( .A(n2191), .B(n2190), .Z(n2198) );
  XNOR U2502 ( .A(n2197), .B(n2198), .Z(n2199) );
  XNOR U2503 ( .A(n2200), .B(n2199), .Z(n2231) );
  XNOR U2504 ( .A(n2231), .B(sreg[294]), .Z(n2233) );
  NAND U2505 ( .A(n2192), .B(sreg[293]), .Z(n2196) );
  OR U2506 ( .A(n2194), .B(n2193), .Z(n2195) );
  AND U2507 ( .A(n2196), .B(n2195), .Z(n2232) );
  XOR U2508 ( .A(n2233), .B(n2232), .Z(c[294]) );
  NANDN U2509 ( .A(n2202), .B(n2201), .Z(n2206) );
  NAND U2510 ( .A(n2204), .B(n2203), .Z(n2205) );
  NAND U2511 ( .A(n2206), .B(n2205), .Z(n2267) );
  NANDN U2512 ( .A(n2208), .B(n2207), .Z(n2212) );
  NAND U2513 ( .A(n2210), .B(n2209), .Z(n2211) );
  NAND U2514 ( .A(n2212), .B(n2211), .Z(n2265) );
  XNOR U2515 ( .A(b[7]), .B(a[41]), .Z(n2252) );
  NANDN U2516 ( .A(n2252), .B(n10545), .Z(n2215) );
  NANDN U2517 ( .A(n2213), .B(n10546), .Z(n2214) );
  NAND U2518 ( .A(n2215), .B(n2214), .Z(n2240) );
  XNOR U2519 ( .A(b[3]), .B(a[45]), .Z(n2255) );
  NANDN U2520 ( .A(n2255), .B(n10398), .Z(n2218) );
  NANDN U2521 ( .A(n2216), .B(n10399), .Z(n2217) );
  AND U2522 ( .A(n2218), .B(n2217), .Z(n2241) );
  XNOR U2523 ( .A(n2240), .B(n2241), .Z(n2242) );
  NANDN U2524 ( .A(n527), .B(a[47]), .Z(n2219) );
  XOR U2525 ( .A(n10434), .B(n2219), .Z(n2221) );
  NANDN U2526 ( .A(b[0]), .B(a[46]), .Z(n2220) );
  AND U2527 ( .A(n2221), .B(n2220), .Z(n2248) );
  XNOR U2528 ( .A(b[5]), .B(a[43]), .Z(n2261) );
  NANDN U2529 ( .A(n2261), .B(n10481), .Z(n2224) );
  NAND U2530 ( .A(n2222), .B(n10482), .Z(n2223) );
  NAND U2531 ( .A(n2224), .B(n2223), .Z(n2246) );
  NANDN U2532 ( .A(n529), .B(a[39]), .Z(n2247) );
  XNOR U2533 ( .A(n2246), .B(n2247), .Z(n2249) );
  XOR U2534 ( .A(n2248), .B(n2249), .Z(n2243) );
  XOR U2535 ( .A(n2242), .B(n2243), .Z(n2264) );
  XOR U2536 ( .A(n2265), .B(n2264), .Z(n2266) );
  XNOR U2537 ( .A(n2267), .B(n2266), .Z(n2236) );
  NAND U2538 ( .A(n2226), .B(n2225), .Z(n2230) );
  NAND U2539 ( .A(n2228), .B(n2227), .Z(n2229) );
  NAND U2540 ( .A(n2230), .B(n2229), .Z(n2237) );
  XNOR U2541 ( .A(n2236), .B(n2237), .Z(n2238) );
  XNOR U2542 ( .A(n2239), .B(n2238), .Z(n2270) );
  XNOR U2543 ( .A(n2270), .B(sreg[295]), .Z(n2272) );
  NAND U2544 ( .A(n2231), .B(sreg[294]), .Z(n2235) );
  OR U2545 ( .A(n2233), .B(n2232), .Z(n2234) );
  AND U2546 ( .A(n2235), .B(n2234), .Z(n2271) );
  XOR U2547 ( .A(n2272), .B(n2271), .Z(c[295]) );
  NANDN U2548 ( .A(n2241), .B(n2240), .Z(n2245) );
  NAND U2549 ( .A(n2243), .B(n2242), .Z(n2244) );
  NAND U2550 ( .A(n2245), .B(n2244), .Z(n2306) );
  NANDN U2551 ( .A(n2247), .B(n2246), .Z(n2251) );
  NAND U2552 ( .A(n2249), .B(n2248), .Z(n2250) );
  NAND U2553 ( .A(n2251), .B(n2250), .Z(n2304) );
  XNOR U2554 ( .A(b[7]), .B(a[42]), .Z(n2291) );
  NANDN U2555 ( .A(n2291), .B(n10545), .Z(n2254) );
  NANDN U2556 ( .A(n2252), .B(n10546), .Z(n2253) );
  NAND U2557 ( .A(n2254), .B(n2253), .Z(n2279) );
  XNOR U2558 ( .A(b[3]), .B(a[46]), .Z(n2294) );
  NANDN U2559 ( .A(n2294), .B(n10398), .Z(n2257) );
  NANDN U2560 ( .A(n2255), .B(n10399), .Z(n2256) );
  AND U2561 ( .A(n2257), .B(n2256), .Z(n2280) );
  XNOR U2562 ( .A(n2279), .B(n2280), .Z(n2281) );
  NANDN U2563 ( .A(n527), .B(a[48]), .Z(n2258) );
  XOR U2564 ( .A(n10434), .B(n2258), .Z(n2260) );
  NANDN U2565 ( .A(b[0]), .B(a[47]), .Z(n2259) );
  AND U2566 ( .A(n2260), .B(n2259), .Z(n2287) );
  XOR U2567 ( .A(b[5]), .B(a[44]), .Z(n2300) );
  NAND U2568 ( .A(n2300), .B(n10481), .Z(n2263) );
  NANDN U2569 ( .A(n2261), .B(n10482), .Z(n2262) );
  NAND U2570 ( .A(n2263), .B(n2262), .Z(n2285) );
  NANDN U2571 ( .A(n529), .B(a[40]), .Z(n2286) );
  XNOR U2572 ( .A(n2285), .B(n2286), .Z(n2288) );
  XOR U2573 ( .A(n2287), .B(n2288), .Z(n2282) );
  XOR U2574 ( .A(n2281), .B(n2282), .Z(n2303) );
  XOR U2575 ( .A(n2304), .B(n2303), .Z(n2305) );
  XNOR U2576 ( .A(n2306), .B(n2305), .Z(n2275) );
  NAND U2577 ( .A(n2265), .B(n2264), .Z(n2269) );
  NAND U2578 ( .A(n2267), .B(n2266), .Z(n2268) );
  NAND U2579 ( .A(n2269), .B(n2268), .Z(n2276) );
  XNOR U2580 ( .A(n2275), .B(n2276), .Z(n2277) );
  XNOR U2581 ( .A(n2278), .B(n2277), .Z(n2309) );
  XNOR U2582 ( .A(n2309), .B(sreg[296]), .Z(n2311) );
  NAND U2583 ( .A(n2270), .B(sreg[295]), .Z(n2274) );
  OR U2584 ( .A(n2272), .B(n2271), .Z(n2273) );
  AND U2585 ( .A(n2274), .B(n2273), .Z(n2310) );
  XOR U2586 ( .A(n2311), .B(n2310), .Z(c[296]) );
  NANDN U2587 ( .A(n2280), .B(n2279), .Z(n2284) );
  NAND U2588 ( .A(n2282), .B(n2281), .Z(n2283) );
  NAND U2589 ( .A(n2284), .B(n2283), .Z(n2345) );
  NANDN U2590 ( .A(n2286), .B(n2285), .Z(n2290) );
  NAND U2591 ( .A(n2288), .B(n2287), .Z(n2289) );
  NAND U2592 ( .A(n2290), .B(n2289), .Z(n2343) );
  XOR U2593 ( .A(b[7]), .B(n2369), .Z(n2330) );
  NANDN U2594 ( .A(n2330), .B(n10545), .Z(n2293) );
  NANDN U2595 ( .A(n2291), .B(n10546), .Z(n2292) );
  NAND U2596 ( .A(n2293), .B(n2292), .Z(n2318) );
  XNOR U2597 ( .A(b[3]), .B(a[47]), .Z(n2333) );
  NANDN U2598 ( .A(n2333), .B(n10398), .Z(n2296) );
  NANDN U2599 ( .A(n2294), .B(n10399), .Z(n2295) );
  AND U2600 ( .A(n2296), .B(n2295), .Z(n2319) );
  XNOR U2601 ( .A(n2318), .B(n2319), .Z(n2320) );
  NANDN U2602 ( .A(n527), .B(a[49]), .Z(n2297) );
  XOR U2603 ( .A(n10434), .B(n2297), .Z(n2299) );
  NANDN U2604 ( .A(b[0]), .B(a[48]), .Z(n2298) );
  AND U2605 ( .A(n2299), .B(n2298), .Z(n2326) );
  XOR U2606 ( .A(b[5]), .B(a[45]), .Z(n2339) );
  NAND U2607 ( .A(n2339), .B(n10481), .Z(n2302) );
  NAND U2608 ( .A(n2300), .B(n10482), .Z(n2301) );
  NAND U2609 ( .A(n2302), .B(n2301), .Z(n2324) );
  NANDN U2610 ( .A(n529), .B(a[41]), .Z(n2325) );
  XNOR U2611 ( .A(n2324), .B(n2325), .Z(n2327) );
  XOR U2612 ( .A(n2326), .B(n2327), .Z(n2321) );
  XOR U2613 ( .A(n2320), .B(n2321), .Z(n2342) );
  XOR U2614 ( .A(n2343), .B(n2342), .Z(n2344) );
  XNOR U2615 ( .A(n2345), .B(n2344), .Z(n2314) );
  NAND U2616 ( .A(n2304), .B(n2303), .Z(n2308) );
  NAND U2617 ( .A(n2306), .B(n2305), .Z(n2307) );
  NAND U2618 ( .A(n2308), .B(n2307), .Z(n2315) );
  XNOR U2619 ( .A(n2314), .B(n2315), .Z(n2316) );
  XNOR U2620 ( .A(n2317), .B(n2316), .Z(n2348) );
  XNOR U2621 ( .A(n2348), .B(sreg[297]), .Z(n2350) );
  NAND U2622 ( .A(n2309), .B(sreg[296]), .Z(n2313) );
  OR U2623 ( .A(n2311), .B(n2310), .Z(n2312) );
  AND U2624 ( .A(n2313), .B(n2312), .Z(n2349) );
  XOR U2625 ( .A(n2350), .B(n2349), .Z(c[297]) );
  NANDN U2626 ( .A(n2319), .B(n2318), .Z(n2323) );
  NAND U2627 ( .A(n2321), .B(n2320), .Z(n2322) );
  NAND U2628 ( .A(n2323), .B(n2322), .Z(n2385) );
  NANDN U2629 ( .A(n2325), .B(n2324), .Z(n2329) );
  NAND U2630 ( .A(n2327), .B(n2326), .Z(n2328) );
  NAND U2631 ( .A(n2329), .B(n2328), .Z(n2383) );
  XNOR U2632 ( .A(b[7]), .B(a[44]), .Z(n2376) );
  NANDN U2633 ( .A(n2376), .B(n10545), .Z(n2332) );
  NANDN U2634 ( .A(n2330), .B(n10546), .Z(n2331) );
  NAND U2635 ( .A(n2332), .B(n2331), .Z(n2357) );
  XNOR U2636 ( .A(b[3]), .B(a[48]), .Z(n2379) );
  NANDN U2637 ( .A(n2379), .B(n10398), .Z(n2335) );
  NANDN U2638 ( .A(n2333), .B(n10399), .Z(n2334) );
  AND U2639 ( .A(n2335), .B(n2334), .Z(n2358) );
  XNOR U2640 ( .A(n2357), .B(n2358), .Z(n2359) );
  NANDN U2641 ( .A(n527), .B(a[50]), .Z(n2336) );
  XOR U2642 ( .A(n10434), .B(n2336), .Z(n2338) );
  NANDN U2643 ( .A(b[0]), .B(a[49]), .Z(n2337) );
  AND U2644 ( .A(n2338), .B(n2337), .Z(n2365) );
  XOR U2645 ( .A(b[5]), .B(a[46]), .Z(n2370) );
  NAND U2646 ( .A(n2370), .B(n10481), .Z(n2341) );
  NAND U2647 ( .A(n2339), .B(n10482), .Z(n2340) );
  NAND U2648 ( .A(n2341), .B(n2340), .Z(n2363) );
  NANDN U2649 ( .A(n529), .B(a[42]), .Z(n2364) );
  XNOR U2650 ( .A(n2363), .B(n2364), .Z(n2366) );
  XOR U2651 ( .A(n2365), .B(n2366), .Z(n2360) );
  XOR U2652 ( .A(n2359), .B(n2360), .Z(n2382) );
  XOR U2653 ( .A(n2383), .B(n2382), .Z(n2384) );
  XNOR U2654 ( .A(n2385), .B(n2384), .Z(n2353) );
  NAND U2655 ( .A(n2343), .B(n2342), .Z(n2347) );
  NAND U2656 ( .A(n2345), .B(n2344), .Z(n2346) );
  NAND U2657 ( .A(n2347), .B(n2346), .Z(n2354) );
  XNOR U2658 ( .A(n2353), .B(n2354), .Z(n2355) );
  XNOR U2659 ( .A(n2356), .B(n2355), .Z(n2388) );
  XNOR U2660 ( .A(n2388), .B(sreg[298]), .Z(n2390) );
  NAND U2661 ( .A(n2348), .B(sreg[297]), .Z(n2352) );
  OR U2662 ( .A(n2350), .B(n2349), .Z(n2351) );
  AND U2663 ( .A(n2352), .B(n2351), .Z(n2389) );
  XOR U2664 ( .A(n2390), .B(n2389), .Z(c[298]) );
  NANDN U2665 ( .A(n2358), .B(n2357), .Z(n2362) );
  NAND U2666 ( .A(n2360), .B(n2359), .Z(n2361) );
  NAND U2667 ( .A(n2362), .B(n2361), .Z(n2424) );
  NANDN U2668 ( .A(n2364), .B(n2363), .Z(n2368) );
  NAND U2669 ( .A(n2366), .B(n2365), .Z(n2367) );
  NAND U2670 ( .A(n2368), .B(n2367), .Z(n2421) );
  ANDN U2671 ( .B(b[7]), .A(n2369), .Z(n2403) );
  XOR U2672 ( .A(b[5]), .B(a[47]), .Z(n2418) );
  NAND U2673 ( .A(n10481), .B(n2418), .Z(n2372) );
  NAND U2674 ( .A(n10482), .B(n2370), .Z(n2371) );
  NAND U2675 ( .A(n2372), .B(n2371), .Z(n2404) );
  XOR U2676 ( .A(n2403), .B(n2404), .Z(n2405) );
  NANDN U2677 ( .A(n527), .B(a[51]), .Z(n2373) );
  XOR U2678 ( .A(n10434), .B(n2373), .Z(n2375) );
  NANDN U2679 ( .A(b[0]), .B(a[50]), .Z(n2374) );
  AND U2680 ( .A(n2375), .B(n2374), .Z(n2406) );
  XOR U2681 ( .A(n2405), .B(n2406), .Z(n2400) );
  XNOR U2682 ( .A(b[7]), .B(a[45]), .Z(n2409) );
  NANDN U2683 ( .A(n2409), .B(n10545), .Z(n2378) );
  NANDN U2684 ( .A(n2376), .B(n10546), .Z(n2377) );
  NAND U2685 ( .A(n2378), .B(n2377), .Z(n2397) );
  XNOR U2686 ( .A(b[3]), .B(a[49]), .Z(n2412) );
  NANDN U2687 ( .A(n2412), .B(n10398), .Z(n2381) );
  NANDN U2688 ( .A(n2379), .B(n10399), .Z(n2380) );
  AND U2689 ( .A(n2381), .B(n2380), .Z(n2398) );
  XNOR U2690 ( .A(n2397), .B(n2398), .Z(n2399) );
  XNOR U2691 ( .A(n2400), .B(n2399), .Z(n2422) );
  XNOR U2692 ( .A(n2421), .B(n2422), .Z(n2423) );
  XNOR U2693 ( .A(n2424), .B(n2423), .Z(n2393) );
  NAND U2694 ( .A(n2383), .B(n2382), .Z(n2387) );
  NAND U2695 ( .A(n2385), .B(n2384), .Z(n2386) );
  NAND U2696 ( .A(n2387), .B(n2386), .Z(n2394) );
  XNOR U2697 ( .A(n2393), .B(n2394), .Z(n2395) );
  XNOR U2698 ( .A(n2396), .B(n2395), .Z(n2427) );
  XNOR U2699 ( .A(n2427), .B(sreg[299]), .Z(n2429) );
  NAND U2700 ( .A(n2388), .B(sreg[298]), .Z(n2392) );
  OR U2701 ( .A(n2390), .B(n2389), .Z(n2391) );
  AND U2702 ( .A(n2392), .B(n2391), .Z(n2428) );
  XOR U2703 ( .A(n2429), .B(n2428), .Z(c[299]) );
  NANDN U2704 ( .A(n2398), .B(n2397), .Z(n2402) );
  NAND U2705 ( .A(n2400), .B(n2399), .Z(n2401) );
  NAND U2706 ( .A(n2402), .B(n2401), .Z(n2463) );
  OR U2707 ( .A(n2404), .B(n2403), .Z(n2408) );
  NANDN U2708 ( .A(n2406), .B(n2405), .Z(n2407) );
  NAND U2709 ( .A(n2408), .B(n2407), .Z(n2461) );
  XNOR U2710 ( .A(b[7]), .B(a[46]), .Z(n2448) );
  NANDN U2711 ( .A(n2448), .B(n10545), .Z(n2411) );
  NANDN U2712 ( .A(n2409), .B(n10546), .Z(n2410) );
  NAND U2713 ( .A(n2411), .B(n2410), .Z(n2436) );
  XNOR U2714 ( .A(b[3]), .B(a[50]), .Z(n2451) );
  NANDN U2715 ( .A(n2451), .B(n10398), .Z(n2414) );
  NANDN U2716 ( .A(n2412), .B(n10399), .Z(n2413) );
  AND U2717 ( .A(n2414), .B(n2413), .Z(n2437) );
  XNOR U2718 ( .A(n2436), .B(n2437), .Z(n2438) );
  NANDN U2719 ( .A(n527), .B(a[52]), .Z(n2415) );
  XOR U2720 ( .A(n10434), .B(n2415), .Z(n2417) );
  NANDN U2721 ( .A(b[0]), .B(a[51]), .Z(n2416) );
  AND U2722 ( .A(n2417), .B(n2416), .Z(n2444) );
  XOR U2723 ( .A(b[5]), .B(a[48]), .Z(n2457) );
  NAND U2724 ( .A(n2457), .B(n10481), .Z(n2420) );
  NAND U2725 ( .A(n2418), .B(n10482), .Z(n2419) );
  NAND U2726 ( .A(n2420), .B(n2419), .Z(n2442) );
  NANDN U2727 ( .A(n529), .B(a[44]), .Z(n2443) );
  XNOR U2728 ( .A(n2442), .B(n2443), .Z(n2445) );
  XOR U2729 ( .A(n2444), .B(n2445), .Z(n2439) );
  XOR U2730 ( .A(n2438), .B(n2439), .Z(n2460) );
  XNOR U2731 ( .A(n2461), .B(n2460), .Z(n2462) );
  XNOR U2732 ( .A(n2463), .B(n2462), .Z(n2432) );
  NANDN U2733 ( .A(n2422), .B(n2421), .Z(n2426) );
  NAND U2734 ( .A(n2424), .B(n2423), .Z(n2425) );
  NAND U2735 ( .A(n2426), .B(n2425), .Z(n2433) );
  XNOR U2736 ( .A(n2432), .B(n2433), .Z(n2434) );
  XNOR U2737 ( .A(n2435), .B(n2434), .Z(n2464) );
  XNOR U2738 ( .A(n2464), .B(sreg[300]), .Z(n2466) );
  NAND U2739 ( .A(n2427), .B(sreg[299]), .Z(n2431) );
  OR U2740 ( .A(n2429), .B(n2428), .Z(n2430) );
  AND U2741 ( .A(n2431), .B(n2430), .Z(n2465) );
  XOR U2742 ( .A(n2466), .B(n2465), .Z(c[300]) );
  NANDN U2743 ( .A(n2437), .B(n2436), .Z(n2441) );
  NAND U2744 ( .A(n2439), .B(n2438), .Z(n2440) );
  NAND U2745 ( .A(n2441), .B(n2440), .Z(n2500) );
  NANDN U2746 ( .A(n2443), .B(n2442), .Z(n2447) );
  NAND U2747 ( .A(n2445), .B(n2444), .Z(n2446) );
  NAND U2748 ( .A(n2447), .B(n2446), .Z(n2498) );
  XNOR U2749 ( .A(b[7]), .B(a[47]), .Z(n2485) );
  NANDN U2750 ( .A(n2485), .B(n10545), .Z(n2450) );
  NANDN U2751 ( .A(n2448), .B(n10546), .Z(n2449) );
  NAND U2752 ( .A(n2450), .B(n2449), .Z(n2473) );
  XNOR U2753 ( .A(b[3]), .B(a[51]), .Z(n2488) );
  NANDN U2754 ( .A(n2488), .B(n10398), .Z(n2453) );
  NANDN U2755 ( .A(n2451), .B(n10399), .Z(n2452) );
  AND U2756 ( .A(n2453), .B(n2452), .Z(n2474) );
  XNOR U2757 ( .A(n2473), .B(n2474), .Z(n2475) );
  NANDN U2758 ( .A(n527), .B(a[53]), .Z(n2454) );
  XOR U2759 ( .A(n10434), .B(n2454), .Z(n2456) );
  NANDN U2760 ( .A(b[0]), .B(a[52]), .Z(n2455) );
  AND U2761 ( .A(n2456), .B(n2455), .Z(n2481) );
  XOR U2762 ( .A(b[5]), .B(a[49]), .Z(n2494) );
  NAND U2763 ( .A(n2494), .B(n10481), .Z(n2459) );
  NAND U2764 ( .A(n2457), .B(n10482), .Z(n2458) );
  NAND U2765 ( .A(n2459), .B(n2458), .Z(n2479) );
  NANDN U2766 ( .A(n529), .B(a[45]), .Z(n2480) );
  XNOR U2767 ( .A(n2479), .B(n2480), .Z(n2482) );
  XOR U2768 ( .A(n2481), .B(n2482), .Z(n2476) );
  XOR U2769 ( .A(n2475), .B(n2476), .Z(n2497) );
  XOR U2770 ( .A(n2498), .B(n2497), .Z(n2499) );
  XNOR U2771 ( .A(n2500), .B(n2499), .Z(n2469) );
  XNOR U2772 ( .A(n2469), .B(n2470), .Z(n2471) );
  XNOR U2773 ( .A(n2472), .B(n2471), .Z(n2503) );
  XNOR U2774 ( .A(n2503), .B(sreg[301]), .Z(n2505) );
  NAND U2775 ( .A(n2464), .B(sreg[300]), .Z(n2468) );
  OR U2776 ( .A(n2466), .B(n2465), .Z(n2467) );
  AND U2777 ( .A(n2468), .B(n2467), .Z(n2504) );
  XOR U2778 ( .A(n2505), .B(n2504), .Z(c[301]) );
  NANDN U2779 ( .A(n2474), .B(n2473), .Z(n2478) );
  NAND U2780 ( .A(n2476), .B(n2475), .Z(n2477) );
  NAND U2781 ( .A(n2478), .B(n2477), .Z(n2539) );
  NANDN U2782 ( .A(n2480), .B(n2479), .Z(n2484) );
  NAND U2783 ( .A(n2482), .B(n2481), .Z(n2483) );
  NAND U2784 ( .A(n2484), .B(n2483), .Z(n2537) );
  XNOR U2785 ( .A(b[7]), .B(a[48]), .Z(n2524) );
  NANDN U2786 ( .A(n2524), .B(n10545), .Z(n2487) );
  NANDN U2787 ( .A(n2485), .B(n10546), .Z(n2486) );
  NAND U2788 ( .A(n2487), .B(n2486), .Z(n2512) );
  XNOR U2789 ( .A(b[3]), .B(a[52]), .Z(n2527) );
  NANDN U2790 ( .A(n2527), .B(n10398), .Z(n2490) );
  NANDN U2791 ( .A(n2488), .B(n10399), .Z(n2489) );
  AND U2792 ( .A(n2490), .B(n2489), .Z(n2513) );
  XNOR U2793 ( .A(n2512), .B(n2513), .Z(n2514) );
  NANDN U2794 ( .A(n527), .B(a[54]), .Z(n2491) );
  XOR U2795 ( .A(n10434), .B(n2491), .Z(n2493) );
  NANDN U2796 ( .A(b[0]), .B(a[53]), .Z(n2492) );
  AND U2797 ( .A(n2493), .B(n2492), .Z(n2520) );
  XOR U2798 ( .A(b[5]), .B(a[50]), .Z(n2533) );
  NAND U2799 ( .A(n2533), .B(n10481), .Z(n2496) );
  NAND U2800 ( .A(n2494), .B(n10482), .Z(n2495) );
  NAND U2801 ( .A(n2496), .B(n2495), .Z(n2518) );
  NANDN U2802 ( .A(n529), .B(a[46]), .Z(n2519) );
  XNOR U2803 ( .A(n2518), .B(n2519), .Z(n2521) );
  XOR U2804 ( .A(n2520), .B(n2521), .Z(n2515) );
  XOR U2805 ( .A(n2514), .B(n2515), .Z(n2536) );
  XOR U2806 ( .A(n2537), .B(n2536), .Z(n2538) );
  XNOR U2807 ( .A(n2539), .B(n2538), .Z(n2508) );
  NAND U2808 ( .A(n2498), .B(n2497), .Z(n2502) );
  NAND U2809 ( .A(n2500), .B(n2499), .Z(n2501) );
  NAND U2810 ( .A(n2502), .B(n2501), .Z(n2509) );
  XNOR U2811 ( .A(n2508), .B(n2509), .Z(n2510) );
  XNOR U2812 ( .A(n2511), .B(n2510), .Z(n2542) );
  XNOR U2813 ( .A(n2542), .B(sreg[302]), .Z(n2544) );
  NAND U2814 ( .A(n2503), .B(sreg[301]), .Z(n2507) );
  OR U2815 ( .A(n2505), .B(n2504), .Z(n2506) );
  AND U2816 ( .A(n2507), .B(n2506), .Z(n2543) );
  XOR U2817 ( .A(n2544), .B(n2543), .Z(c[302]) );
  NANDN U2818 ( .A(n2513), .B(n2512), .Z(n2517) );
  NAND U2819 ( .A(n2515), .B(n2514), .Z(n2516) );
  NAND U2820 ( .A(n2517), .B(n2516), .Z(n2578) );
  NANDN U2821 ( .A(n2519), .B(n2518), .Z(n2523) );
  NAND U2822 ( .A(n2521), .B(n2520), .Z(n2522) );
  NAND U2823 ( .A(n2523), .B(n2522), .Z(n2576) );
  XNOR U2824 ( .A(b[7]), .B(a[49]), .Z(n2563) );
  NANDN U2825 ( .A(n2563), .B(n10545), .Z(n2526) );
  NANDN U2826 ( .A(n2524), .B(n10546), .Z(n2525) );
  NAND U2827 ( .A(n2526), .B(n2525), .Z(n2551) );
  XNOR U2828 ( .A(b[3]), .B(a[53]), .Z(n2566) );
  NANDN U2829 ( .A(n2566), .B(n10398), .Z(n2529) );
  NANDN U2830 ( .A(n2527), .B(n10399), .Z(n2528) );
  AND U2831 ( .A(n2529), .B(n2528), .Z(n2552) );
  XNOR U2832 ( .A(n2551), .B(n2552), .Z(n2553) );
  NANDN U2833 ( .A(n527), .B(a[55]), .Z(n2530) );
  XOR U2834 ( .A(n10434), .B(n2530), .Z(n2532) );
  NANDN U2835 ( .A(b[0]), .B(a[54]), .Z(n2531) );
  AND U2836 ( .A(n2532), .B(n2531), .Z(n2559) );
  XOR U2837 ( .A(b[5]), .B(a[51]), .Z(n2572) );
  NAND U2838 ( .A(n2572), .B(n10481), .Z(n2535) );
  NAND U2839 ( .A(n2533), .B(n10482), .Z(n2534) );
  NAND U2840 ( .A(n2535), .B(n2534), .Z(n2557) );
  NANDN U2841 ( .A(n529), .B(a[47]), .Z(n2558) );
  XNOR U2842 ( .A(n2557), .B(n2558), .Z(n2560) );
  XOR U2843 ( .A(n2559), .B(n2560), .Z(n2554) );
  XOR U2844 ( .A(n2553), .B(n2554), .Z(n2575) );
  XOR U2845 ( .A(n2576), .B(n2575), .Z(n2577) );
  XNOR U2846 ( .A(n2578), .B(n2577), .Z(n2547) );
  NAND U2847 ( .A(n2537), .B(n2536), .Z(n2541) );
  NAND U2848 ( .A(n2539), .B(n2538), .Z(n2540) );
  NAND U2849 ( .A(n2541), .B(n2540), .Z(n2548) );
  XNOR U2850 ( .A(n2547), .B(n2548), .Z(n2549) );
  XNOR U2851 ( .A(n2550), .B(n2549), .Z(n2581) );
  XNOR U2852 ( .A(n2581), .B(sreg[303]), .Z(n2583) );
  NAND U2853 ( .A(n2542), .B(sreg[302]), .Z(n2546) );
  OR U2854 ( .A(n2544), .B(n2543), .Z(n2545) );
  AND U2855 ( .A(n2546), .B(n2545), .Z(n2582) );
  XOR U2856 ( .A(n2583), .B(n2582), .Z(c[303]) );
  NANDN U2857 ( .A(n2552), .B(n2551), .Z(n2556) );
  NAND U2858 ( .A(n2554), .B(n2553), .Z(n2555) );
  NAND U2859 ( .A(n2556), .B(n2555), .Z(n2617) );
  NANDN U2860 ( .A(n2558), .B(n2557), .Z(n2562) );
  NAND U2861 ( .A(n2560), .B(n2559), .Z(n2561) );
  NAND U2862 ( .A(n2562), .B(n2561), .Z(n2615) );
  XNOR U2863 ( .A(b[7]), .B(a[50]), .Z(n2590) );
  NANDN U2864 ( .A(n2590), .B(n10545), .Z(n2565) );
  NANDN U2865 ( .A(n2563), .B(n10546), .Z(n2564) );
  NAND U2866 ( .A(n2565), .B(n2564), .Z(n2608) );
  XNOR U2867 ( .A(b[3]), .B(a[54]), .Z(n2593) );
  NANDN U2868 ( .A(n2593), .B(n10398), .Z(n2568) );
  NANDN U2869 ( .A(n2566), .B(n10399), .Z(n2567) );
  AND U2870 ( .A(n2568), .B(n2567), .Z(n2609) );
  XNOR U2871 ( .A(n2608), .B(n2609), .Z(n2610) );
  NANDN U2872 ( .A(n527), .B(a[56]), .Z(n2569) );
  XOR U2873 ( .A(n10434), .B(n2569), .Z(n2571) );
  NANDN U2874 ( .A(b[0]), .B(a[55]), .Z(n2570) );
  AND U2875 ( .A(n2571), .B(n2570), .Z(n2604) );
  XOR U2876 ( .A(b[5]), .B(a[52]), .Z(n2599) );
  NAND U2877 ( .A(n2599), .B(n10481), .Z(n2574) );
  NAND U2878 ( .A(n2572), .B(n10482), .Z(n2573) );
  NAND U2879 ( .A(n2574), .B(n2573), .Z(n2602) );
  NANDN U2880 ( .A(n529), .B(a[48]), .Z(n2603) );
  XNOR U2881 ( .A(n2602), .B(n2603), .Z(n2605) );
  XOR U2882 ( .A(n2604), .B(n2605), .Z(n2611) );
  XOR U2883 ( .A(n2610), .B(n2611), .Z(n2614) );
  XOR U2884 ( .A(n2615), .B(n2614), .Z(n2616) );
  XNOR U2885 ( .A(n2617), .B(n2616), .Z(n2586) );
  NAND U2886 ( .A(n2576), .B(n2575), .Z(n2580) );
  NAND U2887 ( .A(n2578), .B(n2577), .Z(n2579) );
  NAND U2888 ( .A(n2580), .B(n2579), .Z(n2587) );
  XNOR U2889 ( .A(n2586), .B(n2587), .Z(n2588) );
  XNOR U2890 ( .A(n2589), .B(n2588), .Z(n2620) );
  XNOR U2891 ( .A(n2620), .B(sreg[304]), .Z(n2622) );
  NAND U2892 ( .A(n2581), .B(sreg[303]), .Z(n2585) );
  OR U2893 ( .A(n2583), .B(n2582), .Z(n2584) );
  AND U2894 ( .A(n2585), .B(n2584), .Z(n2621) );
  XOR U2895 ( .A(n2622), .B(n2621), .Z(c[304]) );
  XNOR U2896 ( .A(b[7]), .B(a[51]), .Z(n2641) );
  NANDN U2897 ( .A(n2641), .B(n10545), .Z(n2592) );
  NANDN U2898 ( .A(n2590), .B(n10546), .Z(n2591) );
  NAND U2899 ( .A(n2592), .B(n2591), .Z(n2629) );
  XNOR U2900 ( .A(b[3]), .B(a[55]), .Z(n2644) );
  NANDN U2901 ( .A(n2644), .B(n10398), .Z(n2595) );
  NANDN U2902 ( .A(n2593), .B(n10399), .Z(n2594) );
  AND U2903 ( .A(n2595), .B(n2594), .Z(n2630) );
  XNOR U2904 ( .A(n2629), .B(n2630), .Z(n2631) );
  NANDN U2905 ( .A(n527), .B(a[57]), .Z(n2596) );
  XOR U2906 ( .A(n10434), .B(n2596), .Z(n2598) );
  NANDN U2907 ( .A(b[0]), .B(a[56]), .Z(n2597) );
  AND U2908 ( .A(n2598), .B(n2597), .Z(n2637) );
  XOR U2909 ( .A(b[5]), .B(a[53]), .Z(n2650) );
  NAND U2910 ( .A(n2650), .B(n10481), .Z(n2601) );
  NAND U2911 ( .A(n2599), .B(n10482), .Z(n2600) );
  NAND U2912 ( .A(n2601), .B(n2600), .Z(n2635) );
  NANDN U2913 ( .A(n529), .B(a[49]), .Z(n2636) );
  XNOR U2914 ( .A(n2635), .B(n2636), .Z(n2638) );
  XOR U2915 ( .A(n2637), .B(n2638), .Z(n2632) );
  XOR U2916 ( .A(n2631), .B(n2632), .Z(n2655) );
  NANDN U2917 ( .A(n2603), .B(n2602), .Z(n2607) );
  NAND U2918 ( .A(n2605), .B(n2604), .Z(n2606) );
  NAND U2919 ( .A(n2607), .B(n2606), .Z(n2653) );
  NANDN U2920 ( .A(n2609), .B(n2608), .Z(n2613) );
  NAND U2921 ( .A(n2611), .B(n2610), .Z(n2612) );
  AND U2922 ( .A(n2613), .B(n2612), .Z(n2654) );
  XNOR U2923 ( .A(n2653), .B(n2654), .Z(n2656) );
  XNOR U2924 ( .A(n2655), .B(n2656), .Z(n2625) );
  NAND U2925 ( .A(n2615), .B(n2614), .Z(n2619) );
  NAND U2926 ( .A(n2617), .B(n2616), .Z(n2618) );
  NAND U2927 ( .A(n2619), .B(n2618), .Z(n2626) );
  XNOR U2928 ( .A(n2625), .B(n2626), .Z(n2627) );
  XNOR U2929 ( .A(n2628), .B(n2627), .Z(n2659) );
  XNOR U2930 ( .A(n2659), .B(sreg[305]), .Z(n2661) );
  NAND U2931 ( .A(n2620), .B(sreg[304]), .Z(n2624) );
  OR U2932 ( .A(n2622), .B(n2621), .Z(n2623) );
  AND U2933 ( .A(n2624), .B(n2623), .Z(n2660) );
  XOR U2934 ( .A(n2661), .B(n2660), .Z(c[305]) );
  NANDN U2935 ( .A(n2630), .B(n2629), .Z(n2634) );
  NAND U2936 ( .A(n2632), .B(n2631), .Z(n2633) );
  NAND U2937 ( .A(n2634), .B(n2633), .Z(n2695) );
  NANDN U2938 ( .A(n2636), .B(n2635), .Z(n2640) );
  NAND U2939 ( .A(n2638), .B(n2637), .Z(n2639) );
  NAND U2940 ( .A(n2640), .B(n2639), .Z(n2693) );
  XNOR U2941 ( .A(b[7]), .B(a[52]), .Z(n2680) );
  NANDN U2942 ( .A(n2680), .B(n10545), .Z(n2643) );
  NANDN U2943 ( .A(n2641), .B(n10546), .Z(n2642) );
  NAND U2944 ( .A(n2643), .B(n2642), .Z(n2668) );
  XNOR U2945 ( .A(b[3]), .B(a[56]), .Z(n2683) );
  NANDN U2946 ( .A(n2683), .B(n10398), .Z(n2646) );
  NANDN U2947 ( .A(n2644), .B(n10399), .Z(n2645) );
  AND U2948 ( .A(n2646), .B(n2645), .Z(n2669) );
  XNOR U2949 ( .A(n2668), .B(n2669), .Z(n2670) );
  NANDN U2950 ( .A(n527), .B(a[58]), .Z(n2647) );
  XOR U2951 ( .A(n10434), .B(n2647), .Z(n2649) );
  NANDN U2952 ( .A(b[0]), .B(a[57]), .Z(n2648) );
  AND U2953 ( .A(n2649), .B(n2648), .Z(n2676) );
  XOR U2954 ( .A(b[5]), .B(a[54]), .Z(n2689) );
  NAND U2955 ( .A(n2689), .B(n10481), .Z(n2652) );
  NAND U2956 ( .A(n2650), .B(n10482), .Z(n2651) );
  NAND U2957 ( .A(n2652), .B(n2651), .Z(n2674) );
  NANDN U2958 ( .A(n529), .B(a[50]), .Z(n2675) );
  XNOR U2959 ( .A(n2674), .B(n2675), .Z(n2677) );
  XOR U2960 ( .A(n2676), .B(n2677), .Z(n2671) );
  XOR U2961 ( .A(n2670), .B(n2671), .Z(n2692) );
  XOR U2962 ( .A(n2693), .B(n2692), .Z(n2694) );
  XNOR U2963 ( .A(n2695), .B(n2694), .Z(n2664) );
  NANDN U2964 ( .A(n2654), .B(n2653), .Z(n2658) );
  NAND U2965 ( .A(n2656), .B(n2655), .Z(n2657) );
  NAND U2966 ( .A(n2658), .B(n2657), .Z(n2665) );
  XNOR U2967 ( .A(n2664), .B(n2665), .Z(n2666) );
  XNOR U2968 ( .A(n2667), .B(n2666), .Z(n2698) );
  XNOR U2969 ( .A(n2698), .B(sreg[306]), .Z(n2700) );
  NAND U2970 ( .A(n2659), .B(sreg[305]), .Z(n2663) );
  OR U2971 ( .A(n2661), .B(n2660), .Z(n2662) );
  AND U2972 ( .A(n2663), .B(n2662), .Z(n2699) );
  XOR U2973 ( .A(n2700), .B(n2699), .Z(c[306]) );
  NANDN U2974 ( .A(n2669), .B(n2668), .Z(n2673) );
  NAND U2975 ( .A(n2671), .B(n2670), .Z(n2672) );
  NAND U2976 ( .A(n2673), .B(n2672), .Z(n2734) );
  NANDN U2977 ( .A(n2675), .B(n2674), .Z(n2679) );
  NAND U2978 ( .A(n2677), .B(n2676), .Z(n2678) );
  NAND U2979 ( .A(n2679), .B(n2678), .Z(n2732) );
  XNOR U2980 ( .A(b[7]), .B(a[53]), .Z(n2725) );
  NANDN U2981 ( .A(n2725), .B(n10545), .Z(n2682) );
  NANDN U2982 ( .A(n2680), .B(n10546), .Z(n2681) );
  NAND U2983 ( .A(n2682), .B(n2681), .Z(n2707) );
  XNOR U2984 ( .A(b[3]), .B(a[57]), .Z(n2728) );
  NANDN U2985 ( .A(n2728), .B(n10398), .Z(n2685) );
  NANDN U2986 ( .A(n2683), .B(n10399), .Z(n2684) );
  AND U2987 ( .A(n2685), .B(n2684), .Z(n2708) );
  XNOR U2988 ( .A(n2707), .B(n2708), .Z(n2709) );
  NANDN U2989 ( .A(n527), .B(a[59]), .Z(n2686) );
  XOR U2990 ( .A(n10434), .B(n2686), .Z(n2688) );
  NANDN U2991 ( .A(b[0]), .B(a[58]), .Z(n2687) );
  AND U2992 ( .A(n2688), .B(n2687), .Z(n2715) );
  XOR U2993 ( .A(b[5]), .B(a[55]), .Z(n2719) );
  NAND U2994 ( .A(n2719), .B(n10481), .Z(n2691) );
  NAND U2995 ( .A(n2689), .B(n10482), .Z(n2690) );
  NAND U2996 ( .A(n2691), .B(n2690), .Z(n2713) );
  NANDN U2997 ( .A(n529), .B(a[51]), .Z(n2714) );
  XNOR U2998 ( .A(n2713), .B(n2714), .Z(n2716) );
  XOR U2999 ( .A(n2715), .B(n2716), .Z(n2710) );
  XOR U3000 ( .A(n2709), .B(n2710), .Z(n2731) );
  XOR U3001 ( .A(n2732), .B(n2731), .Z(n2733) );
  XNOR U3002 ( .A(n2734), .B(n2733), .Z(n2703) );
  NAND U3003 ( .A(n2693), .B(n2692), .Z(n2697) );
  NAND U3004 ( .A(n2695), .B(n2694), .Z(n2696) );
  NAND U3005 ( .A(n2697), .B(n2696), .Z(n2704) );
  XNOR U3006 ( .A(n2703), .B(n2704), .Z(n2705) );
  XNOR U3007 ( .A(n2706), .B(n2705), .Z(n2737) );
  XNOR U3008 ( .A(n2737), .B(sreg[307]), .Z(n2739) );
  NAND U3009 ( .A(n2698), .B(sreg[306]), .Z(n2702) );
  OR U3010 ( .A(n2700), .B(n2699), .Z(n2701) );
  AND U3011 ( .A(n2702), .B(n2701), .Z(n2738) );
  XOR U3012 ( .A(n2739), .B(n2738), .Z(c[307]) );
  NANDN U3013 ( .A(n2708), .B(n2707), .Z(n2712) );
  NAND U3014 ( .A(n2710), .B(n2709), .Z(n2711) );
  NAND U3015 ( .A(n2712), .B(n2711), .Z(n2773) );
  NANDN U3016 ( .A(n2714), .B(n2713), .Z(n2718) );
  NAND U3017 ( .A(n2716), .B(n2715), .Z(n2717) );
  NAND U3018 ( .A(n2718), .B(n2717), .Z(n2771) );
  XNOR U3019 ( .A(b[5]), .B(a[56]), .Z(n2746) );
  NANDN U3020 ( .A(n2746), .B(n10481), .Z(n2721) );
  NAND U3021 ( .A(n10482), .B(n2719), .Z(n2720) );
  AND U3022 ( .A(n2721), .B(n2720), .Z(n2764) );
  NANDN U3023 ( .A(n529), .B(a[52]), .Z(n2765) );
  XOR U3024 ( .A(n2764), .B(n2765), .Z(n2767) );
  NANDN U3025 ( .A(n527), .B(a[60]), .Z(n2722) );
  XOR U3026 ( .A(n10434), .B(n2722), .Z(n2724) );
  NANDN U3027 ( .A(b[0]), .B(a[59]), .Z(n2723) );
  AND U3028 ( .A(n2724), .B(n2723), .Z(n2766) );
  XNOR U3029 ( .A(n2767), .B(n2766), .Z(n2761) );
  XNOR U3030 ( .A(b[7]), .B(a[54]), .Z(n2752) );
  NANDN U3031 ( .A(n2752), .B(n10545), .Z(n2727) );
  NANDN U3032 ( .A(n2725), .B(n10546), .Z(n2726) );
  NAND U3033 ( .A(n2727), .B(n2726), .Z(n2758) );
  XNOR U3034 ( .A(b[3]), .B(a[58]), .Z(n2755) );
  NANDN U3035 ( .A(n2755), .B(n10398), .Z(n2730) );
  NANDN U3036 ( .A(n2728), .B(n10399), .Z(n2729) );
  AND U3037 ( .A(n2730), .B(n2729), .Z(n2759) );
  XNOR U3038 ( .A(n2758), .B(n2759), .Z(n2760) );
  XNOR U3039 ( .A(n2761), .B(n2760), .Z(n2770) );
  XOR U3040 ( .A(n2771), .B(n2770), .Z(n2772) );
  XNOR U3041 ( .A(n2773), .B(n2772), .Z(n2742) );
  NAND U3042 ( .A(n2732), .B(n2731), .Z(n2736) );
  NAND U3043 ( .A(n2734), .B(n2733), .Z(n2735) );
  NAND U3044 ( .A(n2736), .B(n2735), .Z(n2743) );
  XNOR U3045 ( .A(n2742), .B(n2743), .Z(n2744) );
  XNOR U3046 ( .A(n2745), .B(n2744), .Z(n2774) );
  XNOR U3047 ( .A(n2774), .B(sreg[308]), .Z(n2776) );
  NAND U3048 ( .A(n2737), .B(sreg[307]), .Z(n2741) );
  OR U3049 ( .A(n2739), .B(n2738), .Z(n2740) );
  AND U3050 ( .A(n2741), .B(n2740), .Z(n2775) );
  XOR U3051 ( .A(n2776), .B(n2775), .Z(c[308]) );
  XOR U3052 ( .A(b[5]), .B(a[57]), .Z(n2794) );
  NAND U3053 ( .A(n10481), .B(n2794), .Z(n2748) );
  NANDN U3054 ( .A(n2746), .B(n10482), .Z(n2747) );
  AND U3055 ( .A(n2748), .B(n2747), .Z(n2803) );
  NANDN U3056 ( .A(n529), .B(a[53]), .Z(n2804) );
  XOR U3057 ( .A(n2803), .B(n2804), .Z(n2806) );
  NANDN U3058 ( .A(n527), .B(a[61]), .Z(n2749) );
  XOR U3059 ( .A(n10434), .B(n2749), .Z(n2751) );
  NANDN U3060 ( .A(b[0]), .B(a[60]), .Z(n2750) );
  AND U3061 ( .A(n2751), .B(n2750), .Z(n2805) );
  XNOR U3062 ( .A(n2806), .B(n2805), .Z(n2800) );
  XNOR U3063 ( .A(b[7]), .B(a[55]), .Z(n2785) );
  NANDN U3064 ( .A(n2785), .B(n10545), .Z(n2754) );
  NANDN U3065 ( .A(n2752), .B(n10546), .Z(n2753) );
  NAND U3066 ( .A(n2754), .B(n2753), .Z(n2797) );
  XNOR U3067 ( .A(b[3]), .B(a[59]), .Z(n2788) );
  NANDN U3068 ( .A(n2788), .B(n10398), .Z(n2757) );
  NANDN U3069 ( .A(n2755), .B(n10399), .Z(n2756) );
  AND U3070 ( .A(n2757), .B(n2756), .Z(n2798) );
  XNOR U3071 ( .A(n2797), .B(n2798), .Z(n2799) );
  XNOR U3072 ( .A(n2800), .B(n2799), .Z(n2811) );
  NANDN U3073 ( .A(n2759), .B(n2758), .Z(n2763) );
  NANDN U3074 ( .A(n2761), .B(n2760), .Z(n2762) );
  NAND U3075 ( .A(n2763), .B(n2762), .Z(n2809) );
  OR U3076 ( .A(n2765), .B(n2764), .Z(n2769) );
  NAND U3077 ( .A(n2767), .B(n2766), .Z(n2768) );
  AND U3078 ( .A(n2769), .B(n2768), .Z(n2810) );
  XNOR U3079 ( .A(n2809), .B(n2810), .Z(n2812) );
  XOR U3080 ( .A(n2811), .B(n2812), .Z(n2779) );
  XOR U3081 ( .A(n2779), .B(n2780), .Z(n2781) );
  XNOR U3082 ( .A(n2782), .B(n2781), .Z(n2813) );
  XNOR U3083 ( .A(n2813), .B(sreg[309]), .Z(n2815) );
  NAND U3084 ( .A(n2774), .B(sreg[308]), .Z(n2778) );
  OR U3085 ( .A(n2776), .B(n2775), .Z(n2777) );
  AND U3086 ( .A(n2778), .B(n2777), .Z(n2814) );
  XOR U3087 ( .A(n2815), .B(n2814), .Z(c[309]) );
  OR U3088 ( .A(n2780), .B(n2779), .Z(n2784) );
  NAND U3089 ( .A(n2782), .B(n2781), .Z(n2783) );
  NAND U3090 ( .A(n2784), .B(n2783), .Z(n2821) );
  XNOR U3091 ( .A(b[7]), .B(a[56]), .Z(n2834) );
  NANDN U3092 ( .A(n2834), .B(n10545), .Z(n2787) );
  NANDN U3093 ( .A(n2785), .B(n10546), .Z(n2786) );
  NAND U3094 ( .A(n2787), .B(n2786), .Z(n2822) );
  XNOR U3095 ( .A(b[3]), .B(a[60]), .Z(n2837) );
  NANDN U3096 ( .A(n2837), .B(n10398), .Z(n2790) );
  NANDN U3097 ( .A(n2788), .B(n10399), .Z(n2789) );
  AND U3098 ( .A(n2790), .B(n2789), .Z(n2823) );
  XNOR U3099 ( .A(n2822), .B(n2823), .Z(n2824) );
  NANDN U3100 ( .A(n527), .B(a[62]), .Z(n2791) );
  XOR U3101 ( .A(n10434), .B(n2791), .Z(n2793) );
  NANDN U3102 ( .A(b[0]), .B(a[61]), .Z(n2792) );
  AND U3103 ( .A(n2793), .B(n2792), .Z(n2830) );
  XOR U3104 ( .A(b[5]), .B(a[58]), .Z(n2843) );
  NAND U3105 ( .A(n2843), .B(n10481), .Z(n2796) );
  NAND U3106 ( .A(n2794), .B(n10482), .Z(n2795) );
  NAND U3107 ( .A(n2796), .B(n2795), .Z(n2828) );
  NANDN U3108 ( .A(n529), .B(a[54]), .Z(n2829) );
  XNOR U3109 ( .A(n2828), .B(n2829), .Z(n2831) );
  XOR U3110 ( .A(n2830), .B(n2831), .Z(n2825) );
  XOR U3111 ( .A(n2824), .B(n2825), .Z(n2848) );
  NANDN U3112 ( .A(n2798), .B(n2797), .Z(n2802) );
  NANDN U3113 ( .A(n2800), .B(n2799), .Z(n2801) );
  NAND U3114 ( .A(n2802), .B(n2801), .Z(n2846) );
  OR U3115 ( .A(n2804), .B(n2803), .Z(n2808) );
  NAND U3116 ( .A(n2806), .B(n2805), .Z(n2807) );
  AND U3117 ( .A(n2808), .B(n2807), .Z(n2847) );
  XNOR U3118 ( .A(n2846), .B(n2847), .Z(n2849) );
  XNOR U3119 ( .A(n2848), .B(n2849), .Z(n2818) );
  XNOR U3120 ( .A(n2818), .B(n2819), .Z(n2820) );
  XNOR U3121 ( .A(n2821), .B(n2820), .Z(n2852) );
  XNOR U3122 ( .A(n2852), .B(sreg[310]), .Z(n2854) );
  NAND U3123 ( .A(n2813), .B(sreg[309]), .Z(n2817) );
  OR U3124 ( .A(n2815), .B(n2814), .Z(n2816) );
  AND U3125 ( .A(n2817), .B(n2816), .Z(n2853) );
  XOR U3126 ( .A(n2854), .B(n2853), .Z(c[310]) );
  NANDN U3127 ( .A(n2823), .B(n2822), .Z(n2827) );
  NAND U3128 ( .A(n2825), .B(n2824), .Z(n2826) );
  NAND U3129 ( .A(n2827), .B(n2826), .Z(n2888) );
  NANDN U3130 ( .A(n2829), .B(n2828), .Z(n2833) );
  NAND U3131 ( .A(n2831), .B(n2830), .Z(n2832) );
  NAND U3132 ( .A(n2833), .B(n2832), .Z(n2886) );
  XNOR U3133 ( .A(b[7]), .B(a[57]), .Z(n2873) );
  NANDN U3134 ( .A(n2873), .B(n10545), .Z(n2836) );
  NANDN U3135 ( .A(n2834), .B(n10546), .Z(n2835) );
  NAND U3136 ( .A(n2836), .B(n2835), .Z(n2861) );
  XNOR U3137 ( .A(b[3]), .B(a[61]), .Z(n2876) );
  NANDN U3138 ( .A(n2876), .B(n10398), .Z(n2839) );
  NANDN U3139 ( .A(n2837), .B(n10399), .Z(n2838) );
  AND U3140 ( .A(n2839), .B(n2838), .Z(n2862) );
  XNOR U3141 ( .A(n2861), .B(n2862), .Z(n2863) );
  NANDN U3142 ( .A(n527), .B(a[63]), .Z(n2840) );
  XOR U3143 ( .A(n10434), .B(n2840), .Z(n2842) );
  NANDN U3144 ( .A(b[0]), .B(a[62]), .Z(n2841) );
  AND U3145 ( .A(n2842), .B(n2841), .Z(n2869) );
  XOR U3146 ( .A(b[5]), .B(a[59]), .Z(n2882) );
  NAND U3147 ( .A(n2882), .B(n10481), .Z(n2845) );
  NAND U3148 ( .A(n2843), .B(n10482), .Z(n2844) );
  NAND U3149 ( .A(n2845), .B(n2844), .Z(n2867) );
  NANDN U3150 ( .A(n529), .B(a[55]), .Z(n2868) );
  XNOR U3151 ( .A(n2867), .B(n2868), .Z(n2870) );
  XOR U3152 ( .A(n2869), .B(n2870), .Z(n2864) );
  XOR U3153 ( .A(n2863), .B(n2864), .Z(n2885) );
  XOR U3154 ( .A(n2886), .B(n2885), .Z(n2887) );
  XNOR U3155 ( .A(n2888), .B(n2887), .Z(n2857) );
  NANDN U3156 ( .A(n2847), .B(n2846), .Z(n2851) );
  NAND U3157 ( .A(n2849), .B(n2848), .Z(n2850) );
  NAND U3158 ( .A(n2851), .B(n2850), .Z(n2858) );
  XNOR U3159 ( .A(n2857), .B(n2858), .Z(n2859) );
  XNOR U3160 ( .A(n2860), .B(n2859), .Z(n2891) );
  XNOR U3161 ( .A(n2891), .B(sreg[311]), .Z(n2893) );
  NAND U3162 ( .A(n2852), .B(sreg[310]), .Z(n2856) );
  OR U3163 ( .A(n2854), .B(n2853), .Z(n2855) );
  AND U3164 ( .A(n2856), .B(n2855), .Z(n2892) );
  XOR U3165 ( .A(n2893), .B(n2892), .Z(c[311]) );
  NANDN U3166 ( .A(n2862), .B(n2861), .Z(n2866) );
  NAND U3167 ( .A(n2864), .B(n2863), .Z(n2865) );
  NAND U3168 ( .A(n2866), .B(n2865), .Z(n2927) );
  NANDN U3169 ( .A(n2868), .B(n2867), .Z(n2872) );
  NAND U3170 ( .A(n2870), .B(n2869), .Z(n2871) );
  NAND U3171 ( .A(n2872), .B(n2871), .Z(n2925) );
  XNOR U3172 ( .A(b[7]), .B(a[58]), .Z(n2912) );
  NANDN U3173 ( .A(n2912), .B(n10545), .Z(n2875) );
  NANDN U3174 ( .A(n2873), .B(n10546), .Z(n2874) );
  NAND U3175 ( .A(n2875), .B(n2874), .Z(n2900) );
  XNOR U3176 ( .A(b[3]), .B(a[62]), .Z(n2915) );
  NANDN U3177 ( .A(n2915), .B(n10398), .Z(n2878) );
  NANDN U3178 ( .A(n2876), .B(n10399), .Z(n2877) );
  AND U3179 ( .A(n2878), .B(n2877), .Z(n2901) );
  XNOR U3180 ( .A(n2900), .B(n2901), .Z(n2902) );
  NANDN U3181 ( .A(n527), .B(a[64]), .Z(n2879) );
  XOR U3182 ( .A(n10434), .B(n2879), .Z(n2881) );
  NANDN U3183 ( .A(b[0]), .B(a[63]), .Z(n2880) );
  AND U3184 ( .A(n2881), .B(n2880), .Z(n2908) );
  XOR U3185 ( .A(b[5]), .B(a[60]), .Z(n2921) );
  NAND U3186 ( .A(n2921), .B(n10481), .Z(n2884) );
  NAND U3187 ( .A(n2882), .B(n10482), .Z(n2883) );
  NAND U3188 ( .A(n2884), .B(n2883), .Z(n2906) );
  NANDN U3189 ( .A(n529), .B(a[56]), .Z(n2907) );
  XNOR U3190 ( .A(n2906), .B(n2907), .Z(n2909) );
  XOR U3191 ( .A(n2908), .B(n2909), .Z(n2903) );
  XOR U3192 ( .A(n2902), .B(n2903), .Z(n2924) );
  XOR U3193 ( .A(n2925), .B(n2924), .Z(n2926) );
  XNOR U3194 ( .A(n2927), .B(n2926), .Z(n2896) );
  NAND U3195 ( .A(n2886), .B(n2885), .Z(n2890) );
  NAND U3196 ( .A(n2888), .B(n2887), .Z(n2889) );
  NAND U3197 ( .A(n2890), .B(n2889), .Z(n2897) );
  XNOR U3198 ( .A(n2896), .B(n2897), .Z(n2898) );
  XNOR U3199 ( .A(n2899), .B(n2898), .Z(n2930) );
  XNOR U3200 ( .A(n2930), .B(sreg[312]), .Z(n2932) );
  NAND U3201 ( .A(n2891), .B(sreg[311]), .Z(n2895) );
  OR U3202 ( .A(n2893), .B(n2892), .Z(n2894) );
  AND U3203 ( .A(n2895), .B(n2894), .Z(n2931) );
  XOR U3204 ( .A(n2932), .B(n2931), .Z(c[312]) );
  NANDN U3205 ( .A(n2901), .B(n2900), .Z(n2905) );
  NAND U3206 ( .A(n2903), .B(n2902), .Z(n2904) );
  NAND U3207 ( .A(n2905), .B(n2904), .Z(n2966) );
  NANDN U3208 ( .A(n2907), .B(n2906), .Z(n2911) );
  NAND U3209 ( .A(n2909), .B(n2908), .Z(n2910) );
  NAND U3210 ( .A(n2911), .B(n2910), .Z(n2964) );
  XNOR U3211 ( .A(b[7]), .B(a[59]), .Z(n2951) );
  NANDN U3212 ( .A(n2951), .B(n10545), .Z(n2914) );
  NANDN U3213 ( .A(n2912), .B(n10546), .Z(n2913) );
  NAND U3214 ( .A(n2914), .B(n2913), .Z(n2939) );
  XNOR U3215 ( .A(b[3]), .B(a[63]), .Z(n2954) );
  NANDN U3216 ( .A(n2954), .B(n10398), .Z(n2917) );
  NANDN U3217 ( .A(n2915), .B(n10399), .Z(n2916) );
  AND U3218 ( .A(n2917), .B(n2916), .Z(n2940) );
  XNOR U3219 ( .A(n2939), .B(n2940), .Z(n2941) );
  NANDN U3220 ( .A(n527), .B(a[65]), .Z(n2918) );
  XOR U3221 ( .A(n10434), .B(n2918), .Z(n2920) );
  NANDN U3222 ( .A(b[0]), .B(a[64]), .Z(n2919) );
  AND U3223 ( .A(n2920), .B(n2919), .Z(n2947) );
  XOR U3224 ( .A(b[5]), .B(a[61]), .Z(n2960) );
  NAND U3225 ( .A(n2960), .B(n10481), .Z(n2923) );
  NAND U3226 ( .A(n2921), .B(n10482), .Z(n2922) );
  NAND U3227 ( .A(n2923), .B(n2922), .Z(n2945) );
  NANDN U3228 ( .A(n529), .B(a[57]), .Z(n2946) );
  XNOR U3229 ( .A(n2945), .B(n2946), .Z(n2948) );
  XOR U3230 ( .A(n2947), .B(n2948), .Z(n2942) );
  XOR U3231 ( .A(n2941), .B(n2942), .Z(n2963) );
  XOR U3232 ( .A(n2964), .B(n2963), .Z(n2965) );
  XNOR U3233 ( .A(n2966), .B(n2965), .Z(n2935) );
  NAND U3234 ( .A(n2925), .B(n2924), .Z(n2929) );
  NAND U3235 ( .A(n2927), .B(n2926), .Z(n2928) );
  NAND U3236 ( .A(n2929), .B(n2928), .Z(n2936) );
  XNOR U3237 ( .A(n2935), .B(n2936), .Z(n2937) );
  XNOR U3238 ( .A(n2938), .B(n2937), .Z(n2969) );
  XNOR U3239 ( .A(n2969), .B(sreg[313]), .Z(n2971) );
  NAND U3240 ( .A(n2930), .B(sreg[312]), .Z(n2934) );
  OR U3241 ( .A(n2932), .B(n2931), .Z(n2933) );
  AND U3242 ( .A(n2934), .B(n2933), .Z(n2970) );
  XOR U3243 ( .A(n2971), .B(n2970), .Z(c[313]) );
  NANDN U3244 ( .A(n2940), .B(n2939), .Z(n2944) );
  NAND U3245 ( .A(n2942), .B(n2941), .Z(n2943) );
  NAND U3246 ( .A(n2944), .B(n2943), .Z(n3005) );
  NANDN U3247 ( .A(n2946), .B(n2945), .Z(n2950) );
  NAND U3248 ( .A(n2948), .B(n2947), .Z(n2949) );
  NAND U3249 ( .A(n2950), .B(n2949), .Z(n3003) );
  XNOR U3250 ( .A(b[7]), .B(a[60]), .Z(n2990) );
  NANDN U3251 ( .A(n2990), .B(n10545), .Z(n2953) );
  NANDN U3252 ( .A(n2951), .B(n10546), .Z(n2952) );
  NAND U3253 ( .A(n2953), .B(n2952), .Z(n2978) );
  XNOR U3254 ( .A(b[3]), .B(a[64]), .Z(n2993) );
  NANDN U3255 ( .A(n2993), .B(n10398), .Z(n2956) );
  NANDN U3256 ( .A(n2954), .B(n10399), .Z(n2955) );
  AND U3257 ( .A(n2956), .B(n2955), .Z(n2979) );
  XNOR U3258 ( .A(n2978), .B(n2979), .Z(n2980) );
  NANDN U3259 ( .A(n527), .B(a[66]), .Z(n2957) );
  XOR U3260 ( .A(n10434), .B(n2957), .Z(n2959) );
  NANDN U3261 ( .A(b[0]), .B(a[65]), .Z(n2958) );
  AND U3262 ( .A(n2959), .B(n2958), .Z(n2986) );
  XOR U3263 ( .A(b[5]), .B(a[62]), .Z(n2999) );
  NAND U3264 ( .A(n2999), .B(n10481), .Z(n2962) );
  NAND U3265 ( .A(n2960), .B(n10482), .Z(n2961) );
  NAND U3266 ( .A(n2962), .B(n2961), .Z(n2984) );
  NANDN U3267 ( .A(n529), .B(a[58]), .Z(n2985) );
  XNOR U3268 ( .A(n2984), .B(n2985), .Z(n2987) );
  XOR U3269 ( .A(n2986), .B(n2987), .Z(n2981) );
  XOR U3270 ( .A(n2980), .B(n2981), .Z(n3002) );
  XOR U3271 ( .A(n3003), .B(n3002), .Z(n3004) );
  XNOR U3272 ( .A(n3005), .B(n3004), .Z(n2974) );
  NAND U3273 ( .A(n2964), .B(n2963), .Z(n2968) );
  NAND U3274 ( .A(n2966), .B(n2965), .Z(n2967) );
  NAND U3275 ( .A(n2968), .B(n2967), .Z(n2975) );
  XNOR U3276 ( .A(n2974), .B(n2975), .Z(n2976) );
  XNOR U3277 ( .A(n2977), .B(n2976), .Z(n3008) );
  XNOR U3278 ( .A(n3008), .B(sreg[314]), .Z(n3010) );
  NAND U3279 ( .A(n2969), .B(sreg[313]), .Z(n2973) );
  OR U3280 ( .A(n2971), .B(n2970), .Z(n2972) );
  AND U3281 ( .A(n2973), .B(n2972), .Z(n3009) );
  XOR U3282 ( .A(n3010), .B(n3009), .Z(c[314]) );
  NANDN U3283 ( .A(n2979), .B(n2978), .Z(n2983) );
  NAND U3284 ( .A(n2981), .B(n2980), .Z(n2982) );
  NAND U3285 ( .A(n2983), .B(n2982), .Z(n3044) );
  NANDN U3286 ( .A(n2985), .B(n2984), .Z(n2989) );
  NAND U3287 ( .A(n2987), .B(n2986), .Z(n2988) );
  NAND U3288 ( .A(n2989), .B(n2988), .Z(n3042) );
  XNOR U3289 ( .A(b[7]), .B(a[61]), .Z(n3029) );
  NANDN U3290 ( .A(n3029), .B(n10545), .Z(n2992) );
  NANDN U3291 ( .A(n2990), .B(n10546), .Z(n2991) );
  NAND U3292 ( .A(n2992), .B(n2991), .Z(n3017) );
  XNOR U3293 ( .A(b[3]), .B(a[65]), .Z(n3032) );
  NANDN U3294 ( .A(n3032), .B(n10398), .Z(n2995) );
  NANDN U3295 ( .A(n2993), .B(n10399), .Z(n2994) );
  AND U3296 ( .A(n2995), .B(n2994), .Z(n3018) );
  XNOR U3297 ( .A(n3017), .B(n3018), .Z(n3019) );
  NANDN U3298 ( .A(n527), .B(a[67]), .Z(n2996) );
  XOR U3299 ( .A(n10434), .B(n2996), .Z(n2998) );
  NANDN U3300 ( .A(b[0]), .B(a[66]), .Z(n2997) );
  AND U3301 ( .A(n2998), .B(n2997), .Z(n3025) );
  XOR U3302 ( .A(b[5]), .B(a[63]), .Z(n3038) );
  NAND U3303 ( .A(n3038), .B(n10481), .Z(n3001) );
  NAND U3304 ( .A(n2999), .B(n10482), .Z(n3000) );
  NAND U3305 ( .A(n3001), .B(n3000), .Z(n3023) );
  NANDN U3306 ( .A(n529), .B(a[59]), .Z(n3024) );
  XNOR U3307 ( .A(n3023), .B(n3024), .Z(n3026) );
  XOR U3308 ( .A(n3025), .B(n3026), .Z(n3020) );
  XOR U3309 ( .A(n3019), .B(n3020), .Z(n3041) );
  XOR U3310 ( .A(n3042), .B(n3041), .Z(n3043) );
  XNOR U3311 ( .A(n3044), .B(n3043), .Z(n3013) );
  NAND U3312 ( .A(n3003), .B(n3002), .Z(n3007) );
  NAND U3313 ( .A(n3005), .B(n3004), .Z(n3006) );
  NAND U3314 ( .A(n3007), .B(n3006), .Z(n3014) );
  XNOR U3315 ( .A(n3013), .B(n3014), .Z(n3015) );
  XNOR U3316 ( .A(n3016), .B(n3015), .Z(n3047) );
  XNOR U3317 ( .A(n3047), .B(sreg[315]), .Z(n3049) );
  NAND U3318 ( .A(n3008), .B(sreg[314]), .Z(n3012) );
  OR U3319 ( .A(n3010), .B(n3009), .Z(n3011) );
  AND U3320 ( .A(n3012), .B(n3011), .Z(n3048) );
  XOR U3321 ( .A(n3049), .B(n3048), .Z(c[315]) );
  NANDN U3322 ( .A(n3018), .B(n3017), .Z(n3022) );
  NAND U3323 ( .A(n3020), .B(n3019), .Z(n3021) );
  NAND U3324 ( .A(n3022), .B(n3021), .Z(n3083) );
  NANDN U3325 ( .A(n3024), .B(n3023), .Z(n3028) );
  NAND U3326 ( .A(n3026), .B(n3025), .Z(n3027) );
  NAND U3327 ( .A(n3028), .B(n3027), .Z(n3081) );
  XNOR U3328 ( .A(b[7]), .B(a[62]), .Z(n3068) );
  NANDN U3329 ( .A(n3068), .B(n10545), .Z(n3031) );
  NANDN U3330 ( .A(n3029), .B(n10546), .Z(n3030) );
  NAND U3331 ( .A(n3031), .B(n3030), .Z(n3056) );
  XNOR U3332 ( .A(b[3]), .B(a[66]), .Z(n3071) );
  NANDN U3333 ( .A(n3071), .B(n10398), .Z(n3034) );
  NANDN U3334 ( .A(n3032), .B(n10399), .Z(n3033) );
  AND U3335 ( .A(n3034), .B(n3033), .Z(n3057) );
  XNOR U3336 ( .A(n3056), .B(n3057), .Z(n3058) );
  NANDN U3337 ( .A(n527), .B(a[68]), .Z(n3035) );
  XOR U3338 ( .A(n10434), .B(n3035), .Z(n3037) );
  NANDN U3339 ( .A(b[0]), .B(a[67]), .Z(n3036) );
  AND U3340 ( .A(n3037), .B(n3036), .Z(n3064) );
  XOR U3341 ( .A(b[5]), .B(a[64]), .Z(n3077) );
  NAND U3342 ( .A(n3077), .B(n10481), .Z(n3040) );
  NAND U3343 ( .A(n3038), .B(n10482), .Z(n3039) );
  NAND U3344 ( .A(n3040), .B(n3039), .Z(n3062) );
  NANDN U3345 ( .A(n529), .B(a[60]), .Z(n3063) );
  XNOR U3346 ( .A(n3062), .B(n3063), .Z(n3065) );
  XOR U3347 ( .A(n3064), .B(n3065), .Z(n3059) );
  XOR U3348 ( .A(n3058), .B(n3059), .Z(n3080) );
  XOR U3349 ( .A(n3081), .B(n3080), .Z(n3082) );
  XNOR U3350 ( .A(n3083), .B(n3082), .Z(n3052) );
  NAND U3351 ( .A(n3042), .B(n3041), .Z(n3046) );
  NAND U3352 ( .A(n3044), .B(n3043), .Z(n3045) );
  NAND U3353 ( .A(n3046), .B(n3045), .Z(n3053) );
  XNOR U3354 ( .A(n3052), .B(n3053), .Z(n3054) );
  XNOR U3355 ( .A(n3055), .B(n3054), .Z(n3086) );
  XNOR U3356 ( .A(n3086), .B(sreg[316]), .Z(n3088) );
  NAND U3357 ( .A(n3047), .B(sreg[315]), .Z(n3051) );
  OR U3358 ( .A(n3049), .B(n3048), .Z(n3050) );
  AND U3359 ( .A(n3051), .B(n3050), .Z(n3087) );
  XOR U3360 ( .A(n3088), .B(n3087), .Z(c[316]) );
  NANDN U3361 ( .A(n3057), .B(n3056), .Z(n3061) );
  NAND U3362 ( .A(n3059), .B(n3058), .Z(n3060) );
  NAND U3363 ( .A(n3061), .B(n3060), .Z(n3122) );
  NANDN U3364 ( .A(n3063), .B(n3062), .Z(n3067) );
  NAND U3365 ( .A(n3065), .B(n3064), .Z(n3066) );
  NAND U3366 ( .A(n3067), .B(n3066), .Z(n3120) );
  XNOR U3367 ( .A(b[7]), .B(a[63]), .Z(n3107) );
  NANDN U3368 ( .A(n3107), .B(n10545), .Z(n3070) );
  NANDN U3369 ( .A(n3068), .B(n10546), .Z(n3069) );
  NAND U3370 ( .A(n3070), .B(n3069), .Z(n3095) );
  XNOR U3371 ( .A(b[3]), .B(a[67]), .Z(n3110) );
  NANDN U3372 ( .A(n3110), .B(n10398), .Z(n3073) );
  NANDN U3373 ( .A(n3071), .B(n10399), .Z(n3072) );
  AND U3374 ( .A(n3073), .B(n3072), .Z(n3096) );
  XNOR U3375 ( .A(n3095), .B(n3096), .Z(n3097) );
  NANDN U3376 ( .A(n527), .B(a[69]), .Z(n3074) );
  XOR U3377 ( .A(n10434), .B(n3074), .Z(n3076) );
  NANDN U3378 ( .A(b[0]), .B(a[68]), .Z(n3075) );
  AND U3379 ( .A(n3076), .B(n3075), .Z(n3103) );
  XOR U3380 ( .A(b[5]), .B(a[65]), .Z(n3116) );
  NAND U3381 ( .A(n3116), .B(n10481), .Z(n3079) );
  NAND U3382 ( .A(n3077), .B(n10482), .Z(n3078) );
  NAND U3383 ( .A(n3079), .B(n3078), .Z(n3101) );
  NANDN U3384 ( .A(n529), .B(a[61]), .Z(n3102) );
  XNOR U3385 ( .A(n3101), .B(n3102), .Z(n3104) );
  XOR U3386 ( .A(n3103), .B(n3104), .Z(n3098) );
  XOR U3387 ( .A(n3097), .B(n3098), .Z(n3119) );
  XOR U3388 ( .A(n3120), .B(n3119), .Z(n3121) );
  XNOR U3389 ( .A(n3122), .B(n3121), .Z(n3091) );
  NAND U3390 ( .A(n3081), .B(n3080), .Z(n3085) );
  NAND U3391 ( .A(n3083), .B(n3082), .Z(n3084) );
  NAND U3392 ( .A(n3085), .B(n3084), .Z(n3092) );
  XNOR U3393 ( .A(n3091), .B(n3092), .Z(n3093) );
  XNOR U3394 ( .A(n3094), .B(n3093), .Z(n3125) );
  XNOR U3395 ( .A(n3125), .B(sreg[317]), .Z(n3127) );
  NAND U3396 ( .A(n3086), .B(sreg[316]), .Z(n3090) );
  OR U3397 ( .A(n3088), .B(n3087), .Z(n3089) );
  AND U3398 ( .A(n3090), .B(n3089), .Z(n3126) );
  XOR U3399 ( .A(n3127), .B(n3126), .Z(c[317]) );
  NANDN U3400 ( .A(n3096), .B(n3095), .Z(n3100) );
  NAND U3401 ( .A(n3098), .B(n3097), .Z(n3099) );
  NAND U3402 ( .A(n3100), .B(n3099), .Z(n3161) );
  NANDN U3403 ( .A(n3102), .B(n3101), .Z(n3106) );
  NAND U3404 ( .A(n3104), .B(n3103), .Z(n3105) );
  NAND U3405 ( .A(n3106), .B(n3105), .Z(n3159) );
  XNOR U3406 ( .A(b[7]), .B(a[64]), .Z(n3146) );
  NANDN U3407 ( .A(n3146), .B(n10545), .Z(n3109) );
  NANDN U3408 ( .A(n3107), .B(n10546), .Z(n3108) );
  NAND U3409 ( .A(n3109), .B(n3108), .Z(n3134) );
  XNOR U3410 ( .A(b[3]), .B(a[68]), .Z(n3149) );
  NANDN U3411 ( .A(n3149), .B(n10398), .Z(n3112) );
  NANDN U3412 ( .A(n3110), .B(n10399), .Z(n3111) );
  AND U3413 ( .A(n3112), .B(n3111), .Z(n3135) );
  XNOR U3414 ( .A(n3134), .B(n3135), .Z(n3136) );
  NANDN U3415 ( .A(n527), .B(a[70]), .Z(n3113) );
  XOR U3416 ( .A(n10434), .B(n3113), .Z(n3115) );
  NANDN U3417 ( .A(b[0]), .B(a[69]), .Z(n3114) );
  AND U3418 ( .A(n3115), .B(n3114), .Z(n3142) );
  XOR U3419 ( .A(b[5]), .B(a[66]), .Z(n3155) );
  NAND U3420 ( .A(n3155), .B(n10481), .Z(n3118) );
  NAND U3421 ( .A(n3116), .B(n10482), .Z(n3117) );
  NAND U3422 ( .A(n3118), .B(n3117), .Z(n3140) );
  NANDN U3423 ( .A(n529), .B(a[62]), .Z(n3141) );
  XNOR U3424 ( .A(n3140), .B(n3141), .Z(n3143) );
  XOR U3425 ( .A(n3142), .B(n3143), .Z(n3137) );
  XOR U3426 ( .A(n3136), .B(n3137), .Z(n3158) );
  XOR U3427 ( .A(n3159), .B(n3158), .Z(n3160) );
  XNOR U3428 ( .A(n3161), .B(n3160), .Z(n3130) );
  NAND U3429 ( .A(n3120), .B(n3119), .Z(n3124) );
  NAND U3430 ( .A(n3122), .B(n3121), .Z(n3123) );
  NAND U3431 ( .A(n3124), .B(n3123), .Z(n3131) );
  XNOR U3432 ( .A(n3130), .B(n3131), .Z(n3132) );
  XNOR U3433 ( .A(n3133), .B(n3132), .Z(n3164) );
  XNOR U3434 ( .A(n3164), .B(sreg[318]), .Z(n3166) );
  NAND U3435 ( .A(n3125), .B(sreg[317]), .Z(n3129) );
  OR U3436 ( .A(n3127), .B(n3126), .Z(n3128) );
  AND U3437 ( .A(n3129), .B(n3128), .Z(n3165) );
  XOR U3438 ( .A(n3166), .B(n3165), .Z(c[318]) );
  NANDN U3439 ( .A(n3135), .B(n3134), .Z(n3139) );
  NAND U3440 ( .A(n3137), .B(n3136), .Z(n3138) );
  NAND U3441 ( .A(n3139), .B(n3138), .Z(n3200) );
  NANDN U3442 ( .A(n3141), .B(n3140), .Z(n3145) );
  NAND U3443 ( .A(n3143), .B(n3142), .Z(n3144) );
  NAND U3444 ( .A(n3145), .B(n3144), .Z(n3198) );
  XNOR U3445 ( .A(b[7]), .B(a[65]), .Z(n3185) );
  NANDN U3446 ( .A(n3185), .B(n10545), .Z(n3148) );
  NANDN U3447 ( .A(n3146), .B(n10546), .Z(n3147) );
  NAND U3448 ( .A(n3148), .B(n3147), .Z(n3173) );
  XNOR U3449 ( .A(b[3]), .B(a[69]), .Z(n3188) );
  NANDN U3450 ( .A(n3188), .B(n10398), .Z(n3151) );
  NANDN U3451 ( .A(n3149), .B(n10399), .Z(n3150) );
  AND U3452 ( .A(n3151), .B(n3150), .Z(n3174) );
  XNOR U3453 ( .A(n3173), .B(n3174), .Z(n3175) );
  NANDN U3454 ( .A(n527), .B(a[71]), .Z(n3152) );
  XOR U3455 ( .A(n10434), .B(n3152), .Z(n3154) );
  NANDN U3456 ( .A(b[0]), .B(a[70]), .Z(n3153) );
  AND U3457 ( .A(n3154), .B(n3153), .Z(n3181) );
  XOR U3458 ( .A(b[5]), .B(a[67]), .Z(n3194) );
  NAND U3459 ( .A(n3194), .B(n10481), .Z(n3157) );
  NAND U3460 ( .A(n3155), .B(n10482), .Z(n3156) );
  NAND U3461 ( .A(n3157), .B(n3156), .Z(n3179) );
  NANDN U3462 ( .A(n529), .B(a[63]), .Z(n3180) );
  XNOR U3463 ( .A(n3179), .B(n3180), .Z(n3182) );
  XOR U3464 ( .A(n3181), .B(n3182), .Z(n3176) );
  XOR U3465 ( .A(n3175), .B(n3176), .Z(n3197) );
  XOR U3466 ( .A(n3198), .B(n3197), .Z(n3199) );
  XNOR U3467 ( .A(n3200), .B(n3199), .Z(n3169) );
  NAND U3468 ( .A(n3159), .B(n3158), .Z(n3163) );
  NAND U3469 ( .A(n3161), .B(n3160), .Z(n3162) );
  NAND U3470 ( .A(n3163), .B(n3162), .Z(n3170) );
  XNOR U3471 ( .A(n3169), .B(n3170), .Z(n3171) );
  XNOR U3472 ( .A(n3172), .B(n3171), .Z(n3203) );
  XNOR U3473 ( .A(n3203), .B(sreg[319]), .Z(n3205) );
  NAND U3474 ( .A(n3164), .B(sreg[318]), .Z(n3168) );
  OR U3475 ( .A(n3166), .B(n3165), .Z(n3167) );
  AND U3476 ( .A(n3168), .B(n3167), .Z(n3204) );
  XOR U3477 ( .A(n3205), .B(n3204), .Z(c[319]) );
  NANDN U3478 ( .A(n3174), .B(n3173), .Z(n3178) );
  NAND U3479 ( .A(n3176), .B(n3175), .Z(n3177) );
  NAND U3480 ( .A(n3178), .B(n3177), .Z(n3239) );
  NANDN U3481 ( .A(n3180), .B(n3179), .Z(n3184) );
  NAND U3482 ( .A(n3182), .B(n3181), .Z(n3183) );
  NAND U3483 ( .A(n3184), .B(n3183), .Z(n3237) );
  XNOR U3484 ( .A(b[7]), .B(a[66]), .Z(n3224) );
  NANDN U3485 ( .A(n3224), .B(n10545), .Z(n3187) );
  NANDN U3486 ( .A(n3185), .B(n10546), .Z(n3186) );
  NAND U3487 ( .A(n3187), .B(n3186), .Z(n3212) );
  XNOR U3488 ( .A(b[3]), .B(a[70]), .Z(n3227) );
  NANDN U3489 ( .A(n3227), .B(n10398), .Z(n3190) );
  NANDN U3490 ( .A(n3188), .B(n10399), .Z(n3189) );
  AND U3491 ( .A(n3190), .B(n3189), .Z(n3213) );
  XNOR U3492 ( .A(n3212), .B(n3213), .Z(n3214) );
  NANDN U3493 ( .A(n527), .B(a[72]), .Z(n3191) );
  XOR U3494 ( .A(n10434), .B(n3191), .Z(n3193) );
  NANDN U3495 ( .A(b[0]), .B(a[71]), .Z(n3192) );
  AND U3496 ( .A(n3193), .B(n3192), .Z(n3220) );
  XOR U3497 ( .A(b[5]), .B(a[68]), .Z(n3233) );
  NAND U3498 ( .A(n3233), .B(n10481), .Z(n3196) );
  NAND U3499 ( .A(n3194), .B(n10482), .Z(n3195) );
  NAND U3500 ( .A(n3196), .B(n3195), .Z(n3218) );
  NANDN U3501 ( .A(n529), .B(a[64]), .Z(n3219) );
  XNOR U3502 ( .A(n3218), .B(n3219), .Z(n3221) );
  XOR U3503 ( .A(n3220), .B(n3221), .Z(n3215) );
  XOR U3504 ( .A(n3214), .B(n3215), .Z(n3236) );
  XOR U3505 ( .A(n3237), .B(n3236), .Z(n3238) );
  XNOR U3506 ( .A(n3239), .B(n3238), .Z(n3208) );
  NAND U3507 ( .A(n3198), .B(n3197), .Z(n3202) );
  NAND U3508 ( .A(n3200), .B(n3199), .Z(n3201) );
  NAND U3509 ( .A(n3202), .B(n3201), .Z(n3209) );
  XNOR U3510 ( .A(n3208), .B(n3209), .Z(n3210) );
  XNOR U3511 ( .A(n3211), .B(n3210), .Z(n3242) );
  XNOR U3512 ( .A(n3242), .B(sreg[320]), .Z(n3244) );
  NAND U3513 ( .A(n3203), .B(sreg[319]), .Z(n3207) );
  OR U3514 ( .A(n3205), .B(n3204), .Z(n3206) );
  AND U3515 ( .A(n3207), .B(n3206), .Z(n3243) );
  XOR U3516 ( .A(n3244), .B(n3243), .Z(c[320]) );
  NANDN U3517 ( .A(n3213), .B(n3212), .Z(n3217) );
  NAND U3518 ( .A(n3215), .B(n3214), .Z(n3216) );
  NAND U3519 ( .A(n3217), .B(n3216), .Z(n3278) );
  NANDN U3520 ( .A(n3219), .B(n3218), .Z(n3223) );
  NAND U3521 ( .A(n3221), .B(n3220), .Z(n3222) );
  NAND U3522 ( .A(n3223), .B(n3222), .Z(n3276) );
  XNOR U3523 ( .A(b[7]), .B(a[67]), .Z(n3263) );
  NANDN U3524 ( .A(n3263), .B(n10545), .Z(n3226) );
  NANDN U3525 ( .A(n3224), .B(n10546), .Z(n3225) );
  NAND U3526 ( .A(n3226), .B(n3225), .Z(n3251) );
  XNOR U3527 ( .A(b[3]), .B(a[71]), .Z(n3266) );
  NANDN U3528 ( .A(n3266), .B(n10398), .Z(n3229) );
  NANDN U3529 ( .A(n3227), .B(n10399), .Z(n3228) );
  AND U3530 ( .A(n3229), .B(n3228), .Z(n3252) );
  XNOR U3531 ( .A(n3251), .B(n3252), .Z(n3253) );
  NANDN U3532 ( .A(n527), .B(a[73]), .Z(n3230) );
  XOR U3533 ( .A(n10434), .B(n3230), .Z(n3232) );
  NANDN U3534 ( .A(b[0]), .B(a[72]), .Z(n3231) );
  AND U3535 ( .A(n3232), .B(n3231), .Z(n3259) );
  XOR U3536 ( .A(b[5]), .B(a[69]), .Z(n3272) );
  NAND U3537 ( .A(n3272), .B(n10481), .Z(n3235) );
  NAND U3538 ( .A(n3233), .B(n10482), .Z(n3234) );
  NAND U3539 ( .A(n3235), .B(n3234), .Z(n3257) );
  NANDN U3540 ( .A(n529), .B(a[65]), .Z(n3258) );
  XNOR U3541 ( .A(n3257), .B(n3258), .Z(n3260) );
  XOR U3542 ( .A(n3259), .B(n3260), .Z(n3254) );
  XOR U3543 ( .A(n3253), .B(n3254), .Z(n3275) );
  XOR U3544 ( .A(n3276), .B(n3275), .Z(n3277) );
  XNOR U3545 ( .A(n3278), .B(n3277), .Z(n3247) );
  NAND U3546 ( .A(n3237), .B(n3236), .Z(n3241) );
  NAND U3547 ( .A(n3239), .B(n3238), .Z(n3240) );
  NAND U3548 ( .A(n3241), .B(n3240), .Z(n3248) );
  XNOR U3549 ( .A(n3247), .B(n3248), .Z(n3249) );
  XNOR U3550 ( .A(n3250), .B(n3249), .Z(n3281) );
  XNOR U3551 ( .A(n3281), .B(sreg[321]), .Z(n3283) );
  NAND U3552 ( .A(n3242), .B(sreg[320]), .Z(n3246) );
  OR U3553 ( .A(n3244), .B(n3243), .Z(n3245) );
  AND U3554 ( .A(n3246), .B(n3245), .Z(n3282) );
  XOR U3555 ( .A(n3283), .B(n3282), .Z(c[321]) );
  NANDN U3556 ( .A(n3252), .B(n3251), .Z(n3256) );
  NAND U3557 ( .A(n3254), .B(n3253), .Z(n3255) );
  NAND U3558 ( .A(n3256), .B(n3255), .Z(n3317) );
  NANDN U3559 ( .A(n3258), .B(n3257), .Z(n3262) );
  NAND U3560 ( .A(n3260), .B(n3259), .Z(n3261) );
  NAND U3561 ( .A(n3262), .B(n3261), .Z(n3315) );
  XNOR U3562 ( .A(b[7]), .B(a[68]), .Z(n3302) );
  NANDN U3563 ( .A(n3302), .B(n10545), .Z(n3265) );
  NANDN U3564 ( .A(n3263), .B(n10546), .Z(n3264) );
  NAND U3565 ( .A(n3265), .B(n3264), .Z(n3290) );
  XNOR U3566 ( .A(b[3]), .B(a[72]), .Z(n3305) );
  NANDN U3567 ( .A(n3305), .B(n10398), .Z(n3268) );
  NANDN U3568 ( .A(n3266), .B(n10399), .Z(n3267) );
  AND U3569 ( .A(n3268), .B(n3267), .Z(n3291) );
  XNOR U3570 ( .A(n3290), .B(n3291), .Z(n3292) );
  NANDN U3571 ( .A(n527), .B(a[74]), .Z(n3269) );
  XOR U3572 ( .A(n10434), .B(n3269), .Z(n3271) );
  NANDN U3573 ( .A(b[0]), .B(a[73]), .Z(n3270) );
  AND U3574 ( .A(n3271), .B(n3270), .Z(n3298) );
  XOR U3575 ( .A(b[5]), .B(a[70]), .Z(n3311) );
  NAND U3576 ( .A(n3311), .B(n10481), .Z(n3274) );
  NAND U3577 ( .A(n3272), .B(n10482), .Z(n3273) );
  NAND U3578 ( .A(n3274), .B(n3273), .Z(n3296) );
  NANDN U3579 ( .A(n529), .B(a[66]), .Z(n3297) );
  XNOR U3580 ( .A(n3296), .B(n3297), .Z(n3299) );
  XOR U3581 ( .A(n3298), .B(n3299), .Z(n3293) );
  XOR U3582 ( .A(n3292), .B(n3293), .Z(n3314) );
  XOR U3583 ( .A(n3315), .B(n3314), .Z(n3316) );
  XNOR U3584 ( .A(n3317), .B(n3316), .Z(n3286) );
  NAND U3585 ( .A(n3276), .B(n3275), .Z(n3280) );
  NAND U3586 ( .A(n3278), .B(n3277), .Z(n3279) );
  NAND U3587 ( .A(n3280), .B(n3279), .Z(n3287) );
  XNOR U3588 ( .A(n3286), .B(n3287), .Z(n3288) );
  XNOR U3589 ( .A(n3289), .B(n3288), .Z(n3320) );
  XNOR U3590 ( .A(n3320), .B(sreg[322]), .Z(n3322) );
  NAND U3591 ( .A(n3281), .B(sreg[321]), .Z(n3285) );
  OR U3592 ( .A(n3283), .B(n3282), .Z(n3284) );
  AND U3593 ( .A(n3285), .B(n3284), .Z(n3321) );
  XOR U3594 ( .A(n3322), .B(n3321), .Z(c[322]) );
  NANDN U3595 ( .A(n3291), .B(n3290), .Z(n3295) );
  NAND U3596 ( .A(n3293), .B(n3292), .Z(n3294) );
  NAND U3597 ( .A(n3295), .B(n3294), .Z(n3356) );
  NANDN U3598 ( .A(n3297), .B(n3296), .Z(n3301) );
  NAND U3599 ( .A(n3299), .B(n3298), .Z(n3300) );
  NAND U3600 ( .A(n3301), .B(n3300), .Z(n3354) );
  XNOR U3601 ( .A(b[7]), .B(a[69]), .Z(n3341) );
  NANDN U3602 ( .A(n3341), .B(n10545), .Z(n3304) );
  NANDN U3603 ( .A(n3302), .B(n10546), .Z(n3303) );
  NAND U3604 ( .A(n3304), .B(n3303), .Z(n3329) );
  XNOR U3605 ( .A(b[3]), .B(a[73]), .Z(n3344) );
  NANDN U3606 ( .A(n3344), .B(n10398), .Z(n3307) );
  NANDN U3607 ( .A(n3305), .B(n10399), .Z(n3306) );
  AND U3608 ( .A(n3307), .B(n3306), .Z(n3330) );
  XNOR U3609 ( .A(n3329), .B(n3330), .Z(n3331) );
  NANDN U3610 ( .A(n527), .B(a[75]), .Z(n3308) );
  XOR U3611 ( .A(n10434), .B(n3308), .Z(n3310) );
  NANDN U3612 ( .A(b[0]), .B(a[74]), .Z(n3309) );
  AND U3613 ( .A(n3310), .B(n3309), .Z(n3337) );
  XOR U3614 ( .A(b[5]), .B(a[71]), .Z(n3350) );
  NAND U3615 ( .A(n3350), .B(n10481), .Z(n3313) );
  NAND U3616 ( .A(n3311), .B(n10482), .Z(n3312) );
  NAND U3617 ( .A(n3313), .B(n3312), .Z(n3335) );
  NANDN U3618 ( .A(n529), .B(a[67]), .Z(n3336) );
  XNOR U3619 ( .A(n3335), .B(n3336), .Z(n3338) );
  XOR U3620 ( .A(n3337), .B(n3338), .Z(n3332) );
  XOR U3621 ( .A(n3331), .B(n3332), .Z(n3353) );
  XOR U3622 ( .A(n3354), .B(n3353), .Z(n3355) );
  XNOR U3623 ( .A(n3356), .B(n3355), .Z(n3325) );
  NAND U3624 ( .A(n3315), .B(n3314), .Z(n3319) );
  NAND U3625 ( .A(n3317), .B(n3316), .Z(n3318) );
  NAND U3626 ( .A(n3319), .B(n3318), .Z(n3326) );
  XNOR U3627 ( .A(n3325), .B(n3326), .Z(n3327) );
  XNOR U3628 ( .A(n3328), .B(n3327), .Z(n3359) );
  XNOR U3629 ( .A(n3359), .B(sreg[323]), .Z(n3361) );
  NAND U3630 ( .A(n3320), .B(sreg[322]), .Z(n3324) );
  OR U3631 ( .A(n3322), .B(n3321), .Z(n3323) );
  AND U3632 ( .A(n3324), .B(n3323), .Z(n3360) );
  XOR U3633 ( .A(n3361), .B(n3360), .Z(c[323]) );
  NANDN U3634 ( .A(n3330), .B(n3329), .Z(n3334) );
  NAND U3635 ( .A(n3332), .B(n3331), .Z(n3333) );
  NAND U3636 ( .A(n3334), .B(n3333), .Z(n3395) );
  NANDN U3637 ( .A(n3336), .B(n3335), .Z(n3340) );
  NAND U3638 ( .A(n3338), .B(n3337), .Z(n3339) );
  NAND U3639 ( .A(n3340), .B(n3339), .Z(n3393) );
  XNOR U3640 ( .A(b[7]), .B(a[70]), .Z(n3380) );
  NANDN U3641 ( .A(n3380), .B(n10545), .Z(n3343) );
  NANDN U3642 ( .A(n3341), .B(n10546), .Z(n3342) );
  NAND U3643 ( .A(n3343), .B(n3342), .Z(n3368) );
  XNOR U3644 ( .A(b[3]), .B(a[74]), .Z(n3383) );
  NANDN U3645 ( .A(n3383), .B(n10398), .Z(n3346) );
  NANDN U3646 ( .A(n3344), .B(n10399), .Z(n3345) );
  AND U3647 ( .A(n3346), .B(n3345), .Z(n3369) );
  XNOR U3648 ( .A(n3368), .B(n3369), .Z(n3370) );
  NANDN U3649 ( .A(n527), .B(a[76]), .Z(n3347) );
  XOR U3650 ( .A(n10434), .B(n3347), .Z(n3349) );
  NANDN U3651 ( .A(b[0]), .B(a[75]), .Z(n3348) );
  AND U3652 ( .A(n3349), .B(n3348), .Z(n3376) );
  XOR U3653 ( .A(b[5]), .B(a[72]), .Z(n3389) );
  NAND U3654 ( .A(n3389), .B(n10481), .Z(n3352) );
  NAND U3655 ( .A(n3350), .B(n10482), .Z(n3351) );
  NAND U3656 ( .A(n3352), .B(n3351), .Z(n3374) );
  NANDN U3657 ( .A(n529), .B(a[68]), .Z(n3375) );
  XNOR U3658 ( .A(n3374), .B(n3375), .Z(n3377) );
  XOR U3659 ( .A(n3376), .B(n3377), .Z(n3371) );
  XOR U3660 ( .A(n3370), .B(n3371), .Z(n3392) );
  XOR U3661 ( .A(n3393), .B(n3392), .Z(n3394) );
  XNOR U3662 ( .A(n3395), .B(n3394), .Z(n3364) );
  NAND U3663 ( .A(n3354), .B(n3353), .Z(n3358) );
  NAND U3664 ( .A(n3356), .B(n3355), .Z(n3357) );
  NAND U3665 ( .A(n3358), .B(n3357), .Z(n3365) );
  XNOR U3666 ( .A(n3364), .B(n3365), .Z(n3366) );
  XNOR U3667 ( .A(n3367), .B(n3366), .Z(n3398) );
  XNOR U3668 ( .A(n3398), .B(sreg[324]), .Z(n3400) );
  NAND U3669 ( .A(n3359), .B(sreg[323]), .Z(n3363) );
  OR U3670 ( .A(n3361), .B(n3360), .Z(n3362) );
  AND U3671 ( .A(n3363), .B(n3362), .Z(n3399) );
  XOR U3672 ( .A(n3400), .B(n3399), .Z(c[324]) );
  NANDN U3673 ( .A(n3369), .B(n3368), .Z(n3373) );
  NAND U3674 ( .A(n3371), .B(n3370), .Z(n3372) );
  NAND U3675 ( .A(n3373), .B(n3372), .Z(n3434) );
  NANDN U3676 ( .A(n3375), .B(n3374), .Z(n3379) );
  NAND U3677 ( .A(n3377), .B(n3376), .Z(n3378) );
  NAND U3678 ( .A(n3379), .B(n3378), .Z(n3432) );
  XNOR U3679 ( .A(b[7]), .B(a[71]), .Z(n3419) );
  NANDN U3680 ( .A(n3419), .B(n10545), .Z(n3382) );
  NANDN U3681 ( .A(n3380), .B(n10546), .Z(n3381) );
  NAND U3682 ( .A(n3382), .B(n3381), .Z(n3407) );
  XNOR U3683 ( .A(b[3]), .B(a[75]), .Z(n3422) );
  NANDN U3684 ( .A(n3422), .B(n10398), .Z(n3385) );
  NANDN U3685 ( .A(n3383), .B(n10399), .Z(n3384) );
  AND U3686 ( .A(n3385), .B(n3384), .Z(n3408) );
  XNOR U3687 ( .A(n3407), .B(n3408), .Z(n3409) );
  NANDN U3688 ( .A(n527), .B(a[77]), .Z(n3386) );
  XOR U3689 ( .A(n10434), .B(n3386), .Z(n3388) );
  NANDN U3690 ( .A(b[0]), .B(a[76]), .Z(n3387) );
  AND U3691 ( .A(n3388), .B(n3387), .Z(n3415) );
  XOR U3692 ( .A(b[5]), .B(a[73]), .Z(n3428) );
  NAND U3693 ( .A(n3428), .B(n10481), .Z(n3391) );
  NAND U3694 ( .A(n3389), .B(n10482), .Z(n3390) );
  NAND U3695 ( .A(n3391), .B(n3390), .Z(n3413) );
  NANDN U3696 ( .A(n529), .B(a[69]), .Z(n3414) );
  XNOR U3697 ( .A(n3413), .B(n3414), .Z(n3416) );
  XOR U3698 ( .A(n3415), .B(n3416), .Z(n3410) );
  XOR U3699 ( .A(n3409), .B(n3410), .Z(n3431) );
  XOR U3700 ( .A(n3432), .B(n3431), .Z(n3433) );
  XNOR U3701 ( .A(n3434), .B(n3433), .Z(n3403) );
  NAND U3702 ( .A(n3393), .B(n3392), .Z(n3397) );
  NAND U3703 ( .A(n3395), .B(n3394), .Z(n3396) );
  NAND U3704 ( .A(n3397), .B(n3396), .Z(n3404) );
  XNOR U3705 ( .A(n3403), .B(n3404), .Z(n3405) );
  XNOR U3706 ( .A(n3406), .B(n3405), .Z(n3437) );
  XNOR U3707 ( .A(n3437), .B(sreg[325]), .Z(n3439) );
  NAND U3708 ( .A(n3398), .B(sreg[324]), .Z(n3402) );
  OR U3709 ( .A(n3400), .B(n3399), .Z(n3401) );
  AND U3710 ( .A(n3402), .B(n3401), .Z(n3438) );
  XOR U3711 ( .A(n3439), .B(n3438), .Z(c[325]) );
  NANDN U3712 ( .A(n3408), .B(n3407), .Z(n3412) );
  NAND U3713 ( .A(n3410), .B(n3409), .Z(n3411) );
  NAND U3714 ( .A(n3412), .B(n3411), .Z(n3473) );
  NANDN U3715 ( .A(n3414), .B(n3413), .Z(n3418) );
  NAND U3716 ( .A(n3416), .B(n3415), .Z(n3417) );
  NAND U3717 ( .A(n3418), .B(n3417), .Z(n3471) );
  XNOR U3718 ( .A(b[7]), .B(a[72]), .Z(n3458) );
  NANDN U3719 ( .A(n3458), .B(n10545), .Z(n3421) );
  NANDN U3720 ( .A(n3419), .B(n10546), .Z(n3420) );
  NAND U3721 ( .A(n3421), .B(n3420), .Z(n3446) );
  XNOR U3722 ( .A(b[3]), .B(a[76]), .Z(n3461) );
  NANDN U3723 ( .A(n3461), .B(n10398), .Z(n3424) );
  NANDN U3724 ( .A(n3422), .B(n10399), .Z(n3423) );
  AND U3725 ( .A(n3424), .B(n3423), .Z(n3447) );
  XNOR U3726 ( .A(n3446), .B(n3447), .Z(n3448) );
  NANDN U3727 ( .A(n527), .B(a[78]), .Z(n3425) );
  XOR U3728 ( .A(n10434), .B(n3425), .Z(n3427) );
  NANDN U3729 ( .A(b[0]), .B(a[77]), .Z(n3426) );
  AND U3730 ( .A(n3427), .B(n3426), .Z(n3454) );
  XOR U3731 ( .A(b[5]), .B(a[74]), .Z(n3467) );
  NAND U3732 ( .A(n3467), .B(n10481), .Z(n3430) );
  NAND U3733 ( .A(n3428), .B(n10482), .Z(n3429) );
  NAND U3734 ( .A(n3430), .B(n3429), .Z(n3452) );
  NANDN U3735 ( .A(n529), .B(a[70]), .Z(n3453) );
  XNOR U3736 ( .A(n3452), .B(n3453), .Z(n3455) );
  XOR U3737 ( .A(n3454), .B(n3455), .Z(n3449) );
  XOR U3738 ( .A(n3448), .B(n3449), .Z(n3470) );
  XOR U3739 ( .A(n3471), .B(n3470), .Z(n3472) );
  XNOR U3740 ( .A(n3473), .B(n3472), .Z(n3442) );
  NAND U3741 ( .A(n3432), .B(n3431), .Z(n3436) );
  NAND U3742 ( .A(n3434), .B(n3433), .Z(n3435) );
  NAND U3743 ( .A(n3436), .B(n3435), .Z(n3443) );
  XNOR U3744 ( .A(n3442), .B(n3443), .Z(n3444) );
  XNOR U3745 ( .A(n3445), .B(n3444), .Z(n3476) );
  XNOR U3746 ( .A(n3476), .B(sreg[326]), .Z(n3478) );
  NAND U3747 ( .A(n3437), .B(sreg[325]), .Z(n3441) );
  OR U3748 ( .A(n3439), .B(n3438), .Z(n3440) );
  AND U3749 ( .A(n3441), .B(n3440), .Z(n3477) );
  XOR U3750 ( .A(n3478), .B(n3477), .Z(c[326]) );
  NANDN U3751 ( .A(n3447), .B(n3446), .Z(n3451) );
  NAND U3752 ( .A(n3449), .B(n3448), .Z(n3450) );
  NAND U3753 ( .A(n3451), .B(n3450), .Z(n3512) );
  NANDN U3754 ( .A(n3453), .B(n3452), .Z(n3457) );
  NAND U3755 ( .A(n3455), .B(n3454), .Z(n3456) );
  NAND U3756 ( .A(n3457), .B(n3456), .Z(n3510) );
  XNOR U3757 ( .A(b[7]), .B(a[73]), .Z(n3497) );
  NANDN U3758 ( .A(n3497), .B(n10545), .Z(n3460) );
  NANDN U3759 ( .A(n3458), .B(n10546), .Z(n3459) );
  NAND U3760 ( .A(n3460), .B(n3459), .Z(n3485) );
  XNOR U3761 ( .A(b[3]), .B(a[77]), .Z(n3500) );
  NANDN U3762 ( .A(n3500), .B(n10398), .Z(n3463) );
  NANDN U3763 ( .A(n3461), .B(n10399), .Z(n3462) );
  AND U3764 ( .A(n3463), .B(n3462), .Z(n3486) );
  XNOR U3765 ( .A(n3485), .B(n3486), .Z(n3487) );
  NANDN U3766 ( .A(n527), .B(a[79]), .Z(n3464) );
  XOR U3767 ( .A(n10434), .B(n3464), .Z(n3466) );
  NANDN U3768 ( .A(b[0]), .B(a[78]), .Z(n3465) );
  AND U3769 ( .A(n3466), .B(n3465), .Z(n3493) );
  XOR U3770 ( .A(b[5]), .B(a[75]), .Z(n3506) );
  NAND U3771 ( .A(n3506), .B(n10481), .Z(n3469) );
  NAND U3772 ( .A(n3467), .B(n10482), .Z(n3468) );
  NAND U3773 ( .A(n3469), .B(n3468), .Z(n3491) );
  NANDN U3774 ( .A(n529), .B(a[71]), .Z(n3492) );
  XNOR U3775 ( .A(n3491), .B(n3492), .Z(n3494) );
  XOR U3776 ( .A(n3493), .B(n3494), .Z(n3488) );
  XOR U3777 ( .A(n3487), .B(n3488), .Z(n3509) );
  XOR U3778 ( .A(n3510), .B(n3509), .Z(n3511) );
  XNOR U3779 ( .A(n3512), .B(n3511), .Z(n3481) );
  NAND U3780 ( .A(n3471), .B(n3470), .Z(n3475) );
  NAND U3781 ( .A(n3473), .B(n3472), .Z(n3474) );
  NAND U3782 ( .A(n3475), .B(n3474), .Z(n3482) );
  XNOR U3783 ( .A(n3481), .B(n3482), .Z(n3483) );
  XNOR U3784 ( .A(n3484), .B(n3483), .Z(n3515) );
  XNOR U3785 ( .A(n3515), .B(sreg[327]), .Z(n3517) );
  NAND U3786 ( .A(n3476), .B(sreg[326]), .Z(n3480) );
  OR U3787 ( .A(n3478), .B(n3477), .Z(n3479) );
  AND U3788 ( .A(n3480), .B(n3479), .Z(n3516) );
  XOR U3789 ( .A(n3517), .B(n3516), .Z(c[327]) );
  NANDN U3790 ( .A(n3486), .B(n3485), .Z(n3490) );
  NAND U3791 ( .A(n3488), .B(n3487), .Z(n3489) );
  NAND U3792 ( .A(n3490), .B(n3489), .Z(n3551) );
  NANDN U3793 ( .A(n3492), .B(n3491), .Z(n3496) );
  NAND U3794 ( .A(n3494), .B(n3493), .Z(n3495) );
  NAND U3795 ( .A(n3496), .B(n3495), .Z(n3549) );
  XNOR U3796 ( .A(b[7]), .B(a[74]), .Z(n3536) );
  NANDN U3797 ( .A(n3536), .B(n10545), .Z(n3499) );
  NANDN U3798 ( .A(n3497), .B(n10546), .Z(n3498) );
  NAND U3799 ( .A(n3499), .B(n3498), .Z(n3524) );
  XNOR U3800 ( .A(b[3]), .B(a[78]), .Z(n3539) );
  NANDN U3801 ( .A(n3539), .B(n10398), .Z(n3502) );
  NANDN U3802 ( .A(n3500), .B(n10399), .Z(n3501) );
  AND U3803 ( .A(n3502), .B(n3501), .Z(n3525) );
  XNOR U3804 ( .A(n3524), .B(n3525), .Z(n3526) );
  NANDN U3805 ( .A(n527), .B(a[80]), .Z(n3503) );
  XOR U3806 ( .A(n10434), .B(n3503), .Z(n3505) );
  NANDN U3807 ( .A(b[0]), .B(a[79]), .Z(n3504) );
  AND U3808 ( .A(n3505), .B(n3504), .Z(n3532) );
  XOR U3809 ( .A(b[5]), .B(a[76]), .Z(n3545) );
  NAND U3810 ( .A(n3545), .B(n10481), .Z(n3508) );
  NAND U3811 ( .A(n3506), .B(n10482), .Z(n3507) );
  NAND U3812 ( .A(n3508), .B(n3507), .Z(n3530) );
  NANDN U3813 ( .A(n529), .B(a[72]), .Z(n3531) );
  XNOR U3814 ( .A(n3530), .B(n3531), .Z(n3533) );
  XOR U3815 ( .A(n3532), .B(n3533), .Z(n3527) );
  XOR U3816 ( .A(n3526), .B(n3527), .Z(n3548) );
  XOR U3817 ( .A(n3549), .B(n3548), .Z(n3550) );
  XNOR U3818 ( .A(n3551), .B(n3550), .Z(n3520) );
  NAND U3819 ( .A(n3510), .B(n3509), .Z(n3514) );
  NAND U3820 ( .A(n3512), .B(n3511), .Z(n3513) );
  NAND U3821 ( .A(n3514), .B(n3513), .Z(n3521) );
  XNOR U3822 ( .A(n3520), .B(n3521), .Z(n3522) );
  XNOR U3823 ( .A(n3523), .B(n3522), .Z(n3554) );
  XNOR U3824 ( .A(n3554), .B(sreg[328]), .Z(n3556) );
  NAND U3825 ( .A(n3515), .B(sreg[327]), .Z(n3519) );
  OR U3826 ( .A(n3517), .B(n3516), .Z(n3518) );
  AND U3827 ( .A(n3519), .B(n3518), .Z(n3555) );
  XOR U3828 ( .A(n3556), .B(n3555), .Z(c[328]) );
  NANDN U3829 ( .A(n3525), .B(n3524), .Z(n3529) );
  NAND U3830 ( .A(n3527), .B(n3526), .Z(n3528) );
  NAND U3831 ( .A(n3529), .B(n3528), .Z(n3590) );
  NANDN U3832 ( .A(n3531), .B(n3530), .Z(n3535) );
  NAND U3833 ( .A(n3533), .B(n3532), .Z(n3534) );
  NAND U3834 ( .A(n3535), .B(n3534), .Z(n3588) );
  XNOR U3835 ( .A(b[7]), .B(a[75]), .Z(n3575) );
  NANDN U3836 ( .A(n3575), .B(n10545), .Z(n3538) );
  NANDN U3837 ( .A(n3536), .B(n10546), .Z(n3537) );
  NAND U3838 ( .A(n3538), .B(n3537), .Z(n3563) );
  XNOR U3839 ( .A(b[3]), .B(a[79]), .Z(n3578) );
  NANDN U3840 ( .A(n3578), .B(n10398), .Z(n3541) );
  NANDN U3841 ( .A(n3539), .B(n10399), .Z(n3540) );
  AND U3842 ( .A(n3541), .B(n3540), .Z(n3564) );
  XNOR U3843 ( .A(n3563), .B(n3564), .Z(n3565) );
  NANDN U3844 ( .A(n527), .B(a[81]), .Z(n3542) );
  XOR U3845 ( .A(n10434), .B(n3542), .Z(n3544) );
  NANDN U3846 ( .A(b[0]), .B(a[80]), .Z(n3543) );
  AND U3847 ( .A(n3544), .B(n3543), .Z(n3571) );
  XOR U3848 ( .A(b[5]), .B(a[77]), .Z(n3584) );
  NAND U3849 ( .A(n3584), .B(n10481), .Z(n3547) );
  NAND U3850 ( .A(n3545), .B(n10482), .Z(n3546) );
  NAND U3851 ( .A(n3547), .B(n3546), .Z(n3569) );
  NANDN U3852 ( .A(n529), .B(a[73]), .Z(n3570) );
  XNOR U3853 ( .A(n3569), .B(n3570), .Z(n3572) );
  XOR U3854 ( .A(n3571), .B(n3572), .Z(n3566) );
  XOR U3855 ( .A(n3565), .B(n3566), .Z(n3587) );
  XOR U3856 ( .A(n3588), .B(n3587), .Z(n3589) );
  XNOR U3857 ( .A(n3590), .B(n3589), .Z(n3559) );
  NAND U3858 ( .A(n3549), .B(n3548), .Z(n3553) );
  NAND U3859 ( .A(n3551), .B(n3550), .Z(n3552) );
  NAND U3860 ( .A(n3553), .B(n3552), .Z(n3560) );
  XNOR U3861 ( .A(n3559), .B(n3560), .Z(n3561) );
  XNOR U3862 ( .A(n3562), .B(n3561), .Z(n3593) );
  XNOR U3863 ( .A(n3593), .B(sreg[329]), .Z(n3595) );
  NAND U3864 ( .A(n3554), .B(sreg[328]), .Z(n3558) );
  OR U3865 ( .A(n3556), .B(n3555), .Z(n3557) );
  AND U3866 ( .A(n3558), .B(n3557), .Z(n3594) );
  XOR U3867 ( .A(n3595), .B(n3594), .Z(c[329]) );
  NANDN U3868 ( .A(n3564), .B(n3563), .Z(n3568) );
  NAND U3869 ( .A(n3566), .B(n3565), .Z(n3567) );
  NAND U3870 ( .A(n3568), .B(n3567), .Z(n3629) );
  NANDN U3871 ( .A(n3570), .B(n3569), .Z(n3574) );
  NAND U3872 ( .A(n3572), .B(n3571), .Z(n3573) );
  NAND U3873 ( .A(n3574), .B(n3573), .Z(n3627) );
  XNOR U3874 ( .A(b[7]), .B(a[76]), .Z(n3614) );
  NANDN U3875 ( .A(n3614), .B(n10545), .Z(n3577) );
  NANDN U3876 ( .A(n3575), .B(n10546), .Z(n3576) );
  NAND U3877 ( .A(n3577), .B(n3576), .Z(n3602) );
  XNOR U3878 ( .A(b[3]), .B(a[80]), .Z(n3617) );
  NANDN U3879 ( .A(n3617), .B(n10398), .Z(n3580) );
  NANDN U3880 ( .A(n3578), .B(n10399), .Z(n3579) );
  AND U3881 ( .A(n3580), .B(n3579), .Z(n3603) );
  XNOR U3882 ( .A(n3602), .B(n3603), .Z(n3604) );
  NANDN U3883 ( .A(n527), .B(a[82]), .Z(n3581) );
  XOR U3884 ( .A(n10434), .B(n3581), .Z(n3583) );
  NANDN U3885 ( .A(b[0]), .B(a[81]), .Z(n3582) );
  AND U3886 ( .A(n3583), .B(n3582), .Z(n3610) );
  XOR U3887 ( .A(b[5]), .B(a[78]), .Z(n3623) );
  NAND U3888 ( .A(n3623), .B(n10481), .Z(n3586) );
  NAND U3889 ( .A(n3584), .B(n10482), .Z(n3585) );
  NAND U3890 ( .A(n3586), .B(n3585), .Z(n3608) );
  NANDN U3891 ( .A(n529), .B(a[74]), .Z(n3609) );
  XNOR U3892 ( .A(n3608), .B(n3609), .Z(n3611) );
  XOR U3893 ( .A(n3610), .B(n3611), .Z(n3605) );
  XOR U3894 ( .A(n3604), .B(n3605), .Z(n3626) );
  XOR U3895 ( .A(n3627), .B(n3626), .Z(n3628) );
  XNOR U3896 ( .A(n3629), .B(n3628), .Z(n3598) );
  NAND U3897 ( .A(n3588), .B(n3587), .Z(n3592) );
  NAND U3898 ( .A(n3590), .B(n3589), .Z(n3591) );
  NAND U3899 ( .A(n3592), .B(n3591), .Z(n3599) );
  XNOR U3900 ( .A(n3598), .B(n3599), .Z(n3600) );
  XNOR U3901 ( .A(n3601), .B(n3600), .Z(n3632) );
  XNOR U3902 ( .A(n3632), .B(sreg[330]), .Z(n3634) );
  NAND U3903 ( .A(n3593), .B(sreg[329]), .Z(n3597) );
  OR U3904 ( .A(n3595), .B(n3594), .Z(n3596) );
  AND U3905 ( .A(n3597), .B(n3596), .Z(n3633) );
  XOR U3906 ( .A(n3634), .B(n3633), .Z(c[330]) );
  NANDN U3907 ( .A(n3603), .B(n3602), .Z(n3607) );
  NAND U3908 ( .A(n3605), .B(n3604), .Z(n3606) );
  NAND U3909 ( .A(n3607), .B(n3606), .Z(n3668) );
  NANDN U3910 ( .A(n3609), .B(n3608), .Z(n3613) );
  NAND U3911 ( .A(n3611), .B(n3610), .Z(n3612) );
  NAND U3912 ( .A(n3613), .B(n3612), .Z(n3666) );
  XNOR U3913 ( .A(b[7]), .B(a[77]), .Z(n3653) );
  NANDN U3914 ( .A(n3653), .B(n10545), .Z(n3616) );
  NANDN U3915 ( .A(n3614), .B(n10546), .Z(n3615) );
  NAND U3916 ( .A(n3616), .B(n3615), .Z(n3641) );
  XNOR U3917 ( .A(b[3]), .B(a[81]), .Z(n3656) );
  NANDN U3918 ( .A(n3656), .B(n10398), .Z(n3619) );
  NANDN U3919 ( .A(n3617), .B(n10399), .Z(n3618) );
  AND U3920 ( .A(n3619), .B(n3618), .Z(n3642) );
  XNOR U3921 ( .A(n3641), .B(n3642), .Z(n3643) );
  NANDN U3922 ( .A(n527), .B(a[83]), .Z(n3620) );
  XOR U3923 ( .A(n10434), .B(n3620), .Z(n3622) );
  NANDN U3924 ( .A(b[0]), .B(a[82]), .Z(n3621) );
  AND U3925 ( .A(n3622), .B(n3621), .Z(n3649) );
  XOR U3926 ( .A(b[5]), .B(a[79]), .Z(n3662) );
  NAND U3927 ( .A(n3662), .B(n10481), .Z(n3625) );
  NAND U3928 ( .A(n3623), .B(n10482), .Z(n3624) );
  NAND U3929 ( .A(n3625), .B(n3624), .Z(n3647) );
  NANDN U3930 ( .A(n529), .B(a[75]), .Z(n3648) );
  XNOR U3931 ( .A(n3647), .B(n3648), .Z(n3650) );
  XOR U3932 ( .A(n3649), .B(n3650), .Z(n3644) );
  XOR U3933 ( .A(n3643), .B(n3644), .Z(n3665) );
  XOR U3934 ( .A(n3666), .B(n3665), .Z(n3667) );
  XNOR U3935 ( .A(n3668), .B(n3667), .Z(n3637) );
  NAND U3936 ( .A(n3627), .B(n3626), .Z(n3631) );
  NAND U3937 ( .A(n3629), .B(n3628), .Z(n3630) );
  NAND U3938 ( .A(n3631), .B(n3630), .Z(n3638) );
  XNOR U3939 ( .A(n3637), .B(n3638), .Z(n3639) );
  XNOR U3940 ( .A(n3640), .B(n3639), .Z(n3671) );
  XNOR U3941 ( .A(n3671), .B(sreg[331]), .Z(n3673) );
  NAND U3942 ( .A(n3632), .B(sreg[330]), .Z(n3636) );
  OR U3943 ( .A(n3634), .B(n3633), .Z(n3635) );
  AND U3944 ( .A(n3636), .B(n3635), .Z(n3672) );
  XOR U3945 ( .A(n3673), .B(n3672), .Z(c[331]) );
  NANDN U3946 ( .A(n3642), .B(n3641), .Z(n3646) );
  NAND U3947 ( .A(n3644), .B(n3643), .Z(n3645) );
  NAND U3948 ( .A(n3646), .B(n3645), .Z(n3707) );
  NANDN U3949 ( .A(n3648), .B(n3647), .Z(n3652) );
  NAND U3950 ( .A(n3650), .B(n3649), .Z(n3651) );
  NAND U3951 ( .A(n3652), .B(n3651), .Z(n3705) );
  XNOR U3952 ( .A(b[7]), .B(a[78]), .Z(n3692) );
  NANDN U3953 ( .A(n3692), .B(n10545), .Z(n3655) );
  NANDN U3954 ( .A(n3653), .B(n10546), .Z(n3654) );
  NAND U3955 ( .A(n3655), .B(n3654), .Z(n3680) );
  XNOR U3956 ( .A(b[3]), .B(a[82]), .Z(n3695) );
  NANDN U3957 ( .A(n3695), .B(n10398), .Z(n3658) );
  NANDN U3958 ( .A(n3656), .B(n10399), .Z(n3657) );
  AND U3959 ( .A(n3658), .B(n3657), .Z(n3681) );
  XNOR U3960 ( .A(n3680), .B(n3681), .Z(n3682) );
  NANDN U3961 ( .A(n527), .B(a[84]), .Z(n3659) );
  XOR U3962 ( .A(n10434), .B(n3659), .Z(n3661) );
  NANDN U3963 ( .A(b[0]), .B(a[83]), .Z(n3660) );
  AND U3964 ( .A(n3661), .B(n3660), .Z(n3688) );
  XOR U3965 ( .A(b[5]), .B(a[80]), .Z(n3701) );
  NAND U3966 ( .A(n3701), .B(n10481), .Z(n3664) );
  NAND U3967 ( .A(n3662), .B(n10482), .Z(n3663) );
  NAND U3968 ( .A(n3664), .B(n3663), .Z(n3686) );
  NANDN U3969 ( .A(n529), .B(a[76]), .Z(n3687) );
  XNOR U3970 ( .A(n3686), .B(n3687), .Z(n3689) );
  XOR U3971 ( .A(n3688), .B(n3689), .Z(n3683) );
  XOR U3972 ( .A(n3682), .B(n3683), .Z(n3704) );
  XOR U3973 ( .A(n3705), .B(n3704), .Z(n3706) );
  XNOR U3974 ( .A(n3707), .B(n3706), .Z(n3676) );
  NAND U3975 ( .A(n3666), .B(n3665), .Z(n3670) );
  NAND U3976 ( .A(n3668), .B(n3667), .Z(n3669) );
  NAND U3977 ( .A(n3670), .B(n3669), .Z(n3677) );
  XNOR U3978 ( .A(n3676), .B(n3677), .Z(n3678) );
  XNOR U3979 ( .A(n3679), .B(n3678), .Z(n3710) );
  XNOR U3980 ( .A(n3710), .B(sreg[332]), .Z(n3712) );
  NAND U3981 ( .A(n3671), .B(sreg[331]), .Z(n3675) );
  OR U3982 ( .A(n3673), .B(n3672), .Z(n3674) );
  AND U3983 ( .A(n3675), .B(n3674), .Z(n3711) );
  XOR U3984 ( .A(n3712), .B(n3711), .Z(c[332]) );
  NANDN U3985 ( .A(n3681), .B(n3680), .Z(n3685) );
  NAND U3986 ( .A(n3683), .B(n3682), .Z(n3684) );
  NAND U3987 ( .A(n3685), .B(n3684), .Z(n3746) );
  NANDN U3988 ( .A(n3687), .B(n3686), .Z(n3691) );
  NAND U3989 ( .A(n3689), .B(n3688), .Z(n3690) );
  NAND U3990 ( .A(n3691), .B(n3690), .Z(n3744) );
  XNOR U3991 ( .A(b[7]), .B(a[79]), .Z(n3731) );
  NANDN U3992 ( .A(n3731), .B(n10545), .Z(n3694) );
  NANDN U3993 ( .A(n3692), .B(n10546), .Z(n3693) );
  NAND U3994 ( .A(n3694), .B(n3693), .Z(n3719) );
  XNOR U3995 ( .A(b[3]), .B(a[83]), .Z(n3734) );
  NANDN U3996 ( .A(n3734), .B(n10398), .Z(n3697) );
  NANDN U3997 ( .A(n3695), .B(n10399), .Z(n3696) );
  AND U3998 ( .A(n3697), .B(n3696), .Z(n3720) );
  XNOR U3999 ( .A(n3719), .B(n3720), .Z(n3721) );
  NANDN U4000 ( .A(n527), .B(a[85]), .Z(n3698) );
  XOR U4001 ( .A(n10434), .B(n3698), .Z(n3700) );
  NANDN U4002 ( .A(b[0]), .B(a[84]), .Z(n3699) );
  AND U4003 ( .A(n3700), .B(n3699), .Z(n3727) );
  XOR U4004 ( .A(b[5]), .B(a[81]), .Z(n3740) );
  NAND U4005 ( .A(n3740), .B(n10481), .Z(n3703) );
  NAND U4006 ( .A(n3701), .B(n10482), .Z(n3702) );
  NAND U4007 ( .A(n3703), .B(n3702), .Z(n3725) );
  NANDN U4008 ( .A(n529), .B(a[77]), .Z(n3726) );
  XNOR U4009 ( .A(n3725), .B(n3726), .Z(n3728) );
  XOR U4010 ( .A(n3727), .B(n3728), .Z(n3722) );
  XOR U4011 ( .A(n3721), .B(n3722), .Z(n3743) );
  XOR U4012 ( .A(n3744), .B(n3743), .Z(n3745) );
  XNOR U4013 ( .A(n3746), .B(n3745), .Z(n3715) );
  NAND U4014 ( .A(n3705), .B(n3704), .Z(n3709) );
  NAND U4015 ( .A(n3707), .B(n3706), .Z(n3708) );
  NAND U4016 ( .A(n3709), .B(n3708), .Z(n3716) );
  XNOR U4017 ( .A(n3715), .B(n3716), .Z(n3717) );
  XNOR U4018 ( .A(n3718), .B(n3717), .Z(n3749) );
  XNOR U4019 ( .A(n3749), .B(sreg[333]), .Z(n3751) );
  NAND U4020 ( .A(n3710), .B(sreg[332]), .Z(n3714) );
  OR U4021 ( .A(n3712), .B(n3711), .Z(n3713) );
  AND U4022 ( .A(n3714), .B(n3713), .Z(n3750) );
  XOR U4023 ( .A(n3751), .B(n3750), .Z(c[333]) );
  NANDN U4024 ( .A(n3720), .B(n3719), .Z(n3724) );
  NAND U4025 ( .A(n3722), .B(n3721), .Z(n3723) );
  NAND U4026 ( .A(n3724), .B(n3723), .Z(n3785) );
  NANDN U4027 ( .A(n3726), .B(n3725), .Z(n3730) );
  NAND U4028 ( .A(n3728), .B(n3727), .Z(n3729) );
  NAND U4029 ( .A(n3730), .B(n3729), .Z(n3783) );
  XNOR U4030 ( .A(b[7]), .B(a[80]), .Z(n3770) );
  NANDN U4031 ( .A(n3770), .B(n10545), .Z(n3733) );
  NANDN U4032 ( .A(n3731), .B(n10546), .Z(n3732) );
  NAND U4033 ( .A(n3733), .B(n3732), .Z(n3758) );
  XNOR U4034 ( .A(b[3]), .B(a[84]), .Z(n3773) );
  NANDN U4035 ( .A(n3773), .B(n10398), .Z(n3736) );
  NANDN U4036 ( .A(n3734), .B(n10399), .Z(n3735) );
  AND U4037 ( .A(n3736), .B(n3735), .Z(n3759) );
  XNOR U4038 ( .A(n3758), .B(n3759), .Z(n3760) );
  NANDN U4039 ( .A(n527), .B(a[86]), .Z(n3737) );
  XOR U4040 ( .A(n10434), .B(n3737), .Z(n3739) );
  NANDN U4041 ( .A(b[0]), .B(a[85]), .Z(n3738) );
  AND U4042 ( .A(n3739), .B(n3738), .Z(n3766) );
  XOR U4043 ( .A(b[5]), .B(a[82]), .Z(n3779) );
  NAND U4044 ( .A(n3779), .B(n10481), .Z(n3742) );
  NAND U4045 ( .A(n3740), .B(n10482), .Z(n3741) );
  NAND U4046 ( .A(n3742), .B(n3741), .Z(n3764) );
  NANDN U4047 ( .A(n529), .B(a[78]), .Z(n3765) );
  XNOR U4048 ( .A(n3764), .B(n3765), .Z(n3767) );
  XOR U4049 ( .A(n3766), .B(n3767), .Z(n3761) );
  XOR U4050 ( .A(n3760), .B(n3761), .Z(n3782) );
  XOR U4051 ( .A(n3783), .B(n3782), .Z(n3784) );
  XNOR U4052 ( .A(n3785), .B(n3784), .Z(n3754) );
  NAND U4053 ( .A(n3744), .B(n3743), .Z(n3748) );
  NAND U4054 ( .A(n3746), .B(n3745), .Z(n3747) );
  NAND U4055 ( .A(n3748), .B(n3747), .Z(n3755) );
  XNOR U4056 ( .A(n3754), .B(n3755), .Z(n3756) );
  XNOR U4057 ( .A(n3757), .B(n3756), .Z(n3788) );
  XNOR U4058 ( .A(n3788), .B(sreg[334]), .Z(n3790) );
  NAND U4059 ( .A(n3749), .B(sreg[333]), .Z(n3753) );
  OR U4060 ( .A(n3751), .B(n3750), .Z(n3752) );
  AND U4061 ( .A(n3753), .B(n3752), .Z(n3789) );
  XOR U4062 ( .A(n3790), .B(n3789), .Z(c[334]) );
  NANDN U4063 ( .A(n3759), .B(n3758), .Z(n3763) );
  NAND U4064 ( .A(n3761), .B(n3760), .Z(n3762) );
  NAND U4065 ( .A(n3763), .B(n3762), .Z(n3824) );
  NANDN U4066 ( .A(n3765), .B(n3764), .Z(n3769) );
  NAND U4067 ( .A(n3767), .B(n3766), .Z(n3768) );
  NAND U4068 ( .A(n3769), .B(n3768), .Z(n3822) );
  XNOR U4069 ( .A(b[7]), .B(a[81]), .Z(n3809) );
  NANDN U4070 ( .A(n3809), .B(n10545), .Z(n3772) );
  NANDN U4071 ( .A(n3770), .B(n10546), .Z(n3771) );
  NAND U4072 ( .A(n3772), .B(n3771), .Z(n3797) );
  XNOR U4073 ( .A(b[3]), .B(a[85]), .Z(n3812) );
  NANDN U4074 ( .A(n3812), .B(n10398), .Z(n3775) );
  NANDN U4075 ( .A(n3773), .B(n10399), .Z(n3774) );
  AND U4076 ( .A(n3775), .B(n3774), .Z(n3798) );
  XNOR U4077 ( .A(n3797), .B(n3798), .Z(n3799) );
  NANDN U4078 ( .A(n527), .B(a[87]), .Z(n3776) );
  XOR U4079 ( .A(n10434), .B(n3776), .Z(n3778) );
  NANDN U4080 ( .A(b[0]), .B(a[86]), .Z(n3777) );
  AND U4081 ( .A(n3778), .B(n3777), .Z(n3805) );
  XOR U4082 ( .A(b[5]), .B(a[83]), .Z(n3818) );
  NAND U4083 ( .A(n3818), .B(n10481), .Z(n3781) );
  NAND U4084 ( .A(n3779), .B(n10482), .Z(n3780) );
  NAND U4085 ( .A(n3781), .B(n3780), .Z(n3803) );
  NANDN U4086 ( .A(n529), .B(a[79]), .Z(n3804) );
  XNOR U4087 ( .A(n3803), .B(n3804), .Z(n3806) );
  XOR U4088 ( .A(n3805), .B(n3806), .Z(n3800) );
  XOR U4089 ( .A(n3799), .B(n3800), .Z(n3821) );
  XOR U4090 ( .A(n3822), .B(n3821), .Z(n3823) );
  XNOR U4091 ( .A(n3824), .B(n3823), .Z(n3793) );
  NAND U4092 ( .A(n3783), .B(n3782), .Z(n3787) );
  NAND U4093 ( .A(n3785), .B(n3784), .Z(n3786) );
  NAND U4094 ( .A(n3787), .B(n3786), .Z(n3794) );
  XNOR U4095 ( .A(n3793), .B(n3794), .Z(n3795) );
  XNOR U4096 ( .A(n3796), .B(n3795), .Z(n3827) );
  XNOR U4097 ( .A(n3827), .B(sreg[335]), .Z(n3829) );
  NAND U4098 ( .A(n3788), .B(sreg[334]), .Z(n3792) );
  OR U4099 ( .A(n3790), .B(n3789), .Z(n3791) );
  AND U4100 ( .A(n3792), .B(n3791), .Z(n3828) );
  XOR U4101 ( .A(n3829), .B(n3828), .Z(c[335]) );
  NANDN U4102 ( .A(n3798), .B(n3797), .Z(n3802) );
  NAND U4103 ( .A(n3800), .B(n3799), .Z(n3801) );
  NAND U4104 ( .A(n3802), .B(n3801), .Z(n3863) );
  NANDN U4105 ( .A(n3804), .B(n3803), .Z(n3808) );
  NAND U4106 ( .A(n3806), .B(n3805), .Z(n3807) );
  NAND U4107 ( .A(n3808), .B(n3807), .Z(n3861) );
  XNOR U4108 ( .A(b[7]), .B(a[82]), .Z(n3848) );
  NANDN U4109 ( .A(n3848), .B(n10545), .Z(n3811) );
  NANDN U4110 ( .A(n3809), .B(n10546), .Z(n3810) );
  NAND U4111 ( .A(n3811), .B(n3810), .Z(n3836) );
  XNOR U4112 ( .A(b[3]), .B(a[86]), .Z(n3851) );
  NANDN U4113 ( .A(n3851), .B(n10398), .Z(n3814) );
  NANDN U4114 ( .A(n3812), .B(n10399), .Z(n3813) );
  AND U4115 ( .A(n3814), .B(n3813), .Z(n3837) );
  XNOR U4116 ( .A(n3836), .B(n3837), .Z(n3838) );
  NANDN U4117 ( .A(n527), .B(a[88]), .Z(n3815) );
  XOR U4118 ( .A(n10434), .B(n3815), .Z(n3817) );
  NANDN U4119 ( .A(b[0]), .B(a[87]), .Z(n3816) );
  AND U4120 ( .A(n3817), .B(n3816), .Z(n3844) );
  XOR U4121 ( .A(b[5]), .B(a[84]), .Z(n3857) );
  NAND U4122 ( .A(n3857), .B(n10481), .Z(n3820) );
  NAND U4123 ( .A(n3818), .B(n10482), .Z(n3819) );
  NAND U4124 ( .A(n3820), .B(n3819), .Z(n3842) );
  NANDN U4125 ( .A(n529), .B(a[80]), .Z(n3843) );
  XNOR U4126 ( .A(n3842), .B(n3843), .Z(n3845) );
  XOR U4127 ( .A(n3844), .B(n3845), .Z(n3839) );
  XOR U4128 ( .A(n3838), .B(n3839), .Z(n3860) );
  XOR U4129 ( .A(n3861), .B(n3860), .Z(n3862) );
  XNOR U4130 ( .A(n3863), .B(n3862), .Z(n3832) );
  NAND U4131 ( .A(n3822), .B(n3821), .Z(n3826) );
  NAND U4132 ( .A(n3824), .B(n3823), .Z(n3825) );
  NAND U4133 ( .A(n3826), .B(n3825), .Z(n3833) );
  XNOR U4134 ( .A(n3832), .B(n3833), .Z(n3834) );
  XNOR U4135 ( .A(n3835), .B(n3834), .Z(n3866) );
  XNOR U4136 ( .A(n3866), .B(sreg[336]), .Z(n3868) );
  NAND U4137 ( .A(n3827), .B(sreg[335]), .Z(n3831) );
  OR U4138 ( .A(n3829), .B(n3828), .Z(n3830) );
  AND U4139 ( .A(n3831), .B(n3830), .Z(n3867) );
  XOR U4140 ( .A(n3868), .B(n3867), .Z(c[336]) );
  NANDN U4141 ( .A(n3837), .B(n3836), .Z(n3841) );
  NAND U4142 ( .A(n3839), .B(n3838), .Z(n3840) );
  NAND U4143 ( .A(n3841), .B(n3840), .Z(n3902) );
  NANDN U4144 ( .A(n3843), .B(n3842), .Z(n3847) );
  NAND U4145 ( .A(n3845), .B(n3844), .Z(n3846) );
  NAND U4146 ( .A(n3847), .B(n3846), .Z(n3900) );
  XNOR U4147 ( .A(b[7]), .B(a[83]), .Z(n3887) );
  NANDN U4148 ( .A(n3887), .B(n10545), .Z(n3850) );
  NANDN U4149 ( .A(n3848), .B(n10546), .Z(n3849) );
  NAND U4150 ( .A(n3850), .B(n3849), .Z(n3875) );
  XNOR U4151 ( .A(b[3]), .B(a[87]), .Z(n3890) );
  NANDN U4152 ( .A(n3890), .B(n10398), .Z(n3853) );
  NANDN U4153 ( .A(n3851), .B(n10399), .Z(n3852) );
  AND U4154 ( .A(n3853), .B(n3852), .Z(n3876) );
  XNOR U4155 ( .A(n3875), .B(n3876), .Z(n3877) );
  NANDN U4156 ( .A(n527), .B(a[89]), .Z(n3854) );
  XOR U4157 ( .A(n10434), .B(n3854), .Z(n3856) );
  NANDN U4158 ( .A(b[0]), .B(a[88]), .Z(n3855) );
  AND U4159 ( .A(n3856), .B(n3855), .Z(n3883) );
  XOR U4160 ( .A(b[5]), .B(a[85]), .Z(n3896) );
  NAND U4161 ( .A(n3896), .B(n10481), .Z(n3859) );
  NAND U4162 ( .A(n3857), .B(n10482), .Z(n3858) );
  NAND U4163 ( .A(n3859), .B(n3858), .Z(n3881) );
  NANDN U4164 ( .A(n529), .B(a[81]), .Z(n3882) );
  XNOR U4165 ( .A(n3881), .B(n3882), .Z(n3884) );
  XOR U4166 ( .A(n3883), .B(n3884), .Z(n3878) );
  XOR U4167 ( .A(n3877), .B(n3878), .Z(n3899) );
  XOR U4168 ( .A(n3900), .B(n3899), .Z(n3901) );
  XNOR U4169 ( .A(n3902), .B(n3901), .Z(n3871) );
  NAND U4170 ( .A(n3861), .B(n3860), .Z(n3865) );
  NAND U4171 ( .A(n3863), .B(n3862), .Z(n3864) );
  NAND U4172 ( .A(n3865), .B(n3864), .Z(n3872) );
  XNOR U4173 ( .A(n3871), .B(n3872), .Z(n3873) );
  XNOR U4174 ( .A(n3874), .B(n3873), .Z(n3905) );
  XNOR U4175 ( .A(n3905), .B(sreg[337]), .Z(n3907) );
  NAND U4176 ( .A(n3866), .B(sreg[336]), .Z(n3870) );
  OR U4177 ( .A(n3868), .B(n3867), .Z(n3869) );
  AND U4178 ( .A(n3870), .B(n3869), .Z(n3906) );
  XOR U4179 ( .A(n3907), .B(n3906), .Z(c[337]) );
  NANDN U4180 ( .A(n3876), .B(n3875), .Z(n3880) );
  NAND U4181 ( .A(n3878), .B(n3877), .Z(n3879) );
  NAND U4182 ( .A(n3880), .B(n3879), .Z(n3941) );
  NANDN U4183 ( .A(n3882), .B(n3881), .Z(n3886) );
  NAND U4184 ( .A(n3884), .B(n3883), .Z(n3885) );
  NAND U4185 ( .A(n3886), .B(n3885), .Z(n3939) );
  XNOR U4186 ( .A(b[7]), .B(a[84]), .Z(n3926) );
  NANDN U4187 ( .A(n3926), .B(n10545), .Z(n3889) );
  NANDN U4188 ( .A(n3887), .B(n10546), .Z(n3888) );
  NAND U4189 ( .A(n3889), .B(n3888), .Z(n3914) );
  XNOR U4190 ( .A(b[3]), .B(a[88]), .Z(n3929) );
  NANDN U4191 ( .A(n3929), .B(n10398), .Z(n3892) );
  NANDN U4192 ( .A(n3890), .B(n10399), .Z(n3891) );
  AND U4193 ( .A(n3892), .B(n3891), .Z(n3915) );
  XNOR U4194 ( .A(n3914), .B(n3915), .Z(n3916) );
  NANDN U4195 ( .A(n527), .B(a[90]), .Z(n3893) );
  XOR U4196 ( .A(n10434), .B(n3893), .Z(n3895) );
  NANDN U4197 ( .A(b[0]), .B(a[89]), .Z(n3894) );
  AND U4198 ( .A(n3895), .B(n3894), .Z(n3922) );
  XOR U4199 ( .A(b[5]), .B(a[86]), .Z(n3935) );
  NAND U4200 ( .A(n3935), .B(n10481), .Z(n3898) );
  NAND U4201 ( .A(n3896), .B(n10482), .Z(n3897) );
  NAND U4202 ( .A(n3898), .B(n3897), .Z(n3920) );
  NANDN U4203 ( .A(n529), .B(a[82]), .Z(n3921) );
  XNOR U4204 ( .A(n3920), .B(n3921), .Z(n3923) );
  XOR U4205 ( .A(n3922), .B(n3923), .Z(n3917) );
  XOR U4206 ( .A(n3916), .B(n3917), .Z(n3938) );
  XOR U4207 ( .A(n3939), .B(n3938), .Z(n3940) );
  XNOR U4208 ( .A(n3941), .B(n3940), .Z(n3910) );
  NAND U4209 ( .A(n3900), .B(n3899), .Z(n3904) );
  NAND U4210 ( .A(n3902), .B(n3901), .Z(n3903) );
  NAND U4211 ( .A(n3904), .B(n3903), .Z(n3911) );
  XNOR U4212 ( .A(n3910), .B(n3911), .Z(n3912) );
  XNOR U4213 ( .A(n3913), .B(n3912), .Z(n3944) );
  XNOR U4214 ( .A(n3944), .B(sreg[338]), .Z(n3946) );
  NAND U4215 ( .A(n3905), .B(sreg[337]), .Z(n3909) );
  OR U4216 ( .A(n3907), .B(n3906), .Z(n3908) );
  AND U4217 ( .A(n3909), .B(n3908), .Z(n3945) );
  XOR U4218 ( .A(n3946), .B(n3945), .Z(c[338]) );
  NANDN U4219 ( .A(n3915), .B(n3914), .Z(n3919) );
  NAND U4220 ( .A(n3917), .B(n3916), .Z(n3918) );
  NAND U4221 ( .A(n3919), .B(n3918), .Z(n3980) );
  NANDN U4222 ( .A(n3921), .B(n3920), .Z(n3925) );
  NAND U4223 ( .A(n3923), .B(n3922), .Z(n3924) );
  NAND U4224 ( .A(n3925), .B(n3924), .Z(n3978) );
  XNOR U4225 ( .A(b[7]), .B(a[85]), .Z(n3965) );
  NANDN U4226 ( .A(n3965), .B(n10545), .Z(n3928) );
  NANDN U4227 ( .A(n3926), .B(n10546), .Z(n3927) );
  NAND U4228 ( .A(n3928), .B(n3927), .Z(n3953) );
  XNOR U4229 ( .A(b[3]), .B(a[89]), .Z(n3968) );
  NANDN U4230 ( .A(n3968), .B(n10398), .Z(n3931) );
  NANDN U4231 ( .A(n3929), .B(n10399), .Z(n3930) );
  AND U4232 ( .A(n3931), .B(n3930), .Z(n3954) );
  XNOR U4233 ( .A(n3953), .B(n3954), .Z(n3955) );
  NANDN U4234 ( .A(n527), .B(a[91]), .Z(n3932) );
  XOR U4235 ( .A(n10434), .B(n3932), .Z(n3934) );
  NANDN U4236 ( .A(b[0]), .B(a[90]), .Z(n3933) );
  AND U4237 ( .A(n3934), .B(n3933), .Z(n3961) );
  XOR U4238 ( .A(b[5]), .B(a[87]), .Z(n3974) );
  NAND U4239 ( .A(n3974), .B(n10481), .Z(n3937) );
  NAND U4240 ( .A(n3935), .B(n10482), .Z(n3936) );
  NAND U4241 ( .A(n3937), .B(n3936), .Z(n3959) );
  NANDN U4242 ( .A(n529), .B(a[83]), .Z(n3960) );
  XNOR U4243 ( .A(n3959), .B(n3960), .Z(n3962) );
  XOR U4244 ( .A(n3961), .B(n3962), .Z(n3956) );
  XOR U4245 ( .A(n3955), .B(n3956), .Z(n3977) );
  XOR U4246 ( .A(n3978), .B(n3977), .Z(n3979) );
  XNOR U4247 ( .A(n3980), .B(n3979), .Z(n3949) );
  NAND U4248 ( .A(n3939), .B(n3938), .Z(n3943) );
  NAND U4249 ( .A(n3941), .B(n3940), .Z(n3942) );
  NAND U4250 ( .A(n3943), .B(n3942), .Z(n3950) );
  XNOR U4251 ( .A(n3949), .B(n3950), .Z(n3951) );
  XNOR U4252 ( .A(n3952), .B(n3951), .Z(n3983) );
  XNOR U4253 ( .A(n3983), .B(sreg[339]), .Z(n3985) );
  NAND U4254 ( .A(n3944), .B(sreg[338]), .Z(n3948) );
  OR U4255 ( .A(n3946), .B(n3945), .Z(n3947) );
  AND U4256 ( .A(n3948), .B(n3947), .Z(n3984) );
  XOR U4257 ( .A(n3985), .B(n3984), .Z(c[339]) );
  NANDN U4258 ( .A(n3954), .B(n3953), .Z(n3958) );
  NAND U4259 ( .A(n3956), .B(n3955), .Z(n3957) );
  NAND U4260 ( .A(n3958), .B(n3957), .Z(n4019) );
  NANDN U4261 ( .A(n3960), .B(n3959), .Z(n3964) );
  NAND U4262 ( .A(n3962), .B(n3961), .Z(n3963) );
  NAND U4263 ( .A(n3964), .B(n3963), .Z(n4017) );
  XNOR U4264 ( .A(b[7]), .B(a[86]), .Z(n4004) );
  NANDN U4265 ( .A(n4004), .B(n10545), .Z(n3967) );
  NANDN U4266 ( .A(n3965), .B(n10546), .Z(n3966) );
  NAND U4267 ( .A(n3967), .B(n3966), .Z(n3992) );
  XNOR U4268 ( .A(b[3]), .B(a[90]), .Z(n4007) );
  NANDN U4269 ( .A(n4007), .B(n10398), .Z(n3970) );
  NANDN U4270 ( .A(n3968), .B(n10399), .Z(n3969) );
  AND U4271 ( .A(n3970), .B(n3969), .Z(n3993) );
  XNOR U4272 ( .A(n3992), .B(n3993), .Z(n3994) );
  NANDN U4273 ( .A(n527), .B(a[92]), .Z(n3971) );
  XOR U4274 ( .A(n10434), .B(n3971), .Z(n3973) );
  NANDN U4275 ( .A(b[0]), .B(a[91]), .Z(n3972) );
  AND U4276 ( .A(n3973), .B(n3972), .Z(n4000) );
  XOR U4277 ( .A(b[5]), .B(a[88]), .Z(n4013) );
  NAND U4278 ( .A(n4013), .B(n10481), .Z(n3976) );
  NAND U4279 ( .A(n3974), .B(n10482), .Z(n3975) );
  NAND U4280 ( .A(n3976), .B(n3975), .Z(n3998) );
  NANDN U4281 ( .A(n529), .B(a[84]), .Z(n3999) );
  XNOR U4282 ( .A(n3998), .B(n3999), .Z(n4001) );
  XOR U4283 ( .A(n4000), .B(n4001), .Z(n3995) );
  XOR U4284 ( .A(n3994), .B(n3995), .Z(n4016) );
  XOR U4285 ( .A(n4017), .B(n4016), .Z(n4018) );
  XNOR U4286 ( .A(n4019), .B(n4018), .Z(n3988) );
  NAND U4287 ( .A(n3978), .B(n3977), .Z(n3982) );
  NAND U4288 ( .A(n3980), .B(n3979), .Z(n3981) );
  NAND U4289 ( .A(n3982), .B(n3981), .Z(n3989) );
  XNOR U4290 ( .A(n3988), .B(n3989), .Z(n3990) );
  XNOR U4291 ( .A(n3991), .B(n3990), .Z(n4022) );
  XNOR U4292 ( .A(n4022), .B(sreg[340]), .Z(n4024) );
  NAND U4293 ( .A(n3983), .B(sreg[339]), .Z(n3987) );
  OR U4294 ( .A(n3985), .B(n3984), .Z(n3986) );
  AND U4295 ( .A(n3987), .B(n3986), .Z(n4023) );
  XOR U4296 ( .A(n4024), .B(n4023), .Z(c[340]) );
  NANDN U4297 ( .A(n3993), .B(n3992), .Z(n3997) );
  NAND U4298 ( .A(n3995), .B(n3994), .Z(n3996) );
  NAND U4299 ( .A(n3997), .B(n3996), .Z(n4058) );
  NANDN U4300 ( .A(n3999), .B(n3998), .Z(n4003) );
  NAND U4301 ( .A(n4001), .B(n4000), .Z(n4002) );
  NAND U4302 ( .A(n4003), .B(n4002), .Z(n4056) );
  XNOR U4303 ( .A(b[7]), .B(a[87]), .Z(n4043) );
  NANDN U4304 ( .A(n4043), .B(n10545), .Z(n4006) );
  NANDN U4305 ( .A(n4004), .B(n10546), .Z(n4005) );
  NAND U4306 ( .A(n4006), .B(n4005), .Z(n4031) );
  XNOR U4307 ( .A(b[3]), .B(a[91]), .Z(n4046) );
  NANDN U4308 ( .A(n4046), .B(n10398), .Z(n4009) );
  NANDN U4309 ( .A(n4007), .B(n10399), .Z(n4008) );
  AND U4310 ( .A(n4009), .B(n4008), .Z(n4032) );
  XNOR U4311 ( .A(n4031), .B(n4032), .Z(n4033) );
  NANDN U4312 ( .A(n527), .B(a[93]), .Z(n4010) );
  XOR U4313 ( .A(n10434), .B(n4010), .Z(n4012) );
  NANDN U4314 ( .A(b[0]), .B(a[92]), .Z(n4011) );
  AND U4315 ( .A(n4012), .B(n4011), .Z(n4039) );
  XOR U4316 ( .A(b[5]), .B(a[89]), .Z(n4052) );
  NAND U4317 ( .A(n4052), .B(n10481), .Z(n4015) );
  NAND U4318 ( .A(n4013), .B(n10482), .Z(n4014) );
  NAND U4319 ( .A(n4015), .B(n4014), .Z(n4037) );
  NANDN U4320 ( .A(n529), .B(a[85]), .Z(n4038) );
  XNOR U4321 ( .A(n4037), .B(n4038), .Z(n4040) );
  XOR U4322 ( .A(n4039), .B(n4040), .Z(n4034) );
  XOR U4323 ( .A(n4033), .B(n4034), .Z(n4055) );
  XOR U4324 ( .A(n4056), .B(n4055), .Z(n4057) );
  XNOR U4325 ( .A(n4058), .B(n4057), .Z(n4027) );
  NAND U4326 ( .A(n4017), .B(n4016), .Z(n4021) );
  NAND U4327 ( .A(n4019), .B(n4018), .Z(n4020) );
  NAND U4328 ( .A(n4021), .B(n4020), .Z(n4028) );
  XNOR U4329 ( .A(n4027), .B(n4028), .Z(n4029) );
  XNOR U4330 ( .A(n4030), .B(n4029), .Z(n4061) );
  XNOR U4331 ( .A(n4061), .B(sreg[341]), .Z(n4063) );
  NAND U4332 ( .A(n4022), .B(sreg[340]), .Z(n4026) );
  OR U4333 ( .A(n4024), .B(n4023), .Z(n4025) );
  AND U4334 ( .A(n4026), .B(n4025), .Z(n4062) );
  XOR U4335 ( .A(n4063), .B(n4062), .Z(c[341]) );
  NANDN U4336 ( .A(n4032), .B(n4031), .Z(n4036) );
  NAND U4337 ( .A(n4034), .B(n4033), .Z(n4035) );
  NAND U4338 ( .A(n4036), .B(n4035), .Z(n4097) );
  NANDN U4339 ( .A(n4038), .B(n4037), .Z(n4042) );
  NAND U4340 ( .A(n4040), .B(n4039), .Z(n4041) );
  NAND U4341 ( .A(n4042), .B(n4041), .Z(n4095) );
  XNOR U4342 ( .A(b[7]), .B(a[88]), .Z(n4082) );
  NANDN U4343 ( .A(n4082), .B(n10545), .Z(n4045) );
  NANDN U4344 ( .A(n4043), .B(n10546), .Z(n4044) );
  NAND U4345 ( .A(n4045), .B(n4044), .Z(n4070) );
  XNOR U4346 ( .A(b[3]), .B(a[92]), .Z(n4085) );
  NANDN U4347 ( .A(n4085), .B(n10398), .Z(n4048) );
  NANDN U4348 ( .A(n4046), .B(n10399), .Z(n4047) );
  AND U4349 ( .A(n4048), .B(n4047), .Z(n4071) );
  XNOR U4350 ( .A(n4070), .B(n4071), .Z(n4072) );
  NANDN U4351 ( .A(n527), .B(a[94]), .Z(n4049) );
  XOR U4352 ( .A(n10434), .B(n4049), .Z(n4051) );
  NANDN U4353 ( .A(b[0]), .B(a[93]), .Z(n4050) );
  AND U4354 ( .A(n4051), .B(n4050), .Z(n4078) );
  XOR U4355 ( .A(b[5]), .B(a[90]), .Z(n4091) );
  NAND U4356 ( .A(n4091), .B(n10481), .Z(n4054) );
  NAND U4357 ( .A(n4052), .B(n10482), .Z(n4053) );
  NAND U4358 ( .A(n4054), .B(n4053), .Z(n4076) );
  NANDN U4359 ( .A(n529), .B(a[86]), .Z(n4077) );
  XNOR U4360 ( .A(n4076), .B(n4077), .Z(n4079) );
  XOR U4361 ( .A(n4078), .B(n4079), .Z(n4073) );
  XOR U4362 ( .A(n4072), .B(n4073), .Z(n4094) );
  XOR U4363 ( .A(n4095), .B(n4094), .Z(n4096) );
  XNOR U4364 ( .A(n4097), .B(n4096), .Z(n4066) );
  NAND U4365 ( .A(n4056), .B(n4055), .Z(n4060) );
  NAND U4366 ( .A(n4058), .B(n4057), .Z(n4059) );
  NAND U4367 ( .A(n4060), .B(n4059), .Z(n4067) );
  XNOR U4368 ( .A(n4066), .B(n4067), .Z(n4068) );
  XNOR U4369 ( .A(n4069), .B(n4068), .Z(n4100) );
  XNOR U4370 ( .A(n4100), .B(sreg[342]), .Z(n4102) );
  NAND U4371 ( .A(n4061), .B(sreg[341]), .Z(n4065) );
  OR U4372 ( .A(n4063), .B(n4062), .Z(n4064) );
  AND U4373 ( .A(n4065), .B(n4064), .Z(n4101) );
  XOR U4374 ( .A(n4102), .B(n4101), .Z(c[342]) );
  NANDN U4375 ( .A(n4071), .B(n4070), .Z(n4075) );
  NAND U4376 ( .A(n4073), .B(n4072), .Z(n4074) );
  NAND U4377 ( .A(n4075), .B(n4074), .Z(n4136) );
  NANDN U4378 ( .A(n4077), .B(n4076), .Z(n4081) );
  NAND U4379 ( .A(n4079), .B(n4078), .Z(n4080) );
  NAND U4380 ( .A(n4081), .B(n4080), .Z(n4134) );
  XNOR U4381 ( .A(b[7]), .B(a[89]), .Z(n4121) );
  NANDN U4382 ( .A(n4121), .B(n10545), .Z(n4084) );
  NANDN U4383 ( .A(n4082), .B(n10546), .Z(n4083) );
  NAND U4384 ( .A(n4084), .B(n4083), .Z(n4109) );
  XNOR U4385 ( .A(b[3]), .B(a[93]), .Z(n4124) );
  NANDN U4386 ( .A(n4124), .B(n10398), .Z(n4087) );
  NANDN U4387 ( .A(n4085), .B(n10399), .Z(n4086) );
  AND U4388 ( .A(n4087), .B(n4086), .Z(n4110) );
  XNOR U4389 ( .A(n4109), .B(n4110), .Z(n4111) );
  NANDN U4390 ( .A(n527), .B(a[95]), .Z(n4088) );
  XOR U4391 ( .A(n10434), .B(n4088), .Z(n4090) );
  NANDN U4392 ( .A(b[0]), .B(a[94]), .Z(n4089) );
  AND U4393 ( .A(n4090), .B(n4089), .Z(n4117) );
  XOR U4394 ( .A(b[5]), .B(a[91]), .Z(n4130) );
  NAND U4395 ( .A(n4130), .B(n10481), .Z(n4093) );
  NAND U4396 ( .A(n4091), .B(n10482), .Z(n4092) );
  NAND U4397 ( .A(n4093), .B(n4092), .Z(n4115) );
  NANDN U4398 ( .A(n529), .B(a[87]), .Z(n4116) );
  XNOR U4399 ( .A(n4115), .B(n4116), .Z(n4118) );
  XOR U4400 ( .A(n4117), .B(n4118), .Z(n4112) );
  XOR U4401 ( .A(n4111), .B(n4112), .Z(n4133) );
  XOR U4402 ( .A(n4134), .B(n4133), .Z(n4135) );
  XNOR U4403 ( .A(n4136), .B(n4135), .Z(n4105) );
  NAND U4404 ( .A(n4095), .B(n4094), .Z(n4099) );
  NAND U4405 ( .A(n4097), .B(n4096), .Z(n4098) );
  NAND U4406 ( .A(n4099), .B(n4098), .Z(n4106) );
  XNOR U4407 ( .A(n4105), .B(n4106), .Z(n4107) );
  XNOR U4408 ( .A(n4108), .B(n4107), .Z(n4139) );
  XNOR U4409 ( .A(n4139), .B(sreg[343]), .Z(n4141) );
  NAND U4410 ( .A(n4100), .B(sreg[342]), .Z(n4104) );
  OR U4411 ( .A(n4102), .B(n4101), .Z(n4103) );
  AND U4412 ( .A(n4104), .B(n4103), .Z(n4140) );
  XOR U4413 ( .A(n4141), .B(n4140), .Z(c[343]) );
  NANDN U4414 ( .A(n4110), .B(n4109), .Z(n4114) );
  NAND U4415 ( .A(n4112), .B(n4111), .Z(n4113) );
  NAND U4416 ( .A(n4114), .B(n4113), .Z(n4175) );
  NANDN U4417 ( .A(n4116), .B(n4115), .Z(n4120) );
  NAND U4418 ( .A(n4118), .B(n4117), .Z(n4119) );
  NAND U4419 ( .A(n4120), .B(n4119), .Z(n4173) );
  XNOR U4420 ( .A(b[7]), .B(a[90]), .Z(n4160) );
  NANDN U4421 ( .A(n4160), .B(n10545), .Z(n4123) );
  NANDN U4422 ( .A(n4121), .B(n10546), .Z(n4122) );
  NAND U4423 ( .A(n4123), .B(n4122), .Z(n4148) );
  XNOR U4424 ( .A(b[3]), .B(a[94]), .Z(n4163) );
  NANDN U4425 ( .A(n4163), .B(n10398), .Z(n4126) );
  NANDN U4426 ( .A(n4124), .B(n10399), .Z(n4125) );
  AND U4427 ( .A(n4126), .B(n4125), .Z(n4149) );
  XNOR U4428 ( .A(n4148), .B(n4149), .Z(n4150) );
  NANDN U4429 ( .A(n527), .B(a[96]), .Z(n4127) );
  XOR U4430 ( .A(n10434), .B(n4127), .Z(n4129) );
  NANDN U4431 ( .A(b[0]), .B(a[95]), .Z(n4128) );
  AND U4432 ( .A(n4129), .B(n4128), .Z(n4156) );
  XOR U4433 ( .A(b[5]), .B(a[92]), .Z(n4169) );
  NAND U4434 ( .A(n4169), .B(n10481), .Z(n4132) );
  NAND U4435 ( .A(n4130), .B(n10482), .Z(n4131) );
  NAND U4436 ( .A(n4132), .B(n4131), .Z(n4154) );
  NANDN U4437 ( .A(n529), .B(a[88]), .Z(n4155) );
  XNOR U4438 ( .A(n4154), .B(n4155), .Z(n4157) );
  XOR U4439 ( .A(n4156), .B(n4157), .Z(n4151) );
  XOR U4440 ( .A(n4150), .B(n4151), .Z(n4172) );
  XOR U4441 ( .A(n4173), .B(n4172), .Z(n4174) );
  XNOR U4442 ( .A(n4175), .B(n4174), .Z(n4144) );
  NAND U4443 ( .A(n4134), .B(n4133), .Z(n4138) );
  NAND U4444 ( .A(n4136), .B(n4135), .Z(n4137) );
  NAND U4445 ( .A(n4138), .B(n4137), .Z(n4145) );
  XNOR U4446 ( .A(n4144), .B(n4145), .Z(n4146) );
  XNOR U4447 ( .A(n4147), .B(n4146), .Z(n4178) );
  XNOR U4448 ( .A(n4178), .B(sreg[344]), .Z(n4180) );
  NAND U4449 ( .A(n4139), .B(sreg[343]), .Z(n4143) );
  OR U4450 ( .A(n4141), .B(n4140), .Z(n4142) );
  AND U4451 ( .A(n4143), .B(n4142), .Z(n4179) );
  XOR U4452 ( .A(n4180), .B(n4179), .Z(c[344]) );
  NANDN U4453 ( .A(n4149), .B(n4148), .Z(n4153) );
  NAND U4454 ( .A(n4151), .B(n4150), .Z(n4152) );
  NAND U4455 ( .A(n4153), .B(n4152), .Z(n4214) );
  NANDN U4456 ( .A(n4155), .B(n4154), .Z(n4159) );
  NAND U4457 ( .A(n4157), .B(n4156), .Z(n4158) );
  NAND U4458 ( .A(n4159), .B(n4158), .Z(n4212) );
  XNOR U4459 ( .A(b[7]), .B(a[91]), .Z(n4199) );
  NANDN U4460 ( .A(n4199), .B(n10545), .Z(n4162) );
  NANDN U4461 ( .A(n4160), .B(n10546), .Z(n4161) );
  NAND U4462 ( .A(n4162), .B(n4161), .Z(n4187) );
  XNOR U4463 ( .A(b[3]), .B(a[95]), .Z(n4202) );
  NANDN U4464 ( .A(n4202), .B(n10398), .Z(n4165) );
  NANDN U4465 ( .A(n4163), .B(n10399), .Z(n4164) );
  AND U4466 ( .A(n4165), .B(n4164), .Z(n4188) );
  XNOR U4467 ( .A(n4187), .B(n4188), .Z(n4189) );
  NANDN U4468 ( .A(n527), .B(a[97]), .Z(n4166) );
  XOR U4469 ( .A(n10434), .B(n4166), .Z(n4168) );
  NANDN U4470 ( .A(b[0]), .B(a[96]), .Z(n4167) );
  AND U4471 ( .A(n4168), .B(n4167), .Z(n4195) );
  XOR U4472 ( .A(b[5]), .B(a[93]), .Z(n4208) );
  NAND U4473 ( .A(n4208), .B(n10481), .Z(n4171) );
  NAND U4474 ( .A(n4169), .B(n10482), .Z(n4170) );
  NAND U4475 ( .A(n4171), .B(n4170), .Z(n4193) );
  NANDN U4476 ( .A(n529), .B(a[89]), .Z(n4194) );
  XNOR U4477 ( .A(n4193), .B(n4194), .Z(n4196) );
  XOR U4478 ( .A(n4195), .B(n4196), .Z(n4190) );
  XOR U4479 ( .A(n4189), .B(n4190), .Z(n4211) );
  XOR U4480 ( .A(n4212), .B(n4211), .Z(n4213) );
  XNOR U4481 ( .A(n4214), .B(n4213), .Z(n4183) );
  NAND U4482 ( .A(n4173), .B(n4172), .Z(n4177) );
  NAND U4483 ( .A(n4175), .B(n4174), .Z(n4176) );
  NAND U4484 ( .A(n4177), .B(n4176), .Z(n4184) );
  XNOR U4485 ( .A(n4183), .B(n4184), .Z(n4185) );
  XNOR U4486 ( .A(n4186), .B(n4185), .Z(n4217) );
  XNOR U4487 ( .A(n4217), .B(sreg[345]), .Z(n4219) );
  NAND U4488 ( .A(n4178), .B(sreg[344]), .Z(n4182) );
  OR U4489 ( .A(n4180), .B(n4179), .Z(n4181) );
  AND U4490 ( .A(n4182), .B(n4181), .Z(n4218) );
  XOR U4491 ( .A(n4219), .B(n4218), .Z(c[345]) );
  NANDN U4492 ( .A(n4188), .B(n4187), .Z(n4192) );
  NAND U4493 ( .A(n4190), .B(n4189), .Z(n4191) );
  NAND U4494 ( .A(n4192), .B(n4191), .Z(n4253) );
  NANDN U4495 ( .A(n4194), .B(n4193), .Z(n4198) );
  NAND U4496 ( .A(n4196), .B(n4195), .Z(n4197) );
  NAND U4497 ( .A(n4198), .B(n4197), .Z(n4251) );
  XNOR U4498 ( .A(b[7]), .B(a[92]), .Z(n4238) );
  NANDN U4499 ( .A(n4238), .B(n10545), .Z(n4201) );
  NANDN U4500 ( .A(n4199), .B(n10546), .Z(n4200) );
  NAND U4501 ( .A(n4201), .B(n4200), .Z(n4226) );
  XNOR U4502 ( .A(b[3]), .B(a[96]), .Z(n4241) );
  NANDN U4503 ( .A(n4241), .B(n10398), .Z(n4204) );
  NANDN U4504 ( .A(n4202), .B(n10399), .Z(n4203) );
  AND U4505 ( .A(n4204), .B(n4203), .Z(n4227) );
  XNOR U4506 ( .A(n4226), .B(n4227), .Z(n4228) );
  NANDN U4507 ( .A(n527), .B(a[98]), .Z(n4205) );
  XOR U4508 ( .A(n10434), .B(n4205), .Z(n4207) );
  NANDN U4509 ( .A(b[0]), .B(a[97]), .Z(n4206) );
  AND U4510 ( .A(n4207), .B(n4206), .Z(n4234) );
  XOR U4511 ( .A(b[5]), .B(a[94]), .Z(n4247) );
  NAND U4512 ( .A(n4247), .B(n10481), .Z(n4210) );
  NAND U4513 ( .A(n4208), .B(n10482), .Z(n4209) );
  NAND U4514 ( .A(n4210), .B(n4209), .Z(n4232) );
  NANDN U4515 ( .A(n529), .B(a[90]), .Z(n4233) );
  XNOR U4516 ( .A(n4232), .B(n4233), .Z(n4235) );
  XOR U4517 ( .A(n4234), .B(n4235), .Z(n4229) );
  XOR U4518 ( .A(n4228), .B(n4229), .Z(n4250) );
  XOR U4519 ( .A(n4251), .B(n4250), .Z(n4252) );
  XNOR U4520 ( .A(n4253), .B(n4252), .Z(n4222) );
  NAND U4521 ( .A(n4212), .B(n4211), .Z(n4216) );
  NAND U4522 ( .A(n4214), .B(n4213), .Z(n4215) );
  NAND U4523 ( .A(n4216), .B(n4215), .Z(n4223) );
  XNOR U4524 ( .A(n4222), .B(n4223), .Z(n4224) );
  XNOR U4525 ( .A(n4225), .B(n4224), .Z(n4256) );
  XNOR U4526 ( .A(n4256), .B(sreg[346]), .Z(n4258) );
  NAND U4527 ( .A(n4217), .B(sreg[345]), .Z(n4221) );
  OR U4528 ( .A(n4219), .B(n4218), .Z(n4220) );
  AND U4529 ( .A(n4221), .B(n4220), .Z(n4257) );
  XOR U4530 ( .A(n4258), .B(n4257), .Z(c[346]) );
  NANDN U4531 ( .A(n4227), .B(n4226), .Z(n4231) );
  NAND U4532 ( .A(n4229), .B(n4228), .Z(n4230) );
  NAND U4533 ( .A(n4231), .B(n4230), .Z(n4292) );
  NANDN U4534 ( .A(n4233), .B(n4232), .Z(n4237) );
  NAND U4535 ( .A(n4235), .B(n4234), .Z(n4236) );
  NAND U4536 ( .A(n4237), .B(n4236), .Z(n4290) );
  XNOR U4537 ( .A(b[7]), .B(a[93]), .Z(n4277) );
  NANDN U4538 ( .A(n4277), .B(n10545), .Z(n4240) );
  NANDN U4539 ( .A(n4238), .B(n10546), .Z(n4239) );
  NAND U4540 ( .A(n4240), .B(n4239), .Z(n4265) );
  XNOR U4541 ( .A(b[3]), .B(a[97]), .Z(n4280) );
  NANDN U4542 ( .A(n4280), .B(n10398), .Z(n4243) );
  NANDN U4543 ( .A(n4241), .B(n10399), .Z(n4242) );
  AND U4544 ( .A(n4243), .B(n4242), .Z(n4266) );
  XNOR U4545 ( .A(n4265), .B(n4266), .Z(n4267) );
  NANDN U4546 ( .A(n527), .B(a[99]), .Z(n4244) );
  XOR U4547 ( .A(n10434), .B(n4244), .Z(n4246) );
  NANDN U4548 ( .A(b[0]), .B(a[98]), .Z(n4245) );
  AND U4549 ( .A(n4246), .B(n4245), .Z(n4273) );
  XOR U4550 ( .A(b[5]), .B(a[95]), .Z(n4286) );
  NAND U4551 ( .A(n4286), .B(n10481), .Z(n4249) );
  NAND U4552 ( .A(n4247), .B(n10482), .Z(n4248) );
  NAND U4553 ( .A(n4249), .B(n4248), .Z(n4271) );
  NANDN U4554 ( .A(n529), .B(a[91]), .Z(n4272) );
  XNOR U4555 ( .A(n4271), .B(n4272), .Z(n4274) );
  XOR U4556 ( .A(n4273), .B(n4274), .Z(n4268) );
  XOR U4557 ( .A(n4267), .B(n4268), .Z(n4289) );
  XOR U4558 ( .A(n4290), .B(n4289), .Z(n4291) );
  XNOR U4559 ( .A(n4292), .B(n4291), .Z(n4261) );
  NAND U4560 ( .A(n4251), .B(n4250), .Z(n4255) );
  NAND U4561 ( .A(n4253), .B(n4252), .Z(n4254) );
  NAND U4562 ( .A(n4255), .B(n4254), .Z(n4262) );
  XNOR U4563 ( .A(n4261), .B(n4262), .Z(n4263) );
  XNOR U4564 ( .A(n4264), .B(n4263), .Z(n4295) );
  XNOR U4565 ( .A(n4295), .B(sreg[347]), .Z(n4297) );
  NAND U4566 ( .A(n4256), .B(sreg[346]), .Z(n4260) );
  OR U4567 ( .A(n4258), .B(n4257), .Z(n4259) );
  AND U4568 ( .A(n4260), .B(n4259), .Z(n4296) );
  XOR U4569 ( .A(n4297), .B(n4296), .Z(c[347]) );
  NANDN U4570 ( .A(n4266), .B(n4265), .Z(n4270) );
  NAND U4571 ( .A(n4268), .B(n4267), .Z(n4269) );
  NAND U4572 ( .A(n4270), .B(n4269), .Z(n4331) );
  NANDN U4573 ( .A(n4272), .B(n4271), .Z(n4276) );
  NAND U4574 ( .A(n4274), .B(n4273), .Z(n4275) );
  NAND U4575 ( .A(n4276), .B(n4275), .Z(n4329) );
  XNOR U4576 ( .A(b[7]), .B(a[94]), .Z(n4316) );
  NANDN U4577 ( .A(n4316), .B(n10545), .Z(n4279) );
  NANDN U4578 ( .A(n4277), .B(n10546), .Z(n4278) );
  NAND U4579 ( .A(n4279), .B(n4278), .Z(n4304) );
  XNOR U4580 ( .A(b[3]), .B(a[98]), .Z(n4319) );
  NANDN U4581 ( .A(n4319), .B(n10398), .Z(n4282) );
  NANDN U4582 ( .A(n4280), .B(n10399), .Z(n4281) );
  AND U4583 ( .A(n4282), .B(n4281), .Z(n4305) );
  XNOR U4584 ( .A(n4304), .B(n4305), .Z(n4306) );
  NANDN U4585 ( .A(n527), .B(a[100]), .Z(n4283) );
  XOR U4586 ( .A(n10434), .B(n4283), .Z(n4285) );
  NANDN U4587 ( .A(b[0]), .B(a[99]), .Z(n4284) );
  AND U4588 ( .A(n4285), .B(n4284), .Z(n4312) );
  XOR U4589 ( .A(b[5]), .B(a[96]), .Z(n4325) );
  NAND U4590 ( .A(n4325), .B(n10481), .Z(n4288) );
  NAND U4591 ( .A(n4286), .B(n10482), .Z(n4287) );
  NAND U4592 ( .A(n4288), .B(n4287), .Z(n4310) );
  NANDN U4593 ( .A(n529), .B(a[92]), .Z(n4311) );
  XNOR U4594 ( .A(n4310), .B(n4311), .Z(n4313) );
  XOR U4595 ( .A(n4312), .B(n4313), .Z(n4307) );
  XOR U4596 ( .A(n4306), .B(n4307), .Z(n4328) );
  XOR U4597 ( .A(n4329), .B(n4328), .Z(n4330) );
  XNOR U4598 ( .A(n4331), .B(n4330), .Z(n4300) );
  NAND U4599 ( .A(n4290), .B(n4289), .Z(n4294) );
  NAND U4600 ( .A(n4292), .B(n4291), .Z(n4293) );
  NAND U4601 ( .A(n4294), .B(n4293), .Z(n4301) );
  XNOR U4602 ( .A(n4300), .B(n4301), .Z(n4302) );
  XNOR U4603 ( .A(n4303), .B(n4302), .Z(n4334) );
  XNOR U4604 ( .A(n4334), .B(sreg[348]), .Z(n4336) );
  NAND U4605 ( .A(n4295), .B(sreg[347]), .Z(n4299) );
  OR U4606 ( .A(n4297), .B(n4296), .Z(n4298) );
  AND U4607 ( .A(n4299), .B(n4298), .Z(n4335) );
  XOR U4608 ( .A(n4336), .B(n4335), .Z(c[348]) );
  NANDN U4609 ( .A(n4305), .B(n4304), .Z(n4309) );
  NAND U4610 ( .A(n4307), .B(n4306), .Z(n4308) );
  NAND U4611 ( .A(n4309), .B(n4308), .Z(n4370) );
  NANDN U4612 ( .A(n4311), .B(n4310), .Z(n4315) );
  NAND U4613 ( .A(n4313), .B(n4312), .Z(n4314) );
  NAND U4614 ( .A(n4315), .B(n4314), .Z(n4368) );
  XNOR U4615 ( .A(b[7]), .B(a[95]), .Z(n4355) );
  NANDN U4616 ( .A(n4355), .B(n10545), .Z(n4318) );
  NANDN U4617 ( .A(n4316), .B(n10546), .Z(n4317) );
  NAND U4618 ( .A(n4318), .B(n4317), .Z(n4343) );
  XNOR U4619 ( .A(b[3]), .B(a[99]), .Z(n4358) );
  NANDN U4620 ( .A(n4358), .B(n10398), .Z(n4321) );
  NANDN U4621 ( .A(n4319), .B(n10399), .Z(n4320) );
  AND U4622 ( .A(n4321), .B(n4320), .Z(n4344) );
  XNOR U4623 ( .A(n4343), .B(n4344), .Z(n4345) );
  NANDN U4624 ( .A(n527), .B(a[101]), .Z(n4322) );
  XOR U4625 ( .A(n10434), .B(n4322), .Z(n4324) );
  NANDN U4626 ( .A(b[0]), .B(a[100]), .Z(n4323) );
  AND U4627 ( .A(n4324), .B(n4323), .Z(n4351) );
  XOR U4628 ( .A(b[5]), .B(a[97]), .Z(n4364) );
  NAND U4629 ( .A(n4364), .B(n10481), .Z(n4327) );
  NAND U4630 ( .A(n4325), .B(n10482), .Z(n4326) );
  NAND U4631 ( .A(n4327), .B(n4326), .Z(n4349) );
  NANDN U4632 ( .A(n529), .B(a[93]), .Z(n4350) );
  XNOR U4633 ( .A(n4349), .B(n4350), .Z(n4352) );
  XOR U4634 ( .A(n4351), .B(n4352), .Z(n4346) );
  XOR U4635 ( .A(n4345), .B(n4346), .Z(n4367) );
  XOR U4636 ( .A(n4368), .B(n4367), .Z(n4369) );
  XNOR U4637 ( .A(n4370), .B(n4369), .Z(n4339) );
  NAND U4638 ( .A(n4329), .B(n4328), .Z(n4333) );
  NAND U4639 ( .A(n4331), .B(n4330), .Z(n4332) );
  NAND U4640 ( .A(n4333), .B(n4332), .Z(n4340) );
  XNOR U4641 ( .A(n4339), .B(n4340), .Z(n4341) );
  XNOR U4642 ( .A(n4342), .B(n4341), .Z(n4373) );
  XNOR U4643 ( .A(n4373), .B(sreg[349]), .Z(n4375) );
  NAND U4644 ( .A(n4334), .B(sreg[348]), .Z(n4338) );
  OR U4645 ( .A(n4336), .B(n4335), .Z(n4337) );
  AND U4646 ( .A(n4338), .B(n4337), .Z(n4374) );
  XOR U4647 ( .A(n4375), .B(n4374), .Z(c[349]) );
  NANDN U4648 ( .A(n4344), .B(n4343), .Z(n4348) );
  NAND U4649 ( .A(n4346), .B(n4345), .Z(n4347) );
  NAND U4650 ( .A(n4348), .B(n4347), .Z(n4409) );
  NANDN U4651 ( .A(n4350), .B(n4349), .Z(n4354) );
  NAND U4652 ( .A(n4352), .B(n4351), .Z(n4353) );
  NAND U4653 ( .A(n4354), .B(n4353), .Z(n4407) );
  XNOR U4654 ( .A(b[7]), .B(a[96]), .Z(n4394) );
  NANDN U4655 ( .A(n4394), .B(n10545), .Z(n4357) );
  NANDN U4656 ( .A(n4355), .B(n10546), .Z(n4356) );
  NAND U4657 ( .A(n4357), .B(n4356), .Z(n4382) );
  XNOR U4658 ( .A(b[3]), .B(a[100]), .Z(n4397) );
  NANDN U4659 ( .A(n4397), .B(n10398), .Z(n4360) );
  NANDN U4660 ( .A(n4358), .B(n10399), .Z(n4359) );
  AND U4661 ( .A(n4360), .B(n4359), .Z(n4383) );
  XNOR U4662 ( .A(n4382), .B(n4383), .Z(n4384) );
  NANDN U4663 ( .A(n527), .B(a[102]), .Z(n4361) );
  XOR U4664 ( .A(n10434), .B(n4361), .Z(n4363) );
  NANDN U4665 ( .A(b[0]), .B(a[101]), .Z(n4362) );
  AND U4666 ( .A(n4363), .B(n4362), .Z(n4390) );
  XOR U4667 ( .A(b[5]), .B(a[98]), .Z(n4403) );
  NAND U4668 ( .A(n4403), .B(n10481), .Z(n4366) );
  NAND U4669 ( .A(n4364), .B(n10482), .Z(n4365) );
  NAND U4670 ( .A(n4366), .B(n4365), .Z(n4388) );
  NANDN U4671 ( .A(n529), .B(a[94]), .Z(n4389) );
  XNOR U4672 ( .A(n4388), .B(n4389), .Z(n4391) );
  XOR U4673 ( .A(n4390), .B(n4391), .Z(n4385) );
  XOR U4674 ( .A(n4384), .B(n4385), .Z(n4406) );
  XOR U4675 ( .A(n4407), .B(n4406), .Z(n4408) );
  XNOR U4676 ( .A(n4409), .B(n4408), .Z(n4378) );
  NAND U4677 ( .A(n4368), .B(n4367), .Z(n4372) );
  NAND U4678 ( .A(n4370), .B(n4369), .Z(n4371) );
  NAND U4679 ( .A(n4372), .B(n4371), .Z(n4379) );
  XNOR U4680 ( .A(n4378), .B(n4379), .Z(n4380) );
  XNOR U4681 ( .A(n4381), .B(n4380), .Z(n4412) );
  XNOR U4682 ( .A(n4412), .B(sreg[350]), .Z(n4414) );
  NAND U4683 ( .A(n4373), .B(sreg[349]), .Z(n4377) );
  OR U4684 ( .A(n4375), .B(n4374), .Z(n4376) );
  AND U4685 ( .A(n4377), .B(n4376), .Z(n4413) );
  XOR U4686 ( .A(n4414), .B(n4413), .Z(c[350]) );
  NANDN U4687 ( .A(n4383), .B(n4382), .Z(n4387) );
  NAND U4688 ( .A(n4385), .B(n4384), .Z(n4386) );
  NAND U4689 ( .A(n4387), .B(n4386), .Z(n4448) );
  NANDN U4690 ( .A(n4389), .B(n4388), .Z(n4393) );
  NAND U4691 ( .A(n4391), .B(n4390), .Z(n4392) );
  NAND U4692 ( .A(n4393), .B(n4392), .Z(n4446) );
  XNOR U4693 ( .A(b[7]), .B(a[97]), .Z(n4433) );
  NANDN U4694 ( .A(n4433), .B(n10545), .Z(n4396) );
  NANDN U4695 ( .A(n4394), .B(n10546), .Z(n4395) );
  NAND U4696 ( .A(n4396), .B(n4395), .Z(n4421) );
  XNOR U4697 ( .A(b[3]), .B(a[101]), .Z(n4436) );
  NANDN U4698 ( .A(n4436), .B(n10398), .Z(n4399) );
  NANDN U4699 ( .A(n4397), .B(n10399), .Z(n4398) );
  AND U4700 ( .A(n4399), .B(n4398), .Z(n4422) );
  XNOR U4701 ( .A(n4421), .B(n4422), .Z(n4423) );
  NANDN U4702 ( .A(n527), .B(a[103]), .Z(n4400) );
  XOR U4703 ( .A(n10434), .B(n4400), .Z(n4402) );
  NANDN U4704 ( .A(b[0]), .B(a[102]), .Z(n4401) );
  AND U4705 ( .A(n4402), .B(n4401), .Z(n4429) );
  XOR U4706 ( .A(b[5]), .B(a[99]), .Z(n4442) );
  NAND U4707 ( .A(n4442), .B(n10481), .Z(n4405) );
  NAND U4708 ( .A(n4403), .B(n10482), .Z(n4404) );
  NAND U4709 ( .A(n4405), .B(n4404), .Z(n4427) );
  NANDN U4710 ( .A(n529), .B(a[95]), .Z(n4428) );
  XNOR U4711 ( .A(n4427), .B(n4428), .Z(n4430) );
  XOR U4712 ( .A(n4429), .B(n4430), .Z(n4424) );
  XOR U4713 ( .A(n4423), .B(n4424), .Z(n4445) );
  XOR U4714 ( .A(n4446), .B(n4445), .Z(n4447) );
  XNOR U4715 ( .A(n4448), .B(n4447), .Z(n4417) );
  NAND U4716 ( .A(n4407), .B(n4406), .Z(n4411) );
  NAND U4717 ( .A(n4409), .B(n4408), .Z(n4410) );
  NAND U4718 ( .A(n4411), .B(n4410), .Z(n4418) );
  XNOR U4719 ( .A(n4417), .B(n4418), .Z(n4419) );
  XNOR U4720 ( .A(n4420), .B(n4419), .Z(n4451) );
  XNOR U4721 ( .A(n4451), .B(sreg[351]), .Z(n4453) );
  NAND U4722 ( .A(n4412), .B(sreg[350]), .Z(n4416) );
  OR U4723 ( .A(n4414), .B(n4413), .Z(n4415) );
  AND U4724 ( .A(n4416), .B(n4415), .Z(n4452) );
  XOR U4725 ( .A(n4453), .B(n4452), .Z(c[351]) );
  NANDN U4726 ( .A(n4422), .B(n4421), .Z(n4426) );
  NAND U4727 ( .A(n4424), .B(n4423), .Z(n4425) );
  NAND U4728 ( .A(n4426), .B(n4425), .Z(n4487) );
  NANDN U4729 ( .A(n4428), .B(n4427), .Z(n4432) );
  NAND U4730 ( .A(n4430), .B(n4429), .Z(n4431) );
  NAND U4731 ( .A(n4432), .B(n4431), .Z(n4485) );
  XNOR U4732 ( .A(b[7]), .B(a[98]), .Z(n4472) );
  NANDN U4733 ( .A(n4472), .B(n10545), .Z(n4435) );
  NANDN U4734 ( .A(n4433), .B(n10546), .Z(n4434) );
  NAND U4735 ( .A(n4435), .B(n4434), .Z(n4460) );
  XNOR U4736 ( .A(b[3]), .B(a[102]), .Z(n4475) );
  NANDN U4737 ( .A(n4475), .B(n10398), .Z(n4438) );
  NANDN U4738 ( .A(n4436), .B(n10399), .Z(n4437) );
  AND U4739 ( .A(n4438), .B(n4437), .Z(n4461) );
  XNOR U4740 ( .A(n4460), .B(n4461), .Z(n4462) );
  NANDN U4741 ( .A(n527), .B(a[104]), .Z(n4439) );
  XOR U4742 ( .A(n10434), .B(n4439), .Z(n4441) );
  NANDN U4743 ( .A(b[0]), .B(a[103]), .Z(n4440) );
  AND U4744 ( .A(n4441), .B(n4440), .Z(n4468) );
  XOR U4745 ( .A(b[5]), .B(a[100]), .Z(n4481) );
  NAND U4746 ( .A(n4481), .B(n10481), .Z(n4444) );
  NAND U4747 ( .A(n4442), .B(n10482), .Z(n4443) );
  NAND U4748 ( .A(n4444), .B(n4443), .Z(n4466) );
  NANDN U4749 ( .A(n529), .B(a[96]), .Z(n4467) );
  XNOR U4750 ( .A(n4466), .B(n4467), .Z(n4469) );
  XOR U4751 ( .A(n4468), .B(n4469), .Z(n4463) );
  XOR U4752 ( .A(n4462), .B(n4463), .Z(n4484) );
  XOR U4753 ( .A(n4485), .B(n4484), .Z(n4486) );
  XNOR U4754 ( .A(n4487), .B(n4486), .Z(n4456) );
  NAND U4755 ( .A(n4446), .B(n4445), .Z(n4450) );
  NAND U4756 ( .A(n4448), .B(n4447), .Z(n4449) );
  NAND U4757 ( .A(n4450), .B(n4449), .Z(n4457) );
  XNOR U4758 ( .A(n4456), .B(n4457), .Z(n4458) );
  XNOR U4759 ( .A(n4459), .B(n4458), .Z(n4490) );
  XNOR U4760 ( .A(n4490), .B(sreg[352]), .Z(n4492) );
  NAND U4761 ( .A(n4451), .B(sreg[351]), .Z(n4455) );
  OR U4762 ( .A(n4453), .B(n4452), .Z(n4454) );
  AND U4763 ( .A(n4455), .B(n4454), .Z(n4491) );
  XOR U4764 ( .A(n4492), .B(n4491), .Z(c[352]) );
  NANDN U4765 ( .A(n4461), .B(n4460), .Z(n4465) );
  NAND U4766 ( .A(n4463), .B(n4462), .Z(n4464) );
  NAND U4767 ( .A(n4465), .B(n4464), .Z(n4526) );
  NANDN U4768 ( .A(n4467), .B(n4466), .Z(n4471) );
  NAND U4769 ( .A(n4469), .B(n4468), .Z(n4470) );
  NAND U4770 ( .A(n4471), .B(n4470), .Z(n4524) );
  XNOR U4771 ( .A(b[7]), .B(a[99]), .Z(n4517) );
  NANDN U4772 ( .A(n4517), .B(n10545), .Z(n4474) );
  NANDN U4773 ( .A(n4472), .B(n10546), .Z(n4473) );
  NAND U4774 ( .A(n4474), .B(n4473), .Z(n4499) );
  XNOR U4775 ( .A(b[3]), .B(a[103]), .Z(n4520) );
  NANDN U4776 ( .A(n4520), .B(n10398), .Z(n4477) );
  NANDN U4777 ( .A(n4475), .B(n10399), .Z(n4476) );
  AND U4778 ( .A(n4477), .B(n4476), .Z(n4500) );
  XNOR U4779 ( .A(n4499), .B(n4500), .Z(n4501) );
  NANDN U4780 ( .A(n527), .B(a[105]), .Z(n4478) );
  XOR U4781 ( .A(n10434), .B(n4478), .Z(n4480) );
  NANDN U4782 ( .A(b[0]), .B(a[104]), .Z(n4479) );
  AND U4783 ( .A(n4480), .B(n4479), .Z(n4507) );
  XOR U4784 ( .A(b[5]), .B(a[101]), .Z(n4514) );
  NAND U4785 ( .A(n4514), .B(n10481), .Z(n4483) );
  NAND U4786 ( .A(n4481), .B(n10482), .Z(n4482) );
  NAND U4787 ( .A(n4483), .B(n4482), .Z(n4505) );
  NANDN U4788 ( .A(n529), .B(a[97]), .Z(n4506) );
  XNOR U4789 ( .A(n4505), .B(n4506), .Z(n4508) );
  XOR U4790 ( .A(n4507), .B(n4508), .Z(n4502) );
  XOR U4791 ( .A(n4501), .B(n4502), .Z(n4523) );
  XOR U4792 ( .A(n4524), .B(n4523), .Z(n4525) );
  XNOR U4793 ( .A(n4526), .B(n4525), .Z(n4495) );
  NAND U4794 ( .A(n4485), .B(n4484), .Z(n4489) );
  NAND U4795 ( .A(n4487), .B(n4486), .Z(n4488) );
  NAND U4796 ( .A(n4489), .B(n4488), .Z(n4496) );
  XNOR U4797 ( .A(n4495), .B(n4496), .Z(n4497) );
  XNOR U4798 ( .A(n4498), .B(n4497), .Z(n4529) );
  XNOR U4799 ( .A(n4529), .B(sreg[353]), .Z(n4531) );
  NAND U4800 ( .A(n4490), .B(sreg[352]), .Z(n4494) );
  OR U4801 ( .A(n4492), .B(n4491), .Z(n4493) );
  AND U4802 ( .A(n4494), .B(n4493), .Z(n4530) );
  XOR U4803 ( .A(n4531), .B(n4530), .Z(c[353]) );
  NANDN U4804 ( .A(n4500), .B(n4499), .Z(n4504) );
  NAND U4805 ( .A(n4502), .B(n4501), .Z(n4503) );
  NAND U4806 ( .A(n4504), .B(n4503), .Z(n4565) );
  NANDN U4807 ( .A(n4506), .B(n4505), .Z(n4510) );
  NAND U4808 ( .A(n4508), .B(n4507), .Z(n4509) );
  NAND U4809 ( .A(n4510), .B(n4509), .Z(n4563) );
  NANDN U4810 ( .A(n527), .B(a[106]), .Z(n4511) );
  XOR U4811 ( .A(n10434), .B(n4511), .Z(n4513) );
  NANDN U4812 ( .A(b[0]), .B(a[105]), .Z(n4512) );
  AND U4813 ( .A(n4513), .B(n4512), .Z(n4546) );
  XOR U4814 ( .A(b[5]), .B(a[102]), .Z(n4559) );
  NAND U4815 ( .A(n4559), .B(n10481), .Z(n4516) );
  NAND U4816 ( .A(n4514), .B(n10482), .Z(n4515) );
  NAND U4817 ( .A(n4516), .B(n4515), .Z(n4544) );
  NANDN U4818 ( .A(n529), .B(a[98]), .Z(n4545) );
  XNOR U4819 ( .A(n4544), .B(n4545), .Z(n4547) );
  XOR U4820 ( .A(n4546), .B(n4547), .Z(n4540) );
  XNOR U4821 ( .A(b[7]), .B(a[100]), .Z(n4550) );
  NANDN U4822 ( .A(n4550), .B(n10545), .Z(n4519) );
  NANDN U4823 ( .A(n4517), .B(n10546), .Z(n4518) );
  NAND U4824 ( .A(n4519), .B(n4518), .Z(n4538) );
  XNOR U4825 ( .A(b[3]), .B(a[104]), .Z(n4553) );
  NANDN U4826 ( .A(n4553), .B(n10398), .Z(n4522) );
  NANDN U4827 ( .A(n4520), .B(n10399), .Z(n4521) );
  AND U4828 ( .A(n4522), .B(n4521), .Z(n4539) );
  XNOR U4829 ( .A(n4538), .B(n4539), .Z(n4541) );
  XOR U4830 ( .A(n4540), .B(n4541), .Z(n4562) );
  XOR U4831 ( .A(n4563), .B(n4562), .Z(n4564) );
  XNOR U4832 ( .A(n4565), .B(n4564), .Z(n4534) );
  NAND U4833 ( .A(n4524), .B(n4523), .Z(n4528) );
  NAND U4834 ( .A(n4526), .B(n4525), .Z(n4527) );
  NAND U4835 ( .A(n4528), .B(n4527), .Z(n4535) );
  XNOR U4836 ( .A(n4534), .B(n4535), .Z(n4536) );
  XNOR U4837 ( .A(n4537), .B(n4536), .Z(n4568) );
  XNOR U4838 ( .A(n4568), .B(sreg[354]), .Z(n4570) );
  NAND U4839 ( .A(n4529), .B(sreg[353]), .Z(n4533) );
  OR U4840 ( .A(n4531), .B(n4530), .Z(n4532) );
  AND U4841 ( .A(n4533), .B(n4532), .Z(n4569) );
  XOR U4842 ( .A(n4570), .B(n4569), .Z(c[354]) );
  NANDN U4843 ( .A(n4539), .B(n4538), .Z(n4543) );
  NAND U4844 ( .A(n4541), .B(n4540), .Z(n4542) );
  NAND U4845 ( .A(n4543), .B(n4542), .Z(n4604) );
  NANDN U4846 ( .A(n4545), .B(n4544), .Z(n4549) );
  NAND U4847 ( .A(n4547), .B(n4546), .Z(n4548) );
  NAND U4848 ( .A(n4549), .B(n4548), .Z(n4602) );
  XNOR U4849 ( .A(b[7]), .B(a[101]), .Z(n4589) );
  NANDN U4850 ( .A(n4589), .B(n10545), .Z(n4552) );
  NANDN U4851 ( .A(n4550), .B(n10546), .Z(n4551) );
  NAND U4852 ( .A(n4552), .B(n4551), .Z(n4577) );
  XNOR U4853 ( .A(b[3]), .B(a[105]), .Z(n4592) );
  NANDN U4854 ( .A(n4592), .B(n10398), .Z(n4555) );
  NANDN U4855 ( .A(n4553), .B(n10399), .Z(n4554) );
  AND U4856 ( .A(n4555), .B(n4554), .Z(n4578) );
  XNOR U4857 ( .A(n4577), .B(n4578), .Z(n4579) );
  NANDN U4858 ( .A(n527), .B(a[107]), .Z(n4556) );
  XOR U4859 ( .A(n10434), .B(n4556), .Z(n4558) );
  NANDN U4860 ( .A(b[0]), .B(a[106]), .Z(n4557) );
  AND U4861 ( .A(n4558), .B(n4557), .Z(n4585) );
  XOR U4862 ( .A(b[5]), .B(a[103]), .Z(n4598) );
  NAND U4863 ( .A(n4598), .B(n10481), .Z(n4561) );
  NAND U4864 ( .A(n4559), .B(n10482), .Z(n4560) );
  NAND U4865 ( .A(n4561), .B(n4560), .Z(n4583) );
  NANDN U4866 ( .A(n529), .B(a[99]), .Z(n4584) );
  XNOR U4867 ( .A(n4583), .B(n4584), .Z(n4586) );
  XOR U4868 ( .A(n4585), .B(n4586), .Z(n4580) );
  XOR U4869 ( .A(n4579), .B(n4580), .Z(n4601) );
  XOR U4870 ( .A(n4602), .B(n4601), .Z(n4603) );
  XNOR U4871 ( .A(n4604), .B(n4603), .Z(n4573) );
  NAND U4872 ( .A(n4563), .B(n4562), .Z(n4567) );
  NAND U4873 ( .A(n4565), .B(n4564), .Z(n4566) );
  NAND U4874 ( .A(n4567), .B(n4566), .Z(n4574) );
  XNOR U4875 ( .A(n4573), .B(n4574), .Z(n4575) );
  XNOR U4876 ( .A(n4576), .B(n4575), .Z(n4607) );
  XNOR U4877 ( .A(n4607), .B(sreg[355]), .Z(n4609) );
  NAND U4878 ( .A(n4568), .B(sreg[354]), .Z(n4572) );
  OR U4879 ( .A(n4570), .B(n4569), .Z(n4571) );
  AND U4880 ( .A(n4572), .B(n4571), .Z(n4608) );
  XOR U4881 ( .A(n4609), .B(n4608), .Z(c[355]) );
  NANDN U4882 ( .A(n4578), .B(n4577), .Z(n4582) );
  NAND U4883 ( .A(n4580), .B(n4579), .Z(n4581) );
  NAND U4884 ( .A(n4582), .B(n4581), .Z(n4643) );
  NANDN U4885 ( .A(n4584), .B(n4583), .Z(n4588) );
  NAND U4886 ( .A(n4586), .B(n4585), .Z(n4587) );
  NAND U4887 ( .A(n4588), .B(n4587), .Z(n4641) );
  XNOR U4888 ( .A(b[7]), .B(a[102]), .Z(n4628) );
  NANDN U4889 ( .A(n4628), .B(n10545), .Z(n4591) );
  NANDN U4890 ( .A(n4589), .B(n10546), .Z(n4590) );
  NAND U4891 ( .A(n4591), .B(n4590), .Z(n4616) );
  XNOR U4892 ( .A(b[3]), .B(a[106]), .Z(n4631) );
  NANDN U4893 ( .A(n4631), .B(n10398), .Z(n4594) );
  NANDN U4894 ( .A(n4592), .B(n10399), .Z(n4593) );
  AND U4895 ( .A(n4594), .B(n4593), .Z(n4617) );
  XNOR U4896 ( .A(n4616), .B(n4617), .Z(n4618) );
  NANDN U4897 ( .A(n527), .B(a[108]), .Z(n4595) );
  XOR U4898 ( .A(n10434), .B(n4595), .Z(n4597) );
  NANDN U4899 ( .A(b[0]), .B(a[107]), .Z(n4596) );
  AND U4900 ( .A(n4597), .B(n4596), .Z(n4624) );
  XOR U4901 ( .A(b[5]), .B(a[104]), .Z(n4637) );
  NAND U4902 ( .A(n4637), .B(n10481), .Z(n4600) );
  NAND U4903 ( .A(n4598), .B(n10482), .Z(n4599) );
  NAND U4904 ( .A(n4600), .B(n4599), .Z(n4622) );
  NANDN U4905 ( .A(n529), .B(a[100]), .Z(n4623) );
  XNOR U4906 ( .A(n4622), .B(n4623), .Z(n4625) );
  XOR U4907 ( .A(n4624), .B(n4625), .Z(n4619) );
  XOR U4908 ( .A(n4618), .B(n4619), .Z(n4640) );
  XOR U4909 ( .A(n4641), .B(n4640), .Z(n4642) );
  XNOR U4910 ( .A(n4643), .B(n4642), .Z(n4612) );
  NAND U4911 ( .A(n4602), .B(n4601), .Z(n4606) );
  NAND U4912 ( .A(n4604), .B(n4603), .Z(n4605) );
  NAND U4913 ( .A(n4606), .B(n4605), .Z(n4613) );
  XNOR U4914 ( .A(n4612), .B(n4613), .Z(n4614) );
  XNOR U4915 ( .A(n4615), .B(n4614), .Z(n4646) );
  XNOR U4916 ( .A(n4646), .B(sreg[356]), .Z(n4648) );
  NAND U4917 ( .A(n4607), .B(sreg[355]), .Z(n4611) );
  OR U4918 ( .A(n4609), .B(n4608), .Z(n4610) );
  AND U4919 ( .A(n4611), .B(n4610), .Z(n4647) );
  XOR U4920 ( .A(n4648), .B(n4647), .Z(c[356]) );
  NANDN U4921 ( .A(n4617), .B(n4616), .Z(n4621) );
  NAND U4922 ( .A(n4619), .B(n4618), .Z(n4620) );
  NAND U4923 ( .A(n4621), .B(n4620), .Z(n4682) );
  NANDN U4924 ( .A(n4623), .B(n4622), .Z(n4627) );
  NAND U4925 ( .A(n4625), .B(n4624), .Z(n4626) );
  NAND U4926 ( .A(n4627), .B(n4626), .Z(n4680) );
  XNOR U4927 ( .A(b[7]), .B(a[103]), .Z(n4667) );
  NANDN U4928 ( .A(n4667), .B(n10545), .Z(n4630) );
  NANDN U4929 ( .A(n4628), .B(n10546), .Z(n4629) );
  NAND U4930 ( .A(n4630), .B(n4629), .Z(n4655) );
  XNOR U4931 ( .A(b[3]), .B(a[107]), .Z(n4670) );
  NANDN U4932 ( .A(n4670), .B(n10398), .Z(n4633) );
  NANDN U4933 ( .A(n4631), .B(n10399), .Z(n4632) );
  AND U4934 ( .A(n4633), .B(n4632), .Z(n4656) );
  XNOR U4935 ( .A(n4655), .B(n4656), .Z(n4657) );
  NANDN U4936 ( .A(n527), .B(a[109]), .Z(n4634) );
  XOR U4937 ( .A(n10434), .B(n4634), .Z(n4636) );
  NANDN U4938 ( .A(b[0]), .B(a[108]), .Z(n4635) );
  AND U4939 ( .A(n4636), .B(n4635), .Z(n4663) );
  XOR U4940 ( .A(b[5]), .B(a[105]), .Z(n4676) );
  NAND U4941 ( .A(n4676), .B(n10481), .Z(n4639) );
  NAND U4942 ( .A(n4637), .B(n10482), .Z(n4638) );
  NAND U4943 ( .A(n4639), .B(n4638), .Z(n4661) );
  NANDN U4944 ( .A(n529), .B(a[101]), .Z(n4662) );
  XNOR U4945 ( .A(n4661), .B(n4662), .Z(n4664) );
  XOR U4946 ( .A(n4663), .B(n4664), .Z(n4658) );
  XOR U4947 ( .A(n4657), .B(n4658), .Z(n4679) );
  XOR U4948 ( .A(n4680), .B(n4679), .Z(n4681) );
  XNOR U4949 ( .A(n4682), .B(n4681), .Z(n4651) );
  NAND U4950 ( .A(n4641), .B(n4640), .Z(n4645) );
  NAND U4951 ( .A(n4643), .B(n4642), .Z(n4644) );
  NAND U4952 ( .A(n4645), .B(n4644), .Z(n4652) );
  XNOR U4953 ( .A(n4651), .B(n4652), .Z(n4653) );
  XNOR U4954 ( .A(n4654), .B(n4653), .Z(n4685) );
  XNOR U4955 ( .A(n4685), .B(sreg[357]), .Z(n4687) );
  NAND U4956 ( .A(n4646), .B(sreg[356]), .Z(n4650) );
  OR U4957 ( .A(n4648), .B(n4647), .Z(n4649) );
  AND U4958 ( .A(n4650), .B(n4649), .Z(n4686) );
  XOR U4959 ( .A(n4687), .B(n4686), .Z(c[357]) );
  NANDN U4960 ( .A(n4656), .B(n4655), .Z(n4660) );
  NAND U4961 ( .A(n4658), .B(n4657), .Z(n4659) );
  NAND U4962 ( .A(n4660), .B(n4659), .Z(n4721) );
  NANDN U4963 ( .A(n4662), .B(n4661), .Z(n4666) );
  NAND U4964 ( .A(n4664), .B(n4663), .Z(n4665) );
  NAND U4965 ( .A(n4666), .B(n4665), .Z(n4719) );
  XNOR U4966 ( .A(b[7]), .B(a[104]), .Z(n4706) );
  NANDN U4967 ( .A(n4706), .B(n10545), .Z(n4669) );
  NANDN U4968 ( .A(n4667), .B(n10546), .Z(n4668) );
  NAND U4969 ( .A(n4669), .B(n4668), .Z(n4694) );
  XNOR U4970 ( .A(b[3]), .B(a[108]), .Z(n4709) );
  NANDN U4971 ( .A(n4709), .B(n10398), .Z(n4672) );
  NANDN U4972 ( .A(n4670), .B(n10399), .Z(n4671) );
  AND U4973 ( .A(n4672), .B(n4671), .Z(n4695) );
  XNOR U4974 ( .A(n4694), .B(n4695), .Z(n4696) );
  NANDN U4975 ( .A(n527), .B(a[110]), .Z(n4673) );
  XOR U4976 ( .A(n10434), .B(n4673), .Z(n4675) );
  NANDN U4977 ( .A(b[0]), .B(a[109]), .Z(n4674) );
  AND U4978 ( .A(n4675), .B(n4674), .Z(n4702) );
  XOR U4979 ( .A(b[5]), .B(a[106]), .Z(n4715) );
  NAND U4980 ( .A(n4715), .B(n10481), .Z(n4678) );
  NAND U4981 ( .A(n4676), .B(n10482), .Z(n4677) );
  NAND U4982 ( .A(n4678), .B(n4677), .Z(n4700) );
  NANDN U4983 ( .A(n529), .B(a[102]), .Z(n4701) );
  XNOR U4984 ( .A(n4700), .B(n4701), .Z(n4703) );
  XOR U4985 ( .A(n4702), .B(n4703), .Z(n4697) );
  XOR U4986 ( .A(n4696), .B(n4697), .Z(n4718) );
  XOR U4987 ( .A(n4719), .B(n4718), .Z(n4720) );
  XNOR U4988 ( .A(n4721), .B(n4720), .Z(n4690) );
  NAND U4989 ( .A(n4680), .B(n4679), .Z(n4684) );
  NAND U4990 ( .A(n4682), .B(n4681), .Z(n4683) );
  NAND U4991 ( .A(n4684), .B(n4683), .Z(n4691) );
  XNOR U4992 ( .A(n4690), .B(n4691), .Z(n4692) );
  XNOR U4993 ( .A(n4693), .B(n4692), .Z(n4724) );
  XNOR U4994 ( .A(n4724), .B(sreg[358]), .Z(n4726) );
  NAND U4995 ( .A(n4685), .B(sreg[357]), .Z(n4689) );
  OR U4996 ( .A(n4687), .B(n4686), .Z(n4688) );
  AND U4997 ( .A(n4689), .B(n4688), .Z(n4725) );
  XOR U4998 ( .A(n4726), .B(n4725), .Z(c[358]) );
  NANDN U4999 ( .A(n4695), .B(n4694), .Z(n4699) );
  NAND U5000 ( .A(n4697), .B(n4696), .Z(n4698) );
  NAND U5001 ( .A(n4699), .B(n4698), .Z(n4760) );
  NANDN U5002 ( .A(n4701), .B(n4700), .Z(n4705) );
  NAND U5003 ( .A(n4703), .B(n4702), .Z(n4704) );
  NAND U5004 ( .A(n4705), .B(n4704), .Z(n4758) );
  XNOR U5005 ( .A(b[7]), .B(a[105]), .Z(n4745) );
  NANDN U5006 ( .A(n4745), .B(n10545), .Z(n4708) );
  NANDN U5007 ( .A(n4706), .B(n10546), .Z(n4707) );
  NAND U5008 ( .A(n4708), .B(n4707), .Z(n4733) );
  XNOR U5009 ( .A(b[3]), .B(a[109]), .Z(n4748) );
  NANDN U5010 ( .A(n4748), .B(n10398), .Z(n4711) );
  NANDN U5011 ( .A(n4709), .B(n10399), .Z(n4710) );
  AND U5012 ( .A(n4711), .B(n4710), .Z(n4734) );
  XNOR U5013 ( .A(n4733), .B(n4734), .Z(n4735) );
  NANDN U5014 ( .A(n527), .B(a[111]), .Z(n4712) );
  XOR U5015 ( .A(n10434), .B(n4712), .Z(n4714) );
  NANDN U5016 ( .A(b[0]), .B(a[110]), .Z(n4713) );
  AND U5017 ( .A(n4714), .B(n4713), .Z(n4741) );
  XOR U5018 ( .A(b[5]), .B(a[107]), .Z(n4754) );
  NAND U5019 ( .A(n4754), .B(n10481), .Z(n4717) );
  NAND U5020 ( .A(n4715), .B(n10482), .Z(n4716) );
  NAND U5021 ( .A(n4717), .B(n4716), .Z(n4739) );
  NANDN U5022 ( .A(n529), .B(a[103]), .Z(n4740) );
  XNOR U5023 ( .A(n4739), .B(n4740), .Z(n4742) );
  XOR U5024 ( .A(n4741), .B(n4742), .Z(n4736) );
  XOR U5025 ( .A(n4735), .B(n4736), .Z(n4757) );
  XOR U5026 ( .A(n4758), .B(n4757), .Z(n4759) );
  XNOR U5027 ( .A(n4760), .B(n4759), .Z(n4729) );
  NAND U5028 ( .A(n4719), .B(n4718), .Z(n4723) );
  NAND U5029 ( .A(n4721), .B(n4720), .Z(n4722) );
  NAND U5030 ( .A(n4723), .B(n4722), .Z(n4730) );
  XNOR U5031 ( .A(n4729), .B(n4730), .Z(n4731) );
  XNOR U5032 ( .A(n4732), .B(n4731), .Z(n4763) );
  XNOR U5033 ( .A(n4763), .B(sreg[359]), .Z(n4765) );
  NAND U5034 ( .A(n4724), .B(sreg[358]), .Z(n4728) );
  OR U5035 ( .A(n4726), .B(n4725), .Z(n4727) );
  AND U5036 ( .A(n4728), .B(n4727), .Z(n4764) );
  XOR U5037 ( .A(n4765), .B(n4764), .Z(c[359]) );
  NANDN U5038 ( .A(n4734), .B(n4733), .Z(n4738) );
  NAND U5039 ( .A(n4736), .B(n4735), .Z(n4737) );
  NAND U5040 ( .A(n4738), .B(n4737), .Z(n4799) );
  NANDN U5041 ( .A(n4740), .B(n4739), .Z(n4744) );
  NAND U5042 ( .A(n4742), .B(n4741), .Z(n4743) );
  NAND U5043 ( .A(n4744), .B(n4743), .Z(n4797) );
  XNOR U5044 ( .A(b[7]), .B(a[106]), .Z(n4784) );
  NANDN U5045 ( .A(n4784), .B(n10545), .Z(n4747) );
  NANDN U5046 ( .A(n4745), .B(n10546), .Z(n4746) );
  NAND U5047 ( .A(n4747), .B(n4746), .Z(n4772) );
  XNOR U5048 ( .A(b[3]), .B(a[110]), .Z(n4787) );
  NANDN U5049 ( .A(n4787), .B(n10398), .Z(n4750) );
  NANDN U5050 ( .A(n4748), .B(n10399), .Z(n4749) );
  AND U5051 ( .A(n4750), .B(n4749), .Z(n4773) );
  XNOR U5052 ( .A(n4772), .B(n4773), .Z(n4774) );
  NANDN U5053 ( .A(n527), .B(a[112]), .Z(n4751) );
  XOR U5054 ( .A(n10434), .B(n4751), .Z(n4753) );
  NANDN U5055 ( .A(b[0]), .B(a[111]), .Z(n4752) );
  AND U5056 ( .A(n4753), .B(n4752), .Z(n4780) );
  XOR U5057 ( .A(b[5]), .B(a[108]), .Z(n4793) );
  NAND U5058 ( .A(n4793), .B(n10481), .Z(n4756) );
  NAND U5059 ( .A(n4754), .B(n10482), .Z(n4755) );
  NAND U5060 ( .A(n4756), .B(n4755), .Z(n4778) );
  NANDN U5061 ( .A(n529), .B(a[104]), .Z(n4779) );
  XNOR U5062 ( .A(n4778), .B(n4779), .Z(n4781) );
  XOR U5063 ( .A(n4780), .B(n4781), .Z(n4775) );
  XOR U5064 ( .A(n4774), .B(n4775), .Z(n4796) );
  XOR U5065 ( .A(n4797), .B(n4796), .Z(n4798) );
  XNOR U5066 ( .A(n4799), .B(n4798), .Z(n4768) );
  NAND U5067 ( .A(n4758), .B(n4757), .Z(n4762) );
  NAND U5068 ( .A(n4760), .B(n4759), .Z(n4761) );
  NAND U5069 ( .A(n4762), .B(n4761), .Z(n4769) );
  XNOR U5070 ( .A(n4768), .B(n4769), .Z(n4770) );
  XNOR U5071 ( .A(n4771), .B(n4770), .Z(n4802) );
  XNOR U5072 ( .A(n4802), .B(sreg[360]), .Z(n4804) );
  NAND U5073 ( .A(n4763), .B(sreg[359]), .Z(n4767) );
  OR U5074 ( .A(n4765), .B(n4764), .Z(n4766) );
  AND U5075 ( .A(n4767), .B(n4766), .Z(n4803) );
  XOR U5076 ( .A(n4804), .B(n4803), .Z(c[360]) );
  NANDN U5077 ( .A(n4773), .B(n4772), .Z(n4777) );
  NAND U5078 ( .A(n4775), .B(n4774), .Z(n4776) );
  NAND U5079 ( .A(n4777), .B(n4776), .Z(n4838) );
  NANDN U5080 ( .A(n4779), .B(n4778), .Z(n4783) );
  NAND U5081 ( .A(n4781), .B(n4780), .Z(n4782) );
  NAND U5082 ( .A(n4783), .B(n4782), .Z(n4836) );
  XNOR U5083 ( .A(b[7]), .B(a[107]), .Z(n4823) );
  NANDN U5084 ( .A(n4823), .B(n10545), .Z(n4786) );
  NANDN U5085 ( .A(n4784), .B(n10546), .Z(n4785) );
  NAND U5086 ( .A(n4786), .B(n4785), .Z(n4811) );
  XNOR U5087 ( .A(b[3]), .B(a[111]), .Z(n4826) );
  NANDN U5088 ( .A(n4826), .B(n10398), .Z(n4789) );
  NANDN U5089 ( .A(n4787), .B(n10399), .Z(n4788) );
  AND U5090 ( .A(n4789), .B(n4788), .Z(n4812) );
  XNOR U5091 ( .A(n4811), .B(n4812), .Z(n4813) );
  NANDN U5092 ( .A(n527), .B(a[113]), .Z(n4790) );
  XOR U5093 ( .A(n10434), .B(n4790), .Z(n4792) );
  NANDN U5094 ( .A(b[0]), .B(a[112]), .Z(n4791) );
  AND U5095 ( .A(n4792), .B(n4791), .Z(n4819) );
  XOR U5096 ( .A(b[5]), .B(a[109]), .Z(n4832) );
  NAND U5097 ( .A(n4832), .B(n10481), .Z(n4795) );
  NAND U5098 ( .A(n4793), .B(n10482), .Z(n4794) );
  NAND U5099 ( .A(n4795), .B(n4794), .Z(n4817) );
  NANDN U5100 ( .A(n529), .B(a[105]), .Z(n4818) );
  XNOR U5101 ( .A(n4817), .B(n4818), .Z(n4820) );
  XOR U5102 ( .A(n4819), .B(n4820), .Z(n4814) );
  XOR U5103 ( .A(n4813), .B(n4814), .Z(n4835) );
  XOR U5104 ( .A(n4836), .B(n4835), .Z(n4837) );
  XNOR U5105 ( .A(n4838), .B(n4837), .Z(n4807) );
  NAND U5106 ( .A(n4797), .B(n4796), .Z(n4801) );
  NAND U5107 ( .A(n4799), .B(n4798), .Z(n4800) );
  NAND U5108 ( .A(n4801), .B(n4800), .Z(n4808) );
  XNOR U5109 ( .A(n4807), .B(n4808), .Z(n4809) );
  XNOR U5110 ( .A(n4810), .B(n4809), .Z(n4841) );
  XNOR U5111 ( .A(n4841), .B(sreg[361]), .Z(n4843) );
  NAND U5112 ( .A(n4802), .B(sreg[360]), .Z(n4806) );
  OR U5113 ( .A(n4804), .B(n4803), .Z(n4805) );
  AND U5114 ( .A(n4806), .B(n4805), .Z(n4842) );
  XOR U5115 ( .A(n4843), .B(n4842), .Z(c[361]) );
  NANDN U5116 ( .A(n4812), .B(n4811), .Z(n4816) );
  NAND U5117 ( .A(n4814), .B(n4813), .Z(n4815) );
  NAND U5118 ( .A(n4816), .B(n4815), .Z(n4877) );
  NANDN U5119 ( .A(n4818), .B(n4817), .Z(n4822) );
  NAND U5120 ( .A(n4820), .B(n4819), .Z(n4821) );
  NAND U5121 ( .A(n4822), .B(n4821), .Z(n4875) );
  XNOR U5122 ( .A(b[7]), .B(a[108]), .Z(n4862) );
  NANDN U5123 ( .A(n4862), .B(n10545), .Z(n4825) );
  NANDN U5124 ( .A(n4823), .B(n10546), .Z(n4824) );
  NAND U5125 ( .A(n4825), .B(n4824), .Z(n4850) );
  XNOR U5126 ( .A(b[3]), .B(a[112]), .Z(n4865) );
  NANDN U5127 ( .A(n4865), .B(n10398), .Z(n4828) );
  NANDN U5128 ( .A(n4826), .B(n10399), .Z(n4827) );
  AND U5129 ( .A(n4828), .B(n4827), .Z(n4851) );
  XNOR U5130 ( .A(n4850), .B(n4851), .Z(n4852) );
  NANDN U5131 ( .A(n527), .B(a[114]), .Z(n4829) );
  XOR U5132 ( .A(n10434), .B(n4829), .Z(n4831) );
  NANDN U5133 ( .A(b[0]), .B(a[113]), .Z(n4830) );
  AND U5134 ( .A(n4831), .B(n4830), .Z(n4858) );
  XOR U5135 ( .A(b[5]), .B(a[110]), .Z(n4871) );
  NAND U5136 ( .A(n4871), .B(n10481), .Z(n4834) );
  NAND U5137 ( .A(n4832), .B(n10482), .Z(n4833) );
  NAND U5138 ( .A(n4834), .B(n4833), .Z(n4856) );
  NANDN U5139 ( .A(n529), .B(a[106]), .Z(n4857) );
  XNOR U5140 ( .A(n4856), .B(n4857), .Z(n4859) );
  XOR U5141 ( .A(n4858), .B(n4859), .Z(n4853) );
  XOR U5142 ( .A(n4852), .B(n4853), .Z(n4874) );
  XOR U5143 ( .A(n4875), .B(n4874), .Z(n4876) );
  XNOR U5144 ( .A(n4877), .B(n4876), .Z(n4846) );
  NAND U5145 ( .A(n4836), .B(n4835), .Z(n4840) );
  NAND U5146 ( .A(n4838), .B(n4837), .Z(n4839) );
  NAND U5147 ( .A(n4840), .B(n4839), .Z(n4847) );
  XNOR U5148 ( .A(n4846), .B(n4847), .Z(n4848) );
  XNOR U5149 ( .A(n4849), .B(n4848), .Z(n4880) );
  XNOR U5150 ( .A(n4880), .B(sreg[362]), .Z(n4882) );
  NAND U5151 ( .A(n4841), .B(sreg[361]), .Z(n4845) );
  OR U5152 ( .A(n4843), .B(n4842), .Z(n4844) );
  AND U5153 ( .A(n4845), .B(n4844), .Z(n4881) );
  XOR U5154 ( .A(n4882), .B(n4881), .Z(c[362]) );
  NANDN U5155 ( .A(n4851), .B(n4850), .Z(n4855) );
  NAND U5156 ( .A(n4853), .B(n4852), .Z(n4854) );
  NAND U5157 ( .A(n4855), .B(n4854), .Z(n4916) );
  NANDN U5158 ( .A(n4857), .B(n4856), .Z(n4861) );
  NAND U5159 ( .A(n4859), .B(n4858), .Z(n4860) );
  NAND U5160 ( .A(n4861), .B(n4860), .Z(n4914) );
  XNOR U5161 ( .A(b[7]), .B(a[109]), .Z(n4901) );
  NANDN U5162 ( .A(n4901), .B(n10545), .Z(n4864) );
  NANDN U5163 ( .A(n4862), .B(n10546), .Z(n4863) );
  NAND U5164 ( .A(n4864), .B(n4863), .Z(n4889) );
  XNOR U5165 ( .A(b[3]), .B(a[113]), .Z(n4904) );
  NANDN U5166 ( .A(n4904), .B(n10398), .Z(n4867) );
  NANDN U5167 ( .A(n4865), .B(n10399), .Z(n4866) );
  AND U5168 ( .A(n4867), .B(n4866), .Z(n4890) );
  XNOR U5169 ( .A(n4889), .B(n4890), .Z(n4891) );
  NANDN U5170 ( .A(n527), .B(a[115]), .Z(n4868) );
  XOR U5171 ( .A(n10434), .B(n4868), .Z(n4870) );
  NANDN U5172 ( .A(b[0]), .B(a[114]), .Z(n4869) );
  AND U5173 ( .A(n4870), .B(n4869), .Z(n4897) );
  XOR U5174 ( .A(b[5]), .B(a[111]), .Z(n4910) );
  NAND U5175 ( .A(n4910), .B(n10481), .Z(n4873) );
  NAND U5176 ( .A(n4871), .B(n10482), .Z(n4872) );
  NAND U5177 ( .A(n4873), .B(n4872), .Z(n4895) );
  NANDN U5178 ( .A(n529), .B(a[107]), .Z(n4896) );
  XNOR U5179 ( .A(n4895), .B(n4896), .Z(n4898) );
  XOR U5180 ( .A(n4897), .B(n4898), .Z(n4892) );
  XOR U5181 ( .A(n4891), .B(n4892), .Z(n4913) );
  XOR U5182 ( .A(n4914), .B(n4913), .Z(n4915) );
  XNOR U5183 ( .A(n4916), .B(n4915), .Z(n4885) );
  NAND U5184 ( .A(n4875), .B(n4874), .Z(n4879) );
  NAND U5185 ( .A(n4877), .B(n4876), .Z(n4878) );
  NAND U5186 ( .A(n4879), .B(n4878), .Z(n4886) );
  XNOR U5187 ( .A(n4885), .B(n4886), .Z(n4887) );
  XNOR U5188 ( .A(n4888), .B(n4887), .Z(n4919) );
  XNOR U5189 ( .A(n4919), .B(sreg[363]), .Z(n4921) );
  NAND U5190 ( .A(n4880), .B(sreg[362]), .Z(n4884) );
  OR U5191 ( .A(n4882), .B(n4881), .Z(n4883) );
  AND U5192 ( .A(n4884), .B(n4883), .Z(n4920) );
  XOR U5193 ( .A(n4921), .B(n4920), .Z(c[363]) );
  NANDN U5194 ( .A(n4890), .B(n4889), .Z(n4894) );
  NAND U5195 ( .A(n4892), .B(n4891), .Z(n4893) );
  NAND U5196 ( .A(n4894), .B(n4893), .Z(n4955) );
  NANDN U5197 ( .A(n4896), .B(n4895), .Z(n4900) );
  NAND U5198 ( .A(n4898), .B(n4897), .Z(n4899) );
  NAND U5199 ( .A(n4900), .B(n4899), .Z(n4953) );
  XNOR U5200 ( .A(b[7]), .B(a[110]), .Z(n4940) );
  NANDN U5201 ( .A(n4940), .B(n10545), .Z(n4903) );
  NANDN U5202 ( .A(n4901), .B(n10546), .Z(n4902) );
  NAND U5203 ( .A(n4903), .B(n4902), .Z(n4928) );
  XNOR U5204 ( .A(b[3]), .B(a[114]), .Z(n4943) );
  NANDN U5205 ( .A(n4943), .B(n10398), .Z(n4906) );
  NANDN U5206 ( .A(n4904), .B(n10399), .Z(n4905) );
  AND U5207 ( .A(n4906), .B(n4905), .Z(n4929) );
  XNOR U5208 ( .A(n4928), .B(n4929), .Z(n4930) );
  NANDN U5209 ( .A(n527), .B(a[116]), .Z(n4907) );
  XOR U5210 ( .A(n10434), .B(n4907), .Z(n4909) );
  NANDN U5211 ( .A(b[0]), .B(a[115]), .Z(n4908) );
  AND U5212 ( .A(n4909), .B(n4908), .Z(n4936) );
  XOR U5213 ( .A(b[5]), .B(a[112]), .Z(n4949) );
  NAND U5214 ( .A(n4949), .B(n10481), .Z(n4912) );
  NAND U5215 ( .A(n4910), .B(n10482), .Z(n4911) );
  NAND U5216 ( .A(n4912), .B(n4911), .Z(n4934) );
  NANDN U5217 ( .A(n529), .B(a[108]), .Z(n4935) );
  XNOR U5218 ( .A(n4934), .B(n4935), .Z(n4937) );
  XOR U5219 ( .A(n4936), .B(n4937), .Z(n4931) );
  XOR U5220 ( .A(n4930), .B(n4931), .Z(n4952) );
  XOR U5221 ( .A(n4953), .B(n4952), .Z(n4954) );
  XNOR U5222 ( .A(n4955), .B(n4954), .Z(n4924) );
  NAND U5223 ( .A(n4914), .B(n4913), .Z(n4918) );
  NAND U5224 ( .A(n4916), .B(n4915), .Z(n4917) );
  NAND U5225 ( .A(n4918), .B(n4917), .Z(n4925) );
  XNOR U5226 ( .A(n4924), .B(n4925), .Z(n4926) );
  XNOR U5227 ( .A(n4927), .B(n4926), .Z(n4958) );
  XNOR U5228 ( .A(n4958), .B(sreg[364]), .Z(n4960) );
  NAND U5229 ( .A(n4919), .B(sreg[363]), .Z(n4923) );
  OR U5230 ( .A(n4921), .B(n4920), .Z(n4922) );
  AND U5231 ( .A(n4923), .B(n4922), .Z(n4959) );
  XOR U5232 ( .A(n4960), .B(n4959), .Z(c[364]) );
  NANDN U5233 ( .A(n4929), .B(n4928), .Z(n4933) );
  NAND U5234 ( .A(n4931), .B(n4930), .Z(n4932) );
  NAND U5235 ( .A(n4933), .B(n4932), .Z(n4994) );
  NANDN U5236 ( .A(n4935), .B(n4934), .Z(n4939) );
  NAND U5237 ( .A(n4937), .B(n4936), .Z(n4938) );
  NAND U5238 ( .A(n4939), .B(n4938), .Z(n4992) );
  XNOR U5239 ( .A(b[7]), .B(a[111]), .Z(n4979) );
  NANDN U5240 ( .A(n4979), .B(n10545), .Z(n4942) );
  NANDN U5241 ( .A(n4940), .B(n10546), .Z(n4941) );
  NAND U5242 ( .A(n4942), .B(n4941), .Z(n4967) );
  XNOR U5243 ( .A(b[3]), .B(a[115]), .Z(n4982) );
  NANDN U5244 ( .A(n4982), .B(n10398), .Z(n4945) );
  NANDN U5245 ( .A(n4943), .B(n10399), .Z(n4944) );
  AND U5246 ( .A(n4945), .B(n4944), .Z(n4968) );
  XNOR U5247 ( .A(n4967), .B(n4968), .Z(n4969) );
  NANDN U5248 ( .A(n527), .B(a[117]), .Z(n4946) );
  XOR U5249 ( .A(n10434), .B(n4946), .Z(n4948) );
  NANDN U5250 ( .A(b[0]), .B(a[116]), .Z(n4947) );
  AND U5251 ( .A(n4948), .B(n4947), .Z(n4975) );
  XOR U5252 ( .A(b[5]), .B(a[113]), .Z(n4988) );
  NAND U5253 ( .A(n4988), .B(n10481), .Z(n4951) );
  NAND U5254 ( .A(n4949), .B(n10482), .Z(n4950) );
  NAND U5255 ( .A(n4951), .B(n4950), .Z(n4973) );
  NANDN U5256 ( .A(n529), .B(a[109]), .Z(n4974) );
  XNOR U5257 ( .A(n4973), .B(n4974), .Z(n4976) );
  XOR U5258 ( .A(n4975), .B(n4976), .Z(n4970) );
  XOR U5259 ( .A(n4969), .B(n4970), .Z(n4991) );
  XOR U5260 ( .A(n4992), .B(n4991), .Z(n4993) );
  XNOR U5261 ( .A(n4994), .B(n4993), .Z(n4963) );
  NAND U5262 ( .A(n4953), .B(n4952), .Z(n4957) );
  NAND U5263 ( .A(n4955), .B(n4954), .Z(n4956) );
  NAND U5264 ( .A(n4957), .B(n4956), .Z(n4964) );
  XNOR U5265 ( .A(n4963), .B(n4964), .Z(n4965) );
  XNOR U5266 ( .A(n4966), .B(n4965), .Z(n4997) );
  XNOR U5267 ( .A(n4997), .B(sreg[365]), .Z(n4999) );
  NAND U5268 ( .A(n4958), .B(sreg[364]), .Z(n4962) );
  OR U5269 ( .A(n4960), .B(n4959), .Z(n4961) );
  AND U5270 ( .A(n4962), .B(n4961), .Z(n4998) );
  XOR U5271 ( .A(n4999), .B(n4998), .Z(c[365]) );
  NANDN U5272 ( .A(n4968), .B(n4967), .Z(n4972) );
  NAND U5273 ( .A(n4970), .B(n4969), .Z(n4971) );
  NAND U5274 ( .A(n4972), .B(n4971), .Z(n5033) );
  NANDN U5275 ( .A(n4974), .B(n4973), .Z(n4978) );
  NAND U5276 ( .A(n4976), .B(n4975), .Z(n4977) );
  NAND U5277 ( .A(n4978), .B(n4977), .Z(n5031) );
  XNOR U5278 ( .A(b[7]), .B(a[112]), .Z(n5018) );
  NANDN U5279 ( .A(n5018), .B(n10545), .Z(n4981) );
  NANDN U5280 ( .A(n4979), .B(n10546), .Z(n4980) );
  NAND U5281 ( .A(n4981), .B(n4980), .Z(n5006) );
  XNOR U5282 ( .A(b[3]), .B(a[116]), .Z(n5021) );
  NANDN U5283 ( .A(n5021), .B(n10398), .Z(n4984) );
  NANDN U5284 ( .A(n4982), .B(n10399), .Z(n4983) );
  AND U5285 ( .A(n4984), .B(n4983), .Z(n5007) );
  XNOR U5286 ( .A(n5006), .B(n5007), .Z(n5008) );
  NANDN U5287 ( .A(n527), .B(a[118]), .Z(n4985) );
  XOR U5288 ( .A(n10434), .B(n4985), .Z(n4987) );
  NANDN U5289 ( .A(b[0]), .B(a[117]), .Z(n4986) );
  AND U5290 ( .A(n4987), .B(n4986), .Z(n5014) );
  XOR U5291 ( .A(b[5]), .B(a[114]), .Z(n5027) );
  NAND U5292 ( .A(n5027), .B(n10481), .Z(n4990) );
  NAND U5293 ( .A(n4988), .B(n10482), .Z(n4989) );
  NAND U5294 ( .A(n4990), .B(n4989), .Z(n5012) );
  NANDN U5295 ( .A(n529), .B(a[110]), .Z(n5013) );
  XNOR U5296 ( .A(n5012), .B(n5013), .Z(n5015) );
  XOR U5297 ( .A(n5014), .B(n5015), .Z(n5009) );
  XOR U5298 ( .A(n5008), .B(n5009), .Z(n5030) );
  XOR U5299 ( .A(n5031), .B(n5030), .Z(n5032) );
  XNOR U5300 ( .A(n5033), .B(n5032), .Z(n5002) );
  NAND U5301 ( .A(n4992), .B(n4991), .Z(n4996) );
  NAND U5302 ( .A(n4994), .B(n4993), .Z(n4995) );
  NAND U5303 ( .A(n4996), .B(n4995), .Z(n5003) );
  XNOR U5304 ( .A(n5002), .B(n5003), .Z(n5004) );
  XNOR U5305 ( .A(n5005), .B(n5004), .Z(n5036) );
  XNOR U5306 ( .A(n5036), .B(sreg[366]), .Z(n5038) );
  NAND U5307 ( .A(n4997), .B(sreg[365]), .Z(n5001) );
  OR U5308 ( .A(n4999), .B(n4998), .Z(n5000) );
  AND U5309 ( .A(n5001), .B(n5000), .Z(n5037) );
  XOR U5310 ( .A(n5038), .B(n5037), .Z(c[366]) );
  NANDN U5311 ( .A(n5007), .B(n5006), .Z(n5011) );
  NAND U5312 ( .A(n5009), .B(n5008), .Z(n5010) );
  NAND U5313 ( .A(n5011), .B(n5010), .Z(n5072) );
  NANDN U5314 ( .A(n5013), .B(n5012), .Z(n5017) );
  NAND U5315 ( .A(n5015), .B(n5014), .Z(n5016) );
  NAND U5316 ( .A(n5017), .B(n5016), .Z(n5070) );
  XNOR U5317 ( .A(b[7]), .B(a[113]), .Z(n5057) );
  NANDN U5318 ( .A(n5057), .B(n10545), .Z(n5020) );
  NANDN U5319 ( .A(n5018), .B(n10546), .Z(n5019) );
  NAND U5320 ( .A(n5020), .B(n5019), .Z(n5045) );
  XNOR U5321 ( .A(b[3]), .B(a[117]), .Z(n5060) );
  NANDN U5322 ( .A(n5060), .B(n10398), .Z(n5023) );
  NANDN U5323 ( .A(n5021), .B(n10399), .Z(n5022) );
  AND U5324 ( .A(n5023), .B(n5022), .Z(n5046) );
  XNOR U5325 ( .A(n5045), .B(n5046), .Z(n5047) );
  NANDN U5326 ( .A(n527), .B(a[119]), .Z(n5024) );
  XOR U5327 ( .A(n10434), .B(n5024), .Z(n5026) );
  NANDN U5328 ( .A(b[0]), .B(a[118]), .Z(n5025) );
  AND U5329 ( .A(n5026), .B(n5025), .Z(n5053) );
  XOR U5330 ( .A(b[5]), .B(a[115]), .Z(n5066) );
  NAND U5331 ( .A(n5066), .B(n10481), .Z(n5029) );
  NAND U5332 ( .A(n5027), .B(n10482), .Z(n5028) );
  NAND U5333 ( .A(n5029), .B(n5028), .Z(n5051) );
  NANDN U5334 ( .A(n529), .B(a[111]), .Z(n5052) );
  XNOR U5335 ( .A(n5051), .B(n5052), .Z(n5054) );
  XOR U5336 ( .A(n5053), .B(n5054), .Z(n5048) );
  XOR U5337 ( .A(n5047), .B(n5048), .Z(n5069) );
  XOR U5338 ( .A(n5070), .B(n5069), .Z(n5071) );
  XNOR U5339 ( .A(n5072), .B(n5071), .Z(n5041) );
  NAND U5340 ( .A(n5031), .B(n5030), .Z(n5035) );
  NAND U5341 ( .A(n5033), .B(n5032), .Z(n5034) );
  NAND U5342 ( .A(n5035), .B(n5034), .Z(n5042) );
  XNOR U5343 ( .A(n5041), .B(n5042), .Z(n5043) );
  XNOR U5344 ( .A(n5044), .B(n5043), .Z(n5075) );
  XNOR U5345 ( .A(n5075), .B(sreg[367]), .Z(n5077) );
  NAND U5346 ( .A(n5036), .B(sreg[366]), .Z(n5040) );
  OR U5347 ( .A(n5038), .B(n5037), .Z(n5039) );
  AND U5348 ( .A(n5040), .B(n5039), .Z(n5076) );
  XOR U5349 ( .A(n5077), .B(n5076), .Z(c[367]) );
  NANDN U5350 ( .A(n5046), .B(n5045), .Z(n5050) );
  NAND U5351 ( .A(n5048), .B(n5047), .Z(n5049) );
  NAND U5352 ( .A(n5050), .B(n5049), .Z(n5111) );
  NANDN U5353 ( .A(n5052), .B(n5051), .Z(n5056) );
  NAND U5354 ( .A(n5054), .B(n5053), .Z(n5055) );
  NAND U5355 ( .A(n5056), .B(n5055), .Z(n5109) );
  XNOR U5356 ( .A(b[7]), .B(a[114]), .Z(n5096) );
  NANDN U5357 ( .A(n5096), .B(n10545), .Z(n5059) );
  NANDN U5358 ( .A(n5057), .B(n10546), .Z(n5058) );
  NAND U5359 ( .A(n5059), .B(n5058), .Z(n5084) );
  XNOR U5360 ( .A(b[3]), .B(a[118]), .Z(n5099) );
  NANDN U5361 ( .A(n5099), .B(n10398), .Z(n5062) );
  NANDN U5362 ( .A(n5060), .B(n10399), .Z(n5061) );
  AND U5363 ( .A(n5062), .B(n5061), .Z(n5085) );
  XNOR U5364 ( .A(n5084), .B(n5085), .Z(n5086) );
  NANDN U5365 ( .A(n527), .B(a[120]), .Z(n5063) );
  XOR U5366 ( .A(n10434), .B(n5063), .Z(n5065) );
  NANDN U5367 ( .A(b[0]), .B(a[119]), .Z(n5064) );
  AND U5368 ( .A(n5065), .B(n5064), .Z(n5092) );
  XOR U5369 ( .A(b[5]), .B(a[116]), .Z(n5105) );
  NAND U5370 ( .A(n5105), .B(n10481), .Z(n5068) );
  NAND U5371 ( .A(n5066), .B(n10482), .Z(n5067) );
  NAND U5372 ( .A(n5068), .B(n5067), .Z(n5090) );
  NANDN U5373 ( .A(n529), .B(a[112]), .Z(n5091) );
  XNOR U5374 ( .A(n5090), .B(n5091), .Z(n5093) );
  XOR U5375 ( .A(n5092), .B(n5093), .Z(n5087) );
  XOR U5376 ( .A(n5086), .B(n5087), .Z(n5108) );
  XOR U5377 ( .A(n5109), .B(n5108), .Z(n5110) );
  XNOR U5378 ( .A(n5111), .B(n5110), .Z(n5080) );
  NAND U5379 ( .A(n5070), .B(n5069), .Z(n5074) );
  NAND U5380 ( .A(n5072), .B(n5071), .Z(n5073) );
  NAND U5381 ( .A(n5074), .B(n5073), .Z(n5081) );
  XNOR U5382 ( .A(n5080), .B(n5081), .Z(n5082) );
  XNOR U5383 ( .A(n5083), .B(n5082), .Z(n5114) );
  XNOR U5384 ( .A(n5114), .B(sreg[368]), .Z(n5116) );
  NAND U5385 ( .A(n5075), .B(sreg[367]), .Z(n5079) );
  OR U5386 ( .A(n5077), .B(n5076), .Z(n5078) );
  AND U5387 ( .A(n5079), .B(n5078), .Z(n5115) );
  XOR U5388 ( .A(n5116), .B(n5115), .Z(c[368]) );
  NANDN U5389 ( .A(n5085), .B(n5084), .Z(n5089) );
  NAND U5390 ( .A(n5087), .B(n5086), .Z(n5088) );
  NAND U5391 ( .A(n5089), .B(n5088), .Z(n5150) );
  NANDN U5392 ( .A(n5091), .B(n5090), .Z(n5095) );
  NAND U5393 ( .A(n5093), .B(n5092), .Z(n5094) );
  NAND U5394 ( .A(n5095), .B(n5094), .Z(n5148) );
  XNOR U5395 ( .A(b[7]), .B(a[115]), .Z(n5135) );
  NANDN U5396 ( .A(n5135), .B(n10545), .Z(n5098) );
  NANDN U5397 ( .A(n5096), .B(n10546), .Z(n5097) );
  NAND U5398 ( .A(n5098), .B(n5097), .Z(n5123) );
  XNOR U5399 ( .A(b[3]), .B(a[119]), .Z(n5138) );
  NANDN U5400 ( .A(n5138), .B(n10398), .Z(n5101) );
  NANDN U5401 ( .A(n5099), .B(n10399), .Z(n5100) );
  AND U5402 ( .A(n5101), .B(n5100), .Z(n5124) );
  XNOR U5403 ( .A(n5123), .B(n5124), .Z(n5125) );
  NANDN U5404 ( .A(n527), .B(a[121]), .Z(n5102) );
  XOR U5405 ( .A(n10434), .B(n5102), .Z(n5104) );
  NANDN U5406 ( .A(b[0]), .B(a[120]), .Z(n5103) );
  AND U5407 ( .A(n5104), .B(n5103), .Z(n5131) );
  XOR U5408 ( .A(b[5]), .B(a[117]), .Z(n5144) );
  NAND U5409 ( .A(n5144), .B(n10481), .Z(n5107) );
  NAND U5410 ( .A(n5105), .B(n10482), .Z(n5106) );
  NAND U5411 ( .A(n5107), .B(n5106), .Z(n5129) );
  NANDN U5412 ( .A(n529), .B(a[113]), .Z(n5130) );
  XNOR U5413 ( .A(n5129), .B(n5130), .Z(n5132) );
  XOR U5414 ( .A(n5131), .B(n5132), .Z(n5126) );
  XOR U5415 ( .A(n5125), .B(n5126), .Z(n5147) );
  XOR U5416 ( .A(n5148), .B(n5147), .Z(n5149) );
  XNOR U5417 ( .A(n5150), .B(n5149), .Z(n5119) );
  NAND U5418 ( .A(n5109), .B(n5108), .Z(n5113) );
  NAND U5419 ( .A(n5111), .B(n5110), .Z(n5112) );
  NAND U5420 ( .A(n5113), .B(n5112), .Z(n5120) );
  XNOR U5421 ( .A(n5119), .B(n5120), .Z(n5121) );
  XNOR U5422 ( .A(n5122), .B(n5121), .Z(n5153) );
  XNOR U5423 ( .A(n5153), .B(sreg[369]), .Z(n5155) );
  NAND U5424 ( .A(n5114), .B(sreg[368]), .Z(n5118) );
  OR U5425 ( .A(n5116), .B(n5115), .Z(n5117) );
  AND U5426 ( .A(n5118), .B(n5117), .Z(n5154) );
  XOR U5427 ( .A(n5155), .B(n5154), .Z(c[369]) );
  NANDN U5428 ( .A(n5124), .B(n5123), .Z(n5128) );
  NAND U5429 ( .A(n5126), .B(n5125), .Z(n5127) );
  NAND U5430 ( .A(n5128), .B(n5127), .Z(n5189) );
  NANDN U5431 ( .A(n5130), .B(n5129), .Z(n5134) );
  NAND U5432 ( .A(n5132), .B(n5131), .Z(n5133) );
  NAND U5433 ( .A(n5134), .B(n5133), .Z(n5187) );
  XNOR U5434 ( .A(b[7]), .B(a[116]), .Z(n5174) );
  NANDN U5435 ( .A(n5174), .B(n10545), .Z(n5137) );
  NANDN U5436 ( .A(n5135), .B(n10546), .Z(n5136) );
  NAND U5437 ( .A(n5137), .B(n5136), .Z(n5162) );
  XNOR U5438 ( .A(b[3]), .B(a[120]), .Z(n5177) );
  NANDN U5439 ( .A(n5177), .B(n10398), .Z(n5140) );
  NANDN U5440 ( .A(n5138), .B(n10399), .Z(n5139) );
  AND U5441 ( .A(n5140), .B(n5139), .Z(n5163) );
  XNOR U5442 ( .A(n5162), .B(n5163), .Z(n5164) );
  NANDN U5443 ( .A(n527), .B(a[122]), .Z(n5141) );
  XOR U5444 ( .A(n10434), .B(n5141), .Z(n5143) );
  NANDN U5445 ( .A(b[0]), .B(a[121]), .Z(n5142) );
  AND U5446 ( .A(n5143), .B(n5142), .Z(n5170) );
  XOR U5447 ( .A(b[5]), .B(a[118]), .Z(n5183) );
  NAND U5448 ( .A(n5183), .B(n10481), .Z(n5146) );
  NAND U5449 ( .A(n5144), .B(n10482), .Z(n5145) );
  NAND U5450 ( .A(n5146), .B(n5145), .Z(n5168) );
  NANDN U5451 ( .A(n529), .B(a[114]), .Z(n5169) );
  XNOR U5452 ( .A(n5168), .B(n5169), .Z(n5171) );
  XOR U5453 ( .A(n5170), .B(n5171), .Z(n5165) );
  XOR U5454 ( .A(n5164), .B(n5165), .Z(n5186) );
  XOR U5455 ( .A(n5187), .B(n5186), .Z(n5188) );
  XNOR U5456 ( .A(n5189), .B(n5188), .Z(n5158) );
  NAND U5457 ( .A(n5148), .B(n5147), .Z(n5152) );
  NAND U5458 ( .A(n5150), .B(n5149), .Z(n5151) );
  NAND U5459 ( .A(n5152), .B(n5151), .Z(n5159) );
  XNOR U5460 ( .A(n5158), .B(n5159), .Z(n5160) );
  XNOR U5461 ( .A(n5161), .B(n5160), .Z(n5192) );
  XNOR U5462 ( .A(n5192), .B(sreg[370]), .Z(n5194) );
  NAND U5463 ( .A(n5153), .B(sreg[369]), .Z(n5157) );
  OR U5464 ( .A(n5155), .B(n5154), .Z(n5156) );
  AND U5465 ( .A(n5157), .B(n5156), .Z(n5193) );
  XOR U5466 ( .A(n5194), .B(n5193), .Z(c[370]) );
  NANDN U5467 ( .A(n5163), .B(n5162), .Z(n5167) );
  NAND U5468 ( .A(n5165), .B(n5164), .Z(n5166) );
  NAND U5469 ( .A(n5167), .B(n5166), .Z(n5228) );
  NANDN U5470 ( .A(n5169), .B(n5168), .Z(n5173) );
  NAND U5471 ( .A(n5171), .B(n5170), .Z(n5172) );
  NAND U5472 ( .A(n5173), .B(n5172), .Z(n5226) );
  XNOR U5473 ( .A(b[7]), .B(a[117]), .Z(n5213) );
  NANDN U5474 ( .A(n5213), .B(n10545), .Z(n5176) );
  NANDN U5475 ( .A(n5174), .B(n10546), .Z(n5175) );
  NAND U5476 ( .A(n5176), .B(n5175), .Z(n5201) );
  XNOR U5477 ( .A(b[3]), .B(a[121]), .Z(n5216) );
  NANDN U5478 ( .A(n5216), .B(n10398), .Z(n5179) );
  NANDN U5479 ( .A(n5177), .B(n10399), .Z(n5178) );
  AND U5480 ( .A(n5179), .B(n5178), .Z(n5202) );
  XNOR U5481 ( .A(n5201), .B(n5202), .Z(n5203) );
  NANDN U5482 ( .A(n527), .B(a[123]), .Z(n5180) );
  XOR U5483 ( .A(n10434), .B(n5180), .Z(n5182) );
  NANDN U5484 ( .A(b[0]), .B(a[122]), .Z(n5181) );
  AND U5485 ( .A(n5182), .B(n5181), .Z(n5209) );
  XOR U5486 ( .A(b[5]), .B(a[119]), .Z(n5222) );
  NAND U5487 ( .A(n5222), .B(n10481), .Z(n5185) );
  NAND U5488 ( .A(n5183), .B(n10482), .Z(n5184) );
  NAND U5489 ( .A(n5185), .B(n5184), .Z(n5207) );
  NANDN U5490 ( .A(n529), .B(a[115]), .Z(n5208) );
  XNOR U5491 ( .A(n5207), .B(n5208), .Z(n5210) );
  XOR U5492 ( .A(n5209), .B(n5210), .Z(n5204) );
  XOR U5493 ( .A(n5203), .B(n5204), .Z(n5225) );
  XOR U5494 ( .A(n5226), .B(n5225), .Z(n5227) );
  XNOR U5495 ( .A(n5228), .B(n5227), .Z(n5197) );
  NAND U5496 ( .A(n5187), .B(n5186), .Z(n5191) );
  NAND U5497 ( .A(n5189), .B(n5188), .Z(n5190) );
  NAND U5498 ( .A(n5191), .B(n5190), .Z(n5198) );
  XNOR U5499 ( .A(n5197), .B(n5198), .Z(n5199) );
  XNOR U5500 ( .A(n5200), .B(n5199), .Z(n5231) );
  XNOR U5501 ( .A(n5231), .B(sreg[371]), .Z(n5233) );
  NAND U5502 ( .A(n5192), .B(sreg[370]), .Z(n5196) );
  OR U5503 ( .A(n5194), .B(n5193), .Z(n5195) );
  AND U5504 ( .A(n5196), .B(n5195), .Z(n5232) );
  XOR U5505 ( .A(n5233), .B(n5232), .Z(c[371]) );
  NANDN U5506 ( .A(n5202), .B(n5201), .Z(n5206) );
  NAND U5507 ( .A(n5204), .B(n5203), .Z(n5205) );
  NAND U5508 ( .A(n5206), .B(n5205), .Z(n5267) );
  NANDN U5509 ( .A(n5208), .B(n5207), .Z(n5212) );
  NAND U5510 ( .A(n5210), .B(n5209), .Z(n5211) );
  NAND U5511 ( .A(n5212), .B(n5211), .Z(n5265) );
  XNOR U5512 ( .A(b[7]), .B(a[118]), .Z(n5252) );
  NANDN U5513 ( .A(n5252), .B(n10545), .Z(n5215) );
  NANDN U5514 ( .A(n5213), .B(n10546), .Z(n5214) );
  NAND U5515 ( .A(n5215), .B(n5214), .Z(n5240) );
  XNOR U5516 ( .A(b[3]), .B(a[122]), .Z(n5255) );
  NANDN U5517 ( .A(n5255), .B(n10398), .Z(n5218) );
  NANDN U5518 ( .A(n5216), .B(n10399), .Z(n5217) );
  AND U5519 ( .A(n5218), .B(n5217), .Z(n5241) );
  XNOR U5520 ( .A(n5240), .B(n5241), .Z(n5242) );
  NANDN U5521 ( .A(n527), .B(a[124]), .Z(n5219) );
  XOR U5522 ( .A(n10434), .B(n5219), .Z(n5221) );
  NANDN U5523 ( .A(b[0]), .B(a[123]), .Z(n5220) );
  AND U5524 ( .A(n5221), .B(n5220), .Z(n5248) );
  XOR U5525 ( .A(b[5]), .B(a[120]), .Z(n5261) );
  NAND U5526 ( .A(n5261), .B(n10481), .Z(n5224) );
  NAND U5527 ( .A(n5222), .B(n10482), .Z(n5223) );
  NAND U5528 ( .A(n5224), .B(n5223), .Z(n5246) );
  NANDN U5529 ( .A(n529), .B(a[116]), .Z(n5247) );
  XNOR U5530 ( .A(n5246), .B(n5247), .Z(n5249) );
  XOR U5531 ( .A(n5248), .B(n5249), .Z(n5243) );
  XOR U5532 ( .A(n5242), .B(n5243), .Z(n5264) );
  XOR U5533 ( .A(n5265), .B(n5264), .Z(n5266) );
  XNOR U5534 ( .A(n5267), .B(n5266), .Z(n5236) );
  NAND U5535 ( .A(n5226), .B(n5225), .Z(n5230) );
  NAND U5536 ( .A(n5228), .B(n5227), .Z(n5229) );
  NAND U5537 ( .A(n5230), .B(n5229), .Z(n5237) );
  XNOR U5538 ( .A(n5236), .B(n5237), .Z(n5238) );
  XNOR U5539 ( .A(n5239), .B(n5238), .Z(n5270) );
  XNOR U5540 ( .A(n5270), .B(sreg[372]), .Z(n5272) );
  NAND U5541 ( .A(n5231), .B(sreg[371]), .Z(n5235) );
  OR U5542 ( .A(n5233), .B(n5232), .Z(n5234) );
  AND U5543 ( .A(n5235), .B(n5234), .Z(n5271) );
  XOR U5544 ( .A(n5272), .B(n5271), .Z(c[372]) );
  NANDN U5545 ( .A(n5241), .B(n5240), .Z(n5245) );
  NAND U5546 ( .A(n5243), .B(n5242), .Z(n5244) );
  NAND U5547 ( .A(n5245), .B(n5244), .Z(n5306) );
  NANDN U5548 ( .A(n5247), .B(n5246), .Z(n5251) );
  NAND U5549 ( .A(n5249), .B(n5248), .Z(n5250) );
  NAND U5550 ( .A(n5251), .B(n5250), .Z(n5304) );
  XNOR U5551 ( .A(b[7]), .B(a[119]), .Z(n5291) );
  NANDN U5552 ( .A(n5291), .B(n10545), .Z(n5254) );
  NANDN U5553 ( .A(n5252), .B(n10546), .Z(n5253) );
  NAND U5554 ( .A(n5254), .B(n5253), .Z(n5279) );
  XNOR U5555 ( .A(b[3]), .B(a[123]), .Z(n5294) );
  NANDN U5556 ( .A(n5294), .B(n10398), .Z(n5257) );
  NANDN U5557 ( .A(n5255), .B(n10399), .Z(n5256) );
  AND U5558 ( .A(n5257), .B(n5256), .Z(n5280) );
  XNOR U5559 ( .A(n5279), .B(n5280), .Z(n5281) );
  NANDN U5560 ( .A(n527), .B(a[125]), .Z(n5258) );
  XOR U5561 ( .A(n10434), .B(n5258), .Z(n5260) );
  NANDN U5562 ( .A(b[0]), .B(a[124]), .Z(n5259) );
  AND U5563 ( .A(n5260), .B(n5259), .Z(n5287) );
  XOR U5564 ( .A(b[5]), .B(a[121]), .Z(n5300) );
  NAND U5565 ( .A(n5300), .B(n10481), .Z(n5263) );
  NAND U5566 ( .A(n5261), .B(n10482), .Z(n5262) );
  NAND U5567 ( .A(n5263), .B(n5262), .Z(n5285) );
  NANDN U5568 ( .A(n529), .B(a[117]), .Z(n5286) );
  XNOR U5569 ( .A(n5285), .B(n5286), .Z(n5288) );
  XOR U5570 ( .A(n5287), .B(n5288), .Z(n5282) );
  XOR U5571 ( .A(n5281), .B(n5282), .Z(n5303) );
  XOR U5572 ( .A(n5304), .B(n5303), .Z(n5305) );
  XNOR U5573 ( .A(n5306), .B(n5305), .Z(n5275) );
  NAND U5574 ( .A(n5265), .B(n5264), .Z(n5269) );
  NAND U5575 ( .A(n5267), .B(n5266), .Z(n5268) );
  NAND U5576 ( .A(n5269), .B(n5268), .Z(n5276) );
  XNOR U5577 ( .A(n5275), .B(n5276), .Z(n5277) );
  XNOR U5578 ( .A(n5278), .B(n5277), .Z(n5309) );
  XNOR U5579 ( .A(n5309), .B(sreg[373]), .Z(n5311) );
  NAND U5580 ( .A(n5270), .B(sreg[372]), .Z(n5274) );
  OR U5581 ( .A(n5272), .B(n5271), .Z(n5273) );
  AND U5582 ( .A(n5274), .B(n5273), .Z(n5310) );
  XOR U5583 ( .A(n5311), .B(n5310), .Z(c[373]) );
  NANDN U5584 ( .A(n5280), .B(n5279), .Z(n5284) );
  NAND U5585 ( .A(n5282), .B(n5281), .Z(n5283) );
  NAND U5586 ( .A(n5284), .B(n5283), .Z(n5345) );
  NANDN U5587 ( .A(n5286), .B(n5285), .Z(n5290) );
  NAND U5588 ( .A(n5288), .B(n5287), .Z(n5289) );
  NAND U5589 ( .A(n5290), .B(n5289), .Z(n5343) );
  XNOR U5590 ( .A(b[7]), .B(a[120]), .Z(n5330) );
  NANDN U5591 ( .A(n5330), .B(n10545), .Z(n5293) );
  NANDN U5592 ( .A(n5291), .B(n10546), .Z(n5292) );
  NAND U5593 ( .A(n5293), .B(n5292), .Z(n5318) );
  XNOR U5594 ( .A(b[3]), .B(a[124]), .Z(n5333) );
  NANDN U5595 ( .A(n5333), .B(n10398), .Z(n5296) );
  NANDN U5596 ( .A(n5294), .B(n10399), .Z(n5295) );
  AND U5597 ( .A(n5296), .B(n5295), .Z(n5319) );
  XNOR U5598 ( .A(n5318), .B(n5319), .Z(n5320) );
  NANDN U5599 ( .A(n527), .B(a[126]), .Z(n5297) );
  XOR U5600 ( .A(n10434), .B(n5297), .Z(n5299) );
  NANDN U5601 ( .A(b[0]), .B(a[125]), .Z(n5298) );
  AND U5602 ( .A(n5299), .B(n5298), .Z(n5326) );
  XOR U5603 ( .A(b[5]), .B(a[122]), .Z(n5339) );
  NAND U5604 ( .A(n5339), .B(n10481), .Z(n5302) );
  NAND U5605 ( .A(n5300), .B(n10482), .Z(n5301) );
  NAND U5606 ( .A(n5302), .B(n5301), .Z(n5324) );
  NANDN U5607 ( .A(n529), .B(a[118]), .Z(n5325) );
  XNOR U5608 ( .A(n5324), .B(n5325), .Z(n5327) );
  XOR U5609 ( .A(n5326), .B(n5327), .Z(n5321) );
  XOR U5610 ( .A(n5320), .B(n5321), .Z(n5342) );
  XOR U5611 ( .A(n5343), .B(n5342), .Z(n5344) );
  XNOR U5612 ( .A(n5345), .B(n5344), .Z(n5314) );
  NAND U5613 ( .A(n5304), .B(n5303), .Z(n5308) );
  NAND U5614 ( .A(n5306), .B(n5305), .Z(n5307) );
  NAND U5615 ( .A(n5308), .B(n5307), .Z(n5315) );
  XNOR U5616 ( .A(n5314), .B(n5315), .Z(n5316) );
  XNOR U5617 ( .A(n5317), .B(n5316), .Z(n5348) );
  XNOR U5618 ( .A(n5348), .B(sreg[374]), .Z(n5350) );
  NAND U5619 ( .A(n5309), .B(sreg[373]), .Z(n5313) );
  OR U5620 ( .A(n5311), .B(n5310), .Z(n5312) );
  AND U5621 ( .A(n5313), .B(n5312), .Z(n5349) );
  XOR U5622 ( .A(n5350), .B(n5349), .Z(c[374]) );
  NANDN U5623 ( .A(n5319), .B(n5318), .Z(n5323) );
  NAND U5624 ( .A(n5321), .B(n5320), .Z(n5322) );
  NAND U5625 ( .A(n5323), .B(n5322), .Z(n5384) );
  NANDN U5626 ( .A(n5325), .B(n5324), .Z(n5329) );
  NAND U5627 ( .A(n5327), .B(n5326), .Z(n5328) );
  NAND U5628 ( .A(n5329), .B(n5328), .Z(n5382) );
  XNOR U5629 ( .A(b[7]), .B(a[121]), .Z(n5369) );
  NANDN U5630 ( .A(n5369), .B(n10545), .Z(n5332) );
  NANDN U5631 ( .A(n5330), .B(n10546), .Z(n5331) );
  NAND U5632 ( .A(n5332), .B(n5331), .Z(n5357) );
  XNOR U5633 ( .A(b[3]), .B(a[125]), .Z(n5372) );
  NANDN U5634 ( .A(n5372), .B(n10398), .Z(n5335) );
  NANDN U5635 ( .A(n5333), .B(n10399), .Z(n5334) );
  AND U5636 ( .A(n5335), .B(n5334), .Z(n5358) );
  XNOR U5637 ( .A(n5357), .B(n5358), .Z(n5359) );
  NANDN U5638 ( .A(n527), .B(a[127]), .Z(n5336) );
  XOR U5639 ( .A(n10434), .B(n5336), .Z(n5338) );
  NANDN U5640 ( .A(b[0]), .B(a[126]), .Z(n5337) );
  AND U5641 ( .A(n5338), .B(n5337), .Z(n5365) );
  XOR U5642 ( .A(b[5]), .B(a[123]), .Z(n5378) );
  NAND U5643 ( .A(n5378), .B(n10481), .Z(n5341) );
  NAND U5644 ( .A(n5339), .B(n10482), .Z(n5340) );
  NAND U5645 ( .A(n5341), .B(n5340), .Z(n5363) );
  NANDN U5646 ( .A(n529), .B(a[119]), .Z(n5364) );
  XNOR U5647 ( .A(n5363), .B(n5364), .Z(n5366) );
  XOR U5648 ( .A(n5365), .B(n5366), .Z(n5360) );
  XOR U5649 ( .A(n5359), .B(n5360), .Z(n5381) );
  XOR U5650 ( .A(n5382), .B(n5381), .Z(n5383) );
  XNOR U5651 ( .A(n5384), .B(n5383), .Z(n5353) );
  NAND U5652 ( .A(n5343), .B(n5342), .Z(n5347) );
  NAND U5653 ( .A(n5345), .B(n5344), .Z(n5346) );
  NAND U5654 ( .A(n5347), .B(n5346), .Z(n5354) );
  XNOR U5655 ( .A(n5353), .B(n5354), .Z(n5355) );
  XNOR U5656 ( .A(n5356), .B(n5355), .Z(n5387) );
  XNOR U5657 ( .A(n5387), .B(sreg[375]), .Z(n5389) );
  NAND U5658 ( .A(n5348), .B(sreg[374]), .Z(n5352) );
  OR U5659 ( .A(n5350), .B(n5349), .Z(n5351) );
  AND U5660 ( .A(n5352), .B(n5351), .Z(n5388) );
  XOR U5661 ( .A(n5389), .B(n5388), .Z(c[375]) );
  NANDN U5662 ( .A(n5358), .B(n5357), .Z(n5362) );
  NAND U5663 ( .A(n5360), .B(n5359), .Z(n5361) );
  NAND U5664 ( .A(n5362), .B(n5361), .Z(n5423) );
  NANDN U5665 ( .A(n5364), .B(n5363), .Z(n5368) );
  NAND U5666 ( .A(n5366), .B(n5365), .Z(n5367) );
  NAND U5667 ( .A(n5368), .B(n5367), .Z(n5421) );
  XNOR U5668 ( .A(b[7]), .B(a[122]), .Z(n5408) );
  NANDN U5669 ( .A(n5408), .B(n10545), .Z(n5371) );
  NANDN U5670 ( .A(n5369), .B(n10546), .Z(n5370) );
  NAND U5671 ( .A(n5371), .B(n5370), .Z(n5396) );
  XNOR U5672 ( .A(b[3]), .B(a[126]), .Z(n5411) );
  NANDN U5673 ( .A(n5411), .B(n10398), .Z(n5374) );
  NANDN U5674 ( .A(n5372), .B(n10399), .Z(n5373) );
  AND U5675 ( .A(n5374), .B(n5373), .Z(n5397) );
  XNOR U5676 ( .A(n5396), .B(n5397), .Z(n5398) );
  NANDN U5677 ( .A(n527), .B(a[128]), .Z(n5375) );
  XOR U5678 ( .A(n10434), .B(n5375), .Z(n5377) );
  NANDN U5679 ( .A(b[0]), .B(a[127]), .Z(n5376) );
  AND U5680 ( .A(n5377), .B(n5376), .Z(n5404) );
  XOR U5681 ( .A(b[5]), .B(a[124]), .Z(n5417) );
  NAND U5682 ( .A(n5417), .B(n10481), .Z(n5380) );
  NAND U5683 ( .A(n5378), .B(n10482), .Z(n5379) );
  NAND U5684 ( .A(n5380), .B(n5379), .Z(n5402) );
  NANDN U5685 ( .A(n529), .B(a[120]), .Z(n5403) );
  XNOR U5686 ( .A(n5402), .B(n5403), .Z(n5405) );
  XOR U5687 ( .A(n5404), .B(n5405), .Z(n5399) );
  XOR U5688 ( .A(n5398), .B(n5399), .Z(n5420) );
  XOR U5689 ( .A(n5421), .B(n5420), .Z(n5422) );
  XNOR U5690 ( .A(n5423), .B(n5422), .Z(n5392) );
  NAND U5691 ( .A(n5382), .B(n5381), .Z(n5386) );
  NAND U5692 ( .A(n5384), .B(n5383), .Z(n5385) );
  NAND U5693 ( .A(n5386), .B(n5385), .Z(n5393) );
  XNOR U5694 ( .A(n5392), .B(n5393), .Z(n5394) );
  XNOR U5695 ( .A(n5395), .B(n5394), .Z(n5426) );
  XNOR U5696 ( .A(n5426), .B(sreg[376]), .Z(n5428) );
  NAND U5697 ( .A(n5387), .B(sreg[375]), .Z(n5391) );
  OR U5698 ( .A(n5389), .B(n5388), .Z(n5390) );
  AND U5699 ( .A(n5391), .B(n5390), .Z(n5427) );
  XOR U5700 ( .A(n5428), .B(n5427), .Z(c[376]) );
  NANDN U5701 ( .A(n5397), .B(n5396), .Z(n5401) );
  NAND U5702 ( .A(n5399), .B(n5398), .Z(n5400) );
  NAND U5703 ( .A(n5401), .B(n5400), .Z(n5462) );
  NANDN U5704 ( .A(n5403), .B(n5402), .Z(n5407) );
  NAND U5705 ( .A(n5405), .B(n5404), .Z(n5406) );
  NAND U5706 ( .A(n5407), .B(n5406), .Z(n5460) );
  XNOR U5707 ( .A(b[7]), .B(a[123]), .Z(n5447) );
  NANDN U5708 ( .A(n5447), .B(n10545), .Z(n5410) );
  NANDN U5709 ( .A(n5408), .B(n10546), .Z(n5409) );
  NAND U5710 ( .A(n5410), .B(n5409), .Z(n5435) );
  XNOR U5711 ( .A(b[3]), .B(a[127]), .Z(n5450) );
  NANDN U5712 ( .A(n5450), .B(n10398), .Z(n5413) );
  NANDN U5713 ( .A(n5411), .B(n10399), .Z(n5412) );
  AND U5714 ( .A(n5413), .B(n5412), .Z(n5436) );
  XNOR U5715 ( .A(n5435), .B(n5436), .Z(n5437) );
  NANDN U5716 ( .A(n527), .B(a[129]), .Z(n5414) );
  XOR U5717 ( .A(n10434), .B(n5414), .Z(n5416) );
  NANDN U5718 ( .A(b[0]), .B(a[128]), .Z(n5415) );
  AND U5719 ( .A(n5416), .B(n5415), .Z(n5443) );
  XOR U5720 ( .A(b[5]), .B(a[125]), .Z(n5456) );
  NAND U5721 ( .A(n5456), .B(n10481), .Z(n5419) );
  NAND U5722 ( .A(n5417), .B(n10482), .Z(n5418) );
  NAND U5723 ( .A(n5419), .B(n5418), .Z(n5441) );
  NANDN U5724 ( .A(n529), .B(a[121]), .Z(n5442) );
  XNOR U5725 ( .A(n5441), .B(n5442), .Z(n5444) );
  XOR U5726 ( .A(n5443), .B(n5444), .Z(n5438) );
  XOR U5727 ( .A(n5437), .B(n5438), .Z(n5459) );
  XOR U5728 ( .A(n5460), .B(n5459), .Z(n5461) );
  XNOR U5729 ( .A(n5462), .B(n5461), .Z(n5431) );
  NAND U5730 ( .A(n5421), .B(n5420), .Z(n5425) );
  NAND U5731 ( .A(n5423), .B(n5422), .Z(n5424) );
  NAND U5732 ( .A(n5425), .B(n5424), .Z(n5432) );
  XNOR U5733 ( .A(n5431), .B(n5432), .Z(n5433) );
  XNOR U5734 ( .A(n5434), .B(n5433), .Z(n5465) );
  XNOR U5735 ( .A(n5465), .B(sreg[377]), .Z(n5467) );
  NAND U5736 ( .A(n5426), .B(sreg[376]), .Z(n5430) );
  OR U5737 ( .A(n5428), .B(n5427), .Z(n5429) );
  AND U5738 ( .A(n5430), .B(n5429), .Z(n5466) );
  XOR U5739 ( .A(n5467), .B(n5466), .Z(c[377]) );
  NANDN U5740 ( .A(n5436), .B(n5435), .Z(n5440) );
  NAND U5741 ( .A(n5438), .B(n5437), .Z(n5439) );
  NAND U5742 ( .A(n5440), .B(n5439), .Z(n5501) );
  NANDN U5743 ( .A(n5442), .B(n5441), .Z(n5446) );
  NAND U5744 ( .A(n5444), .B(n5443), .Z(n5445) );
  NAND U5745 ( .A(n5446), .B(n5445), .Z(n5499) );
  XNOR U5746 ( .A(b[7]), .B(a[124]), .Z(n5486) );
  NANDN U5747 ( .A(n5486), .B(n10545), .Z(n5449) );
  NANDN U5748 ( .A(n5447), .B(n10546), .Z(n5448) );
  NAND U5749 ( .A(n5449), .B(n5448), .Z(n5474) );
  XNOR U5750 ( .A(b[3]), .B(a[128]), .Z(n5489) );
  NANDN U5751 ( .A(n5489), .B(n10398), .Z(n5452) );
  NANDN U5752 ( .A(n5450), .B(n10399), .Z(n5451) );
  AND U5753 ( .A(n5452), .B(n5451), .Z(n5475) );
  XNOR U5754 ( .A(n5474), .B(n5475), .Z(n5476) );
  NANDN U5755 ( .A(n527), .B(a[130]), .Z(n5453) );
  XOR U5756 ( .A(n10434), .B(n5453), .Z(n5455) );
  NANDN U5757 ( .A(b[0]), .B(a[129]), .Z(n5454) );
  AND U5758 ( .A(n5455), .B(n5454), .Z(n5482) );
  XOR U5759 ( .A(b[5]), .B(a[126]), .Z(n5495) );
  NAND U5760 ( .A(n5495), .B(n10481), .Z(n5458) );
  NAND U5761 ( .A(n5456), .B(n10482), .Z(n5457) );
  NAND U5762 ( .A(n5458), .B(n5457), .Z(n5480) );
  NANDN U5763 ( .A(n529), .B(a[122]), .Z(n5481) );
  XNOR U5764 ( .A(n5480), .B(n5481), .Z(n5483) );
  XOR U5765 ( .A(n5482), .B(n5483), .Z(n5477) );
  XOR U5766 ( .A(n5476), .B(n5477), .Z(n5498) );
  XOR U5767 ( .A(n5499), .B(n5498), .Z(n5500) );
  XNOR U5768 ( .A(n5501), .B(n5500), .Z(n5470) );
  NAND U5769 ( .A(n5460), .B(n5459), .Z(n5464) );
  NAND U5770 ( .A(n5462), .B(n5461), .Z(n5463) );
  NAND U5771 ( .A(n5464), .B(n5463), .Z(n5471) );
  XNOR U5772 ( .A(n5470), .B(n5471), .Z(n5472) );
  XNOR U5773 ( .A(n5473), .B(n5472), .Z(n5504) );
  XNOR U5774 ( .A(n5504), .B(sreg[378]), .Z(n5506) );
  NAND U5775 ( .A(n5465), .B(sreg[377]), .Z(n5469) );
  OR U5776 ( .A(n5467), .B(n5466), .Z(n5468) );
  AND U5777 ( .A(n5469), .B(n5468), .Z(n5505) );
  XOR U5778 ( .A(n5506), .B(n5505), .Z(c[378]) );
  NANDN U5779 ( .A(n5475), .B(n5474), .Z(n5479) );
  NAND U5780 ( .A(n5477), .B(n5476), .Z(n5478) );
  NAND U5781 ( .A(n5479), .B(n5478), .Z(n5540) );
  NANDN U5782 ( .A(n5481), .B(n5480), .Z(n5485) );
  NAND U5783 ( .A(n5483), .B(n5482), .Z(n5484) );
  NAND U5784 ( .A(n5485), .B(n5484), .Z(n5538) );
  XNOR U5785 ( .A(b[7]), .B(a[125]), .Z(n5531) );
  NANDN U5786 ( .A(n5531), .B(n10545), .Z(n5488) );
  NANDN U5787 ( .A(n5486), .B(n10546), .Z(n5487) );
  NAND U5788 ( .A(n5488), .B(n5487), .Z(n5513) );
  XNOR U5789 ( .A(b[3]), .B(a[129]), .Z(n5534) );
  NANDN U5790 ( .A(n5534), .B(n10398), .Z(n5491) );
  NANDN U5791 ( .A(n5489), .B(n10399), .Z(n5490) );
  AND U5792 ( .A(n5491), .B(n5490), .Z(n5514) );
  XNOR U5793 ( .A(n5513), .B(n5514), .Z(n5515) );
  NANDN U5794 ( .A(n527), .B(a[131]), .Z(n5492) );
  XOR U5795 ( .A(n10434), .B(n5492), .Z(n5494) );
  NANDN U5796 ( .A(b[0]), .B(a[130]), .Z(n5493) );
  AND U5797 ( .A(n5494), .B(n5493), .Z(n5521) );
  XOR U5798 ( .A(b[5]), .B(a[127]), .Z(n5528) );
  NAND U5799 ( .A(n5528), .B(n10481), .Z(n5497) );
  NAND U5800 ( .A(n5495), .B(n10482), .Z(n5496) );
  NAND U5801 ( .A(n5497), .B(n5496), .Z(n5519) );
  NANDN U5802 ( .A(n529), .B(a[123]), .Z(n5520) );
  XNOR U5803 ( .A(n5519), .B(n5520), .Z(n5522) );
  XOR U5804 ( .A(n5521), .B(n5522), .Z(n5516) );
  XOR U5805 ( .A(n5515), .B(n5516), .Z(n5537) );
  XOR U5806 ( .A(n5538), .B(n5537), .Z(n5539) );
  XNOR U5807 ( .A(n5540), .B(n5539), .Z(n5509) );
  NAND U5808 ( .A(n5499), .B(n5498), .Z(n5503) );
  NAND U5809 ( .A(n5501), .B(n5500), .Z(n5502) );
  NAND U5810 ( .A(n5503), .B(n5502), .Z(n5510) );
  XNOR U5811 ( .A(n5509), .B(n5510), .Z(n5511) );
  XNOR U5812 ( .A(n5512), .B(n5511), .Z(n5543) );
  XNOR U5813 ( .A(n5543), .B(sreg[379]), .Z(n5545) );
  NAND U5814 ( .A(n5504), .B(sreg[378]), .Z(n5508) );
  OR U5815 ( .A(n5506), .B(n5505), .Z(n5507) );
  AND U5816 ( .A(n5508), .B(n5507), .Z(n5544) );
  XOR U5817 ( .A(n5545), .B(n5544), .Z(c[379]) );
  NANDN U5818 ( .A(n5514), .B(n5513), .Z(n5518) );
  NAND U5819 ( .A(n5516), .B(n5515), .Z(n5517) );
  NAND U5820 ( .A(n5518), .B(n5517), .Z(n5579) );
  NANDN U5821 ( .A(n5520), .B(n5519), .Z(n5524) );
  NAND U5822 ( .A(n5522), .B(n5521), .Z(n5523) );
  NAND U5823 ( .A(n5524), .B(n5523), .Z(n5577) );
  NANDN U5824 ( .A(n527), .B(a[132]), .Z(n5525) );
  XOR U5825 ( .A(n10434), .B(n5525), .Z(n5527) );
  NANDN U5826 ( .A(b[0]), .B(a[131]), .Z(n5526) );
  AND U5827 ( .A(n5527), .B(n5526), .Z(n5560) );
  XOR U5828 ( .A(b[5]), .B(a[128]), .Z(n5573) );
  NAND U5829 ( .A(n5573), .B(n10481), .Z(n5530) );
  NAND U5830 ( .A(n5528), .B(n10482), .Z(n5529) );
  NAND U5831 ( .A(n5530), .B(n5529), .Z(n5558) );
  NANDN U5832 ( .A(n529), .B(a[124]), .Z(n5559) );
  XNOR U5833 ( .A(n5558), .B(n5559), .Z(n5561) );
  XOR U5834 ( .A(n5560), .B(n5561), .Z(n5554) );
  XNOR U5835 ( .A(b[7]), .B(a[126]), .Z(n5564) );
  NANDN U5836 ( .A(n5564), .B(n10545), .Z(n5533) );
  NANDN U5837 ( .A(n5531), .B(n10546), .Z(n5532) );
  NAND U5838 ( .A(n5533), .B(n5532), .Z(n5552) );
  XNOR U5839 ( .A(b[3]), .B(a[130]), .Z(n5567) );
  NANDN U5840 ( .A(n5567), .B(n10398), .Z(n5536) );
  NANDN U5841 ( .A(n5534), .B(n10399), .Z(n5535) );
  AND U5842 ( .A(n5536), .B(n5535), .Z(n5553) );
  XNOR U5843 ( .A(n5552), .B(n5553), .Z(n5555) );
  XOR U5844 ( .A(n5554), .B(n5555), .Z(n5576) );
  XOR U5845 ( .A(n5577), .B(n5576), .Z(n5578) );
  XNOR U5846 ( .A(n5579), .B(n5578), .Z(n5548) );
  NAND U5847 ( .A(n5538), .B(n5537), .Z(n5542) );
  NAND U5848 ( .A(n5540), .B(n5539), .Z(n5541) );
  NAND U5849 ( .A(n5542), .B(n5541), .Z(n5549) );
  XNOR U5850 ( .A(n5548), .B(n5549), .Z(n5550) );
  XNOR U5851 ( .A(n5551), .B(n5550), .Z(n5582) );
  XNOR U5852 ( .A(n5582), .B(sreg[380]), .Z(n5584) );
  NAND U5853 ( .A(n5543), .B(sreg[379]), .Z(n5547) );
  OR U5854 ( .A(n5545), .B(n5544), .Z(n5546) );
  AND U5855 ( .A(n5547), .B(n5546), .Z(n5583) );
  XOR U5856 ( .A(n5584), .B(n5583), .Z(c[380]) );
  NANDN U5857 ( .A(n5553), .B(n5552), .Z(n5557) );
  NAND U5858 ( .A(n5555), .B(n5554), .Z(n5556) );
  NAND U5859 ( .A(n5557), .B(n5556), .Z(n5618) );
  NANDN U5860 ( .A(n5559), .B(n5558), .Z(n5563) );
  NAND U5861 ( .A(n5561), .B(n5560), .Z(n5562) );
  NAND U5862 ( .A(n5563), .B(n5562), .Z(n5616) );
  XNOR U5863 ( .A(b[7]), .B(a[127]), .Z(n5603) );
  NANDN U5864 ( .A(n5603), .B(n10545), .Z(n5566) );
  NANDN U5865 ( .A(n5564), .B(n10546), .Z(n5565) );
  NAND U5866 ( .A(n5566), .B(n5565), .Z(n5591) );
  XNOR U5867 ( .A(b[3]), .B(a[131]), .Z(n5606) );
  NANDN U5868 ( .A(n5606), .B(n10398), .Z(n5569) );
  NANDN U5869 ( .A(n5567), .B(n10399), .Z(n5568) );
  AND U5870 ( .A(n5569), .B(n5568), .Z(n5592) );
  XNOR U5871 ( .A(n5591), .B(n5592), .Z(n5593) );
  NANDN U5872 ( .A(n527), .B(a[133]), .Z(n5570) );
  XOR U5873 ( .A(n10434), .B(n5570), .Z(n5572) );
  NANDN U5874 ( .A(b[0]), .B(a[132]), .Z(n5571) );
  AND U5875 ( .A(n5572), .B(n5571), .Z(n5599) );
  XOR U5876 ( .A(b[5]), .B(a[129]), .Z(n5612) );
  NAND U5877 ( .A(n5612), .B(n10481), .Z(n5575) );
  NAND U5878 ( .A(n5573), .B(n10482), .Z(n5574) );
  NAND U5879 ( .A(n5575), .B(n5574), .Z(n5597) );
  NANDN U5880 ( .A(n529), .B(a[125]), .Z(n5598) );
  XNOR U5881 ( .A(n5597), .B(n5598), .Z(n5600) );
  XOR U5882 ( .A(n5599), .B(n5600), .Z(n5594) );
  XOR U5883 ( .A(n5593), .B(n5594), .Z(n5615) );
  XOR U5884 ( .A(n5616), .B(n5615), .Z(n5617) );
  XNOR U5885 ( .A(n5618), .B(n5617), .Z(n5587) );
  NAND U5886 ( .A(n5577), .B(n5576), .Z(n5581) );
  NAND U5887 ( .A(n5579), .B(n5578), .Z(n5580) );
  NAND U5888 ( .A(n5581), .B(n5580), .Z(n5588) );
  XNOR U5889 ( .A(n5587), .B(n5588), .Z(n5589) );
  XNOR U5890 ( .A(n5590), .B(n5589), .Z(n5621) );
  XNOR U5891 ( .A(n5621), .B(sreg[381]), .Z(n5623) );
  NAND U5892 ( .A(n5582), .B(sreg[380]), .Z(n5586) );
  OR U5893 ( .A(n5584), .B(n5583), .Z(n5585) );
  AND U5894 ( .A(n5586), .B(n5585), .Z(n5622) );
  XOR U5895 ( .A(n5623), .B(n5622), .Z(c[381]) );
  NANDN U5896 ( .A(n5592), .B(n5591), .Z(n5596) );
  NAND U5897 ( .A(n5594), .B(n5593), .Z(n5595) );
  NAND U5898 ( .A(n5596), .B(n5595), .Z(n5657) );
  NANDN U5899 ( .A(n5598), .B(n5597), .Z(n5602) );
  NAND U5900 ( .A(n5600), .B(n5599), .Z(n5601) );
  NAND U5901 ( .A(n5602), .B(n5601), .Z(n5655) );
  XNOR U5902 ( .A(b[7]), .B(a[128]), .Z(n5642) );
  NANDN U5903 ( .A(n5642), .B(n10545), .Z(n5605) );
  NANDN U5904 ( .A(n5603), .B(n10546), .Z(n5604) );
  NAND U5905 ( .A(n5605), .B(n5604), .Z(n5630) );
  XNOR U5906 ( .A(b[3]), .B(a[132]), .Z(n5645) );
  NANDN U5907 ( .A(n5645), .B(n10398), .Z(n5608) );
  NANDN U5908 ( .A(n5606), .B(n10399), .Z(n5607) );
  AND U5909 ( .A(n5608), .B(n5607), .Z(n5631) );
  XNOR U5910 ( .A(n5630), .B(n5631), .Z(n5632) );
  NANDN U5911 ( .A(n527), .B(a[134]), .Z(n5609) );
  XOR U5912 ( .A(n10434), .B(n5609), .Z(n5611) );
  NANDN U5913 ( .A(b[0]), .B(a[133]), .Z(n5610) );
  AND U5914 ( .A(n5611), .B(n5610), .Z(n5638) );
  XOR U5915 ( .A(b[5]), .B(a[130]), .Z(n5651) );
  NAND U5916 ( .A(n5651), .B(n10481), .Z(n5614) );
  NAND U5917 ( .A(n5612), .B(n10482), .Z(n5613) );
  NAND U5918 ( .A(n5614), .B(n5613), .Z(n5636) );
  NANDN U5919 ( .A(n529), .B(a[126]), .Z(n5637) );
  XNOR U5920 ( .A(n5636), .B(n5637), .Z(n5639) );
  XOR U5921 ( .A(n5638), .B(n5639), .Z(n5633) );
  XOR U5922 ( .A(n5632), .B(n5633), .Z(n5654) );
  XOR U5923 ( .A(n5655), .B(n5654), .Z(n5656) );
  XNOR U5924 ( .A(n5657), .B(n5656), .Z(n5626) );
  NAND U5925 ( .A(n5616), .B(n5615), .Z(n5620) );
  NAND U5926 ( .A(n5618), .B(n5617), .Z(n5619) );
  NAND U5927 ( .A(n5620), .B(n5619), .Z(n5627) );
  XNOR U5928 ( .A(n5626), .B(n5627), .Z(n5628) );
  XNOR U5929 ( .A(n5629), .B(n5628), .Z(n5660) );
  XNOR U5930 ( .A(n5660), .B(sreg[382]), .Z(n5662) );
  NAND U5931 ( .A(n5621), .B(sreg[381]), .Z(n5625) );
  OR U5932 ( .A(n5623), .B(n5622), .Z(n5624) );
  AND U5933 ( .A(n5625), .B(n5624), .Z(n5661) );
  XOR U5934 ( .A(n5662), .B(n5661), .Z(c[382]) );
  NANDN U5935 ( .A(n5631), .B(n5630), .Z(n5635) );
  NAND U5936 ( .A(n5633), .B(n5632), .Z(n5634) );
  NAND U5937 ( .A(n5635), .B(n5634), .Z(n5696) );
  NANDN U5938 ( .A(n5637), .B(n5636), .Z(n5641) );
  NAND U5939 ( .A(n5639), .B(n5638), .Z(n5640) );
  NAND U5940 ( .A(n5641), .B(n5640), .Z(n5694) );
  XNOR U5941 ( .A(b[7]), .B(a[129]), .Z(n5681) );
  NANDN U5942 ( .A(n5681), .B(n10545), .Z(n5644) );
  NANDN U5943 ( .A(n5642), .B(n10546), .Z(n5643) );
  NAND U5944 ( .A(n5644), .B(n5643), .Z(n5669) );
  XNOR U5945 ( .A(b[3]), .B(a[133]), .Z(n5684) );
  NANDN U5946 ( .A(n5684), .B(n10398), .Z(n5647) );
  NANDN U5947 ( .A(n5645), .B(n10399), .Z(n5646) );
  AND U5948 ( .A(n5647), .B(n5646), .Z(n5670) );
  XNOR U5949 ( .A(n5669), .B(n5670), .Z(n5671) );
  NANDN U5950 ( .A(n527), .B(a[135]), .Z(n5648) );
  XOR U5951 ( .A(n10434), .B(n5648), .Z(n5650) );
  NANDN U5952 ( .A(b[0]), .B(a[134]), .Z(n5649) );
  AND U5953 ( .A(n5650), .B(n5649), .Z(n5677) );
  XOR U5954 ( .A(b[5]), .B(a[131]), .Z(n5690) );
  NAND U5955 ( .A(n5690), .B(n10481), .Z(n5653) );
  NAND U5956 ( .A(n5651), .B(n10482), .Z(n5652) );
  NAND U5957 ( .A(n5653), .B(n5652), .Z(n5675) );
  NANDN U5958 ( .A(n529), .B(a[127]), .Z(n5676) );
  XNOR U5959 ( .A(n5675), .B(n5676), .Z(n5678) );
  XOR U5960 ( .A(n5677), .B(n5678), .Z(n5672) );
  XOR U5961 ( .A(n5671), .B(n5672), .Z(n5693) );
  XOR U5962 ( .A(n5694), .B(n5693), .Z(n5695) );
  XNOR U5963 ( .A(n5696), .B(n5695), .Z(n5665) );
  NAND U5964 ( .A(n5655), .B(n5654), .Z(n5659) );
  NAND U5965 ( .A(n5657), .B(n5656), .Z(n5658) );
  NAND U5966 ( .A(n5659), .B(n5658), .Z(n5666) );
  XNOR U5967 ( .A(n5665), .B(n5666), .Z(n5667) );
  XNOR U5968 ( .A(n5668), .B(n5667), .Z(n5699) );
  XNOR U5969 ( .A(n5699), .B(sreg[383]), .Z(n5701) );
  NAND U5970 ( .A(n5660), .B(sreg[382]), .Z(n5664) );
  OR U5971 ( .A(n5662), .B(n5661), .Z(n5663) );
  AND U5972 ( .A(n5664), .B(n5663), .Z(n5700) );
  XOR U5973 ( .A(n5701), .B(n5700), .Z(c[383]) );
  NANDN U5974 ( .A(n5670), .B(n5669), .Z(n5674) );
  NAND U5975 ( .A(n5672), .B(n5671), .Z(n5673) );
  NAND U5976 ( .A(n5674), .B(n5673), .Z(n5735) );
  NANDN U5977 ( .A(n5676), .B(n5675), .Z(n5680) );
  NAND U5978 ( .A(n5678), .B(n5677), .Z(n5679) );
  NAND U5979 ( .A(n5680), .B(n5679), .Z(n5733) );
  XNOR U5980 ( .A(b[7]), .B(a[130]), .Z(n5720) );
  NANDN U5981 ( .A(n5720), .B(n10545), .Z(n5683) );
  NANDN U5982 ( .A(n5681), .B(n10546), .Z(n5682) );
  NAND U5983 ( .A(n5683), .B(n5682), .Z(n5708) );
  XNOR U5984 ( .A(b[3]), .B(a[134]), .Z(n5723) );
  NANDN U5985 ( .A(n5723), .B(n10398), .Z(n5686) );
  NANDN U5986 ( .A(n5684), .B(n10399), .Z(n5685) );
  AND U5987 ( .A(n5686), .B(n5685), .Z(n5709) );
  XNOR U5988 ( .A(n5708), .B(n5709), .Z(n5710) );
  NANDN U5989 ( .A(n527), .B(a[136]), .Z(n5687) );
  XOR U5990 ( .A(n10434), .B(n5687), .Z(n5689) );
  NANDN U5991 ( .A(b[0]), .B(a[135]), .Z(n5688) );
  AND U5992 ( .A(n5689), .B(n5688), .Z(n5716) );
  XOR U5993 ( .A(b[5]), .B(a[132]), .Z(n5729) );
  NAND U5994 ( .A(n5729), .B(n10481), .Z(n5692) );
  NAND U5995 ( .A(n5690), .B(n10482), .Z(n5691) );
  NAND U5996 ( .A(n5692), .B(n5691), .Z(n5714) );
  NANDN U5997 ( .A(n529), .B(a[128]), .Z(n5715) );
  XNOR U5998 ( .A(n5714), .B(n5715), .Z(n5717) );
  XOR U5999 ( .A(n5716), .B(n5717), .Z(n5711) );
  XOR U6000 ( .A(n5710), .B(n5711), .Z(n5732) );
  XOR U6001 ( .A(n5733), .B(n5732), .Z(n5734) );
  XNOR U6002 ( .A(n5735), .B(n5734), .Z(n5704) );
  NAND U6003 ( .A(n5694), .B(n5693), .Z(n5698) );
  NAND U6004 ( .A(n5696), .B(n5695), .Z(n5697) );
  NAND U6005 ( .A(n5698), .B(n5697), .Z(n5705) );
  XNOR U6006 ( .A(n5704), .B(n5705), .Z(n5706) );
  XNOR U6007 ( .A(n5707), .B(n5706), .Z(n5738) );
  XNOR U6008 ( .A(n5738), .B(sreg[384]), .Z(n5740) );
  NAND U6009 ( .A(n5699), .B(sreg[383]), .Z(n5703) );
  OR U6010 ( .A(n5701), .B(n5700), .Z(n5702) );
  AND U6011 ( .A(n5703), .B(n5702), .Z(n5739) );
  XOR U6012 ( .A(n5740), .B(n5739), .Z(c[384]) );
  NANDN U6013 ( .A(n5709), .B(n5708), .Z(n5713) );
  NAND U6014 ( .A(n5711), .B(n5710), .Z(n5712) );
  NAND U6015 ( .A(n5713), .B(n5712), .Z(n5774) );
  NANDN U6016 ( .A(n5715), .B(n5714), .Z(n5719) );
  NAND U6017 ( .A(n5717), .B(n5716), .Z(n5718) );
  NAND U6018 ( .A(n5719), .B(n5718), .Z(n5772) );
  XNOR U6019 ( .A(b[7]), .B(a[131]), .Z(n5759) );
  NANDN U6020 ( .A(n5759), .B(n10545), .Z(n5722) );
  NANDN U6021 ( .A(n5720), .B(n10546), .Z(n5721) );
  NAND U6022 ( .A(n5722), .B(n5721), .Z(n5747) );
  XNOR U6023 ( .A(b[3]), .B(a[135]), .Z(n5762) );
  NANDN U6024 ( .A(n5762), .B(n10398), .Z(n5725) );
  NANDN U6025 ( .A(n5723), .B(n10399), .Z(n5724) );
  AND U6026 ( .A(n5725), .B(n5724), .Z(n5748) );
  XNOR U6027 ( .A(n5747), .B(n5748), .Z(n5749) );
  NANDN U6028 ( .A(n527), .B(a[137]), .Z(n5726) );
  XOR U6029 ( .A(n10434), .B(n5726), .Z(n5728) );
  NANDN U6030 ( .A(b[0]), .B(a[136]), .Z(n5727) );
  AND U6031 ( .A(n5728), .B(n5727), .Z(n5755) );
  XOR U6032 ( .A(b[5]), .B(a[133]), .Z(n5768) );
  NAND U6033 ( .A(n5768), .B(n10481), .Z(n5731) );
  NAND U6034 ( .A(n5729), .B(n10482), .Z(n5730) );
  NAND U6035 ( .A(n5731), .B(n5730), .Z(n5753) );
  NANDN U6036 ( .A(n529), .B(a[129]), .Z(n5754) );
  XNOR U6037 ( .A(n5753), .B(n5754), .Z(n5756) );
  XOR U6038 ( .A(n5755), .B(n5756), .Z(n5750) );
  XOR U6039 ( .A(n5749), .B(n5750), .Z(n5771) );
  XOR U6040 ( .A(n5772), .B(n5771), .Z(n5773) );
  XNOR U6041 ( .A(n5774), .B(n5773), .Z(n5743) );
  NAND U6042 ( .A(n5733), .B(n5732), .Z(n5737) );
  NAND U6043 ( .A(n5735), .B(n5734), .Z(n5736) );
  NAND U6044 ( .A(n5737), .B(n5736), .Z(n5744) );
  XNOR U6045 ( .A(n5743), .B(n5744), .Z(n5745) );
  XNOR U6046 ( .A(n5746), .B(n5745), .Z(n5777) );
  XNOR U6047 ( .A(n5777), .B(sreg[385]), .Z(n5779) );
  NAND U6048 ( .A(n5738), .B(sreg[384]), .Z(n5742) );
  OR U6049 ( .A(n5740), .B(n5739), .Z(n5741) );
  AND U6050 ( .A(n5742), .B(n5741), .Z(n5778) );
  XOR U6051 ( .A(n5779), .B(n5778), .Z(c[385]) );
  NANDN U6052 ( .A(n5748), .B(n5747), .Z(n5752) );
  NAND U6053 ( .A(n5750), .B(n5749), .Z(n5751) );
  NAND U6054 ( .A(n5752), .B(n5751), .Z(n5813) );
  NANDN U6055 ( .A(n5754), .B(n5753), .Z(n5758) );
  NAND U6056 ( .A(n5756), .B(n5755), .Z(n5757) );
  NAND U6057 ( .A(n5758), .B(n5757), .Z(n5811) );
  XNOR U6058 ( .A(b[7]), .B(a[132]), .Z(n5798) );
  NANDN U6059 ( .A(n5798), .B(n10545), .Z(n5761) );
  NANDN U6060 ( .A(n5759), .B(n10546), .Z(n5760) );
  NAND U6061 ( .A(n5761), .B(n5760), .Z(n5786) );
  XNOR U6062 ( .A(b[3]), .B(a[136]), .Z(n5801) );
  NANDN U6063 ( .A(n5801), .B(n10398), .Z(n5764) );
  NANDN U6064 ( .A(n5762), .B(n10399), .Z(n5763) );
  AND U6065 ( .A(n5764), .B(n5763), .Z(n5787) );
  XNOR U6066 ( .A(n5786), .B(n5787), .Z(n5788) );
  NANDN U6067 ( .A(n527), .B(a[138]), .Z(n5765) );
  XOR U6068 ( .A(n10434), .B(n5765), .Z(n5767) );
  NANDN U6069 ( .A(b[0]), .B(a[137]), .Z(n5766) );
  AND U6070 ( .A(n5767), .B(n5766), .Z(n5794) );
  XOR U6071 ( .A(b[5]), .B(a[134]), .Z(n5807) );
  NAND U6072 ( .A(n5807), .B(n10481), .Z(n5770) );
  NAND U6073 ( .A(n5768), .B(n10482), .Z(n5769) );
  NAND U6074 ( .A(n5770), .B(n5769), .Z(n5792) );
  NANDN U6075 ( .A(n529), .B(a[130]), .Z(n5793) );
  XNOR U6076 ( .A(n5792), .B(n5793), .Z(n5795) );
  XOR U6077 ( .A(n5794), .B(n5795), .Z(n5789) );
  XOR U6078 ( .A(n5788), .B(n5789), .Z(n5810) );
  XOR U6079 ( .A(n5811), .B(n5810), .Z(n5812) );
  XNOR U6080 ( .A(n5813), .B(n5812), .Z(n5782) );
  NAND U6081 ( .A(n5772), .B(n5771), .Z(n5776) );
  NAND U6082 ( .A(n5774), .B(n5773), .Z(n5775) );
  NAND U6083 ( .A(n5776), .B(n5775), .Z(n5783) );
  XNOR U6084 ( .A(n5782), .B(n5783), .Z(n5784) );
  XNOR U6085 ( .A(n5785), .B(n5784), .Z(n5816) );
  XNOR U6086 ( .A(n5816), .B(sreg[386]), .Z(n5818) );
  NAND U6087 ( .A(n5777), .B(sreg[385]), .Z(n5781) );
  OR U6088 ( .A(n5779), .B(n5778), .Z(n5780) );
  AND U6089 ( .A(n5781), .B(n5780), .Z(n5817) );
  XOR U6090 ( .A(n5818), .B(n5817), .Z(c[386]) );
  NANDN U6091 ( .A(n5787), .B(n5786), .Z(n5791) );
  NAND U6092 ( .A(n5789), .B(n5788), .Z(n5790) );
  NAND U6093 ( .A(n5791), .B(n5790), .Z(n5852) );
  NANDN U6094 ( .A(n5793), .B(n5792), .Z(n5797) );
  NAND U6095 ( .A(n5795), .B(n5794), .Z(n5796) );
  NAND U6096 ( .A(n5797), .B(n5796), .Z(n5850) );
  XNOR U6097 ( .A(b[7]), .B(a[133]), .Z(n5837) );
  NANDN U6098 ( .A(n5837), .B(n10545), .Z(n5800) );
  NANDN U6099 ( .A(n5798), .B(n10546), .Z(n5799) );
  NAND U6100 ( .A(n5800), .B(n5799), .Z(n5825) );
  XNOR U6101 ( .A(b[3]), .B(a[137]), .Z(n5840) );
  NANDN U6102 ( .A(n5840), .B(n10398), .Z(n5803) );
  NANDN U6103 ( .A(n5801), .B(n10399), .Z(n5802) );
  AND U6104 ( .A(n5803), .B(n5802), .Z(n5826) );
  XNOR U6105 ( .A(n5825), .B(n5826), .Z(n5827) );
  NANDN U6106 ( .A(n527), .B(a[139]), .Z(n5804) );
  XOR U6107 ( .A(n10434), .B(n5804), .Z(n5806) );
  NANDN U6108 ( .A(b[0]), .B(a[138]), .Z(n5805) );
  AND U6109 ( .A(n5806), .B(n5805), .Z(n5833) );
  XOR U6110 ( .A(b[5]), .B(a[135]), .Z(n5846) );
  NAND U6111 ( .A(n5846), .B(n10481), .Z(n5809) );
  NAND U6112 ( .A(n5807), .B(n10482), .Z(n5808) );
  NAND U6113 ( .A(n5809), .B(n5808), .Z(n5831) );
  NANDN U6114 ( .A(n529), .B(a[131]), .Z(n5832) );
  XNOR U6115 ( .A(n5831), .B(n5832), .Z(n5834) );
  XOR U6116 ( .A(n5833), .B(n5834), .Z(n5828) );
  XOR U6117 ( .A(n5827), .B(n5828), .Z(n5849) );
  XOR U6118 ( .A(n5850), .B(n5849), .Z(n5851) );
  XNOR U6119 ( .A(n5852), .B(n5851), .Z(n5821) );
  NAND U6120 ( .A(n5811), .B(n5810), .Z(n5815) );
  NAND U6121 ( .A(n5813), .B(n5812), .Z(n5814) );
  NAND U6122 ( .A(n5815), .B(n5814), .Z(n5822) );
  XNOR U6123 ( .A(n5821), .B(n5822), .Z(n5823) );
  XNOR U6124 ( .A(n5824), .B(n5823), .Z(n5855) );
  XNOR U6125 ( .A(n5855), .B(sreg[387]), .Z(n5857) );
  NAND U6126 ( .A(n5816), .B(sreg[386]), .Z(n5820) );
  OR U6127 ( .A(n5818), .B(n5817), .Z(n5819) );
  AND U6128 ( .A(n5820), .B(n5819), .Z(n5856) );
  XOR U6129 ( .A(n5857), .B(n5856), .Z(c[387]) );
  NANDN U6130 ( .A(n5826), .B(n5825), .Z(n5830) );
  NAND U6131 ( .A(n5828), .B(n5827), .Z(n5829) );
  NAND U6132 ( .A(n5830), .B(n5829), .Z(n5891) );
  NANDN U6133 ( .A(n5832), .B(n5831), .Z(n5836) );
  NAND U6134 ( .A(n5834), .B(n5833), .Z(n5835) );
  NAND U6135 ( .A(n5836), .B(n5835), .Z(n5889) );
  XNOR U6136 ( .A(b[7]), .B(a[134]), .Z(n5876) );
  NANDN U6137 ( .A(n5876), .B(n10545), .Z(n5839) );
  NANDN U6138 ( .A(n5837), .B(n10546), .Z(n5838) );
  NAND U6139 ( .A(n5839), .B(n5838), .Z(n5864) );
  XNOR U6140 ( .A(b[3]), .B(a[138]), .Z(n5879) );
  NANDN U6141 ( .A(n5879), .B(n10398), .Z(n5842) );
  NANDN U6142 ( .A(n5840), .B(n10399), .Z(n5841) );
  AND U6143 ( .A(n5842), .B(n5841), .Z(n5865) );
  XNOR U6144 ( .A(n5864), .B(n5865), .Z(n5866) );
  NANDN U6145 ( .A(n527), .B(a[140]), .Z(n5843) );
  XOR U6146 ( .A(n10434), .B(n5843), .Z(n5845) );
  NANDN U6147 ( .A(b[0]), .B(a[139]), .Z(n5844) );
  AND U6148 ( .A(n5845), .B(n5844), .Z(n5872) );
  XOR U6149 ( .A(b[5]), .B(a[136]), .Z(n5885) );
  NAND U6150 ( .A(n5885), .B(n10481), .Z(n5848) );
  NAND U6151 ( .A(n5846), .B(n10482), .Z(n5847) );
  NAND U6152 ( .A(n5848), .B(n5847), .Z(n5870) );
  NANDN U6153 ( .A(n529), .B(a[132]), .Z(n5871) );
  XNOR U6154 ( .A(n5870), .B(n5871), .Z(n5873) );
  XOR U6155 ( .A(n5872), .B(n5873), .Z(n5867) );
  XOR U6156 ( .A(n5866), .B(n5867), .Z(n5888) );
  XOR U6157 ( .A(n5889), .B(n5888), .Z(n5890) );
  XNOR U6158 ( .A(n5891), .B(n5890), .Z(n5860) );
  NAND U6159 ( .A(n5850), .B(n5849), .Z(n5854) );
  NAND U6160 ( .A(n5852), .B(n5851), .Z(n5853) );
  NAND U6161 ( .A(n5854), .B(n5853), .Z(n5861) );
  XNOR U6162 ( .A(n5860), .B(n5861), .Z(n5862) );
  XNOR U6163 ( .A(n5863), .B(n5862), .Z(n5894) );
  XNOR U6164 ( .A(n5894), .B(sreg[388]), .Z(n5896) );
  NAND U6165 ( .A(n5855), .B(sreg[387]), .Z(n5859) );
  OR U6166 ( .A(n5857), .B(n5856), .Z(n5858) );
  AND U6167 ( .A(n5859), .B(n5858), .Z(n5895) );
  XOR U6168 ( .A(n5896), .B(n5895), .Z(c[388]) );
  NANDN U6169 ( .A(n5865), .B(n5864), .Z(n5869) );
  NAND U6170 ( .A(n5867), .B(n5866), .Z(n5868) );
  NAND U6171 ( .A(n5869), .B(n5868), .Z(n5930) );
  NANDN U6172 ( .A(n5871), .B(n5870), .Z(n5875) );
  NAND U6173 ( .A(n5873), .B(n5872), .Z(n5874) );
  NAND U6174 ( .A(n5875), .B(n5874), .Z(n5928) );
  XNOR U6175 ( .A(b[7]), .B(a[135]), .Z(n5915) );
  NANDN U6176 ( .A(n5915), .B(n10545), .Z(n5878) );
  NANDN U6177 ( .A(n5876), .B(n10546), .Z(n5877) );
  NAND U6178 ( .A(n5878), .B(n5877), .Z(n5903) );
  XNOR U6179 ( .A(b[3]), .B(a[139]), .Z(n5918) );
  NANDN U6180 ( .A(n5918), .B(n10398), .Z(n5881) );
  NANDN U6181 ( .A(n5879), .B(n10399), .Z(n5880) );
  AND U6182 ( .A(n5881), .B(n5880), .Z(n5904) );
  XNOR U6183 ( .A(n5903), .B(n5904), .Z(n5905) );
  NANDN U6184 ( .A(n527), .B(a[141]), .Z(n5882) );
  XOR U6185 ( .A(n10434), .B(n5882), .Z(n5884) );
  NANDN U6186 ( .A(b[0]), .B(a[140]), .Z(n5883) );
  AND U6187 ( .A(n5884), .B(n5883), .Z(n5911) );
  XOR U6188 ( .A(b[5]), .B(a[137]), .Z(n5924) );
  NAND U6189 ( .A(n5924), .B(n10481), .Z(n5887) );
  NAND U6190 ( .A(n5885), .B(n10482), .Z(n5886) );
  NAND U6191 ( .A(n5887), .B(n5886), .Z(n5909) );
  NANDN U6192 ( .A(n529), .B(a[133]), .Z(n5910) );
  XNOR U6193 ( .A(n5909), .B(n5910), .Z(n5912) );
  XOR U6194 ( .A(n5911), .B(n5912), .Z(n5906) );
  XOR U6195 ( .A(n5905), .B(n5906), .Z(n5927) );
  XOR U6196 ( .A(n5928), .B(n5927), .Z(n5929) );
  XNOR U6197 ( .A(n5930), .B(n5929), .Z(n5899) );
  NAND U6198 ( .A(n5889), .B(n5888), .Z(n5893) );
  NAND U6199 ( .A(n5891), .B(n5890), .Z(n5892) );
  NAND U6200 ( .A(n5893), .B(n5892), .Z(n5900) );
  XNOR U6201 ( .A(n5899), .B(n5900), .Z(n5901) );
  XNOR U6202 ( .A(n5902), .B(n5901), .Z(n5933) );
  XNOR U6203 ( .A(n5933), .B(sreg[389]), .Z(n5935) );
  NAND U6204 ( .A(n5894), .B(sreg[388]), .Z(n5898) );
  OR U6205 ( .A(n5896), .B(n5895), .Z(n5897) );
  AND U6206 ( .A(n5898), .B(n5897), .Z(n5934) );
  XOR U6207 ( .A(n5935), .B(n5934), .Z(c[389]) );
  NANDN U6208 ( .A(n5904), .B(n5903), .Z(n5908) );
  NAND U6209 ( .A(n5906), .B(n5905), .Z(n5907) );
  NAND U6210 ( .A(n5908), .B(n5907), .Z(n5969) );
  NANDN U6211 ( .A(n5910), .B(n5909), .Z(n5914) );
  NAND U6212 ( .A(n5912), .B(n5911), .Z(n5913) );
  NAND U6213 ( .A(n5914), .B(n5913), .Z(n5967) );
  XNOR U6214 ( .A(b[7]), .B(a[136]), .Z(n5954) );
  NANDN U6215 ( .A(n5954), .B(n10545), .Z(n5917) );
  NANDN U6216 ( .A(n5915), .B(n10546), .Z(n5916) );
  NAND U6217 ( .A(n5917), .B(n5916), .Z(n5942) );
  XNOR U6218 ( .A(b[3]), .B(a[140]), .Z(n5957) );
  NANDN U6219 ( .A(n5957), .B(n10398), .Z(n5920) );
  NANDN U6220 ( .A(n5918), .B(n10399), .Z(n5919) );
  AND U6221 ( .A(n5920), .B(n5919), .Z(n5943) );
  XNOR U6222 ( .A(n5942), .B(n5943), .Z(n5944) );
  NANDN U6223 ( .A(n527), .B(a[142]), .Z(n5921) );
  XOR U6224 ( .A(n10434), .B(n5921), .Z(n5923) );
  NANDN U6225 ( .A(b[0]), .B(a[141]), .Z(n5922) );
  AND U6226 ( .A(n5923), .B(n5922), .Z(n5950) );
  XOR U6227 ( .A(b[5]), .B(a[138]), .Z(n5963) );
  NAND U6228 ( .A(n5963), .B(n10481), .Z(n5926) );
  NAND U6229 ( .A(n5924), .B(n10482), .Z(n5925) );
  NAND U6230 ( .A(n5926), .B(n5925), .Z(n5948) );
  NANDN U6231 ( .A(n529), .B(a[134]), .Z(n5949) );
  XNOR U6232 ( .A(n5948), .B(n5949), .Z(n5951) );
  XOR U6233 ( .A(n5950), .B(n5951), .Z(n5945) );
  XOR U6234 ( .A(n5944), .B(n5945), .Z(n5966) );
  XOR U6235 ( .A(n5967), .B(n5966), .Z(n5968) );
  XNOR U6236 ( .A(n5969), .B(n5968), .Z(n5938) );
  NAND U6237 ( .A(n5928), .B(n5927), .Z(n5932) );
  NAND U6238 ( .A(n5930), .B(n5929), .Z(n5931) );
  NAND U6239 ( .A(n5932), .B(n5931), .Z(n5939) );
  XNOR U6240 ( .A(n5938), .B(n5939), .Z(n5940) );
  XNOR U6241 ( .A(n5941), .B(n5940), .Z(n5972) );
  XNOR U6242 ( .A(n5972), .B(sreg[390]), .Z(n5974) );
  NAND U6243 ( .A(n5933), .B(sreg[389]), .Z(n5937) );
  OR U6244 ( .A(n5935), .B(n5934), .Z(n5936) );
  AND U6245 ( .A(n5937), .B(n5936), .Z(n5973) );
  XOR U6246 ( .A(n5974), .B(n5973), .Z(c[390]) );
  NANDN U6247 ( .A(n5943), .B(n5942), .Z(n5947) );
  NAND U6248 ( .A(n5945), .B(n5944), .Z(n5946) );
  NAND U6249 ( .A(n5947), .B(n5946), .Z(n6008) );
  NANDN U6250 ( .A(n5949), .B(n5948), .Z(n5953) );
  NAND U6251 ( .A(n5951), .B(n5950), .Z(n5952) );
  NAND U6252 ( .A(n5953), .B(n5952), .Z(n6006) );
  XNOR U6253 ( .A(b[7]), .B(a[137]), .Z(n5993) );
  NANDN U6254 ( .A(n5993), .B(n10545), .Z(n5956) );
  NANDN U6255 ( .A(n5954), .B(n10546), .Z(n5955) );
  NAND U6256 ( .A(n5956), .B(n5955), .Z(n5981) );
  XNOR U6257 ( .A(b[3]), .B(a[141]), .Z(n5996) );
  NANDN U6258 ( .A(n5996), .B(n10398), .Z(n5959) );
  NANDN U6259 ( .A(n5957), .B(n10399), .Z(n5958) );
  AND U6260 ( .A(n5959), .B(n5958), .Z(n5982) );
  XNOR U6261 ( .A(n5981), .B(n5982), .Z(n5983) );
  NANDN U6262 ( .A(n527), .B(a[143]), .Z(n5960) );
  XOR U6263 ( .A(n10434), .B(n5960), .Z(n5962) );
  NANDN U6264 ( .A(b[0]), .B(a[142]), .Z(n5961) );
  AND U6265 ( .A(n5962), .B(n5961), .Z(n5989) );
  XOR U6266 ( .A(b[5]), .B(a[139]), .Z(n6002) );
  NAND U6267 ( .A(n6002), .B(n10481), .Z(n5965) );
  NAND U6268 ( .A(n5963), .B(n10482), .Z(n5964) );
  NAND U6269 ( .A(n5965), .B(n5964), .Z(n5987) );
  NANDN U6270 ( .A(n529), .B(a[135]), .Z(n5988) );
  XNOR U6271 ( .A(n5987), .B(n5988), .Z(n5990) );
  XOR U6272 ( .A(n5989), .B(n5990), .Z(n5984) );
  XOR U6273 ( .A(n5983), .B(n5984), .Z(n6005) );
  XOR U6274 ( .A(n6006), .B(n6005), .Z(n6007) );
  XNOR U6275 ( .A(n6008), .B(n6007), .Z(n5977) );
  NAND U6276 ( .A(n5967), .B(n5966), .Z(n5971) );
  NAND U6277 ( .A(n5969), .B(n5968), .Z(n5970) );
  NAND U6278 ( .A(n5971), .B(n5970), .Z(n5978) );
  XNOR U6279 ( .A(n5977), .B(n5978), .Z(n5979) );
  XNOR U6280 ( .A(n5980), .B(n5979), .Z(n6011) );
  XNOR U6281 ( .A(n6011), .B(sreg[391]), .Z(n6013) );
  NAND U6282 ( .A(n5972), .B(sreg[390]), .Z(n5976) );
  OR U6283 ( .A(n5974), .B(n5973), .Z(n5975) );
  AND U6284 ( .A(n5976), .B(n5975), .Z(n6012) );
  XOR U6285 ( .A(n6013), .B(n6012), .Z(c[391]) );
  NANDN U6286 ( .A(n5982), .B(n5981), .Z(n5986) );
  NAND U6287 ( .A(n5984), .B(n5983), .Z(n5985) );
  NAND U6288 ( .A(n5986), .B(n5985), .Z(n6047) );
  NANDN U6289 ( .A(n5988), .B(n5987), .Z(n5992) );
  NAND U6290 ( .A(n5990), .B(n5989), .Z(n5991) );
  NAND U6291 ( .A(n5992), .B(n5991), .Z(n6045) );
  XNOR U6292 ( .A(b[7]), .B(a[138]), .Z(n6032) );
  NANDN U6293 ( .A(n6032), .B(n10545), .Z(n5995) );
  NANDN U6294 ( .A(n5993), .B(n10546), .Z(n5994) );
  NAND U6295 ( .A(n5995), .B(n5994), .Z(n6020) );
  XNOR U6296 ( .A(b[3]), .B(a[142]), .Z(n6035) );
  NANDN U6297 ( .A(n6035), .B(n10398), .Z(n5998) );
  NANDN U6298 ( .A(n5996), .B(n10399), .Z(n5997) );
  AND U6299 ( .A(n5998), .B(n5997), .Z(n6021) );
  XNOR U6300 ( .A(n6020), .B(n6021), .Z(n6022) );
  NANDN U6301 ( .A(n527), .B(a[144]), .Z(n5999) );
  XOR U6302 ( .A(n10434), .B(n5999), .Z(n6001) );
  NANDN U6303 ( .A(b[0]), .B(a[143]), .Z(n6000) );
  AND U6304 ( .A(n6001), .B(n6000), .Z(n6028) );
  XOR U6305 ( .A(b[5]), .B(a[140]), .Z(n6041) );
  NAND U6306 ( .A(n6041), .B(n10481), .Z(n6004) );
  NAND U6307 ( .A(n6002), .B(n10482), .Z(n6003) );
  NAND U6308 ( .A(n6004), .B(n6003), .Z(n6026) );
  NANDN U6309 ( .A(n529), .B(a[136]), .Z(n6027) );
  XNOR U6310 ( .A(n6026), .B(n6027), .Z(n6029) );
  XOR U6311 ( .A(n6028), .B(n6029), .Z(n6023) );
  XOR U6312 ( .A(n6022), .B(n6023), .Z(n6044) );
  XOR U6313 ( .A(n6045), .B(n6044), .Z(n6046) );
  XNOR U6314 ( .A(n6047), .B(n6046), .Z(n6016) );
  NAND U6315 ( .A(n6006), .B(n6005), .Z(n6010) );
  NAND U6316 ( .A(n6008), .B(n6007), .Z(n6009) );
  NAND U6317 ( .A(n6010), .B(n6009), .Z(n6017) );
  XNOR U6318 ( .A(n6016), .B(n6017), .Z(n6018) );
  XNOR U6319 ( .A(n6019), .B(n6018), .Z(n6050) );
  XNOR U6320 ( .A(n6050), .B(sreg[392]), .Z(n6052) );
  NAND U6321 ( .A(n6011), .B(sreg[391]), .Z(n6015) );
  OR U6322 ( .A(n6013), .B(n6012), .Z(n6014) );
  AND U6323 ( .A(n6015), .B(n6014), .Z(n6051) );
  XOR U6324 ( .A(n6052), .B(n6051), .Z(c[392]) );
  NANDN U6325 ( .A(n6021), .B(n6020), .Z(n6025) );
  NAND U6326 ( .A(n6023), .B(n6022), .Z(n6024) );
  NAND U6327 ( .A(n6025), .B(n6024), .Z(n6086) );
  NANDN U6328 ( .A(n6027), .B(n6026), .Z(n6031) );
  NAND U6329 ( .A(n6029), .B(n6028), .Z(n6030) );
  NAND U6330 ( .A(n6031), .B(n6030), .Z(n6084) );
  XNOR U6331 ( .A(b[7]), .B(a[139]), .Z(n6071) );
  NANDN U6332 ( .A(n6071), .B(n10545), .Z(n6034) );
  NANDN U6333 ( .A(n6032), .B(n10546), .Z(n6033) );
  NAND U6334 ( .A(n6034), .B(n6033), .Z(n6059) );
  XNOR U6335 ( .A(b[3]), .B(a[143]), .Z(n6074) );
  NANDN U6336 ( .A(n6074), .B(n10398), .Z(n6037) );
  NANDN U6337 ( .A(n6035), .B(n10399), .Z(n6036) );
  AND U6338 ( .A(n6037), .B(n6036), .Z(n6060) );
  XNOR U6339 ( .A(n6059), .B(n6060), .Z(n6061) );
  NANDN U6340 ( .A(n527), .B(a[145]), .Z(n6038) );
  XOR U6341 ( .A(n10434), .B(n6038), .Z(n6040) );
  NANDN U6342 ( .A(b[0]), .B(a[144]), .Z(n6039) );
  AND U6343 ( .A(n6040), .B(n6039), .Z(n6067) );
  XOR U6344 ( .A(b[5]), .B(a[141]), .Z(n6080) );
  NAND U6345 ( .A(n6080), .B(n10481), .Z(n6043) );
  NAND U6346 ( .A(n6041), .B(n10482), .Z(n6042) );
  NAND U6347 ( .A(n6043), .B(n6042), .Z(n6065) );
  NANDN U6348 ( .A(n529), .B(a[137]), .Z(n6066) );
  XNOR U6349 ( .A(n6065), .B(n6066), .Z(n6068) );
  XOR U6350 ( .A(n6067), .B(n6068), .Z(n6062) );
  XOR U6351 ( .A(n6061), .B(n6062), .Z(n6083) );
  XOR U6352 ( .A(n6084), .B(n6083), .Z(n6085) );
  XNOR U6353 ( .A(n6086), .B(n6085), .Z(n6055) );
  NAND U6354 ( .A(n6045), .B(n6044), .Z(n6049) );
  NAND U6355 ( .A(n6047), .B(n6046), .Z(n6048) );
  NAND U6356 ( .A(n6049), .B(n6048), .Z(n6056) );
  XNOR U6357 ( .A(n6055), .B(n6056), .Z(n6057) );
  XNOR U6358 ( .A(n6058), .B(n6057), .Z(n6089) );
  XNOR U6359 ( .A(n6089), .B(sreg[393]), .Z(n6091) );
  NAND U6360 ( .A(n6050), .B(sreg[392]), .Z(n6054) );
  OR U6361 ( .A(n6052), .B(n6051), .Z(n6053) );
  AND U6362 ( .A(n6054), .B(n6053), .Z(n6090) );
  XOR U6363 ( .A(n6091), .B(n6090), .Z(c[393]) );
  NANDN U6364 ( .A(n6060), .B(n6059), .Z(n6064) );
  NAND U6365 ( .A(n6062), .B(n6061), .Z(n6063) );
  NAND U6366 ( .A(n6064), .B(n6063), .Z(n6125) );
  NANDN U6367 ( .A(n6066), .B(n6065), .Z(n6070) );
  NAND U6368 ( .A(n6068), .B(n6067), .Z(n6069) );
  NAND U6369 ( .A(n6070), .B(n6069), .Z(n6123) );
  XNOR U6370 ( .A(b[7]), .B(a[140]), .Z(n6110) );
  NANDN U6371 ( .A(n6110), .B(n10545), .Z(n6073) );
  NANDN U6372 ( .A(n6071), .B(n10546), .Z(n6072) );
  NAND U6373 ( .A(n6073), .B(n6072), .Z(n6098) );
  XNOR U6374 ( .A(b[3]), .B(a[144]), .Z(n6113) );
  NANDN U6375 ( .A(n6113), .B(n10398), .Z(n6076) );
  NANDN U6376 ( .A(n6074), .B(n10399), .Z(n6075) );
  AND U6377 ( .A(n6076), .B(n6075), .Z(n6099) );
  XNOR U6378 ( .A(n6098), .B(n6099), .Z(n6100) );
  NANDN U6379 ( .A(n527), .B(a[146]), .Z(n6077) );
  XOR U6380 ( .A(n10434), .B(n6077), .Z(n6079) );
  NANDN U6381 ( .A(b[0]), .B(a[145]), .Z(n6078) );
  AND U6382 ( .A(n6079), .B(n6078), .Z(n6106) );
  XOR U6383 ( .A(b[5]), .B(a[142]), .Z(n6119) );
  NAND U6384 ( .A(n6119), .B(n10481), .Z(n6082) );
  NAND U6385 ( .A(n6080), .B(n10482), .Z(n6081) );
  NAND U6386 ( .A(n6082), .B(n6081), .Z(n6104) );
  NANDN U6387 ( .A(n529), .B(a[138]), .Z(n6105) );
  XNOR U6388 ( .A(n6104), .B(n6105), .Z(n6107) );
  XOR U6389 ( .A(n6106), .B(n6107), .Z(n6101) );
  XOR U6390 ( .A(n6100), .B(n6101), .Z(n6122) );
  XOR U6391 ( .A(n6123), .B(n6122), .Z(n6124) );
  XNOR U6392 ( .A(n6125), .B(n6124), .Z(n6094) );
  NAND U6393 ( .A(n6084), .B(n6083), .Z(n6088) );
  NAND U6394 ( .A(n6086), .B(n6085), .Z(n6087) );
  NAND U6395 ( .A(n6088), .B(n6087), .Z(n6095) );
  XNOR U6396 ( .A(n6094), .B(n6095), .Z(n6096) );
  XNOR U6397 ( .A(n6097), .B(n6096), .Z(n6128) );
  XNOR U6398 ( .A(n6128), .B(sreg[394]), .Z(n6130) );
  NAND U6399 ( .A(n6089), .B(sreg[393]), .Z(n6093) );
  OR U6400 ( .A(n6091), .B(n6090), .Z(n6092) );
  AND U6401 ( .A(n6093), .B(n6092), .Z(n6129) );
  XOR U6402 ( .A(n6130), .B(n6129), .Z(c[394]) );
  NANDN U6403 ( .A(n6099), .B(n6098), .Z(n6103) );
  NAND U6404 ( .A(n6101), .B(n6100), .Z(n6102) );
  NAND U6405 ( .A(n6103), .B(n6102), .Z(n6164) );
  NANDN U6406 ( .A(n6105), .B(n6104), .Z(n6109) );
  NAND U6407 ( .A(n6107), .B(n6106), .Z(n6108) );
  NAND U6408 ( .A(n6109), .B(n6108), .Z(n6162) );
  XNOR U6409 ( .A(b[7]), .B(a[141]), .Z(n6149) );
  NANDN U6410 ( .A(n6149), .B(n10545), .Z(n6112) );
  NANDN U6411 ( .A(n6110), .B(n10546), .Z(n6111) );
  NAND U6412 ( .A(n6112), .B(n6111), .Z(n6137) );
  XNOR U6413 ( .A(b[3]), .B(a[145]), .Z(n6152) );
  NANDN U6414 ( .A(n6152), .B(n10398), .Z(n6115) );
  NANDN U6415 ( .A(n6113), .B(n10399), .Z(n6114) );
  AND U6416 ( .A(n6115), .B(n6114), .Z(n6138) );
  XNOR U6417 ( .A(n6137), .B(n6138), .Z(n6139) );
  NANDN U6418 ( .A(n527), .B(a[147]), .Z(n6116) );
  XOR U6419 ( .A(n10434), .B(n6116), .Z(n6118) );
  NANDN U6420 ( .A(b[0]), .B(a[146]), .Z(n6117) );
  AND U6421 ( .A(n6118), .B(n6117), .Z(n6145) );
  XOR U6422 ( .A(b[5]), .B(a[143]), .Z(n6158) );
  NAND U6423 ( .A(n6158), .B(n10481), .Z(n6121) );
  NAND U6424 ( .A(n6119), .B(n10482), .Z(n6120) );
  NAND U6425 ( .A(n6121), .B(n6120), .Z(n6143) );
  NANDN U6426 ( .A(n529), .B(a[139]), .Z(n6144) );
  XNOR U6427 ( .A(n6143), .B(n6144), .Z(n6146) );
  XOR U6428 ( .A(n6145), .B(n6146), .Z(n6140) );
  XOR U6429 ( .A(n6139), .B(n6140), .Z(n6161) );
  XOR U6430 ( .A(n6162), .B(n6161), .Z(n6163) );
  XNOR U6431 ( .A(n6164), .B(n6163), .Z(n6133) );
  NAND U6432 ( .A(n6123), .B(n6122), .Z(n6127) );
  NAND U6433 ( .A(n6125), .B(n6124), .Z(n6126) );
  NAND U6434 ( .A(n6127), .B(n6126), .Z(n6134) );
  XNOR U6435 ( .A(n6133), .B(n6134), .Z(n6135) );
  XNOR U6436 ( .A(n6136), .B(n6135), .Z(n6167) );
  XNOR U6437 ( .A(n6167), .B(sreg[395]), .Z(n6169) );
  NAND U6438 ( .A(n6128), .B(sreg[394]), .Z(n6132) );
  OR U6439 ( .A(n6130), .B(n6129), .Z(n6131) );
  AND U6440 ( .A(n6132), .B(n6131), .Z(n6168) );
  XOR U6441 ( .A(n6169), .B(n6168), .Z(c[395]) );
  NANDN U6442 ( .A(n6138), .B(n6137), .Z(n6142) );
  NAND U6443 ( .A(n6140), .B(n6139), .Z(n6141) );
  NAND U6444 ( .A(n6142), .B(n6141), .Z(n6203) );
  NANDN U6445 ( .A(n6144), .B(n6143), .Z(n6148) );
  NAND U6446 ( .A(n6146), .B(n6145), .Z(n6147) );
  NAND U6447 ( .A(n6148), .B(n6147), .Z(n6201) );
  XNOR U6448 ( .A(b[7]), .B(a[142]), .Z(n6188) );
  NANDN U6449 ( .A(n6188), .B(n10545), .Z(n6151) );
  NANDN U6450 ( .A(n6149), .B(n10546), .Z(n6150) );
  NAND U6451 ( .A(n6151), .B(n6150), .Z(n6176) );
  XNOR U6452 ( .A(b[3]), .B(a[146]), .Z(n6191) );
  NANDN U6453 ( .A(n6191), .B(n10398), .Z(n6154) );
  NANDN U6454 ( .A(n6152), .B(n10399), .Z(n6153) );
  AND U6455 ( .A(n6154), .B(n6153), .Z(n6177) );
  XNOR U6456 ( .A(n6176), .B(n6177), .Z(n6178) );
  NANDN U6457 ( .A(n527), .B(a[148]), .Z(n6155) );
  XOR U6458 ( .A(n10434), .B(n6155), .Z(n6157) );
  NANDN U6459 ( .A(b[0]), .B(a[147]), .Z(n6156) );
  AND U6460 ( .A(n6157), .B(n6156), .Z(n6184) );
  XOR U6461 ( .A(b[5]), .B(a[144]), .Z(n6197) );
  NAND U6462 ( .A(n6197), .B(n10481), .Z(n6160) );
  NAND U6463 ( .A(n6158), .B(n10482), .Z(n6159) );
  NAND U6464 ( .A(n6160), .B(n6159), .Z(n6182) );
  NANDN U6465 ( .A(n529), .B(a[140]), .Z(n6183) );
  XNOR U6466 ( .A(n6182), .B(n6183), .Z(n6185) );
  XOR U6467 ( .A(n6184), .B(n6185), .Z(n6179) );
  XOR U6468 ( .A(n6178), .B(n6179), .Z(n6200) );
  XOR U6469 ( .A(n6201), .B(n6200), .Z(n6202) );
  XNOR U6470 ( .A(n6203), .B(n6202), .Z(n6172) );
  NAND U6471 ( .A(n6162), .B(n6161), .Z(n6166) );
  NAND U6472 ( .A(n6164), .B(n6163), .Z(n6165) );
  NAND U6473 ( .A(n6166), .B(n6165), .Z(n6173) );
  XNOR U6474 ( .A(n6172), .B(n6173), .Z(n6174) );
  XNOR U6475 ( .A(n6175), .B(n6174), .Z(n6206) );
  XNOR U6476 ( .A(n6206), .B(sreg[396]), .Z(n6208) );
  NAND U6477 ( .A(n6167), .B(sreg[395]), .Z(n6171) );
  OR U6478 ( .A(n6169), .B(n6168), .Z(n6170) );
  AND U6479 ( .A(n6171), .B(n6170), .Z(n6207) );
  XOR U6480 ( .A(n6208), .B(n6207), .Z(c[396]) );
  NANDN U6481 ( .A(n6177), .B(n6176), .Z(n6181) );
  NAND U6482 ( .A(n6179), .B(n6178), .Z(n6180) );
  NAND U6483 ( .A(n6181), .B(n6180), .Z(n6242) );
  NANDN U6484 ( .A(n6183), .B(n6182), .Z(n6187) );
  NAND U6485 ( .A(n6185), .B(n6184), .Z(n6186) );
  NAND U6486 ( .A(n6187), .B(n6186), .Z(n6240) );
  XNOR U6487 ( .A(b[7]), .B(a[143]), .Z(n6227) );
  NANDN U6488 ( .A(n6227), .B(n10545), .Z(n6190) );
  NANDN U6489 ( .A(n6188), .B(n10546), .Z(n6189) );
  NAND U6490 ( .A(n6190), .B(n6189), .Z(n6215) );
  XNOR U6491 ( .A(b[3]), .B(a[147]), .Z(n6230) );
  NANDN U6492 ( .A(n6230), .B(n10398), .Z(n6193) );
  NANDN U6493 ( .A(n6191), .B(n10399), .Z(n6192) );
  AND U6494 ( .A(n6193), .B(n6192), .Z(n6216) );
  XNOR U6495 ( .A(n6215), .B(n6216), .Z(n6217) );
  NANDN U6496 ( .A(n527), .B(a[149]), .Z(n6194) );
  XOR U6497 ( .A(n10434), .B(n6194), .Z(n6196) );
  NANDN U6498 ( .A(b[0]), .B(a[148]), .Z(n6195) );
  AND U6499 ( .A(n6196), .B(n6195), .Z(n6223) );
  XOR U6500 ( .A(b[5]), .B(a[145]), .Z(n6236) );
  NAND U6501 ( .A(n6236), .B(n10481), .Z(n6199) );
  NAND U6502 ( .A(n6197), .B(n10482), .Z(n6198) );
  NAND U6503 ( .A(n6199), .B(n6198), .Z(n6221) );
  NANDN U6504 ( .A(n529), .B(a[141]), .Z(n6222) );
  XNOR U6505 ( .A(n6221), .B(n6222), .Z(n6224) );
  XOR U6506 ( .A(n6223), .B(n6224), .Z(n6218) );
  XOR U6507 ( .A(n6217), .B(n6218), .Z(n6239) );
  XOR U6508 ( .A(n6240), .B(n6239), .Z(n6241) );
  XNOR U6509 ( .A(n6242), .B(n6241), .Z(n6211) );
  NAND U6510 ( .A(n6201), .B(n6200), .Z(n6205) );
  NAND U6511 ( .A(n6203), .B(n6202), .Z(n6204) );
  NAND U6512 ( .A(n6205), .B(n6204), .Z(n6212) );
  XNOR U6513 ( .A(n6211), .B(n6212), .Z(n6213) );
  XNOR U6514 ( .A(n6214), .B(n6213), .Z(n6245) );
  XNOR U6515 ( .A(n6245), .B(sreg[397]), .Z(n6247) );
  NAND U6516 ( .A(n6206), .B(sreg[396]), .Z(n6210) );
  OR U6517 ( .A(n6208), .B(n6207), .Z(n6209) );
  AND U6518 ( .A(n6210), .B(n6209), .Z(n6246) );
  XOR U6519 ( .A(n6247), .B(n6246), .Z(c[397]) );
  NANDN U6520 ( .A(n6216), .B(n6215), .Z(n6220) );
  NAND U6521 ( .A(n6218), .B(n6217), .Z(n6219) );
  NAND U6522 ( .A(n6220), .B(n6219), .Z(n6281) );
  NANDN U6523 ( .A(n6222), .B(n6221), .Z(n6226) );
  NAND U6524 ( .A(n6224), .B(n6223), .Z(n6225) );
  NAND U6525 ( .A(n6226), .B(n6225), .Z(n6279) );
  XNOR U6526 ( .A(b[7]), .B(a[144]), .Z(n6266) );
  NANDN U6527 ( .A(n6266), .B(n10545), .Z(n6229) );
  NANDN U6528 ( .A(n6227), .B(n10546), .Z(n6228) );
  NAND U6529 ( .A(n6229), .B(n6228), .Z(n6254) );
  XNOR U6530 ( .A(b[3]), .B(a[148]), .Z(n6269) );
  NANDN U6531 ( .A(n6269), .B(n10398), .Z(n6232) );
  NANDN U6532 ( .A(n6230), .B(n10399), .Z(n6231) );
  AND U6533 ( .A(n6232), .B(n6231), .Z(n6255) );
  XNOR U6534 ( .A(n6254), .B(n6255), .Z(n6256) );
  NANDN U6535 ( .A(n527), .B(a[150]), .Z(n6233) );
  XOR U6536 ( .A(n10434), .B(n6233), .Z(n6235) );
  NANDN U6537 ( .A(b[0]), .B(a[149]), .Z(n6234) );
  AND U6538 ( .A(n6235), .B(n6234), .Z(n6262) );
  XOR U6539 ( .A(b[5]), .B(a[146]), .Z(n6275) );
  NAND U6540 ( .A(n6275), .B(n10481), .Z(n6238) );
  NAND U6541 ( .A(n6236), .B(n10482), .Z(n6237) );
  NAND U6542 ( .A(n6238), .B(n6237), .Z(n6260) );
  NANDN U6543 ( .A(n529), .B(a[142]), .Z(n6261) );
  XNOR U6544 ( .A(n6260), .B(n6261), .Z(n6263) );
  XOR U6545 ( .A(n6262), .B(n6263), .Z(n6257) );
  XOR U6546 ( .A(n6256), .B(n6257), .Z(n6278) );
  XOR U6547 ( .A(n6279), .B(n6278), .Z(n6280) );
  XNOR U6548 ( .A(n6281), .B(n6280), .Z(n6250) );
  NAND U6549 ( .A(n6240), .B(n6239), .Z(n6244) );
  NAND U6550 ( .A(n6242), .B(n6241), .Z(n6243) );
  NAND U6551 ( .A(n6244), .B(n6243), .Z(n6251) );
  XNOR U6552 ( .A(n6250), .B(n6251), .Z(n6252) );
  XNOR U6553 ( .A(n6253), .B(n6252), .Z(n6284) );
  XNOR U6554 ( .A(n6284), .B(sreg[398]), .Z(n6286) );
  NAND U6555 ( .A(n6245), .B(sreg[397]), .Z(n6249) );
  OR U6556 ( .A(n6247), .B(n6246), .Z(n6248) );
  AND U6557 ( .A(n6249), .B(n6248), .Z(n6285) );
  XOR U6558 ( .A(n6286), .B(n6285), .Z(c[398]) );
  NANDN U6559 ( .A(n6255), .B(n6254), .Z(n6259) );
  NAND U6560 ( .A(n6257), .B(n6256), .Z(n6258) );
  NAND U6561 ( .A(n6259), .B(n6258), .Z(n6320) );
  NANDN U6562 ( .A(n6261), .B(n6260), .Z(n6265) );
  NAND U6563 ( .A(n6263), .B(n6262), .Z(n6264) );
  NAND U6564 ( .A(n6265), .B(n6264), .Z(n6318) );
  XNOR U6565 ( .A(b[7]), .B(a[145]), .Z(n6305) );
  NANDN U6566 ( .A(n6305), .B(n10545), .Z(n6268) );
  NANDN U6567 ( .A(n6266), .B(n10546), .Z(n6267) );
  NAND U6568 ( .A(n6268), .B(n6267), .Z(n6293) );
  XNOR U6569 ( .A(b[3]), .B(a[149]), .Z(n6308) );
  NANDN U6570 ( .A(n6308), .B(n10398), .Z(n6271) );
  NANDN U6571 ( .A(n6269), .B(n10399), .Z(n6270) );
  AND U6572 ( .A(n6271), .B(n6270), .Z(n6294) );
  XNOR U6573 ( .A(n6293), .B(n6294), .Z(n6295) );
  NANDN U6574 ( .A(n527), .B(a[151]), .Z(n6272) );
  XOR U6575 ( .A(n10434), .B(n6272), .Z(n6274) );
  NANDN U6576 ( .A(b[0]), .B(a[150]), .Z(n6273) );
  AND U6577 ( .A(n6274), .B(n6273), .Z(n6301) );
  XOR U6578 ( .A(b[5]), .B(a[147]), .Z(n6314) );
  NAND U6579 ( .A(n6314), .B(n10481), .Z(n6277) );
  NAND U6580 ( .A(n6275), .B(n10482), .Z(n6276) );
  NAND U6581 ( .A(n6277), .B(n6276), .Z(n6299) );
  NANDN U6582 ( .A(n529), .B(a[143]), .Z(n6300) );
  XNOR U6583 ( .A(n6299), .B(n6300), .Z(n6302) );
  XOR U6584 ( .A(n6301), .B(n6302), .Z(n6296) );
  XOR U6585 ( .A(n6295), .B(n6296), .Z(n6317) );
  XOR U6586 ( .A(n6318), .B(n6317), .Z(n6319) );
  XNOR U6587 ( .A(n6320), .B(n6319), .Z(n6289) );
  NAND U6588 ( .A(n6279), .B(n6278), .Z(n6283) );
  NAND U6589 ( .A(n6281), .B(n6280), .Z(n6282) );
  NAND U6590 ( .A(n6283), .B(n6282), .Z(n6290) );
  XNOR U6591 ( .A(n6289), .B(n6290), .Z(n6291) );
  XNOR U6592 ( .A(n6292), .B(n6291), .Z(n6323) );
  XNOR U6593 ( .A(n6323), .B(sreg[399]), .Z(n6325) );
  NAND U6594 ( .A(n6284), .B(sreg[398]), .Z(n6288) );
  OR U6595 ( .A(n6286), .B(n6285), .Z(n6287) );
  AND U6596 ( .A(n6288), .B(n6287), .Z(n6324) );
  XOR U6597 ( .A(n6325), .B(n6324), .Z(c[399]) );
  NANDN U6598 ( .A(n6294), .B(n6293), .Z(n6298) );
  NAND U6599 ( .A(n6296), .B(n6295), .Z(n6297) );
  NAND U6600 ( .A(n6298), .B(n6297), .Z(n6359) );
  NANDN U6601 ( .A(n6300), .B(n6299), .Z(n6304) );
  NAND U6602 ( .A(n6302), .B(n6301), .Z(n6303) );
  NAND U6603 ( .A(n6304), .B(n6303), .Z(n6357) );
  XNOR U6604 ( .A(b[7]), .B(a[146]), .Z(n6344) );
  NANDN U6605 ( .A(n6344), .B(n10545), .Z(n6307) );
  NANDN U6606 ( .A(n6305), .B(n10546), .Z(n6306) );
  NAND U6607 ( .A(n6307), .B(n6306), .Z(n6332) );
  XNOR U6608 ( .A(b[3]), .B(a[150]), .Z(n6347) );
  NANDN U6609 ( .A(n6347), .B(n10398), .Z(n6310) );
  NANDN U6610 ( .A(n6308), .B(n10399), .Z(n6309) );
  AND U6611 ( .A(n6310), .B(n6309), .Z(n6333) );
  XNOR U6612 ( .A(n6332), .B(n6333), .Z(n6334) );
  NANDN U6613 ( .A(n527), .B(a[152]), .Z(n6311) );
  XOR U6614 ( .A(n10434), .B(n6311), .Z(n6313) );
  NANDN U6615 ( .A(b[0]), .B(a[151]), .Z(n6312) );
  AND U6616 ( .A(n6313), .B(n6312), .Z(n6340) );
  XOR U6617 ( .A(b[5]), .B(a[148]), .Z(n6353) );
  NAND U6618 ( .A(n6353), .B(n10481), .Z(n6316) );
  NAND U6619 ( .A(n6314), .B(n10482), .Z(n6315) );
  NAND U6620 ( .A(n6316), .B(n6315), .Z(n6338) );
  NANDN U6621 ( .A(n529), .B(a[144]), .Z(n6339) );
  XNOR U6622 ( .A(n6338), .B(n6339), .Z(n6341) );
  XOR U6623 ( .A(n6340), .B(n6341), .Z(n6335) );
  XOR U6624 ( .A(n6334), .B(n6335), .Z(n6356) );
  XOR U6625 ( .A(n6357), .B(n6356), .Z(n6358) );
  XNOR U6626 ( .A(n6359), .B(n6358), .Z(n6328) );
  NAND U6627 ( .A(n6318), .B(n6317), .Z(n6322) );
  NAND U6628 ( .A(n6320), .B(n6319), .Z(n6321) );
  NAND U6629 ( .A(n6322), .B(n6321), .Z(n6329) );
  XNOR U6630 ( .A(n6328), .B(n6329), .Z(n6330) );
  XNOR U6631 ( .A(n6331), .B(n6330), .Z(n6362) );
  XNOR U6632 ( .A(n6362), .B(sreg[400]), .Z(n6364) );
  NAND U6633 ( .A(n6323), .B(sreg[399]), .Z(n6327) );
  OR U6634 ( .A(n6325), .B(n6324), .Z(n6326) );
  AND U6635 ( .A(n6327), .B(n6326), .Z(n6363) );
  XOR U6636 ( .A(n6364), .B(n6363), .Z(c[400]) );
  NANDN U6637 ( .A(n6333), .B(n6332), .Z(n6337) );
  NAND U6638 ( .A(n6335), .B(n6334), .Z(n6336) );
  NAND U6639 ( .A(n6337), .B(n6336), .Z(n6398) );
  NANDN U6640 ( .A(n6339), .B(n6338), .Z(n6343) );
  NAND U6641 ( .A(n6341), .B(n6340), .Z(n6342) );
  NAND U6642 ( .A(n6343), .B(n6342), .Z(n6396) );
  XNOR U6643 ( .A(b[7]), .B(a[147]), .Z(n6383) );
  NANDN U6644 ( .A(n6383), .B(n10545), .Z(n6346) );
  NANDN U6645 ( .A(n6344), .B(n10546), .Z(n6345) );
  NAND U6646 ( .A(n6346), .B(n6345), .Z(n6371) );
  XNOR U6647 ( .A(b[3]), .B(a[151]), .Z(n6386) );
  NANDN U6648 ( .A(n6386), .B(n10398), .Z(n6349) );
  NANDN U6649 ( .A(n6347), .B(n10399), .Z(n6348) );
  AND U6650 ( .A(n6349), .B(n6348), .Z(n6372) );
  XNOR U6651 ( .A(n6371), .B(n6372), .Z(n6373) );
  NANDN U6652 ( .A(n527), .B(a[153]), .Z(n6350) );
  XOR U6653 ( .A(n10434), .B(n6350), .Z(n6352) );
  NANDN U6654 ( .A(b[0]), .B(a[152]), .Z(n6351) );
  AND U6655 ( .A(n6352), .B(n6351), .Z(n6379) );
  XOR U6656 ( .A(b[5]), .B(a[149]), .Z(n6392) );
  NAND U6657 ( .A(n6392), .B(n10481), .Z(n6355) );
  NAND U6658 ( .A(n6353), .B(n10482), .Z(n6354) );
  NAND U6659 ( .A(n6355), .B(n6354), .Z(n6377) );
  NANDN U6660 ( .A(n529), .B(a[145]), .Z(n6378) );
  XNOR U6661 ( .A(n6377), .B(n6378), .Z(n6380) );
  XOR U6662 ( .A(n6379), .B(n6380), .Z(n6374) );
  XOR U6663 ( .A(n6373), .B(n6374), .Z(n6395) );
  XOR U6664 ( .A(n6396), .B(n6395), .Z(n6397) );
  XNOR U6665 ( .A(n6398), .B(n6397), .Z(n6367) );
  NAND U6666 ( .A(n6357), .B(n6356), .Z(n6361) );
  NAND U6667 ( .A(n6359), .B(n6358), .Z(n6360) );
  NAND U6668 ( .A(n6361), .B(n6360), .Z(n6368) );
  XNOR U6669 ( .A(n6367), .B(n6368), .Z(n6369) );
  XNOR U6670 ( .A(n6370), .B(n6369), .Z(n6401) );
  XNOR U6671 ( .A(n6401), .B(sreg[401]), .Z(n6403) );
  NAND U6672 ( .A(n6362), .B(sreg[400]), .Z(n6366) );
  OR U6673 ( .A(n6364), .B(n6363), .Z(n6365) );
  AND U6674 ( .A(n6366), .B(n6365), .Z(n6402) );
  XOR U6675 ( .A(n6403), .B(n6402), .Z(c[401]) );
  NANDN U6676 ( .A(n6372), .B(n6371), .Z(n6376) );
  NAND U6677 ( .A(n6374), .B(n6373), .Z(n6375) );
  NAND U6678 ( .A(n6376), .B(n6375), .Z(n6437) );
  NANDN U6679 ( .A(n6378), .B(n6377), .Z(n6382) );
  NAND U6680 ( .A(n6380), .B(n6379), .Z(n6381) );
  NAND U6681 ( .A(n6382), .B(n6381), .Z(n6435) );
  XNOR U6682 ( .A(b[7]), .B(a[148]), .Z(n6422) );
  NANDN U6683 ( .A(n6422), .B(n10545), .Z(n6385) );
  NANDN U6684 ( .A(n6383), .B(n10546), .Z(n6384) );
  NAND U6685 ( .A(n6385), .B(n6384), .Z(n6410) );
  XNOR U6686 ( .A(b[3]), .B(a[152]), .Z(n6425) );
  NANDN U6687 ( .A(n6425), .B(n10398), .Z(n6388) );
  NANDN U6688 ( .A(n6386), .B(n10399), .Z(n6387) );
  AND U6689 ( .A(n6388), .B(n6387), .Z(n6411) );
  XNOR U6690 ( .A(n6410), .B(n6411), .Z(n6412) );
  NANDN U6691 ( .A(n527), .B(a[154]), .Z(n6389) );
  XOR U6692 ( .A(n10434), .B(n6389), .Z(n6391) );
  NANDN U6693 ( .A(b[0]), .B(a[153]), .Z(n6390) );
  AND U6694 ( .A(n6391), .B(n6390), .Z(n6418) );
  XOR U6695 ( .A(b[5]), .B(a[150]), .Z(n6431) );
  NAND U6696 ( .A(n6431), .B(n10481), .Z(n6394) );
  NAND U6697 ( .A(n6392), .B(n10482), .Z(n6393) );
  NAND U6698 ( .A(n6394), .B(n6393), .Z(n6416) );
  NANDN U6699 ( .A(n529), .B(a[146]), .Z(n6417) );
  XNOR U6700 ( .A(n6416), .B(n6417), .Z(n6419) );
  XOR U6701 ( .A(n6418), .B(n6419), .Z(n6413) );
  XOR U6702 ( .A(n6412), .B(n6413), .Z(n6434) );
  XOR U6703 ( .A(n6435), .B(n6434), .Z(n6436) );
  XNOR U6704 ( .A(n6437), .B(n6436), .Z(n6406) );
  NAND U6705 ( .A(n6396), .B(n6395), .Z(n6400) );
  NAND U6706 ( .A(n6398), .B(n6397), .Z(n6399) );
  NAND U6707 ( .A(n6400), .B(n6399), .Z(n6407) );
  XNOR U6708 ( .A(n6406), .B(n6407), .Z(n6408) );
  XNOR U6709 ( .A(n6409), .B(n6408), .Z(n6440) );
  XNOR U6710 ( .A(n6440), .B(sreg[402]), .Z(n6442) );
  NAND U6711 ( .A(n6401), .B(sreg[401]), .Z(n6405) );
  OR U6712 ( .A(n6403), .B(n6402), .Z(n6404) );
  AND U6713 ( .A(n6405), .B(n6404), .Z(n6441) );
  XOR U6714 ( .A(n6442), .B(n6441), .Z(c[402]) );
  NANDN U6715 ( .A(n6411), .B(n6410), .Z(n6415) );
  NAND U6716 ( .A(n6413), .B(n6412), .Z(n6414) );
  NAND U6717 ( .A(n6415), .B(n6414), .Z(n6476) );
  NANDN U6718 ( .A(n6417), .B(n6416), .Z(n6421) );
  NAND U6719 ( .A(n6419), .B(n6418), .Z(n6420) );
  NAND U6720 ( .A(n6421), .B(n6420), .Z(n6474) );
  XNOR U6721 ( .A(b[7]), .B(a[149]), .Z(n6461) );
  NANDN U6722 ( .A(n6461), .B(n10545), .Z(n6424) );
  NANDN U6723 ( .A(n6422), .B(n10546), .Z(n6423) );
  NAND U6724 ( .A(n6424), .B(n6423), .Z(n6449) );
  XNOR U6725 ( .A(b[3]), .B(a[153]), .Z(n6464) );
  NANDN U6726 ( .A(n6464), .B(n10398), .Z(n6427) );
  NANDN U6727 ( .A(n6425), .B(n10399), .Z(n6426) );
  AND U6728 ( .A(n6427), .B(n6426), .Z(n6450) );
  XNOR U6729 ( .A(n6449), .B(n6450), .Z(n6451) );
  NANDN U6730 ( .A(n527), .B(a[155]), .Z(n6428) );
  XOR U6731 ( .A(n10434), .B(n6428), .Z(n6430) );
  NANDN U6732 ( .A(b[0]), .B(a[154]), .Z(n6429) );
  AND U6733 ( .A(n6430), .B(n6429), .Z(n6457) );
  XOR U6734 ( .A(b[5]), .B(a[151]), .Z(n6470) );
  NAND U6735 ( .A(n6470), .B(n10481), .Z(n6433) );
  NAND U6736 ( .A(n6431), .B(n10482), .Z(n6432) );
  NAND U6737 ( .A(n6433), .B(n6432), .Z(n6455) );
  NANDN U6738 ( .A(n529), .B(a[147]), .Z(n6456) );
  XNOR U6739 ( .A(n6455), .B(n6456), .Z(n6458) );
  XOR U6740 ( .A(n6457), .B(n6458), .Z(n6452) );
  XOR U6741 ( .A(n6451), .B(n6452), .Z(n6473) );
  XOR U6742 ( .A(n6474), .B(n6473), .Z(n6475) );
  XNOR U6743 ( .A(n6476), .B(n6475), .Z(n6445) );
  NAND U6744 ( .A(n6435), .B(n6434), .Z(n6439) );
  NAND U6745 ( .A(n6437), .B(n6436), .Z(n6438) );
  NAND U6746 ( .A(n6439), .B(n6438), .Z(n6446) );
  XNOR U6747 ( .A(n6445), .B(n6446), .Z(n6447) );
  XNOR U6748 ( .A(n6448), .B(n6447), .Z(n6479) );
  XNOR U6749 ( .A(n6479), .B(sreg[403]), .Z(n6481) );
  NAND U6750 ( .A(n6440), .B(sreg[402]), .Z(n6444) );
  OR U6751 ( .A(n6442), .B(n6441), .Z(n6443) );
  AND U6752 ( .A(n6444), .B(n6443), .Z(n6480) );
  XOR U6753 ( .A(n6481), .B(n6480), .Z(c[403]) );
  NANDN U6754 ( .A(n6450), .B(n6449), .Z(n6454) );
  NAND U6755 ( .A(n6452), .B(n6451), .Z(n6453) );
  NAND U6756 ( .A(n6454), .B(n6453), .Z(n6515) );
  NANDN U6757 ( .A(n6456), .B(n6455), .Z(n6460) );
  NAND U6758 ( .A(n6458), .B(n6457), .Z(n6459) );
  NAND U6759 ( .A(n6460), .B(n6459), .Z(n6513) );
  XNOR U6760 ( .A(b[7]), .B(a[150]), .Z(n6500) );
  NANDN U6761 ( .A(n6500), .B(n10545), .Z(n6463) );
  NANDN U6762 ( .A(n6461), .B(n10546), .Z(n6462) );
  NAND U6763 ( .A(n6463), .B(n6462), .Z(n6488) );
  XNOR U6764 ( .A(b[3]), .B(a[154]), .Z(n6503) );
  NANDN U6765 ( .A(n6503), .B(n10398), .Z(n6466) );
  NANDN U6766 ( .A(n6464), .B(n10399), .Z(n6465) );
  AND U6767 ( .A(n6466), .B(n6465), .Z(n6489) );
  XNOR U6768 ( .A(n6488), .B(n6489), .Z(n6490) );
  NANDN U6769 ( .A(n527), .B(a[156]), .Z(n6467) );
  XOR U6770 ( .A(n10434), .B(n6467), .Z(n6469) );
  NANDN U6771 ( .A(b[0]), .B(a[155]), .Z(n6468) );
  AND U6772 ( .A(n6469), .B(n6468), .Z(n6496) );
  XOR U6773 ( .A(b[5]), .B(a[152]), .Z(n6509) );
  NAND U6774 ( .A(n6509), .B(n10481), .Z(n6472) );
  NAND U6775 ( .A(n6470), .B(n10482), .Z(n6471) );
  NAND U6776 ( .A(n6472), .B(n6471), .Z(n6494) );
  NANDN U6777 ( .A(n529), .B(a[148]), .Z(n6495) );
  XNOR U6778 ( .A(n6494), .B(n6495), .Z(n6497) );
  XOR U6779 ( .A(n6496), .B(n6497), .Z(n6491) );
  XOR U6780 ( .A(n6490), .B(n6491), .Z(n6512) );
  XOR U6781 ( .A(n6513), .B(n6512), .Z(n6514) );
  XNOR U6782 ( .A(n6515), .B(n6514), .Z(n6484) );
  NAND U6783 ( .A(n6474), .B(n6473), .Z(n6478) );
  NAND U6784 ( .A(n6476), .B(n6475), .Z(n6477) );
  NAND U6785 ( .A(n6478), .B(n6477), .Z(n6485) );
  XNOR U6786 ( .A(n6484), .B(n6485), .Z(n6486) );
  XNOR U6787 ( .A(n6487), .B(n6486), .Z(n6518) );
  XNOR U6788 ( .A(n6518), .B(sreg[404]), .Z(n6520) );
  NAND U6789 ( .A(n6479), .B(sreg[403]), .Z(n6483) );
  OR U6790 ( .A(n6481), .B(n6480), .Z(n6482) );
  AND U6791 ( .A(n6483), .B(n6482), .Z(n6519) );
  XOR U6792 ( .A(n6520), .B(n6519), .Z(c[404]) );
  NANDN U6793 ( .A(n6489), .B(n6488), .Z(n6493) );
  NAND U6794 ( .A(n6491), .B(n6490), .Z(n6492) );
  NAND U6795 ( .A(n6493), .B(n6492), .Z(n6554) );
  NANDN U6796 ( .A(n6495), .B(n6494), .Z(n6499) );
  NAND U6797 ( .A(n6497), .B(n6496), .Z(n6498) );
  NAND U6798 ( .A(n6499), .B(n6498), .Z(n6552) );
  XNOR U6799 ( .A(b[7]), .B(a[151]), .Z(n6545) );
  NANDN U6800 ( .A(n6545), .B(n10545), .Z(n6502) );
  NANDN U6801 ( .A(n6500), .B(n10546), .Z(n6501) );
  NAND U6802 ( .A(n6502), .B(n6501), .Z(n6527) );
  XNOR U6803 ( .A(b[3]), .B(a[155]), .Z(n6548) );
  NANDN U6804 ( .A(n6548), .B(n10398), .Z(n6505) );
  NANDN U6805 ( .A(n6503), .B(n10399), .Z(n6504) );
  AND U6806 ( .A(n6505), .B(n6504), .Z(n6528) );
  XNOR U6807 ( .A(n6527), .B(n6528), .Z(n6529) );
  NANDN U6808 ( .A(n527), .B(a[157]), .Z(n6506) );
  XOR U6809 ( .A(n10434), .B(n6506), .Z(n6508) );
  NANDN U6810 ( .A(b[0]), .B(a[156]), .Z(n6507) );
  AND U6811 ( .A(n6508), .B(n6507), .Z(n6535) );
  XOR U6812 ( .A(b[5]), .B(a[153]), .Z(n6542) );
  NAND U6813 ( .A(n6542), .B(n10481), .Z(n6511) );
  NAND U6814 ( .A(n6509), .B(n10482), .Z(n6510) );
  NAND U6815 ( .A(n6511), .B(n6510), .Z(n6533) );
  NANDN U6816 ( .A(n529), .B(a[149]), .Z(n6534) );
  XNOR U6817 ( .A(n6533), .B(n6534), .Z(n6536) );
  XOR U6818 ( .A(n6535), .B(n6536), .Z(n6530) );
  XOR U6819 ( .A(n6529), .B(n6530), .Z(n6551) );
  XOR U6820 ( .A(n6552), .B(n6551), .Z(n6553) );
  XNOR U6821 ( .A(n6554), .B(n6553), .Z(n6523) );
  NAND U6822 ( .A(n6513), .B(n6512), .Z(n6517) );
  NAND U6823 ( .A(n6515), .B(n6514), .Z(n6516) );
  NAND U6824 ( .A(n6517), .B(n6516), .Z(n6524) );
  XNOR U6825 ( .A(n6523), .B(n6524), .Z(n6525) );
  XNOR U6826 ( .A(n6526), .B(n6525), .Z(n6557) );
  XNOR U6827 ( .A(n6557), .B(sreg[405]), .Z(n6559) );
  NAND U6828 ( .A(n6518), .B(sreg[404]), .Z(n6522) );
  OR U6829 ( .A(n6520), .B(n6519), .Z(n6521) );
  AND U6830 ( .A(n6522), .B(n6521), .Z(n6558) );
  XOR U6831 ( .A(n6559), .B(n6558), .Z(c[405]) );
  NANDN U6832 ( .A(n6528), .B(n6527), .Z(n6532) );
  NAND U6833 ( .A(n6530), .B(n6529), .Z(n6531) );
  NAND U6834 ( .A(n6532), .B(n6531), .Z(n6593) );
  NANDN U6835 ( .A(n6534), .B(n6533), .Z(n6538) );
  NAND U6836 ( .A(n6536), .B(n6535), .Z(n6537) );
  NAND U6837 ( .A(n6538), .B(n6537), .Z(n6591) );
  NANDN U6838 ( .A(n527), .B(a[158]), .Z(n6539) );
  XOR U6839 ( .A(n10434), .B(n6539), .Z(n6541) );
  NANDN U6840 ( .A(b[0]), .B(a[157]), .Z(n6540) );
  AND U6841 ( .A(n6541), .B(n6540), .Z(n6574) );
  XOR U6842 ( .A(b[5]), .B(a[154]), .Z(n6587) );
  NAND U6843 ( .A(n6587), .B(n10481), .Z(n6544) );
  NAND U6844 ( .A(n6542), .B(n10482), .Z(n6543) );
  NAND U6845 ( .A(n6544), .B(n6543), .Z(n6572) );
  NANDN U6846 ( .A(n529), .B(a[150]), .Z(n6573) );
  XNOR U6847 ( .A(n6572), .B(n6573), .Z(n6575) );
  XOR U6848 ( .A(n6574), .B(n6575), .Z(n6568) );
  XNOR U6849 ( .A(b[7]), .B(a[152]), .Z(n6578) );
  NANDN U6850 ( .A(n6578), .B(n10545), .Z(n6547) );
  NANDN U6851 ( .A(n6545), .B(n10546), .Z(n6546) );
  NAND U6852 ( .A(n6547), .B(n6546), .Z(n6566) );
  XNOR U6853 ( .A(b[3]), .B(a[156]), .Z(n6581) );
  NANDN U6854 ( .A(n6581), .B(n10398), .Z(n6550) );
  NANDN U6855 ( .A(n6548), .B(n10399), .Z(n6549) );
  AND U6856 ( .A(n6550), .B(n6549), .Z(n6567) );
  XNOR U6857 ( .A(n6566), .B(n6567), .Z(n6569) );
  XOR U6858 ( .A(n6568), .B(n6569), .Z(n6590) );
  XOR U6859 ( .A(n6591), .B(n6590), .Z(n6592) );
  XNOR U6860 ( .A(n6593), .B(n6592), .Z(n6562) );
  NAND U6861 ( .A(n6552), .B(n6551), .Z(n6556) );
  NAND U6862 ( .A(n6554), .B(n6553), .Z(n6555) );
  NAND U6863 ( .A(n6556), .B(n6555), .Z(n6563) );
  XNOR U6864 ( .A(n6562), .B(n6563), .Z(n6564) );
  XNOR U6865 ( .A(n6565), .B(n6564), .Z(n6596) );
  XNOR U6866 ( .A(n6596), .B(sreg[406]), .Z(n6598) );
  NAND U6867 ( .A(n6557), .B(sreg[405]), .Z(n6561) );
  OR U6868 ( .A(n6559), .B(n6558), .Z(n6560) );
  AND U6869 ( .A(n6561), .B(n6560), .Z(n6597) );
  XOR U6870 ( .A(n6598), .B(n6597), .Z(c[406]) );
  NANDN U6871 ( .A(n6567), .B(n6566), .Z(n6571) );
  NAND U6872 ( .A(n6569), .B(n6568), .Z(n6570) );
  NAND U6873 ( .A(n6571), .B(n6570), .Z(n6632) );
  NANDN U6874 ( .A(n6573), .B(n6572), .Z(n6577) );
  NAND U6875 ( .A(n6575), .B(n6574), .Z(n6576) );
  NAND U6876 ( .A(n6577), .B(n6576), .Z(n6630) );
  XNOR U6877 ( .A(b[7]), .B(a[153]), .Z(n6617) );
  NANDN U6878 ( .A(n6617), .B(n10545), .Z(n6580) );
  NANDN U6879 ( .A(n6578), .B(n10546), .Z(n6579) );
  NAND U6880 ( .A(n6580), .B(n6579), .Z(n6605) );
  XNOR U6881 ( .A(b[3]), .B(a[157]), .Z(n6620) );
  NANDN U6882 ( .A(n6620), .B(n10398), .Z(n6583) );
  NANDN U6883 ( .A(n6581), .B(n10399), .Z(n6582) );
  AND U6884 ( .A(n6583), .B(n6582), .Z(n6606) );
  XNOR U6885 ( .A(n6605), .B(n6606), .Z(n6607) );
  NANDN U6886 ( .A(n527), .B(a[159]), .Z(n6584) );
  XOR U6887 ( .A(n10434), .B(n6584), .Z(n6586) );
  NANDN U6888 ( .A(b[0]), .B(a[158]), .Z(n6585) );
  AND U6889 ( .A(n6586), .B(n6585), .Z(n6613) );
  XOR U6890 ( .A(b[5]), .B(a[155]), .Z(n6626) );
  NAND U6891 ( .A(n6626), .B(n10481), .Z(n6589) );
  NAND U6892 ( .A(n6587), .B(n10482), .Z(n6588) );
  NAND U6893 ( .A(n6589), .B(n6588), .Z(n6611) );
  NANDN U6894 ( .A(n529), .B(a[151]), .Z(n6612) );
  XNOR U6895 ( .A(n6611), .B(n6612), .Z(n6614) );
  XOR U6896 ( .A(n6613), .B(n6614), .Z(n6608) );
  XOR U6897 ( .A(n6607), .B(n6608), .Z(n6629) );
  XOR U6898 ( .A(n6630), .B(n6629), .Z(n6631) );
  XNOR U6899 ( .A(n6632), .B(n6631), .Z(n6601) );
  NAND U6900 ( .A(n6591), .B(n6590), .Z(n6595) );
  NAND U6901 ( .A(n6593), .B(n6592), .Z(n6594) );
  NAND U6902 ( .A(n6595), .B(n6594), .Z(n6602) );
  XNOR U6903 ( .A(n6601), .B(n6602), .Z(n6603) );
  XNOR U6904 ( .A(n6604), .B(n6603), .Z(n6635) );
  XNOR U6905 ( .A(n6635), .B(sreg[407]), .Z(n6637) );
  NAND U6906 ( .A(n6596), .B(sreg[406]), .Z(n6600) );
  OR U6907 ( .A(n6598), .B(n6597), .Z(n6599) );
  AND U6908 ( .A(n6600), .B(n6599), .Z(n6636) );
  XOR U6909 ( .A(n6637), .B(n6636), .Z(c[407]) );
  NANDN U6910 ( .A(n6606), .B(n6605), .Z(n6610) );
  NAND U6911 ( .A(n6608), .B(n6607), .Z(n6609) );
  NAND U6912 ( .A(n6610), .B(n6609), .Z(n6671) );
  NANDN U6913 ( .A(n6612), .B(n6611), .Z(n6616) );
  NAND U6914 ( .A(n6614), .B(n6613), .Z(n6615) );
  NAND U6915 ( .A(n6616), .B(n6615), .Z(n6669) );
  XNOR U6916 ( .A(b[7]), .B(a[154]), .Z(n6656) );
  NANDN U6917 ( .A(n6656), .B(n10545), .Z(n6619) );
  NANDN U6918 ( .A(n6617), .B(n10546), .Z(n6618) );
  NAND U6919 ( .A(n6619), .B(n6618), .Z(n6644) );
  XNOR U6920 ( .A(b[3]), .B(a[158]), .Z(n6659) );
  NANDN U6921 ( .A(n6659), .B(n10398), .Z(n6622) );
  NANDN U6922 ( .A(n6620), .B(n10399), .Z(n6621) );
  AND U6923 ( .A(n6622), .B(n6621), .Z(n6645) );
  XNOR U6924 ( .A(n6644), .B(n6645), .Z(n6646) );
  NANDN U6925 ( .A(n527), .B(a[160]), .Z(n6623) );
  XOR U6926 ( .A(n10434), .B(n6623), .Z(n6625) );
  NANDN U6927 ( .A(b[0]), .B(a[159]), .Z(n6624) );
  AND U6928 ( .A(n6625), .B(n6624), .Z(n6652) );
  XOR U6929 ( .A(b[5]), .B(a[156]), .Z(n6665) );
  NAND U6930 ( .A(n6665), .B(n10481), .Z(n6628) );
  NAND U6931 ( .A(n6626), .B(n10482), .Z(n6627) );
  NAND U6932 ( .A(n6628), .B(n6627), .Z(n6650) );
  NANDN U6933 ( .A(n529), .B(a[152]), .Z(n6651) );
  XNOR U6934 ( .A(n6650), .B(n6651), .Z(n6653) );
  XOR U6935 ( .A(n6652), .B(n6653), .Z(n6647) );
  XOR U6936 ( .A(n6646), .B(n6647), .Z(n6668) );
  XOR U6937 ( .A(n6669), .B(n6668), .Z(n6670) );
  XNOR U6938 ( .A(n6671), .B(n6670), .Z(n6640) );
  NAND U6939 ( .A(n6630), .B(n6629), .Z(n6634) );
  NAND U6940 ( .A(n6632), .B(n6631), .Z(n6633) );
  NAND U6941 ( .A(n6634), .B(n6633), .Z(n6641) );
  XNOR U6942 ( .A(n6640), .B(n6641), .Z(n6642) );
  XNOR U6943 ( .A(n6643), .B(n6642), .Z(n6674) );
  XNOR U6944 ( .A(n6674), .B(sreg[408]), .Z(n6676) );
  NAND U6945 ( .A(n6635), .B(sreg[407]), .Z(n6639) );
  OR U6946 ( .A(n6637), .B(n6636), .Z(n6638) );
  AND U6947 ( .A(n6639), .B(n6638), .Z(n6675) );
  XOR U6948 ( .A(n6676), .B(n6675), .Z(c[408]) );
  NANDN U6949 ( .A(n6645), .B(n6644), .Z(n6649) );
  NAND U6950 ( .A(n6647), .B(n6646), .Z(n6648) );
  NAND U6951 ( .A(n6649), .B(n6648), .Z(n6710) );
  NANDN U6952 ( .A(n6651), .B(n6650), .Z(n6655) );
  NAND U6953 ( .A(n6653), .B(n6652), .Z(n6654) );
  NAND U6954 ( .A(n6655), .B(n6654), .Z(n6708) );
  XNOR U6955 ( .A(b[7]), .B(a[155]), .Z(n6695) );
  NANDN U6956 ( .A(n6695), .B(n10545), .Z(n6658) );
  NANDN U6957 ( .A(n6656), .B(n10546), .Z(n6657) );
  NAND U6958 ( .A(n6658), .B(n6657), .Z(n6683) );
  XNOR U6959 ( .A(b[3]), .B(a[159]), .Z(n6698) );
  NANDN U6960 ( .A(n6698), .B(n10398), .Z(n6661) );
  NANDN U6961 ( .A(n6659), .B(n10399), .Z(n6660) );
  AND U6962 ( .A(n6661), .B(n6660), .Z(n6684) );
  XNOR U6963 ( .A(n6683), .B(n6684), .Z(n6685) );
  NANDN U6964 ( .A(n527), .B(a[161]), .Z(n6662) );
  XOR U6965 ( .A(n10434), .B(n6662), .Z(n6664) );
  NANDN U6966 ( .A(b[0]), .B(a[160]), .Z(n6663) );
  AND U6967 ( .A(n6664), .B(n6663), .Z(n6691) );
  XOR U6968 ( .A(b[5]), .B(a[157]), .Z(n6704) );
  NAND U6969 ( .A(n6704), .B(n10481), .Z(n6667) );
  NAND U6970 ( .A(n6665), .B(n10482), .Z(n6666) );
  NAND U6971 ( .A(n6667), .B(n6666), .Z(n6689) );
  NANDN U6972 ( .A(n529), .B(a[153]), .Z(n6690) );
  XNOR U6973 ( .A(n6689), .B(n6690), .Z(n6692) );
  XOR U6974 ( .A(n6691), .B(n6692), .Z(n6686) );
  XOR U6975 ( .A(n6685), .B(n6686), .Z(n6707) );
  XOR U6976 ( .A(n6708), .B(n6707), .Z(n6709) );
  XNOR U6977 ( .A(n6710), .B(n6709), .Z(n6679) );
  NAND U6978 ( .A(n6669), .B(n6668), .Z(n6673) );
  NAND U6979 ( .A(n6671), .B(n6670), .Z(n6672) );
  NAND U6980 ( .A(n6673), .B(n6672), .Z(n6680) );
  XNOR U6981 ( .A(n6679), .B(n6680), .Z(n6681) );
  XNOR U6982 ( .A(n6682), .B(n6681), .Z(n6713) );
  XNOR U6983 ( .A(n6713), .B(sreg[409]), .Z(n6715) );
  NAND U6984 ( .A(n6674), .B(sreg[408]), .Z(n6678) );
  OR U6985 ( .A(n6676), .B(n6675), .Z(n6677) );
  AND U6986 ( .A(n6678), .B(n6677), .Z(n6714) );
  XOR U6987 ( .A(n6715), .B(n6714), .Z(c[409]) );
  NANDN U6988 ( .A(n6684), .B(n6683), .Z(n6688) );
  NAND U6989 ( .A(n6686), .B(n6685), .Z(n6687) );
  NAND U6990 ( .A(n6688), .B(n6687), .Z(n6749) );
  NANDN U6991 ( .A(n6690), .B(n6689), .Z(n6694) );
  NAND U6992 ( .A(n6692), .B(n6691), .Z(n6693) );
  NAND U6993 ( .A(n6694), .B(n6693), .Z(n6747) );
  XNOR U6994 ( .A(b[7]), .B(a[156]), .Z(n6734) );
  NANDN U6995 ( .A(n6734), .B(n10545), .Z(n6697) );
  NANDN U6996 ( .A(n6695), .B(n10546), .Z(n6696) );
  NAND U6997 ( .A(n6697), .B(n6696), .Z(n6722) );
  XNOR U6998 ( .A(b[3]), .B(a[160]), .Z(n6737) );
  NANDN U6999 ( .A(n6737), .B(n10398), .Z(n6700) );
  NANDN U7000 ( .A(n6698), .B(n10399), .Z(n6699) );
  AND U7001 ( .A(n6700), .B(n6699), .Z(n6723) );
  XNOR U7002 ( .A(n6722), .B(n6723), .Z(n6724) );
  NANDN U7003 ( .A(n527), .B(a[162]), .Z(n6701) );
  XOR U7004 ( .A(n10434), .B(n6701), .Z(n6703) );
  NANDN U7005 ( .A(b[0]), .B(a[161]), .Z(n6702) );
  AND U7006 ( .A(n6703), .B(n6702), .Z(n6730) );
  XOR U7007 ( .A(b[5]), .B(a[158]), .Z(n6743) );
  NAND U7008 ( .A(n6743), .B(n10481), .Z(n6706) );
  NAND U7009 ( .A(n6704), .B(n10482), .Z(n6705) );
  NAND U7010 ( .A(n6706), .B(n6705), .Z(n6728) );
  NANDN U7011 ( .A(n529), .B(a[154]), .Z(n6729) );
  XNOR U7012 ( .A(n6728), .B(n6729), .Z(n6731) );
  XOR U7013 ( .A(n6730), .B(n6731), .Z(n6725) );
  XOR U7014 ( .A(n6724), .B(n6725), .Z(n6746) );
  XOR U7015 ( .A(n6747), .B(n6746), .Z(n6748) );
  XNOR U7016 ( .A(n6749), .B(n6748), .Z(n6718) );
  NAND U7017 ( .A(n6708), .B(n6707), .Z(n6712) );
  NAND U7018 ( .A(n6710), .B(n6709), .Z(n6711) );
  NAND U7019 ( .A(n6712), .B(n6711), .Z(n6719) );
  XNOR U7020 ( .A(n6718), .B(n6719), .Z(n6720) );
  XNOR U7021 ( .A(n6721), .B(n6720), .Z(n6752) );
  XNOR U7022 ( .A(n6752), .B(sreg[410]), .Z(n6754) );
  NAND U7023 ( .A(n6713), .B(sreg[409]), .Z(n6717) );
  OR U7024 ( .A(n6715), .B(n6714), .Z(n6716) );
  AND U7025 ( .A(n6717), .B(n6716), .Z(n6753) );
  XOR U7026 ( .A(n6754), .B(n6753), .Z(c[410]) );
  NANDN U7027 ( .A(n6723), .B(n6722), .Z(n6727) );
  NAND U7028 ( .A(n6725), .B(n6724), .Z(n6726) );
  NAND U7029 ( .A(n6727), .B(n6726), .Z(n6788) );
  NANDN U7030 ( .A(n6729), .B(n6728), .Z(n6733) );
  NAND U7031 ( .A(n6731), .B(n6730), .Z(n6732) );
  NAND U7032 ( .A(n6733), .B(n6732), .Z(n6786) );
  XNOR U7033 ( .A(b[7]), .B(a[157]), .Z(n6773) );
  NANDN U7034 ( .A(n6773), .B(n10545), .Z(n6736) );
  NANDN U7035 ( .A(n6734), .B(n10546), .Z(n6735) );
  NAND U7036 ( .A(n6736), .B(n6735), .Z(n6761) );
  XNOR U7037 ( .A(b[3]), .B(a[161]), .Z(n6776) );
  NANDN U7038 ( .A(n6776), .B(n10398), .Z(n6739) );
  NANDN U7039 ( .A(n6737), .B(n10399), .Z(n6738) );
  AND U7040 ( .A(n6739), .B(n6738), .Z(n6762) );
  XNOR U7041 ( .A(n6761), .B(n6762), .Z(n6763) );
  NANDN U7042 ( .A(n527), .B(a[163]), .Z(n6740) );
  XOR U7043 ( .A(n10434), .B(n6740), .Z(n6742) );
  NANDN U7044 ( .A(b[0]), .B(a[162]), .Z(n6741) );
  AND U7045 ( .A(n6742), .B(n6741), .Z(n6769) );
  XOR U7046 ( .A(b[5]), .B(a[159]), .Z(n6782) );
  NAND U7047 ( .A(n6782), .B(n10481), .Z(n6745) );
  NAND U7048 ( .A(n6743), .B(n10482), .Z(n6744) );
  NAND U7049 ( .A(n6745), .B(n6744), .Z(n6767) );
  NANDN U7050 ( .A(n529), .B(a[155]), .Z(n6768) );
  XNOR U7051 ( .A(n6767), .B(n6768), .Z(n6770) );
  XOR U7052 ( .A(n6769), .B(n6770), .Z(n6764) );
  XOR U7053 ( .A(n6763), .B(n6764), .Z(n6785) );
  XOR U7054 ( .A(n6786), .B(n6785), .Z(n6787) );
  XNOR U7055 ( .A(n6788), .B(n6787), .Z(n6757) );
  NAND U7056 ( .A(n6747), .B(n6746), .Z(n6751) );
  NAND U7057 ( .A(n6749), .B(n6748), .Z(n6750) );
  NAND U7058 ( .A(n6751), .B(n6750), .Z(n6758) );
  XNOR U7059 ( .A(n6757), .B(n6758), .Z(n6759) );
  XNOR U7060 ( .A(n6760), .B(n6759), .Z(n6791) );
  XNOR U7061 ( .A(n6791), .B(sreg[411]), .Z(n6793) );
  NAND U7062 ( .A(n6752), .B(sreg[410]), .Z(n6756) );
  OR U7063 ( .A(n6754), .B(n6753), .Z(n6755) );
  AND U7064 ( .A(n6756), .B(n6755), .Z(n6792) );
  XOR U7065 ( .A(n6793), .B(n6792), .Z(c[411]) );
  NANDN U7066 ( .A(n6762), .B(n6761), .Z(n6766) );
  NAND U7067 ( .A(n6764), .B(n6763), .Z(n6765) );
  NAND U7068 ( .A(n6766), .B(n6765), .Z(n6827) );
  NANDN U7069 ( .A(n6768), .B(n6767), .Z(n6772) );
  NAND U7070 ( .A(n6770), .B(n6769), .Z(n6771) );
  NAND U7071 ( .A(n6772), .B(n6771), .Z(n6825) );
  XNOR U7072 ( .A(b[7]), .B(a[158]), .Z(n6818) );
  NANDN U7073 ( .A(n6818), .B(n10545), .Z(n6775) );
  NANDN U7074 ( .A(n6773), .B(n10546), .Z(n6774) );
  NAND U7075 ( .A(n6775), .B(n6774), .Z(n6800) );
  XNOR U7076 ( .A(b[3]), .B(a[162]), .Z(n6821) );
  NANDN U7077 ( .A(n6821), .B(n10398), .Z(n6778) );
  NANDN U7078 ( .A(n6776), .B(n10399), .Z(n6777) );
  AND U7079 ( .A(n6778), .B(n6777), .Z(n6801) );
  XNOR U7080 ( .A(n6800), .B(n6801), .Z(n6802) );
  NANDN U7081 ( .A(n527), .B(a[164]), .Z(n6779) );
  XOR U7082 ( .A(n10434), .B(n6779), .Z(n6781) );
  NANDN U7083 ( .A(b[0]), .B(a[163]), .Z(n6780) );
  AND U7084 ( .A(n6781), .B(n6780), .Z(n6808) );
  XOR U7085 ( .A(b[5]), .B(a[160]), .Z(n6815) );
  NAND U7086 ( .A(n6815), .B(n10481), .Z(n6784) );
  NAND U7087 ( .A(n6782), .B(n10482), .Z(n6783) );
  NAND U7088 ( .A(n6784), .B(n6783), .Z(n6806) );
  NANDN U7089 ( .A(n529), .B(a[156]), .Z(n6807) );
  XNOR U7090 ( .A(n6806), .B(n6807), .Z(n6809) );
  XOR U7091 ( .A(n6808), .B(n6809), .Z(n6803) );
  XOR U7092 ( .A(n6802), .B(n6803), .Z(n6824) );
  XOR U7093 ( .A(n6825), .B(n6824), .Z(n6826) );
  XNOR U7094 ( .A(n6827), .B(n6826), .Z(n6796) );
  NAND U7095 ( .A(n6786), .B(n6785), .Z(n6790) );
  NAND U7096 ( .A(n6788), .B(n6787), .Z(n6789) );
  NAND U7097 ( .A(n6790), .B(n6789), .Z(n6797) );
  XNOR U7098 ( .A(n6796), .B(n6797), .Z(n6798) );
  XNOR U7099 ( .A(n6799), .B(n6798), .Z(n6830) );
  XNOR U7100 ( .A(n6830), .B(sreg[412]), .Z(n6832) );
  NAND U7101 ( .A(n6791), .B(sreg[411]), .Z(n6795) );
  OR U7102 ( .A(n6793), .B(n6792), .Z(n6794) );
  AND U7103 ( .A(n6795), .B(n6794), .Z(n6831) );
  XOR U7104 ( .A(n6832), .B(n6831), .Z(c[412]) );
  NANDN U7105 ( .A(n6801), .B(n6800), .Z(n6805) );
  NAND U7106 ( .A(n6803), .B(n6802), .Z(n6804) );
  NAND U7107 ( .A(n6805), .B(n6804), .Z(n6866) );
  NANDN U7108 ( .A(n6807), .B(n6806), .Z(n6811) );
  NAND U7109 ( .A(n6809), .B(n6808), .Z(n6810) );
  NAND U7110 ( .A(n6811), .B(n6810), .Z(n6864) );
  NANDN U7111 ( .A(n527), .B(a[165]), .Z(n6812) );
  XOR U7112 ( .A(n10434), .B(n6812), .Z(n6814) );
  NANDN U7113 ( .A(b[0]), .B(a[164]), .Z(n6813) );
  AND U7114 ( .A(n6814), .B(n6813), .Z(n6847) );
  XOR U7115 ( .A(b[5]), .B(a[161]), .Z(n6860) );
  NAND U7116 ( .A(n6860), .B(n10481), .Z(n6817) );
  NAND U7117 ( .A(n6815), .B(n10482), .Z(n6816) );
  NAND U7118 ( .A(n6817), .B(n6816), .Z(n6845) );
  NANDN U7119 ( .A(n529), .B(a[157]), .Z(n6846) );
  XNOR U7120 ( .A(n6845), .B(n6846), .Z(n6848) );
  XOR U7121 ( .A(n6847), .B(n6848), .Z(n6841) );
  XNOR U7122 ( .A(b[7]), .B(a[159]), .Z(n6851) );
  NANDN U7123 ( .A(n6851), .B(n10545), .Z(n6820) );
  NANDN U7124 ( .A(n6818), .B(n10546), .Z(n6819) );
  NAND U7125 ( .A(n6820), .B(n6819), .Z(n6839) );
  XNOR U7126 ( .A(b[3]), .B(a[163]), .Z(n6854) );
  NANDN U7127 ( .A(n6854), .B(n10398), .Z(n6823) );
  NANDN U7128 ( .A(n6821), .B(n10399), .Z(n6822) );
  AND U7129 ( .A(n6823), .B(n6822), .Z(n6840) );
  XNOR U7130 ( .A(n6839), .B(n6840), .Z(n6842) );
  XOR U7131 ( .A(n6841), .B(n6842), .Z(n6863) );
  XOR U7132 ( .A(n6864), .B(n6863), .Z(n6865) );
  XNOR U7133 ( .A(n6866), .B(n6865), .Z(n6835) );
  NAND U7134 ( .A(n6825), .B(n6824), .Z(n6829) );
  NAND U7135 ( .A(n6827), .B(n6826), .Z(n6828) );
  NAND U7136 ( .A(n6829), .B(n6828), .Z(n6836) );
  XNOR U7137 ( .A(n6835), .B(n6836), .Z(n6837) );
  XNOR U7138 ( .A(n6838), .B(n6837), .Z(n6869) );
  XNOR U7139 ( .A(n6869), .B(sreg[413]), .Z(n6871) );
  NAND U7140 ( .A(n6830), .B(sreg[412]), .Z(n6834) );
  OR U7141 ( .A(n6832), .B(n6831), .Z(n6833) );
  AND U7142 ( .A(n6834), .B(n6833), .Z(n6870) );
  XOR U7143 ( .A(n6871), .B(n6870), .Z(c[413]) );
  NANDN U7144 ( .A(n6840), .B(n6839), .Z(n6844) );
  NAND U7145 ( .A(n6842), .B(n6841), .Z(n6843) );
  NAND U7146 ( .A(n6844), .B(n6843), .Z(n6905) );
  NANDN U7147 ( .A(n6846), .B(n6845), .Z(n6850) );
  NAND U7148 ( .A(n6848), .B(n6847), .Z(n6849) );
  NAND U7149 ( .A(n6850), .B(n6849), .Z(n6903) );
  XNOR U7150 ( .A(b[7]), .B(a[160]), .Z(n6890) );
  NANDN U7151 ( .A(n6890), .B(n10545), .Z(n6853) );
  NANDN U7152 ( .A(n6851), .B(n10546), .Z(n6852) );
  NAND U7153 ( .A(n6853), .B(n6852), .Z(n6878) );
  XNOR U7154 ( .A(b[3]), .B(a[164]), .Z(n6893) );
  NANDN U7155 ( .A(n6893), .B(n10398), .Z(n6856) );
  NANDN U7156 ( .A(n6854), .B(n10399), .Z(n6855) );
  AND U7157 ( .A(n6856), .B(n6855), .Z(n6879) );
  XNOR U7158 ( .A(n6878), .B(n6879), .Z(n6880) );
  NANDN U7159 ( .A(n527), .B(a[166]), .Z(n6857) );
  XOR U7160 ( .A(n10434), .B(n6857), .Z(n6859) );
  NANDN U7161 ( .A(b[0]), .B(a[165]), .Z(n6858) );
  AND U7162 ( .A(n6859), .B(n6858), .Z(n6886) );
  XOR U7163 ( .A(b[5]), .B(a[162]), .Z(n6899) );
  NAND U7164 ( .A(n6899), .B(n10481), .Z(n6862) );
  NAND U7165 ( .A(n6860), .B(n10482), .Z(n6861) );
  NAND U7166 ( .A(n6862), .B(n6861), .Z(n6884) );
  NANDN U7167 ( .A(n529), .B(a[158]), .Z(n6885) );
  XNOR U7168 ( .A(n6884), .B(n6885), .Z(n6887) );
  XOR U7169 ( .A(n6886), .B(n6887), .Z(n6881) );
  XOR U7170 ( .A(n6880), .B(n6881), .Z(n6902) );
  XOR U7171 ( .A(n6903), .B(n6902), .Z(n6904) );
  XNOR U7172 ( .A(n6905), .B(n6904), .Z(n6874) );
  NAND U7173 ( .A(n6864), .B(n6863), .Z(n6868) );
  NAND U7174 ( .A(n6866), .B(n6865), .Z(n6867) );
  NAND U7175 ( .A(n6868), .B(n6867), .Z(n6875) );
  XNOR U7176 ( .A(n6874), .B(n6875), .Z(n6876) );
  XNOR U7177 ( .A(n6877), .B(n6876), .Z(n6908) );
  XNOR U7178 ( .A(n6908), .B(sreg[414]), .Z(n6910) );
  NAND U7179 ( .A(n6869), .B(sreg[413]), .Z(n6873) );
  OR U7180 ( .A(n6871), .B(n6870), .Z(n6872) );
  AND U7181 ( .A(n6873), .B(n6872), .Z(n6909) );
  XOR U7182 ( .A(n6910), .B(n6909), .Z(c[414]) );
  NANDN U7183 ( .A(n6879), .B(n6878), .Z(n6883) );
  NAND U7184 ( .A(n6881), .B(n6880), .Z(n6882) );
  NAND U7185 ( .A(n6883), .B(n6882), .Z(n6944) );
  NANDN U7186 ( .A(n6885), .B(n6884), .Z(n6889) );
  NAND U7187 ( .A(n6887), .B(n6886), .Z(n6888) );
  NAND U7188 ( .A(n6889), .B(n6888), .Z(n6942) );
  XNOR U7189 ( .A(b[7]), .B(a[161]), .Z(n6929) );
  NANDN U7190 ( .A(n6929), .B(n10545), .Z(n6892) );
  NANDN U7191 ( .A(n6890), .B(n10546), .Z(n6891) );
  NAND U7192 ( .A(n6892), .B(n6891), .Z(n6917) );
  XNOR U7193 ( .A(b[3]), .B(a[165]), .Z(n6932) );
  NANDN U7194 ( .A(n6932), .B(n10398), .Z(n6895) );
  NANDN U7195 ( .A(n6893), .B(n10399), .Z(n6894) );
  AND U7196 ( .A(n6895), .B(n6894), .Z(n6918) );
  XNOR U7197 ( .A(n6917), .B(n6918), .Z(n6919) );
  NANDN U7198 ( .A(n527), .B(a[167]), .Z(n6896) );
  XOR U7199 ( .A(n10434), .B(n6896), .Z(n6898) );
  NANDN U7200 ( .A(b[0]), .B(a[166]), .Z(n6897) );
  AND U7201 ( .A(n6898), .B(n6897), .Z(n6925) );
  XOR U7202 ( .A(b[5]), .B(a[163]), .Z(n6938) );
  NAND U7203 ( .A(n6938), .B(n10481), .Z(n6901) );
  NAND U7204 ( .A(n6899), .B(n10482), .Z(n6900) );
  NAND U7205 ( .A(n6901), .B(n6900), .Z(n6923) );
  NANDN U7206 ( .A(n529), .B(a[159]), .Z(n6924) );
  XNOR U7207 ( .A(n6923), .B(n6924), .Z(n6926) );
  XOR U7208 ( .A(n6925), .B(n6926), .Z(n6920) );
  XOR U7209 ( .A(n6919), .B(n6920), .Z(n6941) );
  XOR U7210 ( .A(n6942), .B(n6941), .Z(n6943) );
  XNOR U7211 ( .A(n6944), .B(n6943), .Z(n6913) );
  NAND U7212 ( .A(n6903), .B(n6902), .Z(n6907) );
  NAND U7213 ( .A(n6905), .B(n6904), .Z(n6906) );
  NAND U7214 ( .A(n6907), .B(n6906), .Z(n6914) );
  XNOR U7215 ( .A(n6913), .B(n6914), .Z(n6915) );
  XNOR U7216 ( .A(n6916), .B(n6915), .Z(n6947) );
  XNOR U7217 ( .A(n6947), .B(sreg[415]), .Z(n6949) );
  NAND U7218 ( .A(n6908), .B(sreg[414]), .Z(n6912) );
  OR U7219 ( .A(n6910), .B(n6909), .Z(n6911) );
  AND U7220 ( .A(n6912), .B(n6911), .Z(n6948) );
  XOR U7221 ( .A(n6949), .B(n6948), .Z(c[415]) );
  NANDN U7222 ( .A(n6918), .B(n6917), .Z(n6922) );
  NAND U7223 ( .A(n6920), .B(n6919), .Z(n6921) );
  NAND U7224 ( .A(n6922), .B(n6921), .Z(n6983) );
  NANDN U7225 ( .A(n6924), .B(n6923), .Z(n6928) );
  NAND U7226 ( .A(n6926), .B(n6925), .Z(n6927) );
  NAND U7227 ( .A(n6928), .B(n6927), .Z(n6981) );
  XNOR U7228 ( .A(b[7]), .B(a[162]), .Z(n6968) );
  NANDN U7229 ( .A(n6968), .B(n10545), .Z(n6931) );
  NANDN U7230 ( .A(n6929), .B(n10546), .Z(n6930) );
  NAND U7231 ( .A(n6931), .B(n6930), .Z(n6956) );
  XNOR U7232 ( .A(b[3]), .B(a[166]), .Z(n6971) );
  NANDN U7233 ( .A(n6971), .B(n10398), .Z(n6934) );
  NANDN U7234 ( .A(n6932), .B(n10399), .Z(n6933) );
  AND U7235 ( .A(n6934), .B(n6933), .Z(n6957) );
  XNOR U7236 ( .A(n6956), .B(n6957), .Z(n6958) );
  NANDN U7237 ( .A(n527), .B(a[168]), .Z(n6935) );
  XOR U7238 ( .A(n10434), .B(n6935), .Z(n6937) );
  NANDN U7239 ( .A(b[0]), .B(a[167]), .Z(n6936) );
  AND U7240 ( .A(n6937), .B(n6936), .Z(n6964) );
  XOR U7241 ( .A(b[5]), .B(a[164]), .Z(n6977) );
  NAND U7242 ( .A(n6977), .B(n10481), .Z(n6940) );
  NAND U7243 ( .A(n6938), .B(n10482), .Z(n6939) );
  NAND U7244 ( .A(n6940), .B(n6939), .Z(n6962) );
  NANDN U7245 ( .A(n529), .B(a[160]), .Z(n6963) );
  XNOR U7246 ( .A(n6962), .B(n6963), .Z(n6965) );
  XOR U7247 ( .A(n6964), .B(n6965), .Z(n6959) );
  XOR U7248 ( .A(n6958), .B(n6959), .Z(n6980) );
  XOR U7249 ( .A(n6981), .B(n6980), .Z(n6982) );
  XNOR U7250 ( .A(n6983), .B(n6982), .Z(n6952) );
  NAND U7251 ( .A(n6942), .B(n6941), .Z(n6946) );
  NAND U7252 ( .A(n6944), .B(n6943), .Z(n6945) );
  NAND U7253 ( .A(n6946), .B(n6945), .Z(n6953) );
  XNOR U7254 ( .A(n6952), .B(n6953), .Z(n6954) );
  XNOR U7255 ( .A(n6955), .B(n6954), .Z(n6986) );
  XNOR U7256 ( .A(n6986), .B(sreg[416]), .Z(n6988) );
  NAND U7257 ( .A(n6947), .B(sreg[415]), .Z(n6951) );
  OR U7258 ( .A(n6949), .B(n6948), .Z(n6950) );
  AND U7259 ( .A(n6951), .B(n6950), .Z(n6987) );
  XOR U7260 ( .A(n6988), .B(n6987), .Z(c[416]) );
  NANDN U7261 ( .A(n6957), .B(n6956), .Z(n6961) );
  NAND U7262 ( .A(n6959), .B(n6958), .Z(n6960) );
  NAND U7263 ( .A(n6961), .B(n6960), .Z(n7022) );
  NANDN U7264 ( .A(n6963), .B(n6962), .Z(n6967) );
  NAND U7265 ( .A(n6965), .B(n6964), .Z(n6966) );
  NAND U7266 ( .A(n6967), .B(n6966), .Z(n7020) );
  XNOR U7267 ( .A(b[7]), .B(a[163]), .Z(n7007) );
  NANDN U7268 ( .A(n7007), .B(n10545), .Z(n6970) );
  NANDN U7269 ( .A(n6968), .B(n10546), .Z(n6969) );
  NAND U7270 ( .A(n6970), .B(n6969), .Z(n6995) );
  XNOR U7271 ( .A(b[3]), .B(a[167]), .Z(n7010) );
  NANDN U7272 ( .A(n7010), .B(n10398), .Z(n6973) );
  NANDN U7273 ( .A(n6971), .B(n10399), .Z(n6972) );
  AND U7274 ( .A(n6973), .B(n6972), .Z(n6996) );
  XNOR U7275 ( .A(n6995), .B(n6996), .Z(n6997) );
  NANDN U7276 ( .A(n527), .B(a[169]), .Z(n6974) );
  XOR U7277 ( .A(n10434), .B(n6974), .Z(n6976) );
  NANDN U7278 ( .A(b[0]), .B(a[168]), .Z(n6975) );
  AND U7279 ( .A(n6976), .B(n6975), .Z(n7003) );
  XOR U7280 ( .A(b[5]), .B(a[165]), .Z(n7016) );
  NAND U7281 ( .A(n7016), .B(n10481), .Z(n6979) );
  NAND U7282 ( .A(n6977), .B(n10482), .Z(n6978) );
  NAND U7283 ( .A(n6979), .B(n6978), .Z(n7001) );
  NANDN U7284 ( .A(n529), .B(a[161]), .Z(n7002) );
  XNOR U7285 ( .A(n7001), .B(n7002), .Z(n7004) );
  XOR U7286 ( .A(n7003), .B(n7004), .Z(n6998) );
  XOR U7287 ( .A(n6997), .B(n6998), .Z(n7019) );
  XOR U7288 ( .A(n7020), .B(n7019), .Z(n7021) );
  XNOR U7289 ( .A(n7022), .B(n7021), .Z(n6991) );
  NAND U7290 ( .A(n6981), .B(n6980), .Z(n6985) );
  NAND U7291 ( .A(n6983), .B(n6982), .Z(n6984) );
  NAND U7292 ( .A(n6985), .B(n6984), .Z(n6992) );
  XNOR U7293 ( .A(n6991), .B(n6992), .Z(n6993) );
  XNOR U7294 ( .A(n6994), .B(n6993), .Z(n7025) );
  XNOR U7295 ( .A(n7025), .B(sreg[417]), .Z(n7027) );
  NAND U7296 ( .A(n6986), .B(sreg[416]), .Z(n6990) );
  OR U7297 ( .A(n6988), .B(n6987), .Z(n6989) );
  AND U7298 ( .A(n6990), .B(n6989), .Z(n7026) );
  XOR U7299 ( .A(n7027), .B(n7026), .Z(c[417]) );
  NANDN U7300 ( .A(n6996), .B(n6995), .Z(n7000) );
  NAND U7301 ( .A(n6998), .B(n6997), .Z(n6999) );
  NAND U7302 ( .A(n7000), .B(n6999), .Z(n7061) );
  NANDN U7303 ( .A(n7002), .B(n7001), .Z(n7006) );
  NAND U7304 ( .A(n7004), .B(n7003), .Z(n7005) );
  NAND U7305 ( .A(n7006), .B(n7005), .Z(n7059) );
  XNOR U7306 ( .A(b[7]), .B(a[164]), .Z(n7052) );
  NANDN U7307 ( .A(n7052), .B(n10545), .Z(n7009) );
  NANDN U7308 ( .A(n7007), .B(n10546), .Z(n7008) );
  NAND U7309 ( .A(n7009), .B(n7008), .Z(n7034) );
  XNOR U7310 ( .A(b[3]), .B(a[168]), .Z(n7055) );
  NANDN U7311 ( .A(n7055), .B(n10398), .Z(n7012) );
  NANDN U7312 ( .A(n7010), .B(n10399), .Z(n7011) );
  AND U7313 ( .A(n7012), .B(n7011), .Z(n7035) );
  XNOR U7314 ( .A(n7034), .B(n7035), .Z(n7036) );
  NANDN U7315 ( .A(n527), .B(a[170]), .Z(n7013) );
  XOR U7316 ( .A(n10434), .B(n7013), .Z(n7015) );
  NANDN U7317 ( .A(b[0]), .B(a[169]), .Z(n7014) );
  AND U7318 ( .A(n7015), .B(n7014), .Z(n7042) );
  XOR U7319 ( .A(b[5]), .B(a[166]), .Z(n7049) );
  NAND U7320 ( .A(n7049), .B(n10481), .Z(n7018) );
  NAND U7321 ( .A(n7016), .B(n10482), .Z(n7017) );
  NAND U7322 ( .A(n7018), .B(n7017), .Z(n7040) );
  NANDN U7323 ( .A(n529), .B(a[162]), .Z(n7041) );
  XNOR U7324 ( .A(n7040), .B(n7041), .Z(n7043) );
  XOR U7325 ( .A(n7042), .B(n7043), .Z(n7037) );
  XOR U7326 ( .A(n7036), .B(n7037), .Z(n7058) );
  XOR U7327 ( .A(n7059), .B(n7058), .Z(n7060) );
  XNOR U7328 ( .A(n7061), .B(n7060), .Z(n7030) );
  NAND U7329 ( .A(n7020), .B(n7019), .Z(n7024) );
  NAND U7330 ( .A(n7022), .B(n7021), .Z(n7023) );
  NAND U7331 ( .A(n7024), .B(n7023), .Z(n7031) );
  XNOR U7332 ( .A(n7030), .B(n7031), .Z(n7032) );
  XNOR U7333 ( .A(n7033), .B(n7032), .Z(n7064) );
  XNOR U7334 ( .A(n7064), .B(sreg[418]), .Z(n7066) );
  NAND U7335 ( .A(n7025), .B(sreg[417]), .Z(n7029) );
  OR U7336 ( .A(n7027), .B(n7026), .Z(n7028) );
  AND U7337 ( .A(n7029), .B(n7028), .Z(n7065) );
  XOR U7338 ( .A(n7066), .B(n7065), .Z(c[418]) );
  NANDN U7339 ( .A(n7035), .B(n7034), .Z(n7039) );
  NAND U7340 ( .A(n7037), .B(n7036), .Z(n7038) );
  NAND U7341 ( .A(n7039), .B(n7038), .Z(n7100) );
  NANDN U7342 ( .A(n7041), .B(n7040), .Z(n7045) );
  NAND U7343 ( .A(n7043), .B(n7042), .Z(n7044) );
  NAND U7344 ( .A(n7045), .B(n7044), .Z(n7098) );
  NANDN U7345 ( .A(n527), .B(a[171]), .Z(n7046) );
  XOR U7346 ( .A(n10434), .B(n7046), .Z(n7048) );
  NANDN U7347 ( .A(b[0]), .B(a[170]), .Z(n7047) );
  AND U7348 ( .A(n7048), .B(n7047), .Z(n7081) );
  XOR U7349 ( .A(b[5]), .B(a[167]), .Z(n7094) );
  NAND U7350 ( .A(n7094), .B(n10481), .Z(n7051) );
  NAND U7351 ( .A(n7049), .B(n10482), .Z(n7050) );
  NAND U7352 ( .A(n7051), .B(n7050), .Z(n7079) );
  NANDN U7353 ( .A(n529), .B(a[163]), .Z(n7080) );
  XNOR U7354 ( .A(n7079), .B(n7080), .Z(n7082) );
  XOR U7355 ( .A(n7081), .B(n7082), .Z(n7075) );
  XNOR U7356 ( .A(b[7]), .B(a[165]), .Z(n7085) );
  NANDN U7357 ( .A(n7085), .B(n10545), .Z(n7054) );
  NANDN U7358 ( .A(n7052), .B(n10546), .Z(n7053) );
  NAND U7359 ( .A(n7054), .B(n7053), .Z(n7073) );
  XNOR U7360 ( .A(b[3]), .B(a[169]), .Z(n7088) );
  NANDN U7361 ( .A(n7088), .B(n10398), .Z(n7057) );
  NANDN U7362 ( .A(n7055), .B(n10399), .Z(n7056) );
  AND U7363 ( .A(n7057), .B(n7056), .Z(n7074) );
  XNOR U7364 ( .A(n7073), .B(n7074), .Z(n7076) );
  XOR U7365 ( .A(n7075), .B(n7076), .Z(n7097) );
  XOR U7366 ( .A(n7098), .B(n7097), .Z(n7099) );
  XNOR U7367 ( .A(n7100), .B(n7099), .Z(n7069) );
  NAND U7368 ( .A(n7059), .B(n7058), .Z(n7063) );
  NAND U7369 ( .A(n7061), .B(n7060), .Z(n7062) );
  NAND U7370 ( .A(n7063), .B(n7062), .Z(n7070) );
  XNOR U7371 ( .A(n7069), .B(n7070), .Z(n7071) );
  XNOR U7372 ( .A(n7072), .B(n7071), .Z(n7103) );
  XNOR U7373 ( .A(n7103), .B(sreg[419]), .Z(n7105) );
  NAND U7374 ( .A(n7064), .B(sreg[418]), .Z(n7068) );
  OR U7375 ( .A(n7066), .B(n7065), .Z(n7067) );
  AND U7376 ( .A(n7068), .B(n7067), .Z(n7104) );
  XOR U7377 ( .A(n7105), .B(n7104), .Z(c[419]) );
  NANDN U7378 ( .A(n7074), .B(n7073), .Z(n7078) );
  NAND U7379 ( .A(n7076), .B(n7075), .Z(n7077) );
  NAND U7380 ( .A(n7078), .B(n7077), .Z(n7139) );
  NANDN U7381 ( .A(n7080), .B(n7079), .Z(n7084) );
  NAND U7382 ( .A(n7082), .B(n7081), .Z(n7083) );
  NAND U7383 ( .A(n7084), .B(n7083), .Z(n7137) );
  XNOR U7384 ( .A(b[7]), .B(a[166]), .Z(n7124) );
  NANDN U7385 ( .A(n7124), .B(n10545), .Z(n7087) );
  NANDN U7386 ( .A(n7085), .B(n10546), .Z(n7086) );
  NAND U7387 ( .A(n7087), .B(n7086), .Z(n7112) );
  XNOR U7388 ( .A(b[3]), .B(a[170]), .Z(n7127) );
  NANDN U7389 ( .A(n7127), .B(n10398), .Z(n7090) );
  NANDN U7390 ( .A(n7088), .B(n10399), .Z(n7089) );
  AND U7391 ( .A(n7090), .B(n7089), .Z(n7113) );
  XNOR U7392 ( .A(n7112), .B(n7113), .Z(n7114) );
  NANDN U7393 ( .A(n527), .B(a[172]), .Z(n7091) );
  XOR U7394 ( .A(n10434), .B(n7091), .Z(n7093) );
  NANDN U7395 ( .A(b[0]), .B(a[171]), .Z(n7092) );
  AND U7396 ( .A(n7093), .B(n7092), .Z(n7120) );
  XOR U7397 ( .A(b[5]), .B(a[168]), .Z(n7133) );
  NAND U7398 ( .A(n7133), .B(n10481), .Z(n7096) );
  NAND U7399 ( .A(n7094), .B(n10482), .Z(n7095) );
  NAND U7400 ( .A(n7096), .B(n7095), .Z(n7118) );
  NANDN U7401 ( .A(n529), .B(a[164]), .Z(n7119) );
  XNOR U7402 ( .A(n7118), .B(n7119), .Z(n7121) );
  XOR U7403 ( .A(n7120), .B(n7121), .Z(n7115) );
  XOR U7404 ( .A(n7114), .B(n7115), .Z(n7136) );
  XOR U7405 ( .A(n7137), .B(n7136), .Z(n7138) );
  XNOR U7406 ( .A(n7139), .B(n7138), .Z(n7108) );
  NAND U7407 ( .A(n7098), .B(n7097), .Z(n7102) );
  NAND U7408 ( .A(n7100), .B(n7099), .Z(n7101) );
  NAND U7409 ( .A(n7102), .B(n7101), .Z(n7109) );
  XNOR U7410 ( .A(n7108), .B(n7109), .Z(n7110) );
  XNOR U7411 ( .A(n7111), .B(n7110), .Z(n7142) );
  XNOR U7412 ( .A(n7142), .B(sreg[420]), .Z(n7144) );
  NAND U7413 ( .A(n7103), .B(sreg[419]), .Z(n7107) );
  OR U7414 ( .A(n7105), .B(n7104), .Z(n7106) );
  AND U7415 ( .A(n7107), .B(n7106), .Z(n7143) );
  XOR U7416 ( .A(n7144), .B(n7143), .Z(c[420]) );
  NANDN U7417 ( .A(n7113), .B(n7112), .Z(n7117) );
  NAND U7418 ( .A(n7115), .B(n7114), .Z(n7116) );
  NAND U7419 ( .A(n7117), .B(n7116), .Z(n7178) );
  NANDN U7420 ( .A(n7119), .B(n7118), .Z(n7123) );
  NAND U7421 ( .A(n7121), .B(n7120), .Z(n7122) );
  NAND U7422 ( .A(n7123), .B(n7122), .Z(n7176) );
  XNOR U7423 ( .A(b[7]), .B(a[167]), .Z(n7163) );
  NANDN U7424 ( .A(n7163), .B(n10545), .Z(n7126) );
  NANDN U7425 ( .A(n7124), .B(n10546), .Z(n7125) );
  NAND U7426 ( .A(n7126), .B(n7125), .Z(n7151) );
  XNOR U7427 ( .A(b[3]), .B(a[171]), .Z(n7166) );
  NANDN U7428 ( .A(n7166), .B(n10398), .Z(n7129) );
  NANDN U7429 ( .A(n7127), .B(n10399), .Z(n7128) );
  AND U7430 ( .A(n7129), .B(n7128), .Z(n7152) );
  XNOR U7431 ( .A(n7151), .B(n7152), .Z(n7153) );
  NANDN U7432 ( .A(n527), .B(a[173]), .Z(n7130) );
  XOR U7433 ( .A(n10434), .B(n7130), .Z(n7132) );
  NANDN U7434 ( .A(b[0]), .B(a[172]), .Z(n7131) );
  AND U7435 ( .A(n7132), .B(n7131), .Z(n7159) );
  XOR U7436 ( .A(b[5]), .B(a[169]), .Z(n7172) );
  NAND U7437 ( .A(n7172), .B(n10481), .Z(n7135) );
  NAND U7438 ( .A(n7133), .B(n10482), .Z(n7134) );
  NAND U7439 ( .A(n7135), .B(n7134), .Z(n7157) );
  NANDN U7440 ( .A(n529), .B(a[165]), .Z(n7158) );
  XNOR U7441 ( .A(n7157), .B(n7158), .Z(n7160) );
  XOR U7442 ( .A(n7159), .B(n7160), .Z(n7154) );
  XOR U7443 ( .A(n7153), .B(n7154), .Z(n7175) );
  XOR U7444 ( .A(n7176), .B(n7175), .Z(n7177) );
  XNOR U7445 ( .A(n7178), .B(n7177), .Z(n7147) );
  NAND U7446 ( .A(n7137), .B(n7136), .Z(n7141) );
  NAND U7447 ( .A(n7139), .B(n7138), .Z(n7140) );
  NAND U7448 ( .A(n7141), .B(n7140), .Z(n7148) );
  XNOR U7449 ( .A(n7147), .B(n7148), .Z(n7149) );
  XNOR U7450 ( .A(n7150), .B(n7149), .Z(n7181) );
  XNOR U7451 ( .A(n7181), .B(sreg[421]), .Z(n7183) );
  NAND U7452 ( .A(n7142), .B(sreg[420]), .Z(n7146) );
  OR U7453 ( .A(n7144), .B(n7143), .Z(n7145) );
  AND U7454 ( .A(n7146), .B(n7145), .Z(n7182) );
  XOR U7455 ( .A(n7183), .B(n7182), .Z(c[421]) );
  NANDN U7456 ( .A(n7152), .B(n7151), .Z(n7156) );
  NAND U7457 ( .A(n7154), .B(n7153), .Z(n7155) );
  NAND U7458 ( .A(n7156), .B(n7155), .Z(n7217) );
  NANDN U7459 ( .A(n7158), .B(n7157), .Z(n7162) );
  NAND U7460 ( .A(n7160), .B(n7159), .Z(n7161) );
  NAND U7461 ( .A(n7162), .B(n7161), .Z(n7215) );
  XNOR U7462 ( .A(b[7]), .B(a[168]), .Z(n7202) );
  NANDN U7463 ( .A(n7202), .B(n10545), .Z(n7165) );
  NANDN U7464 ( .A(n7163), .B(n10546), .Z(n7164) );
  NAND U7465 ( .A(n7165), .B(n7164), .Z(n7190) );
  XNOR U7466 ( .A(b[3]), .B(a[172]), .Z(n7205) );
  NANDN U7467 ( .A(n7205), .B(n10398), .Z(n7168) );
  NANDN U7468 ( .A(n7166), .B(n10399), .Z(n7167) );
  AND U7469 ( .A(n7168), .B(n7167), .Z(n7191) );
  XNOR U7470 ( .A(n7190), .B(n7191), .Z(n7192) );
  NANDN U7471 ( .A(n527), .B(a[174]), .Z(n7169) );
  XOR U7472 ( .A(n10434), .B(n7169), .Z(n7171) );
  NANDN U7473 ( .A(b[0]), .B(a[173]), .Z(n7170) );
  AND U7474 ( .A(n7171), .B(n7170), .Z(n7198) );
  XOR U7475 ( .A(b[5]), .B(a[170]), .Z(n7211) );
  NAND U7476 ( .A(n7211), .B(n10481), .Z(n7174) );
  NAND U7477 ( .A(n7172), .B(n10482), .Z(n7173) );
  NAND U7478 ( .A(n7174), .B(n7173), .Z(n7196) );
  NANDN U7479 ( .A(n529), .B(a[166]), .Z(n7197) );
  XNOR U7480 ( .A(n7196), .B(n7197), .Z(n7199) );
  XOR U7481 ( .A(n7198), .B(n7199), .Z(n7193) );
  XOR U7482 ( .A(n7192), .B(n7193), .Z(n7214) );
  XOR U7483 ( .A(n7215), .B(n7214), .Z(n7216) );
  XNOR U7484 ( .A(n7217), .B(n7216), .Z(n7186) );
  NAND U7485 ( .A(n7176), .B(n7175), .Z(n7180) );
  NAND U7486 ( .A(n7178), .B(n7177), .Z(n7179) );
  NAND U7487 ( .A(n7180), .B(n7179), .Z(n7187) );
  XNOR U7488 ( .A(n7186), .B(n7187), .Z(n7188) );
  XNOR U7489 ( .A(n7189), .B(n7188), .Z(n7220) );
  XNOR U7490 ( .A(n7220), .B(sreg[422]), .Z(n7222) );
  NAND U7491 ( .A(n7181), .B(sreg[421]), .Z(n7185) );
  OR U7492 ( .A(n7183), .B(n7182), .Z(n7184) );
  AND U7493 ( .A(n7185), .B(n7184), .Z(n7221) );
  XOR U7494 ( .A(n7222), .B(n7221), .Z(c[422]) );
  NANDN U7495 ( .A(n7191), .B(n7190), .Z(n7195) );
  NAND U7496 ( .A(n7193), .B(n7192), .Z(n7194) );
  NAND U7497 ( .A(n7195), .B(n7194), .Z(n7256) );
  NANDN U7498 ( .A(n7197), .B(n7196), .Z(n7201) );
  NAND U7499 ( .A(n7199), .B(n7198), .Z(n7200) );
  NAND U7500 ( .A(n7201), .B(n7200), .Z(n7254) );
  XNOR U7501 ( .A(b[7]), .B(a[169]), .Z(n7241) );
  NANDN U7502 ( .A(n7241), .B(n10545), .Z(n7204) );
  NANDN U7503 ( .A(n7202), .B(n10546), .Z(n7203) );
  NAND U7504 ( .A(n7204), .B(n7203), .Z(n7229) );
  XNOR U7505 ( .A(b[3]), .B(a[173]), .Z(n7244) );
  NANDN U7506 ( .A(n7244), .B(n10398), .Z(n7207) );
  NANDN U7507 ( .A(n7205), .B(n10399), .Z(n7206) );
  AND U7508 ( .A(n7207), .B(n7206), .Z(n7230) );
  XNOR U7509 ( .A(n7229), .B(n7230), .Z(n7231) );
  NANDN U7510 ( .A(n527), .B(a[175]), .Z(n7208) );
  XOR U7511 ( .A(n10434), .B(n7208), .Z(n7210) );
  NANDN U7512 ( .A(b[0]), .B(a[174]), .Z(n7209) );
  AND U7513 ( .A(n7210), .B(n7209), .Z(n7237) );
  XOR U7514 ( .A(b[5]), .B(a[171]), .Z(n7250) );
  NAND U7515 ( .A(n7250), .B(n10481), .Z(n7213) );
  NAND U7516 ( .A(n7211), .B(n10482), .Z(n7212) );
  NAND U7517 ( .A(n7213), .B(n7212), .Z(n7235) );
  NANDN U7518 ( .A(n529), .B(a[167]), .Z(n7236) );
  XNOR U7519 ( .A(n7235), .B(n7236), .Z(n7238) );
  XOR U7520 ( .A(n7237), .B(n7238), .Z(n7232) );
  XOR U7521 ( .A(n7231), .B(n7232), .Z(n7253) );
  XOR U7522 ( .A(n7254), .B(n7253), .Z(n7255) );
  XNOR U7523 ( .A(n7256), .B(n7255), .Z(n7225) );
  NAND U7524 ( .A(n7215), .B(n7214), .Z(n7219) );
  NAND U7525 ( .A(n7217), .B(n7216), .Z(n7218) );
  NAND U7526 ( .A(n7219), .B(n7218), .Z(n7226) );
  XNOR U7527 ( .A(n7225), .B(n7226), .Z(n7227) );
  XNOR U7528 ( .A(n7228), .B(n7227), .Z(n7259) );
  XNOR U7529 ( .A(n7259), .B(sreg[423]), .Z(n7261) );
  NAND U7530 ( .A(n7220), .B(sreg[422]), .Z(n7224) );
  OR U7531 ( .A(n7222), .B(n7221), .Z(n7223) );
  AND U7532 ( .A(n7224), .B(n7223), .Z(n7260) );
  XOR U7533 ( .A(n7261), .B(n7260), .Z(c[423]) );
  NANDN U7534 ( .A(n7230), .B(n7229), .Z(n7234) );
  NAND U7535 ( .A(n7232), .B(n7231), .Z(n7233) );
  NAND U7536 ( .A(n7234), .B(n7233), .Z(n7295) );
  NANDN U7537 ( .A(n7236), .B(n7235), .Z(n7240) );
  NAND U7538 ( .A(n7238), .B(n7237), .Z(n7239) );
  NAND U7539 ( .A(n7240), .B(n7239), .Z(n7293) );
  XNOR U7540 ( .A(b[7]), .B(a[170]), .Z(n7280) );
  NANDN U7541 ( .A(n7280), .B(n10545), .Z(n7243) );
  NANDN U7542 ( .A(n7241), .B(n10546), .Z(n7242) );
  NAND U7543 ( .A(n7243), .B(n7242), .Z(n7268) );
  XNOR U7544 ( .A(b[3]), .B(a[174]), .Z(n7283) );
  NANDN U7545 ( .A(n7283), .B(n10398), .Z(n7246) );
  NANDN U7546 ( .A(n7244), .B(n10399), .Z(n7245) );
  AND U7547 ( .A(n7246), .B(n7245), .Z(n7269) );
  XNOR U7548 ( .A(n7268), .B(n7269), .Z(n7270) );
  NANDN U7549 ( .A(n527), .B(a[176]), .Z(n7247) );
  XOR U7550 ( .A(n10434), .B(n7247), .Z(n7249) );
  NANDN U7551 ( .A(b[0]), .B(a[175]), .Z(n7248) );
  AND U7552 ( .A(n7249), .B(n7248), .Z(n7276) );
  XOR U7553 ( .A(b[5]), .B(a[172]), .Z(n7289) );
  NAND U7554 ( .A(n7289), .B(n10481), .Z(n7252) );
  NAND U7555 ( .A(n7250), .B(n10482), .Z(n7251) );
  NAND U7556 ( .A(n7252), .B(n7251), .Z(n7274) );
  NANDN U7557 ( .A(n529), .B(a[168]), .Z(n7275) );
  XNOR U7558 ( .A(n7274), .B(n7275), .Z(n7277) );
  XOR U7559 ( .A(n7276), .B(n7277), .Z(n7271) );
  XOR U7560 ( .A(n7270), .B(n7271), .Z(n7292) );
  XOR U7561 ( .A(n7293), .B(n7292), .Z(n7294) );
  XNOR U7562 ( .A(n7295), .B(n7294), .Z(n7264) );
  NAND U7563 ( .A(n7254), .B(n7253), .Z(n7258) );
  NAND U7564 ( .A(n7256), .B(n7255), .Z(n7257) );
  NAND U7565 ( .A(n7258), .B(n7257), .Z(n7265) );
  XNOR U7566 ( .A(n7264), .B(n7265), .Z(n7266) );
  XNOR U7567 ( .A(n7267), .B(n7266), .Z(n7298) );
  XNOR U7568 ( .A(n7298), .B(sreg[424]), .Z(n7300) );
  NAND U7569 ( .A(n7259), .B(sreg[423]), .Z(n7263) );
  OR U7570 ( .A(n7261), .B(n7260), .Z(n7262) );
  AND U7571 ( .A(n7263), .B(n7262), .Z(n7299) );
  XOR U7572 ( .A(n7300), .B(n7299), .Z(c[424]) );
  NANDN U7573 ( .A(n7269), .B(n7268), .Z(n7273) );
  NAND U7574 ( .A(n7271), .B(n7270), .Z(n7272) );
  NAND U7575 ( .A(n7273), .B(n7272), .Z(n7334) );
  NANDN U7576 ( .A(n7275), .B(n7274), .Z(n7279) );
  NAND U7577 ( .A(n7277), .B(n7276), .Z(n7278) );
  NAND U7578 ( .A(n7279), .B(n7278), .Z(n7332) );
  XNOR U7579 ( .A(b[7]), .B(a[171]), .Z(n7319) );
  NANDN U7580 ( .A(n7319), .B(n10545), .Z(n7282) );
  NANDN U7581 ( .A(n7280), .B(n10546), .Z(n7281) );
  NAND U7582 ( .A(n7282), .B(n7281), .Z(n7307) );
  XNOR U7583 ( .A(b[3]), .B(a[175]), .Z(n7322) );
  NANDN U7584 ( .A(n7322), .B(n10398), .Z(n7285) );
  NANDN U7585 ( .A(n7283), .B(n10399), .Z(n7284) );
  AND U7586 ( .A(n7285), .B(n7284), .Z(n7308) );
  XNOR U7587 ( .A(n7307), .B(n7308), .Z(n7309) );
  NANDN U7588 ( .A(n527), .B(a[177]), .Z(n7286) );
  XOR U7589 ( .A(n10434), .B(n7286), .Z(n7288) );
  NANDN U7590 ( .A(b[0]), .B(a[176]), .Z(n7287) );
  AND U7591 ( .A(n7288), .B(n7287), .Z(n7315) );
  XOR U7592 ( .A(b[5]), .B(a[173]), .Z(n7328) );
  NAND U7593 ( .A(n7328), .B(n10481), .Z(n7291) );
  NAND U7594 ( .A(n7289), .B(n10482), .Z(n7290) );
  NAND U7595 ( .A(n7291), .B(n7290), .Z(n7313) );
  NANDN U7596 ( .A(n529), .B(a[169]), .Z(n7314) );
  XNOR U7597 ( .A(n7313), .B(n7314), .Z(n7316) );
  XOR U7598 ( .A(n7315), .B(n7316), .Z(n7310) );
  XOR U7599 ( .A(n7309), .B(n7310), .Z(n7331) );
  XOR U7600 ( .A(n7332), .B(n7331), .Z(n7333) );
  XNOR U7601 ( .A(n7334), .B(n7333), .Z(n7303) );
  NAND U7602 ( .A(n7293), .B(n7292), .Z(n7297) );
  NAND U7603 ( .A(n7295), .B(n7294), .Z(n7296) );
  NAND U7604 ( .A(n7297), .B(n7296), .Z(n7304) );
  XNOR U7605 ( .A(n7303), .B(n7304), .Z(n7305) );
  XNOR U7606 ( .A(n7306), .B(n7305), .Z(n7337) );
  XNOR U7607 ( .A(n7337), .B(sreg[425]), .Z(n7339) );
  NAND U7608 ( .A(n7298), .B(sreg[424]), .Z(n7302) );
  OR U7609 ( .A(n7300), .B(n7299), .Z(n7301) );
  AND U7610 ( .A(n7302), .B(n7301), .Z(n7338) );
  XOR U7611 ( .A(n7339), .B(n7338), .Z(c[425]) );
  NANDN U7612 ( .A(n7308), .B(n7307), .Z(n7312) );
  NAND U7613 ( .A(n7310), .B(n7309), .Z(n7311) );
  NAND U7614 ( .A(n7312), .B(n7311), .Z(n7373) );
  NANDN U7615 ( .A(n7314), .B(n7313), .Z(n7318) );
  NAND U7616 ( .A(n7316), .B(n7315), .Z(n7317) );
  NAND U7617 ( .A(n7318), .B(n7317), .Z(n7371) );
  XNOR U7618 ( .A(b[7]), .B(a[172]), .Z(n7358) );
  NANDN U7619 ( .A(n7358), .B(n10545), .Z(n7321) );
  NANDN U7620 ( .A(n7319), .B(n10546), .Z(n7320) );
  NAND U7621 ( .A(n7321), .B(n7320), .Z(n7346) );
  XNOR U7622 ( .A(b[3]), .B(a[176]), .Z(n7361) );
  NANDN U7623 ( .A(n7361), .B(n10398), .Z(n7324) );
  NANDN U7624 ( .A(n7322), .B(n10399), .Z(n7323) );
  AND U7625 ( .A(n7324), .B(n7323), .Z(n7347) );
  XNOR U7626 ( .A(n7346), .B(n7347), .Z(n7348) );
  NANDN U7627 ( .A(n527), .B(a[178]), .Z(n7325) );
  XOR U7628 ( .A(n10434), .B(n7325), .Z(n7327) );
  NANDN U7629 ( .A(b[0]), .B(a[177]), .Z(n7326) );
  AND U7630 ( .A(n7327), .B(n7326), .Z(n7354) );
  XOR U7631 ( .A(b[5]), .B(a[174]), .Z(n7367) );
  NAND U7632 ( .A(n7367), .B(n10481), .Z(n7330) );
  NAND U7633 ( .A(n7328), .B(n10482), .Z(n7329) );
  NAND U7634 ( .A(n7330), .B(n7329), .Z(n7352) );
  NANDN U7635 ( .A(n529), .B(a[170]), .Z(n7353) );
  XNOR U7636 ( .A(n7352), .B(n7353), .Z(n7355) );
  XOR U7637 ( .A(n7354), .B(n7355), .Z(n7349) );
  XOR U7638 ( .A(n7348), .B(n7349), .Z(n7370) );
  XOR U7639 ( .A(n7371), .B(n7370), .Z(n7372) );
  XNOR U7640 ( .A(n7373), .B(n7372), .Z(n7342) );
  NAND U7641 ( .A(n7332), .B(n7331), .Z(n7336) );
  NAND U7642 ( .A(n7334), .B(n7333), .Z(n7335) );
  NAND U7643 ( .A(n7336), .B(n7335), .Z(n7343) );
  XNOR U7644 ( .A(n7342), .B(n7343), .Z(n7344) );
  XNOR U7645 ( .A(n7345), .B(n7344), .Z(n7376) );
  XNOR U7646 ( .A(n7376), .B(sreg[426]), .Z(n7378) );
  NAND U7647 ( .A(n7337), .B(sreg[425]), .Z(n7341) );
  OR U7648 ( .A(n7339), .B(n7338), .Z(n7340) );
  AND U7649 ( .A(n7341), .B(n7340), .Z(n7377) );
  XOR U7650 ( .A(n7378), .B(n7377), .Z(c[426]) );
  NANDN U7651 ( .A(n7347), .B(n7346), .Z(n7351) );
  NAND U7652 ( .A(n7349), .B(n7348), .Z(n7350) );
  NAND U7653 ( .A(n7351), .B(n7350), .Z(n7412) );
  NANDN U7654 ( .A(n7353), .B(n7352), .Z(n7357) );
  NAND U7655 ( .A(n7355), .B(n7354), .Z(n7356) );
  NAND U7656 ( .A(n7357), .B(n7356), .Z(n7410) );
  XNOR U7657 ( .A(b[7]), .B(a[173]), .Z(n7397) );
  NANDN U7658 ( .A(n7397), .B(n10545), .Z(n7360) );
  NANDN U7659 ( .A(n7358), .B(n10546), .Z(n7359) );
  NAND U7660 ( .A(n7360), .B(n7359), .Z(n7385) );
  XNOR U7661 ( .A(b[3]), .B(a[177]), .Z(n7400) );
  NANDN U7662 ( .A(n7400), .B(n10398), .Z(n7363) );
  NANDN U7663 ( .A(n7361), .B(n10399), .Z(n7362) );
  AND U7664 ( .A(n7363), .B(n7362), .Z(n7386) );
  XNOR U7665 ( .A(n7385), .B(n7386), .Z(n7387) );
  NANDN U7666 ( .A(n527), .B(a[179]), .Z(n7364) );
  XOR U7667 ( .A(n10434), .B(n7364), .Z(n7366) );
  NANDN U7668 ( .A(b[0]), .B(a[178]), .Z(n7365) );
  AND U7669 ( .A(n7366), .B(n7365), .Z(n7393) );
  XOR U7670 ( .A(b[5]), .B(a[175]), .Z(n7406) );
  NAND U7671 ( .A(n7406), .B(n10481), .Z(n7369) );
  NAND U7672 ( .A(n7367), .B(n10482), .Z(n7368) );
  NAND U7673 ( .A(n7369), .B(n7368), .Z(n7391) );
  NANDN U7674 ( .A(n529), .B(a[171]), .Z(n7392) );
  XNOR U7675 ( .A(n7391), .B(n7392), .Z(n7394) );
  XOR U7676 ( .A(n7393), .B(n7394), .Z(n7388) );
  XOR U7677 ( .A(n7387), .B(n7388), .Z(n7409) );
  XOR U7678 ( .A(n7410), .B(n7409), .Z(n7411) );
  XNOR U7679 ( .A(n7412), .B(n7411), .Z(n7381) );
  NAND U7680 ( .A(n7371), .B(n7370), .Z(n7375) );
  NAND U7681 ( .A(n7373), .B(n7372), .Z(n7374) );
  NAND U7682 ( .A(n7375), .B(n7374), .Z(n7382) );
  XNOR U7683 ( .A(n7381), .B(n7382), .Z(n7383) );
  XNOR U7684 ( .A(n7384), .B(n7383), .Z(n7415) );
  XNOR U7685 ( .A(n7415), .B(sreg[427]), .Z(n7417) );
  NAND U7686 ( .A(n7376), .B(sreg[426]), .Z(n7380) );
  OR U7687 ( .A(n7378), .B(n7377), .Z(n7379) );
  AND U7688 ( .A(n7380), .B(n7379), .Z(n7416) );
  XOR U7689 ( .A(n7417), .B(n7416), .Z(c[427]) );
  NANDN U7690 ( .A(n7386), .B(n7385), .Z(n7390) );
  NAND U7691 ( .A(n7388), .B(n7387), .Z(n7389) );
  NAND U7692 ( .A(n7390), .B(n7389), .Z(n7451) );
  NANDN U7693 ( .A(n7392), .B(n7391), .Z(n7396) );
  NAND U7694 ( .A(n7394), .B(n7393), .Z(n7395) );
  NAND U7695 ( .A(n7396), .B(n7395), .Z(n7449) );
  XNOR U7696 ( .A(b[7]), .B(a[174]), .Z(n7436) );
  NANDN U7697 ( .A(n7436), .B(n10545), .Z(n7399) );
  NANDN U7698 ( .A(n7397), .B(n10546), .Z(n7398) );
  NAND U7699 ( .A(n7399), .B(n7398), .Z(n7424) );
  XNOR U7700 ( .A(b[3]), .B(a[178]), .Z(n7439) );
  NANDN U7701 ( .A(n7439), .B(n10398), .Z(n7402) );
  NANDN U7702 ( .A(n7400), .B(n10399), .Z(n7401) );
  AND U7703 ( .A(n7402), .B(n7401), .Z(n7425) );
  XNOR U7704 ( .A(n7424), .B(n7425), .Z(n7426) );
  NANDN U7705 ( .A(n527), .B(a[180]), .Z(n7403) );
  XOR U7706 ( .A(n10434), .B(n7403), .Z(n7405) );
  NANDN U7707 ( .A(b[0]), .B(a[179]), .Z(n7404) );
  AND U7708 ( .A(n7405), .B(n7404), .Z(n7432) );
  XOR U7709 ( .A(b[5]), .B(a[176]), .Z(n7445) );
  NAND U7710 ( .A(n7445), .B(n10481), .Z(n7408) );
  NAND U7711 ( .A(n7406), .B(n10482), .Z(n7407) );
  NAND U7712 ( .A(n7408), .B(n7407), .Z(n7430) );
  NANDN U7713 ( .A(n529), .B(a[172]), .Z(n7431) );
  XNOR U7714 ( .A(n7430), .B(n7431), .Z(n7433) );
  XOR U7715 ( .A(n7432), .B(n7433), .Z(n7427) );
  XOR U7716 ( .A(n7426), .B(n7427), .Z(n7448) );
  XOR U7717 ( .A(n7449), .B(n7448), .Z(n7450) );
  XNOR U7718 ( .A(n7451), .B(n7450), .Z(n7420) );
  NAND U7719 ( .A(n7410), .B(n7409), .Z(n7414) );
  NAND U7720 ( .A(n7412), .B(n7411), .Z(n7413) );
  NAND U7721 ( .A(n7414), .B(n7413), .Z(n7421) );
  XNOR U7722 ( .A(n7420), .B(n7421), .Z(n7422) );
  XNOR U7723 ( .A(n7423), .B(n7422), .Z(n7454) );
  XNOR U7724 ( .A(n7454), .B(sreg[428]), .Z(n7456) );
  NAND U7725 ( .A(n7415), .B(sreg[427]), .Z(n7419) );
  OR U7726 ( .A(n7417), .B(n7416), .Z(n7418) );
  AND U7727 ( .A(n7419), .B(n7418), .Z(n7455) );
  XOR U7728 ( .A(n7456), .B(n7455), .Z(c[428]) );
  NANDN U7729 ( .A(n7425), .B(n7424), .Z(n7429) );
  NAND U7730 ( .A(n7427), .B(n7426), .Z(n7428) );
  NAND U7731 ( .A(n7429), .B(n7428), .Z(n7490) );
  NANDN U7732 ( .A(n7431), .B(n7430), .Z(n7435) );
  NAND U7733 ( .A(n7433), .B(n7432), .Z(n7434) );
  NAND U7734 ( .A(n7435), .B(n7434), .Z(n7488) );
  XNOR U7735 ( .A(b[7]), .B(a[175]), .Z(n7475) );
  NANDN U7736 ( .A(n7475), .B(n10545), .Z(n7438) );
  NANDN U7737 ( .A(n7436), .B(n10546), .Z(n7437) );
  NAND U7738 ( .A(n7438), .B(n7437), .Z(n7463) );
  XNOR U7739 ( .A(b[3]), .B(a[179]), .Z(n7478) );
  NANDN U7740 ( .A(n7478), .B(n10398), .Z(n7441) );
  NANDN U7741 ( .A(n7439), .B(n10399), .Z(n7440) );
  AND U7742 ( .A(n7441), .B(n7440), .Z(n7464) );
  XNOR U7743 ( .A(n7463), .B(n7464), .Z(n7465) );
  NANDN U7744 ( .A(n527), .B(a[181]), .Z(n7442) );
  XOR U7745 ( .A(n10434), .B(n7442), .Z(n7444) );
  NANDN U7746 ( .A(b[0]), .B(a[180]), .Z(n7443) );
  AND U7747 ( .A(n7444), .B(n7443), .Z(n7471) );
  XOR U7748 ( .A(b[5]), .B(a[177]), .Z(n7484) );
  NAND U7749 ( .A(n7484), .B(n10481), .Z(n7447) );
  NAND U7750 ( .A(n7445), .B(n10482), .Z(n7446) );
  NAND U7751 ( .A(n7447), .B(n7446), .Z(n7469) );
  NANDN U7752 ( .A(n529), .B(a[173]), .Z(n7470) );
  XNOR U7753 ( .A(n7469), .B(n7470), .Z(n7472) );
  XOR U7754 ( .A(n7471), .B(n7472), .Z(n7466) );
  XOR U7755 ( .A(n7465), .B(n7466), .Z(n7487) );
  XOR U7756 ( .A(n7488), .B(n7487), .Z(n7489) );
  XNOR U7757 ( .A(n7490), .B(n7489), .Z(n7459) );
  NAND U7758 ( .A(n7449), .B(n7448), .Z(n7453) );
  NAND U7759 ( .A(n7451), .B(n7450), .Z(n7452) );
  NAND U7760 ( .A(n7453), .B(n7452), .Z(n7460) );
  XNOR U7761 ( .A(n7459), .B(n7460), .Z(n7461) );
  XNOR U7762 ( .A(n7462), .B(n7461), .Z(n7493) );
  XNOR U7763 ( .A(n7493), .B(sreg[429]), .Z(n7495) );
  NAND U7764 ( .A(n7454), .B(sreg[428]), .Z(n7458) );
  OR U7765 ( .A(n7456), .B(n7455), .Z(n7457) );
  AND U7766 ( .A(n7458), .B(n7457), .Z(n7494) );
  XOR U7767 ( .A(n7495), .B(n7494), .Z(c[429]) );
  NANDN U7768 ( .A(n7464), .B(n7463), .Z(n7468) );
  NAND U7769 ( .A(n7466), .B(n7465), .Z(n7467) );
  NAND U7770 ( .A(n7468), .B(n7467), .Z(n7529) );
  NANDN U7771 ( .A(n7470), .B(n7469), .Z(n7474) );
  NAND U7772 ( .A(n7472), .B(n7471), .Z(n7473) );
  NAND U7773 ( .A(n7474), .B(n7473), .Z(n7527) );
  XNOR U7774 ( .A(b[7]), .B(a[176]), .Z(n7514) );
  NANDN U7775 ( .A(n7514), .B(n10545), .Z(n7477) );
  NANDN U7776 ( .A(n7475), .B(n10546), .Z(n7476) );
  NAND U7777 ( .A(n7477), .B(n7476), .Z(n7502) );
  XNOR U7778 ( .A(b[3]), .B(a[180]), .Z(n7517) );
  NANDN U7779 ( .A(n7517), .B(n10398), .Z(n7480) );
  NANDN U7780 ( .A(n7478), .B(n10399), .Z(n7479) );
  AND U7781 ( .A(n7480), .B(n7479), .Z(n7503) );
  XNOR U7782 ( .A(n7502), .B(n7503), .Z(n7504) );
  NANDN U7783 ( .A(n527), .B(a[182]), .Z(n7481) );
  XOR U7784 ( .A(n10434), .B(n7481), .Z(n7483) );
  NANDN U7785 ( .A(b[0]), .B(a[181]), .Z(n7482) );
  AND U7786 ( .A(n7483), .B(n7482), .Z(n7510) );
  XOR U7787 ( .A(b[5]), .B(a[178]), .Z(n7523) );
  NAND U7788 ( .A(n7523), .B(n10481), .Z(n7486) );
  NAND U7789 ( .A(n7484), .B(n10482), .Z(n7485) );
  NAND U7790 ( .A(n7486), .B(n7485), .Z(n7508) );
  NANDN U7791 ( .A(n529), .B(a[174]), .Z(n7509) );
  XNOR U7792 ( .A(n7508), .B(n7509), .Z(n7511) );
  XOR U7793 ( .A(n7510), .B(n7511), .Z(n7505) );
  XOR U7794 ( .A(n7504), .B(n7505), .Z(n7526) );
  XOR U7795 ( .A(n7527), .B(n7526), .Z(n7528) );
  XNOR U7796 ( .A(n7529), .B(n7528), .Z(n7498) );
  NAND U7797 ( .A(n7488), .B(n7487), .Z(n7492) );
  NAND U7798 ( .A(n7490), .B(n7489), .Z(n7491) );
  NAND U7799 ( .A(n7492), .B(n7491), .Z(n7499) );
  XNOR U7800 ( .A(n7498), .B(n7499), .Z(n7500) );
  XNOR U7801 ( .A(n7501), .B(n7500), .Z(n7532) );
  XNOR U7802 ( .A(n7532), .B(sreg[430]), .Z(n7534) );
  NAND U7803 ( .A(n7493), .B(sreg[429]), .Z(n7497) );
  OR U7804 ( .A(n7495), .B(n7494), .Z(n7496) );
  AND U7805 ( .A(n7497), .B(n7496), .Z(n7533) );
  XOR U7806 ( .A(n7534), .B(n7533), .Z(c[430]) );
  NANDN U7807 ( .A(n7503), .B(n7502), .Z(n7507) );
  NAND U7808 ( .A(n7505), .B(n7504), .Z(n7506) );
  NAND U7809 ( .A(n7507), .B(n7506), .Z(n7568) );
  NANDN U7810 ( .A(n7509), .B(n7508), .Z(n7513) );
  NAND U7811 ( .A(n7511), .B(n7510), .Z(n7512) );
  NAND U7812 ( .A(n7513), .B(n7512), .Z(n7566) );
  XNOR U7813 ( .A(b[7]), .B(a[177]), .Z(n7553) );
  NANDN U7814 ( .A(n7553), .B(n10545), .Z(n7516) );
  NANDN U7815 ( .A(n7514), .B(n10546), .Z(n7515) );
  NAND U7816 ( .A(n7516), .B(n7515), .Z(n7541) );
  XNOR U7817 ( .A(b[3]), .B(a[181]), .Z(n7556) );
  NANDN U7818 ( .A(n7556), .B(n10398), .Z(n7519) );
  NANDN U7819 ( .A(n7517), .B(n10399), .Z(n7518) );
  AND U7820 ( .A(n7519), .B(n7518), .Z(n7542) );
  XNOR U7821 ( .A(n7541), .B(n7542), .Z(n7543) );
  NANDN U7822 ( .A(n527), .B(a[183]), .Z(n7520) );
  XOR U7823 ( .A(n10434), .B(n7520), .Z(n7522) );
  NANDN U7824 ( .A(b[0]), .B(a[182]), .Z(n7521) );
  AND U7825 ( .A(n7522), .B(n7521), .Z(n7549) );
  XOR U7826 ( .A(b[5]), .B(a[179]), .Z(n7562) );
  NAND U7827 ( .A(n7562), .B(n10481), .Z(n7525) );
  NAND U7828 ( .A(n7523), .B(n10482), .Z(n7524) );
  NAND U7829 ( .A(n7525), .B(n7524), .Z(n7547) );
  NANDN U7830 ( .A(n529), .B(a[175]), .Z(n7548) );
  XNOR U7831 ( .A(n7547), .B(n7548), .Z(n7550) );
  XOR U7832 ( .A(n7549), .B(n7550), .Z(n7544) );
  XOR U7833 ( .A(n7543), .B(n7544), .Z(n7565) );
  XOR U7834 ( .A(n7566), .B(n7565), .Z(n7567) );
  XNOR U7835 ( .A(n7568), .B(n7567), .Z(n7537) );
  NAND U7836 ( .A(n7527), .B(n7526), .Z(n7531) );
  NAND U7837 ( .A(n7529), .B(n7528), .Z(n7530) );
  NAND U7838 ( .A(n7531), .B(n7530), .Z(n7538) );
  XNOR U7839 ( .A(n7537), .B(n7538), .Z(n7539) );
  XNOR U7840 ( .A(n7540), .B(n7539), .Z(n7571) );
  XNOR U7841 ( .A(n7571), .B(sreg[431]), .Z(n7573) );
  NAND U7842 ( .A(n7532), .B(sreg[430]), .Z(n7536) );
  OR U7843 ( .A(n7534), .B(n7533), .Z(n7535) );
  AND U7844 ( .A(n7536), .B(n7535), .Z(n7572) );
  XOR U7845 ( .A(n7573), .B(n7572), .Z(c[431]) );
  NANDN U7846 ( .A(n7542), .B(n7541), .Z(n7546) );
  NAND U7847 ( .A(n7544), .B(n7543), .Z(n7545) );
  NAND U7848 ( .A(n7546), .B(n7545), .Z(n7607) );
  NANDN U7849 ( .A(n7548), .B(n7547), .Z(n7552) );
  NAND U7850 ( .A(n7550), .B(n7549), .Z(n7551) );
  NAND U7851 ( .A(n7552), .B(n7551), .Z(n7605) );
  XNOR U7852 ( .A(b[7]), .B(a[178]), .Z(n7592) );
  NANDN U7853 ( .A(n7592), .B(n10545), .Z(n7555) );
  NANDN U7854 ( .A(n7553), .B(n10546), .Z(n7554) );
  NAND U7855 ( .A(n7555), .B(n7554), .Z(n7580) );
  XNOR U7856 ( .A(b[3]), .B(a[182]), .Z(n7595) );
  NANDN U7857 ( .A(n7595), .B(n10398), .Z(n7558) );
  NANDN U7858 ( .A(n7556), .B(n10399), .Z(n7557) );
  AND U7859 ( .A(n7558), .B(n7557), .Z(n7581) );
  XNOR U7860 ( .A(n7580), .B(n7581), .Z(n7582) );
  NANDN U7861 ( .A(n527), .B(a[184]), .Z(n7559) );
  XOR U7862 ( .A(n10434), .B(n7559), .Z(n7561) );
  NANDN U7863 ( .A(b[0]), .B(a[183]), .Z(n7560) );
  AND U7864 ( .A(n7561), .B(n7560), .Z(n7588) );
  XOR U7865 ( .A(b[5]), .B(a[180]), .Z(n7601) );
  NAND U7866 ( .A(n7601), .B(n10481), .Z(n7564) );
  NAND U7867 ( .A(n7562), .B(n10482), .Z(n7563) );
  NAND U7868 ( .A(n7564), .B(n7563), .Z(n7586) );
  NANDN U7869 ( .A(n529), .B(a[176]), .Z(n7587) );
  XNOR U7870 ( .A(n7586), .B(n7587), .Z(n7589) );
  XOR U7871 ( .A(n7588), .B(n7589), .Z(n7583) );
  XOR U7872 ( .A(n7582), .B(n7583), .Z(n7604) );
  XOR U7873 ( .A(n7605), .B(n7604), .Z(n7606) );
  XNOR U7874 ( .A(n7607), .B(n7606), .Z(n7576) );
  NAND U7875 ( .A(n7566), .B(n7565), .Z(n7570) );
  NAND U7876 ( .A(n7568), .B(n7567), .Z(n7569) );
  NAND U7877 ( .A(n7570), .B(n7569), .Z(n7577) );
  XNOR U7878 ( .A(n7576), .B(n7577), .Z(n7578) );
  XNOR U7879 ( .A(n7579), .B(n7578), .Z(n7610) );
  XNOR U7880 ( .A(n7610), .B(sreg[432]), .Z(n7612) );
  NAND U7881 ( .A(n7571), .B(sreg[431]), .Z(n7575) );
  OR U7882 ( .A(n7573), .B(n7572), .Z(n7574) );
  AND U7883 ( .A(n7575), .B(n7574), .Z(n7611) );
  XOR U7884 ( .A(n7612), .B(n7611), .Z(c[432]) );
  NANDN U7885 ( .A(n7581), .B(n7580), .Z(n7585) );
  NAND U7886 ( .A(n7583), .B(n7582), .Z(n7584) );
  NAND U7887 ( .A(n7585), .B(n7584), .Z(n7646) );
  NANDN U7888 ( .A(n7587), .B(n7586), .Z(n7591) );
  NAND U7889 ( .A(n7589), .B(n7588), .Z(n7590) );
  NAND U7890 ( .A(n7591), .B(n7590), .Z(n7644) );
  XNOR U7891 ( .A(b[7]), .B(a[179]), .Z(n7631) );
  NANDN U7892 ( .A(n7631), .B(n10545), .Z(n7594) );
  NANDN U7893 ( .A(n7592), .B(n10546), .Z(n7593) );
  NAND U7894 ( .A(n7594), .B(n7593), .Z(n7619) );
  XNOR U7895 ( .A(b[3]), .B(a[183]), .Z(n7634) );
  NANDN U7896 ( .A(n7634), .B(n10398), .Z(n7597) );
  NANDN U7897 ( .A(n7595), .B(n10399), .Z(n7596) );
  AND U7898 ( .A(n7597), .B(n7596), .Z(n7620) );
  XNOR U7899 ( .A(n7619), .B(n7620), .Z(n7621) );
  NANDN U7900 ( .A(n527), .B(a[185]), .Z(n7598) );
  XOR U7901 ( .A(n10434), .B(n7598), .Z(n7600) );
  NANDN U7902 ( .A(b[0]), .B(a[184]), .Z(n7599) );
  AND U7903 ( .A(n7600), .B(n7599), .Z(n7627) );
  XOR U7904 ( .A(b[5]), .B(a[181]), .Z(n7640) );
  NAND U7905 ( .A(n7640), .B(n10481), .Z(n7603) );
  NAND U7906 ( .A(n7601), .B(n10482), .Z(n7602) );
  NAND U7907 ( .A(n7603), .B(n7602), .Z(n7625) );
  NANDN U7908 ( .A(n529), .B(a[177]), .Z(n7626) );
  XNOR U7909 ( .A(n7625), .B(n7626), .Z(n7628) );
  XOR U7910 ( .A(n7627), .B(n7628), .Z(n7622) );
  XOR U7911 ( .A(n7621), .B(n7622), .Z(n7643) );
  XOR U7912 ( .A(n7644), .B(n7643), .Z(n7645) );
  XNOR U7913 ( .A(n7646), .B(n7645), .Z(n7615) );
  NAND U7914 ( .A(n7605), .B(n7604), .Z(n7609) );
  NAND U7915 ( .A(n7607), .B(n7606), .Z(n7608) );
  NAND U7916 ( .A(n7609), .B(n7608), .Z(n7616) );
  XNOR U7917 ( .A(n7615), .B(n7616), .Z(n7617) );
  XNOR U7918 ( .A(n7618), .B(n7617), .Z(n7649) );
  XNOR U7919 ( .A(n7649), .B(sreg[433]), .Z(n7651) );
  NAND U7920 ( .A(n7610), .B(sreg[432]), .Z(n7614) );
  OR U7921 ( .A(n7612), .B(n7611), .Z(n7613) );
  AND U7922 ( .A(n7614), .B(n7613), .Z(n7650) );
  XOR U7923 ( .A(n7651), .B(n7650), .Z(c[433]) );
  NANDN U7924 ( .A(n7620), .B(n7619), .Z(n7624) );
  NAND U7925 ( .A(n7622), .B(n7621), .Z(n7623) );
  NAND U7926 ( .A(n7624), .B(n7623), .Z(n7685) );
  NANDN U7927 ( .A(n7626), .B(n7625), .Z(n7630) );
  NAND U7928 ( .A(n7628), .B(n7627), .Z(n7629) );
  NAND U7929 ( .A(n7630), .B(n7629), .Z(n7683) );
  XNOR U7930 ( .A(b[7]), .B(a[180]), .Z(n7670) );
  NANDN U7931 ( .A(n7670), .B(n10545), .Z(n7633) );
  NANDN U7932 ( .A(n7631), .B(n10546), .Z(n7632) );
  NAND U7933 ( .A(n7633), .B(n7632), .Z(n7658) );
  XNOR U7934 ( .A(b[3]), .B(a[184]), .Z(n7673) );
  NANDN U7935 ( .A(n7673), .B(n10398), .Z(n7636) );
  NANDN U7936 ( .A(n7634), .B(n10399), .Z(n7635) );
  AND U7937 ( .A(n7636), .B(n7635), .Z(n7659) );
  XNOR U7938 ( .A(n7658), .B(n7659), .Z(n7660) );
  NANDN U7939 ( .A(n527), .B(a[186]), .Z(n7637) );
  XOR U7940 ( .A(n10434), .B(n7637), .Z(n7639) );
  NANDN U7941 ( .A(b[0]), .B(a[185]), .Z(n7638) );
  AND U7942 ( .A(n7639), .B(n7638), .Z(n7666) );
  XOR U7943 ( .A(b[5]), .B(a[182]), .Z(n7679) );
  NAND U7944 ( .A(n7679), .B(n10481), .Z(n7642) );
  NAND U7945 ( .A(n7640), .B(n10482), .Z(n7641) );
  NAND U7946 ( .A(n7642), .B(n7641), .Z(n7664) );
  NANDN U7947 ( .A(n529), .B(a[178]), .Z(n7665) );
  XNOR U7948 ( .A(n7664), .B(n7665), .Z(n7667) );
  XOR U7949 ( .A(n7666), .B(n7667), .Z(n7661) );
  XOR U7950 ( .A(n7660), .B(n7661), .Z(n7682) );
  XOR U7951 ( .A(n7683), .B(n7682), .Z(n7684) );
  XNOR U7952 ( .A(n7685), .B(n7684), .Z(n7654) );
  NAND U7953 ( .A(n7644), .B(n7643), .Z(n7648) );
  NAND U7954 ( .A(n7646), .B(n7645), .Z(n7647) );
  NAND U7955 ( .A(n7648), .B(n7647), .Z(n7655) );
  XNOR U7956 ( .A(n7654), .B(n7655), .Z(n7656) );
  XNOR U7957 ( .A(n7657), .B(n7656), .Z(n7688) );
  XNOR U7958 ( .A(n7688), .B(sreg[434]), .Z(n7690) );
  NAND U7959 ( .A(n7649), .B(sreg[433]), .Z(n7653) );
  OR U7960 ( .A(n7651), .B(n7650), .Z(n7652) );
  AND U7961 ( .A(n7653), .B(n7652), .Z(n7689) );
  XOR U7962 ( .A(n7690), .B(n7689), .Z(c[434]) );
  NANDN U7963 ( .A(n7659), .B(n7658), .Z(n7663) );
  NAND U7964 ( .A(n7661), .B(n7660), .Z(n7662) );
  NAND U7965 ( .A(n7663), .B(n7662), .Z(n7724) );
  NANDN U7966 ( .A(n7665), .B(n7664), .Z(n7669) );
  NAND U7967 ( .A(n7667), .B(n7666), .Z(n7668) );
  NAND U7968 ( .A(n7669), .B(n7668), .Z(n7722) );
  XNOR U7969 ( .A(b[7]), .B(a[181]), .Z(n7709) );
  NANDN U7970 ( .A(n7709), .B(n10545), .Z(n7672) );
  NANDN U7971 ( .A(n7670), .B(n10546), .Z(n7671) );
  NAND U7972 ( .A(n7672), .B(n7671), .Z(n7697) );
  XNOR U7973 ( .A(b[3]), .B(a[185]), .Z(n7712) );
  NANDN U7974 ( .A(n7712), .B(n10398), .Z(n7675) );
  NANDN U7975 ( .A(n7673), .B(n10399), .Z(n7674) );
  AND U7976 ( .A(n7675), .B(n7674), .Z(n7698) );
  XNOR U7977 ( .A(n7697), .B(n7698), .Z(n7699) );
  NANDN U7978 ( .A(n527), .B(a[187]), .Z(n7676) );
  XOR U7979 ( .A(n10434), .B(n7676), .Z(n7678) );
  NANDN U7980 ( .A(b[0]), .B(a[186]), .Z(n7677) );
  AND U7981 ( .A(n7678), .B(n7677), .Z(n7705) );
  XOR U7982 ( .A(b[5]), .B(a[183]), .Z(n7718) );
  NAND U7983 ( .A(n7718), .B(n10481), .Z(n7681) );
  NAND U7984 ( .A(n7679), .B(n10482), .Z(n7680) );
  NAND U7985 ( .A(n7681), .B(n7680), .Z(n7703) );
  NANDN U7986 ( .A(n529), .B(a[179]), .Z(n7704) );
  XNOR U7987 ( .A(n7703), .B(n7704), .Z(n7706) );
  XOR U7988 ( .A(n7705), .B(n7706), .Z(n7700) );
  XOR U7989 ( .A(n7699), .B(n7700), .Z(n7721) );
  XOR U7990 ( .A(n7722), .B(n7721), .Z(n7723) );
  XNOR U7991 ( .A(n7724), .B(n7723), .Z(n7693) );
  NAND U7992 ( .A(n7683), .B(n7682), .Z(n7687) );
  NAND U7993 ( .A(n7685), .B(n7684), .Z(n7686) );
  NAND U7994 ( .A(n7687), .B(n7686), .Z(n7694) );
  XNOR U7995 ( .A(n7693), .B(n7694), .Z(n7695) );
  XNOR U7996 ( .A(n7696), .B(n7695), .Z(n7727) );
  XNOR U7997 ( .A(n7727), .B(sreg[435]), .Z(n7729) );
  NAND U7998 ( .A(n7688), .B(sreg[434]), .Z(n7692) );
  OR U7999 ( .A(n7690), .B(n7689), .Z(n7691) );
  AND U8000 ( .A(n7692), .B(n7691), .Z(n7728) );
  XOR U8001 ( .A(n7729), .B(n7728), .Z(c[435]) );
  NANDN U8002 ( .A(n7698), .B(n7697), .Z(n7702) );
  NAND U8003 ( .A(n7700), .B(n7699), .Z(n7701) );
  NAND U8004 ( .A(n7702), .B(n7701), .Z(n7763) );
  NANDN U8005 ( .A(n7704), .B(n7703), .Z(n7708) );
  NAND U8006 ( .A(n7706), .B(n7705), .Z(n7707) );
  NAND U8007 ( .A(n7708), .B(n7707), .Z(n7761) );
  XNOR U8008 ( .A(b[7]), .B(a[182]), .Z(n7748) );
  NANDN U8009 ( .A(n7748), .B(n10545), .Z(n7711) );
  NANDN U8010 ( .A(n7709), .B(n10546), .Z(n7710) );
  NAND U8011 ( .A(n7711), .B(n7710), .Z(n7736) );
  XNOR U8012 ( .A(b[3]), .B(a[186]), .Z(n7751) );
  NANDN U8013 ( .A(n7751), .B(n10398), .Z(n7714) );
  NANDN U8014 ( .A(n7712), .B(n10399), .Z(n7713) );
  AND U8015 ( .A(n7714), .B(n7713), .Z(n7737) );
  XNOR U8016 ( .A(n7736), .B(n7737), .Z(n7738) );
  NANDN U8017 ( .A(n527), .B(a[188]), .Z(n7715) );
  XOR U8018 ( .A(n10434), .B(n7715), .Z(n7717) );
  NANDN U8019 ( .A(b[0]), .B(a[187]), .Z(n7716) );
  AND U8020 ( .A(n7717), .B(n7716), .Z(n7744) );
  XOR U8021 ( .A(b[5]), .B(a[184]), .Z(n7757) );
  NAND U8022 ( .A(n7757), .B(n10481), .Z(n7720) );
  NAND U8023 ( .A(n7718), .B(n10482), .Z(n7719) );
  NAND U8024 ( .A(n7720), .B(n7719), .Z(n7742) );
  NANDN U8025 ( .A(n529), .B(a[180]), .Z(n7743) );
  XNOR U8026 ( .A(n7742), .B(n7743), .Z(n7745) );
  XOR U8027 ( .A(n7744), .B(n7745), .Z(n7739) );
  XOR U8028 ( .A(n7738), .B(n7739), .Z(n7760) );
  XOR U8029 ( .A(n7761), .B(n7760), .Z(n7762) );
  XNOR U8030 ( .A(n7763), .B(n7762), .Z(n7732) );
  NAND U8031 ( .A(n7722), .B(n7721), .Z(n7726) );
  NAND U8032 ( .A(n7724), .B(n7723), .Z(n7725) );
  NAND U8033 ( .A(n7726), .B(n7725), .Z(n7733) );
  XNOR U8034 ( .A(n7732), .B(n7733), .Z(n7734) );
  XNOR U8035 ( .A(n7735), .B(n7734), .Z(n7766) );
  XNOR U8036 ( .A(n7766), .B(sreg[436]), .Z(n7768) );
  NAND U8037 ( .A(n7727), .B(sreg[435]), .Z(n7731) );
  OR U8038 ( .A(n7729), .B(n7728), .Z(n7730) );
  AND U8039 ( .A(n7731), .B(n7730), .Z(n7767) );
  XOR U8040 ( .A(n7768), .B(n7767), .Z(c[436]) );
  NANDN U8041 ( .A(n7737), .B(n7736), .Z(n7741) );
  NAND U8042 ( .A(n7739), .B(n7738), .Z(n7740) );
  NAND U8043 ( .A(n7741), .B(n7740), .Z(n7802) );
  NANDN U8044 ( .A(n7743), .B(n7742), .Z(n7747) );
  NAND U8045 ( .A(n7745), .B(n7744), .Z(n7746) );
  NAND U8046 ( .A(n7747), .B(n7746), .Z(n7800) );
  XNOR U8047 ( .A(b[7]), .B(a[183]), .Z(n7787) );
  NANDN U8048 ( .A(n7787), .B(n10545), .Z(n7750) );
  NANDN U8049 ( .A(n7748), .B(n10546), .Z(n7749) );
  NAND U8050 ( .A(n7750), .B(n7749), .Z(n7775) );
  XNOR U8051 ( .A(b[3]), .B(a[187]), .Z(n7790) );
  NANDN U8052 ( .A(n7790), .B(n10398), .Z(n7753) );
  NANDN U8053 ( .A(n7751), .B(n10399), .Z(n7752) );
  AND U8054 ( .A(n7753), .B(n7752), .Z(n7776) );
  XNOR U8055 ( .A(n7775), .B(n7776), .Z(n7777) );
  NANDN U8056 ( .A(n527), .B(a[189]), .Z(n7754) );
  XOR U8057 ( .A(n10434), .B(n7754), .Z(n7756) );
  NANDN U8058 ( .A(b[0]), .B(a[188]), .Z(n7755) );
  AND U8059 ( .A(n7756), .B(n7755), .Z(n7783) );
  XOR U8060 ( .A(b[5]), .B(a[185]), .Z(n7796) );
  NAND U8061 ( .A(n7796), .B(n10481), .Z(n7759) );
  NAND U8062 ( .A(n7757), .B(n10482), .Z(n7758) );
  NAND U8063 ( .A(n7759), .B(n7758), .Z(n7781) );
  NANDN U8064 ( .A(n529), .B(a[181]), .Z(n7782) );
  XNOR U8065 ( .A(n7781), .B(n7782), .Z(n7784) );
  XOR U8066 ( .A(n7783), .B(n7784), .Z(n7778) );
  XOR U8067 ( .A(n7777), .B(n7778), .Z(n7799) );
  XOR U8068 ( .A(n7800), .B(n7799), .Z(n7801) );
  XNOR U8069 ( .A(n7802), .B(n7801), .Z(n7771) );
  NAND U8070 ( .A(n7761), .B(n7760), .Z(n7765) );
  NAND U8071 ( .A(n7763), .B(n7762), .Z(n7764) );
  NAND U8072 ( .A(n7765), .B(n7764), .Z(n7772) );
  XNOR U8073 ( .A(n7771), .B(n7772), .Z(n7773) );
  XNOR U8074 ( .A(n7774), .B(n7773), .Z(n7805) );
  XNOR U8075 ( .A(n7805), .B(sreg[437]), .Z(n7807) );
  NAND U8076 ( .A(n7766), .B(sreg[436]), .Z(n7770) );
  OR U8077 ( .A(n7768), .B(n7767), .Z(n7769) );
  AND U8078 ( .A(n7770), .B(n7769), .Z(n7806) );
  XOR U8079 ( .A(n7807), .B(n7806), .Z(c[437]) );
  NANDN U8080 ( .A(n7776), .B(n7775), .Z(n7780) );
  NAND U8081 ( .A(n7778), .B(n7777), .Z(n7779) );
  NAND U8082 ( .A(n7780), .B(n7779), .Z(n7841) );
  NANDN U8083 ( .A(n7782), .B(n7781), .Z(n7786) );
  NAND U8084 ( .A(n7784), .B(n7783), .Z(n7785) );
  NAND U8085 ( .A(n7786), .B(n7785), .Z(n7839) );
  XNOR U8086 ( .A(b[7]), .B(a[184]), .Z(n7832) );
  NANDN U8087 ( .A(n7832), .B(n10545), .Z(n7789) );
  NANDN U8088 ( .A(n7787), .B(n10546), .Z(n7788) );
  NAND U8089 ( .A(n7789), .B(n7788), .Z(n7814) );
  XNOR U8090 ( .A(b[3]), .B(a[188]), .Z(n7835) );
  NANDN U8091 ( .A(n7835), .B(n10398), .Z(n7792) );
  NANDN U8092 ( .A(n7790), .B(n10399), .Z(n7791) );
  AND U8093 ( .A(n7792), .B(n7791), .Z(n7815) );
  XNOR U8094 ( .A(n7814), .B(n7815), .Z(n7816) );
  NANDN U8095 ( .A(n527), .B(a[190]), .Z(n7793) );
  XOR U8096 ( .A(n10434), .B(n7793), .Z(n7795) );
  NANDN U8097 ( .A(b[0]), .B(a[189]), .Z(n7794) );
  AND U8098 ( .A(n7795), .B(n7794), .Z(n7822) );
  XOR U8099 ( .A(b[5]), .B(a[186]), .Z(n7829) );
  NAND U8100 ( .A(n7829), .B(n10481), .Z(n7798) );
  NAND U8101 ( .A(n7796), .B(n10482), .Z(n7797) );
  NAND U8102 ( .A(n7798), .B(n7797), .Z(n7820) );
  NANDN U8103 ( .A(n529), .B(a[182]), .Z(n7821) );
  XNOR U8104 ( .A(n7820), .B(n7821), .Z(n7823) );
  XOR U8105 ( .A(n7822), .B(n7823), .Z(n7817) );
  XOR U8106 ( .A(n7816), .B(n7817), .Z(n7838) );
  XOR U8107 ( .A(n7839), .B(n7838), .Z(n7840) );
  XNOR U8108 ( .A(n7841), .B(n7840), .Z(n7810) );
  NAND U8109 ( .A(n7800), .B(n7799), .Z(n7804) );
  NAND U8110 ( .A(n7802), .B(n7801), .Z(n7803) );
  NAND U8111 ( .A(n7804), .B(n7803), .Z(n7811) );
  XNOR U8112 ( .A(n7810), .B(n7811), .Z(n7812) );
  XNOR U8113 ( .A(n7813), .B(n7812), .Z(n7844) );
  XNOR U8114 ( .A(n7844), .B(sreg[438]), .Z(n7846) );
  NAND U8115 ( .A(n7805), .B(sreg[437]), .Z(n7809) );
  OR U8116 ( .A(n7807), .B(n7806), .Z(n7808) );
  AND U8117 ( .A(n7809), .B(n7808), .Z(n7845) );
  XOR U8118 ( .A(n7846), .B(n7845), .Z(c[438]) );
  NANDN U8119 ( .A(n7815), .B(n7814), .Z(n7819) );
  NAND U8120 ( .A(n7817), .B(n7816), .Z(n7818) );
  NAND U8121 ( .A(n7819), .B(n7818), .Z(n7880) );
  NANDN U8122 ( .A(n7821), .B(n7820), .Z(n7825) );
  NAND U8123 ( .A(n7823), .B(n7822), .Z(n7824) );
  NAND U8124 ( .A(n7825), .B(n7824), .Z(n7878) );
  NANDN U8125 ( .A(n527), .B(a[191]), .Z(n7826) );
  XOR U8126 ( .A(n10434), .B(n7826), .Z(n7828) );
  NANDN U8127 ( .A(b[0]), .B(a[190]), .Z(n7827) );
  AND U8128 ( .A(n7828), .B(n7827), .Z(n7861) );
  XOR U8129 ( .A(b[5]), .B(a[187]), .Z(n7874) );
  NAND U8130 ( .A(n7874), .B(n10481), .Z(n7831) );
  NAND U8131 ( .A(n7829), .B(n10482), .Z(n7830) );
  NAND U8132 ( .A(n7831), .B(n7830), .Z(n7859) );
  NANDN U8133 ( .A(n529), .B(a[183]), .Z(n7860) );
  XNOR U8134 ( .A(n7859), .B(n7860), .Z(n7862) );
  XOR U8135 ( .A(n7861), .B(n7862), .Z(n7855) );
  XNOR U8136 ( .A(b[7]), .B(a[185]), .Z(n7865) );
  NANDN U8137 ( .A(n7865), .B(n10545), .Z(n7834) );
  NANDN U8138 ( .A(n7832), .B(n10546), .Z(n7833) );
  NAND U8139 ( .A(n7834), .B(n7833), .Z(n7853) );
  XNOR U8140 ( .A(b[3]), .B(a[189]), .Z(n7868) );
  NANDN U8141 ( .A(n7868), .B(n10398), .Z(n7837) );
  NANDN U8142 ( .A(n7835), .B(n10399), .Z(n7836) );
  AND U8143 ( .A(n7837), .B(n7836), .Z(n7854) );
  XNOR U8144 ( .A(n7853), .B(n7854), .Z(n7856) );
  XOR U8145 ( .A(n7855), .B(n7856), .Z(n7877) );
  XOR U8146 ( .A(n7878), .B(n7877), .Z(n7879) );
  XNOR U8147 ( .A(n7880), .B(n7879), .Z(n7849) );
  NAND U8148 ( .A(n7839), .B(n7838), .Z(n7843) );
  NAND U8149 ( .A(n7841), .B(n7840), .Z(n7842) );
  NAND U8150 ( .A(n7843), .B(n7842), .Z(n7850) );
  XNOR U8151 ( .A(n7849), .B(n7850), .Z(n7851) );
  XNOR U8152 ( .A(n7852), .B(n7851), .Z(n7883) );
  XNOR U8153 ( .A(n7883), .B(sreg[439]), .Z(n7885) );
  NAND U8154 ( .A(n7844), .B(sreg[438]), .Z(n7848) );
  OR U8155 ( .A(n7846), .B(n7845), .Z(n7847) );
  AND U8156 ( .A(n7848), .B(n7847), .Z(n7884) );
  XOR U8157 ( .A(n7885), .B(n7884), .Z(c[439]) );
  NANDN U8158 ( .A(n7854), .B(n7853), .Z(n7858) );
  NAND U8159 ( .A(n7856), .B(n7855), .Z(n7857) );
  NAND U8160 ( .A(n7858), .B(n7857), .Z(n7919) );
  NANDN U8161 ( .A(n7860), .B(n7859), .Z(n7864) );
  NAND U8162 ( .A(n7862), .B(n7861), .Z(n7863) );
  NAND U8163 ( .A(n7864), .B(n7863), .Z(n7917) );
  XNOR U8164 ( .A(b[7]), .B(a[186]), .Z(n7904) );
  NANDN U8165 ( .A(n7904), .B(n10545), .Z(n7867) );
  NANDN U8166 ( .A(n7865), .B(n10546), .Z(n7866) );
  NAND U8167 ( .A(n7867), .B(n7866), .Z(n7892) );
  XNOR U8168 ( .A(b[3]), .B(a[190]), .Z(n7907) );
  NANDN U8169 ( .A(n7907), .B(n10398), .Z(n7870) );
  NANDN U8170 ( .A(n7868), .B(n10399), .Z(n7869) );
  AND U8171 ( .A(n7870), .B(n7869), .Z(n7893) );
  XNOR U8172 ( .A(n7892), .B(n7893), .Z(n7894) );
  NANDN U8173 ( .A(n527), .B(a[192]), .Z(n7871) );
  XOR U8174 ( .A(n10434), .B(n7871), .Z(n7873) );
  NANDN U8175 ( .A(b[0]), .B(a[191]), .Z(n7872) );
  AND U8176 ( .A(n7873), .B(n7872), .Z(n7900) );
  XOR U8177 ( .A(b[5]), .B(a[188]), .Z(n7913) );
  NAND U8178 ( .A(n7913), .B(n10481), .Z(n7876) );
  NAND U8179 ( .A(n7874), .B(n10482), .Z(n7875) );
  NAND U8180 ( .A(n7876), .B(n7875), .Z(n7898) );
  NANDN U8181 ( .A(n529), .B(a[184]), .Z(n7899) );
  XNOR U8182 ( .A(n7898), .B(n7899), .Z(n7901) );
  XOR U8183 ( .A(n7900), .B(n7901), .Z(n7895) );
  XOR U8184 ( .A(n7894), .B(n7895), .Z(n7916) );
  XOR U8185 ( .A(n7917), .B(n7916), .Z(n7918) );
  XNOR U8186 ( .A(n7919), .B(n7918), .Z(n7888) );
  NAND U8187 ( .A(n7878), .B(n7877), .Z(n7882) );
  NAND U8188 ( .A(n7880), .B(n7879), .Z(n7881) );
  NAND U8189 ( .A(n7882), .B(n7881), .Z(n7889) );
  XNOR U8190 ( .A(n7888), .B(n7889), .Z(n7890) );
  XNOR U8191 ( .A(n7891), .B(n7890), .Z(n7922) );
  XNOR U8192 ( .A(n7922), .B(sreg[440]), .Z(n7924) );
  NAND U8193 ( .A(n7883), .B(sreg[439]), .Z(n7887) );
  OR U8194 ( .A(n7885), .B(n7884), .Z(n7886) );
  AND U8195 ( .A(n7887), .B(n7886), .Z(n7923) );
  XOR U8196 ( .A(n7924), .B(n7923), .Z(c[440]) );
  NANDN U8197 ( .A(n7893), .B(n7892), .Z(n7897) );
  NAND U8198 ( .A(n7895), .B(n7894), .Z(n7896) );
  NAND U8199 ( .A(n7897), .B(n7896), .Z(n7958) );
  NANDN U8200 ( .A(n7899), .B(n7898), .Z(n7903) );
  NAND U8201 ( .A(n7901), .B(n7900), .Z(n7902) );
  NAND U8202 ( .A(n7903), .B(n7902), .Z(n7956) );
  XNOR U8203 ( .A(b[7]), .B(a[187]), .Z(n7943) );
  NANDN U8204 ( .A(n7943), .B(n10545), .Z(n7906) );
  NANDN U8205 ( .A(n7904), .B(n10546), .Z(n7905) );
  NAND U8206 ( .A(n7906), .B(n7905), .Z(n7931) );
  XNOR U8207 ( .A(b[3]), .B(a[191]), .Z(n7946) );
  NANDN U8208 ( .A(n7946), .B(n10398), .Z(n7909) );
  NANDN U8209 ( .A(n7907), .B(n10399), .Z(n7908) );
  AND U8210 ( .A(n7909), .B(n7908), .Z(n7932) );
  XNOR U8211 ( .A(n7931), .B(n7932), .Z(n7933) );
  NANDN U8212 ( .A(n527), .B(a[193]), .Z(n7910) );
  XOR U8213 ( .A(n10434), .B(n7910), .Z(n7912) );
  NANDN U8214 ( .A(b[0]), .B(a[192]), .Z(n7911) );
  AND U8215 ( .A(n7912), .B(n7911), .Z(n7939) );
  XOR U8216 ( .A(b[5]), .B(a[189]), .Z(n7952) );
  NAND U8217 ( .A(n7952), .B(n10481), .Z(n7915) );
  NAND U8218 ( .A(n7913), .B(n10482), .Z(n7914) );
  NAND U8219 ( .A(n7915), .B(n7914), .Z(n7937) );
  NANDN U8220 ( .A(n529), .B(a[185]), .Z(n7938) );
  XNOR U8221 ( .A(n7937), .B(n7938), .Z(n7940) );
  XOR U8222 ( .A(n7939), .B(n7940), .Z(n7934) );
  XOR U8223 ( .A(n7933), .B(n7934), .Z(n7955) );
  XOR U8224 ( .A(n7956), .B(n7955), .Z(n7957) );
  XNOR U8225 ( .A(n7958), .B(n7957), .Z(n7927) );
  NAND U8226 ( .A(n7917), .B(n7916), .Z(n7921) );
  NAND U8227 ( .A(n7919), .B(n7918), .Z(n7920) );
  NAND U8228 ( .A(n7921), .B(n7920), .Z(n7928) );
  XNOR U8229 ( .A(n7927), .B(n7928), .Z(n7929) );
  XNOR U8230 ( .A(n7930), .B(n7929), .Z(n7961) );
  XNOR U8231 ( .A(n7961), .B(sreg[441]), .Z(n7963) );
  NAND U8232 ( .A(n7922), .B(sreg[440]), .Z(n7926) );
  OR U8233 ( .A(n7924), .B(n7923), .Z(n7925) );
  AND U8234 ( .A(n7926), .B(n7925), .Z(n7962) );
  XOR U8235 ( .A(n7963), .B(n7962), .Z(c[441]) );
  NANDN U8236 ( .A(n7932), .B(n7931), .Z(n7936) );
  NAND U8237 ( .A(n7934), .B(n7933), .Z(n7935) );
  NAND U8238 ( .A(n7936), .B(n7935), .Z(n7997) );
  NANDN U8239 ( .A(n7938), .B(n7937), .Z(n7942) );
  NAND U8240 ( .A(n7940), .B(n7939), .Z(n7941) );
  NAND U8241 ( .A(n7942), .B(n7941), .Z(n7995) );
  XNOR U8242 ( .A(b[7]), .B(a[188]), .Z(n7988) );
  NANDN U8243 ( .A(n7988), .B(n10545), .Z(n7945) );
  NANDN U8244 ( .A(n7943), .B(n10546), .Z(n7944) );
  NAND U8245 ( .A(n7945), .B(n7944), .Z(n7970) );
  XNOR U8246 ( .A(b[3]), .B(a[192]), .Z(n7991) );
  NANDN U8247 ( .A(n7991), .B(n10398), .Z(n7948) );
  NANDN U8248 ( .A(n7946), .B(n10399), .Z(n7947) );
  AND U8249 ( .A(n7948), .B(n7947), .Z(n7971) );
  XNOR U8250 ( .A(n7970), .B(n7971), .Z(n7972) );
  NANDN U8251 ( .A(n527), .B(a[194]), .Z(n7949) );
  XOR U8252 ( .A(n10434), .B(n7949), .Z(n7951) );
  NANDN U8253 ( .A(b[0]), .B(a[193]), .Z(n7950) );
  AND U8254 ( .A(n7951), .B(n7950), .Z(n7978) );
  XOR U8255 ( .A(b[5]), .B(a[190]), .Z(n7985) );
  NAND U8256 ( .A(n7985), .B(n10481), .Z(n7954) );
  NAND U8257 ( .A(n7952), .B(n10482), .Z(n7953) );
  NAND U8258 ( .A(n7954), .B(n7953), .Z(n7976) );
  NANDN U8259 ( .A(n529), .B(a[186]), .Z(n7977) );
  XNOR U8260 ( .A(n7976), .B(n7977), .Z(n7979) );
  XOR U8261 ( .A(n7978), .B(n7979), .Z(n7973) );
  XOR U8262 ( .A(n7972), .B(n7973), .Z(n7994) );
  XOR U8263 ( .A(n7995), .B(n7994), .Z(n7996) );
  XNOR U8264 ( .A(n7997), .B(n7996), .Z(n7966) );
  NAND U8265 ( .A(n7956), .B(n7955), .Z(n7960) );
  NAND U8266 ( .A(n7958), .B(n7957), .Z(n7959) );
  NAND U8267 ( .A(n7960), .B(n7959), .Z(n7967) );
  XNOR U8268 ( .A(n7966), .B(n7967), .Z(n7968) );
  XNOR U8269 ( .A(n7969), .B(n7968), .Z(n8000) );
  XNOR U8270 ( .A(n8000), .B(sreg[442]), .Z(n8002) );
  NAND U8271 ( .A(n7961), .B(sreg[441]), .Z(n7965) );
  OR U8272 ( .A(n7963), .B(n7962), .Z(n7964) );
  AND U8273 ( .A(n7965), .B(n7964), .Z(n8001) );
  XOR U8274 ( .A(n8002), .B(n8001), .Z(c[442]) );
  NANDN U8275 ( .A(n7971), .B(n7970), .Z(n7975) );
  NAND U8276 ( .A(n7973), .B(n7972), .Z(n7974) );
  NAND U8277 ( .A(n7975), .B(n7974), .Z(n8036) );
  NANDN U8278 ( .A(n7977), .B(n7976), .Z(n7981) );
  NAND U8279 ( .A(n7979), .B(n7978), .Z(n7980) );
  NAND U8280 ( .A(n7981), .B(n7980), .Z(n8034) );
  NANDN U8281 ( .A(n527), .B(a[195]), .Z(n7982) );
  XOR U8282 ( .A(n10434), .B(n7982), .Z(n7984) );
  NANDN U8283 ( .A(b[0]), .B(a[194]), .Z(n7983) );
  AND U8284 ( .A(n7984), .B(n7983), .Z(n8017) );
  XOR U8285 ( .A(b[5]), .B(a[191]), .Z(n8030) );
  NAND U8286 ( .A(n8030), .B(n10481), .Z(n7987) );
  NAND U8287 ( .A(n7985), .B(n10482), .Z(n7986) );
  NAND U8288 ( .A(n7987), .B(n7986), .Z(n8015) );
  NANDN U8289 ( .A(n529), .B(a[187]), .Z(n8016) );
  XNOR U8290 ( .A(n8015), .B(n8016), .Z(n8018) );
  XOR U8291 ( .A(n8017), .B(n8018), .Z(n8011) );
  XNOR U8292 ( .A(b[7]), .B(a[189]), .Z(n8021) );
  NANDN U8293 ( .A(n8021), .B(n10545), .Z(n7990) );
  NANDN U8294 ( .A(n7988), .B(n10546), .Z(n7989) );
  NAND U8295 ( .A(n7990), .B(n7989), .Z(n8009) );
  XNOR U8296 ( .A(b[3]), .B(a[193]), .Z(n8024) );
  NANDN U8297 ( .A(n8024), .B(n10398), .Z(n7993) );
  NANDN U8298 ( .A(n7991), .B(n10399), .Z(n7992) );
  AND U8299 ( .A(n7993), .B(n7992), .Z(n8010) );
  XNOR U8300 ( .A(n8009), .B(n8010), .Z(n8012) );
  XOR U8301 ( .A(n8011), .B(n8012), .Z(n8033) );
  XOR U8302 ( .A(n8034), .B(n8033), .Z(n8035) );
  XNOR U8303 ( .A(n8036), .B(n8035), .Z(n8005) );
  NAND U8304 ( .A(n7995), .B(n7994), .Z(n7999) );
  NAND U8305 ( .A(n7997), .B(n7996), .Z(n7998) );
  NAND U8306 ( .A(n7999), .B(n7998), .Z(n8006) );
  XNOR U8307 ( .A(n8005), .B(n8006), .Z(n8007) );
  XNOR U8308 ( .A(n8008), .B(n8007), .Z(n8039) );
  XNOR U8309 ( .A(n8039), .B(sreg[443]), .Z(n8041) );
  NAND U8310 ( .A(n8000), .B(sreg[442]), .Z(n8004) );
  OR U8311 ( .A(n8002), .B(n8001), .Z(n8003) );
  AND U8312 ( .A(n8004), .B(n8003), .Z(n8040) );
  XOR U8313 ( .A(n8041), .B(n8040), .Z(c[443]) );
  NANDN U8314 ( .A(n8010), .B(n8009), .Z(n8014) );
  NAND U8315 ( .A(n8012), .B(n8011), .Z(n8013) );
  NAND U8316 ( .A(n8014), .B(n8013), .Z(n8075) );
  NANDN U8317 ( .A(n8016), .B(n8015), .Z(n8020) );
  NAND U8318 ( .A(n8018), .B(n8017), .Z(n8019) );
  NAND U8319 ( .A(n8020), .B(n8019), .Z(n8073) );
  XNOR U8320 ( .A(b[7]), .B(a[190]), .Z(n8060) );
  NANDN U8321 ( .A(n8060), .B(n10545), .Z(n8023) );
  NANDN U8322 ( .A(n8021), .B(n10546), .Z(n8022) );
  NAND U8323 ( .A(n8023), .B(n8022), .Z(n8048) );
  XNOR U8324 ( .A(b[3]), .B(a[194]), .Z(n8063) );
  NANDN U8325 ( .A(n8063), .B(n10398), .Z(n8026) );
  NANDN U8326 ( .A(n8024), .B(n10399), .Z(n8025) );
  AND U8327 ( .A(n8026), .B(n8025), .Z(n8049) );
  XNOR U8328 ( .A(n8048), .B(n8049), .Z(n8050) );
  NANDN U8329 ( .A(n527), .B(a[196]), .Z(n8027) );
  XOR U8330 ( .A(n10434), .B(n8027), .Z(n8029) );
  NANDN U8331 ( .A(b[0]), .B(a[195]), .Z(n8028) );
  AND U8332 ( .A(n8029), .B(n8028), .Z(n8056) );
  XOR U8333 ( .A(b[5]), .B(a[192]), .Z(n8069) );
  NAND U8334 ( .A(n8069), .B(n10481), .Z(n8032) );
  NAND U8335 ( .A(n8030), .B(n10482), .Z(n8031) );
  NAND U8336 ( .A(n8032), .B(n8031), .Z(n8054) );
  NANDN U8337 ( .A(n529), .B(a[188]), .Z(n8055) );
  XNOR U8338 ( .A(n8054), .B(n8055), .Z(n8057) );
  XOR U8339 ( .A(n8056), .B(n8057), .Z(n8051) );
  XOR U8340 ( .A(n8050), .B(n8051), .Z(n8072) );
  XOR U8341 ( .A(n8073), .B(n8072), .Z(n8074) );
  XNOR U8342 ( .A(n8075), .B(n8074), .Z(n8044) );
  NAND U8343 ( .A(n8034), .B(n8033), .Z(n8038) );
  NAND U8344 ( .A(n8036), .B(n8035), .Z(n8037) );
  NAND U8345 ( .A(n8038), .B(n8037), .Z(n8045) );
  XNOR U8346 ( .A(n8044), .B(n8045), .Z(n8046) );
  XNOR U8347 ( .A(n8047), .B(n8046), .Z(n8078) );
  XNOR U8348 ( .A(n8078), .B(sreg[444]), .Z(n8080) );
  NAND U8349 ( .A(n8039), .B(sreg[443]), .Z(n8043) );
  OR U8350 ( .A(n8041), .B(n8040), .Z(n8042) );
  AND U8351 ( .A(n8043), .B(n8042), .Z(n8079) );
  XOR U8352 ( .A(n8080), .B(n8079), .Z(c[444]) );
  NANDN U8353 ( .A(n8049), .B(n8048), .Z(n8053) );
  NAND U8354 ( .A(n8051), .B(n8050), .Z(n8052) );
  NAND U8355 ( .A(n8053), .B(n8052), .Z(n8114) );
  NANDN U8356 ( .A(n8055), .B(n8054), .Z(n8059) );
  NAND U8357 ( .A(n8057), .B(n8056), .Z(n8058) );
  NAND U8358 ( .A(n8059), .B(n8058), .Z(n8112) );
  XNOR U8359 ( .A(b[7]), .B(a[191]), .Z(n8099) );
  NANDN U8360 ( .A(n8099), .B(n10545), .Z(n8062) );
  NANDN U8361 ( .A(n8060), .B(n10546), .Z(n8061) );
  NAND U8362 ( .A(n8062), .B(n8061), .Z(n8087) );
  XNOR U8363 ( .A(b[3]), .B(a[195]), .Z(n8102) );
  NANDN U8364 ( .A(n8102), .B(n10398), .Z(n8065) );
  NANDN U8365 ( .A(n8063), .B(n10399), .Z(n8064) );
  AND U8366 ( .A(n8065), .B(n8064), .Z(n8088) );
  XNOR U8367 ( .A(n8087), .B(n8088), .Z(n8089) );
  NANDN U8368 ( .A(n527), .B(a[197]), .Z(n8066) );
  XOR U8369 ( .A(n10434), .B(n8066), .Z(n8068) );
  NANDN U8370 ( .A(b[0]), .B(a[196]), .Z(n8067) );
  AND U8371 ( .A(n8068), .B(n8067), .Z(n8095) );
  XOR U8372 ( .A(b[5]), .B(a[193]), .Z(n8108) );
  NAND U8373 ( .A(n8108), .B(n10481), .Z(n8071) );
  NAND U8374 ( .A(n8069), .B(n10482), .Z(n8070) );
  NAND U8375 ( .A(n8071), .B(n8070), .Z(n8093) );
  NANDN U8376 ( .A(n529), .B(a[189]), .Z(n8094) );
  XNOR U8377 ( .A(n8093), .B(n8094), .Z(n8096) );
  XOR U8378 ( .A(n8095), .B(n8096), .Z(n8090) );
  XOR U8379 ( .A(n8089), .B(n8090), .Z(n8111) );
  XOR U8380 ( .A(n8112), .B(n8111), .Z(n8113) );
  XNOR U8381 ( .A(n8114), .B(n8113), .Z(n8083) );
  NAND U8382 ( .A(n8073), .B(n8072), .Z(n8077) );
  NAND U8383 ( .A(n8075), .B(n8074), .Z(n8076) );
  NAND U8384 ( .A(n8077), .B(n8076), .Z(n8084) );
  XNOR U8385 ( .A(n8083), .B(n8084), .Z(n8085) );
  XNOR U8386 ( .A(n8086), .B(n8085), .Z(n8117) );
  XNOR U8387 ( .A(n8117), .B(sreg[445]), .Z(n8119) );
  NAND U8388 ( .A(n8078), .B(sreg[444]), .Z(n8082) );
  OR U8389 ( .A(n8080), .B(n8079), .Z(n8081) );
  AND U8390 ( .A(n8082), .B(n8081), .Z(n8118) );
  XOR U8391 ( .A(n8119), .B(n8118), .Z(c[445]) );
  NANDN U8392 ( .A(n8088), .B(n8087), .Z(n8092) );
  NAND U8393 ( .A(n8090), .B(n8089), .Z(n8091) );
  NAND U8394 ( .A(n8092), .B(n8091), .Z(n8153) );
  NANDN U8395 ( .A(n8094), .B(n8093), .Z(n8098) );
  NAND U8396 ( .A(n8096), .B(n8095), .Z(n8097) );
  NAND U8397 ( .A(n8098), .B(n8097), .Z(n8151) );
  XNOR U8398 ( .A(b[7]), .B(a[192]), .Z(n8138) );
  NANDN U8399 ( .A(n8138), .B(n10545), .Z(n8101) );
  NANDN U8400 ( .A(n8099), .B(n10546), .Z(n8100) );
  NAND U8401 ( .A(n8101), .B(n8100), .Z(n8126) );
  XNOR U8402 ( .A(b[3]), .B(a[196]), .Z(n8141) );
  NANDN U8403 ( .A(n8141), .B(n10398), .Z(n8104) );
  NANDN U8404 ( .A(n8102), .B(n10399), .Z(n8103) );
  AND U8405 ( .A(n8104), .B(n8103), .Z(n8127) );
  XNOR U8406 ( .A(n8126), .B(n8127), .Z(n8128) );
  NANDN U8407 ( .A(n527), .B(a[198]), .Z(n8105) );
  XOR U8408 ( .A(n10434), .B(n8105), .Z(n8107) );
  NANDN U8409 ( .A(b[0]), .B(a[197]), .Z(n8106) );
  AND U8410 ( .A(n8107), .B(n8106), .Z(n8134) );
  XOR U8411 ( .A(b[5]), .B(a[194]), .Z(n8147) );
  NAND U8412 ( .A(n8147), .B(n10481), .Z(n8110) );
  NAND U8413 ( .A(n8108), .B(n10482), .Z(n8109) );
  NAND U8414 ( .A(n8110), .B(n8109), .Z(n8132) );
  NANDN U8415 ( .A(n529), .B(a[190]), .Z(n8133) );
  XNOR U8416 ( .A(n8132), .B(n8133), .Z(n8135) );
  XOR U8417 ( .A(n8134), .B(n8135), .Z(n8129) );
  XOR U8418 ( .A(n8128), .B(n8129), .Z(n8150) );
  XOR U8419 ( .A(n8151), .B(n8150), .Z(n8152) );
  XNOR U8420 ( .A(n8153), .B(n8152), .Z(n8122) );
  NAND U8421 ( .A(n8112), .B(n8111), .Z(n8116) );
  NAND U8422 ( .A(n8114), .B(n8113), .Z(n8115) );
  NAND U8423 ( .A(n8116), .B(n8115), .Z(n8123) );
  XNOR U8424 ( .A(n8122), .B(n8123), .Z(n8124) );
  XNOR U8425 ( .A(n8125), .B(n8124), .Z(n8156) );
  XNOR U8426 ( .A(n8156), .B(sreg[446]), .Z(n8158) );
  NAND U8427 ( .A(n8117), .B(sreg[445]), .Z(n8121) );
  OR U8428 ( .A(n8119), .B(n8118), .Z(n8120) );
  AND U8429 ( .A(n8121), .B(n8120), .Z(n8157) );
  XOR U8430 ( .A(n8158), .B(n8157), .Z(c[446]) );
  NANDN U8431 ( .A(n8127), .B(n8126), .Z(n8131) );
  NAND U8432 ( .A(n8129), .B(n8128), .Z(n8130) );
  NAND U8433 ( .A(n8131), .B(n8130), .Z(n8192) );
  NANDN U8434 ( .A(n8133), .B(n8132), .Z(n8137) );
  NAND U8435 ( .A(n8135), .B(n8134), .Z(n8136) );
  NAND U8436 ( .A(n8137), .B(n8136), .Z(n8190) );
  XNOR U8437 ( .A(b[7]), .B(a[193]), .Z(n8177) );
  NANDN U8438 ( .A(n8177), .B(n10545), .Z(n8140) );
  NANDN U8439 ( .A(n8138), .B(n10546), .Z(n8139) );
  NAND U8440 ( .A(n8140), .B(n8139), .Z(n8165) );
  XNOR U8441 ( .A(b[3]), .B(a[197]), .Z(n8180) );
  NANDN U8442 ( .A(n8180), .B(n10398), .Z(n8143) );
  NANDN U8443 ( .A(n8141), .B(n10399), .Z(n8142) );
  AND U8444 ( .A(n8143), .B(n8142), .Z(n8166) );
  XNOR U8445 ( .A(n8165), .B(n8166), .Z(n8167) );
  NANDN U8446 ( .A(n527), .B(a[199]), .Z(n8144) );
  XOR U8447 ( .A(n10434), .B(n8144), .Z(n8146) );
  NANDN U8448 ( .A(b[0]), .B(a[198]), .Z(n8145) );
  AND U8449 ( .A(n8146), .B(n8145), .Z(n8173) );
  XOR U8450 ( .A(b[5]), .B(a[195]), .Z(n8186) );
  NAND U8451 ( .A(n8186), .B(n10481), .Z(n8149) );
  NAND U8452 ( .A(n8147), .B(n10482), .Z(n8148) );
  NAND U8453 ( .A(n8149), .B(n8148), .Z(n8171) );
  NANDN U8454 ( .A(n529), .B(a[191]), .Z(n8172) );
  XNOR U8455 ( .A(n8171), .B(n8172), .Z(n8174) );
  XOR U8456 ( .A(n8173), .B(n8174), .Z(n8168) );
  XOR U8457 ( .A(n8167), .B(n8168), .Z(n8189) );
  XOR U8458 ( .A(n8190), .B(n8189), .Z(n8191) );
  XNOR U8459 ( .A(n8192), .B(n8191), .Z(n8161) );
  NAND U8460 ( .A(n8151), .B(n8150), .Z(n8155) );
  NAND U8461 ( .A(n8153), .B(n8152), .Z(n8154) );
  NAND U8462 ( .A(n8155), .B(n8154), .Z(n8162) );
  XNOR U8463 ( .A(n8161), .B(n8162), .Z(n8163) );
  XNOR U8464 ( .A(n8164), .B(n8163), .Z(n8195) );
  XNOR U8465 ( .A(n8195), .B(sreg[447]), .Z(n8197) );
  NAND U8466 ( .A(n8156), .B(sreg[446]), .Z(n8160) );
  OR U8467 ( .A(n8158), .B(n8157), .Z(n8159) );
  AND U8468 ( .A(n8160), .B(n8159), .Z(n8196) );
  XOR U8469 ( .A(n8197), .B(n8196), .Z(c[447]) );
  NANDN U8470 ( .A(n8166), .B(n8165), .Z(n8170) );
  NAND U8471 ( .A(n8168), .B(n8167), .Z(n8169) );
  NAND U8472 ( .A(n8170), .B(n8169), .Z(n8231) );
  NANDN U8473 ( .A(n8172), .B(n8171), .Z(n8176) );
  NAND U8474 ( .A(n8174), .B(n8173), .Z(n8175) );
  NAND U8475 ( .A(n8176), .B(n8175), .Z(n8229) );
  XNOR U8476 ( .A(b[7]), .B(a[194]), .Z(n8216) );
  NANDN U8477 ( .A(n8216), .B(n10545), .Z(n8179) );
  NANDN U8478 ( .A(n8177), .B(n10546), .Z(n8178) );
  NAND U8479 ( .A(n8179), .B(n8178), .Z(n8204) );
  XNOR U8480 ( .A(b[3]), .B(a[198]), .Z(n8219) );
  NANDN U8481 ( .A(n8219), .B(n10398), .Z(n8182) );
  NANDN U8482 ( .A(n8180), .B(n10399), .Z(n8181) );
  AND U8483 ( .A(n8182), .B(n8181), .Z(n8205) );
  XNOR U8484 ( .A(n8204), .B(n8205), .Z(n8206) );
  NANDN U8485 ( .A(n527), .B(a[200]), .Z(n8183) );
  XOR U8486 ( .A(n10434), .B(n8183), .Z(n8185) );
  NANDN U8487 ( .A(b[0]), .B(a[199]), .Z(n8184) );
  AND U8488 ( .A(n8185), .B(n8184), .Z(n8212) );
  XOR U8489 ( .A(b[5]), .B(a[196]), .Z(n8225) );
  NAND U8490 ( .A(n8225), .B(n10481), .Z(n8188) );
  NAND U8491 ( .A(n8186), .B(n10482), .Z(n8187) );
  NAND U8492 ( .A(n8188), .B(n8187), .Z(n8210) );
  NANDN U8493 ( .A(n529), .B(a[192]), .Z(n8211) );
  XNOR U8494 ( .A(n8210), .B(n8211), .Z(n8213) );
  XOR U8495 ( .A(n8212), .B(n8213), .Z(n8207) );
  XOR U8496 ( .A(n8206), .B(n8207), .Z(n8228) );
  XOR U8497 ( .A(n8229), .B(n8228), .Z(n8230) );
  XNOR U8498 ( .A(n8231), .B(n8230), .Z(n8200) );
  NAND U8499 ( .A(n8190), .B(n8189), .Z(n8194) );
  NAND U8500 ( .A(n8192), .B(n8191), .Z(n8193) );
  NAND U8501 ( .A(n8194), .B(n8193), .Z(n8201) );
  XNOR U8502 ( .A(n8200), .B(n8201), .Z(n8202) );
  XNOR U8503 ( .A(n8203), .B(n8202), .Z(n8234) );
  XNOR U8504 ( .A(n8234), .B(sreg[448]), .Z(n8236) );
  NAND U8505 ( .A(n8195), .B(sreg[447]), .Z(n8199) );
  OR U8506 ( .A(n8197), .B(n8196), .Z(n8198) );
  AND U8507 ( .A(n8199), .B(n8198), .Z(n8235) );
  XOR U8508 ( .A(n8236), .B(n8235), .Z(c[448]) );
  NANDN U8509 ( .A(n8205), .B(n8204), .Z(n8209) );
  NAND U8510 ( .A(n8207), .B(n8206), .Z(n8208) );
  NAND U8511 ( .A(n8209), .B(n8208), .Z(n8270) );
  NANDN U8512 ( .A(n8211), .B(n8210), .Z(n8215) );
  NAND U8513 ( .A(n8213), .B(n8212), .Z(n8214) );
  NAND U8514 ( .A(n8215), .B(n8214), .Z(n8268) );
  XNOR U8515 ( .A(b[7]), .B(a[195]), .Z(n8255) );
  NANDN U8516 ( .A(n8255), .B(n10545), .Z(n8218) );
  NANDN U8517 ( .A(n8216), .B(n10546), .Z(n8217) );
  NAND U8518 ( .A(n8218), .B(n8217), .Z(n8243) );
  XNOR U8519 ( .A(b[3]), .B(a[199]), .Z(n8258) );
  NANDN U8520 ( .A(n8258), .B(n10398), .Z(n8221) );
  NANDN U8521 ( .A(n8219), .B(n10399), .Z(n8220) );
  AND U8522 ( .A(n8221), .B(n8220), .Z(n8244) );
  XNOR U8523 ( .A(n8243), .B(n8244), .Z(n8245) );
  NANDN U8524 ( .A(n527), .B(a[201]), .Z(n8222) );
  XOR U8525 ( .A(n10434), .B(n8222), .Z(n8224) );
  NANDN U8526 ( .A(b[0]), .B(a[200]), .Z(n8223) );
  AND U8527 ( .A(n8224), .B(n8223), .Z(n8251) );
  XOR U8528 ( .A(b[5]), .B(a[197]), .Z(n8264) );
  NAND U8529 ( .A(n8264), .B(n10481), .Z(n8227) );
  NAND U8530 ( .A(n8225), .B(n10482), .Z(n8226) );
  NAND U8531 ( .A(n8227), .B(n8226), .Z(n8249) );
  NANDN U8532 ( .A(n529), .B(a[193]), .Z(n8250) );
  XNOR U8533 ( .A(n8249), .B(n8250), .Z(n8252) );
  XOR U8534 ( .A(n8251), .B(n8252), .Z(n8246) );
  XOR U8535 ( .A(n8245), .B(n8246), .Z(n8267) );
  XOR U8536 ( .A(n8268), .B(n8267), .Z(n8269) );
  XNOR U8537 ( .A(n8270), .B(n8269), .Z(n8239) );
  NAND U8538 ( .A(n8229), .B(n8228), .Z(n8233) );
  NAND U8539 ( .A(n8231), .B(n8230), .Z(n8232) );
  NAND U8540 ( .A(n8233), .B(n8232), .Z(n8240) );
  XNOR U8541 ( .A(n8239), .B(n8240), .Z(n8241) );
  XNOR U8542 ( .A(n8242), .B(n8241), .Z(n8273) );
  XNOR U8543 ( .A(n8273), .B(sreg[449]), .Z(n8275) );
  NAND U8544 ( .A(n8234), .B(sreg[448]), .Z(n8238) );
  OR U8545 ( .A(n8236), .B(n8235), .Z(n8237) );
  AND U8546 ( .A(n8238), .B(n8237), .Z(n8274) );
  XOR U8547 ( .A(n8275), .B(n8274), .Z(c[449]) );
  NANDN U8548 ( .A(n8244), .B(n8243), .Z(n8248) );
  NAND U8549 ( .A(n8246), .B(n8245), .Z(n8247) );
  NAND U8550 ( .A(n8248), .B(n8247), .Z(n8309) );
  NANDN U8551 ( .A(n8250), .B(n8249), .Z(n8254) );
  NAND U8552 ( .A(n8252), .B(n8251), .Z(n8253) );
  NAND U8553 ( .A(n8254), .B(n8253), .Z(n8307) );
  XNOR U8554 ( .A(b[7]), .B(a[196]), .Z(n8294) );
  NANDN U8555 ( .A(n8294), .B(n10545), .Z(n8257) );
  NANDN U8556 ( .A(n8255), .B(n10546), .Z(n8256) );
  NAND U8557 ( .A(n8257), .B(n8256), .Z(n8282) );
  XNOR U8558 ( .A(b[3]), .B(a[200]), .Z(n8297) );
  NANDN U8559 ( .A(n8297), .B(n10398), .Z(n8260) );
  NANDN U8560 ( .A(n8258), .B(n10399), .Z(n8259) );
  AND U8561 ( .A(n8260), .B(n8259), .Z(n8283) );
  XNOR U8562 ( .A(n8282), .B(n8283), .Z(n8284) );
  NANDN U8563 ( .A(n527), .B(a[202]), .Z(n8261) );
  XOR U8564 ( .A(n10434), .B(n8261), .Z(n8263) );
  NANDN U8565 ( .A(b[0]), .B(a[201]), .Z(n8262) );
  AND U8566 ( .A(n8263), .B(n8262), .Z(n8290) );
  XOR U8567 ( .A(b[5]), .B(a[198]), .Z(n8303) );
  NAND U8568 ( .A(n8303), .B(n10481), .Z(n8266) );
  NAND U8569 ( .A(n8264), .B(n10482), .Z(n8265) );
  NAND U8570 ( .A(n8266), .B(n8265), .Z(n8288) );
  NANDN U8571 ( .A(n529), .B(a[194]), .Z(n8289) );
  XNOR U8572 ( .A(n8288), .B(n8289), .Z(n8291) );
  XOR U8573 ( .A(n8290), .B(n8291), .Z(n8285) );
  XOR U8574 ( .A(n8284), .B(n8285), .Z(n8306) );
  XOR U8575 ( .A(n8307), .B(n8306), .Z(n8308) );
  XNOR U8576 ( .A(n8309), .B(n8308), .Z(n8278) );
  NAND U8577 ( .A(n8268), .B(n8267), .Z(n8272) );
  NAND U8578 ( .A(n8270), .B(n8269), .Z(n8271) );
  NAND U8579 ( .A(n8272), .B(n8271), .Z(n8279) );
  XNOR U8580 ( .A(n8278), .B(n8279), .Z(n8280) );
  XNOR U8581 ( .A(n8281), .B(n8280), .Z(n8312) );
  XNOR U8582 ( .A(n8312), .B(sreg[450]), .Z(n8314) );
  NAND U8583 ( .A(n8273), .B(sreg[449]), .Z(n8277) );
  OR U8584 ( .A(n8275), .B(n8274), .Z(n8276) );
  AND U8585 ( .A(n8277), .B(n8276), .Z(n8313) );
  XOR U8586 ( .A(n8314), .B(n8313), .Z(c[450]) );
  NANDN U8587 ( .A(n8283), .B(n8282), .Z(n8287) );
  NAND U8588 ( .A(n8285), .B(n8284), .Z(n8286) );
  NAND U8589 ( .A(n8287), .B(n8286), .Z(n8348) );
  NANDN U8590 ( .A(n8289), .B(n8288), .Z(n8293) );
  NAND U8591 ( .A(n8291), .B(n8290), .Z(n8292) );
  NAND U8592 ( .A(n8293), .B(n8292), .Z(n8346) );
  XNOR U8593 ( .A(b[7]), .B(a[197]), .Z(n8339) );
  NANDN U8594 ( .A(n8339), .B(n10545), .Z(n8296) );
  NANDN U8595 ( .A(n8294), .B(n10546), .Z(n8295) );
  NAND U8596 ( .A(n8296), .B(n8295), .Z(n8321) );
  XNOR U8597 ( .A(b[3]), .B(a[201]), .Z(n8342) );
  NANDN U8598 ( .A(n8342), .B(n10398), .Z(n8299) );
  NANDN U8599 ( .A(n8297), .B(n10399), .Z(n8298) );
  AND U8600 ( .A(n8299), .B(n8298), .Z(n8322) );
  XNOR U8601 ( .A(n8321), .B(n8322), .Z(n8323) );
  NANDN U8602 ( .A(n527), .B(a[203]), .Z(n8300) );
  XOR U8603 ( .A(n10434), .B(n8300), .Z(n8302) );
  NANDN U8604 ( .A(b[0]), .B(a[202]), .Z(n8301) );
  AND U8605 ( .A(n8302), .B(n8301), .Z(n8329) );
  XOR U8606 ( .A(b[5]), .B(a[199]), .Z(n8336) );
  NAND U8607 ( .A(n8336), .B(n10481), .Z(n8305) );
  NAND U8608 ( .A(n8303), .B(n10482), .Z(n8304) );
  NAND U8609 ( .A(n8305), .B(n8304), .Z(n8327) );
  NANDN U8610 ( .A(n529), .B(a[195]), .Z(n8328) );
  XNOR U8611 ( .A(n8327), .B(n8328), .Z(n8330) );
  XOR U8612 ( .A(n8329), .B(n8330), .Z(n8324) );
  XOR U8613 ( .A(n8323), .B(n8324), .Z(n8345) );
  XOR U8614 ( .A(n8346), .B(n8345), .Z(n8347) );
  XNOR U8615 ( .A(n8348), .B(n8347), .Z(n8317) );
  NAND U8616 ( .A(n8307), .B(n8306), .Z(n8311) );
  NAND U8617 ( .A(n8309), .B(n8308), .Z(n8310) );
  NAND U8618 ( .A(n8311), .B(n8310), .Z(n8318) );
  XNOR U8619 ( .A(n8317), .B(n8318), .Z(n8319) );
  XNOR U8620 ( .A(n8320), .B(n8319), .Z(n8351) );
  XNOR U8621 ( .A(n8351), .B(sreg[451]), .Z(n8353) );
  NAND U8622 ( .A(n8312), .B(sreg[450]), .Z(n8316) );
  OR U8623 ( .A(n8314), .B(n8313), .Z(n8315) );
  AND U8624 ( .A(n8316), .B(n8315), .Z(n8352) );
  XOR U8625 ( .A(n8353), .B(n8352), .Z(c[451]) );
  NANDN U8626 ( .A(n8322), .B(n8321), .Z(n8326) );
  NAND U8627 ( .A(n8324), .B(n8323), .Z(n8325) );
  NAND U8628 ( .A(n8326), .B(n8325), .Z(n8387) );
  NANDN U8629 ( .A(n8328), .B(n8327), .Z(n8332) );
  NAND U8630 ( .A(n8330), .B(n8329), .Z(n8331) );
  NAND U8631 ( .A(n8332), .B(n8331), .Z(n8385) );
  NANDN U8632 ( .A(n527), .B(a[204]), .Z(n8333) );
  XOR U8633 ( .A(n10434), .B(n8333), .Z(n8335) );
  NANDN U8634 ( .A(b[0]), .B(a[203]), .Z(n8334) );
  AND U8635 ( .A(n8335), .B(n8334), .Z(n8368) );
  XOR U8636 ( .A(b[5]), .B(a[200]), .Z(n8381) );
  NAND U8637 ( .A(n8381), .B(n10481), .Z(n8338) );
  NAND U8638 ( .A(n8336), .B(n10482), .Z(n8337) );
  NAND U8639 ( .A(n8338), .B(n8337), .Z(n8366) );
  NANDN U8640 ( .A(n529), .B(a[196]), .Z(n8367) );
  XNOR U8641 ( .A(n8366), .B(n8367), .Z(n8369) );
  XOR U8642 ( .A(n8368), .B(n8369), .Z(n8362) );
  XNOR U8643 ( .A(b[7]), .B(a[198]), .Z(n8372) );
  NANDN U8644 ( .A(n8372), .B(n10545), .Z(n8341) );
  NANDN U8645 ( .A(n8339), .B(n10546), .Z(n8340) );
  NAND U8646 ( .A(n8341), .B(n8340), .Z(n8360) );
  XNOR U8647 ( .A(b[3]), .B(a[202]), .Z(n8375) );
  NANDN U8648 ( .A(n8375), .B(n10398), .Z(n8344) );
  NANDN U8649 ( .A(n8342), .B(n10399), .Z(n8343) );
  AND U8650 ( .A(n8344), .B(n8343), .Z(n8361) );
  XNOR U8651 ( .A(n8360), .B(n8361), .Z(n8363) );
  XOR U8652 ( .A(n8362), .B(n8363), .Z(n8384) );
  XOR U8653 ( .A(n8385), .B(n8384), .Z(n8386) );
  XNOR U8654 ( .A(n8387), .B(n8386), .Z(n8356) );
  NAND U8655 ( .A(n8346), .B(n8345), .Z(n8350) );
  NAND U8656 ( .A(n8348), .B(n8347), .Z(n8349) );
  NAND U8657 ( .A(n8350), .B(n8349), .Z(n8357) );
  XNOR U8658 ( .A(n8356), .B(n8357), .Z(n8358) );
  XNOR U8659 ( .A(n8359), .B(n8358), .Z(n8390) );
  XNOR U8660 ( .A(n8390), .B(sreg[452]), .Z(n8392) );
  NAND U8661 ( .A(n8351), .B(sreg[451]), .Z(n8355) );
  OR U8662 ( .A(n8353), .B(n8352), .Z(n8354) );
  AND U8663 ( .A(n8355), .B(n8354), .Z(n8391) );
  XOR U8664 ( .A(n8392), .B(n8391), .Z(c[452]) );
  NANDN U8665 ( .A(n8361), .B(n8360), .Z(n8365) );
  NAND U8666 ( .A(n8363), .B(n8362), .Z(n8364) );
  NAND U8667 ( .A(n8365), .B(n8364), .Z(n8426) );
  NANDN U8668 ( .A(n8367), .B(n8366), .Z(n8371) );
  NAND U8669 ( .A(n8369), .B(n8368), .Z(n8370) );
  NAND U8670 ( .A(n8371), .B(n8370), .Z(n8424) );
  XNOR U8671 ( .A(b[7]), .B(a[199]), .Z(n8411) );
  NANDN U8672 ( .A(n8411), .B(n10545), .Z(n8374) );
  NANDN U8673 ( .A(n8372), .B(n10546), .Z(n8373) );
  NAND U8674 ( .A(n8374), .B(n8373), .Z(n8399) );
  XNOR U8675 ( .A(b[3]), .B(a[203]), .Z(n8414) );
  NANDN U8676 ( .A(n8414), .B(n10398), .Z(n8377) );
  NANDN U8677 ( .A(n8375), .B(n10399), .Z(n8376) );
  AND U8678 ( .A(n8377), .B(n8376), .Z(n8400) );
  XNOR U8679 ( .A(n8399), .B(n8400), .Z(n8401) );
  NANDN U8680 ( .A(n527), .B(a[205]), .Z(n8378) );
  XOR U8681 ( .A(n10434), .B(n8378), .Z(n8380) );
  IV U8682 ( .A(a[204]), .Z(n8645) );
  NANDN U8683 ( .A(n8645), .B(n527), .Z(n8379) );
  AND U8684 ( .A(n8380), .B(n8379), .Z(n8407) );
  XOR U8685 ( .A(b[5]), .B(a[201]), .Z(n8420) );
  NAND U8686 ( .A(n8420), .B(n10481), .Z(n8383) );
  NAND U8687 ( .A(n8381), .B(n10482), .Z(n8382) );
  NAND U8688 ( .A(n8383), .B(n8382), .Z(n8405) );
  NANDN U8689 ( .A(n529), .B(a[197]), .Z(n8406) );
  XNOR U8690 ( .A(n8405), .B(n8406), .Z(n8408) );
  XOR U8691 ( .A(n8407), .B(n8408), .Z(n8402) );
  XOR U8692 ( .A(n8401), .B(n8402), .Z(n8423) );
  XOR U8693 ( .A(n8424), .B(n8423), .Z(n8425) );
  XNOR U8694 ( .A(n8426), .B(n8425), .Z(n8395) );
  NAND U8695 ( .A(n8385), .B(n8384), .Z(n8389) );
  NAND U8696 ( .A(n8387), .B(n8386), .Z(n8388) );
  NAND U8697 ( .A(n8389), .B(n8388), .Z(n8396) );
  XNOR U8698 ( .A(n8395), .B(n8396), .Z(n8397) );
  XNOR U8699 ( .A(n8398), .B(n8397), .Z(n8429) );
  XNOR U8700 ( .A(n8429), .B(sreg[453]), .Z(n8431) );
  NAND U8701 ( .A(n8390), .B(sreg[452]), .Z(n8394) );
  OR U8702 ( .A(n8392), .B(n8391), .Z(n8393) );
  AND U8703 ( .A(n8394), .B(n8393), .Z(n8430) );
  XOR U8704 ( .A(n8431), .B(n8430), .Z(c[453]) );
  NANDN U8705 ( .A(n8400), .B(n8399), .Z(n8404) );
  NAND U8706 ( .A(n8402), .B(n8401), .Z(n8403) );
  NAND U8707 ( .A(n8404), .B(n8403), .Z(n8465) );
  NANDN U8708 ( .A(n8406), .B(n8405), .Z(n8410) );
  NAND U8709 ( .A(n8408), .B(n8407), .Z(n8409) );
  NAND U8710 ( .A(n8410), .B(n8409), .Z(n8463) );
  XNOR U8711 ( .A(b[7]), .B(a[200]), .Z(n8450) );
  NANDN U8712 ( .A(n8450), .B(n10545), .Z(n8413) );
  NANDN U8713 ( .A(n8411), .B(n10546), .Z(n8412) );
  NAND U8714 ( .A(n8413), .B(n8412), .Z(n8438) );
  XOR U8715 ( .A(b[3]), .B(n8645), .Z(n8453) );
  NANDN U8716 ( .A(n8453), .B(n10398), .Z(n8416) );
  NANDN U8717 ( .A(n8414), .B(n10399), .Z(n8415) );
  AND U8718 ( .A(n8416), .B(n8415), .Z(n8439) );
  XNOR U8719 ( .A(n8438), .B(n8439), .Z(n8440) );
  NANDN U8720 ( .A(n527), .B(a[206]), .Z(n8417) );
  XOR U8721 ( .A(n10434), .B(n8417), .Z(n8419) );
  NANDN U8722 ( .A(b[0]), .B(a[205]), .Z(n8418) );
  AND U8723 ( .A(n8419), .B(n8418), .Z(n8446) );
  XOR U8724 ( .A(b[5]), .B(a[202]), .Z(n8459) );
  NAND U8725 ( .A(n8459), .B(n10481), .Z(n8422) );
  NAND U8726 ( .A(n8420), .B(n10482), .Z(n8421) );
  NAND U8727 ( .A(n8422), .B(n8421), .Z(n8444) );
  NANDN U8728 ( .A(n529), .B(a[198]), .Z(n8445) );
  XNOR U8729 ( .A(n8444), .B(n8445), .Z(n8447) );
  XOR U8730 ( .A(n8446), .B(n8447), .Z(n8441) );
  XOR U8731 ( .A(n8440), .B(n8441), .Z(n8462) );
  XOR U8732 ( .A(n8463), .B(n8462), .Z(n8464) );
  XNOR U8733 ( .A(n8465), .B(n8464), .Z(n8434) );
  NAND U8734 ( .A(n8424), .B(n8423), .Z(n8428) );
  NAND U8735 ( .A(n8426), .B(n8425), .Z(n8427) );
  NAND U8736 ( .A(n8428), .B(n8427), .Z(n8435) );
  XNOR U8737 ( .A(n8434), .B(n8435), .Z(n8436) );
  XNOR U8738 ( .A(n8437), .B(n8436), .Z(n8468) );
  XNOR U8739 ( .A(n8468), .B(sreg[454]), .Z(n8470) );
  NAND U8740 ( .A(n8429), .B(sreg[453]), .Z(n8433) );
  OR U8741 ( .A(n8431), .B(n8430), .Z(n8432) );
  AND U8742 ( .A(n8433), .B(n8432), .Z(n8469) );
  XOR U8743 ( .A(n8470), .B(n8469), .Z(c[454]) );
  NANDN U8744 ( .A(n8439), .B(n8438), .Z(n8443) );
  NAND U8745 ( .A(n8441), .B(n8440), .Z(n8442) );
  NAND U8746 ( .A(n8443), .B(n8442), .Z(n8504) );
  NANDN U8747 ( .A(n8445), .B(n8444), .Z(n8449) );
  NAND U8748 ( .A(n8447), .B(n8446), .Z(n8448) );
  NAND U8749 ( .A(n8449), .B(n8448), .Z(n8502) );
  XNOR U8750 ( .A(b[7]), .B(a[201]), .Z(n8489) );
  NANDN U8751 ( .A(n8489), .B(n10545), .Z(n8452) );
  NANDN U8752 ( .A(n8450), .B(n10546), .Z(n8451) );
  NAND U8753 ( .A(n8452), .B(n8451), .Z(n8477) );
  XNOR U8754 ( .A(b[3]), .B(a[205]), .Z(n8492) );
  NANDN U8755 ( .A(n8492), .B(n10398), .Z(n8455) );
  NANDN U8756 ( .A(n8453), .B(n10399), .Z(n8454) );
  AND U8757 ( .A(n8455), .B(n8454), .Z(n8478) );
  XNOR U8758 ( .A(n8477), .B(n8478), .Z(n8479) );
  NANDN U8759 ( .A(n527), .B(a[207]), .Z(n8456) );
  XOR U8760 ( .A(n10434), .B(n8456), .Z(n8458) );
  NANDN U8761 ( .A(b[0]), .B(a[206]), .Z(n8457) );
  AND U8762 ( .A(n8458), .B(n8457), .Z(n8485) );
  XOR U8763 ( .A(b[5]), .B(a[203]), .Z(n8498) );
  NAND U8764 ( .A(n8498), .B(n10481), .Z(n8461) );
  NAND U8765 ( .A(n8459), .B(n10482), .Z(n8460) );
  NAND U8766 ( .A(n8461), .B(n8460), .Z(n8483) );
  NANDN U8767 ( .A(n529), .B(a[199]), .Z(n8484) );
  XNOR U8768 ( .A(n8483), .B(n8484), .Z(n8486) );
  XOR U8769 ( .A(n8485), .B(n8486), .Z(n8480) );
  XOR U8770 ( .A(n8479), .B(n8480), .Z(n8501) );
  XOR U8771 ( .A(n8502), .B(n8501), .Z(n8503) );
  XNOR U8772 ( .A(n8504), .B(n8503), .Z(n8473) );
  NAND U8773 ( .A(n8463), .B(n8462), .Z(n8467) );
  NAND U8774 ( .A(n8465), .B(n8464), .Z(n8466) );
  NAND U8775 ( .A(n8467), .B(n8466), .Z(n8474) );
  XNOR U8776 ( .A(n8473), .B(n8474), .Z(n8475) );
  XNOR U8777 ( .A(n8476), .B(n8475), .Z(n8507) );
  XNOR U8778 ( .A(n8507), .B(sreg[455]), .Z(n8509) );
  NAND U8779 ( .A(n8468), .B(sreg[454]), .Z(n8472) );
  OR U8780 ( .A(n8470), .B(n8469), .Z(n8471) );
  AND U8781 ( .A(n8472), .B(n8471), .Z(n8508) );
  XOR U8782 ( .A(n8509), .B(n8508), .Z(c[455]) );
  NANDN U8783 ( .A(n8478), .B(n8477), .Z(n8482) );
  NAND U8784 ( .A(n8480), .B(n8479), .Z(n8481) );
  NAND U8785 ( .A(n8482), .B(n8481), .Z(n8543) );
  NANDN U8786 ( .A(n8484), .B(n8483), .Z(n8488) );
  NAND U8787 ( .A(n8486), .B(n8485), .Z(n8487) );
  NAND U8788 ( .A(n8488), .B(n8487), .Z(n8541) );
  XNOR U8789 ( .A(b[7]), .B(a[202]), .Z(n8528) );
  NANDN U8790 ( .A(n8528), .B(n10545), .Z(n8491) );
  NANDN U8791 ( .A(n8489), .B(n10546), .Z(n8490) );
  NAND U8792 ( .A(n8491), .B(n8490), .Z(n8516) );
  XNOR U8793 ( .A(b[3]), .B(a[206]), .Z(n8531) );
  NANDN U8794 ( .A(n8531), .B(n10398), .Z(n8494) );
  NANDN U8795 ( .A(n8492), .B(n10399), .Z(n8493) );
  AND U8796 ( .A(n8494), .B(n8493), .Z(n8517) );
  XNOR U8797 ( .A(n8516), .B(n8517), .Z(n8518) );
  NANDN U8798 ( .A(n527), .B(a[208]), .Z(n8495) );
  XOR U8799 ( .A(n10434), .B(n8495), .Z(n8497) );
  NANDN U8800 ( .A(b[0]), .B(a[207]), .Z(n8496) );
  AND U8801 ( .A(n8497), .B(n8496), .Z(n8524) );
  XNOR U8802 ( .A(b[5]), .B(a[204]), .Z(n8537) );
  NANDN U8803 ( .A(n8537), .B(n10481), .Z(n8500) );
  NAND U8804 ( .A(n8498), .B(n10482), .Z(n8499) );
  NAND U8805 ( .A(n8500), .B(n8499), .Z(n8522) );
  NANDN U8806 ( .A(n529), .B(a[200]), .Z(n8523) );
  XNOR U8807 ( .A(n8522), .B(n8523), .Z(n8525) );
  XOR U8808 ( .A(n8524), .B(n8525), .Z(n8519) );
  XOR U8809 ( .A(n8518), .B(n8519), .Z(n8540) );
  XOR U8810 ( .A(n8541), .B(n8540), .Z(n8542) );
  XNOR U8811 ( .A(n8543), .B(n8542), .Z(n8512) );
  NAND U8812 ( .A(n8502), .B(n8501), .Z(n8506) );
  NAND U8813 ( .A(n8504), .B(n8503), .Z(n8505) );
  NAND U8814 ( .A(n8506), .B(n8505), .Z(n8513) );
  XNOR U8815 ( .A(n8512), .B(n8513), .Z(n8514) );
  XNOR U8816 ( .A(n8515), .B(n8514), .Z(n8546) );
  XNOR U8817 ( .A(n8546), .B(sreg[456]), .Z(n8548) );
  NAND U8818 ( .A(n8507), .B(sreg[455]), .Z(n8511) );
  OR U8819 ( .A(n8509), .B(n8508), .Z(n8510) );
  AND U8820 ( .A(n8511), .B(n8510), .Z(n8547) );
  XOR U8821 ( .A(n8548), .B(n8547), .Z(c[456]) );
  NANDN U8822 ( .A(n8517), .B(n8516), .Z(n8521) );
  NAND U8823 ( .A(n8519), .B(n8518), .Z(n8520) );
  NAND U8824 ( .A(n8521), .B(n8520), .Z(n8582) );
  NANDN U8825 ( .A(n8523), .B(n8522), .Z(n8527) );
  NAND U8826 ( .A(n8525), .B(n8524), .Z(n8526) );
  NAND U8827 ( .A(n8527), .B(n8526), .Z(n8580) );
  XNOR U8828 ( .A(b[7]), .B(a[203]), .Z(n8567) );
  NANDN U8829 ( .A(n8567), .B(n10545), .Z(n8530) );
  NANDN U8830 ( .A(n8528), .B(n10546), .Z(n8529) );
  NAND U8831 ( .A(n8530), .B(n8529), .Z(n8555) );
  XNOR U8832 ( .A(b[3]), .B(a[207]), .Z(n8570) );
  NANDN U8833 ( .A(n8570), .B(n10398), .Z(n8533) );
  NANDN U8834 ( .A(n8531), .B(n10399), .Z(n8532) );
  AND U8835 ( .A(n8533), .B(n8532), .Z(n8556) );
  XNOR U8836 ( .A(n8555), .B(n8556), .Z(n8557) );
  NANDN U8837 ( .A(n527), .B(a[209]), .Z(n8534) );
  XOR U8838 ( .A(n10434), .B(n8534), .Z(n8536) );
  NANDN U8839 ( .A(b[0]), .B(a[208]), .Z(n8535) );
  AND U8840 ( .A(n8536), .B(n8535), .Z(n8563) );
  XOR U8841 ( .A(b[5]), .B(a[205]), .Z(n8576) );
  NAND U8842 ( .A(n8576), .B(n10481), .Z(n8539) );
  NANDN U8843 ( .A(n8537), .B(n10482), .Z(n8538) );
  NAND U8844 ( .A(n8539), .B(n8538), .Z(n8561) );
  NANDN U8845 ( .A(n529), .B(a[201]), .Z(n8562) );
  XNOR U8846 ( .A(n8561), .B(n8562), .Z(n8564) );
  XOR U8847 ( .A(n8563), .B(n8564), .Z(n8558) );
  XOR U8848 ( .A(n8557), .B(n8558), .Z(n8579) );
  XOR U8849 ( .A(n8580), .B(n8579), .Z(n8581) );
  XNOR U8850 ( .A(n8582), .B(n8581), .Z(n8551) );
  NAND U8851 ( .A(n8541), .B(n8540), .Z(n8545) );
  NAND U8852 ( .A(n8543), .B(n8542), .Z(n8544) );
  NAND U8853 ( .A(n8545), .B(n8544), .Z(n8552) );
  XNOR U8854 ( .A(n8551), .B(n8552), .Z(n8553) );
  XNOR U8855 ( .A(n8554), .B(n8553), .Z(n8585) );
  XNOR U8856 ( .A(n8585), .B(sreg[457]), .Z(n8587) );
  NAND U8857 ( .A(n8546), .B(sreg[456]), .Z(n8550) );
  OR U8858 ( .A(n8548), .B(n8547), .Z(n8549) );
  AND U8859 ( .A(n8550), .B(n8549), .Z(n8586) );
  XOR U8860 ( .A(n8587), .B(n8586), .Z(c[457]) );
  NANDN U8861 ( .A(n8556), .B(n8555), .Z(n8560) );
  NAND U8862 ( .A(n8558), .B(n8557), .Z(n8559) );
  NAND U8863 ( .A(n8560), .B(n8559), .Z(n8621) );
  NANDN U8864 ( .A(n8562), .B(n8561), .Z(n8566) );
  NAND U8865 ( .A(n8564), .B(n8563), .Z(n8565) );
  NAND U8866 ( .A(n8566), .B(n8565), .Z(n8619) );
  XOR U8867 ( .A(b[7]), .B(n8645), .Z(n8606) );
  NANDN U8868 ( .A(n8606), .B(n10545), .Z(n8569) );
  NANDN U8869 ( .A(n8567), .B(n10546), .Z(n8568) );
  NAND U8870 ( .A(n8569), .B(n8568), .Z(n8594) );
  XNOR U8871 ( .A(b[3]), .B(a[208]), .Z(n8609) );
  NANDN U8872 ( .A(n8609), .B(n10398), .Z(n8572) );
  NANDN U8873 ( .A(n8570), .B(n10399), .Z(n8571) );
  AND U8874 ( .A(n8572), .B(n8571), .Z(n8595) );
  XNOR U8875 ( .A(n8594), .B(n8595), .Z(n8596) );
  NANDN U8876 ( .A(n527), .B(a[210]), .Z(n8573) );
  XOR U8877 ( .A(n10434), .B(n8573), .Z(n8575) );
  NANDN U8878 ( .A(b[0]), .B(a[209]), .Z(n8574) );
  AND U8879 ( .A(n8575), .B(n8574), .Z(n8602) );
  XOR U8880 ( .A(b[5]), .B(a[206]), .Z(n8615) );
  NAND U8881 ( .A(n8615), .B(n10481), .Z(n8578) );
  NAND U8882 ( .A(n8576), .B(n10482), .Z(n8577) );
  NAND U8883 ( .A(n8578), .B(n8577), .Z(n8600) );
  NANDN U8884 ( .A(n529), .B(a[202]), .Z(n8601) );
  XNOR U8885 ( .A(n8600), .B(n8601), .Z(n8603) );
  XOR U8886 ( .A(n8602), .B(n8603), .Z(n8597) );
  XOR U8887 ( .A(n8596), .B(n8597), .Z(n8618) );
  XOR U8888 ( .A(n8619), .B(n8618), .Z(n8620) );
  XNOR U8889 ( .A(n8621), .B(n8620), .Z(n8590) );
  NAND U8890 ( .A(n8580), .B(n8579), .Z(n8584) );
  NAND U8891 ( .A(n8582), .B(n8581), .Z(n8583) );
  NAND U8892 ( .A(n8584), .B(n8583), .Z(n8591) );
  XNOR U8893 ( .A(n8590), .B(n8591), .Z(n8592) );
  XNOR U8894 ( .A(n8593), .B(n8592), .Z(n8624) );
  XNOR U8895 ( .A(n8624), .B(sreg[458]), .Z(n8626) );
  NAND U8896 ( .A(n8585), .B(sreg[457]), .Z(n8589) );
  OR U8897 ( .A(n8587), .B(n8586), .Z(n8588) );
  AND U8898 ( .A(n8589), .B(n8588), .Z(n8625) );
  XOR U8899 ( .A(n8626), .B(n8625), .Z(c[458]) );
  NANDN U8900 ( .A(n8595), .B(n8594), .Z(n8599) );
  NAND U8901 ( .A(n8597), .B(n8596), .Z(n8598) );
  NAND U8902 ( .A(n8599), .B(n8598), .Z(n8661) );
  NANDN U8903 ( .A(n8601), .B(n8600), .Z(n8605) );
  NAND U8904 ( .A(n8603), .B(n8602), .Z(n8604) );
  NAND U8905 ( .A(n8605), .B(n8604), .Z(n8659) );
  XNOR U8906 ( .A(b[7]), .B(a[205]), .Z(n8652) );
  NANDN U8907 ( .A(n8652), .B(n10545), .Z(n8608) );
  NANDN U8908 ( .A(n8606), .B(n10546), .Z(n8607) );
  NAND U8909 ( .A(n8608), .B(n8607), .Z(n8633) );
  XNOR U8910 ( .A(b[3]), .B(a[209]), .Z(n8655) );
  NANDN U8911 ( .A(n8655), .B(n10398), .Z(n8611) );
  NANDN U8912 ( .A(n8609), .B(n10399), .Z(n8610) );
  AND U8913 ( .A(n8611), .B(n8610), .Z(n8634) );
  XNOR U8914 ( .A(n8633), .B(n8634), .Z(n8635) );
  NANDN U8915 ( .A(n527), .B(a[211]), .Z(n8612) );
  XOR U8916 ( .A(n10434), .B(n8612), .Z(n8614) );
  NANDN U8917 ( .A(b[0]), .B(a[210]), .Z(n8613) );
  AND U8918 ( .A(n8614), .B(n8613), .Z(n8641) );
  XOR U8919 ( .A(b[5]), .B(a[207]), .Z(n8646) );
  NAND U8920 ( .A(n8646), .B(n10481), .Z(n8617) );
  NAND U8921 ( .A(n8615), .B(n10482), .Z(n8616) );
  NAND U8922 ( .A(n8617), .B(n8616), .Z(n8639) );
  NANDN U8923 ( .A(n529), .B(a[203]), .Z(n8640) );
  XNOR U8924 ( .A(n8639), .B(n8640), .Z(n8642) );
  XOR U8925 ( .A(n8641), .B(n8642), .Z(n8636) );
  XOR U8926 ( .A(n8635), .B(n8636), .Z(n8658) );
  XOR U8927 ( .A(n8659), .B(n8658), .Z(n8660) );
  XNOR U8928 ( .A(n8661), .B(n8660), .Z(n8629) );
  NAND U8929 ( .A(n8619), .B(n8618), .Z(n8623) );
  NAND U8930 ( .A(n8621), .B(n8620), .Z(n8622) );
  NAND U8931 ( .A(n8623), .B(n8622), .Z(n8630) );
  XNOR U8932 ( .A(n8629), .B(n8630), .Z(n8631) );
  XNOR U8933 ( .A(n8632), .B(n8631), .Z(n8664) );
  XNOR U8934 ( .A(n8664), .B(sreg[459]), .Z(n8666) );
  NAND U8935 ( .A(n8624), .B(sreg[458]), .Z(n8628) );
  OR U8936 ( .A(n8626), .B(n8625), .Z(n8627) );
  AND U8937 ( .A(n8628), .B(n8627), .Z(n8665) );
  XOR U8938 ( .A(n8666), .B(n8665), .Z(c[459]) );
  NANDN U8939 ( .A(n8634), .B(n8633), .Z(n8638) );
  NAND U8940 ( .A(n8636), .B(n8635), .Z(n8637) );
  NAND U8941 ( .A(n8638), .B(n8637), .Z(n8700) );
  NANDN U8942 ( .A(n8640), .B(n8639), .Z(n8644) );
  NAND U8943 ( .A(n8642), .B(n8641), .Z(n8643) );
  NAND U8944 ( .A(n8644), .B(n8643), .Z(n8697) );
  ANDN U8945 ( .B(b[7]), .A(n8645), .Z(n8679) );
  XOR U8946 ( .A(b[5]), .B(a[208]), .Z(n8694) );
  NAND U8947 ( .A(n10481), .B(n8694), .Z(n8648) );
  NAND U8948 ( .A(n10482), .B(n8646), .Z(n8647) );
  NAND U8949 ( .A(n8648), .B(n8647), .Z(n8680) );
  XOR U8950 ( .A(n8679), .B(n8680), .Z(n8681) );
  NANDN U8951 ( .A(n527), .B(a[212]), .Z(n8649) );
  XOR U8952 ( .A(n10434), .B(n8649), .Z(n8651) );
  NANDN U8953 ( .A(b[0]), .B(a[211]), .Z(n8650) );
  AND U8954 ( .A(n8651), .B(n8650), .Z(n8682) );
  XOR U8955 ( .A(n8681), .B(n8682), .Z(n8676) );
  XNOR U8956 ( .A(b[7]), .B(a[206]), .Z(n8685) );
  NANDN U8957 ( .A(n8685), .B(n10545), .Z(n8654) );
  NANDN U8958 ( .A(n8652), .B(n10546), .Z(n8653) );
  NAND U8959 ( .A(n8654), .B(n8653), .Z(n8673) );
  XNOR U8960 ( .A(b[3]), .B(a[210]), .Z(n8688) );
  NANDN U8961 ( .A(n8688), .B(n10398), .Z(n8657) );
  NANDN U8962 ( .A(n8655), .B(n10399), .Z(n8656) );
  AND U8963 ( .A(n8657), .B(n8656), .Z(n8674) );
  XNOR U8964 ( .A(n8673), .B(n8674), .Z(n8675) );
  XNOR U8965 ( .A(n8676), .B(n8675), .Z(n8698) );
  XNOR U8966 ( .A(n8697), .B(n8698), .Z(n8699) );
  XNOR U8967 ( .A(n8700), .B(n8699), .Z(n8669) );
  NAND U8968 ( .A(n8659), .B(n8658), .Z(n8663) );
  NAND U8969 ( .A(n8661), .B(n8660), .Z(n8662) );
  NAND U8970 ( .A(n8663), .B(n8662), .Z(n8670) );
  XNOR U8971 ( .A(n8669), .B(n8670), .Z(n8671) );
  XNOR U8972 ( .A(n8672), .B(n8671), .Z(n8703) );
  XNOR U8973 ( .A(n8703), .B(sreg[460]), .Z(n8705) );
  NAND U8974 ( .A(n8664), .B(sreg[459]), .Z(n8668) );
  OR U8975 ( .A(n8666), .B(n8665), .Z(n8667) );
  AND U8976 ( .A(n8668), .B(n8667), .Z(n8704) );
  XOR U8977 ( .A(n8705), .B(n8704), .Z(c[460]) );
  NANDN U8978 ( .A(n8674), .B(n8673), .Z(n8678) );
  NAND U8979 ( .A(n8676), .B(n8675), .Z(n8677) );
  NAND U8980 ( .A(n8678), .B(n8677), .Z(n8739) );
  OR U8981 ( .A(n8680), .B(n8679), .Z(n8684) );
  NANDN U8982 ( .A(n8682), .B(n8681), .Z(n8683) );
  NAND U8983 ( .A(n8684), .B(n8683), .Z(n8737) );
  XNOR U8984 ( .A(b[7]), .B(a[207]), .Z(n8724) );
  NANDN U8985 ( .A(n8724), .B(n10545), .Z(n8687) );
  NANDN U8986 ( .A(n8685), .B(n10546), .Z(n8686) );
  NAND U8987 ( .A(n8687), .B(n8686), .Z(n8712) );
  XNOR U8988 ( .A(b[3]), .B(a[211]), .Z(n8727) );
  NANDN U8989 ( .A(n8727), .B(n10398), .Z(n8690) );
  NANDN U8990 ( .A(n8688), .B(n10399), .Z(n8689) );
  AND U8991 ( .A(n8690), .B(n8689), .Z(n8713) );
  XNOR U8992 ( .A(n8712), .B(n8713), .Z(n8714) );
  NANDN U8993 ( .A(n527), .B(a[213]), .Z(n8691) );
  XOR U8994 ( .A(n10434), .B(n8691), .Z(n8693) );
  NANDN U8995 ( .A(b[0]), .B(a[212]), .Z(n8692) );
  AND U8996 ( .A(n8693), .B(n8692), .Z(n8720) );
  XOR U8997 ( .A(b[5]), .B(a[209]), .Z(n8733) );
  NAND U8998 ( .A(n8733), .B(n10481), .Z(n8696) );
  NAND U8999 ( .A(n8694), .B(n10482), .Z(n8695) );
  NAND U9000 ( .A(n8696), .B(n8695), .Z(n8718) );
  NANDN U9001 ( .A(n529), .B(a[205]), .Z(n8719) );
  XNOR U9002 ( .A(n8718), .B(n8719), .Z(n8721) );
  XOR U9003 ( .A(n8720), .B(n8721), .Z(n8715) );
  XOR U9004 ( .A(n8714), .B(n8715), .Z(n8736) );
  XNOR U9005 ( .A(n8737), .B(n8736), .Z(n8738) );
  XNOR U9006 ( .A(n8739), .B(n8738), .Z(n8708) );
  NANDN U9007 ( .A(n8698), .B(n8697), .Z(n8702) );
  NAND U9008 ( .A(n8700), .B(n8699), .Z(n8701) );
  NAND U9009 ( .A(n8702), .B(n8701), .Z(n8709) );
  XNOR U9010 ( .A(n8708), .B(n8709), .Z(n8710) );
  XNOR U9011 ( .A(n8711), .B(n8710), .Z(n8740) );
  XNOR U9012 ( .A(n8740), .B(sreg[461]), .Z(n8742) );
  NAND U9013 ( .A(n8703), .B(sreg[460]), .Z(n8707) );
  OR U9014 ( .A(n8705), .B(n8704), .Z(n8706) );
  AND U9015 ( .A(n8707), .B(n8706), .Z(n8741) );
  XOR U9016 ( .A(n8742), .B(n8741), .Z(c[461]) );
  NANDN U9017 ( .A(n8713), .B(n8712), .Z(n8717) );
  NAND U9018 ( .A(n8715), .B(n8714), .Z(n8716) );
  NAND U9019 ( .A(n8717), .B(n8716), .Z(n8776) );
  NANDN U9020 ( .A(n8719), .B(n8718), .Z(n8723) );
  NAND U9021 ( .A(n8721), .B(n8720), .Z(n8722) );
  NAND U9022 ( .A(n8723), .B(n8722), .Z(n8774) );
  XNOR U9023 ( .A(b[7]), .B(a[208]), .Z(n8761) );
  NANDN U9024 ( .A(n8761), .B(n10545), .Z(n8726) );
  NANDN U9025 ( .A(n8724), .B(n10546), .Z(n8725) );
  NAND U9026 ( .A(n8726), .B(n8725), .Z(n8749) );
  XNOR U9027 ( .A(b[3]), .B(a[212]), .Z(n8764) );
  NANDN U9028 ( .A(n8764), .B(n10398), .Z(n8729) );
  NANDN U9029 ( .A(n8727), .B(n10399), .Z(n8728) );
  AND U9030 ( .A(n8729), .B(n8728), .Z(n8750) );
  XNOR U9031 ( .A(n8749), .B(n8750), .Z(n8751) );
  NANDN U9032 ( .A(n527), .B(a[214]), .Z(n8730) );
  XOR U9033 ( .A(n10434), .B(n8730), .Z(n8732) );
  NANDN U9034 ( .A(b[0]), .B(a[213]), .Z(n8731) );
  AND U9035 ( .A(n8732), .B(n8731), .Z(n8757) );
  XOR U9036 ( .A(b[5]), .B(a[210]), .Z(n8770) );
  NAND U9037 ( .A(n8770), .B(n10481), .Z(n8735) );
  NAND U9038 ( .A(n8733), .B(n10482), .Z(n8734) );
  NAND U9039 ( .A(n8735), .B(n8734), .Z(n8755) );
  NANDN U9040 ( .A(n529), .B(a[206]), .Z(n8756) );
  XNOR U9041 ( .A(n8755), .B(n8756), .Z(n8758) );
  XOR U9042 ( .A(n8757), .B(n8758), .Z(n8752) );
  XOR U9043 ( .A(n8751), .B(n8752), .Z(n8773) );
  XOR U9044 ( .A(n8774), .B(n8773), .Z(n8775) );
  XNOR U9045 ( .A(n8776), .B(n8775), .Z(n8745) );
  XNOR U9046 ( .A(n8745), .B(n8746), .Z(n8747) );
  XNOR U9047 ( .A(n8748), .B(n8747), .Z(n8779) );
  XNOR U9048 ( .A(n8779), .B(sreg[462]), .Z(n8781) );
  NAND U9049 ( .A(n8740), .B(sreg[461]), .Z(n8744) );
  OR U9050 ( .A(n8742), .B(n8741), .Z(n8743) );
  AND U9051 ( .A(n8744), .B(n8743), .Z(n8780) );
  XOR U9052 ( .A(n8781), .B(n8780), .Z(c[462]) );
  NANDN U9053 ( .A(n8750), .B(n8749), .Z(n8754) );
  NAND U9054 ( .A(n8752), .B(n8751), .Z(n8753) );
  NAND U9055 ( .A(n8754), .B(n8753), .Z(n8815) );
  NANDN U9056 ( .A(n8756), .B(n8755), .Z(n8760) );
  NAND U9057 ( .A(n8758), .B(n8757), .Z(n8759) );
  NAND U9058 ( .A(n8760), .B(n8759), .Z(n8813) );
  XNOR U9059 ( .A(b[7]), .B(a[209]), .Z(n8800) );
  NANDN U9060 ( .A(n8800), .B(n10545), .Z(n8763) );
  NANDN U9061 ( .A(n8761), .B(n10546), .Z(n8762) );
  NAND U9062 ( .A(n8763), .B(n8762), .Z(n8788) );
  XNOR U9063 ( .A(b[3]), .B(a[213]), .Z(n8803) );
  NANDN U9064 ( .A(n8803), .B(n10398), .Z(n8766) );
  NANDN U9065 ( .A(n8764), .B(n10399), .Z(n8765) );
  AND U9066 ( .A(n8766), .B(n8765), .Z(n8789) );
  XNOR U9067 ( .A(n8788), .B(n8789), .Z(n8790) );
  NANDN U9068 ( .A(n527), .B(a[215]), .Z(n8767) );
  XOR U9069 ( .A(n10434), .B(n8767), .Z(n8769) );
  NANDN U9070 ( .A(b[0]), .B(a[214]), .Z(n8768) );
  AND U9071 ( .A(n8769), .B(n8768), .Z(n8796) );
  XOR U9072 ( .A(b[5]), .B(a[211]), .Z(n8809) );
  NAND U9073 ( .A(n8809), .B(n10481), .Z(n8772) );
  NAND U9074 ( .A(n8770), .B(n10482), .Z(n8771) );
  NAND U9075 ( .A(n8772), .B(n8771), .Z(n8794) );
  NANDN U9076 ( .A(n529), .B(a[207]), .Z(n8795) );
  XNOR U9077 ( .A(n8794), .B(n8795), .Z(n8797) );
  XOR U9078 ( .A(n8796), .B(n8797), .Z(n8791) );
  XOR U9079 ( .A(n8790), .B(n8791), .Z(n8812) );
  XOR U9080 ( .A(n8813), .B(n8812), .Z(n8814) );
  XNOR U9081 ( .A(n8815), .B(n8814), .Z(n8784) );
  NAND U9082 ( .A(n8774), .B(n8773), .Z(n8778) );
  NAND U9083 ( .A(n8776), .B(n8775), .Z(n8777) );
  NAND U9084 ( .A(n8778), .B(n8777), .Z(n8785) );
  XNOR U9085 ( .A(n8784), .B(n8785), .Z(n8786) );
  XNOR U9086 ( .A(n8787), .B(n8786), .Z(n8818) );
  XNOR U9087 ( .A(n8818), .B(sreg[463]), .Z(n8820) );
  NAND U9088 ( .A(n8779), .B(sreg[462]), .Z(n8783) );
  OR U9089 ( .A(n8781), .B(n8780), .Z(n8782) );
  AND U9090 ( .A(n8783), .B(n8782), .Z(n8819) );
  XOR U9091 ( .A(n8820), .B(n8819), .Z(c[463]) );
  NANDN U9092 ( .A(n8789), .B(n8788), .Z(n8793) );
  NAND U9093 ( .A(n8791), .B(n8790), .Z(n8792) );
  NAND U9094 ( .A(n8793), .B(n8792), .Z(n8854) );
  NANDN U9095 ( .A(n8795), .B(n8794), .Z(n8799) );
  NAND U9096 ( .A(n8797), .B(n8796), .Z(n8798) );
  NAND U9097 ( .A(n8799), .B(n8798), .Z(n8852) );
  XNOR U9098 ( .A(b[7]), .B(a[210]), .Z(n8839) );
  NANDN U9099 ( .A(n8839), .B(n10545), .Z(n8802) );
  NANDN U9100 ( .A(n8800), .B(n10546), .Z(n8801) );
  NAND U9101 ( .A(n8802), .B(n8801), .Z(n8827) );
  XNOR U9102 ( .A(b[3]), .B(a[214]), .Z(n8842) );
  NANDN U9103 ( .A(n8842), .B(n10398), .Z(n8805) );
  NANDN U9104 ( .A(n8803), .B(n10399), .Z(n8804) );
  AND U9105 ( .A(n8805), .B(n8804), .Z(n8828) );
  XNOR U9106 ( .A(n8827), .B(n8828), .Z(n8829) );
  NANDN U9107 ( .A(n527), .B(a[216]), .Z(n8806) );
  XOR U9108 ( .A(n10434), .B(n8806), .Z(n8808) );
  NANDN U9109 ( .A(b[0]), .B(a[215]), .Z(n8807) );
  AND U9110 ( .A(n8808), .B(n8807), .Z(n8835) );
  XOR U9111 ( .A(b[5]), .B(a[212]), .Z(n8848) );
  NAND U9112 ( .A(n8848), .B(n10481), .Z(n8811) );
  NAND U9113 ( .A(n8809), .B(n10482), .Z(n8810) );
  NAND U9114 ( .A(n8811), .B(n8810), .Z(n8833) );
  NANDN U9115 ( .A(n529), .B(a[208]), .Z(n8834) );
  XNOR U9116 ( .A(n8833), .B(n8834), .Z(n8836) );
  XOR U9117 ( .A(n8835), .B(n8836), .Z(n8830) );
  XOR U9118 ( .A(n8829), .B(n8830), .Z(n8851) );
  XOR U9119 ( .A(n8852), .B(n8851), .Z(n8853) );
  XNOR U9120 ( .A(n8854), .B(n8853), .Z(n8823) );
  NAND U9121 ( .A(n8813), .B(n8812), .Z(n8817) );
  NAND U9122 ( .A(n8815), .B(n8814), .Z(n8816) );
  NAND U9123 ( .A(n8817), .B(n8816), .Z(n8824) );
  XNOR U9124 ( .A(n8823), .B(n8824), .Z(n8825) );
  XNOR U9125 ( .A(n8826), .B(n8825), .Z(n8857) );
  XNOR U9126 ( .A(n8857), .B(sreg[464]), .Z(n8859) );
  NAND U9127 ( .A(n8818), .B(sreg[463]), .Z(n8822) );
  OR U9128 ( .A(n8820), .B(n8819), .Z(n8821) );
  AND U9129 ( .A(n8822), .B(n8821), .Z(n8858) );
  XOR U9130 ( .A(n8859), .B(n8858), .Z(c[464]) );
  NANDN U9131 ( .A(n8828), .B(n8827), .Z(n8832) );
  NAND U9132 ( .A(n8830), .B(n8829), .Z(n8831) );
  NAND U9133 ( .A(n8832), .B(n8831), .Z(n8893) );
  NANDN U9134 ( .A(n8834), .B(n8833), .Z(n8838) );
  NAND U9135 ( .A(n8836), .B(n8835), .Z(n8837) );
  NAND U9136 ( .A(n8838), .B(n8837), .Z(n8891) );
  XNOR U9137 ( .A(b[7]), .B(a[211]), .Z(n8878) );
  NANDN U9138 ( .A(n8878), .B(n10545), .Z(n8841) );
  NANDN U9139 ( .A(n8839), .B(n10546), .Z(n8840) );
  NAND U9140 ( .A(n8841), .B(n8840), .Z(n8866) );
  XNOR U9141 ( .A(b[3]), .B(a[215]), .Z(n8881) );
  NANDN U9142 ( .A(n8881), .B(n10398), .Z(n8844) );
  NANDN U9143 ( .A(n8842), .B(n10399), .Z(n8843) );
  AND U9144 ( .A(n8844), .B(n8843), .Z(n8867) );
  XNOR U9145 ( .A(n8866), .B(n8867), .Z(n8868) );
  NANDN U9146 ( .A(n527), .B(a[217]), .Z(n8845) );
  XOR U9147 ( .A(n10434), .B(n8845), .Z(n8847) );
  NANDN U9148 ( .A(b[0]), .B(a[216]), .Z(n8846) );
  AND U9149 ( .A(n8847), .B(n8846), .Z(n8874) );
  XOR U9150 ( .A(b[5]), .B(a[213]), .Z(n8887) );
  NAND U9151 ( .A(n8887), .B(n10481), .Z(n8850) );
  NAND U9152 ( .A(n8848), .B(n10482), .Z(n8849) );
  NAND U9153 ( .A(n8850), .B(n8849), .Z(n8872) );
  NANDN U9154 ( .A(n529), .B(a[209]), .Z(n8873) );
  XNOR U9155 ( .A(n8872), .B(n8873), .Z(n8875) );
  XOR U9156 ( .A(n8874), .B(n8875), .Z(n8869) );
  XOR U9157 ( .A(n8868), .B(n8869), .Z(n8890) );
  XOR U9158 ( .A(n8891), .B(n8890), .Z(n8892) );
  XNOR U9159 ( .A(n8893), .B(n8892), .Z(n8862) );
  NAND U9160 ( .A(n8852), .B(n8851), .Z(n8856) );
  NAND U9161 ( .A(n8854), .B(n8853), .Z(n8855) );
  NAND U9162 ( .A(n8856), .B(n8855), .Z(n8863) );
  XNOR U9163 ( .A(n8862), .B(n8863), .Z(n8864) );
  XNOR U9164 ( .A(n8865), .B(n8864), .Z(n8896) );
  XNOR U9165 ( .A(n8896), .B(sreg[465]), .Z(n8898) );
  NAND U9166 ( .A(n8857), .B(sreg[464]), .Z(n8861) );
  OR U9167 ( .A(n8859), .B(n8858), .Z(n8860) );
  AND U9168 ( .A(n8861), .B(n8860), .Z(n8897) );
  XOR U9169 ( .A(n8898), .B(n8897), .Z(c[465]) );
  NANDN U9170 ( .A(n8867), .B(n8866), .Z(n8871) );
  NAND U9171 ( .A(n8869), .B(n8868), .Z(n8870) );
  NAND U9172 ( .A(n8871), .B(n8870), .Z(n8932) );
  NANDN U9173 ( .A(n8873), .B(n8872), .Z(n8877) );
  NAND U9174 ( .A(n8875), .B(n8874), .Z(n8876) );
  NAND U9175 ( .A(n8877), .B(n8876), .Z(n8930) );
  XNOR U9176 ( .A(b[7]), .B(a[212]), .Z(n8917) );
  NANDN U9177 ( .A(n8917), .B(n10545), .Z(n8880) );
  NANDN U9178 ( .A(n8878), .B(n10546), .Z(n8879) );
  NAND U9179 ( .A(n8880), .B(n8879), .Z(n8905) );
  XNOR U9180 ( .A(b[3]), .B(a[216]), .Z(n8920) );
  NANDN U9181 ( .A(n8920), .B(n10398), .Z(n8883) );
  NANDN U9182 ( .A(n8881), .B(n10399), .Z(n8882) );
  AND U9183 ( .A(n8883), .B(n8882), .Z(n8906) );
  XNOR U9184 ( .A(n8905), .B(n8906), .Z(n8907) );
  NANDN U9185 ( .A(n527), .B(a[218]), .Z(n8884) );
  XOR U9186 ( .A(n10434), .B(n8884), .Z(n8886) );
  NANDN U9187 ( .A(b[0]), .B(a[217]), .Z(n8885) );
  AND U9188 ( .A(n8886), .B(n8885), .Z(n8913) );
  XOR U9189 ( .A(b[5]), .B(a[214]), .Z(n8926) );
  NAND U9190 ( .A(n8926), .B(n10481), .Z(n8889) );
  NAND U9191 ( .A(n8887), .B(n10482), .Z(n8888) );
  NAND U9192 ( .A(n8889), .B(n8888), .Z(n8911) );
  NANDN U9193 ( .A(n529), .B(a[210]), .Z(n8912) );
  XNOR U9194 ( .A(n8911), .B(n8912), .Z(n8914) );
  XOR U9195 ( .A(n8913), .B(n8914), .Z(n8908) );
  XOR U9196 ( .A(n8907), .B(n8908), .Z(n8929) );
  XOR U9197 ( .A(n8930), .B(n8929), .Z(n8931) );
  XNOR U9198 ( .A(n8932), .B(n8931), .Z(n8901) );
  NAND U9199 ( .A(n8891), .B(n8890), .Z(n8895) );
  NAND U9200 ( .A(n8893), .B(n8892), .Z(n8894) );
  NAND U9201 ( .A(n8895), .B(n8894), .Z(n8902) );
  XNOR U9202 ( .A(n8901), .B(n8902), .Z(n8903) );
  XNOR U9203 ( .A(n8904), .B(n8903), .Z(n8935) );
  XNOR U9204 ( .A(n8935), .B(sreg[466]), .Z(n8937) );
  NAND U9205 ( .A(n8896), .B(sreg[465]), .Z(n8900) );
  OR U9206 ( .A(n8898), .B(n8897), .Z(n8899) );
  AND U9207 ( .A(n8900), .B(n8899), .Z(n8936) );
  XOR U9208 ( .A(n8937), .B(n8936), .Z(c[466]) );
  NANDN U9209 ( .A(n8906), .B(n8905), .Z(n8910) );
  NAND U9210 ( .A(n8908), .B(n8907), .Z(n8909) );
  NAND U9211 ( .A(n8910), .B(n8909), .Z(n8971) );
  NANDN U9212 ( .A(n8912), .B(n8911), .Z(n8916) );
  NAND U9213 ( .A(n8914), .B(n8913), .Z(n8915) );
  NAND U9214 ( .A(n8916), .B(n8915), .Z(n8969) );
  XNOR U9215 ( .A(b[7]), .B(a[213]), .Z(n8956) );
  NANDN U9216 ( .A(n8956), .B(n10545), .Z(n8919) );
  NANDN U9217 ( .A(n8917), .B(n10546), .Z(n8918) );
  NAND U9218 ( .A(n8919), .B(n8918), .Z(n8944) );
  XNOR U9219 ( .A(b[3]), .B(a[217]), .Z(n8959) );
  NANDN U9220 ( .A(n8959), .B(n10398), .Z(n8922) );
  NANDN U9221 ( .A(n8920), .B(n10399), .Z(n8921) );
  AND U9222 ( .A(n8922), .B(n8921), .Z(n8945) );
  XNOR U9223 ( .A(n8944), .B(n8945), .Z(n8946) );
  NANDN U9224 ( .A(n527), .B(a[219]), .Z(n8923) );
  XOR U9225 ( .A(n10434), .B(n8923), .Z(n8925) );
  NANDN U9226 ( .A(b[0]), .B(a[218]), .Z(n8924) );
  AND U9227 ( .A(n8925), .B(n8924), .Z(n8952) );
  XOR U9228 ( .A(b[5]), .B(a[215]), .Z(n8965) );
  NAND U9229 ( .A(n8965), .B(n10481), .Z(n8928) );
  NAND U9230 ( .A(n8926), .B(n10482), .Z(n8927) );
  NAND U9231 ( .A(n8928), .B(n8927), .Z(n8950) );
  NANDN U9232 ( .A(n529), .B(a[211]), .Z(n8951) );
  XNOR U9233 ( .A(n8950), .B(n8951), .Z(n8953) );
  XOR U9234 ( .A(n8952), .B(n8953), .Z(n8947) );
  XOR U9235 ( .A(n8946), .B(n8947), .Z(n8968) );
  XOR U9236 ( .A(n8969), .B(n8968), .Z(n8970) );
  XNOR U9237 ( .A(n8971), .B(n8970), .Z(n8940) );
  NAND U9238 ( .A(n8930), .B(n8929), .Z(n8934) );
  NAND U9239 ( .A(n8932), .B(n8931), .Z(n8933) );
  NAND U9240 ( .A(n8934), .B(n8933), .Z(n8941) );
  XNOR U9241 ( .A(n8940), .B(n8941), .Z(n8942) );
  XNOR U9242 ( .A(n8943), .B(n8942), .Z(n8974) );
  XNOR U9243 ( .A(n8974), .B(sreg[467]), .Z(n8976) );
  NAND U9244 ( .A(n8935), .B(sreg[466]), .Z(n8939) );
  OR U9245 ( .A(n8937), .B(n8936), .Z(n8938) );
  AND U9246 ( .A(n8939), .B(n8938), .Z(n8975) );
  XOR U9247 ( .A(n8976), .B(n8975), .Z(c[467]) );
  NANDN U9248 ( .A(n8945), .B(n8944), .Z(n8949) );
  NAND U9249 ( .A(n8947), .B(n8946), .Z(n8948) );
  NAND U9250 ( .A(n8949), .B(n8948), .Z(n9010) );
  NANDN U9251 ( .A(n8951), .B(n8950), .Z(n8955) );
  NAND U9252 ( .A(n8953), .B(n8952), .Z(n8954) );
  NAND U9253 ( .A(n8955), .B(n8954), .Z(n9008) );
  XNOR U9254 ( .A(b[7]), .B(a[214]), .Z(n8995) );
  NANDN U9255 ( .A(n8995), .B(n10545), .Z(n8958) );
  NANDN U9256 ( .A(n8956), .B(n10546), .Z(n8957) );
  NAND U9257 ( .A(n8958), .B(n8957), .Z(n8983) );
  XNOR U9258 ( .A(b[3]), .B(a[218]), .Z(n8998) );
  NANDN U9259 ( .A(n8998), .B(n10398), .Z(n8961) );
  NANDN U9260 ( .A(n8959), .B(n10399), .Z(n8960) );
  AND U9261 ( .A(n8961), .B(n8960), .Z(n8984) );
  XNOR U9262 ( .A(n8983), .B(n8984), .Z(n8985) );
  NANDN U9263 ( .A(n527), .B(a[220]), .Z(n8962) );
  XOR U9264 ( .A(n10434), .B(n8962), .Z(n8964) );
  NANDN U9265 ( .A(b[0]), .B(a[219]), .Z(n8963) );
  AND U9266 ( .A(n8964), .B(n8963), .Z(n8991) );
  XOR U9267 ( .A(b[5]), .B(a[216]), .Z(n9004) );
  NAND U9268 ( .A(n9004), .B(n10481), .Z(n8967) );
  NAND U9269 ( .A(n8965), .B(n10482), .Z(n8966) );
  NAND U9270 ( .A(n8967), .B(n8966), .Z(n8989) );
  NANDN U9271 ( .A(n529), .B(a[212]), .Z(n8990) );
  XNOR U9272 ( .A(n8989), .B(n8990), .Z(n8992) );
  XOR U9273 ( .A(n8991), .B(n8992), .Z(n8986) );
  XOR U9274 ( .A(n8985), .B(n8986), .Z(n9007) );
  XOR U9275 ( .A(n9008), .B(n9007), .Z(n9009) );
  XNOR U9276 ( .A(n9010), .B(n9009), .Z(n8979) );
  NAND U9277 ( .A(n8969), .B(n8968), .Z(n8973) );
  NAND U9278 ( .A(n8971), .B(n8970), .Z(n8972) );
  NAND U9279 ( .A(n8973), .B(n8972), .Z(n8980) );
  XNOR U9280 ( .A(n8979), .B(n8980), .Z(n8981) );
  XNOR U9281 ( .A(n8982), .B(n8981), .Z(n9013) );
  XNOR U9282 ( .A(n9013), .B(sreg[468]), .Z(n9015) );
  NAND U9283 ( .A(n8974), .B(sreg[467]), .Z(n8978) );
  OR U9284 ( .A(n8976), .B(n8975), .Z(n8977) );
  AND U9285 ( .A(n8978), .B(n8977), .Z(n9014) );
  XOR U9286 ( .A(n9015), .B(n9014), .Z(c[468]) );
  NANDN U9287 ( .A(n8984), .B(n8983), .Z(n8988) );
  NAND U9288 ( .A(n8986), .B(n8985), .Z(n8987) );
  NAND U9289 ( .A(n8988), .B(n8987), .Z(n9049) );
  NANDN U9290 ( .A(n8990), .B(n8989), .Z(n8994) );
  NAND U9291 ( .A(n8992), .B(n8991), .Z(n8993) );
  NAND U9292 ( .A(n8994), .B(n8993), .Z(n9047) );
  XNOR U9293 ( .A(b[7]), .B(a[215]), .Z(n9034) );
  NANDN U9294 ( .A(n9034), .B(n10545), .Z(n8997) );
  NANDN U9295 ( .A(n8995), .B(n10546), .Z(n8996) );
  NAND U9296 ( .A(n8997), .B(n8996), .Z(n9022) );
  XNOR U9297 ( .A(b[3]), .B(a[219]), .Z(n9037) );
  NANDN U9298 ( .A(n9037), .B(n10398), .Z(n9000) );
  NANDN U9299 ( .A(n8998), .B(n10399), .Z(n8999) );
  AND U9300 ( .A(n9000), .B(n8999), .Z(n9023) );
  XNOR U9301 ( .A(n9022), .B(n9023), .Z(n9024) );
  NANDN U9302 ( .A(n527), .B(a[221]), .Z(n9001) );
  XOR U9303 ( .A(n10434), .B(n9001), .Z(n9003) );
  NANDN U9304 ( .A(b[0]), .B(a[220]), .Z(n9002) );
  AND U9305 ( .A(n9003), .B(n9002), .Z(n9030) );
  XOR U9306 ( .A(b[5]), .B(a[217]), .Z(n9043) );
  NAND U9307 ( .A(n9043), .B(n10481), .Z(n9006) );
  NAND U9308 ( .A(n9004), .B(n10482), .Z(n9005) );
  NAND U9309 ( .A(n9006), .B(n9005), .Z(n9028) );
  NANDN U9310 ( .A(n529), .B(a[213]), .Z(n9029) );
  XNOR U9311 ( .A(n9028), .B(n9029), .Z(n9031) );
  XOR U9312 ( .A(n9030), .B(n9031), .Z(n9025) );
  XOR U9313 ( .A(n9024), .B(n9025), .Z(n9046) );
  XOR U9314 ( .A(n9047), .B(n9046), .Z(n9048) );
  XNOR U9315 ( .A(n9049), .B(n9048), .Z(n9018) );
  NAND U9316 ( .A(n9008), .B(n9007), .Z(n9012) );
  NAND U9317 ( .A(n9010), .B(n9009), .Z(n9011) );
  NAND U9318 ( .A(n9012), .B(n9011), .Z(n9019) );
  XNOR U9319 ( .A(n9018), .B(n9019), .Z(n9020) );
  XNOR U9320 ( .A(n9021), .B(n9020), .Z(n9052) );
  XNOR U9321 ( .A(n9052), .B(sreg[469]), .Z(n9054) );
  NAND U9322 ( .A(n9013), .B(sreg[468]), .Z(n9017) );
  OR U9323 ( .A(n9015), .B(n9014), .Z(n9016) );
  AND U9324 ( .A(n9017), .B(n9016), .Z(n9053) );
  XOR U9325 ( .A(n9054), .B(n9053), .Z(c[469]) );
  NANDN U9326 ( .A(n9023), .B(n9022), .Z(n9027) );
  NAND U9327 ( .A(n9025), .B(n9024), .Z(n9026) );
  NAND U9328 ( .A(n9027), .B(n9026), .Z(n9088) );
  NANDN U9329 ( .A(n9029), .B(n9028), .Z(n9033) );
  NAND U9330 ( .A(n9031), .B(n9030), .Z(n9032) );
  NAND U9331 ( .A(n9033), .B(n9032), .Z(n9086) );
  XNOR U9332 ( .A(b[7]), .B(a[216]), .Z(n9079) );
  NANDN U9333 ( .A(n9079), .B(n10545), .Z(n9036) );
  NANDN U9334 ( .A(n9034), .B(n10546), .Z(n9035) );
  NAND U9335 ( .A(n9036), .B(n9035), .Z(n9061) );
  XNOR U9336 ( .A(b[3]), .B(a[220]), .Z(n9082) );
  NANDN U9337 ( .A(n9082), .B(n10398), .Z(n9039) );
  NANDN U9338 ( .A(n9037), .B(n10399), .Z(n9038) );
  AND U9339 ( .A(n9039), .B(n9038), .Z(n9062) );
  XNOR U9340 ( .A(n9061), .B(n9062), .Z(n9063) );
  NANDN U9341 ( .A(n527), .B(a[222]), .Z(n9040) );
  XOR U9342 ( .A(n10434), .B(n9040), .Z(n9042) );
  NANDN U9343 ( .A(b[0]), .B(a[221]), .Z(n9041) );
  AND U9344 ( .A(n9042), .B(n9041), .Z(n9069) );
  XOR U9345 ( .A(b[5]), .B(a[218]), .Z(n9076) );
  NAND U9346 ( .A(n9076), .B(n10481), .Z(n9045) );
  NAND U9347 ( .A(n9043), .B(n10482), .Z(n9044) );
  NAND U9348 ( .A(n9045), .B(n9044), .Z(n9067) );
  NANDN U9349 ( .A(n529), .B(a[214]), .Z(n9068) );
  XNOR U9350 ( .A(n9067), .B(n9068), .Z(n9070) );
  XOR U9351 ( .A(n9069), .B(n9070), .Z(n9064) );
  XOR U9352 ( .A(n9063), .B(n9064), .Z(n9085) );
  XOR U9353 ( .A(n9086), .B(n9085), .Z(n9087) );
  XNOR U9354 ( .A(n9088), .B(n9087), .Z(n9057) );
  NAND U9355 ( .A(n9047), .B(n9046), .Z(n9051) );
  NAND U9356 ( .A(n9049), .B(n9048), .Z(n9050) );
  NAND U9357 ( .A(n9051), .B(n9050), .Z(n9058) );
  XNOR U9358 ( .A(n9057), .B(n9058), .Z(n9059) );
  XNOR U9359 ( .A(n9060), .B(n9059), .Z(n9091) );
  XNOR U9360 ( .A(n9091), .B(sreg[470]), .Z(n9093) );
  NAND U9361 ( .A(n9052), .B(sreg[469]), .Z(n9056) );
  OR U9362 ( .A(n9054), .B(n9053), .Z(n9055) );
  AND U9363 ( .A(n9056), .B(n9055), .Z(n9092) );
  XOR U9364 ( .A(n9093), .B(n9092), .Z(c[470]) );
  NANDN U9365 ( .A(n9062), .B(n9061), .Z(n9066) );
  NAND U9366 ( .A(n9064), .B(n9063), .Z(n9065) );
  NAND U9367 ( .A(n9066), .B(n9065), .Z(n9127) );
  NANDN U9368 ( .A(n9068), .B(n9067), .Z(n9072) );
  NAND U9369 ( .A(n9070), .B(n9069), .Z(n9071) );
  NAND U9370 ( .A(n9072), .B(n9071), .Z(n9125) );
  NANDN U9371 ( .A(n527), .B(a[223]), .Z(n9073) );
  XOR U9372 ( .A(n10434), .B(n9073), .Z(n9075) );
  NANDN U9373 ( .A(b[0]), .B(a[222]), .Z(n9074) );
  AND U9374 ( .A(n9075), .B(n9074), .Z(n9108) );
  XOR U9375 ( .A(b[5]), .B(a[219]), .Z(n9121) );
  NAND U9376 ( .A(n9121), .B(n10481), .Z(n9078) );
  NAND U9377 ( .A(n9076), .B(n10482), .Z(n9077) );
  NAND U9378 ( .A(n9078), .B(n9077), .Z(n9106) );
  NANDN U9379 ( .A(n529), .B(a[215]), .Z(n9107) );
  XNOR U9380 ( .A(n9106), .B(n9107), .Z(n9109) );
  XOR U9381 ( .A(n9108), .B(n9109), .Z(n9102) );
  XNOR U9382 ( .A(b[7]), .B(a[217]), .Z(n9112) );
  NANDN U9383 ( .A(n9112), .B(n10545), .Z(n9081) );
  NANDN U9384 ( .A(n9079), .B(n10546), .Z(n9080) );
  NAND U9385 ( .A(n9081), .B(n9080), .Z(n9100) );
  XNOR U9386 ( .A(b[3]), .B(a[221]), .Z(n9115) );
  NANDN U9387 ( .A(n9115), .B(n10398), .Z(n9084) );
  NANDN U9388 ( .A(n9082), .B(n10399), .Z(n9083) );
  AND U9389 ( .A(n9084), .B(n9083), .Z(n9101) );
  XNOR U9390 ( .A(n9100), .B(n9101), .Z(n9103) );
  XOR U9391 ( .A(n9102), .B(n9103), .Z(n9124) );
  XOR U9392 ( .A(n9125), .B(n9124), .Z(n9126) );
  XNOR U9393 ( .A(n9127), .B(n9126), .Z(n9096) );
  NAND U9394 ( .A(n9086), .B(n9085), .Z(n9090) );
  NAND U9395 ( .A(n9088), .B(n9087), .Z(n9089) );
  NAND U9396 ( .A(n9090), .B(n9089), .Z(n9097) );
  XNOR U9397 ( .A(n9096), .B(n9097), .Z(n9098) );
  XNOR U9398 ( .A(n9099), .B(n9098), .Z(n9130) );
  XNOR U9399 ( .A(n9130), .B(sreg[471]), .Z(n9132) );
  NAND U9400 ( .A(n9091), .B(sreg[470]), .Z(n9095) );
  OR U9401 ( .A(n9093), .B(n9092), .Z(n9094) );
  AND U9402 ( .A(n9095), .B(n9094), .Z(n9131) );
  XOR U9403 ( .A(n9132), .B(n9131), .Z(c[471]) );
  NANDN U9404 ( .A(n9101), .B(n9100), .Z(n9105) );
  NAND U9405 ( .A(n9103), .B(n9102), .Z(n9104) );
  NAND U9406 ( .A(n9105), .B(n9104), .Z(n9166) );
  NANDN U9407 ( .A(n9107), .B(n9106), .Z(n9111) );
  NAND U9408 ( .A(n9109), .B(n9108), .Z(n9110) );
  NAND U9409 ( .A(n9111), .B(n9110), .Z(n9164) );
  XNOR U9410 ( .A(b[7]), .B(a[218]), .Z(n9151) );
  NANDN U9411 ( .A(n9151), .B(n10545), .Z(n9114) );
  NANDN U9412 ( .A(n9112), .B(n10546), .Z(n9113) );
  NAND U9413 ( .A(n9114), .B(n9113), .Z(n9139) );
  XNOR U9414 ( .A(b[3]), .B(a[222]), .Z(n9154) );
  NANDN U9415 ( .A(n9154), .B(n10398), .Z(n9117) );
  NANDN U9416 ( .A(n9115), .B(n10399), .Z(n9116) );
  AND U9417 ( .A(n9117), .B(n9116), .Z(n9140) );
  XNOR U9418 ( .A(n9139), .B(n9140), .Z(n9141) );
  NANDN U9419 ( .A(n527), .B(a[224]), .Z(n9118) );
  XOR U9420 ( .A(n10434), .B(n9118), .Z(n9120) );
  NANDN U9421 ( .A(b[0]), .B(a[223]), .Z(n9119) );
  AND U9422 ( .A(n9120), .B(n9119), .Z(n9147) );
  XOR U9423 ( .A(b[5]), .B(a[220]), .Z(n9160) );
  NAND U9424 ( .A(n9160), .B(n10481), .Z(n9123) );
  NAND U9425 ( .A(n9121), .B(n10482), .Z(n9122) );
  NAND U9426 ( .A(n9123), .B(n9122), .Z(n9145) );
  NANDN U9427 ( .A(n529), .B(a[216]), .Z(n9146) );
  XNOR U9428 ( .A(n9145), .B(n9146), .Z(n9148) );
  XOR U9429 ( .A(n9147), .B(n9148), .Z(n9142) );
  XOR U9430 ( .A(n9141), .B(n9142), .Z(n9163) );
  XOR U9431 ( .A(n9164), .B(n9163), .Z(n9165) );
  XNOR U9432 ( .A(n9166), .B(n9165), .Z(n9135) );
  NAND U9433 ( .A(n9125), .B(n9124), .Z(n9129) );
  NAND U9434 ( .A(n9127), .B(n9126), .Z(n9128) );
  NAND U9435 ( .A(n9129), .B(n9128), .Z(n9136) );
  XNOR U9436 ( .A(n9135), .B(n9136), .Z(n9137) );
  XNOR U9437 ( .A(n9138), .B(n9137), .Z(n9169) );
  XNOR U9438 ( .A(n9169), .B(sreg[472]), .Z(n9171) );
  NAND U9439 ( .A(n9130), .B(sreg[471]), .Z(n9134) );
  OR U9440 ( .A(n9132), .B(n9131), .Z(n9133) );
  AND U9441 ( .A(n9134), .B(n9133), .Z(n9170) );
  XOR U9442 ( .A(n9171), .B(n9170), .Z(c[472]) );
  NANDN U9443 ( .A(n9140), .B(n9139), .Z(n9144) );
  NAND U9444 ( .A(n9142), .B(n9141), .Z(n9143) );
  NAND U9445 ( .A(n9144), .B(n9143), .Z(n9205) );
  NANDN U9446 ( .A(n9146), .B(n9145), .Z(n9150) );
  NAND U9447 ( .A(n9148), .B(n9147), .Z(n9149) );
  NAND U9448 ( .A(n9150), .B(n9149), .Z(n9203) );
  XNOR U9449 ( .A(b[7]), .B(a[219]), .Z(n9190) );
  NANDN U9450 ( .A(n9190), .B(n10545), .Z(n9153) );
  NANDN U9451 ( .A(n9151), .B(n10546), .Z(n9152) );
  NAND U9452 ( .A(n9153), .B(n9152), .Z(n9178) );
  XNOR U9453 ( .A(b[3]), .B(a[223]), .Z(n9193) );
  NANDN U9454 ( .A(n9193), .B(n10398), .Z(n9156) );
  NANDN U9455 ( .A(n9154), .B(n10399), .Z(n9155) );
  AND U9456 ( .A(n9156), .B(n9155), .Z(n9179) );
  XNOR U9457 ( .A(n9178), .B(n9179), .Z(n9180) );
  NANDN U9458 ( .A(n527), .B(a[225]), .Z(n9157) );
  XOR U9459 ( .A(n10434), .B(n9157), .Z(n9159) );
  NANDN U9460 ( .A(b[0]), .B(a[224]), .Z(n9158) );
  AND U9461 ( .A(n9159), .B(n9158), .Z(n9186) );
  XOR U9462 ( .A(b[5]), .B(a[221]), .Z(n9199) );
  NAND U9463 ( .A(n9199), .B(n10481), .Z(n9162) );
  NAND U9464 ( .A(n9160), .B(n10482), .Z(n9161) );
  NAND U9465 ( .A(n9162), .B(n9161), .Z(n9184) );
  NANDN U9466 ( .A(n529), .B(a[217]), .Z(n9185) );
  XNOR U9467 ( .A(n9184), .B(n9185), .Z(n9187) );
  XOR U9468 ( .A(n9186), .B(n9187), .Z(n9181) );
  XOR U9469 ( .A(n9180), .B(n9181), .Z(n9202) );
  XOR U9470 ( .A(n9203), .B(n9202), .Z(n9204) );
  XNOR U9471 ( .A(n9205), .B(n9204), .Z(n9174) );
  NAND U9472 ( .A(n9164), .B(n9163), .Z(n9168) );
  NAND U9473 ( .A(n9166), .B(n9165), .Z(n9167) );
  NAND U9474 ( .A(n9168), .B(n9167), .Z(n9175) );
  XNOR U9475 ( .A(n9174), .B(n9175), .Z(n9176) );
  XNOR U9476 ( .A(n9177), .B(n9176), .Z(n9208) );
  XNOR U9477 ( .A(n9208), .B(sreg[473]), .Z(n9210) );
  NAND U9478 ( .A(n9169), .B(sreg[472]), .Z(n9173) );
  OR U9479 ( .A(n9171), .B(n9170), .Z(n9172) );
  AND U9480 ( .A(n9173), .B(n9172), .Z(n9209) );
  XOR U9481 ( .A(n9210), .B(n9209), .Z(c[473]) );
  NANDN U9482 ( .A(n9179), .B(n9178), .Z(n9183) );
  NAND U9483 ( .A(n9181), .B(n9180), .Z(n9182) );
  NAND U9484 ( .A(n9183), .B(n9182), .Z(n9244) );
  NANDN U9485 ( .A(n9185), .B(n9184), .Z(n9189) );
  NAND U9486 ( .A(n9187), .B(n9186), .Z(n9188) );
  NAND U9487 ( .A(n9189), .B(n9188), .Z(n9242) );
  XNOR U9488 ( .A(b[7]), .B(a[220]), .Z(n9229) );
  NANDN U9489 ( .A(n9229), .B(n10545), .Z(n9192) );
  NANDN U9490 ( .A(n9190), .B(n10546), .Z(n9191) );
  NAND U9491 ( .A(n9192), .B(n9191), .Z(n9217) );
  XNOR U9492 ( .A(b[3]), .B(a[224]), .Z(n9232) );
  NANDN U9493 ( .A(n9232), .B(n10398), .Z(n9195) );
  NANDN U9494 ( .A(n9193), .B(n10399), .Z(n9194) );
  AND U9495 ( .A(n9195), .B(n9194), .Z(n9218) );
  XNOR U9496 ( .A(n9217), .B(n9218), .Z(n9219) );
  NANDN U9497 ( .A(n527), .B(a[226]), .Z(n9196) );
  XOR U9498 ( .A(n10434), .B(n9196), .Z(n9198) );
  NANDN U9499 ( .A(b[0]), .B(a[225]), .Z(n9197) );
  AND U9500 ( .A(n9198), .B(n9197), .Z(n9225) );
  XOR U9501 ( .A(b[5]), .B(a[222]), .Z(n9238) );
  NAND U9502 ( .A(n9238), .B(n10481), .Z(n9201) );
  NAND U9503 ( .A(n9199), .B(n10482), .Z(n9200) );
  NAND U9504 ( .A(n9201), .B(n9200), .Z(n9223) );
  NANDN U9505 ( .A(n529), .B(a[218]), .Z(n9224) );
  XNOR U9506 ( .A(n9223), .B(n9224), .Z(n9226) );
  XOR U9507 ( .A(n9225), .B(n9226), .Z(n9220) );
  XOR U9508 ( .A(n9219), .B(n9220), .Z(n9241) );
  XOR U9509 ( .A(n9242), .B(n9241), .Z(n9243) );
  XNOR U9510 ( .A(n9244), .B(n9243), .Z(n9213) );
  NAND U9511 ( .A(n9203), .B(n9202), .Z(n9207) );
  NAND U9512 ( .A(n9205), .B(n9204), .Z(n9206) );
  NAND U9513 ( .A(n9207), .B(n9206), .Z(n9214) );
  XNOR U9514 ( .A(n9213), .B(n9214), .Z(n9215) );
  XNOR U9515 ( .A(n9216), .B(n9215), .Z(n9247) );
  XNOR U9516 ( .A(n9247), .B(sreg[474]), .Z(n9249) );
  NAND U9517 ( .A(n9208), .B(sreg[473]), .Z(n9212) );
  OR U9518 ( .A(n9210), .B(n9209), .Z(n9211) );
  AND U9519 ( .A(n9212), .B(n9211), .Z(n9248) );
  XOR U9520 ( .A(n9249), .B(n9248), .Z(c[474]) );
  NANDN U9521 ( .A(n9218), .B(n9217), .Z(n9222) );
  NAND U9522 ( .A(n9220), .B(n9219), .Z(n9221) );
  NAND U9523 ( .A(n9222), .B(n9221), .Z(n9283) );
  NANDN U9524 ( .A(n9224), .B(n9223), .Z(n9228) );
  NAND U9525 ( .A(n9226), .B(n9225), .Z(n9227) );
  NAND U9526 ( .A(n9228), .B(n9227), .Z(n9281) );
  XNOR U9527 ( .A(b[7]), .B(a[221]), .Z(n9274) );
  NANDN U9528 ( .A(n9274), .B(n10545), .Z(n9231) );
  NANDN U9529 ( .A(n9229), .B(n10546), .Z(n9230) );
  NAND U9530 ( .A(n9231), .B(n9230), .Z(n9256) );
  XNOR U9531 ( .A(b[3]), .B(a[225]), .Z(n9277) );
  NANDN U9532 ( .A(n9277), .B(n10398), .Z(n9234) );
  NANDN U9533 ( .A(n9232), .B(n10399), .Z(n9233) );
  AND U9534 ( .A(n9234), .B(n9233), .Z(n9257) );
  XNOR U9535 ( .A(n9256), .B(n9257), .Z(n9258) );
  NANDN U9536 ( .A(n527), .B(a[227]), .Z(n9235) );
  XOR U9537 ( .A(n10434), .B(n9235), .Z(n9237) );
  NANDN U9538 ( .A(b[0]), .B(a[226]), .Z(n9236) );
  AND U9539 ( .A(n9237), .B(n9236), .Z(n9264) );
  XOR U9540 ( .A(b[5]), .B(a[223]), .Z(n9271) );
  NAND U9541 ( .A(n9271), .B(n10481), .Z(n9240) );
  NAND U9542 ( .A(n9238), .B(n10482), .Z(n9239) );
  NAND U9543 ( .A(n9240), .B(n9239), .Z(n9262) );
  NANDN U9544 ( .A(n529), .B(a[219]), .Z(n9263) );
  XNOR U9545 ( .A(n9262), .B(n9263), .Z(n9265) );
  XOR U9546 ( .A(n9264), .B(n9265), .Z(n9259) );
  XOR U9547 ( .A(n9258), .B(n9259), .Z(n9280) );
  XOR U9548 ( .A(n9281), .B(n9280), .Z(n9282) );
  XNOR U9549 ( .A(n9283), .B(n9282), .Z(n9252) );
  NAND U9550 ( .A(n9242), .B(n9241), .Z(n9246) );
  NAND U9551 ( .A(n9244), .B(n9243), .Z(n9245) );
  NAND U9552 ( .A(n9246), .B(n9245), .Z(n9253) );
  XNOR U9553 ( .A(n9252), .B(n9253), .Z(n9254) );
  XNOR U9554 ( .A(n9255), .B(n9254), .Z(n9286) );
  XNOR U9555 ( .A(n9286), .B(sreg[475]), .Z(n9288) );
  NAND U9556 ( .A(n9247), .B(sreg[474]), .Z(n9251) );
  OR U9557 ( .A(n9249), .B(n9248), .Z(n9250) );
  AND U9558 ( .A(n9251), .B(n9250), .Z(n9287) );
  XOR U9559 ( .A(n9288), .B(n9287), .Z(c[475]) );
  NANDN U9560 ( .A(n9257), .B(n9256), .Z(n9261) );
  NAND U9561 ( .A(n9259), .B(n9258), .Z(n9260) );
  NAND U9562 ( .A(n9261), .B(n9260), .Z(n9322) );
  NANDN U9563 ( .A(n9263), .B(n9262), .Z(n9267) );
  NAND U9564 ( .A(n9265), .B(n9264), .Z(n9266) );
  NAND U9565 ( .A(n9267), .B(n9266), .Z(n9320) );
  NANDN U9566 ( .A(n527), .B(a[228]), .Z(n9268) );
  XOR U9567 ( .A(n10434), .B(n9268), .Z(n9270) );
  NANDN U9568 ( .A(b[0]), .B(a[227]), .Z(n9269) );
  AND U9569 ( .A(n9270), .B(n9269), .Z(n9303) );
  XOR U9570 ( .A(b[5]), .B(a[224]), .Z(n9316) );
  NAND U9571 ( .A(n9316), .B(n10481), .Z(n9273) );
  NAND U9572 ( .A(n9271), .B(n10482), .Z(n9272) );
  NAND U9573 ( .A(n9273), .B(n9272), .Z(n9301) );
  NANDN U9574 ( .A(n529), .B(a[220]), .Z(n9302) );
  XNOR U9575 ( .A(n9301), .B(n9302), .Z(n9304) );
  XOR U9576 ( .A(n9303), .B(n9304), .Z(n9297) );
  XNOR U9577 ( .A(b[7]), .B(a[222]), .Z(n9307) );
  NANDN U9578 ( .A(n9307), .B(n10545), .Z(n9276) );
  NANDN U9579 ( .A(n9274), .B(n10546), .Z(n9275) );
  NAND U9580 ( .A(n9276), .B(n9275), .Z(n9295) );
  XNOR U9581 ( .A(b[3]), .B(a[226]), .Z(n9310) );
  NANDN U9582 ( .A(n9310), .B(n10398), .Z(n9279) );
  NANDN U9583 ( .A(n9277), .B(n10399), .Z(n9278) );
  AND U9584 ( .A(n9279), .B(n9278), .Z(n9296) );
  XNOR U9585 ( .A(n9295), .B(n9296), .Z(n9298) );
  XOR U9586 ( .A(n9297), .B(n9298), .Z(n9319) );
  XOR U9587 ( .A(n9320), .B(n9319), .Z(n9321) );
  XNOR U9588 ( .A(n9322), .B(n9321), .Z(n9291) );
  NAND U9589 ( .A(n9281), .B(n9280), .Z(n9285) );
  NAND U9590 ( .A(n9283), .B(n9282), .Z(n9284) );
  NAND U9591 ( .A(n9285), .B(n9284), .Z(n9292) );
  XNOR U9592 ( .A(n9291), .B(n9292), .Z(n9293) );
  XNOR U9593 ( .A(n9294), .B(n9293), .Z(n9325) );
  XNOR U9594 ( .A(n9325), .B(sreg[476]), .Z(n9327) );
  NAND U9595 ( .A(n9286), .B(sreg[475]), .Z(n9290) );
  OR U9596 ( .A(n9288), .B(n9287), .Z(n9289) );
  AND U9597 ( .A(n9290), .B(n9289), .Z(n9326) );
  XOR U9598 ( .A(n9327), .B(n9326), .Z(c[476]) );
  NANDN U9599 ( .A(n9296), .B(n9295), .Z(n9300) );
  NAND U9600 ( .A(n9298), .B(n9297), .Z(n9299) );
  NAND U9601 ( .A(n9300), .B(n9299), .Z(n9361) );
  NANDN U9602 ( .A(n9302), .B(n9301), .Z(n9306) );
  NAND U9603 ( .A(n9304), .B(n9303), .Z(n9305) );
  NAND U9604 ( .A(n9306), .B(n9305), .Z(n9359) );
  XNOR U9605 ( .A(b[7]), .B(a[223]), .Z(n9346) );
  NANDN U9606 ( .A(n9346), .B(n10545), .Z(n9309) );
  NANDN U9607 ( .A(n9307), .B(n10546), .Z(n9308) );
  NAND U9608 ( .A(n9309), .B(n9308), .Z(n9334) );
  XNOR U9609 ( .A(b[3]), .B(a[227]), .Z(n9349) );
  NANDN U9610 ( .A(n9349), .B(n10398), .Z(n9312) );
  NANDN U9611 ( .A(n9310), .B(n10399), .Z(n9311) );
  AND U9612 ( .A(n9312), .B(n9311), .Z(n9335) );
  XNOR U9613 ( .A(n9334), .B(n9335), .Z(n9336) );
  NANDN U9614 ( .A(n527), .B(a[229]), .Z(n9313) );
  XOR U9615 ( .A(n10434), .B(n9313), .Z(n9315) );
  NANDN U9616 ( .A(b[0]), .B(a[228]), .Z(n9314) );
  AND U9617 ( .A(n9315), .B(n9314), .Z(n9342) );
  XOR U9618 ( .A(b[5]), .B(a[225]), .Z(n9355) );
  NAND U9619 ( .A(n9355), .B(n10481), .Z(n9318) );
  NAND U9620 ( .A(n9316), .B(n10482), .Z(n9317) );
  NAND U9621 ( .A(n9318), .B(n9317), .Z(n9340) );
  NANDN U9622 ( .A(n529), .B(a[221]), .Z(n9341) );
  XNOR U9623 ( .A(n9340), .B(n9341), .Z(n9343) );
  XOR U9624 ( .A(n9342), .B(n9343), .Z(n9337) );
  XOR U9625 ( .A(n9336), .B(n9337), .Z(n9358) );
  XOR U9626 ( .A(n9359), .B(n9358), .Z(n9360) );
  XNOR U9627 ( .A(n9361), .B(n9360), .Z(n9330) );
  NAND U9628 ( .A(n9320), .B(n9319), .Z(n9324) );
  NAND U9629 ( .A(n9322), .B(n9321), .Z(n9323) );
  NAND U9630 ( .A(n9324), .B(n9323), .Z(n9331) );
  XNOR U9631 ( .A(n9330), .B(n9331), .Z(n9332) );
  XNOR U9632 ( .A(n9333), .B(n9332), .Z(n9364) );
  XNOR U9633 ( .A(n9364), .B(sreg[477]), .Z(n9366) );
  NAND U9634 ( .A(n9325), .B(sreg[476]), .Z(n9329) );
  OR U9635 ( .A(n9327), .B(n9326), .Z(n9328) );
  AND U9636 ( .A(n9329), .B(n9328), .Z(n9365) );
  XOR U9637 ( .A(n9366), .B(n9365), .Z(c[477]) );
  NANDN U9638 ( .A(n9335), .B(n9334), .Z(n9339) );
  NAND U9639 ( .A(n9337), .B(n9336), .Z(n9338) );
  NAND U9640 ( .A(n9339), .B(n9338), .Z(n9400) );
  NANDN U9641 ( .A(n9341), .B(n9340), .Z(n9345) );
  NAND U9642 ( .A(n9343), .B(n9342), .Z(n9344) );
  NAND U9643 ( .A(n9345), .B(n9344), .Z(n9398) );
  XNOR U9644 ( .A(b[7]), .B(a[224]), .Z(n9385) );
  NANDN U9645 ( .A(n9385), .B(n10545), .Z(n9348) );
  NANDN U9646 ( .A(n9346), .B(n10546), .Z(n9347) );
  NAND U9647 ( .A(n9348), .B(n9347), .Z(n9373) );
  XNOR U9648 ( .A(b[3]), .B(a[228]), .Z(n9388) );
  NANDN U9649 ( .A(n9388), .B(n10398), .Z(n9351) );
  NANDN U9650 ( .A(n9349), .B(n10399), .Z(n9350) );
  AND U9651 ( .A(n9351), .B(n9350), .Z(n9374) );
  XNOR U9652 ( .A(n9373), .B(n9374), .Z(n9375) );
  NANDN U9653 ( .A(n527), .B(a[230]), .Z(n9352) );
  XOR U9654 ( .A(n10434), .B(n9352), .Z(n9354) );
  NANDN U9655 ( .A(b[0]), .B(a[229]), .Z(n9353) );
  AND U9656 ( .A(n9354), .B(n9353), .Z(n9381) );
  XOR U9657 ( .A(b[5]), .B(a[226]), .Z(n9394) );
  NAND U9658 ( .A(n9394), .B(n10481), .Z(n9357) );
  NAND U9659 ( .A(n9355), .B(n10482), .Z(n9356) );
  NAND U9660 ( .A(n9357), .B(n9356), .Z(n9379) );
  NANDN U9661 ( .A(n529), .B(a[222]), .Z(n9380) );
  XNOR U9662 ( .A(n9379), .B(n9380), .Z(n9382) );
  XOR U9663 ( .A(n9381), .B(n9382), .Z(n9376) );
  XOR U9664 ( .A(n9375), .B(n9376), .Z(n9397) );
  XOR U9665 ( .A(n9398), .B(n9397), .Z(n9399) );
  XNOR U9666 ( .A(n9400), .B(n9399), .Z(n9369) );
  NAND U9667 ( .A(n9359), .B(n9358), .Z(n9363) );
  NAND U9668 ( .A(n9361), .B(n9360), .Z(n9362) );
  NAND U9669 ( .A(n9363), .B(n9362), .Z(n9370) );
  XNOR U9670 ( .A(n9369), .B(n9370), .Z(n9371) );
  XNOR U9671 ( .A(n9372), .B(n9371), .Z(n9403) );
  XNOR U9672 ( .A(n9403), .B(sreg[478]), .Z(n9405) );
  NAND U9673 ( .A(n9364), .B(sreg[477]), .Z(n9368) );
  OR U9674 ( .A(n9366), .B(n9365), .Z(n9367) );
  AND U9675 ( .A(n9368), .B(n9367), .Z(n9404) );
  XOR U9676 ( .A(n9405), .B(n9404), .Z(c[478]) );
  NANDN U9677 ( .A(n9374), .B(n9373), .Z(n9378) );
  NAND U9678 ( .A(n9376), .B(n9375), .Z(n9377) );
  NAND U9679 ( .A(n9378), .B(n9377), .Z(n9439) );
  NANDN U9680 ( .A(n9380), .B(n9379), .Z(n9384) );
  NAND U9681 ( .A(n9382), .B(n9381), .Z(n9383) );
  NAND U9682 ( .A(n9384), .B(n9383), .Z(n9437) );
  XNOR U9683 ( .A(b[7]), .B(a[225]), .Z(n9424) );
  NANDN U9684 ( .A(n9424), .B(n10545), .Z(n9387) );
  NANDN U9685 ( .A(n9385), .B(n10546), .Z(n9386) );
  NAND U9686 ( .A(n9387), .B(n9386), .Z(n9412) );
  XNOR U9687 ( .A(b[3]), .B(a[229]), .Z(n9427) );
  NANDN U9688 ( .A(n9427), .B(n10398), .Z(n9390) );
  NANDN U9689 ( .A(n9388), .B(n10399), .Z(n9389) );
  AND U9690 ( .A(n9390), .B(n9389), .Z(n9413) );
  XNOR U9691 ( .A(n9412), .B(n9413), .Z(n9414) );
  NANDN U9692 ( .A(n527), .B(a[231]), .Z(n9391) );
  XOR U9693 ( .A(n10434), .B(n9391), .Z(n9393) );
  NANDN U9694 ( .A(b[0]), .B(a[230]), .Z(n9392) );
  AND U9695 ( .A(n9393), .B(n9392), .Z(n9420) );
  XOR U9696 ( .A(b[5]), .B(a[227]), .Z(n9433) );
  NAND U9697 ( .A(n9433), .B(n10481), .Z(n9396) );
  NAND U9698 ( .A(n9394), .B(n10482), .Z(n9395) );
  NAND U9699 ( .A(n9396), .B(n9395), .Z(n9418) );
  NANDN U9700 ( .A(n529), .B(a[223]), .Z(n9419) );
  XNOR U9701 ( .A(n9418), .B(n9419), .Z(n9421) );
  XOR U9702 ( .A(n9420), .B(n9421), .Z(n9415) );
  XOR U9703 ( .A(n9414), .B(n9415), .Z(n9436) );
  XOR U9704 ( .A(n9437), .B(n9436), .Z(n9438) );
  XNOR U9705 ( .A(n9439), .B(n9438), .Z(n9408) );
  NAND U9706 ( .A(n9398), .B(n9397), .Z(n9402) );
  NAND U9707 ( .A(n9400), .B(n9399), .Z(n9401) );
  NAND U9708 ( .A(n9402), .B(n9401), .Z(n9409) );
  XNOR U9709 ( .A(n9408), .B(n9409), .Z(n9410) );
  XNOR U9710 ( .A(n9411), .B(n9410), .Z(n9442) );
  XNOR U9711 ( .A(n9442), .B(sreg[479]), .Z(n9444) );
  NAND U9712 ( .A(n9403), .B(sreg[478]), .Z(n9407) );
  OR U9713 ( .A(n9405), .B(n9404), .Z(n9406) );
  AND U9714 ( .A(n9407), .B(n9406), .Z(n9443) );
  XOR U9715 ( .A(n9444), .B(n9443), .Z(c[479]) );
  NANDN U9716 ( .A(n9413), .B(n9412), .Z(n9417) );
  NAND U9717 ( .A(n9415), .B(n9414), .Z(n9416) );
  NAND U9718 ( .A(n9417), .B(n9416), .Z(n9478) );
  NANDN U9719 ( .A(n9419), .B(n9418), .Z(n9423) );
  NAND U9720 ( .A(n9421), .B(n9420), .Z(n9422) );
  NAND U9721 ( .A(n9423), .B(n9422), .Z(n9476) );
  XNOR U9722 ( .A(b[7]), .B(a[226]), .Z(n9463) );
  NANDN U9723 ( .A(n9463), .B(n10545), .Z(n9426) );
  NANDN U9724 ( .A(n9424), .B(n10546), .Z(n9425) );
  NAND U9725 ( .A(n9426), .B(n9425), .Z(n9451) );
  XNOR U9726 ( .A(b[3]), .B(a[230]), .Z(n9466) );
  NANDN U9727 ( .A(n9466), .B(n10398), .Z(n9429) );
  NANDN U9728 ( .A(n9427), .B(n10399), .Z(n9428) );
  AND U9729 ( .A(n9429), .B(n9428), .Z(n9452) );
  XNOR U9730 ( .A(n9451), .B(n9452), .Z(n9453) );
  NANDN U9731 ( .A(n527), .B(a[232]), .Z(n9430) );
  XOR U9732 ( .A(n10434), .B(n9430), .Z(n9432) );
  NANDN U9733 ( .A(b[0]), .B(a[231]), .Z(n9431) );
  AND U9734 ( .A(n9432), .B(n9431), .Z(n9459) );
  XOR U9735 ( .A(b[5]), .B(a[228]), .Z(n9472) );
  NAND U9736 ( .A(n9472), .B(n10481), .Z(n9435) );
  NAND U9737 ( .A(n9433), .B(n10482), .Z(n9434) );
  NAND U9738 ( .A(n9435), .B(n9434), .Z(n9457) );
  NANDN U9739 ( .A(n529), .B(a[224]), .Z(n9458) );
  XNOR U9740 ( .A(n9457), .B(n9458), .Z(n9460) );
  XOR U9741 ( .A(n9459), .B(n9460), .Z(n9454) );
  XOR U9742 ( .A(n9453), .B(n9454), .Z(n9475) );
  XOR U9743 ( .A(n9476), .B(n9475), .Z(n9477) );
  XNOR U9744 ( .A(n9478), .B(n9477), .Z(n9447) );
  NAND U9745 ( .A(n9437), .B(n9436), .Z(n9441) );
  NAND U9746 ( .A(n9439), .B(n9438), .Z(n9440) );
  NAND U9747 ( .A(n9441), .B(n9440), .Z(n9448) );
  XNOR U9748 ( .A(n9447), .B(n9448), .Z(n9449) );
  XNOR U9749 ( .A(n9450), .B(n9449), .Z(n9481) );
  XNOR U9750 ( .A(n9481), .B(sreg[480]), .Z(n9483) );
  NAND U9751 ( .A(n9442), .B(sreg[479]), .Z(n9446) );
  OR U9752 ( .A(n9444), .B(n9443), .Z(n9445) );
  AND U9753 ( .A(n9446), .B(n9445), .Z(n9482) );
  XOR U9754 ( .A(n9483), .B(n9482), .Z(c[480]) );
  NANDN U9755 ( .A(n9452), .B(n9451), .Z(n9456) );
  NAND U9756 ( .A(n9454), .B(n9453), .Z(n9455) );
  NAND U9757 ( .A(n9456), .B(n9455), .Z(n9517) );
  NANDN U9758 ( .A(n9458), .B(n9457), .Z(n9462) );
  NAND U9759 ( .A(n9460), .B(n9459), .Z(n9461) );
  NAND U9760 ( .A(n9462), .B(n9461), .Z(n9515) );
  XNOR U9761 ( .A(b[7]), .B(a[227]), .Z(n9502) );
  NANDN U9762 ( .A(n9502), .B(n10545), .Z(n9465) );
  NANDN U9763 ( .A(n9463), .B(n10546), .Z(n9464) );
  NAND U9764 ( .A(n9465), .B(n9464), .Z(n9490) );
  XNOR U9765 ( .A(b[3]), .B(a[231]), .Z(n9505) );
  NANDN U9766 ( .A(n9505), .B(n10398), .Z(n9468) );
  NANDN U9767 ( .A(n9466), .B(n10399), .Z(n9467) );
  AND U9768 ( .A(n9468), .B(n9467), .Z(n9491) );
  XNOR U9769 ( .A(n9490), .B(n9491), .Z(n9492) );
  NANDN U9770 ( .A(n527), .B(a[233]), .Z(n9469) );
  XOR U9771 ( .A(n10434), .B(n9469), .Z(n9471) );
  NANDN U9772 ( .A(b[0]), .B(a[232]), .Z(n9470) );
  AND U9773 ( .A(n9471), .B(n9470), .Z(n9498) );
  XOR U9774 ( .A(b[5]), .B(a[229]), .Z(n9511) );
  NAND U9775 ( .A(n9511), .B(n10481), .Z(n9474) );
  NAND U9776 ( .A(n9472), .B(n10482), .Z(n9473) );
  NAND U9777 ( .A(n9474), .B(n9473), .Z(n9496) );
  NANDN U9778 ( .A(n529), .B(a[225]), .Z(n9497) );
  XNOR U9779 ( .A(n9496), .B(n9497), .Z(n9499) );
  XOR U9780 ( .A(n9498), .B(n9499), .Z(n9493) );
  XOR U9781 ( .A(n9492), .B(n9493), .Z(n9514) );
  XOR U9782 ( .A(n9515), .B(n9514), .Z(n9516) );
  XNOR U9783 ( .A(n9517), .B(n9516), .Z(n9486) );
  NAND U9784 ( .A(n9476), .B(n9475), .Z(n9480) );
  NAND U9785 ( .A(n9478), .B(n9477), .Z(n9479) );
  NAND U9786 ( .A(n9480), .B(n9479), .Z(n9487) );
  XNOR U9787 ( .A(n9486), .B(n9487), .Z(n9488) );
  XNOR U9788 ( .A(n9489), .B(n9488), .Z(n9520) );
  XNOR U9789 ( .A(n9520), .B(sreg[481]), .Z(n9522) );
  NAND U9790 ( .A(n9481), .B(sreg[480]), .Z(n9485) );
  OR U9791 ( .A(n9483), .B(n9482), .Z(n9484) );
  AND U9792 ( .A(n9485), .B(n9484), .Z(n9521) );
  XOR U9793 ( .A(n9522), .B(n9521), .Z(c[481]) );
  NANDN U9794 ( .A(n9491), .B(n9490), .Z(n9495) );
  NAND U9795 ( .A(n9493), .B(n9492), .Z(n9494) );
  NAND U9796 ( .A(n9495), .B(n9494), .Z(n9556) );
  NANDN U9797 ( .A(n9497), .B(n9496), .Z(n9501) );
  NAND U9798 ( .A(n9499), .B(n9498), .Z(n9500) );
  NAND U9799 ( .A(n9501), .B(n9500), .Z(n9554) );
  XNOR U9800 ( .A(b[7]), .B(a[228]), .Z(n9541) );
  NANDN U9801 ( .A(n9541), .B(n10545), .Z(n9504) );
  NANDN U9802 ( .A(n9502), .B(n10546), .Z(n9503) );
  NAND U9803 ( .A(n9504), .B(n9503), .Z(n9529) );
  XNOR U9804 ( .A(b[3]), .B(a[232]), .Z(n9544) );
  NANDN U9805 ( .A(n9544), .B(n10398), .Z(n9507) );
  NANDN U9806 ( .A(n9505), .B(n10399), .Z(n9506) );
  AND U9807 ( .A(n9507), .B(n9506), .Z(n9530) );
  XNOR U9808 ( .A(n9529), .B(n9530), .Z(n9531) );
  NANDN U9809 ( .A(n527), .B(a[234]), .Z(n9508) );
  XOR U9810 ( .A(n10434), .B(n9508), .Z(n9510) );
  NANDN U9811 ( .A(b[0]), .B(a[233]), .Z(n9509) );
  AND U9812 ( .A(n9510), .B(n9509), .Z(n9537) );
  XOR U9813 ( .A(b[5]), .B(a[230]), .Z(n9550) );
  NAND U9814 ( .A(n9550), .B(n10481), .Z(n9513) );
  NAND U9815 ( .A(n9511), .B(n10482), .Z(n9512) );
  NAND U9816 ( .A(n9513), .B(n9512), .Z(n9535) );
  NANDN U9817 ( .A(n529), .B(a[226]), .Z(n9536) );
  XNOR U9818 ( .A(n9535), .B(n9536), .Z(n9538) );
  XOR U9819 ( .A(n9537), .B(n9538), .Z(n9532) );
  XOR U9820 ( .A(n9531), .B(n9532), .Z(n9553) );
  XOR U9821 ( .A(n9554), .B(n9553), .Z(n9555) );
  XNOR U9822 ( .A(n9556), .B(n9555), .Z(n9525) );
  NAND U9823 ( .A(n9515), .B(n9514), .Z(n9519) );
  NAND U9824 ( .A(n9517), .B(n9516), .Z(n9518) );
  NAND U9825 ( .A(n9519), .B(n9518), .Z(n9526) );
  XNOR U9826 ( .A(n9525), .B(n9526), .Z(n9527) );
  XNOR U9827 ( .A(n9528), .B(n9527), .Z(n9559) );
  XNOR U9828 ( .A(n9559), .B(sreg[482]), .Z(n9561) );
  NAND U9829 ( .A(n9520), .B(sreg[481]), .Z(n9524) );
  OR U9830 ( .A(n9522), .B(n9521), .Z(n9523) );
  AND U9831 ( .A(n9524), .B(n9523), .Z(n9560) );
  XOR U9832 ( .A(n9561), .B(n9560), .Z(c[482]) );
  NANDN U9833 ( .A(n9530), .B(n9529), .Z(n9534) );
  NAND U9834 ( .A(n9532), .B(n9531), .Z(n9533) );
  NAND U9835 ( .A(n9534), .B(n9533), .Z(n9595) );
  NANDN U9836 ( .A(n9536), .B(n9535), .Z(n9540) );
  NAND U9837 ( .A(n9538), .B(n9537), .Z(n9539) );
  NAND U9838 ( .A(n9540), .B(n9539), .Z(n9593) );
  XNOR U9839 ( .A(b[7]), .B(a[229]), .Z(n9586) );
  NANDN U9840 ( .A(n9586), .B(n10545), .Z(n9543) );
  NANDN U9841 ( .A(n9541), .B(n10546), .Z(n9542) );
  NAND U9842 ( .A(n9543), .B(n9542), .Z(n9568) );
  XNOR U9843 ( .A(b[3]), .B(a[233]), .Z(n9589) );
  NANDN U9844 ( .A(n9589), .B(n10398), .Z(n9546) );
  NANDN U9845 ( .A(n9544), .B(n10399), .Z(n9545) );
  AND U9846 ( .A(n9546), .B(n9545), .Z(n9569) );
  XNOR U9847 ( .A(n9568), .B(n9569), .Z(n9570) );
  NANDN U9848 ( .A(n527), .B(a[235]), .Z(n9547) );
  XOR U9849 ( .A(n10434), .B(n9547), .Z(n9549) );
  NANDN U9850 ( .A(b[0]), .B(a[234]), .Z(n9548) );
  AND U9851 ( .A(n9549), .B(n9548), .Z(n9576) );
  XOR U9852 ( .A(b[5]), .B(a[231]), .Z(n9583) );
  NAND U9853 ( .A(n9583), .B(n10481), .Z(n9552) );
  NAND U9854 ( .A(n9550), .B(n10482), .Z(n9551) );
  NAND U9855 ( .A(n9552), .B(n9551), .Z(n9574) );
  NANDN U9856 ( .A(n529), .B(a[227]), .Z(n9575) );
  XNOR U9857 ( .A(n9574), .B(n9575), .Z(n9577) );
  XOR U9858 ( .A(n9576), .B(n9577), .Z(n9571) );
  XOR U9859 ( .A(n9570), .B(n9571), .Z(n9592) );
  XOR U9860 ( .A(n9593), .B(n9592), .Z(n9594) );
  XNOR U9861 ( .A(n9595), .B(n9594), .Z(n9564) );
  NAND U9862 ( .A(n9554), .B(n9553), .Z(n9558) );
  NAND U9863 ( .A(n9556), .B(n9555), .Z(n9557) );
  NAND U9864 ( .A(n9558), .B(n9557), .Z(n9565) );
  XNOR U9865 ( .A(n9564), .B(n9565), .Z(n9566) );
  XNOR U9866 ( .A(n9567), .B(n9566), .Z(n9598) );
  XNOR U9867 ( .A(n9598), .B(sreg[483]), .Z(n9600) );
  NAND U9868 ( .A(n9559), .B(sreg[482]), .Z(n9563) );
  OR U9869 ( .A(n9561), .B(n9560), .Z(n9562) );
  AND U9870 ( .A(n9563), .B(n9562), .Z(n9599) );
  XOR U9871 ( .A(n9600), .B(n9599), .Z(c[483]) );
  NANDN U9872 ( .A(n9569), .B(n9568), .Z(n9573) );
  NAND U9873 ( .A(n9571), .B(n9570), .Z(n9572) );
  NAND U9874 ( .A(n9573), .B(n9572), .Z(n9634) );
  NANDN U9875 ( .A(n9575), .B(n9574), .Z(n9579) );
  NAND U9876 ( .A(n9577), .B(n9576), .Z(n9578) );
  NAND U9877 ( .A(n9579), .B(n9578), .Z(n9632) );
  NANDN U9878 ( .A(n527), .B(a[236]), .Z(n9580) );
  XOR U9879 ( .A(n10434), .B(n9580), .Z(n9582) );
  NANDN U9880 ( .A(b[0]), .B(a[235]), .Z(n9581) );
  AND U9881 ( .A(n9582), .B(n9581), .Z(n9615) );
  XOR U9882 ( .A(b[5]), .B(a[232]), .Z(n9622) );
  NAND U9883 ( .A(n9622), .B(n10481), .Z(n9585) );
  NAND U9884 ( .A(n9583), .B(n10482), .Z(n9584) );
  NAND U9885 ( .A(n9585), .B(n9584), .Z(n9613) );
  NANDN U9886 ( .A(n529), .B(a[228]), .Z(n9614) );
  XNOR U9887 ( .A(n9613), .B(n9614), .Z(n9616) );
  XOR U9888 ( .A(n9615), .B(n9616), .Z(n9609) );
  XNOR U9889 ( .A(b[7]), .B(a[230]), .Z(n9625) );
  NANDN U9890 ( .A(n9625), .B(n10545), .Z(n9588) );
  NANDN U9891 ( .A(n9586), .B(n10546), .Z(n9587) );
  NAND U9892 ( .A(n9588), .B(n9587), .Z(n9607) );
  XNOR U9893 ( .A(b[3]), .B(a[234]), .Z(n9628) );
  NANDN U9894 ( .A(n9628), .B(n10398), .Z(n9591) );
  NANDN U9895 ( .A(n9589), .B(n10399), .Z(n9590) );
  AND U9896 ( .A(n9591), .B(n9590), .Z(n9608) );
  XNOR U9897 ( .A(n9607), .B(n9608), .Z(n9610) );
  XOR U9898 ( .A(n9609), .B(n9610), .Z(n9631) );
  XOR U9899 ( .A(n9632), .B(n9631), .Z(n9633) );
  XNOR U9900 ( .A(n9634), .B(n9633), .Z(n9603) );
  NAND U9901 ( .A(n9593), .B(n9592), .Z(n9597) );
  NAND U9902 ( .A(n9595), .B(n9594), .Z(n9596) );
  NAND U9903 ( .A(n9597), .B(n9596), .Z(n9604) );
  XNOR U9904 ( .A(n9603), .B(n9604), .Z(n9605) );
  XNOR U9905 ( .A(n9606), .B(n9605), .Z(n9637) );
  XNOR U9906 ( .A(n9637), .B(sreg[484]), .Z(n9639) );
  NAND U9907 ( .A(n9598), .B(sreg[483]), .Z(n9602) );
  OR U9908 ( .A(n9600), .B(n9599), .Z(n9601) );
  AND U9909 ( .A(n9602), .B(n9601), .Z(n9638) );
  XOR U9910 ( .A(n9639), .B(n9638), .Z(c[484]) );
  NANDN U9911 ( .A(n9608), .B(n9607), .Z(n9612) );
  NAND U9912 ( .A(n9610), .B(n9609), .Z(n9611) );
  NAND U9913 ( .A(n9612), .B(n9611), .Z(n9673) );
  NANDN U9914 ( .A(n9614), .B(n9613), .Z(n9618) );
  NAND U9915 ( .A(n9616), .B(n9615), .Z(n9617) );
  NAND U9916 ( .A(n9618), .B(n9617), .Z(n9671) );
  NANDN U9917 ( .A(n527), .B(a[237]), .Z(n9619) );
  XOR U9918 ( .A(n10434), .B(n9619), .Z(n9621) );
  NANDN U9919 ( .A(b[0]), .B(a[236]), .Z(n9620) );
  AND U9920 ( .A(n9621), .B(n9620), .Z(n9654) );
  XOR U9921 ( .A(b[5]), .B(a[233]), .Z(n9667) );
  NAND U9922 ( .A(n9667), .B(n10481), .Z(n9624) );
  NAND U9923 ( .A(n9622), .B(n10482), .Z(n9623) );
  NAND U9924 ( .A(n9624), .B(n9623), .Z(n9652) );
  NANDN U9925 ( .A(n529), .B(a[229]), .Z(n9653) );
  XNOR U9926 ( .A(n9652), .B(n9653), .Z(n9655) );
  XOR U9927 ( .A(n9654), .B(n9655), .Z(n9648) );
  XNOR U9928 ( .A(b[7]), .B(a[231]), .Z(n9658) );
  NANDN U9929 ( .A(n9658), .B(n10545), .Z(n9627) );
  NANDN U9930 ( .A(n9625), .B(n10546), .Z(n9626) );
  NAND U9931 ( .A(n9627), .B(n9626), .Z(n9646) );
  XNOR U9932 ( .A(b[3]), .B(a[235]), .Z(n9661) );
  NANDN U9933 ( .A(n9661), .B(n10398), .Z(n9630) );
  NANDN U9934 ( .A(n9628), .B(n10399), .Z(n9629) );
  AND U9935 ( .A(n9630), .B(n9629), .Z(n9647) );
  XNOR U9936 ( .A(n9646), .B(n9647), .Z(n9649) );
  XOR U9937 ( .A(n9648), .B(n9649), .Z(n9670) );
  XOR U9938 ( .A(n9671), .B(n9670), .Z(n9672) );
  XNOR U9939 ( .A(n9673), .B(n9672), .Z(n9642) );
  NAND U9940 ( .A(n9632), .B(n9631), .Z(n9636) );
  NAND U9941 ( .A(n9634), .B(n9633), .Z(n9635) );
  NAND U9942 ( .A(n9636), .B(n9635), .Z(n9643) );
  XNOR U9943 ( .A(n9642), .B(n9643), .Z(n9644) );
  XNOR U9944 ( .A(n9645), .B(n9644), .Z(n9676) );
  XNOR U9945 ( .A(n9676), .B(sreg[485]), .Z(n9678) );
  NAND U9946 ( .A(n9637), .B(sreg[484]), .Z(n9641) );
  OR U9947 ( .A(n9639), .B(n9638), .Z(n9640) );
  AND U9948 ( .A(n9641), .B(n9640), .Z(n9677) );
  XOR U9949 ( .A(n9678), .B(n9677), .Z(c[485]) );
  NANDN U9950 ( .A(n9647), .B(n9646), .Z(n9651) );
  NAND U9951 ( .A(n9649), .B(n9648), .Z(n9650) );
  NAND U9952 ( .A(n9651), .B(n9650), .Z(n9712) );
  NANDN U9953 ( .A(n9653), .B(n9652), .Z(n9657) );
  NAND U9954 ( .A(n9655), .B(n9654), .Z(n9656) );
  NAND U9955 ( .A(n9657), .B(n9656), .Z(n9710) );
  XNOR U9956 ( .A(b[7]), .B(a[232]), .Z(n9697) );
  NANDN U9957 ( .A(n9697), .B(n10545), .Z(n9660) );
  NANDN U9958 ( .A(n9658), .B(n10546), .Z(n9659) );
  NAND U9959 ( .A(n9660), .B(n9659), .Z(n9685) );
  XNOR U9960 ( .A(b[3]), .B(a[236]), .Z(n9700) );
  NANDN U9961 ( .A(n9700), .B(n10398), .Z(n9663) );
  NANDN U9962 ( .A(n9661), .B(n10399), .Z(n9662) );
  AND U9963 ( .A(n9663), .B(n9662), .Z(n9686) );
  XNOR U9964 ( .A(n9685), .B(n9686), .Z(n9687) );
  NANDN U9965 ( .A(n527), .B(a[238]), .Z(n9664) );
  XOR U9966 ( .A(n10434), .B(n9664), .Z(n9666) );
  NANDN U9967 ( .A(b[0]), .B(a[237]), .Z(n9665) );
  AND U9968 ( .A(n9666), .B(n9665), .Z(n9693) );
  XOR U9969 ( .A(b[5]), .B(a[234]), .Z(n9706) );
  NAND U9970 ( .A(n9706), .B(n10481), .Z(n9669) );
  NAND U9971 ( .A(n9667), .B(n10482), .Z(n9668) );
  NAND U9972 ( .A(n9669), .B(n9668), .Z(n9691) );
  NANDN U9973 ( .A(n529), .B(a[230]), .Z(n9692) );
  XNOR U9974 ( .A(n9691), .B(n9692), .Z(n9694) );
  XOR U9975 ( .A(n9693), .B(n9694), .Z(n9688) );
  XOR U9976 ( .A(n9687), .B(n9688), .Z(n9709) );
  XOR U9977 ( .A(n9710), .B(n9709), .Z(n9711) );
  XNOR U9978 ( .A(n9712), .B(n9711), .Z(n9681) );
  NAND U9979 ( .A(n9671), .B(n9670), .Z(n9675) );
  NAND U9980 ( .A(n9673), .B(n9672), .Z(n9674) );
  NAND U9981 ( .A(n9675), .B(n9674), .Z(n9682) );
  XNOR U9982 ( .A(n9681), .B(n9682), .Z(n9683) );
  XNOR U9983 ( .A(n9684), .B(n9683), .Z(n9715) );
  XNOR U9984 ( .A(n9715), .B(sreg[486]), .Z(n9717) );
  NAND U9985 ( .A(n9676), .B(sreg[485]), .Z(n9680) );
  OR U9986 ( .A(n9678), .B(n9677), .Z(n9679) );
  AND U9987 ( .A(n9680), .B(n9679), .Z(n9716) );
  XOR U9988 ( .A(n9717), .B(n9716), .Z(c[486]) );
  NANDN U9989 ( .A(n9686), .B(n9685), .Z(n9690) );
  NAND U9990 ( .A(n9688), .B(n9687), .Z(n9689) );
  NAND U9991 ( .A(n9690), .B(n9689), .Z(n9751) );
  NANDN U9992 ( .A(n9692), .B(n9691), .Z(n9696) );
  NAND U9993 ( .A(n9694), .B(n9693), .Z(n9695) );
  NAND U9994 ( .A(n9696), .B(n9695), .Z(n9749) );
  XNOR U9995 ( .A(b[7]), .B(a[233]), .Z(n9736) );
  NANDN U9996 ( .A(n9736), .B(n10545), .Z(n9699) );
  NANDN U9997 ( .A(n9697), .B(n10546), .Z(n9698) );
  NAND U9998 ( .A(n9699), .B(n9698), .Z(n9724) );
  XNOR U9999 ( .A(b[3]), .B(a[237]), .Z(n9739) );
  NANDN U10000 ( .A(n9739), .B(n10398), .Z(n9702) );
  NANDN U10001 ( .A(n9700), .B(n10399), .Z(n9701) );
  AND U10002 ( .A(n9702), .B(n9701), .Z(n9725) );
  XNOR U10003 ( .A(n9724), .B(n9725), .Z(n9726) );
  NANDN U10004 ( .A(n527), .B(a[239]), .Z(n9703) );
  XOR U10005 ( .A(n10434), .B(n9703), .Z(n9705) );
  NANDN U10006 ( .A(b[0]), .B(a[238]), .Z(n9704) );
  AND U10007 ( .A(n9705), .B(n9704), .Z(n9732) );
  XOR U10008 ( .A(b[5]), .B(a[235]), .Z(n9745) );
  NAND U10009 ( .A(n9745), .B(n10481), .Z(n9708) );
  NAND U10010 ( .A(n9706), .B(n10482), .Z(n9707) );
  NAND U10011 ( .A(n9708), .B(n9707), .Z(n9730) );
  NANDN U10012 ( .A(n529), .B(a[231]), .Z(n9731) );
  XNOR U10013 ( .A(n9730), .B(n9731), .Z(n9733) );
  XOR U10014 ( .A(n9732), .B(n9733), .Z(n9727) );
  XOR U10015 ( .A(n9726), .B(n9727), .Z(n9748) );
  XOR U10016 ( .A(n9749), .B(n9748), .Z(n9750) );
  XNOR U10017 ( .A(n9751), .B(n9750), .Z(n9720) );
  NAND U10018 ( .A(n9710), .B(n9709), .Z(n9714) );
  NAND U10019 ( .A(n9712), .B(n9711), .Z(n9713) );
  NAND U10020 ( .A(n9714), .B(n9713), .Z(n9721) );
  XNOR U10021 ( .A(n9720), .B(n9721), .Z(n9722) );
  XNOR U10022 ( .A(n9723), .B(n9722), .Z(n9754) );
  XNOR U10023 ( .A(n9754), .B(sreg[487]), .Z(n9756) );
  NAND U10024 ( .A(n9715), .B(sreg[486]), .Z(n9719) );
  OR U10025 ( .A(n9717), .B(n9716), .Z(n9718) );
  AND U10026 ( .A(n9719), .B(n9718), .Z(n9755) );
  XOR U10027 ( .A(n9756), .B(n9755), .Z(c[487]) );
  NANDN U10028 ( .A(n9725), .B(n9724), .Z(n9729) );
  NAND U10029 ( .A(n9727), .B(n9726), .Z(n9728) );
  NAND U10030 ( .A(n9729), .B(n9728), .Z(n9790) );
  NANDN U10031 ( .A(n9731), .B(n9730), .Z(n9735) );
  NAND U10032 ( .A(n9733), .B(n9732), .Z(n9734) );
  NAND U10033 ( .A(n9735), .B(n9734), .Z(n9788) );
  XNOR U10034 ( .A(b[7]), .B(a[234]), .Z(n9775) );
  NANDN U10035 ( .A(n9775), .B(n10545), .Z(n9738) );
  NANDN U10036 ( .A(n9736), .B(n10546), .Z(n9737) );
  NAND U10037 ( .A(n9738), .B(n9737), .Z(n9763) );
  XNOR U10038 ( .A(b[3]), .B(a[238]), .Z(n9778) );
  NANDN U10039 ( .A(n9778), .B(n10398), .Z(n9741) );
  NANDN U10040 ( .A(n9739), .B(n10399), .Z(n9740) );
  AND U10041 ( .A(n9741), .B(n9740), .Z(n9764) );
  XNOR U10042 ( .A(n9763), .B(n9764), .Z(n9765) );
  NANDN U10043 ( .A(n527), .B(a[240]), .Z(n9742) );
  XOR U10044 ( .A(n10434), .B(n9742), .Z(n9744) );
  NANDN U10045 ( .A(b[0]), .B(a[239]), .Z(n9743) );
  AND U10046 ( .A(n9744), .B(n9743), .Z(n9771) );
  XOR U10047 ( .A(b[5]), .B(a[236]), .Z(n9784) );
  NAND U10048 ( .A(n9784), .B(n10481), .Z(n9747) );
  NAND U10049 ( .A(n9745), .B(n10482), .Z(n9746) );
  NAND U10050 ( .A(n9747), .B(n9746), .Z(n9769) );
  NANDN U10051 ( .A(n529), .B(a[232]), .Z(n9770) );
  XNOR U10052 ( .A(n9769), .B(n9770), .Z(n9772) );
  XOR U10053 ( .A(n9771), .B(n9772), .Z(n9766) );
  XOR U10054 ( .A(n9765), .B(n9766), .Z(n9787) );
  XOR U10055 ( .A(n9788), .B(n9787), .Z(n9789) );
  XNOR U10056 ( .A(n9790), .B(n9789), .Z(n9759) );
  NAND U10057 ( .A(n9749), .B(n9748), .Z(n9753) );
  NAND U10058 ( .A(n9751), .B(n9750), .Z(n9752) );
  NAND U10059 ( .A(n9753), .B(n9752), .Z(n9760) );
  XNOR U10060 ( .A(n9759), .B(n9760), .Z(n9761) );
  XNOR U10061 ( .A(n9762), .B(n9761), .Z(n9793) );
  XNOR U10062 ( .A(n9793), .B(sreg[488]), .Z(n9795) );
  NAND U10063 ( .A(n9754), .B(sreg[487]), .Z(n9758) );
  OR U10064 ( .A(n9756), .B(n9755), .Z(n9757) );
  AND U10065 ( .A(n9758), .B(n9757), .Z(n9794) );
  XOR U10066 ( .A(n9795), .B(n9794), .Z(c[488]) );
  NANDN U10067 ( .A(n9764), .B(n9763), .Z(n9768) );
  NAND U10068 ( .A(n9766), .B(n9765), .Z(n9767) );
  NAND U10069 ( .A(n9768), .B(n9767), .Z(n9829) );
  NANDN U10070 ( .A(n9770), .B(n9769), .Z(n9774) );
  NAND U10071 ( .A(n9772), .B(n9771), .Z(n9773) );
  NAND U10072 ( .A(n9774), .B(n9773), .Z(n9827) );
  XNOR U10073 ( .A(b[7]), .B(a[235]), .Z(n9814) );
  NANDN U10074 ( .A(n9814), .B(n10545), .Z(n9777) );
  NANDN U10075 ( .A(n9775), .B(n10546), .Z(n9776) );
  NAND U10076 ( .A(n9777), .B(n9776), .Z(n9802) );
  XNOR U10077 ( .A(b[3]), .B(a[239]), .Z(n9817) );
  NANDN U10078 ( .A(n9817), .B(n10398), .Z(n9780) );
  NANDN U10079 ( .A(n9778), .B(n10399), .Z(n9779) );
  AND U10080 ( .A(n9780), .B(n9779), .Z(n9803) );
  XNOR U10081 ( .A(n9802), .B(n9803), .Z(n9804) );
  NANDN U10082 ( .A(n527), .B(a[241]), .Z(n9781) );
  XOR U10083 ( .A(n10434), .B(n9781), .Z(n9783) );
  NANDN U10084 ( .A(b[0]), .B(a[240]), .Z(n9782) );
  AND U10085 ( .A(n9783), .B(n9782), .Z(n9810) );
  XOR U10086 ( .A(b[5]), .B(a[237]), .Z(n9823) );
  NAND U10087 ( .A(n9823), .B(n10481), .Z(n9786) );
  NAND U10088 ( .A(n9784), .B(n10482), .Z(n9785) );
  NAND U10089 ( .A(n9786), .B(n9785), .Z(n9808) );
  NANDN U10090 ( .A(n529), .B(a[233]), .Z(n9809) );
  XNOR U10091 ( .A(n9808), .B(n9809), .Z(n9811) );
  XOR U10092 ( .A(n9810), .B(n9811), .Z(n9805) );
  XOR U10093 ( .A(n9804), .B(n9805), .Z(n9826) );
  XOR U10094 ( .A(n9827), .B(n9826), .Z(n9828) );
  XNOR U10095 ( .A(n9829), .B(n9828), .Z(n9798) );
  NAND U10096 ( .A(n9788), .B(n9787), .Z(n9792) );
  NAND U10097 ( .A(n9790), .B(n9789), .Z(n9791) );
  NAND U10098 ( .A(n9792), .B(n9791), .Z(n9799) );
  XNOR U10099 ( .A(n9798), .B(n9799), .Z(n9800) );
  XNOR U10100 ( .A(n9801), .B(n9800), .Z(n9832) );
  XNOR U10101 ( .A(n9832), .B(sreg[489]), .Z(n9834) );
  NAND U10102 ( .A(n9793), .B(sreg[488]), .Z(n9797) );
  OR U10103 ( .A(n9795), .B(n9794), .Z(n9796) );
  AND U10104 ( .A(n9797), .B(n9796), .Z(n9833) );
  XOR U10105 ( .A(n9834), .B(n9833), .Z(c[489]) );
  NANDN U10106 ( .A(n9803), .B(n9802), .Z(n9807) );
  NAND U10107 ( .A(n9805), .B(n9804), .Z(n9806) );
  NAND U10108 ( .A(n9807), .B(n9806), .Z(n9868) );
  NANDN U10109 ( .A(n9809), .B(n9808), .Z(n9813) );
  NAND U10110 ( .A(n9811), .B(n9810), .Z(n9812) );
  NAND U10111 ( .A(n9813), .B(n9812), .Z(n9866) );
  XNOR U10112 ( .A(b[7]), .B(a[236]), .Z(n9853) );
  NANDN U10113 ( .A(n9853), .B(n10545), .Z(n9816) );
  NANDN U10114 ( .A(n9814), .B(n10546), .Z(n9815) );
  NAND U10115 ( .A(n9816), .B(n9815), .Z(n9841) );
  XNOR U10116 ( .A(b[3]), .B(a[240]), .Z(n9856) );
  NANDN U10117 ( .A(n9856), .B(n10398), .Z(n9819) );
  NANDN U10118 ( .A(n9817), .B(n10399), .Z(n9818) );
  AND U10119 ( .A(n9819), .B(n9818), .Z(n9842) );
  XNOR U10120 ( .A(n9841), .B(n9842), .Z(n9843) );
  NANDN U10121 ( .A(n527), .B(a[242]), .Z(n9820) );
  XOR U10122 ( .A(n10434), .B(n9820), .Z(n9822) );
  NANDN U10123 ( .A(b[0]), .B(a[241]), .Z(n9821) );
  AND U10124 ( .A(n9822), .B(n9821), .Z(n9849) );
  XOR U10125 ( .A(b[5]), .B(a[238]), .Z(n9862) );
  NAND U10126 ( .A(n9862), .B(n10481), .Z(n9825) );
  NAND U10127 ( .A(n9823), .B(n10482), .Z(n9824) );
  NAND U10128 ( .A(n9825), .B(n9824), .Z(n9847) );
  NANDN U10129 ( .A(n529), .B(a[234]), .Z(n9848) );
  XNOR U10130 ( .A(n9847), .B(n9848), .Z(n9850) );
  XOR U10131 ( .A(n9849), .B(n9850), .Z(n9844) );
  XOR U10132 ( .A(n9843), .B(n9844), .Z(n9865) );
  XOR U10133 ( .A(n9866), .B(n9865), .Z(n9867) );
  XNOR U10134 ( .A(n9868), .B(n9867), .Z(n9837) );
  NAND U10135 ( .A(n9827), .B(n9826), .Z(n9831) );
  NAND U10136 ( .A(n9829), .B(n9828), .Z(n9830) );
  NAND U10137 ( .A(n9831), .B(n9830), .Z(n9838) );
  XNOR U10138 ( .A(n9837), .B(n9838), .Z(n9839) );
  XNOR U10139 ( .A(n9840), .B(n9839), .Z(n9871) );
  XNOR U10140 ( .A(n9871), .B(sreg[490]), .Z(n9873) );
  NAND U10141 ( .A(n9832), .B(sreg[489]), .Z(n9836) );
  OR U10142 ( .A(n9834), .B(n9833), .Z(n9835) );
  AND U10143 ( .A(n9836), .B(n9835), .Z(n9872) );
  XOR U10144 ( .A(n9873), .B(n9872), .Z(c[490]) );
  NANDN U10145 ( .A(n9842), .B(n9841), .Z(n9846) );
  NAND U10146 ( .A(n9844), .B(n9843), .Z(n9845) );
  NAND U10147 ( .A(n9846), .B(n9845), .Z(n9907) );
  NANDN U10148 ( .A(n9848), .B(n9847), .Z(n9852) );
  NAND U10149 ( .A(n9850), .B(n9849), .Z(n9851) );
  NAND U10150 ( .A(n9852), .B(n9851), .Z(n9905) );
  XNOR U10151 ( .A(b[7]), .B(a[237]), .Z(n9892) );
  NANDN U10152 ( .A(n9892), .B(n10545), .Z(n9855) );
  NANDN U10153 ( .A(n9853), .B(n10546), .Z(n9854) );
  NAND U10154 ( .A(n9855), .B(n9854), .Z(n9880) );
  XNOR U10155 ( .A(b[3]), .B(a[241]), .Z(n9895) );
  NANDN U10156 ( .A(n9895), .B(n10398), .Z(n9858) );
  NANDN U10157 ( .A(n9856), .B(n10399), .Z(n9857) );
  AND U10158 ( .A(n9858), .B(n9857), .Z(n9881) );
  XNOR U10159 ( .A(n9880), .B(n9881), .Z(n9882) );
  NANDN U10160 ( .A(n527), .B(a[243]), .Z(n9859) );
  XOR U10161 ( .A(n10434), .B(n9859), .Z(n9861) );
  NANDN U10162 ( .A(b[0]), .B(a[242]), .Z(n9860) );
  AND U10163 ( .A(n9861), .B(n9860), .Z(n9888) );
  XOR U10164 ( .A(b[5]), .B(a[239]), .Z(n9901) );
  NAND U10165 ( .A(n9901), .B(n10481), .Z(n9864) );
  NAND U10166 ( .A(n9862), .B(n10482), .Z(n9863) );
  NAND U10167 ( .A(n9864), .B(n9863), .Z(n9886) );
  NANDN U10168 ( .A(n529), .B(a[235]), .Z(n9887) );
  XNOR U10169 ( .A(n9886), .B(n9887), .Z(n9889) );
  XOR U10170 ( .A(n9888), .B(n9889), .Z(n9883) );
  XOR U10171 ( .A(n9882), .B(n9883), .Z(n9904) );
  XOR U10172 ( .A(n9905), .B(n9904), .Z(n9906) );
  XNOR U10173 ( .A(n9907), .B(n9906), .Z(n9876) );
  NAND U10174 ( .A(n9866), .B(n9865), .Z(n9870) );
  NAND U10175 ( .A(n9868), .B(n9867), .Z(n9869) );
  NAND U10176 ( .A(n9870), .B(n9869), .Z(n9877) );
  XNOR U10177 ( .A(n9876), .B(n9877), .Z(n9878) );
  XNOR U10178 ( .A(n9879), .B(n9878), .Z(n9910) );
  XNOR U10179 ( .A(n9910), .B(sreg[491]), .Z(n9912) );
  NAND U10180 ( .A(n9871), .B(sreg[490]), .Z(n9875) );
  OR U10181 ( .A(n9873), .B(n9872), .Z(n9874) );
  AND U10182 ( .A(n9875), .B(n9874), .Z(n9911) );
  XOR U10183 ( .A(n9912), .B(n9911), .Z(c[491]) );
  NANDN U10184 ( .A(n9881), .B(n9880), .Z(n9885) );
  NAND U10185 ( .A(n9883), .B(n9882), .Z(n9884) );
  NAND U10186 ( .A(n9885), .B(n9884), .Z(n9946) );
  NANDN U10187 ( .A(n9887), .B(n9886), .Z(n9891) );
  NAND U10188 ( .A(n9889), .B(n9888), .Z(n9890) );
  NAND U10189 ( .A(n9891), .B(n9890), .Z(n9944) );
  XNOR U10190 ( .A(b[7]), .B(a[238]), .Z(n9931) );
  NANDN U10191 ( .A(n9931), .B(n10545), .Z(n9894) );
  NANDN U10192 ( .A(n9892), .B(n10546), .Z(n9893) );
  NAND U10193 ( .A(n9894), .B(n9893), .Z(n9919) );
  XNOR U10194 ( .A(b[3]), .B(a[242]), .Z(n9934) );
  NANDN U10195 ( .A(n9934), .B(n10398), .Z(n9897) );
  NANDN U10196 ( .A(n9895), .B(n10399), .Z(n9896) );
  AND U10197 ( .A(n9897), .B(n9896), .Z(n9920) );
  XNOR U10198 ( .A(n9919), .B(n9920), .Z(n9921) );
  NANDN U10199 ( .A(n527), .B(a[244]), .Z(n9898) );
  XOR U10200 ( .A(n10434), .B(n9898), .Z(n9900) );
  NANDN U10201 ( .A(b[0]), .B(a[243]), .Z(n9899) );
  AND U10202 ( .A(n9900), .B(n9899), .Z(n9927) );
  XOR U10203 ( .A(b[5]), .B(a[240]), .Z(n9940) );
  NAND U10204 ( .A(n9940), .B(n10481), .Z(n9903) );
  NAND U10205 ( .A(n9901), .B(n10482), .Z(n9902) );
  NAND U10206 ( .A(n9903), .B(n9902), .Z(n9925) );
  NANDN U10207 ( .A(n529), .B(a[236]), .Z(n9926) );
  XNOR U10208 ( .A(n9925), .B(n9926), .Z(n9928) );
  XOR U10209 ( .A(n9927), .B(n9928), .Z(n9922) );
  XOR U10210 ( .A(n9921), .B(n9922), .Z(n9943) );
  XOR U10211 ( .A(n9944), .B(n9943), .Z(n9945) );
  XNOR U10212 ( .A(n9946), .B(n9945), .Z(n9915) );
  NAND U10213 ( .A(n9905), .B(n9904), .Z(n9909) );
  NAND U10214 ( .A(n9907), .B(n9906), .Z(n9908) );
  NAND U10215 ( .A(n9909), .B(n9908), .Z(n9916) );
  XNOR U10216 ( .A(n9915), .B(n9916), .Z(n9917) );
  XNOR U10217 ( .A(n9918), .B(n9917), .Z(n9949) );
  XNOR U10218 ( .A(n9949), .B(sreg[492]), .Z(n9951) );
  NAND U10219 ( .A(n9910), .B(sreg[491]), .Z(n9914) );
  OR U10220 ( .A(n9912), .B(n9911), .Z(n9913) );
  AND U10221 ( .A(n9914), .B(n9913), .Z(n9950) );
  XOR U10222 ( .A(n9951), .B(n9950), .Z(c[492]) );
  NANDN U10223 ( .A(n9920), .B(n9919), .Z(n9924) );
  NAND U10224 ( .A(n9922), .B(n9921), .Z(n9923) );
  NAND U10225 ( .A(n9924), .B(n9923), .Z(n9985) );
  NANDN U10226 ( .A(n9926), .B(n9925), .Z(n9930) );
  NAND U10227 ( .A(n9928), .B(n9927), .Z(n9929) );
  NAND U10228 ( .A(n9930), .B(n9929), .Z(n9983) );
  XNOR U10229 ( .A(b[7]), .B(a[239]), .Z(n9970) );
  NANDN U10230 ( .A(n9970), .B(n10545), .Z(n9933) );
  NANDN U10231 ( .A(n9931), .B(n10546), .Z(n9932) );
  NAND U10232 ( .A(n9933), .B(n9932), .Z(n9958) );
  XNOR U10233 ( .A(b[3]), .B(a[243]), .Z(n9973) );
  NANDN U10234 ( .A(n9973), .B(n10398), .Z(n9936) );
  NANDN U10235 ( .A(n9934), .B(n10399), .Z(n9935) );
  AND U10236 ( .A(n9936), .B(n9935), .Z(n9959) );
  XNOR U10237 ( .A(n9958), .B(n9959), .Z(n9960) );
  NANDN U10238 ( .A(n527), .B(a[245]), .Z(n9937) );
  XOR U10239 ( .A(n10434), .B(n9937), .Z(n9939) );
  NANDN U10240 ( .A(b[0]), .B(a[244]), .Z(n9938) );
  AND U10241 ( .A(n9939), .B(n9938), .Z(n9966) );
  XOR U10242 ( .A(b[5]), .B(a[241]), .Z(n9979) );
  NAND U10243 ( .A(n9979), .B(n10481), .Z(n9942) );
  NAND U10244 ( .A(n9940), .B(n10482), .Z(n9941) );
  NAND U10245 ( .A(n9942), .B(n9941), .Z(n9964) );
  NANDN U10246 ( .A(n529), .B(a[237]), .Z(n9965) );
  XNOR U10247 ( .A(n9964), .B(n9965), .Z(n9967) );
  XOR U10248 ( .A(n9966), .B(n9967), .Z(n9961) );
  XOR U10249 ( .A(n9960), .B(n9961), .Z(n9982) );
  XOR U10250 ( .A(n9983), .B(n9982), .Z(n9984) );
  XNOR U10251 ( .A(n9985), .B(n9984), .Z(n9954) );
  NAND U10252 ( .A(n9944), .B(n9943), .Z(n9948) );
  NAND U10253 ( .A(n9946), .B(n9945), .Z(n9947) );
  NAND U10254 ( .A(n9948), .B(n9947), .Z(n9955) );
  XNOR U10255 ( .A(n9954), .B(n9955), .Z(n9956) );
  XNOR U10256 ( .A(n9957), .B(n9956), .Z(n9988) );
  XNOR U10257 ( .A(n9988), .B(sreg[493]), .Z(n9990) );
  NAND U10258 ( .A(n9949), .B(sreg[492]), .Z(n9953) );
  OR U10259 ( .A(n9951), .B(n9950), .Z(n9952) );
  AND U10260 ( .A(n9953), .B(n9952), .Z(n9989) );
  XOR U10261 ( .A(n9990), .B(n9989), .Z(c[493]) );
  NANDN U10262 ( .A(n9959), .B(n9958), .Z(n9963) );
  NAND U10263 ( .A(n9961), .B(n9960), .Z(n9962) );
  NAND U10264 ( .A(n9963), .B(n9962), .Z(n10024) );
  NANDN U10265 ( .A(n9965), .B(n9964), .Z(n9969) );
  NAND U10266 ( .A(n9967), .B(n9966), .Z(n9968) );
  NAND U10267 ( .A(n9969), .B(n9968), .Z(n10022) );
  XNOR U10268 ( .A(b[7]), .B(a[240]), .Z(n10009) );
  NANDN U10269 ( .A(n10009), .B(n10545), .Z(n9972) );
  NANDN U10270 ( .A(n9970), .B(n10546), .Z(n9971) );
  NAND U10271 ( .A(n9972), .B(n9971), .Z(n9997) );
  XNOR U10272 ( .A(b[3]), .B(a[244]), .Z(n10012) );
  NANDN U10273 ( .A(n10012), .B(n10398), .Z(n9975) );
  NANDN U10274 ( .A(n9973), .B(n10399), .Z(n9974) );
  AND U10275 ( .A(n9975), .B(n9974), .Z(n9998) );
  XNOR U10276 ( .A(n9997), .B(n9998), .Z(n9999) );
  NANDN U10277 ( .A(n527), .B(a[246]), .Z(n9976) );
  XOR U10278 ( .A(n10434), .B(n9976), .Z(n9978) );
  NANDN U10279 ( .A(b[0]), .B(a[245]), .Z(n9977) );
  AND U10280 ( .A(n9978), .B(n9977), .Z(n10005) );
  XOR U10281 ( .A(b[5]), .B(a[242]), .Z(n10018) );
  NAND U10282 ( .A(n10018), .B(n10481), .Z(n9981) );
  NAND U10283 ( .A(n9979), .B(n10482), .Z(n9980) );
  NAND U10284 ( .A(n9981), .B(n9980), .Z(n10003) );
  NANDN U10285 ( .A(n529), .B(a[238]), .Z(n10004) );
  XNOR U10286 ( .A(n10003), .B(n10004), .Z(n10006) );
  XOR U10287 ( .A(n10005), .B(n10006), .Z(n10000) );
  XOR U10288 ( .A(n9999), .B(n10000), .Z(n10021) );
  XOR U10289 ( .A(n10022), .B(n10021), .Z(n10023) );
  XNOR U10290 ( .A(n10024), .B(n10023), .Z(n9993) );
  NAND U10291 ( .A(n9983), .B(n9982), .Z(n9987) );
  NAND U10292 ( .A(n9985), .B(n9984), .Z(n9986) );
  NAND U10293 ( .A(n9987), .B(n9986), .Z(n9994) );
  XNOR U10294 ( .A(n9993), .B(n9994), .Z(n9995) );
  XNOR U10295 ( .A(n9996), .B(n9995), .Z(n10027) );
  XNOR U10296 ( .A(n10027), .B(sreg[494]), .Z(n10029) );
  NAND U10297 ( .A(n9988), .B(sreg[493]), .Z(n9992) );
  OR U10298 ( .A(n9990), .B(n9989), .Z(n9991) );
  AND U10299 ( .A(n9992), .B(n9991), .Z(n10028) );
  XOR U10300 ( .A(n10029), .B(n10028), .Z(c[494]) );
  NANDN U10301 ( .A(n9998), .B(n9997), .Z(n10002) );
  NAND U10302 ( .A(n10000), .B(n9999), .Z(n10001) );
  NAND U10303 ( .A(n10002), .B(n10001), .Z(n10063) );
  NANDN U10304 ( .A(n10004), .B(n10003), .Z(n10008) );
  NAND U10305 ( .A(n10006), .B(n10005), .Z(n10007) );
  NAND U10306 ( .A(n10008), .B(n10007), .Z(n10061) );
  XNOR U10307 ( .A(b[7]), .B(a[241]), .Z(n10048) );
  NANDN U10308 ( .A(n10048), .B(n10545), .Z(n10011) );
  NANDN U10309 ( .A(n10009), .B(n10546), .Z(n10010) );
  NAND U10310 ( .A(n10011), .B(n10010), .Z(n10036) );
  XNOR U10311 ( .A(b[3]), .B(a[245]), .Z(n10051) );
  NANDN U10312 ( .A(n10051), .B(n10398), .Z(n10014) );
  NANDN U10313 ( .A(n10012), .B(n10399), .Z(n10013) );
  AND U10314 ( .A(n10014), .B(n10013), .Z(n10037) );
  XNOR U10315 ( .A(n10036), .B(n10037), .Z(n10038) );
  NANDN U10316 ( .A(n527), .B(a[247]), .Z(n10015) );
  XOR U10317 ( .A(n10434), .B(n10015), .Z(n10017) );
  NANDN U10318 ( .A(b[0]), .B(a[246]), .Z(n10016) );
  AND U10319 ( .A(n10017), .B(n10016), .Z(n10044) );
  XOR U10320 ( .A(b[5]), .B(a[243]), .Z(n10057) );
  NAND U10321 ( .A(n10057), .B(n10481), .Z(n10020) );
  NAND U10322 ( .A(n10018), .B(n10482), .Z(n10019) );
  NAND U10323 ( .A(n10020), .B(n10019), .Z(n10042) );
  NANDN U10324 ( .A(n529), .B(a[239]), .Z(n10043) );
  XNOR U10325 ( .A(n10042), .B(n10043), .Z(n10045) );
  XOR U10326 ( .A(n10044), .B(n10045), .Z(n10039) );
  XOR U10327 ( .A(n10038), .B(n10039), .Z(n10060) );
  XOR U10328 ( .A(n10061), .B(n10060), .Z(n10062) );
  XNOR U10329 ( .A(n10063), .B(n10062), .Z(n10032) );
  NAND U10330 ( .A(n10022), .B(n10021), .Z(n10026) );
  NAND U10331 ( .A(n10024), .B(n10023), .Z(n10025) );
  NAND U10332 ( .A(n10026), .B(n10025), .Z(n10033) );
  XNOR U10333 ( .A(n10032), .B(n10033), .Z(n10034) );
  XNOR U10334 ( .A(n10035), .B(n10034), .Z(n10066) );
  XNOR U10335 ( .A(n10066), .B(sreg[495]), .Z(n10068) );
  NAND U10336 ( .A(n10027), .B(sreg[494]), .Z(n10031) );
  OR U10337 ( .A(n10029), .B(n10028), .Z(n10030) );
  AND U10338 ( .A(n10031), .B(n10030), .Z(n10067) );
  XOR U10339 ( .A(n10068), .B(n10067), .Z(c[495]) );
  NANDN U10340 ( .A(n10037), .B(n10036), .Z(n10041) );
  NAND U10341 ( .A(n10039), .B(n10038), .Z(n10040) );
  NAND U10342 ( .A(n10041), .B(n10040), .Z(n10102) );
  NANDN U10343 ( .A(n10043), .B(n10042), .Z(n10047) );
  NAND U10344 ( .A(n10045), .B(n10044), .Z(n10046) );
  NAND U10345 ( .A(n10047), .B(n10046), .Z(n10100) );
  XNOR U10346 ( .A(b[7]), .B(a[242]), .Z(n10087) );
  NANDN U10347 ( .A(n10087), .B(n10545), .Z(n10050) );
  NANDN U10348 ( .A(n10048), .B(n10546), .Z(n10049) );
  NAND U10349 ( .A(n10050), .B(n10049), .Z(n10075) );
  XNOR U10350 ( .A(b[3]), .B(a[246]), .Z(n10090) );
  NANDN U10351 ( .A(n10090), .B(n10398), .Z(n10053) );
  NANDN U10352 ( .A(n10051), .B(n10399), .Z(n10052) );
  AND U10353 ( .A(n10053), .B(n10052), .Z(n10076) );
  XNOR U10354 ( .A(n10075), .B(n10076), .Z(n10077) );
  NANDN U10355 ( .A(n527), .B(a[248]), .Z(n10054) );
  XOR U10356 ( .A(n10434), .B(n10054), .Z(n10056) );
  IV U10357 ( .A(a[247]), .Z(n10321) );
  NANDN U10358 ( .A(n10321), .B(n527), .Z(n10055) );
  AND U10359 ( .A(n10056), .B(n10055), .Z(n10083) );
  XOR U10360 ( .A(b[5]), .B(a[244]), .Z(n10096) );
  NAND U10361 ( .A(n10096), .B(n10481), .Z(n10059) );
  NAND U10362 ( .A(n10057), .B(n10482), .Z(n10058) );
  NAND U10363 ( .A(n10059), .B(n10058), .Z(n10081) );
  NANDN U10364 ( .A(n529), .B(a[240]), .Z(n10082) );
  XNOR U10365 ( .A(n10081), .B(n10082), .Z(n10084) );
  XOR U10366 ( .A(n10083), .B(n10084), .Z(n10078) );
  XOR U10367 ( .A(n10077), .B(n10078), .Z(n10099) );
  XOR U10368 ( .A(n10100), .B(n10099), .Z(n10101) );
  XNOR U10369 ( .A(n10102), .B(n10101), .Z(n10071) );
  NAND U10370 ( .A(n10061), .B(n10060), .Z(n10065) );
  NAND U10371 ( .A(n10063), .B(n10062), .Z(n10064) );
  NAND U10372 ( .A(n10065), .B(n10064), .Z(n10072) );
  XNOR U10373 ( .A(n10071), .B(n10072), .Z(n10073) );
  XNOR U10374 ( .A(n10074), .B(n10073), .Z(n10105) );
  XNOR U10375 ( .A(n10105), .B(sreg[496]), .Z(n10107) );
  NAND U10376 ( .A(n10066), .B(sreg[495]), .Z(n10070) );
  OR U10377 ( .A(n10068), .B(n10067), .Z(n10069) );
  AND U10378 ( .A(n10070), .B(n10069), .Z(n10106) );
  XOR U10379 ( .A(n10107), .B(n10106), .Z(c[496]) );
  NANDN U10380 ( .A(n10076), .B(n10075), .Z(n10080) );
  NAND U10381 ( .A(n10078), .B(n10077), .Z(n10079) );
  NAND U10382 ( .A(n10080), .B(n10079), .Z(n10141) );
  NANDN U10383 ( .A(n10082), .B(n10081), .Z(n10086) );
  NAND U10384 ( .A(n10084), .B(n10083), .Z(n10085) );
  NAND U10385 ( .A(n10086), .B(n10085), .Z(n10139) );
  XNOR U10386 ( .A(b[7]), .B(a[243]), .Z(n10126) );
  NANDN U10387 ( .A(n10126), .B(n10545), .Z(n10089) );
  NANDN U10388 ( .A(n10087), .B(n10546), .Z(n10088) );
  NAND U10389 ( .A(n10089), .B(n10088), .Z(n10114) );
  XOR U10390 ( .A(b[3]), .B(n10321), .Z(n10129) );
  NANDN U10391 ( .A(n10129), .B(n10398), .Z(n10092) );
  NANDN U10392 ( .A(n10090), .B(n10399), .Z(n10091) );
  AND U10393 ( .A(n10092), .B(n10091), .Z(n10115) );
  XNOR U10394 ( .A(n10114), .B(n10115), .Z(n10116) );
  NANDN U10395 ( .A(n527), .B(a[249]), .Z(n10093) );
  XOR U10396 ( .A(n10434), .B(n10093), .Z(n10095) );
  NANDN U10397 ( .A(b[0]), .B(a[248]), .Z(n10094) );
  AND U10398 ( .A(n10095), .B(n10094), .Z(n10122) );
  XOR U10399 ( .A(b[5]), .B(a[245]), .Z(n10135) );
  NAND U10400 ( .A(n10135), .B(n10481), .Z(n10098) );
  NAND U10401 ( .A(n10096), .B(n10482), .Z(n10097) );
  NAND U10402 ( .A(n10098), .B(n10097), .Z(n10120) );
  NANDN U10403 ( .A(n529), .B(a[241]), .Z(n10121) );
  XNOR U10404 ( .A(n10120), .B(n10121), .Z(n10123) );
  XOR U10405 ( .A(n10122), .B(n10123), .Z(n10117) );
  XOR U10406 ( .A(n10116), .B(n10117), .Z(n10138) );
  XOR U10407 ( .A(n10139), .B(n10138), .Z(n10140) );
  XNOR U10408 ( .A(n10141), .B(n10140), .Z(n10110) );
  NAND U10409 ( .A(n10100), .B(n10099), .Z(n10104) );
  NAND U10410 ( .A(n10102), .B(n10101), .Z(n10103) );
  NAND U10411 ( .A(n10104), .B(n10103), .Z(n10111) );
  XNOR U10412 ( .A(n10110), .B(n10111), .Z(n10112) );
  XNOR U10413 ( .A(n10113), .B(n10112), .Z(n10144) );
  XNOR U10414 ( .A(n10144), .B(sreg[497]), .Z(n10146) );
  NAND U10415 ( .A(n10105), .B(sreg[496]), .Z(n10109) );
  OR U10416 ( .A(n10107), .B(n10106), .Z(n10108) );
  AND U10417 ( .A(n10109), .B(n10108), .Z(n10145) );
  XOR U10418 ( .A(n10146), .B(n10145), .Z(c[497]) );
  NANDN U10419 ( .A(n10115), .B(n10114), .Z(n10119) );
  NAND U10420 ( .A(n10117), .B(n10116), .Z(n10118) );
  NAND U10421 ( .A(n10119), .B(n10118), .Z(n10180) );
  NANDN U10422 ( .A(n10121), .B(n10120), .Z(n10125) );
  NAND U10423 ( .A(n10123), .B(n10122), .Z(n10124) );
  NAND U10424 ( .A(n10125), .B(n10124), .Z(n10178) );
  XNOR U10425 ( .A(b[7]), .B(a[244]), .Z(n10165) );
  NANDN U10426 ( .A(n10165), .B(n10545), .Z(n10128) );
  NANDN U10427 ( .A(n10126), .B(n10546), .Z(n10127) );
  NAND U10428 ( .A(n10128), .B(n10127), .Z(n10153) );
  XNOR U10429 ( .A(b[3]), .B(a[248]), .Z(n10168) );
  NANDN U10430 ( .A(n10168), .B(n10398), .Z(n10131) );
  NANDN U10431 ( .A(n10129), .B(n10399), .Z(n10130) );
  AND U10432 ( .A(n10131), .B(n10130), .Z(n10154) );
  XNOR U10433 ( .A(n10153), .B(n10154), .Z(n10155) );
  NANDN U10434 ( .A(n527), .B(a[250]), .Z(n10132) );
  XOR U10435 ( .A(n10434), .B(n10132), .Z(n10134) );
  IV U10436 ( .A(a[249]), .Z(n10331) );
  NANDN U10437 ( .A(n10331), .B(n527), .Z(n10133) );
  AND U10438 ( .A(n10134), .B(n10133), .Z(n10161) );
  XOR U10439 ( .A(b[5]), .B(a[246]), .Z(n10174) );
  NAND U10440 ( .A(n10174), .B(n10481), .Z(n10137) );
  NAND U10441 ( .A(n10135), .B(n10482), .Z(n10136) );
  NAND U10442 ( .A(n10137), .B(n10136), .Z(n10159) );
  NANDN U10443 ( .A(n529), .B(a[242]), .Z(n10160) );
  XNOR U10444 ( .A(n10159), .B(n10160), .Z(n10162) );
  XOR U10445 ( .A(n10161), .B(n10162), .Z(n10156) );
  XOR U10446 ( .A(n10155), .B(n10156), .Z(n10177) );
  XOR U10447 ( .A(n10178), .B(n10177), .Z(n10179) );
  XNOR U10448 ( .A(n10180), .B(n10179), .Z(n10149) );
  NAND U10449 ( .A(n10139), .B(n10138), .Z(n10143) );
  NAND U10450 ( .A(n10141), .B(n10140), .Z(n10142) );
  NAND U10451 ( .A(n10143), .B(n10142), .Z(n10150) );
  XNOR U10452 ( .A(n10149), .B(n10150), .Z(n10151) );
  XNOR U10453 ( .A(n10152), .B(n10151), .Z(n10183) );
  XNOR U10454 ( .A(n10183), .B(sreg[498]), .Z(n10185) );
  NAND U10455 ( .A(n10144), .B(sreg[497]), .Z(n10148) );
  OR U10456 ( .A(n10146), .B(n10145), .Z(n10147) );
  AND U10457 ( .A(n10148), .B(n10147), .Z(n10184) );
  XOR U10458 ( .A(n10185), .B(n10184), .Z(c[498]) );
  NANDN U10459 ( .A(n10154), .B(n10153), .Z(n10158) );
  NAND U10460 ( .A(n10156), .B(n10155), .Z(n10157) );
  NAND U10461 ( .A(n10158), .B(n10157), .Z(n10219) );
  NANDN U10462 ( .A(n10160), .B(n10159), .Z(n10164) );
  NAND U10463 ( .A(n10162), .B(n10161), .Z(n10163) );
  NAND U10464 ( .A(n10164), .B(n10163), .Z(n10217) );
  XNOR U10465 ( .A(b[7]), .B(a[245]), .Z(n10204) );
  NANDN U10466 ( .A(n10204), .B(n10545), .Z(n10167) );
  NANDN U10467 ( .A(n10165), .B(n10546), .Z(n10166) );
  NAND U10468 ( .A(n10167), .B(n10166), .Z(n10192) );
  XOR U10469 ( .A(b[3]), .B(n10331), .Z(n10207) );
  NANDN U10470 ( .A(n10207), .B(n10398), .Z(n10170) );
  NANDN U10471 ( .A(n10168), .B(n10399), .Z(n10169) );
  AND U10472 ( .A(n10170), .B(n10169), .Z(n10193) );
  XNOR U10473 ( .A(n10192), .B(n10193), .Z(n10194) );
  NANDN U10474 ( .A(n527), .B(a[251]), .Z(n10171) );
  XOR U10475 ( .A(n10434), .B(n10171), .Z(n10173) );
  NANDN U10476 ( .A(b[0]), .B(a[250]), .Z(n10172) );
  AND U10477 ( .A(n10173), .B(n10172), .Z(n10200) );
  XNOR U10478 ( .A(b[5]), .B(a[247]), .Z(n10213) );
  NANDN U10479 ( .A(n10213), .B(n10481), .Z(n10176) );
  NAND U10480 ( .A(n10174), .B(n10482), .Z(n10175) );
  NAND U10481 ( .A(n10176), .B(n10175), .Z(n10198) );
  NANDN U10482 ( .A(n529), .B(a[243]), .Z(n10199) );
  XNOR U10483 ( .A(n10198), .B(n10199), .Z(n10201) );
  XOR U10484 ( .A(n10200), .B(n10201), .Z(n10195) );
  XOR U10485 ( .A(n10194), .B(n10195), .Z(n10216) );
  XOR U10486 ( .A(n10217), .B(n10216), .Z(n10218) );
  XNOR U10487 ( .A(n10219), .B(n10218), .Z(n10188) );
  NAND U10488 ( .A(n10178), .B(n10177), .Z(n10182) );
  NAND U10489 ( .A(n10180), .B(n10179), .Z(n10181) );
  NAND U10490 ( .A(n10182), .B(n10181), .Z(n10189) );
  XNOR U10491 ( .A(n10188), .B(n10189), .Z(n10190) );
  XNOR U10492 ( .A(n10191), .B(n10190), .Z(n10222) );
  XNOR U10493 ( .A(n10222), .B(sreg[499]), .Z(n10224) );
  NAND U10494 ( .A(n10183), .B(sreg[498]), .Z(n10187) );
  OR U10495 ( .A(n10185), .B(n10184), .Z(n10186) );
  AND U10496 ( .A(n10187), .B(n10186), .Z(n10223) );
  XOR U10497 ( .A(n10224), .B(n10223), .Z(c[499]) );
  NANDN U10498 ( .A(n10193), .B(n10192), .Z(n10197) );
  NAND U10499 ( .A(n10195), .B(n10194), .Z(n10196) );
  NAND U10500 ( .A(n10197), .B(n10196), .Z(n10258) );
  NANDN U10501 ( .A(n10199), .B(n10198), .Z(n10203) );
  NAND U10502 ( .A(n10201), .B(n10200), .Z(n10202) );
  NAND U10503 ( .A(n10203), .B(n10202), .Z(n10256) );
  XNOR U10504 ( .A(b[7]), .B(a[246]), .Z(n10243) );
  NANDN U10505 ( .A(n10243), .B(n10545), .Z(n10206) );
  NANDN U10506 ( .A(n10204), .B(n10546), .Z(n10205) );
  NAND U10507 ( .A(n10206), .B(n10205), .Z(n10231) );
  XNOR U10508 ( .A(b[3]), .B(a[250]), .Z(n10246) );
  NANDN U10509 ( .A(n10246), .B(n10398), .Z(n10209) );
  NANDN U10510 ( .A(n10207), .B(n10399), .Z(n10208) );
  AND U10511 ( .A(n10209), .B(n10208), .Z(n10232) );
  XNOR U10512 ( .A(n10231), .B(n10232), .Z(n10233) );
  NANDN U10513 ( .A(n527), .B(a[252]), .Z(n10210) );
  XOR U10514 ( .A(n10434), .B(n10210), .Z(n10212) );
  NANDN U10515 ( .A(b[0]), .B(a[251]), .Z(n10211) );
  AND U10516 ( .A(n10212), .B(n10211), .Z(n10239) );
  XOR U10517 ( .A(b[5]), .B(a[248]), .Z(n10252) );
  NAND U10518 ( .A(n10252), .B(n10481), .Z(n10215) );
  NANDN U10519 ( .A(n10213), .B(n10482), .Z(n10214) );
  NAND U10520 ( .A(n10215), .B(n10214), .Z(n10237) );
  NANDN U10521 ( .A(n529), .B(a[244]), .Z(n10238) );
  XNOR U10522 ( .A(n10237), .B(n10238), .Z(n10240) );
  XOR U10523 ( .A(n10239), .B(n10240), .Z(n10234) );
  XOR U10524 ( .A(n10233), .B(n10234), .Z(n10255) );
  XOR U10525 ( .A(n10256), .B(n10255), .Z(n10257) );
  XNOR U10526 ( .A(n10258), .B(n10257), .Z(n10227) );
  NAND U10527 ( .A(n10217), .B(n10216), .Z(n10221) );
  NAND U10528 ( .A(n10219), .B(n10218), .Z(n10220) );
  NAND U10529 ( .A(n10221), .B(n10220), .Z(n10228) );
  XNOR U10530 ( .A(n10227), .B(n10228), .Z(n10229) );
  XNOR U10531 ( .A(n10230), .B(n10229), .Z(n10261) );
  XNOR U10532 ( .A(n10261), .B(sreg[500]), .Z(n10263) );
  NAND U10533 ( .A(n10222), .B(sreg[499]), .Z(n10226) );
  OR U10534 ( .A(n10224), .B(n10223), .Z(n10225) );
  AND U10535 ( .A(n10226), .B(n10225), .Z(n10262) );
  XOR U10536 ( .A(n10263), .B(n10262), .Z(c[500]) );
  NANDN U10537 ( .A(n10232), .B(n10231), .Z(n10236) );
  NAND U10538 ( .A(n10234), .B(n10233), .Z(n10235) );
  NAND U10539 ( .A(n10236), .B(n10235), .Z(n10297) );
  NANDN U10540 ( .A(n10238), .B(n10237), .Z(n10242) );
  NAND U10541 ( .A(n10240), .B(n10239), .Z(n10241) );
  NAND U10542 ( .A(n10242), .B(n10241), .Z(n10295) );
  XOR U10543 ( .A(b[7]), .B(n10321), .Z(n10282) );
  NANDN U10544 ( .A(n10282), .B(n10545), .Z(n10245) );
  NANDN U10545 ( .A(n10243), .B(n10546), .Z(n10244) );
  NAND U10546 ( .A(n10245), .B(n10244), .Z(n10270) );
  XNOR U10547 ( .A(b[3]), .B(a[251]), .Z(n10285) );
  NANDN U10548 ( .A(n10285), .B(n10398), .Z(n10248) );
  NANDN U10549 ( .A(n10246), .B(n10399), .Z(n10247) );
  AND U10550 ( .A(n10248), .B(n10247), .Z(n10271) );
  XNOR U10551 ( .A(n10270), .B(n10271), .Z(n10272) );
  NANDN U10552 ( .A(n527), .B(a[253]), .Z(n10249) );
  XOR U10553 ( .A(n10434), .B(n10249), .Z(n10251) );
  IV U10554 ( .A(a[252]), .Z(n10439) );
  NANDN U10555 ( .A(n10439), .B(n527), .Z(n10250) );
  AND U10556 ( .A(n10251), .B(n10250), .Z(n10278) );
  XNOR U10557 ( .A(b[5]), .B(a[249]), .Z(n10291) );
  NANDN U10558 ( .A(n10291), .B(n10481), .Z(n10254) );
  NAND U10559 ( .A(n10252), .B(n10482), .Z(n10253) );
  NAND U10560 ( .A(n10254), .B(n10253), .Z(n10276) );
  NANDN U10561 ( .A(n529), .B(a[245]), .Z(n10277) );
  XNOR U10562 ( .A(n10276), .B(n10277), .Z(n10279) );
  XOR U10563 ( .A(n10278), .B(n10279), .Z(n10273) );
  XOR U10564 ( .A(n10272), .B(n10273), .Z(n10294) );
  XOR U10565 ( .A(n10295), .B(n10294), .Z(n10296) );
  XNOR U10566 ( .A(n10297), .B(n10296), .Z(n10266) );
  NAND U10567 ( .A(n10256), .B(n10255), .Z(n10260) );
  NAND U10568 ( .A(n10258), .B(n10257), .Z(n10259) );
  NAND U10569 ( .A(n10260), .B(n10259), .Z(n10267) );
  XNOR U10570 ( .A(n10266), .B(n10267), .Z(n10268) );
  XNOR U10571 ( .A(n10269), .B(n10268), .Z(n10300) );
  XNOR U10572 ( .A(n10300), .B(sreg[501]), .Z(n10302) );
  NAND U10573 ( .A(n10261), .B(sreg[500]), .Z(n10265) );
  OR U10574 ( .A(n10263), .B(n10262), .Z(n10264) );
  AND U10575 ( .A(n10265), .B(n10264), .Z(n10301) );
  XOR U10576 ( .A(n10302), .B(n10301), .Z(c[501]) );
  NANDN U10577 ( .A(n10271), .B(n10270), .Z(n10275) );
  NAND U10578 ( .A(n10273), .B(n10272), .Z(n10274) );
  NAND U10579 ( .A(n10275), .B(n10274), .Z(n10338) );
  NANDN U10580 ( .A(n10277), .B(n10276), .Z(n10281) );
  NAND U10581 ( .A(n10279), .B(n10278), .Z(n10280) );
  NAND U10582 ( .A(n10281), .B(n10280), .Z(n10336) );
  XNOR U10583 ( .A(b[7]), .B(a[248]), .Z(n10332) );
  NANDN U10584 ( .A(n10332), .B(n10545), .Z(n10284) );
  NANDN U10585 ( .A(n10282), .B(n10546), .Z(n10283) );
  NAND U10586 ( .A(n10284), .B(n10283), .Z(n10309) );
  XOR U10587 ( .A(b[3]), .B(n10439), .Z(n10328) );
  NANDN U10588 ( .A(n10328), .B(n10398), .Z(n10287) );
  NANDN U10589 ( .A(n10285), .B(n10399), .Z(n10286) );
  AND U10590 ( .A(n10287), .B(n10286), .Z(n10310) );
  XNOR U10591 ( .A(n10309), .B(n10310), .Z(n10311) );
  NANDN U10592 ( .A(n527), .B(a[254]), .Z(n10288) );
  XOR U10593 ( .A(n10434), .B(n10288), .Z(n10290) );
  NANDN U10594 ( .A(b[0]), .B(a[253]), .Z(n10289) );
  AND U10595 ( .A(n10290), .B(n10289), .Z(n10317) );
  XOR U10596 ( .A(b[5]), .B(a[250]), .Z(n10325) );
  NAND U10597 ( .A(n10325), .B(n10481), .Z(n10293) );
  NANDN U10598 ( .A(n10291), .B(n10482), .Z(n10292) );
  NAND U10599 ( .A(n10293), .B(n10292), .Z(n10315) );
  NANDN U10600 ( .A(n529), .B(a[246]), .Z(n10316) );
  XNOR U10601 ( .A(n10315), .B(n10316), .Z(n10318) );
  XOR U10602 ( .A(n10317), .B(n10318), .Z(n10312) );
  XOR U10603 ( .A(n10311), .B(n10312), .Z(n10335) );
  XOR U10604 ( .A(n10336), .B(n10335), .Z(n10337) );
  XNOR U10605 ( .A(n10338), .B(n10337), .Z(n10305) );
  NAND U10606 ( .A(n10295), .B(n10294), .Z(n10299) );
  NAND U10607 ( .A(n10297), .B(n10296), .Z(n10298) );
  NAND U10608 ( .A(n10299), .B(n10298), .Z(n10306) );
  XNOR U10609 ( .A(n10305), .B(n10306), .Z(n10307) );
  XNOR U10610 ( .A(n10308), .B(n10307), .Z(n10341) );
  XNOR U10611 ( .A(n10341), .B(sreg[502]), .Z(n10343) );
  NAND U10612 ( .A(n10300), .B(sreg[501]), .Z(n10304) );
  OR U10613 ( .A(n10302), .B(n10301), .Z(n10303) );
  AND U10614 ( .A(n10304), .B(n10303), .Z(n10342) );
  XOR U10615 ( .A(n10343), .B(n10342), .Z(c[502]) );
  NANDN U10616 ( .A(n10310), .B(n10309), .Z(n10314) );
  NAND U10617 ( .A(n10312), .B(n10311), .Z(n10313) );
  NAND U10618 ( .A(n10314), .B(n10313), .Z(n10353) );
  NANDN U10619 ( .A(n10316), .B(n10315), .Z(n10320) );
  NAND U10620 ( .A(n10318), .B(n10317), .Z(n10319) );
  NAND U10621 ( .A(n10320), .B(n10319), .Z(n10351) );
  ANDN U10622 ( .B(b[7]), .A(n10321), .Z(n10365) );
  IV U10623 ( .A(a[255]), .Z(n10480) );
  NANDN U10624 ( .A(n10480), .B(b[0]), .Z(n10322) );
  XOR U10625 ( .A(n10434), .B(n10322), .Z(n10324) );
  NANDN U10626 ( .A(b[0]), .B(a[254]), .Z(n10323) );
  AND U10627 ( .A(n10324), .B(n10323), .Z(n10363) );
  XNOR U10628 ( .A(b[5]), .B(a[251]), .Z(n10376) );
  NANDN U10629 ( .A(n10376), .B(n10481), .Z(n10327) );
  NAND U10630 ( .A(n10482), .B(n10325), .Z(n10326) );
  AND U10631 ( .A(n10327), .B(n10326), .Z(n10362) );
  XNOR U10632 ( .A(n10363), .B(n10362), .Z(n10364) );
  XOR U10633 ( .A(n10365), .B(n10364), .Z(n10359) );
  XNOR U10634 ( .A(b[3]), .B(a[253]), .Z(n10371) );
  NANDN U10635 ( .A(n10371), .B(n10398), .Z(n10330) );
  NANDN U10636 ( .A(n10328), .B(n10399), .Z(n10329) );
  NAND U10637 ( .A(n10330), .B(n10329), .Z(n10356) );
  XOR U10638 ( .A(b[7]), .B(n10331), .Z(n10368) );
  NANDN U10639 ( .A(n10368), .B(n10545), .Z(n10334) );
  NANDN U10640 ( .A(n10332), .B(n10546), .Z(n10333) );
  AND U10641 ( .A(n10334), .B(n10333), .Z(n10357) );
  XNOR U10642 ( .A(n10356), .B(n10357), .Z(n10358) );
  XOR U10643 ( .A(n10359), .B(n10358), .Z(n10350) );
  XOR U10644 ( .A(n10351), .B(n10350), .Z(n10352) );
  XNOR U10645 ( .A(n10353), .B(n10352), .Z(n10346) );
  NAND U10646 ( .A(n10336), .B(n10335), .Z(n10340) );
  NAND U10647 ( .A(n10338), .B(n10337), .Z(n10339) );
  NAND U10648 ( .A(n10340), .B(n10339), .Z(n10347) );
  XNOR U10649 ( .A(n10346), .B(n10347), .Z(n10348) );
  XNOR U10650 ( .A(n10349), .B(n10348), .Z(n10379) );
  XNOR U10651 ( .A(n10379), .B(sreg[503]), .Z(n10381) );
  NAND U10652 ( .A(n10341), .B(sreg[502]), .Z(n10345) );
  OR U10653 ( .A(n10343), .B(n10342), .Z(n10344) );
  AND U10654 ( .A(n10345), .B(n10344), .Z(n10380) );
  XOR U10655 ( .A(n10381), .B(n10380), .Z(c[503]) );
  NAND U10656 ( .A(n10351), .B(n10350), .Z(n10355) );
  NAND U10657 ( .A(n10353), .B(n10352), .Z(n10354) );
  NAND U10658 ( .A(n10355), .B(n10354), .Z(n10386) );
  NANDN U10659 ( .A(n10357), .B(n10356), .Z(n10361) );
  NAND U10660 ( .A(n10359), .B(n10358), .Z(n10360) );
  NAND U10661 ( .A(n10361), .B(n10360), .Z(n10418) );
  NANDN U10662 ( .A(n10363), .B(n10362), .Z(n10367) );
  NANDN U10663 ( .A(n10365), .B(n10364), .Z(n10366) );
  NAND U10664 ( .A(n10367), .B(n10366), .Z(n10415) );
  XNOR U10665 ( .A(n529), .B(a[250]), .Z(n10392) );
  NAND U10666 ( .A(n10392), .B(n10545), .Z(n10370) );
  NANDN U10667 ( .A(n10368), .B(n10546), .Z(n10369) );
  NAND U10668 ( .A(n10370), .B(n10369), .Z(n10406) );
  XNOR U10669 ( .A(b[3]), .B(a[254]), .Z(n10400) );
  NANDN U10670 ( .A(n10400), .B(n10398), .Z(n10373) );
  NANDN U10671 ( .A(n10371), .B(n10399), .Z(n10372) );
  NAND U10672 ( .A(n10373), .B(n10372), .Z(n10403) );
  NANDN U10673 ( .A(n10434), .B(n10480), .Z(n10375) );
  NANDN U10674 ( .A(n527), .B(b[1]), .Z(n10374) );
  AND U10675 ( .A(n10375), .B(n10374), .Z(n10409) );
  NANDN U10676 ( .A(n529), .B(a[248]), .Z(n10410) );
  XNOR U10677 ( .A(n10409), .B(n10410), .Z(n10411) );
  XOR U10678 ( .A(b[5]), .B(n10439), .Z(n10395) );
  NANDN U10679 ( .A(n10395), .B(n10481), .Z(n10378) );
  NANDN U10680 ( .A(n10376), .B(n10482), .Z(n10377) );
  AND U10681 ( .A(n10378), .B(n10377), .Z(n10412) );
  XNOR U10682 ( .A(n10403), .B(n10404), .Z(n10405) );
  XOR U10683 ( .A(n10406), .B(n10405), .Z(n10416) );
  XNOR U10684 ( .A(n10415), .B(n10416), .Z(n10417) );
  XOR U10685 ( .A(n10418), .B(n10417), .Z(n10387) );
  XOR U10686 ( .A(n10386), .B(n10387), .Z(n10388) );
  XOR U10687 ( .A(n10389), .B(n10388), .Z(n10385) );
  NAND U10688 ( .A(n10379), .B(sreg[503]), .Z(n10383) );
  OR U10689 ( .A(n10381), .B(n10380), .Z(n10382) );
  AND U10690 ( .A(n10383), .B(n10382), .Z(n10384) );
  XOR U10691 ( .A(n10385), .B(n10384), .Z(c[504]) );
  OR U10692 ( .A(n10385), .B(n10384), .Z(n10422) );
  OR U10693 ( .A(n10387), .B(n10386), .Z(n10391) );
  NAND U10694 ( .A(n10389), .B(n10388), .Z(n10390) );
  NAND U10695 ( .A(n10391), .B(n10390), .Z(n10426) );
  ANDN U10696 ( .B(a[249]), .A(n529), .Z(n10489) );
  IV U10697 ( .A(n10489), .Z(n10514) );
  XNOR U10698 ( .A(b[7]), .B(a[251]), .Z(n10440) );
  NANDN U10699 ( .A(n10440), .B(n10545), .Z(n10394) );
  NAND U10700 ( .A(n10546), .B(n10392), .Z(n10393) );
  AND U10701 ( .A(n10394), .B(n10393), .Z(n10446) );
  XOR U10702 ( .A(n10514), .B(n10446), .Z(n10448) );
  XOR U10703 ( .A(b[5]), .B(a[253]), .Z(n10443) );
  NAND U10704 ( .A(n10481), .B(n10443), .Z(n10397) );
  NANDN U10705 ( .A(n10395), .B(n10482), .Z(n10396) );
  NAND U10706 ( .A(n10397), .B(n10396), .Z(n10447) );
  XNOR U10707 ( .A(n10448), .B(n10447), .Z(n10431) );
  XNOR U10708 ( .A(n528), .B(a[255]), .Z(n10436) );
  NAND U10709 ( .A(n10436), .B(n10398), .Z(n10402) );
  NANDN U10710 ( .A(n10400), .B(n10399), .Z(n10401) );
  AND U10711 ( .A(n10402), .B(n10401), .Z(n10429) );
  XNOR U10712 ( .A(n10434), .B(n10429), .Z(n10430) );
  XNOR U10713 ( .A(n10431), .B(n10430), .Z(n10454) );
  NANDN U10714 ( .A(n10404), .B(n10403), .Z(n10408) );
  NAND U10715 ( .A(n10406), .B(n10405), .Z(n10407) );
  NAND U10716 ( .A(n10408), .B(n10407), .Z(n10451) );
  OR U10717 ( .A(n10410), .B(n10409), .Z(n10414) );
  OR U10718 ( .A(n10412), .B(n10411), .Z(n10413) );
  AND U10719 ( .A(n10414), .B(n10413), .Z(n10452) );
  XNOR U10720 ( .A(n10451), .B(n10452), .Z(n10453) );
  XOR U10721 ( .A(n10454), .B(n10453), .Z(n10423) );
  NANDN U10722 ( .A(n10416), .B(n10415), .Z(n10420) );
  NANDN U10723 ( .A(n10418), .B(n10417), .Z(n10419) );
  AND U10724 ( .A(n10420), .B(n10419), .Z(n10424) );
  XNOR U10725 ( .A(n10423), .B(n10424), .Z(n10425) );
  XOR U10726 ( .A(n10426), .B(n10425), .Z(n10421) );
  XOR U10727 ( .A(n10422), .B(n10421), .Z(c[505]) );
  OR U10728 ( .A(n10422), .B(n10421), .Z(n10458) );
  NANDN U10729 ( .A(n10424), .B(n10423), .Z(n10428) );
  NAND U10730 ( .A(n10426), .B(n10425), .Z(n10427) );
  NAND U10731 ( .A(n10428), .B(n10427), .Z(n10462) );
  OR U10732 ( .A(n10429), .B(b[1]), .Z(n10433) );
  NAND U10733 ( .A(n10431), .B(n10430), .Z(n10432) );
  NAND U10734 ( .A(n10433), .B(n10432), .Z(n10468) );
  NANDN U10735 ( .A(n10434), .B(b[2]), .Z(n10486) );
  XOR U10736 ( .A(n528), .B(n10486), .Z(n10438) );
  XOR U10737 ( .A(b[2]), .B(n10434), .Z(n10435) );
  NANDN U10738 ( .A(n10436), .B(n10435), .Z(n10437) );
  AND U10739 ( .A(n10438), .B(n10437), .Z(n10487) );
  NANDN U10740 ( .A(n529), .B(a[250]), .Z(n10488) );
  XOR U10741 ( .A(n10487), .B(n10488), .Z(n10490) );
  XOR U10742 ( .A(n10489), .B(n10490), .Z(n10473) );
  XOR U10743 ( .A(b[7]), .B(n10439), .Z(n10477) );
  NANDN U10744 ( .A(n10477), .B(n10545), .Z(n10442) );
  NANDN U10745 ( .A(n10440), .B(n10546), .Z(n10441) );
  AND U10746 ( .A(n10442), .B(n10441), .Z(n10471) );
  XOR U10747 ( .A(b[5]), .B(a[254]), .Z(n10483) );
  NAND U10748 ( .A(n10483), .B(n10481), .Z(n10445) );
  NAND U10749 ( .A(n10443), .B(n10482), .Z(n10444) );
  AND U10750 ( .A(n10445), .B(n10444), .Z(n10472) );
  XOR U10751 ( .A(n10473), .B(n10474), .Z(n10465) );
  NANDN U10752 ( .A(n10514), .B(n10446), .Z(n10450) );
  OR U10753 ( .A(n10448), .B(n10447), .Z(n10449) );
  AND U10754 ( .A(n10450), .B(n10449), .Z(n10466) );
  XOR U10755 ( .A(n10465), .B(n10466), .Z(n10467) );
  XOR U10756 ( .A(n10468), .B(n10467), .Z(n10460) );
  NANDN U10757 ( .A(n10452), .B(n10451), .Z(n10456) );
  NANDN U10758 ( .A(n10454), .B(n10453), .Z(n10455) );
  AND U10759 ( .A(n10456), .B(n10455), .Z(n10459) );
  XNOR U10760 ( .A(n10460), .B(n10459), .Z(n10461) );
  XOR U10761 ( .A(n10462), .B(n10461), .Z(n10457) );
  XOR U10762 ( .A(n10458), .B(n10457), .Z(c[506]) );
  OR U10763 ( .A(n10458), .B(n10457), .Z(n10528) );
  NANDN U10764 ( .A(n10460), .B(n10459), .Z(n10464) );
  NAND U10765 ( .A(n10462), .B(n10461), .Z(n10463) );
  NAND U10766 ( .A(n10464), .B(n10463), .Z(n10496) );
  OR U10767 ( .A(n10466), .B(n10465), .Z(n10470) );
  NANDN U10768 ( .A(n10468), .B(n10467), .Z(n10469) );
  NAND U10769 ( .A(n10470), .B(n10469), .Z(n10493) );
  OR U10770 ( .A(n10472), .B(n10471), .Z(n10476) );
  NAND U10771 ( .A(n10474), .B(n10473), .Z(n10475) );
  NAND U10772 ( .A(n10476), .B(n10475), .Z(n10502) );
  XNOR U10773 ( .A(b[7]), .B(a[253]), .Z(n10517) );
  NANDN U10774 ( .A(n10517), .B(n10545), .Z(n10479) );
  NANDN U10775 ( .A(n10477), .B(n10546), .Z(n10478) );
  NAND U10776 ( .A(n10479), .B(n10478), .Z(n10505) );
  XNOR U10777 ( .A(b[5]), .B(n10480), .Z(n10523) );
  NAND U10778 ( .A(n10523), .B(n10481), .Z(n10485) );
  NAND U10779 ( .A(n10483), .B(n10482), .Z(n10484) );
  AND U10780 ( .A(n10485), .B(n10484), .Z(n10506) );
  XNOR U10781 ( .A(n10505), .B(n10506), .Z(n10507) );
  ANDN U10782 ( .B(n10486), .A(n528), .Z(n10512) );
  NANDN U10783 ( .A(n529), .B(a[251]), .Z(n10511) );
  XOR U10784 ( .A(n10512), .B(n10511), .Z(n10513) );
  XOR U10785 ( .A(n10514), .B(n10513), .Z(n10508) );
  XNOR U10786 ( .A(n10507), .B(n10508), .Z(n10499) );
  NANDN U10787 ( .A(n10488), .B(n10487), .Z(n10492) );
  OR U10788 ( .A(n10490), .B(n10489), .Z(n10491) );
  NAND U10789 ( .A(n10492), .B(n10491), .Z(n10500) );
  XOR U10790 ( .A(n10502), .B(n10501), .Z(n10494) );
  XNOR U10791 ( .A(n10493), .B(n10494), .Z(n10495) );
  XOR U10792 ( .A(n10496), .B(n10495), .Z(n10527) );
  XOR U10793 ( .A(n10528), .B(n10527), .Z(c[507]) );
  NANDN U10794 ( .A(n10494), .B(n10493), .Z(n10498) );
  NAND U10795 ( .A(n10496), .B(n10495), .Z(n10497) );
  NAND U10796 ( .A(n10498), .B(n10497), .Z(n10533) );
  OR U10797 ( .A(n10500), .B(n10499), .Z(n10504) );
  NANDN U10798 ( .A(n10502), .B(n10501), .Z(n10503) );
  NAND U10799 ( .A(n10504), .B(n10503), .Z(n10532) );
  NANDN U10800 ( .A(n10506), .B(n10505), .Z(n10510) );
  NANDN U10801 ( .A(n10508), .B(n10507), .Z(n10509) );
  NAND U10802 ( .A(n10510), .B(n10509), .Z(n10536) );
  OR U10803 ( .A(n10512), .B(n10511), .Z(n10516) );
  NANDN U10804 ( .A(n10514), .B(n10513), .Z(n10515) );
  NAND U10805 ( .A(n10516), .B(n10515), .Z(n10535) );
  AND U10806 ( .A(b[7]), .B(a[252]), .Z(n10554) );
  XNOR U10807 ( .A(b[7]), .B(a[254]), .Z(n10547) );
  NANDN U10808 ( .A(n10547), .B(n10545), .Z(n10519) );
  NANDN U10809 ( .A(n10517), .B(n10546), .Z(n10518) );
  AND U10810 ( .A(n10519), .B(n10518), .Z(n10540) );
  XOR U10811 ( .A(n10554), .B(n10540), .Z(n10541) );
  XNOR U10812 ( .A(b[5]), .B(n10520), .Z(n10525) );
  XOR U10813 ( .A(n10521), .B(b[3]), .Z(n10522) );
  NANDN U10814 ( .A(n10523), .B(n10522), .Z(n10524) );
  NAND U10815 ( .A(n10525), .B(n10524), .Z(n10542) );
  XNOR U10816 ( .A(n10535), .B(n10534), .Z(n10537) );
  XNOR U10817 ( .A(n10536), .B(n10537), .Z(n10531) );
  XOR U10818 ( .A(n10532), .B(n10531), .Z(n10526) );
  XNOR U10819 ( .A(n10533), .B(n10526), .Z(n10530) );
  OR U10820 ( .A(n10528), .B(n10527), .Z(n10529) );
  XOR U10821 ( .A(n10530), .B(n10529), .Z(c[508]) );
  OR U10822 ( .A(n10530), .B(n10529), .Z(n10573) );
  NAND U10823 ( .A(n10535), .B(n10534), .Z(n10539) );
  NANDN U10824 ( .A(n10537), .B(n10536), .Z(n10538) );
  AND U10825 ( .A(n10539), .B(n10538), .Z(n10563) );
  NANDN U10826 ( .A(n529), .B(a[253]), .Z(n10551) );
  XOR U10827 ( .A(n10552), .B(n10551), .Z(n10553) );
  XNOR U10828 ( .A(n10554), .B(n10553), .Z(n10568) );
  OR U10829 ( .A(n10540), .B(n10554), .Z(n10544) );
  NANDN U10830 ( .A(n10542), .B(n10541), .Z(n10543) );
  AND U10831 ( .A(n10544), .B(n10543), .Z(n10565) );
  XNOR U10832 ( .A(n529), .B(a[255]), .Z(n10558) );
  NAND U10833 ( .A(n10558), .B(n10545), .Z(n10549) );
  NANDN U10834 ( .A(n10547), .B(n10546), .Z(n10548) );
  AND U10835 ( .A(n10549), .B(n10548), .Z(n10566) );
  XNOR U10836 ( .A(n10565), .B(n10566), .Z(n10567) );
  XNOR U10837 ( .A(n10563), .B(n10562), .Z(n10550) );
  XOR U10838 ( .A(n10564), .B(n10550), .Z(n10572) );
  XNOR U10839 ( .A(n10573), .B(n10572), .Z(c[509]) );
  AND U10840 ( .A(a[254]), .B(b[7]), .Z(n10577) );
  IV U10841 ( .A(n10577), .Z(n10575) );
  OR U10842 ( .A(n10552), .B(n10551), .Z(n10556) );
  NAND U10843 ( .A(n10554), .B(n10553), .Z(n10555) );
  NAND U10844 ( .A(n10556), .B(n10555), .Z(n10574) );
  AND U10845 ( .A(b[5]), .B(b[6]), .Z(n10581) );
  XOR U10846 ( .A(b[7]), .B(n10581), .Z(n10560) );
  NANDN U10847 ( .A(n10558), .B(n10557), .Z(n10559) );
  AND U10848 ( .A(n10560), .B(n10559), .Z(n10576) );
  XNOR U10849 ( .A(n10574), .B(n10576), .Z(n10561) );
  XNOR U10850 ( .A(n10575), .B(n10561), .Z(n10579) );
  OR U10851 ( .A(n10566), .B(n10565), .Z(n10570) );
  OR U10852 ( .A(n10568), .B(n10567), .Z(n10569) );
  NAND U10853 ( .A(n10570), .B(n10569), .Z(n10580) );
  XOR U10854 ( .A(n10578), .B(n10580), .Z(n10571) );
  XNOR U10855 ( .A(n10579), .B(n10571), .Z(n10582) );
  NANDN U10856 ( .A(n10573), .B(n10572), .Z(n10583) );
  XNOR U10857 ( .A(n10582), .B(n10583), .Z(c[510]) );
endmodule

