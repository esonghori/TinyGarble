
module mult_N256_CC16 ( clk, rst, a, b, c );
  input [255:0] a;
  input [15:0] b;
  output [511:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159;
  wire   [511:0] sreg;

  DFF \sreg_reg[495]  ( .D(c[511]), .CLK(clk), .RST(rst), .Q(sreg[495]) );
  DFF \sreg_reg[494]  ( .D(c[510]), .CLK(clk), .RST(rst), .Q(sreg[494]) );
  DFF \sreg_reg[493]  ( .D(c[509]), .CLK(clk), .RST(rst), .Q(sreg[493]) );
  DFF \sreg_reg[492]  ( .D(c[508]), .CLK(clk), .RST(rst), .Q(sreg[492]) );
  DFF \sreg_reg[491]  ( .D(c[507]), .CLK(clk), .RST(rst), .Q(sreg[491]) );
  DFF \sreg_reg[490]  ( .D(c[506]), .CLK(clk), .RST(rst), .Q(sreg[490]) );
  DFF \sreg_reg[489]  ( .D(c[505]), .CLK(clk), .RST(rst), .Q(sreg[489]) );
  DFF \sreg_reg[488]  ( .D(c[504]), .CLK(clk), .RST(rst), .Q(sreg[488]) );
  DFF \sreg_reg[487]  ( .D(c[503]), .CLK(clk), .RST(rst), .Q(sreg[487]) );
  DFF \sreg_reg[486]  ( .D(c[502]), .CLK(clk), .RST(rst), .Q(sreg[486]) );
  DFF \sreg_reg[485]  ( .D(c[501]), .CLK(clk), .RST(rst), .Q(sreg[485]) );
  DFF \sreg_reg[484]  ( .D(c[500]), .CLK(clk), .RST(rst), .Q(sreg[484]) );
  DFF \sreg_reg[483]  ( .D(c[499]), .CLK(clk), .RST(rst), .Q(sreg[483]) );
  DFF \sreg_reg[482]  ( .D(c[498]), .CLK(clk), .RST(rst), .Q(sreg[482]) );
  DFF \sreg_reg[481]  ( .D(c[497]), .CLK(clk), .RST(rst), .Q(sreg[481]) );
  DFF \sreg_reg[480]  ( .D(c[496]), .CLK(clk), .RST(rst), .Q(sreg[480]) );
  DFF \sreg_reg[479]  ( .D(c[495]), .CLK(clk), .RST(rst), .Q(sreg[479]) );
  DFF \sreg_reg[478]  ( .D(c[494]), .CLK(clk), .RST(rst), .Q(sreg[478]) );
  DFF \sreg_reg[477]  ( .D(c[493]), .CLK(clk), .RST(rst), .Q(sreg[477]) );
  DFF \sreg_reg[476]  ( .D(c[492]), .CLK(clk), .RST(rst), .Q(sreg[476]) );
  DFF \sreg_reg[475]  ( .D(c[491]), .CLK(clk), .RST(rst), .Q(sreg[475]) );
  DFF \sreg_reg[474]  ( .D(c[490]), .CLK(clk), .RST(rst), .Q(sreg[474]) );
  DFF \sreg_reg[473]  ( .D(c[489]), .CLK(clk), .RST(rst), .Q(sreg[473]) );
  DFF \sreg_reg[472]  ( .D(c[488]), .CLK(clk), .RST(rst), .Q(sreg[472]) );
  DFF \sreg_reg[471]  ( .D(c[487]), .CLK(clk), .RST(rst), .Q(sreg[471]) );
  DFF \sreg_reg[470]  ( .D(c[486]), .CLK(clk), .RST(rst), .Q(sreg[470]) );
  DFF \sreg_reg[469]  ( .D(c[485]), .CLK(clk), .RST(rst), .Q(sreg[469]) );
  DFF \sreg_reg[468]  ( .D(c[484]), .CLK(clk), .RST(rst), .Q(sreg[468]) );
  DFF \sreg_reg[467]  ( .D(c[483]), .CLK(clk), .RST(rst), .Q(sreg[467]) );
  DFF \sreg_reg[466]  ( .D(c[482]), .CLK(clk), .RST(rst), .Q(sreg[466]) );
  DFF \sreg_reg[465]  ( .D(c[481]), .CLK(clk), .RST(rst), .Q(sreg[465]) );
  DFF \sreg_reg[464]  ( .D(c[480]), .CLK(clk), .RST(rst), .Q(sreg[464]) );
  DFF \sreg_reg[463]  ( .D(c[479]), .CLK(clk), .RST(rst), .Q(sreg[463]) );
  DFF \sreg_reg[462]  ( .D(c[478]), .CLK(clk), .RST(rst), .Q(sreg[462]) );
  DFF \sreg_reg[461]  ( .D(c[477]), .CLK(clk), .RST(rst), .Q(sreg[461]) );
  DFF \sreg_reg[460]  ( .D(c[476]), .CLK(clk), .RST(rst), .Q(sreg[460]) );
  DFF \sreg_reg[459]  ( .D(c[475]), .CLK(clk), .RST(rst), .Q(sreg[459]) );
  DFF \sreg_reg[458]  ( .D(c[474]), .CLK(clk), .RST(rst), .Q(sreg[458]) );
  DFF \sreg_reg[457]  ( .D(c[473]), .CLK(clk), .RST(rst), .Q(sreg[457]) );
  DFF \sreg_reg[456]  ( .D(c[472]), .CLK(clk), .RST(rst), .Q(sreg[456]) );
  DFF \sreg_reg[455]  ( .D(c[471]), .CLK(clk), .RST(rst), .Q(sreg[455]) );
  DFF \sreg_reg[454]  ( .D(c[470]), .CLK(clk), .RST(rst), .Q(sreg[454]) );
  DFF \sreg_reg[453]  ( .D(c[469]), .CLK(clk), .RST(rst), .Q(sreg[453]) );
  DFF \sreg_reg[452]  ( .D(c[468]), .CLK(clk), .RST(rst), .Q(sreg[452]) );
  DFF \sreg_reg[451]  ( .D(c[467]), .CLK(clk), .RST(rst), .Q(sreg[451]) );
  DFF \sreg_reg[450]  ( .D(c[466]), .CLK(clk), .RST(rst), .Q(sreg[450]) );
  DFF \sreg_reg[449]  ( .D(c[465]), .CLK(clk), .RST(rst), .Q(sreg[449]) );
  DFF \sreg_reg[448]  ( .D(c[464]), .CLK(clk), .RST(rst), .Q(sreg[448]) );
  DFF \sreg_reg[447]  ( .D(c[463]), .CLK(clk), .RST(rst), .Q(sreg[447]) );
  DFF \sreg_reg[446]  ( .D(c[462]), .CLK(clk), .RST(rst), .Q(sreg[446]) );
  DFF \sreg_reg[445]  ( .D(c[461]), .CLK(clk), .RST(rst), .Q(sreg[445]) );
  DFF \sreg_reg[444]  ( .D(c[460]), .CLK(clk), .RST(rst), .Q(sreg[444]) );
  DFF \sreg_reg[443]  ( .D(c[459]), .CLK(clk), .RST(rst), .Q(sreg[443]) );
  DFF \sreg_reg[442]  ( .D(c[458]), .CLK(clk), .RST(rst), .Q(sreg[442]) );
  DFF \sreg_reg[441]  ( .D(c[457]), .CLK(clk), .RST(rst), .Q(sreg[441]) );
  DFF \sreg_reg[440]  ( .D(c[456]), .CLK(clk), .RST(rst), .Q(sreg[440]) );
  DFF \sreg_reg[439]  ( .D(c[455]), .CLK(clk), .RST(rst), .Q(sreg[439]) );
  DFF \sreg_reg[438]  ( .D(c[454]), .CLK(clk), .RST(rst), .Q(sreg[438]) );
  DFF \sreg_reg[437]  ( .D(c[453]), .CLK(clk), .RST(rst), .Q(sreg[437]) );
  DFF \sreg_reg[436]  ( .D(c[452]), .CLK(clk), .RST(rst), .Q(sreg[436]) );
  DFF \sreg_reg[435]  ( .D(c[451]), .CLK(clk), .RST(rst), .Q(sreg[435]) );
  DFF \sreg_reg[434]  ( .D(c[450]), .CLK(clk), .RST(rst), .Q(sreg[434]) );
  DFF \sreg_reg[433]  ( .D(c[449]), .CLK(clk), .RST(rst), .Q(sreg[433]) );
  DFF \sreg_reg[432]  ( .D(c[448]), .CLK(clk), .RST(rst), .Q(sreg[432]) );
  DFF \sreg_reg[431]  ( .D(c[447]), .CLK(clk), .RST(rst), .Q(sreg[431]) );
  DFF \sreg_reg[430]  ( .D(c[446]), .CLK(clk), .RST(rst), .Q(sreg[430]) );
  DFF \sreg_reg[429]  ( .D(c[445]), .CLK(clk), .RST(rst), .Q(sreg[429]) );
  DFF \sreg_reg[428]  ( .D(c[444]), .CLK(clk), .RST(rst), .Q(sreg[428]) );
  DFF \sreg_reg[427]  ( .D(c[443]), .CLK(clk), .RST(rst), .Q(sreg[427]) );
  DFF \sreg_reg[426]  ( .D(c[442]), .CLK(clk), .RST(rst), .Q(sreg[426]) );
  DFF \sreg_reg[425]  ( .D(c[441]), .CLK(clk), .RST(rst), .Q(sreg[425]) );
  DFF \sreg_reg[424]  ( .D(c[440]), .CLK(clk), .RST(rst), .Q(sreg[424]) );
  DFF \sreg_reg[423]  ( .D(c[439]), .CLK(clk), .RST(rst), .Q(sreg[423]) );
  DFF \sreg_reg[422]  ( .D(c[438]), .CLK(clk), .RST(rst), .Q(sreg[422]) );
  DFF \sreg_reg[421]  ( .D(c[437]), .CLK(clk), .RST(rst), .Q(sreg[421]) );
  DFF \sreg_reg[420]  ( .D(c[436]), .CLK(clk), .RST(rst), .Q(sreg[420]) );
  DFF \sreg_reg[419]  ( .D(c[435]), .CLK(clk), .RST(rst), .Q(sreg[419]) );
  DFF \sreg_reg[418]  ( .D(c[434]), .CLK(clk), .RST(rst), .Q(sreg[418]) );
  DFF \sreg_reg[417]  ( .D(c[433]), .CLK(clk), .RST(rst), .Q(sreg[417]) );
  DFF \sreg_reg[416]  ( .D(c[432]), .CLK(clk), .RST(rst), .Q(sreg[416]) );
  DFF \sreg_reg[415]  ( .D(c[431]), .CLK(clk), .RST(rst), .Q(sreg[415]) );
  DFF \sreg_reg[414]  ( .D(c[430]), .CLK(clk), .RST(rst), .Q(sreg[414]) );
  DFF \sreg_reg[413]  ( .D(c[429]), .CLK(clk), .RST(rst), .Q(sreg[413]) );
  DFF \sreg_reg[412]  ( .D(c[428]), .CLK(clk), .RST(rst), .Q(sreg[412]) );
  DFF \sreg_reg[411]  ( .D(c[427]), .CLK(clk), .RST(rst), .Q(sreg[411]) );
  DFF \sreg_reg[410]  ( .D(c[426]), .CLK(clk), .RST(rst), .Q(sreg[410]) );
  DFF \sreg_reg[409]  ( .D(c[425]), .CLK(clk), .RST(rst), .Q(sreg[409]) );
  DFF \sreg_reg[408]  ( .D(c[424]), .CLK(clk), .RST(rst), .Q(sreg[408]) );
  DFF \sreg_reg[407]  ( .D(c[423]), .CLK(clk), .RST(rst), .Q(sreg[407]) );
  DFF \sreg_reg[406]  ( .D(c[422]), .CLK(clk), .RST(rst), .Q(sreg[406]) );
  DFF \sreg_reg[405]  ( .D(c[421]), .CLK(clk), .RST(rst), .Q(sreg[405]) );
  DFF \sreg_reg[404]  ( .D(c[420]), .CLK(clk), .RST(rst), .Q(sreg[404]) );
  DFF \sreg_reg[403]  ( .D(c[419]), .CLK(clk), .RST(rst), .Q(sreg[403]) );
  DFF \sreg_reg[402]  ( .D(c[418]), .CLK(clk), .RST(rst), .Q(sreg[402]) );
  DFF \sreg_reg[401]  ( .D(c[417]), .CLK(clk), .RST(rst), .Q(sreg[401]) );
  DFF \sreg_reg[400]  ( .D(c[416]), .CLK(clk), .RST(rst), .Q(sreg[400]) );
  DFF \sreg_reg[399]  ( .D(c[415]), .CLK(clk), .RST(rst), .Q(sreg[399]) );
  DFF \sreg_reg[398]  ( .D(c[414]), .CLK(clk), .RST(rst), .Q(sreg[398]) );
  DFF \sreg_reg[397]  ( .D(c[413]), .CLK(clk), .RST(rst), .Q(sreg[397]) );
  DFF \sreg_reg[396]  ( .D(c[412]), .CLK(clk), .RST(rst), .Q(sreg[396]) );
  DFF \sreg_reg[395]  ( .D(c[411]), .CLK(clk), .RST(rst), .Q(sreg[395]) );
  DFF \sreg_reg[394]  ( .D(c[410]), .CLK(clk), .RST(rst), .Q(sreg[394]) );
  DFF \sreg_reg[393]  ( .D(c[409]), .CLK(clk), .RST(rst), .Q(sreg[393]) );
  DFF \sreg_reg[392]  ( .D(c[408]), .CLK(clk), .RST(rst), .Q(sreg[392]) );
  DFF \sreg_reg[391]  ( .D(c[407]), .CLK(clk), .RST(rst), .Q(sreg[391]) );
  DFF \sreg_reg[390]  ( .D(c[406]), .CLK(clk), .RST(rst), .Q(sreg[390]) );
  DFF \sreg_reg[389]  ( .D(c[405]), .CLK(clk), .RST(rst), .Q(sreg[389]) );
  DFF \sreg_reg[388]  ( .D(c[404]), .CLK(clk), .RST(rst), .Q(sreg[388]) );
  DFF \sreg_reg[387]  ( .D(c[403]), .CLK(clk), .RST(rst), .Q(sreg[387]) );
  DFF \sreg_reg[386]  ( .D(c[402]), .CLK(clk), .RST(rst), .Q(sreg[386]) );
  DFF \sreg_reg[385]  ( .D(c[401]), .CLK(clk), .RST(rst), .Q(sreg[385]) );
  DFF \sreg_reg[384]  ( .D(c[400]), .CLK(clk), .RST(rst), .Q(sreg[384]) );
  DFF \sreg_reg[383]  ( .D(c[399]), .CLK(clk), .RST(rst), .Q(sreg[383]) );
  DFF \sreg_reg[382]  ( .D(c[398]), .CLK(clk), .RST(rst), .Q(sreg[382]) );
  DFF \sreg_reg[381]  ( .D(c[397]), .CLK(clk), .RST(rst), .Q(sreg[381]) );
  DFF \sreg_reg[380]  ( .D(c[396]), .CLK(clk), .RST(rst), .Q(sreg[380]) );
  DFF \sreg_reg[379]  ( .D(c[395]), .CLK(clk), .RST(rst), .Q(sreg[379]) );
  DFF \sreg_reg[378]  ( .D(c[394]), .CLK(clk), .RST(rst), .Q(sreg[378]) );
  DFF \sreg_reg[377]  ( .D(c[393]), .CLK(clk), .RST(rst), .Q(sreg[377]) );
  DFF \sreg_reg[376]  ( .D(c[392]), .CLK(clk), .RST(rst), .Q(sreg[376]) );
  DFF \sreg_reg[375]  ( .D(c[391]), .CLK(clk), .RST(rst), .Q(sreg[375]) );
  DFF \sreg_reg[374]  ( .D(c[390]), .CLK(clk), .RST(rst), .Q(sreg[374]) );
  DFF \sreg_reg[373]  ( .D(c[389]), .CLK(clk), .RST(rst), .Q(sreg[373]) );
  DFF \sreg_reg[372]  ( .D(c[388]), .CLK(clk), .RST(rst), .Q(sreg[372]) );
  DFF \sreg_reg[371]  ( .D(c[387]), .CLK(clk), .RST(rst), .Q(sreg[371]) );
  DFF \sreg_reg[370]  ( .D(c[386]), .CLK(clk), .RST(rst), .Q(sreg[370]) );
  DFF \sreg_reg[369]  ( .D(c[385]), .CLK(clk), .RST(rst), .Q(sreg[369]) );
  DFF \sreg_reg[368]  ( .D(c[384]), .CLK(clk), .RST(rst), .Q(sreg[368]) );
  DFF \sreg_reg[367]  ( .D(c[383]), .CLK(clk), .RST(rst), .Q(sreg[367]) );
  DFF \sreg_reg[366]  ( .D(c[382]), .CLK(clk), .RST(rst), .Q(sreg[366]) );
  DFF \sreg_reg[365]  ( .D(c[381]), .CLK(clk), .RST(rst), .Q(sreg[365]) );
  DFF \sreg_reg[364]  ( .D(c[380]), .CLK(clk), .RST(rst), .Q(sreg[364]) );
  DFF \sreg_reg[363]  ( .D(c[379]), .CLK(clk), .RST(rst), .Q(sreg[363]) );
  DFF \sreg_reg[362]  ( .D(c[378]), .CLK(clk), .RST(rst), .Q(sreg[362]) );
  DFF \sreg_reg[361]  ( .D(c[377]), .CLK(clk), .RST(rst), .Q(sreg[361]) );
  DFF \sreg_reg[360]  ( .D(c[376]), .CLK(clk), .RST(rst), .Q(sreg[360]) );
  DFF \sreg_reg[359]  ( .D(c[375]), .CLK(clk), .RST(rst), .Q(sreg[359]) );
  DFF \sreg_reg[358]  ( .D(c[374]), .CLK(clk), .RST(rst), .Q(sreg[358]) );
  DFF \sreg_reg[357]  ( .D(c[373]), .CLK(clk), .RST(rst), .Q(sreg[357]) );
  DFF \sreg_reg[356]  ( .D(c[372]), .CLK(clk), .RST(rst), .Q(sreg[356]) );
  DFF \sreg_reg[355]  ( .D(c[371]), .CLK(clk), .RST(rst), .Q(sreg[355]) );
  DFF \sreg_reg[354]  ( .D(c[370]), .CLK(clk), .RST(rst), .Q(sreg[354]) );
  DFF \sreg_reg[353]  ( .D(c[369]), .CLK(clk), .RST(rst), .Q(sreg[353]) );
  DFF \sreg_reg[352]  ( .D(c[368]), .CLK(clk), .RST(rst), .Q(sreg[352]) );
  DFF \sreg_reg[351]  ( .D(c[367]), .CLK(clk), .RST(rst), .Q(sreg[351]) );
  DFF \sreg_reg[350]  ( .D(c[366]), .CLK(clk), .RST(rst), .Q(sreg[350]) );
  DFF \sreg_reg[349]  ( .D(c[365]), .CLK(clk), .RST(rst), .Q(sreg[349]) );
  DFF \sreg_reg[348]  ( .D(c[364]), .CLK(clk), .RST(rst), .Q(sreg[348]) );
  DFF \sreg_reg[347]  ( .D(c[363]), .CLK(clk), .RST(rst), .Q(sreg[347]) );
  DFF \sreg_reg[346]  ( .D(c[362]), .CLK(clk), .RST(rst), .Q(sreg[346]) );
  DFF \sreg_reg[345]  ( .D(c[361]), .CLK(clk), .RST(rst), .Q(sreg[345]) );
  DFF \sreg_reg[344]  ( .D(c[360]), .CLK(clk), .RST(rst), .Q(sreg[344]) );
  DFF \sreg_reg[343]  ( .D(c[359]), .CLK(clk), .RST(rst), .Q(sreg[343]) );
  DFF \sreg_reg[342]  ( .D(c[358]), .CLK(clk), .RST(rst), .Q(sreg[342]) );
  DFF \sreg_reg[341]  ( .D(c[357]), .CLK(clk), .RST(rst), .Q(sreg[341]) );
  DFF \sreg_reg[340]  ( .D(c[356]), .CLK(clk), .RST(rst), .Q(sreg[340]) );
  DFF \sreg_reg[339]  ( .D(c[355]), .CLK(clk), .RST(rst), .Q(sreg[339]) );
  DFF \sreg_reg[338]  ( .D(c[354]), .CLK(clk), .RST(rst), .Q(sreg[338]) );
  DFF \sreg_reg[337]  ( .D(c[353]), .CLK(clk), .RST(rst), .Q(sreg[337]) );
  DFF \sreg_reg[336]  ( .D(c[352]), .CLK(clk), .RST(rst), .Q(sreg[336]) );
  DFF \sreg_reg[335]  ( .D(c[351]), .CLK(clk), .RST(rst), .Q(sreg[335]) );
  DFF \sreg_reg[334]  ( .D(c[350]), .CLK(clk), .RST(rst), .Q(sreg[334]) );
  DFF \sreg_reg[333]  ( .D(c[349]), .CLK(clk), .RST(rst), .Q(sreg[333]) );
  DFF \sreg_reg[332]  ( .D(c[348]), .CLK(clk), .RST(rst), .Q(sreg[332]) );
  DFF \sreg_reg[331]  ( .D(c[347]), .CLK(clk), .RST(rst), .Q(sreg[331]) );
  DFF \sreg_reg[330]  ( .D(c[346]), .CLK(clk), .RST(rst), .Q(sreg[330]) );
  DFF \sreg_reg[329]  ( .D(c[345]), .CLK(clk), .RST(rst), .Q(sreg[329]) );
  DFF \sreg_reg[328]  ( .D(c[344]), .CLK(clk), .RST(rst), .Q(sreg[328]) );
  DFF \sreg_reg[327]  ( .D(c[343]), .CLK(clk), .RST(rst), .Q(sreg[327]) );
  DFF \sreg_reg[326]  ( .D(c[342]), .CLK(clk), .RST(rst), .Q(sreg[326]) );
  DFF \sreg_reg[325]  ( .D(c[341]), .CLK(clk), .RST(rst), .Q(sreg[325]) );
  DFF \sreg_reg[324]  ( .D(c[340]), .CLK(clk), .RST(rst), .Q(sreg[324]) );
  DFF \sreg_reg[323]  ( .D(c[339]), .CLK(clk), .RST(rst), .Q(sreg[323]) );
  DFF \sreg_reg[322]  ( .D(c[338]), .CLK(clk), .RST(rst), .Q(sreg[322]) );
  DFF \sreg_reg[321]  ( .D(c[337]), .CLK(clk), .RST(rst), .Q(sreg[321]) );
  DFF \sreg_reg[320]  ( .D(c[336]), .CLK(clk), .RST(rst), .Q(sreg[320]) );
  DFF \sreg_reg[319]  ( .D(c[335]), .CLK(clk), .RST(rst), .Q(sreg[319]) );
  DFF \sreg_reg[318]  ( .D(c[334]), .CLK(clk), .RST(rst), .Q(sreg[318]) );
  DFF \sreg_reg[317]  ( .D(c[333]), .CLK(clk), .RST(rst), .Q(sreg[317]) );
  DFF \sreg_reg[316]  ( .D(c[332]), .CLK(clk), .RST(rst), .Q(sreg[316]) );
  DFF \sreg_reg[315]  ( .D(c[331]), .CLK(clk), .RST(rst), .Q(sreg[315]) );
  DFF \sreg_reg[314]  ( .D(c[330]), .CLK(clk), .RST(rst), .Q(sreg[314]) );
  DFF \sreg_reg[313]  ( .D(c[329]), .CLK(clk), .RST(rst), .Q(sreg[313]) );
  DFF \sreg_reg[312]  ( .D(c[328]), .CLK(clk), .RST(rst), .Q(sreg[312]) );
  DFF \sreg_reg[311]  ( .D(c[327]), .CLK(clk), .RST(rst), .Q(sreg[311]) );
  DFF \sreg_reg[310]  ( .D(c[326]), .CLK(clk), .RST(rst), .Q(sreg[310]) );
  DFF \sreg_reg[309]  ( .D(c[325]), .CLK(clk), .RST(rst), .Q(sreg[309]) );
  DFF \sreg_reg[308]  ( .D(c[324]), .CLK(clk), .RST(rst), .Q(sreg[308]) );
  DFF \sreg_reg[307]  ( .D(c[323]), .CLK(clk), .RST(rst), .Q(sreg[307]) );
  DFF \sreg_reg[306]  ( .D(c[322]), .CLK(clk), .RST(rst), .Q(sreg[306]) );
  DFF \sreg_reg[305]  ( .D(c[321]), .CLK(clk), .RST(rst), .Q(sreg[305]) );
  DFF \sreg_reg[304]  ( .D(c[320]), .CLK(clk), .RST(rst), .Q(sreg[304]) );
  DFF \sreg_reg[303]  ( .D(c[319]), .CLK(clk), .RST(rst), .Q(sreg[303]) );
  DFF \sreg_reg[302]  ( .D(c[318]), .CLK(clk), .RST(rst), .Q(sreg[302]) );
  DFF \sreg_reg[301]  ( .D(c[317]), .CLK(clk), .RST(rst), .Q(sreg[301]) );
  DFF \sreg_reg[300]  ( .D(c[316]), .CLK(clk), .RST(rst), .Q(sreg[300]) );
  DFF \sreg_reg[299]  ( .D(c[315]), .CLK(clk), .RST(rst), .Q(sreg[299]) );
  DFF \sreg_reg[298]  ( .D(c[314]), .CLK(clk), .RST(rst), .Q(sreg[298]) );
  DFF \sreg_reg[297]  ( .D(c[313]), .CLK(clk), .RST(rst), .Q(sreg[297]) );
  DFF \sreg_reg[296]  ( .D(c[312]), .CLK(clk), .RST(rst), .Q(sreg[296]) );
  DFF \sreg_reg[295]  ( .D(c[311]), .CLK(clk), .RST(rst), .Q(sreg[295]) );
  DFF \sreg_reg[294]  ( .D(c[310]), .CLK(clk), .RST(rst), .Q(sreg[294]) );
  DFF \sreg_reg[293]  ( .D(c[309]), .CLK(clk), .RST(rst), .Q(sreg[293]) );
  DFF \sreg_reg[292]  ( .D(c[308]), .CLK(clk), .RST(rst), .Q(sreg[292]) );
  DFF \sreg_reg[291]  ( .D(c[307]), .CLK(clk), .RST(rst), .Q(sreg[291]) );
  DFF \sreg_reg[290]  ( .D(c[306]), .CLK(clk), .RST(rst), .Q(sreg[290]) );
  DFF \sreg_reg[289]  ( .D(c[305]), .CLK(clk), .RST(rst), .Q(sreg[289]) );
  DFF \sreg_reg[288]  ( .D(c[304]), .CLK(clk), .RST(rst), .Q(sreg[288]) );
  DFF \sreg_reg[287]  ( .D(c[303]), .CLK(clk), .RST(rst), .Q(sreg[287]) );
  DFF \sreg_reg[286]  ( .D(c[302]), .CLK(clk), .RST(rst), .Q(sreg[286]) );
  DFF \sreg_reg[285]  ( .D(c[301]), .CLK(clk), .RST(rst), .Q(sreg[285]) );
  DFF \sreg_reg[284]  ( .D(c[300]), .CLK(clk), .RST(rst), .Q(sreg[284]) );
  DFF \sreg_reg[283]  ( .D(c[299]), .CLK(clk), .RST(rst), .Q(sreg[283]) );
  DFF \sreg_reg[282]  ( .D(c[298]), .CLK(clk), .RST(rst), .Q(sreg[282]) );
  DFF \sreg_reg[281]  ( .D(c[297]), .CLK(clk), .RST(rst), .Q(sreg[281]) );
  DFF \sreg_reg[280]  ( .D(c[296]), .CLK(clk), .RST(rst), .Q(sreg[280]) );
  DFF \sreg_reg[279]  ( .D(c[295]), .CLK(clk), .RST(rst), .Q(sreg[279]) );
  DFF \sreg_reg[278]  ( .D(c[294]), .CLK(clk), .RST(rst), .Q(sreg[278]) );
  DFF \sreg_reg[277]  ( .D(c[293]), .CLK(clk), .RST(rst), .Q(sreg[277]) );
  DFF \sreg_reg[276]  ( .D(c[292]), .CLK(clk), .RST(rst), .Q(sreg[276]) );
  DFF \sreg_reg[275]  ( .D(c[291]), .CLK(clk), .RST(rst), .Q(sreg[275]) );
  DFF \sreg_reg[274]  ( .D(c[290]), .CLK(clk), .RST(rst), .Q(sreg[274]) );
  DFF \sreg_reg[273]  ( .D(c[289]), .CLK(clk), .RST(rst), .Q(sreg[273]) );
  DFF \sreg_reg[272]  ( .D(c[288]), .CLK(clk), .RST(rst), .Q(sreg[272]) );
  DFF \sreg_reg[271]  ( .D(c[287]), .CLK(clk), .RST(rst), .Q(sreg[271]) );
  DFF \sreg_reg[270]  ( .D(c[286]), .CLK(clk), .RST(rst), .Q(sreg[270]) );
  DFF \sreg_reg[269]  ( .D(c[285]), .CLK(clk), .RST(rst), .Q(sreg[269]) );
  DFF \sreg_reg[268]  ( .D(c[284]), .CLK(clk), .RST(rst), .Q(sreg[268]) );
  DFF \sreg_reg[267]  ( .D(c[283]), .CLK(clk), .RST(rst), .Q(sreg[267]) );
  DFF \sreg_reg[266]  ( .D(c[282]), .CLK(clk), .RST(rst), .Q(sreg[266]) );
  DFF \sreg_reg[265]  ( .D(c[281]), .CLK(clk), .RST(rst), .Q(sreg[265]) );
  DFF \sreg_reg[264]  ( .D(c[280]), .CLK(clk), .RST(rst), .Q(sreg[264]) );
  DFF \sreg_reg[263]  ( .D(c[279]), .CLK(clk), .RST(rst), .Q(sreg[263]) );
  DFF \sreg_reg[262]  ( .D(c[278]), .CLK(clk), .RST(rst), .Q(sreg[262]) );
  DFF \sreg_reg[261]  ( .D(c[277]), .CLK(clk), .RST(rst), .Q(sreg[261]) );
  DFF \sreg_reg[260]  ( .D(c[276]), .CLK(clk), .RST(rst), .Q(sreg[260]) );
  DFF \sreg_reg[259]  ( .D(c[275]), .CLK(clk), .RST(rst), .Q(sreg[259]) );
  DFF \sreg_reg[258]  ( .D(c[274]), .CLK(clk), .RST(rst), .Q(sreg[258]) );
  DFF \sreg_reg[257]  ( .D(c[273]), .CLK(clk), .RST(rst), .Q(sreg[257]) );
  DFF \sreg_reg[256]  ( .D(c[272]), .CLK(clk), .RST(rst), .Q(sreg[256]) );
  DFF \sreg_reg[255]  ( .D(c[271]), .CLK(clk), .RST(rst), .Q(sreg[255]) );
  DFF \sreg_reg[254]  ( .D(c[270]), .CLK(clk), .RST(rst), .Q(sreg[254]) );
  DFF \sreg_reg[253]  ( .D(c[269]), .CLK(clk), .RST(rst), .Q(sreg[253]) );
  DFF \sreg_reg[252]  ( .D(c[268]), .CLK(clk), .RST(rst), .Q(sreg[252]) );
  DFF \sreg_reg[251]  ( .D(c[267]), .CLK(clk), .RST(rst), .Q(sreg[251]) );
  DFF \sreg_reg[250]  ( .D(c[266]), .CLK(clk), .RST(rst), .Q(sreg[250]) );
  DFF \sreg_reg[249]  ( .D(c[265]), .CLK(clk), .RST(rst), .Q(sreg[249]) );
  DFF \sreg_reg[248]  ( .D(c[264]), .CLK(clk), .RST(rst), .Q(sreg[248]) );
  DFF \sreg_reg[247]  ( .D(c[263]), .CLK(clk), .RST(rst), .Q(sreg[247]) );
  DFF \sreg_reg[246]  ( .D(c[262]), .CLK(clk), .RST(rst), .Q(sreg[246]) );
  DFF \sreg_reg[245]  ( .D(c[261]), .CLK(clk), .RST(rst), .Q(sreg[245]) );
  DFF \sreg_reg[244]  ( .D(c[260]), .CLK(clk), .RST(rst), .Q(sreg[244]) );
  DFF \sreg_reg[243]  ( .D(c[259]), .CLK(clk), .RST(rst), .Q(sreg[243]) );
  DFF \sreg_reg[242]  ( .D(c[258]), .CLK(clk), .RST(rst), .Q(sreg[242]) );
  DFF \sreg_reg[241]  ( .D(c[257]), .CLK(clk), .RST(rst), .Q(sreg[241]) );
  DFF \sreg_reg[240]  ( .D(c[256]), .CLK(clk), .RST(rst), .Q(sreg[240]) );
  DFF \sreg_reg[239]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(c[239]) );
  DFF \sreg_reg[238]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(c[238]) );
  DFF \sreg_reg[237]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(c[237]) );
  DFF \sreg_reg[236]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(c[236]) );
  DFF \sreg_reg[235]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(c[235]) );
  DFF \sreg_reg[234]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(c[234]) );
  DFF \sreg_reg[233]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(c[233]) );
  DFF \sreg_reg[232]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(c[232]) );
  DFF \sreg_reg[231]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(c[231]) );
  DFF \sreg_reg[230]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(c[230]) );
  DFF \sreg_reg[229]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(c[229]) );
  DFF \sreg_reg[228]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(c[228]) );
  DFF \sreg_reg[227]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(c[227]) );
  DFF \sreg_reg[226]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(c[226]) );
  DFF \sreg_reg[225]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(c[225]) );
  DFF \sreg_reg[224]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(c[224]) );
  DFF \sreg_reg[223]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(c[223]) );
  DFF \sreg_reg[222]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(c[222]) );
  DFF \sreg_reg[221]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(c[221]) );
  DFF \sreg_reg[220]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(c[220]) );
  DFF \sreg_reg[219]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(c[219]) );
  DFF \sreg_reg[218]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(c[218]) );
  DFF \sreg_reg[217]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(c[217]) );
  DFF \sreg_reg[216]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(c[216]) );
  DFF \sreg_reg[215]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(c[215]) );
  DFF \sreg_reg[214]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(c[214]) );
  DFF \sreg_reg[213]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(c[213]) );
  DFF \sreg_reg[212]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(c[212]) );
  DFF \sreg_reg[211]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(c[211]) );
  DFF \sreg_reg[210]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(c[210]) );
  DFF \sreg_reg[209]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(c[209]) );
  DFF \sreg_reg[208]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(c[208]) );
  DFF \sreg_reg[207]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(c[207]) );
  DFF \sreg_reg[206]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(c[206]) );
  DFF \sreg_reg[205]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(c[205]) );
  DFF \sreg_reg[204]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(c[204]) );
  DFF \sreg_reg[203]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(c[203]) );
  DFF \sreg_reg[202]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(c[202]) );
  DFF \sreg_reg[201]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(c[201]) );
  DFF \sreg_reg[200]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(c[200]) );
  DFF \sreg_reg[199]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(c[199]) );
  DFF \sreg_reg[198]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(c[198]) );
  DFF \sreg_reg[197]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(c[197]) );
  DFF \sreg_reg[196]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(c[196]) );
  DFF \sreg_reg[195]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(c[195]) );
  DFF \sreg_reg[194]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(c[194]) );
  DFF \sreg_reg[193]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(c[193]) );
  DFF \sreg_reg[192]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(c[192]) );
  DFF \sreg_reg[191]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(c[191]) );
  DFF \sreg_reg[190]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(c[190]) );
  DFF \sreg_reg[189]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(c[189]) );
  DFF \sreg_reg[188]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(c[188]) );
  DFF \sreg_reg[187]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(c[187]) );
  DFF \sreg_reg[186]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(c[186]) );
  DFF \sreg_reg[185]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(c[185]) );
  DFF \sreg_reg[184]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(c[184]) );
  DFF \sreg_reg[183]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(c[183]) );
  DFF \sreg_reg[182]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(c[182]) );
  DFF \sreg_reg[181]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(c[181]) );
  DFF \sreg_reg[180]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(c[180]) );
  DFF \sreg_reg[179]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(c[179]) );
  DFF \sreg_reg[178]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(c[178]) );
  DFF \sreg_reg[177]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(c[177]) );
  DFF \sreg_reg[176]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(c[176]) );
  DFF \sreg_reg[175]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(c[175]) );
  DFF \sreg_reg[174]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(c[174]) );
  DFF \sreg_reg[173]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(c[173]) );
  DFF \sreg_reg[172]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(c[172]) );
  DFF \sreg_reg[171]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(c[171]) );
  DFF \sreg_reg[170]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(c[170]) );
  DFF \sreg_reg[169]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(c[169]) );
  DFF \sreg_reg[168]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(c[168]) );
  DFF \sreg_reg[167]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(c[167]) );
  DFF \sreg_reg[166]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(c[166]) );
  DFF \sreg_reg[165]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(c[165]) );
  DFF \sreg_reg[164]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(c[164]) );
  DFF \sreg_reg[163]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(c[163]) );
  DFF \sreg_reg[162]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(c[162]) );
  DFF \sreg_reg[161]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(c[161]) );
  DFF \sreg_reg[160]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(c[160]) );
  DFF \sreg_reg[159]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(c[159]) );
  DFF \sreg_reg[158]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(c[158]) );
  DFF \sreg_reg[157]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(c[157]) );
  DFF \sreg_reg[156]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(c[156]) );
  DFF \sreg_reg[155]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(c[155]) );
  DFF \sreg_reg[154]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(c[154]) );
  DFF \sreg_reg[153]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(c[153]) );
  DFF \sreg_reg[152]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(c[152]) );
  DFF \sreg_reg[151]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(c[151]) );
  DFF \sreg_reg[150]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(c[150]) );
  DFF \sreg_reg[149]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(c[149]) );
  DFF \sreg_reg[148]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(c[148]) );
  DFF \sreg_reg[147]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(c[147]) );
  DFF \sreg_reg[146]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(c[146]) );
  DFF \sreg_reg[145]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(c[145]) );
  DFF \sreg_reg[144]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(c[144]) );
  DFF \sreg_reg[143]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(c[143]) );
  DFF \sreg_reg[142]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(c[142]) );
  DFF \sreg_reg[141]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(c[141]) );
  DFF \sreg_reg[140]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(c[140]) );
  DFF \sreg_reg[139]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(c[139]) );
  DFF \sreg_reg[138]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(c[138]) );
  DFF \sreg_reg[137]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(c[137]) );
  DFF \sreg_reg[136]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(c[136]) );
  DFF \sreg_reg[135]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(c[135]) );
  DFF \sreg_reg[134]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(c[134]) );
  DFF \sreg_reg[133]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(c[133]) );
  DFF \sreg_reg[132]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(c[132]) );
  DFF \sreg_reg[131]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(c[131]) );
  DFF \sreg_reg[130]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(c[130]) );
  DFF \sreg_reg[129]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(c[129]) );
  DFF \sreg_reg[128]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(c[128]) );
  DFF \sreg_reg[127]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(c[127]) );
  DFF \sreg_reg[126]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(c[126]) );
  DFF \sreg_reg[125]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(c[125]) );
  DFF \sreg_reg[124]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(c[124]) );
  DFF \sreg_reg[123]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(c[123]) );
  DFF \sreg_reg[122]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(c[122]) );
  DFF \sreg_reg[121]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(c[121]) );
  DFF \sreg_reg[120]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(c[120]) );
  DFF \sreg_reg[119]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[118]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[117]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[116]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[115]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[114]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[113]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[112]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[111]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[110]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[109]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[108]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[107]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[106]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[105]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[104]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[103]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[102]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[101]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[100]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[99]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[98]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[97]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[96]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[95]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[94]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[93]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[92]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[91]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[90]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[89]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[88]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[87]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[86]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[85]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[84]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[83]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[82]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[81]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[80]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[79]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[78]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[77]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[76]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[75]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[74]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[73]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[72]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[71]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[70]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[69]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[68]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[67]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[66]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[65]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[64]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[63]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[62]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[0]) );
  XNOR U19 ( .A(n20144), .B(n20145), .Z(n20139) );
  OR U20 ( .A(n19508), .B(n19507), .Z(n1) );
  NANDN U21 ( .A(n19510), .B(n19509), .Z(n2) );
  NAND U22 ( .A(n1), .B(n2), .Z(n19594) );
  OR U23 ( .A(n19695), .B(n19694), .Z(n3) );
  NANDN U24 ( .A(n19697), .B(n19696), .Z(n4) );
  NAND U25 ( .A(n3), .B(n4), .Z(n19789) );
  NAND U26 ( .A(n19995), .B(n19994), .Z(n5) );
  XOR U27 ( .A(n19994), .B(n19995), .Z(n6) );
  NAND U28 ( .A(n6), .B(n19993), .Z(n7) );
  NAND U29 ( .A(n5), .B(n7), .Z(n20001) );
  NAND U30 ( .A(n20107), .B(n20105), .Z(n8) );
  XOR U31 ( .A(n20105), .B(n20107), .Z(n9) );
  NANDN U32 ( .A(n20106), .B(n9), .Z(n10) );
  NAND U33 ( .A(n8), .B(n10), .Z(n20141) );
  NANDN U34 ( .A(n728), .B(n727), .Z(n11) );
  NANDN U35 ( .A(n725), .B(n726), .Z(n12) );
  NAND U36 ( .A(n11), .B(n12), .Z(n838) );
  NANDN U37 ( .A(n934), .B(n935), .Z(n13) );
  NANDN U38 ( .A(n933), .B(n932), .Z(n14) );
  NAND U39 ( .A(n13), .B(n14), .Z(n1070) );
  XNOR U40 ( .A(n19549), .B(n19550), .Z(n19544) );
  OR U41 ( .A(n19690), .B(n19691), .Z(n15) );
  NANDN U42 ( .A(n19692), .B(n19693), .Z(n16) );
  NAND U43 ( .A(n15), .B(n16), .Z(n19791) );
  OR U44 ( .A(n273), .B(n274), .Z(n17) );
  NAND U45 ( .A(n276), .B(n275), .Z(n18) );
  NAND U46 ( .A(n17), .B(n18), .Z(n332) );
  OR U47 ( .A(n19594), .B(n19595), .Z(n19) );
  NANDN U48 ( .A(n19597), .B(n19596), .Z(n20) );
  AND U49 ( .A(n19), .B(n20), .Z(n19672) );
  XOR U50 ( .A(n19912), .B(n19911), .Z(n21) );
  NANDN U51 ( .A(n19910), .B(n21), .Z(n22) );
  NAND U52 ( .A(n19912), .B(n19911), .Z(n23) );
  AND U53 ( .A(n22), .B(n23), .Z(n19995) );
  OR U54 ( .A(n19989), .B(n19990), .Z(n24) );
  NAND U55 ( .A(n19991), .B(n19992), .Z(n25) );
  AND U56 ( .A(n24), .B(n25), .Z(n19999) );
  NAND U57 ( .A(n20141), .B(n20139), .Z(n26) );
  XOR U58 ( .A(n20139), .B(n20141), .Z(n27) );
  NANDN U59 ( .A(n20140), .B(n27), .Z(n28) );
  NAND U60 ( .A(n26), .B(n28), .Z(n20152) );
  NANDN U61 ( .A(n904), .B(n905), .Z(n29) );
  NANDN U62 ( .A(n903), .B(n902), .Z(n30) );
  NAND U63 ( .A(n29), .B(n30), .Z(n960) );
  NAND U64 ( .A(n1760), .B(n1759), .Z(n31) );
  NANDN U65 ( .A(n1757), .B(n1758), .Z(n32) );
  NAND U66 ( .A(n31), .B(n32), .Z(n1785) );
  NAND U67 ( .A(n5870), .B(n5869), .Z(n33) );
  NANDN U68 ( .A(n5867), .B(n5868), .Z(n34) );
  NAND U69 ( .A(n33), .B(n34), .Z(n5917) );
  NAND U70 ( .A(n9946), .B(n9945), .Z(n35) );
  NANDN U71 ( .A(n9943), .B(n9944), .Z(n36) );
  NAND U72 ( .A(n35), .B(n36), .Z(n9971) );
  NAND U73 ( .A(n15171), .B(n15170), .Z(n37) );
  NANDN U74 ( .A(n15168), .B(n15169), .Z(n38) );
  NAND U75 ( .A(n37), .B(n38), .Z(n15196) );
  NAND U76 ( .A(n15247), .B(n15246), .Z(n39) );
  NANDN U77 ( .A(n15244), .B(n15245), .Z(n40) );
  NAND U78 ( .A(n39), .B(n40), .Z(n15272) );
  XOR U79 ( .A(n19289), .B(n19290), .Z(n19292) );
  OR U80 ( .A(b[0]), .B(n20120), .Z(n41) );
  AND U81 ( .A(b[1]), .B(n41), .Z(n19527) );
  NANDN U82 ( .A(n641), .B(n642), .Z(n42) );
  NANDN U83 ( .A(n640), .B(n639), .Z(n43) );
  NAND U84 ( .A(n42), .B(n43), .Z(n719) );
  XNOR U85 ( .A(n623), .B(n624), .Z(n618) );
  NANDN U86 ( .A(n771), .B(n770), .Z(n44) );
  NANDN U87 ( .A(n772), .B(n773), .Z(n45) );
  AND U88 ( .A(n44), .B(n45), .Z(n780) );
  OR U89 ( .A(n836), .B(n835), .Z(n46) );
  NANDN U90 ( .A(n838), .B(n837), .Z(n47) );
  NAND U91 ( .A(n46), .B(n47), .Z(n856) );
  NANDN U92 ( .A(n19374), .B(n19375), .Z(n48) );
  NANDN U93 ( .A(n19373), .B(n19372), .Z(n49) );
  NAND U94 ( .A(n48), .B(n49), .Z(n19404) );
  XOR U95 ( .A(n19415), .B(n19416), .Z(n19418) );
  OR U96 ( .A(n19706), .B(n19707), .Z(n50) );
  NANDN U97 ( .A(n19704), .B(n19705), .Z(n51) );
  NAND U98 ( .A(n50), .B(n51), .Z(n19792) );
  NANDN U99 ( .A(n233), .B(n234), .Z(n52) );
  NANDN U100 ( .A(n232), .B(n231), .Z(n53) );
  NAND U101 ( .A(n52), .B(n53), .Z(n268) );
  OR U102 ( .A(n511), .B(n510), .Z(n54) );
  NANDN U103 ( .A(n513), .B(n512), .Z(n55) );
  NAND U104 ( .A(n54), .B(n55), .Z(n574) );
  OR U105 ( .A(n19592), .B(n19593), .Z(n56) );
  NANDN U106 ( .A(n19590), .B(n19591), .Z(n57) );
  NAND U107 ( .A(n56), .B(n57), .Z(n19673) );
  XOR U108 ( .A(n19668), .B(n19669), .Z(n19663) );
  OR U109 ( .A(n19789), .B(n19788), .Z(n58) );
  NANDN U110 ( .A(n19791), .B(n19790), .Z(n59) );
  NAND U111 ( .A(n58), .B(n59), .Z(n19843) );
  NANDN U112 ( .A(n19785), .B(n19810), .Z(n60) );
  NANDN U113 ( .A(n19786), .B(n19787), .Z(n61) );
  AND U114 ( .A(n60), .B(n61), .Z(n19802) );
  OR U115 ( .A(n180), .B(n181), .Z(n62) );
  NANDN U116 ( .A(n183), .B(n182), .Z(n63) );
  AND U117 ( .A(n62), .B(n63), .Z(n192) );
  NANDN U118 ( .A(n1004), .B(n1005), .Z(n64) );
  NANDN U119 ( .A(n1003), .B(n1002), .Z(n65) );
  NAND U120 ( .A(n64), .B(n65), .Z(n1081) );
  OR U121 ( .A(n19800), .B(n19801), .Z(n66) );
  NANDN U122 ( .A(n19798), .B(n19799), .Z(n67) );
  NAND U123 ( .A(n66), .B(n67), .Z(n19901) );
  NANDN U124 ( .A(n20049), .B(n20050), .Z(n68) );
  NANDN U125 ( .A(n20048), .B(n20084), .Z(n69) );
  NAND U126 ( .A(n68), .B(n69), .Z(n20076) );
  NANDN U127 ( .A(n347), .B(n348), .Z(n70) );
  NANDN U128 ( .A(n346), .B(n345), .Z(n71) );
  NAND U129 ( .A(n70), .B(n71), .Z(n387) );
  NANDN U130 ( .A(n709), .B(n710), .Z(n72) );
  NANDN U131 ( .A(n711), .B(n712), .Z(n73) );
  NAND U132 ( .A(n72), .B(n73), .Z(n777) );
  NANDN U133 ( .A(n19395), .B(n19396), .Z(n74) );
  NANDN U134 ( .A(n19394), .B(n19393), .Z(n75) );
  NAND U135 ( .A(n74), .B(n75), .Z(n19471) );
  NAND U136 ( .A(n19747), .B(n19745), .Z(n76) );
  XOR U137 ( .A(n19745), .B(n19747), .Z(n77) );
  NANDN U138 ( .A(n19746), .B(n77), .Z(n78) );
  NAND U139 ( .A(n76), .B(n78), .Z(n19851) );
  NAND U140 ( .A(n20001), .B(n19999), .Z(n79) );
  XOR U141 ( .A(n19999), .B(n20001), .Z(n80) );
  NANDN U142 ( .A(n20000), .B(n80), .Z(n81) );
  NAND U143 ( .A(n79), .B(n81), .Z(n20039) );
  NANDN U144 ( .A(n20154), .B(b[15]), .Z(n82) );
  XNOR U145 ( .A(b[15]), .B(n20154), .Z(n83) );
  NAND U146 ( .A(n83), .B(b[14]), .Z(n84) );
  NAND U147 ( .A(n82), .B(n84), .Z(n85) );
  AND U148 ( .A(a[255]), .B(n85), .Z(n86) );
  NANDN U149 ( .A(n20152), .B(n20151), .Z(n87) );
  XNOR U150 ( .A(n20152), .B(n20151), .Z(n88) );
  NAND U151 ( .A(n88), .B(n20153), .Z(n89) );
  AND U152 ( .A(n87), .B(n89), .Z(n90) );
  XNOR U153 ( .A(n86), .B(n90), .Z(n91) );
  NAND U154 ( .A(n20156), .B(n20155), .Z(n92) );
  XOR U155 ( .A(n20156), .B(n20155), .Z(n93) );
  NAND U156 ( .A(n93), .B(n20157), .Z(n94) );
  AND U157 ( .A(n92), .B(n94), .Z(n95) );
  XNOR U158 ( .A(n91), .B(n95), .Z(n96) );
  NANDN U159 ( .A(n20159), .B(n20158), .Z(n97) );
  XNOR U160 ( .A(n96), .B(n97), .Z(c[511]) );
  IV U161 ( .A(b[0]), .Z(n98) );
  IV U162 ( .A(b[1]), .Z(n99) );
  IV U163 ( .A(b[3]), .Z(n100) );
  IV U164 ( .A(b[5]), .Z(n101) );
  IV U165 ( .A(b[15]), .Z(n102) );
  NAND U166 ( .A(b[0]), .B(a[0]), .Z(n104) );
  XNOR U167 ( .A(n104), .B(sreg[240]), .Z(c[240]) );
  AND U168 ( .A(a[1]), .B(b[0]), .Z(n108) );
  NAND U169 ( .A(b[1]), .B(a[0]), .Z(n103) );
  XNOR U170 ( .A(n108), .B(n103), .Z(n110) );
  XNOR U171 ( .A(sreg[241]), .B(n110), .Z(n112) );
  NANDN U172 ( .A(n104), .B(sreg[240]), .Z(n111) );
  XOR U173 ( .A(n112), .B(n111), .Z(c[241]) );
  NAND U174 ( .A(b[0]), .B(a[2]), .Z(n105) );
  XNOR U175 ( .A(b[1]), .B(n105), .Z(n107) );
  NAND U176 ( .A(n98), .B(a[1]), .Z(n106) );
  AND U177 ( .A(n107), .B(n106), .Z(n115) );
  XOR U178 ( .A(n99), .B(b[2]), .Z(n19521) );
  IV U179 ( .A(a[0]), .Z(n685) );
  OR U180 ( .A(n19521), .B(n685), .Z(n116) );
  XNOR U181 ( .A(n115), .B(n116), .Z(n117) );
  AND U182 ( .A(n685), .B(b[1]), .Z(n109) );
  ANDN U183 ( .B(n109), .A(n108), .Z(n118) );
  XNOR U184 ( .A(n117), .B(n118), .Z(n134) );
  NAND U185 ( .A(sreg[241]), .B(n110), .Z(n114) );
  OR U186 ( .A(n112), .B(n111), .Z(n113) );
  NAND U187 ( .A(n114), .B(n113), .Z(n132) );
  XNOR U188 ( .A(n132), .B(sreg[242]), .Z(n133) );
  XOR U189 ( .A(n134), .B(n133), .Z(c[242]) );
  NANDN U190 ( .A(n116), .B(n115), .Z(n120) );
  NAND U191 ( .A(n118), .B(n117), .Z(n119) );
  NAND U192 ( .A(n120), .B(n119), .Z(n144) );
  NOR U193 ( .A(n100), .B(n19521), .Z(n19556) );
  NAND U194 ( .A(n685), .B(n19556), .Z(n123) );
  AND U195 ( .A(n99), .B(b[3]), .Z(n121) );
  NANDN U196 ( .A(b[2]), .B(n121), .Z(n122) );
  AND U197 ( .A(n123), .B(n122), .Z(n143) );
  XNOR U198 ( .A(a[0]), .B(b[1]), .Z(n125) );
  XNOR U199 ( .A(b[1]), .B(b[2]), .Z(n124) );
  NAND U200 ( .A(n125), .B(n124), .Z(n126) );
  XNOR U201 ( .A(b[3]), .B(b[2]), .Z(n153) );
  OR U202 ( .A(n126), .B(n153), .Z(n128) );
  XOR U203 ( .A(n100), .B(a[1]), .Z(n155) );
  OR U204 ( .A(n155), .B(n19521), .Z(n127) );
  NAND U205 ( .A(n128), .B(n127), .Z(n149) );
  NAND U206 ( .A(b[0]), .B(a[3]), .Z(n129) );
  XNOR U207 ( .A(b[1]), .B(n129), .Z(n131) );
  NAND U208 ( .A(a[2]), .B(n98), .Z(n130) );
  AND U209 ( .A(n131), .B(n130), .Z(n148) );
  XOR U210 ( .A(n149), .B(n148), .Z(n142) );
  XOR U211 ( .A(n143), .B(n142), .Z(n145) );
  XNOR U212 ( .A(n144), .B(n145), .Z(n137) );
  XNOR U213 ( .A(sreg[243]), .B(n137), .Z(n139) );
  NAND U214 ( .A(n132), .B(sreg[242]), .Z(n136) );
  OR U215 ( .A(n134), .B(n133), .Z(n135) );
  AND U216 ( .A(n136), .B(n135), .Z(n138) );
  XOR U217 ( .A(n139), .B(n138), .Z(c[243]) );
  NAND U218 ( .A(sreg[243]), .B(n137), .Z(n141) );
  OR U219 ( .A(n139), .B(n138), .Z(n140) );
  NAND U220 ( .A(n141), .B(n140), .Z(n184) );
  XNOR U221 ( .A(n184), .B(sreg[244]), .Z(n186) );
  NANDN U222 ( .A(n143), .B(n142), .Z(n147) );
  NANDN U223 ( .A(n145), .B(n144), .Z(n146) );
  NAND U224 ( .A(n147), .B(n146), .Z(n183) );
  AND U225 ( .A(n149), .B(n148), .Z(n180) );
  XOR U226 ( .A(n100), .B(b[4]), .Z(n19640) );
  OR U227 ( .A(n19640), .B(n685), .Z(n177) );
  NAND U228 ( .A(b[0]), .B(a[4]), .Z(n150) );
  XNOR U229 ( .A(b[1]), .B(n150), .Z(n152) );
  NAND U230 ( .A(a[3]), .B(n98), .Z(n151) );
  AND U231 ( .A(n152), .B(n151), .Z(n175) );
  XNOR U232 ( .A(b[3]), .B(a[2]), .Z(n171) );
  OR U233 ( .A(n171), .B(n19521), .Z(n157) );
  XOR U234 ( .A(b[3]), .B(b[1]), .Z(n154) );
  ANDN U235 ( .B(n154), .A(n153), .Z(n19554) );
  NANDN U236 ( .A(n155), .B(n19554), .Z(n156) );
  AND U237 ( .A(n157), .B(n156), .Z(n174) );
  XNOR U238 ( .A(n175), .B(n174), .Z(n176) );
  XNOR U239 ( .A(n177), .B(n176), .Z(n181) );
  XOR U240 ( .A(n180), .B(n181), .Z(n182) );
  XNOR U241 ( .A(n183), .B(n182), .Z(n185) );
  XOR U242 ( .A(n186), .B(n185), .Z(c[244]) );
  NAND U243 ( .A(b[0]), .B(a[5]), .Z(n158) );
  XNOR U244 ( .A(b[1]), .B(n158), .Z(n160) );
  NAND U245 ( .A(a[4]), .B(n98), .Z(n159) );
  AND U246 ( .A(n160), .B(n159), .Z(n196) );
  XOR U247 ( .A(b[5]), .B(a[0]), .Z(n164) );
  XOR U248 ( .A(b[5]), .B(b[3]), .Z(n162) );
  IV U249 ( .A(b[4]), .Z(n167) );
  XNOR U250 ( .A(b[5]), .B(n167), .Z(n161) );
  AND U251 ( .A(n162), .B(n161), .Z(n163) );
  NAND U252 ( .A(n164), .B(n163), .Z(n166) );
  XOR U253 ( .A(n101), .B(a[1]), .Z(n205) );
  OR U254 ( .A(n205), .B(n19640), .Z(n165) );
  AND U255 ( .A(n166), .B(n165), .Z(n195) );
  XNOR U256 ( .A(n196), .B(n195), .Z(n211) );
  NAND U257 ( .A(b[5]), .B(n167), .Z(n168) );
  NANDN U258 ( .A(n168), .B(n100), .Z(n170) );
  NOR U259 ( .A(n101), .B(n19640), .Z(n19724) );
  NAND U260 ( .A(n685), .B(n19724), .Z(n169) );
  NAND U261 ( .A(n170), .B(n169), .Z(n209) );
  IV U262 ( .A(a[3]), .Z(n795) );
  XNOR U263 ( .A(n100), .B(n795), .Z(n197) );
  OR U264 ( .A(n197), .B(n19521), .Z(n173) );
  NANDN U265 ( .A(n171), .B(n19554), .Z(n172) );
  AND U266 ( .A(n173), .B(n172), .Z(n208) );
  XNOR U267 ( .A(n209), .B(n208), .Z(n210) );
  XNOR U268 ( .A(n211), .B(n210), .Z(n189) );
  NANDN U269 ( .A(n175), .B(n174), .Z(n179) );
  NAND U270 ( .A(n177), .B(n176), .Z(n178) );
  NAND U271 ( .A(n179), .B(n178), .Z(n190) );
  XOR U272 ( .A(n189), .B(n190), .Z(n191) );
  XOR U273 ( .A(n191), .B(n192), .Z(n214) );
  XNOR U274 ( .A(sreg[245]), .B(n214), .Z(n216) );
  NAND U275 ( .A(n184), .B(sreg[244]), .Z(n188) );
  OR U276 ( .A(n186), .B(n185), .Z(n187) );
  AND U277 ( .A(n188), .B(n187), .Z(n215) );
  XOR U278 ( .A(n216), .B(n215), .Z(c[245]) );
  OR U279 ( .A(n190), .B(n189), .Z(n194) );
  NAND U280 ( .A(n192), .B(n191), .Z(n193) );
  NAND U281 ( .A(n194), .B(n193), .Z(n222) );
  ANDN U282 ( .B(n196), .A(n195), .Z(n228) );
  NANDN U283 ( .A(n197), .B(n19554), .Z(n199) );
  IV U284 ( .A(a[4]), .Z(n877) );
  XNOR U285 ( .A(b[3]), .B(n877), .Z(n235) );
  NANDN U286 ( .A(n19521), .B(n235), .Z(n198) );
  NAND U287 ( .A(n199), .B(n198), .Z(n234) );
  XNOR U288 ( .A(n101), .B(b[6]), .Z(n19766) );
  NAND U289 ( .A(a[0]), .B(n19766), .Z(n232) );
  NAND U290 ( .A(b[0]), .B(a[6]), .Z(n200) );
  XNOR U291 ( .A(b[1]), .B(n200), .Z(n202) );
  NAND U292 ( .A(a[5]), .B(n98), .Z(n201) );
  AND U293 ( .A(n202), .B(n201), .Z(n231) );
  XOR U294 ( .A(n232), .B(n231), .Z(n233) );
  XOR U295 ( .A(n234), .B(n233), .Z(n225) );
  XOR U296 ( .A(b[5]), .B(b[4]), .Z(n204) );
  XNOR U297 ( .A(b[5]), .B(b[3]), .Z(n203) );
  ANDN U298 ( .B(n204), .A(n203), .Z(n19722) );
  NANDN U299 ( .A(n205), .B(n19722), .Z(n207) );
  XOR U300 ( .A(b[5]), .B(a[2]), .Z(n238) );
  NANDN U301 ( .A(n19640), .B(n238), .Z(n206) );
  NAND U302 ( .A(n207), .B(n206), .Z(n226) );
  XNOR U303 ( .A(n225), .B(n226), .Z(n227) );
  XOR U304 ( .A(n228), .B(n227), .Z(n219) );
  NANDN U305 ( .A(n209), .B(n208), .Z(n213) );
  NANDN U306 ( .A(n211), .B(n210), .Z(n212) );
  NAND U307 ( .A(n213), .B(n212), .Z(n220) );
  XNOR U308 ( .A(n219), .B(n220), .Z(n221) );
  XNOR U309 ( .A(n222), .B(n221), .Z(n253) );
  NAND U310 ( .A(sreg[245]), .B(n214), .Z(n218) );
  OR U311 ( .A(n216), .B(n215), .Z(n217) );
  NAND U312 ( .A(n218), .B(n217), .Z(n251) );
  XNOR U313 ( .A(n251), .B(sreg[246]), .Z(n252) );
  XOR U314 ( .A(n253), .B(n252), .Z(c[246]) );
  NANDN U315 ( .A(n220), .B(n219), .Z(n224) );
  NAND U316 ( .A(n222), .B(n221), .Z(n223) );
  NAND U317 ( .A(n224), .B(n223), .Z(n264) );
  NANDN U318 ( .A(n226), .B(n225), .Z(n230) );
  NANDN U319 ( .A(n228), .B(n227), .Z(n229) );
  NAND U320 ( .A(n230), .B(n229), .Z(n262) );
  IV U321 ( .A(a[5]), .Z(n966) );
  XNOR U322 ( .A(n100), .B(n966), .Z(n280) );
  OR U323 ( .A(n280), .B(n19521), .Z(n237) );
  NAND U324 ( .A(n19554), .B(n235), .Z(n236) );
  AND U325 ( .A(n237), .B(n236), .Z(n267) );
  XNOR U326 ( .A(n268), .B(n267), .Z(n269) );
  NAND U327 ( .A(n238), .B(n19722), .Z(n240) );
  XNOR U328 ( .A(n101), .B(n795), .Z(n288) );
  OR U329 ( .A(n288), .B(n19640), .Z(n239) );
  NAND U330 ( .A(n240), .B(n239), .Z(n283) );
  XOR U331 ( .A(b[7]), .B(a[0]), .Z(n243) );
  XOR U332 ( .A(b[7]), .B(b[5]), .Z(n242) );
  XOR U333 ( .A(b[7]), .B(b[6]), .Z(n241) );
  AND U334 ( .A(n242), .B(n241), .Z(n19767) );
  NAND U335 ( .A(n243), .B(n19767), .Z(n245) );
  XOR U336 ( .A(b[7]), .B(a[1]), .Z(n277) );
  NAND U337 ( .A(n277), .B(n19766), .Z(n244) );
  NAND U338 ( .A(n245), .B(n244), .Z(n284) );
  XNOR U339 ( .A(n283), .B(n284), .Z(n276) );
  OR U340 ( .A(b[6]), .B(b[5]), .Z(n246) );
  NAND U341 ( .A(a[0]), .B(n246), .Z(n247) );
  NAND U342 ( .A(b[5]), .B(b[6]), .Z(n19829) );
  IV U343 ( .A(b[7]), .Z(n19714) );
  ANDN U344 ( .B(n19829), .A(n19714), .Z(n19926) );
  AND U345 ( .A(n247), .B(n19926), .Z(n273) );
  NAND U346 ( .A(b[0]), .B(a[7]), .Z(n248) );
  XNOR U347 ( .A(b[1]), .B(n248), .Z(n250) );
  NAND U348 ( .A(a[6]), .B(n98), .Z(n249) );
  AND U349 ( .A(n250), .B(n249), .Z(n274) );
  XOR U350 ( .A(n273), .B(n274), .Z(n275) );
  XOR U351 ( .A(n276), .B(n275), .Z(n270) );
  XOR U352 ( .A(n269), .B(n270), .Z(n261) );
  XNOR U353 ( .A(n262), .B(n261), .Z(n263) );
  XNOR U354 ( .A(n264), .B(n263), .Z(n256) );
  XNOR U355 ( .A(n256), .B(sreg[247]), .Z(n258) );
  NAND U356 ( .A(n251), .B(sreg[246]), .Z(n255) );
  OR U357 ( .A(n253), .B(n252), .Z(n254) );
  AND U358 ( .A(n255), .B(n254), .Z(n257) );
  XOR U359 ( .A(n258), .B(n257), .Z(c[247]) );
  NAND U360 ( .A(n256), .B(sreg[247]), .Z(n260) );
  OR U361 ( .A(n258), .B(n257), .Z(n259) );
  NAND U362 ( .A(n260), .B(n259), .Z(n335) );
  XNOR U363 ( .A(n335), .B(sreg[248]), .Z(n337) );
  NAND U364 ( .A(n262), .B(n261), .Z(n266) );
  OR U365 ( .A(n264), .B(n263), .Z(n265) );
  NAND U366 ( .A(n266), .B(n265), .Z(n294) );
  NANDN U367 ( .A(n268), .B(n267), .Z(n272) );
  NAND U368 ( .A(n270), .B(n269), .Z(n271) );
  NAND U369 ( .A(n272), .B(n271), .Z(n291) );
  IV U370 ( .A(a[2]), .Z(n744) );
  XNOR U371 ( .A(n19714), .B(n744), .Z(n309) );
  NANDN U372 ( .A(n309), .B(n19766), .Z(n279) );
  NAND U373 ( .A(n277), .B(n19767), .Z(n278) );
  NAND U374 ( .A(n279), .B(n278), .Z(n297) );
  NANDN U375 ( .A(n280), .B(n19554), .Z(n282) );
  IV U376 ( .A(a[6]), .Z(n1042) );
  XNOR U377 ( .A(b[3]), .B(n1042), .Z(n306) );
  NANDN U378 ( .A(n19521), .B(n306), .Z(n281) );
  AND U379 ( .A(n282), .B(n281), .Z(n298) );
  XNOR U380 ( .A(n297), .B(n298), .Z(n299) );
  NAND U381 ( .A(n284), .B(n283), .Z(n300) );
  XOR U382 ( .A(n299), .B(n300), .Z(n329) );
  XOR U383 ( .A(b[7]), .B(b[8]), .Z(n19883) );
  NANDN U384 ( .A(n685), .B(n19883), .Z(n326) );
  NAND U385 ( .A(b[0]), .B(a[8]), .Z(n285) );
  XNOR U386 ( .A(b[1]), .B(n285), .Z(n287) );
  NAND U387 ( .A(a[7]), .B(n98), .Z(n286) );
  AND U388 ( .A(n287), .B(n286), .Z(n324) );
  NANDN U389 ( .A(n288), .B(n19722), .Z(n290) );
  XOR U390 ( .A(b[5]), .B(a[4]), .Z(n320) );
  NANDN U391 ( .A(n19640), .B(n320), .Z(n289) );
  AND U392 ( .A(n290), .B(n289), .Z(n323) );
  XNOR U393 ( .A(n324), .B(n323), .Z(n325) );
  XNOR U394 ( .A(n326), .B(n325), .Z(n330) );
  XNOR U395 ( .A(n329), .B(n330), .Z(n331) );
  XNOR U396 ( .A(n332), .B(n331), .Z(n292) );
  XNOR U397 ( .A(n291), .B(n292), .Z(n293) );
  XOR U398 ( .A(n294), .B(n293), .Z(n336) );
  XOR U399 ( .A(n337), .B(n336), .Z(c[248]) );
  NANDN U400 ( .A(n292), .B(n291), .Z(n296) );
  NAND U401 ( .A(n294), .B(n293), .Z(n295) );
  NAND U402 ( .A(n296), .B(n295), .Z(n348) );
  NANDN U403 ( .A(n298), .B(n297), .Z(n302) );
  NANDN U404 ( .A(n300), .B(n299), .Z(n301) );
  NAND U405 ( .A(n302), .B(n301), .Z(n352) );
  NAND U406 ( .A(b[0]), .B(a[9]), .Z(n303) );
  XNOR U407 ( .A(b[1]), .B(n303), .Z(n305) );
  NAND U408 ( .A(a[8]), .B(n98), .Z(n304) );
  AND U409 ( .A(n305), .B(n304), .Z(n362) );
  XNOR U410 ( .A(b[3]), .B(a[7]), .Z(n375) );
  OR U411 ( .A(n375), .B(n19521), .Z(n308) );
  NAND U412 ( .A(n19554), .B(n306), .Z(n307) );
  AND U413 ( .A(n308), .B(n307), .Z(n361) );
  XNOR U414 ( .A(n362), .B(n361), .Z(n363) );
  XNOR U415 ( .A(n19714), .B(n795), .Z(n381) );
  NANDN U416 ( .A(n381), .B(n19766), .Z(n311) );
  NANDN U417 ( .A(n309), .B(n19767), .Z(n310) );
  NAND U418 ( .A(n311), .B(n310), .Z(n367) );
  XOR U419 ( .A(b[9]), .B(a[0]), .Z(n314) );
  XOR U420 ( .A(b[9]), .B(b[7]), .Z(n313) );
  XOR U421 ( .A(b[9]), .B(b[8]), .Z(n312) );
  AND U422 ( .A(n313), .B(n312), .Z(n19937) );
  NAND U423 ( .A(n314), .B(n19937), .Z(n316) );
  XOR U424 ( .A(b[9]), .B(a[1]), .Z(n369) );
  AND U425 ( .A(n369), .B(n19883), .Z(n315) );
  ANDN U426 ( .B(n316), .A(n315), .Z(n368) );
  XNOR U427 ( .A(n367), .B(n368), .Z(n358) );
  ANDN U428 ( .B(n19714), .A(b[8]), .Z(n317) );
  NAND U429 ( .A(b[9]), .B(n317), .Z(n319) );
  AND U430 ( .A(n19883), .B(b[9]), .Z(n19939) );
  NAND U431 ( .A(n685), .B(n19939), .Z(n318) );
  NAND U432 ( .A(n319), .B(n318), .Z(n356) );
  NAND U433 ( .A(n320), .B(n19722), .Z(n322) );
  XNOR U434 ( .A(n101), .B(n966), .Z(n372) );
  OR U435 ( .A(n372), .B(n19640), .Z(n321) );
  NAND U436 ( .A(n322), .B(n321), .Z(n355) );
  XOR U437 ( .A(n356), .B(n355), .Z(n357) );
  XOR U438 ( .A(n358), .B(n357), .Z(n364) );
  XOR U439 ( .A(n363), .B(n364), .Z(n349) );
  NANDN U440 ( .A(n324), .B(n323), .Z(n328) );
  NAND U441 ( .A(n326), .B(n325), .Z(n327) );
  NAND U442 ( .A(n328), .B(n327), .Z(n350) );
  XNOR U443 ( .A(n349), .B(n350), .Z(n351) );
  XNOR U444 ( .A(n352), .B(n351), .Z(n345) );
  NANDN U445 ( .A(n330), .B(n329), .Z(n334) );
  NAND U446 ( .A(n332), .B(n331), .Z(n333) );
  AND U447 ( .A(n334), .B(n333), .Z(n346) );
  XOR U448 ( .A(n345), .B(n346), .Z(n347) );
  XOR U449 ( .A(n348), .B(n347), .Z(n340) );
  XNOR U450 ( .A(n340), .B(sreg[249]), .Z(n342) );
  NAND U451 ( .A(n335), .B(sreg[248]), .Z(n339) );
  OR U452 ( .A(n337), .B(n336), .Z(n338) );
  AND U453 ( .A(n339), .B(n338), .Z(n341) );
  XOR U454 ( .A(n342), .B(n341), .Z(c[249]) );
  NAND U455 ( .A(n340), .B(sreg[249]), .Z(n344) );
  OR U456 ( .A(n342), .B(n341), .Z(n343) );
  NAND U457 ( .A(n344), .B(n343), .Z(n438) );
  XNOR U458 ( .A(n438), .B(sreg[250]), .Z(n440) );
  NANDN U459 ( .A(n350), .B(n349), .Z(n354) );
  NAND U460 ( .A(n352), .B(n351), .Z(n353) );
  NAND U461 ( .A(n354), .B(n353), .Z(n385) );
  OR U462 ( .A(n356), .B(n355), .Z(n360) );
  NANDN U463 ( .A(n358), .B(n357), .Z(n359) );
  NAND U464 ( .A(n360), .B(n359), .Z(n392) );
  NANDN U465 ( .A(n362), .B(n361), .Z(n366) );
  NANDN U466 ( .A(n364), .B(n363), .Z(n365) );
  NAND U467 ( .A(n366), .B(n365), .Z(n391) );
  NANDN U468 ( .A(n368), .B(n367), .Z(n411) );
  NAND U469 ( .A(n19937), .B(n369), .Z(n371) );
  XOR U470 ( .A(b[9]), .B(a[2]), .Z(n424) );
  NAND U471 ( .A(n19883), .B(n424), .Z(n370) );
  NAND U472 ( .A(n371), .B(n370), .Z(n409) );
  NANDN U473 ( .A(n372), .B(n19722), .Z(n374) );
  XNOR U474 ( .A(n101), .B(n1042), .Z(n435) );
  OR U475 ( .A(n435), .B(n19640), .Z(n373) );
  AND U476 ( .A(n374), .B(n373), .Z(n408) );
  XNOR U477 ( .A(n409), .B(n408), .Z(n410) );
  XNOR U478 ( .A(n411), .B(n410), .Z(n397) );
  IV U479 ( .A(a[8]), .Z(n1171) );
  XNOR U480 ( .A(n100), .B(n1171), .Z(n421) );
  OR U481 ( .A(n421), .B(n19521), .Z(n377) );
  NANDN U482 ( .A(n375), .B(n19554), .Z(n376) );
  AND U483 ( .A(n377), .B(n376), .Z(n396) );
  XNOR U484 ( .A(n397), .B(n396), .Z(n398) );
  XNOR U485 ( .A(b[9]), .B(b[10]), .Z(n20020) );
  ANDN U486 ( .B(a[0]), .A(n20020), .Z(n405) );
  NAND U487 ( .A(b[0]), .B(a[10]), .Z(n378) );
  XNOR U488 ( .A(b[1]), .B(n378), .Z(n380) );
  NAND U489 ( .A(a[9]), .B(n98), .Z(n379) );
  AND U490 ( .A(n380), .B(n379), .Z(n403) );
  NANDN U491 ( .A(n381), .B(n19767), .Z(n383) );
  XNOR U492 ( .A(b[7]), .B(a[4]), .Z(n414) );
  NANDN U493 ( .A(n414), .B(n19766), .Z(n382) );
  AND U494 ( .A(n383), .B(n382), .Z(n402) );
  XNOR U495 ( .A(n403), .B(n402), .Z(n404) );
  XOR U496 ( .A(n405), .B(n404), .Z(n399) );
  XNOR U497 ( .A(n398), .B(n399), .Z(n390) );
  XNOR U498 ( .A(n391), .B(n390), .Z(n393) );
  XNOR U499 ( .A(n392), .B(n393), .Z(n384) );
  XNOR U500 ( .A(n385), .B(n384), .Z(n386) );
  XOR U501 ( .A(n387), .B(n386), .Z(n439) );
  XOR U502 ( .A(n440), .B(n439), .Z(c[250]) );
  NANDN U503 ( .A(n385), .B(n384), .Z(n389) );
  NAND U504 ( .A(n387), .B(n386), .Z(n388) );
  NAND U505 ( .A(n389), .B(n388), .Z(n451) );
  NAND U506 ( .A(n391), .B(n390), .Z(n395) );
  NANDN U507 ( .A(n393), .B(n392), .Z(n394) );
  NAND U508 ( .A(n395), .B(n394), .Z(n449) );
  NANDN U509 ( .A(n397), .B(n396), .Z(n401) );
  NANDN U510 ( .A(n399), .B(n398), .Z(n400) );
  NAND U511 ( .A(n401), .B(n400), .Z(n456) );
  NANDN U512 ( .A(n403), .B(n402), .Z(n407) );
  NANDN U513 ( .A(n405), .B(n404), .Z(n406) );
  NAND U514 ( .A(n407), .B(n406), .Z(n455) );
  NANDN U515 ( .A(n409), .B(n408), .Z(n413) );
  NAND U516 ( .A(n411), .B(n410), .Z(n412) );
  NAND U517 ( .A(n413), .B(n412), .Z(n493) );
  NANDN U518 ( .A(n414), .B(n19767), .Z(n416) );
  XNOR U519 ( .A(b[7]), .B(a[5]), .Z(n474) );
  NANDN U520 ( .A(n474), .B(n19766), .Z(n415) );
  NAND U521 ( .A(n416), .B(n415), .Z(n463) );
  NAND U522 ( .A(a[0]), .B(b[9]), .Z(n417) );
  AND U523 ( .A(n417), .B(b[11]), .Z(n420) );
  IV U524 ( .A(b[9]), .Z(n19975) );
  AND U525 ( .A(n685), .B(n19975), .Z(n418) );
  NANDN U526 ( .A(n418), .B(b[10]), .Z(n419) );
  AND U527 ( .A(n420), .B(n419), .Z(n460) );
  NANDN U528 ( .A(n421), .B(n19554), .Z(n423) );
  IV U529 ( .A(a[9]), .Z(n1276) );
  XNOR U530 ( .A(b[3]), .B(n1276), .Z(n477) );
  NANDN U531 ( .A(n19521), .B(n477), .Z(n422) );
  NAND U532 ( .A(n423), .B(n422), .Z(n461) );
  XNOR U533 ( .A(n460), .B(n461), .Z(n462) );
  XOR U534 ( .A(n463), .B(n462), .Z(n492) );
  XNOR U535 ( .A(n493), .B(n492), .Z(n495) );
  XNOR U536 ( .A(n19975), .B(n795), .Z(n483) );
  NANDN U537 ( .A(n483), .B(n19883), .Z(n426) );
  NAND U538 ( .A(n424), .B(n19937), .Z(n425) );
  NAND U539 ( .A(n426), .B(n425), .Z(n473) );
  XOR U540 ( .A(b[11]), .B(a[0]), .Z(n429) );
  XOR U541 ( .A(b[11]), .B(b[9]), .Z(n428) );
  XOR U542 ( .A(b[11]), .B(b[10]), .Z(n427) );
  AND U543 ( .A(n428), .B(n427), .Z(n19960) );
  NAND U544 ( .A(n429), .B(n19960), .Z(n431) );
  IV U545 ( .A(b[11]), .Z(n20052) );
  XOR U546 ( .A(n20052), .B(a[1]), .Z(n469) );
  OR U547 ( .A(n469), .B(n20020), .Z(n430) );
  NAND U548 ( .A(n431), .B(n430), .Z(n472) );
  XNOR U549 ( .A(n473), .B(n472), .Z(n489) );
  NAND U550 ( .A(b[0]), .B(a[11]), .Z(n432) );
  XNOR U551 ( .A(b[1]), .B(n432), .Z(n434) );
  NAND U552 ( .A(a[10]), .B(n98), .Z(n433) );
  AND U553 ( .A(n434), .B(n433), .Z(n487) );
  NANDN U554 ( .A(n435), .B(n19722), .Z(n437) );
  IV U555 ( .A(a[7]), .Z(n1093) );
  XNOR U556 ( .A(b[5]), .B(n1093), .Z(n466) );
  NANDN U557 ( .A(n19640), .B(n466), .Z(n436) );
  AND U558 ( .A(n437), .B(n436), .Z(n486) );
  XNOR U559 ( .A(n487), .B(n486), .Z(n488) );
  XOR U560 ( .A(n489), .B(n488), .Z(n494) );
  XNOR U561 ( .A(n495), .B(n494), .Z(n454) );
  XNOR U562 ( .A(n455), .B(n454), .Z(n457) );
  XNOR U563 ( .A(n456), .B(n457), .Z(n448) );
  XOR U564 ( .A(n449), .B(n448), .Z(n450) );
  XNOR U565 ( .A(n451), .B(n450), .Z(n443) );
  XNOR U566 ( .A(n443), .B(sreg[251]), .Z(n445) );
  NAND U567 ( .A(n438), .B(sreg[250]), .Z(n442) );
  OR U568 ( .A(n440), .B(n439), .Z(n441) );
  AND U569 ( .A(n442), .B(n441), .Z(n444) );
  XOR U570 ( .A(n445), .B(n444), .Z(c[251]) );
  NAND U571 ( .A(n443), .B(sreg[251]), .Z(n447) );
  OR U572 ( .A(n445), .B(n444), .Z(n446) );
  NAND U573 ( .A(n447), .B(n446), .Z(n558) );
  XNOR U574 ( .A(n558), .B(sreg[252]), .Z(n560) );
  NAND U575 ( .A(n449), .B(n448), .Z(n453) );
  NAND U576 ( .A(n451), .B(n450), .Z(n452) );
  NAND U577 ( .A(n453), .B(n452), .Z(n501) );
  NAND U578 ( .A(n455), .B(n454), .Z(n459) );
  NANDN U579 ( .A(n457), .B(n456), .Z(n458) );
  NAND U580 ( .A(n459), .B(n458), .Z(n498) );
  OR U581 ( .A(n461), .B(n460), .Z(n465) );
  OR U582 ( .A(n463), .B(n462), .Z(n464) );
  NAND U583 ( .A(n465), .B(n464), .Z(n507) );
  NAND U584 ( .A(n19722), .B(n466), .Z(n468) );
  XNOR U585 ( .A(n101), .B(n1171), .Z(n541) );
  OR U586 ( .A(n541), .B(n19640), .Z(n467) );
  NAND U587 ( .A(n468), .B(n467), .Z(n511) );
  XNOR U588 ( .A(n20052), .B(n744), .Z(n544) );
  OR U589 ( .A(n544), .B(n20020), .Z(n471) );
  NANDN U590 ( .A(n469), .B(n19960), .Z(n470) );
  NAND U591 ( .A(n471), .B(n470), .Z(n510) );
  XOR U592 ( .A(n511), .B(n510), .Z(n512) );
  NAND U593 ( .A(n473), .B(n472), .Z(n523) );
  NANDN U594 ( .A(n474), .B(n19767), .Z(n476) );
  XNOR U595 ( .A(b[7]), .B(a[6]), .Z(n555) );
  NANDN U596 ( .A(n555), .B(n19766), .Z(n475) );
  NAND U597 ( .A(n476), .B(n475), .Z(n521) );
  IV U598 ( .A(a[10]), .Z(n1354) );
  XNOR U599 ( .A(n100), .B(n1354), .Z(n535) );
  OR U600 ( .A(n535), .B(n19521), .Z(n479) );
  NAND U601 ( .A(n19554), .B(n477), .Z(n478) );
  AND U602 ( .A(n479), .B(n478), .Z(n520) );
  XNOR U603 ( .A(n521), .B(n520), .Z(n522) );
  XNOR U604 ( .A(n523), .B(n522), .Z(n513) );
  XNOR U605 ( .A(n512), .B(n513), .Z(n516) );
  XNOR U606 ( .A(b[11]), .B(b[12]), .Z(n20057) );
  ANDN U607 ( .B(a[0]), .A(n20057), .Z(n529) );
  NAND U608 ( .A(b[0]), .B(a[12]), .Z(n480) );
  XNOR U609 ( .A(b[1]), .B(n480), .Z(n482) );
  NAND U610 ( .A(a[11]), .B(n98), .Z(n481) );
  AND U611 ( .A(n482), .B(n481), .Z(n527) );
  NANDN U612 ( .A(n483), .B(n19937), .Z(n485) );
  XOR U613 ( .A(b[9]), .B(a[4]), .Z(n538) );
  NAND U614 ( .A(n19883), .B(n538), .Z(n484) );
  AND U615 ( .A(n485), .B(n484), .Z(n526) );
  XNOR U616 ( .A(n527), .B(n526), .Z(n528) );
  XOR U617 ( .A(n529), .B(n528), .Z(n514) );
  NANDN U618 ( .A(n487), .B(n486), .Z(n491) );
  NAND U619 ( .A(n489), .B(n488), .Z(n490) );
  NAND U620 ( .A(n491), .B(n490), .Z(n515) );
  XOR U621 ( .A(n514), .B(n515), .Z(n517) );
  XOR U622 ( .A(n516), .B(n517), .Z(n505) );
  NAND U623 ( .A(n493), .B(n492), .Z(n497) );
  NANDN U624 ( .A(n495), .B(n494), .Z(n496) );
  AND U625 ( .A(n497), .B(n496), .Z(n504) );
  XOR U626 ( .A(n505), .B(n504), .Z(n506) );
  XNOR U627 ( .A(n507), .B(n506), .Z(n499) );
  XNOR U628 ( .A(n498), .B(n499), .Z(n500) );
  XOR U629 ( .A(n501), .B(n500), .Z(n559) );
  XOR U630 ( .A(n560), .B(n559), .Z(c[252]) );
  NANDN U631 ( .A(n499), .B(n498), .Z(n503) );
  NAND U632 ( .A(n501), .B(n500), .Z(n502) );
  NAND U633 ( .A(n503), .B(n502), .Z(n571) );
  OR U634 ( .A(n505), .B(n504), .Z(n509) );
  NAND U635 ( .A(n507), .B(n506), .Z(n508) );
  NAND U636 ( .A(n509), .B(n508), .Z(n569) );
  NANDN U637 ( .A(n515), .B(n514), .Z(n519) );
  OR U638 ( .A(n517), .B(n516), .Z(n518) );
  NAND U639 ( .A(n519), .B(n518), .Z(n575) );
  XNOR U640 ( .A(n574), .B(n575), .Z(n576) );
  NANDN U641 ( .A(n521), .B(n520), .Z(n525) );
  NAND U642 ( .A(n523), .B(n522), .Z(n524) );
  NAND U643 ( .A(n525), .B(n524), .Z(n615) );
  NANDN U644 ( .A(n527), .B(n526), .Z(n531) );
  NANDN U645 ( .A(n529), .B(n528), .Z(n530) );
  AND U646 ( .A(n531), .B(n530), .Z(n616) );
  XNOR U647 ( .A(n615), .B(n616), .Z(n617) );
  ANDN U648 ( .B(n20052), .A(b[12]), .Z(n532) );
  NAND U649 ( .A(b[13]), .B(n532), .Z(n534) );
  IV U650 ( .A(b[13]), .Z(n20154) );
  NOR U651 ( .A(n20154), .B(n20057), .Z(n20100) );
  NAND U652 ( .A(n685), .B(n20100), .Z(n533) );
  NAND U653 ( .A(n534), .B(n533), .Z(n596) );
  NANDN U654 ( .A(n535), .B(n19554), .Z(n537) );
  IV U655 ( .A(a[11]), .Z(n1432) );
  XNOR U656 ( .A(b[3]), .B(n1432), .Z(n612) );
  NANDN U657 ( .A(n19521), .B(n612), .Z(n536) );
  NAND U658 ( .A(n537), .B(n536), .Z(n594) );
  XNOR U659 ( .A(b[9]), .B(n966), .Z(n582) );
  NAND U660 ( .A(n19883), .B(n582), .Z(n540) );
  NAND U661 ( .A(n538), .B(n19937), .Z(n539) );
  AND U662 ( .A(n540), .B(n539), .Z(n595) );
  XNOR U663 ( .A(n594), .B(n595), .Z(n597) );
  XOR U664 ( .A(n596), .B(n597), .Z(n621) );
  NANDN U665 ( .A(n541), .B(n19722), .Z(n543) );
  XOR U666 ( .A(b[5]), .B(a[9]), .Z(n606) );
  NANDN U667 ( .A(n19640), .B(n606), .Z(n542) );
  NAND U668 ( .A(n543), .B(n542), .Z(n622) );
  XNOR U669 ( .A(n621), .B(n622), .Z(n624) );
  XOR U670 ( .A(b[11]), .B(a[3]), .Z(n603) );
  NANDN U671 ( .A(n20020), .B(n603), .Z(n546) );
  NANDN U672 ( .A(n544), .B(n19960), .Z(n545) );
  NAND U673 ( .A(n546), .B(n545), .Z(n581) );
  XOR U674 ( .A(b[13]), .B(a[1]), .Z(n585) );
  ANDN U675 ( .B(n585), .A(n20057), .Z(n551) );
  XOR U676 ( .A(b[13]), .B(a[0]), .Z(n549) );
  XOR U677 ( .A(b[13]), .B(b[11]), .Z(n548) );
  XOR U678 ( .A(b[13]), .B(b[12]), .Z(n547) );
  AND U679 ( .A(n548), .B(n547), .Z(n20098) );
  NAND U680 ( .A(n549), .B(n20098), .Z(n550) );
  NANDN U681 ( .A(n551), .B(n550), .Z(n580) );
  XNOR U682 ( .A(n581), .B(n580), .Z(n591) );
  NAND U683 ( .A(b[0]), .B(a[13]), .Z(n552) );
  XNOR U684 ( .A(b[1]), .B(n552), .Z(n554) );
  NAND U685 ( .A(a[12]), .B(n98), .Z(n553) );
  AND U686 ( .A(n554), .B(n553), .Z(n589) );
  NANDN U687 ( .A(n555), .B(n19767), .Z(n557) );
  XNOR U688 ( .A(n19714), .B(n1093), .Z(n609) );
  NANDN U689 ( .A(n609), .B(n19766), .Z(n556) );
  AND U690 ( .A(n557), .B(n556), .Z(n588) );
  XNOR U691 ( .A(n589), .B(n588), .Z(n590) );
  XOR U692 ( .A(n591), .B(n590), .Z(n623) );
  XOR U693 ( .A(n617), .B(n618), .Z(n577) );
  XOR U694 ( .A(n576), .B(n577), .Z(n568) );
  XOR U695 ( .A(n569), .B(n568), .Z(n570) );
  XNOR U696 ( .A(n571), .B(n570), .Z(n563) );
  XNOR U697 ( .A(n563), .B(sreg[253]), .Z(n565) );
  NAND U698 ( .A(n558), .B(sreg[252]), .Z(n562) );
  OR U699 ( .A(n560), .B(n559), .Z(n561) );
  AND U700 ( .A(n562), .B(n561), .Z(n564) );
  XOR U701 ( .A(n565), .B(n564), .Z(c[253]) );
  NAND U702 ( .A(n563), .B(sreg[253]), .Z(n567) );
  OR U703 ( .A(n565), .B(n564), .Z(n566) );
  NAND U704 ( .A(n567), .B(n566), .Z(n699) );
  XNOR U705 ( .A(n699), .B(sreg[254]), .Z(n701) );
  NAND U706 ( .A(n569), .B(n568), .Z(n573) );
  NAND U707 ( .A(n571), .B(n570), .Z(n572) );
  NAND U708 ( .A(n573), .B(n572), .Z(n630) );
  NANDN U709 ( .A(n575), .B(n574), .Z(n579) );
  NAND U710 ( .A(n577), .B(n576), .Z(n578) );
  NAND U711 ( .A(n579), .B(n578), .Z(n627) );
  AND U712 ( .A(n581), .B(n580), .Z(n641) );
  NAND U713 ( .A(n19937), .B(n582), .Z(n584) );
  XNOR U714 ( .A(b[9]), .B(n1042), .Z(n673) );
  NAND U715 ( .A(n19883), .B(n673), .Z(n583) );
  NAND U716 ( .A(n584), .B(n583), .Z(n640) );
  NAND U717 ( .A(n20098), .B(n585), .Z(n587) );
  XOR U718 ( .A(b[13]), .B(a[2]), .Z(n661) );
  NANDN U719 ( .A(n20057), .B(n661), .Z(n586) );
  AND U720 ( .A(n587), .B(n586), .Z(n639) );
  XNOR U721 ( .A(n640), .B(n639), .Z(n642) );
  XOR U722 ( .A(n641), .B(n642), .Z(n693) );
  NANDN U723 ( .A(n589), .B(n588), .Z(n593) );
  NAND U724 ( .A(n591), .B(n590), .Z(n592) );
  NAND U725 ( .A(n593), .B(n592), .Z(n694) );
  XOR U726 ( .A(n693), .B(n694), .Z(n696) );
  NANDN U727 ( .A(n595), .B(n594), .Z(n599) );
  NAND U728 ( .A(n597), .B(n596), .Z(n598) );
  NAND U729 ( .A(n599), .B(n598), .Z(n652) );
  XOR U730 ( .A(n20154), .B(b[14]), .Z(n20121) );
  ANDN U731 ( .B(a[0]), .A(n20121), .Z(n646) );
  NAND U732 ( .A(b[0]), .B(a[14]), .Z(n600) );
  XNOR U733 ( .A(b[1]), .B(n600), .Z(n602) );
  NAND U734 ( .A(a[13]), .B(n98), .Z(n601) );
  AND U735 ( .A(n602), .B(n601), .Z(n644) );
  NAND U736 ( .A(n603), .B(n19960), .Z(n605) );
  XNOR U737 ( .A(n20052), .B(n877), .Z(n676) );
  OR U738 ( .A(n676), .B(n20020), .Z(n604) );
  AND U739 ( .A(n605), .B(n604), .Z(n643) );
  XNOR U740 ( .A(n644), .B(n643), .Z(n645) );
  XOR U741 ( .A(n646), .B(n645), .Z(n649) );
  NAND U742 ( .A(n606), .B(n19722), .Z(n608) );
  XNOR U743 ( .A(n101), .B(n1354), .Z(n679) );
  OR U744 ( .A(n679), .B(n19640), .Z(n607) );
  NAND U745 ( .A(n608), .B(n607), .Z(n658) );
  XNOR U746 ( .A(b[7]), .B(n1171), .Z(n690) );
  NAND U747 ( .A(n690), .B(n19766), .Z(n611) );
  NANDN U748 ( .A(n609), .B(n19767), .Z(n610) );
  NAND U749 ( .A(n611), .B(n610), .Z(n655) );
  NAND U750 ( .A(n19554), .B(n612), .Z(n614) );
  IV U751 ( .A(a[12]), .Z(n1495) );
  XNOR U752 ( .A(b[3]), .B(n1495), .Z(n682) );
  NANDN U753 ( .A(n19521), .B(n682), .Z(n613) );
  AND U754 ( .A(n614), .B(n613), .Z(n656) );
  XNOR U755 ( .A(n655), .B(n656), .Z(n657) );
  XNOR U756 ( .A(n658), .B(n657), .Z(n650) );
  XNOR U757 ( .A(n649), .B(n650), .Z(n651) );
  XNOR U758 ( .A(n652), .B(n651), .Z(n695) );
  XNOR U759 ( .A(n696), .B(n695), .Z(n636) );
  NANDN U760 ( .A(n616), .B(n615), .Z(n620) );
  NAND U761 ( .A(n618), .B(n617), .Z(n619) );
  NAND U762 ( .A(n620), .B(n619), .Z(n633) );
  OR U763 ( .A(n622), .B(n621), .Z(n626) );
  NANDN U764 ( .A(n624), .B(n623), .Z(n625) );
  AND U765 ( .A(n626), .B(n625), .Z(n634) );
  XNOR U766 ( .A(n633), .B(n634), .Z(n635) );
  XNOR U767 ( .A(n636), .B(n635), .Z(n628) );
  XNOR U768 ( .A(n627), .B(n628), .Z(n629) );
  XOR U769 ( .A(n630), .B(n629), .Z(n700) );
  XOR U770 ( .A(n701), .B(n700), .Z(c[254]) );
  NANDN U771 ( .A(n628), .B(n627), .Z(n632) );
  NAND U772 ( .A(n630), .B(n629), .Z(n631) );
  NAND U773 ( .A(n632), .B(n631), .Z(n712) );
  NANDN U774 ( .A(n634), .B(n633), .Z(n638) );
  NAND U775 ( .A(n636), .B(n635), .Z(n637) );
  NAND U776 ( .A(n638), .B(n637), .Z(n710) );
  NANDN U777 ( .A(n644), .B(n643), .Z(n648) );
  NANDN U778 ( .A(n646), .B(n645), .Z(n647) );
  AND U779 ( .A(n648), .B(n647), .Z(n720) );
  XNOR U780 ( .A(n719), .B(n720), .Z(n721) );
  NANDN U781 ( .A(n650), .B(n649), .Z(n654) );
  NAND U782 ( .A(n652), .B(n651), .Z(n653) );
  AND U783 ( .A(n654), .B(n653), .Z(n722) );
  XNOR U784 ( .A(n721), .B(n722), .Z(n716) );
  NANDN U785 ( .A(n656), .B(n655), .Z(n660) );
  NAND U786 ( .A(n658), .B(n657), .Z(n659) );
  NAND U787 ( .A(n660), .B(n659), .Z(n771) );
  XNOR U788 ( .A(n20154), .B(n795), .Z(n735) );
  OR U789 ( .A(n735), .B(n20057), .Z(n663) );
  NAND U790 ( .A(n661), .B(n20098), .Z(n662) );
  NAND U791 ( .A(n663), .B(n662), .Z(n757) );
  XNOR U792 ( .A(b[13]), .B(n102), .Z(n665) );
  XNOR U793 ( .A(a[0]), .B(b[14]), .Z(n664) );
  AND U794 ( .A(n665), .B(n664), .Z(n667) );
  XNOR U795 ( .A(b[13]), .B(a[0]), .Z(n666) );
  NAND U796 ( .A(n667), .B(n666), .Z(n669) );
  XOR U797 ( .A(b[15]), .B(a[1]), .Z(n747) );
  NANDN U798 ( .A(n20121), .B(n747), .Z(n668) );
  NAND U799 ( .A(n669), .B(n668), .Z(n756) );
  XNOR U800 ( .A(n757), .B(n756), .Z(n732) );
  AND U801 ( .A(a[15]), .B(b[0]), .Z(n670) );
  XOR U802 ( .A(b[1]), .B(n670), .Z(n672) );
  NAND U803 ( .A(a[14]), .B(n98), .Z(n671) );
  NAND U804 ( .A(n672), .B(n671), .Z(n729) );
  NAND U805 ( .A(n19937), .B(n673), .Z(n675) );
  XNOR U806 ( .A(b[9]), .B(n1093), .Z(n761) );
  NAND U807 ( .A(n19883), .B(n761), .Z(n674) );
  NAND U808 ( .A(n675), .B(n674), .Z(n730) );
  XNOR U809 ( .A(n729), .B(n730), .Z(n731) );
  XOR U810 ( .A(n732), .B(n731), .Z(n770) );
  XOR U811 ( .A(n771), .B(n770), .Z(n772) );
  NANDN U812 ( .A(n676), .B(n19960), .Z(n678) );
  XOR U813 ( .A(b[11]), .B(a[5]), .Z(n741) );
  NANDN U814 ( .A(n20020), .B(n741), .Z(n677) );
  NAND U815 ( .A(n678), .B(n677), .Z(n727) );
  NANDN U816 ( .A(n679), .B(n19722), .Z(n681) );
  XOR U817 ( .A(b[5]), .B(a[11]), .Z(n750) );
  NANDN U818 ( .A(n19640), .B(n750), .Z(n680) );
  AND U819 ( .A(n681), .B(n680), .Z(n725) );
  XNOR U820 ( .A(b[3]), .B(a[13]), .Z(n758) );
  OR U821 ( .A(n758), .B(n19521), .Z(n684) );
  NAND U822 ( .A(n19554), .B(n682), .Z(n683) );
  NAND U823 ( .A(n684), .B(n683), .Z(n726) );
  XOR U824 ( .A(n725), .B(n726), .Z(n728) );
  XOR U825 ( .A(n727), .B(n728), .Z(n767) );
  NAND U826 ( .A(n685), .B(n20154), .Z(n686) );
  NAND U827 ( .A(b[14]), .B(n686), .Z(n688) );
  AND U828 ( .A(a[0]), .B(b[13]), .Z(n687) );
  ANDN U829 ( .B(n688), .A(n687), .Z(n689) );
  ANDN U830 ( .B(n689), .A(n102), .Z(n764) );
  NAND U831 ( .A(n19767), .B(n690), .Z(n692) );
  XNOR U832 ( .A(b[7]), .B(a[9]), .Z(n753) );
  NANDN U833 ( .A(n753), .B(n19766), .Z(n691) );
  NAND U834 ( .A(n692), .B(n691), .Z(n765) );
  XOR U835 ( .A(n764), .B(n765), .Z(n766) );
  XOR U836 ( .A(n767), .B(n766), .Z(n773) );
  XNOR U837 ( .A(n772), .B(n773), .Z(n713) );
  NANDN U838 ( .A(n694), .B(n693), .Z(n698) );
  OR U839 ( .A(n696), .B(n695), .Z(n697) );
  AND U840 ( .A(n698), .B(n697), .Z(n714) );
  XOR U841 ( .A(n713), .B(n714), .Z(n715) );
  XOR U842 ( .A(n716), .B(n715), .Z(n709) );
  XOR U843 ( .A(n710), .B(n709), .Z(n711) );
  XOR U844 ( .A(n712), .B(n711), .Z(n704) );
  XNOR U845 ( .A(n704), .B(sreg[255]), .Z(n706) );
  NAND U846 ( .A(n699), .B(sreg[254]), .Z(n703) );
  OR U847 ( .A(n701), .B(n700), .Z(n702) );
  AND U848 ( .A(n703), .B(n702), .Z(n705) );
  XOR U849 ( .A(n706), .B(n705), .Z(c[255]) );
  NAND U850 ( .A(n704), .B(sreg[255]), .Z(n708) );
  OR U851 ( .A(n706), .B(n705), .Z(n707) );
  NAND U852 ( .A(n708), .B(n707), .Z(n845) );
  XNOR U853 ( .A(n845), .B(sreg[256]), .Z(n847) );
  NAND U854 ( .A(n714), .B(n713), .Z(n718) );
  NANDN U855 ( .A(n716), .B(n715), .Z(n717) );
  NAND U856 ( .A(n718), .B(n717), .Z(n774) );
  NANDN U857 ( .A(n720), .B(n719), .Z(n724) );
  NAND U858 ( .A(n722), .B(n721), .Z(n723) );
  NAND U859 ( .A(n724), .B(n723), .Z(n783) );
  NANDN U860 ( .A(n730), .B(n729), .Z(n734) );
  NAND U861 ( .A(n732), .B(n731), .Z(n733) );
  AND U862 ( .A(n734), .B(n733), .Z(n835) );
  XNOR U863 ( .A(n20154), .B(n877), .Z(n817) );
  OR U864 ( .A(n817), .B(n20057), .Z(n737) );
  NANDN U865 ( .A(n735), .B(n20098), .Z(n736) );
  NAND U866 ( .A(n737), .B(n736), .Z(n826) );
  NAND U867 ( .A(b[0]), .B(a[16]), .Z(n738) );
  XNOR U868 ( .A(b[1]), .B(n738), .Z(n740) );
  NAND U869 ( .A(a[15]), .B(n98), .Z(n739) );
  AND U870 ( .A(n740), .B(n739), .Z(n823) );
  NAND U871 ( .A(b[15]), .B(a[0]), .Z(n824) );
  XNOR U872 ( .A(n823), .B(n824), .Z(n825) );
  XOR U873 ( .A(n826), .B(n825), .Z(n836) );
  XOR U874 ( .A(n835), .B(n836), .Z(n837) );
  XNOR U875 ( .A(n838), .B(n837), .Z(n842) );
  XNOR U876 ( .A(n20052), .B(n1042), .Z(n792) );
  OR U877 ( .A(n792), .B(n20020), .Z(n743) );
  NAND U878 ( .A(n741), .B(n19960), .Z(n742) );
  NAND U879 ( .A(n743), .B(n742), .Z(n805) );
  XNOR U880 ( .A(n102), .B(n744), .Z(n796) );
  OR U881 ( .A(n796), .B(n20121), .Z(n749) );
  XOR U882 ( .A(b[15]), .B(b[13]), .Z(n746) );
  XOR U883 ( .A(b[15]), .B(b[14]), .Z(n745) );
  AND U884 ( .A(n746), .B(n745), .Z(n20122) );
  NAND U885 ( .A(n747), .B(n20122), .Z(n748) );
  NAND U886 ( .A(n749), .B(n748), .Z(n802) );
  NAND U887 ( .A(n750), .B(n19722), .Z(n752) );
  XNOR U888 ( .A(b[5]), .B(n1495), .Z(n808) );
  NANDN U889 ( .A(n19640), .B(n808), .Z(n751) );
  AND U890 ( .A(n752), .B(n751), .Z(n803) );
  XNOR U891 ( .A(n802), .B(n803), .Z(n804) );
  XNOR U892 ( .A(n805), .B(n804), .Z(n829) );
  NANDN U893 ( .A(n753), .B(n19767), .Z(n755) );
  XNOR U894 ( .A(n19714), .B(n1354), .Z(n811) );
  NANDN U895 ( .A(n811), .B(n19766), .Z(n754) );
  NAND U896 ( .A(n755), .B(n754), .Z(n830) );
  XOR U897 ( .A(n829), .B(n830), .Z(n832) );
  NAND U898 ( .A(n757), .B(n756), .Z(n789) );
  IV U899 ( .A(a[14]), .Z(n1639) );
  XNOR U900 ( .A(n100), .B(n1639), .Z(n814) );
  OR U901 ( .A(n814), .B(n19521), .Z(n760) );
  NANDN U902 ( .A(n758), .B(n19554), .Z(n759) );
  NAND U903 ( .A(n760), .B(n759), .Z(n787) );
  NAND U904 ( .A(n19937), .B(n761), .Z(n763) );
  XOR U905 ( .A(b[9]), .B(a[8]), .Z(n799) );
  NAND U906 ( .A(n19883), .B(n799), .Z(n762) );
  AND U907 ( .A(n763), .B(n762), .Z(n786) );
  XNOR U908 ( .A(n787), .B(n786), .Z(n788) );
  XNOR U909 ( .A(n789), .B(n788), .Z(n831) );
  XNOR U910 ( .A(n832), .B(n831), .Z(n839) );
  OR U911 ( .A(n765), .B(n764), .Z(n769) );
  NAND U912 ( .A(n767), .B(n766), .Z(n768) );
  NAND U913 ( .A(n769), .B(n768), .Z(n840) );
  XNOR U914 ( .A(n839), .B(n840), .Z(n841) );
  XNOR U915 ( .A(n842), .B(n841), .Z(n781) );
  XOR U916 ( .A(n781), .B(n780), .Z(n782) );
  XNOR U917 ( .A(n783), .B(n782), .Z(n775) );
  XNOR U918 ( .A(n774), .B(n775), .Z(n776) );
  XOR U919 ( .A(n777), .B(n776), .Z(n846) );
  XOR U920 ( .A(n847), .B(n846), .Z(c[256]) );
  NANDN U921 ( .A(n775), .B(n774), .Z(n779) );
  NAND U922 ( .A(n777), .B(n776), .Z(n778) );
  NAND U923 ( .A(n779), .B(n778), .Z(n853) );
  OR U924 ( .A(n781), .B(n780), .Z(n785) );
  NAND U925 ( .A(n783), .B(n782), .Z(n784) );
  NAND U926 ( .A(n785), .B(n784), .Z(n851) );
  NANDN U927 ( .A(n787), .B(n786), .Z(n791) );
  NAND U928 ( .A(n789), .B(n788), .Z(n790) );
  NAND U929 ( .A(n791), .B(n790), .Z(n868) );
  XNOR U930 ( .A(n20052), .B(n1093), .Z(n874) );
  OR U931 ( .A(n874), .B(n20020), .Z(n794) );
  NANDN U932 ( .A(n792), .B(n19960), .Z(n793) );
  NAND U933 ( .A(n794), .B(n793), .Z(n887) );
  XNOR U934 ( .A(n102), .B(n795), .Z(n878) );
  OR U935 ( .A(n878), .B(n20121), .Z(n798) );
  NANDN U936 ( .A(n796), .B(n20122), .Z(n797) );
  NAND U937 ( .A(n798), .B(n797), .Z(n884) );
  XNOR U938 ( .A(n19975), .B(n1276), .Z(n881) );
  NANDN U939 ( .A(n881), .B(n19883), .Z(n801) );
  NAND U940 ( .A(n799), .B(n19937), .Z(n800) );
  AND U941 ( .A(n801), .B(n800), .Z(n885) );
  XNOR U942 ( .A(n884), .B(n885), .Z(n886) );
  XOR U943 ( .A(n887), .B(n886), .Z(n869) );
  XNOR U944 ( .A(n868), .B(n869), .Z(n870) );
  NANDN U945 ( .A(n803), .B(n802), .Z(n807) );
  NAND U946 ( .A(n805), .B(n804), .Z(n806) );
  NAND U947 ( .A(n807), .B(n806), .Z(n871) );
  XOR U948 ( .A(n870), .B(n871), .Z(n865) );
  NAND U949 ( .A(n19722), .B(n808), .Z(n810) );
  IV U950 ( .A(a[13]), .Z(n1561) );
  XNOR U951 ( .A(b[5]), .B(n1561), .Z(n912) );
  NANDN U952 ( .A(n19640), .B(n912), .Z(n809) );
  NAND U953 ( .A(n810), .B(n809), .Z(n893) );
  XNOR U954 ( .A(n19714), .B(n1432), .Z(n915) );
  NANDN U955 ( .A(n915), .B(n19766), .Z(n813) );
  NANDN U956 ( .A(n811), .B(n19767), .Z(n812) );
  NAND U957 ( .A(n813), .B(n812), .Z(n890) );
  NANDN U958 ( .A(n814), .B(n19554), .Z(n816) );
  IV U959 ( .A(a[15]), .Z(n1717) );
  XNOR U960 ( .A(b[3]), .B(n1717), .Z(n918) );
  NANDN U961 ( .A(n19521), .B(n918), .Z(n815) );
  AND U962 ( .A(n816), .B(n815), .Z(n891) );
  XNOR U963 ( .A(n890), .B(n891), .Z(n892) );
  XNOR U964 ( .A(n893), .B(n892), .Z(n899) );
  XNOR U965 ( .A(n20154), .B(n966), .Z(n906) );
  OR U966 ( .A(n906), .B(n20057), .Z(n819) );
  NANDN U967 ( .A(n817), .B(n20098), .Z(n818) );
  NAND U968 ( .A(n819), .B(n818), .Z(n905) );
  NAND U969 ( .A(b[0]), .B(a[17]), .Z(n820) );
  XNOR U970 ( .A(b[1]), .B(n820), .Z(n822) );
  NAND U971 ( .A(a[16]), .B(n98), .Z(n821) );
  AND U972 ( .A(n822), .B(n821), .Z(n902) );
  NAND U973 ( .A(b[15]), .B(a[1]), .Z(n903) );
  XOR U974 ( .A(n902), .B(n903), .Z(n904) );
  XOR U975 ( .A(n905), .B(n904), .Z(n896) );
  NANDN U976 ( .A(n824), .B(n823), .Z(n828) );
  NAND U977 ( .A(n826), .B(n825), .Z(n827) );
  NAND U978 ( .A(n828), .B(n827), .Z(n897) );
  XNOR U979 ( .A(n896), .B(n897), .Z(n898) );
  XOR U980 ( .A(n899), .B(n898), .Z(n862) );
  NANDN U981 ( .A(n830), .B(n829), .Z(n834) );
  OR U982 ( .A(n832), .B(n831), .Z(n833) );
  NAND U983 ( .A(n834), .B(n833), .Z(n863) );
  XOR U984 ( .A(n862), .B(n863), .Z(n864) );
  XNOR U985 ( .A(n865), .B(n864), .Z(n859) );
  NANDN U986 ( .A(n840), .B(n839), .Z(n844) );
  NANDN U987 ( .A(n842), .B(n841), .Z(n843) );
  NAND U988 ( .A(n844), .B(n843), .Z(n857) );
  XNOR U989 ( .A(n856), .B(n857), .Z(n858) );
  XOR U990 ( .A(n859), .B(n858), .Z(n850) );
  XOR U991 ( .A(n851), .B(n850), .Z(n852) );
  XNOR U992 ( .A(n853), .B(n852), .Z(n921) );
  XNOR U993 ( .A(n921), .B(sreg[257]), .Z(n923) );
  NAND U994 ( .A(n845), .B(sreg[256]), .Z(n849) );
  OR U995 ( .A(n847), .B(n846), .Z(n848) );
  AND U996 ( .A(n849), .B(n848), .Z(n922) );
  XOR U997 ( .A(n923), .B(n922), .Z(c[257]) );
  NAND U998 ( .A(n851), .B(n850), .Z(n855) );
  NAND U999 ( .A(n853), .B(n852), .Z(n854) );
  NAND U1000 ( .A(n855), .B(n854), .Z(n929) );
  NANDN U1001 ( .A(n857), .B(n856), .Z(n861) );
  NAND U1002 ( .A(n859), .B(n858), .Z(n860) );
  NAND U1003 ( .A(n861), .B(n860), .Z(n926) );
  OR U1004 ( .A(n863), .B(n862), .Z(n867) );
  NAND U1005 ( .A(n865), .B(n864), .Z(n866) );
  NAND U1006 ( .A(n867), .B(n866), .Z(n994) );
  NANDN U1007 ( .A(n869), .B(n868), .Z(n873) );
  NANDN U1008 ( .A(n871), .B(n870), .Z(n872) );
  NAND U1009 ( .A(n873), .B(n872), .Z(n991) );
  XNOR U1010 ( .A(n20052), .B(n1171), .Z(n963) );
  OR U1011 ( .A(n963), .B(n20020), .Z(n876) );
  NANDN U1012 ( .A(n874), .B(n19960), .Z(n875) );
  NAND U1013 ( .A(n876), .B(n875), .Z(n976) );
  XNOR U1014 ( .A(n102), .B(n877), .Z(n967) );
  OR U1015 ( .A(n967), .B(n20121), .Z(n880) );
  NANDN U1016 ( .A(n878), .B(n20122), .Z(n879) );
  NAND U1017 ( .A(n880), .B(n879), .Z(n973) );
  XNOR U1018 ( .A(n19975), .B(n1354), .Z(n970) );
  NANDN U1019 ( .A(n970), .B(n19883), .Z(n883) );
  NANDN U1020 ( .A(n881), .B(n19937), .Z(n882) );
  AND U1021 ( .A(n883), .B(n882), .Z(n974) );
  XNOR U1022 ( .A(n973), .B(n974), .Z(n975) );
  XNOR U1023 ( .A(n976), .B(n975), .Z(n985) );
  NANDN U1024 ( .A(n885), .B(n884), .Z(n889) );
  NAND U1025 ( .A(n887), .B(n886), .Z(n888) );
  NAND U1026 ( .A(n889), .B(n888), .Z(n986) );
  XOR U1027 ( .A(n985), .B(n986), .Z(n988) );
  NANDN U1028 ( .A(n891), .B(n890), .Z(n895) );
  NAND U1029 ( .A(n893), .B(n892), .Z(n894) );
  NAND U1030 ( .A(n895), .B(n894), .Z(n987) );
  XNOR U1031 ( .A(n988), .B(n987), .Z(n935) );
  NANDN U1032 ( .A(n897), .B(n896), .Z(n901) );
  NAND U1033 ( .A(n899), .B(n898), .Z(n900) );
  NAND U1034 ( .A(n901), .B(n900), .Z(n933) );
  XNOR U1035 ( .A(n20154), .B(n1042), .Z(n945) );
  OR U1036 ( .A(n945), .B(n20057), .Z(n908) );
  NANDN U1037 ( .A(n906), .B(n20098), .Z(n907) );
  AND U1038 ( .A(n908), .B(n907), .Z(n937) );
  NAND U1039 ( .A(b[0]), .B(a[18]), .Z(n909) );
  XNOR U1040 ( .A(b[1]), .B(n909), .Z(n911) );
  NAND U1041 ( .A(a[17]), .B(n98), .Z(n910) );
  AND U1042 ( .A(n911), .B(n910), .Z(n936) );
  XOR U1043 ( .A(n937), .B(n936), .Z(n939) );
  NAND U1044 ( .A(a[2]), .B(b[15]), .Z(n938) );
  XOR U1045 ( .A(n939), .B(n938), .Z(n957) );
  NAND U1046 ( .A(n19722), .B(n912), .Z(n914) );
  XNOR U1047 ( .A(b[5]), .B(n1639), .Z(n948) );
  NANDN U1048 ( .A(n19640), .B(n948), .Z(n913) );
  NAND U1049 ( .A(n914), .B(n913), .Z(n982) );
  XNOR U1050 ( .A(n19714), .B(n1495), .Z(n951) );
  NANDN U1051 ( .A(n951), .B(n19766), .Z(n917) );
  NANDN U1052 ( .A(n915), .B(n19767), .Z(n916) );
  NAND U1053 ( .A(n917), .B(n916), .Z(n979) );
  NAND U1054 ( .A(n19554), .B(n918), .Z(n920) );
  IV U1055 ( .A(a[16]), .Z(n1793) );
  XNOR U1056 ( .A(b[3]), .B(n1793), .Z(n954) );
  NANDN U1057 ( .A(n19521), .B(n954), .Z(n919) );
  AND U1058 ( .A(n920), .B(n919), .Z(n980) );
  XNOR U1059 ( .A(n979), .B(n980), .Z(n981) );
  XOR U1060 ( .A(n982), .B(n981), .Z(n958) );
  XOR U1061 ( .A(n957), .B(n958), .Z(n959) );
  XOR U1062 ( .A(n960), .B(n959), .Z(n932) );
  XOR U1063 ( .A(n933), .B(n932), .Z(n934) );
  XOR U1064 ( .A(n935), .B(n934), .Z(n992) );
  XOR U1065 ( .A(n991), .B(n992), .Z(n993) );
  XOR U1066 ( .A(n994), .B(n993), .Z(n927) );
  XNOR U1067 ( .A(n926), .B(n927), .Z(n928) );
  XNOR U1068 ( .A(n929), .B(n928), .Z(n997) );
  XNOR U1069 ( .A(n997), .B(sreg[258]), .Z(n999) );
  NAND U1070 ( .A(n921), .B(sreg[257]), .Z(n925) );
  OR U1071 ( .A(n923), .B(n922), .Z(n924) );
  AND U1072 ( .A(n925), .B(n924), .Z(n998) );
  XOR U1073 ( .A(n999), .B(n998), .Z(c[258]) );
  NANDN U1074 ( .A(n927), .B(n926), .Z(n931) );
  NAND U1075 ( .A(n929), .B(n928), .Z(n930) );
  NAND U1076 ( .A(n931), .B(n930), .Z(n1005) );
  NANDN U1077 ( .A(n937), .B(n936), .Z(n941) );
  OR U1078 ( .A(n939), .B(n938), .Z(n940) );
  NAND U1079 ( .A(n941), .B(n940), .Z(n1036) );
  NAND U1080 ( .A(b[0]), .B(a[19]), .Z(n942) );
  XNOR U1081 ( .A(b[1]), .B(n942), .Z(n944) );
  NAND U1082 ( .A(a[18]), .B(n98), .Z(n943) );
  AND U1083 ( .A(n944), .B(n943), .Z(n1012) );
  XNOR U1084 ( .A(n20154), .B(n1093), .Z(n1021) );
  OR U1085 ( .A(n1021), .B(n20057), .Z(n947) );
  NANDN U1086 ( .A(n945), .B(n20098), .Z(n946) );
  AND U1087 ( .A(n947), .B(n946), .Z(n1013) );
  XOR U1088 ( .A(n1012), .B(n1013), .Z(n1015) );
  NAND U1089 ( .A(a[3]), .B(b[15]), .Z(n1014) );
  XOR U1090 ( .A(n1015), .B(n1014), .Z(n1033) );
  NAND U1091 ( .A(n19722), .B(n948), .Z(n950) );
  XNOR U1092 ( .A(b[5]), .B(n1717), .Z(n1024) );
  NANDN U1093 ( .A(n19640), .B(n1024), .Z(n949) );
  NAND U1094 ( .A(n950), .B(n949), .Z(n1058) );
  XNOR U1095 ( .A(n19714), .B(n1561), .Z(n1027) );
  NANDN U1096 ( .A(n1027), .B(n19766), .Z(n953) );
  NANDN U1097 ( .A(n951), .B(n19767), .Z(n952) );
  NAND U1098 ( .A(n953), .B(n952), .Z(n1055) );
  NAND U1099 ( .A(n19554), .B(n954), .Z(n956) );
  IV U1100 ( .A(a[17]), .Z(n1871) );
  XNOR U1101 ( .A(b[3]), .B(n1871), .Z(n1030) );
  NANDN U1102 ( .A(n19521), .B(n1030), .Z(n955) );
  AND U1103 ( .A(n956), .B(n955), .Z(n1056) );
  XNOR U1104 ( .A(n1055), .B(n1056), .Z(n1057) );
  XOR U1105 ( .A(n1058), .B(n1057), .Z(n1034) );
  XOR U1106 ( .A(n1033), .B(n1034), .Z(n1035) );
  XNOR U1107 ( .A(n1036), .B(n1035), .Z(n1006) );
  NAND U1108 ( .A(n958), .B(n957), .Z(n962) );
  NAND U1109 ( .A(n960), .B(n959), .Z(n961) );
  NAND U1110 ( .A(n962), .B(n961), .Z(n1007) );
  XOR U1111 ( .A(n1006), .B(n1007), .Z(n1009) );
  XNOR U1112 ( .A(n20052), .B(n1276), .Z(n1039) );
  OR U1113 ( .A(n1039), .B(n20020), .Z(n965) );
  NANDN U1114 ( .A(n963), .B(n19960), .Z(n964) );
  NAND U1115 ( .A(n965), .B(n964), .Z(n1052) );
  XNOR U1116 ( .A(n102), .B(n966), .Z(n1043) );
  OR U1117 ( .A(n1043), .B(n20121), .Z(n969) );
  NANDN U1118 ( .A(n967), .B(n20122), .Z(n968) );
  NAND U1119 ( .A(n969), .B(n968), .Z(n1049) );
  XNOR U1120 ( .A(n19975), .B(n1432), .Z(n1046) );
  NANDN U1121 ( .A(n1046), .B(n19883), .Z(n972) );
  NANDN U1122 ( .A(n970), .B(n19937), .Z(n971) );
  AND U1123 ( .A(n972), .B(n971), .Z(n1050) );
  XNOR U1124 ( .A(n1049), .B(n1050), .Z(n1051) );
  XNOR U1125 ( .A(n1052), .B(n1051), .Z(n1061) );
  NANDN U1126 ( .A(n974), .B(n973), .Z(n978) );
  NAND U1127 ( .A(n976), .B(n975), .Z(n977) );
  NAND U1128 ( .A(n978), .B(n977), .Z(n1062) );
  XNOR U1129 ( .A(n1061), .B(n1062), .Z(n1063) );
  NANDN U1130 ( .A(n980), .B(n979), .Z(n984) );
  NAND U1131 ( .A(n982), .B(n981), .Z(n983) );
  AND U1132 ( .A(n984), .B(n983), .Z(n1064) );
  XNOR U1133 ( .A(n1063), .B(n1064), .Z(n1008) );
  XNOR U1134 ( .A(n1009), .B(n1008), .Z(n1067) );
  NANDN U1135 ( .A(n986), .B(n985), .Z(n990) );
  OR U1136 ( .A(n988), .B(n987), .Z(n989) );
  NAND U1137 ( .A(n990), .B(n989), .Z(n1068) );
  XNOR U1138 ( .A(n1067), .B(n1068), .Z(n1069) );
  XNOR U1139 ( .A(n1070), .B(n1069), .Z(n1002) );
  OR U1140 ( .A(n992), .B(n991), .Z(n996) );
  NAND U1141 ( .A(n994), .B(n993), .Z(n995) );
  NAND U1142 ( .A(n996), .B(n995), .Z(n1003) );
  XOR U1143 ( .A(n1002), .B(n1003), .Z(n1004) );
  XOR U1144 ( .A(n1005), .B(n1004), .Z(n1073) );
  XNOR U1145 ( .A(n1073), .B(sreg[259]), .Z(n1075) );
  NAND U1146 ( .A(n997), .B(sreg[258]), .Z(n1001) );
  OR U1147 ( .A(n999), .B(n998), .Z(n1000) );
  AND U1148 ( .A(n1001), .B(n1000), .Z(n1074) );
  XOR U1149 ( .A(n1075), .B(n1074), .Z(c[259]) );
  NANDN U1150 ( .A(n1007), .B(n1006), .Z(n1011) );
  OR U1151 ( .A(n1009), .B(n1008), .Z(n1010) );
  NAND U1152 ( .A(n1011), .B(n1010), .Z(n1148) );
  NANDN U1153 ( .A(n1013), .B(n1012), .Z(n1017) );
  OR U1154 ( .A(n1015), .B(n1014), .Z(n1016) );
  NAND U1155 ( .A(n1017), .B(n1016), .Z(n1136) );
  NAND U1156 ( .A(b[0]), .B(a[20]), .Z(n1018) );
  XNOR U1157 ( .A(b[1]), .B(n1018), .Z(n1020) );
  NAND U1158 ( .A(a[19]), .B(n98), .Z(n1019) );
  AND U1159 ( .A(n1020), .B(n1019), .Z(n1112) );
  XNOR U1160 ( .A(n20154), .B(n1171), .Z(n1121) );
  OR U1161 ( .A(n1121), .B(n20057), .Z(n1023) );
  NANDN U1162 ( .A(n1021), .B(n20098), .Z(n1022) );
  AND U1163 ( .A(n1023), .B(n1022), .Z(n1113) );
  XOR U1164 ( .A(n1112), .B(n1113), .Z(n1115) );
  NAND U1165 ( .A(a[4]), .B(b[15]), .Z(n1114) );
  XOR U1166 ( .A(n1115), .B(n1114), .Z(n1133) );
  NAND U1167 ( .A(n19722), .B(n1024), .Z(n1026) );
  XNOR U1168 ( .A(b[5]), .B(n1793), .Z(n1124) );
  NANDN U1169 ( .A(n19640), .B(n1124), .Z(n1025) );
  NAND U1170 ( .A(n1026), .B(n1025), .Z(n1109) );
  XNOR U1171 ( .A(n19714), .B(n1639), .Z(n1127) );
  NANDN U1172 ( .A(n1127), .B(n19766), .Z(n1029) );
  NANDN U1173 ( .A(n1027), .B(n19767), .Z(n1028) );
  NAND U1174 ( .A(n1029), .B(n1028), .Z(n1106) );
  NAND U1175 ( .A(n19554), .B(n1030), .Z(n1032) );
  IV U1176 ( .A(a[18]), .Z(n1976) );
  XNOR U1177 ( .A(b[3]), .B(n1976), .Z(n1130) );
  NANDN U1178 ( .A(n19521), .B(n1130), .Z(n1031) );
  AND U1179 ( .A(n1032), .B(n1031), .Z(n1107) );
  XNOR U1180 ( .A(n1106), .B(n1107), .Z(n1108) );
  XOR U1181 ( .A(n1109), .B(n1108), .Z(n1134) );
  XOR U1182 ( .A(n1133), .B(n1134), .Z(n1135) );
  XNOR U1183 ( .A(n1136), .B(n1135), .Z(n1084) );
  NAND U1184 ( .A(n1034), .B(n1033), .Z(n1038) );
  NAND U1185 ( .A(n1036), .B(n1035), .Z(n1037) );
  NAND U1186 ( .A(n1038), .B(n1037), .Z(n1085) );
  XOR U1187 ( .A(n1084), .B(n1085), .Z(n1087) );
  XNOR U1188 ( .A(n20052), .B(n1354), .Z(n1090) );
  OR U1189 ( .A(n1090), .B(n20020), .Z(n1041) );
  NANDN U1190 ( .A(n1039), .B(n19960), .Z(n1040) );
  NAND U1191 ( .A(n1041), .B(n1040), .Z(n1103) );
  XNOR U1192 ( .A(n102), .B(n1042), .Z(n1094) );
  OR U1193 ( .A(n1094), .B(n20121), .Z(n1045) );
  NANDN U1194 ( .A(n1043), .B(n20122), .Z(n1044) );
  NAND U1195 ( .A(n1045), .B(n1044), .Z(n1100) );
  XNOR U1196 ( .A(n19975), .B(n1495), .Z(n1097) );
  NANDN U1197 ( .A(n1097), .B(n19883), .Z(n1048) );
  NANDN U1198 ( .A(n1046), .B(n19937), .Z(n1047) );
  AND U1199 ( .A(n1048), .B(n1047), .Z(n1101) );
  XNOR U1200 ( .A(n1100), .B(n1101), .Z(n1102) );
  XNOR U1201 ( .A(n1103), .B(n1102), .Z(n1139) );
  NANDN U1202 ( .A(n1050), .B(n1049), .Z(n1054) );
  NAND U1203 ( .A(n1052), .B(n1051), .Z(n1053) );
  NAND U1204 ( .A(n1054), .B(n1053), .Z(n1140) );
  XNOR U1205 ( .A(n1139), .B(n1140), .Z(n1141) );
  NANDN U1206 ( .A(n1056), .B(n1055), .Z(n1060) );
  NAND U1207 ( .A(n1058), .B(n1057), .Z(n1059) );
  AND U1208 ( .A(n1060), .B(n1059), .Z(n1142) );
  XNOR U1209 ( .A(n1141), .B(n1142), .Z(n1086) );
  XNOR U1210 ( .A(n1087), .B(n1086), .Z(n1145) );
  NANDN U1211 ( .A(n1062), .B(n1061), .Z(n1066) );
  NAND U1212 ( .A(n1064), .B(n1063), .Z(n1065) );
  NAND U1213 ( .A(n1066), .B(n1065), .Z(n1146) );
  XNOR U1214 ( .A(n1145), .B(n1146), .Z(n1147) );
  XOR U1215 ( .A(n1148), .B(n1147), .Z(n1078) );
  NANDN U1216 ( .A(n1068), .B(n1067), .Z(n1072) );
  NAND U1217 ( .A(n1070), .B(n1069), .Z(n1071) );
  NAND U1218 ( .A(n1072), .B(n1071), .Z(n1079) );
  XNOR U1219 ( .A(n1078), .B(n1079), .Z(n1080) );
  XNOR U1220 ( .A(n1081), .B(n1080), .Z(n1151) );
  XNOR U1221 ( .A(n1151), .B(sreg[260]), .Z(n1153) );
  NAND U1222 ( .A(n1073), .B(sreg[259]), .Z(n1077) );
  OR U1223 ( .A(n1075), .B(n1074), .Z(n1076) );
  AND U1224 ( .A(n1077), .B(n1076), .Z(n1152) );
  XOR U1225 ( .A(n1153), .B(n1152), .Z(c[260]) );
  NANDN U1226 ( .A(n1079), .B(n1078), .Z(n1083) );
  NAND U1227 ( .A(n1081), .B(n1080), .Z(n1082) );
  NAND U1228 ( .A(n1083), .B(n1082), .Z(n1159) );
  NANDN U1229 ( .A(n1085), .B(n1084), .Z(n1089) );
  OR U1230 ( .A(n1087), .B(n1086), .Z(n1088) );
  NAND U1231 ( .A(n1089), .B(n1088), .Z(n1226) );
  XNOR U1232 ( .A(n20052), .B(n1432), .Z(n1168) );
  OR U1233 ( .A(n1168), .B(n20020), .Z(n1092) );
  NANDN U1234 ( .A(n1090), .B(n19960), .Z(n1091) );
  NAND U1235 ( .A(n1092), .B(n1091), .Z(n1181) );
  XNOR U1236 ( .A(n102), .B(n1093), .Z(n1172) );
  OR U1237 ( .A(n1172), .B(n20121), .Z(n1096) );
  NANDN U1238 ( .A(n1094), .B(n20122), .Z(n1095) );
  NAND U1239 ( .A(n1096), .B(n1095), .Z(n1178) );
  XNOR U1240 ( .A(n19975), .B(n1561), .Z(n1175) );
  NANDN U1241 ( .A(n1175), .B(n19883), .Z(n1099) );
  NANDN U1242 ( .A(n1097), .B(n19937), .Z(n1098) );
  AND U1243 ( .A(n1099), .B(n1098), .Z(n1179) );
  XNOR U1244 ( .A(n1178), .B(n1179), .Z(n1180) );
  XNOR U1245 ( .A(n1181), .B(n1180), .Z(n1217) );
  NANDN U1246 ( .A(n1101), .B(n1100), .Z(n1105) );
  NAND U1247 ( .A(n1103), .B(n1102), .Z(n1104) );
  NAND U1248 ( .A(n1105), .B(n1104), .Z(n1218) );
  XNOR U1249 ( .A(n1217), .B(n1218), .Z(n1219) );
  NANDN U1250 ( .A(n1107), .B(n1106), .Z(n1111) );
  NAND U1251 ( .A(n1109), .B(n1108), .Z(n1110) );
  AND U1252 ( .A(n1111), .B(n1110), .Z(n1220) );
  XNOR U1253 ( .A(n1219), .B(n1220), .Z(n1164) );
  NANDN U1254 ( .A(n1113), .B(n1112), .Z(n1117) );
  OR U1255 ( .A(n1115), .B(n1114), .Z(n1116) );
  NAND U1256 ( .A(n1117), .B(n1116), .Z(n1214) );
  NAND U1257 ( .A(b[0]), .B(a[21]), .Z(n1118) );
  XNOR U1258 ( .A(b[1]), .B(n1118), .Z(n1120) );
  NAND U1259 ( .A(a[20]), .B(n98), .Z(n1119) );
  AND U1260 ( .A(n1120), .B(n1119), .Z(n1190) );
  XNOR U1261 ( .A(n20154), .B(n1276), .Z(n1196) );
  OR U1262 ( .A(n1196), .B(n20057), .Z(n1123) );
  NANDN U1263 ( .A(n1121), .B(n20098), .Z(n1122) );
  AND U1264 ( .A(n1123), .B(n1122), .Z(n1191) );
  XOR U1265 ( .A(n1190), .B(n1191), .Z(n1193) );
  NAND U1266 ( .A(a[5]), .B(b[15]), .Z(n1192) );
  XOR U1267 ( .A(n1193), .B(n1192), .Z(n1211) );
  NAND U1268 ( .A(n19722), .B(n1124), .Z(n1126) );
  XNOR U1269 ( .A(b[5]), .B(n1871), .Z(n1202) );
  NANDN U1270 ( .A(n19640), .B(n1202), .Z(n1125) );
  NAND U1271 ( .A(n1126), .B(n1125), .Z(n1187) );
  XNOR U1272 ( .A(n19714), .B(n1717), .Z(n1205) );
  NANDN U1273 ( .A(n1205), .B(n19766), .Z(n1129) );
  NANDN U1274 ( .A(n1127), .B(n19767), .Z(n1128) );
  NAND U1275 ( .A(n1129), .B(n1128), .Z(n1184) );
  NAND U1276 ( .A(n19554), .B(n1130), .Z(n1132) );
  IV U1277 ( .A(a[19]), .Z(n2027) );
  XNOR U1278 ( .A(b[3]), .B(n2027), .Z(n1208) );
  NANDN U1279 ( .A(n19521), .B(n1208), .Z(n1131) );
  AND U1280 ( .A(n1132), .B(n1131), .Z(n1185) );
  XNOR U1281 ( .A(n1184), .B(n1185), .Z(n1186) );
  XOR U1282 ( .A(n1187), .B(n1186), .Z(n1212) );
  XOR U1283 ( .A(n1211), .B(n1212), .Z(n1213) );
  XNOR U1284 ( .A(n1214), .B(n1213), .Z(n1162) );
  NAND U1285 ( .A(n1134), .B(n1133), .Z(n1138) );
  NAND U1286 ( .A(n1136), .B(n1135), .Z(n1137) );
  NAND U1287 ( .A(n1138), .B(n1137), .Z(n1163) );
  XOR U1288 ( .A(n1162), .B(n1163), .Z(n1165) );
  XNOR U1289 ( .A(n1164), .B(n1165), .Z(n1223) );
  NANDN U1290 ( .A(n1140), .B(n1139), .Z(n1144) );
  NAND U1291 ( .A(n1142), .B(n1141), .Z(n1143) );
  NAND U1292 ( .A(n1144), .B(n1143), .Z(n1224) );
  XNOR U1293 ( .A(n1223), .B(n1224), .Z(n1225) );
  XOR U1294 ( .A(n1226), .B(n1225), .Z(n1156) );
  NANDN U1295 ( .A(n1146), .B(n1145), .Z(n1150) );
  NANDN U1296 ( .A(n1148), .B(n1147), .Z(n1149) );
  NAND U1297 ( .A(n1150), .B(n1149), .Z(n1157) );
  XNOR U1298 ( .A(n1156), .B(n1157), .Z(n1158) );
  XNOR U1299 ( .A(n1159), .B(n1158), .Z(n1229) );
  XNOR U1300 ( .A(n1229), .B(sreg[261]), .Z(n1231) );
  NAND U1301 ( .A(n1151), .B(sreg[260]), .Z(n1155) );
  OR U1302 ( .A(n1153), .B(n1152), .Z(n1154) );
  AND U1303 ( .A(n1155), .B(n1154), .Z(n1230) );
  XOR U1304 ( .A(n1231), .B(n1230), .Z(c[261]) );
  NANDN U1305 ( .A(n1157), .B(n1156), .Z(n1161) );
  NAND U1306 ( .A(n1159), .B(n1158), .Z(n1160) );
  NAND U1307 ( .A(n1161), .B(n1160), .Z(n1237) );
  NANDN U1308 ( .A(n1163), .B(n1162), .Z(n1167) );
  OR U1309 ( .A(n1165), .B(n1164), .Z(n1166) );
  NAND U1310 ( .A(n1167), .B(n1166), .Z(n1304) );
  XNOR U1311 ( .A(n20052), .B(n1495), .Z(n1273) );
  OR U1312 ( .A(n1273), .B(n20020), .Z(n1170) );
  NANDN U1313 ( .A(n1168), .B(n19960), .Z(n1169) );
  NAND U1314 ( .A(n1170), .B(n1169), .Z(n1286) );
  XNOR U1315 ( .A(n102), .B(n1171), .Z(n1277) );
  OR U1316 ( .A(n1277), .B(n20121), .Z(n1174) );
  NANDN U1317 ( .A(n1172), .B(n20122), .Z(n1173) );
  NAND U1318 ( .A(n1174), .B(n1173), .Z(n1283) );
  XNOR U1319 ( .A(n19975), .B(n1639), .Z(n1280) );
  NANDN U1320 ( .A(n1280), .B(n19883), .Z(n1177) );
  NANDN U1321 ( .A(n1175), .B(n19937), .Z(n1176) );
  AND U1322 ( .A(n1177), .B(n1176), .Z(n1284) );
  XNOR U1323 ( .A(n1283), .B(n1284), .Z(n1285) );
  XNOR U1324 ( .A(n1286), .B(n1285), .Z(n1295) );
  NANDN U1325 ( .A(n1179), .B(n1178), .Z(n1183) );
  NAND U1326 ( .A(n1181), .B(n1180), .Z(n1182) );
  NAND U1327 ( .A(n1183), .B(n1182), .Z(n1296) );
  XNOR U1328 ( .A(n1295), .B(n1296), .Z(n1297) );
  NANDN U1329 ( .A(n1185), .B(n1184), .Z(n1189) );
  NAND U1330 ( .A(n1187), .B(n1186), .Z(n1188) );
  AND U1331 ( .A(n1189), .B(n1188), .Z(n1298) );
  XNOR U1332 ( .A(n1297), .B(n1298), .Z(n1242) );
  NANDN U1333 ( .A(n1191), .B(n1190), .Z(n1195) );
  OR U1334 ( .A(n1193), .B(n1192), .Z(n1194) );
  NAND U1335 ( .A(n1195), .B(n1194), .Z(n1270) );
  XNOR U1336 ( .A(n20154), .B(n1354), .Z(n1255) );
  OR U1337 ( .A(n1255), .B(n20057), .Z(n1198) );
  NANDN U1338 ( .A(n1196), .B(n20098), .Z(n1197) );
  AND U1339 ( .A(n1198), .B(n1197), .Z(n1247) );
  NAND U1340 ( .A(b[0]), .B(a[22]), .Z(n1199) );
  XNOR U1341 ( .A(b[1]), .B(n1199), .Z(n1201) );
  NAND U1342 ( .A(a[21]), .B(n98), .Z(n1200) );
  AND U1343 ( .A(n1201), .B(n1200), .Z(n1246) );
  XOR U1344 ( .A(n1247), .B(n1246), .Z(n1249) );
  NAND U1345 ( .A(a[6]), .B(b[15]), .Z(n1248) );
  XOR U1346 ( .A(n1249), .B(n1248), .Z(n1267) );
  NAND U1347 ( .A(n19722), .B(n1202), .Z(n1204) );
  XNOR U1348 ( .A(b[5]), .B(n1976), .Z(n1258) );
  NANDN U1349 ( .A(n19640), .B(n1258), .Z(n1203) );
  NAND U1350 ( .A(n1204), .B(n1203), .Z(n1292) );
  XNOR U1351 ( .A(n19714), .B(n1793), .Z(n1261) );
  NANDN U1352 ( .A(n1261), .B(n19766), .Z(n1207) );
  NANDN U1353 ( .A(n1205), .B(n19767), .Z(n1206) );
  NAND U1354 ( .A(n1207), .B(n1206), .Z(n1289) );
  NAND U1355 ( .A(n19554), .B(n1208), .Z(n1210) );
  IV U1356 ( .A(a[20]), .Z(n2105) );
  XNOR U1357 ( .A(b[3]), .B(n2105), .Z(n1264) );
  NANDN U1358 ( .A(n19521), .B(n1264), .Z(n1209) );
  AND U1359 ( .A(n1210), .B(n1209), .Z(n1290) );
  XNOR U1360 ( .A(n1289), .B(n1290), .Z(n1291) );
  XOR U1361 ( .A(n1292), .B(n1291), .Z(n1268) );
  XOR U1362 ( .A(n1267), .B(n1268), .Z(n1269) );
  XNOR U1363 ( .A(n1270), .B(n1269), .Z(n1240) );
  NAND U1364 ( .A(n1212), .B(n1211), .Z(n1216) );
  NAND U1365 ( .A(n1214), .B(n1213), .Z(n1215) );
  NAND U1366 ( .A(n1216), .B(n1215), .Z(n1241) );
  XOR U1367 ( .A(n1240), .B(n1241), .Z(n1243) );
  XNOR U1368 ( .A(n1242), .B(n1243), .Z(n1301) );
  NANDN U1369 ( .A(n1218), .B(n1217), .Z(n1222) );
  NAND U1370 ( .A(n1220), .B(n1219), .Z(n1221) );
  NAND U1371 ( .A(n1222), .B(n1221), .Z(n1302) );
  XNOR U1372 ( .A(n1301), .B(n1302), .Z(n1303) );
  XOR U1373 ( .A(n1304), .B(n1303), .Z(n1234) );
  NANDN U1374 ( .A(n1224), .B(n1223), .Z(n1228) );
  NANDN U1375 ( .A(n1226), .B(n1225), .Z(n1227) );
  NAND U1376 ( .A(n1228), .B(n1227), .Z(n1235) );
  XNOR U1377 ( .A(n1234), .B(n1235), .Z(n1236) );
  XNOR U1378 ( .A(n1237), .B(n1236), .Z(n1307) );
  XNOR U1379 ( .A(n1307), .B(sreg[262]), .Z(n1309) );
  NAND U1380 ( .A(n1229), .B(sreg[261]), .Z(n1233) );
  OR U1381 ( .A(n1231), .B(n1230), .Z(n1232) );
  AND U1382 ( .A(n1233), .B(n1232), .Z(n1308) );
  XOR U1383 ( .A(n1309), .B(n1308), .Z(c[262]) );
  NANDN U1384 ( .A(n1235), .B(n1234), .Z(n1239) );
  NAND U1385 ( .A(n1237), .B(n1236), .Z(n1238) );
  NAND U1386 ( .A(n1239), .B(n1238), .Z(n1315) );
  NANDN U1387 ( .A(n1241), .B(n1240), .Z(n1245) );
  OR U1388 ( .A(n1243), .B(n1242), .Z(n1244) );
  NAND U1389 ( .A(n1245), .B(n1244), .Z(n1382) );
  NANDN U1390 ( .A(n1247), .B(n1246), .Z(n1251) );
  OR U1391 ( .A(n1249), .B(n1248), .Z(n1250) );
  NAND U1392 ( .A(n1251), .B(n1250), .Z(n1348) );
  NAND U1393 ( .A(b[0]), .B(a[23]), .Z(n1252) );
  XNOR U1394 ( .A(b[1]), .B(n1252), .Z(n1254) );
  NAND U1395 ( .A(a[22]), .B(n98), .Z(n1253) );
  AND U1396 ( .A(n1254), .B(n1253), .Z(n1324) );
  XNOR U1397 ( .A(n20154), .B(n1432), .Z(n1333) );
  OR U1398 ( .A(n1333), .B(n20057), .Z(n1257) );
  NANDN U1399 ( .A(n1255), .B(n20098), .Z(n1256) );
  AND U1400 ( .A(n1257), .B(n1256), .Z(n1325) );
  XOR U1401 ( .A(n1324), .B(n1325), .Z(n1327) );
  NAND U1402 ( .A(a[7]), .B(b[15]), .Z(n1326) );
  XOR U1403 ( .A(n1327), .B(n1326), .Z(n1345) );
  NAND U1404 ( .A(n19722), .B(n1258), .Z(n1260) );
  XNOR U1405 ( .A(b[5]), .B(n2027), .Z(n1336) );
  NANDN U1406 ( .A(n19640), .B(n1336), .Z(n1259) );
  NAND U1407 ( .A(n1260), .B(n1259), .Z(n1370) );
  XNOR U1408 ( .A(n19714), .B(n1871), .Z(n1339) );
  NANDN U1409 ( .A(n1339), .B(n19766), .Z(n1263) );
  NANDN U1410 ( .A(n1261), .B(n19767), .Z(n1262) );
  NAND U1411 ( .A(n1263), .B(n1262), .Z(n1367) );
  NAND U1412 ( .A(n19554), .B(n1264), .Z(n1266) );
  IV U1413 ( .A(a[21]), .Z(n2195) );
  XNOR U1414 ( .A(b[3]), .B(n2195), .Z(n1342) );
  NANDN U1415 ( .A(n19521), .B(n1342), .Z(n1265) );
  AND U1416 ( .A(n1266), .B(n1265), .Z(n1368) );
  XNOR U1417 ( .A(n1367), .B(n1368), .Z(n1369) );
  XOR U1418 ( .A(n1370), .B(n1369), .Z(n1346) );
  XOR U1419 ( .A(n1345), .B(n1346), .Z(n1347) );
  XNOR U1420 ( .A(n1348), .B(n1347), .Z(n1318) );
  NAND U1421 ( .A(n1268), .B(n1267), .Z(n1272) );
  NAND U1422 ( .A(n1270), .B(n1269), .Z(n1271) );
  NAND U1423 ( .A(n1272), .B(n1271), .Z(n1319) );
  XOR U1424 ( .A(n1318), .B(n1319), .Z(n1321) );
  XNOR U1425 ( .A(n20052), .B(n1561), .Z(n1351) );
  OR U1426 ( .A(n1351), .B(n20020), .Z(n1275) );
  NANDN U1427 ( .A(n1273), .B(n19960), .Z(n1274) );
  NAND U1428 ( .A(n1275), .B(n1274), .Z(n1364) );
  XNOR U1429 ( .A(n102), .B(n1276), .Z(n1355) );
  OR U1430 ( .A(n1355), .B(n20121), .Z(n1279) );
  NANDN U1431 ( .A(n1277), .B(n20122), .Z(n1278) );
  NAND U1432 ( .A(n1279), .B(n1278), .Z(n1361) );
  XNOR U1433 ( .A(n19975), .B(n1717), .Z(n1358) );
  NANDN U1434 ( .A(n1358), .B(n19883), .Z(n1282) );
  NANDN U1435 ( .A(n1280), .B(n19937), .Z(n1281) );
  AND U1436 ( .A(n1282), .B(n1281), .Z(n1362) );
  XNOR U1437 ( .A(n1361), .B(n1362), .Z(n1363) );
  XNOR U1438 ( .A(n1364), .B(n1363), .Z(n1373) );
  NANDN U1439 ( .A(n1284), .B(n1283), .Z(n1288) );
  NAND U1440 ( .A(n1286), .B(n1285), .Z(n1287) );
  NAND U1441 ( .A(n1288), .B(n1287), .Z(n1374) );
  XNOR U1442 ( .A(n1373), .B(n1374), .Z(n1375) );
  NANDN U1443 ( .A(n1290), .B(n1289), .Z(n1294) );
  NAND U1444 ( .A(n1292), .B(n1291), .Z(n1293) );
  AND U1445 ( .A(n1294), .B(n1293), .Z(n1376) );
  XNOR U1446 ( .A(n1375), .B(n1376), .Z(n1320) );
  XNOR U1447 ( .A(n1321), .B(n1320), .Z(n1379) );
  NANDN U1448 ( .A(n1296), .B(n1295), .Z(n1300) );
  NAND U1449 ( .A(n1298), .B(n1297), .Z(n1299) );
  NAND U1450 ( .A(n1300), .B(n1299), .Z(n1380) );
  XNOR U1451 ( .A(n1379), .B(n1380), .Z(n1381) );
  XOR U1452 ( .A(n1382), .B(n1381), .Z(n1312) );
  NANDN U1453 ( .A(n1302), .B(n1301), .Z(n1306) );
  NANDN U1454 ( .A(n1304), .B(n1303), .Z(n1305) );
  NAND U1455 ( .A(n1306), .B(n1305), .Z(n1313) );
  XNOR U1456 ( .A(n1312), .B(n1313), .Z(n1314) );
  XNOR U1457 ( .A(n1315), .B(n1314), .Z(n1385) );
  XNOR U1458 ( .A(n1385), .B(sreg[263]), .Z(n1387) );
  NAND U1459 ( .A(n1307), .B(sreg[262]), .Z(n1311) );
  OR U1460 ( .A(n1309), .B(n1308), .Z(n1310) );
  AND U1461 ( .A(n1311), .B(n1310), .Z(n1386) );
  XOR U1462 ( .A(n1387), .B(n1386), .Z(c[263]) );
  NANDN U1463 ( .A(n1313), .B(n1312), .Z(n1317) );
  NAND U1464 ( .A(n1315), .B(n1314), .Z(n1316) );
  NAND U1465 ( .A(n1317), .B(n1316), .Z(n1393) );
  NANDN U1466 ( .A(n1319), .B(n1318), .Z(n1323) );
  OR U1467 ( .A(n1321), .B(n1320), .Z(n1322) );
  NAND U1468 ( .A(n1323), .B(n1322), .Z(n1460) );
  NANDN U1469 ( .A(n1325), .B(n1324), .Z(n1329) );
  OR U1470 ( .A(n1327), .B(n1326), .Z(n1328) );
  NAND U1471 ( .A(n1329), .B(n1328), .Z(n1426) );
  NAND U1472 ( .A(b[0]), .B(a[24]), .Z(n1330) );
  XNOR U1473 ( .A(b[1]), .B(n1330), .Z(n1332) );
  NAND U1474 ( .A(a[23]), .B(n98), .Z(n1331) );
  AND U1475 ( .A(n1332), .B(n1331), .Z(n1402) );
  XNOR U1476 ( .A(n20154), .B(n1495), .Z(n1411) );
  OR U1477 ( .A(n1411), .B(n20057), .Z(n1335) );
  NANDN U1478 ( .A(n1333), .B(n20098), .Z(n1334) );
  AND U1479 ( .A(n1335), .B(n1334), .Z(n1403) );
  XOR U1480 ( .A(n1402), .B(n1403), .Z(n1405) );
  NAND U1481 ( .A(a[8]), .B(b[15]), .Z(n1404) );
  XOR U1482 ( .A(n1405), .B(n1404), .Z(n1423) );
  NAND U1483 ( .A(n19722), .B(n1336), .Z(n1338) );
  XNOR U1484 ( .A(b[5]), .B(n2105), .Z(n1414) );
  NANDN U1485 ( .A(n19640), .B(n1414), .Z(n1337) );
  NAND U1486 ( .A(n1338), .B(n1337), .Z(n1448) );
  XNOR U1487 ( .A(n19714), .B(n1976), .Z(n1417) );
  NANDN U1488 ( .A(n1417), .B(n19766), .Z(n1341) );
  NANDN U1489 ( .A(n1339), .B(n19767), .Z(n1340) );
  NAND U1490 ( .A(n1341), .B(n1340), .Z(n1445) );
  NAND U1491 ( .A(n19554), .B(n1342), .Z(n1344) );
  IV U1492 ( .A(a[22]), .Z(n2261) );
  XNOR U1493 ( .A(b[3]), .B(n2261), .Z(n1420) );
  NANDN U1494 ( .A(n19521), .B(n1420), .Z(n1343) );
  AND U1495 ( .A(n1344), .B(n1343), .Z(n1446) );
  XNOR U1496 ( .A(n1445), .B(n1446), .Z(n1447) );
  XOR U1497 ( .A(n1448), .B(n1447), .Z(n1424) );
  XOR U1498 ( .A(n1423), .B(n1424), .Z(n1425) );
  XNOR U1499 ( .A(n1426), .B(n1425), .Z(n1396) );
  NAND U1500 ( .A(n1346), .B(n1345), .Z(n1350) );
  NAND U1501 ( .A(n1348), .B(n1347), .Z(n1349) );
  NAND U1502 ( .A(n1350), .B(n1349), .Z(n1397) );
  XOR U1503 ( .A(n1396), .B(n1397), .Z(n1399) );
  XNOR U1504 ( .A(n20052), .B(n1639), .Z(n1429) );
  OR U1505 ( .A(n1429), .B(n20020), .Z(n1353) );
  NANDN U1506 ( .A(n1351), .B(n19960), .Z(n1352) );
  NAND U1507 ( .A(n1353), .B(n1352), .Z(n1442) );
  XNOR U1508 ( .A(n102), .B(n1354), .Z(n1433) );
  OR U1509 ( .A(n1433), .B(n20121), .Z(n1357) );
  NANDN U1510 ( .A(n1355), .B(n20122), .Z(n1356) );
  NAND U1511 ( .A(n1357), .B(n1356), .Z(n1439) );
  XNOR U1512 ( .A(n19975), .B(n1793), .Z(n1436) );
  NANDN U1513 ( .A(n1436), .B(n19883), .Z(n1360) );
  NANDN U1514 ( .A(n1358), .B(n19937), .Z(n1359) );
  AND U1515 ( .A(n1360), .B(n1359), .Z(n1440) );
  XNOR U1516 ( .A(n1439), .B(n1440), .Z(n1441) );
  XNOR U1517 ( .A(n1442), .B(n1441), .Z(n1451) );
  NANDN U1518 ( .A(n1362), .B(n1361), .Z(n1366) );
  NAND U1519 ( .A(n1364), .B(n1363), .Z(n1365) );
  NAND U1520 ( .A(n1366), .B(n1365), .Z(n1452) );
  XNOR U1521 ( .A(n1451), .B(n1452), .Z(n1453) );
  NANDN U1522 ( .A(n1368), .B(n1367), .Z(n1372) );
  NAND U1523 ( .A(n1370), .B(n1369), .Z(n1371) );
  AND U1524 ( .A(n1372), .B(n1371), .Z(n1454) );
  XNOR U1525 ( .A(n1453), .B(n1454), .Z(n1398) );
  XNOR U1526 ( .A(n1399), .B(n1398), .Z(n1457) );
  NANDN U1527 ( .A(n1374), .B(n1373), .Z(n1378) );
  NAND U1528 ( .A(n1376), .B(n1375), .Z(n1377) );
  NAND U1529 ( .A(n1378), .B(n1377), .Z(n1458) );
  XNOR U1530 ( .A(n1457), .B(n1458), .Z(n1459) );
  XOR U1531 ( .A(n1460), .B(n1459), .Z(n1390) );
  NANDN U1532 ( .A(n1380), .B(n1379), .Z(n1384) );
  NANDN U1533 ( .A(n1382), .B(n1381), .Z(n1383) );
  NAND U1534 ( .A(n1384), .B(n1383), .Z(n1391) );
  XNOR U1535 ( .A(n1390), .B(n1391), .Z(n1392) );
  XNOR U1536 ( .A(n1393), .B(n1392), .Z(n1463) );
  XNOR U1537 ( .A(n1463), .B(sreg[264]), .Z(n1465) );
  NAND U1538 ( .A(n1385), .B(sreg[263]), .Z(n1389) );
  OR U1539 ( .A(n1387), .B(n1386), .Z(n1388) );
  AND U1540 ( .A(n1389), .B(n1388), .Z(n1464) );
  XOR U1541 ( .A(n1465), .B(n1464), .Z(c[264]) );
  NANDN U1542 ( .A(n1391), .B(n1390), .Z(n1395) );
  NAND U1543 ( .A(n1393), .B(n1392), .Z(n1394) );
  NAND U1544 ( .A(n1395), .B(n1394), .Z(n1471) );
  NANDN U1545 ( .A(n1397), .B(n1396), .Z(n1401) );
  OR U1546 ( .A(n1399), .B(n1398), .Z(n1400) );
  NAND U1547 ( .A(n1401), .B(n1400), .Z(n1538) );
  NANDN U1548 ( .A(n1403), .B(n1402), .Z(n1407) );
  OR U1549 ( .A(n1405), .B(n1404), .Z(n1406) );
  NAND U1550 ( .A(n1407), .B(n1406), .Z(n1526) );
  NAND U1551 ( .A(b[0]), .B(a[25]), .Z(n1408) );
  XNOR U1552 ( .A(b[1]), .B(n1408), .Z(n1410) );
  NAND U1553 ( .A(a[24]), .B(n98), .Z(n1409) );
  AND U1554 ( .A(n1410), .B(n1409), .Z(n1502) );
  XNOR U1555 ( .A(n20154), .B(n1561), .Z(n1511) );
  OR U1556 ( .A(n1511), .B(n20057), .Z(n1413) );
  NANDN U1557 ( .A(n1411), .B(n20098), .Z(n1412) );
  AND U1558 ( .A(n1413), .B(n1412), .Z(n1503) );
  XOR U1559 ( .A(n1502), .B(n1503), .Z(n1505) );
  NAND U1560 ( .A(a[9]), .B(b[15]), .Z(n1504) );
  XOR U1561 ( .A(n1505), .B(n1504), .Z(n1523) );
  NAND U1562 ( .A(n19722), .B(n1414), .Z(n1416) );
  XNOR U1563 ( .A(b[5]), .B(n2195), .Z(n1514) );
  NANDN U1564 ( .A(n19640), .B(n1514), .Z(n1415) );
  NAND U1565 ( .A(n1416), .B(n1415), .Z(n1483) );
  XNOR U1566 ( .A(n19714), .B(n2027), .Z(n1517) );
  NANDN U1567 ( .A(n1517), .B(n19766), .Z(n1419) );
  NANDN U1568 ( .A(n1417), .B(n19767), .Z(n1418) );
  NAND U1569 ( .A(n1419), .B(n1418), .Z(n1480) );
  NAND U1570 ( .A(n19554), .B(n1420), .Z(n1422) );
  IV U1571 ( .A(a[23]), .Z(n2366) );
  XNOR U1572 ( .A(b[3]), .B(n2366), .Z(n1520) );
  NANDN U1573 ( .A(n19521), .B(n1520), .Z(n1421) );
  AND U1574 ( .A(n1422), .B(n1421), .Z(n1481) );
  XNOR U1575 ( .A(n1480), .B(n1481), .Z(n1482) );
  XOR U1576 ( .A(n1483), .B(n1482), .Z(n1524) );
  XOR U1577 ( .A(n1523), .B(n1524), .Z(n1525) );
  XNOR U1578 ( .A(n1526), .B(n1525), .Z(n1474) );
  NAND U1579 ( .A(n1424), .B(n1423), .Z(n1428) );
  NAND U1580 ( .A(n1426), .B(n1425), .Z(n1427) );
  NAND U1581 ( .A(n1428), .B(n1427), .Z(n1475) );
  XOR U1582 ( .A(n1474), .B(n1475), .Z(n1477) );
  XNOR U1583 ( .A(n20052), .B(n1717), .Z(n1492) );
  OR U1584 ( .A(n1492), .B(n20020), .Z(n1431) );
  NANDN U1585 ( .A(n1429), .B(n19960), .Z(n1430) );
  NAND U1586 ( .A(n1431), .B(n1430), .Z(n1489) );
  XNOR U1587 ( .A(n102), .B(n1432), .Z(n1496) );
  OR U1588 ( .A(n1496), .B(n20121), .Z(n1435) );
  NANDN U1589 ( .A(n1433), .B(n20122), .Z(n1434) );
  NAND U1590 ( .A(n1435), .B(n1434), .Z(n1486) );
  XNOR U1591 ( .A(n19975), .B(n1871), .Z(n1499) );
  NANDN U1592 ( .A(n1499), .B(n19883), .Z(n1438) );
  NANDN U1593 ( .A(n1436), .B(n19937), .Z(n1437) );
  AND U1594 ( .A(n1438), .B(n1437), .Z(n1487) );
  XNOR U1595 ( .A(n1486), .B(n1487), .Z(n1488) );
  XNOR U1596 ( .A(n1489), .B(n1488), .Z(n1529) );
  NANDN U1597 ( .A(n1440), .B(n1439), .Z(n1444) );
  NAND U1598 ( .A(n1442), .B(n1441), .Z(n1443) );
  NAND U1599 ( .A(n1444), .B(n1443), .Z(n1530) );
  XNOR U1600 ( .A(n1529), .B(n1530), .Z(n1531) );
  NANDN U1601 ( .A(n1446), .B(n1445), .Z(n1450) );
  NAND U1602 ( .A(n1448), .B(n1447), .Z(n1449) );
  AND U1603 ( .A(n1450), .B(n1449), .Z(n1532) );
  XNOR U1604 ( .A(n1531), .B(n1532), .Z(n1476) );
  XNOR U1605 ( .A(n1477), .B(n1476), .Z(n1535) );
  NANDN U1606 ( .A(n1452), .B(n1451), .Z(n1456) );
  NAND U1607 ( .A(n1454), .B(n1453), .Z(n1455) );
  NAND U1608 ( .A(n1456), .B(n1455), .Z(n1536) );
  XNOR U1609 ( .A(n1535), .B(n1536), .Z(n1537) );
  XOR U1610 ( .A(n1538), .B(n1537), .Z(n1468) );
  NANDN U1611 ( .A(n1458), .B(n1457), .Z(n1462) );
  NANDN U1612 ( .A(n1460), .B(n1459), .Z(n1461) );
  NAND U1613 ( .A(n1462), .B(n1461), .Z(n1469) );
  XNOR U1614 ( .A(n1468), .B(n1469), .Z(n1470) );
  XNOR U1615 ( .A(n1471), .B(n1470), .Z(n1541) );
  XNOR U1616 ( .A(n1541), .B(sreg[265]), .Z(n1543) );
  NAND U1617 ( .A(n1463), .B(sreg[264]), .Z(n1467) );
  OR U1618 ( .A(n1465), .B(n1464), .Z(n1466) );
  AND U1619 ( .A(n1467), .B(n1466), .Z(n1542) );
  XOR U1620 ( .A(n1543), .B(n1542), .Z(c[265]) );
  NANDN U1621 ( .A(n1469), .B(n1468), .Z(n1473) );
  NAND U1622 ( .A(n1471), .B(n1470), .Z(n1472) );
  NAND U1623 ( .A(n1473), .B(n1472), .Z(n1549) );
  NANDN U1624 ( .A(n1475), .B(n1474), .Z(n1479) );
  OR U1625 ( .A(n1477), .B(n1476), .Z(n1478) );
  NAND U1626 ( .A(n1479), .B(n1478), .Z(n1616) );
  NANDN U1627 ( .A(n1481), .B(n1480), .Z(n1485) );
  NAND U1628 ( .A(n1483), .B(n1482), .Z(n1484) );
  NAND U1629 ( .A(n1485), .B(n1484), .Z(n1610) );
  NANDN U1630 ( .A(n1487), .B(n1486), .Z(n1491) );
  NAND U1631 ( .A(n1489), .B(n1488), .Z(n1490) );
  NAND U1632 ( .A(n1491), .B(n1490), .Z(n1607) );
  XNOR U1633 ( .A(n20052), .B(n1793), .Z(n1558) );
  OR U1634 ( .A(n1558), .B(n20020), .Z(n1494) );
  NANDN U1635 ( .A(n1492), .B(n19960), .Z(n1493) );
  NAND U1636 ( .A(n1494), .B(n1493), .Z(n1571) );
  XNOR U1637 ( .A(n102), .B(n1495), .Z(n1562) );
  OR U1638 ( .A(n1562), .B(n20121), .Z(n1498) );
  NANDN U1639 ( .A(n1496), .B(n20122), .Z(n1497) );
  NAND U1640 ( .A(n1498), .B(n1497), .Z(n1568) );
  XNOR U1641 ( .A(n19975), .B(n1976), .Z(n1565) );
  NANDN U1642 ( .A(n1565), .B(n19883), .Z(n1501) );
  NANDN U1643 ( .A(n1499), .B(n19937), .Z(n1500) );
  AND U1644 ( .A(n1501), .B(n1500), .Z(n1569) );
  XNOR U1645 ( .A(n1568), .B(n1569), .Z(n1570) );
  XNOR U1646 ( .A(n1571), .B(n1570), .Z(n1608) );
  XNOR U1647 ( .A(n1607), .B(n1608), .Z(n1609) );
  XNOR U1648 ( .A(n1610), .B(n1609), .Z(n1555) );
  NANDN U1649 ( .A(n1503), .B(n1502), .Z(n1507) );
  OR U1650 ( .A(n1505), .B(n1504), .Z(n1506) );
  NAND U1651 ( .A(n1507), .B(n1506), .Z(n1604) );
  NAND U1652 ( .A(b[0]), .B(a[26]), .Z(n1508) );
  XNOR U1653 ( .A(b[1]), .B(n1508), .Z(n1510) );
  NAND U1654 ( .A(a[25]), .B(n98), .Z(n1509) );
  AND U1655 ( .A(n1510), .B(n1509), .Z(n1580) );
  XNOR U1656 ( .A(n20154), .B(n1639), .Z(n1589) );
  OR U1657 ( .A(n1589), .B(n20057), .Z(n1513) );
  NANDN U1658 ( .A(n1511), .B(n20098), .Z(n1512) );
  AND U1659 ( .A(n1513), .B(n1512), .Z(n1581) );
  XOR U1660 ( .A(n1580), .B(n1581), .Z(n1583) );
  NAND U1661 ( .A(a[10]), .B(b[15]), .Z(n1582) );
  XOR U1662 ( .A(n1583), .B(n1582), .Z(n1601) );
  NAND U1663 ( .A(n19722), .B(n1514), .Z(n1516) );
  XNOR U1664 ( .A(b[5]), .B(n2261), .Z(n1592) );
  NANDN U1665 ( .A(n19640), .B(n1592), .Z(n1515) );
  NAND U1666 ( .A(n1516), .B(n1515), .Z(n1577) );
  XNOR U1667 ( .A(n19714), .B(n2105), .Z(n1595) );
  NANDN U1668 ( .A(n1595), .B(n19766), .Z(n1519) );
  NANDN U1669 ( .A(n1517), .B(n19767), .Z(n1518) );
  NAND U1670 ( .A(n1519), .B(n1518), .Z(n1574) );
  NAND U1671 ( .A(n19554), .B(n1520), .Z(n1522) );
  IV U1672 ( .A(a[24]), .Z(n2417) );
  XNOR U1673 ( .A(b[3]), .B(n2417), .Z(n1598) );
  NANDN U1674 ( .A(n19521), .B(n1598), .Z(n1521) );
  AND U1675 ( .A(n1522), .B(n1521), .Z(n1575) );
  XNOR U1676 ( .A(n1574), .B(n1575), .Z(n1576) );
  XOR U1677 ( .A(n1577), .B(n1576), .Z(n1602) );
  XOR U1678 ( .A(n1601), .B(n1602), .Z(n1603) );
  XNOR U1679 ( .A(n1604), .B(n1603), .Z(n1552) );
  NAND U1680 ( .A(n1524), .B(n1523), .Z(n1528) );
  NAND U1681 ( .A(n1526), .B(n1525), .Z(n1527) );
  NAND U1682 ( .A(n1528), .B(n1527), .Z(n1553) );
  XNOR U1683 ( .A(n1552), .B(n1553), .Z(n1554) );
  XOR U1684 ( .A(n1555), .B(n1554), .Z(n1613) );
  NANDN U1685 ( .A(n1530), .B(n1529), .Z(n1534) );
  NAND U1686 ( .A(n1532), .B(n1531), .Z(n1533) );
  NAND U1687 ( .A(n1534), .B(n1533), .Z(n1614) );
  XOR U1688 ( .A(n1613), .B(n1614), .Z(n1615) );
  XOR U1689 ( .A(n1616), .B(n1615), .Z(n1546) );
  NANDN U1690 ( .A(n1536), .B(n1535), .Z(n1540) );
  NANDN U1691 ( .A(n1538), .B(n1537), .Z(n1539) );
  NAND U1692 ( .A(n1540), .B(n1539), .Z(n1547) );
  XNOR U1693 ( .A(n1546), .B(n1547), .Z(n1548) );
  XNOR U1694 ( .A(n1549), .B(n1548), .Z(n1619) );
  XNOR U1695 ( .A(n1619), .B(sreg[266]), .Z(n1621) );
  NAND U1696 ( .A(n1541), .B(sreg[265]), .Z(n1545) );
  OR U1697 ( .A(n1543), .B(n1542), .Z(n1544) );
  AND U1698 ( .A(n1545), .B(n1544), .Z(n1620) );
  XOR U1699 ( .A(n1621), .B(n1620), .Z(c[266]) );
  NANDN U1700 ( .A(n1547), .B(n1546), .Z(n1551) );
  NAND U1701 ( .A(n1549), .B(n1548), .Z(n1550) );
  NAND U1702 ( .A(n1551), .B(n1550), .Z(n1627) );
  NANDN U1703 ( .A(n1553), .B(n1552), .Z(n1557) );
  NAND U1704 ( .A(n1555), .B(n1554), .Z(n1556) );
  NAND U1705 ( .A(n1557), .B(n1556), .Z(n1694) );
  XNOR U1706 ( .A(n20052), .B(n1871), .Z(n1636) );
  OR U1707 ( .A(n1636), .B(n20020), .Z(n1560) );
  NANDN U1708 ( .A(n1558), .B(n19960), .Z(n1559) );
  NAND U1709 ( .A(n1560), .B(n1559), .Z(n1649) );
  XNOR U1710 ( .A(n102), .B(n1561), .Z(n1640) );
  OR U1711 ( .A(n1640), .B(n20121), .Z(n1564) );
  NANDN U1712 ( .A(n1562), .B(n20122), .Z(n1563) );
  NAND U1713 ( .A(n1564), .B(n1563), .Z(n1646) );
  XNOR U1714 ( .A(n19975), .B(n2027), .Z(n1643) );
  NANDN U1715 ( .A(n1643), .B(n19883), .Z(n1567) );
  NANDN U1716 ( .A(n1565), .B(n19937), .Z(n1566) );
  AND U1717 ( .A(n1567), .B(n1566), .Z(n1647) );
  XNOR U1718 ( .A(n1646), .B(n1647), .Z(n1648) );
  XNOR U1719 ( .A(n1649), .B(n1648), .Z(n1685) );
  NANDN U1720 ( .A(n1569), .B(n1568), .Z(n1573) );
  NAND U1721 ( .A(n1571), .B(n1570), .Z(n1572) );
  NAND U1722 ( .A(n1573), .B(n1572), .Z(n1686) );
  XNOR U1723 ( .A(n1685), .B(n1686), .Z(n1687) );
  NANDN U1724 ( .A(n1575), .B(n1574), .Z(n1579) );
  NAND U1725 ( .A(n1577), .B(n1576), .Z(n1578) );
  AND U1726 ( .A(n1579), .B(n1578), .Z(n1688) );
  XNOR U1727 ( .A(n1687), .B(n1688), .Z(n1632) );
  NANDN U1728 ( .A(n1581), .B(n1580), .Z(n1585) );
  OR U1729 ( .A(n1583), .B(n1582), .Z(n1584) );
  NAND U1730 ( .A(n1585), .B(n1584), .Z(n1682) );
  NAND U1731 ( .A(b[0]), .B(a[27]), .Z(n1586) );
  XNOR U1732 ( .A(b[1]), .B(n1586), .Z(n1588) );
  NAND U1733 ( .A(a[26]), .B(n98), .Z(n1587) );
  AND U1734 ( .A(n1588), .B(n1587), .Z(n1658) );
  XNOR U1735 ( .A(n20154), .B(n1717), .Z(n1664) );
  OR U1736 ( .A(n1664), .B(n20057), .Z(n1591) );
  NANDN U1737 ( .A(n1589), .B(n20098), .Z(n1590) );
  AND U1738 ( .A(n1591), .B(n1590), .Z(n1659) );
  XOR U1739 ( .A(n1658), .B(n1659), .Z(n1661) );
  NAND U1740 ( .A(a[11]), .B(b[15]), .Z(n1660) );
  XOR U1741 ( .A(n1661), .B(n1660), .Z(n1679) );
  NAND U1742 ( .A(n19722), .B(n1592), .Z(n1594) );
  XNOR U1743 ( .A(b[5]), .B(n2366), .Z(n1670) );
  NANDN U1744 ( .A(n19640), .B(n1670), .Z(n1593) );
  NAND U1745 ( .A(n1594), .B(n1593), .Z(n1655) );
  XNOR U1746 ( .A(n19714), .B(n2195), .Z(n1673) );
  NANDN U1747 ( .A(n1673), .B(n19766), .Z(n1597) );
  NANDN U1748 ( .A(n1595), .B(n19767), .Z(n1596) );
  NAND U1749 ( .A(n1597), .B(n1596), .Z(n1652) );
  NAND U1750 ( .A(n19554), .B(n1598), .Z(n1600) );
  IV U1751 ( .A(a[25]), .Z(n2495) );
  XNOR U1752 ( .A(b[3]), .B(n2495), .Z(n1676) );
  NANDN U1753 ( .A(n19521), .B(n1676), .Z(n1599) );
  AND U1754 ( .A(n1600), .B(n1599), .Z(n1653) );
  XNOR U1755 ( .A(n1652), .B(n1653), .Z(n1654) );
  XOR U1756 ( .A(n1655), .B(n1654), .Z(n1680) );
  XOR U1757 ( .A(n1679), .B(n1680), .Z(n1681) );
  XNOR U1758 ( .A(n1682), .B(n1681), .Z(n1630) );
  NAND U1759 ( .A(n1602), .B(n1601), .Z(n1606) );
  NAND U1760 ( .A(n1604), .B(n1603), .Z(n1605) );
  NAND U1761 ( .A(n1606), .B(n1605), .Z(n1631) );
  XOR U1762 ( .A(n1630), .B(n1631), .Z(n1633) );
  XNOR U1763 ( .A(n1632), .B(n1633), .Z(n1691) );
  NANDN U1764 ( .A(n1608), .B(n1607), .Z(n1612) );
  NAND U1765 ( .A(n1610), .B(n1609), .Z(n1611) );
  AND U1766 ( .A(n1612), .B(n1611), .Z(n1692) );
  XNOR U1767 ( .A(n1691), .B(n1692), .Z(n1693) );
  XOR U1768 ( .A(n1694), .B(n1693), .Z(n1624) );
  OR U1769 ( .A(n1614), .B(n1613), .Z(n1618) );
  NANDN U1770 ( .A(n1616), .B(n1615), .Z(n1617) );
  NAND U1771 ( .A(n1618), .B(n1617), .Z(n1625) );
  XNOR U1772 ( .A(n1624), .B(n1625), .Z(n1626) );
  XNOR U1773 ( .A(n1627), .B(n1626), .Z(n1697) );
  XNOR U1774 ( .A(n1697), .B(sreg[267]), .Z(n1699) );
  NAND U1775 ( .A(n1619), .B(sreg[266]), .Z(n1623) );
  OR U1776 ( .A(n1621), .B(n1620), .Z(n1622) );
  AND U1777 ( .A(n1623), .B(n1622), .Z(n1698) );
  XOR U1778 ( .A(n1699), .B(n1698), .Z(c[267]) );
  NANDN U1779 ( .A(n1625), .B(n1624), .Z(n1629) );
  NAND U1780 ( .A(n1627), .B(n1626), .Z(n1628) );
  NAND U1781 ( .A(n1629), .B(n1628), .Z(n1705) );
  NANDN U1782 ( .A(n1631), .B(n1630), .Z(n1635) );
  OR U1783 ( .A(n1633), .B(n1632), .Z(n1634) );
  NAND U1784 ( .A(n1635), .B(n1634), .Z(n1770) );
  XNOR U1785 ( .A(n20052), .B(n1976), .Z(n1714) );
  OR U1786 ( .A(n1714), .B(n20020), .Z(n1638) );
  NANDN U1787 ( .A(n1636), .B(n19960), .Z(n1637) );
  NAND U1788 ( .A(n1638), .B(n1637), .Z(n1727) );
  XNOR U1789 ( .A(n102), .B(n1639), .Z(n1718) );
  OR U1790 ( .A(n1718), .B(n20121), .Z(n1642) );
  NANDN U1791 ( .A(n1640), .B(n20122), .Z(n1641) );
  NAND U1792 ( .A(n1642), .B(n1641), .Z(n1724) );
  XNOR U1793 ( .A(n19975), .B(n2105), .Z(n1721) );
  NANDN U1794 ( .A(n1721), .B(n19883), .Z(n1645) );
  NANDN U1795 ( .A(n1643), .B(n19937), .Z(n1644) );
  AND U1796 ( .A(n1645), .B(n1644), .Z(n1725) );
  XNOR U1797 ( .A(n1724), .B(n1725), .Z(n1726) );
  XNOR U1798 ( .A(n1727), .B(n1726), .Z(n1761) );
  NANDN U1799 ( .A(n1647), .B(n1646), .Z(n1651) );
  NAND U1800 ( .A(n1649), .B(n1648), .Z(n1650) );
  NAND U1801 ( .A(n1651), .B(n1650), .Z(n1762) );
  XNOR U1802 ( .A(n1761), .B(n1762), .Z(n1763) );
  NANDN U1803 ( .A(n1653), .B(n1652), .Z(n1657) );
  NAND U1804 ( .A(n1655), .B(n1654), .Z(n1656) );
  AND U1805 ( .A(n1657), .B(n1656), .Z(n1764) );
  XNOR U1806 ( .A(n1763), .B(n1764), .Z(n1710) );
  NANDN U1807 ( .A(n1659), .B(n1658), .Z(n1663) );
  OR U1808 ( .A(n1661), .B(n1660), .Z(n1662) );
  NAND U1809 ( .A(n1663), .B(n1662), .Z(n1760) );
  XNOR U1810 ( .A(n20154), .B(n1793), .Z(n1745) );
  OR U1811 ( .A(n1745), .B(n20057), .Z(n1666) );
  NANDN U1812 ( .A(n1664), .B(n20098), .Z(n1665) );
  NAND U1813 ( .A(n1666), .B(n1665), .Z(n1736) );
  AND U1814 ( .A(a[28]), .B(b[0]), .Z(n1667) );
  XOR U1815 ( .A(b[1]), .B(n1667), .Z(n1669) );
  NAND U1816 ( .A(a[27]), .B(n98), .Z(n1668) );
  NAND U1817 ( .A(n1669), .B(n1668), .Z(n1737) );
  XNOR U1818 ( .A(n1736), .B(n1737), .Z(n1738) );
  NAND U1819 ( .A(a[12]), .B(b[15]), .Z(n1739) );
  XOR U1820 ( .A(n1738), .B(n1739), .Z(n1757) );
  NAND U1821 ( .A(n19722), .B(n1670), .Z(n1672) );
  XNOR U1822 ( .A(b[5]), .B(n2417), .Z(n1748) );
  NANDN U1823 ( .A(n19640), .B(n1748), .Z(n1671) );
  NAND U1824 ( .A(n1672), .B(n1671), .Z(n1733) );
  XNOR U1825 ( .A(n19714), .B(n2261), .Z(n1751) );
  NANDN U1826 ( .A(n1751), .B(n19766), .Z(n1675) );
  NANDN U1827 ( .A(n1673), .B(n19767), .Z(n1674) );
  NAND U1828 ( .A(n1675), .B(n1674), .Z(n1730) );
  NAND U1829 ( .A(n19554), .B(n1676), .Z(n1678) );
  IV U1830 ( .A(a[26]), .Z(n2600) );
  XNOR U1831 ( .A(b[3]), .B(n2600), .Z(n1754) );
  NANDN U1832 ( .A(n19521), .B(n1754), .Z(n1677) );
  AND U1833 ( .A(n1678), .B(n1677), .Z(n1731) );
  XNOR U1834 ( .A(n1730), .B(n1731), .Z(n1732) );
  XOR U1835 ( .A(n1733), .B(n1732), .Z(n1758) );
  XNOR U1836 ( .A(n1757), .B(n1758), .Z(n1759) );
  XNOR U1837 ( .A(n1760), .B(n1759), .Z(n1708) );
  NAND U1838 ( .A(n1680), .B(n1679), .Z(n1684) );
  NAND U1839 ( .A(n1682), .B(n1681), .Z(n1683) );
  NAND U1840 ( .A(n1684), .B(n1683), .Z(n1709) );
  XOR U1841 ( .A(n1708), .B(n1709), .Z(n1711) );
  XNOR U1842 ( .A(n1710), .B(n1711), .Z(n1767) );
  NANDN U1843 ( .A(n1686), .B(n1685), .Z(n1690) );
  NAND U1844 ( .A(n1688), .B(n1687), .Z(n1689) );
  NAND U1845 ( .A(n1690), .B(n1689), .Z(n1768) );
  XNOR U1846 ( .A(n1767), .B(n1768), .Z(n1769) );
  XOR U1847 ( .A(n1770), .B(n1769), .Z(n1702) );
  NANDN U1848 ( .A(n1692), .B(n1691), .Z(n1696) );
  NANDN U1849 ( .A(n1694), .B(n1693), .Z(n1695) );
  NAND U1850 ( .A(n1696), .B(n1695), .Z(n1703) );
  XNOR U1851 ( .A(n1702), .B(n1703), .Z(n1704) );
  XNOR U1852 ( .A(n1705), .B(n1704), .Z(n1773) );
  XNOR U1853 ( .A(n1773), .B(sreg[268]), .Z(n1775) );
  NAND U1854 ( .A(n1697), .B(sreg[267]), .Z(n1701) );
  OR U1855 ( .A(n1699), .B(n1698), .Z(n1700) );
  AND U1856 ( .A(n1701), .B(n1700), .Z(n1774) );
  XOR U1857 ( .A(n1775), .B(n1774), .Z(c[268]) );
  NANDN U1858 ( .A(n1703), .B(n1702), .Z(n1707) );
  NAND U1859 ( .A(n1705), .B(n1704), .Z(n1706) );
  NAND U1860 ( .A(n1707), .B(n1706), .Z(n1781) );
  NANDN U1861 ( .A(n1709), .B(n1708), .Z(n1713) );
  OR U1862 ( .A(n1711), .B(n1710), .Z(n1712) );
  NAND U1863 ( .A(n1713), .B(n1712), .Z(n1848) );
  XNOR U1864 ( .A(n20052), .B(n2027), .Z(n1790) );
  OR U1865 ( .A(n1790), .B(n20020), .Z(n1716) );
  NANDN U1866 ( .A(n1714), .B(n19960), .Z(n1715) );
  NAND U1867 ( .A(n1716), .B(n1715), .Z(n1803) );
  XNOR U1868 ( .A(n102), .B(n1717), .Z(n1794) );
  OR U1869 ( .A(n1794), .B(n20121), .Z(n1720) );
  NANDN U1870 ( .A(n1718), .B(n20122), .Z(n1719) );
  NAND U1871 ( .A(n1720), .B(n1719), .Z(n1800) );
  XNOR U1872 ( .A(n19975), .B(n2195), .Z(n1797) );
  NANDN U1873 ( .A(n1797), .B(n19883), .Z(n1723) );
  NANDN U1874 ( .A(n1721), .B(n19937), .Z(n1722) );
  AND U1875 ( .A(n1723), .B(n1722), .Z(n1801) );
  XNOR U1876 ( .A(n1800), .B(n1801), .Z(n1802) );
  XNOR U1877 ( .A(n1803), .B(n1802), .Z(n1839) );
  NANDN U1878 ( .A(n1725), .B(n1724), .Z(n1729) );
  NAND U1879 ( .A(n1727), .B(n1726), .Z(n1728) );
  NAND U1880 ( .A(n1729), .B(n1728), .Z(n1840) );
  XNOR U1881 ( .A(n1839), .B(n1840), .Z(n1841) );
  NANDN U1882 ( .A(n1731), .B(n1730), .Z(n1735) );
  NAND U1883 ( .A(n1733), .B(n1732), .Z(n1734) );
  AND U1884 ( .A(n1735), .B(n1734), .Z(n1842) );
  XNOR U1885 ( .A(n1841), .B(n1842), .Z(n1786) );
  NANDN U1886 ( .A(n1737), .B(n1736), .Z(n1741) );
  NANDN U1887 ( .A(n1739), .B(n1738), .Z(n1740) );
  NAND U1888 ( .A(n1741), .B(n1740), .Z(n1836) );
  NAND U1889 ( .A(b[0]), .B(a[29]), .Z(n1742) );
  XNOR U1890 ( .A(b[1]), .B(n1742), .Z(n1744) );
  NAND U1891 ( .A(a[28]), .B(n98), .Z(n1743) );
  AND U1892 ( .A(n1744), .B(n1743), .Z(n1812) );
  XNOR U1893 ( .A(n20154), .B(n1871), .Z(n1821) );
  OR U1894 ( .A(n1821), .B(n20057), .Z(n1747) );
  NANDN U1895 ( .A(n1745), .B(n20098), .Z(n1746) );
  AND U1896 ( .A(n1747), .B(n1746), .Z(n1813) );
  XOR U1897 ( .A(n1812), .B(n1813), .Z(n1815) );
  NAND U1898 ( .A(a[13]), .B(b[15]), .Z(n1814) );
  XOR U1899 ( .A(n1815), .B(n1814), .Z(n1833) );
  NAND U1900 ( .A(n19722), .B(n1748), .Z(n1750) );
  XNOR U1901 ( .A(b[5]), .B(n2495), .Z(n1824) );
  NANDN U1902 ( .A(n19640), .B(n1824), .Z(n1749) );
  NAND U1903 ( .A(n1750), .B(n1749), .Z(n1809) );
  XNOR U1904 ( .A(n19714), .B(n2366), .Z(n1827) );
  NANDN U1905 ( .A(n1827), .B(n19766), .Z(n1753) );
  NANDN U1906 ( .A(n1751), .B(n19767), .Z(n1752) );
  NAND U1907 ( .A(n1753), .B(n1752), .Z(n1806) );
  NAND U1908 ( .A(n19554), .B(n1754), .Z(n1756) );
  IV U1909 ( .A(a[27]), .Z(n2651) );
  XNOR U1910 ( .A(b[3]), .B(n2651), .Z(n1830) );
  NANDN U1911 ( .A(n19521), .B(n1830), .Z(n1755) );
  AND U1912 ( .A(n1756), .B(n1755), .Z(n1807) );
  XNOR U1913 ( .A(n1806), .B(n1807), .Z(n1808) );
  XOR U1914 ( .A(n1809), .B(n1808), .Z(n1834) );
  XOR U1915 ( .A(n1833), .B(n1834), .Z(n1835) );
  XNOR U1916 ( .A(n1836), .B(n1835), .Z(n1784) );
  XOR U1917 ( .A(n1784), .B(n1785), .Z(n1787) );
  XNOR U1918 ( .A(n1786), .B(n1787), .Z(n1845) );
  NANDN U1919 ( .A(n1762), .B(n1761), .Z(n1766) );
  NAND U1920 ( .A(n1764), .B(n1763), .Z(n1765) );
  NAND U1921 ( .A(n1766), .B(n1765), .Z(n1846) );
  XNOR U1922 ( .A(n1845), .B(n1846), .Z(n1847) );
  XOR U1923 ( .A(n1848), .B(n1847), .Z(n1778) );
  NANDN U1924 ( .A(n1768), .B(n1767), .Z(n1772) );
  NANDN U1925 ( .A(n1770), .B(n1769), .Z(n1771) );
  NAND U1926 ( .A(n1772), .B(n1771), .Z(n1779) );
  XNOR U1927 ( .A(n1778), .B(n1779), .Z(n1780) );
  XNOR U1928 ( .A(n1781), .B(n1780), .Z(n1851) );
  XNOR U1929 ( .A(n1851), .B(sreg[269]), .Z(n1853) );
  NAND U1930 ( .A(n1773), .B(sreg[268]), .Z(n1777) );
  OR U1931 ( .A(n1775), .B(n1774), .Z(n1776) );
  AND U1932 ( .A(n1777), .B(n1776), .Z(n1852) );
  XOR U1933 ( .A(n1853), .B(n1852), .Z(c[269]) );
  NANDN U1934 ( .A(n1779), .B(n1778), .Z(n1783) );
  NAND U1935 ( .A(n1781), .B(n1780), .Z(n1782) );
  NAND U1936 ( .A(n1783), .B(n1782), .Z(n1859) );
  NANDN U1937 ( .A(n1785), .B(n1784), .Z(n1789) );
  OR U1938 ( .A(n1787), .B(n1786), .Z(n1788) );
  NAND U1939 ( .A(n1789), .B(n1788), .Z(n1926) );
  XNOR U1940 ( .A(n20052), .B(n2105), .Z(n1868) );
  OR U1941 ( .A(n1868), .B(n20020), .Z(n1792) );
  NANDN U1942 ( .A(n1790), .B(n19960), .Z(n1791) );
  NAND U1943 ( .A(n1792), .B(n1791), .Z(n1881) );
  XNOR U1944 ( .A(n102), .B(n1793), .Z(n1872) );
  OR U1945 ( .A(n1872), .B(n20121), .Z(n1796) );
  NANDN U1946 ( .A(n1794), .B(n20122), .Z(n1795) );
  NAND U1947 ( .A(n1796), .B(n1795), .Z(n1878) );
  XNOR U1948 ( .A(n19975), .B(n2261), .Z(n1875) );
  NANDN U1949 ( .A(n1875), .B(n19883), .Z(n1799) );
  NANDN U1950 ( .A(n1797), .B(n19937), .Z(n1798) );
  AND U1951 ( .A(n1799), .B(n1798), .Z(n1879) );
  XNOR U1952 ( .A(n1878), .B(n1879), .Z(n1880) );
  XNOR U1953 ( .A(n1881), .B(n1880), .Z(n1917) );
  NANDN U1954 ( .A(n1801), .B(n1800), .Z(n1805) );
  NAND U1955 ( .A(n1803), .B(n1802), .Z(n1804) );
  NAND U1956 ( .A(n1805), .B(n1804), .Z(n1918) );
  XNOR U1957 ( .A(n1917), .B(n1918), .Z(n1919) );
  NANDN U1958 ( .A(n1807), .B(n1806), .Z(n1811) );
  NAND U1959 ( .A(n1809), .B(n1808), .Z(n1810) );
  AND U1960 ( .A(n1811), .B(n1810), .Z(n1920) );
  XNOR U1961 ( .A(n1919), .B(n1920), .Z(n1864) );
  NANDN U1962 ( .A(n1813), .B(n1812), .Z(n1817) );
  OR U1963 ( .A(n1815), .B(n1814), .Z(n1816) );
  NAND U1964 ( .A(n1817), .B(n1816), .Z(n1914) );
  NAND U1965 ( .A(b[0]), .B(a[30]), .Z(n1818) );
  XNOR U1966 ( .A(b[1]), .B(n1818), .Z(n1820) );
  NAND U1967 ( .A(a[29]), .B(n98), .Z(n1819) );
  AND U1968 ( .A(n1820), .B(n1819), .Z(n1890) );
  XNOR U1969 ( .A(n20154), .B(n1976), .Z(n1899) );
  OR U1970 ( .A(n1899), .B(n20057), .Z(n1823) );
  NANDN U1971 ( .A(n1821), .B(n20098), .Z(n1822) );
  AND U1972 ( .A(n1823), .B(n1822), .Z(n1891) );
  XOR U1973 ( .A(n1890), .B(n1891), .Z(n1893) );
  NAND U1974 ( .A(a[14]), .B(b[15]), .Z(n1892) );
  XOR U1975 ( .A(n1893), .B(n1892), .Z(n1911) );
  NAND U1976 ( .A(n19722), .B(n1824), .Z(n1826) );
  XNOR U1977 ( .A(b[5]), .B(n2600), .Z(n1902) );
  NANDN U1978 ( .A(n19640), .B(n1902), .Z(n1825) );
  NAND U1979 ( .A(n1826), .B(n1825), .Z(n1887) );
  XNOR U1980 ( .A(n19714), .B(n2417), .Z(n1905) );
  NANDN U1981 ( .A(n1905), .B(n19766), .Z(n1829) );
  NANDN U1982 ( .A(n1827), .B(n19767), .Z(n1828) );
  NAND U1983 ( .A(n1829), .B(n1828), .Z(n1884) );
  NAND U1984 ( .A(n19554), .B(n1830), .Z(n1832) );
  IV U1985 ( .A(a[28]), .Z(n2729) );
  XNOR U1986 ( .A(b[3]), .B(n2729), .Z(n1908) );
  NANDN U1987 ( .A(n19521), .B(n1908), .Z(n1831) );
  AND U1988 ( .A(n1832), .B(n1831), .Z(n1885) );
  XNOR U1989 ( .A(n1884), .B(n1885), .Z(n1886) );
  XOR U1990 ( .A(n1887), .B(n1886), .Z(n1912) );
  XOR U1991 ( .A(n1911), .B(n1912), .Z(n1913) );
  XNOR U1992 ( .A(n1914), .B(n1913), .Z(n1862) );
  NAND U1993 ( .A(n1834), .B(n1833), .Z(n1838) );
  NAND U1994 ( .A(n1836), .B(n1835), .Z(n1837) );
  NAND U1995 ( .A(n1838), .B(n1837), .Z(n1863) );
  XOR U1996 ( .A(n1862), .B(n1863), .Z(n1865) );
  XNOR U1997 ( .A(n1864), .B(n1865), .Z(n1923) );
  NANDN U1998 ( .A(n1840), .B(n1839), .Z(n1844) );
  NAND U1999 ( .A(n1842), .B(n1841), .Z(n1843) );
  NAND U2000 ( .A(n1844), .B(n1843), .Z(n1924) );
  XNOR U2001 ( .A(n1923), .B(n1924), .Z(n1925) );
  XOR U2002 ( .A(n1926), .B(n1925), .Z(n1856) );
  NANDN U2003 ( .A(n1846), .B(n1845), .Z(n1850) );
  NANDN U2004 ( .A(n1848), .B(n1847), .Z(n1849) );
  NAND U2005 ( .A(n1850), .B(n1849), .Z(n1857) );
  XNOR U2006 ( .A(n1856), .B(n1857), .Z(n1858) );
  XNOR U2007 ( .A(n1859), .B(n1858), .Z(n1929) );
  XNOR U2008 ( .A(n1929), .B(sreg[270]), .Z(n1931) );
  NAND U2009 ( .A(n1851), .B(sreg[269]), .Z(n1855) );
  OR U2010 ( .A(n1853), .B(n1852), .Z(n1854) );
  AND U2011 ( .A(n1855), .B(n1854), .Z(n1930) );
  XOR U2012 ( .A(n1931), .B(n1930), .Z(c[270]) );
  NANDN U2013 ( .A(n1857), .B(n1856), .Z(n1861) );
  NAND U2014 ( .A(n1859), .B(n1858), .Z(n1860) );
  NAND U2015 ( .A(n1861), .B(n1860), .Z(n1937) );
  NANDN U2016 ( .A(n1863), .B(n1862), .Z(n1867) );
  OR U2017 ( .A(n1865), .B(n1864), .Z(n1866) );
  NAND U2018 ( .A(n1867), .B(n1866), .Z(n2004) );
  XNOR U2019 ( .A(n20052), .B(n2195), .Z(n1973) );
  OR U2020 ( .A(n1973), .B(n20020), .Z(n1870) );
  NANDN U2021 ( .A(n1868), .B(n19960), .Z(n1869) );
  NAND U2022 ( .A(n1870), .B(n1869), .Z(n1986) );
  XNOR U2023 ( .A(n102), .B(n1871), .Z(n1977) );
  OR U2024 ( .A(n1977), .B(n20121), .Z(n1874) );
  NANDN U2025 ( .A(n1872), .B(n20122), .Z(n1873) );
  NAND U2026 ( .A(n1874), .B(n1873), .Z(n1983) );
  XNOR U2027 ( .A(n19975), .B(n2366), .Z(n1980) );
  NANDN U2028 ( .A(n1980), .B(n19883), .Z(n1877) );
  NANDN U2029 ( .A(n1875), .B(n19937), .Z(n1876) );
  AND U2030 ( .A(n1877), .B(n1876), .Z(n1984) );
  XNOR U2031 ( .A(n1983), .B(n1984), .Z(n1985) );
  XNOR U2032 ( .A(n1986), .B(n1985), .Z(n1995) );
  NANDN U2033 ( .A(n1879), .B(n1878), .Z(n1883) );
  NAND U2034 ( .A(n1881), .B(n1880), .Z(n1882) );
  NAND U2035 ( .A(n1883), .B(n1882), .Z(n1996) );
  XNOR U2036 ( .A(n1995), .B(n1996), .Z(n1997) );
  NANDN U2037 ( .A(n1885), .B(n1884), .Z(n1889) );
  NAND U2038 ( .A(n1887), .B(n1886), .Z(n1888) );
  AND U2039 ( .A(n1889), .B(n1888), .Z(n1998) );
  XNOR U2040 ( .A(n1997), .B(n1998), .Z(n1942) );
  NANDN U2041 ( .A(n1891), .B(n1890), .Z(n1895) );
  OR U2042 ( .A(n1893), .B(n1892), .Z(n1894) );
  NAND U2043 ( .A(n1895), .B(n1894), .Z(n1970) );
  NAND U2044 ( .A(b[0]), .B(a[31]), .Z(n1896) );
  XNOR U2045 ( .A(b[1]), .B(n1896), .Z(n1898) );
  NAND U2046 ( .A(a[30]), .B(n98), .Z(n1897) );
  AND U2047 ( .A(n1898), .B(n1897), .Z(n1946) );
  XNOR U2048 ( .A(n20154), .B(n2027), .Z(n1955) );
  OR U2049 ( .A(n1955), .B(n20057), .Z(n1901) );
  NANDN U2050 ( .A(n1899), .B(n20098), .Z(n1900) );
  AND U2051 ( .A(n1901), .B(n1900), .Z(n1947) );
  XOR U2052 ( .A(n1946), .B(n1947), .Z(n1949) );
  NAND U2053 ( .A(a[15]), .B(b[15]), .Z(n1948) );
  XOR U2054 ( .A(n1949), .B(n1948), .Z(n1967) );
  NAND U2055 ( .A(n19722), .B(n1902), .Z(n1904) );
  XNOR U2056 ( .A(b[5]), .B(n2651), .Z(n1958) );
  NANDN U2057 ( .A(n19640), .B(n1958), .Z(n1903) );
  NAND U2058 ( .A(n1904), .B(n1903), .Z(n1992) );
  XNOR U2059 ( .A(n19714), .B(n2495), .Z(n1961) );
  NANDN U2060 ( .A(n1961), .B(n19766), .Z(n1907) );
  NANDN U2061 ( .A(n1905), .B(n19767), .Z(n1906) );
  NAND U2062 ( .A(n1907), .B(n1906), .Z(n1989) );
  NAND U2063 ( .A(n19554), .B(n1908), .Z(n1910) );
  IV U2064 ( .A(a[29]), .Z(n2807) );
  XNOR U2065 ( .A(b[3]), .B(n2807), .Z(n1964) );
  NANDN U2066 ( .A(n19521), .B(n1964), .Z(n1909) );
  AND U2067 ( .A(n1910), .B(n1909), .Z(n1990) );
  XNOR U2068 ( .A(n1989), .B(n1990), .Z(n1991) );
  XOR U2069 ( .A(n1992), .B(n1991), .Z(n1968) );
  XOR U2070 ( .A(n1967), .B(n1968), .Z(n1969) );
  XNOR U2071 ( .A(n1970), .B(n1969), .Z(n1940) );
  NAND U2072 ( .A(n1912), .B(n1911), .Z(n1916) );
  NAND U2073 ( .A(n1914), .B(n1913), .Z(n1915) );
  NAND U2074 ( .A(n1916), .B(n1915), .Z(n1941) );
  XOR U2075 ( .A(n1940), .B(n1941), .Z(n1943) );
  XNOR U2076 ( .A(n1942), .B(n1943), .Z(n2001) );
  NANDN U2077 ( .A(n1918), .B(n1917), .Z(n1922) );
  NAND U2078 ( .A(n1920), .B(n1919), .Z(n1921) );
  NAND U2079 ( .A(n1922), .B(n1921), .Z(n2002) );
  XNOR U2080 ( .A(n2001), .B(n2002), .Z(n2003) );
  XOR U2081 ( .A(n2004), .B(n2003), .Z(n1934) );
  NANDN U2082 ( .A(n1924), .B(n1923), .Z(n1928) );
  NANDN U2083 ( .A(n1926), .B(n1925), .Z(n1927) );
  NAND U2084 ( .A(n1928), .B(n1927), .Z(n1935) );
  XNOR U2085 ( .A(n1934), .B(n1935), .Z(n1936) );
  XNOR U2086 ( .A(n1937), .B(n1936), .Z(n2007) );
  XNOR U2087 ( .A(n2007), .B(sreg[271]), .Z(n2009) );
  NAND U2088 ( .A(n1929), .B(sreg[270]), .Z(n1933) );
  OR U2089 ( .A(n1931), .B(n1930), .Z(n1932) );
  AND U2090 ( .A(n1933), .B(n1932), .Z(n2008) );
  XOR U2091 ( .A(n2009), .B(n2008), .Z(c[271]) );
  NANDN U2092 ( .A(n1935), .B(n1934), .Z(n1939) );
  NAND U2093 ( .A(n1937), .B(n1936), .Z(n1938) );
  NAND U2094 ( .A(n1939), .B(n1938), .Z(n2015) );
  NANDN U2095 ( .A(n1941), .B(n1940), .Z(n1945) );
  OR U2096 ( .A(n1943), .B(n1942), .Z(n1944) );
  NAND U2097 ( .A(n1945), .B(n1944), .Z(n2082) );
  NANDN U2098 ( .A(n1947), .B(n1946), .Z(n1951) );
  OR U2099 ( .A(n1949), .B(n1948), .Z(n1950) );
  NAND U2100 ( .A(n1951), .B(n1950), .Z(n2070) );
  NAND U2101 ( .A(b[0]), .B(a[32]), .Z(n1952) );
  XNOR U2102 ( .A(b[1]), .B(n1952), .Z(n1954) );
  NAND U2103 ( .A(a[31]), .B(n98), .Z(n1953) );
  AND U2104 ( .A(n1954), .B(n1953), .Z(n2046) );
  XNOR U2105 ( .A(n20154), .B(n2105), .Z(n2055) );
  OR U2106 ( .A(n2055), .B(n20057), .Z(n1957) );
  NANDN U2107 ( .A(n1955), .B(n20098), .Z(n1956) );
  AND U2108 ( .A(n1957), .B(n1956), .Z(n2047) );
  XOR U2109 ( .A(n2046), .B(n2047), .Z(n2049) );
  NAND U2110 ( .A(a[16]), .B(b[15]), .Z(n2048) );
  XOR U2111 ( .A(n2049), .B(n2048), .Z(n2067) );
  NAND U2112 ( .A(n19722), .B(n1958), .Z(n1960) );
  XNOR U2113 ( .A(b[5]), .B(n2729), .Z(n2058) );
  NANDN U2114 ( .A(n19640), .B(n2058), .Z(n1959) );
  NAND U2115 ( .A(n1960), .B(n1959), .Z(n2043) );
  XNOR U2116 ( .A(n19714), .B(n2600), .Z(n2061) );
  NANDN U2117 ( .A(n2061), .B(n19766), .Z(n1963) );
  NANDN U2118 ( .A(n1961), .B(n19767), .Z(n1962) );
  NAND U2119 ( .A(n1963), .B(n1962), .Z(n2040) );
  NAND U2120 ( .A(n19554), .B(n1964), .Z(n1966) );
  IV U2121 ( .A(a[30]), .Z(n2885) );
  XNOR U2122 ( .A(b[3]), .B(n2885), .Z(n2064) );
  NANDN U2123 ( .A(n19521), .B(n2064), .Z(n1965) );
  AND U2124 ( .A(n1966), .B(n1965), .Z(n2041) );
  XNOR U2125 ( .A(n2040), .B(n2041), .Z(n2042) );
  XOR U2126 ( .A(n2043), .B(n2042), .Z(n2068) );
  XOR U2127 ( .A(n2067), .B(n2068), .Z(n2069) );
  XNOR U2128 ( .A(n2070), .B(n2069), .Z(n2018) );
  NAND U2129 ( .A(n1968), .B(n1967), .Z(n1972) );
  NAND U2130 ( .A(n1970), .B(n1969), .Z(n1971) );
  NAND U2131 ( .A(n1972), .B(n1971), .Z(n2019) );
  XOR U2132 ( .A(n2018), .B(n2019), .Z(n2021) );
  XNOR U2133 ( .A(n20052), .B(n2261), .Z(n2024) );
  OR U2134 ( .A(n2024), .B(n20020), .Z(n1975) );
  NANDN U2135 ( .A(n1973), .B(n19960), .Z(n1974) );
  NAND U2136 ( .A(n1975), .B(n1974), .Z(n2037) );
  XNOR U2137 ( .A(n102), .B(n1976), .Z(n2028) );
  OR U2138 ( .A(n2028), .B(n20121), .Z(n1979) );
  NANDN U2139 ( .A(n1977), .B(n20122), .Z(n1978) );
  NAND U2140 ( .A(n1979), .B(n1978), .Z(n2034) );
  XNOR U2141 ( .A(n19975), .B(n2417), .Z(n2031) );
  NANDN U2142 ( .A(n2031), .B(n19883), .Z(n1982) );
  NANDN U2143 ( .A(n1980), .B(n19937), .Z(n1981) );
  AND U2144 ( .A(n1982), .B(n1981), .Z(n2035) );
  XNOR U2145 ( .A(n2034), .B(n2035), .Z(n2036) );
  XNOR U2146 ( .A(n2037), .B(n2036), .Z(n2073) );
  NANDN U2147 ( .A(n1984), .B(n1983), .Z(n1988) );
  NAND U2148 ( .A(n1986), .B(n1985), .Z(n1987) );
  NAND U2149 ( .A(n1988), .B(n1987), .Z(n2074) );
  XNOR U2150 ( .A(n2073), .B(n2074), .Z(n2075) );
  NANDN U2151 ( .A(n1990), .B(n1989), .Z(n1994) );
  NAND U2152 ( .A(n1992), .B(n1991), .Z(n1993) );
  AND U2153 ( .A(n1994), .B(n1993), .Z(n2076) );
  XNOR U2154 ( .A(n2075), .B(n2076), .Z(n2020) );
  XNOR U2155 ( .A(n2021), .B(n2020), .Z(n2079) );
  NANDN U2156 ( .A(n1996), .B(n1995), .Z(n2000) );
  NAND U2157 ( .A(n1998), .B(n1997), .Z(n1999) );
  NAND U2158 ( .A(n2000), .B(n1999), .Z(n2080) );
  XNOR U2159 ( .A(n2079), .B(n2080), .Z(n2081) );
  XOR U2160 ( .A(n2082), .B(n2081), .Z(n2012) );
  NANDN U2161 ( .A(n2002), .B(n2001), .Z(n2006) );
  NANDN U2162 ( .A(n2004), .B(n2003), .Z(n2005) );
  NAND U2163 ( .A(n2006), .B(n2005), .Z(n2013) );
  XNOR U2164 ( .A(n2012), .B(n2013), .Z(n2014) );
  XNOR U2165 ( .A(n2015), .B(n2014), .Z(n2085) );
  XNOR U2166 ( .A(n2085), .B(sreg[272]), .Z(n2087) );
  NAND U2167 ( .A(n2007), .B(sreg[271]), .Z(n2011) );
  OR U2168 ( .A(n2009), .B(n2008), .Z(n2010) );
  AND U2169 ( .A(n2011), .B(n2010), .Z(n2086) );
  XOR U2170 ( .A(n2087), .B(n2086), .Z(c[272]) );
  NANDN U2171 ( .A(n2013), .B(n2012), .Z(n2017) );
  NAND U2172 ( .A(n2015), .B(n2014), .Z(n2016) );
  NAND U2173 ( .A(n2017), .B(n2016), .Z(n2093) );
  NANDN U2174 ( .A(n2019), .B(n2018), .Z(n2023) );
  OR U2175 ( .A(n2021), .B(n2020), .Z(n2022) );
  NAND U2176 ( .A(n2023), .B(n2022), .Z(n2160) );
  XNOR U2177 ( .A(n20052), .B(n2366), .Z(n2102) );
  OR U2178 ( .A(n2102), .B(n20020), .Z(n2026) );
  NANDN U2179 ( .A(n2024), .B(n19960), .Z(n2025) );
  NAND U2180 ( .A(n2026), .B(n2025), .Z(n2115) );
  XNOR U2181 ( .A(n102), .B(n2027), .Z(n2106) );
  OR U2182 ( .A(n2106), .B(n20121), .Z(n2030) );
  NANDN U2183 ( .A(n2028), .B(n20122), .Z(n2029) );
  NAND U2184 ( .A(n2030), .B(n2029), .Z(n2112) );
  XNOR U2185 ( .A(n19975), .B(n2495), .Z(n2109) );
  NANDN U2186 ( .A(n2109), .B(n19883), .Z(n2033) );
  NANDN U2187 ( .A(n2031), .B(n19937), .Z(n2032) );
  AND U2188 ( .A(n2033), .B(n2032), .Z(n2113) );
  XNOR U2189 ( .A(n2112), .B(n2113), .Z(n2114) );
  XNOR U2190 ( .A(n2115), .B(n2114), .Z(n2151) );
  NANDN U2191 ( .A(n2035), .B(n2034), .Z(n2039) );
  NAND U2192 ( .A(n2037), .B(n2036), .Z(n2038) );
  NAND U2193 ( .A(n2039), .B(n2038), .Z(n2152) );
  XNOR U2194 ( .A(n2151), .B(n2152), .Z(n2153) );
  NANDN U2195 ( .A(n2041), .B(n2040), .Z(n2045) );
  NAND U2196 ( .A(n2043), .B(n2042), .Z(n2044) );
  AND U2197 ( .A(n2045), .B(n2044), .Z(n2154) );
  XNOR U2198 ( .A(n2153), .B(n2154), .Z(n2098) );
  NANDN U2199 ( .A(n2047), .B(n2046), .Z(n2051) );
  OR U2200 ( .A(n2049), .B(n2048), .Z(n2050) );
  NAND U2201 ( .A(n2051), .B(n2050), .Z(n2148) );
  NAND U2202 ( .A(b[0]), .B(a[33]), .Z(n2052) );
  XNOR U2203 ( .A(b[1]), .B(n2052), .Z(n2054) );
  NAND U2204 ( .A(a[32]), .B(n98), .Z(n2053) );
  AND U2205 ( .A(n2054), .B(n2053), .Z(n2124) );
  XNOR U2206 ( .A(n20154), .B(n2195), .Z(n2133) );
  OR U2207 ( .A(n2133), .B(n20057), .Z(n2057) );
  NANDN U2208 ( .A(n2055), .B(n20098), .Z(n2056) );
  AND U2209 ( .A(n2057), .B(n2056), .Z(n2125) );
  XOR U2210 ( .A(n2124), .B(n2125), .Z(n2127) );
  NAND U2211 ( .A(a[17]), .B(b[15]), .Z(n2126) );
  XOR U2212 ( .A(n2127), .B(n2126), .Z(n2145) );
  NAND U2213 ( .A(n19722), .B(n2058), .Z(n2060) );
  XNOR U2214 ( .A(b[5]), .B(n2807), .Z(n2136) );
  NANDN U2215 ( .A(n19640), .B(n2136), .Z(n2059) );
  NAND U2216 ( .A(n2060), .B(n2059), .Z(n2121) );
  XNOR U2217 ( .A(n19714), .B(n2651), .Z(n2139) );
  NANDN U2218 ( .A(n2139), .B(n19766), .Z(n2063) );
  NANDN U2219 ( .A(n2061), .B(n19767), .Z(n2062) );
  NAND U2220 ( .A(n2063), .B(n2062), .Z(n2118) );
  NAND U2221 ( .A(n19554), .B(n2064), .Z(n2066) );
  IV U2222 ( .A(a[31]), .Z(n2963) );
  XNOR U2223 ( .A(b[3]), .B(n2963), .Z(n2142) );
  NANDN U2224 ( .A(n19521), .B(n2142), .Z(n2065) );
  AND U2225 ( .A(n2066), .B(n2065), .Z(n2119) );
  XNOR U2226 ( .A(n2118), .B(n2119), .Z(n2120) );
  XOR U2227 ( .A(n2121), .B(n2120), .Z(n2146) );
  XOR U2228 ( .A(n2145), .B(n2146), .Z(n2147) );
  XNOR U2229 ( .A(n2148), .B(n2147), .Z(n2096) );
  NAND U2230 ( .A(n2068), .B(n2067), .Z(n2072) );
  NAND U2231 ( .A(n2070), .B(n2069), .Z(n2071) );
  NAND U2232 ( .A(n2072), .B(n2071), .Z(n2097) );
  XOR U2233 ( .A(n2096), .B(n2097), .Z(n2099) );
  XNOR U2234 ( .A(n2098), .B(n2099), .Z(n2157) );
  NANDN U2235 ( .A(n2074), .B(n2073), .Z(n2078) );
  NAND U2236 ( .A(n2076), .B(n2075), .Z(n2077) );
  NAND U2237 ( .A(n2078), .B(n2077), .Z(n2158) );
  XNOR U2238 ( .A(n2157), .B(n2158), .Z(n2159) );
  XOR U2239 ( .A(n2160), .B(n2159), .Z(n2090) );
  NANDN U2240 ( .A(n2080), .B(n2079), .Z(n2084) );
  NANDN U2241 ( .A(n2082), .B(n2081), .Z(n2083) );
  NAND U2242 ( .A(n2084), .B(n2083), .Z(n2091) );
  XNOR U2243 ( .A(n2090), .B(n2091), .Z(n2092) );
  XNOR U2244 ( .A(n2093), .B(n2092), .Z(n2163) );
  XNOR U2245 ( .A(n2163), .B(sreg[273]), .Z(n2165) );
  NAND U2246 ( .A(n2085), .B(sreg[272]), .Z(n2089) );
  OR U2247 ( .A(n2087), .B(n2086), .Z(n2088) );
  AND U2248 ( .A(n2089), .B(n2088), .Z(n2164) );
  XOR U2249 ( .A(n2165), .B(n2164), .Z(c[273]) );
  NANDN U2250 ( .A(n2091), .B(n2090), .Z(n2095) );
  NAND U2251 ( .A(n2093), .B(n2092), .Z(n2094) );
  NAND U2252 ( .A(n2095), .B(n2094), .Z(n2171) );
  NANDN U2253 ( .A(n2097), .B(n2096), .Z(n2101) );
  OR U2254 ( .A(n2099), .B(n2098), .Z(n2100) );
  NAND U2255 ( .A(n2101), .B(n2100), .Z(n2238) );
  XNOR U2256 ( .A(n20052), .B(n2417), .Z(n2192) );
  OR U2257 ( .A(n2192), .B(n20020), .Z(n2104) );
  NANDN U2258 ( .A(n2102), .B(n19960), .Z(n2103) );
  NAND U2259 ( .A(n2104), .B(n2103), .Z(n2189) );
  XNOR U2260 ( .A(n102), .B(n2105), .Z(n2196) );
  OR U2261 ( .A(n2196), .B(n20121), .Z(n2108) );
  NANDN U2262 ( .A(n2106), .B(n20122), .Z(n2107) );
  NAND U2263 ( .A(n2108), .B(n2107), .Z(n2186) );
  XNOR U2264 ( .A(n19975), .B(n2600), .Z(n2199) );
  NANDN U2265 ( .A(n2199), .B(n19883), .Z(n2111) );
  NANDN U2266 ( .A(n2109), .B(n19937), .Z(n2110) );
  AND U2267 ( .A(n2111), .B(n2110), .Z(n2187) );
  XNOR U2268 ( .A(n2186), .B(n2187), .Z(n2188) );
  XNOR U2269 ( .A(n2189), .B(n2188), .Z(n2229) );
  NANDN U2270 ( .A(n2113), .B(n2112), .Z(n2117) );
  NAND U2271 ( .A(n2115), .B(n2114), .Z(n2116) );
  NAND U2272 ( .A(n2117), .B(n2116), .Z(n2230) );
  XNOR U2273 ( .A(n2229), .B(n2230), .Z(n2231) );
  NANDN U2274 ( .A(n2119), .B(n2118), .Z(n2123) );
  NAND U2275 ( .A(n2121), .B(n2120), .Z(n2122) );
  AND U2276 ( .A(n2123), .B(n2122), .Z(n2232) );
  XNOR U2277 ( .A(n2231), .B(n2232), .Z(n2176) );
  NANDN U2278 ( .A(n2125), .B(n2124), .Z(n2129) );
  OR U2279 ( .A(n2127), .B(n2126), .Z(n2128) );
  NAND U2280 ( .A(n2129), .B(n2128), .Z(n2226) );
  NAND U2281 ( .A(b[0]), .B(a[34]), .Z(n2130) );
  XNOR U2282 ( .A(b[1]), .B(n2130), .Z(n2132) );
  NAND U2283 ( .A(a[33]), .B(n98), .Z(n2131) );
  AND U2284 ( .A(n2132), .B(n2131), .Z(n2202) );
  XNOR U2285 ( .A(n20154), .B(n2261), .Z(n2211) );
  OR U2286 ( .A(n2211), .B(n20057), .Z(n2135) );
  NANDN U2287 ( .A(n2133), .B(n20098), .Z(n2134) );
  AND U2288 ( .A(n2135), .B(n2134), .Z(n2203) );
  XOR U2289 ( .A(n2202), .B(n2203), .Z(n2205) );
  NAND U2290 ( .A(a[18]), .B(b[15]), .Z(n2204) );
  XOR U2291 ( .A(n2205), .B(n2204), .Z(n2223) );
  NAND U2292 ( .A(n19722), .B(n2136), .Z(n2138) );
  XNOR U2293 ( .A(b[5]), .B(n2885), .Z(n2214) );
  NANDN U2294 ( .A(n19640), .B(n2214), .Z(n2137) );
  NAND U2295 ( .A(n2138), .B(n2137), .Z(n2183) );
  XNOR U2296 ( .A(n19714), .B(n2729), .Z(n2217) );
  NANDN U2297 ( .A(n2217), .B(n19766), .Z(n2141) );
  NANDN U2298 ( .A(n2139), .B(n19767), .Z(n2140) );
  NAND U2299 ( .A(n2141), .B(n2140), .Z(n2180) );
  NAND U2300 ( .A(n19554), .B(n2142), .Z(n2144) );
  IV U2301 ( .A(a[32]), .Z(n3068) );
  XNOR U2302 ( .A(b[3]), .B(n3068), .Z(n2220) );
  NANDN U2303 ( .A(n19521), .B(n2220), .Z(n2143) );
  AND U2304 ( .A(n2144), .B(n2143), .Z(n2181) );
  XNOR U2305 ( .A(n2180), .B(n2181), .Z(n2182) );
  XOR U2306 ( .A(n2183), .B(n2182), .Z(n2224) );
  XOR U2307 ( .A(n2223), .B(n2224), .Z(n2225) );
  XNOR U2308 ( .A(n2226), .B(n2225), .Z(n2174) );
  NAND U2309 ( .A(n2146), .B(n2145), .Z(n2150) );
  NAND U2310 ( .A(n2148), .B(n2147), .Z(n2149) );
  NAND U2311 ( .A(n2150), .B(n2149), .Z(n2175) );
  XOR U2312 ( .A(n2174), .B(n2175), .Z(n2177) );
  XNOR U2313 ( .A(n2176), .B(n2177), .Z(n2235) );
  NANDN U2314 ( .A(n2152), .B(n2151), .Z(n2156) );
  NAND U2315 ( .A(n2154), .B(n2153), .Z(n2155) );
  NAND U2316 ( .A(n2156), .B(n2155), .Z(n2236) );
  XNOR U2317 ( .A(n2235), .B(n2236), .Z(n2237) );
  XOR U2318 ( .A(n2238), .B(n2237), .Z(n2168) );
  NANDN U2319 ( .A(n2158), .B(n2157), .Z(n2162) );
  NANDN U2320 ( .A(n2160), .B(n2159), .Z(n2161) );
  NAND U2321 ( .A(n2162), .B(n2161), .Z(n2169) );
  XNOR U2322 ( .A(n2168), .B(n2169), .Z(n2170) );
  XNOR U2323 ( .A(n2171), .B(n2170), .Z(n2241) );
  XNOR U2324 ( .A(n2241), .B(sreg[274]), .Z(n2243) );
  NAND U2325 ( .A(n2163), .B(sreg[273]), .Z(n2167) );
  OR U2326 ( .A(n2165), .B(n2164), .Z(n2166) );
  AND U2327 ( .A(n2167), .B(n2166), .Z(n2242) );
  XOR U2328 ( .A(n2243), .B(n2242), .Z(c[274]) );
  NANDN U2329 ( .A(n2169), .B(n2168), .Z(n2173) );
  NAND U2330 ( .A(n2171), .B(n2170), .Z(n2172) );
  NAND U2331 ( .A(n2173), .B(n2172), .Z(n2249) );
  NANDN U2332 ( .A(n2175), .B(n2174), .Z(n2179) );
  OR U2333 ( .A(n2177), .B(n2176), .Z(n2178) );
  NAND U2334 ( .A(n2179), .B(n2178), .Z(n2316) );
  NANDN U2335 ( .A(n2181), .B(n2180), .Z(n2185) );
  NAND U2336 ( .A(n2183), .B(n2182), .Z(n2184) );
  NAND U2337 ( .A(n2185), .B(n2184), .Z(n2310) );
  NANDN U2338 ( .A(n2187), .B(n2186), .Z(n2191) );
  NAND U2339 ( .A(n2189), .B(n2188), .Z(n2190) );
  NAND U2340 ( .A(n2191), .B(n2190), .Z(n2307) );
  XNOR U2341 ( .A(n20052), .B(n2495), .Z(n2258) );
  OR U2342 ( .A(n2258), .B(n20020), .Z(n2194) );
  NANDN U2343 ( .A(n2192), .B(n19960), .Z(n2193) );
  NAND U2344 ( .A(n2194), .B(n2193), .Z(n2271) );
  XNOR U2345 ( .A(n102), .B(n2195), .Z(n2262) );
  OR U2346 ( .A(n2262), .B(n20121), .Z(n2198) );
  NANDN U2347 ( .A(n2196), .B(n20122), .Z(n2197) );
  NAND U2348 ( .A(n2198), .B(n2197), .Z(n2268) );
  XNOR U2349 ( .A(n19975), .B(n2651), .Z(n2265) );
  NANDN U2350 ( .A(n2265), .B(n19883), .Z(n2201) );
  NANDN U2351 ( .A(n2199), .B(n19937), .Z(n2200) );
  AND U2352 ( .A(n2201), .B(n2200), .Z(n2269) );
  XNOR U2353 ( .A(n2268), .B(n2269), .Z(n2270) );
  XNOR U2354 ( .A(n2271), .B(n2270), .Z(n2308) );
  XNOR U2355 ( .A(n2307), .B(n2308), .Z(n2309) );
  XNOR U2356 ( .A(n2310), .B(n2309), .Z(n2255) );
  NANDN U2357 ( .A(n2203), .B(n2202), .Z(n2207) );
  OR U2358 ( .A(n2205), .B(n2204), .Z(n2206) );
  NAND U2359 ( .A(n2207), .B(n2206), .Z(n2304) );
  NAND U2360 ( .A(b[0]), .B(a[35]), .Z(n2208) );
  XNOR U2361 ( .A(b[1]), .B(n2208), .Z(n2210) );
  NAND U2362 ( .A(a[34]), .B(n98), .Z(n2209) );
  AND U2363 ( .A(n2210), .B(n2209), .Z(n2280) );
  XNOR U2364 ( .A(n20154), .B(n2366), .Z(n2289) );
  OR U2365 ( .A(n2289), .B(n20057), .Z(n2213) );
  NANDN U2366 ( .A(n2211), .B(n20098), .Z(n2212) );
  AND U2367 ( .A(n2213), .B(n2212), .Z(n2281) );
  XOR U2368 ( .A(n2280), .B(n2281), .Z(n2283) );
  NAND U2369 ( .A(a[19]), .B(b[15]), .Z(n2282) );
  XOR U2370 ( .A(n2283), .B(n2282), .Z(n2301) );
  NAND U2371 ( .A(n19722), .B(n2214), .Z(n2216) );
  XNOR U2372 ( .A(b[5]), .B(n2963), .Z(n2292) );
  NANDN U2373 ( .A(n19640), .B(n2292), .Z(n2215) );
  NAND U2374 ( .A(n2216), .B(n2215), .Z(n2277) );
  XNOR U2375 ( .A(n19714), .B(n2807), .Z(n2295) );
  NANDN U2376 ( .A(n2295), .B(n19766), .Z(n2219) );
  NANDN U2377 ( .A(n2217), .B(n19767), .Z(n2218) );
  NAND U2378 ( .A(n2219), .B(n2218), .Z(n2274) );
  NAND U2379 ( .A(n19554), .B(n2220), .Z(n2222) );
  IV U2380 ( .A(a[33]), .Z(n3146) );
  XNOR U2381 ( .A(b[3]), .B(n3146), .Z(n2298) );
  NANDN U2382 ( .A(n19521), .B(n2298), .Z(n2221) );
  AND U2383 ( .A(n2222), .B(n2221), .Z(n2275) );
  XNOR U2384 ( .A(n2274), .B(n2275), .Z(n2276) );
  XOR U2385 ( .A(n2277), .B(n2276), .Z(n2302) );
  XOR U2386 ( .A(n2301), .B(n2302), .Z(n2303) );
  XNOR U2387 ( .A(n2304), .B(n2303), .Z(n2252) );
  NAND U2388 ( .A(n2224), .B(n2223), .Z(n2228) );
  NAND U2389 ( .A(n2226), .B(n2225), .Z(n2227) );
  NAND U2390 ( .A(n2228), .B(n2227), .Z(n2253) );
  XNOR U2391 ( .A(n2252), .B(n2253), .Z(n2254) );
  XOR U2392 ( .A(n2255), .B(n2254), .Z(n2313) );
  NANDN U2393 ( .A(n2230), .B(n2229), .Z(n2234) );
  NAND U2394 ( .A(n2232), .B(n2231), .Z(n2233) );
  NAND U2395 ( .A(n2234), .B(n2233), .Z(n2314) );
  XOR U2396 ( .A(n2313), .B(n2314), .Z(n2315) );
  XOR U2397 ( .A(n2316), .B(n2315), .Z(n2246) );
  NANDN U2398 ( .A(n2236), .B(n2235), .Z(n2240) );
  NANDN U2399 ( .A(n2238), .B(n2237), .Z(n2239) );
  NAND U2400 ( .A(n2240), .B(n2239), .Z(n2247) );
  XNOR U2401 ( .A(n2246), .B(n2247), .Z(n2248) );
  XNOR U2402 ( .A(n2249), .B(n2248), .Z(n2319) );
  XNOR U2403 ( .A(n2319), .B(sreg[275]), .Z(n2321) );
  NAND U2404 ( .A(n2241), .B(sreg[274]), .Z(n2245) );
  OR U2405 ( .A(n2243), .B(n2242), .Z(n2244) );
  AND U2406 ( .A(n2245), .B(n2244), .Z(n2320) );
  XOR U2407 ( .A(n2321), .B(n2320), .Z(c[275]) );
  NANDN U2408 ( .A(n2247), .B(n2246), .Z(n2251) );
  NAND U2409 ( .A(n2249), .B(n2248), .Z(n2250) );
  NAND U2410 ( .A(n2251), .B(n2250), .Z(n2327) );
  NANDN U2411 ( .A(n2253), .B(n2252), .Z(n2257) );
  NAND U2412 ( .A(n2255), .B(n2254), .Z(n2256) );
  NAND U2413 ( .A(n2257), .B(n2256), .Z(n2394) );
  XNOR U2414 ( .A(n20052), .B(n2600), .Z(n2363) );
  OR U2415 ( .A(n2363), .B(n20020), .Z(n2260) );
  NANDN U2416 ( .A(n2258), .B(n19960), .Z(n2259) );
  NAND U2417 ( .A(n2260), .B(n2259), .Z(n2376) );
  XNOR U2418 ( .A(n102), .B(n2261), .Z(n2367) );
  OR U2419 ( .A(n2367), .B(n20121), .Z(n2264) );
  NANDN U2420 ( .A(n2262), .B(n20122), .Z(n2263) );
  NAND U2421 ( .A(n2264), .B(n2263), .Z(n2373) );
  XNOR U2422 ( .A(n19975), .B(n2729), .Z(n2370) );
  NANDN U2423 ( .A(n2370), .B(n19883), .Z(n2267) );
  NANDN U2424 ( .A(n2265), .B(n19937), .Z(n2266) );
  AND U2425 ( .A(n2267), .B(n2266), .Z(n2374) );
  XNOR U2426 ( .A(n2373), .B(n2374), .Z(n2375) );
  XNOR U2427 ( .A(n2376), .B(n2375), .Z(n2385) );
  NANDN U2428 ( .A(n2269), .B(n2268), .Z(n2273) );
  NAND U2429 ( .A(n2271), .B(n2270), .Z(n2272) );
  NAND U2430 ( .A(n2273), .B(n2272), .Z(n2386) );
  XNOR U2431 ( .A(n2385), .B(n2386), .Z(n2387) );
  NANDN U2432 ( .A(n2275), .B(n2274), .Z(n2279) );
  NAND U2433 ( .A(n2277), .B(n2276), .Z(n2278) );
  AND U2434 ( .A(n2279), .B(n2278), .Z(n2388) );
  XNOR U2435 ( .A(n2387), .B(n2388), .Z(n2332) );
  NANDN U2436 ( .A(n2281), .B(n2280), .Z(n2285) );
  OR U2437 ( .A(n2283), .B(n2282), .Z(n2284) );
  NAND U2438 ( .A(n2285), .B(n2284), .Z(n2360) );
  NAND U2439 ( .A(b[0]), .B(a[36]), .Z(n2286) );
  XNOR U2440 ( .A(b[1]), .B(n2286), .Z(n2288) );
  NAND U2441 ( .A(a[35]), .B(n98), .Z(n2287) );
  AND U2442 ( .A(n2288), .B(n2287), .Z(n2336) );
  XNOR U2443 ( .A(n20154), .B(n2417), .Z(n2345) );
  OR U2444 ( .A(n2345), .B(n20057), .Z(n2291) );
  NANDN U2445 ( .A(n2289), .B(n20098), .Z(n2290) );
  AND U2446 ( .A(n2291), .B(n2290), .Z(n2337) );
  XOR U2447 ( .A(n2336), .B(n2337), .Z(n2339) );
  NAND U2448 ( .A(a[20]), .B(b[15]), .Z(n2338) );
  XOR U2449 ( .A(n2339), .B(n2338), .Z(n2357) );
  NAND U2450 ( .A(n19722), .B(n2292), .Z(n2294) );
  XNOR U2451 ( .A(b[5]), .B(n3068), .Z(n2348) );
  NANDN U2452 ( .A(n19640), .B(n2348), .Z(n2293) );
  NAND U2453 ( .A(n2294), .B(n2293), .Z(n2382) );
  XNOR U2454 ( .A(n19714), .B(n2885), .Z(n2351) );
  NANDN U2455 ( .A(n2351), .B(n19766), .Z(n2297) );
  NANDN U2456 ( .A(n2295), .B(n19767), .Z(n2296) );
  NAND U2457 ( .A(n2297), .B(n2296), .Z(n2379) );
  NAND U2458 ( .A(n19554), .B(n2298), .Z(n2300) );
  IV U2459 ( .A(a[34]), .Z(n3224) );
  XNOR U2460 ( .A(b[3]), .B(n3224), .Z(n2354) );
  NANDN U2461 ( .A(n19521), .B(n2354), .Z(n2299) );
  AND U2462 ( .A(n2300), .B(n2299), .Z(n2380) );
  XNOR U2463 ( .A(n2379), .B(n2380), .Z(n2381) );
  XOR U2464 ( .A(n2382), .B(n2381), .Z(n2358) );
  XOR U2465 ( .A(n2357), .B(n2358), .Z(n2359) );
  XNOR U2466 ( .A(n2360), .B(n2359), .Z(n2330) );
  NAND U2467 ( .A(n2302), .B(n2301), .Z(n2306) );
  NAND U2468 ( .A(n2304), .B(n2303), .Z(n2305) );
  NAND U2469 ( .A(n2306), .B(n2305), .Z(n2331) );
  XOR U2470 ( .A(n2330), .B(n2331), .Z(n2333) );
  XNOR U2471 ( .A(n2332), .B(n2333), .Z(n2391) );
  NANDN U2472 ( .A(n2308), .B(n2307), .Z(n2312) );
  NAND U2473 ( .A(n2310), .B(n2309), .Z(n2311) );
  AND U2474 ( .A(n2312), .B(n2311), .Z(n2392) );
  XNOR U2475 ( .A(n2391), .B(n2392), .Z(n2393) );
  XOR U2476 ( .A(n2394), .B(n2393), .Z(n2324) );
  OR U2477 ( .A(n2314), .B(n2313), .Z(n2318) );
  NANDN U2478 ( .A(n2316), .B(n2315), .Z(n2317) );
  NAND U2479 ( .A(n2318), .B(n2317), .Z(n2325) );
  XNOR U2480 ( .A(n2324), .B(n2325), .Z(n2326) );
  XNOR U2481 ( .A(n2327), .B(n2326), .Z(n2397) );
  XNOR U2482 ( .A(n2397), .B(sreg[276]), .Z(n2399) );
  NAND U2483 ( .A(n2319), .B(sreg[275]), .Z(n2323) );
  OR U2484 ( .A(n2321), .B(n2320), .Z(n2322) );
  AND U2485 ( .A(n2323), .B(n2322), .Z(n2398) );
  XOR U2486 ( .A(n2399), .B(n2398), .Z(c[276]) );
  NANDN U2487 ( .A(n2325), .B(n2324), .Z(n2329) );
  NAND U2488 ( .A(n2327), .B(n2326), .Z(n2328) );
  NAND U2489 ( .A(n2329), .B(n2328), .Z(n2405) );
  NANDN U2490 ( .A(n2331), .B(n2330), .Z(n2335) );
  OR U2491 ( .A(n2333), .B(n2332), .Z(n2334) );
  NAND U2492 ( .A(n2335), .B(n2334), .Z(n2472) );
  NANDN U2493 ( .A(n2337), .B(n2336), .Z(n2341) );
  OR U2494 ( .A(n2339), .B(n2338), .Z(n2340) );
  NAND U2495 ( .A(n2341), .B(n2340), .Z(n2460) );
  NAND U2496 ( .A(b[0]), .B(a[37]), .Z(n2342) );
  XNOR U2497 ( .A(b[1]), .B(n2342), .Z(n2344) );
  NAND U2498 ( .A(a[36]), .B(n98), .Z(n2343) );
  AND U2499 ( .A(n2344), .B(n2343), .Z(n2436) );
  XNOR U2500 ( .A(n20154), .B(n2495), .Z(n2445) );
  OR U2501 ( .A(n2445), .B(n20057), .Z(n2347) );
  NANDN U2502 ( .A(n2345), .B(n20098), .Z(n2346) );
  AND U2503 ( .A(n2347), .B(n2346), .Z(n2437) );
  XOR U2504 ( .A(n2436), .B(n2437), .Z(n2439) );
  NAND U2505 ( .A(a[21]), .B(b[15]), .Z(n2438) );
  XOR U2506 ( .A(n2439), .B(n2438), .Z(n2457) );
  NAND U2507 ( .A(n19722), .B(n2348), .Z(n2350) );
  XNOR U2508 ( .A(b[5]), .B(n3146), .Z(n2448) );
  NANDN U2509 ( .A(n19640), .B(n2448), .Z(n2349) );
  NAND U2510 ( .A(n2350), .B(n2349), .Z(n2433) );
  XNOR U2511 ( .A(n19714), .B(n2963), .Z(n2451) );
  NANDN U2512 ( .A(n2451), .B(n19766), .Z(n2353) );
  NANDN U2513 ( .A(n2351), .B(n19767), .Z(n2352) );
  NAND U2514 ( .A(n2353), .B(n2352), .Z(n2430) );
  NAND U2515 ( .A(n19554), .B(n2354), .Z(n2356) );
  IV U2516 ( .A(a[35]), .Z(n3275) );
  XNOR U2517 ( .A(b[3]), .B(n3275), .Z(n2454) );
  NANDN U2518 ( .A(n19521), .B(n2454), .Z(n2355) );
  AND U2519 ( .A(n2356), .B(n2355), .Z(n2431) );
  XNOR U2520 ( .A(n2430), .B(n2431), .Z(n2432) );
  XOR U2521 ( .A(n2433), .B(n2432), .Z(n2458) );
  XOR U2522 ( .A(n2457), .B(n2458), .Z(n2459) );
  XNOR U2523 ( .A(n2460), .B(n2459), .Z(n2408) );
  NAND U2524 ( .A(n2358), .B(n2357), .Z(n2362) );
  NAND U2525 ( .A(n2360), .B(n2359), .Z(n2361) );
  NAND U2526 ( .A(n2362), .B(n2361), .Z(n2409) );
  XOR U2527 ( .A(n2408), .B(n2409), .Z(n2411) );
  XNOR U2528 ( .A(n20052), .B(n2651), .Z(n2414) );
  OR U2529 ( .A(n2414), .B(n20020), .Z(n2365) );
  NANDN U2530 ( .A(n2363), .B(n19960), .Z(n2364) );
  NAND U2531 ( .A(n2365), .B(n2364), .Z(n2427) );
  XNOR U2532 ( .A(n102), .B(n2366), .Z(n2418) );
  OR U2533 ( .A(n2418), .B(n20121), .Z(n2369) );
  NANDN U2534 ( .A(n2367), .B(n20122), .Z(n2368) );
  NAND U2535 ( .A(n2369), .B(n2368), .Z(n2424) );
  XNOR U2536 ( .A(n19975), .B(n2807), .Z(n2421) );
  NANDN U2537 ( .A(n2421), .B(n19883), .Z(n2372) );
  NANDN U2538 ( .A(n2370), .B(n19937), .Z(n2371) );
  AND U2539 ( .A(n2372), .B(n2371), .Z(n2425) );
  XNOR U2540 ( .A(n2424), .B(n2425), .Z(n2426) );
  XNOR U2541 ( .A(n2427), .B(n2426), .Z(n2463) );
  NANDN U2542 ( .A(n2374), .B(n2373), .Z(n2378) );
  NAND U2543 ( .A(n2376), .B(n2375), .Z(n2377) );
  NAND U2544 ( .A(n2378), .B(n2377), .Z(n2464) );
  XNOR U2545 ( .A(n2463), .B(n2464), .Z(n2465) );
  NANDN U2546 ( .A(n2380), .B(n2379), .Z(n2384) );
  NAND U2547 ( .A(n2382), .B(n2381), .Z(n2383) );
  AND U2548 ( .A(n2384), .B(n2383), .Z(n2466) );
  XNOR U2549 ( .A(n2465), .B(n2466), .Z(n2410) );
  XNOR U2550 ( .A(n2411), .B(n2410), .Z(n2469) );
  NANDN U2551 ( .A(n2386), .B(n2385), .Z(n2390) );
  NAND U2552 ( .A(n2388), .B(n2387), .Z(n2389) );
  NAND U2553 ( .A(n2390), .B(n2389), .Z(n2470) );
  XNOR U2554 ( .A(n2469), .B(n2470), .Z(n2471) );
  XOR U2555 ( .A(n2472), .B(n2471), .Z(n2402) );
  NANDN U2556 ( .A(n2392), .B(n2391), .Z(n2396) );
  NANDN U2557 ( .A(n2394), .B(n2393), .Z(n2395) );
  NAND U2558 ( .A(n2396), .B(n2395), .Z(n2403) );
  XNOR U2559 ( .A(n2402), .B(n2403), .Z(n2404) );
  XNOR U2560 ( .A(n2405), .B(n2404), .Z(n2475) );
  XNOR U2561 ( .A(n2475), .B(sreg[277]), .Z(n2477) );
  NAND U2562 ( .A(n2397), .B(sreg[276]), .Z(n2401) );
  OR U2563 ( .A(n2399), .B(n2398), .Z(n2400) );
  AND U2564 ( .A(n2401), .B(n2400), .Z(n2476) );
  XOR U2565 ( .A(n2477), .B(n2476), .Z(c[277]) );
  NANDN U2566 ( .A(n2403), .B(n2402), .Z(n2407) );
  NAND U2567 ( .A(n2405), .B(n2404), .Z(n2406) );
  NAND U2568 ( .A(n2407), .B(n2406), .Z(n2483) );
  NANDN U2569 ( .A(n2409), .B(n2408), .Z(n2413) );
  OR U2570 ( .A(n2411), .B(n2410), .Z(n2412) );
  NAND U2571 ( .A(n2413), .B(n2412), .Z(n2550) );
  XNOR U2572 ( .A(n20052), .B(n2729), .Z(n2492) );
  OR U2573 ( .A(n2492), .B(n20020), .Z(n2416) );
  NANDN U2574 ( .A(n2414), .B(n19960), .Z(n2415) );
  NAND U2575 ( .A(n2416), .B(n2415), .Z(n2505) );
  XNOR U2576 ( .A(n102), .B(n2417), .Z(n2496) );
  OR U2577 ( .A(n2496), .B(n20121), .Z(n2420) );
  NANDN U2578 ( .A(n2418), .B(n20122), .Z(n2419) );
  NAND U2579 ( .A(n2420), .B(n2419), .Z(n2502) );
  XNOR U2580 ( .A(n19975), .B(n2885), .Z(n2499) );
  NANDN U2581 ( .A(n2499), .B(n19883), .Z(n2423) );
  NANDN U2582 ( .A(n2421), .B(n19937), .Z(n2422) );
  AND U2583 ( .A(n2423), .B(n2422), .Z(n2503) );
  XNOR U2584 ( .A(n2502), .B(n2503), .Z(n2504) );
  XNOR U2585 ( .A(n2505), .B(n2504), .Z(n2541) );
  NANDN U2586 ( .A(n2425), .B(n2424), .Z(n2429) );
  NAND U2587 ( .A(n2427), .B(n2426), .Z(n2428) );
  NAND U2588 ( .A(n2429), .B(n2428), .Z(n2542) );
  XNOR U2589 ( .A(n2541), .B(n2542), .Z(n2543) );
  NANDN U2590 ( .A(n2431), .B(n2430), .Z(n2435) );
  NAND U2591 ( .A(n2433), .B(n2432), .Z(n2434) );
  AND U2592 ( .A(n2435), .B(n2434), .Z(n2544) );
  XNOR U2593 ( .A(n2543), .B(n2544), .Z(n2488) );
  NANDN U2594 ( .A(n2437), .B(n2436), .Z(n2441) );
  OR U2595 ( .A(n2439), .B(n2438), .Z(n2440) );
  NAND U2596 ( .A(n2441), .B(n2440), .Z(n2538) );
  NAND U2597 ( .A(b[0]), .B(a[38]), .Z(n2442) );
  XNOR U2598 ( .A(b[1]), .B(n2442), .Z(n2444) );
  NAND U2599 ( .A(a[37]), .B(n98), .Z(n2443) );
  AND U2600 ( .A(n2444), .B(n2443), .Z(n2514) );
  XNOR U2601 ( .A(n20154), .B(n2600), .Z(n2523) );
  OR U2602 ( .A(n2523), .B(n20057), .Z(n2447) );
  NANDN U2603 ( .A(n2445), .B(n20098), .Z(n2446) );
  AND U2604 ( .A(n2447), .B(n2446), .Z(n2515) );
  XOR U2605 ( .A(n2514), .B(n2515), .Z(n2517) );
  NAND U2606 ( .A(a[22]), .B(b[15]), .Z(n2516) );
  XOR U2607 ( .A(n2517), .B(n2516), .Z(n2535) );
  NAND U2608 ( .A(n19722), .B(n2448), .Z(n2450) );
  XNOR U2609 ( .A(b[5]), .B(n3224), .Z(n2526) );
  NANDN U2610 ( .A(n19640), .B(n2526), .Z(n2449) );
  NAND U2611 ( .A(n2450), .B(n2449), .Z(n2511) );
  XNOR U2612 ( .A(n19714), .B(n3068), .Z(n2529) );
  NANDN U2613 ( .A(n2529), .B(n19766), .Z(n2453) );
  NANDN U2614 ( .A(n2451), .B(n19767), .Z(n2452) );
  NAND U2615 ( .A(n2453), .B(n2452), .Z(n2508) );
  NAND U2616 ( .A(n19554), .B(n2454), .Z(n2456) );
  IV U2617 ( .A(a[36]), .Z(n3353) );
  XNOR U2618 ( .A(b[3]), .B(n3353), .Z(n2532) );
  NANDN U2619 ( .A(n19521), .B(n2532), .Z(n2455) );
  AND U2620 ( .A(n2456), .B(n2455), .Z(n2509) );
  XNOR U2621 ( .A(n2508), .B(n2509), .Z(n2510) );
  XOR U2622 ( .A(n2511), .B(n2510), .Z(n2536) );
  XOR U2623 ( .A(n2535), .B(n2536), .Z(n2537) );
  XNOR U2624 ( .A(n2538), .B(n2537), .Z(n2486) );
  NAND U2625 ( .A(n2458), .B(n2457), .Z(n2462) );
  NAND U2626 ( .A(n2460), .B(n2459), .Z(n2461) );
  NAND U2627 ( .A(n2462), .B(n2461), .Z(n2487) );
  XOR U2628 ( .A(n2486), .B(n2487), .Z(n2489) );
  XNOR U2629 ( .A(n2488), .B(n2489), .Z(n2547) );
  NANDN U2630 ( .A(n2464), .B(n2463), .Z(n2468) );
  NAND U2631 ( .A(n2466), .B(n2465), .Z(n2467) );
  NAND U2632 ( .A(n2468), .B(n2467), .Z(n2548) );
  XNOR U2633 ( .A(n2547), .B(n2548), .Z(n2549) );
  XOR U2634 ( .A(n2550), .B(n2549), .Z(n2480) );
  NANDN U2635 ( .A(n2470), .B(n2469), .Z(n2474) );
  NANDN U2636 ( .A(n2472), .B(n2471), .Z(n2473) );
  NAND U2637 ( .A(n2474), .B(n2473), .Z(n2481) );
  XNOR U2638 ( .A(n2480), .B(n2481), .Z(n2482) );
  XNOR U2639 ( .A(n2483), .B(n2482), .Z(n2553) );
  XNOR U2640 ( .A(n2553), .B(sreg[278]), .Z(n2555) );
  NAND U2641 ( .A(n2475), .B(sreg[277]), .Z(n2479) );
  OR U2642 ( .A(n2477), .B(n2476), .Z(n2478) );
  AND U2643 ( .A(n2479), .B(n2478), .Z(n2554) );
  XOR U2644 ( .A(n2555), .B(n2554), .Z(c[278]) );
  NANDN U2645 ( .A(n2481), .B(n2480), .Z(n2485) );
  NAND U2646 ( .A(n2483), .B(n2482), .Z(n2484) );
  NAND U2647 ( .A(n2485), .B(n2484), .Z(n2561) );
  NANDN U2648 ( .A(n2487), .B(n2486), .Z(n2491) );
  OR U2649 ( .A(n2489), .B(n2488), .Z(n2490) );
  NAND U2650 ( .A(n2491), .B(n2490), .Z(n2628) );
  XNOR U2651 ( .A(n20052), .B(n2807), .Z(n2597) );
  OR U2652 ( .A(n2597), .B(n20020), .Z(n2494) );
  NANDN U2653 ( .A(n2492), .B(n19960), .Z(n2493) );
  NAND U2654 ( .A(n2494), .B(n2493), .Z(n2610) );
  XNOR U2655 ( .A(n102), .B(n2495), .Z(n2601) );
  OR U2656 ( .A(n2601), .B(n20121), .Z(n2498) );
  NANDN U2657 ( .A(n2496), .B(n20122), .Z(n2497) );
  NAND U2658 ( .A(n2498), .B(n2497), .Z(n2607) );
  XNOR U2659 ( .A(n19975), .B(n2963), .Z(n2604) );
  NANDN U2660 ( .A(n2604), .B(n19883), .Z(n2501) );
  NANDN U2661 ( .A(n2499), .B(n19937), .Z(n2500) );
  AND U2662 ( .A(n2501), .B(n2500), .Z(n2608) );
  XNOR U2663 ( .A(n2607), .B(n2608), .Z(n2609) );
  XNOR U2664 ( .A(n2610), .B(n2609), .Z(n2619) );
  NANDN U2665 ( .A(n2503), .B(n2502), .Z(n2507) );
  NAND U2666 ( .A(n2505), .B(n2504), .Z(n2506) );
  NAND U2667 ( .A(n2507), .B(n2506), .Z(n2620) );
  XNOR U2668 ( .A(n2619), .B(n2620), .Z(n2621) );
  NANDN U2669 ( .A(n2509), .B(n2508), .Z(n2513) );
  NAND U2670 ( .A(n2511), .B(n2510), .Z(n2512) );
  AND U2671 ( .A(n2513), .B(n2512), .Z(n2622) );
  XNOR U2672 ( .A(n2621), .B(n2622), .Z(n2566) );
  NANDN U2673 ( .A(n2515), .B(n2514), .Z(n2519) );
  OR U2674 ( .A(n2517), .B(n2516), .Z(n2518) );
  NAND U2675 ( .A(n2519), .B(n2518), .Z(n2594) );
  NAND U2676 ( .A(b[0]), .B(a[39]), .Z(n2520) );
  XNOR U2677 ( .A(b[1]), .B(n2520), .Z(n2522) );
  NAND U2678 ( .A(a[38]), .B(n98), .Z(n2521) );
  AND U2679 ( .A(n2522), .B(n2521), .Z(n2570) );
  XNOR U2680 ( .A(n20154), .B(n2651), .Z(n2579) );
  OR U2681 ( .A(n2579), .B(n20057), .Z(n2525) );
  NANDN U2682 ( .A(n2523), .B(n20098), .Z(n2524) );
  AND U2683 ( .A(n2525), .B(n2524), .Z(n2571) );
  XOR U2684 ( .A(n2570), .B(n2571), .Z(n2573) );
  NAND U2685 ( .A(a[23]), .B(b[15]), .Z(n2572) );
  XOR U2686 ( .A(n2573), .B(n2572), .Z(n2591) );
  NAND U2687 ( .A(n19722), .B(n2526), .Z(n2528) );
  XNOR U2688 ( .A(b[5]), .B(n3275), .Z(n2582) );
  NANDN U2689 ( .A(n19640), .B(n2582), .Z(n2527) );
  NAND U2690 ( .A(n2528), .B(n2527), .Z(n2616) );
  XNOR U2691 ( .A(n19714), .B(n3146), .Z(n2585) );
  NANDN U2692 ( .A(n2585), .B(n19766), .Z(n2531) );
  NANDN U2693 ( .A(n2529), .B(n19767), .Z(n2530) );
  NAND U2694 ( .A(n2531), .B(n2530), .Z(n2613) );
  NAND U2695 ( .A(n19554), .B(n2532), .Z(n2534) );
  IV U2696 ( .A(a[37]), .Z(n3458) );
  XNOR U2697 ( .A(b[3]), .B(n3458), .Z(n2588) );
  NANDN U2698 ( .A(n19521), .B(n2588), .Z(n2533) );
  AND U2699 ( .A(n2534), .B(n2533), .Z(n2614) );
  XNOR U2700 ( .A(n2613), .B(n2614), .Z(n2615) );
  XOR U2701 ( .A(n2616), .B(n2615), .Z(n2592) );
  XOR U2702 ( .A(n2591), .B(n2592), .Z(n2593) );
  XNOR U2703 ( .A(n2594), .B(n2593), .Z(n2564) );
  NAND U2704 ( .A(n2536), .B(n2535), .Z(n2540) );
  NAND U2705 ( .A(n2538), .B(n2537), .Z(n2539) );
  NAND U2706 ( .A(n2540), .B(n2539), .Z(n2565) );
  XOR U2707 ( .A(n2564), .B(n2565), .Z(n2567) );
  XNOR U2708 ( .A(n2566), .B(n2567), .Z(n2625) );
  NANDN U2709 ( .A(n2542), .B(n2541), .Z(n2546) );
  NAND U2710 ( .A(n2544), .B(n2543), .Z(n2545) );
  NAND U2711 ( .A(n2546), .B(n2545), .Z(n2626) );
  XNOR U2712 ( .A(n2625), .B(n2626), .Z(n2627) );
  XOR U2713 ( .A(n2628), .B(n2627), .Z(n2558) );
  NANDN U2714 ( .A(n2548), .B(n2547), .Z(n2552) );
  NANDN U2715 ( .A(n2550), .B(n2549), .Z(n2551) );
  NAND U2716 ( .A(n2552), .B(n2551), .Z(n2559) );
  XNOR U2717 ( .A(n2558), .B(n2559), .Z(n2560) );
  XNOR U2718 ( .A(n2561), .B(n2560), .Z(n2631) );
  XNOR U2719 ( .A(n2631), .B(sreg[279]), .Z(n2633) );
  NAND U2720 ( .A(n2553), .B(sreg[278]), .Z(n2557) );
  OR U2721 ( .A(n2555), .B(n2554), .Z(n2556) );
  AND U2722 ( .A(n2557), .B(n2556), .Z(n2632) );
  XOR U2723 ( .A(n2633), .B(n2632), .Z(c[279]) );
  NANDN U2724 ( .A(n2559), .B(n2558), .Z(n2563) );
  NAND U2725 ( .A(n2561), .B(n2560), .Z(n2562) );
  NAND U2726 ( .A(n2563), .B(n2562), .Z(n2639) );
  NANDN U2727 ( .A(n2565), .B(n2564), .Z(n2569) );
  OR U2728 ( .A(n2567), .B(n2566), .Z(n2568) );
  NAND U2729 ( .A(n2569), .B(n2568), .Z(n2706) );
  NANDN U2730 ( .A(n2571), .B(n2570), .Z(n2575) );
  OR U2731 ( .A(n2573), .B(n2572), .Z(n2574) );
  NAND U2732 ( .A(n2575), .B(n2574), .Z(n2694) );
  NAND U2733 ( .A(b[0]), .B(a[40]), .Z(n2576) );
  XNOR U2734 ( .A(b[1]), .B(n2576), .Z(n2578) );
  NAND U2735 ( .A(a[39]), .B(n98), .Z(n2577) );
  AND U2736 ( .A(n2578), .B(n2577), .Z(n2670) );
  XNOR U2737 ( .A(n20154), .B(n2729), .Z(n2676) );
  OR U2738 ( .A(n2676), .B(n20057), .Z(n2581) );
  NANDN U2739 ( .A(n2579), .B(n20098), .Z(n2580) );
  AND U2740 ( .A(n2581), .B(n2580), .Z(n2671) );
  XOR U2741 ( .A(n2670), .B(n2671), .Z(n2673) );
  NAND U2742 ( .A(a[24]), .B(b[15]), .Z(n2672) );
  XOR U2743 ( .A(n2673), .B(n2672), .Z(n2691) );
  NAND U2744 ( .A(n19722), .B(n2582), .Z(n2584) );
  XNOR U2745 ( .A(b[5]), .B(n3353), .Z(n2682) );
  NANDN U2746 ( .A(n19640), .B(n2682), .Z(n2583) );
  NAND U2747 ( .A(n2584), .B(n2583), .Z(n2667) );
  XNOR U2748 ( .A(n19714), .B(n3224), .Z(n2685) );
  NANDN U2749 ( .A(n2685), .B(n19766), .Z(n2587) );
  NANDN U2750 ( .A(n2585), .B(n19767), .Z(n2586) );
  NAND U2751 ( .A(n2587), .B(n2586), .Z(n2664) );
  NAND U2752 ( .A(n19554), .B(n2588), .Z(n2590) );
  IV U2753 ( .A(a[38]), .Z(n3536) );
  XNOR U2754 ( .A(b[3]), .B(n3536), .Z(n2688) );
  NANDN U2755 ( .A(n19521), .B(n2688), .Z(n2589) );
  AND U2756 ( .A(n2590), .B(n2589), .Z(n2665) );
  XNOR U2757 ( .A(n2664), .B(n2665), .Z(n2666) );
  XOR U2758 ( .A(n2667), .B(n2666), .Z(n2692) );
  XOR U2759 ( .A(n2691), .B(n2692), .Z(n2693) );
  XNOR U2760 ( .A(n2694), .B(n2693), .Z(n2642) );
  NAND U2761 ( .A(n2592), .B(n2591), .Z(n2596) );
  NAND U2762 ( .A(n2594), .B(n2593), .Z(n2595) );
  NAND U2763 ( .A(n2596), .B(n2595), .Z(n2643) );
  XOR U2764 ( .A(n2642), .B(n2643), .Z(n2645) );
  XNOR U2765 ( .A(n20052), .B(n2885), .Z(n2648) );
  OR U2766 ( .A(n2648), .B(n20020), .Z(n2599) );
  NANDN U2767 ( .A(n2597), .B(n19960), .Z(n2598) );
  NAND U2768 ( .A(n2599), .B(n2598), .Z(n2661) );
  XNOR U2769 ( .A(n102), .B(n2600), .Z(n2652) );
  OR U2770 ( .A(n2652), .B(n20121), .Z(n2603) );
  NANDN U2771 ( .A(n2601), .B(n20122), .Z(n2602) );
  NAND U2772 ( .A(n2603), .B(n2602), .Z(n2658) );
  XNOR U2773 ( .A(n19975), .B(n3068), .Z(n2655) );
  NANDN U2774 ( .A(n2655), .B(n19883), .Z(n2606) );
  NANDN U2775 ( .A(n2604), .B(n19937), .Z(n2605) );
  AND U2776 ( .A(n2606), .B(n2605), .Z(n2659) );
  XNOR U2777 ( .A(n2658), .B(n2659), .Z(n2660) );
  XNOR U2778 ( .A(n2661), .B(n2660), .Z(n2697) );
  NANDN U2779 ( .A(n2608), .B(n2607), .Z(n2612) );
  NAND U2780 ( .A(n2610), .B(n2609), .Z(n2611) );
  NAND U2781 ( .A(n2612), .B(n2611), .Z(n2698) );
  XNOR U2782 ( .A(n2697), .B(n2698), .Z(n2699) );
  NANDN U2783 ( .A(n2614), .B(n2613), .Z(n2618) );
  NAND U2784 ( .A(n2616), .B(n2615), .Z(n2617) );
  AND U2785 ( .A(n2618), .B(n2617), .Z(n2700) );
  XNOR U2786 ( .A(n2699), .B(n2700), .Z(n2644) );
  XNOR U2787 ( .A(n2645), .B(n2644), .Z(n2703) );
  NANDN U2788 ( .A(n2620), .B(n2619), .Z(n2624) );
  NAND U2789 ( .A(n2622), .B(n2621), .Z(n2623) );
  NAND U2790 ( .A(n2624), .B(n2623), .Z(n2704) );
  XNOR U2791 ( .A(n2703), .B(n2704), .Z(n2705) );
  XOR U2792 ( .A(n2706), .B(n2705), .Z(n2636) );
  NANDN U2793 ( .A(n2626), .B(n2625), .Z(n2630) );
  NANDN U2794 ( .A(n2628), .B(n2627), .Z(n2629) );
  NAND U2795 ( .A(n2630), .B(n2629), .Z(n2637) );
  XNOR U2796 ( .A(n2636), .B(n2637), .Z(n2638) );
  XNOR U2797 ( .A(n2639), .B(n2638), .Z(n2709) );
  XNOR U2798 ( .A(n2709), .B(sreg[280]), .Z(n2711) );
  NAND U2799 ( .A(n2631), .B(sreg[279]), .Z(n2635) );
  OR U2800 ( .A(n2633), .B(n2632), .Z(n2634) );
  AND U2801 ( .A(n2635), .B(n2634), .Z(n2710) );
  XOR U2802 ( .A(n2711), .B(n2710), .Z(c[280]) );
  NANDN U2803 ( .A(n2637), .B(n2636), .Z(n2641) );
  NAND U2804 ( .A(n2639), .B(n2638), .Z(n2640) );
  NAND U2805 ( .A(n2641), .B(n2640), .Z(n2717) );
  NANDN U2806 ( .A(n2643), .B(n2642), .Z(n2647) );
  OR U2807 ( .A(n2645), .B(n2644), .Z(n2646) );
  NAND U2808 ( .A(n2647), .B(n2646), .Z(n2784) );
  XNOR U2809 ( .A(n20052), .B(n2963), .Z(n2726) );
  OR U2810 ( .A(n2726), .B(n20020), .Z(n2650) );
  NANDN U2811 ( .A(n2648), .B(n19960), .Z(n2649) );
  NAND U2812 ( .A(n2650), .B(n2649), .Z(n2739) );
  XNOR U2813 ( .A(n102), .B(n2651), .Z(n2730) );
  OR U2814 ( .A(n2730), .B(n20121), .Z(n2654) );
  NANDN U2815 ( .A(n2652), .B(n20122), .Z(n2653) );
  NAND U2816 ( .A(n2654), .B(n2653), .Z(n2736) );
  XNOR U2817 ( .A(n19975), .B(n3146), .Z(n2733) );
  NANDN U2818 ( .A(n2733), .B(n19883), .Z(n2657) );
  NANDN U2819 ( .A(n2655), .B(n19937), .Z(n2656) );
  AND U2820 ( .A(n2657), .B(n2656), .Z(n2737) );
  XNOR U2821 ( .A(n2736), .B(n2737), .Z(n2738) );
  XNOR U2822 ( .A(n2739), .B(n2738), .Z(n2775) );
  NANDN U2823 ( .A(n2659), .B(n2658), .Z(n2663) );
  NAND U2824 ( .A(n2661), .B(n2660), .Z(n2662) );
  NAND U2825 ( .A(n2663), .B(n2662), .Z(n2776) );
  XNOR U2826 ( .A(n2775), .B(n2776), .Z(n2777) );
  NANDN U2827 ( .A(n2665), .B(n2664), .Z(n2669) );
  NAND U2828 ( .A(n2667), .B(n2666), .Z(n2668) );
  AND U2829 ( .A(n2669), .B(n2668), .Z(n2778) );
  XNOR U2830 ( .A(n2777), .B(n2778), .Z(n2722) );
  NANDN U2831 ( .A(n2671), .B(n2670), .Z(n2675) );
  OR U2832 ( .A(n2673), .B(n2672), .Z(n2674) );
  NAND U2833 ( .A(n2675), .B(n2674), .Z(n2772) );
  XNOR U2834 ( .A(n20154), .B(n2807), .Z(n2757) );
  OR U2835 ( .A(n2757), .B(n20057), .Z(n2678) );
  NANDN U2836 ( .A(n2676), .B(n20098), .Z(n2677) );
  AND U2837 ( .A(n2678), .B(n2677), .Z(n2749) );
  NAND U2838 ( .A(b[0]), .B(a[41]), .Z(n2679) );
  XNOR U2839 ( .A(b[1]), .B(n2679), .Z(n2681) );
  NAND U2840 ( .A(a[40]), .B(n98), .Z(n2680) );
  AND U2841 ( .A(n2681), .B(n2680), .Z(n2748) );
  XOR U2842 ( .A(n2749), .B(n2748), .Z(n2751) );
  NAND U2843 ( .A(a[25]), .B(b[15]), .Z(n2750) );
  XOR U2844 ( .A(n2751), .B(n2750), .Z(n2769) );
  NAND U2845 ( .A(n19722), .B(n2682), .Z(n2684) );
  XNOR U2846 ( .A(b[5]), .B(n3458), .Z(n2760) );
  NANDN U2847 ( .A(n19640), .B(n2760), .Z(n2683) );
  NAND U2848 ( .A(n2684), .B(n2683), .Z(n2745) );
  XNOR U2849 ( .A(n19714), .B(n3275), .Z(n2763) );
  NANDN U2850 ( .A(n2763), .B(n19766), .Z(n2687) );
  NANDN U2851 ( .A(n2685), .B(n19767), .Z(n2686) );
  NAND U2852 ( .A(n2687), .B(n2686), .Z(n2742) );
  NAND U2853 ( .A(n19554), .B(n2688), .Z(n2690) );
  IV U2854 ( .A(a[39]), .Z(n3587) );
  XNOR U2855 ( .A(b[3]), .B(n3587), .Z(n2766) );
  NANDN U2856 ( .A(n19521), .B(n2766), .Z(n2689) );
  AND U2857 ( .A(n2690), .B(n2689), .Z(n2743) );
  XNOR U2858 ( .A(n2742), .B(n2743), .Z(n2744) );
  XOR U2859 ( .A(n2745), .B(n2744), .Z(n2770) );
  XOR U2860 ( .A(n2769), .B(n2770), .Z(n2771) );
  XNOR U2861 ( .A(n2772), .B(n2771), .Z(n2720) );
  NAND U2862 ( .A(n2692), .B(n2691), .Z(n2696) );
  NAND U2863 ( .A(n2694), .B(n2693), .Z(n2695) );
  NAND U2864 ( .A(n2696), .B(n2695), .Z(n2721) );
  XOR U2865 ( .A(n2720), .B(n2721), .Z(n2723) );
  XNOR U2866 ( .A(n2722), .B(n2723), .Z(n2781) );
  NANDN U2867 ( .A(n2698), .B(n2697), .Z(n2702) );
  NAND U2868 ( .A(n2700), .B(n2699), .Z(n2701) );
  NAND U2869 ( .A(n2702), .B(n2701), .Z(n2782) );
  XNOR U2870 ( .A(n2781), .B(n2782), .Z(n2783) );
  XOR U2871 ( .A(n2784), .B(n2783), .Z(n2714) );
  NANDN U2872 ( .A(n2704), .B(n2703), .Z(n2708) );
  NANDN U2873 ( .A(n2706), .B(n2705), .Z(n2707) );
  NAND U2874 ( .A(n2708), .B(n2707), .Z(n2715) );
  XNOR U2875 ( .A(n2714), .B(n2715), .Z(n2716) );
  XNOR U2876 ( .A(n2717), .B(n2716), .Z(n2787) );
  XNOR U2877 ( .A(n2787), .B(sreg[281]), .Z(n2789) );
  NAND U2878 ( .A(n2709), .B(sreg[280]), .Z(n2713) );
  OR U2879 ( .A(n2711), .B(n2710), .Z(n2712) );
  AND U2880 ( .A(n2713), .B(n2712), .Z(n2788) );
  XOR U2881 ( .A(n2789), .B(n2788), .Z(c[281]) );
  NANDN U2882 ( .A(n2715), .B(n2714), .Z(n2719) );
  NAND U2883 ( .A(n2717), .B(n2716), .Z(n2718) );
  NAND U2884 ( .A(n2719), .B(n2718), .Z(n2795) );
  NANDN U2885 ( .A(n2721), .B(n2720), .Z(n2725) );
  OR U2886 ( .A(n2723), .B(n2722), .Z(n2724) );
  NAND U2887 ( .A(n2725), .B(n2724), .Z(n2862) );
  XNOR U2888 ( .A(n20052), .B(n3068), .Z(n2804) );
  OR U2889 ( .A(n2804), .B(n20020), .Z(n2728) );
  NANDN U2890 ( .A(n2726), .B(n19960), .Z(n2727) );
  NAND U2891 ( .A(n2728), .B(n2727), .Z(n2817) );
  XNOR U2892 ( .A(n102), .B(n2729), .Z(n2808) );
  OR U2893 ( .A(n2808), .B(n20121), .Z(n2732) );
  NANDN U2894 ( .A(n2730), .B(n20122), .Z(n2731) );
  NAND U2895 ( .A(n2732), .B(n2731), .Z(n2814) );
  XNOR U2896 ( .A(n19975), .B(n3224), .Z(n2811) );
  NANDN U2897 ( .A(n2811), .B(n19883), .Z(n2735) );
  NANDN U2898 ( .A(n2733), .B(n19937), .Z(n2734) );
  AND U2899 ( .A(n2735), .B(n2734), .Z(n2815) );
  XNOR U2900 ( .A(n2814), .B(n2815), .Z(n2816) );
  XNOR U2901 ( .A(n2817), .B(n2816), .Z(n2853) );
  NANDN U2902 ( .A(n2737), .B(n2736), .Z(n2741) );
  NAND U2903 ( .A(n2739), .B(n2738), .Z(n2740) );
  NAND U2904 ( .A(n2741), .B(n2740), .Z(n2854) );
  XNOR U2905 ( .A(n2853), .B(n2854), .Z(n2855) );
  NANDN U2906 ( .A(n2743), .B(n2742), .Z(n2747) );
  NAND U2907 ( .A(n2745), .B(n2744), .Z(n2746) );
  AND U2908 ( .A(n2747), .B(n2746), .Z(n2856) );
  XNOR U2909 ( .A(n2855), .B(n2856), .Z(n2800) );
  NANDN U2910 ( .A(n2749), .B(n2748), .Z(n2753) );
  OR U2911 ( .A(n2751), .B(n2750), .Z(n2752) );
  NAND U2912 ( .A(n2753), .B(n2752), .Z(n2850) );
  NAND U2913 ( .A(b[0]), .B(a[42]), .Z(n2754) );
  XNOR U2914 ( .A(b[1]), .B(n2754), .Z(n2756) );
  NAND U2915 ( .A(a[41]), .B(n98), .Z(n2755) );
  AND U2916 ( .A(n2756), .B(n2755), .Z(n2826) );
  XNOR U2917 ( .A(n20154), .B(n2885), .Z(n2835) );
  OR U2918 ( .A(n2835), .B(n20057), .Z(n2759) );
  NANDN U2919 ( .A(n2757), .B(n20098), .Z(n2758) );
  AND U2920 ( .A(n2759), .B(n2758), .Z(n2827) );
  XOR U2921 ( .A(n2826), .B(n2827), .Z(n2829) );
  NAND U2922 ( .A(a[26]), .B(b[15]), .Z(n2828) );
  XOR U2923 ( .A(n2829), .B(n2828), .Z(n2847) );
  NAND U2924 ( .A(n19722), .B(n2760), .Z(n2762) );
  XNOR U2925 ( .A(b[5]), .B(n3536), .Z(n2838) );
  NANDN U2926 ( .A(n19640), .B(n2838), .Z(n2761) );
  NAND U2927 ( .A(n2762), .B(n2761), .Z(n2823) );
  XNOR U2928 ( .A(n19714), .B(n3353), .Z(n2841) );
  NANDN U2929 ( .A(n2841), .B(n19766), .Z(n2765) );
  NANDN U2930 ( .A(n2763), .B(n19767), .Z(n2764) );
  NAND U2931 ( .A(n2765), .B(n2764), .Z(n2820) );
  NAND U2932 ( .A(n19554), .B(n2766), .Z(n2768) );
  IV U2933 ( .A(a[40]), .Z(n3692) );
  XNOR U2934 ( .A(b[3]), .B(n3692), .Z(n2844) );
  NANDN U2935 ( .A(n19521), .B(n2844), .Z(n2767) );
  AND U2936 ( .A(n2768), .B(n2767), .Z(n2821) );
  XNOR U2937 ( .A(n2820), .B(n2821), .Z(n2822) );
  XOR U2938 ( .A(n2823), .B(n2822), .Z(n2848) );
  XOR U2939 ( .A(n2847), .B(n2848), .Z(n2849) );
  XNOR U2940 ( .A(n2850), .B(n2849), .Z(n2798) );
  NAND U2941 ( .A(n2770), .B(n2769), .Z(n2774) );
  NAND U2942 ( .A(n2772), .B(n2771), .Z(n2773) );
  NAND U2943 ( .A(n2774), .B(n2773), .Z(n2799) );
  XOR U2944 ( .A(n2798), .B(n2799), .Z(n2801) );
  XNOR U2945 ( .A(n2800), .B(n2801), .Z(n2859) );
  NANDN U2946 ( .A(n2776), .B(n2775), .Z(n2780) );
  NAND U2947 ( .A(n2778), .B(n2777), .Z(n2779) );
  NAND U2948 ( .A(n2780), .B(n2779), .Z(n2860) );
  XNOR U2949 ( .A(n2859), .B(n2860), .Z(n2861) );
  XOR U2950 ( .A(n2862), .B(n2861), .Z(n2792) );
  NANDN U2951 ( .A(n2782), .B(n2781), .Z(n2786) );
  NANDN U2952 ( .A(n2784), .B(n2783), .Z(n2785) );
  NAND U2953 ( .A(n2786), .B(n2785), .Z(n2793) );
  XNOR U2954 ( .A(n2792), .B(n2793), .Z(n2794) );
  XNOR U2955 ( .A(n2795), .B(n2794), .Z(n2865) );
  XNOR U2956 ( .A(n2865), .B(sreg[282]), .Z(n2867) );
  NAND U2957 ( .A(n2787), .B(sreg[281]), .Z(n2791) );
  OR U2958 ( .A(n2789), .B(n2788), .Z(n2790) );
  AND U2959 ( .A(n2791), .B(n2790), .Z(n2866) );
  XOR U2960 ( .A(n2867), .B(n2866), .Z(c[282]) );
  NANDN U2961 ( .A(n2793), .B(n2792), .Z(n2797) );
  NAND U2962 ( .A(n2795), .B(n2794), .Z(n2796) );
  NAND U2963 ( .A(n2797), .B(n2796), .Z(n2873) );
  NANDN U2964 ( .A(n2799), .B(n2798), .Z(n2803) );
  OR U2965 ( .A(n2801), .B(n2800), .Z(n2802) );
  NAND U2966 ( .A(n2803), .B(n2802), .Z(n2940) );
  XNOR U2967 ( .A(n20052), .B(n3146), .Z(n2882) );
  OR U2968 ( .A(n2882), .B(n20020), .Z(n2806) );
  NANDN U2969 ( .A(n2804), .B(n19960), .Z(n2805) );
  NAND U2970 ( .A(n2806), .B(n2805), .Z(n2895) );
  XNOR U2971 ( .A(n102), .B(n2807), .Z(n2886) );
  OR U2972 ( .A(n2886), .B(n20121), .Z(n2810) );
  NANDN U2973 ( .A(n2808), .B(n20122), .Z(n2809) );
  NAND U2974 ( .A(n2810), .B(n2809), .Z(n2892) );
  XNOR U2975 ( .A(n19975), .B(n3275), .Z(n2889) );
  NANDN U2976 ( .A(n2889), .B(n19883), .Z(n2813) );
  NANDN U2977 ( .A(n2811), .B(n19937), .Z(n2812) );
  AND U2978 ( .A(n2813), .B(n2812), .Z(n2893) );
  XNOR U2979 ( .A(n2892), .B(n2893), .Z(n2894) );
  XNOR U2980 ( .A(n2895), .B(n2894), .Z(n2931) );
  NANDN U2981 ( .A(n2815), .B(n2814), .Z(n2819) );
  NAND U2982 ( .A(n2817), .B(n2816), .Z(n2818) );
  NAND U2983 ( .A(n2819), .B(n2818), .Z(n2932) );
  XNOR U2984 ( .A(n2931), .B(n2932), .Z(n2933) );
  NANDN U2985 ( .A(n2821), .B(n2820), .Z(n2825) );
  NAND U2986 ( .A(n2823), .B(n2822), .Z(n2824) );
  AND U2987 ( .A(n2825), .B(n2824), .Z(n2934) );
  XNOR U2988 ( .A(n2933), .B(n2934), .Z(n2878) );
  NANDN U2989 ( .A(n2827), .B(n2826), .Z(n2831) );
  OR U2990 ( .A(n2829), .B(n2828), .Z(n2830) );
  NAND U2991 ( .A(n2831), .B(n2830), .Z(n2928) );
  NAND U2992 ( .A(b[0]), .B(a[43]), .Z(n2832) );
  XNOR U2993 ( .A(b[1]), .B(n2832), .Z(n2834) );
  NAND U2994 ( .A(a[42]), .B(n98), .Z(n2833) );
  AND U2995 ( .A(n2834), .B(n2833), .Z(n2904) );
  XNOR U2996 ( .A(n20154), .B(n2963), .Z(n2910) );
  OR U2997 ( .A(n2910), .B(n20057), .Z(n2837) );
  NANDN U2998 ( .A(n2835), .B(n20098), .Z(n2836) );
  AND U2999 ( .A(n2837), .B(n2836), .Z(n2905) );
  XOR U3000 ( .A(n2904), .B(n2905), .Z(n2907) );
  NAND U3001 ( .A(a[27]), .B(b[15]), .Z(n2906) );
  XOR U3002 ( .A(n2907), .B(n2906), .Z(n2925) );
  NAND U3003 ( .A(n19722), .B(n2838), .Z(n2840) );
  XNOR U3004 ( .A(b[5]), .B(n3587), .Z(n2916) );
  NANDN U3005 ( .A(n19640), .B(n2916), .Z(n2839) );
  NAND U3006 ( .A(n2840), .B(n2839), .Z(n2901) );
  XNOR U3007 ( .A(n19714), .B(n3458), .Z(n2919) );
  NANDN U3008 ( .A(n2919), .B(n19766), .Z(n2843) );
  NANDN U3009 ( .A(n2841), .B(n19767), .Z(n2842) );
  NAND U3010 ( .A(n2843), .B(n2842), .Z(n2898) );
  NAND U3011 ( .A(n19554), .B(n2844), .Z(n2846) );
  IV U3012 ( .A(a[41]), .Z(n3743) );
  XNOR U3013 ( .A(b[3]), .B(n3743), .Z(n2922) );
  NANDN U3014 ( .A(n19521), .B(n2922), .Z(n2845) );
  AND U3015 ( .A(n2846), .B(n2845), .Z(n2899) );
  XNOR U3016 ( .A(n2898), .B(n2899), .Z(n2900) );
  XOR U3017 ( .A(n2901), .B(n2900), .Z(n2926) );
  XOR U3018 ( .A(n2925), .B(n2926), .Z(n2927) );
  XNOR U3019 ( .A(n2928), .B(n2927), .Z(n2876) );
  NAND U3020 ( .A(n2848), .B(n2847), .Z(n2852) );
  NAND U3021 ( .A(n2850), .B(n2849), .Z(n2851) );
  NAND U3022 ( .A(n2852), .B(n2851), .Z(n2877) );
  XOR U3023 ( .A(n2876), .B(n2877), .Z(n2879) );
  XNOR U3024 ( .A(n2878), .B(n2879), .Z(n2937) );
  NANDN U3025 ( .A(n2854), .B(n2853), .Z(n2858) );
  NAND U3026 ( .A(n2856), .B(n2855), .Z(n2857) );
  NAND U3027 ( .A(n2858), .B(n2857), .Z(n2938) );
  XNOR U3028 ( .A(n2937), .B(n2938), .Z(n2939) );
  XOR U3029 ( .A(n2940), .B(n2939), .Z(n2870) );
  NANDN U3030 ( .A(n2860), .B(n2859), .Z(n2864) );
  NANDN U3031 ( .A(n2862), .B(n2861), .Z(n2863) );
  NAND U3032 ( .A(n2864), .B(n2863), .Z(n2871) );
  XNOR U3033 ( .A(n2870), .B(n2871), .Z(n2872) );
  XNOR U3034 ( .A(n2873), .B(n2872), .Z(n2943) );
  XNOR U3035 ( .A(n2943), .B(sreg[283]), .Z(n2945) );
  NAND U3036 ( .A(n2865), .B(sreg[282]), .Z(n2869) );
  OR U3037 ( .A(n2867), .B(n2866), .Z(n2868) );
  AND U3038 ( .A(n2869), .B(n2868), .Z(n2944) );
  XOR U3039 ( .A(n2945), .B(n2944), .Z(c[283]) );
  NANDN U3040 ( .A(n2871), .B(n2870), .Z(n2875) );
  NAND U3041 ( .A(n2873), .B(n2872), .Z(n2874) );
  NAND U3042 ( .A(n2875), .B(n2874), .Z(n2951) );
  NANDN U3043 ( .A(n2877), .B(n2876), .Z(n2881) );
  OR U3044 ( .A(n2879), .B(n2878), .Z(n2880) );
  NAND U3045 ( .A(n2881), .B(n2880), .Z(n3018) );
  XNOR U3046 ( .A(n20052), .B(n3224), .Z(n2960) );
  OR U3047 ( .A(n2960), .B(n20020), .Z(n2884) );
  NANDN U3048 ( .A(n2882), .B(n19960), .Z(n2883) );
  NAND U3049 ( .A(n2884), .B(n2883), .Z(n2973) );
  XNOR U3050 ( .A(n102), .B(n2885), .Z(n2964) );
  OR U3051 ( .A(n2964), .B(n20121), .Z(n2888) );
  NANDN U3052 ( .A(n2886), .B(n20122), .Z(n2887) );
  NAND U3053 ( .A(n2888), .B(n2887), .Z(n2970) );
  XNOR U3054 ( .A(n19975), .B(n3353), .Z(n2967) );
  NANDN U3055 ( .A(n2967), .B(n19883), .Z(n2891) );
  NANDN U3056 ( .A(n2889), .B(n19937), .Z(n2890) );
  AND U3057 ( .A(n2891), .B(n2890), .Z(n2971) );
  XNOR U3058 ( .A(n2970), .B(n2971), .Z(n2972) );
  XNOR U3059 ( .A(n2973), .B(n2972), .Z(n3009) );
  NANDN U3060 ( .A(n2893), .B(n2892), .Z(n2897) );
  NAND U3061 ( .A(n2895), .B(n2894), .Z(n2896) );
  NAND U3062 ( .A(n2897), .B(n2896), .Z(n3010) );
  XNOR U3063 ( .A(n3009), .B(n3010), .Z(n3011) );
  NANDN U3064 ( .A(n2899), .B(n2898), .Z(n2903) );
  NAND U3065 ( .A(n2901), .B(n2900), .Z(n2902) );
  AND U3066 ( .A(n2903), .B(n2902), .Z(n3012) );
  XNOR U3067 ( .A(n3011), .B(n3012), .Z(n2956) );
  NANDN U3068 ( .A(n2905), .B(n2904), .Z(n2909) );
  OR U3069 ( .A(n2907), .B(n2906), .Z(n2908) );
  NAND U3070 ( .A(n2909), .B(n2908), .Z(n3006) );
  XNOR U3071 ( .A(n20154), .B(n3068), .Z(n2991) );
  OR U3072 ( .A(n2991), .B(n20057), .Z(n2912) );
  NANDN U3073 ( .A(n2910), .B(n20098), .Z(n2911) );
  AND U3074 ( .A(n2912), .B(n2911), .Z(n2983) );
  NAND U3075 ( .A(b[0]), .B(a[44]), .Z(n2913) );
  XNOR U3076 ( .A(b[1]), .B(n2913), .Z(n2915) );
  NAND U3077 ( .A(a[43]), .B(n98), .Z(n2914) );
  AND U3078 ( .A(n2915), .B(n2914), .Z(n2982) );
  XOR U3079 ( .A(n2983), .B(n2982), .Z(n2985) );
  NAND U3080 ( .A(a[28]), .B(b[15]), .Z(n2984) );
  XOR U3081 ( .A(n2985), .B(n2984), .Z(n3003) );
  NAND U3082 ( .A(n19722), .B(n2916), .Z(n2918) );
  XNOR U3083 ( .A(b[5]), .B(n3692), .Z(n2994) );
  NANDN U3084 ( .A(n19640), .B(n2994), .Z(n2917) );
  NAND U3085 ( .A(n2918), .B(n2917), .Z(n2979) );
  XNOR U3086 ( .A(n19714), .B(n3536), .Z(n2997) );
  NANDN U3087 ( .A(n2997), .B(n19766), .Z(n2921) );
  NANDN U3088 ( .A(n2919), .B(n19767), .Z(n2920) );
  NAND U3089 ( .A(n2921), .B(n2920), .Z(n2976) );
  NAND U3090 ( .A(n19554), .B(n2922), .Z(n2924) );
  IV U3091 ( .A(a[42]), .Z(n3848) );
  XNOR U3092 ( .A(b[3]), .B(n3848), .Z(n3000) );
  NANDN U3093 ( .A(n19521), .B(n3000), .Z(n2923) );
  AND U3094 ( .A(n2924), .B(n2923), .Z(n2977) );
  XNOR U3095 ( .A(n2976), .B(n2977), .Z(n2978) );
  XOR U3096 ( .A(n2979), .B(n2978), .Z(n3004) );
  XOR U3097 ( .A(n3003), .B(n3004), .Z(n3005) );
  XNOR U3098 ( .A(n3006), .B(n3005), .Z(n2954) );
  NAND U3099 ( .A(n2926), .B(n2925), .Z(n2930) );
  NAND U3100 ( .A(n2928), .B(n2927), .Z(n2929) );
  NAND U3101 ( .A(n2930), .B(n2929), .Z(n2955) );
  XOR U3102 ( .A(n2954), .B(n2955), .Z(n2957) );
  XNOR U3103 ( .A(n2956), .B(n2957), .Z(n3015) );
  NANDN U3104 ( .A(n2932), .B(n2931), .Z(n2936) );
  NAND U3105 ( .A(n2934), .B(n2933), .Z(n2935) );
  NAND U3106 ( .A(n2936), .B(n2935), .Z(n3016) );
  XNOR U3107 ( .A(n3015), .B(n3016), .Z(n3017) );
  XOR U3108 ( .A(n3018), .B(n3017), .Z(n2948) );
  NANDN U3109 ( .A(n2938), .B(n2937), .Z(n2942) );
  NANDN U3110 ( .A(n2940), .B(n2939), .Z(n2941) );
  NAND U3111 ( .A(n2942), .B(n2941), .Z(n2949) );
  XNOR U3112 ( .A(n2948), .B(n2949), .Z(n2950) );
  XNOR U3113 ( .A(n2951), .B(n2950), .Z(n3021) );
  XNOR U3114 ( .A(n3021), .B(sreg[284]), .Z(n3023) );
  NAND U3115 ( .A(n2943), .B(sreg[283]), .Z(n2947) );
  OR U3116 ( .A(n2945), .B(n2944), .Z(n2946) );
  AND U3117 ( .A(n2947), .B(n2946), .Z(n3022) );
  XOR U3118 ( .A(n3023), .B(n3022), .Z(c[284]) );
  NANDN U3119 ( .A(n2949), .B(n2948), .Z(n2953) );
  NAND U3120 ( .A(n2951), .B(n2950), .Z(n2952) );
  NAND U3121 ( .A(n2953), .B(n2952), .Z(n3029) );
  NANDN U3122 ( .A(n2955), .B(n2954), .Z(n2959) );
  OR U3123 ( .A(n2957), .B(n2956), .Z(n2958) );
  NAND U3124 ( .A(n2959), .B(n2958), .Z(n3096) );
  XNOR U3125 ( .A(n20052), .B(n3275), .Z(n3065) );
  OR U3126 ( .A(n3065), .B(n20020), .Z(n2962) );
  NANDN U3127 ( .A(n2960), .B(n19960), .Z(n2961) );
  NAND U3128 ( .A(n2962), .B(n2961), .Z(n3078) );
  XNOR U3129 ( .A(n102), .B(n2963), .Z(n3069) );
  OR U3130 ( .A(n3069), .B(n20121), .Z(n2966) );
  NANDN U3131 ( .A(n2964), .B(n20122), .Z(n2965) );
  NAND U3132 ( .A(n2966), .B(n2965), .Z(n3075) );
  XNOR U3133 ( .A(n19975), .B(n3458), .Z(n3072) );
  NANDN U3134 ( .A(n3072), .B(n19883), .Z(n2969) );
  NANDN U3135 ( .A(n2967), .B(n19937), .Z(n2968) );
  AND U3136 ( .A(n2969), .B(n2968), .Z(n3076) );
  XNOR U3137 ( .A(n3075), .B(n3076), .Z(n3077) );
  XNOR U3138 ( .A(n3078), .B(n3077), .Z(n3087) );
  NANDN U3139 ( .A(n2971), .B(n2970), .Z(n2975) );
  NAND U3140 ( .A(n2973), .B(n2972), .Z(n2974) );
  NAND U3141 ( .A(n2975), .B(n2974), .Z(n3088) );
  XNOR U3142 ( .A(n3087), .B(n3088), .Z(n3089) );
  NANDN U3143 ( .A(n2977), .B(n2976), .Z(n2981) );
  NAND U3144 ( .A(n2979), .B(n2978), .Z(n2980) );
  AND U3145 ( .A(n2981), .B(n2980), .Z(n3090) );
  XNOR U3146 ( .A(n3089), .B(n3090), .Z(n3034) );
  NANDN U3147 ( .A(n2983), .B(n2982), .Z(n2987) );
  OR U3148 ( .A(n2985), .B(n2984), .Z(n2986) );
  NAND U3149 ( .A(n2987), .B(n2986), .Z(n3062) );
  NAND U3150 ( .A(b[0]), .B(a[45]), .Z(n2988) );
  XNOR U3151 ( .A(b[1]), .B(n2988), .Z(n2990) );
  NAND U3152 ( .A(a[44]), .B(n98), .Z(n2989) );
  AND U3153 ( .A(n2990), .B(n2989), .Z(n3038) );
  XNOR U3154 ( .A(n20154), .B(n3146), .Z(n3047) );
  OR U3155 ( .A(n3047), .B(n20057), .Z(n2993) );
  NANDN U3156 ( .A(n2991), .B(n20098), .Z(n2992) );
  AND U3157 ( .A(n2993), .B(n2992), .Z(n3039) );
  XOR U3158 ( .A(n3038), .B(n3039), .Z(n3041) );
  NAND U3159 ( .A(a[29]), .B(b[15]), .Z(n3040) );
  XOR U3160 ( .A(n3041), .B(n3040), .Z(n3059) );
  NAND U3161 ( .A(n19722), .B(n2994), .Z(n2996) );
  XNOR U3162 ( .A(b[5]), .B(n3743), .Z(n3050) );
  NANDN U3163 ( .A(n19640), .B(n3050), .Z(n2995) );
  NAND U3164 ( .A(n2996), .B(n2995), .Z(n3084) );
  XNOR U3165 ( .A(n19714), .B(n3587), .Z(n3053) );
  NANDN U3166 ( .A(n3053), .B(n19766), .Z(n2999) );
  NANDN U3167 ( .A(n2997), .B(n19767), .Z(n2998) );
  NAND U3168 ( .A(n2999), .B(n2998), .Z(n3081) );
  NAND U3169 ( .A(n19554), .B(n3000), .Z(n3002) );
  IV U3170 ( .A(a[43]), .Z(n3926) );
  XNOR U3171 ( .A(b[3]), .B(n3926), .Z(n3056) );
  NANDN U3172 ( .A(n19521), .B(n3056), .Z(n3001) );
  AND U3173 ( .A(n3002), .B(n3001), .Z(n3082) );
  XNOR U3174 ( .A(n3081), .B(n3082), .Z(n3083) );
  XOR U3175 ( .A(n3084), .B(n3083), .Z(n3060) );
  XOR U3176 ( .A(n3059), .B(n3060), .Z(n3061) );
  XNOR U3177 ( .A(n3062), .B(n3061), .Z(n3032) );
  NAND U3178 ( .A(n3004), .B(n3003), .Z(n3008) );
  NAND U3179 ( .A(n3006), .B(n3005), .Z(n3007) );
  NAND U3180 ( .A(n3008), .B(n3007), .Z(n3033) );
  XOR U3181 ( .A(n3032), .B(n3033), .Z(n3035) );
  XNOR U3182 ( .A(n3034), .B(n3035), .Z(n3093) );
  NANDN U3183 ( .A(n3010), .B(n3009), .Z(n3014) );
  NAND U3184 ( .A(n3012), .B(n3011), .Z(n3013) );
  NAND U3185 ( .A(n3014), .B(n3013), .Z(n3094) );
  XNOR U3186 ( .A(n3093), .B(n3094), .Z(n3095) );
  XOR U3187 ( .A(n3096), .B(n3095), .Z(n3026) );
  NANDN U3188 ( .A(n3016), .B(n3015), .Z(n3020) );
  NANDN U3189 ( .A(n3018), .B(n3017), .Z(n3019) );
  NAND U3190 ( .A(n3020), .B(n3019), .Z(n3027) );
  XNOR U3191 ( .A(n3026), .B(n3027), .Z(n3028) );
  XNOR U3192 ( .A(n3029), .B(n3028), .Z(n3099) );
  XNOR U3193 ( .A(n3099), .B(sreg[285]), .Z(n3101) );
  NAND U3194 ( .A(n3021), .B(sreg[284]), .Z(n3025) );
  OR U3195 ( .A(n3023), .B(n3022), .Z(n3024) );
  AND U3196 ( .A(n3025), .B(n3024), .Z(n3100) );
  XOR U3197 ( .A(n3101), .B(n3100), .Z(c[285]) );
  NANDN U3198 ( .A(n3027), .B(n3026), .Z(n3031) );
  NAND U3199 ( .A(n3029), .B(n3028), .Z(n3030) );
  NAND U3200 ( .A(n3031), .B(n3030), .Z(n3107) );
  NANDN U3201 ( .A(n3033), .B(n3032), .Z(n3037) );
  OR U3202 ( .A(n3035), .B(n3034), .Z(n3036) );
  NAND U3203 ( .A(n3037), .B(n3036), .Z(n3174) );
  NANDN U3204 ( .A(n3039), .B(n3038), .Z(n3043) );
  OR U3205 ( .A(n3041), .B(n3040), .Z(n3042) );
  NAND U3206 ( .A(n3043), .B(n3042), .Z(n3140) );
  NAND U3207 ( .A(b[0]), .B(a[46]), .Z(n3044) );
  XNOR U3208 ( .A(b[1]), .B(n3044), .Z(n3046) );
  NAND U3209 ( .A(a[45]), .B(n98), .Z(n3045) );
  AND U3210 ( .A(n3046), .B(n3045), .Z(n3116) );
  XNOR U3211 ( .A(n20154), .B(n3224), .Z(n3125) );
  OR U3212 ( .A(n3125), .B(n20057), .Z(n3049) );
  NANDN U3213 ( .A(n3047), .B(n20098), .Z(n3048) );
  AND U3214 ( .A(n3049), .B(n3048), .Z(n3117) );
  XOR U3215 ( .A(n3116), .B(n3117), .Z(n3119) );
  NAND U3216 ( .A(a[30]), .B(b[15]), .Z(n3118) );
  XOR U3217 ( .A(n3119), .B(n3118), .Z(n3137) );
  NAND U3218 ( .A(n19722), .B(n3050), .Z(n3052) );
  XNOR U3219 ( .A(b[5]), .B(n3848), .Z(n3128) );
  NANDN U3220 ( .A(n19640), .B(n3128), .Z(n3051) );
  NAND U3221 ( .A(n3052), .B(n3051), .Z(n3162) );
  XNOR U3222 ( .A(n19714), .B(n3692), .Z(n3131) );
  NANDN U3223 ( .A(n3131), .B(n19766), .Z(n3055) );
  NANDN U3224 ( .A(n3053), .B(n19767), .Z(n3054) );
  NAND U3225 ( .A(n3055), .B(n3054), .Z(n3159) );
  NAND U3226 ( .A(n19554), .B(n3056), .Z(n3058) );
  IV U3227 ( .A(a[44]), .Z(n3977) );
  XNOR U3228 ( .A(b[3]), .B(n3977), .Z(n3134) );
  NANDN U3229 ( .A(n19521), .B(n3134), .Z(n3057) );
  AND U3230 ( .A(n3058), .B(n3057), .Z(n3160) );
  XNOR U3231 ( .A(n3159), .B(n3160), .Z(n3161) );
  XOR U3232 ( .A(n3162), .B(n3161), .Z(n3138) );
  XOR U3233 ( .A(n3137), .B(n3138), .Z(n3139) );
  XNOR U3234 ( .A(n3140), .B(n3139), .Z(n3110) );
  NAND U3235 ( .A(n3060), .B(n3059), .Z(n3064) );
  NAND U3236 ( .A(n3062), .B(n3061), .Z(n3063) );
  NAND U3237 ( .A(n3064), .B(n3063), .Z(n3111) );
  XOR U3238 ( .A(n3110), .B(n3111), .Z(n3113) );
  XNOR U3239 ( .A(n20052), .B(n3353), .Z(n3143) );
  OR U3240 ( .A(n3143), .B(n20020), .Z(n3067) );
  NANDN U3241 ( .A(n3065), .B(n19960), .Z(n3066) );
  NAND U3242 ( .A(n3067), .B(n3066), .Z(n3156) );
  XNOR U3243 ( .A(n102), .B(n3068), .Z(n3147) );
  OR U3244 ( .A(n3147), .B(n20121), .Z(n3071) );
  NANDN U3245 ( .A(n3069), .B(n20122), .Z(n3070) );
  NAND U3246 ( .A(n3071), .B(n3070), .Z(n3153) );
  XNOR U3247 ( .A(n19975), .B(n3536), .Z(n3150) );
  NANDN U3248 ( .A(n3150), .B(n19883), .Z(n3074) );
  NANDN U3249 ( .A(n3072), .B(n19937), .Z(n3073) );
  AND U3250 ( .A(n3074), .B(n3073), .Z(n3154) );
  XNOR U3251 ( .A(n3153), .B(n3154), .Z(n3155) );
  XNOR U3252 ( .A(n3156), .B(n3155), .Z(n3165) );
  NANDN U3253 ( .A(n3076), .B(n3075), .Z(n3080) );
  NAND U3254 ( .A(n3078), .B(n3077), .Z(n3079) );
  NAND U3255 ( .A(n3080), .B(n3079), .Z(n3166) );
  XNOR U3256 ( .A(n3165), .B(n3166), .Z(n3167) );
  NANDN U3257 ( .A(n3082), .B(n3081), .Z(n3086) );
  NAND U3258 ( .A(n3084), .B(n3083), .Z(n3085) );
  AND U3259 ( .A(n3086), .B(n3085), .Z(n3168) );
  XNOR U3260 ( .A(n3167), .B(n3168), .Z(n3112) );
  XNOR U3261 ( .A(n3113), .B(n3112), .Z(n3171) );
  NANDN U3262 ( .A(n3088), .B(n3087), .Z(n3092) );
  NAND U3263 ( .A(n3090), .B(n3089), .Z(n3091) );
  NAND U3264 ( .A(n3092), .B(n3091), .Z(n3172) );
  XNOR U3265 ( .A(n3171), .B(n3172), .Z(n3173) );
  XOR U3266 ( .A(n3174), .B(n3173), .Z(n3104) );
  NANDN U3267 ( .A(n3094), .B(n3093), .Z(n3098) );
  NANDN U3268 ( .A(n3096), .B(n3095), .Z(n3097) );
  NAND U3269 ( .A(n3098), .B(n3097), .Z(n3105) );
  XNOR U3270 ( .A(n3104), .B(n3105), .Z(n3106) );
  XNOR U3271 ( .A(n3107), .B(n3106), .Z(n3177) );
  XNOR U3272 ( .A(n3177), .B(sreg[286]), .Z(n3179) );
  NAND U3273 ( .A(n3099), .B(sreg[285]), .Z(n3103) );
  OR U3274 ( .A(n3101), .B(n3100), .Z(n3102) );
  AND U3275 ( .A(n3103), .B(n3102), .Z(n3178) );
  XOR U3276 ( .A(n3179), .B(n3178), .Z(c[286]) );
  NANDN U3277 ( .A(n3105), .B(n3104), .Z(n3109) );
  NAND U3278 ( .A(n3107), .B(n3106), .Z(n3108) );
  NAND U3279 ( .A(n3109), .B(n3108), .Z(n3185) );
  NANDN U3280 ( .A(n3111), .B(n3110), .Z(n3115) );
  OR U3281 ( .A(n3113), .B(n3112), .Z(n3114) );
  NAND U3282 ( .A(n3115), .B(n3114), .Z(n3252) );
  NANDN U3283 ( .A(n3117), .B(n3116), .Z(n3121) );
  OR U3284 ( .A(n3119), .B(n3118), .Z(n3120) );
  NAND U3285 ( .A(n3121), .B(n3120), .Z(n3218) );
  NAND U3286 ( .A(b[0]), .B(a[47]), .Z(n3122) );
  XNOR U3287 ( .A(b[1]), .B(n3122), .Z(n3124) );
  NAND U3288 ( .A(a[46]), .B(n98), .Z(n3123) );
  AND U3289 ( .A(n3124), .B(n3123), .Z(n3194) );
  XNOR U3290 ( .A(n20154), .B(n3275), .Z(n3203) );
  OR U3291 ( .A(n3203), .B(n20057), .Z(n3127) );
  NANDN U3292 ( .A(n3125), .B(n20098), .Z(n3126) );
  AND U3293 ( .A(n3127), .B(n3126), .Z(n3195) );
  XOR U3294 ( .A(n3194), .B(n3195), .Z(n3197) );
  NAND U3295 ( .A(a[31]), .B(b[15]), .Z(n3196) );
  XOR U3296 ( .A(n3197), .B(n3196), .Z(n3215) );
  NAND U3297 ( .A(n19722), .B(n3128), .Z(n3130) );
  XNOR U3298 ( .A(b[5]), .B(n3926), .Z(n3206) );
  NANDN U3299 ( .A(n19640), .B(n3206), .Z(n3129) );
  NAND U3300 ( .A(n3130), .B(n3129), .Z(n3240) );
  XNOR U3301 ( .A(n19714), .B(n3743), .Z(n3209) );
  NANDN U3302 ( .A(n3209), .B(n19766), .Z(n3133) );
  NANDN U3303 ( .A(n3131), .B(n19767), .Z(n3132) );
  NAND U3304 ( .A(n3133), .B(n3132), .Z(n3237) );
  NAND U3305 ( .A(n19554), .B(n3134), .Z(n3136) );
  IV U3306 ( .A(a[45]), .Z(n4055) );
  XNOR U3307 ( .A(b[3]), .B(n4055), .Z(n3212) );
  NANDN U3308 ( .A(n19521), .B(n3212), .Z(n3135) );
  AND U3309 ( .A(n3136), .B(n3135), .Z(n3238) );
  XNOR U3310 ( .A(n3237), .B(n3238), .Z(n3239) );
  XOR U3311 ( .A(n3240), .B(n3239), .Z(n3216) );
  XOR U3312 ( .A(n3215), .B(n3216), .Z(n3217) );
  XNOR U3313 ( .A(n3218), .B(n3217), .Z(n3188) );
  NAND U3314 ( .A(n3138), .B(n3137), .Z(n3142) );
  NAND U3315 ( .A(n3140), .B(n3139), .Z(n3141) );
  NAND U3316 ( .A(n3142), .B(n3141), .Z(n3189) );
  XOR U3317 ( .A(n3188), .B(n3189), .Z(n3191) );
  XNOR U3318 ( .A(n20052), .B(n3458), .Z(n3221) );
  OR U3319 ( .A(n3221), .B(n20020), .Z(n3145) );
  NANDN U3320 ( .A(n3143), .B(n19960), .Z(n3144) );
  NAND U3321 ( .A(n3145), .B(n3144), .Z(n3234) );
  XNOR U3322 ( .A(n102), .B(n3146), .Z(n3225) );
  OR U3323 ( .A(n3225), .B(n20121), .Z(n3149) );
  NANDN U3324 ( .A(n3147), .B(n20122), .Z(n3148) );
  NAND U3325 ( .A(n3149), .B(n3148), .Z(n3231) );
  XNOR U3326 ( .A(n19975), .B(n3587), .Z(n3228) );
  NANDN U3327 ( .A(n3228), .B(n19883), .Z(n3152) );
  NANDN U3328 ( .A(n3150), .B(n19937), .Z(n3151) );
  AND U3329 ( .A(n3152), .B(n3151), .Z(n3232) );
  XNOR U3330 ( .A(n3231), .B(n3232), .Z(n3233) );
  XNOR U3331 ( .A(n3234), .B(n3233), .Z(n3243) );
  NANDN U3332 ( .A(n3154), .B(n3153), .Z(n3158) );
  NAND U3333 ( .A(n3156), .B(n3155), .Z(n3157) );
  NAND U3334 ( .A(n3158), .B(n3157), .Z(n3244) );
  XNOR U3335 ( .A(n3243), .B(n3244), .Z(n3245) );
  NANDN U3336 ( .A(n3160), .B(n3159), .Z(n3164) );
  NAND U3337 ( .A(n3162), .B(n3161), .Z(n3163) );
  AND U3338 ( .A(n3164), .B(n3163), .Z(n3246) );
  XNOR U3339 ( .A(n3245), .B(n3246), .Z(n3190) );
  XNOR U3340 ( .A(n3191), .B(n3190), .Z(n3249) );
  NANDN U3341 ( .A(n3166), .B(n3165), .Z(n3170) );
  NAND U3342 ( .A(n3168), .B(n3167), .Z(n3169) );
  NAND U3343 ( .A(n3170), .B(n3169), .Z(n3250) );
  XNOR U3344 ( .A(n3249), .B(n3250), .Z(n3251) );
  XOR U3345 ( .A(n3252), .B(n3251), .Z(n3182) );
  NANDN U3346 ( .A(n3172), .B(n3171), .Z(n3176) );
  NANDN U3347 ( .A(n3174), .B(n3173), .Z(n3175) );
  NAND U3348 ( .A(n3176), .B(n3175), .Z(n3183) );
  XNOR U3349 ( .A(n3182), .B(n3183), .Z(n3184) );
  XNOR U3350 ( .A(n3185), .B(n3184), .Z(n3255) );
  XNOR U3351 ( .A(n3255), .B(sreg[287]), .Z(n3257) );
  NAND U3352 ( .A(n3177), .B(sreg[286]), .Z(n3181) );
  OR U3353 ( .A(n3179), .B(n3178), .Z(n3180) );
  AND U3354 ( .A(n3181), .B(n3180), .Z(n3256) );
  XOR U3355 ( .A(n3257), .B(n3256), .Z(c[287]) );
  NANDN U3356 ( .A(n3183), .B(n3182), .Z(n3187) );
  NAND U3357 ( .A(n3185), .B(n3184), .Z(n3186) );
  NAND U3358 ( .A(n3187), .B(n3186), .Z(n3263) );
  NANDN U3359 ( .A(n3189), .B(n3188), .Z(n3193) );
  OR U3360 ( .A(n3191), .B(n3190), .Z(n3192) );
  NAND U3361 ( .A(n3193), .B(n3192), .Z(n3330) );
  NANDN U3362 ( .A(n3195), .B(n3194), .Z(n3199) );
  OR U3363 ( .A(n3197), .B(n3196), .Z(n3198) );
  NAND U3364 ( .A(n3199), .B(n3198), .Z(n3318) );
  NAND U3365 ( .A(b[0]), .B(a[48]), .Z(n3200) );
  XNOR U3366 ( .A(b[1]), .B(n3200), .Z(n3202) );
  NAND U3367 ( .A(a[47]), .B(n98), .Z(n3201) );
  AND U3368 ( .A(n3202), .B(n3201), .Z(n3294) );
  XNOR U3369 ( .A(n20154), .B(n3353), .Z(n3303) );
  OR U3370 ( .A(n3303), .B(n20057), .Z(n3205) );
  NANDN U3371 ( .A(n3203), .B(n20098), .Z(n3204) );
  AND U3372 ( .A(n3205), .B(n3204), .Z(n3295) );
  XOR U3373 ( .A(n3294), .B(n3295), .Z(n3297) );
  NAND U3374 ( .A(a[32]), .B(b[15]), .Z(n3296) );
  XOR U3375 ( .A(n3297), .B(n3296), .Z(n3315) );
  NAND U3376 ( .A(n19722), .B(n3206), .Z(n3208) );
  XNOR U3377 ( .A(b[5]), .B(n3977), .Z(n3306) );
  NANDN U3378 ( .A(n19640), .B(n3306), .Z(n3207) );
  NAND U3379 ( .A(n3208), .B(n3207), .Z(n3291) );
  XNOR U3380 ( .A(n19714), .B(n3848), .Z(n3309) );
  NANDN U3381 ( .A(n3309), .B(n19766), .Z(n3211) );
  NANDN U3382 ( .A(n3209), .B(n19767), .Z(n3210) );
  NAND U3383 ( .A(n3211), .B(n3210), .Z(n3288) );
  NAND U3384 ( .A(n19554), .B(n3212), .Z(n3214) );
  IV U3385 ( .A(a[46]), .Z(n4133) );
  XNOR U3386 ( .A(b[3]), .B(n4133), .Z(n3312) );
  NANDN U3387 ( .A(n19521), .B(n3312), .Z(n3213) );
  AND U3388 ( .A(n3214), .B(n3213), .Z(n3289) );
  XNOR U3389 ( .A(n3288), .B(n3289), .Z(n3290) );
  XOR U3390 ( .A(n3291), .B(n3290), .Z(n3316) );
  XOR U3391 ( .A(n3315), .B(n3316), .Z(n3317) );
  XNOR U3392 ( .A(n3318), .B(n3317), .Z(n3266) );
  NAND U3393 ( .A(n3216), .B(n3215), .Z(n3220) );
  NAND U3394 ( .A(n3218), .B(n3217), .Z(n3219) );
  NAND U3395 ( .A(n3220), .B(n3219), .Z(n3267) );
  XOR U3396 ( .A(n3266), .B(n3267), .Z(n3269) );
  XNOR U3397 ( .A(n20052), .B(n3536), .Z(n3272) );
  OR U3398 ( .A(n3272), .B(n20020), .Z(n3223) );
  NANDN U3399 ( .A(n3221), .B(n19960), .Z(n3222) );
  NAND U3400 ( .A(n3223), .B(n3222), .Z(n3285) );
  XNOR U3401 ( .A(n102), .B(n3224), .Z(n3276) );
  OR U3402 ( .A(n3276), .B(n20121), .Z(n3227) );
  NANDN U3403 ( .A(n3225), .B(n20122), .Z(n3226) );
  NAND U3404 ( .A(n3227), .B(n3226), .Z(n3282) );
  XNOR U3405 ( .A(n19975), .B(n3692), .Z(n3279) );
  NANDN U3406 ( .A(n3279), .B(n19883), .Z(n3230) );
  NANDN U3407 ( .A(n3228), .B(n19937), .Z(n3229) );
  AND U3408 ( .A(n3230), .B(n3229), .Z(n3283) );
  XNOR U3409 ( .A(n3282), .B(n3283), .Z(n3284) );
  XNOR U3410 ( .A(n3285), .B(n3284), .Z(n3321) );
  NANDN U3411 ( .A(n3232), .B(n3231), .Z(n3236) );
  NAND U3412 ( .A(n3234), .B(n3233), .Z(n3235) );
  NAND U3413 ( .A(n3236), .B(n3235), .Z(n3322) );
  XNOR U3414 ( .A(n3321), .B(n3322), .Z(n3323) );
  NANDN U3415 ( .A(n3238), .B(n3237), .Z(n3242) );
  NAND U3416 ( .A(n3240), .B(n3239), .Z(n3241) );
  AND U3417 ( .A(n3242), .B(n3241), .Z(n3324) );
  XNOR U3418 ( .A(n3323), .B(n3324), .Z(n3268) );
  XNOR U3419 ( .A(n3269), .B(n3268), .Z(n3327) );
  NANDN U3420 ( .A(n3244), .B(n3243), .Z(n3248) );
  NAND U3421 ( .A(n3246), .B(n3245), .Z(n3247) );
  NAND U3422 ( .A(n3248), .B(n3247), .Z(n3328) );
  XNOR U3423 ( .A(n3327), .B(n3328), .Z(n3329) );
  XOR U3424 ( .A(n3330), .B(n3329), .Z(n3260) );
  NANDN U3425 ( .A(n3250), .B(n3249), .Z(n3254) );
  NANDN U3426 ( .A(n3252), .B(n3251), .Z(n3253) );
  NAND U3427 ( .A(n3254), .B(n3253), .Z(n3261) );
  XNOR U3428 ( .A(n3260), .B(n3261), .Z(n3262) );
  XNOR U3429 ( .A(n3263), .B(n3262), .Z(n3333) );
  XNOR U3430 ( .A(n3333), .B(sreg[288]), .Z(n3335) );
  NAND U3431 ( .A(n3255), .B(sreg[287]), .Z(n3259) );
  OR U3432 ( .A(n3257), .B(n3256), .Z(n3258) );
  AND U3433 ( .A(n3259), .B(n3258), .Z(n3334) );
  XOR U3434 ( .A(n3335), .B(n3334), .Z(c[288]) );
  NANDN U3435 ( .A(n3261), .B(n3260), .Z(n3265) );
  NAND U3436 ( .A(n3263), .B(n3262), .Z(n3264) );
  NAND U3437 ( .A(n3265), .B(n3264), .Z(n3341) );
  NANDN U3438 ( .A(n3267), .B(n3266), .Z(n3271) );
  OR U3439 ( .A(n3269), .B(n3268), .Z(n3270) );
  NAND U3440 ( .A(n3271), .B(n3270), .Z(n3408) );
  XNOR U3441 ( .A(n20052), .B(n3587), .Z(n3350) );
  OR U3442 ( .A(n3350), .B(n20020), .Z(n3274) );
  NANDN U3443 ( .A(n3272), .B(n19960), .Z(n3273) );
  NAND U3444 ( .A(n3274), .B(n3273), .Z(n3363) );
  XNOR U3445 ( .A(n102), .B(n3275), .Z(n3354) );
  OR U3446 ( .A(n3354), .B(n20121), .Z(n3278) );
  NANDN U3447 ( .A(n3276), .B(n20122), .Z(n3277) );
  NAND U3448 ( .A(n3278), .B(n3277), .Z(n3360) );
  XNOR U3449 ( .A(n19975), .B(n3743), .Z(n3357) );
  NANDN U3450 ( .A(n3357), .B(n19883), .Z(n3281) );
  NANDN U3451 ( .A(n3279), .B(n19937), .Z(n3280) );
  AND U3452 ( .A(n3281), .B(n3280), .Z(n3361) );
  XNOR U3453 ( .A(n3360), .B(n3361), .Z(n3362) );
  XNOR U3454 ( .A(n3363), .B(n3362), .Z(n3399) );
  NANDN U3455 ( .A(n3283), .B(n3282), .Z(n3287) );
  NAND U3456 ( .A(n3285), .B(n3284), .Z(n3286) );
  NAND U3457 ( .A(n3287), .B(n3286), .Z(n3400) );
  XNOR U3458 ( .A(n3399), .B(n3400), .Z(n3401) );
  NANDN U3459 ( .A(n3289), .B(n3288), .Z(n3293) );
  NAND U3460 ( .A(n3291), .B(n3290), .Z(n3292) );
  AND U3461 ( .A(n3293), .B(n3292), .Z(n3402) );
  XNOR U3462 ( .A(n3401), .B(n3402), .Z(n3346) );
  NANDN U3463 ( .A(n3295), .B(n3294), .Z(n3299) );
  OR U3464 ( .A(n3297), .B(n3296), .Z(n3298) );
  NAND U3465 ( .A(n3299), .B(n3298), .Z(n3396) );
  NAND U3466 ( .A(b[0]), .B(a[49]), .Z(n3300) );
  XNOR U3467 ( .A(b[1]), .B(n3300), .Z(n3302) );
  NAND U3468 ( .A(a[48]), .B(n98), .Z(n3301) );
  AND U3469 ( .A(n3302), .B(n3301), .Z(n3372) );
  XNOR U3470 ( .A(n20154), .B(n3458), .Z(n3378) );
  OR U3471 ( .A(n3378), .B(n20057), .Z(n3305) );
  NANDN U3472 ( .A(n3303), .B(n20098), .Z(n3304) );
  AND U3473 ( .A(n3305), .B(n3304), .Z(n3373) );
  XOR U3474 ( .A(n3372), .B(n3373), .Z(n3375) );
  NAND U3475 ( .A(a[33]), .B(b[15]), .Z(n3374) );
  XOR U3476 ( .A(n3375), .B(n3374), .Z(n3393) );
  NAND U3477 ( .A(n19722), .B(n3306), .Z(n3308) );
  XNOR U3478 ( .A(b[5]), .B(n4055), .Z(n3384) );
  NANDN U3479 ( .A(n19640), .B(n3384), .Z(n3307) );
  NAND U3480 ( .A(n3308), .B(n3307), .Z(n3369) );
  XNOR U3481 ( .A(n19714), .B(n3926), .Z(n3387) );
  NANDN U3482 ( .A(n3387), .B(n19766), .Z(n3311) );
  NANDN U3483 ( .A(n3309), .B(n19767), .Z(n3310) );
  NAND U3484 ( .A(n3311), .B(n3310), .Z(n3366) );
  NAND U3485 ( .A(n19554), .B(n3312), .Z(n3314) );
  IV U3486 ( .A(a[47]), .Z(n4211) );
  XNOR U3487 ( .A(b[3]), .B(n4211), .Z(n3390) );
  NANDN U3488 ( .A(n19521), .B(n3390), .Z(n3313) );
  AND U3489 ( .A(n3314), .B(n3313), .Z(n3367) );
  XNOR U3490 ( .A(n3366), .B(n3367), .Z(n3368) );
  XOR U3491 ( .A(n3369), .B(n3368), .Z(n3394) );
  XOR U3492 ( .A(n3393), .B(n3394), .Z(n3395) );
  XNOR U3493 ( .A(n3396), .B(n3395), .Z(n3344) );
  NAND U3494 ( .A(n3316), .B(n3315), .Z(n3320) );
  NAND U3495 ( .A(n3318), .B(n3317), .Z(n3319) );
  NAND U3496 ( .A(n3320), .B(n3319), .Z(n3345) );
  XOR U3497 ( .A(n3344), .B(n3345), .Z(n3347) );
  XNOR U3498 ( .A(n3346), .B(n3347), .Z(n3405) );
  NANDN U3499 ( .A(n3322), .B(n3321), .Z(n3326) );
  NAND U3500 ( .A(n3324), .B(n3323), .Z(n3325) );
  NAND U3501 ( .A(n3326), .B(n3325), .Z(n3406) );
  XNOR U3502 ( .A(n3405), .B(n3406), .Z(n3407) );
  XOR U3503 ( .A(n3408), .B(n3407), .Z(n3338) );
  NANDN U3504 ( .A(n3328), .B(n3327), .Z(n3332) );
  NANDN U3505 ( .A(n3330), .B(n3329), .Z(n3331) );
  NAND U3506 ( .A(n3332), .B(n3331), .Z(n3339) );
  XNOR U3507 ( .A(n3338), .B(n3339), .Z(n3340) );
  XNOR U3508 ( .A(n3341), .B(n3340), .Z(n3411) );
  XNOR U3509 ( .A(n3411), .B(sreg[289]), .Z(n3413) );
  NAND U3510 ( .A(n3333), .B(sreg[288]), .Z(n3337) );
  OR U3511 ( .A(n3335), .B(n3334), .Z(n3336) );
  AND U3512 ( .A(n3337), .B(n3336), .Z(n3412) );
  XOR U3513 ( .A(n3413), .B(n3412), .Z(c[289]) );
  NANDN U3514 ( .A(n3339), .B(n3338), .Z(n3343) );
  NAND U3515 ( .A(n3341), .B(n3340), .Z(n3342) );
  NAND U3516 ( .A(n3343), .B(n3342), .Z(n3419) );
  NANDN U3517 ( .A(n3345), .B(n3344), .Z(n3349) );
  OR U3518 ( .A(n3347), .B(n3346), .Z(n3348) );
  NAND U3519 ( .A(n3349), .B(n3348), .Z(n3486) );
  XNOR U3520 ( .A(n20052), .B(n3692), .Z(n3455) );
  OR U3521 ( .A(n3455), .B(n20020), .Z(n3352) );
  NANDN U3522 ( .A(n3350), .B(n19960), .Z(n3351) );
  NAND U3523 ( .A(n3352), .B(n3351), .Z(n3468) );
  XNOR U3524 ( .A(n102), .B(n3353), .Z(n3459) );
  OR U3525 ( .A(n3459), .B(n20121), .Z(n3356) );
  NANDN U3526 ( .A(n3354), .B(n20122), .Z(n3355) );
  NAND U3527 ( .A(n3356), .B(n3355), .Z(n3465) );
  XNOR U3528 ( .A(n19975), .B(n3848), .Z(n3462) );
  NANDN U3529 ( .A(n3462), .B(n19883), .Z(n3359) );
  NANDN U3530 ( .A(n3357), .B(n19937), .Z(n3358) );
  AND U3531 ( .A(n3359), .B(n3358), .Z(n3466) );
  XNOR U3532 ( .A(n3465), .B(n3466), .Z(n3467) );
  XNOR U3533 ( .A(n3468), .B(n3467), .Z(n3477) );
  NANDN U3534 ( .A(n3361), .B(n3360), .Z(n3365) );
  NAND U3535 ( .A(n3363), .B(n3362), .Z(n3364) );
  NAND U3536 ( .A(n3365), .B(n3364), .Z(n3478) );
  XNOR U3537 ( .A(n3477), .B(n3478), .Z(n3479) );
  NANDN U3538 ( .A(n3367), .B(n3366), .Z(n3371) );
  NAND U3539 ( .A(n3369), .B(n3368), .Z(n3370) );
  AND U3540 ( .A(n3371), .B(n3370), .Z(n3480) );
  XNOR U3541 ( .A(n3479), .B(n3480), .Z(n3424) );
  NANDN U3542 ( .A(n3373), .B(n3372), .Z(n3377) );
  OR U3543 ( .A(n3375), .B(n3374), .Z(n3376) );
  NAND U3544 ( .A(n3377), .B(n3376), .Z(n3452) );
  XNOR U3545 ( .A(n20154), .B(n3536), .Z(n3434) );
  OR U3546 ( .A(n3434), .B(n20057), .Z(n3380) );
  NANDN U3547 ( .A(n3378), .B(n20098), .Z(n3379) );
  AND U3548 ( .A(n3380), .B(n3379), .Z(n3429) );
  NAND U3549 ( .A(b[0]), .B(a[50]), .Z(n3381) );
  XNOR U3550 ( .A(b[1]), .B(n3381), .Z(n3383) );
  NAND U3551 ( .A(a[49]), .B(n98), .Z(n3382) );
  AND U3552 ( .A(n3383), .B(n3382), .Z(n3428) );
  XOR U3553 ( .A(n3429), .B(n3428), .Z(n3431) );
  NAND U3554 ( .A(a[34]), .B(b[15]), .Z(n3430) );
  XOR U3555 ( .A(n3431), .B(n3430), .Z(n3449) );
  NAND U3556 ( .A(n19722), .B(n3384), .Z(n3386) );
  XNOR U3557 ( .A(b[5]), .B(n4133), .Z(n3440) );
  NANDN U3558 ( .A(n19640), .B(n3440), .Z(n3385) );
  NAND U3559 ( .A(n3386), .B(n3385), .Z(n3474) );
  XNOR U3560 ( .A(n19714), .B(n3977), .Z(n3443) );
  NANDN U3561 ( .A(n3443), .B(n19766), .Z(n3389) );
  NANDN U3562 ( .A(n3387), .B(n19767), .Z(n3388) );
  NAND U3563 ( .A(n3389), .B(n3388), .Z(n3471) );
  NAND U3564 ( .A(n19554), .B(n3390), .Z(n3392) );
  IV U3565 ( .A(a[48]), .Z(n4289) );
  XNOR U3566 ( .A(b[3]), .B(n4289), .Z(n3446) );
  NANDN U3567 ( .A(n19521), .B(n3446), .Z(n3391) );
  AND U3568 ( .A(n3392), .B(n3391), .Z(n3472) );
  XNOR U3569 ( .A(n3471), .B(n3472), .Z(n3473) );
  XOR U3570 ( .A(n3474), .B(n3473), .Z(n3450) );
  XOR U3571 ( .A(n3449), .B(n3450), .Z(n3451) );
  XNOR U3572 ( .A(n3452), .B(n3451), .Z(n3422) );
  NAND U3573 ( .A(n3394), .B(n3393), .Z(n3398) );
  NAND U3574 ( .A(n3396), .B(n3395), .Z(n3397) );
  NAND U3575 ( .A(n3398), .B(n3397), .Z(n3423) );
  XOR U3576 ( .A(n3422), .B(n3423), .Z(n3425) );
  XNOR U3577 ( .A(n3424), .B(n3425), .Z(n3483) );
  NANDN U3578 ( .A(n3400), .B(n3399), .Z(n3404) );
  NAND U3579 ( .A(n3402), .B(n3401), .Z(n3403) );
  NAND U3580 ( .A(n3404), .B(n3403), .Z(n3484) );
  XNOR U3581 ( .A(n3483), .B(n3484), .Z(n3485) );
  XOR U3582 ( .A(n3486), .B(n3485), .Z(n3416) );
  NANDN U3583 ( .A(n3406), .B(n3405), .Z(n3410) );
  NANDN U3584 ( .A(n3408), .B(n3407), .Z(n3409) );
  NAND U3585 ( .A(n3410), .B(n3409), .Z(n3417) );
  XNOR U3586 ( .A(n3416), .B(n3417), .Z(n3418) );
  XNOR U3587 ( .A(n3419), .B(n3418), .Z(n3489) );
  XNOR U3588 ( .A(n3489), .B(sreg[290]), .Z(n3491) );
  NAND U3589 ( .A(n3411), .B(sreg[289]), .Z(n3415) );
  OR U3590 ( .A(n3413), .B(n3412), .Z(n3414) );
  AND U3591 ( .A(n3415), .B(n3414), .Z(n3490) );
  XOR U3592 ( .A(n3491), .B(n3490), .Z(c[290]) );
  NANDN U3593 ( .A(n3417), .B(n3416), .Z(n3421) );
  NAND U3594 ( .A(n3419), .B(n3418), .Z(n3420) );
  NAND U3595 ( .A(n3421), .B(n3420), .Z(n3497) );
  NANDN U3596 ( .A(n3423), .B(n3422), .Z(n3427) );
  OR U3597 ( .A(n3425), .B(n3424), .Z(n3426) );
  NAND U3598 ( .A(n3427), .B(n3426), .Z(n3564) );
  NANDN U3599 ( .A(n3429), .B(n3428), .Z(n3433) );
  OR U3600 ( .A(n3431), .B(n3430), .Z(n3432) );
  NAND U3601 ( .A(n3433), .B(n3432), .Z(n3530) );
  XNOR U3602 ( .A(n20154), .B(n3587), .Z(n3515) );
  OR U3603 ( .A(n3515), .B(n20057), .Z(n3436) );
  NANDN U3604 ( .A(n3434), .B(n20098), .Z(n3435) );
  AND U3605 ( .A(n3436), .B(n3435), .Z(n3507) );
  NAND U3606 ( .A(b[0]), .B(a[51]), .Z(n3437) );
  XNOR U3607 ( .A(b[1]), .B(n3437), .Z(n3439) );
  NAND U3608 ( .A(a[50]), .B(n98), .Z(n3438) );
  AND U3609 ( .A(n3439), .B(n3438), .Z(n3506) );
  XOR U3610 ( .A(n3507), .B(n3506), .Z(n3509) );
  NAND U3611 ( .A(a[35]), .B(b[15]), .Z(n3508) );
  XOR U3612 ( .A(n3509), .B(n3508), .Z(n3527) );
  NAND U3613 ( .A(n19722), .B(n3440), .Z(n3442) );
  XNOR U3614 ( .A(b[5]), .B(n4211), .Z(n3518) );
  NANDN U3615 ( .A(n19640), .B(n3518), .Z(n3441) );
  NAND U3616 ( .A(n3442), .B(n3441), .Z(n3552) );
  XNOR U3617 ( .A(n19714), .B(n4055), .Z(n3521) );
  NANDN U3618 ( .A(n3521), .B(n19766), .Z(n3445) );
  NANDN U3619 ( .A(n3443), .B(n19767), .Z(n3444) );
  NAND U3620 ( .A(n3445), .B(n3444), .Z(n3549) );
  NAND U3621 ( .A(n19554), .B(n3446), .Z(n3448) );
  IV U3622 ( .A(a[49]), .Z(n4367) );
  XNOR U3623 ( .A(b[3]), .B(n4367), .Z(n3524) );
  NANDN U3624 ( .A(n19521), .B(n3524), .Z(n3447) );
  AND U3625 ( .A(n3448), .B(n3447), .Z(n3550) );
  XNOR U3626 ( .A(n3549), .B(n3550), .Z(n3551) );
  XOR U3627 ( .A(n3552), .B(n3551), .Z(n3528) );
  XOR U3628 ( .A(n3527), .B(n3528), .Z(n3529) );
  XNOR U3629 ( .A(n3530), .B(n3529), .Z(n3500) );
  NAND U3630 ( .A(n3450), .B(n3449), .Z(n3454) );
  NAND U3631 ( .A(n3452), .B(n3451), .Z(n3453) );
  NAND U3632 ( .A(n3454), .B(n3453), .Z(n3501) );
  XOR U3633 ( .A(n3500), .B(n3501), .Z(n3503) );
  XNOR U3634 ( .A(n20052), .B(n3743), .Z(n3533) );
  OR U3635 ( .A(n3533), .B(n20020), .Z(n3457) );
  NANDN U3636 ( .A(n3455), .B(n19960), .Z(n3456) );
  NAND U3637 ( .A(n3457), .B(n3456), .Z(n3546) );
  XNOR U3638 ( .A(n102), .B(n3458), .Z(n3537) );
  OR U3639 ( .A(n3537), .B(n20121), .Z(n3461) );
  NANDN U3640 ( .A(n3459), .B(n20122), .Z(n3460) );
  NAND U3641 ( .A(n3461), .B(n3460), .Z(n3543) );
  XNOR U3642 ( .A(n19975), .B(n3926), .Z(n3540) );
  NANDN U3643 ( .A(n3540), .B(n19883), .Z(n3464) );
  NANDN U3644 ( .A(n3462), .B(n19937), .Z(n3463) );
  AND U3645 ( .A(n3464), .B(n3463), .Z(n3544) );
  XNOR U3646 ( .A(n3543), .B(n3544), .Z(n3545) );
  XNOR U3647 ( .A(n3546), .B(n3545), .Z(n3555) );
  NANDN U3648 ( .A(n3466), .B(n3465), .Z(n3470) );
  NAND U3649 ( .A(n3468), .B(n3467), .Z(n3469) );
  NAND U3650 ( .A(n3470), .B(n3469), .Z(n3556) );
  XNOR U3651 ( .A(n3555), .B(n3556), .Z(n3557) );
  NANDN U3652 ( .A(n3472), .B(n3471), .Z(n3476) );
  NAND U3653 ( .A(n3474), .B(n3473), .Z(n3475) );
  AND U3654 ( .A(n3476), .B(n3475), .Z(n3558) );
  XNOR U3655 ( .A(n3557), .B(n3558), .Z(n3502) );
  XNOR U3656 ( .A(n3503), .B(n3502), .Z(n3561) );
  NANDN U3657 ( .A(n3478), .B(n3477), .Z(n3482) );
  NAND U3658 ( .A(n3480), .B(n3479), .Z(n3481) );
  NAND U3659 ( .A(n3482), .B(n3481), .Z(n3562) );
  XNOR U3660 ( .A(n3561), .B(n3562), .Z(n3563) );
  XOR U3661 ( .A(n3564), .B(n3563), .Z(n3494) );
  NANDN U3662 ( .A(n3484), .B(n3483), .Z(n3488) );
  NANDN U3663 ( .A(n3486), .B(n3485), .Z(n3487) );
  NAND U3664 ( .A(n3488), .B(n3487), .Z(n3495) );
  XNOR U3665 ( .A(n3494), .B(n3495), .Z(n3496) );
  XNOR U3666 ( .A(n3497), .B(n3496), .Z(n3567) );
  XNOR U3667 ( .A(n3567), .B(sreg[291]), .Z(n3569) );
  NAND U3668 ( .A(n3489), .B(sreg[290]), .Z(n3493) );
  OR U3669 ( .A(n3491), .B(n3490), .Z(n3492) );
  AND U3670 ( .A(n3493), .B(n3492), .Z(n3568) );
  XOR U3671 ( .A(n3569), .B(n3568), .Z(c[291]) );
  NANDN U3672 ( .A(n3495), .B(n3494), .Z(n3499) );
  NAND U3673 ( .A(n3497), .B(n3496), .Z(n3498) );
  NAND U3674 ( .A(n3499), .B(n3498), .Z(n3575) );
  NANDN U3675 ( .A(n3501), .B(n3500), .Z(n3505) );
  OR U3676 ( .A(n3503), .B(n3502), .Z(n3504) );
  NAND U3677 ( .A(n3505), .B(n3504), .Z(n3642) );
  NANDN U3678 ( .A(n3507), .B(n3506), .Z(n3511) );
  OR U3679 ( .A(n3509), .B(n3508), .Z(n3510) );
  NAND U3680 ( .A(n3511), .B(n3510), .Z(n3630) );
  NAND U3681 ( .A(b[0]), .B(a[52]), .Z(n3512) );
  XNOR U3682 ( .A(b[1]), .B(n3512), .Z(n3514) );
  NAND U3683 ( .A(a[51]), .B(n98), .Z(n3513) );
  AND U3684 ( .A(n3514), .B(n3513), .Z(n3606) );
  XNOR U3685 ( .A(n20154), .B(n3692), .Z(n3615) );
  OR U3686 ( .A(n3615), .B(n20057), .Z(n3517) );
  NANDN U3687 ( .A(n3515), .B(n20098), .Z(n3516) );
  AND U3688 ( .A(n3517), .B(n3516), .Z(n3607) );
  XOR U3689 ( .A(n3606), .B(n3607), .Z(n3609) );
  NAND U3690 ( .A(a[36]), .B(b[15]), .Z(n3608) );
  XOR U3691 ( .A(n3609), .B(n3608), .Z(n3627) );
  NAND U3692 ( .A(n19722), .B(n3518), .Z(n3520) );
  XNOR U3693 ( .A(b[5]), .B(n4289), .Z(n3618) );
  NANDN U3694 ( .A(n19640), .B(n3618), .Z(n3519) );
  NAND U3695 ( .A(n3520), .B(n3519), .Z(n3603) );
  XNOR U3696 ( .A(n19714), .B(n4133), .Z(n3621) );
  NANDN U3697 ( .A(n3621), .B(n19766), .Z(n3523) );
  NANDN U3698 ( .A(n3521), .B(n19767), .Z(n3522) );
  NAND U3699 ( .A(n3523), .B(n3522), .Z(n3600) );
  NAND U3700 ( .A(n19554), .B(n3524), .Z(n3526) );
  IV U3701 ( .A(a[50]), .Z(n4472) );
  XNOR U3702 ( .A(b[3]), .B(n4472), .Z(n3624) );
  NANDN U3703 ( .A(n19521), .B(n3624), .Z(n3525) );
  AND U3704 ( .A(n3526), .B(n3525), .Z(n3601) );
  XNOR U3705 ( .A(n3600), .B(n3601), .Z(n3602) );
  XOR U3706 ( .A(n3603), .B(n3602), .Z(n3628) );
  XOR U3707 ( .A(n3627), .B(n3628), .Z(n3629) );
  XNOR U3708 ( .A(n3630), .B(n3629), .Z(n3578) );
  NAND U3709 ( .A(n3528), .B(n3527), .Z(n3532) );
  NAND U3710 ( .A(n3530), .B(n3529), .Z(n3531) );
  NAND U3711 ( .A(n3532), .B(n3531), .Z(n3579) );
  XOR U3712 ( .A(n3578), .B(n3579), .Z(n3581) );
  XNOR U3713 ( .A(n20052), .B(n3848), .Z(n3584) );
  OR U3714 ( .A(n3584), .B(n20020), .Z(n3535) );
  NANDN U3715 ( .A(n3533), .B(n19960), .Z(n3534) );
  NAND U3716 ( .A(n3535), .B(n3534), .Z(n3597) );
  XNOR U3717 ( .A(n102), .B(n3536), .Z(n3588) );
  OR U3718 ( .A(n3588), .B(n20121), .Z(n3539) );
  NANDN U3719 ( .A(n3537), .B(n20122), .Z(n3538) );
  NAND U3720 ( .A(n3539), .B(n3538), .Z(n3594) );
  XNOR U3721 ( .A(n19975), .B(n3977), .Z(n3591) );
  NANDN U3722 ( .A(n3591), .B(n19883), .Z(n3542) );
  NANDN U3723 ( .A(n3540), .B(n19937), .Z(n3541) );
  AND U3724 ( .A(n3542), .B(n3541), .Z(n3595) );
  XNOR U3725 ( .A(n3594), .B(n3595), .Z(n3596) );
  XNOR U3726 ( .A(n3597), .B(n3596), .Z(n3633) );
  NANDN U3727 ( .A(n3544), .B(n3543), .Z(n3548) );
  NAND U3728 ( .A(n3546), .B(n3545), .Z(n3547) );
  NAND U3729 ( .A(n3548), .B(n3547), .Z(n3634) );
  XNOR U3730 ( .A(n3633), .B(n3634), .Z(n3635) );
  NANDN U3731 ( .A(n3550), .B(n3549), .Z(n3554) );
  NAND U3732 ( .A(n3552), .B(n3551), .Z(n3553) );
  AND U3733 ( .A(n3554), .B(n3553), .Z(n3636) );
  XNOR U3734 ( .A(n3635), .B(n3636), .Z(n3580) );
  XNOR U3735 ( .A(n3581), .B(n3580), .Z(n3639) );
  NANDN U3736 ( .A(n3556), .B(n3555), .Z(n3560) );
  NAND U3737 ( .A(n3558), .B(n3557), .Z(n3559) );
  NAND U3738 ( .A(n3560), .B(n3559), .Z(n3640) );
  XNOR U3739 ( .A(n3639), .B(n3640), .Z(n3641) );
  XOR U3740 ( .A(n3642), .B(n3641), .Z(n3572) );
  NANDN U3741 ( .A(n3562), .B(n3561), .Z(n3566) );
  NANDN U3742 ( .A(n3564), .B(n3563), .Z(n3565) );
  NAND U3743 ( .A(n3566), .B(n3565), .Z(n3573) );
  XNOR U3744 ( .A(n3572), .B(n3573), .Z(n3574) );
  XNOR U3745 ( .A(n3575), .B(n3574), .Z(n3645) );
  XNOR U3746 ( .A(n3645), .B(sreg[292]), .Z(n3647) );
  NAND U3747 ( .A(n3567), .B(sreg[291]), .Z(n3571) );
  OR U3748 ( .A(n3569), .B(n3568), .Z(n3570) );
  AND U3749 ( .A(n3571), .B(n3570), .Z(n3646) );
  XOR U3750 ( .A(n3647), .B(n3646), .Z(c[292]) );
  NANDN U3751 ( .A(n3573), .B(n3572), .Z(n3577) );
  NAND U3752 ( .A(n3575), .B(n3574), .Z(n3576) );
  NAND U3753 ( .A(n3577), .B(n3576), .Z(n3653) );
  NANDN U3754 ( .A(n3579), .B(n3578), .Z(n3583) );
  OR U3755 ( .A(n3581), .B(n3580), .Z(n3582) );
  NAND U3756 ( .A(n3583), .B(n3582), .Z(n3720) );
  XNOR U3757 ( .A(n20052), .B(n3926), .Z(n3689) );
  OR U3758 ( .A(n3689), .B(n20020), .Z(n3586) );
  NANDN U3759 ( .A(n3584), .B(n19960), .Z(n3585) );
  NAND U3760 ( .A(n3586), .B(n3585), .Z(n3702) );
  XNOR U3761 ( .A(n102), .B(n3587), .Z(n3693) );
  OR U3762 ( .A(n3693), .B(n20121), .Z(n3590) );
  NANDN U3763 ( .A(n3588), .B(n20122), .Z(n3589) );
  NAND U3764 ( .A(n3590), .B(n3589), .Z(n3699) );
  XNOR U3765 ( .A(n19975), .B(n4055), .Z(n3696) );
  NANDN U3766 ( .A(n3696), .B(n19883), .Z(n3593) );
  NANDN U3767 ( .A(n3591), .B(n19937), .Z(n3592) );
  AND U3768 ( .A(n3593), .B(n3592), .Z(n3700) );
  XNOR U3769 ( .A(n3699), .B(n3700), .Z(n3701) );
  XNOR U3770 ( .A(n3702), .B(n3701), .Z(n3711) );
  NANDN U3771 ( .A(n3595), .B(n3594), .Z(n3599) );
  NAND U3772 ( .A(n3597), .B(n3596), .Z(n3598) );
  NAND U3773 ( .A(n3599), .B(n3598), .Z(n3712) );
  XNOR U3774 ( .A(n3711), .B(n3712), .Z(n3713) );
  NANDN U3775 ( .A(n3601), .B(n3600), .Z(n3605) );
  NAND U3776 ( .A(n3603), .B(n3602), .Z(n3604) );
  AND U3777 ( .A(n3605), .B(n3604), .Z(n3714) );
  XNOR U3778 ( .A(n3713), .B(n3714), .Z(n3658) );
  NANDN U3779 ( .A(n3607), .B(n3606), .Z(n3611) );
  OR U3780 ( .A(n3609), .B(n3608), .Z(n3610) );
  NAND U3781 ( .A(n3611), .B(n3610), .Z(n3686) );
  NAND U3782 ( .A(b[0]), .B(a[53]), .Z(n3612) );
  XNOR U3783 ( .A(b[1]), .B(n3612), .Z(n3614) );
  NAND U3784 ( .A(a[52]), .B(n98), .Z(n3613) );
  AND U3785 ( .A(n3614), .B(n3613), .Z(n3662) );
  XNOR U3786 ( .A(n20154), .B(n3743), .Z(n3668) );
  OR U3787 ( .A(n3668), .B(n20057), .Z(n3617) );
  NANDN U3788 ( .A(n3615), .B(n20098), .Z(n3616) );
  AND U3789 ( .A(n3617), .B(n3616), .Z(n3663) );
  XOR U3790 ( .A(n3662), .B(n3663), .Z(n3665) );
  NAND U3791 ( .A(a[37]), .B(b[15]), .Z(n3664) );
  XOR U3792 ( .A(n3665), .B(n3664), .Z(n3683) );
  NAND U3793 ( .A(n19722), .B(n3618), .Z(n3620) );
  XNOR U3794 ( .A(b[5]), .B(n4367), .Z(n3674) );
  NANDN U3795 ( .A(n19640), .B(n3674), .Z(n3619) );
  NAND U3796 ( .A(n3620), .B(n3619), .Z(n3708) );
  XNOR U3797 ( .A(n19714), .B(n4211), .Z(n3677) );
  NANDN U3798 ( .A(n3677), .B(n19766), .Z(n3623) );
  NANDN U3799 ( .A(n3621), .B(n19767), .Z(n3622) );
  NAND U3800 ( .A(n3623), .B(n3622), .Z(n3705) );
  NAND U3801 ( .A(n19554), .B(n3624), .Z(n3626) );
  IV U3802 ( .A(a[51]), .Z(n4523) );
  XNOR U3803 ( .A(b[3]), .B(n4523), .Z(n3680) );
  NANDN U3804 ( .A(n19521), .B(n3680), .Z(n3625) );
  AND U3805 ( .A(n3626), .B(n3625), .Z(n3706) );
  XNOR U3806 ( .A(n3705), .B(n3706), .Z(n3707) );
  XOR U3807 ( .A(n3708), .B(n3707), .Z(n3684) );
  XOR U3808 ( .A(n3683), .B(n3684), .Z(n3685) );
  XNOR U3809 ( .A(n3686), .B(n3685), .Z(n3656) );
  NAND U3810 ( .A(n3628), .B(n3627), .Z(n3632) );
  NAND U3811 ( .A(n3630), .B(n3629), .Z(n3631) );
  NAND U3812 ( .A(n3632), .B(n3631), .Z(n3657) );
  XOR U3813 ( .A(n3656), .B(n3657), .Z(n3659) );
  XNOR U3814 ( .A(n3658), .B(n3659), .Z(n3717) );
  NANDN U3815 ( .A(n3634), .B(n3633), .Z(n3638) );
  NAND U3816 ( .A(n3636), .B(n3635), .Z(n3637) );
  NAND U3817 ( .A(n3638), .B(n3637), .Z(n3718) );
  XNOR U3818 ( .A(n3717), .B(n3718), .Z(n3719) );
  XOR U3819 ( .A(n3720), .B(n3719), .Z(n3650) );
  NANDN U3820 ( .A(n3640), .B(n3639), .Z(n3644) );
  NANDN U3821 ( .A(n3642), .B(n3641), .Z(n3643) );
  NAND U3822 ( .A(n3644), .B(n3643), .Z(n3651) );
  XNOR U3823 ( .A(n3650), .B(n3651), .Z(n3652) );
  XNOR U3824 ( .A(n3653), .B(n3652), .Z(n3723) );
  XNOR U3825 ( .A(n3723), .B(sreg[293]), .Z(n3725) );
  NAND U3826 ( .A(n3645), .B(sreg[292]), .Z(n3649) );
  OR U3827 ( .A(n3647), .B(n3646), .Z(n3648) );
  AND U3828 ( .A(n3649), .B(n3648), .Z(n3724) );
  XOR U3829 ( .A(n3725), .B(n3724), .Z(c[293]) );
  NANDN U3830 ( .A(n3651), .B(n3650), .Z(n3655) );
  NAND U3831 ( .A(n3653), .B(n3652), .Z(n3654) );
  NAND U3832 ( .A(n3655), .B(n3654), .Z(n3731) );
  NANDN U3833 ( .A(n3657), .B(n3656), .Z(n3661) );
  OR U3834 ( .A(n3659), .B(n3658), .Z(n3660) );
  NAND U3835 ( .A(n3661), .B(n3660), .Z(n3798) );
  NANDN U3836 ( .A(n3663), .B(n3662), .Z(n3667) );
  OR U3837 ( .A(n3665), .B(n3664), .Z(n3666) );
  NAND U3838 ( .A(n3667), .B(n3666), .Z(n3786) );
  XNOR U3839 ( .A(n20154), .B(n3848), .Z(n3771) );
  OR U3840 ( .A(n3771), .B(n20057), .Z(n3670) );
  NANDN U3841 ( .A(n3668), .B(n20098), .Z(n3669) );
  AND U3842 ( .A(n3670), .B(n3669), .Z(n3763) );
  NAND U3843 ( .A(b[0]), .B(a[54]), .Z(n3671) );
  XNOR U3844 ( .A(b[1]), .B(n3671), .Z(n3673) );
  NAND U3845 ( .A(a[53]), .B(n98), .Z(n3672) );
  AND U3846 ( .A(n3673), .B(n3672), .Z(n3762) );
  XOR U3847 ( .A(n3763), .B(n3762), .Z(n3765) );
  NAND U3848 ( .A(a[38]), .B(b[15]), .Z(n3764) );
  XOR U3849 ( .A(n3765), .B(n3764), .Z(n3783) );
  NAND U3850 ( .A(n19722), .B(n3674), .Z(n3676) );
  XNOR U3851 ( .A(b[5]), .B(n4472), .Z(n3774) );
  NANDN U3852 ( .A(n19640), .B(n3774), .Z(n3675) );
  NAND U3853 ( .A(n3676), .B(n3675), .Z(n3759) );
  XNOR U3854 ( .A(n19714), .B(n4289), .Z(n3777) );
  NANDN U3855 ( .A(n3777), .B(n19766), .Z(n3679) );
  NANDN U3856 ( .A(n3677), .B(n19767), .Z(n3678) );
  NAND U3857 ( .A(n3679), .B(n3678), .Z(n3756) );
  NAND U3858 ( .A(n19554), .B(n3680), .Z(n3682) );
  IV U3859 ( .A(a[52]), .Z(n4601) );
  XNOR U3860 ( .A(b[3]), .B(n4601), .Z(n3780) );
  NANDN U3861 ( .A(n19521), .B(n3780), .Z(n3681) );
  AND U3862 ( .A(n3682), .B(n3681), .Z(n3757) );
  XNOR U3863 ( .A(n3756), .B(n3757), .Z(n3758) );
  XOR U3864 ( .A(n3759), .B(n3758), .Z(n3784) );
  XOR U3865 ( .A(n3783), .B(n3784), .Z(n3785) );
  XNOR U3866 ( .A(n3786), .B(n3785), .Z(n3734) );
  NAND U3867 ( .A(n3684), .B(n3683), .Z(n3688) );
  NAND U3868 ( .A(n3686), .B(n3685), .Z(n3687) );
  NAND U3869 ( .A(n3688), .B(n3687), .Z(n3735) );
  XOR U3870 ( .A(n3734), .B(n3735), .Z(n3737) );
  XNOR U3871 ( .A(n20052), .B(n3977), .Z(n3740) );
  OR U3872 ( .A(n3740), .B(n20020), .Z(n3691) );
  NANDN U3873 ( .A(n3689), .B(n19960), .Z(n3690) );
  NAND U3874 ( .A(n3691), .B(n3690), .Z(n3753) );
  XNOR U3875 ( .A(n102), .B(n3692), .Z(n3744) );
  OR U3876 ( .A(n3744), .B(n20121), .Z(n3695) );
  NANDN U3877 ( .A(n3693), .B(n20122), .Z(n3694) );
  NAND U3878 ( .A(n3695), .B(n3694), .Z(n3750) );
  XNOR U3879 ( .A(n19975), .B(n4133), .Z(n3747) );
  NANDN U3880 ( .A(n3747), .B(n19883), .Z(n3698) );
  NANDN U3881 ( .A(n3696), .B(n19937), .Z(n3697) );
  AND U3882 ( .A(n3698), .B(n3697), .Z(n3751) );
  XNOR U3883 ( .A(n3750), .B(n3751), .Z(n3752) );
  XNOR U3884 ( .A(n3753), .B(n3752), .Z(n3789) );
  NANDN U3885 ( .A(n3700), .B(n3699), .Z(n3704) );
  NAND U3886 ( .A(n3702), .B(n3701), .Z(n3703) );
  NAND U3887 ( .A(n3704), .B(n3703), .Z(n3790) );
  XNOR U3888 ( .A(n3789), .B(n3790), .Z(n3791) );
  NANDN U3889 ( .A(n3706), .B(n3705), .Z(n3710) );
  NAND U3890 ( .A(n3708), .B(n3707), .Z(n3709) );
  AND U3891 ( .A(n3710), .B(n3709), .Z(n3792) );
  XNOR U3892 ( .A(n3791), .B(n3792), .Z(n3736) );
  XNOR U3893 ( .A(n3737), .B(n3736), .Z(n3795) );
  NANDN U3894 ( .A(n3712), .B(n3711), .Z(n3716) );
  NAND U3895 ( .A(n3714), .B(n3713), .Z(n3715) );
  NAND U3896 ( .A(n3716), .B(n3715), .Z(n3796) );
  XNOR U3897 ( .A(n3795), .B(n3796), .Z(n3797) );
  XOR U3898 ( .A(n3798), .B(n3797), .Z(n3728) );
  NANDN U3899 ( .A(n3718), .B(n3717), .Z(n3722) );
  NANDN U3900 ( .A(n3720), .B(n3719), .Z(n3721) );
  NAND U3901 ( .A(n3722), .B(n3721), .Z(n3729) );
  XNOR U3902 ( .A(n3728), .B(n3729), .Z(n3730) );
  XNOR U3903 ( .A(n3731), .B(n3730), .Z(n3801) );
  XNOR U3904 ( .A(n3801), .B(sreg[294]), .Z(n3803) );
  NAND U3905 ( .A(n3723), .B(sreg[293]), .Z(n3727) );
  OR U3906 ( .A(n3725), .B(n3724), .Z(n3726) );
  AND U3907 ( .A(n3727), .B(n3726), .Z(n3802) );
  XOR U3908 ( .A(n3803), .B(n3802), .Z(c[294]) );
  NANDN U3909 ( .A(n3729), .B(n3728), .Z(n3733) );
  NAND U3910 ( .A(n3731), .B(n3730), .Z(n3732) );
  NAND U3911 ( .A(n3733), .B(n3732), .Z(n3809) );
  NANDN U3912 ( .A(n3735), .B(n3734), .Z(n3739) );
  OR U3913 ( .A(n3737), .B(n3736), .Z(n3738) );
  NAND U3914 ( .A(n3739), .B(n3738), .Z(n3876) );
  XNOR U3915 ( .A(n20052), .B(n4055), .Z(n3845) );
  OR U3916 ( .A(n3845), .B(n20020), .Z(n3742) );
  NANDN U3917 ( .A(n3740), .B(n19960), .Z(n3741) );
  NAND U3918 ( .A(n3742), .B(n3741), .Z(n3858) );
  XNOR U3919 ( .A(n102), .B(n3743), .Z(n3849) );
  OR U3920 ( .A(n3849), .B(n20121), .Z(n3746) );
  NANDN U3921 ( .A(n3744), .B(n20122), .Z(n3745) );
  NAND U3922 ( .A(n3746), .B(n3745), .Z(n3855) );
  XNOR U3923 ( .A(n19975), .B(n4211), .Z(n3852) );
  NANDN U3924 ( .A(n3852), .B(n19883), .Z(n3749) );
  NANDN U3925 ( .A(n3747), .B(n19937), .Z(n3748) );
  AND U3926 ( .A(n3749), .B(n3748), .Z(n3856) );
  XNOR U3927 ( .A(n3855), .B(n3856), .Z(n3857) );
  XNOR U3928 ( .A(n3858), .B(n3857), .Z(n3867) );
  NANDN U3929 ( .A(n3751), .B(n3750), .Z(n3755) );
  NAND U3930 ( .A(n3753), .B(n3752), .Z(n3754) );
  NAND U3931 ( .A(n3755), .B(n3754), .Z(n3868) );
  XNOR U3932 ( .A(n3867), .B(n3868), .Z(n3869) );
  NANDN U3933 ( .A(n3757), .B(n3756), .Z(n3761) );
  NAND U3934 ( .A(n3759), .B(n3758), .Z(n3760) );
  AND U3935 ( .A(n3761), .B(n3760), .Z(n3870) );
  XNOR U3936 ( .A(n3869), .B(n3870), .Z(n3814) );
  NANDN U3937 ( .A(n3763), .B(n3762), .Z(n3767) );
  OR U3938 ( .A(n3765), .B(n3764), .Z(n3766) );
  NAND U3939 ( .A(n3767), .B(n3766), .Z(n3842) );
  NAND U3940 ( .A(b[0]), .B(a[55]), .Z(n3768) );
  XNOR U3941 ( .A(b[1]), .B(n3768), .Z(n3770) );
  NAND U3942 ( .A(a[54]), .B(n98), .Z(n3769) );
  AND U3943 ( .A(n3770), .B(n3769), .Z(n3818) );
  XNOR U3944 ( .A(n20154), .B(n3926), .Z(n3827) );
  OR U3945 ( .A(n3827), .B(n20057), .Z(n3773) );
  NANDN U3946 ( .A(n3771), .B(n20098), .Z(n3772) );
  AND U3947 ( .A(n3773), .B(n3772), .Z(n3819) );
  XOR U3948 ( .A(n3818), .B(n3819), .Z(n3821) );
  NAND U3949 ( .A(a[39]), .B(b[15]), .Z(n3820) );
  XOR U3950 ( .A(n3821), .B(n3820), .Z(n3839) );
  NAND U3951 ( .A(n19722), .B(n3774), .Z(n3776) );
  XNOR U3952 ( .A(b[5]), .B(n4523), .Z(n3830) );
  NANDN U3953 ( .A(n19640), .B(n3830), .Z(n3775) );
  NAND U3954 ( .A(n3776), .B(n3775), .Z(n3864) );
  XNOR U3955 ( .A(n19714), .B(n4367), .Z(n3833) );
  NANDN U3956 ( .A(n3833), .B(n19766), .Z(n3779) );
  NANDN U3957 ( .A(n3777), .B(n19767), .Z(n3778) );
  NAND U3958 ( .A(n3779), .B(n3778), .Z(n3861) );
  NAND U3959 ( .A(n19554), .B(n3780), .Z(n3782) );
  IV U3960 ( .A(a[53]), .Z(n4679) );
  XNOR U3961 ( .A(b[3]), .B(n4679), .Z(n3836) );
  NANDN U3962 ( .A(n19521), .B(n3836), .Z(n3781) );
  AND U3963 ( .A(n3782), .B(n3781), .Z(n3862) );
  XNOR U3964 ( .A(n3861), .B(n3862), .Z(n3863) );
  XOR U3965 ( .A(n3864), .B(n3863), .Z(n3840) );
  XOR U3966 ( .A(n3839), .B(n3840), .Z(n3841) );
  XNOR U3967 ( .A(n3842), .B(n3841), .Z(n3812) );
  NAND U3968 ( .A(n3784), .B(n3783), .Z(n3788) );
  NAND U3969 ( .A(n3786), .B(n3785), .Z(n3787) );
  NAND U3970 ( .A(n3788), .B(n3787), .Z(n3813) );
  XOR U3971 ( .A(n3812), .B(n3813), .Z(n3815) );
  XNOR U3972 ( .A(n3814), .B(n3815), .Z(n3873) );
  NANDN U3973 ( .A(n3790), .B(n3789), .Z(n3794) );
  NAND U3974 ( .A(n3792), .B(n3791), .Z(n3793) );
  NAND U3975 ( .A(n3794), .B(n3793), .Z(n3874) );
  XNOR U3976 ( .A(n3873), .B(n3874), .Z(n3875) );
  XOR U3977 ( .A(n3876), .B(n3875), .Z(n3806) );
  NANDN U3978 ( .A(n3796), .B(n3795), .Z(n3800) );
  NANDN U3979 ( .A(n3798), .B(n3797), .Z(n3799) );
  NAND U3980 ( .A(n3800), .B(n3799), .Z(n3807) );
  XNOR U3981 ( .A(n3806), .B(n3807), .Z(n3808) );
  XNOR U3982 ( .A(n3809), .B(n3808), .Z(n3879) );
  XNOR U3983 ( .A(n3879), .B(sreg[295]), .Z(n3881) );
  NAND U3984 ( .A(n3801), .B(sreg[294]), .Z(n3805) );
  OR U3985 ( .A(n3803), .B(n3802), .Z(n3804) );
  AND U3986 ( .A(n3805), .B(n3804), .Z(n3880) );
  XOR U3987 ( .A(n3881), .B(n3880), .Z(c[295]) );
  NANDN U3988 ( .A(n3807), .B(n3806), .Z(n3811) );
  NAND U3989 ( .A(n3809), .B(n3808), .Z(n3810) );
  NAND U3990 ( .A(n3811), .B(n3810), .Z(n3887) );
  NANDN U3991 ( .A(n3813), .B(n3812), .Z(n3817) );
  OR U3992 ( .A(n3815), .B(n3814), .Z(n3816) );
  NAND U3993 ( .A(n3817), .B(n3816), .Z(n3954) );
  NANDN U3994 ( .A(n3819), .B(n3818), .Z(n3823) );
  OR U3995 ( .A(n3821), .B(n3820), .Z(n3822) );
  NAND U3996 ( .A(n3823), .B(n3822), .Z(n3920) );
  NAND U3997 ( .A(b[0]), .B(a[56]), .Z(n3824) );
  XNOR U3998 ( .A(b[1]), .B(n3824), .Z(n3826) );
  NAND U3999 ( .A(a[55]), .B(n98), .Z(n3825) );
  AND U4000 ( .A(n3826), .B(n3825), .Z(n3896) );
  XNOR U4001 ( .A(n20154), .B(n3977), .Z(n3902) );
  OR U4002 ( .A(n3902), .B(n20057), .Z(n3829) );
  NANDN U4003 ( .A(n3827), .B(n20098), .Z(n3828) );
  AND U4004 ( .A(n3829), .B(n3828), .Z(n3897) );
  XOR U4005 ( .A(n3896), .B(n3897), .Z(n3899) );
  NAND U4006 ( .A(a[40]), .B(b[15]), .Z(n3898) );
  XOR U4007 ( .A(n3899), .B(n3898), .Z(n3917) );
  NAND U4008 ( .A(n19722), .B(n3830), .Z(n3832) );
  XNOR U4009 ( .A(b[5]), .B(n4601), .Z(n3908) );
  NANDN U4010 ( .A(n19640), .B(n3908), .Z(n3831) );
  NAND U4011 ( .A(n3832), .B(n3831), .Z(n3942) );
  XNOR U4012 ( .A(n19714), .B(n4472), .Z(n3911) );
  NANDN U4013 ( .A(n3911), .B(n19766), .Z(n3835) );
  NANDN U4014 ( .A(n3833), .B(n19767), .Z(n3834) );
  NAND U4015 ( .A(n3835), .B(n3834), .Z(n3939) );
  NAND U4016 ( .A(n19554), .B(n3836), .Z(n3838) );
  IV U4017 ( .A(a[54]), .Z(n4757) );
  XNOR U4018 ( .A(b[3]), .B(n4757), .Z(n3914) );
  NANDN U4019 ( .A(n19521), .B(n3914), .Z(n3837) );
  AND U4020 ( .A(n3838), .B(n3837), .Z(n3940) );
  XNOR U4021 ( .A(n3939), .B(n3940), .Z(n3941) );
  XOR U4022 ( .A(n3942), .B(n3941), .Z(n3918) );
  XOR U4023 ( .A(n3917), .B(n3918), .Z(n3919) );
  XNOR U4024 ( .A(n3920), .B(n3919), .Z(n3890) );
  NAND U4025 ( .A(n3840), .B(n3839), .Z(n3844) );
  NAND U4026 ( .A(n3842), .B(n3841), .Z(n3843) );
  NAND U4027 ( .A(n3844), .B(n3843), .Z(n3891) );
  XOR U4028 ( .A(n3890), .B(n3891), .Z(n3893) );
  XNOR U4029 ( .A(n20052), .B(n4133), .Z(n3923) );
  OR U4030 ( .A(n3923), .B(n20020), .Z(n3847) );
  NANDN U4031 ( .A(n3845), .B(n19960), .Z(n3846) );
  NAND U4032 ( .A(n3847), .B(n3846), .Z(n3936) );
  XNOR U4033 ( .A(n102), .B(n3848), .Z(n3927) );
  OR U4034 ( .A(n3927), .B(n20121), .Z(n3851) );
  NANDN U4035 ( .A(n3849), .B(n20122), .Z(n3850) );
  NAND U4036 ( .A(n3851), .B(n3850), .Z(n3933) );
  XNOR U4037 ( .A(n19975), .B(n4289), .Z(n3930) );
  NANDN U4038 ( .A(n3930), .B(n19883), .Z(n3854) );
  NANDN U4039 ( .A(n3852), .B(n19937), .Z(n3853) );
  AND U4040 ( .A(n3854), .B(n3853), .Z(n3934) );
  XNOR U4041 ( .A(n3933), .B(n3934), .Z(n3935) );
  XNOR U4042 ( .A(n3936), .B(n3935), .Z(n3945) );
  NANDN U4043 ( .A(n3856), .B(n3855), .Z(n3860) );
  NAND U4044 ( .A(n3858), .B(n3857), .Z(n3859) );
  NAND U4045 ( .A(n3860), .B(n3859), .Z(n3946) );
  XNOR U4046 ( .A(n3945), .B(n3946), .Z(n3947) );
  NANDN U4047 ( .A(n3862), .B(n3861), .Z(n3866) );
  NAND U4048 ( .A(n3864), .B(n3863), .Z(n3865) );
  AND U4049 ( .A(n3866), .B(n3865), .Z(n3948) );
  XNOR U4050 ( .A(n3947), .B(n3948), .Z(n3892) );
  XNOR U4051 ( .A(n3893), .B(n3892), .Z(n3951) );
  NANDN U4052 ( .A(n3868), .B(n3867), .Z(n3872) );
  NAND U4053 ( .A(n3870), .B(n3869), .Z(n3871) );
  NAND U4054 ( .A(n3872), .B(n3871), .Z(n3952) );
  XNOR U4055 ( .A(n3951), .B(n3952), .Z(n3953) );
  XOR U4056 ( .A(n3954), .B(n3953), .Z(n3884) );
  NANDN U4057 ( .A(n3874), .B(n3873), .Z(n3878) );
  NANDN U4058 ( .A(n3876), .B(n3875), .Z(n3877) );
  NAND U4059 ( .A(n3878), .B(n3877), .Z(n3885) );
  XNOR U4060 ( .A(n3884), .B(n3885), .Z(n3886) );
  XNOR U4061 ( .A(n3887), .B(n3886), .Z(n3957) );
  XNOR U4062 ( .A(n3957), .B(sreg[296]), .Z(n3959) );
  NAND U4063 ( .A(n3879), .B(sreg[295]), .Z(n3883) );
  OR U4064 ( .A(n3881), .B(n3880), .Z(n3882) );
  AND U4065 ( .A(n3883), .B(n3882), .Z(n3958) );
  XOR U4066 ( .A(n3959), .B(n3958), .Z(c[296]) );
  NANDN U4067 ( .A(n3885), .B(n3884), .Z(n3889) );
  NAND U4068 ( .A(n3887), .B(n3886), .Z(n3888) );
  NAND U4069 ( .A(n3889), .B(n3888), .Z(n3965) );
  NANDN U4070 ( .A(n3891), .B(n3890), .Z(n3895) );
  OR U4071 ( .A(n3893), .B(n3892), .Z(n3894) );
  NAND U4072 ( .A(n3895), .B(n3894), .Z(n4032) );
  NANDN U4073 ( .A(n3897), .B(n3896), .Z(n3901) );
  OR U4074 ( .A(n3899), .B(n3898), .Z(n3900) );
  NAND U4075 ( .A(n3901), .B(n3900), .Z(n4020) );
  XNOR U4076 ( .A(n20154), .B(n4055), .Z(n4005) );
  OR U4077 ( .A(n4005), .B(n20057), .Z(n3904) );
  NANDN U4078 ( .A(n3902), .B(n20098), .Z(n3903) );
  AND U4079 ( .A(n3904), .B(n3903), .Z(n3997) );
  NAND U4080 ( .A(b[0]), .B(a[57]), .Z(n3905) );
  XNOR U4081 ( .A(b[1]), .B(n3905), .Z(n3907) );
  NAND U4082 ( .A(a[56]), .B(n98), .Z(n3906) );
  AND U4083 ( .A(n3907), .B(n3906), .Z(n3996) );
  XOR U4084 ( .A(n3997), .B(n3996), .Z(n3999) );
  NAND U4085 ( .A(a[41]), .B(b[15]), .Z(n3998) );
  XOR U4086 ( .A(n3999), .B(n3998), .Z(n4017) );
  NAND U4087 ( .A(n19722), .B(n3908), .Z(n3910) );
  XNOR U4088 ( .A(b[5]), .B(n4679), .Z(n4008) );
  NANDN U4089 ( .A(n19640), .B(n4008), .Z(n3909) );
  NAND U4090 ( .A(n3910), .B(n3909), .Z(n3993) );
  XNOR U4091 ( .A(n19714), .B(n4523), .Z(n4011) );
  NANDN U4092 ( .A(n4011), .B(n19766), .Z(n3913) );
  NANDN U4093 ( .A(n3911), .B(n19767), .Z(n3912) );
  NAND U4094 ( .A(n3913), .B(n3912), .Z(n3990) );
  NAND U4095 ( .A(n19554), .B(n3914), .Z(n3916) );
  IV U4096 ( .A(a[55]), .Z(n4835) );
  XNOR U4097 ( .A(b[3]), .B(n4835), .Z(n4014) );
  NANDN U4098 ( .A(n19521), .B(n4014), .Z(n3915) );
  AND U4099 ( .A(n3916), .B(n3915), .Z(n3991) );
  XNOR U4100 ( .A(n3990), .B(n3991), .Z(n3992) );
  XOR U4101 ( .A(n3993), .B(n3992), .Z(n4018) );
  XOR U4102 ( .A(n4017), .B(n4018), .Z(n4019) );
  XNOR U4103 ( .A(n4020), .B(n4019), .Z(n3968) );
  NAND U4104 ( .A(n3918), .B(n3917), .Z(n3922) );
  NAND U4105 ( .A(n3920), .B(n3919), .Z(n3921) );
  NAND U4106 ( .A(n3922), .B(n3921), .Z(n3969) );
  XOR U4107 ( .A(n3968), .B(n3969), .Z(n3971) );
  XNOR U4108 ( .A(n20052), .B(n4211), .Z(n3974) );
  OR U4109 ( .A(n3974), .B(n20020), .Z(n3925) );
  NANDN U4110 ( .A(n3923), .B(n19960), .Z(n3924) );
  NAND U4111 ( .A(n3925), .B(n3924), .Z(n3987) );
  XNOR U4112 ( .A(n102), .B(n3926), .Z(n3978) );
  OR U4113 ( .A(n3978), .B(n20121), .Z(n3929) );
  NANDN U4114 ( .A(n3927), .B(n20122), .Z(n3928) );
  NAND U4115 ( .A(n3929), .B(n3928), .Z(n3984) );
  XNOR U4116 ( .A(n19975), .B(n4367), .Z(n3981) );
  NANDN U4117 ( .A(n3981), .B(n19883), .Z(n3932) );
  NANDN U4118 ( .A(n3930), .B(n19937), .Z(n3931) );
  AND U4119 ( .A(n3932), .B(n3931), .Z(n3985) );
  XNOR U4120 ( .A(n3984), .B(n3985), .Z(n3986) );
  XNOR U4121 ( .A(n3987), .B(n3986), .Z(n4023) );
  NANDN U4122 ( .A(n3934), .B(n3933), .Z(n3938) );
  NAND U4123 ( .A(n3936), .B(n3935), .Z(n3937) );
  NAND U4124 ( .A(n3938), .B(n3937), .Z(n4024) );
  XNOR U4125 ( .A(n4023), .B(n4024), .Z(n4025) );
  NANDN U4126 ( .A(n3940), .B(n3939), .Z(n3944) );
  NAND U4127 ( .A(n3942), .B(n3941), .Z(n3943) );
  AND U4128 ( .A(n3944), .B(n3943), .Z(n4026) );
  XNOR U4129 ( .A(n4025), .B(n4026), .Z(n3970) );
  XNOR U4130 ( .A(n3971), .B(n3970), .Z(n4029) );
  NANDN U4131 ( .A(n3946), .B(n3945), .Z(n3950) );
  NAND U4132 ( .A(n3948), .B(n3947), .Z(n3949) );
  NAND U4133 ( .A(n3950), .B(n3949), .Z(n4030) );
  XNOR U4134 ( .A(n4029), .B(n4030), .Z(n4031) );
  XOR U4135 ( .A(n4032), .B(n4031), .Z(n3962) );
  NANDN U4136 ( .A(n3952), .B(n3951), .Z(n3956) );
  NANDN U4137 ( .A(n3954), .B(n3953), .Z(n3955) );
  NAND U4138 ( .A(n3956), .B(n3955), .Z(n3963) );
  XNOR U4139 ( .A(n3962), .B(n3963), .Z(n3964) );
  XNOR U4140 ( .A(n3965), .B(n3964), .Z(n4035) );
  XNOR U4141 ( .A(n4035), .B(sreg[297]), .Z(n4037) );
  NAND U4142 ( .A(n3957), .B(sreg[296]), .Z(n3961) );
  OR U4143 ( .A(n3959), .B(n3958), .Z(n3960) );
  AND U4144 ( .A(n3961), .B(n3960), .Z(n4036) );
  XOR U4145 ( .A(n4037), .B(n4036), .Z(c[297]) );
  NANDN U4146 ( .A(n3963), .B(n3962), .Z(n3967) );
  NAND U4147 ( .A(n3965), .B(n3964), .Z(n3966) );
  NAND U4148 ( .A(n3967), .B(n3966), .Z(n4043) );
  NANDN U4149 ( .A(n3969), .B(n3968), .Z(n3973) );
  OR U4150 ( .A(n3971), .B(n3970), .Z(n3972) );
  NAND U4151 ( .A(n3973), .B(n3972), .Z(n4110) );
  XNOR U4152 ( .A(n20052), .B(n4289), .Z(n4052) );
  OR U4153 ( .A(n4052), .B(n20020), .Z(n3976) );
  NANDN U4154 ( .A(n3974), .B(n19960), .Z(n3975) );
  NAND U4155 ( .A(n3976), .B(n3975), .Z(n4065) );
  XNOR U4156 ( .A(n102), .B(n3977), .Z(n4056) );
  OR U4157 ( .A(n4056), .B(n20121), .Z(n3980) );
  NANDN U4158 ( .A(n3978), .B(n20122), .Z(n3979) );
  NAND U4159 ( .A(n3980), .B(n3979), .Z(n4062) );
  XNOR U4160 ( .A(n19975), .B(n4472), .Z(n4059) );
  NANDN U4161 ( .A(n4059), .B(n19883), .Z(n3983) );
  NANDN U4162 ( .A(n3981), .B(n19937), .Z(n3982) );
  AND U4163 ( .A(n3983), .B(n3982), .Z(n4063) );
  XNOR U4164 ( .A(n4062), .B(n4063), .Z(n4064) );
  XNOR U4165 ( .A(n4065), .B(n4064), .Z(n4101) );
  NANDN U4166 ( .A(n3985), .B(n3984), .Z(n3989) );
  NAND U4167 ( .A(n3987), .B(n3986), .Z(n3988) );
  NAND U4168 ( .A(n3989), .B(n3988), .Z(n4102) );
  XNOR U4169 ( .A(n4101), .B(n4102), .Z(n4103) );
  NANDN U4170 ( .A(n3991), .B(n3990), .Z(n3995) );
  NAND U4171 ( .A(n3993), .B(n3992), .Z(n3994) );
  AND U4172 ( .A(n3995), .B(n3994), .Z(n4104) );
  XNOR U4173 ( .A(n4103), .B(n4104), .Z(n4048) );
  NANDN U4174 ( .A(n3997), .B(n3996), .Z(n4001) );
  OR U4175 ( .A(n3999), .B(n3998), .Z(n4000) );
  NAND U4176 ( .A(n4001), .B(n4000), .Z(n4098) );
  NAND U4177 ( .A(b[0]), .B(a[58]), .Z(n4002) );
  XNOR U4178 ( .A(b[1]), .B(n4002), .Z(n4004) );
  NAND U4179 ( .A(a[57]), .B(n98), .Z(n4003) );
  AND U4180 ( .A(n4004), .B(n4003), .Z(n4074) );
  XNOR U4181 ( .A(n20154), .B(n4133), .Z(n4083) );
  OR U4182 ( .A(n4083), .B(n20057), .Z(n4007) );
  NANDN U4183 ( .A(n4005), .B(n20098), .Z(n4006) );
  AND U4184 ( .A(n4007), .B(n4006), .Z(n4075) );
  XOR U4185 ( .A(n4074), .B(n4075), .Z(n4077) );
  NAND U4186 ( .A(a[42]), .B(b[15]), .Z(n4076) );
  XOR U4187 ( .A(n4077), .B(n4076), .Z(n4095) );
  NAND U4188 ( .A(n19722), .B(n4008), .Z(n4010) );
  XNOR U4189 ( .A(b[5]), .B(n4757), .Z(n4086) );
  NANDN U4190 ( .A(n19640), .B(n4086), .Z(n4009) );
  NAND U4191 ( .A(n4010), .B(n4009), .Z(n4071) );
  XNOR U4192 ( .A(n19714), .B(n4601), .Z(n4089) );
  NANDN U4193 ( .A(n4089), .B(n19766), .Z(n4013) );
  NANDN U4194 ( .A(n4011), .B(n19767), .Z(n4012) );
  NAND U4195 ( .A(n4013), .B(n4012), .Z(n4068) );
  NAND U4196 ( .A(n19554), .B(n4014), .Z(n4016) );
  IV U4197 ( .A(a[56]), .Z(n4913) );
  XNOR U4198 ( .A(b[3]), .B(n4913), .Z(n4092) );
  NANDN U4199 ( .A(n19521), .B(n4092), .Z(n4015) );
  AND U4200 ( .A(n4016), .B(n4015), .Z(n4069) );
  XNOR U4201 ( .A(n4068), .B(n4069), .Z(n4070) );
  XOR U4202 ( .A(n4071), .B(n4070), .Z(n4096) );
  XOR U4203 ( .A(n4095), .B(n4096), .Z(n4097) );
  XNOR U4204 ( .A(n4098), .B(n4097), .Z(n4046) );
  NAND U4205 ( .A(n4018), .B(n4017), .Z(n4022) );
  NAND U4206 ( .A(n4020), .B(n4019), .Z(n4021) );
  NAND U4207 ( .A(n4022), .B(n4021), .Z(n4047) );
  XOR U4208 ( .A(n4046), .B(n4047), .Z(n4049) );
  XNOR U4209 ( .A(n4048), .B(n4049), .Z(n4107) );
  NANDN U4210 ( .A(n4024), .B(n4023), .Z(n4028) );
  NAND U4211 ( .A(n4026), .B(n4025), .Z(n4027) );
  NAND U4212 ( .A(n4028), .B(n4027), .Z(n4108) );
  XNOR U4213 ( .A(n4107), .B(n4108), .Z(n4109) );
  XOR U4214 ( .A(n4110), .B(n4109), .Z(n4040) );
  NANDN U4215 ( .A(n4030), .B(n4029), .Z(n4034) );
  NANDN U4216 ( .A(n4032), .B(n4031), .Z(n4033) );
  NAND U4217 ( .A(n4034), .B(n4033), .Z(n4041) );
  XNOR U4218 ( .A(n4040), .B(n4041), .Z(n4042) );
  XNOR U4219 ( .A(n4043), .B(n4042), .Z(n4113) );
  XNOR U4220 ( .A(n4113), .B(sreg[298]), .Z(n4115) );
  NAND U4221 ( .A(n4035), .B(sreg[297]), .Z(n4039) );
  OR U4222 ( .A(n4037), .B(n4036), .Z(n4038) );
  AND U4223 ( .A(n4039), .B(n4038), .Z(n4114) );
  XOR U4224 ( .A(n4115), .B(n4114), .Z(c[298]) );
  NANDN U4225 ( .A(n4041), .B(n4040), .Z(n4045) );
  NAND U4226 ( .A(n4043), .B(n4042), .Z(n4044) );
  NAND U4227 ( .A(n4045), .B(n4044), .Z(n4121) );
  NANDN U4228 ( .A(n4047), .B(n4046), .Z(n4051) );
  OR U4229 ( .A(n4049), .B(n4048), .Z(n4050) );
  NAND U4230 ( .A(n4051), .B(n4050), .Z(n4188) );
  XNOR U4231 ( .A(n20052), .B(n4367), .Z(n4130) );
  OR U4232 ( .A(n4130), .B(n20020), .Z(n4054) );
  NANDN U4233 ( .A(n4052), .B(n19960), .Z(n4053) );
  NAND U4234 ( .A(n4054), .B(n4053), .Z(n4143) );
  XNOR U4235 ( .A(n102), .B(n4055), .Z(n4134) );
  OR U4236 ( .A(n4134), .B(n20121), .Z(n4058) );
  NANDN U4237 ( .A(n4056), .B(n20122), .Z(n4057) );
  NAND U4238 ( .A(n4058), .B(n4057), .Z(n4140) );
  XNOR U4239 ( .A(n19975), .B(n4523), .Z(n4137) );
  NANDN U4240 ( .A(n4137), .B(n19883), .Z(n4061) );
  NANDN U4241 ( .A(n4059), .B(n19937), .Z(n4060) );
  AND U4242 ( .A(n4061), .B(n4060), .Z(n4141) );
  XNOR U4243 ( .A(n4140), .B(n4141), .Z(n4142) );
  XNOR U4244 ( .A(n4143), .B(n4142), .Z(n4179) );
  NANDN U4245 ( .A(n4063), .B(n4062), .Z(n4067) );
  NAND U4246 ( .A(n4065), .B(n4064), .Z(n4066) );
  NAND U4247 ( .A(n4067), .B(n4066), .Z(n4180) );
  XNOR U4248 ( .A(n4179), .B(n4180), .Z(n4181) );
  NANDN U4249 ( .A(n4069), .B(n4068), .Z(n4073) );
  NAND U4250 ( .A(n4071), .B(n4070), .Z(n4072) );
  AND U4251 ( .A(n4073), .B(n4072), .Z(n4182) );
  XNOR U4252 ( .A(n4181), .B(n4182), .Z(n4126) );
  NANDN U4253 ( .A(n4075), .B(n4074), .Z(n4079) );
  OR U4254 ( .A(n4077), .B(n4076), .Z(n4078) );
  NAND U4255 ( .A(n4079), .B(n4078), .Z(n4176) );
  NAND U4256 ( .A(b[0]), .B(a[59]), .Z(n4080) );
  XNOR U4257 ( .A(b[1]), .B(n4080), .Z(n4082) );
  NAND U4258 ( .A(a[58]), .B(n98), .Z(n4081) );
  AND U4259 ( .A(n4082), .B(n4081), .Z(n4152) );
  XNOR U4260 ( .A(n20154), .B(n4211), .Z(n4161) );
  OR U4261 ( .A(n4161), .B(n20057), .Z(n4085) );
  NANDN U4262 ( .A(n4083), .B(n20098), .Z(n4084) );
  AND U4263 ( .A(n4085), .B(n4084), .Z(n4153) );
  XOR U4264 ( .A(n4152), .B(n4153), .Z(n4155) );
  NAND U4265 ( .A(a[43]), .B(b[15]), .Z(n4154) );
  XOR U4266 ( .A(n4155), .B(n4154), .Z(n4173) );
  NAND U4267 ( .A(n19722), .B(n4086), .Z(n4088) );
  XNOR U4268 ( .A(b[5]), .B(n4835), .Z(n4164) );
  NANDN U4269 ( .A(n19640), .B(n4164), .Z(n4087) );
  NAND U4270 ( .A(n4088), .B(n4087), .Z(n4149) );
  XNOR U4271 ( .A(n19714), .B(n4679), .Z(n4167) );
  NANDN U4272 ( .A(n4167), .B(n19766), .Z(n4091) );
  NANDN U4273 ( .A(n4089), .B(n19767), .Z(n4090) );
  NAND U4274 ( .A(n4091), .B(n4090), .Z(n4146) );
  NAND U4275 ( .A(n19554), .B(n4092), .Z(n4094) );
  IV U4276 ( .A(a[57]), .Z(n4991) );
  XNOR U4277 ( .A(b[3]), .B(n4991), .Z(n4170) );
  NANDN U4278 ( .A(n19521), .B(n4170), .Z(n4093) );
  AND U4279 ( .A(n4094), .B(n4093), .Z(n4147) );
  XNOR U4280 ( .A(n4146), .B(n4147), .Z(n4148) );
  XOR U4281 ( .A(n4149), .B(n4148), .Z(n4174) );
  XOR U4282 ( .A(n4173), .B(n4174), .Z(n4175) );
  XNOR U4283 ( .A(n4176), .B(n4175), .Z(n4124) );
  NAND U4284 ( .A(n4096), .B(n4095), .Z(n4100) );
  NAND U4285 ( .A(n4098), .B(n4097), .Z(n4099) );
  NAND U4286 ( .A(n4100), .B(n4099), .Z(n4125) );
  XOR U4287 ( .A(n4124), .B(n4125), .Z(n4127) );
  XNOR U4288 ( .A(n4126), .B(n4127), .Z(n4185) );
  NANDN U4289 ( .A(n4102), .B(n4101), .Z(n4106) );
  NAND U4290 ( .A(n4104), .B(n4103), .Z(n4105) );
  NAND U4291 ( .A(n4106), .B(n4105), .Z(n4186) );
  XNOR U4292 ( .A(n4185), .B(n4186), .Z(n4187) );
  XOR U4293 ( .A(n4188), .B(n4187), .Z(n4118) );
  NANDN U4294 ( .A(n4108), .B(n4107), .Z(n4112) );
  NANDN U4295 ( .A(n4110), .B(n4109), .Z(n4111) );
  NAND U4296 ( .A(n4112), .B(n4111), .Z(n4119) );
  XNOR U4297 ( .A(n4118), .B(n4119), .Z(n4120) );
  XNOR U4298 ( .A(n4121), .B(n4120), .Z(n4191) );
  XNOR U4299 ( .A(n4191), .B(sreg[299]), .Z(n4193) );
  NAND U4300 ( .A(n4113), .B(sreg[298]), .Z(n4117) );
  OR U4301 ( .A(n4115), .B(n4114), .Z(n4116) );
  AND U4302 ( .A(n4117), .B(n4116), .Z(n4192) );
  XOR U4303 ( .A(n4193), .B(n4192), .Z(c[299]) );
  NANDN U4304 ( .A(n4119), .B(n4118), .Z(n4123) );
  NAND U4305 ( .A(n4121), .B(n4120), .Z(n4122) );
  NAND U4306 ( .A(n4123), .B(n4122), .Z(n4199) );
  NANDN U4307 ( .A(n4125), .B(n4124), .Z(n4129) );
  OR U4308 ( .A(n4127), .B(n4126), .Z(n4128) );
  NAND U4309 ( .A(n4129), .B(n4128), .Z(n4266) );
  XNOR U4310 ( .A(n20052), .B(n4472), .Z(n4208) );
  OR U4311 ( .A(n4208), .B(n20020), .Z(n4132) );
  NANDN U4312 ( .A(n4130), .B(n19960), .Z(n4131) );
  NAND U4313 ( .A(n4132), .B(n4131), .Z(n4221) );
  XNOR U4314 ( .A(n102), .B(n4133), .Z(n4212) );
  OR U4315 ( .A(n4212), .B(n20121), .Z(n4136) );
  NANDN U4316 ( .A(n4134), .B(n20122), .Z(n4135) );
  NAND U4317 ( .A(n4136), .B(n4135), .Z(n4218) );
  XNOR U4318 ( .A(n19975), .B(n4601), .Z(n4215) );
  NANDN U4319 ( .A(n4215), .B(n19883), .Z(n4139) );
  NANDN U4320 ( .A(n4137), .B(n19937), .Z(n4138) );
  AND U4321 ( .A(n4139), .B(n4138), .Z(n4219) );
  XNOR U4322 ( .A(n4218), .B(n4219), .Z(n4220) );
  XNOR U4323 ( .A(n4221), .B(n4220), .Z(n4257) );
  NANDN U4324 ( .A(n4141), .B(n4140), .Z(n4145) );
  NAND U4325 ( .A(n4143), .B(n4142), .Z(n4144) );
  NAND U4326 ( .A(n4145), .B(n4144), .Z(n4258) );
  XNOR U4327 ( .A(n4257), .B(n4258), .Z(n4259) );
  NANDN U4328 ( .A(n4147), .B(n4146), .Z(n4151) );
  NAND U4329 ( .A(n4149), .B(n4148), .Z(n4150) );
  AND U4330 ( .A(n4151), .B(n4150), .Z(n4260) );
  XNOR U4331 ( .A(n4259), .B(n4260), .Z(n4204) );
  NANDN U4332 ( .A(n4153), .B(n4152), .Z(n4157) );
  OR U4333 ( .A(n4155), .B(n4154), .Z(n4156) );
  NAND U4334 ( .A(n4157), .B(n4156), .Z(n4254) );
  NAND U4335 ( .A(b[0]), .B(a[60]), .Z(n4158) );
  XNOR U4336 ( .A(b[1]), .B(n4158), .Z(n4160) );
  NAND U4337 ( .A(a[59]), .B(n98), .Z(n4159) );
  AND U4338 ( .A(n4160), .B(n4159), .Z(n4230) );
  XNOR U4339 ( .A(n20154), .B(n4289), .Z(n4239) );
  OR U4340 ( .A(n4239), .B(n20057), .Z(n4163) );
  NANDN U4341 ( .A(n4161), .B(n20098), .Z(n4162) );
  AND U4342 ( .A(n4163), .B(n4162), .Z(n4231) );
  XOR U4343 ( .A(n4230), .B(n4231), .Z(n4233) );
  NAND U4344 ( .A(a[44]), .B(b[15]), .Z(n4232) );
  XOR U4345 ( .A(n4233), .B(n4232), .Z(n4251) );
  NAND U4346 ( .A(n19722), .B(n4164), .Z(n4166) );
  XNOR U4347 ( .A(b[5]), .B(n4913), .Z(n4242) );
  NANDN U4348 ( .A(n19640), .B(n4242), .Z(n4165) );
  NAND U4349 ( .A(n4166), .B(n4165), .Z(n4227) );
  XNOR U4350 ( .A(n19714), .B(n4757), .Z(n4245) );
  NANDN U4351 ( .A(n4245), .B(n19766), .Z(n4169) );
  NANDN U4352 ( .A(n4167), .B(n19767), .Z(n4168) );
  NAND U4353 ( .A(n4169), .B(n4168), .Z(n4224) );
  NAND U4354 ( .A(n19554), .B(n4170), .Z(n4172) );
  IV U4355 ( .A(a[58]), .Z(n5069) );
  XNOR U4356 ( .A(b[3]), .B(n5069), .Z(n4248) );
  NANDN U4357 ( .A(n19521), .B(n4248), .Z(n4171) );
  AND U4358 ( .A(n4172), .B(n4171), .Z(n4225) );
  XNOR U4359 ( .A(n4224), .B(n4225), .Z(n4226) );
  XOR U4360 ( .A(n4227), .B(n4226), .Z(n4252) );
  XOR U4361 ( .A(n4251), .B(n4252), .Z(n4253) );
  XNOR U4362 ( .A(n4254), .B(n4253), .Z(n4202) );
  NAND U4363 ( .A(n4174), .B(n4173), .Z(n4178) );
  NAND U4364 ( .A(n4176), .B(n4175), .Z(n4177) );
  NAND U4365 ( .A(n4178), .B(n4177), .Z(n4203) );
  XOR U4366 ( .A(n4202), .B(n4203), .Z(n4205) );
  XNOR U4367 ( .A(n4204), .B(n4205), .Z(n4263) );
  NANDN U4368 ( .A(n4180), .B(n4179), .Z(n4184) );
  NAND U4369 ( .A(n4182), .B(n4181), .Z(n4183) );
  NAND U4370 ( .A(n4184), .B(n4183), .Z(n4264) );
  XNOR U4371 ( .A(n4263), .B(n4264), .Z(n4265) );
  XOR U4372 ( .A(n4266), .B(n4265), .Z(n4196) );
  NANDN U4373 ( .A(n4186), .B(n4185), .Z(n4190) );
  NANDN U4374 ( .A(n4188), .B(n4187), .Z(n4189) );
  NAND U4375 ( .A(n4190), .B(n4189), .Z(n4197) );
  XNOR U4376 ( .A(n4196), .B(n4197), .Z(n4198) );
  XNOR U4377 ( .A(n4199), .B(n4198), .Z(n4269) );
  XNOR U4378 ( .A(n4269), .B(sreg[300]), .Z(n4271) );
  NAND U4379 ( .A(n4191), .B(sreg[299]), .Z(n4195) );
  OR U4380 ( .A(n4193), .B(n4192), .Z(n4194) );
  AND U4381 ( .A(n4195), .B(n4194), .Z(n4270) );
  XOR U4382 ( .A(n4271), .B(n4270), .Z(c[300]) );
  NANDN U4383 ( .A(n4197), .B(n4196), .Z(n4201) );
  NAND U4384 ( .A(n4199), .B(n4198), .Z(n4200) );
  NAND U4385 ( .A(n4201), .B(n4200), .Z(n4277) );
  NANDN U4386 ( .A(n4203), .B(n4202), .Z(n4207) );
  OR U4387 ( .A(n4205), .B(n4204), .Z(n4206) );
  NAND U4388 ( .A(n4207), .B(n4206), .Z(n4344) );
  XNOR U4389 ( .A(n20052), .B(n4523), .Z(n4286) );
  OR U4390 ( .A(n4286), .B(n20020), .Z(n4210) );
  NANDN U4391 ( .A(n4208), .B(n19960), .Z(n4209) );
  NAND U4392 ( .A(n4210), .B(n4209), .Z(n4299) );
  XNOR U4393 ( .A(n102), .B(n4211), .Z(n4290) );
  OR U4394 ( .A(n4290), .B(n20121), .Z(n4214) );
  NANDN U4395 ( .A(n4212), .B(n20122), .Z(n4213) );
  NAND U4396 ( .A(n4214), .B(n4213), .Z(n4296) );
  XNOR U4397 ( .A(n19975), .B(n4679), .Z(n4293) );
  NANDN U4398 ( .A(n4293), .B(n19883), .Z(n4217) );
  NANDN U4399 ( .A(n4215), .B(n19937), .Z(n4216) );
  AND U4400 ( .A(n4217), .B(n4216), .Z(n4297) );
  XNOR U4401 ( .A(n4296), .B(n4297), .Z(n4298) );
  XNOR U4402 ( .A(n4299), .B(n4298), .Z(n4335) );
  NANDN U4403 ( .A(n4219), .B(n4218), .Z(n4223) );
  NAND U4404 ( .A(n4221), .B(n4220), .Z(n4222) );
  NAND U4405 ( .A(n4223), .B(n4222), .Z(n4336) );
  XNOR U4406 ( .A(n4335), .B(n4336), .Z(n4337) );
  NANDN U4407 ( .A(n4225), .B(n4224), .Z(n4229) );
  NAND U4408 ( .A(n4227), .B(n4226), .Z(n4228) );
  AND U4409 ( .A(n4229), .B(n4228), .Z(n4338) );
  XNOR U4410 ( .A(n4337), .B(n4338), .Z(n4282) );
  NANDN U4411 ( .A(n4231), .B(n4230), .Z(n4235) );
  OR U4412 ( .A(n4233), .B(n4232), .Z(n4234) );
  NAND U4413 ( .A(n4235), .B(n4234), .Z(n4332) );
  NAND U4414 ( .A(b[0]), .B(a[61]), .Z(n4236) );
  XNOR U4415 ( .A(b[1]), .B(n4236), .Z(n4238) );
  NAND U4416 ( .A(a[60]), .B(n98), .Z(n4237) );
  AND U4417 ( .A(n4238), .B(n4237), .Z(n4308) );
  XNOR U4418 ( .A(n20154), .B(n4367), .Z(n4314) );
  OR U4419 ( .A(n4314), .B(n20057), .Z(n4241) );
  NANDN U4420 ( .A(n4239), .B(n20098), .Z(n4240) );
  AND U4421 ( .A(n4241), .B(n4240), .Z(n4309) );
  XOR U4422 ( .A(n4308), .B(n4309), .Z(n4311) );
  NAND U4423 ( .A(a[45]), .B(b[15]), .Z(n4310) );
  XOR U4424 ( .A(n4311), .B(n4310), .Z(n4329) );
  NAND U4425 ( .A(n19722), .B(n4242), .Z(n4244) );
  XNOR U4426 ( .A(b[5]), .B(n4991), .Z(n4320) );
  NANDN U4427 ( .A(n19640), .B(n4320), .Z(n4243) );
  NAND U4428 ( .A(n4244), .B(n4243), .Z(n4305) );
  XNOR U4429 ( .A(n19714), .B(n4835), .Z(n4323) );
  NANDN U4430 ( .A(n4323), .B(n19766), .Z(n4247) );
  NANDN U4431 ( .A(n4245), .B(n19767), .Z(n4246) );
  NAND U4432 ( .A(n4247), .B(n4246), .Z(n4302) );
  NAND U4433 ( .A(n19554), .B(n4248), .Z(n4250) );
  IV U4434 ( .A(a[59]), .Z(n5147) );
  XNOR U4435 ( .A(b[3]), .B(n5147), .Z(n4326) );
  NANDN U4436 ( .A(n19521), .B(n4326), .Z(n4249) );
  AND U4437 ( .A(n4250), .B(n4249), .Z(n4303) );
  XNOR U4438 ( .A(n4302), .B(n4303), .Z(n4304) );
  XOR U4439 ( .A(n4305), .B(n4304), .Z(n4330) );
  XOR U4440 ( .A(n4329), .B(n4330), .Z(n4331) );
  XNOR U4441 ( .A(n4332), .B(n4331), .Z(n4280) );
  NAND U4442 ( .A(n4252), .B(n4251), .Z(n4256) );
  NAND U4443 ( .A(n4254), .B(n4253), .Z(n4255) );
  NAND U4444 ( .A(n4256), .B(n4255), .Z(n4281) );
  XOR U4445 ( .A(n4280), .B(n4281), .Z(n4283) );
  XNOR U4446 ( .A(n4282), .B(n4283), .Z(n4341) );
  NANDN U4447 ( .A(n4258), .B(n4257), .Z(n4262) );
  NAND U4448 ( .A(n4260), .B(n4259), .Z(n4261) );
  NAND U4449 ( .A(n4262), .B(n4261), .Z(n4342) );
  XNOR U4450 ( .A(n4341), .B(n4342), .Z(n4343) );
  XOR U4451 ( .A(n4344), .B(n4343), .Z(n4274) );
  NANDN U4452 ( .A(n4264), .B(n4263), .Z(n4268) );
  NANDN U4453 ( .A(n4266), .B(n4265), .Z(n4267) );
  NAND U4454 ( .A(n4268), .B(n4267), .Z(n4275) );
  XNOR U4455 ( .A(n4274), .B(n4275), .Z(n4276) );
  XNOR U4456 ( .A(n4277), .B(n4276), .Z(n4347) );
  XNOR U4457 ( .A(n4347), .B(sreg[301]), .Z(n4349) );
  NAND U4458 ( .A(n4269), .B(sreg[300]), .Z(n4273) );
  OR U4459 ( .A(n4271), .B(n4270), .Z(n4272) );
  AND U4460 ( .A(n4273), .B(n4272), .Z(n4348) );
  XOR U4461 ( .A(n4349), .B(n4348), .Z(c[301]) );
  NANDN U4462 ( .A(n4275), .B(n4274), .Z(n4279) );
  NAND U4463 ( .A(n4277), .B(n4276), .Z(n4278) );
  NAND U4464 ( .A(n4279), .B(n4278), .Z(n4355) );
  NANDN U4465 ( .A(n4281), .B(n4280), .Z(n4285) );
  OR U4466 ( .A(n4283), .B(n4282), .Z(n4284) );
  NAND U4467 ( .A(n4285), .B(n4284), .Z(n4422) );
  XNOR U4468 ( .A(n20052), .B(n4601), .Z(n4364) );
  OR U4469 ( .A(n4364), .B(n20020), .Z(n4288) );
  NANDN U4470 ( .A(n4286), .B(n19960), .Z(n4287) );
  NAND U4471 ( .A(n4288), .B(n4287), .Z(n4377) );
  XNOR U4472 ( .A(n102), .B(n4289), .Z(n4368) );
  OR U4473 ( .A(n4368), .B(n20121), .Z(n4292) );
  NANDN U4474 ( .A(n4290), .B(n20122), .Z(n4291) );
  NAND U4475 ( .A(n4292), .B(n4291), .Z(n4374) );
  XNOR U4476 ( .A(n19975), .B(n4757), .Z(n4371) );
  NANDN U4477 ( .A(n4371), .B(n19883), .Z(n4295) );
  NANDN U4478 ( .A(n4293), .B(n19937), .Z(n4294) );
  AND U4479 ( .A(n4295), .B(n4294), .Z(n4375) );
  XNOR U4480 ( .A(n4374), .B(n4375), .Z(n4376) );
  XNOR U4481 ( .A(n4377), .B(n4376), .Z(n4413) );
  NANDN U4482 ( .A(n4297), .B(n4296), .Z(n4301) );
  NAND U4483 ( .A(n4299), .B(n4298), .Z(n4300) );
  NAND U4484 ( .A(n4301), .B(n4300), .Z(n4414) );
  XNOR U4485 ( .A(n4413), .B(n4414), .Z(n4415) );
  NANDN U4486 ( .A(n4303), .B(n4302), .Z(n4307) );
  NAND U4487 ( .A(n4305), .B(n4304), .Z(n4306) );
  AND U4488 ( .A(n4307), .B(n4306), .Z(n4416) );
  XNOR U4489 ( .A(n4415), .B(n4416), .Z(n4360) );
  NANDN U4490 ( .A(n4309), .B(n4308), .Z(n4313) );
  OR U4491 ( .A(n4311), .B(n4310), .Z(n4312) );
  NAND U4492 ( .A(n4313), .B(n4312), .Z(n4410) );
  XNOR U4493 ( .A(n20154), .B(n4472), .Z(n4392) );
  OR U4494 ( .A(n4392), .B(n20057), .Z(n4316) );
  NANDN U4495 ( .A(n4314), .B(n20098), .Z(n4315) );
  AND U4496 ( .A(n4316), .B(n4315), .Z(n4387) );
  NAND U4497 ( .A(b[0]), .B(a[62]), .Z(n4317) );
  XNOR U4498 ( .A(b[1]), .B(n4317), .Z(n4319) );
  NAND U4499 ( .A(a[61]), .B(n98), .Z(n4318) );
  AND U4500 ( .A(n4319), .B(n4318), .Z(n4386) );
  XOR U4501 ( .A(n4387), .B(n4386), .Z(n4389) );
  NAND U4502 ( .A(a[46]), .B(b[15]), .Z(n4388) );
  XOR U4503 ( .A(n4389), .B(n4388), .Z(n4407) );
  NAND U4504 ( .A(n19722), .B(n4320), .Z(n4322) );
  XNOR U4505 ( .A(b[5]), .B(n5069), .Z(n4398) );
  NANDN U4506 ( .A(n19640), .B(n4398), .Z(n4321) );
  NAND U4507 ( .A(n4322), .B(n4321), .Z(n4383) );
  XNOR U4508 ( .A(n19714), .B(n4913), .Z(n4401) );
  NANDN U4509 ( .A(n4401), .B(n19766), .Z(n4325) );
  NANDN U4510 ( .A(n4323), .B(n19767), .Z(n4324) );
  NAND U4511 ( .A(n4325), .B(n4324), .Z(n4380) );
  NAND U4512 ( .A(n19554), .B(n4326), .Z(n4328) );
  IV U4513 ( .A(a[60]), .Z(n5225) );
  XNOR U4514 ( .A(b[3]), .B(n5225), .Z(n4404) );
  NANDN U4515 ( .A(n19521), .B(n4404), .Z(n4327) );
  AND U4516 ( .A(n4328), .B(n4327), .Z(n4381) );
  XNOR U4517 ( .A(n4380), .B(n4381), .Z(n4382) );
  XOR U4518 ( .A(n4383), .B(n4382), .Z(n4408) );
  XOR U4519 ( .A(n4407), .B(n4408), .Z(n4409) );
  XNOR U4520 ( .A(n4410), .B(n4409), .Z(n4358) );
  NAND U4521 ( .A(n4330), .B(n4329), .Z(n4334) );
  NAND U4522 ( .A(n4332), .B(n4331), .Z(n4333) );
  NAND U4523 ( .A(n4334), .B(n4333), .Z(n4359) );
  XOR U4524 ( .A(n4358), .B(n4359), .Z(n4361) );
  XNOR U4525 ( .A(n4360), .B(n4361), .Z(n4419) );
  NANDN U4526 ( .A(n4336), .B(n4335), .Z(n4340) );
  NAND U4527 ( .A(n4338), .B(n4337), .Z(n4339) );
  NAND U4528 ( .A(n4340), .B(n4339), .Z(n4420) );
  XNOR U4529 ( .A(n4419), .B(n4420), .Z(n4421) );
  XOR U4530 ( .A(n4422), .B(n4421), .Z(n4352) );
  NANDN U4531 ( .A(n4342), .B(n4341), .Z(n4346) );
  NANDN U4532 ( .A(n4344), .B(n4343), .Z(n4345) );
  NAND U4533 ( .A(n4346), .B(n4345), .Z(n4353) );
  XNOR U4534 ( .A(n4352), .B(n4353), .Z(n4354) );
  XNOR U4535 ( .A(n4355), .B(n4354), .Z(n4425) );
  XNOR U4536 ( .A(n4425), .B(sreg[302]), .Z(n4427) );
  NAND U4537 ( .A(n4347), .B(sreg[301]), .Z(n4351) );
  OR U4538 ( .A(n4349), .B(n4348), .Z(n4350) );
  AND U4539 ( .A(n4351), .B(n4350), .Z(n4426) );
  XOR U4540 ( .A(n4427), .B(n4426), .Z(c[302]) );
  NANDN U4541 ( .A(n4353), .B(n4352), .Z(n4357) );
  NAND U4542 ( .A(n4355), .B(n4354), .Z(n4356) );
  NAND U4543 ( .A(n4357), .B(n4356), .Z(n4433) );
  NANDN U4544 ( .A(n4359), .B(n4358), .Z(n4363) );
  OR U4545 ( .A(n4361), .B(n4360), .Z(n4362) );
  NAND U4546 ( .A(n4363), .B(n4362), .Z(n4500) );
  XNOR U4547 ( .A(n20052), .B(n4679), .Z(n4469) );
  OR U4548 ( .A(n4469), .B(n20020), .Z(n4366) );
  NANDN U4549 ( .A(n4364), .B(n19960), .Z(n4365) );
  NAND U4550 ( .A(n4366), .B(n4365), .Z(n4482) );
  XNOR U4551 ( .A(n102), .B(n4367), .Z(n4473) );
  OR U4552 ( .A(n4473), .B(n20121), .Z(n4370) );
  NANDN U4553 ( .A(n4368), .B(n20122), .Z(n4369) );
  NAND U4554 ( .A(n4370), .B(n4369), .Z(n4479) );
  XNOR U4555 ( .A(n19975), .B(n4835), .Z(n4476) );
  NANDN U4556 ( .A(n4476), .B(n19883), .Z(n4373) );
  NANDN U4557 ( .A(n4371), .B(n19937), .Z(n4372) );
  AND U4558 ( .A(n4373), .B(n4372), .Z(n4480) );
  XNOR U4559 ( .A(n4479), .B(n4480), .Z(n4481) );
  XNOR U4560 ( .A(n4482), .B(n4481), .Z(n4491) );
  NANDN U4561 ( .A(n4375), .B(n4374), .Z(n4379) );
  NAND U4562 ( .A(n4377), .B(n4376), .Z(n4378) );
  NAND U4563 ( .A(n4379), .B(n4378), .Z(n4492) );
  XNOR U4564 ( .A(n4491), .B(n4492), .Z(n4493) );
  NANDN U4565 ( .A(n4381), .B(n4380), .Z(n4385) );
  NAND U4566 ( .A(n4383), .B(n4382), .Z(n4384) );
  AND U4567 ( .A(n4385), .B(n4384), .Z(n4494) );
  XNOR U4568 ( .A(n4493), .B(n4494), .Z(n4438) );
  NANDN U4569 ( .A(n4387), .B(n4386), .Z(n4391) );
  OR U4570 ( .A(n4389), .B(n4388), .Z(n4390) );
  NAND U4571 ( .A(n4391), .B(n4390), .Z(n4466) );
  XNOR U4572 ( .A(n20154), .B(n4523), .Z(n4451) );
  OR U4573 ( .A(n4451), .B(n20057), .Z(n4394) );
  NANDN U4574 ( .A(n4392), .B(n20098), .Z(n4393) );
  AND U4575 ( .A(n4394), .B(n4393), .Z(n4443) );
  NAND U4576 ( .A(b[0]), .B(a[63]), .Z(n4395) );
  XNOR U4577 ( .A(b[1]), .B(n4395), .Z(n4397) );
  NAND U4578 ( .A(a[62]), .B(n98), .Z(n4396) );
  AND U4579 ( .A(n4397), .B(n4396), .Z(n4442) );
  XOR U4580 ( .A(n4443), .B(n4442), .Z(n4445) );
  NAND U4581 ( .A(a[47]), .B(b[15]), .Z(n4444) );
  XOR U4582 ( .A(n4445), .B(n4444), .Z(n4463) );
  NAND U4583 ( .A(n19722), .B(n4398), .Z(n4400) );
  XNOR U4584 ( .A(b[5]), .B(n5147), .Z(n4454) );
  NANDN U4585 ( .A(n19640), .B(n4454), .Z(n4399) );
  NAND U4586 ( .A(n4400), .B(n4399), .Z(n4488) );
  XNOR U4587 ( .A(n19714), .B(n4991), .Z(n4457) );
  NANDN U4588 ( .A(n4457), .B(n19766), .Z(n4403) );
  NANDN U4589 ( .A(n4401), .B(n19767), .Z(n4402) );
  NAND U4590 ( .A(n4403), .B(n4402), .Z(n4485) );
  NAND U4591 ( .A(n19554), .B(n4404), .Z(n4406) );
  IV U4592 ( .A(a[61]), .Z(n5303) );
  XNOR U4593 ( .A(b[3]), .B(n5303), .Z(n4460) );
  NANDN U4594 ( .A(n19521), .B(n4460), .Z(n4405) );
  AND U4595 ( .A(n4406), .B(n4405), .Z(n4486) );
  XNOR U4596 ( .A(n4485), .B(n4486), .Z(n4487) );
  XOR U4597 ( .A(n4488), .B(n4487), .Z(n4464) );
  XOR U4598 ( .A(n4463), .B(n4464), .Z(n4465) );
  XNOR U4599 ( .A(n4466), .B(n4465), .Z(n4436) );
  NAND U4600 ( .A(n4408), .B(n4407), .Z(n4412) );
  NAND U4601 ( .A(n4410), .B(n4409), .Z(n4411) );
  NAND U4602 ( .A(n4412), .B(n4411), .Z(n4437) );
  XOR U4603 ( .A(n4436), .B(n4437), .Z(n4439) );
  XNOR U4604 ( .A(n4438), .B(n4439), .Z(n4497) );
  NANDN U4605 ( .A(n4414), .B(n4413), .Z(n4418) );
  NAND U4606 ( .A(n4416), .B(n4415), .Z(n4417) );
  NAND U4607 ( .A(n4418), .B(n4417), .Z(n4498) );
  XNOR U4608 ( .A(n4497), .B(n4498), .Z(n4499) );
  XOR U4609 ( .A(n4500), .B(n4499), .Z(n4430) );
  NANDN U4610 ( .A(n4420), .B(n4419), .Z(n4424) );
  NANDN U4611 ( .A(n4422), .B(n4421), .Z(n4423) );
  NAND U4612 ( .A(n4424), .B(n4423), .Z(n4431) );
  XNOR U4613 ( .A(n4430), .B(n4431), .Z(n4432) );
  XNOR U4614 ( .A(n4433), .B(n4432), .Z(n4503) );
  XNOR U4615 ( .A(n4503), .B(sreg[303]), .Z(n4505) );
  NAND U4616 ( .A(n4425), .B(sreg[302]), .Z(n4429) );
  OR U4617 ( .A(n4427), .B(n4426), .Z(n4428) );
  AND U4618 ( .A(n4429), .B(n4428), .Z(n4504) );
  XOR U4619 ( .A(n4505), .B(n4504), .Z(c[303]) );
  NANDN U4620 ( .A(n4431), .B(n4430), .Z(n4435) );
  NAND U4621 ( .A(n4433), .B(n4432), .Z(n4434) );
  NAND U4622 ( .A(n4435), .B(n4434), .Z(n4511) );
  NANDN U4623 ( .A(n4437), .B(n4436), .Z(n4441) );
  OR U4624 ( .A(n4439), .B(n4438), .Z(n4440) );
  NAND U4625 ( .A(n4441), .B(n4440), .Z(n4578) );
  NANDN U4626 ( .A(n4443), .B(n4442), .Z(n4447) );
  OR U4627 ( .A(n4445), .B(n4444), .Z(n4446) );
  NAND U4628 ( .A(n4447), .B(n4446), .Z(n4566) );
  NAND U4629 ( .A(b[0]), .B(a[64]), .Z(n4448) );
  XNOR U4630 ( .A(b[1]), .B(n4448), .Z(n4450) );
  NAND U4631 ( .A(a[63]), .B(n98), .Z(n4449) );
  AND U4632 ( .A(n4450), .B(n4449), .Z(n4542) );
  XNOR U4633 ( .A(n20154), .B(n4601), .Z(n4551) );
  OR U4634 ( .A(n4551), .B(n20057), .Z(n4453) );
  NANDN U4635 ( .A(n4451), .B(n20098), .Z(n4452) );
  AND U4636 ( .A(n4453), .B(n4452), .Z(n4543) );
  XOR U4637 ( .A(n4542), .B(n4543), .Z(n4545) );
  NAND U4638 ( .A(a[48]), .B(b[15]), .Z(n4544) );
  XOR U4639 ( .A(n4545), .B(n4544), .Z(n4563) );
  NAND U4640 ( .A(n19722), .B(n4454), .Z(n4456) );
  XNOR U4641 ( .A(b[5]), .B(n5225), .Z(n4554) );
  NANDN U4642 ( .A(n19640), .B(n4554), .Z(n4455) );
  NAND U4643 ( .A(n4456), .B(n4455), .Z(n4539) );
  XNOR U4644 ( .A(n19714), .B(n5069), .Z(n4557) );
  NANDN U4645 ( .A(n4557), .B(n19766), .Z(n4459) );
  NANDN U4646 ( .A(n4457), .B(n19767), .Z(n4458) );
  NAND U4647 ( .A(n4459), .B(n4458), .Z(n4536) );
  NAND U4648 ( .A(n19554), .B(n4460), .Z(n4462) );
  IV U4649 ( .A(a[62]), .Z(n5381) );
  XNOR U4650 ( .A(b[3]), .B(n5381), .Z(n4560) );
  NANDN U4651 ( .A(n19521), .B(n4560), .Z(n4461) );
  AND U4652 ( .A(n4462), .B(n4461), .Z(n4537) );
  XNOR U4653 ( .A(n4536), .B(n4537), .Z(n4538) );
  XOR U4654 ( .A(n4539), .B(n4538), .Z(n4564) );
  XOR U4655 ( .A(n4563), .B(n4564), .Z(n4565) );
  XNOR U4656 ( .A(n4566), .B(n4565), .Z(n4514) );
  NAND U4657 ( .A(n4464), .B(n4463), .Z(n4468) );
  NAND U4658 ( .A(n4466), .B(n4465), .Z(n4467) );
  NAND U4659 ( .A(n4468), .B(n4467), .Z(n4515) );
  XOR U4660 ( .A(n4514), .B(n4515), .Z(n4517) );
  XNOR U4661 ( .A(n20052), .B(n4757), .Z(n4520) );
  OR U4662 ( .A(n4520), .B(n20020), .Z(n4471) );
  NANDN U4663 ( .A(n4469), .B(n19960), .Z(n4470) );
  NAND U4664 ( .A(n4471), .B(n4470), .Z(n4533) );
  XNOR U4665 ( .A(n102), .B(n4472), .Z(n4524) );
  OR U4666 ( .A(n4524), .B(n20121), .Z(n4475) );
  NANDN U4667 ( .A(n4473), .B(n20122), .Z(n4474) );
  NAND U4668 ( .A(n4475), .B(n4474), .Z(n4530) );
  XNOR U4669 ( .A(n19975), .B(n4913), .Z(n4527) );
  NANDN U4670 ( .A(n4527), .B(n19883), .Z(n4478) );
  NANDN U4671 ( .A(n4476), .B(n19937), .Z(n4477) );
  AND U4672 ( .A(n4478), .B(n4477), .Z(n4531) );
  XNOR U4673 ( .A(n4530), .B(n4531), .Z(n4532) );
  XNOR U4674 ( .A(n4533), .B(n4532), .Z(n4569) );
  NANDN U4675 ( .A(n4480), .B(n4479), .Z(n4484) );
  NAND U4676 ( .A(n4482), .B(n4481), .Z(n4483) );
  NAND U4677 ( .A(n4484), .B(n4483), .Z(n4570) );
  XNOR U4678 ( .A(n4569), .B(n4570), .Z(n4571) );
  NANDN U4679 ( .A(n4486), .B(n4485), .Z(n4490) );
  NAND U4680 ( .A(n4488), .B(n4487), .Z(n4489) );
  AND U4681 ( .A(n4490), .B(n4489), .Z(n4572) );
  XNOR U4682 ( .A(n4571), .B(n4572), .Z(n4516) );
  XNOR U4683 ( .A(n4517), .B(n4516), .Z(n4575) );
  NANDN U4684 ( .A(n4492), .B(n4491), .Z(n4496) );
  NAND U4685 ( .A(n4494), .B(n4493), .Z(n4495) );
  NAND U4686 ( .A(n4496), .B(n4495), .Z(n4576) );
  XNOR U4687 ( .A(n4575), .B(n4576), .Z(n4577) );
  XOR U4688 ( .A(n4578), .B(n4577), .Z(n4508) );
  NANDN U4689 ( .A(n4498), .B(n4497), .Z(n4502) );
  NANDN U4690 ( .A(n4500), .B(n4499), .Z(n4501) );
  NAND U4691 ( .A(n4502), .B(n4501), .Z(n4509) );
  XNOR U4692 ( .A(n4508), .B(n4509), .Z(n4510) );
  XNOR U4693 ( .A(n4511), .B(n4510), .Z(n4581) );
  XNOR U4694 ( .A(n4581), .B(sreg[304]), .Z(n4583) );
  NAND U4695 ( .A(n4503), .B(sreg[303]), .Z(n4507) );
  OR U4696 ( .A(n4505), .B(n4504), .Z(n4506) );
  AND U4697 ( .A(n4507), .B(n4506), .Z(n4582) );
  XOR U4698 ( .A(n4583), .B(n4582), .Z(c[304]) );
  NANDN U4699 ( .A(n4509), .B(n4508), .Z(n4513) );
  NAND U4700 ( .A(n4511), .B(n4510), .Z(n4512) );
  NAND U4701 ( .A(n4513), .B(n4512), .Z(n4589) );
  NANDN U4702 ( .A(n4515), .B(n4514), .Z(n4519) );
  OR U4703 ( .A(n4517), .B(n4516), .Z(n4518) );
  NAND U4704 ( .A(n4519), .B(n4518), .Z(n4656) );
  XNOR U4705 ( .A(n20052), .B(n4835), .Z(n4598) );
  OR U4706 ( .A(n4598), .B(n20020), .Z(n4522) );
  NANDN U4707 ( .A(n4520), .B(n19960), .Z(n4521) );
  NAND U4708 ( .A(n4522), .B(n4521), .Z(n4611) );
  XNOR U4709 ( .A(n102), .B(n4523), .Z(n4602) );
  OR U4710 ( .A(n4602), .B(n20121), .Z(n4526) );
  NANDN U4711 ( .A(n4524), .B(n20122), .Z(n4525) );
  NAND U4712 ( .A(n4526), .B(n4525), .Z(n4608) );
  XNOR U4713 ( .A(n19975), .B(n4991), .Z(n4605) );
  NANDN U4714 ( .A(n4605), .B(n19883), .Z(n4529) );
  NANDN U4715 ( .A(n4527), .B(n19937), .Z(n4528) );
  AND U4716 ( .A(n4529), .B(n4528), .Z(n4609) );
  XNOR U4717 ( .A(n4608), .B(n4609), .Z(n4610) );
  XNOR U4718 ( .A(n4611), .B(n4610), .Z(n4647) );
  NANDN U4719 ( .A(n4531), .B(n4530), .Z(n4535) );
  NAND U4720 ( .A(n4533), .B(n4532), .Z(n4534) );
  NAND U4721 ( .A(n4535), .B(n4534), .Z(n4648) );
  XNOR U4722 ( .A(n4647), .B(n4648), .Z(n4649) );
  NANDN U4723 ( .A(n4537), .B(n4536), .Z(n4541) );
  NAND U4724 ( .A(n4539), .B(n4538), .Z(n4540) );
  AND U4725 ( .A(n4541), .B(n4540), .Z(n4650) );
  XNOR U4726 ( .A(n4649), .B(n4650), .Z(n4594) );
  NANDN U4727 ( .A(n4543), .B(n4542), .Z(n4547) );
  OR U4728 ( .A(n4545), .B(n4544), .Z(n4546) );
  NAND U4729 ( .A(n4547), .B(n4546), .Z(n4644) );
  NAND U4730 ( .A(b[0]), .B(a[65]), .Z(n4548) );
  XNOR U4731 ( .A(b[1]), .B(n4548), .Z(n4550) );
  NAND U4732 ( .A(a[64]), .B(n98), .Z(n4549) );
  AND U4733 ( .A(n4550), .B(n4549), .Z(n4620) );
  XNOR U4734 ( .A(n20154), .B(n4679), .Z(n4629) );
  OR U4735 ( .A(n4629), .B(n20057), .Z(n4553) );
  NANDN U4736 ( .A(n4551), .B(n20098), .Z(n4552) );
  AND U4737 ( .A(n4553), .B(n4552), .Z(n4621) );
  XOR U4738 ( .A(n4620), .B(n4621), .Z(n4623) );
  NAND U4739 ( .A(a[49]), .B(b[15]), .Z(n4622) );
  XOR U4740 ( .A(n4623), .B(n4622), .Z(n4641) );
  NAND U4741 ( .A(n19722), .B(n4554), .Z(n4556) );
  XNOR U4742 ( .A(b[5]), .B(n5303), .Z(n4632) );
  NANDN U4743 ( .A(n19640), .B(n4632), .Z(n4555) );
  NAND U4744 ( .A(n4556), .B(n4555), .Z(n4617) );
  XNOR U4745 ( .A(n19714), .B(n5147), .Z(n4635) );
  NANDN U4746 ( .A(n4635), .B(n19766), .Z(n4559) );
  NANDN U4747 ( .A(n4557), .B(n19767), .Z(n4558) );
  NAND U4748 ( .A(n4559), .B(n4558), .Z(n4614) );
  NAND U4749 ( .A(n19554), .B(n4560), .Z(n4562) );
  IV U4750 ( .A(a[63]), .Z(n5459) );
  XNOR U4751 ( .A(b[3]), .B(n5459), .Z(n4638) );
  NANDN U4752 ( .A(n19521), .B(n4638), .Z(n4561) );
  AND U4753 ( .A(n4562), .B(n4561), .Z(n4615) );
  XNOR U4754 ( .A(n4614), .B(n4615), .Z(n4616) );
  XOR U4755 ( .A(n4617), .B(n4616), .Z(n4642) );
  XOR U4756 ( .A(n4641), .B(n4642), .Z(n4643) );
  XNOR U4757 ( .A(n4644), .B(n4643), .Z(n4592) );
  NAND U4758 ( .A(n4564), .B(n4563), .Z(n4568) );
  NAND U4759 ( .A(n4566), .B(n4565), .Z(n4567) );
  NAND U4760 ( .A(n4568), .B(n4567), .Z(n4593) );
  XOR U4761 ( .A(n4592), .B(n4593), .Z(n4595) );
  XNOR U4762 ( .A(n4594), .B(n4595), .Z(n4653) );
  NANDN U4763 ( .A(n4570), .B(n4569), .Z(n4574) );
  NAND U4764 ( .A(n4572), .B(n4571), .Z(n4573) );
  NAND U4765 ( .A(n4574), .B(n4573), .Z(n4654) );
  XNOR U4766 ( .A(n4653), .B(n4654), .Z(n4655) );
  XOR U4767 ( .A(n4656), .B(n4655), .Z(n4586) );
  NANDN U4768 ( .A(n4576), .B(n4575), .Z(n4580) );
  NANDN U4769 ( .A(n4578), .B(n4577), .Z(n4579) );
  NAND U4770 ( .A(n4580), .B(n4579), .Z(n4587) );
  XNOR U4771 ( .A(n4586), .B(n4587), .Z(n4588) );
  XNOR U4772 ( .A(n4589), .B(n4588), .Z(n4659) );
  XNOR U4773 ( .A(n4659), .B(sreg[305]), .Z(n4661) );
  NAND U4774 ( .A(n4581), .B(sreg[304]), .Z(n4585) );
  OR U4775 ( .A(n4583), .B(n4582), .Z(n4584) );
  AND U4776 ( .A(n4585), .B(n4584), .Z(n4660) );
  XOR U4777 ( .A(n4661), .B(n4660), .Z(c[305]) );
  NANDN U4778 ( .A(n4587), .B(n4586), .Z(n4591) );
  NAND U4779 ( .A(n4589), .B(n4588), .Z(n4590) );
  NAND U4780 ( .A(n4591), .B(n4590), .Z(n4667) );
  NANDN U4781 ( .A(n4593), .B(n4592), .Z(n4597) );
  OR U4782 ( .A(n4595), .B(n4594), .Z(n4596) );
  NAND U4783 ( .A(n4597), .B(n4596), .Z(n4734) );
  XNOR U4784 ( .A(n20052), .B(n4913), .Z(n4676) );
  OR U4785 ( .A(n4676), .B(n20020), .Z(n4600) );
  NANDN U4786 ( .A(n4598), .B(n19960), .Z(n4599) );
  NAND U4787 ( .A(n4600), .B(n4599), .Z(n4689) );
  XNOR U4788 ( .A(n102), .B(n4601), .Z(n4680) );
  OR U4789 ( .A(n4680), .B(n20121), .Z(n4604) );
  NANDN U4790 ( .A(n4602), .B(n20122), .Z(n4603) );
  NAND U4791 ( .A(n4604), .B(n4603), .Z(n4686) );
  XNOR U4792 ( .A(n19975), .B(n5069), .Z(n4683) );
  NANDN U4793 ( .A(n4683), .B(n19883), .Z(n4607) );
  NANDN U4794 ( .A(n4605), .B(n19937), .Z(n4606) );
  AND U4795 ( .A(n4607), .B(n4606), .Z(n4687) );
  XNOR U4796 ( .A(n4686), .B(n4687), .Z(n4688) );
  XNOR U4797 ( .A(n4689), .B(n4688), .Z(n4725) );
  NANDN U4798 ( .A(n4609), .B(n4608), .Z(n4613) );
  NAND U4799 ( .A(n4611), .B(n4610), .Z(n4612) );
  NAND U4800 ( .A(n4613), .B(n4612), .Z(n4726) );
  XNOR U4801 ( .A(n4725), .B(n4726), .Z(n4727) );
  NANDN U4802 ( .A(n4615), .B(n4614), .Z(n4619) );
  NAND U4803 ( .A(n4617), .B(n4616), .Z(n4618) );
  AND U4804 ( .A(n4619), .B(n4618), .Z(n4728) );
  XNOR U4805 ( .A(n4727), .B(n4728), .Z(n4672) );
  NANDN U4806 ( .A(n4621), .B(n4620), .Z(n4625) );
  OR U4807 ( .A(n4623), .B(n4622), .Z(n4624) );
  NAND U4808 ( .A(n4625), .B(n4624), .Z(n4722) );
  NAND U4809 ( .A(b[0]), .B(a[66]), .Z(n4626) );
  XNOR U4810 ( .A(b[1]), .B(n4626), .Z(n4628) );
  NAND U4811 ( .A(a[65]), .B(n98), .Z(n4627) );
  AND U4812 ( .A(n4628), .B(n4627), .Z(n4698) );
  XNOR U4813 ( .A(n20154), .B(n4757), .Z(n4707) );
  OR U4814 ( .A(n4707), .B(n20057), .Z(n4631) );
  NANDN U4815 ( .A(n4629), .B(n20098), .Z(n4630) );
  AND U4816 ( .A(n4631), .B(n4630), .Z(n4699) );
  XOR U4817 ( .A(n4698), .B(n4699), .Z(n4701) );
  NAND U4818 ( .A(a[50]), .B(b[15]), .Z(n4700) );
  XOR U4819 ( .A(n4701), .B(n4700), .Z(n4719) );
  NAND U4820 ( .A(n19722), .B(n4632), .Z(n4634) );
  XNOR U4821 ( .A(b[5]), .B(n5381), .Z(n4710) );
  NANDN U4822 ( .A(n19640), .B(n4710), .Z(n4633) );
  NAND U4823 ( .A(n4634), .B(n4633), .Z(n4695) );
  XNOR U4824 ( .A(n19714), .B(n5225), .Z(n4713) );
  NANDN U4825 ( .A(n4713), .B(n19766), .Z(n4637) );
  NANDN U4826 ( .A(n4635), .B(n19767), .Z(n4636) );
  NAND U4827 ( .A(n4637), .B(n4636), .Z(n4692) );
  NAND U4828 ( .A(n19554), .B(n4638), .Z(n4640) );
  IV U4829 ( .A(a[64]), .Z(n5549) );
  XNOR U4830 ( .A(b[3]), .B(n5549), .Z(n4716) );
  NANDN U4831 ( .A(n19521), .B(n4716), .Z(n4639) );
  AND U4832 ( .A(n4640), .B(n4639), .Z(n4693) );
  XNOR U4833 ( .A(n4692), .B(n4693), .Z(n4694) );
  XOR U4834 ( .A(n4695), .B(n4694), .Z(n4720) );
  XOR U4835 ( .A(n4719), .B(n4720), .Z(n4721) );
  XNOR U4836 ( .A(n4722), .B(n4721), .Z(n4670) );
  NAND U4837 ( .A(n4642), .B(n4641), .Z(n4646) );
  NAND U4838 ( .A(n4644), .B(n4643), .Z(n4645) );
  NAND U4839 ( .A(n4646), .B(n4645), .Z(n4671) );
  XOR U4840 ( .A(n4670), .B(n4671), .Z(n4673) );
  XNOR U4841 ( .A(n4672), .B(n4673), .Z(n4731) );
  NANDN U4842 ( .A(n4648), .B(n4647), .Z(n4652) );
  NAND U4843 ( .A(n4650), .B(n4649), .Z(n4651) );
  NAND U4844 ( .A(n4652), .B(n4651), .Z(n4732) );
  XNOR U4845 ( .A(n4731), .B(n4732), .Z(n4733) );
  XOR U4846 ( .A(n4734), .B(n4733), .Z(n4664) );
  NANDN U4847 ( .A(n4654), .B(n4653), .Z(n4658) );
  NANDN U4848 ( .A(n4656), .B(n4655), .Z(n4657) );
  NAND U4849 ( .A(n4658), .B(n4657), .Z(n4665) );
  XNOR U4850 ( .A(n4664), .B(n4665), .Z(n4666) );
  XNOR U4851 ( .A(n4667), .B(n4666), .Z(n4737) );
  XNOR U4852 ( .A(n4737), .B(sreg[306]), .Z(n4739) );
  NAND U4853 ( .A(n4659), .B(sreg[305]), .Z(n4663) );
  OR U4854 ( .A(n4661), .B(n4660), .Z(n4662) );
  AND U4855 ( .A(n4663), .B(n4662), .Z(n4738) );
  XOR U4856 ( .A(n4739), .B(n4738), .Z(c[306]) );
  NANDN U4857 ( .A(n4665), .B(n4664), .Z(n4669) );
  NAND U4858 ( .A(n4667), .B(n4666), .Z(n4668) );
  NAND U4859 ( .A(n4669), .B(n4668), .Z(n4745) );
  NANDN U4860 ( .A(n4671), .B(n4670), .Z(n4675) );
  OR U4861 ( .A(n4673), .B(n4672), .Z(n4674) );
  NAND U4862 ( .A(n4675), .B(n4674), .Z(n4812) );
  XNOR U4863 ( .A(n20052), .B(n4991), .Z(n4754) );
  OR U4864 ( .A(n4754), .B(n20020), .Z(n4678) );
  NANDN U4865 ( .A(n4676), .B(n19960), .Z(n4677) );
  NAND U4866 ( .A(n4678), .B(n4677), .Z(n4767) );
  XNOR U4867 ( .A(n102), .B(n4679), .Z(n4758) );
  OR U4868 ( .A(n4758), .B(n20121), .Z(n4682) );
  NANDN U4869 ( .A(n4680), .B(n20122), .Z(n4681) );
  NAND U4870 ( .A(n4682), .B(n4681), .Z(n4764) );
  XNOR U4871 ( .A(n19975), .B(n5147), .Z(n4761) );
  NANDN U4872 ( .A(n4761), .B(n19883), .Z(n4685) );
  NANDN U4873 ( .A(n4683), .B(n19937), .Z(n4684) );
  AND U4874 ( .A(n4685), .B(n4684), .Z(n4765) );
  XNOR U4875 ( .A(n4764), .B(n4765), .Z(n4766) );
  XNOR U4876 ( .A(n4767), .B(n4766), .Z(n4803) );
  NANDN U4877 ( .A(n4687), .B(n4686), .Z(n4691) );
  NAND U4878 ( .A(n4689), .B(n4688), .Z(n4690) );
  NAND U4879 ( .A(n4691), .B(n4690), .Z(n4804) );
  XNOR U4880 ( .A(n4803), .B(n4804), .Z(n4805) );
  NANDN U4881 ( .A(n4693), .B(n4692), .Z(n4697) );
  NAND U4882 ( .A(n4695), .B(n4694), .Z(n4696) );
  AND U4883 ( .A(n4697), .B(n4696), .Z(n4806) );
  XNOR U4884 ( .A(n4805), .B(n4806), .Z(n4750) );
  NANDN U4885 ( .A(n4699), .B(n4698), .Z(n4703) );
  OR U4886 ( .A(n4701), .B(n4700), .Z(n4702) );
  NAND U4887 ( .A(n4703), .B(n4702), .Z(n4800) );
  NAND U4888 ( .A(b[0]), .B(a[67]), .Z(n4704) );
  XNOR U4889 ( .A(b[1]), .B(n4704), .Z(n4706) );
  NAND U4890 ( .A(a[66]), .B(n98), .Z(n4705) );
  AND U4891 ( .A(n4706), .B(n4705), .Z(n4776) );
  XNOR U4892 ( .A(n20154), .B(n4835), .Z(n4782) );
  OR U4893 ( .A(n4782), .B(n20057), .Z(n4709) );
  NANDN U4894 ( .A(n4707), .B(n20098), .Z(n4708) );
  AND U4895 ( .A(n4709), .B(n4708), .Z(n4777) );
  XOR U4896 ( .A(n4776), .B(n4777), .Z(n4779) );
  NAND U4897 ( .A(a[51]), .B(b[15]), .Z(n4778) );
  XOR U4898 ( .A(n4779), .B(n4778), .Z(n4797) );
  NAND U4899 ( .A(n19722), .B(n4710), .Z(n4712) );
  XNOR U4900 ( .A(b[5]), .B(n5459), .Z(n4788) );
  NANDN U4901 ( .A(n19640), .B(n4788), .Z(n4711) );
  NAND U4902 ( .A(n4712), .B(n4711), .Z(n4773) );
  XNOR U4903 ( .A(n19714), .B(n5303), .Z(n4791) );
  NANDN U4904 ( .A(n4791), .B(n19766), .Z(n4715) );
  NANDN U4905 ( .A(n4713), .B(n19767), .Z(n4714) );
  NAND U4906 ( .A(n4715), .B(n4714), .Z(n4770) );
  NAND U4907 ( .A(n19554), .B(n4716), .Z(n4718) );
  IV U4908 ( .A(a[65]), .Z(n5615) );
  XNOR U4909 ( .A(b[3]), .B(n5615), .Z(n4794) );
  NANDN U4910 ( .A(n19521), .B(n4794), .Z(n4717) );
  AND U4911 ( .A(n4718), .B(n4717), .Z(n4771) );
  XNOR U4912 ( .A(n4770), .B(n4771), .Z(n4772) );
  XOR U4913 ( .A(n4773), .B(n4772), .Z(n4798) );
  XOR U4914 ( .A(n4797), .B(n4798), .Z(n4799) );
  XNOR U4915 ( .A(n4800), .B(n4799), .Z(n4748) );
  NAND U4916 ( .A(n4720), .B(n4719), .Z(n4724) );
  NAND U4917 ( .A(n4722), .B(n4721), .Z(n4723) );
  NAND U4918 ( .A(n4724), .B(n4723), .Z(n4749) );
  XOR U4919 ( .A(n4748), .B(n4749), .Z(n4751) );
  XNOR U4920 ( .A(n4750), .B(n4751), .Z(n4809) );
  NANDN U4921 ( .A(n4726), .B(n4725), .Z(n4730) );
  NAND U4922 ( .A(n4728), .B(n4727), .Z(n4729) );
  NAND U4923 ( .A(n4730), .B(n4729), .Z(n4810) );
  XNOR U4924 ( .A(n4809), .B(n4810), .Z(n4811) );
  XOR U4925 ( .A(n4812), .B(n4811), .Z(n4742) );
  NANDN U4926 ( .A(n4732), .B(n4731), .Z(n4736) );
  NANDN U4927 ( .A(n4734), .B(n4733), .Z(n4735) );
  NAND U4928 ( .A(n4736), .B(n4735), .Z(n4743) );
  XNOR U4929 ( .A(n4742), .B(n4743), .Z(n4744) );
  XNOR U4930 ( .A(n4745), .B(n4744), .Z(n4815) );
  XNOR U4931 ( .A(n4815), .B(sreg[307]), .Z(n4817) );
  NAND U4932 ( .A(n4737), .B(sreg[306]), .Z(n4741) );
  OR U4933 ( .A(n4739), .B(n4738), .Z(n4740) );
  AND U4934 ( .A(n4741), .B(n4740), .Z(n4816) );
  XOR U4935 ( .A(n4817), .B(n4816), .Z(c[307]) );
  NANDN U4936 ( .A(n4743), .B(n4742), .Z(n4747) );
  NAND U4937 ( .A(n4745), .B(n4744), .Z(n4746) );
  NAND U4938 ( .A(n4747), .B(n4746), .Z(n4823) );
  NANDN U4939 ( .A(n4749), .B(n4748), .Z(n4753) );
  OR U4940 ( .A(n4751), .B(n4750), .Z(n4752) );
  NAND U4941 ( .A(n4753), .B(n4752), .Z(n4890) );
  XNOR U4942 ( .A(n20052), .B(n5069), .Z(n4832) );
  OR U4943 ( .A(n4832), .B(n20020), .Z(n4756) );
  NANDN U4944 ( .A(n4754), .B(n19960), .Z(n4755) );
  NAND U4945 ( .A(n4756), .B(n4755), .Z(n4845) );
  XNOR U4946 ( .A(n102), .B(n4757), .Z(n4836) );
  OR U4947 ( .A(n4836), .B(n20121), .Z(n4760) );
  NANDN U4948 ( .A(n4758), .B(n20122), .Z(n4759) );
  NAND U4949 ( .A(n4760), .B(n4759), .Z(n4842) );
  XNOR U4950 ( .A(n19975), .B(n5225), .Z(n4839) );
  NANDN U4951 ( .A(n4839), .B(n19883), .Z(n4763) );
  NANDN U4952 ( .A(n4761), .B(n19937), .Z(n4762) );
  AND U4953 ( .A(n4763), .B(n4762), .Z(n4843) );
  XNOR U4954 ( .A(n4842), .B(n4843), .Z(n4844) );
  XNOR U4955 ( .A(n4845), .B(n4844), .Z(n4881) );
  NANDN U4956 ( .A(n4765), .B(n4764), .Z(n4769) );
  NAND U4957 ( .A(n4767), .B(n4766), .Z(n4768) );
  NAND U4958 ( .A(n4769), .B(n4768), .Z(n4882) );
  XNOR U4959 ( .A(n4881), .B(n4882), .Z(n4883) );
  NANDN U4960 ( .A(n4771), .B(n4770), .Z(n4775) );
  NAND U4961 ( .A(n4773), .B(n4772), .Z(n4774) );
  AND U4962 ( .A(n4775), .B(n4774), .Z(n4884) );
  XNOR U4963 ( .A(n4883), .B(n4884), .Z(n4828) );
  NANDN U4964 ( .A(n4777), .B(n4776), .Z(n4781) );
  OR U4965 ( .A(n4779), .B(n4778), .Z(n4780) );
  NAND U4966 ( .A(n4781), .B(n4780), .Z(n4878) );
  XNOR U4967 ( .A(n20154), .B(n4913), .Z(n4863) );
  OR U4968 ( .A(n4863), .B(n20057), .Z(n4784) );
  NANDN U4969 ( .A(n4782), .B(n20098), .Z(n4783) );
  AND U4970 ( .A(n4784), .B(n4783), .Z(n4855) );
  NAND U4971 ( .A(b[0]), .B(a[68]), .Z(n4785) );
  XNOR U4972 ( .A(b[1]), .B(n4785), .Z(n4787) );
  NAND U4973 ( .A(a[67]), .B(n98), .Z(n4786) );
  AND U4974 ( .A(n4787), .B(n4786), .Z(n4854) );
  XOR U4975 ( .A(n4855), .B(n4854), .Z(n4857) );
  NAND U4976 ( .A(a[52]), .B(b[15]), .Z(n4856) );
  XOR U4977 ( .A(n4857), .B(n4856), .Z(n4875) );
  NAND U4978 ( .A(n19722), .B(n4788), .Z(n4790) );
  XNOR U4979 ( .A(b[5]), .B(n5549), .Z(n4866) );
  NANDN U4980 ( .A(n19640), .B(n4866), .Z(n4789) );
  NAND U4981 ( .A(n4790), .B(n4789), .Z(n4851) );
  XNOR U4982 ( .A(n19714), .B(n5381), .Z(n4869) );
  NANDN U4983 ( .A(n4869), .B(n19766), .Z(n4793) );
  NANDN U4984 ( .A(n4791), .B(n19767), .Z(n4792) );
  NAND U4985 ( .A(n4793), .B(n4792), .Z(n4848) );
  NAND U4986 ( .A(n19554), .B(n4794), .Z(n4796) );
  IV U4987 ( .A(a[66]), .Z(n5693) );
  XNOR U4988 ( .A(b[3]), .B(n5693), .Z(n4872) );
  NANDN U4989 ( .A(n19521), .B(n4872), .Z(n4795) );
  AND U4990 ( .A(n4796), .B(n4795), .Z(n4849) );
  XNOR U4991 ( .A(n4848), .B(n4849), .Z(n4850) );
  XOR U4992 ( .A(n4851), .B(n4850), .Z(n4876) );
  XOR U4993 ( .A(n4875), .B(n4876), .Z(n4877) );
  XNOR U4994 ( .A(n4878), .B(n4877), .Z(n4826) );
  NAND U4995 ( .A(n4798), .B(n4797), .Z(n4802) );
  NAND U4996 ( .A(n4800), .B(n4799), .Z(n4801) );
  NAND U4997 ( .A(n4802), .B(n4801), .Z(n4827) );
  XOR U4998 ( .A(n4826), .B(n4827), .Z(n4829) );
  XNOR U4999 ( .A(n4828), .B(n4829), .Z(n4887) );
  NANDN U5000 ( .A(n4804), .B(n4803), .Z(n4808) );
  NAND U5001 ( .A(n4806), .B(n4805), .Z(n4807) );
  NAND U5002 ( .A(n4808), .B(n4807), .Z(n4888) );
  XNOR U5003 ( .A(n4887), .B(n4888), .Z(n4889) );
  XOR U5004 ( .A(n4890), .B(n4889), .Z(n4820) );
  NANDN U5005 ( .A(n4810), .B(n4809), .Z(n4814) );
  NANDN U5006 ( .A(n4812), .B(n4811), .Z(n4813) );
  NAND U5007 ( .A(n4814), .B(n4813), .Z(n4821) );
  XNOR U5008 ( .A(n4820), .B(n4821), .Z(n4822) );
  XNOR U5009 ( .A(n4823), .B(n4822), .Z(n4893) );
  XNOR U5010 ( .A(n4893), .B(sreg[308]), .Z(n4895) );
  NAND U5011 ( .A(n4815), .B(sreg[307]), .Z(n4819) );
  OR U5012 ( .A(n4817), .B(n4816), .Z(n4818) );
  AND U5013 ( .A(n4819), .B(n4818), .Z(n4894) );
  XOR U5014 ( .A(n4895), .B(n4894), .Z(c[308]) );
  NANDN U5015 ( .A(n4821), .B(n4820), .Z(n4825) );
  NAND U5016 ( .A(n4823), .B(n4822), .Z(n4824) );
  NAND U5017 ( .A(n4825), .B(n4824), .Z(n4901) );
  NANDN U5018 ( .A(n4827), .B(n4826), .Z(n4831) );
  OR U5019 ( .A(n4829), .B(n4828), .Z(n4830) );
  NAND U5020 ( .A(n4831), .B(n4830), .Z(n4968) );
  XNOR U5021 ( .A(n20052), .B(n5147), .Z(n4910) );
  OR U5022 ( .A(n4910), .B(n20020), .Z(n4834) );
  NANDN U5023 ( .A(n4832), .B(n19960), .Z(n4833) );
  NAND U5024 ( .A(n4834), .B(n4833), .Z(n4923) );
  XNOR U5025 ( .A(n102), .B(n4835), .Z(n4914) );
  OR U5026 ( .A(n4914), .B(n20121), .Z(n4838) );
  NANDN U5027 ( .A(n4836), .B(n20122), .Z(n4837) );
  NAND U5028 ( .A(n4838), .B(n4837), .Z(n4920) );
  XNOR U5029 ( .A(n19975), .B(n5303), .Z(n4917) );
  NANDN U5030 ( .A(n4917), .B(n19883), .Z(n4841) );
  NANDN U5031 ( .A(n4839), .B(n19937), .Z(n4840) );
  AND U5032 ( .A(n4841), .B(n4840), .Z(n4921) );
  XNOR U5033 ( .A(n4920), .B(n4921), .Z(n4922) );
  XNOR U5034 ( .A(n4923), .B(n4922), .Z(n4959) );
  NANDN U5035 ( .A(n4843), .B(n4842), .Z(n4847) );
  NAND U5036 ( .A(n4845), .B(n4844), .Z(n4846) );
  NAND U5037 ( .A(n4847), .B(n4846), .Z(n4960) );
  XNOR U5038 ( .A(n4959), .B(n4960), .Z(n4961) );
  NANDN U5039 ( .A(n4849), .B(n4848), .Z(n4853) );
  NAND U5040 ( .A(n4851), .B(n4850), .Z(n4852) );
  AND U5041 ( .A(n4853), .B(n4852), .Z(n4962) );
  XNOR U5042 ( .A(n4961), .B(n4962), .Z(n4906) );
  NANDN U5043 ( .A(n4855), .B(n4854), .Z(n4859) );
  OR U5044 ( .A(n4857), .B(n4856), .Z(n4858) );
  NAND U5045 ( .A(n4859), .B(n4858), .Z(n4956) );
  NAND U5046 ( .A(b[0]), .B(a[69]), .Z(n4860) );
  XNOR U5047 ( .A(b[1]), .B(n4860), .Z(n4862) );
  NAND U5048 ( .A(a[68]), .B(n98), .Z(n4861) );
  AND U5049 ( .A(n4862), .B(n4861), .Z(n4932) );
  XNOR U5050 ( .A(n20154), .B(n4991), .Z(n4941) );
  OR U5051 ( .A(n4941), .B(n20057), .Z(n4865) );
  NANDN U5052 ( .A(n4863), .B(n20098), .Z(n4864) );
  AND U5053 ( .A(n4865), .B(n4864), .Z(n4933) );
  XOR U5054 ( .A(n4932), .B(n4933), .Z(n4935) );
  NAND U5055 ( .A(a[53]), .B(b[15]), .Z(n4934) );
  XOR U5056 ( .A(n4935), .B(n4934), .Z(n4953) );
  NAND U5057 ( .A(n19722), .B(n4866), .Z(n4868) );
  XNOR U5058 ( .A(b[5]), .B(n5615), .Z(n4944) );
  NANDN U5059 ( .A(n19640), .B(n4944), .Z(n4867) );
  NAND U5060 ( .A(n4868), .B(n4867), .Z(n4929) );
  XNOR U5061 ( .A(n19714), .B(n5459), .Z(n4947) );
  NANDN U5062 ( .A(n4947), .B(n19766), .Z(n4871) );
  NANDN U5063 ( .A(n4869), .B(n19767), .Z(n4870) );
  NAND U5064 ( .A(n4871), .B(n4870), .Z(n4926) );
  NAND U5065 ( .A(n19554), .B(n4872), .Z(n4874) );
  IV U5066 ( .A(a[67]), .Z(n5771) );
  XNOR U5067 ( .A(b[3]), .B(n5771), .Z(n4950) );
  NANDN U5068 ( .A(n19521), .B(n4950), .Z(n4873) );
  AND U5069 ( .A(n4874), .B(n4873), .Z(n4927) );
  XNOR U5070 ( .A(n4926), .B(n4927), .Z(n4928) );
  XOR U5071 ( .A(n4929), .B(n4928), .Z(n4954) );
  XOR U5072 ( .A(n4953), .B(n4954), .Z(n4955) );
  XNOR U5073 ( .A(n4956), .B(n4955), .Z(n4904) );
  NAND U5074 ( .A(n4876), .B(n4875), .Z(n4880) );
  NAND U5075 ( .A(n4878), .B(n4877), .Z(n4879) );
  NAND U5076 ( .A(n4880), .B(n4879), .Z(n4905) );
  XOR U5077 ( .A(n4904), .B(n4905), .Z(n4907) );
  XNOR U5078 ( .A(n4906), .B(n4907), .Z(n4965) );
  NANDN U5079 ( .A(n4882), .B(n4881), .Z(n4886) );
  NAND U5080 ( .A(n4884), .B(n4883), .Z(n4885) );
  NAND U5081 ( .A(n4886), .B(n4885), .Z(n4966) );
  XNOR U5082 ( .A(n4965), .B(n4966), .Z(n4967) );
  XOR U5083 ( .A(n4968), .B(n4967), .Z(n4898) );
  NANDN U5084 ( .A(n4888), .B(n4887), .Z(n4892) );
  NANDN U5085 ( .A(n4890), .B(n4889), .Z(n4891) );
  NAND U5086 ( .A(n4892), .B(n4891), .Z(n4899) );
  XNOR U5087 ( .A(n4898), .B(n4899), .Z(n4900) );
  XNOR U5088 ( .A(n4901), .B(n4900), .Z(n4971) );
  XNOR U5089 ( .A(n4971), .B(sreg[309]), .Z(n4973) );
  NAND U5090 ( .A(n4893), .B(sreg[308]), .Z(n4897) );
  OR U5091 ( .A(n4895), .B(n4894), .Z(n4896) );
  AND U5092 ( .A(n4897), .B(n4896), .Z(n4972) );
  XOR U5093 ( .A(n4973), .B(n4972), .Z(c[309]) );
  NANDN U5094 ( .A(n4899), .B(n4898), .Z(n4903) );
  NAND U5095 ( .A(n4901), .B(n4900), .Z(n4902) );
  NAND U5096 ( .A(n4903), .B(n4902), .Z(n4979) );
  NANDN U5097 ( .A(n4905), .B(n4904), .Z(n4909) );
  OR U5098 ( .A(n4907), .B(n4906), .Z(n4908) );
  NAND U5099 ( .A(n4909), .B(n4908), .Z(n5046) );
  XNOR U5100 ( .A(n20052), .B(n5225), .Z(n4988) );
  OR U5101 ( .A(n4988), .B(n20020), .Z(n4912) );
  NANDN U5102 ( .A(n4910), .B(n19960), .Z(n4911) );
  NAND U5103 ( .A(n4912), .B(n4911), .Z(n5001) );
  XNOR U5104 ( .A(n102), .B(n4913), .Z(n4992) );
  OR U5105 ( .A(n4992), .B(n20121), .Z(n4916) );
  NANDN U5106 ( .A(n4914), .B(n20122), .Z(n4915) );
  NAND U5107 ( .A(n4916), .B(n4915), .Z(n4998) );
  XNOR U5108 ( .A(n19975), .B(n5381), .Z(n4995) );
  NANDN U5109 ( .A(n4995), .B(n19883), .Z(n4919) );
  NANDN U5110 ( .A(n4917), .B(n19937), .Z(n4918) );
  AND U5111 ( .A(n4919), .B(n4918), .Z(n4999) );
  XNOR U5112 ( .A(n4998), .B(n4999), .Z(n5000) );
  XNOR U5113 ( .A(n5001), .B(n5000), .Z(n5037) );
  NANDN U5114 ( .A(n4921), .B(n4920), .Z(n4925) );
  NAND U5115 ( .A(n4923), .B(n4922), .Z(n4924) );
  NAND U5116 ( .A(n4925), .B(n4924), .Z(n5038) );
  XNOR U5117 ( .A(n5037), .B(n5038), .Z(n5039) );
  NANDN U5118 ( .A(n4927), .B(n4926), .Z(n4931) );
  NAND U5119 ( .A(n4929), .B(n4928), .Z(n4930) );
  AND U5120 ( .A(n4931), .B(n4930), .Z(n5040) );
  XNOR U5121 ( .A(n5039), .B(n5040), .Z(n4984) );
  NANDN U5122 ( .A(n4933), .B(n4932), .Z(n4937) );
  OR U5123 ( .A(n4935), .B(n4934), .Z(n4936) );
  NAND U5124 ( .A(n4937), .B(n4936), .Z(n5034) );
  NAND U5125 ( .A(b[0]), .B(a[70]), .Z(n4938) );
  XNOR U5126 ( .A(b[1]), .B(n4938), .Z(n4940) );
  NAND U5127 ( .A(a[69]), .B(n98), .Z(n4939) );
  AND U5128 ( .A(n4940), .B(n4939), .Z(n5010) );
  XNOR U5129 ( .A(n20154), .B(n5069), .Z(n5019) );
  OR U5130 ( .A(n5019), .B(n20057), .Z(n4943) );
  NANDN U5131 ( .A(n4941), .B(n20098), .Z(n4942) );
  AND U5132 ( .A(n4943), .B(n4942), .Z(n5011) );
  XOR U5133 ( .A(n5010), .B(n5011), .Z(n5013) );
  NAND U5134 ( .A(a[54]), .B(b[15]), .Z(n5012) );
  XOR U5135 ( .A(n5013), .B(n5012), .Z(n5031) );
  NAND U5136 ( .A(n19722), .B(n4944), .Z(n4946) );
  XNOR U5137 ( .A(b[5]), .B(n5693), .Z(n5022) );
  NANDN U5138 ( .A(n19640), .B(n5022), .Z(n4945) );
  NAND U5139 ( .A(n4946), .B(n4945), .Z(n5007) );
  XNOR U5140 ( .A(n19714), .B(n5549), .Z(n5025) );
  NANDN U5141 ( .A(n5025), .B(n19766), .Z(n4949) );
  NANDN U5142 ( .A(n4947), .B(n19767), .Z(n4948) );
  NAND U5143 ( .A(n4949), .B(n4948), .Z(n5004) );
  NAND U5144 ( .A(n19554), .B(n4950), .Z(n4952) );
  IV U5145 ( .A(a[68]), .Z(n5874) );
  XNOR U5146 ( .A(b[3]), .B(n5874), .Z(n5028) );
  NANDN U5147 ( .A(n19521), .B(n5028), .Z(n4951) );
  AND U5148 ( .A(n4952), .B(n4951), .Z(n5005) );
  XNOR U5149 ( .A(n5004), .B(n5005), .Z(n5006) );
  XOR U5150 ( .A(n5007), .B(n5006), .Z(n5032) );
  XOR U5151 ( .A(n5031), .B(n5032), .Z(n5033) );
  XNOR U5152 ( .A(n5034), .B(n5033), .Z(n4982) );
  NAND U5153 ( .A(n4954), .B(n4953), .Z(n4958) );
  NAND U5154 ( .A(n4956), .B(n4955), .Z(n4957) );
  NAND U5155 ( .A(n4958), .B(n4957), .Z(n4983) );
  XOR U5156 ( .A(n4982), .B(n4983), .Z(n4985) );
  XNOR U5157 ( .A(n4984), .B(n4985), .Z(n5043) );
  NANDN U5158 ( .A(n4960), .B(n4959), .Z(n4964) );
  NAND U5159 ( .A(n4962), .B(n4961), .Z(n4963) );
  NAND U5160 ( .A(n4964), .B(n4963), .Z(n5044) );
  XNOR U5161 ( .A(n5043), .B(n5044), .Z(n5045) );
  XOR U5162 ( .A(n5046), .B(n5045), .Z(n4976) );
  NANDN U5163 ( .A(n4966), .B(n4965), .Z(n4970) );
  NANDN U5164 ( .A(n4968), .B(n4967), .Z(n4969) );
  NAND U5165 ( .A(n4970), .B(n4969), .Z(n4977) );
  XNOR U5166 ( .A(n4976), .B(n4977), .Z(n4978) );
  XNOR U5167 ( .A(n4979), .B(n4978), .Z(n5049) );
  XNOR U5168 ( .A(n5049), .B(sreg[310]), .Z(n5051) );
  NAND U5169 ( .A(n4971), .B(sreg[309]), .Z(n4975) );
  OR U5170 ( .A(n4973), .B(n4972), .Z(n4974) );
  AND U5171 ( .A(n4975), .B(n4974), .Z(n5050) );
  XOR U5172 ( .A(n5051), .B(n5050), .Z(c[310]) );
  NANDN U5173 ( .A(n4977), .B(n4976), .Z(n4981) );
  NAND U5174 ( .A(n4979), .B(n4978), .Z(n4980) );
  NAND U5175 ( .A(n4981), .B(n4980), .Z(n5057) );
  NANDN U5176 ( .A(n4983), .B(n4982), .Z(n4987) );
  OR U5177 ( .A(n4985), .B(n4984), .Z(n4986) );
  NAND U5178 ( .A(n4987), .B(n4986), .Z(n5124) );
  XNOR U5179 ( .A(n20052), .B(n5303), .Z(n5066) );
  OR U5180 ( .A(n5066), .B(n20020), .Z(n4990) );
  NANDN U5181 ( .A(n4988), .B(n19960), .Z(n4989) );
  NAND U5182 ( .A(n4990), .B(n4989), .Z(n5079) );
  XNOR U5183 ( .A(n102), .B(n4991), .Z(n5070) );
  OR U5184 ( .A(n5070), .B(n20121), .Z(n4994) );
  NANDN U5185 ( .A(n4992), .B(n20122), .Z(n4993) );
  NAND U5186 ( .A(n4994), .B(n4993), .Z(n5076) );
  XNOR U5187 ( .A(n19975), .B(n5459), .Z(n5073) );
  NANDN U5188 ( .A(n5073), .B(n19883), .Z(n4997) );
  NANDN U5189 ( .A(n4995), .B(n19937), .Z(n4996) );
  AND U5190 ( .A(n4997), .B(n4996), .Z(n5077) );
  XNOR U5191 ( .A(n5076), .B(n5077), .Z(n5078) );
  XNOR U5192 ( .A(n5079), .B(n5078), .Z(n5115) );
  NANDN U5193 ( .A(n4999), .B(n4998), .Z(n5003) );
  NAND U5194 ( .A(n5001), .B(n5000), .Z(n5002) );
  NAND U5195 ( .A(n5003), .B(n5002), .Z(n5116) );
  XNOR U5196 ( .A(n5115), .B(n5116), .Z(n5117) );
  NANDN U5197 ( .A(n5005), .B(n5004), .Z(n5009) );
  NAND U5198 ( .A(n5007), .B(n5006), .Z(n5008) );
  AND U5199 ( .A(n5009), .B(n5008), .Z(n5118) );
  XNOR U5200 ( .A(n5117), .B(n5118), .Z(n5062) );
  NANDN U5201 ( .A(n5011), .B(n5010), .Z(n5015) );
  OR U5202 ( .A(n5013), .B(n5012), .Z(n5014) );
  NAND U5203 ( .A(n5015), .B(n5014), .Z(n5112) );
  NAND U5204 ( .A(b[0]), .B(a[71]), .Z(n5016) );
  XNOR U5205 ( .A(b[1]), .B(n5016), .Z(n5018) );
  NAND U5206 ( .A(a[70]), .B(n98), .Z(n5017) );
  AND U5207 ( .A(n5018), .B(n5017), .Z(n5088) );
  XNOR U5208 ( .A(n20154), .B(n5147), .Z(n5097) );
  OR U5209 ( .A(n5097), .B(n20057), .Z(n5021) );
  NANDN U5210 ( .A(n5019), .B(n20098), .Z(n5020) );
  AND U5211 ( .A(n5021), .B(n5020), .Z(n5089) );
  XOR U5212 ( .A(n5088), .B(n5089), .Z(n5091) );
  NAND U5213 ( .A(a[55]), .B(b[15]), .Z(n5090) );
  XOR U5214 ( .A(n5091), .B(n5090), .Z(n5109) );
  NAND U5215 ( .A(n19722), .B(n5022), .Z(n5024) );
  XNOR U5216 ( .A(b[5]), .B(n5771), .Z(n5100) );
  NANDN U5217 ( .A(n19640), .B(n5100), .Z(n5023) );
  NAND U5218 ( .A(n5024), .B(n5023), .Z(n5085) );
  XNOR U5219 ( .A(n19714), .B(n5615), .Z(n5103) );
  NANDN U5220 ( .A(n5103), .B(n19766), .Z(n5027) );
  NANDN U5221 ( .A(n5025), .B(n19767), .Z(n5026) );
  NAND U5222 ( .A(n5027), .B(n5026), .Z(n5082) );
  NAND U5223 ( .A(n19554), .B(n5028), .Z(n5030) );
  IV U5224 ( .A(a[69]), .Z(n5925) );
  XNOR U5225 ( .A(b[3]), .B(n5925), .Z(n5106) );
  NANDN U5226 ( .A(n19521), .B(n5106), .Z(n5029) );
  AND U5227 ( .A(n5030), .B(n5029), .Z(n5083) );
  XNOR U5228 ( .A(n5082), .B(n5083), .Z(n5084) );
  XOR U5229 ( .A(n5085), .B(n5084), .Z(n5110) );
  XOR U5230 ( .A(n5109), .B(n5110), .Z(n5111) );
  XNOR U5231 ( .A(n5112), .B(n5111), .Z(n5060) );
  NAND U5232 ( .A(n5032), .B(n5031), .Z(n5036) );
  NAND U5233 ( .A(n5034), .B(n5033), .Z(n5035) );
  NAND U5234 ( .A(n5036), .B(n5035), .Z(n5061) );
  XOR U5235 ( .A(n5060), .B(n5061), .Z(n5063) );
  XNOR U5236 ( .A(n5062), .B(n5063), .Z(n5121) );
  NANDN U5237 ( .A(n5038), .B(n5037), .Z(n5042) );
  NAND U5238 ( .A(n5040), .B(n5039), .Z(n5041) );
  NAND U5239 ( .A(n5042), .B(n5041), .Z(n5122) );
  XNOR U5240 ( .A(n5121), .B(n5122), .Z(n5123) );
  XOR U5241 ( .A(n5124), .B(n5123), .Z(n5054) );
  NANDN U5242 ( .A(n5044), .B(n5043), .Z(n5048) );
  NANDN U5243 ( .A(n5046), .B(n5045), .Z(n5047) );
  NAND U5244 ( .A(n5048), .B(n5047), .Z(n5055) );
  XNOR U5245 ( .A(n5054), .B(n5055), .Z(n5056) );
  XNOR U5246 ( .A(n5057), .B(n5056), .Z(n5127) );
  XNOR U5247 ( .A(n5127), .B(sreg[311]), .Z(n5129) );
  NAND U5248 ( .A(n5049), .B(sreg[310]), .Z(n5053) );
  OR U5249 ( .A(n5051), .B(n5050), .Z(n5052) );
  AND U5250 ( .A(n5053), .B(n5052), .Z(n5128) );
  XOR U5251 ( .A(n5129), .B(n5128), .Z(c[311]) );
  NANDN U5252 ( .A(n5055), .B(n5054), .Z(n5059) );
  NAND U5253 ( .A(n5057), .B(n5056), .Z(n5058) );
  NAND U5254 ( .A(n5059), .B(n5058), .Z(n5135) );
  NANDN U5255 ( .A(n5061), .B(n5060), .Z(n5065) );
  OR U5256 ( .A(n5063), .B(n5062), .Z(n5064) );
  NAND U5257 ( .A(n5065), .B(n5064), .Z(n5202) );
  XNOR U5258 ( .A(n20052), .B(n5381), .Z(n5144) );
  OR U5259 ( .A(n5144), .B(n20020), .Z(n5068) );
  NANDN U5260 ( .A(n5066), .B(n19960), .Z(n5067) );
  NAND U5261 ( .A(n5068), .B(n5067), .Z(n5157) );
  XNOR U5262 ( .A(n102), .B(n5069), .Z(n5148) );
  OR U5263 ( .A(n5148), .B(n20121), .Z(n5072) );
  NANDN U5264 ( .A(n5070), .B(n20122), .Z(n5071) );
  NAND U5265 ( .A(n5072), .B(n5071), .Z(n5154) );
  XNOR U5266 ( .A(n19975), .B(n5549), .Z(n5151) );
  NANDN U5267 ( .A(n5151), .B(n19883), .Z(n5075) );
  NANDN U5268 ( .A(n5073), .B(n19937), .Z(n5074) );
  AND U5269 ( .A(n5075), .B(n5074), .Z(n5155) );
  XNOR U5270 ( .A(n5154), .B(n5155), .Z(n5156) );
  XNOR U5271 ( .A(n5157), .B(n5156), .Z(n5193) );
  NANDN U5272 ( .A(n5077), .B(n5076), .Z(n5081) );
  NAND U5273 ( .A(n5079), .B(n5078), .Z(n5080) );
  NAND U5274 ( .A(n5081), .B(n5080), .Z(n5194) );
  XNOR U5275 ( .A(n5193), .B(n5194), .Z(n5195) );
  NANDN U5276 ( .A(n5083), .B(n5082), .Z(n5087) );
  NAND U5277 ( .A(n5085), .B(n5084), .Z(n5086) );
  AND U5278 ( .A(n5087), .B(n5086), .Z(n5196) );
  XNOR U5279 ( .A(n5195), .B(n5196), .Z(n5140) );
  NANDN U5280 ( .A(n5089), .B(n5088), .Z(n5093) );
  OR U5281 ( .A(n5091), .B(n5090), .Z(n5092) );
  NAND U5282 ( .A(n5093), .B(n5092), .Z(n5190) );
  NAND U5283 ( .A(b[0]), .B(a[72]), .Z(n5094) );
  XNOR U5284 ( .A(b[1]), .B(n5094), .Z(n5096) );
  NAND U5285 ( .A(a[71]), .B(n98), .Z(n5095) );
  AND U5286 ( .A(n5096), .B(n5095), .Z(n5166) );
  XNOR U5287 ( .A(n20154), .B(n5225), .Z(n5175) );
  OR U5288 ( .A(n5175), .B(n20057), .Z(n5099) );
  NANDN U5289 ( .A(n5097), .B(n20098), .Z(n5098) );
  AND U5290 ( .A(n5099), .B(n5098), .Z(n5167) );
  XOR U5291 ( .A(n5166), .B(n5167), .Z(n5169) );
  NAND U5292 ( .A(a[56]), .B(b[15]), .Z(n5168) );
  XOR U5293 ( .A(n5169), .B(n5168), .Z(n5187) );
  NAND U5294 ( .A(n19722), .B(n5100), .Z(n5102) );
  XNOR U5295 ( .A(b[5]), .B(n5874), .Z(n5178) );
  NANDN U5296 ( .A(n19640), .B(n5178), .Z(n5101) );
  NAND U5297 ( .A(n5102), .B(n5101), .Z(n5163) );
  XNOR U5298 ( .A(n19714), .B(n5693), .Z(n5181) );
  NANDN U5299 ( .A(n5181), .B(n19766), .Z(n5105) );
  NANDN U5300 ( .A(n5103), .B(n19767), .Z(n5104) );
  NAND U5301 ( .A(n5105), .B(n5104), .Z(n5160) );
  NAND U5302 ( .A(n19554), .B(n5106), .Z(n5108) );
  IV U5303 ( .A(a[70]), .Z(n6030) );
  XNOR U5304 ( .A(b[3]), .B(n6030), .Z(n5184) );
  NANDN U5305 ( .A(n19521), .B(n5184), .Z(n5107) );
  AND U5306 ( .A(n5108), .B(n5107), .Z(n5161) );
  XNOR U5307 ( .A(n5160), .B(n5161), .Z(n5162) );
  XOR U5308 ( .A(n5163), .B(n5162), .Z(n5188) );
  XOR U5309 ( .A(n5187), .B(n5188), .Z(n5189) );
  XNOR U5310 ( .A(n5190), .B(n5189), .Z(n5138) );
  NAND U5311 ( .A(n5110), .B(n5109), .Z(n5114) );
  NAND U5312 ( .A(n5112), .B(n5111), .Z(n5113) );
  NAND U5313 ( .A(n5114), .B(n5113), .Z(n5139) );
  XOR U5314 ( .A(n5138), .B(n5139), .Z(n5141) );
  XNOR U5315 ( .A(n5140), .B(n5141), .Z(n5199) );
  NANDN U5316 ( .A(n5116), .B(n5115), .Z(n5120) );
  NAND U5317 ( .A(n5118), .B(n5117), .Z(n5119) );
  NAND U5318 ( .A(n5120), .B(n5119), .Z(n5200) );
  XNOR U5319 ( .A(n5199), .B(n5200), .Z(n5201) );
  XOR U5320 ( .A(n5202), .B(n5201), .Z(n5132) );
  NANDN U5321 ( .A(n5122), .B(n5121), .Z(n5126) );
  NANDN U5322 ( .A(n5124), .B(n5123), .Z(n5125) );
  NAND U5323 ( .A(n5126), .B(n5125), .Z(n5133) );
  XNOR U5324 ( .A(n5132), .B(n5133), .Z(n5134) );
  XNOR U5325 ( .A(n5135), .B(n5134), .Z(n5205) );
  XNOR U5326 ( .A(n5205), .B(sreg[312]), .Z(n5207) );
  NAND U5327 ( .A(n5127), .B(sreg[311]), .Z(n5131) );
  OR U5328 ( .A(n5129), .B(n5128), .Z(n5130) );
  AND U5329 ( .A(n5131), .B(n5130), .Z(n5206) );
  XOR U5330 ( .A(n5207), .B(n5206), .Z(c[312]) );
  NANDN U5331 ( .A(n5133), .B(n5132), .Z(n5137) );
  NAND U5332 ( .A(n5135), .B(n5134), .Z(n5136) );
  NAND U5333 ( .A(n5137), .B(n5136), .Z(n5213) );
  NANDN U5334 ( .A(n5139), .B(n5138), .Z(n5143) );
  OR U5335 ( .A(n5141), .B(n5140), .Z(n5142) );
  NAND U5336 ( .A(n5143), .B(n5142), .Z(n5280) );
  XNOR U5337 ( .A(n20052), .B(n5459), .Z(n5222) );
  OR U5338 ( .A(n5222), .B(n20020), .Z(n5146) );
  NANDN U5339 ( .A(n5144), .B(n19960), .Z(n5145) );
  NAND U5340 ( .A(n5146), .B(n5145), .Z(n5235) );
  XNOR U5341 ( .A(n102), .B(n5147), .Z(n5226) );
  OR U5342 ( .A(n5226), .B(n20121), .Z(n5150) );
  NANDN U5343 ( .A(n5148), .B(n20122), .Z(n5149) );
  NAND U5344 ( .A(n5150), .B(n5149), .Z(n5232) );
  XNOR U5345 ( .A(n19975), .B(n5615), .Z(n5229) );
  NANDN U5346 ( .A(n5229), .B(n19883), .Z(n5153) );
  NANDN U5347 ( .A(n5151), .B(n19937), .Z(n5152) );
  AND U5348 ( .A(n5153), .B(n5152), .Z(n5233) );
  XNOR U5349 ( .A(n5232), .B(n5233), .Z(n5234) );
  XNOR U5350 ( .A(n5235), .B(n5234), .Z(n5271) );
  NANDN U5351 ( .A(n5155), .B(n5154), .Z(n5159) );
  NAND U5352 ( .A(n5157), .B(n5156), .Z(n5158) );
  NAND U5353 ( .A(n5159), .B(n5158), .Z(n5272) );
  XNOR U5354 ( .A(n5271), .B(n5272), .Z(n5273) );
  NANDN U5355 ( .A(n5161), .B(n5160), .Z(n5165) );
  NAND U5356 ( .A(n5163), .B(n5162), .Z(n5164) );
  AND U5357 ( .A(n5165), .B(n5164), .Z(n5274) );
  XNOR U5358 ( .A(n5273), .B(n5274), .Z(n5218) );
  NANDN U5359 ( .A(n5167), .B(n5166), .Z(n5171) );
  OR U5360 ( .A(n5169), .B(n5168), .Z(n5170) );
  NAND U5361 ( .A(n5171), .B(n5170), .Z(n5268) );
  NAND U5362 ( .A(b[0]), .B(a[73]), .Z(n5172) );
  XNOR U5363 ( .A(b[1]), .B(n5172), .Z(n5174) );
  NAND U5364 ( .A(a[72]), .B(n98), .Z(n5173) );
  AND U5365 ( .A(n5174), .B(n5173), .Z(n5244) );
  XNOR U5366 ( .A(n20154), .B(n5303), .Z(n5250) );
  OR U5367 ( .A(n5250), .B(n20057), .Z(n5177) );
  NANDN U5368 ( .A(n5175), .B(n20098), .Z(n5176) );
  AND U5369 ( .A(n5177), .B(n5176), .Z(n5245) );
  XOR U5370 ( .A(n5244), .B(n5245), .Z(n5247) );
  NAND U5371 ( .A(a[57]), .B(b[15]), .Z(n5246) );
  XOR U5372 ( .A(n5247), .B(n5246), .Z(n5265) );
  NAND U5373 ( .A(n19722), .B(n5178), .Z(n5180) );
  XNOR U5374 ( .A(b[5]), .B(n5925), .Z(n5256) );
  NANDN U5375 ( .A(n19640), .B(n5256), .Z(n5179) );
  NAND U5376 ( .A(n5180), .B(n5179), .Z(n5241) );
  XNOR U5377 ( .A(n19714), .B(n5771), .Z(n5259) );
  NANDN U5378 ( .A(n5259), .B(n19766), .Z(n5183) );
  NANDN U5379 ( .A(n5181), .B(n19767), .Z(n5182) );
  NAND U5380 ( .A(n5183), .B(n5182), .Z(n5238) );
  NAND U5381 ( .A(n19554), .B(n5184), .Z(n5186) );
  IV U5382 ( .A(a[71]), .Z(n6108) );
  XNOR U5383 ( .A(b[3]), .B(n6108), .Z(n5262) );
  NANDN U5384 ( .A(n19521), .B(n5262), .Z(n5185) );
  AND U5385 ( .A(n5186), .B(n5185), .Z(n5239) );
  XNOR U5386 ( .A(n5238), .B(n5239), .Z(n5240) );
  XOR U5387 ( .A(n5241), .B(n5240), .Z(n5266) );
  XOR U5388 ( .A(n5265), .B(n5266), .Z(n5267) );
  XNOR U5389 ( .A(n5268), .B(n5267), .Z(n5216) );
  NAND U5390 ( .A(n5188), .B(n5187), .Z(n5192) );
  NAND U5391 ( .A(n5190), .B(n5189), .Z(n5191) );
  NAND U5392 ( .A(n5192), .B(n5191), .Z(n5217) );
  XOR U5393 ( .A(n5216), .B(n5217), .Z(n5219) );
  XNOR U5394 ( .A(n5218), .B(n5219), .Z(n5277) );
  NANDN U5395 ( .A(n5194), .B(n5193), .Z(n5198) );
  NAND U5396 ( .A(n5196), .B(n5195), .Z(n5197) );
  NAND U5397 ( .A(n5198), .B(n5197), .Z(n5278) );
  XNOR U5398 ( .A(n5277), .B(n5278), .Z(n5279) );
  XOR U5399 ( .A(n5280), .B(n5279), .Z(n5210) );
  NANDN U5400 ( .A(n5200), .B(n5199), .Z(n5204) );
  NANDN U5401 ( .A(n5202), .B(n5201), .Z(n5203) );
  NAND U5402 ( .A(n5204), .B(n5203), .Z(n5211) );
  XNOR U5403 ( .A(n5210), .B(n5211), .Z(n5212) );
  XNOR U5404 ( .A(n5213), .B(n5212), .Z(n5283) );
  XNOR U5405 ( .A(n5283), .B(sreg[313]), .Z(n5285) );
  NAND U5406 ( .A(n5205), .B(sreg[312]), .Z(n5209) );
  OR U5407 ( .A(n5207), .B(n5206), .Z(n5208) );
  AND U5408 ( .A(n5209), .B(n5208), .Z(n5284) );
  XOR U5409 ( .A(n5285), .B(n5284), .Z(c[313]) );
  NANDN U5410 ( .A(n5211), .B(n5210), .Z(n5215) );
  NAND U5411 ( .A(n5213), .B(n5212), .Z(n5214) );
  NAND U5412 ( .A(n5215), .B(n5214), .Z(n5291) );
  NANDN U5413 ( .A(n5217), .B(n5216), .Z(n5221) );
  OR U5414 ( .A(n5219), .B(n5218), .Z(n5220) );
  NAND U5415 ( .A(n5221), .B(n5220), .Z(n5358) );
  XNOR U5416 ( .A(n20052), .B(n5549), .Z(n5300) );
  OR U5417 ( .A(n5300), .B(n20020), .Z(n5224) );
  NANDN U5418 ( .A(n5222), .B(n19960), .Z(n5223) );
  NAND U5419 ( .A(n5224), .B(n5223), .Z(n5313) );
  XNOR U5420 ( .A(n102), .B(n5225), .Z(n5304) );
  OR U5421 ( .A(n5304), .B(n20121), .Z(n5228) );
  NANDN U5422 ( .A(n5226), .B(n20122), .Z(n5227) );
  NAND U5423 ( .A(n5228), .B(n5227), .Z(n5310) );
  XNOR U5424 ( .A(n19975), .B(n5693), .Z(n5307) );
  NANDN U5425 ( .A(n5307), .B(n19883), .Z(n5231) );
  NANDN U5426 ( .A(n5229), .B(n19937), .Z(n5230) );
  AND U5427 ( .A(n5231), .B(n5230), .Z(n5311) );
  XNOR U5428 ( .A(n5310), .B(n5311), .Z(n5312) );
  XNOR U5429 ( .A(n5313), .B(n5312), .Z(n5349) );
  NANDN U5430 ( .A(n5233), .B(n5232), .Z(n5237) );
  NAND U5431 ( .A(n5235), .B(n5234), .Z(n5236) );
  NAND U5432 ( .A(n5237), .B(n5236), .Z(n5350) );
  XNOR U5433 ( .A(n5349), .B(n5350), .Z(n5351) );
  NANDN U5434 ( .A(n5239), .B(n5238), .Z(n5243) );
  NAND U5435 ( .A(n5241), .B(n5240), .Z(n5242) );
  AND U5436 ( .A(n5243), .B(n5242), .Z(n5352) );
  XNOR U5437 ( .A(n5351), .B(n5352), .Z(n5296) );
  NANDN U5438 ( .A(n5245), .B(n5244), .Z(n5249) );
  OR U5439 ( .A(n5247), .B(n5246), .Z(n5248) );
  NAND U5440 ( .A(n5249), .B(n5248), .Z(n5346) );
  XNOR U5441 ( .A(n20154), .B(n5381), .Z(n5331) );
  OR U5442 ( .A(n5331), .B(n20057), .Z(n5252) );
  NANDN U5443 ( .A(n5250), .B(n20098), .Z(n5251) );
  AND U5444 ( .A(n5252), .B(n5251), .Z(n5323) );
  NAND U5445 ( .A(b[0]), .B(a[74]), .Z(n5253) );
  XNOR U5446 ( .A(b[1]), .B(n5253), .Z(n5255) );
  NAND U5447 ( .A(a[73]), .B(n98), .Z(n5254) );
  AND U5448 ( .A(n5255), .B(n5254), .Z(n5322) );
  XOR U5449 ( .A(n5323), .B(n5322), .Z(n5325) );
  NAND U5450 ( .A(a[58]), .B(b[15]), .Z(n5324) );
  XOR U5451 ( .A(n5325), .B(n5324), .Z(n5343) );
  NAND U5452 ( .A(n19722), .B(n5256), .Z(n5258) );
  XNOR U5453 ( .A(b[5]), .B(n6030), .Z(n5334) );
  NANDN U5454 ( .A(n19640), .B(n5334), .Z(n5257) );
  NAND U5455 ( .A(n5258), .B(n5257), .Z(n5319) );
  XNOR U5456 ( .A(n19714), .B(n5874), .Z(n5337) );
  NANDN U5457 ( .A(n5337), .B(n19766), .Z(n5261) );
  NANDN U5458 ( .A(n5259), .B(n19767), .Z(n5260) );
  NAND U5459 ( .A(n5261), .B(n5260), .Z(n5316) );
  NAND U5460 ( .A(n19554), .B(n5262), .Z(n5264) );
  IV U5461 ( .A(a[72]), .Z(n6186) );
  XNOR U5462 ( .A(b[3]), .B(n6186), .Z(n5340) );
  NANDN U5463 ( .A(n19521), .B(n5340), .Z(n5263) );
  AND U5464 ( .A(n5264), .B(n5263), .Z(n5317) );
  XNOR U5465 ( .A(n5316), .B(n5317), .Z(n5318) );
  XOR U5466 ( .A(n5319), .B(n5318), .Z(n5344) );
  XOR U5467 ( .A(n5343), .B(n5344), .Z(n5345) );
  XNOR U5468 ( .A(n5346), .B(n5345), .Z(n5294) );
  NAND U5469 ( .A(n5266), .B(n5265), .Z(n5270) );
  NAND U5470 ( .A(n5268), .B(n5267), .Z(n5269) );
  NAND U5471 ( .A(n5270), .B(n5269), .Z(n5295) );
  XOR U5472 ( .A(n5294), .B(n5295), .Z(n5297) );
  XNOR U5473 ( .A(n5296), .B(n5297), .Z(n5355) );
  NANDN U5474 ( .A(n5272), .B(n5271), .Z(n5276) );
  NAND U5475 ( .A(n5274), .B(n5273), .Z(n5275) );
  NAND U5476 ( .A(n5276), .B(n5275), .Z(n5356) );
  XNOR U5477 ( .A(n5355), .B(n5356), .Z(n5357) );
  XOR U5478 ( .A(n5358), .B(n5357), .Z(n5288) );
  NANDN U5479 ( .A(n5278), .B(n5277), .Z(n5282) );
  NANDN U5480 ( .A(n5280), .B(n5279), .Z(n5281) );
  NAND U5481 ( .A(n5282), .B(n5281), .Z(n5289) );
  XNOR U5482 ( .A(n5288), .B(n5289), .Z(n5290) );
  XNOR U5483 ( .A(n5291), .B(n5290), .Z(n5361) );
  XNOR U5484 ( .A(n5361), .B(sreg[314]), .Z(n5363) );
  NAND U5485 ( .A(n5283), .B(sreg[313]), .Z(n5287) );
  OR U5486 ( .A(n5285), .B(n5284), .Z(n5286) );
  AND U5487 ( .A(n5287), .B(n5286), .Z(n5362) );
  XOR U5488 ( .A(n5363), .B(n5362), .Z(c[314]) );
  NANDN U5489 ( .A(n5289), .B(n5288), .Z(n5293) );
  NAND U5490 ( .A(n5291), .B(n5290), .Z(n5292) );
  NAND U5491 ( .A(n5293), .B(n5292), .Z(n5369) );
  NANDN U5492 ( .A(n5295), .B(n5294), .Z(n5299) );
  OR U5493 ( .A(n5297), .B(n5296), .Z(n5298) );
  NAND U5494 ( .A(n5299), .B(n5298), .Z(n5436) );
  XNOR U5495 ( .A(n20052), .B(n5615), .Z(n5378) );
  OR U5496 ( .A(n5378), .B(n20020), .Z(n5302) );
  NANDN U5497 ( .A(n5300), .B(n19960), .Z(n5301) );
  NAND U5498 ( .A(n5302), .B(n5301), .Z(n5391) );
  XNOR U5499 ( .A(n102), .B(n5303), .Z(n5382) );
  OR U5500 ( .A(n5382), .B(n20121), .Z(n5306) );
  NANDN U5501 ( .A(n5304), .B(n20122), .Z(n5305) );
  NAND U5502 ( .A(n5306), .B(n5305), .Z(n5388) );
  XNOR U5503 ( .A(n19975), .B(n5771), .Z(n5385) );
  NANDN U5504 ( .A(n5385), .B(n19883), .Z(n5309) );
  NANDN U5505 ( .A(n5307), .B(n19937), .Z(n5308) );
  AND U5506 ( .A(n5309), .B(n5308), .Z(n5389) );
  XNOR U5507 ( .A(n5388), .B(n5389), .Z(n5390) );
  XNOR U5508 ( .A(n5391), .B(n5390), .Z(n5427) );
  NANDN U5509 ( .A(n5311), .B(n5310), .Z(n5315) );
  NAND U5510 ( .A(n5313), .B(n5312), .Z(n5314) );
  NAND U5511 ( .A(n5315), .B(n5314), .Z(n5428) );
  XNOR U5512 ( .A(n5427), .B(n5428), .Z(n5429) );
  NANDN U5513 ( .A(n5317), .B(n5316), .Z(n5321) );
  NAND U5514 ( .A(n5319), .B(n5318), .Z(n5320) );
  AND U5515 ( .A(n5321), .B(n5320), .Z(n5430) );
  XNOR U5516 ( .A(n5429), .B(n5430), .Z(n5374) );
  NANDN U5517 ( .A(n5323), .B(n5322), .Z(n5327) );
  OR U5518 ( .A(n5325), .B(n5324), .Z(n5326) );
  NAND U5519 ( .A(n5327), .B(n5326), .Z(n5424) );
  NAND U5520 ( .A(b[0]), .B(a[75]), .Z(n5328) );
  XNOR U5521 ( .A(b[1]), .B(n5328), .Z(n5330) );
  NAND U5522 ( .A(a[74]), .B(n98), .Z(n5329) );
  AND U5523 ( .A(n5330), .B(n5329), .Z(n5400) );
  XNOR U5524 ( .A(n20154), .B(n5459), .Z(n5409) );
  OR U5525 ( .A(n5409), .B(n20057), .Z(n5333) );
  NANDN U5526 ( .A(n5331), .B(n20098), .Z(n5332) );
  AND U5527 ( .A(n5333), .B(n5332), .Z(n5401) );
  XOR U5528 ( .A(n5400), .B(n5401), .Z(n5403) );
  NAND U5529 ( .A(a[59]), .B(b[15]), .Z(n5402) );
  XOR U5530 ( .A(n5403), .B(n5402), .Z(n5421) );
  NAND U5531 ( .A(n19722), .B(n5334), .Z(n5336) );
  XNOR U5532 ( .A(b[5]), .B(n6108), .Z(n5412) );
  NANDN U5533 ( .A(n19640), .B(n5412), .Z(n5335) );
  NAND U5534 ( .A(n5336), .B(n5335), .Z(n5397) );
  XNOR U5535 ( .A(n19714), .B(n5925), .Z(n5415) );
  NANDN U5536 ( .A(n5415), .B(n19766), .Z(n5339) );
  NANDN U5537 ( .A(n5337), .B(n19767), .Z(n5338) );
  NAND U5538 ( .A(n5339), .B(n5338), .Z(n5394) );
  NAND U5539 ( .A(n19554), .B(n5340), .Z(n5342) );
  IV U5540 ( .A(a[73]), .Z(n6237) );
  XNOR U5541 ( .A(b[3]), .B(n6237), .Z(n5418) );
  NANDN U5542 ( .A(n19521), .B(n5418), .Z(n5341) );
  AND U5543 ( .A(n5342), .B(n5341), .Z(n5395) );
  XNOR U5544 ( .A(n5394), .B(n5395), .Z(n5396) );
  XOR U5545 ( .A(n5397), .B(n5396), .Z(n5422) );
  XOR U5546 ( .A(n5421), .B(n5422), .Z(n5423) );
  XNOR U5547 ( .A(n5424), .B(n5423), .Z(n5372) );
  NAND U5548 ( .A(n5344), .B(n5343), .Z(n5348) );
  NAND U5549 ( .A(n5346), .B(n5345), .Z(n5347) );
  NAND U5550 ( .A(n5348), .B(n5347), .Z(n5373) );
  XOR U5551 ( .A(n5372), .B(n5373), .Z(n5375) );
  XNOR U5552 ( .A(n5374), .B(n5375), .Z(n5433) );
  NANDN U5553 ( .A(n5350), .B(n5349), .Z(n5354) );
  NAND U5554 ( .A(n5352), .B(n5351), .Z(n5353) );
  NAND U5555 ( .A(n5354), .B(n5353), .Z(n5434) );
  XNOR U5556 ( .A(n5433), .B(n5434), .Z(n5435) );
  XOR U5557 ( .A(n5436), .B(n5435), .Z(n5366) );
  NANDN U5558 ( .A(n5356), .B(n5355), .Z(n5360) );
  NANDN U5559 ( .A(n5358), .B(n5357), .Z(n5359) );
  NAND U5560 ( .A(n5360), .B(n5359), .Z(n5367) );
  XNOR U5561 ( .A(n5366), .B(n5367), .Z(n5368) );
  XNOR U5562 ( .A(n5369), .B(n5368), .Z(n5439) );
  XNOR U5563 ( .A(n5439), .B(sreg[315]), .Z(n5441) );
  NAND U5564 ( .A(n5361), .B(sreg[314]), .Z(n5365) );
  OR U5565 ( .A(n5363), .B(n5362), .Z(n5364) );
  AND U5566 ( .A(n5365), .B(n5364), .Z(n5440) );
  XOR U5567 ( .A(n5441), .B(n5440), .Z(c[315]) );
  NANDN U5568 ( .A(n5367), .B(n5366), .Z(n5371) );
  NAND U5569 ( .A(n5369), .B(n5368), .Z(n5370) );
  NAND U5570 ( .A(n5371), .B(n5370), .Z(n5447) );
  NANDN U5571 ( .A(n5373), .B(n5372), .Z(n5377) );
  OR U5572 ( .A(n5375), .B(n5374), .Z(n5376) );
  NAND U5573 ( .A(n5377), .B(n5376), .Z(n5514) );
  XNOR U5574 ( .A(n20052), .B(n5693), .Z(n5456) );
  OR U5575 ( .A(n5456), .B(n20020), .Z(n5380) );
  NANDN U5576 ( .A(n5378), .B(n19960), .Z(n5379) );
  NAND U5577 ( .A(n5380), .B(n5379), .Z(n5469) );
  XNOR U5578 ( .A(n102), .B(n5381), .Z(n5460) );
  OR U5579 ( .A(n5460), .B(n20121), .Z(n5384) );
  NANDN U5580 ( .A(n5382), .B(n20122), .Z(n5383) );
  NAND U5581 ( .A(n5384), .B(n5383), .Z(n5466) );
  XNOR U5582 ( .A(n19975), .B(n5874), .Z(n5463) );
  NANDN U5583 ( .A(n5463), .B(n19883), .Z(n5387) );
  NANDN U5584 ( .A(n5385), .B(n19937), .Z(n5386) );
  AND U5585 ( .A(n5387), .B(n5386), .Z(n5467) );
  XNOR U5586 ( .A(n5466), .B(n5467), .Z(n5468) );
  XNOR U5587 ( .A(n5469), .B(n5468), .Z(n5505) );
  NANDN U5588 ( .A(n5389), .B(n5388), .Z(n5393) );
  NAND U5589 ( .A(n5391), .B(n5390), .Z(n5392) );
  NAND U5590 ( .A(n5393), .B(n5392), .Z(n5506) );
  XNOR U5591 ( .A(n5505), .B(n5506), .Z(n5507) );
  NANDN U5592 ( .A(n5395), .B(n5394), .Z(n5399) );
  NAND U5593 ( .A(n5397), .B(n5396), .Z(n5398) );
  AND U5594 ( .A(n5399), .B(n5398), .Z(n5508) );
  XNOR U5595 ( .A(n5507), .B(n5508), .Z(n5452) );
  NANDN U5596 ( .A(n5401), .B(n5400), .Z(n5405) );
  OR U5597 ( .A(n5403), .B(n5402), .Z(n5404) );
  NAND U5598 ( .A(n5405), .B(n5404), .Z(n5502) );
  NAND U5599 ( .A(b[0]), .B(a[76]), .Z(n5406) );
  XNOR U5600 ( .A(b[1]), .B(n5406), .Z(n5408) );
  NAND U5601 ( .A(a[75]), .B(n98), .Z(n5407) );
  AND U5602 ( .A(n5408), .B(n5407), .Z(n5478) );
  XNOR U5603 ( .A(n20154), .B(n5549), .Z(n5487) );
  OR U5604 ( .A(n5487), .B(n20057), .Z(n5411) );
  NANDN U5605 ( .A(n5409), .B(n20098), .Z(n5410) );
  AND U5606 ( .A(n5411), .B(n5410), .Z(n5479) );
  XOR U5607 ( .A(n5478), .B(n5479), .Z(n5481) );
  NAND U5608 ( .A(a[60]), .B(b[15]), .Z(n5480) );
  XOR U5609 ( .A(n5481), .B(n5480), .Z(n5499) );
  NAND U5610 ( .A(n19722), .B(n5412), .Z(n5414) );
  XNOR U5611 ( .A(b[5]), .B(n6186), .Z(n5490) );
  NANDN U5612 ( .A(n19640), .B(n5490), .Z(n5413) );
  NAND U5613 ( .A(n5414), .B(n5413), .Z(n5475) );
  XNOR U5614 ( .A(n19714), .B(n6030), .Z(n5493) );
  NANDN U5615 ( .A(n5493), .B(n19766), .Z(n5417) );
  NANDN U5616 ( .A(n5415), .B(n19767), .Z(n5416) );
  NAND U5617 ( .A(n5417), .B(n5416), .Z(n5472) );
  NAND U5618 ( .A(n19554), .B(n5418), .Z(n5420) );
  IV U5619 ( .A(a[74]), .Z(n6315) );
  XNOR U5620 ( .A(b[3]), .B(n6315), .Z(n5496) );
  NANDN U5621 ( .A(n19521), .B(n5496), .Z(n5419) );
  AND U5622 ( .A(n5420), .B(n5419), .Z(n5473) );
  XNOR U5623 ( .A(n5472), .B(n5473), .Z(n5474) );
  XOR U5624 ( .A(n5475), .B(n5474), .Z(n5500) );
  XOR U5625 ( .A(n5499), .B(n5500), .Z(n5501) );
  XNOR U5626 ( .A(n5502), .B(n5501), .Z(n5450) );
  NAND U5627 ( .A(n5422), .B(n5421), .Z(n5426) );
  NAND U5628 ( .A(n5424), .B(n5423), .Z(n5425) );
  NAND U5629 ( .A(n5426), .B(n5425), .Z(n5451) );
  XOR U5630 ( .A(n5450), .B(n5451), .Z(n5453) );
  XNOR U5631 ( .A(n5452), .B(n5453), .Z(n5511) );
  NANDN U5632 ( .A(n5428), .B(n5427), .Z(n5432) );
  NAND U5633 ( .A(n5430), .B(n5429), .Z(n5431) );
  NAND U5634 ( .A(n5432), .B(n5431), .Z(n5512) );
  XNOR U5635 ( .A(n5511), .B(n5512), .Z(n5513) );
  XOR U5636 ( .A(n5514), .B(n5513), .Z(n5444) );
  NANDN U5637 ( .A(n5434), .B(n5433), .Z(n5438) );
  NANDN U5638 ( .A(n5436), .B(n5435), .Z(n5437) );
  NAND U5639 ( .A(n5438), .B(n5437), .Z(n5445) );
  XNOR U5640 ( .A(n5444), .B(n5445), .Z(n5446) );
  XNOR U5641 ( .A(n5447), .B(n5446), .Z(n5517) );
  XNOR U5642 ( .A(n5517), .B(sreg[316]), .Z(n5519) );
  NAND U5643 ( .A(n5439), .B(sreg[315]), .Z(n5443) );
  OR U5644 ( .A(n5441), .B(n5440), .Z(n5442) );
  AND U5645 ( .A(n5443), .B(n5442), .Z(n5518) );
  XOR U5646 ( .A(n5519), .B(n5518), .Z(c[316]) );
  NANDN U5647 ( .A(n5445), .B(n5444), .Z(n5449) );
  NAND U5648 ( .A(n5447), .B(n5446), .Z(n5448) );
  NAND U5649 ( .A(n5449), .B(n5448), .Z(n5525) );
  NANDN U5650 ( .A(n5451), .B(n5450), .Z(n5455) );
  OR U5651 ( .A(n5453), .B(n5452), .Z(n5454) );
  NAND U5652 ( .A(n5455), .B(n5454), .Z(n5592) );
  XNOR U5653 ( .A(n20052), .B(n5771), .Z(n5546) );
  OR U5654 ( .A(n5546), .B(n20020), .Z(n5458) );
  NANDN U5655 ( .A(n5456), .B(n19960), .Z(n5457) );
  NAND U5656 ( .A(n5458), .B(n5457), .Z(n5543) );
  XNOR U5657 ( .A(n102), .B(n5459), .Z(n5550) );
  OR U5658 ( .A(n5550), .B(n20121), .Z(n5462) );
  NANDN U5659 ( .A(n5460), .B(n20122), .Z(n5461) );
  NAND U5660 ( .A(n5462), .B(n5461), .Z(n5540) );
  XNOR U5661 ( .A(n19975), .B(n5925), .Z(n5553) );
  NANDN U5662 ( .A(n5553), .B(n19883), .Z(n5465) );
  NANDN U5663 ( .A(n5463), .B(n19937), .Z(n5464) );
  AND U5664 ( .A(n5465), .B(n5464), .Z(n5541) );
  XNOR U5665 ( .A(n5540), .B(n5541), .Z(n5542) );
  XNOR U5666 ( .A(n5543), .B(n5542), .Z(n5583) );
  NANDN U5667 ( .A(n5467), .B(n5466), .Z(n5471) );
  NAND U5668 ( .A(n5469), .B(n5468), .Z(n5470) );
  NAND U5669 ( .A(n5471), .B(n5470), .Z(n5584) );
  XNOR U5670 ( .A(n5583), .B(n5584), .Z(n5585) );
  NANDN U5671 ( .A(n5473), .B(n5472), .Z(n5477) );
  NAND U5672 ( .A(n5475), .B(n5474), .Z(n5476) );
  AND U5673 ( .A(n5477), .B(n5476), .Z(n5586) );
  XNOR U5674 ( .A(n5585), .B(n5586), .Z(n5530) );
  NANDN U5675 ( .A(n5479), .B(n5478), .Z(n5483) );
  OR U5676 ( .A(n5481), .B(n5480), .Z(n5482) );
  NAND U5677 ( .A(n5483), .B(n5482), .Z(n5580) );
  NAND U5678 ( .A(b[0]), .B(a[77]), .Z(n5484) );
  XNOR U5679 ( .A(b[1]), .B(n5484), .Z(n5486) );
  NAND U5680 ( .A(a[76]), .B(n98), .Z(n5485) );
  AND U5681 ( .A(n5486), .B(n5485), .Z(n5556) );
  XNOR U5682 ( .A(n20154), .B(n5615), .Z(n5565) );
  OR U5683 ( .A(n5565), .B(n20057), .Z(n5489) );
  NANDN U5684 ( .A(n5487), .B(n20098), .Z(n5488) );
  AND U5685 ( .A(n5489), .B(n5488), .Z(n5557) );
  XOR U5686 ( .A(n5556), .B(n5557), .Z(n5559) );
  NAND U5687 ( .A(a[61]), .B(b[15]), .Z(n5558) );
  XOR U5688 ( .A(n5559), .B(n5558), .Z(n5577) );
  NAND U5689 ( .A(n19722), .B(n5490), .Z(n5492) );
  XNOR U5690 ( .A(b[5]), .B(n6237), .Z(n5568) );
  NANDN U5691 ( .A(n19640), .B(n5568), .Z(n5491) );
  NAND U5692 ( .A(n5492), .B(n5491), .Z(n5537) );
  XNOR U5693 ( .A(n19714), .B(n6108), .Z(n5571) );
  NANDN U5694 ( .A(n5571), .B(n19766), .Z(n5495) );
  NANDN U5695 ( .A(n5493), .B(n19767), .Z(n5494) );
  NAND U5696 ( .A(n5495), .B(n5494), .Z(n5534) );
  NAND U5697 ( .A(n19554), .B(n5496), .Z(n5498) );
  IV U5698 ( .A(a[75]), .Z(n6393) );
  XNOR U5699 ( .A(b[3]), .B(n6393), .Z(n5574) );
  NANDN U5700 ( .A(n19521), .B(n5574), .Z(n5497) );
  AND U5701 ( .A(n5498), .B(n5497), .Z(n5535) );
  XNOR U5702 ( .A(n5534), .B(n5535), .Z(n5536) );
  XOR U5703 ( .A(n5537), .B(n5536), .Z(n5578) );
  XOR U5704 ( .A(n5577), .B(n5578), .Z(n5579) );
  XNOR U5705 ( .A(n5580), .B(n5579), .Z(n5528) );
  NAND U5706 ( .A(n5500), .B(n5499), .Z(n5504) );
  NAND U5707 ( .A(n5502), .B(n5501), .Z(n5503) );
  NAND U5708 ( .A(n5504), .B(n5503), .Z(n5529) );
  XOR U5709 ( .A(n5528), .B(n5529), .Z(n5531) );
  XNOR U5710 ( .A(n5530), .B(n5531), .Z(n5589) );
  NANDN U5711 ( .A(n5506), .B(n5505), .Z(n5510) );
  NAND U5712 ( .A(n5508), .B(n5507), .Z(n5509) );
  NAND U5713 ( .A(n5510), .B(n5509), .Z(n5590) );
  XNOR U5714 ( .A(n5589), .B(n5590), .Z(n5591) );
  XOR U5715 ( .A(n5592), .B(n5591), .Z(n5522) );
  NANDN U5716 ( .A(n5512), .B(n5511), .Z(n5516) );
  NANDN U5717 ( .A(n5514), .B(n5513), .Z(n5515) );
  NAND U5718 ( .A(n5516), .B(n5515), .Z(n5523) );
  XNOR U5719 ( .A(n5522), .B(n5523), .Z(n5524) );
  XNOR U5720 ( .A(n5525), .B(n5524), .Z(n5595) );
  XNOR U5721 ( .A(n5595), .B(sreg[317]), .Z(n5597) );
  NAND U5722 ( .A(n5517), .B(sreg[316]), .Z(n5521) );
  OR U5723 ( .A(n5519), .B(n5518), .Z(n5520) );
  AND U5724 ( .A(n5521), .B(n5520), .Z(n5596) );
  XOR U5725 ( .A(n5597), .B(n5596), .Z(c[317]) );
  NANDN U5726 ( .A(n5523), .B(n5522), .Z(n5527) );
  NAND U5727 ( .A(n5525), .B(n5524), .Z(n5526) );
  NAND U5728 ( .A(n5527), .B(n5526), .Z(n5603) );
  NANDN U5729 ( .A(n5529), .B(n5528), .Z(n5533) );
  OR U5730 ( .A(n5531), .B(n5530), .Z(n5532) );
  NAND U5731 ( .A(n5533), .B(n5532), .Z(n5670) );
  NANDN U5732 ( .A(n5535), .B(n5534), .Z(n5539) );
  NAND U5733 ( .A(n5537), .B(n5536), .Z(n5538) );
  NAND U5734 ( .A(n5539), .B(n5538), .Z(n5664) );
  NANDN U5735 ( .A(n5541), .B(n5540), .Z(n5545) );
  NAND U5736 ( .A(n5543), .B(n5542), .Z(n5544) );
  NAND U5737 ( .A(n5545), .B(n5544), .Z(n5661) );
  XNOR U5738 ( .A(n20052), .B(n5874), .Z(n5612) );
  OR U5739 ( .A(n5612), .B(n20020), .Z(n5548) );
  NANDN U5740 ( .A(n5546), .B(n19960), .Z(n5547) );
  NAND U5741 ( .A(n5548), .B(n5547), .Z(n5625) );
  XNOR U5742 ( .A(n102), .B(n5549), .Z(n5616) );
  OR U5743 ( .A(n5616), .B(n20121), .Z(n5552) );
  NANDN U5744 ( .A(n5550), .B(n20122), .Z(n5551) );
  NAND U5745 ( .A(n5552), .B(n5551), .Z(n5622) );
  XNOR U5746 ( .A(n19975), .B(n6030), .Z(n5619) );
  NANDN U5747 ( .A(n5619), .B(n19883), .Z(n5555) );
  NANDN U5748 ( .A(n5553), .B(n19937), .Z(n5554) );
  AND U5749 ( .A(n5555), .B(n5554), .Z(n5623) );
  XNOR U5750 ( .A(n5622), .B(n5623), .Z(n5624) );
  XNOR U5751 ( .A(n5625), .B(n5624), .Z(n5662) );
  XNOR U5752 ( .A(n5661), .B(n5662), .Z(n5663) );
  XNOR U5753 ( .A(n5664), .B(n5663), .Z(n5609) );
  NANDN U5754 ( .A(n5557), .B(n5556), .Z(n5561) );
  OR U5755 ( .A(n5559), .B(n5558), .Z(n5560) );
  NAND U5756 ( .A(n5561), .B(n5560), .Z(n5658) );
  NAND U5757 ( .A(b[0]), .B(a[78]), .Z(n5562) );
  XNOR U5758 ( .A(b[1]), .B(n5562), .Z(n5564) );
  NAND U5759 ( .A(a[77]), .B(n98), .Z(n5563) );
  AND U5760 ( .A(n5564), .B(n5563), .Z(n5634) );
  XNOR U5761 ( .A(n20154), .B(n5693), .Z(n5643) );
  OR U5762 ( .A(n5643), .B(n20057), .Z(n5567) );
  NANDN U5763 ( .A(n5565), .B(n20098), .Z(n5566) );
  AND U5764 ( .A(n5567), .B(n5566), .Z(n5635) );
  XOR U5765 ( .A(n5634), .B(n5635), .Z(n5637) );
  NAND U5766 ( .A(a[62]), .B(b[15]), .Z(n5636) );
  XOR U5767 ( .A(n5637), .B(n5636), .Z(n5655) );
  NAND U5768 ( .A(n19722), .B(n5568), .Z(n5570) );
  XNOR U5769 ( .A(b[5]), .B(n6315), .Z(n5646) );
  NANDN U5770 ( .A(n19640), .B(n5646), .Z(n5569) );
  NAND U5771 ( .A(n5570), .B(n5569), .Z(n5631) );
  XNOR U5772 ( .A(n19714), .B(n6186), .Z(n5649) );
  NANDN U5773 ( .A(n5649), .B(n19766), .Z(n5573) );
  NANDN U5774 ( .A(n5571), .B(n19767), .Z(n5572) );
  NAND U5775 ( .A(n5573), .B(n5572), .Z(n5628) );
  NAND U5776 ( .A(n19554), .B(n5574), .Z(n5576) );
  IV U5777 ( .A(a[76]), .Z(n6471) );
  XNOR U5778 ( .A(b[3]), .B(n6471), .Z(n5652) );
  NANDN U5779 ( .A(n19521), .B(n5652), .Z(n5575) );
  AND U5780 ( .A(n5576), .B(n5575), .Z(n5629) );
  XNOR U5781 ( .A(n5628), .B(n5629), .Z(n5630) );
  XOR U5782 ( .A(n5631), .B(n5630), .Z(n5656) );
  XOR U5783 ( .A(n5655), .B(n5656), .Z(n5657) );
  XNOR U5784 ( .A(n5658), .B(n5657), .Z(n5606) );
  NAND U5785 ( .A(n5578), .B(n5577), .Z(n5582) );
  NAND U5786 ( .A(n5580), .B(n5579), .Z(n5581) );
  NAND U5787 ( .A(n5582), .B(n5581), .Z(n5607) );
  XNOR U5788 ( .A(n5606), .B(n5607), .Z(n5608) );
  XOR U5789 ( .A(n5609), .B(n5608), .Z(n5667) );
  NANDN U5790 ( .A(n5584), .B(n5583), .Z(n5588) );
  NAND U5791 ( .A(n5586), .B(n5585), .Z(n5587) );
  NAND U5792 ( .A(n5588), .B(n5587), .Z(n5668) );
  XOR U5793 ( .A(n5667), .B(n5668), .Z(n5669) );
  XOR U5794 ( .A(n5670), .B(n5669), .Z(n5600) );
  NANDN U5795 ( .A(n5590), .B(n5589), .Z(n5594) );
  NANDN U5796 ( .A(n5592), .B(n5591), .Z(n5593) );
  NAND U5797 ( .A(n5594), .B(n5593), .Z(n5601) );
  XNOR U5798 ( .A(n5600), .B(n5601), .Z(n5602) );
  XNOR U5799 ( .A(n5603), .B(n5602), .Z(n5673) );
  XNOR U5800 ( .A(n5673), .B(sreg[318]), .Z(n5675) );
  NAND U5801 ( .A(n5595), .B(sreg[317]), .Z(n5599) );
  OR U5802 ( .A(n5597), .B(n5596), .Z(n5598) );
  AND U5803 ( .A(n5599), .B(n5598), .Z(n5674) );
  XOR U5804 ( .A(n5675), .B(n5674), .Z(c[318]) );
  NANDN U5805 ( .A(n5601), .B(n5600), .Z(n5605) );
  NAND U5806 ( .A(n5603), .B(n5602), .Z(n5604) );
  NAND U5807 ( .A(n5605), .B(n5604), .Z(n5681) );
  NANDN U5808 ( .A(n5607), .B(n5606), .Z(n5611) );
  NAND U5809 ( .A(n5609), .B(n5608), .Z(n5610) );
  NAND U5810 ( .A(n5611), .B(n5610), .Z(n5748) );
  XNOR U5811 ( .A(n20052), .B(n5925), .Z(n5690) );
  OR U5812 ( .A(n5690), .B(n20020), .Z(n5614) );
  NANDN U5813 ( .A(n5612), .B(n19960), .Z(n5613) );
  NAND U5814 ( .A(n5614), .B(n5613), .Z(n5703) );
  XNOR U5815 ( .A(n102), .B(n5615), .Z(n5694) );
  OR U5816 ( .A(n5694), .B(n20121), .Z(n5618) );
  NANDN U5817 ( .A(n5616), .B(n20122), .Z(n5617) );
  NAND U5818 ( .A(n5618), .B(n5617), .Z(n5700) );
  XNOR U5819 ( .A(n19975), .B(n6108), .Z(n5697) );
  NANDN U5820 ( .A(n5697), .B(n19883), .Z(n5621) );
  NANDN U5821 ( .A(n5619), .B(n19937), .Z(n5620) );
  AND U5822 ( .A(n5621), .B(n5620), .Z(n5701) );
  XNOR U5823 ( .A(n5700), .B(n5701), .Z(n5702) );
  XNOR U5824 ( .A(n5703), .B(n5702), .Z(n5739) );
  NANDN U5825 ( .A(n5623), .B(n5622), .Z(n5627) );
  NAND U5826 ( .A(n5625), .B(n5624), .Z(n5626) );
  NAND U5827 ( .A(n5627), .B(n5626), .Z(n5740) );
  XNOR U5828 ( .A(n5739), .B(n5740), .Z(n5741) );
  NANDN U5829 ( .A(n5629), .B(n5628), .Z(n5633) );
  NAND U5830 ( .A(n5631), .B(n5630), .Z(n5632) );
  AND U5831 ( .A(n5633), .B(n5632), .Z(n5742) );
  XNOR U5832 ( .A(n5741), .B(n5742), .Z(n5686) );
  NANDN U5833 ( .A(n5635), .B(n5634), .Z(n5639) );
  OR U5834 ( .A(n5637), .B(n5636), .Z(n5638) );
  NAND U5835 ( .A(n5639), .B(n5638), .Z(n5736) );
  NAND U5836 ( .A(b[0]), .B(a[79]), .Z(n5640) );
  XNOR U5837 ( .A(b[1]), .B(n5640), .Z(n5642) );
  NAND U5838 ( .A(a[78]), .B(n98), .Z(n5641) );
  AND U5839 ( .A(n5642), .B(n5641), .Z(n5712) );
  XNOR U5840 ( .A(n20154), .B(n5771), .Z(n5718) );
  OR U5841 ( .A(n5718), .B(n20057), .Z(n5645) );
  NANDN U5842 ( .A(n5643), .B(n20098), .Z(n5644) );
  AND U5843 ( .A(n5645), .B(n5644), .Z(n5713) );
  XOR U5844 ( .A(n5712), .B(n5713), .Z(n5715) );
  NAND U5845 ( .A(a[63]), .B(b[15]), .Z(n5714) );
  XOR U5846 ( .A(n5715), .B(n5714), .Z(n5733) );
  NAND U5847 ( .A(n19722), .B(n5646), .Z(n5648) );
  XNOR U5848 ( .A(b[5]), .B(n6393), .Z(n5724) );
  NANDN U5849 ( .A(n19640), .B(n5724), .Z(n5647) );
  NAND U5850 ( .A(n5648), .B(n5647), .Z(n5709) );
  XNOR U5851 ( .A(n19714), .B(n6237), .Z(n5727) );
  NANDN U5852 ( .A(n5727), .B(n19766), .Z(n5651) );
  NANDN U5853 ( .A(n5649), .B(n19767), .Z(n5650) );
  NAND U5854 ( .A(n5651), .B(n5650), .Z(n5706) );
  NAND U5855 ( .A(n19554), .B(n5652), .Z(n5654) );
  IV U5856 ( .A(a[77]), .Z(n6549) );
  XNOR U5857 ( .A(b[3]), .B(n6549), .Z(n5730) );
  NANDN U5858 ( .A(n19521), .B(n5730), .Z(n5653) );
  AND U5859 ( .A(n5654), .B(n5653), .Z(n5707) );
  XNOR U5860 ( .A(n5706), .B(n5707), .Z(n5708) );
  XOR U5861 ( .A(n5709), .B(n5708), .Z(n5734) );
  XOR U5862 ( .A(n5733), .B(n5734), .Z(n5735) );
  XNOR U5863 ( .A(n5736), .B(n5735), .Z(n5684) );
  NAND U5864 ( .A(n5656), .B(n5655), .Z(n5660) );
  NAND U5865 ( .A(n5658), .B(n5657), .Z(n5659) );
  NAND U5866 ( .A(n5660), .B(n5659), .Z(n5685) );
  XOR U5867 ( .A(n5684), .B(n5685), .Z(n5687) );
  XNOR U5868 ( .A(n5686), .B(n5687), .Z(n5745) );
  NANDN U5869 ( .A(n5662), .B(n5661), .Z(n5666) );
  NAND U5870 ( .A(n5664), .B(n5663), .Z(n5665) );
  AND U5871 ( .A(n5666), .B(n5665), .Z(n5746) );
  XNOR U5872 ( .A(n5745), .B(n5746), .Z(n5747) );
  XOR U5873 ( .A(n5748), .B(n5747), .Z(n5678) );
  OR U5874 ( .A(n5668), .B(n5667), .Z(n5672) );
  NANDN U5875 ( .A(n5670), .B(n5669), .Z(n5671) );
  NAND U5876 ( .A(n5672), .B(n5671), .Z(n5679) );
  XNOR U5877 ( .A(n5678), .B(n5679), .Z(n5680) );
  XNOR U5878 ( .A(n5681), .B(n5680), .Z(n5751) );
  XNOR U5879 ( .A(n5751), .B(sreg[319]), .Z(n5753) );
  NAND U5880 ( .A(n5673), .B(sreg[318]), .Z(n5677) );
  OR U5881 ( .A(n5675), .B(n5674), .Z(n5676) );
  AND U5882 ( .A(n5677), .B(n5676), .Z(n5752) );
  XOR U5883 ( .A(n5753), .B(n5752), .Z(c[319]) );
  NANDN U5884 ( .A(n5679), .B(n5678), .Z(n5683) );
  NAND U5885 ( .A(n5681), .B(n5680), .Z(n5682) );
  NAND U5886 ( .A(n5683), .B(n5682), .Z(n5759) );
  NANDN U5887 ( .A(n5685), .B(n5684), .Z(n5689) );
  OR U5888 ( .A(n5687), .B(n5686), .Z(n5688) );
  NAND U5889 ( .A(n5689), .B(n5688), .Z(n5826) );
  XNOR U5890 ( .A(n20052), .B(n6030), .Z(n5768) );
  OR U5891 ( .A(n5768), .B(n20020), .Z(n5692) );
  NANDN U5892 ( .A(n5690), .B(n19960), .Z(n5691) );
  NAND U5893 ( .A(n5692), .B(n5691), .Z(n5781) );
  XNOR U5894 ( .A(n102), .B(n5693), .Z(n5772) );
  OR U5895 ( .A(n5772), .B(n20121), .Z(n5696) );
  NANDN U5896 ( .A(n5694), .B(n20122), .Z(n5695) );
  NAND U5897 ( .A(n5696), .B(n5695), .Z(n5778) );
  XNOR U5898 ( .A(n19975), .B(n6186), .Z(n5775) );
  NANDN U5899 ( .A(n5775), .B(n19883), .Z(n5699) );
  NANDN U5900 ( .A(n5697), .B(n19937), .Z(n5698) );
  AND U5901 ( .A(n5699), .B(n5698), .Z(n5779) );
  XNOR U5902 ( .A(n5778), .B(n5779), .Z(n5780) );
  XNOR U5903 ( .A(n5781), .B(n5780), .Z(n5817) );
  NANDN U5904 ( .A(n5701), .B(n5700), .Z(n5705) );
  NAND U5905 ( .A(n5703), .B(n5702), .Z(n5704) );
  NAND U5906 ( .A(n5705), .B(n5704), .Z(n5818) );
  XNOR U5907 ( .A(n5817), .B(n5818), .Z(n5819) );
  NANDN U5908 ( .A(n5707), .B(n5706), .Z(n5711) );
  NAND U5909 ( .A(n5709), .B(n5708), .Z(n5710) );
  AND U5910 ( .A(n5711), .B(n5710), .Z(n5820) );
  XNOR U5911 ( .A(n5819), .B(n5820), .Z(n5764) );
  NANDN U5912 ( .A(n5713), .B(n5712), .Z(n5717) );
  OR U5913 ( .A(n5715), .B(n5714), .Z(n5716) );
  NAND U5914 ( .A(n5717), .B(n5716), .Z(n5814) );
  XNOR U5915 ( .A(n20154), .B(n5874), .Z(n5796) );
  OR U5916 ( .A(n5796), .B(n20057), .Z(n5720) );
  NANDN U5917 ( .A(n5718), .B(n20098), .Z(n5719) );
  AND U5918 ( .A(n5720), .B(n5719), .Z(n5791) );
  NAND U5919 ( .A(b[0]), .B(a[80]), .Z(n5721) );
  XNOR U5920 ( .A(b[1]), .B(n5721), .Z(n5723) );
  NAND U5921 ( .A(a[79]), .B(n98), .Z(n5722) );
  AND U5922 ( .A(n5723), .B(n5722), .Z(n5790) );
  XOR U5923 ( .A(n5791), .B(n5790), .Z(n5793) );
  NAND U5924 ( .A(a[64]), .B(b[15]), .Z(n5792) );
  XOR U5925 ( .A(n5793), .B(n5792), .Z(n5811) );
  NAND U5926 ( .A(n19722), .B(n5724), .Z(n5726) );
  XNOR U5927 ( .A(b[5]), .B(n6471), .Z(n5802) );
  NANDN U5928 ( .A(n19640), .B(n5802), .Z(n5725) );
  NAND U5929 ( .A(n5726), .B(n5725), .Z(n5787) );
  XNOR U5930 ( .A(n19714), .B(n6315), .Z(n5805) );
  NANDN U5931 ( .A(n5805), .B(n19766), .Z(n5729) );
  NANDN U5932 ( .A(n5727), .B(n19767), .Z(n5728) );
  NAND U5933 ( .A(n5729), .B(n5728), .Z(n5784) );
  NAND U5934 ( .A(n19554), .B(n5730), .Z(n5732) );
  IV U5935 ( .A(a[78]), .Z(n6627) );
  XNOR U5936 ( .A(b[3]), .B(n6627), .Z(n5808) );
  NANDN U5937 ( .A(n19521), .B(n5808), .Z(n5731) );
  AND U5938 ( .A(n5732), .B(n5731), .Z(n5785) );
  XNOR U5939 ( .A(n5784), .B(n5785), .Z(n5786) );
  XOR U5940 ( .A(n5787), .B(n5786), .Z(n5812) );
  XOR U5941 ( .A(n5811), .B(n5812), .Z(n5813) );
  XNOR U5942 ( .A(n5814), .B(n5813), .Z(n5762) );
  NAND U5943 ( .A(n5734), .B(n5733), .Z(n5738) );
  NAND U5944 ( .A(n5736), .B(n5735), .Z(n5737) );
  NAND U5945 ( .A(n5738), .B(n5737), .Z(n5763) );
  XOR U5946 ( .A(n5762), .B(n5763), .Z(n5765) );
  XNOR U5947 ( .A(n5764), .B(n5765), .Z(n5823) );
  NANDN U5948 ( .A(n5740), .B(n5739), .Z(n5744) );
  NAND U5949 ( .A(n5742), .B(n5741), .Z(n5743) );
  NAND U5950 ( .A(n5744), .B(n5743), .Z(n5824) );
  XNOR U5951 ( .A(n5823), .B(n5824), .Z(n5825) );
  XOR U5952 ( .A(n5826), .B(n5825), .Z(n5756) );
  NANDN U5953 ( .A(n5746), .B(n5745), .Z(n5750) );
  NANDN U5954 ( .A(n5748), .B(n5747), .Z(n5749) );
  NAND U5955 ( .A(n5750), .B(n5749), .Z(n5757) );
  XNOR U5956 ( .A(n5756), .B(n5757), .Z(n5758) );
  XNOR U5957 ( .A(n5759), .B(n5758), .Z(n5829) );
  XNOR U5958 ( .A(n5829), .B(sreg[320]), .Z(n5831) );
  NAND U5959 ( .A(n5751), .B(sreg[319]), .Z(n5755) );
  OR U5960 ( .A(n5753), .B(n5752), .Z(n5754) );
  AND U5961 ( .A(n5755), .B(n5754), .Z(n5830) );
  XOR U5962 ( .A(n5831), .B(n5830), .Z(c[320]) );
  NANDN U5963 ( .A(n5757), .B(n5756), .Z(n5761) );
  NAND U5964 ( .A(n5759), .B(n5758), .Z(n5760) );
  NAND U5965 ( .A(n5761), .B(n5760), .Z(n5837) );
  NANDN U5966 ( .A(n5763), .B(n5762), .Z(n5767) );
  OR U5967 ( .A(n5765), .B(n5764), .Z(n5766) );
  NAND U5968 ( .A(n5767), .B(n5766), .Z(n5902) );
  XNOR U5969 ( .A(n20052), .B(n6108), .Z(n5871) );
  OR U5970 ( .A(n5871), .B(n20020), .Z(n5770) );
  NANDN U5971 ( .A(n5768), .B(n19960), .Z(n5769) );
  NAND U5972 ( .A(n5770), .B(n5769), .Z(n5884) );
  XNOR U5973 ( .A(n102), .B(n5771), .Z(n5875) );
  OR U5974 ( .A(n5875), .B(n20121), .Z(n5774) );
  NANDN U5975 ( .A(n5772), .B(n20122), .Z(n5773) );
  NAND U5976 ( .A(n5774), .B(n5773), .Z(n5881) );
  XNOR U5977 ( .A(n19975), .B(n6237), .Z(n5878) );
  NANDN U5978 ( .A(n5878), .B(n19883), .Z(n5777) );
  NANDN U5979 ( .A(n5775), .B(n19937), .Z(n5776) );
  AND U5980 ( .A(n5777), .B(n5776), .Z(n5882) );
  XNOR U5981 ( .A(n5881), .B(n5882), .Z(n5883) );
  XNOR U5982 ( .A(n5884), .B(n5883), .Z(n5893) );
  NANDN U5983 ( .A(n5779), .B(n5778), .Z(n5783) );
  NAND U5984 ( .A(n5781), .B(n5780), .Z(n5782) );
  NAND U5985 ( .A(n5783), .B(n5782), .Z(n5894) );
  XNOR U5986 ( .A(n5893), .B(n5894), .Z(n5895) );
  NANDN U5987 ( .A(n5785), .B(n5784), .Z(n5789) );
  NAND U5988 ( .A(n5787), .B(n5786), .Z(n5788) );
  AND U5989 ( .A(n5789), .B(n5788), .Z(n5896) );
  XNOR U5990 ( .A(n5895), .B(n5896), .Z(n5842) );
  NANDN U5991 ( .A(n5791), .B(n5790), .Z(n5795) );
  OR U5992 ( .A(n5793), .B(n5792), .Z(n5794) );
  NAND U5993 ( .A(n5795), .B(n5794), .Z(n5870) );
  XNOR U5994 ( .A(n20154), .B(n5925), .Z(n5855) );
  OR U5995 ( .A(n5855), .B(n20057), .Z(n5798) );
  NANDN U5996 ( .A(n5796), .B(n20098), .Z(n5797) );
  NAND U5997 ( .A(n5798), .B(n5797), .Z(n5846) );
  AND U5998 ( .A(a[81]), .B(b[0]), .Z(n5799) );
  XOR U5999 ( .A(b[1]), .B(n5799), .Z(n5801) );
  NAND U6000 ( .A(b[1]), .B(n98), .Z(n15156) );
  NANDN U6001 ( .A(n15156), .B(a[80]), .Z(n5800) );
  NAND U6002 ( .A(n5801), .B(n5800), .Z(n5847) );
  XNOR U6003 ( .A(n5846), .B(n5847), .Z(n5848) );
  NAND U6004 ( .A(a[65]), .B(b[15]), .Z(n5849) );
  XOR U6005 ( .A(n5848), .B(n5849), .Z(n5867) );
  NAND U6006 ( .A(n19722), .B(n5802), .Z(n5804) );
  XNOR U6007 ( .A(b[5]), .B(n6549), .Z(n5858) );
  NANDN U6008 ( .A(n19640), .B(n5858), .Z(n5803) );
  NAND U6009 ( .A(n5804), .B(n5803), .Z(n5890) );
  XNOR U6010 ( .A(n19714), .B(n6393), .Z(n5861) );
  NANDN U6011 ( .A(n5861), .B(n19766), .Z(n5807) );
  NANDN U6012 ( .A(n5805), .B(n19767), .Z(n5806) );
  NAND U6013 ( .A(n5807), .B(n5806), .Z(n5887) );
  NAND U6014 ( .A(n19554), .B(n5808), .Z(n5810) );
  IV U6015 ( .A(a[79]), .Z(n6705) );
  XNOR U6016 ( .A(b[3]), .B(n6705), .Z(n5864) );
  NANDN U6017 ( .A(n19521), .B(n5864), .Z(n5809) );
  AND U6018 ( .A(n5810), .B(n5809), .Z(n5888) );
  XNOR U6019 ( .A(n5887), .B(n5888), .Z(n5889) );
  XOR U6020 ( .A(n5890), .B(n5889), .Z(n5868) );
  XNOR U6021 ( .A(n5867), .B(n5868), .Z(n5869) );
  XNOR U6022 ( .A(n5870), .B(n5869), .Z(n5840) );
  NAND U6023 ( .A(n5812), .B(n5811), .Z(n5816) );
  NAND U6024 ( .A(n5814), .B(n5813), .Z(n5815) );
  NAND U6025 ( .A(n5816), .B(n5815), .Z(n5841) );
  XOR U6026 ( .A(n5840), .B(n5841), .Z(n5843) );
  XNOR U6027 ( .A(n5842), .B(n5843), .Z(n5899) );
  NANDN U6028 ( .A(n5818), .B(n5817), .Z(n5822) );
  NAND U6029 ( .A(n5820), .B(n5819), .Z(n5821) );
  NAND U6030 ( .A(n5822), .B(n5821), .Z(n5900) );
  XNOR U6031 ( .A(n5899), .B(n5900), .Z(n5901) );
  XOR U6032 ( .A(n5902), .B(n5901), .Z(n5834) );
  NANDN U6033 ( .A(n5824), .B(n5823), .Z(n5828) );
  NANDN U6034 ( .A(n5826), .B(n5825), .Z(n5827) );
  NAND U6035 ( .A(n5828), .B(n5827), .Z(n5835) );
  XNOR U6036 ( .A(n5834), .B(n5835), .Z(n5836) );
  XNOR U6037 ( .A(n5837), .B(n5836), .Z(n5905) );
  XNOR U6038 ( .A(n5905), .B(sreg[321]), .Z(n5907) );
  NAND U6039 ( .A(n5829), .B(sreg[320]), .Z(n5833) );
  OR U6040 ( .A(n5831), .B(n5830), .Z(n5832) );
  AND U6041 ( .A(n5833), .B(n5832), .Z(n5906) );
  XOR U6042 ( .A(n5907), .B(n5906), .Z(c[321]) );
  NANDN U6043 ( .A(n5835), .B(n5834), .Z(n5839) );
  NAND U6044 ( .A(n5837), .B(n5836), .Z(n5838) );
  NAND U6045 ( .A(n5839), .B(n5838), .Z(n5913) );
  NANDN U6046 ( .A(n5841), .B(n5840), .Z(n5845) );
  OR U6047 ( .A(n5843), .B(n5842), .Z(n5844) );
  NAND U6048 ( .A(n5845), .B(n5844), .Z(n5980) );
  NANDN U6049 ( .A(n5847), .B(n5846), .Z(n5851) );
  NANDN U6050 ( .A(n5849), .B(n5848), .Z(n5850) );
  NAND U6051 ( .A(n5851), .B(n5850), .Z(n5968) );
  NAND U6052 ( .A(b[0]), .B(a[82]), .Z(n5852) );
  XNOR U6053 ( .A(b[1]), .B(n5852), .Z(n5854) );
  NAND U6054 ( .A(a[81]), .B(n98), .Z(n5853) );
  AND U6055 ( .A(n5854), .B(n5853), .Z(n5944) );
  XNOR U6056 ( .A(n20154), .B(n6030), .Z(n5953) );
  OR U6057 ( .A(n5953), .B(n20057), .Z(n5857) );
  NANDN U6058 ( .A(n5855), .B(n20098), .Z(n5856) );
  AND U6059 ( .A(n5857), .B(n5856), .Z(n5945) );
  XOR U6060 ( .A(n5944), .B(n5945), .Z(n5947) );
  NAND U6061 ( .A(a[66]), .B(b[15]), .Z(n5946) );
  XOR U6062 ( .A(n5947), .B(n5946), .Z(n5965) );
  NAND U6063 ( .A(n19722), .B(n5858), .Z(n5860) );
  XNOR U6064 ( .A(b[5]), .B(n6627), .Z(n5956) );
  NANDN U6065 ( .A(n19640), .B(n5956), .Z(n5859) );
  NAND U6066 ( .A(n5860), .B(n5859), .Z(n5941) );
  XNOR U6067 ( .A(n19714), .B(n6471), .Z(n5959) );
  NANDN U6068 ( .A(n5959), .B(n19766), .Z(n5863) );
  NANDN U6069 ( .A(n5861), .B(n19767), .Z(n5862) );
  NAND U6070 ( .A(n5863), .B(n5862), .Z(n5938) );
  NAND U6071 ( .A(n19554), .B(n5864), .Z(n5866) );
  IV U6072 ( .A(a[80]), .Z(n6783) );
  XNOR U6073 ( .A(b[3]), .B(n6783), .Z(n5962) );
  NANDN U6074 ( .A(n19521), .B(n5962), .Z(n5865) );
  AND U6075 ( .A(n5866), .B(n5865), .Z(n5939) );
  XNOR U6076 ( .A(n5938), .B(n5939), .Z(n5940) );
  XOR U6077 ( .A(n5941), .B(n5940), .Z(n5966) );
  XOR U6078 ( .A(n5965), .B(n5966), .Z(n5967) );
  XNOR U6079 ( .A(n5968), .B(n5967), .Z(n5916) );
  XOR U6080 ( .A(n5916), .B(n5917), .Z(n5919) );
  XNOR U6081 ( .A(n20052), .B(n6186), .Z(n5922) );
  OR U6082 ( .A(n5922), .B(n20020), .Z(n5873) );
  NANDN U6083 ( .A(n5871), .B(n19960), .Z(n5872) );
  NAND U6084 ( .A(n5873), .B(n5872), .Z(n5935) );
  XNOR U6085 ( .A(n102), .B(n5874), .Z(n5926) );
  OR U6086 ( .A(n5926), .B(n20121), .Z(n5877) );
  NANDN U6087 ( .A(n5875), .B(n20122), .Z(n5876) );
  NAND U6088 ( .A(n5877), .B(n5876), .Z(n5932) );
  XNOR U6089 ( .A(n19975), .B(n6315), .Z(n5929) );
  NANDN U6090 ( .A(n5929), .B(n19883), .Z(n5880) );
  NANDN U6091 ( .A(n5878), .B(n19937), .Z(n5879) );
  AND U6092 ( .A(n5880), .B(n5879), .Z(n5933) );
  XNOR U6093 ( .A(n5932), .B(n5933), .Z(n5934) );
  XNOR U6094 ( .A(n5935), .B(n5934), .Z(n5971) );
  NANDN U6095 ( .A(n5882), .B(n5881), .Z(n5886) );
  NAND U6096 ( .A(n5884), .B(n5883), .Z(n5885) );
  NAND U6097 ( .A(n5886), .B(n5885), .Z(n5972) );
  XNOR U6098 ( .A(n5971), .B(n5972), .Z(n5973) );
  NANDN U6099 ( .A(n5888), .B(n5887), .Z(n5892) );
  NAND U6100 ( .A(n5890), .B(n5889), .Z(n5891) );
  AND U6101 ( .A(n5892), .B(n5891), .Z(n5974) );
  XNOR U6102 ( .A(n5973), .B(n5974), .Z(n5918) );
  XNOR U6103 ( .A(n5919), .B(n5918), .Z(n5977) );
  NANDN U6104 ( .A(n5894), .B(n5893), .Z(n5898) );
  NAND U6105 ( .A(n5896), .B(n5895), .Z(n5897) );
  NAND U6106 ( .A(n5898), .B(n5897), .Z(n5978) );
  XNOR U6107 ( .A(n5977), .B(n5978), .Z(n5979) );
  XOR U6108 ( .A(n5980), .B(n5979), .Z(n5910) );
  NANDN U6109 ( .A(n5900), .B(n5899), .Z(n5904) );
  NANDN U6110 ( .A(n5902), .B(n5901), .Z(n5903) );
  NAND U6111 ( .A(n5904), .B(n5903), .Z(n5911) );
  XNOR U6112 ( .A(n5910), .B(n5911), .Z(n5912) );
  XNOR U6113 ( .A(n5913), .B(n5912), .Z(n5983) );
  XNOR U6114 ( .A(n5983), .B(sreg[322]), .Z(n5985) );
  NAND U6115 ( .A(n5905), .B(sreg[321]), .Z(n5909) );
  OR U6116 ( .A(n5907), .B(n5906), .Z(n5908) );
  AND U6117 ( .A(n5909), .B(n5908), .Z(n5984) );
  XOR U6118 ( .A(n5985), .B(n5984), .Z(c[322]) );
  NANDN U6119 ( .A(n5911), .B(n5910), .Z(n5915) );
  NAND U6120 ( .A(n5913), .B(n5912), .Z(n5914) );
  NAND U6121 ( .A(n5915), .B(n5914), .Z(n5991) );
  NANDN U6122 ( .A(n5917), .B(n5916), .Z(n5921) );
  OR U6123 ( .A(n5919), .B(n5918), .Z(n5920) );
  NAND U6124 ( .A(n5921), .B(n5920), .Z(n6058) );
  XNOR U6125 ( .A(n20052), .B(n6237), .Z(n6027) );
  OR U6126 ( .A(n6027), .B(n20020), .Z(n5924) );
  NANDN U6127 ( .A(n5922), .B(n19960), .Z(n5923) );
  NAND U6128 ( .A(n5924), .B(n5923), .Z(n6040) );
  XNOR U6129 ( .A(n102), .B(n5925), .Z(n6031) );
  OR U6130 ( .A(n6031), .B(n20121), .Z(n5928) );
  NANDN U6131 ( .A(n5926), .B(n20122), .Z(n5927) );
  NAND U6132 ( .A(n5928), .B(n5927), .Z(n6037) );
  XNOR U6133 ( .A(n19975), .B(n6393), .Z(n6034) );
  NANDN U6134 ( .A(n6034), .B(n19883), .Z(n5931) );
  NANDN U6135 ( .A(n5929), .B(n19937), .Z(n5930) );
  AND U6136 ( .A(n5931), .B(n5930), .Z(n6038) );
  XNOR U6137 ( .A(n6037), .B(n6038), .Z(n6039) );
  XNOR U6138 ( .A(n6040), .B(n6039), .Z(n6049) );
  NANDN U6139 ( .A(n5933), .B(n5932), .Z(n5937) );
  NAND U6140 ( .A(n5935), .B(n5934), .Z(n5936) );
  NAND U6141 ( .A(n5937), .B(n5936), .Z(n6050) );
  XNOR U6142 ( .A(n6049), .B(n6050), .Z(n6051) );
  NANDN U6143 ( .A(n5939), .B(n5938), .Z(n5943) );
  NAND U6144 ( .A(n5941), .B(n5940), .Z(n5942) );
  AND U6145 ( .A(n5943), .B(n5942), .Z(n6052) );
  XNOR U6146 ( .A(n6051), .B(n6052), .Z(n5996) );
  NANDN U6147 ( .A(n5945), .B(n5944), .Z(n5949) );
  OR U6148 ( .A(n5947), .B(n5946), .Z(n5948) );
  NAND U6149 ( .A(n5949), .B(n5948), .Z(n6024) );
  NAND U6150 ( .A(b[0]), .B(a[83]), .Z(n5950) );
  XNOR U6151 ( .A(b[1]), .B(n5950), .Z(n5952) );
  NAND U6152 ( .A(a[82]), .B(n98), .Z(n5951) );
  AND U6153 ( .A(n5952), .B(n5951), .Z(n6000) );
  XNOR U6154 ( .A(n20154), .B(n6108), .Z(n6009) );
  OR U6155 ( .A(n6009), .B(n20057), .Z(n5955) );
  NANDN U6156 ( .A(n5953), .B(n20098), .Z(n5954) );
  AND U6157 ( .A(n5955), .B(n5954), .Z(n6001) );
  XOR U6158 ( .A(n6000), .B(n6001), .Z(n6003) );
  NAND U6159 ( .A(a[67]), .B(b[15]), .Z(n6002) );
  XOR U6160 ( .A(n6003), .B(n6002), .Z(n6021) );
  NAND U6161 ( .A(n19722), .B(n5956), .Z(n5958) );
  XNOR U6162 ( .A(b[5]), .B(n6705), .Z(n6012) );
  NANDN U6163 ( .A(n19640), .B(n6012), .Z(n5957) );
  NAND U6164 ( .A(n5958), .B(n5957), .Z(n6046) );
  XNOR U6165 ( .A(n19714), .B(n6549), .Z(n6015) );
  NANDN U6166 ( .A(n6015), .B(n19766), .Z(n5961) );
  NANDN U6167 ( .A(n5959), .B(n19767), .Z(n5960) );
  NAND U6168 ( .A(n5961), .B(n5960), .Z(n6043) );
  NAND U6169 ( .A(n19554), .B(n5962), .Z(n5964) );
  IV U6170 ( .A(a[81]), .Z(n6888) );
  XNOR U6171 ( .A(b[3]), .B(n6888), .Z(n6018) );
  NANDN U6172 ( .A(n19521), .B(n6018), .Z(n5963) );
  AND U6173 ( .A(n5964), .B(n5963), .Z(n6044) );
  XNOR U6174 ( .A(n6043), .B(n6044), .Z(n6045) );
  XOR U6175 ( .A(n6046), .B(n6045), .Z(n6022) );
  XOR U6176 ( .A(n6021), .B(n6022), .Z(n6023) );
  XNOR U6177 ( .A(n6024), .B(n6023), .Z(n5994) );
  NAND U6178 ( .A(n5966), .B(n5965), .Z(n5970) );
  NAND U6179 ( .A(n5968), .B(n5967), .Z(n5969) );
  NAND U6180 ( .A(n5970), .B(n5969), .Z(n5995) );
  XOR U6181 ( .A(n5994), .B(n5995), .Z(n5997) );
  XNOR U6182 ( .A(n5996), .B(n5997), .Z(n6055) );
  NANDN U6183 ( .A(n5972), .B(n5971), .Z(n5976) );
  NAND U6184 ( .A(n5974), .B(n5973), .Z(n5975) );
  NAND U6185 ( .A(n5976), .B(n5975), .Z(n6056) );
  XNOR U6186 ( .A(n6055), .B(n6056), .Z(n6057) );
  XOR U6187 ( .A(n6058), .B(n6057), .Z(n5988) );
  NANDN U6188 ( .A(n5978), .B(n5977), .Z(n5982) );
  NANDN U6189 ( .A(n5980), .B(n5979), .Z(n5981) );
  NAND U6190 ( .A(n5982), .B(n5981), .Z(n5989) );
  XNOR U6191 ( .A(n5988), .B(n5989), .Z(n5990) );
  XNOR U6192 ( .A(n5991), .B(n5990), .Z(n6061) );
  XNOR U6193 ( .A(n6061), .B(sreg[323]), .Z(n6063) );
  NAND U6194 ( .A(n5983), .B(sreg[322]), .Z(n5987) );
  OR U6195 ( .A(n5985), .B(n5984), .Z(n5986) );
  AND U6196 ( .A(n5987), .B(n5986), .Z(n6062) );
  XOR U6197 ( .A(n6063), .B(n6062), .Z(c[323]) );
  NANDN U6198 ( .A(n5989), .B(n5988), .Z(n5993) );
  NAND U6199 ( .A(n5991), .B(n5990), .Z(n5992) );
  NAND U6200 ( .A(n5993), .B(n5992), .Z(n6069) );
  NANDN U6201 ( .A(n5995), .B(n5994), .Z(n5999) );
  OR U6202 ( .A(n5997), .B(n5996), .Z(n5998) );
  NAND U6203 ( .A(n5999), .B(n5998), .Z(n6136) );
  NANDN U6204 ( .A(n6001), .B(n6000), .Z(n6005) );
  OR U6205 ( .A(n6003), .B(n6002), .Z(n6004) );
  NAND U6206 ( .A(n6005), .B(n6004), .Z(n6102) );
  NAND U6207 ( .A(b[0]), .B(a[84]), .Z(n6006) );
  XNOR U6208 ( .A(b[1]), .B(n6006), .Z(n6008) );
  NAND U6209 ( .A(a[83]), .B(n98), .Z(n6007) );
  AND U6210 ( .A(n6008), .B(n6007), .Z(n6078) );
  XNOR U6211 ( .A(n20154), .B(n6186), .Z(n6087) );
  OR U6212 ( .A(n6087), .B(n20057), .Z(n6011) );
  NANDN U6213 ( .A(n6009), .B(n20098), .Z(n6010) );
  AND U6214 ( .A(n6011), .B(n6010), .Z(n6079) );
  XOR U6215 ( .A(n6078), .B(n6079), .Z(n6081) );
  NAND U6216 ( .A(a[68]), .B(b[15]), .Z(n6080) );
  XOR U6217 ( .A(n6081), .B(n6080), .Z(n6099) );
  NAND U6218 ( .A(n19722), .B(n6012), .Z(n6014) );
  XNOR U6219 ( .A(b[5]), .B(n6783), .Z(n6090) );
  NANDN U6220 ( .A(n19640), .B(n6090), .Z(n6013) );
  NAND U6221 ( .A(n6014), .B(n6013), .Z(n6124) );
  XNOR U6222 ( .A(n19714), .B(n6627), .Z(n6093) );
  NANDN U6223 ( .A(n6093), .B(n19766), .Z(n6017) );
  NANDN U6224 ( .A(n6015), .B(n19767), .Z(n6016) );
  NAND U6225 ( .A(n6017), .B(n6016), .Z(n6121) );
  NAND U6226 ( .A(n19554), .B(n6018), .Z(n6020) );
  IV U6227 ( .A(a[82]), .Z(n6951) );
  XNOR U6228 ( .A(b[3]), .B(n6951), .Z(n6096) );
  NANDN U6229 ( .A(n19521), .B(n6096), .Z(n6019) );
  AND U6230 ( .A(n6020), .B(n6019), .Z(n6122) );
  XNOR U6231 ( .A(n6121), .B(n6122), .Z(n6123) );
  XOR U6232 ( .A(n6124), .B(n6123), .Z(n6100) );
  XOR U6233 ( .A(n6099), .B(n6100), .Z(n6101) );
  XNOR U6234 ( .A(n6102), .B(n6101), .Z(n6072) );
  NAND U6235 ( .A(n6022), .B(n6021), .Z(n6026) );
  NAND U6236 ( .A(n6024), .B(n6023), .Z(n6025) );
  NAND U6237 ( .A(n6026), .B(n6025), .Z(n6073) );
  XOR U6238 ( .A(n6072), .B(n6073), .Z(n6075) );
  XNOR U6239 ( .A(n20052), .B(n6315), .Z(n6105) );
  OR U6240 ( .A(n6105), .B(n20020), .Z(n6029) );
  NANDN U6241 ( .A(n6027), .B(n19960), .Z(n6028) );
  NAND U6242 ( .A(n6029), .B(n6028), .Z(n6118) );
  XNOR U6243 ( .A(n102), .B(n6030), .Z(n6109) );
  OR U6244 ( .A(n6109), .B(n20121), .Z(n6033) );
  NANDN U6245 ( .A(n6031), .B(n20122), .Z(n6032) );
  NAND U6246 ( .A(n6033), .B(n6032), .Z(n6115) );
  XNOR U6247 ( .A(n19975), .B(n6471), .Z(n6112) );
  NANDN U6248 ( .A(n6112), .B(n19883), .Z(n6036) );
  NANDN U6249 ( .A(n6034), .B(n19937), .Z(n6035) );
  AND U6250 ( .A(n6036), .B(n6035), .Z(n6116) );
  XNOR U6251 ( .A(n6115), .B(n6116), .Z(n6117) );
  XNOR U6252 ( .A(n6118), .B(n6117), .Z(n6127) );
  NANDN U6253 ( .A(n6038), .B(n6037), .Z(n6042) );
  NAND U6254 ( .A(n6040), .B(n6039), .Z(n6041) );
  NAND U6255 ( .A(n6042), .B(n6041), .Z(n6128) );
  XNOR U6256 ( .A(n6127), .B(n6128), .Z(n6129) );
  NANDN U6257 ( .A(n6044), .B(n6043), .Z(n6048) );
  NAND U6258 ( .A(n6046), .B(n6045), .Z(n6047) );
  AND U6259 ( .A(n6048), .B(n6047), .Z(n6130) );
  XNOR U6260 ( .A(n6129), .B(n6130), .Z(n6074) );
  XNOR U6261 ( .A(n6075), .B(n6074), .Z(n6133) );
  NANDN U6262 ( .A(n6050), .B(n6049), .Z(n6054) );
  NAND U6263 ( .A(n6052), .B(n6051), .Z(n6053) );
  NAND U6264 ( .A(n6054), .B(n6053), .Z(n6134) );
  XNOR U6265 ( .A(n6133), .B(n6134), .Z(n6135) );
  XOR U6266 ( .A(n6136), .B(n6135), .Z(n6066) );
  NANDN U6267 ( .A(n6056), .B(n6055), .Z(n6060) );
  NANDN U6268 ( .A(n6058), .B(n6057), .Z(n6059) );
  NAND U6269 ( .A(n6060), .B(n6059), .Z(n6067) );
  XNOR U6270 ( .A(n6066), .B(n6067), .Z(n6068) );
  XNOR U6271 ( .A(n6069), .B(n6068), .Z(n6139) );
  XNOR U6272 ( .A(n6139), .B(sreg[324]), .Z(n6141) );
  NAND U6273 ( .A(n6061), .B(sreg[323]), .Z(n6065) );
  OR U6274 ( .A(n6063), .B(n6062), .Z(n6064) );
  AND U6275 ( .A(n6065), .B(n6064), .Z(n6140) );
  XOR U6276 ( .A(n6141), .B(n6140), .Z(c[324]) );
  NANDN U6277 ( .A(n6067), .B(n6066), .Z(n6071) );
  NAND U6278 ( .A(n6069), .B(n6068), .Z(n6070) );
  NAND U6279 ( .A(n6071), .B(n6070), .Z(n6147) );
  NANDN U6280 ( .A(n6073), .B(n6072), .Z(n6077) );
  OR U6281 ( .A(n6075), .B(n6074), .Z(n6076) );
  NAND U6282 ( .A(n6077), .B(n6076), .Z(n6214) );
  NANDN U6283 ( .A(n6079), .B(n6078), .Z(n6083) );
  OR U6284 ( .A(n6081), .B(n6080), .Z(n6082) );
  NAND U6285 ( .A(n6083), .B(n6082), .Z(n6180) );
  NAND U6286 ( .A(b[0]), .B(a[85]), .Z(n6084) );
  XNOR U6287 ( .A(b[1]), .B(n6084), .Z(n6086) );
  NAND U6288 ( .A(a[84]), .B(n98), .Z(n6085) );
  AND U6289 ( .A(n6086), .B(n6085), .Z(n6156) );
  XNOR U6290 ( .A(n20154), .B(n6237), .Z(n6165) );
  OR U6291 ( .A(n6165), .B(n20057), .Z(n6089) );
  NANDN U6292 ( .A(n6087), .B(n20098), .Z(n6088) );
  AND U6293 ( .A(n6089), .B(n6088), .Z(n6157) );
  XOR U6294 ( .A(n6156), .B(n6157), .Z(n6159) );
  NAND U6295 ( .A(a[69]), .B(b[15]), .Z(n6158) );
  XOR U6296 ( .A(n6159), .B(n6158), .Z(n6177) );
  NAND U6297 ( .A(n19722), .B(n6090), .Z(n6092) );
  XNOR U6298 ( .A(b[5]), .B(n6888), .Z(n6168) );
  NANDN U6299 ( .A(n19640), .B(n6168), .Z(n6091) );
  NAND U6300 ( .A(n6092), .B(n6091), .Z(n6202) );
  XNOR U6301 ( .A(n19714), .B(n6705), .Z(n6171) );
  NANDN U6302 ( .A(n6171), .B(n19766), .Z(n6095) );
  NANDN U6303 ( .A(n6093), .B(n19767), .Z(n6094) );
  NAND U6304 ( .A(n6095), .B(n6094), .Z(n6199) );
  NAND U6305 ( .A(n19554), .B(n6096), .Z(n6098) );
  IV U6306 ( .A(a[83]), .Z(n7044) );
  XNOR U6307 ( .A(b[3]), .B(n7044), .Z(n6174) );
  NANDN U6308 ( .A(n19521), .B(n6174), .Z(n6097) );
  AND U6309 ( .A(n6098), .B(n6097), .Z(n6200) );
  XNOR U6310 ( .A(n6199), .B(n6200), .Z(n6201) );
  XOR U6311 ( .A(n6202), .B(n6201), .Z(n6178) );
  XOR U6312 ( .A(n6177), .B(n6178), .Z(n6179) );
  XNOR U6313 ( .A(n6180), .B(n6179), .Z(n6150) );
  NAND U6314 ( .A(n6100), .B(n6099), .Z(n6104) );
  NAND U6315 ( .A(n6102), .B(n6101), .Z(n6103) );
  NAND U6316 ( .A(n6104), .B(n6103), .Z(n6151) );
  XOR U6317 ( .A(n6150), .B(n6151), .Z(n6153) );
  XNOR U6318 ( .A(n20052), .B(n6393), .Z(n6183) );
  OR U6319 ( .A(n6183), .B(n20020), .Z(n6107) );
  NANDN U6320 ( .A(n6105), .B(n19960), .Z(n6106) );
  NAND U6321 ( .A(n6107), .B(n6106), .Z(n6196) );
  XNOR U6322 ( .A(n102), .B(n6108), .Z(n6187) );
  OR U6323 ( .A(n6187), .B(n20121), .Z(n6111) );
  NANDN U6324 ( .A(n6109), .B(n20122), .Z(n6110) );
  NAND U6325 ( .A(n6111), .B(n6110), .Z(n6193) );
  XNOR U6326 ( .A(n19975), .B(n6549), .Z(n6190) );
  NANDN U6327 ( .A(n6190), .B(n19883), .Z(n6114) );
  NANDN U6328 ( .A(n6112), .B(n19937), .Z(n6113) );
  AND U6329 ( .A(n6114), .B(n6113), .Z(n6194) );
  XNOR U6330 ( .A(n6193), .B(n6194), .Z(n6195) );
  XNOR U6331 ( .A(n6196), .B(n6195), .Z(n6205) );
  NANDN U6332 ( .A(n6116), .B(n6115), .Z(n6120) );
  NAND U6333 ( .A(n6118), .B(n6117), .Z(n6119) );
  NAND U6334 ( .A(n6120), .B(n6119), .Z(n6206) );
  XNOR U6335 ( .A(n6205), .B(n6206), .Z(n6207) );
  NANDN U6336 ( .A(n6122), .B(n6121), .Z(n6126) );
  NAND U6337 ( .A(n6124), .B(n6123), .Z(n6125) );
  AND U6338 ( .A(n6126), .B(n6125), .Z(n6208) );
  XNOR U6339 ( .A(n6207), .B(n6208), .Z(n6152) );
  XNOR U6340 ( .A(n6153), .B(n6152), .Z(n6211) );
  NANDN U6341 ( .A(n6128), .B(n6127), .Z(n6132) );
  NAND U6342 ( .A(n6130), .B(n6129), .Z(n6131) );
  NAND U6343 ( .A(n6132), .B(n6131), .Z(n6212) );
  XNOR U6344 ( .A(n6211), .B(n6212), .Z(n6213) );
  XOR U6345 ( .A(n6214), .B(n6213), .Z(n6144) );
  NANDN U6346 ( .A(n6134), .B(n6133), .Z(n6138) );
  NANDN U6347 ( .A(n6136), .B(n6135), .Z(n6137) );
  NAND U6348 ( .A(n6138), .B(n6137), .Z(n6145) );
  XNOR U6349 ( .A(n6144), .B(n6145), .Z(n6146) );
  XNOR U6350 ( .A(n6147), .B(n6146), .Z(n6217) );
  XNOR U6351 ( .A(n6217), .B(sreg[325]), .Z(n6219) );
  NAND U6352 ( .A(n6139), .B(sreg[324]), .Z(n6143) );
  OR U6353 ( .A(n6141), .B(n6140), .Z(n6142) );
  AND U6354 ( .A(n6143), .B(n6142), .Z(n6218) );
  XOR U6355 ( .A(n6219), .B(n6218), .Z(c[325]) );
  NANDN U6356 ( .A(n6145), .B(n6144), .Z(n6149) );
  NAND U6357 ( .A(n6147), .B(n6146), .Z(n6148) );
  NAND U6358 ( .A(n6149), .B(n6148), .Z(n6225) );
  NANDN U6359 ( .A(n6151), .B(n6150), .Z(n6155) );
  OR U6360 ( .A(n6153), .B(n6152), .Z(n6154) );
  NAND U6361 ( .A(n6155), .B(n6154), .Z(n6292) );
  NANDN U6362 ( .A(n6157), .B(n6156), .Z(n6161) );
  OR U6363 ( .A(n6159), .B(n6158), .Z(n6160) );
  NAND U6364 ( .A(n6161), .B(n6160), .Z(n6280) );
  NAND U6365 ( .A(b[0]), .B(a[86]), .Z(n6162) );
  XNOR U6366 ( .A(b[1]), .B(n6162), .Z(n6164) );
  NAND U6367 ( .A(a[85]), .B(n98), .Z(n6163) );
  AND U6368 ( .A(n6164), .B(n6163), .Z(n6256) );
  XNOR U6369 ( .A(n20154), .B(n6315), .Z(n6265) );
  OR U6370 ( .A(n6265), .B(n20057), .Z(n6167) );
  NANDN U6371 ( .A(n6165), .B(n20098), .Z(n6166) );
  AND U6372 ( .A(n6167), .B(n6166), .Z(n6257) );
  XOR U6373 ( .A(n6256), .B(n6257), .Z(n6259) );
  NAND U6374 ( .A(a[70]), .B(b[15]), .Z(n6258) );
  XOR U6375 ( .A(n6259), .B(n6258), .Z(n6277) );
  NAND U6376 ( .A(n19722), .B(n6168), .Z(n6170) );
  XNOR U6377 ( .A(b[5]), .B(n6951), .Z(n6268) );
  NANDN U6378 ( .A(n19640), .B(n6268), .Z(n6169) );
  NAND U6379 ( .A(n6170), .B(n6169), .Z(n6253) );
  XNOR U6380 ( .A(n19714), .B(n6783), .Z(n6271) );
  NANDN U6381 ( .A(n6271), .B(n19766), .Z(n6173) );
  NANDN U6382 ( .A(n6171), .B(n19767), .Z(n6172) );
  NAND U6383 ( .A(n6173), .B(n6172), .Z(n6250) );
  NAND U6384 ( .A(n19554), .B(n6174), .Z(n6176) );
  IV U6385 ( .A(a[84]), .Z(n7095) );
  XNOR U6386 ( .A(b[3]), .B(n7095), .Z(n6274) );
  NANDN U6387 ( .A(n19521), .B(n6274), .Z(n6175) );
  AND U6388 ( .A(n6176), .B(n6175), .Z(n6251) );
  XNOR U6389 ( .A(n6250), .B(n6251), .Z(n6252) );
  XOR U6390 ( .A(n6253), .B(n6252), .Z(n6278) );
  XOR U6391 ( .A(n6277), .B(n6278), .Z(n6279) );
  XNOR U6392 ( .A(n6280), .B(n6279), .Z(n6228) );
  NAND U6393 ( .A(n6178), .B(n6177), .Z(n6182) );
  NAND U6394 ( .A(n6180), .B(n6179), .Z(n6181) );
  NAND U6395 ( .A(n6182), .B(n6181), .Z(n6229) );
  XOR U6396 ( .A(n6228), .B(n6229), .Z(n6231) );
  XNOR U6397 ( .A(n20052), .B(n6471), .Z(n6234) );
  OR U6398 ( .A(n6234), .B(n20020), .Z(n6185) );
  NANDN U6399 ( .A(n6183), .B(n19960), .Z(n6184) );
  NAND U6400 ( .A(n6185), .B(n6184), .Z(n6247) );
  XNOR U6401 ( .A(n102), .B(n6186), .Z(n6238) );
  OR U6402 ( .A(n6238), .B(n20121), .Z(n6189) );
  NANDN U6403 ( .A(n6187), .B(n20122), .Z(n6188) );
  NAND U6404 ( .A(n6189), .B(n6188), .Z(n6244) );
  XNOR U6405 ( .A(n19975), .B(n6627), .Z(n6241) );
  NANDN U6406 ( .A(n6241), .B(n19883), .Z(n6192) );
  NANDN U6407 ( .A(n6190), .B(n19937), .Z(n6191) );
  AND U6408 ( .A(n6192), .B(n6191), .Z(n6245) );
  XNOR U6409 ( .A(n6244), .B(n6245), .Z(n6246) );
  XNOR U6410 ( .A(n6247), .B(n6246), .Z(n6283) );
  NANDN U6411 ( .A(n6194), .B(n6193), .Z(n6198) );
  NAND U6412 ( .A(n6196), .B(n6195), .Z(n6197) );
  NAND U6413 ( .A(n6198), .B(n6197), .Z(n6284) );
  XNOR U6414 ( .A(n6283), .B(n6284), .Z(n6285) );
  NANDN U6415 ( .A(n6200), .B(n6199), .Z(n6204) );
  NAND U6416 ( .A(n6202), .B(n6201), .Z(n6203) );
  AND U6417 ( .A(n6204), .B(n6203), .Z(n6286) );
  XNOR U6418 ( .A(n6285), .B(n6286), .Z(n6230) );
  XNOR U6419 ( .A(n6231), .B(n6230), .Z(n6289) );
  NANDN U6420 ( .A(n6206), .B(n6205), .Z(n6210) );
  NAND U6421 ( .A(n6208), .B(n6207), .Z(n6209) );
  NAND U6422 ( .A(n6210), .B(n6209), .Z(n6290) );
  XNOR U6423 ( .A(n6289), .B(n6290), .Z(n6291) );
  XOR U6424 ( .A(n6292), .B(n6291), .Z(n6222) );
  NANDN U6425 ( .A(n6212), .B(n6211), .Z(n6216) );
  NANDN U6426 ( .A(n6214), .B(n6213), .Z(n6215) );
  NAND U6427 ( .A(n6216), .B(n6215), .Z(n6223) );
  XNOR U6428 ( .A(n6222), .B(n6223), .Z(n6224) );
  XNOR U6429 ( .A(n6225), .B(n6224), .Z(n6295) );
  XNOR U6430 ( .A(n6295), .B(sreg[326]), .Z(n6297) );
  NAND U6431 ( .A(n6217), .B(sreg[325]), .Z(n6221) );
  OR U6432 ( .A(n6219), .B(n6218), .Z(n6220) );
  AND U6433 ( .A(n6221), .B(n6220), .Z(n6296) );
  XOR U6434 ( .A(n6297), .B(n6296), .Z(c[326]) );
  NANDN U6435 ( .A(n6223), .B(n6222), .Z(n6227) );
  NAND U6436 ( .A(n6225), .B(n6224), .Z(n6226) );
  NAND U6437 ( .A(n6227), .B(n6226), .Z(n6303) );
  NANDN U6438 ( .A(n6229), .B(n6228), .Z(n6233) );
  OR U6439 ( .A(n6231), .B(n6230), .Z(n6232) );
  NAND U6440 ( .A(n6233), .B(n6232), .Z(n6370) );
  XNOR U6441 ( .A(n20052), .B(n6549), .Z(n6312) );
  OR U6442 ( .A(n6312), .B(n20020), .Z(n6236) );
  NANDN U6443 ( .A(n6234), .B(n19960), .Z(n6235) );
  NAND U6444 ( .A(n6236), .B(n6235), .Z(n6325) );
  XNOR U6445 ( .A(n102), .B(n6237), .Z(n6316) );
  OR U6446 ( .A(n6316), .B(n20121), .Z(n6240) );
  NANDN U6447 ( .A(n6238), .B(n20122), .Z(n6239) );
  NAND U6448 ( .A(n6240), .B(n6239), .Z(n6322) );
  XNOR U6449 ( .A(n19975), .B(n6705), .Z(n6319) );
  NANDN U6450 ( .A(n6319), .B(n19883), .Z(n6243) );
  NANDN U6451 ( .A(n6241), .B(n19937), .Z(n6242) );
  AND U6452 ( .A(n6243), .B(n6242), .Z(n6323) );
  XNOR U6453 ( .A(n6322), .B(n6323), .Z(n6324) );
  XNOR U6454 ( .A(n6325), .B(n6324), .Z(n6361) );
  NANDN U6455 ( .A(n6245), .B(n6244), .Z(n6249) );
  NAND U6456 ( .A(n6247), .B(n6246), .Z(n6248) );
  NAND U6457 ( .A(n6249), .B(n6248), .Z(n6362) );
  XNOR U6458 ( .A(n6361), .B(n6362), .Z(n6363) );
  NANDN U6459 ( .A(n6251), .B(n6250), .Z(n6255) );
  NAND U6460 ( .A(n6253), .B(n6252), .Z(n6254) );
  AND U6461 ( .A(n6255), .B(n6254), .Z(n6364) );
  XNOR U6462 ( .A(n6363), .B(n6364), .Z(n6308) );
  NANDN U6463 ( .A(n6257), .B(n6256), .Z(n6261) );
  OR U6464 ( .A(n6259), .B(n6258), .Z(n6260) );
  NAND U6465 ( .A(n6261), .B(n6260), .Z(n6358) );
  NAND U6466 ( .A(b[0]), .B(a[87]), .Z(n6262) );
  XNOR U6467 ( .A(b[1]), .B(n6262), .Z(n6264) );
  NAND U6468 ( .A(a[86]), .B(n98), .Z(n6263) );
  AND U6469 ( .A(n6264), .B(n6263), .Z(n6334) );
  XNOR U6470 ( .A(n20154), .B(n6393), .Z(n6343) );
  OR U6471 ( .A(n6343), .B(n20057), .Z(n6267) );
  NANDN U6472 ( .A(n6265), .B(n20098), .Z(n6266) );
  AND U6473 ( .A(n6267), .B(n6266), .Z(n6335) );
  XOR U6474 ( .A(n6334), .B(n6335), .Z(n6337) );
  NAND U6475 ( .A(a[71]), .B(b[15]), .Z(n6336) );
  XOR U6476 ( .A(n6337), .B(n6336), .Z(n6355) );
  NAND U6477 ( .A(n19722), .B(n6268), .Z(n6270) );
  XNOR U6478 ( .A(b[5]), .B(n7044), .Z(n6346) );
  NANDN U6479 ( .A(n19640), .B(n6346), .Z(n6269) );
  NAND U6480 ( .A(n6270), .B(n6269), .Z(n6331) );
  XNOR U6481 ( .A(n19714), .B(n6888), .Z(n6349) );
  NANDN U6482 ( .A(n6349), .B(n19766), .Z(n6273) );
  NANDN U6483 ( .A(n6271), .B(n19767), .Z(n6272) );
  NAND U6484 ( .A(n6273), .B(n6272), .Z(n6328) );
  NAND U6485 ( .A(n19554), .B(n6274), .Z(n6276) );
  IV U6486 ( .A(a[85]), .Z(n7173) );
  XNOR U6487 ( .A(b[3]), .B(n7173), .Z(n6352) );
  NANDN U6488 ( .A(n19521), .B(n6352), .Z(n6275) );
  AND U6489 ( .A(n6276), .B(n6275), .Z(n6329) );
  XNOR U6490 ( .A(n6328), .B(n6329), .Z(n6330) );
  XOR U6491 ( .A(n6331), .B(n6330), .Z(n6356) );
  XOR U6492 ( .A(n6355), .B(n6356), .Z(n6357) );
  XNOR U6493 ( .A(n6358), .B(n6357), .Z(n6306) );
  NAND U6494 ( .A(n6278), .B(n6277), .Z(n6282) );
  NAND U6495 ( .A(n6280), .B(n6279), .Z(n6281) );
  NAND U6496 ( .A(n6282), .B(n6281), .Z(n6307) );
  XOR U6497 ( .A(n6306), .B(n6307), .Z(n6309) );
  XNOR U6498 ( .A(n6308), .B(n6309), .Z(n6367) );
  NANDN U6499 ( .A(n6284), .B(n6283), .Z(n6288) );
  NAND U6500 ( .A(n6286), .B(n6285), .Z(n6287) );
  NAND U6501 ( .A(n6288), .B(n6287), .Z(n6368) );
  XNOR U6502 ( .A(n6367), .B(n6368), .Z(n6369) );
  XOR U6503 ( .A(n6370), .B(n6369), .Z(n6300) );
  NANDN U6504 ( .A(n6290), .B(n6289), .Z(n6294) );
  NANDN U6505 ( .A(n6292), .B(n6291), .Z(n6293) );
  NAND U6506 ( .A(n6294), .B(n6293), .Z(n6301) );
  XNOR U6507 ( .A(n6300), .B(n6301), .Z(n6302) );
  XNOR U6508 ( .A(n6303), .B(n6302), .Z(n6373) );
  XNOR U6509 ( .A(n6373), .B(sreg[327]), .Z(n6375) );
  NAND U6510 ( .A(n6295), .B(sreg[326]), .Z(n6299) );
  OR U6511 ( .A(n6297), .B(n6296), .Z(n6298) );
  AND U6512 ( .A(n6299), .B(n6298), .Z(n6374) );
  XOR U6513 ( .A(n6375), .B(n6374), .Z(c[327]) );
  NANDN U6514 ( .A(n6301), .B(n6300), .Z(n6305) );
  NAND U6515 ( .A(n6303), .B(n6302), .Z(n6304) );
  NAND U6516 ( .A(n6305), .B(n6304), .Z(n6381) );
  NANDN U6517 ( .A(n6307), .B(n6306), .Z(n6311) );
  OR U6518 ( .A(n6309), .B(n6308), .Z(n6310) );
  NAND U6519 ( .A(n6311), .B(n6310), .Z(n6448) );
  XNOR U6520 ( .A(n20052), .B(n6627), .Z(n6390) );
  OR U6521 ( .A(n6390), .B(n20020), .Z(n6314) );
  NANDN U6522 ( .A(n6312), .B(n19960), .Z(n6313) );
  NAND U6523 ( .A(n6314), .B(n6313), .Z(n6403) );
  XNOR U6524 ( .A(n102), .B(n6315), .Z(n6394) );
  OR U6525 ( .A(n6394), .B(n20121), .Z(n6318) );
  NANDN U6526 ( .A(n6316), .B(n20122), .Z(n6317) );
  NAND U6527 ( .A(n6318), .B(n6317), .Z(n6400) );
  XNOR U6528 ( .A(n19975), .B(n6783), .Z(n6397) );
  NANDN U6529 ( .A(n6397), .B(n19883), .Z(n6321) );
  NANDN U6530 ( .A(n6319), .B(n19937), .Z(n6320) );
  AND U6531 ( .A(n6321), .B(n6320), .Z(n6401) );
  XNOR U6532 ( .A(n6400), .B(n6401), .Z(n6402) );
  XNOR U6533 ( .A(n6403), .B(n6402), .Z(n6439) );
  NANDN U6534 ( .A(n6323), .B(n6322), .Z(n6327) );
  NAND U6535 ( .A(n6325), .B(n6324), .Z(n6326) );
  NAND U6536 ( .A(n6327), .B(n6326), .Z(n6440) );
  XNOR U6537 ( .A(n6439), .B(n6440), .Z(n6441) );
  NANDN U6538 ( .A(n6329), .B(n6328), .Z(n6333) );
  NAND U6539 ( .A(n6331), .B(n6330), .Z(n6332) );
  AND U6540 ( .A(n6333), .B(n6332), .Z(n6442) );
  XNOR U6541 ( .A(n6441), .B(n6442), .Z(n6386) );
  NANDN U6542 ( .A(n6335), .B(n6334), .Z(n6339) );
  OR U6543 ( .A(n6337), .B(n6336), .Z(n6338) );
  NAND U6544 ( .A(n6339), .B(n6338), .Z(n6436) );
  NAND U6545 ( .A(b[0]), .B(a[88]), .Z(n6340) );
  XNOR U6546 ( .A(b[1]), .B(n6340), .Z(n6342) );
  NAND U6547 ( .A(a[87]), .B(n98), .Z(n6341) );
  AND U6548 ( .A(n6342), .B(n6341), .Z(n6412) );
  XNOR U6549 ( .A(n20154), .B(n6471), .Z(n6421) );
  OR U6550 ( .A(n6421), .B(n20057), .Z(n6345) );
  NANDN U6551 ( .A(n6343), .B(n20098), .Z(n6344) );
  AND U6552 ( .A(n6345), .B(n6344), .Z(n6413) );
  XOR U6553 ( .A(n6412), .B(n6413), .Z(n6415) );
  NAND U6554 ( .A(a[72]), .B(b[15]), .Z(n6414) );
  XOR U6555 ( .A(n6415), .B(n6414), .Z(n6433) );
  NAND U6556 ( .A(n19722), .B(n6346), .Z(n6348) );
  XNOR U6557 ( .A(b[5]), .B(n7095), .Z(n6424) );
  NANDN U6558 ( .A(n19640), .B(n6424), .Z(n6347) );
  NAND U6559 ( .A(n6348), .B(n6347), .Z(n6409) );
  XNOR U6560 ( .A(n19714), .B(n6951), .Z(n6427) );
  NANDN U6561 ( .A(n6427), .B(n19766), .Z(n6351) );
  NANDN U6562 ( .A(n6349), .B(n19767), .Z(n6350) );
  NAND U6563 ( .A(n6351), .B(n6350), .Z(n6406) );
  NAND U6564 ( .A(n19554), .B(n6352), .Z(n6354) );
  IV U6565 ( .A(a[86]), .Z(n7251) );
  XNOR U6566 ( .A(b[3]), .B(n7251), .Z(n6430) );
  NANDN U6567 ( .A(n19521), .B(n6430), .Z(n6353) );
  AND U6568 ( .A(n6354), .B(n6353), .Z(n6407) );
  XNOR U6569 ( .A(n6406), .B(n6407), .Z(n6408) );
  XOR U6570 ( .A(n6409), .B(n6408), .Z(n6434) );
  XOR U6571 ( .A(n6433), .B(n6434), .Z(n6435) );
  XNOR U6572 ( .A(n6436), .B(n6435), .Z(n6384) );
  NAND U6573 ( .A(n6356), .B(n6355), .Z(n6360) );
  NAND U6574 ( .A(n6358), .B(n6357), .Z(n6359) );
  NAND U6575 ( .A(n6360), .B(n6359), .Z(n6385) );
  XOR U6576 ( .A(n6384), .B(n6385), .Z(n6387) );
  XNOR U6577 ( .A(n6386), .B(n6387), .Z(n6445) );
  NANDN U6578 ( .A(n6362), .B(n6361), .Z(n6366) );
  NAND U6579 ( .A(n6364), .B(n6363), .Z(n6365) );
  NAND U6580 ( .A(n6366), .B(n6365), .Z(n6446) );
  XNOR U6581 ( .A(n6445), .B(n6446), .Z(n6447) );
  XOR U6582 ( .A(n6448), .B(n6447), .Z(n6378) );
  NANDN U6583 ( .A(n6368), .B(n6367), .Z(n6372) );
  NANDN U6584 ( .A(n6370), .B(n6369), .Z(n6371) );
  NAND U6585 ( .A(n6372), .B(n6371), .Z(n6379) );
  XNOR U6586 ( .A(n6378), .B(n6379), .Z(n6380) );
  XNOR U6587 ( .A(n6381), .B(n6380), .Z(n6451) );
  XNOR U6588 ( .A(n6451), .B(sreg[328]), .Z(n6453) );
  NAND U6589 ( .A(n6373), .B(sreg[327]), .Z(n6377) );
  OR U6590 ( .A(n6375), .B(n6374), .Z(n6376) );
  AND U6591 ( .A(n6377), .B(n6376), .Z(n6452) );
  XOR U6592 ( .A(n6453), .B(n6452), .Z(c[328]) );
  NANDN U6593 ( .A(n6379), .B(n6378), .Z(n6383) );
  NAND U6594 ( .A(n6381), .B(n6380), .Z(n6382) );
  NAND U6595 ( .A(n6383), .B(n6382), .Z(n6459) );
  NANDN U6596 ( .A(n6385), .B(n6384), .Z(n6389) );
  OR U6597 ( .A(n6387), .B(n6386), .Z(n6388) );
  NAND U6598 ( .A(n6389), .B(n6388), .Z(n6526) );
  XNOR U6599 ( .A(n20052), .B(n6705), .Z(n6468) );
  OR U6600 ( .A(n6468), .B(n20020), .Z(n6392) );
  NANDN U6601 ( .A(n6390), .B(n19960), .Z(n6391) );
  NAND U6602 ( .A(n6392), .B(n6391), .Z(n6481) );
  XNOR U6603 ( .A(n102), .B(n6393), .Z(n6472) );
  OR U6604 ( .A(n6472), .B(n20121), .Z(n6396) );
  NANDN U6605 ( .A(n6394), .B(n20122), .Z(n6395) );
  NAND U6606 ( .A(n6396), .B(n6395), .Z(n6478) );
  XNOR U6607 ( .A(n19975), .B(n6888), .Z(n6475) );
  NANDN U6608 ( .A(n6475), .B(n19883), .Z(n6399) );
  NANDN U6609 ( .A(n6397), .B(n19937), .Z(n6398) );
  AND U6610 ( .A(n6399), .B(n6398), .Z(n6479) );
  XNOR U6611 ( .A(n6478), .B(n6479), .Z(n6480) );
  XNOR U6612 ( .A(n6481), .B(n6480), .Z(n6517) );
  NANDN U6613 ( .A(n6401), .B(n6400), .Z(n6405) );
  NAND U6614 ( .A(n6403), .B(n6402), .Z(n6404) );
  NAND U6615 ( .A(n6405), .B(n6404), .Z(n6518) );
  XNOR U6616 ( .A(n6517), .B(n6518), .Z(n6519) );
  NANDN U6617 ( .A(n6407), .B(n6406), .Z(n6411) );
  NAND U6618 ( .A(n6409), .B(n6408), .Z(n6410) );
  AND U6619 ( .A(n6411), .B(n6410), .Z(n6520) );
  XNOR U6620 ( .A(n6519), .B(n6520), .Z(n6464) );
  NANDN U6621 ( .A(n6413), .B(n6412), .Z(n6417) );
  OR U6622 ( .A(n6415), .B(n6414), .Z(n6416) );
  NAND U6623 ( .A(n6417), .B(n6416), .Z(n6514) );
  NAND U6624 ( .A(b[0]), .B(a[89]), .Z(n6418) );
  XNOR U6625 ( .A(b[1]), .B(n6418), .Z(n6420) );
  NAND U6626 ( .A(a[88]), .B(n98), .Z(n6419) );
  AND U6627 ( .A(n6420), .B(n6419), .Z(n6490) );
  XNOR U6628 ( .A(n20154), .B(n6549), .Z(n6499) );
  OR U6629 ( .A(n6499), .B(n20057), .Z(n6423) );
  NANDN U6630 ( .A(n6421), .B(n20098), .Z(n6422) );
  AND U6631 ( .A(n6423), .B(n6422), .Z(n6491) );
  XOR U6632 ( .A(n6490), .B(n6491), .Z(n6493) );
  NAND U6633 ( .A(a[73]), .B(b[15]), .Z(n6492) );
  XOR U6634 ( .A(n6493), .B(n6492), .Z(n6511) );
  NAND U6635 ( .A(n19722), .B(n6424), .Z(n6426) );
  XNOR U6636 ( .A(b[5]), .B(n7173), .Z(n6502) );
  NANDN U6637 ( .A(n19640), .B(n6502), .Z(n6425) );
  NAND U6638 ( .A(n6426), .B(n6425), .Z(n6487) );
  XNOR U6639 ( .A(n19714), .B(n7044), .Z(n6505) );
  NANDN U6640 ( .A(n6505), .B(n19766), .Z(n6429) );
  NANDN U6641 ( .A(n6427), .B(n19767), .Z(n6428) );
  NAND U6642 ( .A(n6429), .B(n6428), .Z(n6484) );
  NAND U6643 ( .A(n19554), .B(n6430), .Z(n6432) );
  IV U6644 ( .A(a[87]), .Z(n7329) );
  XNOR U6645 ( .A(b[3]), .B(n7329), .Z(n6508) );
  NANDN U6646 ( .A(n19521), .B(n6508), .Z(n6431) );
  AND U6647 ( .A(n6432), .B(n6431), .Z(n6485) );
  XNOR U6648 ( .A(n6484), .B(n6485), .Z(n6486) );
  XOR U6649 ( .A(n6487), .B(n6486), .Z(n6512) );
  XOR U6650 ( .A(n6511), .B(n6512), .Z(n6513) );
  XNOR U6651 ( .A(n6514), .B(n6513), .Z(n6462) );
  NAND U6652 ( .A(n6434), .B(n6433), .Z(n6438) );
  NAND U6653 ( .A(n6436), .B(n6435), .Z(n6437) );
  NAND U6654 ( .A(n6438), .B(n6437), .Z(n6463) );
  XOR U6655 ( .A(n6462), .B(n6463), .Z(n6465) );
  XNOR U6656 ( .A(n6464), .B(n6465), .Z(n6523) );
  NANDN U6657 ( .A(n6440), .B(n6439), .Z(n6444) );
  NAND U6658 ( .A(n6442), .B(n6441), .Z(n6443) );
  NAND U6659 ( .A(n6444), .B(n6443), .Z(n6524) );
  XNOR U6660 ( .A(n6523), .B(n6524), .Z(n6525) );
  XOR U6661 ( .A(n6526), .B(n6525), .Z(n6456) );
  NANDN U6662 ( .A(n6446), .B(n6445), .Z(n6450) );
  NANDN U6663 ( .A(n6448), .B(n6447), .Z(n6449) );
  NAND U6664 ( .A(n6450), .B(n6449), .Z(n6457) );
  XNOR U6665 ( .A(n6456), .B(n6457), .Z(n6458) );
  XNOR U6666 ( .A(n6459), .B(n6458), .Z(n6529) );
  XNOR U6667 ( .A(n6529), .B(sreg[329]), .Z(n6531) );
  NAND U6668 ( .A(n6451), .B(sreg[328]), .Z(n6455) );
  OR U6669 ( .A(n6453), .B(n6452), .Z(n6454) );
  AND U6670 ( .A(n6455), .B(n6454), .Z(n6530) );
  XOR U6671 ( .A(n6531), .B(n6530), .Z(c[329]) );
  NANDN U6672 ( .A(n6457), .B(n6456), .Z(n6461) );
  NAND U6673 ( .A(n6459), .B(n6458), .Z(n6460) );
  NAND U6674 ( .A(n6461), .B(n6460), .Z(n6537) );
  NANDN U6675 ( .A(n6463), .B(n6462), .Z(n6467) );
  OR U6676 ( .A(n6465), .B(n6464), .Z(n6466) );
  NAND U6677 ( .A(n6467), .B(n6466), .Z(n6604) );
  XNOR U6678 ( .A(n20052), .B(n6783), .Z(n6546) );
  OR U6679 ( .A(n6546), .B(n20020), .Z(n6470) );
  NANDN U6680 ( .A(n6468), .B(n19960), .Z(n6469) );
  NAND U6681 ( .A(n6470), .B(n6469), .Z(n6559) );
  XNOR U6682 ( .A(n102), .B(n6471), .Z(n6550) );
  OR U6683 ( .A(n6550), .B(n20121), .Z(n6474) );
  NANDN U6684 ( .A(n6472), .B(n20122), .Z(n6473) );
  NAND U6685 ( .A(n6474), .B(n6473), .Z(n6556) );
  XNOR U6686 ( .A(n19975), .B(n6951), .Z(n6553) );
  NANDN U6687 ( .A(n6553), .B(n19883), .Z(n6477) );
  NANDN U6688 ( .A(n6475), .B(n19937), .Z(n6476) );
  AND U6689 ( .A(n6477), .B(n6476), .Z(n6557) );
  XNOR U6690 ( .A(n6556), .B(n6557), .Z(n6558) );
  XNOR U6691 ( .A(n6559), .B(n6558), .Z(n6595) );
  NANDN U6692 ( .A(n6479), .B(n6478), .Z(n6483) );
  NAND U6693 ( .A(n6481), .B(n6480), .Z(n6482) );
  NAND U6694 ( .A(n6483), .B(n6482), .Z(n6596) );
  XNOR U6695 ( .A(n6595), .B(n6596), .Z(n6597) );
  NANDN U6696 ( .A(n6485), .B(n6484), .Z(n6489) );
  NAND U6697 ( .A(n6487), .B(n6486), .Z(n6488) );
  AND U6698 ( .A(n6489), .B(n6488), .Z(n6598) );
  XNOR U6699 ( .A(n6597), .B(n6598), .Z(n6542) );
  NANDN U6700 ( .A(n6491), .B(n6490), .Z(n6495) );
  OR U6701 ( .A(n6493), .B(n6492), .Z(n6494) );
  NAND U6702 ( .A(n6495), .B(n6494), .Z(n6592) );
  NAND U6703 ( .A(b[0]), .B(a[90]), .Z(n6496) );
  XNOR U6704 ( .A(b[1]), .B(n6496), .Z(n6498) );
  NAND U6705 ( .A(a[89]), .B(n98), .Z(n6497) );
  AND U6706 ( .A(n6498), .B(n6497), .Z(n6568) );
  XNOR U6707 ( .A(n20154), .B(n6627), .Z(n6577) );
  OR U6708 ( .A(n6577), .B(n20057), .Z(n6501) );
  NANDN U6709 ( .A(n6499), .B(n20098), .Z(n6500) );
  AND U6710 ( .A(n6501), .B(n6500), .Z(n6569) );
  XOR U6711 ( .A(n6568), .B(n6569), .Z(n6571) );
  NAND U6712 ( .A(a[74]), .B(b[15]), .Z(n6570) );
  XOR U6713 ( .A(n6571), .B(n6570), .Z(n6589) );
  NAND U6714 ( .A(n19722), .B(n6502), .Z(n6504) );
  XNOR U6715 ( .A(b[5]), .B(n7251), .Z(n6580) );
  NANDN U6716 ( .A(n19640), .B(n6580), .Z(n6503) );
  NAND U6717 ( .A(n6504), .B(n6503), .Z(n6565) );
  XNOR U6718 ( .A(n19714), .B(n7095), .Z(n6583) );
  NANDN U6719 ( .A(n6583), .B(n19766), .Z(n6507) );
  NANDN U6720 ( .A(n6505), .B(n19767), .Z(n6506) );
  NAND U6721 ( .A(n6507), .B(n6506), .Z(n6562) );
  NAND U6722 ( .A(n19554), .B(n6508), .Z(n6510) );
  IV U6723 ( .A(a[88]), .Z(n7407) );
  XNOR U6724 ( .A(b[3]), .B(n7407), .Z(n6586) );
  NANDN U6725 ( .A(n19521), .B(n6586), .Z(n6509) );
  AND U6726 ( .A(n6510), .B(n6509), .Z(n6563) );
  XNOR U6727 ( .A(n6562), .B(n6563), .Z(n6564) );
  XOR U6728 ( .A(n6565), .B(n6564), .Z(n6590) );
  XOR U6729 ( .A(n6589), .B(n6590), .Z(n6591) );
  XNOR U6730 ( .A(n6592), .B(n6591), .Z(n6540) );
  NAND U6731 ( .A(n6512), .B(n6511), .Z(n6516) );
  NAND U6732 ( .A(n6514), .B(n6513), .Z(n6515) );
  NAND U6733 ( .A(n6516), .B(n6515), .Z(n6541) );
  XOR U6734 ( .A(n6540), .B(n6541), .Z(n6543) );
  XNOR U6735 ( .A(n6542), .B(n6543), .Z(n6601) );
  NANDN U6736 ( .A(n6518), .B(n6517), .Z(n6522) );
  NAND U6737 ( .A(n6520), .B(n6519), .Z(n6521) );
  NAND U6738 ( .A(n6522), .B(n6521), .Z(n6602) );
  XNOR U6739 ( .A(n6601), .B(n6602), .Z(n6603) );
  XOR U6740 ( .A(n6604), .B(n6603), .Z(n6534) );
  NANDN U6741 ( .A(n6524), .B(n6523), .Z(n6528) );
  NANDN U6742 ( .A(n6526), .B(n6525), .Z(n6527) );
  NAND U6743 ( .A(n6528), .B(n6527), .Z(n6535) );
  XNOR U6744 ( .A(n6534), .B(n6535), .Z(n6536) );
  XNOR U6745 ( .A(n6537), .B(n6536), .Z(n6607) );
  XNOR U6746 ( .A(n6607), .B(sreg[330]), .Z(n6609) );
  NAND U6747 ( .A(n6529), .B(sreg[329]), .Z(n6533) );
  OR U6748 ( .A(n6531), .B(n6530), .Z(n6532) );
  AND U6749 ( .A(n6533), .B(n6532), .Z(n6608) );
  XOR U6750 ( .A(n6609), .B(n6608), .Z(c[330]) );
  NANDN U6751 ( .A(n6535), .B(n6534), .Z(n6539) );
  NAND U6752 ( .A(n6537), .B(n6536), .Z(n6538) );
  NAND U6753 ( .A(n6539), .B(n6538), .Z(n6615) );
  NANDN U6754 ( .A(n6541), .B(n6540), .Z(n6545) );
  OR U6755 ( .A(n6543), .B(n6542), .Z(n6544) );
  NAND U6756 ( .A(n6545), .B(n6544), .Z(n6682) );
  XNOR U6757 ( .A(n20052), .B(n6888), .Z(n6624) );
  OR U6758 ( .A(n6624), .B(n20020), .Z(n6548) );
  NANDN U6759 ( .A(n6546), .B(n19960), .Z(n6547) );
  NAND U6760 ( .A(n6548), .B(n6547), .Z(n6637) );
  XNOR U6761 ( .A(n102), .B(n6549), .Z(n6628) );
  OR U6762 ( .A(n6628), .B(n20121), .Z(n6552) );
  NANDN U6763 ( .A(n6550), .B(n20122), .Z(n6551) );
  NAND U6764 ( .A(n6552), .B(n6551), .Z(n6634) );
  XNOR U6765 ( .A(n19975), .B(n7044), .Z(n6631) );
  NANDN U6766 ( .A(n6631), .B(n19883), .Z(n6555) );
  NANDN U6767 ( .A(n6553), .B(n19937), .Z(n6554) );
  AND U6768 ( .A(n6555), .B(n6554), .Z(n6635) );
  XNOR U6769 ( .A(n6634), .B(n6635), .Z(n6636) );
  XNOR U6770 ( .A(n6637), .B(n6636), .Z(n6673) );
  NANDN U6771 ( .A(n6557), .B(n6556), .Z(n6561) );
  NAND U6772 ( .A(n6559), .B(n6558), .Z(n6560) );
  NAND U6773 ( .A(n6561), .B(n6560), .Z(n6674) );
  XNOR U6774 ( .A(n6673), .B(n6674), .Z(n6675) );
  NANDN U6775 ( .A(n6563), .B(n6562), .Z(n6567) );
  NAND U6776 ( .A(n6565), .B(n6564), .Z(n6566) );
  AND U6777 ( .A(n6567), .B(n6566), .Z(n6676) );
  XNOR U6778 ( .A(n6675), .B(n6676), .Z(n6620) );
  NANDN U6779 ( .A(n6569), .B(n6568), .Z(n6573) );
  OR U6780 ( .A(n6571), .B(n6570), .Z(n6572) );
  NAND U6781 ( .A(n6573), .B(n6572), .Z(n6670) );
  NAND U6782 ( .A(b[0]), .B(a[91]), .Z(n6574) );
  XNOR U6783 ( .A(b[1]), .B(n6574), .Z(n6576) );
  NAND U6784 ( .A(a[90]), .B(n98), .Z(n6575) );
  AND U6785 ( .A(n6576), .B(n6575), .Z(n6646) );
  XNOR U6786 ( .A(n20154), .B(n6705), .Z(n6652) );
  OR U6787 ( .A(n6652), .B(n20057), .Z(n6579) );
  NANDN U6788 ( .A(n6577), .B(n20098), .Z(n6578) );
  AND U6789 ( .A(n6579), .B(n6578), .Z(n6647) );
  XOR U6790 ( .A(n6646), .B(n6647), .Z(n6649) );
  NAND U6791 ( .A(a[75]), .B(b[15]), .Z(n6648) );
  XOR U6792 ( .A(n6649), .B(n6648), .Z(n6667) );
  NAND U6793 ( .A(n19722), .B(n6580), .Z(n6582) );
  XNOR U6794 ( .A(b[5]), .B(n7329), .Z(n6658) );
  NANDN U6795 ( .A(n19640), .B(n6658), .Z(n6581) );
  NAND U6796 ( .A(n6582), .B(n6581), .Z(n6643) );
  XNOR U6797 ( .A(n19714), .B(n7173), .Z(n6661) );
  NANDN U6798 ( .A(n6661), .B(n19766), .Z(n6585) );
  NANDN U6799 ( .A(n6583), .B(n19767), .Z(n6584) );
  NAND U6800 ( .A(n6585), .B(n6584), .Z(n6640) );
  NAND U6801 ( .A(n19554), .B(n6586), .Z(n6588) );
  IV U6802 ( .A(a[89]), .Z(n7485) );
  XNOR U6803 ( .A(b[3]), .B(n7485), .Z(n6664) );
  NANDN U6804 ( .A(n19521), .B(n6664), .Z(n6587) );
  AND U6805 ( .A(n6588), .B(n6587), .Z(n6641) );
  XNOR U6806 ( .A(n6640), .B(n6641), .Z(n6642) );
  XOR U6807 ( .A(n6643), .B(n6642), .Z(n6668) );
  XOR U6808 ( .A(n6667), .B(n6668), .Z(n6669) );
  XNOR U6809 ( .A(n6670), .B(n6669), .Z(n6618) );
  NAND U6810 ( .A(n6590), .B(n6589), .Z(n6594) );
  NAND U6811 ( .A(n6592), .B(n6591), .Z(n6593) );
  NAND U6812 ( .A(n6594), .B(n6593), .Z(n6619) );
  XOR U6813 ( .A(n6618), .B(n6619), .Z(n6621) );
  XNOR U6814 ( .A(n6620), .B(n6621), .Z(n6679) );
  NANDN U6815 ( .A(n6596), .B(n6595), .Z(n6600) );
  NAND U6816 ( .A(n6598), .B(n6597), .Z(n6599) );
  NAND U6817 ( .A(n6600), .B(n6599), .Z(n6680) );
  XNOR U6818 ( .A(n6679), .B(n6680), .Z(n6681) );
  XOR U6819 ( .A(n6682), .B(n6681), .Z(n6612) );
  NANDN U6820 ( .A(n6602), .B(n6601), .Z(n6606) );
  NANDN U6821 ( .A(n6604), .B(n6603), .Z(n6605) );
  NAND U6822 ( .A(n6606), .B(n6605), .Z(n6613) );
  XNOR U6823 ( .A(n6612), .B(n6613), .Z(n6614) );
  XNOR U6824 ( .A(n6615), .B(n6614), .Z(n6685) );
  XNOR U6825 ( .A(n6685), .B(sreg[331]), .Z(n6687) );
  NAND U6826 ( .A(n6607), .B(sreg[330]), .Z(n6611) );
  OR U6827 ( .A(n6609), .B(n6608), .Z(n6610) );
  AND U6828 ( .A(n6611), .B(n6610), .Z(n6686) );
  XOR U6829 ( .A(n6687), .B(n6686), .Z(c[331]) );
  NANDN U6830 ( .A(n6613), .B(n6612), .Z(n6617) );
  NAND U6831 ( .A(n6615), .B(n6614), .Z(n6616) );
  NAND U6832 ( .A(n6617), .B(n6616), .Z(n6693) );
  NANDN U6833 ( .A(n6619), .B(n6618), .Z(n6623) );
  OR U6834 ( .A(n6621), .B(n6620), .Z(n6622) );
  NAND U6835 ( .A(n6623), .B(n6622), .Z(n6760) );
  XNOR U6836 ( .A(n20052), .B(n6951), .Z(n6702) );
  OR U6837 ( .A(n6702), .B(n20020), .Z(n6626) );
  NANDN U6838 ( .A(n6624), .B(n19960), .Z(n6625) );
  NAND U6839 ( .A(n6626), .B(n6625), .Z(n6715) );
  XNOR U6840 ( .A(n102), .B(n6627), .Z(n6706) );
  OR U6841 ( .A(n6706), .B(n20121), .Z(n6630) );
  NANDN U6842 ( .A(n6628), .B(n20122), .Z(n6629) );
  NAND U6843 ( .A(n6630), .B(n6629), .Z(n6712) );
  XNOR U6844 ( .A(n19975), .B(n7095), .Z(n6709) );
  NANDN U6845 ( .A(n6709), .B(n19883), .Z(n6633) );
  NANDN U6846 ( .A(n6631), .B(n19937), .Z(n6632) );
  AND U6847 ( .A(n6633), .B(n6632), .Z(n6713) );
  XNOR U6848 ( .A(n6712), .B(n6713), .Z(n6714) );
  XNOR U6849 ( .A(n6715), .B(n6714), .Z(n6751) );
  NANDN U6850 ( .A(n6635), .B(n6634), .Z(n6639) );
  NAND U6851 ( .A(n6637), .B(n6636), .Z(n6638) );
  NAND U6852 ( .A(n6639), .B(n6638), .Z(n6752) );
  XNOR U6853 ( .A(n6751), .B(n6752), .Z(n6753) );
  NANDN U6854 ( .A(n6641), .B(n6640), .Z(n6645) );
  NAND U6855 ( .A(n6643), .B(n6642), .Z(n6644) );
  AND U6856 ( .A(n6645), .B(n6644), .Z(n6754) );
  XNOR U6857 ( .A(n6753), .B(n6754), .Z(n6698) );
  NANDN U6858 ( .A(n6647), .B(n6646), .Z(n6651) );
  OR U6859 ( .A(n6649), .B(n6648), .Z(n6650) );
  NAND U6860 ( .A(n6651), .B(n6650), .Z(n6748) );
  XNOR U6861 ( .A(n20154), .B(n6783), .Z(n6733) );
  OR U6862 ( .A(n6733), .B(n20057), .Z(n6654) );
  NANDN U6863 ( .A(n6652), .B(n20098), .Z(n6653) );
  AND U6864 ( .A(n6654), .B(n6653), .Z(n6725) );
  NAND U6865 ( .A(b[0]), .B(a[92]), .Z(n6655) );
  XNOR U6866 ( .A(b[1]), .B(n6655), .Z(n6657) );
  NAND U6867 ( .A(a[91]), .B(n98), .Z(n6656) );
  AND U6868 ( .A(n6657), .B(n6656), .Z(n6724) );
  XOR U6869 ( .A(n6725), .B(n6724), .Z(n6727) );
  NAND U6870 ( .A(a[76]), .B(b[15]), .Z(n6726) );
  XOR U6871 ( .A(n6727), .B(n6726), .Z(n6745) );
  NAND U6872 ( .A(n19722), .B(n6658), .Z(n6660) );
  XNOR U6873 ( .A(b[5]), .B(n7407), .Z(n6736) );
  NANDN U6874 ( .A(n19640), .B(n6736), .Z(n6659) );
  NAND U6875 ( .A(n6660), .B(n6659), .Z(n6721) );
  XNOR U6876 ( .A(n19714), .B(n7251), .Z(n6739) );
  NANDN U6877 ( .A(n6739), .B(n19766), .Z(n6663) );
  NANDN U6878 ( .A(n6661), .B(n19767), .Z(n6662) );
  NAND U6879 ( .A(n6663), .B(n6662), .Z(n6718) );
  NAND U6880 ( .A(n19554), .B(n6664), .Z(n6666) );
  IV U6881 ( .A(a[90]), .Z(n7563) );
  XNOR U6882 ( .A(b[3]), .B(n7563), .Z(n6742) );
  NANDN U6883 ( .A(n19521), .B(n6742), .Z(n6665) );
  AND U6884 ( .A(n6666), .B(n6665), .Z(n6719) );
  XNOR U6885 ( .A(n6718), .B(n6719), .Z(n6720) );
  XOR U6886 ( .A(n6721), .B(n6720), .Z(n6746) );
  XOR U6887 ( .A(n6745), .B(n6746), .Z(n6747) );
  XNOR U6888 ( .A(n6748), .B(n6747), .Z(n6696) );
  NAND U6889 ( .A(n6668), .B(n6667), .Z(n6672) );
  NAND U6890 ( .A(n6670), .B(n6669), .Z(n6671) );
  NAND U6891 ( .A(n6672), .B(n6671), .Z(n6697) );
  XOR U6892 ( .A(n6696), .B(n6697), .Z(n6699) );
  XNOR U6893 ( .A(n6698), .B(n6699), .Z(n6757) );
  NANDN U6894 ( .A(n6674), .B(n6673), .Z(n6678) );
  NAND U6895 ( .A(n6676), .B(n6675), .Z(n6677) );
  NAND U6896 ( .A(n6678), .B(n6677), .Z(n6758) );
  XNOR U6897 ( .A(n6757), .B(n6758), .Z(n6759) );
  XOR U6898 ( .A(n6760), .B(n6759), .Z(n6690) );
  NANDN U6899 ( .A(n6680), .B(n6679), .Z(n6684) );
  NANDN U6900 ( .A(n6682), .B(n6681), .Z(n6683) );
  NAND U6901 ( .A(n6684), .B(n6683), .Z(n6691) );
  XNOR U6902 ( .A(n6690), .B(n6691), .Z(n6692) );
  XNOR U6903 ( .A(n6693), .B(n6692), .Z(n6763) );
  XNOR U6904 ( .A(n6763), .B(sreg[332]), .Z(n6765) );
  NAND U6905 ( .A(n6685), .B(sreg[331]), .Z(n6689) );
  OR U6906 ( .A(n6687), .B(n6686), .Z(n6688) );
  AND U6907 ( .A(n6689), .B(n6688), .Z(n6764) );
  XOR U6908 ( .A(n6765), .B(n6764), .Z(c[332]) );
  NANDN U6909 ( .A(n6691), .B(n6690), .Z(n6695) );
  NAND U6910 ( .A(n6693), .B(n6692), .Z(n6694) );
  NAND U6911 ( .A(n6695), .B(n6694), .Z(n6771) );
  NANDN U6912 ( .A(n6697), .B(n6696), .Z(n6701) );
  OR U6913 ( .A(n6699), .B(n6698), .Z(n6700) );
  NAND U6914 ( .A(n6701), .B(n6700), .Z(n6838) );
  XNOR U6915 ( .A(n20052), .B(n7044), .Z(n6780) );
  OR U6916 ( .A(n6780), .B(n20020), .Z(n6704) );
  NANDN U6917 ( .A(n6702), .B(n19960), .Z(n6703) );
  NAND U6918 ( .A(n6704), .B(n6703), .Z(n6793) );
  XNOR U6919 ( .A(n102), .B(n6705), .Z(n6784) );
  OR U6920 ( .A(n6784), .B(n20121), .Z(n6708) );
  NANDN U6921 ( .A(n6706), .B(n20122), .Z(n6707) );
  NAND U6922 ( .A(n6708), .B(n6707), .Z(n6790) );
  XNOR U6923 ( .A(n19975), .B(n7173), .Z(n6787) );
  NANDN U6924 ( .A(n6787), .B(n19883), .Z(n6711) );
  NANDN U6925 ( .A(n6709), .B(n19937), .Z(n6710) );
  AND U6926 ( .A(n6711), .B(n6710), .Z(n6791) );
  XNOR U6927 ( .A(n6790), .B(n6791), .Z(n6792) );
  XNOR U6928 ( .A(n6793), .B(n6792), .Z(n6829) );
  NANDN U6929 ( .A(n6713), .B(n6712), .Z(n6717) );
  NAND U6930 ( .A(n6715), .B(n6714), .Z(n6716) );
  NAND U6931 ( .A(n6717), .B(n6716), .Z(n6830) );
  XNOR U6932 ( .A(n6829), .B(n6830), .Z(n6831) );
  NANDN U6933 ( .A(n6719), .B(n6718), .Z(n6723) );
  NAND U6934 ( .A(n6721), .B(n6720), .Z(n6722) );
  AND U6935 ( .A(n6723), .B(n6722), .Z(n6832) );
  XNOR U6936 ( .A(n6831), .B(n6832), .Z(n6776) );
  NANDN U6937 ( .A(n6725), .B(n6724), .Z(n6729) );
  OR U6938 ( .A(n6727), .B(n6726), .Z(n6728) );
  NAND U6939 ( .A(n6729), .B(n6728), .Z(n6826) );
  NAND U6940 ( .A(b[0]), .B(a[93]), .Z(n6730) );
  XNOR U6941 ( .A(b[1]), .B(n6730), .Z(n6732) );
  NAND U6942 ( .A(a[92]), .B(n98), .Z(n6731) );
  AND U6943 ( .A(n6732), .B(n6731), .Z(n6802) );
  XNOR U6944 ( .A(n20154), .B(n6888), .Z(n6811) );
  OR U6945 ( .A(n6811), .B(n20057), .Z(n6735) );
  NANDN U6946 ( .A(n6733), .B(n20098), .Z(n6734) );
  AND U6947 ( .A(n6735), .B(n6734), .Z(n6803) );
  XOR U6948 ( .A(n6802), .B(n6803), .Z(n6805) );
  NAND U6949 ( .A(a[77]), .B(b[15]), .Z(n6804) );
  XOR U6950 ( .A(n6805), .B(n6804), .Z(n6823) );
  NAND U6951 ( .A(n19722), .B(n6736), .Z(n6738) );
  XNOR U6952 ( .A(b[5]), .B(n7485), .Z(n6814) );
  NANDN U6953 ( .A(n19640), .B(n6814), .Z(n6737) );
  NAND U6954 ( .A(n6738), .B(n6737), .Z(n6799) );
  XNOR U6955 ( .A(n19714), .B(n7329), .Z(n6817) );
  NANDN U6956 ( .A(n6817), .B(n19766), .Z(n6741) );
  NANDN U6957 ( .A(n6739), .B(n19767), .Z(n6740) );
  NAND U6958 ( .A(n6741), .B(n6740), .Z(n6796) );
  NAND U6959 ( .A(n19554), .B(n6742), .Z(n6744) );
  IV U6960 ( .A(a[91]), .Z(n7641) );
  XNOR U6961 ( .A(b[3]), .B(n7641), .Z(n6820) );
  NANDN U6962 ( .A(n19521), .B(n6820), .Z(n6743) );
  AND U6963 ( .A(n6744), .B(n6743), .Z(n6797) );
  XNOR U6964 ( .A(n6796), .B(n6797), .Z(n6798) );
  XOR U6965 ( .A(n6799), .B(n6798), .Z(n6824) );
  XOR U6966 ( .A(n6823), .B(n6824), .Z(n6825) );
  XNOR U6967 ( .A(n6826), .B(n6825), .Z(n6774) );
  NAND U6968 ( .A(n6746), .B(n6745), .Z(n6750) );
  NAND U6969 ( .A(n6748), .B(n6747), .Z(n6749) );
  NAND U6970 ( .A(n6750), .B(n6749), .Z(n6775) );
  XOR U6971 ( .A(n6774), .B(n6775), .Z(n6777) );
  XNOR U6972 ( .A(n6776), .B(n6777), .Z(n6835) );
  NANDN U6973 ( .A(n6752), .B(n6751), .Z(n6756) );
  NAND U6974 ( .A(n6754), .B(n6753), .Z(n6755) );
  NAND U6975 ( .A(n6756), .B(n6755), .Z(n6836) );
  XNOR U6976 ( .A(n6835), .B(n6836), .Z(n6837) );
  XOR U6977 ( .A(n6838), .B(n6837), .Z(n6768) );
  NANDN U6978 ( .A(n6758), .B(n6757), .Z(n6762) );
  NANDN U6979 ( .A(n6760), .B(n6759), .Z(n6761) );
  NAND U6980 ( .A(n6762), .B(n6761), .Z(n6769) );
  XNOR U6981 ( .A(n6768), .B(n6769), .Z(n6770) );
  XNOR U6982 ( .A(n6771), .B(n6770), .Z(n6841) );
  XNOR U6983 ( .A(n6841), .B(sreg[333]), .Z(n6843) );
  NAND U6984 ( .A(n6763), .B(sreg[332]), .Z(n6767) );
  OR U6985 ( .A(n6765), .B(n6764), .Z(n6766) );
  AND U6986 ( .A(n6767), .B(n6766), .Z(n6842) );
  XOR U6987 ( .A(n6843), .B(n6842), .Z(c[333]) );
  NANDN U6988 ( .A(n6769), .B(n6768), .Z(n6773) );
  NAND U6989 ( .A(n6771), .B(n6770), .Z(n6772) );
  NAND U6990 ( .A(n6773), .B(n6772), .Z(n6849) );
  NANDN U6991 ( .A(n6775), .B(n6774), .Z(n6779) );
  OR U6992 ( .A(n6777), .B(n6776), .Z(n6778) );
  NAND U6993 ( .A(n6779), .B(n6778), .Z(n6916) );
  XNOR U6994 ( .A(n20052), .B(n7095), .Z(n6885) );
  OR U6995 ( .A(n6885), .B(n20020), .Z(n6782) );
  NANDN U6996 ( .A(n6780), .B(n19960), .Z(n6781) );
  NAND U6997 ( .A(n6782), .B(n6781), .Z(n6898) );
  XNOR U6998 ( .A(n102), .B(n6783), .Z(n6889) );
  OR U6999 ( .A(n6889), .B(n20121), .Z(n6786) );
  NANDN U7000 ( .A(n6784), .B(n20122), .Z(n6785) );
  NAND U7001 ( .A(n6786), .B(n6785), .Z(n6895) );
  XNOR U7002 ( .A(n19975), .B(n7251), .Z(n6892) );
  NANDN U7003 ( .A(n6892), .B(n19883), .Z(n6789) );
  NANDN U7004 ( .A(n6787), .B(n19937), .Z(n6788) );
  AND U7005 ( .A(n6789), .B(n6788), .Z(n6896) );
  XNOR U7006 ( .A(n6895), .B(n6896), .Z(n6897) );
  XNOR U7007 ( .A(n6898), .B(n6897), .Z(n6907) );
  NANDN U7008 ( .A(n6791), .B(n6790), .Z(n6795) );
  NAND U7009 ( .A(n6793), .B(n6792), .Z(n6794) );
  NAND U7010 ( .A(n6795), .B(n6794), .Z(n6908) );
  XNOR U7011 ( .A(n6907), .B(n6908), .Z(n6909) );
  NANDN U7012 ( .A(n6797), .B(n6796), .Z(n6801) );
  NAND U7013 ( .A(n6799), .B(n6798), .Z(n6800) );
  AND U7014 ( .A(n6801), .B(n6800), .Z(n6910) );
  XNOR U7015 ( .A(n6909), .B(n6910), .Z(n6854) );
  NANDN U7016 ( .A(n6803), .B(n6802), .Z(n6807) );
  OR U7017 ( .A(n6805), .B(n6804), .Z(n6806) );
  NAND U7018 ( .A(n6807), .B(n6806), .Z(n6882) );
  NAND U7019 ( .A(b[0]), .B(a[94]), .Z(n6808) );
  XNOR U7020 ( .A(b[1]), .B(n6808), .Z(n6810) );
  NAND U7021 ( .A(a[93]), .B(n98), .Z(n6809) );
  AND U7022 ( .A(n6810), .B(n6809), .Z(n6858) );
  XNOR U7023 ( .A(n20154), .B(n6951), .Z(n6867) );
  OR U7024 ( .A(n6867), .B(n20057), .Z(n6813) );
  NANDN U7025 ( .A(n6811), .B(n20098), .Z(n6812) );
  AND U7026 ( .A(n6813), .B(n6812), .Z(n6859) );
  XOR U7027 ( .A(n6858), .B(n6859), .Z(n6861) );
  NAND U7028 ( .A(a[78]), .B(b[15]), .Z(n6860) );
  XOR U7029 ( .A(n6861), .B(n6860), .Z(n6879) );
  NAND U7030 ( .A(n19722), .B(n6814), .Z(n6816) );
  XNOR U7031 ( .A(b[5]), .B(n7563), .Z(n6870) );
  NANDN U7032 ( .A(n19640), .B(n6870), .Z(n6815) );
  NAND U7033 ( .A(n6816), .B(n6815), .Z(n6904) );
  XNOR U7034 ( .A(n19714), .B(n7407), .Z(n6873) );
  NANDN U7035 ( .A(n6873), .B(n19766), .Z(n6819) );
  NANDN U7036 ( .A(n6817), .B(n19767), .Z(n6818) );
  NAND U7037 ( .A(n6819), .B(n6818), .Z(n6901) );
  NAND U7038 ( .A(n19554), .B(n6820), .Z(n6822) );
  IV U7039 ( .A(a[92]), .Z(n7731) );
  XNOR U7040 ( .A(b[3]), .B(n7731), .Z(n6876) );
  NANDN U7041 ( .A(n19521), .B(n6876), .Z(n6821) );
  AND U7042 ( .A(n6822), .B(n6821), .Z(n6902) );
  XNOR U7043 ( .A(n6901), .B(n6902), .Z(n6903) );
  XOR U7044 ( .A(n6904), .B(n6903), .Z(n6880) );
  XOR U7045 ( .A(n6879), .B(n6880), .Z(n6881) );
  XNOR U7046 ( .A(n6882), .B(n6881), .Z(n6852) );
  NAND U7047 ( .A(n6824), .B(n6823), .Z(n6828) );
  NAND U7048 ( .A(n6826), .B(n6825), .Z(n6827) );
  NAND U7049 ( .A(n6828), .B(n6827), .Z(n6853) );
  XOR U7050 ( .A(n6852), .B(n6853), .Z(n6855) );
  XNOR U7051 ( .A(n6854), .B(n6855), .Z(n6913) );
  NANDN U7052 ( .A(n6830), .B(n6829), .Z(n6834) );
  NAND U7053 ( .A(n6832), .B(n6831), .Z(n6833) );
  NAND U7054 ( .A(n6834), .B(n6833), .Z(n6914) );
  XNOR U7055 ( .A(n6913), .B(n6914), .Z(n6915) );
  XOR U7056 ( .A(n6916), .B(n6915), .Z(n6846) );
  NANDN U7057 ( .A(n6836), .B(n6835), .Z(n6840) );
  NANDN U7058 ( .A(n6838), .B(n6837), .Z(n6839) );
  NAND U7059 ( .A(n6840), .B(n6839), .Z(n6847) );
  XNOR U7060 ( .A(n6846), .B(n6847), .Z(n6848) );
  XNOR U7061 ( .A(n6849), .B(n6848), .Z(n6919) );
  XNOR U7062 ( .A(n6919), .B(sreg[334]), .Z(n6921) );
  NAND U7063 ( .A(n6841), .B(sreg[333]), .Z(n6845) );
  OR U7064 ( .A(n6843), .B(n6842), .Z(n6844) );
  AND U7065 ( .A(n6845), .B(n6844), .Z(n6920) );
  XOR U7066 ( .A(n6921), .B(n6920), .Z(c[334]) );
  NANDN U7067 ( .A(n6847), .B(n6846), .Z(n6851) );
  NAND U7068 ( .A(n6849), .B(n6848), .Z(n6850) );
  NAND U7069 ( .A(n6851), .B(n6850), .Z(n6927) );
  NANDN U7070 ( .A(n6853), .B(n6852), .Z(n6857) );
  OR U7071 ( .A(n6855), .B(n6854), .Z(n6856) );
  NAND U7072 ( .A(n6857), .B(n6856), .Z(n6994) );
  NANDN U7073 ( .A(n6859), .B(n6858), .Z(n6863) );
  OR U7074 ( .A(n6861), .B(n6860), .Z(n6862) );
  NAND U7075 ( .A(n6863), .B(n6862), .Z(n6982) );
  NAND U7076 ( .A(b[0]), .B(a[95]), .Z(n6864) );
  XNOR U7077 ( .A(b[1]), .B(n6864), .Z(n6866) );
  NAND U7078 ( .A(a[94]), .B(n98), .Z(n6865) );
  AND U7079 ( .A(n6866), .B(n6865), .Z(n6958) );
  XNOR U7080 ( .A(n20154), .B(n7044), .Z(n6964) );
  OR U7081 ( .A(n6964), .B(n20057), .Z(n6869) );
  NANDN U7082 ( .A(n6867), .B(n20098), .Z(n6868) );
  AND U7083 ( .A(n6869), .B(n6868), .Z(n6959) );
  XOR U7084 ( .A(n6958), .B(n6959), .Z(n6961) );
  NAND U7085 ( .A(a[79]), .B(b[15]), .Z(n6960) );
  XOR U7086 ( .A(n6961), .B(n6960), .Z(n6979) );
  NAND U7087 ( .A(n19722), .B(n6870), .Z(n6872) );
  XNOR U7088 ( .A(b[5]), .B(n7641), .Z(n6970) );
  NANDN U7089 ( .A(n19640), .B(n6970), .Z(n6871) );
  NAND U7090 ( .A(n6872), .B(n6871), .Z(n6939) );
  XNOR U7091 ( .A(n19714), .B(n7485), .Z(n6973) );
  NANDN U7092 ( .A(n6973), .B(n19766), .Z(n6875) );
  NANDN U7093 ( .A(n6873), .B(n19767), .Z(n6874) );
  NAND U7094 ( .A(n6875), .B(n6874), .Z(n6936) );
  NAND U7095 ( .A(n19554), .B(n6876), .Z(n6878) );
  IV U7096 ( .A(a[93]), .Z(n7797) );
  XNOR U7097 ( .A(b[3]), .B(n7797), .Z(n6976) );
  NANDN U7098 ( .A(n19521), .B(n6976), .Z(n6877) );
  AND U7099 ( .A(n6878), .B(n6877), .Z(n6937) );
  XNOR U7100 ( .A(n6936), .B(n6937), .Z(n6938) );
  XOR U7101 ( .A(n6939), .B(n6938), .Z(n6980) );
  XOR U7102 ( .A(n6979), .B(n6980), .Z(n6981) );
  XNOR U7103 ( .A(n6982), .B(n6981), .Z(n6930) );
  NAND U7104 ( .A(n6880), .B(n6879), .Z(n6884) );
  NAND U7105 ( .A(n6882), .B(n6881), .Z(n6883) );
  NAND U7106 ( .A(n6884), .B(n6883), .Z(n6931) );
  XOR U7107 ( .A(n6930), .B(n6931), .Z(n6933) );
  XNOR U7108 ( .A(n20052), .B(n7173), .Z(n6948) );
  OR U7109 ( .A(n6948), .B(n20020), .Z(n6887) );
  NANDN U7110 ( .A(n6885), .B(n19960), .Z(n6886) );
  NAND U7111 ( .A(n6887), .B(n6886), .Z(n6945) );
  XNOR U7112 ( .A(n102), .B(n6888), .Z(n6952) );
  OR U7113 ( .A(n6952), .B(n20121), .Z(n6891) );
  NANDN U7114 ( .A(n6889), .B(n20122), .Z(n6890) );
  NAND U7115 ( .A(n6891), .B(n6890), .Z(n6942) );
  XNOR U7116 ( .A(n19975), .B(n7329), .Z(n6955) );
  NANDN U7117 ( .A(n6955), .B(n19883), .Z(n6894) );
  NANDN U7118 ( .A(n6892), .B(n19937), .Z(n6893) );
  AND U7119 ( .A(n6894), .B(n6893), .Z(n6943) );
  XNOR U7120 ( .A(n6942), .B(n6943), .Z(n6944) );
  XNOR U7121 ( .A(n6945), .B(n6944), .Z(n6985) );
  NANDN U7122 ( .A(n6896), .B(n6895), .Z(n6900) );
  NAND U7123 ( .A(n6898), .B(n6897), .Z(n6899) );
  NAND U7124 ( .A(n6900), .B(n6899), .Z(n6986) );
  XNOR U7125 ( .A(n6985), .B(n6986), .Z(n6987) );
  NANDN U7126 ( .A(n6902), .B(n6901), .Z(n6906) );
  NAND U7127 ( .A(n6904), .B(n6903), .Z(n6905) );
  AND U7128 ( .A(n6906), .B(n6905), .Z(n6988) );
  XNOR U7129 ( .A(n6987), .B(n6988), .Z(n6932) );
  XNOR U7130 ( .A(n6933), .B(n6932), .Z(n6991) );
  NANDN U7131 ( .A(n6908), .B(n6907), .Z(n6912) );
  NAND U7132 ( .A(n6910), .B(n6909), .Z(n6911) );
  NAND U7133 ( .A(n6912), .B(n6911), .Z(n6992) );
  XNOR U7134 ( .A(n6991), .B(n6992), .Z(n6993) );
  XOR U7135 ( .A(n6994), .B(n6993), .Z(n6924) );
  NANDN U7136 ( .A(n6914), .B(n6913), .Z(n6918) );
  NANDN U7137 ( .A(n6916), .B(n6915), .Z(n6917) );
  NAND U7138 ( .A(n6918), .B(n6917), .Z(n6925) );
  XNOR U7139 ( .A(n6924), .B(n6925), .Z(n6926) );
  XNOR U7140 ( .A(n6927), .B(n6926), .Z(n6997) );
  XNOR U7141 ( .A(n6997), .B(sreg[335]), .Z(n6999) );
  NAND U7142 ( .A(n6919), .B(sreg[334]), .Z(n6923) );
  OR U7143 ( .A(n6921), .B(n6920), .Z(n6922) );
  AND U7144 ( .A(n6923), .B(n6922), .Z(n6998) );
  XOR U7145 ( .A(n6999), .B(n6998), .Z(c[335]) );
  NANDN U7146 ( .A(n6925), .B(n6924), .Z(n6929) );
  NAND U7147 ( .A(n6927), .B(n6926), .Z(n6928) );
  NAND U7148 ( .A(n6929), .B(n6928), .Z(n7005) );
  NANDN U7149 ( .A(n6931), .B(n6930), .Z(n6935) );
  OR U7150 ( .A(n6933), .B(n6932), .Z(n6934) );
  NAND U7151 ( .A(n6935), .B(n6934), .Z(n7072) );
  NANDN U7152 ( .A(n6937), .B(n6936), .Z(n6941) );
  NAND U7153 ( .A(n6939), .B(n6938), .Z(n6940) );
  NAND U7154 ( .A(n6941), .B(n6940), .Z(n7066) );
  NANDN U7155 ( .A(n6943), .B(n6942), .Z(n6947) );
  NAND U7156 ( .A(n6945), .B(n6944), .Z(n6946) );
  NAND U7157 ( .A(n6947), .B(n6946), .Z(n7063) );
  XNOR U7158 ( .A(n20052), .B(n7251), .Z(n7041) );
  OR U7159 ( .A(n7041), .B(n20020), .Z(n6950) );
  NANDN U7160 ( .A(n6948), .B(n19960), .Z(n6949) );
  NAND U7161 ( .A(n6950), .B(n6949), .Z(n7054) );
  XNOR U7162 ( .A(n102), .B(n6951), .Z(n7045) );
  OR U7163 ( .A(n7045), .B(n20121), .Z(n6954) );
  NANDN U7164 ( .A(n6952), .B(n20122), .Z(n6953) );
  NAND U7165 ( .A(n6954), .B(n6953), .Z(n7051) );
  XNOR U7166 ( .A(n19975), .B(n7407), .Z(n7048) );
  NANDN U7167 ( .A(n7048), .B(n19883), .Z(n6957) );
  NANDN U7168 ( .A(n6955), .B(n19937), .Z(n6956) );
  AND U7169 ( .A(n6957), .B(n6956), .Z(n7052) );
  XNOR U7170 ( .A(n7051), .B(n7052), .Z(n7053) );
  XNOR U7171 ( .A(n7054), .B(n7053), .Z(n7064) );
  XNOR U7172 ( .A(n7063), .B(n7064), .Z(n7065) );
  XNOR U7173 ( .A(n7066), .B(n7065), .Z(n7011) );
  NANDN U7174 ( .A(n6959), .B(n6958), .Z(n6963) );
  OR U7175 ( .A(n6961), .B(n6960), .Z(n6962) );
  NAND U7176 ( .A(n6963), .B(n6962), .Z(n7038) );
  XNOR U7177 ( .A(n20154), .B(n7095), .Z(n7023) );
  OR U7178 ( .A(n7023), .B(n20057), .Z(n6966) );
  NANDN U7179 ( .A(n6964), .B(n20098), .Z(n6965) );
  AND U7180 ( .A(n6966), .B(n6965), .Z(n7015) );
  NAND U7181 ( .A(b[0]), .B(a[96]), .Z(n6967) );
  XNOR U7182 ( .A(b[1]), .B(n6967), .Z(n6969) );
  NAND U7183 ( .A(a[95]), .B(n98), .Z(n6968) );
  AND U7184 ( .A(n6969), .B(n6968), .Z(n7014) );
  XOR U7185 ( .A(n7015), .B(n7014), .Z(n7017) );
  NAND U7186 ( .A(a[80]), .B(b[15]), .Z(n7016) );
  XOR U7187 ( .A(n7017), .B(n7016), .Z(n7035) );
  NAND U7188 ( .A(n19722), .B(n6970), .Z(n6972) );
  XNOR U7189 ( .A(b[5]), .B(n7731), .Z(n7026) );
  NANDN U7190 ( .A(n19640), .B(n7026), .Z(n6971) );
  NAND U7191 ( .A(n6972), .B(n6971), .Z(n7060) );
  XNOR U7192 ( .A(n19714), .B(n7563), .Z(n7029) );
  NANDN U7193 ( .A(n7029), .B(n19766), .Z(n6975) );
  NANDN U7194 ( .A(n6973), .B(n19767), .Z(n6974) );
  NAND U7195 ( .A(n6975), .B(n6974), .Z(n7057) );
  NAND U7196 ( .A(n19554), .B(n6976), .Z(n6978) );
  IV U7197 ( .A(a[94]), .Z(n7875) );
  XNOR U7198 ( .A(b[3]), .B(n7875), .Z(n7032) );
  NANDN U7199 ( .A(n19521), .B(n7032), .Z(n6977) );
  AND U7200 ( .A(n6978), .B(n6977), .Z(n7058) );
  XNOR U7201 ( .A(n7057), .B(n7058), .Z(n7059) );
  XOR U7202 ( .A(n7060), .B(n7059), .Z(n7036) );
  XOR U7203 ( .A(n7035), .B(n7036), .Z(n7037) );
  XNOR U7204 ( .A(n7038), .B(n7037), .Z(n7008) );
  NAND U7205 ( .A(n6980), .B(n6979), .Z(n6984) );
  NAND U7206 ( .A(n6982), .B(n6981), .Z(n6983) );
  NAND U7207 ( .A(n6984), .B(n6983), .Z(n7009) );
  XNOR U7208 ( .A(n7008), .B(n7009), .Z(n7010) );
  XOR U7209 ( .A(n7011), .B(n7010), .Z(n7069) );
  NANDN U7210 ( .A(n6986), .B(n6985), .Z(n6990) );
  NAND U7211 ( .A(n6988), .B(n6987), .Z(n6989) );
  NAND U7212 ( .A(n6990), .B(n6989), .Z(n7070) );
  XOR U7213 ( .A(n7069), .B(n7070), .Z(n7071) );
  XOR U7214 ( .A(n7072), .B(n7071), .Z(n7002) );
  NANDN U7215 ( .A(n6992), .B(n6991), .Z(n6996) );
  NANDN U7216 ( .A(n6994), .B(n6993), .Z(n6995) );
  NAND U7217 ( .A(n6996), .B(n6995), .Z(n7003) );
  XNOR U7218 ( .A(n7002), .B(n7003), .Z(n7004) );
  XNOR U7219 ( .A(n7005), .B(n7004), .Z(n7075) );
  XNOR U7220 ( .A(n7075), .B(sreg[336]), .Z(n7077) );
  NAND U7221 ( .A(n6997), .B(sreg[335]), .Z(n7001) );
  OR U7222 ( .A(n6999), .B(n6998), .Z(n7000) );
  AND U7223 ( .A(n7001), .B(n7000), .Z(n7076) );
  XOR U7224 ( .A(n7077), .B(n7076), .Z(c[336]) );
  NANDN U7225 ( .A(n7003), .B(n7002), .Z(n7007) );
  NAND U7226 ( .A(n7005), .B(n7004), .Z(n7006) );
  NAND U7227 ( .A(n7007), .B(n7006), .Z(n7083) );
  NANDN U7228 ( .A(n7009), .B(n7008), .Z(n7013) );
  NAND U7229 ( .A(n7011), .B(n7010), .Z(n7012) );
  NAND U7230 ( .A(n7013), .B(n7012), .Z(n7150) );
  NANDN U7231 ( .A(n7015), .B(n7014), .Z(n7019) );
  OR U7232 ( .A(n7017), .B(n7016), .Z(n7018) );
  NAND U7233 ( .A(n7019), .B(n7018), .Z(n7138) );
  NAND U7234 ( .A(b[0]), .B(a[97]), .Z(n7020) );
  XNOR U7235 ( .A(b[1]), .B(n7020), .Z(n7022) );
  NAND U7236 ( .A(a[96]), .B(n98), .Z(n7021) );
  AND U7237 ( .A(n7022), .B(n7021), .Z(n7114) );
  XNOR U7238 ( .A(n20154), .B(n7173), .Z(n7123) );
  OR U7239 ( .A(n7123), .B(n20057), .Z(n7025) );
  NANDN U7240 ( .A(n7023), .B(n20098), .Z(n7024) );
  AND U7241 ( .A(n7025), .B(n7024), .Z(n7115) );
  XOR U7242 ( .A(n7114), .B(n7115), .Z(n7117) );
  NAND U7243 ( .A(a[81]), .B(b[15]), .Z(n7116) );
  XOR U7244 ( .A(n7117), .B(n7116), .Z(n7135) );
  NAND U7245 ( .A(n19722), .B(n7026), .Z(n7028) );
  XNOR U7246 ( .A(b[5]), .B(n7797), .Z(n7126) );
  NANDN U7247 ( .A(n19640), .B(n7126), .Z(n7027) );
  NAND U7248 ( .A(n7028), .B(n7027), .Z(n7111) );
  XNOR U7249 ( .A(n19714), .B(n7641), .Z(n7129) );
  NANDN U7250 ( .A(n7129), .B(n19766), .Z(n7031) );
  NANDN U7251 ( .A(n7029), .B(n19767), .Z(n7030) );
  NAND U7252 ( .A(n7031), .B(n7030), .Z(n7108) );
  NAND U7253 ( .A(n19554), .B(n7032), .Z(n7034) );
  IV U7254 ( .A(a[95]), .Z(n7980) );
  XNOR U7255 ( .A(b[3]), .B(n7980), .Z(n7132) );
  NANDN U7256 ( .A(n19521), .B(n7132), .Z(n7033) );
  AND U7257 ( .A(n7034), .B(n7033), .Z(n7109) );
  XNOR U7258 ( .A(n7108), .B(n7109), .Z(n7110) );
  XOR U7259 ( .A(n7111), .B(n7110), .Z(n7136) );
  XOR U7260 ( .A(n7135), .B(n7136), .Z(n7137) );
  XNOR U7261 ( .A(n7138), .B(n7137), .Z(n7086) );
  NAND U7262 ( .A(n7036), .B(n7035), .Z(n7040) );
  NAND U7263 ( .A(n7038), .B(n7037), .Z(n7039) );
  NAND U7264 ( .A(n7040), .B(n7039), .Z(n7087) );
  XOR U7265 ( .A(n7086), .B(n7087), .Z(n7089) );
  XNOR U7266 ( .A(n20052), .B(n7329), .Z(n7092) );
  OR U7267 ( .A(n7092), .B(n20020), .Z(n7043) );
  NANDN U7268 ( .A(n7041), .B(n19960), .Z(n7042) );
  NAND U7269 ( .A(n7043), .B(n7042), .Z(n7105) );
  XNOR U7270 ( .A(n102), .B(n7044), .Z(n7096) );
  OR U7271 ( .A(n7096), .B(n20121), .Z(n7047) );
  NANDN U7272 ( .A(n7045), .B(n20122), .Z(n7046) );
  NAND U7273 ( .A(n7047), .B(n7046), .Z(n7102) );
  XNOR U7274 ( .A(n19975), .B(n7485), .Z(n7099) );
  NANDN U7275 ( .A(n7099), .B(n19883), .Z(n7050) );
  NANDN U7276 ( .A(n7048), .B(n19937), .Z(n7049) );
  AND U7277 ( .A(n7050), .B(n7049), .Z(n7103) );
  XNOR U7278 ( .A(n7102), .B(n7103), .Z(n7104) );
  XNOR U7279 ( .A(n7105), .B(n7104), .Z(n7141) );
  NANDN U7280 ( .A(n7052), .B(n7051), .Z(n7056) );
  NAND U7281 ( .A(n7054), .B(n7053), .Z(n7055) );
  NAND U7282 ( .A(n7056), .B(n7055), .Z(n7142) );
  XNOR U7283 ( .A(n7141), .B(n7142), .Z(n7143) );
  NANDN U7284 ( .A(n7058), .B(n7057), .Z(n7062) );
  NAND U7285 ( .A(n7060), .B(n7059), .Z(n7061) );
  AND U7286 ( .A(n7062), .B(n7061), .Z(n7144) );
  XNOR U7287 ( .A(n7143), .B(n7144), .Z(n7088) );
  XNOR U7288 ( .A(n7089), .B(n7088), .Z(n7147) );
  NANDN U7289 ( .A(n7064), .B(n7063), .Z(n7068) );
  NAND U7290 ( .A(n7066), .B(n7065), .Z(n7067) );
  AND U7291 ( .A(n7068), .B(n7067), .Z(n7148) );
  XNOR U7292 ( .A(n7147), .B(n7148), .Z(n7149) );
  XOR U7293 ( .A(n7150), .B(n7149), .Z(n7080) );
  OR U7294 ( .A(n7070), .B(n7069), .Z(n7074) );
  NANDN U7295 ( .A(n7072), .B(n7071), .Z(n7073) );
  NAND U7296 ( .A(n7074), .B(n7073), .Z(n7081) );
  XNOR U7297 ( .A(n7080), .B(n7081), .Z(n7082) );
  XNOR U7298 ( .A(n7083), .B(n7082), .Z(n7153) );
  XNOR U7299 ( .A(n7153), .B(sreg[337]), .Z(n7155) );
  NAND U7300 ( .A(n7075), .B(sreg[336]), .Z(n7079) );
  OR U7301 ( .A(n7077), .B(n7076), .Z(n7078) );
  AND U7302 ( .A(n7079), .B(n7078), .Z(n7154) );
  XOR U7303 ( .A(n7155), .B(n7154), .Z(c[337]) );
  NANDN U7304 ( .A(n7081), .B(n7080), .Z(n7085) );
  NAND U7305 ( .A(n7083), .B(n7082), .Z(n7084) );
  NAND U7306 ( .A(n7085), .B(n7084), .Z(n7161) );
  NANDN U7307 ( .A(n7087), .B(n7086), .Z(n7091) );
  OR U7308 ( .A(n7089), .B(n7088), .Z(n7090) );
  NAND U7309 ( .A(n7091), .B(n7090), .Z(n7228) );
  XNOR U7310 ( .A(n20052), .B(n7407), .Z(n7170) );
  OR U7311 ( .A(n7170), .B(n20020), .Z(n7094) );
  NANDN U7312 ( .A(n7092), .B(n19960), .Z(n7093) );
  NAND U7313 ( .A(n7094), .B(n7093), .Z(n7183) );
  XNOR U7314 ( .A(n102), .B(n7095), .Z(n7174) );
  OR U7315 ( .A(n7174), .B(n20121), .Z(n7098) );
  NANDN U7316 ( .A(n7096), .B(n20122), .Z(n7097) );
  NAND U7317 ( .A(n7098), .B(n7097), .Z(n7180) );
  XNOR U7318 ( .A(n19975), .B(n7563), .Z(n7177) );
  NANDN U7319 ( .A(n7177), .B(n19883), .Z(n7101) );
  NANDN U7320 ( .A(n7099), .B(n19937), .Z(n7100) );
  AND U7321 ( .A(n7101), .B(n7100), .Z(n7181) );
  XNOR U7322 ( .A(n7180), .B(n7181), .Z(n7182) );
  XNOR U7323 ( .A(n7183), .B(n7182), .Z(n7219) );
  NANDN U7324 ( .A(n7103), .B(n7102), .Z(n7107) );
  NAND U7325 ( .A(n7105), .B(n7104), .Z(n7106) );
  NAND U7326 ( .A(n7107), .B(n7106), .Z(n7220) );
  XNOR U7327 ( .A(n7219), .B(n7220), .Z(n7221) );
  NANDN U7328 ( .A(n7109), .B(n7108), .Z(n7113) );
  NAND U7329 ( .A(n7111), .B(n7110), .Z(n7112) );
  AND U7330 ( .A(n7113), .B(n7112), .Z(n7222) );
  XNOR U7331 ( .A(n7221), .B(n7222), .Z(n7166) );
  NANDN U7332 ( .A(n7115), .B(n7114), .Z(n7119) );
  OR U7333 ( .A(n7117), .B(n7116), .Z(n7118) );
  NAND U7334 ( .A(n7119), .B(n7118), .Z(n7216) );
  NAND U7335 ( .A(b[0]), .B(a[98]), .Z(n7120) );
  XNOR U7336 ( .A(b[1]), .B(n7120), .Z(n7122) );
  NAND U7337 ( .A(a[97]), .B(n98), .Z(n7121) );
  AND U7338 ( .A(n7122), .B(n7121), .Z(n7192) );
  XNOR U7339 ( .A(n20154), .B(n7251), .Z(n7201) );
  OR U7340 ( .A(n7201), .B(n20057), .Z(n7125) );
  NANDN U7341 ( .A(n7123), .B(n20098), .Z(n7124) );
  AND U7342 ( .A(n7125), .B(n7124), .Z(n7193) );
  XOR U7343 ( .A(n7192), .B(n7193), .Z(n7195) );
  NAND U7344 ( .A(a[82]), .B(b[15]), .Z(n7194) );
  XOR U7345 ( .A(n7195), .B(n7194), .Z(n7213) );
  NAND U7346 ( .A(n19722), .B(n7126), .Z(n7128) );
  XNOR U7347 ( .A(b[5]), .B(n7875), .Z(n7204) );
  NANDN U7348 ( .A(n19640), .B(n7204), .Z(n7127) );
  NAND U7349 ( .A(n7128), .B(n7127), .Z(n7189) );
  XNOR U7350 ( .A(n19714), .B(n7731), .Z(n7207) );
  NANDN U7351 ( .A(n7207), .B(n19766), .Z(n7131) );
  NANDN U7352 ( .A(n7129), .B(n19767), .Z(n7130) );
  NAND U7353 ( .A(n7131), .B(n7130), .Z(n7186) );
  NAND U7354 ( .A(n19554), .B(n7132), .Z(n7134) );
  IV U7355 ( .A(a[96]), .Z(n8031) );
  XNOR U7356 ( .A(b[3]), .B(n8031), .Z(n7210) );
  NANDN U7357 ( .A(n19521), .B(n7210), .Z(n7133) );
  AND U7358 ( .A(n7134), .B(n7133), .Z(n7187) );
  XNOR U7359 ( .A(n7186), .B(n7187), .Z(n7188) );
  XOR U7360 ( .A(n7189), .B(n7188), .Z(n7214) );
  XOR U7361 ( .A(n7213), .B(n7214), .Z(n7215) );
  XNOR U7362 ( .A(n7216), .B(n7215), .Z(n7164) );
  NAND U7363 ( .A(n7136), .B(n7135), .Z(n7140) );
  NAND U7364 ( .A(n7138), .B(n7137), .Z(n7139) );
  NAND U7365 ( .A(n7140), .B(n7139), .Z(n7165) );
  XOR U7366 ( .A(n7164), .B(n7165), .Z(n7167) );
  XNOR U7367 ( .A(n7166), .B(n7167), .Z(n7225) );
  NANDN U7368 ( .A(n7142), .B(n7141), .Z(n7146) );
  NAND U7369 ( .A(n7144), .B(n7143), .Z(n7145) );
  NAND U7370 ( .A(n7146), .B(n7145), .Z(n7226) );
  XNOR U7371 ( .A(n7225), .B(n7226), .Z(n7227) );
  XOR U7372 ( .A(n7228), .B(n7227), .Z(n7158) );
  NANDN U7373 ( .A(n7148), .B(n7147), .Z(n7152) );
  NANDN U7374 ( .A(n7150), .B(n7149), .Z(n7151) );
  NAND U7375 ( .A(n7152), .B(n7151), .Z(n7159) );
  XNOR U7376 ( .A(n7158), .B(n7159), .Z(n7160) );
  XNOR U7377 ( .A(n7161), .B(n7160), .Z(n7231) );
  XNOR U7378 ( .A(n7231), .B(sreg[338]), .Z(n7233) );
  NAND U7379 ( .A(n7153), .B(sreg[337]), .Z(n7157) );
  OR U7380 ( .A(n7155), .B(n7154), .Z(n7156) );
  AND U7381 ( .A(n7157), .B(n7156), .Z(n7232) );
  XOR U7382 ( .A(n7233), .B(n7232), .Z(c[338]) );
  NANDN U7383 ( .A(n7159), .B(n7158), .Z(n7163) );
  NAND U7384 ( .A(n7161), .B(n7160), .Z(n7162) );
  NAND U7385 ( .A(n7163), .B(n7162), .Z(n7239) );
  NANDN U7386 ( .A(n7165), .B(n7164), .Z(n7169) );
  OR U7387 ( .A(n7167), .B(n7166), .Z(n7168) );
  NAND U7388 ( .A(n7169), .B(n7168), .Z(n7306) );
  XNOR U7389 ( .A(n20052), .B(n7485), .Z(n7248) );
  OR U7390 ( .A(n7248), .B(n20020), .Z(n7172) );
  NANDN U7391 ( .A(n7170), .B(n19960), .Z(n7171) );
  NAND U7392 ( .A(n7172), .B(n7171), .Z(n7261) );
  XNOR U7393 ( .A(n102), .B(n7173), .Z(n7252) );
  OR U7394 ( .A(n7252), .B(n20121), .Z(n7176) );
  NANDN U7395 ( .A(n7174), .B(n20122), .Z(n7175) );
  NAND U7396 ( .A(n7176), .B(n7175), .Z(n7258) );
  XNOR U7397 ( .A(n19975), .B(n7641), .Z(n7255) );
  NANDN U7398 ( .A(n7255), .B(n19883), .Z(n7179) );
  NANDN U7399 ( .A(n7177), .B(n19937), .Z(n7178) );
  AND U7400 ( .A(n7179), .B(n7178), .Z(n7259) );
  XNOR U7401 ( .A(n7258), .B(n7259), .Z(n7260) );
  XNOR U7402 ( .A(n7261), .B(n7260), .Z(n7297) );
  NANDN U7403 ( .A(n7181), .B(n7180), .Z(n7185) );
  NAND U7404 ( .A(n7183), .B(n7182), .Z(n7184) );
  NAND U7405 ( .A(n7185), .B(n7184), .Z(n7298) );
  XNOR U7406 ( .A(n7297), .B(n7298), .Z(n7299) );
  NANDN U7407 ( .A(n7187), .B(n7186), .Z(n7191) );
  NAND U7408 ( .A(n7189), .B(n7188), .Z(n7190) );
  AND U7409 ( .A(n7191), .B(n7190), .Z(n7300) );
  XNOR U7410 ( .A(n7299), .B(n7300), .Z(n7244) );
  NANDN U7411 ( .A(n7193), .B(n7192), .Z(n7197) );
  OR U7412 ( .A(n7195), .B(n7194), .Z(n7196) );
  NAND U7413 ( .A(n7197), .B(n7196), .Z(n7294) );
  NAND U7414 ( .A(b[0]), .B(a[99]), .Z(n7198) );
  XNOR U7415 ( .A(b[1]), .B(n7198), .Z(n7200) );
  NAND U7416 ( .A(a[98]), .B(n98), .Z(n7199) );
  AND U7417 ( .A(n7200), .B(n7199), .Z(n7270) );
  XNOR U7418 ( .A(n20154), .B(n7329), .Z(n7276) );
  OR U7419 ( .A(n7276), .B(n20057), .Z(n7203) );
  NANDN U7420 ( .A(n7201), .B(n20098), .Z(n7202) );
  AND U7421 ( .A(n7203), .B(n7202), .Z(n7271) );
  XOR U7422 ( .A(n7270), .B(n7271), .Z(n7273) );
  NAND U7423 ( .A(a[83]), .B(b[15]), .Z(n7272) );
  XOR U7424 ( .A(n7273), .B(n7272), .Z(n7291) );
  NAND U7425 ( .A(n19722), .B(n7204), .Z(n7206) );
  XNOR U7426 ( .A(b[5]), .B(n7980), .Z(n7282) );
  NANDN U7427 ( .A(n19640), .B(n7282), .Z(n7205) );
  NAND U7428 ( .A(n7206), .B(n7205), .Z(n7267) );
  XNOR U7429 ( .A(n19714), .B(n7797), .Z(n7285) );
  NANDN U7430 ( .A(n7285), .B(n19766), .Z(n7209) );
  NANDN U7431 ( .A(n7207), .B(n19767), .Z(n7208) );
  NAND U7432 ( .A(n7209), .B(n7208), .Z(n7264) );
  NAND U7433 ( .A(n19554), .B(n7210), .Z(n7212) );
  IV U7434 ( .A(a[97]), .Z(n8136) );
  XNOR U7435 ( .A(b[3]), .B(n8136), .Z(n7288) );
  NANDN U7436 ( .A(n19521), .B(n7288), .Z(n7211) );
  AND U7437 ( .A(n7212), .B(n7211), .Z(n7265) );
  XNOR U7438 ( .A(n7264), .B(n7265), .Z(n7266) );
  XOR U7439 ( .A(n7267), .B(n7266), .Z(n7292) );
  XOR U7440 ( .A(n7291), .B(n7292), .Z(n7293) );
  XNOR U7441 ( .A(n7294), .B(n7293), .Z(n7242) );
  NAND U7442 ( .A(n7214), .B(n7213), .Z(n7218) );
  NAND U7443 ( .A(n7216), .B(n7215), .Z(n7217) );
  NAND U7444 ( .A(n7218), .B(n7217), .Z(n7243) );
  XOR U7445 ( .A(n7242), .B(n7243), .Z(n7245) );
  XNOR U7446 ( .A(n7244), .B(n7245), .Z(n7303) );
  NANDN U7447 ( .A(n7220), .B(n7219), .Z(n7224) );
  NAND U7448 ( .A(n7222), .B(n7221), .Z(n7223) );
  NAND U7449 ( .A(n7224), .B(n7223), .Z(n7304) );
  XNOR U7450 ( .A(n7303), .B(n7304), .Z(n7305) );
  XOR U7451 ( .A(n7306), .B(n7305), .Z(n7236) );
  NANDN U7452 ( .A(n7226), .B(n7225), .Z(n7230) );
  NANDN U7453 ( .A(n7228), .B(n7227), .Z(n7229) );
  NAND U7454 ( .A(n7230), .B(n7229), .Z(n7237) );
  XNOR U7455 ( .A(n7236), .B(n7237), .Z(n7238) );
  XNOR U7456 ( .A(n7239), .B(n7238), .Z(n7309) );
  XNOR U7457 ( .A(n7309), .B(sreg[339]), .Z(n7311) );
  NAND U7458 ( .A(n7231), .B(sreg[338]), .Z(n7235) );
  OR U7459 ( .A(n7233), .B(n7232), .Z(n7234) );
  AND U7460 ( .A(n7235), .B(n7234), .Z(n7310) );
  XOR U7461 ( .A(n7311), .B(n7310), .Z(c[339]) );
  NANDN U7462 ( .A(n7237), .B(n7236), .Z(n7241) );
  NAND U7463 ( .A(n7239), .B(n7238), .Z(n7240) );
  NAND U7464 ( .A(n7241), .B(n7240), .Z(n7317) );
  NANDN U7465 ( .A(n7243), .B(n7242), .Z(n7247) );
  OR U7466 ( .A(n7245), .B(n7244), .Z(n7246) );
  NAND U7467 ( .A(n7247), .B(n7246), .Z(n7384) );
  XNOR U7468 ( .A(n20052), .B(n7563), .Z(n7326) );
  OR U7469 ( .A(n7326), .B(n20020), .Z(n7250) );
  NANDN U7470 ( .A(n7248), .B(n19960), .Z(n7249) );
  NAND U7471 ( .A(n7250), .B(n7249), .Z(n7339) );
  XNOR U7472 ( .A(n102), .B(n7251), .Z(n7330) );
  OR U7473 ( .A(n7330), .B(n20121), .Z(n7254) );
  NANDN U7474 ( .A(n7252), .B(n20122), .Z(n7253) );
  NAND U7475 ( .A(n7254), .B(n7253), .Z(n7336) );
  XNOR U7476 ( .A(n19975), .B(n7731), .Z(n7333) );
  NANDN U7477 ( .A(n7333), .B(n19883), .Z(n7257) );
  NANDN U7478 ( .A(n7255), .B(n19937), .Z(n7256) );
  AND U7479 ( .A(n7257), .B(n7256), .Z(n7337) );
  XNOR U7480 ( .A(n7336), .B(n7337), .Z(n7338) );
  XNOR U7481 ( .A(n7339), .B(n7338), .Z(n7375) );
  NANDN U7482 ( .A(n7259), .B(n7258), .Z(n7263) );
  NAND U7483 ( .A(n7261), .B(n7260), .Z(n7262) );
  NAND U7484 ( .A(n7263), .B(n7262), .Z(n7376) );
  XNOR U7485 ( .A(n7375), .B(n7376), .Z(n7377) );
  NANDN U7486 ( .A(n7265), .B(n7264), .Z(n7269) );
  NAND U7487 ( .A(n7267), .B(n7266), .Z(n7268) );
  AND U7488 ( .A(n7269), .B(n7268), .Z(n7378) );
  XNOR U7489 ( .A(n7377), .B(n7378), .Z(n7322) );
  NANDN U7490 ( .A(n7271), .B(n7270), .Z(n7275) );
  OR U7491 ( .A(n7273), .B(n7272), .Z(n7274) );
  NAND U7492 ( .A(n7275), .B(n7274), .Z(n7372) );
  XNOR U7493 ( .A(n20154), .B(n7407), .Z(n7354) );
  OR U7494 ( .A(n7354), .B(n20057), .Z(n7278) );
  NANDN U7495 ( .A(n7276), .B(n20098), .Z(n7277) );
  AND U7496 ( .A(n7278), .B(n7277), .Z(n7349) );
  NAND U7497 ( .A(b[0]), .B(a[100]), .Z(n7279) );
  XNOR U7498 ( .A(b[1]), .B(n7279), .Z(n7281) );
  NAND U7499 ( .A(a[99]), .B(n98), .Z(n7280) );
  AND U7500 ( .A(n7281), .B(n7280), .Z(n7348) );
  XOR U7501 ( .A(n7349), .B(n7348), .Z(n7351) );
  NAND U7502 ( .A(a[84]), .B(b[15]), .Z(n7350) );
  XOR U7503 ( .A(n7351), .B(n7350), .Z(n7369) );
  NAND U7504 ( .A(n19722), .B(n7282), .Z(n7284) );
  XNOR U7505 ( .A(b[5]), .B(n8031), .Z(n7360) );
  NANDN U7506 ( .A(n19640), .B(n7360), .Z(n7283) );
  NAND U7507 ( .A(n7284), .B(n7283), .Z(n7345) );
  XNOR U7508 ( .A(n19714), .B(n7875), .Z(n7363) );
  NANDN U7509 ( .A(n7363), .B(n19766), .Z(n7287) );
  NANDN U7510 ( .A(n7285), .B(n19767), .Z(n7286) );
  NAND U7511 ( .A(n7287), .B(n7286), .Z(n7342) );
  NAND U7512 ( .A(n19554), .B(n7288), .Z(n7290) );
  IV U7513 ( .A(a[98]), .Z(n8214) );
  XNOR U7514 ( .A(b[3]), .B(n8214), .Z(n7366) );
  NANDN U7515 ( .A(n19521), .B(n7366), .Z(n7289) );
  AND U7516 ( .A(n7290), .B(n7289), .Z(n7343) );
  XNOR U7517 ( .A(n7342), .B(n7343), .Z(n7344) );
  XOR U7518 ( .A(n7345), .B(n7344), .Z(n7370) );
  XOR U7519 ( .A(n7369), .B(n7370), .Z(n7371) );
  XNOR U7520 ( .A(n7372), .B(n7371), .Z(n7320) );
  NAND U7521 ( .A(n7292), .B(n7291), .Z(n7296) );
  NAND U7522 ( .A(n7294), .B(n7293), .Z(n7295) );
  NAND U7523 ( .A(n7296), .B(n7295), .Z(n7321) );
  XOR U7524 ( .A(n7320), .B(n7321), .Z(n7323) );
  XNOR U7525 ( .A(n7322), .B(n7323), .Z(n7381) );
  NANDN U7526 ( .A(n7298), .B(n7297), .Z(n7302) );
  NAND U7527 ( .A(n7300), .B(n7299), .Z(n7301) );
  NAND U7528 ( .A(n7302), .B(n7301), .Z(n7382) );
  XNOR U7529 ( .A(n7381), .B(n7382), .Z(n7383) );
  XOR U7530 ( .A(n7384), .B(n7383), .Z(n7314) );
  NANDN U7531 ( .A(n7304), .B(n7303), .Z(n7308) );
  NANDN U7532 ( .A(n7306), .B(n7305), .Z(n7307) );
  NAND U7533 ( .A(n7308), .B(n7307), .Z(n7315) );
  XNOR U7534 ( .A(n7314), .B(n7315), .Z(n7316) );
  XNOR U7535 ( .A(n7317), .B(n7316), .Z(n7387) );
  XNOR U7536 ( .A(n7387), .B(sreg[340]), .Z(n7389) );
  NAND U7537 ( .A(n7309), .B(sreg[339]), .Z(n7313) );
  OR U7538 ( .A(n7311), .B(n7310), .Z(n7312) );
  AND U7539 ( .A(n7313), .B(n7312), .Z(n7388) );
  XOR U7540 ( .A(n7389), .B(n7388), .Z(c[340]) );
  NANDN U7541 ( .A(n7315), .B(n7314), .Z(n7319) );
  NAND U7542 ( .A(n7317), .B(n7316), .Z(n7318) );
  NAND U7543 ( .A(n7319), .B(n7318), .Z(n7395) );
  NANDN U7544 ( .A(n7321), .B(n7320), .Z(n7325) );
  OR U7545 ( .A(n7323), .B(n7322), .Z(n7324) );
  NAND U7546 ( .A(n7325), .B(n7324), .Z(n7462) );
  XNOR U7547 ( .A(n20052), .B(n7641), .Z(n7404) );
  OR U7548 ( .A(n7404), .B(n20020), .Z(n7328) );
  NANDN U7549 ( .A(n7326), .B(n19960), .Z(n7327) );
  NAND U7550 ( .A(n7328), .B(n7327), .Z(n7417) );
  XNOR U7551 ( .A(n102), .B(n7329), .Z(n7408) );
  OR U7552 ( .A(n7408), .B(n20121), .Z(n7332) );
  NANDN U7553 ( .A(n7330), .B(n20122), .Z(n7331) );
  NAND U7554 ( .A(n7332), .B(n7331), .Z(n7414) );
  XNOR U7555 ( .A(n19975), .B(n7797), .Z(n7411) );
  NANDN U7556 ( .A(n7411), .B(n19883), .Z(n7335) );
  NANDN U7557 ( .A(n7333), .B(n19937), .Z(n7334) );
  AND U7558 ( .A(n7335), .B(n7334), .Z(n7415) );
  XNOR U7559 ( .A(n7414), .B(n7415), .Z(n7416) );
  XNOR U7560 ( .A(n7417), .B(n7416), .Z(n7453) );
  NANDN U7561 ( .A(n7337), .B(n7336), .Z(n7341) );
  NAND U7562 ( .A(n7339), .B(n7338), .Z(n7340) );
  NAND U7563 ( .A(n7341), .B(n7340), .Z(n7454) );
  XNOR U7564 ( .A(n7453), .B(n7454), .Z(n7455) );
  NANDN U7565 ( .A(n7343), .B(n7342), .Z(n7347) );
  NAND U7566 ( .A(n7345), .B(n7344), .Z(n7346) );
  AND U7567 ( .A(n7347), .B(n7346), .Z(n7456) );
  XNOR U7568 ( .A(n7455), .B(n7456), .Z(n7400) );
  NANDN U7569 ( .A(n7349), .B(n7348), .Z(n7353) );
  OR U7570 ( .A(n7351), .B(n7350), .Z(n7352) );
  NAND U7571 ( .A(n7353), .B(n7352), .Z(n7450) );
  XNOR U7572 ( .A(n20154), .B(n7485), .Z(n7435) );
  OR U7573 ( .A(n7435), .B(n20057), .Z(n7356) );
  NANDN U7574 ( .A(n7354), .B(n20098), .Z(n7355) );
  AND U7575 ( .A(n7356), .B(n7355), .Z(n7427) );
  NAND U7576 ( .A(b[0]), .B(a[101]), .Z(n7357) );
  XNOR U7577 ( .A(b[1]), .B(n7357), .Z(n7359) );
  NAND U7578 ( .A(a[100]), .B(n98), .Z(n7358) );
  AND U7579 ( .A(n7359), .B(n7358), .Z(n7426) );
  XOR U7580 ( .A(n7427), .B(n7426), .Z(n7429) );
  NAND U7581 ( .A(a[85]), .B(b[15]), .Z(n7428) );
  XOR U7582 ( .A(n7429), .B(n7428), .Z(n7447) );
  NAND U7583 ( .A(n19722), .B(n7360), .Z(n7362) );
  XNOR U7584 ( .A(b[5]), .B(n8136), .Z(n7438) );
  NANDN U7585 ( .A(n19640), .B(n7438), .Z(n7361) );
  NAND U7586 ( .A(n7362), .B(n7361), .Z(n7423) );
  XNOR U7587 ( .A(n19714), .B(n7980), .Z(n7441) );
  NANDN U7588 ( .A(n7441), .B(n19766), .Z(n7365) );
  NANDN U7589 ( .A(n7363), .B(n19767), .Z(n7364) );
  NAND U7590 ( .A(n7365), .B(n7364), .Z(n7420) );
  NAND U7591 ( .A(n19554), .B(n7366), .Z(n7368) );
  IV U7592 ( .A(a[99]), .Z(n8265) );
  XNOR U7593 ( .A(b[3]), .B(n8265), .Z(n7444) );
  NANDN U7594 ( .A(n19521), .B(n7444), .Z(n7367) );
  AND U7595 ( .A(n7368), .B(n7367), .Z(n7421) );
  XNOR U7596 ( .A(n7420), .B(n7421), .Z(n7422) );
  XOR U7597 ( .A(n7423), .B(n7422), .Z(n7448) );
  XOR U7598 ( .A(n7447), .B(n7448), .Z(n7449) );
  XNOR U7599 ( .A(n7450), .B(n7449), .Z(n7398) );
  NAND U7600 ( .A(n7370), .B(n7369), .Z(n7374) );
  NAND U7601 ( .A(n7372), .B(n7371), .Z(n7373) );
  NAND U7602 ( .A(n7374), .B(n7373), .Z(n7399) );
  XOR U7603 ( .A(n7398), .B(n7399), .Z(n7401) );
  XNOR U7604 ( .A(n7400), .B(n7401), .Z(n7459) );
  NANDN U7605 ( .A(n7376), .B(n7375), .Z(n7380) );
  NAND U7606 ( .A(n7378), .B(n7377), .Z(n7379) );
  NAND U7607 ( .A(n7380), .B(n7379), .Z(n7460) );
  XNOR U7608 ( .A(n7459), .B(n7460), .Z(n7461) );
  XOR U7609 ( .A(n7462), .B(n7461), .Z(n7392) );
  NANDN U7610 ( .A(n7382), .B(n7381), .Z(n7386) );
  NANDN U7611 ( .A(n7384), .B(n7383), .Z(n7385) );
  NAND U7612 ( .A(n7386), .B(n7385), .Z(n7393) );
  XNOR U7613 ( .A(n7392), .B(n7393), .Z(n7394) );
  XNOR U7614 ( .A(n7395), .B(n7394), .Z(n7465) );
  XNOR U7615 ( .A(n7465), .B(sreg[341]), .Z(n7467) );
  NAND U7616 ( .A(n7387), .B(sreg[340]), .Z(n7391) );
  OR U7617 ( .A(n7389), .B(n7388), .Z(n7390) );
  AND U7618 ( .A(n7391), .B(n7390), .Z(n7466) );
  XOR U7619 ( .A(n7467), .B(n7466), .Z(c[341]) );
  NANDN U7620 ( .A(n7393), .B(n7392), .Z(n7397) );
  NAND U7621 ( .A(n7395), .B(n7394), .Z(n7396) );
  NAND U7622 ( .A(n7397), .B(n7396), .Z(n7473) );
  NANDN U7623 ( .A(n7399), .B(n7398), .Z(n7403) );
  OR U7624 ( .A(n7401), .B(n7400), .Z(n7402) );
  NAND U7625 ( .A(n7403), .B(n7402), .Z(n7540) );
  XNOR U7626 ( .A(n20052), .B(n7731), .Z(n7482) );
  OR U7627 ( .A(n7482), .B(n20020), .Z(n7406) );
  NANDN U7628 ( .A(n7404), .B(n19960), .Z(n7405) );
  NAND U7629 ( .A(n7406), .B(n7405), .Z(n7495) );
  XNOR U7630 ( .A(n102), .B(n7407), .Z(n7486) );
  OR U7631 ( .A(n7486), .B(n20121), .Z(n7410) );
  NANDN U7632 ( .A(n7408), .B(n20122), .Z(n7409) );
  NAND U7633 ( .A(n7410), .B(n7409), .Z(n7492) );
  XNOR U7634 ( .A(n19975), .B(n7875), .Z(n7489) );
  NANDN U7635 ( .A(n7489), .B(n19883), .Z(n7413) );
  NANDN U7636 ( .A(n7411), .B(n19937), .Z(n7412) );
  AND U7637 ( .A(n7413), .B(n7412), .Z(n7493) );
  XNOR U7638 ( .A(n7492), .B(n7493), .Z(n7494) );
  XNOR U7639 ( .A(n7495), .B(n7494), .Z(n7531) );
  NANDN U7640 ( .A(n7415), .B(n7414), .Z(n7419) );
  NAND U7641 ( .A(n7417), .B(n7416), .Z(n7418) );
  NAND U7642 ( .A(n7419), .B(n7418), .Z(n7532) );
  XNOR U7643 ( .A(n7531), .B(n7532), .Z(n7533) );
  NANDN U7644 ( .A(n7421), .B(n7420), .Z(n7425) );
  NAND U7645 ( .A(n7423), .B(n7422), .Z(n7424) );
  AND U7646 ( .A(n7425), .B(n7424), .Z(n7534) );
  XNOR U7647 ( .A(n7533), .B(n7534), .Z(n7478) );
  NANDN U7648 ( .A(n7427), .B(n7426), .Z(n7431) );
  OR U7649 ( .A(n7429), .B(n7428), .Z(n7430) );
  NAND U7650 ( .A(n7431), .B(n7430), .Z(n7528) );
  NAND U7651 ( .A(b[0]), .B(a[102]), .Z(n7432) );
  XNOR U7652 ( .A(b[1]), .B(n7432), .Z(n7434) );
  NAND U7653 ( .A(a[101]), .B(n98), .Z(n7433) );
  AND U7654 ( .A(n7434), .B(n7433), .Z(n7504) );
  XNOR U7655 ( .A(n20154), .B(n7563), .Z(n7513) );
  OR U7656 ( .A(n7513), .B(n20057), .Z(n7437) );
  NANDN U7657 ( .A(n7435), .B(n20098), .Z(n7436) );
  AND U7658 ( .A(n7437), .B(n7436), .Z(n7505) );
  XOR U7659 ( .A(n7504), .B(n7505), .Z(n7507) );
  NAND U7660 ( .A(a[86]), .B(b[15]), .Z(n7506) );
  XOR U7661 ( .A(n7507), .B(n7506), .Z(n7525) );
  NAND U7662 ( .A(n19722), .B(n7438), .Z(n7440) );
  XNOR U7663 ( .A(b[5]), .B(n8214), .Z(n7516) );
  NANDN U7664 ( .A(n19640), .B(n7516), .Z(n7439) );
  NAND U7665 ( .A(n7440), .B(n7439), .Z(n7501) );
  XNOR U7666 ( .A(n19714), .B(n8031), .Z(n7519) );
  NANDN U7667 ( .A(n7519), .B(n19766), .Z(n7443) );
  NANDN U7668 ( .A(n7441), .B(n19767), .Z(n7442) );
  NAND U7669 ( .A(n7443), .B(n7442), .Z(n7498) );
  NAND U7670 ( .A(n19554), .B(n7444), .Z(n7446) );
  IV U7671 ( .A(a[100]), .Z(n8343) );
  XNOR U7672 ( .A(b[3]), .B(n8343), .Z(n7522) );
  NANDN U7673 ( .A(n19521), .B(n7522), .Z(n7445) );
  AND U7674 ( .A(n7446), .B(n7445), .Z(n7499) );
  XNOR U7675 ( .A(n7498), .B(n7499), .Z(n7500) );
  XOR U7676 ( .A(n7501), .B(n7500), .Z(n7526) );
  XOR U7677 ( .A(n7525), .B(n7526), .Z(n7527) );
  XNOR U7678 ( .A(n7528), .B(n7527), .Z(n7476) );
  NAND U7679 ( .A(n7448), .B(n7447), .Z(n7452) );
  NAND U7680 ( .A(n7450), .B(n7449), .Z(n7451) );
  NAND U7681 ( .A(n7452), .B(n7451), .Z(n7477) );
  XOR U7682 ( .A(n7476), .B(n7477), .Z(n7479) );
  XNOR U7683 ( .A(n7478), .B(n7479), .Z(n7537) );
  NANDN U7684 ( .A(n7454), .B(n7453), .Z(n7458) );
  NAND U7685 ( .A(n7456), .B(n7455), .Z(n7457) );
  NAND U7686 ( .A(n7458), .B(n7457), .Z(n7538) );
  XNOR U7687 ( .A(n7537), .B(n7538), .Z(n7539) );
  XOR U7688 ( .A(n7540), .B(n7539), .Z(n7470) );
  NANDN U7689 ( .A(n7460), .B(n7459), .Z(n7464) );
  NANDN U7690 ( .A(n7462), .B(n7461), .Z(n7463) );
  NAND U7691 ( .A(n7464), .B(n7463), .Z(n7471) );
  XNOR U7692 ( .A(n7470), .B(n7471), .Z(n7472) );
  XNOR U7693 ( .A(n7473), .B(n7472), .Z(n7543) );
  XNOR U7694 ( .A(n7543), .B(sreg[342]), .Z(n7545) );
  NAND U7695 ( .A(n7465), .B(sreg[341]), .Z(n7469) );
  OR U7696 ( .A(n7467), .B(n7466), .Z(n7468) );
  AND U7697 ( .A(n7469), .B(n7468), .Z(n7544) );
  XOR U7698 ( .A(n7545), .B(n7544), .Z(c[342]) );
  NANDN U7699 ( .A(n7471), .B(n7470), .Z(n7475) );
  NAND U7700 ( .A(n7473), .B(n7472), .Z(n7474) );
  NAND U7701 ( .A(n7475), .B(n7474), .Z(n7551) );
  NANDN U7702 ( .A(n7477), .B(n7476), .Z(n7481) );
  OR U7703 ( .A(n7479), .B(n7478), .Z(n7480) );
  NAND U7704 ( .A(n7481), .B(n7480), .Z(n7618) );
  XNOR U7705 ( .A(n20052), .B(n7797), .Z(n7560) );
  OR U7706 ( .A(n7560), .B(n20020), .Z(n7484) );
  NANDN U7707 ( .A(n7482), .B(n19960), .Z(n7483) );
  NAND U7708 ( .A(n7484), .B(n7483), .Z(n7573) );
  XNOR U7709 ( .A(n102), .B(n7485), .Z(n7564) );
  OR U7710 ( .A(n7564), .B(n20121), .Z(n7488) );
  NANDN U7711 ( .A(n7486), .B(n20122), .Z(n7487) );
  NAND U7712 ( .A(n7488), .B(n7487), .Z(n7570) );
  XNOR U7713 ( .A(n19975), .B(n7980), .Z(n7567) );
  NANDN U7714 ( .A(n7567), .B(n19883), .Z(n7491) );
  NANDN U7715 ( .A(n7489), .B(n19937), .Z(n7490) );
  AND U7716 ( .A(n7491), .B(n7490), .Z(n7571) );
  XNOR U7717 ( .A(n7570), .B(n7571), .Z(n7572) );
  XNOR U7718 ( .A(n7573), .B(n7572), .Z(n7609) );
  NANDN U7719 ( .A(n7493), .B(n7492), .Z(n7497) );
  NAND U7720 ( .A(n7495), .B(n7494), .Z(n7496) );
  NAND U7721 ( .A(n7497), .B(n7496), .Z(n7610) );
  XNOR U7722 ( .A(n7609), .B(n7610), .Z(n7611) );
  NANDN U7723 ( .A(n7499), .B(n7498), .Z(n7503) );
  NAND U7724 ( .A(n7501), .B(n7500), .Z(n7502) );
  AND U7725 ( .A(n7503), .B(n7502), .Z(n7612) );
  XNOR U7726 ( .A(n7611), .B(n7612), .Z(n7556) );
  NANDN U7727 ( .A(n7505), .B(n7504), .Z(n7509) );
  OR U7728 ( .A(n7507), .B(n7506), .Z(n7508) );
  NAND U7729 ( .A(n7509), .B(n7508), .Z(n7606) );
  NAND U7730 ( .A(b[0]), .B(a[103]), .Z(n7510) );
  XNOR U7731 ( .A(b[1]), .B(n7510), .Z(n7512) );
  NAND U7732 ( .A(a[102]), .B(n98), .Z(n7511) );
  AND U7733 ( .A(n7512), .B(n7511), .Z(n7582) );
  XNOR U7734 ( .A(n20154), .B(n7641), .Z(n7591) );
  OR U7735 ( .A(n7591), .B(n20057), .Z(n7515) );
  NANDN U7736 ( .A(n7513), .B(n20098), .Z(n7514) );
  AND U7737 ( .A(n7515), .B(n7514), .Z(n7583) );
  XOR U7738 ( .A(n7582), .B(n7583), .Z(n7585) );
  NAND U7739 ( .A(a[87]), .B(b[15]), .Z(n7584) );
  XOR U7740 ( .A(n7585), .B(n7584), .Z(n7603) );
  NAND U7741 ( .A(n19722), .B(n7516), .Z(n7518) );
  XNOR U7742 ( .A(b[5]), .B(n8265), .Z(n7594) );
  NANDN U7743 ( .A(n19640), .B(n7594), .Z(n7517) );
  NAND U7744 ( .A(n7518), .B(n7517), .Z(n7579) );
  XNOR U7745 ( .A(n19714), .B(n8136), .Z(n7597) );
  NANDN U7746 ( .A(n7597), .B(n19766), .Z(n7521) );
  NANDN U7747 ( .A(n7519), .B(n19767), .Z(n7520) );
  NAND U7748 ( .A(n7521), .B(n7520), .Z(n7576) );
  NAND U7749 ( .A(n19554), .B(n7522), .Z(n7524) );
  IV U7750 ( .A(a[101]), .Z(n8448) );
  XNOR U7751 ( .A(b[3]), .B(n8448), .Z(n7600) );
  NANDN U7752 ( .A(n19521), .B(n7600), .Z(n7523) );
  AND U7753 ( .A(n7524), .B(n7523), .Z(n7577) );
  XNOR U7754 ( .A(n7576), .B(n7577), .Z(n7578) );
  XOR U7755 ( .A(n7579), .B(n7578), .Z(n7604) );
  XOR U7756 ( .A(n7603), .B(n7604), .Z(n7605) );
  XNOR U7757 ( .A(n7606), .B(n7605), .Z(n7554) );
  NAND U7758 ( .A(n7526), .B(n7525), .Z(n7530) );
  NAND U7759 ( .A(n7528), .B(n7527), .Z(n7529) );
  NAND U7760 ( .A(n7530), .B(n7529), .Z(n7555) );
  XOR U7761 ( .A(n7554), .B(n7555), .Z(n7557) );
  XNOR U7762 ( .A(n7556), .B(n7557), .Z(n7615) );
  NANDN U7763 ( .A(n7532), .B(n7531), .Z(n7536) );
  NAND U7764 ( .A(n7534), .B(n7533), .Z(n7535) );
  NAND U7765 ( .A(n7536), .B(n7535), .Z(n7616) );
  XNOR U7766 ( .A(n7615), .B(n7616), .Z(n7617) );
  XOR U7767 ( .A(n7618), .B(n7617), .Z(n7548) );
  NANDN U7768 ( .A(n7538), .B(n7537), .Z(n7542) );
  NANDN U7769 ( .A(n7540), .B(n7539), .Z(n7541) );
  NAND U7770 ( .A(n7542), .B(n7541), .Z(n7549) );
  XNOR U7771 ( .A(n7548), .B(n7549), .Z(n7550) );
  XNOR U7772 ( .A(n7551), .B(n7550), .Z(n7621) );
  XNOR U7773 ( .A(n7621), .B(sreg[343]), .Z(n7623) );
  NAND U7774 ( .A(n7543), .B(sreg[342]), .Z(n7547) );
  OR U7775 ( .A(n7545), .B(n7544), .Z(n7546) );
  AND U7776 ( .A(n7547), .B(n7546), .Z(n7622) );
  XOR U7777 ( .A(n7623), .B(n7622), .Z(c[343]) );
  NANDN U7778 ( .A(n7549), .B(n7548), .Z(n7553) );
  NAND U7779 ( .A(n7551), .B(n7550), .Z(n7552) );
  NAND U7780 ( .A(n7553), .B(n7552), .Z(n7629) );
  NANDN U7781 ( .A(n7555), .B(n7554), .Z(n7559) );
  OR U7782 ( .A(n7557), .B(n7556), .Z(n7558) );
  NAND U7783 ( .A(n7559), .B(n7558), .Z(n7696) );
  XNOR U7784 ( .A(n20052), .B(n7875), .Z(n7638) );
  OR U7785 ( .A(n7638), .B(n20020), .Z(n7562) );
  NANDN U7786 ( .A(n7560), .B(n19960), .Z(n7561) );
  NAND U7787 ( .A(n7562), .B(n7561), .Z(n7651) );
  XNOR U7788 ( .A(n102), .B(n7563), .Z(n7642) );
  OR U7789 ( .A(n7642), .B(n20121), .Z(n7566) );
  NANDN U7790 ( .A(n7564), .B(n20122), .Z(n7565) );
  NAND U7791 ( .A(n7566), .B(n7565), .Z(n7648) );
  XNOR U7792 ( .A(n19975), .B(n8031), .Z(n7645) );
  NANDN U7793 ( .A(n7645), .B(n19883), .Z(n7569) );
  NANDN U7794 ( .A(n7567), .B(n19937), .Z(n7568) );
  AND U7795 ( .A(n7569), .B(n7568), .Z(n7649) );
  XNOR U7796 ( .A(n7648), .B(n7649), .Z(n7650) );
  XNOR U7797 ( .A(n7651), .B(n7650), .Z(n7687) );
  NANDN U7798 ( .A(n7571), .B(n7570), .Z(n7575) );
  NAND U7799 ( .A(n7573), .B(n7572), .Z(n7574) );
  NAND U7800 ( .A(n7575), .B(n7574), .Z(n7688) );
  XNOR U7801 ( .A(n7687), .B(n7688), .Z(n7689) );
  NANDN U7802 ( .A(n7577), .B(n7576), .Z(n7581) );
  NAND U7803 ( .A(n7579), .B(n7578), .Z(n7580) );
  AND U7804 ( .A(n7581), .B(n7580), .Z(n7690) );
  XNOR U7805 ( .A(n7689), .B(n7690), .Z(n7634) );
  NANDN U7806 ( .A(n7583), .B(n7582), .Z(n7587) );
  OR U7807 ( .A(n7585), .B(n7584), .Z(n7586) );
  NAND U7808 ( .A(n7587), .B(n7586), .Z(n7684) );
  NAND U7809 ( .A(b[0]), .B(a[104]), .Z(n7588) );
  XNOR U7810 ( .A(b[1]), .B(n7588), .Z(n7590) );
  NAND U7811 ( .A(a[103]), .B(n98), .Z(n7589) );
  AND U7812 ( .A(n7590), .B(n7589), .Z(n7660) );
  XNOR U7813 ( .A(n20154), .B(n7731), .Z(n7669) );
  OR U7814 ( .A(n7669), .B(n20057), .Z(n7593) );
  NANDN U7815 ( .A(n7591), .B(n20098), .Z(n7592) );
  AND U7816 ( .A(n7593), .B(n7592), .Z(n7661) );
  XOR U7817 ( .A(n7660), .B(n7661), .Z(n7663) );
  NAND U7818 ( .A(a[88]), .B(b[15]), .Z(n7662) );
  XOR U7819 ( .A(n7663), .B(n7662), .Z(n7681) );
  NAND U7820 ( .A(n19722), .B(n7594), .Z(n7596) );
  XNOR U7821 ( .A(b[5]), .B(n8343), .Z(n7672) );
  NANDN U7822 ( .A(n19640), .B(n7672), .Z(n7595) );
  NAND U7823 ( .A(n7596), .B(n7595), .Z(n7657) );
  XNOR U7824 ( .A(n19714), .B(n8214), .Z(n7675) );
  NANDN U7825 ( .A(n7675), .B(n19766), .Z(n7599) );
  NANDN U7826 ( .A(n7597), .B(n19767), .Z(n7598) );
  NAND U7827 ( .A(n7599), .B(n7598), .Z(n7654) );
  NAND U7828 ( .A(n19554), .B(n7600), .Z(n7602) );
  IV U7829 ( .A(a[102]), .Z(n8499) );
  XNOR U7830 ( .A(b[3]), .B(n8499), .Z(n7678) );
  NANDN U7831 ( .A(n19521), .B(n7678), .Z(n7601) );
  AND U7832 ( .A(n7602), .B(n7601), .Z(n7655) );
  XNOR U7833 ( .A(n7654), .B(n7655), .Z(n7656) );
  XOR U7834 ( .A(n7657), .B(n7656), .Z(n7682) );
  XOR U7835 ( .A(n7681), .B(n7682), .Z(n7683) );
  XNOR U7836 ( .A(n7684), .B(n7683), .Z(n7632) );
  NAND U7837 ( .A(n7604), .B(n7603), .Z(n7608) );
  NAND U7838 ( .A(n7606), .B(n7605), .Z(n7607) );
  NAND U7839 ( .A(n7608), .B(n7607), .Z(n7633) );
  XOR U7840 ( .A(n7632), .B(n7633), .Z(n7635) );
  XNOR U7841 ( .A(n7634), .B(n7635), .Z(n7693) );
  NANDN U7842 ( .A(n7610), .B(n7609), .Z(n7614) );
  NAND U7843 ( .A(n7612), .B(n7611), .Z(n7613) );
  NAND U7844 ( .A(n7614), .B(n7613), .Z(n7694) );
  XNOR U7845 ( .A(n7693), .B(n7694), .Z(n7695) );
  XOR U7846 ( .A(n7696), .B(n7695), .Z(n7626) );
  NANDN U7847 ( .A(n7616), .B(n7615), .Z(n7620) );
  NANDN U7848 ( .A(n7618), .B(n7617), .Z(n7619) );
  NAND U7849 ( .A(n7620), .B(n7619), .Z(n7627) );
  XNOR U7850 ( .A(n7626), .B(n7627), .Z(n7628) );
  XNOR U7851 ( .A(n7629), .B(n7628), .Z(n7699) );
  XNOR U7852 ( .A(n7699), .B(sreg[344]), .Z(n7701) );
  NAND U7853 ( .A(n7621), .B(sreg[343]), .Z(n7625) );
  OR U7854 ( .A(n7623), .B(n7622), .Z(n7624) );
  AND U7855 ( .A(n7625), .B(n7624), .Z(n7700) );
  XOR U7856 ( .A(n7701), .B(n7700), .Z(c[344]) );
  NANDN U7857 ( .A(n7627), .B(n7626), .Z(n7631) );
  NAND U7858 ( .A(n7629), .B(n7628), .Z(n7630) );
  NAND U7859 ( .A(n7631), .B(n7630), .Z(n7707) );
  NANDN U7860 ( .A(n7633), .B(n7632), .Z(n7637) );
  OR U7861 ( .A(n7635), .B(n7634), .Z(n7636) );
  NAND U7862 ( .A(n7637), .B(n7636), .Z(n7774) );
  XNOR U7863 ( .A(n20052), .B(n7980), .Z(n7728) );
  OR U7864 ( .A(n7728), .B(n20020), .Z(n7640) );
  NANDN U7865 ( .A(n7638), .B(n19960), .Z(n7639) );
  NAND U7866 ( .A(n7640), .B(n7639), .Z(n7725) );
  XNOR U7867 ( .A(n102), .B(n7641), .Z(n7732) );
  OR U7868 ( .A(n7732), .B(n20121), .Z(n7644) );
  NANDN U7869 ( .A(n7642), .B(n20122), .Z(n7643) );
  NAND U7870 ( .A(n7644), .B(n7643), .Z(n7722) );
  XNOR U7871 ( .A(n19975), .B(n8136), .Z(n7735) );
  NANDN U7872 ( .A(n7735), .B(n19883), .Z(n7647) );
  NANDN U7873 ( .A(n7645), .B(n19937), .Z(n7646) );
  AND U7874 ( .A(n7647), .B(n7646), .Z(n7723) );
  XNOR U7875 ( .A(n7722), .B(n7723), .Z(n7724) );
  XNOR U7876 ( .A(n7725), .B(n7724), .Z(n7765) );
  NANDN U7877 ( .A(n7649), .B(n7648), .Z(n7653) );
  NAND U7878 ( .A(n7651), .B(n7650), .Z(n7652) );
  NAND U7879 ( .A(n7653), .B(n7652), .Z(n7766) );
  XNOR U7880 ( .A(n7765), .B(n7766), .Z(n7767) );
  NANDN U7881 ( .A(n7655), .B(n7654), .Z(n7659) );
  NAND U7882 ( .A(n7657), .B(n7656), .Z(n7658) );
  AND U7883 ( .A(n7659), .B(n7658), .Z(n7768) );
  XNOR U7884 ( .A(n7767), .B(n7768), .Z(n7712) );
  NANDN U7885 ( .A(n7661), .B(n7660), .Z(n7665) );
  OR U7886 ( .A(n7663), .B(n7662), .Z(n7664) );
  NAND U7887 ( .A(n7665), .B(n7664), .Z(n7762) );
  NAND U7888 ( .A(b[0]), .B(a[105]), .Z(n7666) );
  XNOR U7889 ( .A(b[1]), .B(n7666), .Z(n7668) );
  NAND U7890 ( .A(a[104]), .B(n98), .Z(n7667) );
  AND U7891 ( .A(n7668), .B(n7667), .Z(n7738) );
  XNOR U7892 ( .A(n20154), .B(n7797), .Z(n7747) );
  OR U7893 ( .A(n7747), .B(n20057), .Z(n7671) );
  NANDN U7894 ( .A(n7669), .B(n20098), .Z(n7670) );
  AND U7895 ( .A(n7671), .B(n7670), .Z(n7739) );
  XOR U7896 ( .A(n7738), .B(n7739), .Z(n7741) );
  NAND U7897 ( .A(a[89]), .B(b[15]), .Z(n7740) );
  XOR U7898 ( .A(n7741), .B(n7740), .Z(n7759) );
  NAND U7899 ( .A(n19722), .B(n7672), .Z(n7674) );
  XNOR U7900 ( .A(b[5]), .B(n8448), .Z(n7750) );
  NANDN U7901 ( .A(n19640), .B(n7750), .Z(n7673) );
  NAND U7902 ( .A(n7674), .B(n7673), .Z(n7719) );
  XNOR U7903 ( .A(n19714), .B(n8265), .Z(n7753) );
  NANDN U7904 ( .A(n7753), .B(n19766), .Z(n7677) );
  NANDN U7905 ( .A(n7675), .B(n19767), .Z(n7676) );
  NAND U7906 ( .A(n7677), .B(n7676), .Z(n7716) );
  NAND U7907 ( .A(n19554), .B(n7678), .Z(n7680) );
  IV U7908 ( .A(a[103]), .Z(n8577) );
  XNOR U7909 ( .A(b[3]), .B(n8577), .Z(n7756) );
  NANDN U7910 ( .A(n19521), .B(n7756), .Z(n7679) );
  AND U7911 ( .A(n7680), .B(n7679), .Z(n7717) );
  XNOR U7912 ( .A(n7716), .B(n7717), .Z(n7718) );
  XOR U7913 ( .A(n7719), .B(n7718), .Z(n7760) );
  XOR U7914 ( .A(n7759), .B(n7760), .Z(n7761) );
  XNOR U7915 ( .A(n7762), .B(n7761), .Z(n7710) );
  NAND U7916 ( .A(n7682), .B(n7681), .Z(n7686) );
  NAND U7917 ( .A(n7684), .B(n7683), .Z(n7685) );
  NAND U7918 ( .A(n7686), .B(n7685), .Z(n7711) );
  XOR U7919 ( .A(n7710), .B(n7711), .Z(n7713) );
  XNOR U7920 ( .A(n7712), .B(n7713), .Z(n7771) );
  NANDN U7921 ( .A(n7688), .B(n7687), .Z(n7692) );
  NAND U7922 ( .A(n7690), .B(n7689), .Z(n7691) );
  NAND U7923 ( .A(n7692), .B(n7691), .Z(n7772) );
  XNOR U7924 ( .A(n7771), .B(n7772), .Z(n7773) );
  XOR U7925 ( .A(n7774), .B(n7773), .Z(n7704) );
  NANDN U7926 ( .A(n7694), .B(n7693), .Z(n7698) );
  NANDN U7927 ( .A(n7696), .B(n7695), .Z(n7697) );
  NAND U7928 ( .A(n7698), .B(n7697), .Z(n7705) );
  XNOR U7929 ( .A(n7704), .B(n7705), .Z(n7706) );
  XNOR U7930 ( .A(n7707), .B(n7706), .Z(n7777) );
  XNOR U7931 ( .A(n7777), .B(sreg[345]), .Z(n7779) );
  NAND U7932 ( .A(n7699), .B(sreg[344]), .Z(n7703) );
  OR U7933 ( .A(n7701), .B(n7700), .Z(n7702) );
  AND U7934 ( .A(n7703), .B(n7702), .Z(n7778) );
  XOR U7935 ( .A(n7779), .B(n7778), .Z(c[345]) );
  NANDN U7936 ( .A(n7705), .B(n7704), .Z(n7709) );
  NAND U7937 ( .A(n7707), .B(n7706), .Z(n7708) );
  NAND U7938 ( .A(n7709), .B(n7708), .Z(n7785) );
  NANDN U7939 ( .A(n7711), .B(n7710), .Z(n7715) );
  OR U7940 ( .A(n7713), .B(n7712), .Z(n7714) );
  NAND U7941 ( .A(n7715), .B(n7714), .Z(n7852) );
  NANDN U7942 ( .A(n7717), .B(n7716), .Z(n7721) );
  NAND U7943 ( .A(n7719), .B(n7718), .Z(n7720) );
  NAND U7944 ( .A(n7721), .B(n7720), .Z(n7846) );
  NANDN U7945 ( .A(n7723), .B(n7722), .Z(n7727) );
  NAND U7946 ( .A(n7725), .B(n7724), .Z(n7726) );
  NAND U7947 ( .A(n7727), .B(n7726), .Z(n7843) );
  XNOR U7948 ( .A(n20052), .B(n8031), .Z(n7794) );
  OR U7949 ( .A(n7794), .B(n20020), .Z(n7730) );
  NANDN U7950 ( .A(n7728), .B(n19960), .Z(n7729) );
  NAND U7951 ( .A(n7730), .B(n7729), .Z(n7807) );
  XNOR U7952 ( .A(n102), .B(n7731), .Z(n7798) );
  OR U7953 ( .A(n7798), .B(n20121), .Z(n7734) );
  NANDN U7954 ( .A(n7732), .B(n20122), .Z(n7733) );
  NAND U7955 ( .A(n7734), .B(n7733), .Z(n7804) );
  XNOR U7956 ( .A(n19975), .B(n8214), .Z(n7801) );
  NANDN U7957 ( .A(n7801), .B(n19883), .Z(n7737) );
  NANDN U7958 ( .A(n7735), .B(n19937), .Z(n7736) );
  AND U7959 ( .A(n7737), .B(n7736), .Z(n7805) );
  XNOR U7960 ( .A(n7804), .B(n7805), .Z(n7806) );
  XNOR U7961 ( .A(n7807), .B(n7806), .Z(n7844) );
  XNOR U7962 ( .A(n7843), .B(n7844), .Z(n7845) );
  XNOR U7963 ( .A(n7846), .B(n7845), .Z(n7791) );
  NANDN U7964 ( .A(n7739), .B(n7738), .Z(n7743) );
  OR U7965 ( .A(n7741), .B(n7740), .Z(n7742) );
  NAND U7966 ( .A(n7743), .B(n7742), .Z(n7840) );
  NAND U7967 ( .A(b[0]), .B(a[106]), .Z(n7744) );
  XNOR U7968 ( .A(b[1]), .B(n7744), .Z(n7746) );
  NAND U7969 ( .A(a[105]), .B(n98), .Z(n7745) );
  AND U7970 ( .A(n7746), .B(n7745), .Z(n7816) );
  XNOR U7971 ( .A(n20154), .B(n7875), .Z(n7825) );
  OR U7972 ( .A(n7825), .B(n20057), .Z(n7749) );
  NANDN U7973 ( .A(n7747), .B(n20098), .Z(n7748) );
  AND U7974 ( .A(n7749), .B(n7748), .Z(n7817) );
  XOR U7975 ( .A(n7816), .B(n7817), .Z(n7819) );
  NAND U7976 ( .A(a[90]), .B(b[15]), .Z(n7818) );
  XOR U7977 ( .A(n7819), .B(n7818), .Z(n7837) );
  NAND U7978 ( .A(n19722), .B(n7750), .Z(n7752) );
  XNOR U7979 ( .A(b[5]), .B(n8499), .Z(n7828) );
  NANDN U7980 ( .A(n19640), .B(n7828), .Z(n7751) );
  NAND U7981 ( .A(n7752), .B(n7751), .Z(n7813) );
  XNOR U7982 ( .A(n19714), .B(n8343), .Z(n7831) );
  NANDN U7983 ( .A(n7831), .B(n19766), .Z(n7755) );
  NANDN U7984 ( .A(n7753), .B(n19767), .Z(n7754) );
  NAND U7985 ( .A(n7755), .B(n7754), .Z(n7810) );
  NAND U7986 ( .A(n19554), .B(n7756), .Z(n7758) );
  IV U7987 ( .A(a[104]), .Z(n8682) );
  XNOR U7988 ( .A(b[3]), .B(n8682), .Z(n7834) );
  NANDN U7989 ( .A(n19521), .B(n7834), .Z(n7757) );
  AND U7990 ( .A(n7758), .B(n7757), .Z(n7811) );
  XNOR U7991 ( .A(n7810), .B(n7811), .Z(n7812) );
  XOR U7992 ( .A(n7813), .B(n7812), .Z(n7838) );
  XOR U7993 ( .A(n7837), .B(n7838), .Z(n7839) );
  XNOR U7994 ( .A(n7840), .B(n7839), .Z(n7788) );
  NAND U7995 ( .A(n7760), .B(n7759), .Z(n7764) );
  NAND U7996 ( .A(n7762), .B(n7761), .Z(n7763) );
  NAND U7997 ( .A(n7764), .B(n7763), .Z(n7789) );
  XNOR U7998 ( .A(n7788), .B(n7789), .Z(n7790) );
  XOR U7999 ( .A(n7791), .B(n7790), .Z(n7849) );
  NANDN U8000 ( .A(n7766), .B(n7765), .Z(n7770) );
  NAND U8001 ( .A(n7768), .B(n7767), .Z(n7769) );
  NAND U8002 ( .A(n7770), .B(n7769), .Z(n7850) );
  XOR U8003 ( .A(n7849), .B(n7850), .Z(n7851) );
  XOR U8004 ( .A(n7852), .B(n7851), .Z(n7782) );
  NANDN U8005 ( .A(n7772), .B(n7771), .Z(n7776) );
  NANDN U8006 ( .A(n7774), .B(n7773), .Z(n7775) );
  NAND U8007 ( .A(n7776), .B(n7775), .Z(n7783) );
  XNOR U8008 ( .A(n7782), .B(n7783), .Z(n7784) );
  XNOR U8009 ( .A(n7785), .B(n7784), .Z(n7855) );
  XNOR U8010 ( .A(n7855), .B(sreg[346]), .Z(n7857) );
  NAND U8011 ( .A(n7777), .B(sreg[345]), .Z(n7781) );
  OR U8012 ( .A(n7779), .B(n7778), .Z(n7780) );
  AND U8013 ( .A(n7781), .B(n7780), .Z(n7856) );
  XOR U8014 ( .A(n7857), .B(n7856), .Z(c[346]) );
  NANDN U8015 ( .A(n7783), .B(n7782), .Z(n7787) );
  NAND U8016 ( .A(n7785), .B(n7784), .Z(n7786) );
  NAND U8017 ( .A(n7787), .B(n7786), .Z(n7863) );
  NANDN U8018 ( .A(n7789), .B(n7788), .Z(n7793) );
  NAND U8019 ( .A(n7791), .B(n7790), .Z(n7792) );
  NAND U8020 ( .A(n7793), .B(n7792), .Z(n7930) );
  XNOR U8021 ( .A(n20052), .B(n8136), .Z(n7872) );
  OR U8022 ( .A(n7872), .B(n20020), .Z(n7796) );
  NANDN U8023 ( .A(n7794), .B(n19960), .Z(n7795) );
  NAND U8024 ( .A(n7796), .B(n7795), .Z(n7885) );
  XNOR U8025 ( .A(n102), .B(n7797), .Z(n7876) );
  OR U8026 ( .A(n7876), .B(n20121), .Z(n7800) );
  NANDN U8027 ( .A(n7798), .B(n20122), .Z(n7799) );
  NAND U8028 ( .A(n7800), .B(n7799), .Z(n7882) );
  XNOR U8029 ( .A(n19975), .B(n8265), .Z(n7879) );
  NANDN U8030 ( .A(n7879), .B(n19883), .Z(n7803) );
  NANDN U8031 ( .A(n7801), .B(n19937), .Z(n7802) );
  AND U8032 ( .A(n7803), .B(n7802), .Z(n7883) );
  XNOR U8033 ( .A(n7882), .B(n7883), .Z(n7884) );
  XNOR U8034 ( .A(n7885), .B(n7884), .Z(n7921) );
  NANDN U8035 ( .A(n7805), .B(n7804), .Z(n7809) );
  NAND U8036 ( .A(n7807), .B(n7806), .Z(n7808) );
  NAND U8037 ( .A(n7809), .B(n7808), .Z(n7922) );
  XNOR U8038 ( .A(n7921), .B(n7922), .Z(n7923) );
  NANDN U8039 ( .A(n7811), .B(n7810), .Z(n7815) );
  NAND U8040 ( .A(n7813), .B(n7812), .Z(n7814) );
  AND U8041 ( .A(n7815), .B(n7814), .Z(n7924) );
  XNOR U8042 ( .A(n7923), .B(n7924), .Z(n7868) );
  NANDN U8043 ( .A(n7817), .B(n7816), .Z(n7821) );
  OR U8044 ( .A(n7819), .B(n7818), .Z(n7820) );
  NAND U8045 ( .A(n7821), .B(n7820), .Z(n7918) );
  NAND U8046 ( .A(b[0]), .B(a[107]), .Z(n7822) );
  XNOR U8047 ( .A(b[1]), .B(n7822), .Z(n7824) );
  NAND U8048 ( .A(a[106]), .B(n98), .Z(n7823) );
  AND U8049 ( .A(n7824), .B(n7823), .Z(n7894) );
  XNOR U8050 ( .A(n20154), .B(n7980), .Z(n7903) );
  OR U8051 ( .A(n7903), .B(n20057), .Z(n7827) );
  NANDN U8052 ( .A(n7825), .B(n20098), .Z(n7826) );
  AND U8053 ( .A(n7827), .B(n7826), .Z(n7895) );
  XOR U8054 ( .A(n7894), .B(n7895), .Z(n7897) );
  NAND U8055 ( .A(a[91]), .B(b[15]), .Z(n7896) );
  XOR U8056 ( .A(n7897), .B(n7896), .Z(n7915) );
  NAND U8057 ( .A(n19722), .B(n7828), .Z(n7830) );
  XNOR U8058 ( .A(b[5]), .B(n8577), .Z(n7906) );
  NANDN U8059 ( .A(n19640), .B(n7906), .Z(n7829) );
  NAND U8060 ( .A(n7830), .B(n7829), .Z(n7891) );
  XNOR U8061 ( .A(n19714), .B(n8448), .Z(n7909) );
  NANDN U8062 ( .A(n7909), .B(n19766), .Z(n7833) );
  NANDN U8063 ( .A(n7831), .B(n19767), .Z(n7832) );
  NAND U8064 ( .A(n7833), .B(n7832), .Z(n7888) );
  NAND U8065 ( .A(n19554), .B(n7834), .Z(n7836) );
  IV U8066 ( .A(a[105]), .Z(n8733) );
  XNOR U8067 ( .A(b[3]), .B(n8733), .Z(n7912) );
  NANDN U8068 ( .A(n19521), .B(n7912), .Z(n7835) );
  AND U8069 ( .A(n7836), .B(n7835), .Z(n7889) );
  XNOR U8070 ( .A(n7888), .B(n7889), .Z(n7890) );
  XOR U8071 ( .A(n7891), .B(n7890), .Z(n7916) );
  XOR U8072 ( .A(n7915), .B(n7916), .Z(n7917) );
  XNOR U8073 ( .A(n7918), .B(n7917), .Z(n7866) );
  NAND U8074 ( .A(n7838), .B(n7837), .Z(n7842) );
  NAND U8075 ( .A(n7840), .B(n7839), .Z(n7841) );
  NAND U8076 ( .A(n7842), .B(n7841), .Z(n7867) );
  XOR U8077 ( .A(n7866), .B(n7867), .Z(n7869) );
  XNOR U8078 ( .A(n7868), .B(n7869), .Z(n7927) );
  NANDN U8079 ( .A(n7844), .B(n7843), .Z(n7848) );
  NAND U8080 ( .A(n7846), .B(n7845), .Z(n7847) );
  AND U8081 ( .A(n7848), .B(n7847), .Z(n7928) );
  XNOR U8082 ( .A(n7927), .B(n7928), .Z(n7929) );
  XOR U8083 ( .A(n7930), .B(n7929), .Z(n7860) );
  OR U8084 ( .A(n7850), .B(n7849), .Z(n7854) );
  NANDN U8085 ( .A(n7852), .B(n7851), .Z(n7853) );
  NAND U8086 ( .A(n7854), .B(n7853), .Z(n7861) );
  XNOR U8087 ( .A(n7860), .B(n7861), .Z(n7862) );
  XNOR U8088 ( .A(n7863), .B(n7862), .Z(n7933) );
  XNOR U8089 ( .A(n7933), .B(sreg[347]), .Z(n7935) );
  NAND U8090 ( .A(n7855), .B(sreg[346]), .Z(n7859) );
  OR U8091 ( .A(n7857), .B(n7856), .Z(n7858) );
  AND U8092 ( .A(n7859), .B(n7858), .Z(n7934) );
  XOR U8093 ( .A(n7935), .B(n7934), .Z(c[347]) );
  NANDN U8094 ( .A(n7861), .B(n7860), .Z(n7865) );
  NAND U8095 ( .A(n7863), .B(n7862), .Z(n7864) );
  NAND U8096 ( .A(n7865), .B(n7864), .Z(n7941) );
  NANDN U8097 ( .A(n7867), .B(n7866), .Z(n7871) );
  OR U8098 ( .A(n7869), .B(n7868), .Z(n7870) );
  NAND U8099 ( .A(n7871), .B(n7870), .Z(n8008) );
  XNOR U8100 ( .A(n20052), .B(n8214), .Z(n7977) );
  OR U8101 ( .A(n7977), .B(n20020), .Z(n7874) );
  NANDN U8102 ( .A(n7872), .B(n19960), .Z(n7873) );
  NAND U8103 ( .A(n7874), .B(n7873), .Z(n7990) );
  XNOR U8104 ( .A(n102), .B(n7875), .Z(n7981) );
  OR U8105 ( .A(n7981), .B(n20121), .Z(n7878) );
  NANDN U8106 ( .A(n7876), .B(n20122), .Z(n7877) );
  NAND U8107 ( .A(n7878), .B(n7877), .Z(n7987) );
  XNOR U8108 ( .A(n19975), .B(n8343), .Z(n7984) );
  NANDN U8109 ( .A(n7984), .B(n19883), .Z(n7881) );
  NANDN U8110 ( .A(n7879), .B(n19937), .Z(n7880) );
  AND U8111 ( .A(n7881), .B(n7880), .Z(n7988) );
  XNOR U8112 ( .A(n7987), .B(n7988), .Z(n7989) );
  XNOR U8113 ( .A(n7990), .B(n7989), .Z(n7999) );
  NANDN U8114 ( .A(n7883), .B(n7882), .Z(n7887) );
  NAND U8115 ( .A(n7885), .B(n7884), .Z(n7886) );
  NAND U8116 ( .A(n7887), .B(n7886), .Z(n8000) );
  XNOR U8117 ( .A(n7999), .B(n8000), .Z(n8001) );
  NANDN U8118 ( .A(n7889), .B(n7888), .Z(n7893) );
  NAND U8119 ( .A(n7891), .B(n7890), .Z(n7892) );
  AND U8120 ( .A(n7893), .B(n7892), .Z(n8002) );
  XNOR U8121 ( .A(n8001), .B(n8002), .Z(n7946) );
  NANDN U8122 ( .A(n7895), .B(n7894), .Z(n7899) );
  OR U8123 ( .A(n7897), .B(n7896), .Z(n7898) );
  NAND U8124 ( .A(n7899), .B(n7898), .Z(n7974) );
  NAND U8125 ( .A(b[0]), .B(a[108]), .Z(n7900) );
  XNOR U8126 ( .A(b[1]), .B(n7900), .Z(n7902) );
  NAND U8127 ( .A(a[107]), .B(n98), .Z(n7901) );
  AND U8128 ( .A(n7902), .B(n7901), .Z(n7950) );
  XNOR U8129 ( .A(n20154), .B(n8031), .Z(n7956) );
  OR U8130 ( .A(n7956), .B(n20057), .Z(n7905) );
  NANDN U8131 ( .A(n7903), .B(n20098), .Z(n7904) );
  AND U8132 ( .A(n7905), .B(n7904), .Z(n7951) );
  XOR U8133 ( .A(n7950), .B(n7951), .Z(n7953) );
  NAND U8134 ( .A(a[92]), .B(b[15]), .Z(n7952) );
  XOR U8135 ( .A(n7953), .B(n7952), .Z(n7971) );
  NAND U8136 ( .A(n19722), .B(n7906), .Z(n7908) );
  XNOR U8137 ( .A(b[5]), .B(n8682), .Z(n7962) );
  NANDN U8138 ( .A(n19640), .B(n7962), .Z(n7907) );
  NAND U8139 ( .A(n7908), .B(n7907), .Z(n7996) );
  XNOR U8140 ( .A(n19714), .B(n8499), .Z(n7965) );
  NANDN U8141 ( .A(n7965), .B(n19766), .Z(n7911) );
  NANDN U8142 ( .A(n7909), .B(n19767), .Z(n7910) );
  NAND U8143 ( .A(n7911), .B(n7910), .Z(n7993) );
  NAND U8144 ( .A(n19554), .B(n7912), .Z(n7914) );
  IV U8145 ( .A(a[106]), .Z(n8838) );
  XNOR U8146 ( .A(b[3]), .B(n8838), .Z(n7968) );
  NANDN U8147 ( .A(n19521), .B(n7968), .Z(n7913) );
  AND U8148 ( .A(n7914), .B(n7913), .Z(n7994) );
  XNOR U8149 ( .A(n7993), .B(n7994), .Z(n7995) );
  XOR U8150 ( .A(n7996), .B(n7995), .Z(n7972) );
  XOR U8151 ( .A(n7971), .B(n7972), .Z(n7973) );
  XNOR U8152 ( .A(n7974), .B(n7973), .Z(n7944) );
  NAND U8153 ( .A(n7916), .B(n7915), .Z(n7920) );
  NAND U8154 ( .A(n7918), .B(n7917), .Z(n7919) );
  NAND U8155 ( .A(n7920), .B(n7919), .Z(n7945) );
  XOR U8156 ( .A(n7944), .B(n7945), .Z(n7947) );
  XNOR U8157 ( .A(n7946), .B(n7947), .Z(n8005) );
  NANDN U8158 ( .A(n7922), .B(n7921), .Z(n7926) );
  NAND U8159 ( .A(n7924), .B(n7923), .Z(n7925) );
  NAND U8160 ( .A(n7926), .B(n7925), .Z(n8006) );
  XNOR U8161 ( .A(n8005), .B(n8006), .Z(n8007) );
  XOR U8162 ( .A(n8008), .B(n8007), .Z(n7938) );
  NANDN U8163 ( .A(n7928), .B(n7927), .Z(n7932) );
  NANDN U8164 ( .A(n7930), .B(n7929), .Z(n7931) );
  NAND U8165 ( .A(n7932), .B(n7931), .Z(n7939) );
  XNOR U8166 ( .A(n7938), .B(n7939), .Z(n7940) );
  XNOR U8167 ( .A(n7941), .B(n7940), .Z(n8011) );
  XNOR U8168 ( .A(n8011), .B(sreg[348]), .Z(n8013) );
  NAND U8169 ( .A(n7933), .B(sreg[347]), .Z(n7937) );
  OR U8170 ( .A(n7935), .B(n7934), .Z(n7936) );
  AND U8171 ( .A(n7937), .B(n7936), .Z(n8012) );
  XOR U8172 ( .A(n8013), .B(n8012), .Z(c[348]) );
  NANDN U8173 ( .A(n7939), .B(n7938), .Z(n7943) );
  NAND U8174 ( .A(n7941), .B(n7940), .Z(n7942) );
  NAND U8175 ( .A(n7943), .B(n7942), .Z(n8019) );
  NANDN U8176 ( .A(n7945), .B(n7944), .Z(n7949) );
  OR U8177 ( .A(n7947), .B(n7946), .Z(n7948) );
  NAND U8178 ( .A(n7949), .B(n7948), .Z(n8086) );
  NANDN U8179 ( .A(n7951), .B(n7950), .Z(n7955) );
  OR U8180 ( .A(n7953), .B(n7952), .Z(n7954) );
  NAND U8181 ( .A(n7955), .B(n7954), .Z(n8074) );
  XNOR U8182 ( .A(n20154), .B(n8136), .Z(n8059) );
  OR U8183 ( .A(n8059), .B(n20057), .Z(n7958) );
  NANDN U8184 ( .A(n7956), .B(n20098), .Z(n7957) );
  AND U8185 ( .A(n7958), .B(n7957), .Z(n8051) );
  NAND U8186 ( .A(b[0]), .B(a[109]), .Z(n7959) );
  XNOR U8187 ( .A(b[1]), .B(n7959), .Z(n7961) );
  NAND U8188 ( .A(a[108]), .B(n98), .Z(n7960) );
  AND U8189 ( .A(n7961), .B(n7960), .Z(n8050) );
  XOR U8190 ( .A(n8051), .B(n8050), .Z(n8053) );
  NAND U8191 ( .A(a[93]), .B(b[15]), .Z(n8052) );
  XOR U8192 ( .A(n8053), .B(n8052), .Z(n8071) );
  NAND U8193 ( .A(n19722), .B(n7962), .Z(n7964) );
  XNOR U8194 ( .A(b[5]), .B(n8733), .Z(n8062) );
  NANDN U8195 ( .A(n19640), .B(n8062), .Z(n7963) );
  NAND U8196 ( .A(n7964), .B(n7963), .Z(n8047) );
  XNOR U8197 ( .A(n19714), .B(n8577), .Z(n8065) );
  NANDN U8198 ( .A(n8065), .B(n19766), .Z(n7967) );
  NANDN U8199 ( .A(n7965), .B(n19767), .Z(n7966) );
  NAND U8200 ( .A(n7967), .B(n7966), .Z(n8044) );
  NAND U8201 ( .A(n19554), .B(n7968), .Z(n7970) );
  IV U8202 ( .A(a[107]), .Z(n8916) );
  XNOR U8203 ( .A(b[3]), .B(n8916), .Z(n8068) );
  NANDN U8204 ( .A(n19521), .B(n8068), .Z(n7969) );
  AND U8205 ( .A(n7970), .B(n7969), .Z(n8045) );
  XNOR U8206 ( .A(n8044), .B(n8045), .Z(n8046) );
  XOR U8207 ( .A(n8047), .B(n8046), .Z(n8072) );
  XOR U8208 ( .A(n8071), .B(n8072), .Z(n8073) );
  XNOR U8209 ( .A(n8074), .B(n8073), .Z(n8022) );
  NAND U8210 ( .A(n7972), .B(n7971), .Z(n7976) );
  NAND U8211 ( .A(n7974), .B(n7973), .Z(n7975) );
  NAND U8212 ( .A(n7976), .B(n7975), .Z(n8023) );
  XOR U8213 ( .A(n8022), .B(n8023), .Z(n8025) );
  XNOR U8214 ( .A(n20052), .B(n8265), .Z(n8028) );
  OR U8215 ( .A(n8028), .B(n20020), .Z(n7979) );
  NANDN U8216 ( .A(n7977), .B(n19960), .Z(n7978) );
  NAND U8217 ( .A(n7979), .B(n7978), .Z(n8041) );
  XNOR U8218 ( .A(n102), .B(n7980), .Z(n8032) );
  OR U8219 ( .A(n8032), .B(n20121), .Z(n7983) );
  NANDN U8220 ( .A(n7981), .B(n20122), .Z(n7982) );
  NAND U8221 ( .A(n7983), .B(n7982), .Z(n8038) );
  XNOR U8222 ( .A(n19975), .B(n8448), .Z(n8035) );
  NANDN U8223 ( .A(n8035), .B(n19883), .Z(n7986) );
  NANDN U8224 ( .A(n7984), .B(n19937), .Z(n7985) );
  AND U8225 ( .A(n7986), .B(n7985), .Z(n8039) );
  XNOR U8226 ( .A(n8038), .B(n8039), .Z(n8040) );
  XNOR U8227 ( .A(n8041), .B(n8040), .Z(n8077) );
  NANDN U8228 ( .A(n7988), .B(n7987), .Z(n7992) );
  NAND U8229 ( .A(n7990), .B(n7989), .Z(n7991) );
  NAND U8230 ( .A(n7992), .B(n7991), .Z(n8078) );
  XNOR U8231 ( .A(n8077), .B(n8078), .Z(n8079) );
  NANDN U8232 ( .A(n7994), .B(n7993), .Z(n7998) );
  NAND U8233 ( .A(n7996), .B(n7995), .Z(n7997) );
  AND U8234 ( .A(n7998), .B(n7997), .Z(n8080) );
  XNOR U8235 ( .A(n8079), .B(n8080), .Z(n8024) );
  XNOR U8236 ( .A(n8025), .B(n8024), .Z(n8083) );
  NANDN U8237 ( .A(n8000), .B(n7999), .Z(n8004) );
  NAND U8238 ( .A(n8002), .B(n8001), .Z(n8003) );
  NAND U8239 ( .A(n8004), .B(n8003), .Z(n8084) );
  XNOR U8240 ( .A(n8083), .B(n8084), .Z(n8085) );
  XOR U8241 ( .A(n8086), .B(n8085), .Z(n8016) );
  NANDN U8242 ( .A(n8006), .B(n8005), .Z(n8010) );
  NANDN U8243 ( .A(n8008), .B(n8007), .Z(n8009) );
  NAND U8244 ( .A(n8010), .B(n8009), .Z(n8017) );
  XNOR U8245 ( .A(n8016), .B(n8017), .Z(n8018) );
  XNOR U8246 ( .A(n8019), .B(n8018), .Z(n8089) );
  XNOR U8247 ( .A(n8089), .B(sreg[349]), .Z(n8091) );
  NAND U8248 ( .A(n8011), .B(sreg[348]), .Z(n8015) );
  OR U8249 ( .A(n8013), .B(n8012), .Z(n8014) );
  AND U8250 ( .A(n8015), .B(n8014), .Z(n8090) );
  XOR U8251 ( .A(n8091), .B(n8090), .Z(c[349]) );
  NANDN U8252 ( .A(n8017), .B(n8016), .Z(n8021) );
  NAND U8253 ( .A(n8019), .B(n8018), .Z(n8020) );
  NAND U8254 ( .A(n8021), .B(n8020), .Z(n8097) );
  NANDN U8255 ( .A(n8023), .B(n8022), .Z(n8027) );
  OR U8256 ( .A(n8025), .B(n8024), .Z(n8026) );
  NAND U8257 ( .A(n8027), .B(n8026), .Z(n8164) );
  XNOR U8258 ( .A(n20052), .B(n8343), .Z(n8133) );
  OR U8259 ( .A(n8133), .B(n20020), .Z(n8030) );
  NANDN U8260 ( .A(n8028), .B(n19960), .Z(n8029) );
  NAND U8261 ( .A(n8030), .B(n8029), .Z(n8146) );
  XNOR U8262 ( .A(n102), .B(n8031), .Z(n8137) );
  OR U8263 ( .A(n8137), .B(n20121), .Z(n8034) );
  NANDN U8264 ( .A(n8032), .B(n20122), .Z(n8033) );
  NAND U8265 ( .A(n8034), .B(n8033), .Z(n8143) );
  XNOR U8266 ( .A(n19975), .B(n8499), .Z(n8140) );
  NANDN U8267 ( .A(n8140), .B(n19883), .Z(n8037) );
  NANDN U8268 ( .A(n8035), .B(n19937), .Z(n8036) );
  AND U8269 ( .A(n8037), .B(n8036), .Z(n8144) );
  XNOR U8270 ( .A(n8143), .B(n8144), .Z(n8145) );
  XNOR U8271 ( .A(n8146), .B(n8145), .Z(n8155) );
  NANDN U8272 ( .A(n8039), .B(n8038), .Z(n8043) );
  NAND U8273 ( .A(n8041), .B(n8040), .Z(n8042) );
  NAND U8274 ( .A(n8043), .B(n8042), .Z(n8156) );
  XNOR U8275 ( .A(n8155), .B(n8156), .Z(n8157) );
  NANDN U8276 ( .A(n8045), .B(n8044), .Z(n8049) );
  NAND U8277 ( .A(n8047), .B(n8046), .Z(n8048) );
  AND U8278 ( .A(n8049), .B(n8048), .Z(n8158) );
  XNOR U8279 ( .A(n8157), .B(n8158), .Z(n8102) );
  NANDN U8280 ( .A(n8051), .B(n8050), .Z(n8055) );
  OR U8281 ( .A(n8053), .B(n8052), .Z(n8054) );
  NAND U8282 ( .A(n8055), .B(n8054), .Z(n8130) );
  NAND U8283 ( .A(b[0]), .B(a[110]), .Z(n8056) );
  XNOR U8284 ( .A(b[1]), .B(n8056), .Z(n8058) );
  NAND U8285 ( .A(a[109]), .B(n98), .Z(n8057) );
  AND U8286 ( .A(n8058), .B(n8057), .Z(n8106) );
  XNOR U8287 ( .A(n20154), .B(n8214), .Z(n8115) );
  OR U8288 ( .A(n8115), .B(n20057), .Z(n8061) );
  NANDN U8289 ( .A(n8059), .B(n20098), .Z(n8060) );
  AND U8290 ( .A(n8061), .B(n8060), .Z(n8107) );
  XOR U8291 ( .A(n8106), .B(n8107), .Z(n8109) );
  NAND U8292 ( .A(a[94]), .B(b[15]), .Z(n8108) );
  XOR U8293 ( .A(n8109), .B(n8108), .Z(n8127) );
  NAND U8294 ( .A(n19722), .B(n8062), .Z(n8064) );
  XNOR U8295 ( .A(b[5]), .B(n8838), .Z(n8118) );
  NANDN U8296 ( .A(n19640), .B(n8118), .Z(n8063) );
  NAND U8297 ( .A(n8064), .B(n8063), .Z(n8152) );
  XNOR U8298 ( .A(n19714), .B(n8682), .Z(n8121) );
  NANDN U8299 ( .A(n8121), .B(n19766), .Z(n8067) );
  NANDN U8300 ( .A(n8065), .B(n19767), .Z(n8066) );
  NAND U8301 ( .A(n8067), .B(n8066), .Z(n8149) );
  NAND U8302 ( .A(n19554), .B(n8068), .Z(n8070) );
  IV U8303 ( .A(a[108]), .Z(n8967) );
  XNOR U8304 ( .A(b[3]), .B(n8967), .Z(n8124) );
  NANDN U8305 ( .A(n19521), .B(n8124), .Z(n8069) );
  AND U8306 ( .A(n8070), .B(n8069), .Z(n8150) );
  XNOR U8307 ( .A(n8149), .B(n8150), .Z(n8151) );
  XOR U8308 ( .A(n8152), .B(n8151), .Z(n8128) );
  XOR U8309 ( .A(n8127), .B(n8128), .Z(n8129) );
  XNOR U8310 ( .A(n8130), .B(n8129), .Z(n8100) );
  NAND U8311 ( .A(n8072), .B(n8071), .Z(n8076) );
  NAND U8312 ( .A(n8074), .B(n8073), .Z(n8075) );
  NAND U8313 ( .A(n8076), .B(n8075), .Z(n8101) );
  XOR U8314 ( .A(n8100), .B(n8101), .Z(n8103) );
  XNOR U8315 ( .A(n8102), .B(n8103), .Z(n8161) );
  NANDN U8316 ( .A(n8078), .B(n8077), .Z(n8082) );
  NAND U8317 ( .A(n8080), .B(n8079), .Z(n8081) );
  NAND U8318 ( .A(n8082), .B(n8081), .Z(n8162) );
  XNOR U8319 ( .A(n8161), .B(n8162), .Z(n8163) );
  XOR U8320 ( .A(n8164), .B(n8163), .Z(n8094) );
  NANDN U8321 ( .A(n8084), .B(n8083), .Z(n8088) );
  NANDN U8322 ( .A(n8086), .B(n8085), .Z(n8087) );
  NAND U8323 ( .A(n8088), .B(n8087), .Z(n8095) );
  XNOR U8324 ( .A(n8094), .B(n8095), .Z(n8096) );
  XNOR U8325 ( .A(n8097), .B(n8096), .Z(n8167) );
  XNOR U8326 ( .A(n8167), .B(sreg[350]), .Z(n8169) );
  NAND U8327 ( .A(n8089), .B(sreg[349]), .Z(n8093) );
  OR U8328 ( .A(n8091), .B(n8090), .Z(n8092) );
  AND U8329 ( .A(n8093), .B(n8092), .Z(n8168) );
  XOR U8330 ( .A(n8169), .B(n8168), .Z(c[350]) );
  NANDN U8331 ( .A(n8095), .B(n8094), .Z(n8099) );
  NAND U8332 ( .A(n8097), .B(n8096), .Z(n8098) );
  NAND U8333 ( .A(n8099), .B(n8098), .Z(n8175) );
  NANDN U8334 ( .A(n8101), .B(n8100), .Z(n8105) );
  OR U8335 ( .A(n8103), .B(n8102), .Z(n8104) );
  NAND U8336 ( .A(n8105), .B(n8104), .Z(n8242) );
  NANDN U8337 ( .A(n8107), .B(n8106), .Z(n8111) );
  OR U8338 ( .A(n8109), .B(n8108), .Z(n8110) );
  NAND U8339 ( .A(n8111), .B(n8110), .Z(n8208) );
  NAND U8340 ( .A(b[0]), .B(a[111]), .Z(n8112) );
  XNOR U8341 ( .A(b[1]), .B(n8112), .Z(n8114) );
  NAND U8342 ( .A(a[110]), .B(n98), .Z(n8113) );
  AND U8343 ( .A(n8114), .B(n8113), .Z(n8184) );
  XNOR U8344 ( .A(n20154), .B(n8265), .Z(n8193) );
  OR U8345 ( .A(n8193), .B(n20057), .Z(n8117) );
  NANDN U8346 ( .A(n8115), .B(n20098), .Z(n8116) );
  AND U8347 ( .A(n8117), .B(n8116), .Z(n8185) );
  XOR U8348 ( .A(n8184), .B(n8185), .Z(n8187) );
  NAND U8349 ( .A(a[95]), .B(b[15]), .Z(n8186) );
  XOR U8350 ( .A(n8187), .B(n8186), .Z(n8205) );
  NAND U8351 ( .A(n19722), .B(n8118), .Z(n8120) );
  XNOR U8352 ( .A(b[5]), .B(n8916), .Z(n8196) );
  NANDN U8353 ( .A(n19640), .B(n8196), .Z(n8119) );
  NAND U8354 ( .A(n8120), .B(n8119), .Z(n8230) );
  XNOR U8355 ( .A(n19714), .B(n8733), .Z(n8199) );
  NANDN U8356 ( .A(n8199), .B(n19766), .Z(n8123) );
  NANDN U8357 ( .A(n8121), .B(n19767), .Z(n8122) );
  NAND U8358 ( .A(n8123), .B(n8122), .Z(n8227) );
  NAND U8359 ( .A(n19554), .B(n8124), .Z(n8126) );
  IV U8360 ( .A(a[109]), .Z(n9045) );
  XNOR U8361 ( .A(b[3]), .B(n9045), .Z(n8202) );
  NANDN U8362 ( .A(n19521), .B(n8202), .Z(n8125) );
  AND U8363 ( .A(n8126), .B(n8125), .Z(n8228) );
  XNOR U8364 ( .A(n8227), .B(n8228), .Z(n8229) );
  XOR U8365 ( .A(n8230), .B(n8229), .Z(n8206) );
  XOR U8366 ( .A(n8205), .B(n8206), .Z(n8207) );
  XNOR U8367 ( .A(n8208), .B(n8207), .Z(n8178) );
  NAND U8368 ( .A(n8128), .B(n8127), .Z(n8132) );
  NAND U8369 ( .A(n8130), .B(n8129), .Z(n8131) );
  NAND U8370 ( .A(n8132), .B(n8131), .Z(n8179) );
  XOR U8371 ( .A(n8178), .B(n8179), .Z(n8181) );
  XNOR U8372 ( .A(n20052), .B(n8448), .Z(n8211) );
  OR U8373 ( .A(n8211), .B(n20020), .Z(n8135) );
  NANDN U8374 ( .A(n8133), .B(n19960), .Z(n8134) );
  NAND U8375 ( .A(n8135), .B(n8134), .Z(n8224) );
  XNOR U8376 ( .A(n102), .B(n8136), .Z(n8215) );
  OR U8377 ( .A(n8215), .B(n20121), .Z(n8139) );
  NANDN U8378 ( .A(n8137), .B(n20122), .Z(n8138) );
  NAND U8379 ( .A(n8139), .B(n8138), .Z(n8221) );
  XNOR U8380 ( .A(n19975), .B(n8577), .Z(n8218) );
  NANDN U8381 ( .A(n8218), .B(n19883), .Z(n8142) );
  NANDN U8382 ( .A(n8140), .B(n19937), .Z(n8141) );
  AND U8383 ( .A(n8142), .B(n8141), .Z(n8222) );
  XNOR U8384 ( .A(n8221), .B(n8222), .Z(n8223) );
  XNOR U8385 ( .A(n8224), .B(n8223), .Z(n8233) );
  NANDN U8386 ( .A(n8144), .B(n8143), .Z(n8148) );
  NAND U8387 ( .A(n8146), .B(n8145), .Z(n8147) );
  NAND U8388 ( .A(n8148), .B(n8147), .Z(n8234) );
  XNOR U8389 ( .A(n8233), .B(n8234), .Z(n8235) );
  NANDN U8390 ( .A(n8150), .B(n8149), .Z(n8154) );
  NAND U8391 ( .A(n8152), .B(n8151), .Z(n8153) );
  AND U8392 ( .A(n8154), .B(n8153), .Z(n8236) );
  XNOR U8393 ( .A(n8235), .B(n8236), .Z(n8180) );
  XNOR U8394 ( .A(n8181), .B(n8180), .Z(n8239) );
  NANDN U8395 ( .A(n8156), .B(n8155), .Z(n8160) );
  NAND U8396 ( .A(n8158), .B(n8157), .Z(n8159) );
  NAND U8397 ( .A(n8160), .B(n8159), .Z(n8240) );
  XNOR U8398 ( .A(n8239), .B(n8240), .Z(n8241) );
  XOR U8399 ( .A(n8242), .B(n8241), .Z(n8172) );
  NANDN U8400 ( .A(n8162), .B(n8161), .Z(n8166) );
  NANDN U8401 ( .A(n8164), .B(n8163), .Z(n8165) );
  NAND U8402 ( .A(n8166), .B(n8165), .Z(n8173) );
  XNOR U8403 ( .A(n8172), .B(n8173), .Z(n8174) );
  XNOR U8404 ( .A(n8175), .B(n8174), .Z(n8245) );
  XNOR U8405 ( .A(n8245), .B(sreg[351]), .Z(n8247) );
  NAND U8406 ( .A(n8167), .B(sreg[350]), .Z(n8171) );
  OR U8407 ( .A(n8169), .B(n8168), .Z(n8170) );
  AND U8408 ( .A(n8171), .B(n8170), .Z(n8246) );
  XOR U8409 ( .A(n8247), .B(n8246), .Z(c[351]) );
  NANDN U8410 ( .A(n8173), .B(n8172), .Z(n8177) );
  NAND U8411 ( .A(n8175), .B(n8174), .Z(n8176) );
  NAND U8412 ( .A(n8177), .B(n8176), .Z(n8253) );
  NANDN U8413 ( .A(n8179), .B(n8178), .Z(n8183) );
  OR U8414 ( .A(n8181), .B(n8180), .Z(n8182) );
  NAND U8415 ( .A(n8183), .B(n8182), .Z(n8320) );
  NANDN U8416 ( .A(n8185), .B(n8184), .Z(n8189) );
  OR U8417 ( .A(n8187), .B(n8186), .Z(n8188) );
  NAND U8418 ( .A(n8189), .B(n8188), .Z(n8308) );
  NAND U8419 ( .A(b[0]), .B(a[112]), .Z(n8190) );
  XNOR U8420 ( .A(b[1]), .B(n8190), .Z(n8192) );
  NAND U8421 ( .A(a[111]), .B(n98), .Z(n8191) );
  AND U8422 ( .A(n8192), .B(n8191), .Z(n8284) );
  XNOR U8423 ( .A(n20154), .B(n8343), .Z(n8290) );
  OR U8424 ( .A(n8290), .B(n20057), .Z(n8195) );
  NANDN U8425 ( .A(n8193), .B(n20098), .Z(n8194) );
  AND U8426 ( .A(n8195), .B(n8194), .Z(n8285) );
  XOR U8427 ( .A(n8284), .B(n8285), .Z(n8287) );
  NAND U8428 ( .A(a[96]), .B(b[15]), .Z(n8286) );
  XOR U8429 ( .A(n8287), .B(n8286), .Z(n8305) );
  NAND U8430 ( .A(n19722), .B(n8196), .Z(n8198) );
  XNOR U8431 ( .A(b[5]), .B(n8967), .Z(n8296) );
  NANDN U8432 ( .A(n19640), .B(n8296), .Z(n8197) );
  NAND U8433 ( .A(n8198), .B(n8197), .Z(n8281) );
  XNOR U8434 ( .A(n19714), .B(n8838), .Z(n8299) );
  NANDN U8435 ( .A(n8299), .B(n19766), .Z(n8201) );
  NANDN U8436 ( .A(n8199), .B(n19767), .Z(n8200) );
  NAND U8437 ( .A(n8201), .B(n8200), .Z(n8278) );
  NAND U8438 ( .A(n19554), .B(n8202), .Z(n8204) );
  IV U8439 ( .A(a[110]), .Z(n9123) );
  XNOR U8440 ( .A(b[3]), .B(n9123), .Z(n8302) );
  NANDN U8441 ( .A(n19521), .B(n8302), .Z(n8203) );
  AND U8442 ( .A(n8204), .B(n8203), .Z(n8279) );
  XNOR U8443 ( .A(n8278), .B(n8279), .Z(n8280) );
  XOR U8444 ( .A(n8281), .B(n8280), .Z(n8306) );
  XOR U8445 ( .A(n8305), .B(n8306), .Z(n8307) );
  XNOR U8446 ( .A(n8308), .B(n8307), .Z(n8256) );
  NAND U8447 ( .A(n8206), .B(n8205), .Z(n8210) );
  NAND U8448 ( .A(n8208), .B(n8207), .Z(n8209) );
  NAND U8449 ( .A(n8210), .B(n8209), .Z(n8257) );
  XOR U8450 ( .A(n8256), .B(n8257), .Z(n8259) );
  XNOR U8451 ( .A(n20052), .B(n8499), .Z(n8262) );
  OR U8452 ( .A(n8262), .B(n20020), .Z(n8213) );
  NANDN U8453 ( .A(n8211), .B(n19960), .Z(n8212) );
  NAND U8454 ( .A(n8213), .B(n8212), .Z(n8275) );
  XNOR U8455 ( .A(n102), .B(n8214), .Z(n8266) );
  OR U8456 ( .A(n8266), .B(n20121), .Z(n8217) );
  NANDN U8457 ( .A(n8215), .B(n20122), .Z(n8216) );
  NAND U8458 ( .A(n8217), .B(n8216), .Z(n8272) );
  XNOR U8459 ( .A(n19975), .B(n8682), .Z(n8269) );
  NANDN U8460 ( .A(n8269), .B(n19883), .Z(n8220) );
  NANDN U8461 ( .A(n8218), .B(n19937), .Z(n8219) );
  AND U8462 ( .A(n8220), .B(n8219), .Z(n8273) );
  XNOR U8463 ( .A(n8272), .B(n8273), .Z(n8274) );
  XNOR U8464 ( .A(n8275), .B(n8274), .Z(n8311) );
  NANDN U8465 ( .A(n8222), .B(n8221), .Z(n8226) );
  NAND U8466 ( .A(n8224), .B(n8223), .Z(n8225) );
  NAND U8467 ( .A(n8226), .B(n8225), .Z(n8312) );
  XNOR U8468 ( .A(n8311), .B(n8312), .Z(n8313) );
  NANDN U8469 ( .A(n8228), .B(n8227), .Z(n8232) );
  NAND U8470 ( .A(n8230), .B(n8229), .Z(n8231) );
  AND U8471 ( .A(n8232), .B(n8231), .Z(n8314) );
  XNOR U8472 ( .A(n8313), .B(n8314), .Z(n8258) );
  XNOR U8473 ( .A(n8259), .B(n8258), .Z(n8317) );
  NANDN U8474 ( .A(n8234), .B(n8233), .Z(n8238) );
  NAND U8475 ( .A(n8236), .B(n8235), .Z(n8237) );
  NAND U8476 ( .A(n8238), .B(n8237), .Z(n8318) );
  XNOR U8477 ( .A(n8317), .B(n8318), .Z(n8319) );
  XOR U8478 ( .A(n8320), .B(n8319), .Z(n8250) );
  NANDN U8479 ( .A(n8240), .B(n8239), .Z(n8244) );
  NANDN U8480 ( .A(n8242), .B(n8241), .Z(n8243) );
  NAND U8481 ( .A(n8244), .B(n8243), .Z(n8251) );
  XNOR U8482 ( .A(n8250), .B(n8251), .Z(n8252) );
  XNOR U8483 ( .A(n8253), .B(n8252), .Z(n8323) );
  XNOR U8484 ( .A(n8323), .B(sreg[352]), .Z(n8325) );
  NAND U8485 ( .A(n8245), .B(sreg[351]), .Z(n8249) );
  OR U8486 ( .A(n8247), .B(n8246), .Z(n8248) );
  AND U8487 ( .A(n8249), .B(n8248), .Z(n8324) );
  XOR U8488 ( .A(n8325), .B(n8324), .Z(c[352]) );
  NANDN U8489 ( .A(n8251), .B(n8250), .Z(n8255) );
  NAND U8490 ( .A(n8253), .B(n8252), .Z(n8254) );
  NAND U8491 ( .A(n8255), .B(n8254), .Z(n8331) );
  NANDN U8492 ( .A(n8257), .B(n8256), .Z(n8261) );
  OR U8493 ( .A(n8259), .B(n8258), .Z(n8260) );
  NAND U8494 ( .A(n8261), .B(n8260), .Z(n8398) );
  XNOR U8495 ( .A(n20052), .B(n8577), .Z(n8340) );
  OR U8496 ( .A(n8340), .B(n20020), .Z(n8264) );
  NANDN U8497 ( .A(n8262), .B(n19960), .Z(n8263) );
  NAND U8498 ( .A(n8264), .B(n8263), .Z(n8353) );
  XNOR U8499 ( .A(n102), .B(n8265), .Z(n8344) );
  OR U8500 ( .A(n8344), .B(n20121), .Z(n8268) );
  NANDN U8501 ( .A(n8266), .B(n20122), .Z(n8267) );
  NAND U8502 ( .A(n8268), .B(n8267), .Z(n8350) );
  XNOR U8503 ( .A(n19975), .B(n8733), .Z(n8347) );
  NANDN U8504 ( .A(n8347), .B(n19883), .Z(n8271) );
  NANDN U8505 ( .A(n8269), .B(n19937), .Z(n8270) );
  AND U8506 ( .A(n8271), .B(n8270), .Z(n8351) );
  XNOR U8507 ( .A(n8350), .B(n8351), .Z(n8352) );
  XNOR U8508 ( .A(n8353), .B(n8352), .Z(n8389) );
  NANDN U8509 ( .A(n8273), .B(n8272), .Z(n8277) );
  NAND U8510 ( .A(n8275), .B(n8274), .Z(n8276) );
  NAND U8511 ( .A(n8277), .B(n8276), .Z(n8390) );
  XNOR U8512 ( .A(n8389), .B(n8390), .Z(n8391) );
  NANDN U8513 ( .A(n8279), .B(n8278), .Z(n8283) );
  NAND U8514 ( .A(n8281), .B(n8280), .Z(n8282) );
  AND U8515 ( .A(n8283), .B(n8282), .Z(n8392) );
  XNOR U8516 ( .A(n8391), .B(n8392), .Z(n8336) );
  NANDN U8517 ( .A(n8285), .B(n8284), .Z(n8289) );
  OR U8518 ( .A(n8287), .B(n8286), .Z(n8288) );
  NAND U8519 ( .A(n8289), .B(n8288), .Z(n8386) );
  XNOR U8520 ( .A(n20154), .B(n8448), .Z(n8371) );
  OR U8521 ( .A(n8371), .B(n20057), .Z(n8292) );
  NANDN U8522 ( .A(n8290), .B(n20098), .Z(n8291) );
  AND U8523 ( .A(n8292), .B(n8291), .Z(n8363) );
  NAND U8524 ( .A(b[0]), .B(a[113]), .Z(n8293) );
  XNOR U8525 ( .A(b[1]), .B(n8293), .Z(n8295) );
  NAND U8526 ( .A(a[112]), .B(n98), .Z(n8294) );
  AND U8527 ( .A(n8295), .B(n8294), .Z(n8362) );
  XOR U8528 ( .A(n8363), .B(n8362), .Z(n8365) );
  NAND U8529 ( .A(a[97]), .B(b[15]), .Z(n8364) );
  XOR U8530 ( .A(n8365), .B(n8364), .Z(n8383) );
  NAND U8531 ( .A(n19722), .B(n8296), .Z(n8298) );
  XNOR U8532 ( .A(b[5]), .B(n9045), .Z(n8374) );
  NANDN U8533 ( .A(n19640), .B(n8374), .Z(n8297) );
  NAND U8534 ( .A(n8298), .B(n8297), .Z(n8359) );
  XNOR U8535 ( .A(n19714), .B(n8916), .Z(n8377) );
  NANDN U8536 ( .A(n8377), .B(n19766), .Z(n8301) );
  NANDN U8537 ( .A(n8299), .B(n19767), .Z(n8300) );
  NAND U8538 ( .A(n8301), .B(n8300), .Z(n8356) );
  NAND U8539 ( .A(n19554), .B(n8302), .Z(n8304) );
  IV U8540 ( .A(a[111]), .Z(n9201) );
  XNOR U8541 ( .A(b[3]), .B(n9201), .Z(n8380) );
  NANDN U8542 ( .A(n19521), .B(n8380), .Z(n8303) );
  AND U8543 ( .A(n8304), .B(n8303), .Z(n8357) );
  XNOR U8544 ( .A(n8356), .B(n8357), .Z(n8358) );
  XOR U8545 ( .A(n8359), .B(n8358), .Z(n8384) );
  XOR U8546 ( .A(n8383), .B(n8384), .Z(n8385) );
  XNOR U8547 ( .A(n8386), .B(n8385), .Z(n8334) );
  NAND U8548 ( .A(n8306), .B(n8305), .Z(n8310) );
  NAND U8549 ( .A(n8308), .B(n8307), .Z(n8309) );
  NAND U8550 ( .A(n8310), .B(n8309), .Z(n8335) );
  XOR U8551 ( .A(n8334), .B(n8335), .Z(n8337) );
  XNOR U8552 ( .A(n8336), .B(n8337), .Z(n8395) );
  NANDN U8553 ( .A(n8312), .B(n8311), .Z(n8316) );
  NAND U8554 ( .A(n8314), .B(n8313), .Z(n8315) );
  NAND U8555 ( .A(n8316), .B(n8315), .Z(n8396) );
  XNOR U8556 ( .A(n8395), .B(n8396), .Z(n8397) );
  XOR U8557 ( .A(n8398), .B(n8397), .Z(n8328) );
  NANDN U8558 ( .A(n8318), .B(n8317), .Z(n8322) );
  NANDN U8559 ( .A(n8320), .B(n8319), .Z(n8321) );
  NAND U8560 ( .A(n8322), .B(n8321), .Z(n8329) );
  XNOR U8561 ( .A(n8328), .B(n8329), .Z(n8330) );
  XNOR U8562 ( .A(n8331), .B(n8330), .Z(n8401) );
  XNOR U8563 ( .A(n8401), .B(sreg[353]), .Z(n8403) );
  NAND U8564 ( .A(n8323), .B(sreg[352]), .Z(n8327) );
  OR U8565 ( .A(n8325), .B(n8324), .Z(n8326) );
  AND U8566 ( .A(n8327), .B(n8326), .Z(n8402) );
  XOR U8567 ( .A(n8403), .B(n8402), .Z(c[353]) );
  NANDN U8568 ( .A(n8329), .B(n8328), .Z(n8333) );
  NAND U8569 ( .A(n8331), .B(n8330), .Z(n8332) );
  NAND U8570 ( .A(n8333), .B(n8332), .Z(n8409) );
  NANDN U8571 ( .A(n8335), .B(n8334), .Z(n8339) );
  OR U8572 ( .A(n8337), .B(n8336), .Z(n8338) );
  NAND U8573 ( .A(n8339), .B(n8338), .Z(n8476) );
  XNOR U8574 ( .A(n20052), .B(n8682), .Z(n8445) );
  OR U8575 ( .A(n8445), .B(n20020), .Z(n8342) );
  NANDN U8576 ( .A(n8340), .B(n19960), .Z(n8341) );
  NAND U8577 ( .A(n8342), .B(n8341), .Z(n8458) );
  XNOR U8578 ( .A(n102), .B(n8343), .Z(n8449) );
  OR U8579 ( .A(n8449), .B(n20121), .Z(n8346) );
  NANDN U8580 ( .A(n8344), .B(n20122), .Z(n8345) );
  NAND U8581 ( .A(n8346), .B(n8345), .Z(n8455) );
  XNOR U8582 ( .A(n19975), .B(n8838), .Z(n8452) );
  NANDN U8583 ( .A(n8452), .B(n19883), .Z(n8349) );
  NANDN U8584 ( .A(n8347), .B(n19937), .Z(n8348) );
  AND U8585 ( .A(n8349), .B(n8348), .Z(n8456) );
  XNOR U8586 ( .A(n8455), .B(n8456), .Z(n8457) );
  XNOR U8587 ( .A(n8458), .B(n8457), .Z(n8467) );
  NANDN U8588 ( .A(n8351), .B(n8350), .Z(n8355) );
  NAND U8589 ( .A(n8353), .B(n8352), .Z(n8354) );
  NAND U8590 ( .A(n8355), .B(n8354), .Z(n8468) );
  XNOR U8591 ( .A(n8467), .B(n8468), .Z(n8469) );
  NANDN U8592 ( .A(n8357), .B(n8356), .Z(n8361) );
  NAND U8593 ( .A(n8359), .B(n8358), .Z(n8360) );
  AND U8594 ( .A(n8361), .B(n8360), .Z(n8470) );
  XNOR U8595 ( .A(n8469), .B(n8470), .Z(n8414) );
  NANDN U8596 ( .A(n8363), .B(n8362), .Z(n8367) );
  OR U8597 ( .A(n8365), .B(n8364), .Z(n8366) );
  NAND U8598 ( .A(n8367), .B(n8366), .Z(n8442) );
  NAND U8599 ( .A(b[0]), .B(a[114]), .Z(n8368) );
  XNOR U8600 ( .A(b[1]), .B(n8368), .Z(n8370) );
  NAND U8601 ( .A(a[113]), .B(n98), .Z(n8369) );
  AND U8602 ( .A(n8370), .B(n8369), .Z(n8418) );
  XNOR U8603 ( .A(n20154), .B(n8499), .Z(n8427) );
  OR U8604 ( .A(n8427), .B(n20057), .Z(n8373) );
  NANDN U8605 ( .A(n8371), .B(n20098), .Z(n8372) );
  AND U8606 ( .A(n8373), .B(n8372), .Z(n8419) );
  XOR U8607 ( .A(n8418), .B(n8419), .Z(n8421) );
  NAND U8608 ( .A(a[98]), .B(b[15]), .Z(n8420) );
  XOR U8609 ( .A(n8421), .B(n8420), .Z(n8439) );
  NAND U8610 ( .A(n19722), .B(n8374), .Z(n8376) );
  XNOR U8611 ( .A(b[5]), .B(n9123), .Z(n8430) );
  NANDN U8612 ( .A(n19640), .B(n8430), .Z(n8375) );
  NAND U8613 ( .A(n8376), .B(n8375), .Z(n8464) );
  XNOR U8614 ( .A(n19714), .B(n8967), .Z(n8433) );
  NANDN U8615 ( .A(n8433), .B(n19766), .Z(n8379) );
  NANDN U8616 ( .A(n8377), .B(n19767), .Z(n8378) );
  NAND U8617 ( .A(n8379), .B(n8378), .Z(n8461) );
  NAND U8618 ( .A(n19554), .B(n8380), .Z(n8382) );
  IV U8619 ( .A(a[112]), .Z(n9279) );
  XNOR U8620 ( .A(b[3]), .B(n9279), .Z(n8436) );
  NANDN U8621 ( .A(n19521), .B(n8436), .Z(n8381) );
  AND U8622 ( .A(n8382), .B(n8381), .Z(n8462) );
  XNOR U8623 ( .A(n8461), .B(n8462), .Z(n8463) );
  XOR U8624 ( .A(n8464), .B(n8463), .Z(n8440) );
  XOR U8625 ( .A(n8439), .B(n8440), .Z(n8441) );
  XNOR U8626 ( .A(n8442), .B(n8441), .Z(n8412) );
  NAND U8627 ( .A(n8384), .B(n8383), .Z(n8388) );
  NAND U8628 ( .A(n8386), .B(n8385), .Z(n8387) );
  NAND U8629 ( .A(n8388), .B(n8387), .Z(n8413) );
  XOR U8630 ( .A(n8412), .B(n8413), .Z(n8415) );
  XNOR U8631 ( .A(n8414), .B(n8415), .Z(n8473) );
  NANDN U8632 ( .A(n8390), .B(n8389), .Z(n8394) );
  NAND U8633 ( .A(n8392), .B(n8391), .Z(n8393) );
  NAND U8634 ( .A(n8394), .B(n8393), .Z(n8474) );
  XNOR U8635 ( .A(n8473), .B(n8474), .Z(n8475) );
  XOR U8636 ( .A(n8476), .B(n8475), .Z(n8406) );
  NANDN U8637 ( .A(n8396), .B(n8395), .Z(n8400) );
  NANDN U8638 ( .A(n8398), .B(n8397), .Z(n8399) );
  NAND U8639 ( .A(n8400), .B(n8399), .Z(n8407) );
  XNOR U8640 ( .A(n8406), .B(n8407), .Z(n8408) );
  XNOR U8641 ( .A(n8409), .B(n8408), .Z(n8479) );
  XNOR U8642 ( .A(n8479), .B(sreg[354]), .Z(n8481) );
  NAND U8643 ( .A(n8401), .B(sreg[353]), .Z(n8405) );
  OR U8644 ( .A(n8403), .B(n8402), .Z(n8404) );
  AND U8645 ( .A(n8405), .B(n8404), .Z(n8480) );
  XOR U8646 ( .A(n8481), .B(n8480), .Z(c[354]) );
  NANDN U8647 ( .A(n8407), .B(n8406), .Z(n8411) );
  NAND U8648 ( .A(n8409), .B(n8408), .Z(n8410) );
  NAND U8649 ( .A(n8411), .B(n8410), .Z(n8487) );
  NANDN U8650 ( .A(n8413), .B(n8412), .Z(n8417) );
  OR U8651 ( .A(n8415), .B(n8414), .Z(n8416) );
  NAND U8652 ( .A(n8417), .B(n8416), .Z(n8554) );
  NANDN U8653 ( .A(n8419), .B(n8418), .Z(n8423) );
  OR U8654 ( .A(n8421), .B(n8420), .Z(n8422) );
  NAND U8655 ( .A(n8423), .B(n8422), .Z(n8542) );
  NAND U8656 ( .A(b[0]), .B(a[115]), .Z(n8424) );
  XNOR U8657 ( .A(b[1]), .B(n8424), .Z(n8426) );
  NAND U8658 ( .A(a[114]), .B(n98), .Z(n8425) );
  AND U8659 ( .A(n8426), .B(n8425), .Z(n8518) );
  XNOR U8660 ( .A(n20154), .B(n8577), .Z(n8524) );
  OR U8661 ( .A(n8524), .B(n20057), .Z(n8429) );
  NANDN U8662 ( .A(n8427), .B(n20098), .Z(n8428) );
  AND U8663 ( .A(n8429), .B(n8428), .Z(n8519) );
  XOR U8664 ( .A(n8518), .B(n8519), .Z(n8521) );
  NAND U8665 ( .A(a[99]), .B(b[15]), .Z(n8520) );
  XOR U8666 ( .A(n8521), .B(n8520), .Z(n8539) );
  NAND U8667 ( .A(n19722), .B(n8430), .Z(n8432) );
  XNOR U8668 ( .A(b[5]), .B(n9201), .Z(n8530) );
  NANDN U8669 ( .A(n19640), .B(n8530), .Z(n8431) );
  NAND U8670 ( .A(n8432), .B(n8431), .Z(n8515) );
  XNOR U8671 ( .A(n19714), .B(n9045), .Z(n8533) );
  NANDN U8672 ( .A(n8533), .B(n19766), .Z(n8435) );
  NANDN U8673 ( .A(n8433), .B(n19767), .Z(n8434) );
  NAND U8674 ( .A(n8435), .B(n8434), .Z(n8512) );
  NAND U8675 ( .A(n19554), .B(n8436), .Z(n8438) );
  IV U8676 ( .A(a[113]), .Z(n9357) );
  XNOR U8677 ( .A(b[3]), .B(n9357), .Z(n8536) );
  NANDN U8678 ( .A(n19521), .B(n8536), .Z(n8437) );
  AND U8679 ( .A(n8438), .B(n8437), .Z(n8513) );
  XNOR U8680 ( .A(n8512), .B(n8513), .Z(n8514) );
  XOR U8681 ( .A(n8515), .B(n8514), .Z(n8540) );
  XOR U8682 ( .A(n8539), .B(n8540), .Z(n8541) );
  XNOR U8683 ( .A(n8542), .B(n8541), .Z(n8490) );
  NAND U8684 ( .A(n8440), .B(n8439), .Z(n8444) );
  NAND U8685 ( .A(n8442), .B(n8441), .Z(n8443) );
  NAND U8686 ( .A(n8444), .B(n8443), .Z(n8491) );
  XOR U8687 ( .A(n8490), .B(n8491), .Z(n8493) );
  XNOR U8688 ( .A(n20052), .B(n8733), .Z(n8496) );
  OR U8689 ( .A(n8496), .B(n20020), .Z(n8447) );
  NANDN U8690 ( .A(n8445), .B(n19960), .Z(n8446) );
  NAND U8691 ( .A(n8447), .B(n8446), .Z(n8509) );
  XNOR U8692 ( .A(n102), .B(n8448), .Z(n8500) );
  OR U8693 ( .A(n8500), .B(n20121), .Z(n8451) );
  NANDN U8694 ( .A(n8449), .B(n20122), .Z(n8450) );
  NAND U8695 ( .A(n8451), .B(n8450), .Z(n8506) );
  XNOR U8696 ( .A(n19975), .B(n8916), .Z(n8503) );
  NANDN U8697 ( .A(n8503), .B(n19883), .Z(n8454) );
  NANDN U8698 ( .A(n8452), .B(n19937), .Z(n8453) );
  AND U8699 ( .A(n8454), .B(n8453), .Z(n8507) );
  XNOR U8700 ( .A(n8506), .B(n8507), .Z(n8508) );
  XNOR U8701 ( .A(n8509), .B(n8508), .Z(n8545) );
  NANDN U8702 ( .A(n8456), .B(n8455), .Z(n8460) );
  NAND U8703 ( .A(n8458), .B(n8457), .Z(n8459) );
  NAND U8704 ( .A(n8460), .B(n8459), .Z(n8546) );
  XNOR U8705 ( .A(n8545), .B(n8546), .Z(n8547) );
  NANDN U8706 ( .A(n8462), .B(n8461), .Z(n8466) );
  NAND U8707 ( .A(n8464), .B(n8463), .Z(n8465) );
  AND U8708 ( .A(n8466), .B(n8465), .Z(n8548) );
  XNOR U8709 ( .A(n8547), .B(n8548), .Z(n8492) );
  XNOR U8710 ( .A(n8493), .B(n8492), .Z(n8551) );
  NANDN U8711 ( .A(n8468), .B(n8467), .Z(n8472) );
  NAND U8712 ( .A(n8470), .B(n8469), .Z(n8471) );
  NAND U8713 ( .A(n8472), .B(n8471), .Z(n8552) );
  XNOR U8714 ( .A(n8551), .B(n8552), .Z(n8553) );
  XOR U8715 ( .A(n8554), .B(n8553), .Z(n8484) );
  NANDN U8716 ( .A(n8474), .B(n8473), .Z(n8478) );
  NANDN U8717 ( .A(n8476), .B(n8475), .Z(n8477) );
  NAND U8718 ( .A(n8478), .B(n8477), .Z(n8485) );
  XNOR U8719 ( .A(n8484), .B(n8485), .Z(n8486) );
  XNOR U8720 ( .A(n8487), .B(n8486), .Z(n8557) );
  XNOR U8721 ( .A(n8557), .B(sreg[355]), .Z(n8559) );
  NAND U8722 ( .A(n8479), .B(sreg[354]), .Z(n8483) );
  OR U8723 ( .A(n8481), .B(n8480), .Z(n8482) );
  AND U8724 ( .A(n8483), .B(n8482), .Z(n8558) );
  XOR U8725 ( .A(n8559), .B(n8558), .Z(c[355]) );
  NANDN U8726 ( .A(n8485), .B(n8484), .Z(n8489) );
  NAND U8727 ( .A(n8487), .B(n8486), .Z(n8488) );
  NAND U8728 ( .A(n8489), .B(n8488), .Z(n8565) );
  NANDN U8729 ( .A(n8491), .B(n8490), .Z(n8495) );
  OR U8730 ( .A(n8493), .B(n8492), .Z(n8494) );
  NAND U8731 ( .A(n8495), .B(n8494), .Z(n8632) );
  XNOR U8732 ( .A(n20052), .B(n8838), .Z(n8574) );
  OR U8733 ( .A(n8574), .B(n20020), .Z(n8498) );
  NANDN U8734 ( .A(n8496), .B(n19960), .Z(n8497) );
  NAND U8735 ( .A(n8498), .B(n8497), .Z(n8587) );
  XNOR U8736 ( .A(n102), .B(n8499), .Z(n8578) );
  OR U8737 ( .A(n8578), .B(n20121), .Z(n8502) );
  NANDN U8738 ( .A(n8500), .B(n20122), .Z(n8501) );
  NAND U8739 ( .A(n8502), .B(n8501), .Z(n8584) );
  XNOR U8740 ( .A(n19975), .B(n8967), .Z(n8581) );
  NANDN U8741 ( .A(n8581), .B(n19883), .Z(n8505) );
  NANDN U8742 ( .A(n8503), .B(n19937), .Z(n8504) );
  AND U8743 ( .A(n8505), .B(n8504), .Z(n8585) );
  XNOR U8744 ( .A(n8584), .B(n8585), .Z(n8586) );
  XNOR U8745 ( .A(n8587), .B(n8586), .Z(n8623) );
  NANDN U8746 ( .A(n8507), .B(n8506), .Z(n8511) );
  NAND U8747 ( .A(n8509), .B(n8508), .Z(n8510) );
  NAND U8748 ( .A(n8511), .B(n8510), .Z(n8624) );
  XNOR U8749 ( .A(n8623), .B(n8624), .Z(n8625) );
  NANDN U8750 ( .A(n8513), .B(n8512), .Z(n8517) );
  NAND U8751 ( .A(n8515), .B(n8514), .Z(n8516) );
  AND U8752 ( .A(n8517), .B(n8516), .Z(n8626) );
  XNOR U8753 ( .A(n8625), .B(n8626), .Z(n8570) );
  NANDN U8754 ( .A(n8519), .B(n8518), .Z(n8523) );
  OR U8755 ( .A(n8521), .B(n8520), .Z(n8522) );
  NAND U8756 ( .A(n8523), .B(n8522), .Z(n8620) );
  XNOR U8757 ( .A(n20154), .B(n8682), .Z(n8602) );
  OR U8758 ( .A(n8602), .B(n20057), .Z(n8526) );
  NANDN U8759 ( .A(n8524), .B(n20098), .Z(n8525) );
  AND U8760 ( .A(n8526), .B(n8525), .Z(n8597) );
  NAND U8761 ( .A(b[0]), .B(a[116]), .Z(n8527) );
  XNOR U8762 ( .A(b[1]), .B(n8527), .Z(n8529) );
  NAND U8763 ( .A(a[115]), .B(n98), .Z(n8528) );
  AND U8764 ( .A(n8529), .B(n8528), .Z(n8596) );
  XOR U8765 ( .A(n8597), .B(n8596), .Z(n8599) );
  NAND U8766 ( .A(a[100]), .B(b[15]), .Z(n8598) );
  XOR U8767 ( .A(n8599), .B(n8598), .Z(n8617) );
  NAND U8768 ( .A(n19722), .B(n8530), .Z(n8532) );
  XNOR U8769 ( .A(b[5]), .B(n9279), .Z(n8608) );
  NANDN U8770 ( .A(n19640), .B(n8608), .Z(n8531) );
  NAND U8771 ( .A(n8532), .B(n8531), .Z(n8593) );
  XNOR U8772 ( .A(n19714), .B(n9123), .Z(n8611) );
  NANDN U8773 ( .A(n8611), .B(n19766), .Z(n8535) );
  NANDN U8774 ( .A(n8533), .B(n19767), .Z(n8534) );
  NAND U8775 ( .A(n8535), .B(n8534), .Z(n8590) );
  NAND U8776 ( .A(n19554), .B(n8536), .Z(n8538) );
  IV U8777 ( .A(a[114]), .Z(n9435) );
  XNOR U8778 ( .A(b[3]), .B(n9435), .Z(n8614) );
  NANDN U8779 ( .A(n19521), .B(n8614), .Z(n8537) );
  AND U8780 ( .A(n8538), .B(n8537), .Z(n8591) );
  XNOR U8781 ( .A(n8590), .B(n8591), .Z(n8592) );
  XOR U8782 ( .A(n8593), .B(n8592), .Z(n8618) );
  XOR U8783 ( .A(n8617), .B(n8618), .Z(n8619) );
  XNOR U8784 ( .A(n8620), .B(n8619), .Z(n8568) );
  NAND U8785 ( .A(n8540), .B(n8539), .Z(n8544) );
  NAND U8786 ( .A(n8542), .B(n8541), .Z(n8543) );
  NAND U8787 ( .A(n8544), .B(n8543), .Z(n8569) );
  XOR U8788 ( .A(n8568), .B(n8569), .Z(n8571) );
  XNOR U8789 ( .A(n8570), .B(n8571), .Z(n8629) );
  NANDN U8790 ( .A(n8546), .B(n8545), .Z(n8550) );
  NAND U8791 ( .A(n8548), .B(n8547), .Z(n8549) );
  NAND U8792 ( .A(n8550), .B(n8549), .Z(n8630) );
  XNOR U8793 ( .A(n8629), .B(n8630), .Z(n8631) );
  XOR U8794 ( .A(n8632), .B(n8631), .Z(n8562) );
  NANDN U8795 ( .A(n8552), .B(n8551), .Z(n8556) );
  NANDN U8796 ( .A(n8554), .B(n8553), .Z(n8555) );
  NAND U8797 ( .A(n8556), .B(n8555), .Z(n8563) );
  XNOR U8798 ( .A(n8562), .B(n8563), .Z(n8564) );
  XNOR U8799 ( .A(n8565), .B(n8564), .Z(n8635) );
  XNOR U8800 ( .A(n8635), .B(sreg[356]), .Z(n8637) );
  NAND U8801 ( .A(n8557), .B(sreg[355]), .Z(n8561) );
  OR U8802 ( .A(n8559), .B(n8558), .Z(n8560) );
  AND U8803 ( .A(n8561), .B(n8560), .Z(n8636) );
  XOR U8804 ( .A(n8637), .B(n8636), .Z(c[356]) );
  NANDN U8805 ( .A(n8563), .B(n8562), .Z(n8567) );
  NAND U8806 ( .A(n8565), .B(n8564), .Z(n8566) );
  NAND U8807 ( .A(n8567), .B(n8566), .Z(n8643) );
  NANDN U8808 ( .A(n8569), .B(n8568), .Z(n8573) );
  OR U8809 ( .A(n8571), .B(n8570), .Z(n8572) );
  NAND U8810 ( .A(n8573), .B(n8572), .Z(n8710) );
  XNOR U8811 ( .A(n20052), .B(n8916), .Z(n8679) );
  OR U8812 ( .A(n8679), .B(n20020), .Z(n8576) );
  NANDN U8813 ( .A(n8574), .B(n19960), .Z(n8575) );
  NAND U8814 ( .A(n8576), .B(n8575), .Z(n8692) );
  XNOR U8815 ( .A(n102), .B(n8577), .Z(n8683) );
  OR U8816 ( .A(n8683), .B(n20121), .Z(n8580) );
  NANDN U8817 ( .A(n8578), .B(n20122), .Z(n8579) );
  NAND U8818 ( .A(n8580), .B(n8579), .Z(n8689) );
  XNOR U8819 ( .A(n19975), .B(n9045), .Z(n8686) );
  NANDN U8820 ( .A(n8686), .B(n19883), .Z(n8583) );
  NANDN U8821 ( .A(n8581), .B(n19937), .Z(n8582) );
  AND U8822 ( .A(n8583), .B(n8582), .Z(n8690) );
  XNOR U8823 ( .A(n8689), .B(n8690), .Z(n8691) );
  XNOR U8824 ( .A(n8692), .B(n8691), .Z(n8701) );
  NANDN U8825 ( .A(n8585), .B(n8584), .Z(n8589) );
  NAND U8826 ( .A(n8587), .B(n8586), .Z(n8588) );
  NAND U8827 ( .A(n8589), .B(n8588), .Z(n8702) );
  XNOR U8828 ( .A(n8701), .B(n8702), .Z(n8703) );
  NANDN U8829 ( .A(n8591), .B(n8590), .Z(n8595) );
  NAND U8830 ( .A(n8593), .B(n8592), .Z(n8594) );
  AND U8831 ( .A(n8595), .B(n8594), .Z(n8704) );
  XNOR U8832 ( .A(n8703), .B(n8704), .Z(n8648) );
  NANDN U8833 ( .A(n8597), .B(n8596), .Z(n8601) );
  OR U8834 ( .A(n8599), .B(n8598), .Z(n8600) );
  NAND U8835 ( .A(n8601), .B(n8600), .Z(n8676) );
  XNOR U8836 ( .A(n20154), .B(n8733), .Z(n8661) );
  OR U8837 ( .A(n8661), .B(n20057), .Z(n8604) );
  NANDN U8838 ( .A(n8602), .B(n20098), .Z(n8603) );
  AND U8839 ( .A(n8604), .B(n8603), .Z(n8653) );
  NAND U8840 ( .A(b[0]), .B(a[117]), .Z(n8605) );
  XNOR U8841 ( .A(b[1]), .B(n8605), .Z(n8607) );
  NAND U8842 ( .A(a[116]), .B(n98), .Z(n8606) );
  AND U8843 ( .A(n8607), .B(n8606), .Z(n8652) );
  XOR U8844 ( .A(n8653), .B(n8652), .Z(n8655) );
  NAND U8845 ( .A(a[101]), .B(b[15]), .Z(n8654) );
  XOR U8846 ( .A(n8655), .B(n8654), .Z(n8673) );
  NAND U8847 ( .A(n19722), .B(n8608), .Z(n8610) );
  XNOR U8848 ( .A(b[5]), .B(n9357), .Z(n8664) );
  NANDN U8849 ( .A(n19640), .B(n8664), .Z(n8609) );
  NAND U8850 ( .A(n8610), .B(n8609), .Z(n8698) );
  XNOR U8851 ( .A(n19714), .B(n9201), .Z(n8667) );
  NANDN U8852 ( .A(n8667), .B(n19766), .Z(n8613) );
  NANDN U8853 ( .A(n8611), .B(n19767), .Z(n8612) );
  NAND U8854 ( .A(n8613), .B(n8612), .Z(n8695) );
  NAND U8855 ( .A(n19554), .B(n8614), .Z(n8616) );
  IV U8856 ( .A(a[115]), .Z(n9513) );
  XNOR U8857 ( .A(b[3]), .B(n9513), .Z(n8670) );
  NANDN U8858 ( .A(n19521), .B(n8670), .Z(n8615) );
  AND U8859 ( .A(n8616), .B(n8615), .Z(n8696) );
  XNOR U8860 ( .A(n8695), .B(n8696), .Z(n8697) );
  XOR U8861 ( .A(n8698), .B(n8697), .Z(n8674) );
  XOR U8862 ( .A(n8673), .B(n8674), .Z(n8675) );
  XNOR U8863 ( .A(n8676), .B(n8675), .Z(n8646) );
  NAND U8864 ( .A(n8618), .B(n8617), .Z(n8622) );
  NAND U8865 ( .A(n8620), .B(n8619), .Z(n8621) );
  NAND U8866 ( .A(n8622), .B(n8621), .Z(n8647) );
  XOR U8867 ( .A(n8646), .B(n8647), .Z(n8649) );
  XNOR U8868 ( .A(n8648), .B(n8649), .Z(n8707) );
  NANDN U8869 ( .A(n8624), .B(n8623), .Z(n8628) );
  NAND U8870 ( .A(n8626), .B(n8625), .Z(n8627) );
  NAND U8871 ( .A(n8628), .B(n8627), .Z(n8708) );
  XNOR U8872 ( .A(n8707), .B(n8708), .Z(n8709) );
  XOR U8873 ( .A(n8710), .B(n8709), .Z(n8640) );
  NANDN U8874 ( .A(n8630), .B(n8629), .Z(n8634) );
  NANDN U8875 ( .A(n8632), .B(n8631), .Z(n8633) );
  NAND U8876 ( .A(n8634), .B(n8633), .Z(n8641) );
  XNOR U8877 ( .A(n8640), .B(n8641), .Z(n8642) );
  XNOR U8878 ( .A(n8643), .B(n8642), .Z(n8713) );
  XNOR U8879 ( .A(n8713), .B(sreg[357]), .Z(n8715) );
  NAND U8880 ( .A(n8635), .B(sreg[356]), .Z(n8639) );
  OR U8881 ( .A(n8637), .B(n8636), .Z(n8638) );
  AND U8882 ( .A(n8639), .B(n8638), .Z(n8714) );
  XOR U8883 ( .A(n8715), .B(n8714), .Z(c[357]) );
  NANDN U8884 ( .A(n8641), .B(n8640), .Z(n8645) );
  NAND U8885 ( .A(n8643), .B(n8642), .Z(n8644) );
  NAND U8886 ( .A(n8645), .B(n8644), .Z(n8721) );
  NANDN U8887 ( .A(n8647), .B(n8646), .Z(n8651) );
  OR U8888 ( .A(n8649), .B(n8648), .Z(n8650) );
  NAND U8889 ( .A(n8651), .B(n8650), .Z(n8788) );
  NANDN U8890 ( .A(n8653), .B(n8652), .Z(n8657) );
  OR U8891 ( .A(n8655), .B(n8654), .Z(n8656) );
  NAND U8892 ( .A(n8657), .B(n8656), .Z(n8776) );
  NAND U8893 ( .A(b[0]), .B(a[118]), .Z(n8658) );
  XNOR U8894 ( .A(b[1]), .B(n8658), .Z(n8660) );
  NAND U8895 ( .A(a[117]), .B(n98), .Z(n8659) );
  AND U8896 ( .A(n8660), .B(n8659), .Z(n8752) );
  XNOR U8897 ( .A(n20154), .B(n8838), .Z(n8761) );
  OR U8898 ( .A(n8761), .B(n20057), .Z(n8663) );
  NANDN U8899 ( .A(n8661), .B(n20098), .Z(n8662) );
  AND U8900 ( .A(n8663), .B(n8662), .Z(n8753) );
  XOR U8901 ( .A(n8752), .B(n8753), .Z(n8755) );
  NAND U8902 ( .A(a[102]), .B(b[15]), .Z(n8754) );
  XOR U8903 ( .A(n8755), .B(n8754), .Z(n8773) );
  NAND U8904 ( .A(n19722), .B(n8664), .Z(n8666) );
  XNOR U8905 ( .A(b[5]), .B(n9435), .Z(n8764) );
  NANDN U8906 ( .A(n19640), .B(n8764), .Z(n8665) );
  NAND U8907 ( .A(n8666), .B(n8665), .Z(n8749) );
  XNOR U8908 ( .A(n19714), .B(n9279), .Z(n8767) );
  NANDN U8909 ( .A(n8767), .B(n19766), .Z(n8669) );
  NANDN U8910 ( .A(n8667), .B(n19767), .Z(n8668) );
  NAND U8911 ( .A(n8669), .B(n8668), .Z(n8746) );
  NAND U8912 ( .A(n19554), .B(n8670), .Z(n8672) );
  IV U8913 ( .A(a[116]), .Z(n9591) );
  XNOR U8914 ( .A(b[3]), .B(n9591), .Z(n8770) );
  NANDN U8915 ( .A(n19521), .B(n8770), .Z(n8671) );
  AND U8916 ( .A(n8672), .B(n8671), .Z(n8747) );
  XNOR U8917 ( .A(n8746), .B(n8747), .Z(n8748) );
  XOR U8918 ( .A(n8749), .B(n8748), .Z(n8774) );
  XOR U8919 ( .A(n8773), .B(n8774), .Z(n8775) );
  XNOR U8920 ( .A(n8776), .B(n8775), .Z(n8724) );
  NAND U8921 ( .A(n8674), .B(n8673), .Z(n8678) );
  NAND U8922 ( .A(n8676), .B(n8675), .Z(n8677) );
  NAND U8923 ( .A(n8678), .B(n8677), .Z(n8725) );
  XOR U8924 ( .A(n8724), .B(n8725), .Z(n8727) );
  XNOR U8925 ( .A(n20052), .B(n8967), .Z(n8730) );
  OR U8926 ( .A(n8730), .B(n20020), .Z(n8681) );
  NANDN U8927 ( .A(n8679), .B(n19960), .Z(n8680) );
  NAND U8928 ( .A(n8681), .B(n8680), .Z(n8743) );
  XNOR U8929 ( .A(n102), .B(n8682), .Z(n8734) );
  OR U8930 ( .A(n8734), .B(n20121), .Z(n8685) );
  NANDN U8931 ( .A(n8683), .B(n20122), .Z(n8684) );
  NAND U8932 ( .A(n8685), .B(n8684), .Z(n8740) );
  XNOR U8933 ( .A(n19975), .B(n9123), .Z(n8737) );
  NANDN U8934 ( .A(n8737), .B(n19883), .Z(n8688) );
  NANDN U8935 ( .A(n8686), .B(n19937), .Z(n8687) );
  AND U8936 ( .A(n8688), .B(n8687), .Z(n8741) );
  XNOR U8937 ( .A(n8740), .B(n8741), .Z(n8742) );
  XNOR U8938 ( .A(n8743), .B(n8742), .Z(n8779) );
  NANDN U8939 ( .A(n8690), .B(n8689), .Z(n8694) );
  NAND U8940 ( .A(n8692), .B(n8691), .Z(n8693) );
  NAND U8941 ( .A(n8694), .B(n8693), .Z(n8780) );
  XNOR U8942 ( .A(n8779), .B(n8780), .Z(n8781) );
  NANDN U8943 ( .A(n8696), .B(n8695), .Z(n8700) );
  NAND U8944 ( .A(n8698), .B(n8697), .Z(n8699) );
  AND U8945 ( .A(n8700), .B(n8699), .Z(n8782) );
  XNOR U8946 ( .A(n8781), .B(n8782), .Z(n8726) );
  XNOR U8947 ( .A(n8727), .B(n8726), .Z(n8785) );
  NANDN U8948 ( .A(n8702), .B(n8701), .Z(n8706) );
  NAND U8949 ( .A(n8704), .B(n8703), .Z(n8705) );
  NAND U8950 ( .A(n8706), .B(n8705), .Z(n8786) );
  XNOR U8951 ( .A(n8785), .B(n8786), .Z(n8787) );
  XOR U8952 ( .A(n8788), .B(n8787), .Z(n8718) );
  NANDN U8953 ( .A(n8708), .B(n8707), .Z(n8712) );
  NANDN U8954 ( .A(n8710), .B(n8709), .Z(n8711) );
  NAND U8955 ( .A(n8712), .B(n8711), .Z(n8719) );
  XNOR U8956 ( .A(n8718), .B(n8719), .Z(n8720) );
  XNOR U8957 ( .A(n8721), .B(n8720), .Z(n8791) );
  XNOR U8958 ( .A(n8791), .B(sreg[358]), .Z(n8793) );
  NAND U8959 ( .A(n8713), .B(sreg[357]), .Z(n8717) );
  OR U8960 ( .A(n8715), .B(n8714), .Z(n8716) );
  AND U8961 ( .A(n8717), .B(n8716), .Z(n8792) );
  XOR U8962 ( .A(n8793), .B(n8792), .Z(c[358]) );
  NANDN U8963 ( .A(n8719), .B(n8718), .Z(n8723) );
  NAND U8964 ( .A(n8721), .B(n8720), .Z(n8722) );
  NAND U8965 ( .A(n8723), .B(n8722), .Z(n8799) );
  NANDN U8966 ( .A(n8725), .B(n8724), .Z(n8729) );
  OR U8967 ( .A(n8727), .B(n8726), .Z(n8728) );
  NAND U8968 ( .A(n8729), .B(n8728), .Z(n8866) );
  XNOR U8969 ( .A(n20052), .B(n9045), .Z(n8835) );
  OR U8970 ( .A(n8835), .B(n20020), .Z(n8732) );
  NANDN U8971 ( .A(n8730), .B(n19960), .Z(n8731) );
  NAND U8972 ( .A(n8732), .B(n8731), .Z(n8848) );
  XNOR U8973 ( .A(n102), .B(n8733), .Z(n8839) );
  OR U8974 ( .A(n8839), .B(n20121), .Z(n8736) );
  NANDN U8975 ( .A(n8734), .B(n20122), .Z(n8735) );
  NAND U8976 ( .A(n8736), .B(n8735), .Z(n8845) );
  XNOR U8977 ( .A(n19975), .B(n9201), .Z(n8842) );
  NANDN U8978 ( .A(n8842), .B(n19883), .Z(n8739) );
  NANDN U8979 ( .A(n8737), .B(n19937), .Z(n8738) );
  AND U8980 ( .A(n8739), .B(n8738), .Z(n8846) );
  XNOR U8981 ( .A(n8845), .B(n8846), .Z(n8847) );
  XNOR U8982 ( .A(n8848), .B(n8847), .Z(n8857) );
  NANDN U8983 ( .A(n8741), .B(n8740), .Z(n8745) );
  NAND U8984 ( .A(n8743), .B(n8742), .Z(n8744) );
  NAND U8985 ( .A(n8745), .B(n8744), .Z(n8858) );
  XNOR U8986 ( .A(n8857), .B(n8858), .Z(n8859) );
  NANDN U8987 ( .A(n8747), .B(n8746), .Z(n8751) );
  NAND U8988 ( .A(n8749), .B(n8748), .Z(n8750) );
  AND U8989 ( .A(n8751), .B(n8750), .Z(n8860) );
  XNOR U8990 ( .A(n8859), .B(n8860), .Z(n8804) );
  NANDN U8991 ( .A(n8753), .B(n8752), .Z(n8757) );
  OR U8992 ( .A(n8755), .B(n8754), .Z(n8756) );
  NAND U8993 ( .A(n8757), .B(n8756), .Z(n8832) );
  NAND U8994 ( .A(b[0]), .B(a[119]), .Z(n8758) );
  XNOR U8995 ( .A(b[1]), .B(n8758), .Z(n8760) );
  NAND U8996 ( .A(a[118]), .B(n98), .Z(n8759) );
  AND U8997 ( .A(n8760), .B(n8759), .Z(n8808) );
  XNOR U8998 ( .A(n20154), .B(n8916), .Z(n8814) );
  OR U8999 ( .A(n8814), .B(n20057), .Z(n8763) );
  NANDN U9000 ( .A(n8761), .B(n20098), .Z(n8762) );
  AND U9001 ( .A(n8763), .B(n8762), .Z(n8809) );
  XOR U9002 ( .A(n8808), .B(n8809), .Z(n8811) );
  NAND U9003 ( .A(a[103]), .B(b[15]), .Z(n8810) );
  XOR U9004 ( .A(n8811), .B(n8810), .Z(n8829) );
  NAND U9005 ( .A(n19722), .B(n8764), .Z(n8766) );
  XNOR U9006 ( .A(b[5]), .B(n9513), .Z(n8820) );
  NANDN U9007 ( .A(n19640), .B(n8820), .Z(n8765) );
  NAND U9008 ( .A(n8766), .B(n8765), .Z(n8854) );
  XNOR U9009 ( .A(n19714), .B(n9357), .Z(n8823) );
  NANDN U9010 ( .A(n8823), .B(n19766), .Z(n8769) );
  NANDN U9011 ( .A(n8767), .B(n19767), .Z(n8768) );
  NAND U9012 ( .A(n8769), .B(n8768), .Z(n8851) );
  NAND U9013 ( .A(n19554), .B(n8770), .Z(n8772) );
  IV U9014 ( .A(a[117]), .Z(n9669) );
  XNOR U9015 ( .A(b[3]), .B(n9669), .Z(n8826) );
  NANDN U9016 ( .A(n19521), .B(n8826), .Z(n8771) );
  AND U9017 ( .A(n8772), .B(n8771), .Z(n8852) );
  XNOR U9018 ( .A(n8851), .B(n8852), .Z(n8853) );
  XOR U9019 ( .A(n8854), .B(n8853), .Z(n8830) );
  XOR U9020 ( .A(n8829), .B(n8830), .Z(n8831) );
  XNOR U9021 ( .A(n8832), .B(n8831), .Z(n8802) );
  NAND U9022 ( .A(n8774), .B(n8773), .Z(n8778) );
  NAND U9023 ( .A(n8776), .B(n8775), .Z(n8777) );
  NAND U9024 ( .A(n8778), .B(n8777), .Z(n8803) );
  XOR U9025 ( .A(n8802), .B(n8803), .Z(n8805) );
  XNOR U9026 ( .A(n8804), .B(n8805), .Z(n8863) );
  NANDN U9027 ( .A(n8780), .B(n8779), .Z(n8784) );
  NAND U9028 ( .A(n8782), .B(n8781), .Z(n8783) );
  NAND U9029 ( .A(n8784), .B(n8783), .Z(n8864) );
  XNOR U9030 ( .A(n8863), .B(n8864), .Z(n8865) );
  XOR U9031 ( .A(n8866), .B(n8865), .Z(n8796) );
  NANDN U9032 ( .A(n8786), .B(n8785), .Z(n8790) );
  NANDN U9033 ( .A(n8788), .B(n8787), .Z(n8789) );
  NAND U9034 ( .A(n8790), .B(n8789), .Z(n8797) );
  XNOR U9035 ( .A(n8796), .B(n8797), .Z(n8798) );
  XNOR U9036 ( .A(n8799), .B(n8798), .Z(n8869) );
  XNOR U9037 ( .A(n8869), .B(sreg[359]), .Z(n8871) );
  NAND U9038 ( .A(n8791), .B(sreg[358]), .Z(n8795) );
  OR U9039 ( .A(n8793), .B(n8792), .Z(n8794) );
  AND U9040 ( .A(n8795), .B(n8794), .Z(n8870) );
  XOR U9041 ( .A(n8871), .B(n8870), .Z(c[359]) );
  NANDN U9042 ( .A(n8797), .B(n8796), .Z(n8801) );
  NAND U9043 ( .A(n8799), .B(n8798), .Z(n8800) );
  NAND U9044 ( .A(n8801), .B(n8800), .Z(n8877) );
  NANDN U9045 ( .A(n8803), .B(n8802), .Z(n8807) );
  OR U9046 ( .A(n8805), .B(n8804), .Z(n8806) );
  NAND U9047 ( .A(n8807), .B(n8806), .Z(n8944) );
  NANDN U9048 ( .A(n8809), .B(n8808), .Z(n8813) );
  OR U9049 ( .A(n8811), .B(n8810), .Z(n8812) );
  NAND U9050 ( .A(n8813), .B(n8812), .Z(n8910) );
  XNOR U9051 ( .A(n20154), .B(n8967), .Z(n8892) );
  OR U9052 ( .A(n8892), .B(n20057), .Z(n8816) );
  NANDN U9053 ( .A(n8814), .B(n20098), .Z(n8815) );
  AND U9054 ( .A(n8816), .B(n8815), .Z(n8887) );
  NAND U9055 ( .A(b[0]), .B(a[120]), .Z(n8817) );
  XNOR U9056 ( .A(b[1]), .B(n8817), .Z(n8819) );
  NAND U9057 ( .A(a[119]), .B(n98), .Z(n8818) );
  AND U9058 ( .A(n8819), .B(n8818), .Z(n8886) );
  XOR U9059 ( .A(n8887), .B(n8886), .Z(n8889) );
  NAND U9060 ( .A(a[104]), .B(b[15]), .Z(n8888) );
  XOR U9061 ( .A(n8889), .B(n8888), .Z(n8907) );
  NAND U9062 ( .A(n19722), .B(n8820), .Z(n8822) );
  XNOR U9063 ( .A(b[5]), .B(n9591), .Z(n8898) );
  NANDN U9064 ( .A(n19640), .B(n8898), .Z(n8821) );
  NAND U9065 ( .A(n8822), .B(n8821), .Z(n8932) );
  XNOR U9066 ( .A(n19714), .B(n9435), .Z(n8901) );
  NANDN U9067 ( .A(n8901), .B(n19766), .Z(n8825) );
  NANDN U9068 ( .A(n8823), .B(n19767), .Z(n8824) );
  NAND U9069 ( .A(n8825), .B(n8824), .Z(n8929) );
  NAND U9070 ( .A(n19554), .B(n8826), .Z(n8828) );
  IV U9071 ( .A(a[118]), .Z(n9747) );
  XNOR U9072 ( .A(b[3]), .B(n9747), .Z(n8904) );
  NANDN U9073 ( .A(n19521), .B(n8904), .Z(n8827) );
  AND U9074 ( .A(n8828), .B(n8827), .Z(n8930) );
  XNOR U9075 ( .A(n8929), .B(n8930), .Z(n8931) );
  XOR U9076 ( .A(n8932), .B(n8931), .Z(n8908) );
  XOR U9077 ( .A(n8907), .B(n8908), .Z(n8909) );
  XNOR U9078 ( .A(n8910), .B(n8909), .Z(n8880) );
  NAND U9079 ( .A(n8830), .B(n8829), .Z(n8834) );
  NAND U9080 ( .A(n8832), .B(n8831), .Z(n8833) );
  NAND U9081 ( .A(n8834), .B(n8833), .Z(n8881) );
  XOR U9082 ( .A(n8880), .B(n8881), .Z(n8883) );
  XNOR U9083 ( .A(n20052), .B(n9123), .Z(n8913) );
  OR U9084 ( .A(n8913), .B(n20020), .Z(n8837) );
  NANDN U9085 ( .A(n8835), .B(n19960), .Z(n8836) );
  NAND U9086 ( .A(n8837), .B(n8836), .Z(n8926) );
  XNOR U9087 ( .A(n102), .B(n8838), .Z(n8917) );
  OR U9088 ( .A(n8917), .B(n20121), .Z(n8841) );
  NANDN U9089 ( .A(n8839), .B(n20122), .Z(n8840) );
  NAND U9090 ( .A(n8841), .B(n8840), .Z(n8923) );
  XNOR U9091 ( .A(n19975), .B(n9279), .Z(n8920) );
  NANDN U9092 ( .A(n8920), .B(n19883), .Z(n8844) );
  NANDN U9093 ( .A(n8842), .B(n19937), .Z(n8843) );
  AND U9094 ( .A(n8844), .B(n8843), .Z(n8924) );
  XNOR U9095 ( .A(n8923), .B(n8924), .Z(n8925) );
  XNOR U9096 ( .A(n8926), .B(n8925), .Z(n8935) );
  NANDN U9097 ( .A(n8846), .B(n8845), .Z(n8850) );
  NAND U9098 ( .A(n8848), .B(n8847), .Z(n8849) );
  NAND U9099 ( .A(n8850), .B(n8849), .Z(n8936) );
  XNOR U9100 ( .A(n8935), .B(n8936), .Z(n8937) );
  NANDN U9101 ( .A(n8852), .B(n8851), .Z(n8856) );
  NAND U9102 ( .A(n8854), .B(n8853), .Z(n8855) );
  AND U9103 ( .A(n8856), .B(n8855), .Z(n8938) );
  XNOR U9104 ( .A(n8937), .B(n8938), .Z(n8882) );
  XNOR U9105 ( .A(n8883), .B(n8882), .Z(n8941) );
  NANDN U9106 ( .A(n8858), .B(n8857), .Z(n8862) );
  NAND U9107 ( .A(n8860), .B(n8859), .Z(n8861) );
  NAND U9108 ( .A(n8862), .B(n8861), .Z(n8942) );
  XNOR U9109 ( .A(n8941), .B(n8942), .Z(n8943) );
  XOR U9110 ( .A(n8944), .B(n8943), .Z(n8874) );
  NANDN U9111 ( .A(n8864), .B(n8863), .Z(n8868) );
  NANDN U9112 ( .A(n8866), .B(n8865), .Z(n8867) );
  NAND U9113 ( .A(n8868), .B(n8867), .Z(n8875) );
  XNOR U9114 ( .A(n8874), .B(n8875), .Z(n8876) );
  XNOR U9115 ( .A(n8877), .B(n8876), .Z(n8947) );
  XNOR U9116 ( .A(n8947), .B(sreg[360]), .Z(n8949) );
  NAND U9117 ( .A(n8869), .B(sreg[359]), .Z(n8873) );
  OR U9118 ( .A(n8871), .B(n8870), .Z(n8872) );
  AND U9119 ( .A(n8873), .B(n8872), .Z(n8948) );
  XOR U9120 ( .A(n8949), .B(n8948), .Z(c[360]) );
  NANDN U9121 ( .A(n8875), .B(n8874), .Z(n8879) );
  NAND U9122 ( .A(n8877), .B(n8876), .Z(n8878) );
  NAND U9123 ( .A(n8879), .B(n8878), .Z(n8955) );
  NANDN U9124 ( .A(n8881), .B(n8880), .Z(n8885) );
  OR U9125 ( .A(n8883), .B(n8882), .Z(n8884) );
  NAND U9126 ( .A(n8885), .B(n8884), .Z(n9022) );
  NANDN U9127 ( .A(n8887), .B(n8886), .Z(n8891) );
  OR U9128 ( .A(n8889), .B(n8888), .Z(n8890) );
  NAND U9129 ( .A(n8891), .B(n8890), .Z(n9010) );
  XNOR U9130 ( .A(n20154), .B(n9045), .Z(n8995) );
  OR U9131 ( .A(n8995), .B(n20057), .Z(n8894) );
  NANDN U9132 ( .A(n8892), .B(n20098), .Z(n8893) );
  AND U9133 ( .A(n8894), .B(n8893), .Z(n8987) );
  NAND U9134 ( .A(b[0]), .B(a[121]), .Z(n8895) );
  XNOR U9135 ( .A(b[1]), .B(n8895), .Z(n8897) );
  NAND U9136 ( .A(a[120]), .B(n98), .Z(n8896) );
  AND U9137 ( .A(n8897), .B(n8896), .Z(n8986) );
  XOR U9138 ( .A(n8987), .B(n8986), .Z(n8989) );
  NAND U9139 ( .A(a[105]), .B(b[15]), .Z(n8988) );
  XOR U9140 ( .A(n8989), .B(n8988), .Z(n9007) );
  NAND U9141 ( .A(n19722), .B(n8898), .Z(n8900) );
  XNOR U9142 ( .A(b[5]), .B(n9669), .Z(n8998) );
  NANDN U9143 ( .A(n19640), .B(n8998), .Z(n8899) );
  NAND U9144 ( .A(n8900), .B(n8899), .Z(n8983) );
  XNOR U9145 ( .A(n19714), .B(n9513), .Z(n9001) );
  NANDN U9146 ( .A(n9001), .B(n19766), .Z(n8903) );
  NANDN U9147 ( .A(n8901), .B(n19767), .Z(n8902) );
  NAND U9148 ( .A(n8903), .B(n8902), .Z(n8980) );
  NAND U9149 ( .A(n19554), .B(n8904), .Z(n8906) );
  IV U9150 ( .A(a[119]), .Z(n9852) );
  XNOR U9151 ( .A(b[3]), .B(n9852), .Z(n9004) );
  NANDN U9152 ( .A(n19521), .B(n9004), .Z(n8905) );
  AND U9153 ( .A(n8906), .B(n8905), .Z(n8981) );
  XNOR U9154 ( .A(n8980), .B(n8981), .Z(n8982) );
  XOR U9155 ( .A(n8983), .B(n8982), .Z(n9008) );
  XOR U9156 ( .A(n9007), .B(n9008), .Z(n9009) );
  XNOR U9157 ( .A(n9010), .B(n9009), .Z(n8958) );
  NAND U9158 ( .A(n8908), .B(n8907), .Z(n8912) );
  NAND U9159 ( .A(n8910), .B(n8909), .Z(n8911) );
  NAND U9160 ( .A(n8912), .B(n8911), .Z(n8959) );
  XOR U9161 ( .A(n8958), .B(n8959), .Z(n8961) );
  XNOR U9162 ( .A(n20052), .B(n9201), .Z(n8964) );
  OR U9163 ( .A(n8964), .B(n20020), .Z(n8915) );
  NANDN U9164 ( .A(n8913), .B(n19960), .Z(n8914) );
  NAND U9165 ( .A(n8915), .B(n8914), .Z(n8977) );
  XNOR U9166 ( .A(n102), .B(n8916), .Z(n8968) );
  OR U9167 ( .A(n8968), .B(n20121), .Z(n8919) );
  NANDN U9168 ( .A(n8917), .B(n20122), .Z(n8918) );
  NAND U9169 ( .A(n8919), .B(n8918), .Z(n8974) );
  XNOR U9170 ( .A(n19975), .B(n9357), .Z(n8971) );
  NANDN U9171 ( .A(n8971), .B(n19883), .Z(n8922) );
  NANDN U9172 ( .A(n8920), .B(n19937), .Z(n8921) );
  AND U9173 ( .A(n8922), .B(n8921), .Z(n8975) );
  XNOR U9174 ( .A(n8974), .B(n8975), .Z(n8976) );
  XNOR U9175 ( .A(n8977), .B(n8976), .Z(n9013) );
  NANDN U9176 ( .A(n8924), .B(n8923), .Z(n8928) );
  NAND U9177 ( .A(n8926), .B(n8925), .Z(n8927) );
  NAND U9178 ( .A(n8928), .B(n8927), .Z(n9014) );
  XNOR U9179 ( .A(n9013), .B(n9014), .Z(n9015) );
  NANDN U9180 ( .A(n8930), .B(n8929), .Z(n8934) );
  NAND U9181 ( .A(n8932), .B(n8931), .Z(n8933) );
  AND U9182 ( .A(n8934), .B(n8933), .Z(n9016) );
  XNOR U9183 ( .A(n9015), .B(n9016), .Z(n8960) );
  XNOR U9184 ( .A(n8961), .B(n8960), .Z(n9019) );
  NANDN U9185 ( .A(n8936), .B(n8935), .Z(n8940) );
  NAND U9186 ( .A(n8938), .B(n8937), .Z(n8939) );
  NAND U9187 ( .A(n8940), .B(n8939), .Z(n9020) );
  XNOR U9188 ( .A(n9019), .B(n9020), .Z(n9021) );
  XOR U9189 ( .A(n9022), .B(n9021), .Z(n8952) );
  NANDN U9190 ( .A(n8942), .B(n8941), .Z(n8946) );
  NANDN U9191 ( .A(n8944), .B(n8943), .Z(n8945) );
  NAND U9192 ( .A(n8946), .B(n8945), .Z(n8953) );
  XNOR U9193 ( .A(n8952), .B(n8953), .Z(n8954) );
  XNOR U9194 ( .A(n8955), .B(n8954), .Z(n9025) );
  XNOR U9195 ( .A(n9025), .B(sreg[361]), .Z(n9027) );
  NAND U9196 ( .A(n8947), .B(sreg[360]), .Z(n8951) );
  OR U9197 ( .A(n8949), .B(n8948), .Z(n8950) );
  AND U9198 ( .A(n8951), .B(n8950), .Z(n9026) );
  XOR U9199 ( .A(n9027), .B(n9026), .Z(c[361]) );
  NANDN U9200 ( .A(n8953), .B(n8952), .Z(n8957) );
  NAND U9201 ( .A(n8955), .B(n8954), .Z(n8956) );
  NAND U9202 ( .A(n8957), .B(n8956), .Z(n9033) );
  NANDN U9203 ( .A(n8959), .B(n8958), .Z(n8963) );
  OR U9204 ( .A(n8961), .B(n8960), .Z(n8962) );
  NAND U9205 ( .A(n8963), .B(n8962), .Z(n9100) );
  XNOR U9206 ( .A(n20052), .B(n9279), .Z(n9042) );
  OR U9207 ( .A(n9042), .B(n20020), .Z(n8966) );
  NANDN U9208 ( .A(n8964), .B(n19960), .Z(n8965) );
  NAND U9209 ( .A(n8966), .B(n8965), .Z(n9055) );
  XNOR U9210 ( .A(n102), .B(n8967), .Z(n9046) );
  OR U9211 ( .A(n9046), .B(n20121), .Z(n8970) );
  NANDN U9212 ( .A(n8968), .B(n20122), .Z(n8969) );
  NAND U9213 ( .A(n8970), .B(n8969), .Z(n9052) );
  XNOR U9214 ( .A(n19975), .B(n9435), .Z(n9049) );
  NANDN U9215 ( .A(n9049), .B(n19883), .Z(n8973) );
  NANDN U9216 ( .A(n8971), .B(n19937), .Z(n8972) );
  AND U9217 ( .A(n8973), .B(n8972), .Z(n9053) );
  XNOR U9218 ( .A(n9052), .B(n9053), .Z(n9054) );
  XNOR U9219 ( .A(n9055), .B(n9054), .Z(n9091) );
  NANDN U9220 ( .A(n8975), .B(n8974), .Z(n8979) );
  NAND U9221 ( .A(n8977), .B(n8976), .Z(n8978) );
  NAND U9222 ( .A(n8979), .B(n8978), .Z(n9092) );
  XNOR U9223 ( .A(n9091), .B(n9092), .Z(n9093) );
  NANDN U9224 ( .A(n8981), .B(n8980), .Z(n8985) );
  NAND U9225 ( .A(n8983), .B(n8982), .Z(n8984) );
  AND U9226 ( .A(n8985), .B(n8984), .Z(n9094) );
  XNOR U9227 ( .A(n9093), .B(n9094), .Z(n9038) );
  NANDN U9228 ( .A(n8987), .B(n8986), .Z(n8991) );
  OR U9229 ( .A(n8989), .B(n8988), .Z(n8990) );
  NAND U9230 ( .A(n8991), .B(n8990), .Z(n9088) );
  NAND U9231 ( .A(b[0]), .B(a[122]), .Z(n8992) );
  XNOR U9232 ( .A(b[1]), .B(n8992), .Z(n8994) );
  NAND U9233 ( .A(a[121]), .B(n98), .Z(n8993) );
  AND U9234 ( .A(n8994), .B(n8993), .Z(n9064) );
  XNOR U9235 ( .A(n20154), .B(n9123), .Z(n9070) );
  OR U9236 ( .A(n9070), .B(n20057), .Z(n8997) );
  NANDN U9237 ( .A(n8995), .B(n20098), .Z(n8996) );
  AND U9238 ( .A(n8997), .B(n8996), .Z(n9065) );
  XOR U9239 ( .A(n9064), .B(n9065), .Z(n9067) );
  NAND U9240 ( .A(a[106]), .B(b[15]), .Z(n9066) );
  XOR U9241 ( .A(n9067), .B(n9066), .Z(n9085) );
  NAND U9242 ( .A(n19722), .B(n8998), .Z(n9000) );
  XNOR U9243 ( .A(b[5]), .B(n9747), .Z(n9076) );
  NANDN U9244 ( .A(n19640), .B(n9076), .Z(n8999) );
  NAND U9245 ( .A(n9000), .B(n8999), .Z(n9061) );
  XNOR U9246 ( .A(n19714), .B(n9591), .Z(n9079) );
  NANDN U9247 ( .A(n9079), .B(n19766), .Z(n9003) );
  NANDN U9248 ( .A(n9001), .B(n19767), .Z(n9002) );
  NAND U9249 ( .A(n9003), .B(n9002), .Z(n9058) );
  NAND U9250 ( .A(n19554), .B(n9004), .Z(n9006) );
  IV U9251 ( .A(a[120]), .Z(n9903) );
  XNOR U9252 ( .A(b[3]), .B(n9903), .Z(n9082) );
  NANDN U9253 ( .A(n19521), .B(n9082), .Z(n9005) );
  AND U9254 ( .A(n9006), .B(n9005), .Z(n9059) );
  XNOR U9255 ( .A(n9058), .B(n9059), .Z(n9060) );
  XOR U9256 ( .A(n9061), .B(n9060), .Z(n9086) );
  XOR U9257 ( .A(n9085), .B(n9086), .Z(n9087) );
  XNOR U9258 ( .A(n9088), .B(n9087), .Z(n9036) );
  NAND U9259 ( .A(n9008), .B(n9007), .Z(n9012) );
  NAND U9260 ( .A(n9010), .B(n9009), .Z(n9011) );
  NAND U9261 ( .A(n9012), .B(n9011), .Z(n9037) );
  XOR U9262 ( .A(n9036), .B(n9037), .Z(n9039) );
  XNOR U9263 ( .A(n9038), .B(n9039), .Z(n9097) );
  NANDN U9264 ( .A(n9014), .B(n9013), .Z(n9018) );
  NAND U9265 ( .A(n9016), .B(n9015), .Z(n9017) );
  NAND U9266 ( .A(n9018), .B(n9017), .Z(n9098) );
  XNOR U9267 ( .A(n9097), .B(n9098), .Z(n9099) );
  XOR U9268 ( .A(n9100), .B(n9099), .Z(n9030) );
  NANDN U9269 ( .A(n9020), .B(n9019), .Z(n9024) );
  NANDN U9270 ( .A(n9022), .B(n9021), .Z(n9023) );
  NAND U9271 ( .A(n9024), .B(n9023), .Z(n9031) );
  XNOR U9272 ( .A(n9030), .B(n9031), .Z(n9032) );
  XNOR U9273 ( .A(n9033), .B(n9032), .Z(n9103) );
  XNOR U9274 ( .A(n9103), .B(sreg[362]), .Z(n9105) );
  NAND U9275 ( .A(n9025), .B(sreg[361]), .Z(n9029) );
  OR U9276 ( .A(n9027), .B(n9026), .Z(n9028) );
  AND U9277 ( .A(n9029), .B(n9028), .Z(n9104) );
  XOR U9278 ( .A(n9105), .B(n9104), .Z(c[362]) );
  NANDN U9279 ( .A(n9031), .B(n9030), .Z(n9035) );
  NAND U9280 ( .A(n9033), .B(n9032), .Z(n9034) );
  NAND U9281 ( .A(n9035), .B(n9034), .Z(n9111) );
  NANDN U9282 ( .A(n9037), .B(n9036), .Z(n9041) );
  OR U9283 ( .A(n9039), .B(n9038), .Z(n9040) );
  NAND U9284 ( .A(n9041), .B(n9040), .Z(n9178) );
  XNOR U9285 ( .A(n20052), .B(n9357), .Z(n9120) );
  OR U9286 ( .A(n9120), .B(n20020), .Z(n9044) );
  NANDN U9287 ( .A(n9042), .B(n19960), .Z(n9043) );
  NAND U9288 ( .A(n9044), .B(n9043), .Z(n9133) );
  XNOR U9289 ( .A(n102), .B(n9045), .Z(n9124) );
  OR U9290 ( .A(n9124), .B(n20121), .Z(n9048) );
  NANDN U9291 ( .A(n9046), .B(n20122), .Z(n9047) );
  NAND U9292 ( .A(n9048), .B(n9047), .Z(n9130) );
  XNOR U9293 ( .A(n19975), .B(n9513), .Z(n9127) );
  NANDN U9294 ( .A(n9127), .B(n19883), .Z(n9051) );
  NANDN U9295 ( .A(n9049), .B(n19937), .Z(n9050) );
  AND U9296 ( .A(n9051), .B(n9050), .Z(n9131) );
  XNOR U9297 ( .A(n9130), .B(n9131), .Z(n9132) );
  XNOR U9298 ( .A(n9133), .B(n9132), .Z(n9169) );
  NANDN U9299 ( .A(n9053), .B(n9052), .Z(n9057) );
  NAND U9300 ( .A(n9055), .B(n9054), .Z(n9056) );
  NAND U9301 ( .A(n9057), .B(n9056), .Z(n9170) );
  XNOR U9302 ( .A(n9169), .B(n9170), .Z(n9171) );
  NANDN U9303 ( .A(n9059), .B(n9058), .Z(n9063) );
  NAND U9304 ( .A(n9061), .B(n9060), .Z(n9062) );
  AND U9305 ( .A(n9063), .B(n9062), .Z(n9172) );
  XNOR U9306 ( .A(n9171), .B(n9172), .Z(n9116) );
  NANDN U9307 ( .A(n9065), .B(n9064), .Z(n9069) );
  OR U9308 ( .A(n9067), .B(n9066), .Z(n9068) );
  NAND U9309 ( .A(n9069), .B(n9068), .Z(n9166) );
  XNOR U9310 ( .A(n20154), .B(n9201), .Z(n9151) );
  OR U9311 ( .A(n9151), .B(n20057), .Z(n9072) );
  NANDN U9312 ( .A(n9070), .B(n20098), .Z(n9071) );
  AND U9313 ( .A(n9072), .B(n9071), .Z(n9143) );
  NAND U9314 ( .A(b[0]), .B(a[123]), .Z(n9073) );
  XNOR U9315 ( .A(b[1]), .B(n9073), .Z(n9075) );
  NAND U9316 ( .A(a[122]), .B(n98), .Z(n9074) );
  AND U9317 ( .A(n9075), .B(n9074), .Z(n9142) );
  XOR U9318 ( .A(n9143), .B(n9142), .Z(n9145) );
  NAND U9319 ( .A(a[107]), .B(b[15]), .Z(n9144) );
  XOR U9320 ( .A(n9145), .B(n9144), .Z(n9163) );
  NAND U9321 ( .A(n19722), .B(n9076), .Z(n9078) );
  XNOR U9322 ( .A(b[5]), .B(n9852), .Z(n9154) );
  NANDN U9323 ( .A(n19640), .B(n9154), .Z(n9077) );
  NAND U9324 ( .A(n9078), .B(n9077), .Z(n9139) );
  XNOR U9325 ( .A(n19714), .B(n9669), .Z(n9157) );
  NANDN U9326 ( .A(n9157), .B(n19766), .Z(n9081) );
  NANDN U9327 ( .A(n9079), .B(n19767), .Z(n9080) );
  NAND U9328 ( .A(n9081), .B(n9080), .Z(n9136) );
  NAND U9329 ( .A(n19554), .B(n9082), .Z(n9084) );
  IV U9330 ( .A(a[121]), .Z(n10006) );
  XNOR U9331 ( .A(b[3]), .B(n10006), .Z(n9160) );
  NANDN U9332 ( .A(n19521), .B(n9160), .Z(n9083) );
  AND U9333 ( .A(n9084), .B(n9083), .Z(n9137) );
  XNOR U9334 ( .A(n9136), .B(n9137), .Z(n9138) );
  XOR U9335 ( .A(n9139), .B(n9138), .Z(n9164) );
  XOR U9336 ( .A(n9163), .B(n9164), .Z(n9165) );
  XNOR U9337 ( .A(n9166), .B(n9165), .Z(n9114) );
  NAND U9338 ( .A(n9086), .B(n9085), .Z(n9090) );
  NAND U9339 ( .A(n9088), .B(n9087), .Z(n9089) );
  NAND U9340 ( .A(n9090), .B(n9089), .Z(n9115) );
  XOR U9341 ( .A(n9114), .B(n9115), .Z(n9117) );
  XNOR U9342 ( .A(n9116), .B(n9117), .Z(n9175) );
  NANDN U9343 ( .A(n9092), .B(n9091), .Z(n9096) );
  NAND U9344 ( .A(n9094), .B(n9093), .Z(n9095) );
  NAND U9345 ( .A(n9096), .B(n9095), .Z(n9176) );
  XNOR U9346 ( .A(n9175), .B(n9176), .Z(n9177) );
  XOR U9347 ( .A(n9178), .B(n9177), .Z(n9108) );
  NANDN U9348 ( .A(n9098), .B(n9097), .Z(n9102) );
  NANDN U9349 ( .A(n9100), .B(n9099), .Z(n9101) );
  NAND U9350 ( .A(n9102), .B(n9101), .Z(n9109) );
  XNOR U9351 ( .A(n9108), .B(n9109), .Z(n9110) );
  XNOR U9352 ( .A(n9111), .B(n9110), .Z(n9181) );
  XNOR U9353 ( .A(n9181), .B(sreg[363]), .Z(n9183) );
  NAND U9354 ( .A(n9103), .B(sreg[362]), .Z(n9107) );
  OR U9355 ( .A(n9105), .B(n9104), .Z(n9106) );
  AND U9356 ( .A(n9107), .B(n9106), .Z(n9182) );
  XOR U9357 ( .A(n9183), .B(n9182), .Z(c[363]) );
  NANDN U9358 ( .A(n9109), .B(n9108), .Z(n9113) );
  NAND U9359 ( .A(n9111), .B(n9110), .Z(n9112) );
  NAND U9360 ( .A(n9113), .B(n9112), .Z(n9189) );
  NANDN U9361 ( .A(n9115), .B(n9114), .Z(n9119) );
  OR U9362 ( .A(n9117), .B(n9116), .Z(n9118) );
  NAND U9363 ( .A(n9119), .B(n9118), .Z(n9256) );
  XNOR U9364 ( .A(n20052), .B(n9435), .Z(n9198) );
  OR U9365 ( .A(n9198), .B(n20020), .Z(n9122) );
  NANDN U9366 ( .A(n9120), .B(n19960), .Z(n9121) );
  NAND U9367 ( .A(n9122), .B(n9121), .Z(n9211) );
  XNOR U9368 ( .A(n102), .B(n9123), .Z(n9202) );
  OR U9369 ( .A(n9202), .B(n20121), .Z(n9126) );
  NANDN U9370 ( .A(n9124), .B(n20122), .Z(n9125) );
  NAND U9371 ( .A(n9126), .B(n9125), .Z(n9208) );
  XNOR U9372 ( .A(n19975), .B(n9591), .Z(n9205) );
  NANDN U9373 ( .A(n9205), .B(n19883), .Z(n9129) );
  NANDN U9374 ( .A(n9127), .B(n19937), .Z(n9128) );
  AND U9375 ( .A(n9129), .B(n9128), .Z(n9209) );
  XNOR U9376 ( .A(n9208), .B(n9209), .Z(n9210) );
  XNOR U9377 ( .A(n9211), .B(n9210), .Z(n9247) );
  NANDN U9378 ( .A(n9131), .B(n9130), .Z(n9135) );
  NAND U9379 ( .A(n9133), .B(n9132), .Z(n9134) );
  NAND U9380 ( .A(n9135), .B(n9134), .Z(n9248) );
  XNOR U9381 ( .A(n9247), .B(n9248), .Z(n9249) );
  NANDN U9382 ( .A(n9137), .B(n9136), .Z(n9141) );
  NAND U9383 ( .A(n9139), .B(n9138), .Z(n9140) );
  AND U9384 ( .A(n9141), .B(n9140), .Z(n9250) );
  XNOR U9385 ( .A(n9249), .B(n9250), .Z(n9194) );
  NANDN U9386 ( .A(n9143), .B(n9142), .Z(n9147) );
  OR U9387 ( .A(n9145), .B(n9144), .Z(n9146) );
  NAND U9388 ( .A(n9147), .B(n9146), .Z(n9244) );
  NAND U9389 ( .A(b[0]), .B(a[124]), .Z(n9148) );
  XNOR U9390 ( .A(b[1]), .B(n9148), .Z(n9150) );
  NAND U9391 ( .A(a[123]), .B(n98), .Z(n9149) );
  AND U9392 ( .A(n9150), .B(n9149), .Z(n9220) );
  XNOR U9393 ( .A(n20154), .B(n9279), .Z(n9229) );
  OR U9394 ( .A(n9229), .B(n20057), .Z(n9153) );
  NANDN U9395 ( .A(n9151), .B(n20098), .Z(n9152) );
  AND U9396 ( .A(n9153), .B(n9152), .Z(n9221) );
  XOR U9397 ( .A(n9220), .B(n9221), .Z(n9223) );
  NAND U9398 ( .A(a[108]), .B(b[15]), .Z(n9222) );
  XOR U9399 ( .A(n9223), .B(n9222), .Z(n9241) );
  NAND U9400 ( .A(n19722), .B(n9154), .Z(n9156) );
  XNOR U9401 ( .A(b[5]), .B(n9903), .Z(n9232) );
  NANDN U9402 ( .A(n19640), .B(n9232), .Z(n9155) );
  NAND U9403 ( .A(n9156), .B(n9155), .Z(n9217) );
  XNOR U9404 ( .A(n19714), .B(n9747), .Z(n9235) );
  NANDN U9405 ( .A(n9235), .B(n19766), .Z(n9159) );
  NANDN U9406 ( .A(n9157), .B(n19767), .Z(n9158) );
  NAND U9407 ( .A(n9159), .B(n9158), .Z(n9214) );
  NAND U9408 ( .A(n19554), .B(n9160), .Z(n9162) );
  IV U9409 ( .A(a[122]), .Z(n10084) );
  XNOR U9410 ( .A(b[3]), .B(n10084), .Z(n9238) );
  NANDN U9411 ( .A(n19521), .B(n9238), .Z(n9161) );
  AND U9412 ( .A(n9162), .B(n9161), .Z(n9215) );
  XNOR U9413 ( .A(n9214), .B(n9215), .Z(n9216) );
  XOR U9414 ( .A(n9217), .B(n9216), .Z(n9242) );
  XOR U9415 ( .A(n9241), .B(n9242), .Z(n9243) );
  XNOR U9416 ( .A(n9244), .B(n9243), .Z(n9192) );
  NAND U9417 ( .A(n9164), .B(n9163), .Z(n9168) );
  NAND U9418 ( .A(n9166), .B(n9165), .Z(n9167) );
  NAND U9419 ( .A(n9168), .B(n9167), .Z(n9193) );
  XOR U9420 ( .A(n9192), .B(n9193), .Z(n9195) );
  XNOR U9421 ( .A(n9194), .B(n9195), .Z(n9253) );
  NANDN U9422 ( .A(n9170), .B(n9169), .Z(n9174) );
  NAND U9423 ( .A(n9172), .B(n9171), .Z(n9173) );
  NAND U9424 ( .A(n9174), .B(n9173), .Z(n9254) );
  XNOR U9425 ( .A(n9253), .B(n9254), .Z(n9255) );
  XOR U9426 ( .A(n9256), .B(n9255), .Z(n9186) );
  NANDN U9427 ( .A(n9176), .B(n9175), .Z(n9180) );
  NANDN U9428 ( .A(n9178), .B(n9177), .Z(n9179) );
  NAND U9429 ( .A(n9180), .B(n9179), .Z(n9187) );
  XNOR U9430 ( .A(n9186), .B(n9187), .Z(n9188) );
  XNOR U9431 ( .A(n9189), .B(n9188), .Z(n9259) );
  XNOR U9432 ( .A(n9259), .B(sreg[364]), .Z(n9261) );
  NAND U9433 ( .A(n9181), .B(sreg[363]), .Z(n9185) );
  OR U9434 ( .A(n9183), .B(n9182), .Z(n9184) );
  AND U9435 ( .A(n9185), .B(n9184), .Z(n9260) );
  XOR U9436 ( .A(n9261), .B(n9260), .Z(c[364]) );
  NANDN U9437 ( .A(n9187), .B(n9186), .Z(n9191) );
  NAND U9438 ( .A(n9189), .B(n9188), .Z(n9190) );
  NAND U9439 ( .A(n9191), .B(n9190), .Z(n9267) );
  NANDN U9440 ( .A(n9193), .B(n9192), .Z(n9197) );
  OR U9441 ( .A(n9195), .B(n9194), .Z(n9196) );
  NAND U9442 ( .A(n9197), .B(n9196), .Z(n9334) );
  XNOR U9443 ( .A(n20052), .B(n9513), .Z(n9276) );
  OR U9444 ( .A(n9276), .B(n20020), .Z(n9200) );
  NANDN U9445 ( .A(n9198), .B(n19960), .Z(n9199) );
  NAND U9446 ( .A(n9200), .B(n9199), .Z(n9289) );
  XNOR U9447 ( .A(n102), .B(n9201), .Z(n9280) );
  OR U9448 ( .A(n9280), .B(n20121), .Z(n9204) );
  NANDN U9449 ( .A(n9202), .B(n20122), .Z(n9203) );
  NAND U9450 ( .A(n9204), .B(n9203), .Z(n9286) );
  XNOR U9451 ( .A(n19975), .B(n9669), .Z(n9283) );
  NANDN U9452 ( .A(n9283), .B(n19883), .Z(n9207) );
  NANDN U9453 ( .A(n9205), .B(n19937), .Z(n9206) );
  AND U9454 ( .A(n9207), .B(n9206), .Z(n9287) );
  XNOR U9455 ( .A(n9286), .B(n9287), .Z(n9288) );
  XNOR U9456 ( .A(n9289), .B(n9288), .Z(n9325) );
  NANDN U9457 ( .A(n9209), .B(n9208), .Z(n9213) );
  NAND U9458 ( .A(n9211), .B(n9210), .Z(n9212) );
  NAND U9459 ( .A(n9213), .B(n9212), .Z(n9326) );
  XNOR U9460 ( .A(n9325), .B(n9326), .Z(n9327) );
  NANDN U9461 ( .A(n9215), .B(n9214), .Z(n9219) );
  NAND U9462 ( .A(n9217), .B(n9216), .Z(n9218) );
  AND U9463 ( .A(n9219), .B(n9218), .Z(n9328) );
  XNOR U9464 ( .A(n9327), .B(n9328), .Z(n9272) );
  NANDN U9465 ( .A(n9221), .B(n9220), .Z(n9225) );
  OR U9466 ( .A(n9223), .B(n9222), .Z(n9224) );
  NAND U9467 ( .A(n9225), .B(n9224), .Z(n9322) );
  NAND U9468 ( .A(b[0]), .B(a[125]), .Z(n9226) );
  XNOR U9469 ( .A(b[1]), .B(n9226), .Z(n9228) );
  NAND U9470 ( .A(a[124]), .B(n98), .Z(n9227) );
  AND U9471 ( .A(n9228), .B(n9227), .Z(n9298) );
  XNOR U9472 ( .A(n20154), .B(n9357), .Z(n9307) );
  OR U9473 ( .A(n9307), .B(n20057), .Z(n9231) );
  NANDN U9474 ( .A(n9229), .B(n20098), .Z(n9230) );
  AND U9475 ( .A(n9231), .B(n9230), .Z(n9299) );
  XOR U9476 ( .A(n9298), .B(n9299), .Z(n9301) );
  NAND U9477 ( .A(a[109]), .B(b[15]), .Z(n9300) );
  XOR U9478 ( .A(n9301), .B(n9300), .Z(n9319) );
  NAND U9479 ( .A(n19722), .B(n9232), .Z(n9234) );
  XNOR U9480 ( .A(b[5]), .B(n10006), .Z(n9310) );
  NANDN U9481 ( .A(n19640), .B(n9310), .Z(n9233) );
  NAND U9482 ( .A(n9234), .B(n9233), .Z(n9295) );
  XNOR U9483 ( .A(n19714), .B(n9852), .Z(n9313) );
  NANDN U9484 ( .A(n9313), .B(n19766), .Z(n9237) );
  NANDN U9485 ( .A(n9235), .B(n19767), .Z(n9236) );
  NAND U9486 ( .A(n9237), .B(n9236), .Z(n9292) );
  NAND U9487 ( .A(n19554), .B(n9238), .Z(n9240) );
  IV U9488 ( .A(a[123]), .Z(n10135) );
  XNOR U9489 ( .A(b[3]), .B(n10135), .Z(n9316) );
  NANDN U9490 ( .A(n19521), .B(n9316), .Z(n9239) );
  AND U9491 ( .A(n9240), .B(n9239), .Z(n9293) );
  XNOR U9492 ( .A(n9292), .B(n9293), .Z(n9294) );
  XOR U9493 ( .A(n9295), .B(n9294), .Z(n9320) );
  XOR U9494 ( .A(n9319), .B(n9320), .Z(n9321) );
  XNOR U9495 ( .A(n9322), .B(n9321), .Z(n9270) );
  NAND U9496 ( .A(n9242), .B(n9241), .Z(n9246) );
  NAND U9497 ( .A(n9244), .B(n9243), .Z(n9245) );
  NAND U9498 ( .A(n9246), .B(n9245), .Z(n9271) );
  XOR U9499 ( .A(n9270), .B(n9271), .Z(n9273) );
  XNOR U9500 ( .A(n9272), .B(n9273), .Z(n9331) );
  NANDN U9501 ( .A(n9248), .B(n9247), .Z(n9252) );
  NAND U9502 ( .A(n9250), .B(n9249), .Z(n9251) );
  NAND U9503 ( .A(n9252), .B(n9251), .Z(n9332) );
  XNOR U9504 ( .A(n9331), .B(n9332), .Z(n9333) );
  XOR U9505 ( .A(n9334), .B(n9333), .Z(n9264) );
  NANDN U9506 ( .A(n9254), .B(n9253), .Z(n9258) );
  NANDN U9507 ( .A(n9256), .B(n9255), .Z(n9257) );
  NAND U9508 ( .A(n9258), .B(n9257), .Z(n9265) );
  XNOR U9509 ( .A(n9264), .B(n9265), .Z(n9266) );
  XNOR U9510 ( .A(n9267), .B(n9266), .Z(n9337) );
  XNOR U9511 ( .A(n9337), .B(sreg[365]), .Z(n9339) );
  NAND U9512 ( .A(n9259), .B(sreg[364]), .Z(n9263) );
  OR U9513 ( .A(n9261), .B(n9260), .Z(n9262) );
  AND U9514 ( .A(n9263), .B(n9262), .Z(n9338) );
  XOR U9515 ( .A(n9339), .B(n9338), .Z(c[365]) );
  NANDN U9516 ( .A(n9265), .B(n9264), .Z(n9269) );
  NAND U9517 ( .A(n9267), .B(n9266), .Z(n9268) );
  NAND U9518 ( .A(n9269), .B(n9268), .Z(n9345) );
  NANDN U9519 ( .A(n9271), .B(n9270), .Z(n9275) );
  OR U9520 ( .A(n9273), .B(n9272), .Z(n9274) );
  NAND U9521 ( .A(n9275), .B(n9274), .Z(n9412) );
  XNOR U9522 ( .A(n20052), .B(n9591), .Z(n9354) );
  OR U9523 ( .A(n9354), .B(n20020), .Z(n9278) );
  NANDN U9524 ( .A(n9276), .B(n19960), .Z(n9277) );
  NAND U9525 ( .A(n9278), .B(n9277), .Z(n9367) );
  XNOR U9526 ( .A(n102), .B(n9279), .Z(n9358) );
  OR U9527 ( .A(n9358), .B(n20121), .Z(n9282) );
  NANDN U9528 ( .A(n9280), .B(n20122), .Z(n9281) );
  NAND U9529 ( .A(n9282), .B(n9281), .Z(n9364) );
  XNOR U9530 ( .A(n19975), .B(n9747), .Z(n9361) );
  NANDN U9531 ( .A(n9361), .B(n19883), .Z(n9285) );
  NANDN U9532 ( .A(n9283), .B(n19937), .Z(n9284) );
  AND U9533 ( .A(n9285), .B(n9284), .Z(n9365) );
  XNOR U9534 ( .A(n9364), .B(n9365), .Z(n9366) );
  XNOR U9535 ( .A(n9367), .B(n9366), .Z(n9403) );
  NANDN U9536 ( .A(n9287), .B(n9286), .Z(n9291) );
  NAND U9537 ( .A(n9289), .B(n9288), .Z(n9290) );
  NAND U9538 ( .A(n9291), .B(n9290), .Z(n9404) );
  XNOR U9539 ( .A(n9403), .B(n9404), .Z(n9405) );
  NANDN U9540 ( .A(n9293), .B(n9292), .Z(n9297) );
  NAND U9541 ( .A(n9295), .B(n9294), .Z(n9296) );
  AND U9542 ( .A(n9297), .B(n9296), .Z(n9406) );
  XNOR U9543 ( .A(n9405), .B(n9406), .Z(n9350) );
  NANDN U9544 ( .A(n9299), .B(n9298), .Z(n9303) );
  OR U9545 ( .A(n9301), .B(n9300), .Z(n9302) );
  NAND U9546 ( .A(n9303), .B(n9302), .Z(n9400) );
  NAND U9547 ( .A(b[0]), .B(a[126]), .Z(n9304) );
  XNOR U9548 ( .A(b[1]), .B(n9304), .Z(n9306) );
  NAND U9549 ( .A(a[125]), .B(n98), .Z(n9305) );
  AND U9550 ( .A(n9306), .B(n9305), .Z(n9376) );
  XNOR U9551 ( .A(n20154), .B(n9435), .Z(n9382) );
  OR U9552 ( .A(n9382), .B(n20057), .Z(n9309) );
  NANDN U9553 ( .A(n9307), .B(n20098), .Z(n9308) );
  AND U9554 ( .A(n9309), .B(n9308), .Z(n9377) );
  XOR U9555 ( .A(n9376), .B(n9377), .Z(n9379) );
  NAND U9556 ( .A(a[110]), .B(b[15]), .Z(n9378) );
  XOR U9557 ( .A(n9379), .B(n9378), .Z(n9397) );
  NAND U9558 ( .A(n19722), .B(n9310), .Z(n9312) );
  XNOR U9559 ( .A(b[5]), .B(n10084), .Z(n9388) );
  NANDN U9560 ( .A(n19640), .B(n9388), .Z(n9311) );
  NAND U9561 ( .A(n9312), .B(n9311), .Z(n9373) );
  XNOR U9562 ( .A(n19714), .B(n9903), .Z(n9391) );
  NANDN U9563 ( .A(n9391), .B(n19766), .Z(n9315) );
  NANDN U9564 ( .A(n9313), .B(n19767), .Z(n9314) );
  NAND U9565 ( .A(n9315), .B(n9314), .Z(n9370) );
  NAND U9566 ( .A(n19554), .B(n9316), .Z(n9318) );
  IV U9567 ( .A(a[124]), .Z(n10213) );
  XNOR U9568 ( .A(b[3]), .B(n10213), .Z(n9394) );
  NANDN U9569 ( .A(n19521), .B(n9394), .Z(n9317) );
  AND U9570 ( .A(n9318), .B(n9317), .Z(n9371) );
  XNOR U9571 ( .A(n9370), .B(n9371), .Z(n9372) );
  XOR U9572 ( .A(n9373), .B(n9372), .Z(n9398) );
  XOR U9573 ( .A(n9397), .B(n9398), .Z(n9399) );
  XNOR U9574 ( .A(n9400), .B(n9399), .Z(n9348) );
  NAND U9575 ( .A(n9320), .B(n9319), .Z(n9324) );
  NAND U9576 ( .A(n9322), .B(n9321), .Z(n9323) );
  NAND U9577 ( .A(n9324), .B(n9323), .Z(n9349) );
  XOR U9578 ( .A(n9348), .B(n9349), .Z(n9351) );
  XNOR U9579 ( .A(n9350), .B(n9351), .Z(n9409) );
  NANDN U9580 ( .A(n9326), .B(n9325), .Z(n9330) );
  NAND U9581 ( .A(n9328), .B(n9327), .Z(n9329) );
  NAND U9582 ( .A(n9330), .B(n9329), .Z(n9410) );
  XNOR U9583 ( .A(n9409), .B(n9410), .Z(n9411) );
  XOR U9584 ( .A(n9412), .B(n9411), .Z(n9342) );
  NANDN U9585 ( .A(n9332), .B(n9331), .Z(n9336) );
  NANDN U9586 ( .A(n9334), .B(n9333), .Z(n9335) );
  NAND U9587 ( .A(n9336), .B(n9335), .Z(n9343) );
  XNOR U9588 ( .A(n9342), .B(n9343), .Z(n9344) );
  XNOR U9589 ( .A(n9345), .B(n9344), .Z(n9415) );
  XNOR U9590 ( .A(n9415), .B(sreg[366]), .Z(n9417) );
  NAND U9591 ( .A(n9337), .B(sreg[365]), .Z(n9341) );
  OR U9592 ( .A(n9339), .B(n9338), .Z(n9340) );
  AND U9593 ( .A(n9341), .B(n9340), .Z(n9416) );
  XOR U9594 ( .A(n9417), .B(n9416), .Z(c[366]) );
  NANDN U9595 ( .A(n9343), .B(n9342), .Z(n9347) );
  NAND U9596 ( .A(n9345), .B(n9344), .Z(n9346) );
  NAND U9597 ( .A(n9347), .B(n9346), .Z(n9423) );
  NANDN U9598 ( .A(n9349), .B(n9348), .Z(n9353) );
  OR U9599 ( .A(n9351), .B(n9350), .Z(n9352) );
  NAND U9600 ( .A(n9353), .B(n9352), .Z(n9490) );
  XNOR U9601 ( .A(n20052), .B(n9669), .Z(n9432) );
  OR U9602 ( .A(n9432), .B(n20020), .Z(n9356) );
  NANDN U9603 ( .A(n9354), .B(n19960), .Z(n9355) );
  NAND U9604 ( .A(n9356), .B(n9355), .Z(n9445) );
  XNOR U9605 ( .A(n102), .B(n9357), .Z(n9436) );
  OR U9606 ( .A(n9436), .B(n20121), .Z(n9360) );
  NANDN U9607 ( .A(n9358), .B(n20122), .Z(n9359) );
  NAND U9608 ( .A(n9360), .B(n9359), .Z(n9442) );
  XNOR U9609 ( .A(n19975), .B(n9852), .Z(n9439) );
  NANDN U9610 ( .A(n9439), .B(n19883), .Z(n9363) );
  NANDN U9611 ( .A(n9361), .B(n19937), .Z(n9362) );
  AND U9612 ( .A(n9363), .B(n9362), .Z(n9443) );
  XNOR U9613 ( .A(n9442), .B(n9443), .Z(n9444) );
  XNOR U9614 ( .A(n9445), .B(n9444), .Z(n9481) );
  NANDN U9615 ( .A(n9365), .B(n9364), .Z(n9369) );
  NAND U9616 ( .A(n9367), .B(n9366), .Z(n9368) );
  NAND U9617 ( .A(n9369), .B(n9368), .Z(n9482) );
  XNOR U9618 ( .A(n9481), .B(n9482), .Z(n9483) );
  NANDN U9619 ( .A(n9371), .B(n9370), .Z(n9375) );
  NAND U9620 ( .A(n9373), .B(n9372), .Z(n9374) );
  AND U9621 ( .A(n9375), .B(n9374), .Z(n9484) );
  XNOR U9622 ( .A(n9483), .B(n9484), .Z(n9428) );
  NANDN U9623 ( .A(n9377), .B(n9376), .Z(n9381) );
  OR U9624 ( .A(n9379), .B(n9378), .Z(n9380) );
  NAND U9625 ( .A(n9381), .B(n9380), .Z(n9478) );
  XNOR U9626 ( .A(n20154), .B(n9513), .Z(n9463) );
  OR U9627 ( .A(n9463), .B(n20057), .Z(n9384) );
  NANDN U9628 ( .A(n9382), .B(n20098), .Z(n9383) );
  AND U9629 ( .A(n9384), .B(n9383), .Z(n9455) );
  NAND U9630 ( .A(b[0]), .B(a[127]), .Z(n9385) );
  XNOR U9631 ( .A(b[1]), .B(n9385), .Z(n9387) );
  NAND U9632 ( .A(a[126]), .B(n98), .Z(n9386) );
  AND U9633 ( .A(n9387), .B(n9386), .Z(n9454) );
  XOR U9634 ( .A(n9455), .B(n9454), .Z(n9457) );
  NAND U9635 ( .A(a[111]), .B(b[15]), .Z(n9456) );
  XOR U9636 ( .A(n9457), .B(n9456), .Z(n9475) );
  NAND U9637 ( .A(n19722), .B(n9388), .Z(n9390) );
  XNOR U9638 ( .A(b[5]), .B(n10135), .Z(n9466) );
  NANDN U9639 ( .A(n19640), .B(n9466), .Z(n9389) );
  NAND U9640 ( .A(n9390), .B(n9389), .Z(n9451) );
  XNOR U9641 ( .A(n19714), .B(n10006), .Z(n9469) );
  NANDN U9642 ( .A(n9469), .B(n19766), .Z(n9393) );
  NANDN U9643 ( .A(n9391), .B(n19767), .Z(n9392) );
  NAND U9644 ( .A(n9393), .B(n9392), .Z(n9448) );
  NAND U9645 ( .A(n19554), .B(n9394), .Z(n9396) );
  IV U9646 ( .A(a[125]), .Z(n10291) );
  XNOR U9647 ( .A(b[3]), .B(n10291), .Z(n9472) );
  NANDN U9648 ( .A(n19521), .B(n9472), .Z(n9395) );
  AND U9649 ( .A(n9396), .B(n9395), .Z(n9449) );
  XNOR U9650 ( .A(n9448), .B(n9449), .Z(n9450) );
  XOR U9651 ( .A(n9451), .B(n9450), .Z(n9476) );
  XOR U9652 ( .A(n9475), .B(n9476), .Z(n9477) );
  XNOR U9653 ( .A(n9478), .B(n9477), .Z(n9426) );
  NAND U9654 ( .A(n9398), .B(n9397), .Z(n9402) );
  NAND U9655 ( .A(n9400), .B(n9399), .Z(n9401) );
  NAND U9656 ( .A(n9402), .B(n9401), .Z(n9427) );
  XOR U9657 ( .A(n9426), .B(n9427), .Z(n9429) );
  XNOR U9658 ( .A(n9428), .B(n9429), .Z(n9487) );
  NANDN U9659 ( .A(n9404), .B(n9403), .Z(n9408) );
  NAND U9660 ( .A(n9406), .B(n9405), .Z(n9407) );
  NAND U9661 ( .A(n9408), .B(n9407), .Z(n9488) );
  XNOR U9662 ( .A(n9487), .B(n9488), .Z(n9489) );
  XOR U9663 ( .A(n9490), .B(n9489), .Z(n9420) );
  NANDN U9664 ( .A(n9410), .B(n9409), .Z(n9414) );
  NANDN U9665 ( .A(n9412), .B(n9411), .Z(n9413) );
  NAND U9666 ( .A(n9414), .B(n9413), .Z(n9421) );
  XNOR U9667 ( .A(n9420), .B(n9421), .Z(n9422) );
  XNOR U9668 ( .A(n9423), .B(n9422), .Z(n9493) );
  XNOR U9669 ( .A(n9493), .B(sreg[367]), .Z(n9495) );
  NAND U9670 ( .A(n9415), .B(sreg[366]), .Z(n9419) );
  OR U9671 ( .A(n9417), .B(n9416), .Z(n9418) );
  AND U9672 ( .A(n9419), .B(n9418), .Z(n9494) );
  XOR U9673 ( .A(n9495), .B(n9494), .Z(c[367]) );
  NANDN U9674 ( .A(n9421), .B(n9420), .Z(n9425) );
  NAND U9675 ( .A(n9423), .B(n9422), .Z(n9424) );
  NAND U9676 ( .A(n9425), .B(n9424), .Z(n9501) );
  NANDN U9677 ( .A(n9427), .B(n9426), .Z(n9431) );
  OR U9678 ( .A(n9429), .B(n9428), .Z(n9430) );
  NAND U9679 ( .A(n9431), .B(n9430), .Z(n9568) );
  XNOR U9680 ( .A(n20052), .B(n9747), .Z(n9510) );
  OR U9681 ( .A(n9510), .B(n20020), .Z(n9434) );
  NANDN U9682 ( .A(n9432), .B(n19960), .Z(n9433) );
  NAND U9683 ( .A(n9434), .B(n9433), .Z(n9523) );
  XNOR U9684 ( .A(n102), .B(n9435), .Z(n9514) );
  OR U9685 ( .A(n9514), .B(n20121), .Z(n9438) );
  NANDN U9686 ( .A(n9436), .B(n20122), .Z(n9437) );
  NAND U9687 ( .A(n9438), .B(n9437), .Z(n9520) );
  XNOR U9688 ( .A(n19975), .B(n9903), .Z(n9517) );
  NANDN U9689 ( .A(n9517), .B(n19883), .Z(n9441) );
  NANDN U9690 ( .A(n9439), .B(n19937), .Z(n9440) );
  AND U9691 ( .A(n9441), .B(n9440), .Z(n9521) );
  XNOR U9692 ( .A(n9520), .B(n9521), .Z(n9522) );
  XNOR U9693 ( .A(n9523), .B(n9522), .Z(n9559) );
  NANDN U9694 ( .A(n9443), .B(n9442), .Z(n9447) );
  NAND U9695 ( .A(n9445), .B(n9444), .Z(n9446) );
  NAND U9696 ( .A(n9447), .B(n9446), .Z(n9560) );
  XNOR U9697 ( .A(n9559), .B(n9560), .Z(n9561) );
  NANDN U9698 ( .A(n9449), .B(n9448), .Z(n9453) );
  NAND U9699 ( .A(n9451), .B(n9450), .Z(n9452) );
  AND U9700 ( .A(n9453), .B(n9452), .Z(n9562) );
  XNOR U9701 ( .A(n9561), .B(n9562), .Z(n9506) );
  NANDN U9702 ( .A(n9455), .B(n9454), .Z(n9459) );
  OR U9703 ( .A(n9457), .B(n9456), .Z(n9458) );
  NAND U9704 ( .A(n9459), .B(n9458), .Z(n9556) );
  NAND U9705 ( .A(b[0]), .B(a[128]), .Z(n9460) );
  XNOR U9706 ( .A(b[1]), .B(n9460), .Z(n9462) );
  NAND U9707 ( .A(a[127]), .B(n98), .Z(n9461) );
  AND U9708 ( .A(n9462), .B(n9461), .Z(n9532) );
  XNOR U9709 ( .A(n20154), .B(n9591), .Z(n9541) );
  OR U9710 ( .A(n9541), .B(n20057), .Z(n9465) );
  NANDN U9711 ( .A(n9463), .B(n20098), .Z(n9464) );
  AND U9712 ( .A(n9465), .B(n9464), .Z(n9533) );
  XOR U9713 ( .A(n9532), .B(n9533), .Z(n9535) );
  NAND U9714 ( .A(a[112]), .B(b[15]), .Z(n9534) );
  XOR U9715 ( .A(n9535), .B(n9534), .Z(n9553) );
  NAND U9716 ( .A(n19722), .B(n9466), .Z(n9468) );
  XNOR U9717 ( .A(b[5]), .B(n10213), .Z(n9544) );
  NANDN U9718 ( .A(n19640), .B(n9544), .Z(n9467) );
  NAND U9719 ( .A(n9468), .B(n9467), .Z(n9529) );
  XNOR U9720 ( .A(n19714), .B(n10084), .Z(n9547) );
  NANDN U9721 ( .A(n9547), .B(n19766), .Z(n9471) );
  NANDN U9722 ( .A(n9469), .B(n19767), .Z(n9470) );
  NAND U9723 ( .A(n9471), .B(n9470), .Z(n9526) );
  NAND U9724 ( .A(n19554), .B(n9472), .Z(n9474) );
  IV U9725 ( .A(a[126]), .Z(n10369) );
  XNOR U9726 ( .A(b[3]), .B(n10369), .Z(n9550) );
  NANDN U9727 ( .A(n19521), .B(n9550), .Z(n9473) );
  AND U9728 ( .A(n9474), .B(n9473), .Z(n9527) );
  XNOR U9729 ( .A(n9526), .B(n9527), .Z(n9528) );
  XOR U9730 ( .A(n9529), .B(n9528), .Z(n9554) );
  XOR U9731 ( .A(n9553), .B(n9554), .Z(n9555) );
  XNOR U9732 ( .A(n9556), .B(n9555), .Z(n9504) );
  NAND U9733 ( .A(n9476), .B(n9475), .Z(n9480) );
  NAND U9734 ( .A(n9478), .B(n9477), .Z(n9479) );
  NAND U9735 ( .A(n9480), .B(n9479), .Z(n9505) );
  XOR U9736 ( .A(n9504), .B(n9505), .Z(n9507) );
  XNOR U9737 ( .A(n9506), .B(n9507), .Z(n9565) );
  NANDN U9738 ( .A(n9482), .B(n9481), .Z(n9486) );
  NAND U9739 ( .A(n9484), .B(n9483), .Z(n9485) );
  NAND U9740 ( .A(n9486), .B(n9485), .Z(n9566) );
  XNOR U9741 ( .A(n9565), .B(n9566), .Z(n9567) );
  XOR U9742 ( .A(n9568), .B(n9567), .Z(n9498) );
  NANDN U9743 ( .A(n9488), .B(n9487), .Z(n9492) );
  NANDN U9744 ( .A(n9490), .B(n9489), .Z(n9491) );
  NAND U9745 ( .A(n9492), .B(n9491), .Z(n9499) );
  XNOR U9746 ( .A(n9498), .B(n9499), .Z(n9500) );
  XNOR U9747 ( .A(n9501), .B(n9500), .Z(n9571) );
  XNOR U9748 ( .A(n9571), .B(sreg[368]), .Z(n9573) );
  NAND U9749 ( .A(n9493), .B(sreg[367]), .Z(n9497) );
  OR U9750 ( .A(n9495), .B(n9494), .Z(n9496) );
  AND U9751 ( .A(n9497), .B(n9496), .Z(n9572) );
  XOR U9752 ( .A(n9573), .B(n9572), .Z(c[368]) );
  NANDN U9753 ( .A(n9499), .B(n9498), .Z(n9503) );
  NAND U9754 ( .A(n9501), .B(n9500), .Z(n9502) );
  NAND U9755 ( .A(n9503), .B(n9502), .Z(n9579) );
  NANDN U9756 ( .A(n9505), .B(n9504), .Z(n9509) );
  OR U9757 ( .A(n9507), .B(n9506), .Z(n9508) );
  NAND U9758 ( .A(n9509), .B(n9508), .Z(n9646) );
  XNOR U9759 ( .A(n20052), .B(n9852), .Z(n9588) );
  OR U9760 ( .A(n9588), .B(n20020), .Z(n9512) );
  NANDN U9761 ( .A(n9510), .B(n19960), .Z(n9511) );
  NAND U9762 ( .A(n9512), .B(n9511), .Z(n9601) );
  XNOR U9763 ( .A(n102), .B(n9513), .Z(n9592) );
  OR U9764 ( .A(n9592), .B(n20121), .Z(n9516) );
  NANDN U9765 ( .A(n9514), .B(n20122), .Z(n9515) );
  NAND U9766 ( .A(n9516), .B(n9515), .Z(n9598) );
  XNOR U9767 ( .A(n19975), .B(n10006), .Z(n9595) );
  NANDN U9768 ( .A(n9595), .B(n19883), .Z(n9519) );
  NANDN U9769 ( .A(n9517), .B(n19937), .Z(n9518) );
  AND U9770 ( .A(n9519), .B(n9518), .Z(n9599) );
  XNOR U9771 ( .A(n9598), .B(n9599), .Z(n9600) );
  XNOR U9772 ( .A(n9601), .B(n9600), .Z(n9637) );
  NANDN U9773 ( .A(n9521), .B(n9520), .Z(n9525) );
  NAND U9774 ( .A(n9523), .B(n9522), .Z(n9524) );
  NAND U9775 ( .A(n9525), .B(n9524), .Z(n9638) );
  XNOR U9776 ( .A(n9637), .B(n9638), .Z(n9639) );
  NANDN U9777 ( .A(n9527), .B(n9526), .Z(n9531) );
  NAND U9778 ( .A(n9529), .B(n9528), .Z(n9530) );
  AND U9779 ( .A(n9531), .B(n9530), .Z(n9640) );
  XNOR U9780 ( .A(n9639), .B(n9640), .Z(n9584) );
  NANDN U9781 ( .A(n9533), .B(n9532), .Z(n9537) );
  OR U9782 ( .A(n9535), .B(n9534), .Z(n9536) );
  NAND U9783 ( .A(n9537), .B(n9536), .Z(n9634) );
  NAND U9784 ( .A(b[0]), .B(a[129]), .Z(n9538) );
  XNOR U9785 ( .A(b[1]), .B(n9538), .Z(n9540) );
  NAND U9786 ( .A(a[128]), .B(n98), .Z(n9539) );
  AND U9787 ( .A(n9540), .B(n9539), .Z(n9610) );
  XNOR U9788 ( .A(n20154), .B(n9669), .Z(n9619) );
  OR U9789 ( .A(n9619), .B(n20057), .Z(n9543) );
  NANDN U9790 ( .A(n9541), .B(n20098), .Z(n9542) );
  AND U9791 ( .A(n9543), .B(n9542), .Z(n9611) );
  XOR U9792 ( .A(n9610), .B(n9611), .Z(n9613) );
  NAND U9793 ( .A(a[113]), .B(b[15]), .Z(n9612) );
  XOR U9794 ( .A(n9613), .B(n9612), .Z(n9631) );
  NAND U9795 ( .A(n19722), .B(n9544), .Z(n9546) );
  XNOR U9796 ( .A(b[5]), .B(n10291), .Z(n9622) );
  NANDN U9797 ( .A(n19640), .B(n9622), .Z(n9545) );
  NAND U9798 ( .A(n9546), .B(n9545), .Z(n9607) );
  XNOR U9799 ( .A(n19714), .B(n10135), .Z(n9625) );
  NANDN U9800 ( .A(n9625), .B(n19766), .Z(n9549) );
  NANDN U9801 ( .A(n9547), .B(n19767), .Z(n9548) );
  NAND U9802 ( .A(n9549), .B(n9548), .Z(n9604) );
  NAND U9803 ( .A(n19554), .B(n9550), .Z(n9552) );
  IV U9804 ( .A(a[127]), .Z(n10474) );
  XNOR U9805 ( .A(b[3]), .B(n10474), .Z(n9628) );
  NANDN U9806 ( .A(n19521), .B(n9628), .Z(n9551) );
  AND U9807 ( .A(n9552), .B(n9551), .Z(n9605) );
  XNOR U9808 ( .A(n9604), .B(n9605), .Z(n9606) );
  XOR U9809 ( .A(n9607), .B(n9606), .Z(n9632) );
  XOR U9810 ( .A(n9631), .B(n9632), .Z(n9633) );
  XNOR U9811 ( .A(n9634), .B(n9633), .Z(n9582) );
  NAND U9812 ( .A(n9554), .B(n9553), .Z(n9558) );
  NAND U9813 ( .A(n9556), .B(n9555), .Z(n9557) );
  NAND U9814 ( .A(n9558), .B(n9557), .Z(n9583) );
  XOR U9815 ( .A(n9582), .B(n9583), .Z(n9585) );
  XNOR U9816 ( .A(n9584), .B(n9585), .Z(n9643) );
  NANDN U9817 ( .A(n9560), .B(n9559), .Z(n9564) );
  NAND U9818 ( .A(n9562), .B(n9561), .Z(n9563) );
  NAND U9819 ( .A(n9564), .B(n9563), .Z(n9644) );
  XNOR U9820 ( .A(n9643), .B(n9644), .Z(n9645) );
  XOR U9821 ( .A(n9646), .B(n9645), .Z(n9576) );
  NANDN U9822 ( .A(n9566), .B(n9565), .Z(n9570) );
  NANDN U9823 ( .A(n9568), .B(n9567), .Z(n9569) );
  NAND U9824 ( .A(n9570), .B(n9569), .Z(n9577) );
  XNOR U9825 ( .A(n9576), .B(n9577), .Z(n9578) );
  XNOR U9826 ( .A(n9579), .B(n9578), .Z(n9649) );
  XNOR U9827 ( .A(n9649), .B(sreg[369]), .Z(n9651) );
  NAND U9828 ( .A(n9571), .B(sreg[368]), .Z(n9575) );
  OR U9829 ( .A(n9573), .B(n9572), .Z(n9574) );
  AND U9830 ( .A(n9575), .B(n9574), .Z(n9650) );
  XOR U9831 ( .A(n9651), .B(n9650), .Z(c[369]) );
  NANDN U9832 ( .A(n9577), .B(n9576), .Z(n9581) );
  NAND U9833 ( .A(n9579), .B(n9578), .Z(n9580) );
  NAND U9834 ( .A(n9581), .B(n9580), .Z(n9657) );
  NANDN U9835 ( .A(n9583), .B(n9582), .Z(n9587) );
  OR U9836 ( .A(n9585), .B(n9584), .Z(n9586) );
  NAND U9837 ( .A(n9587), .B(n9586), .Z(n9724) );
  XNOR U9838 ( .A(n20052), .B(n9903), .Z(n9666) );
  OR U9839 ( .A(n9666), .B(n20020), .Z(n9590) );
  NANDN U9840 ( .A(n9588), .B(n19960), .Z(n9589) );
  NAND U9841 ( .A(n9590), .B(n9589), .Z(n9679) );
  XNOR U9842 ( .A(n102), .B(n9591), .Z(n9670) );
  OR U9843 ( .A(n9670), .B(n20121), .Z(n9594) );
  NANDN U9844 ( .A(n9592), .B(n20122), .Z(n9593) );
  NAND U9845 ( .A(n9594), .B(n9593), .Z(n9676) );
  XNOR U9846 ( .A(n19975), .B(n10084), .Z(n9673) );
  NANDN U9847 ( .A(n9673), .B(n19883), .Z(n9597) );
  NANDN U9848 ( .A(n9595), .B(n19937), .Z(n9596) );
  AND U9849 ( .A(n9597), .B(n9596), .Z(n9677) );
  XNOR U9850 ( .A(n9676), .B(n9677), .Z(n9678) );
  XNOR U9851 ( .A(n9679), .B(n9678), .Z(n9715) );
  NANDN U9852 ( .A(n9599), .B(n9598), .Z(n9603) );
  NAND U9853 ( .A(n9601), .B(n9600), .Z(n9602) );
  NAND U9854 ( .A(n9603), .B(n9602), .Z(n9716) );
  XNOR U9855 ( .A(n9715), .B(n9716), .Z(n9717) );
  NANDN U9856 ( .A(n9605), .B(n9604), .Z(n9609) );
  NAND U9857 ( .A(n9607), .B(n9606), .Z(n9608) );
  AND U9858 ( .A(n9609), .B(n9608), .Z(n9718) );
  XNOR U9859 ( .A(n9717), .B(n9718), .Z(n9662) );
  NANDN U9860 ( .A(n9611), .B(n9610), .Z(n9615) );
  OR U9861 ( .A(n9613), .B(n9612), .Z(n9614) );
  NAND U9862 ( .A(n9615), .B(n9614), .Z(n9712) );
  NAND U9863 ( .A(b[0]), .B(a[130]), .Z(n9616) );
  XNOR U9864 ( .A(b[1]), .B(n9616), .Z(n9618) );
  NAND U9865 ( .A(a[129]), .B(n98), .Z(n9617) );
  AND U9866 ( .A(n9618), .B(n9617), .Z(n9688) );
  XNOR U9867 ( .A(n20154), .B(n9747), .Z(n9694) );
  OR U9868 ( .A(n9694), .B(n20057), .Z(n9621) );
  NANDN U9869 ( .A(n9619), .B(n20098), .Z(n9620) );
  AND U9870 ( .A(n9621), .B(n9620), .Z(n9689) );
  XOR U9871 ( .A(n9688), .B(n9689), .Z(n9691) );
  NAND U9872 ( .A(a[114]), .B(b[15]), .Z(n9690) );
  XOR U9873 ( .A(n9691), .B(n9690), .Z(n9709) );
  NAND U9874 ( .A(n19722), .B(n9622), .Z(n9624) );
  XNOR U9875 ( .A(b[5]), .B(n10369), .Z(n9700) );
  NANDN U9876 ( .A(n19640), .B(n9700), .Z(n9623) );
  NAND U9877 ( .A(n9624), .B(n9623), .Z(n9685) );
  XNOR U9878 ( .A(n19714), .B(n10213), .Z(n9703) );
  NANDN U9879 ( .A(n9703), .B(n19766), .Z(n9627) );
  NANDN U9880 ( .A(n9625), .B(n19767), .Z(n9626) );
  NAND U9881 ( .A(n9627), .B(n9626), .Z(n9682) );
  NAND U9882 ( .A(n19554), .B(n9628), .Z(n9630) );
  IV U9883 ( .A(a[128]), .Z(n10525) );
  XNOR U9884 ( .A(b[3]), .B(n10525), .Z(n9706) );
  NANDN U9885 ( .A(n19521), .B(n9706), .Z(n9629) );
  AND U9886 ( .A(n9630), .B(n9629), .Z(n9683) );
  XNOR U9887 ( .A(n9682), .B(n9683), .Z(n9684) );
  XOR U9888 ( .A(n9685), .B(n9684), .Z(n9710) );
  XOR U9889 ( .A(n9709), .B(n9710), .Z(n9711) );
  XNOR U9890 ( .A(n9712), .B(n9711), .Z(n9660) );
  NAND U9891 ( .A(n9632), .B(n9631), .Z(n9636) );
  NAND U9892 ( .A(n9634), .B(n9633), .Z(n9635) );
  NAND U9893 ( .A(n9636), .B(n9635), .Z(n9661) );
  XOR U9894 ( .A(n9660), .B(n9661), .Z(n9663) );
  XNOR U9895 ( .A(n9662), .B(n9663), .Z(n9721) );
  NANDN U9896 ( .A(n9638), .B(n9637), .Z(n9642) );
  NAND U9897 ( .A(n9640), .B(n9639), .Z(n9641) );
  NAND U9898 ( .A(n9642), .B(n9641), .Z(n9722) );
  XNOR U9899 ( .A(n9721), .B(n9722), .Z(n9723) );
  XOR U9900 ( .A(n9724), .B(n9723), .Z(n9654) );
  NANDN U9901 ( .A(n9644), .B(n9643), .Z(n9648) );
  NANDN U9902 ( .A(n9646), .B(n9645), .Z(n9647) );
  NAND U9903 ( .A(n9648), .B(n9647), .Z(n9655) );
  XNOR U9904 ( .A(n9654), .B(n9655), .Z(n9656) );
  XNOR U9905 ( .A(n9657), .B(n9656), .Z(n9727) );
  XNOR U9906 ( .A(n9727), .B(sreg[370]), .Z(n9729) );
  NAND U9907 ( .A(n9649), .B(sreg[369]), .Z(n9653) );
  OR U9908 ( .A(n9651), .B(n9650), .Z(n9652) );
  AND U9909 ( .A(n9653), .B(n9652), .Z(n9728) );
  XOR U9910 ( .A(n9729), .B(n9728), .Z(c[370]) );
  NANDN U9911 ( .A(n9655), .B(n9654), .Z(n9659) );
  NAND U9912 ( .A(n9657), .B(n9656), .Z(n9658) );
  NAND U9913 ( .A(n9659), .B(n9658), .Z(n9735) );
  NANDN U9914 ( .A(n9661), .B(n9660), .Z(n9665) );
  OR U9915 ( .A(n9663), .B(n9662), .Z(n9664) );
  NAND U9916 ( .A(n9665), .B(n9664), .Z(n9802) );
  XNOR U9917 ( .A(n20052), .B(n10006), .Z(n9744) );
  OR U9918 ( .A(n9744), .B(n20020), .Z(n9668) );
  NANDN U9919 ( .A(n9666), .B(n19960), .Z(n9667) );
  NAND U9920 ( .A(n9668), .B(n9667), .Z(n9757) );
  XNOR U9921 ( .A(n102), .B(n9669), .Z(n9748) );
  OR U9922 ( .A(n9748), .B(n20121), .Z(n9672) );
  NANDN U9923 ( .A(n9670), .B(n20122), .Z(n9671) );
  NAND U9924 ( .A(n9672), .B(n9671), .Z(n9754) );
  XNOR U9925 ( .A(n19975), .B(n10135), .Z(n9751) );
  NANDN U9926 ( .A(n9751), .B(n19883), .Z(n9675) );
  NANDN U9927 ( .A(n9673), .B(n19937), .Z(n9674) );
  AND U9928 ( .A(n9675), .B(n9674), .Z(n9755) );
  XNOR U9929 ( .A(n9754), .B(n9755), .Z(n9756) );
  XNOR U9930 ( .A(n9757), .B(n9756), .Z(n9793) );
  NANDN U9931 ( .A(n9677), .B(n9676), .Z(n9681) );
  NAND U9932 ( .A(n9679), .B(n9678), .Z(n9680) );
  NAND U9933 ( .A(n9681), .B(n9680), .Z(n9794) );
  XNOR U9934 ( .A(n9793), .B(n9794), .Z(n9795) );
  NANDN U9935 ( .A(n9683), .B(n9682), .Z(n9687) );
  NAND U9936 ( .A(n9685), .B(n9684), .Z(n9686) );
  AND U9937 ( .A(n9687), .B(n9686), .Z(n9796) );
  XNOR U9938 ( .A(n9795), .B(n9796), .Z(n9740) );
  NANDN U9939 ( .A(n9689), .B(n9688), .Z(n9693) );
  OR U9940 ( .A(n9691), .B(n9690), .Z(n9692) );
  NAND U9941 ( .A(n9693), .B(n9692), .Z(n9790) );
  XNOR U9942 ( .A(n20154), .B(n9852), .Z(n9772) );
  OR U9943 ( .A(n9772), .B(n20057), .Z(n9696) );
  NANDN U9944 ( .A(n9694), .B(n20098), .Z(n9695) );
  AND U9945 ( .A(n9696), .B(n9695), .Z(n9767) );
  NAND U9946 ( .A(b[0]), .B(a[131]), .Z(n9697) );
  XNOR U9947 ( .A(b[1]), .B(n9697), .Z(n9699) );
  NAND U9948 ( .A(a[130]), .B(n98), .Z(n9698) );
  AND U9949 ( .A(n9699), .B(n9698), .Z(n9766) );
  XOR U9950 ( .A(n9767), .B(n9766), .Z(n9769) );
  NAND U9951 ( .A(a[115]), .B(b[15]), .Z(n9768) );
  XOR U9952 ( .A(n9769), .B(n9768), .Z(n9787) );
  NAND U9953 ( .A(n19722), .B(n9700), .Z(n9702) );
  XNOR U9954 ( .A(b[5]), .B(n10474), .Z(n9778) );
  NANDN U9955 ( .A(n19640), .B(n9778), .Z(n9701) );
  NAND U9956 ( .A(n9702), .B(n9701), .Z(n9763) );
  XNOR U9957 ( .A(n19714), .B(n10291), .Z(n9781) );
  NANDN U9958 ( .A(n9781), .B(n19766), .Z(n9705) );
  NANDN U9959 ( .A(n9703), .B(n19767), .Z(n9704) );
  NAND U9960 ( .A(n9705), .B(n9704), .Z(n9760) );
  NAND U9961 ( .A(n19554), .B(n9706), .Z(n9708) );
  IV U9962 ( .A(a[129]), .Z(n10630) );
  XNOR U9963 ( .A(b[3]), .B(n10630), .Z(n9784) );
  NANDN U9964 ( .A(n19521), .B(n9784), .Z(n9707) );
  AND U9965 ( .A(n9708), .B(n9707), .Z(n9761) );
  XNOR U9966 ( .A(n9760), .B(n9761), .Z(n9762) );
  XOR U9967 ( .A(n9763), .B(n9762), .Z(n9788) );
  XOR U9968 ( .A(n9787), .B(n9788), .Z(n9789) );
  XNOR U9969 ( .A(n9790), .B(n9789), .Z(n9738) );
  NAND U9970 ( .A(n9710), .B(n9709), .Z(n9714) );
  NAND U9971 ( .A(n9712), .B(n9711), .Z(n9713) );
  NAND U9972 ( .A(n9714), .B(n9713), .Z(n9739) );
  XOR U9973 ( .A(n9738), .B(n9739), .Z(n9741) );
  XNOR U9974 ( .A(n9740), .B(n9741), .Z(n9799) );
  NANDN U9975 ( .A(n9716), .B(n9715), .Z(n9720) );
  NAND U9976 ( .A(n9718), .B(n9717), .Z(n9719) );
  NAND U9977 ( .A(n9720), .B(n9719), .Z(n9800) );
  XNOR U9978 ( .A(n9799), .B(n9800), .Z(n9801) );
  XOR U9979 ( .A(n9802), .B(n9801), .Z(n9732) );
  NANDN U9980 ( .A(n9722), .B(n9721), .Z(n9726) );
  NANDN U9981 ( .A(n9724), .B(n9723), .Z(n9725) );
  NAND U9982 ( .A(n9726), .B(n9725), .Z(n9733) );
  XNOR U9983 ( .A(n9732), .B(n9733), .Z(n9734) );
  XNOR U9984 ( .A(n9735), .B(n9734), .Z(n9805) );
  XNOR U9985 ( .A(n9805), .B(sreg[371]), .Z(n9807) );
  NAND U9986 ( .A(n9727), .B(sreg[370]), .Z(n9731) );
  OR U9987 ( .A(n9729), .B(n9728), .Z(n9730) );
  AND U9988 ( .A(n9731), .B(n9730), .Z(n9806) );
  XOR U9989 ( .A(n9807), .B(n9806), .Z(c[371]) );
  NANDN U9990 ( .A(n9733), .B(n9732), .Z(n9737) );
  NAND U9991 ( .A(n9735), .B(n9734), .Z(n9736) );
  NAND U9992 ( .A(n9737), .B(n9736), .Z(n9813) );
  NANDN U9993 ( .A(n9739), .B(n9738), .Z(n9743) );
  OR U9994 ( .A(n9741), .B(n9740), .Z(n9742) );
  NAND U9995 ( .A(n9743), .B(n9742), .Z(n9880) );
  XNOR U9996 ( .A(n20052), .B(n10084), .Z(n9849) );
  OR U9997 ( .A(n9849), .B(n20020), .Z(n9746) );
  NANDN U9998 ( .A(n9744), .B(n19960), .Z(n9745) );
  NAND U9999 ( .A(n9746), .B(n9745), .Z(n9862) );
  XNOR U10000 ( .A(n102), .B(n9747), .Z(n9853) );
  OR U10001 ( .A(n9853), .B(n20121), .Z(n9750) );
  NANDN U10002 ( .A(n9748), .B(n20122), .Z(n9749) );
  NAND U10003 ( .A(n9750), .B(n9749), .Z(n9859) );
  XNOR U10004 ( .A(n19975), .B(n10213), .Z(n9856) );
  NANDN U10005 ( .A(n9856), .B(n19883), .Z(n9753) );
  NANDN U10006 ( .A(n9751), .B(n19937), .Z(n9752) );
  AND U10007 ( .A(n9753), .B(n9752), .Z(n9860) );
  XNOR U10008 ( .A(n9859), .B(n9860), .Z(n9861) );
  XNOR U10009 ( .A(n9862), .B(n9861), .Z(n9871) );
  NANDN U10010 ( .A(n9755), .B(n9754), .Z(n9759) );
  NAND U10011 ( .A(n9757), .B(n9756), .Z(n9758) );
  NAND U10012 ( .A(n9759), .B(n9758), .Z(n9872) );
  XNOR U10013 ( .A(n9871), .B(n9872), .Z(n9873) );
  NANDN U10014 ( .A(n9761), .B(n9760), .Z(n9765) );
  NAND U10015 ( .A(n9763), .B(n9762), .Z(n9764) );
  AND U10016 ( .A(n9765), .B(n9764), .Z(n9874) );
  XNOR U10017 ( .A(n9873), .B(n9874), .Z(n9818) );
  NANDN U10018 ( .A(n9767), .B(n9766), .Z(n9771) );
  OR U10019 ( .A(n9769), .B(n9768), .Z(n9770) );
  NAND U10020 ( .A(n9771), .B(n9770), .Z(n9846) );
  XNOR U10021 ( .A(n20154), .B(n9903), .Z(n9828) );
  OR U10022 ( .A(n9828), .B(n20057), .Z(n9774) );
  NANDN U10023 ( .A(n9772), .B(n20098), .Z(n9773) );
  AND U10024 ( .A(n9774), .B(n9773), .Z(n9823) );
  NAND U10025 ( .A(b[0]), .B(a[132]), .Z(n9775) );
  XNOR U10026 ( .A(b[1]), .B(n9775), .Z(n9777) );
  NAND U10027 ( .A(a[131]), .B(n98), .Z(n9776) );
  AND U10028 ( .A(n9777), .B(n9776), .Z(n9822) );
  XOR U10029 ( .A(n9823), .B(n9822), .Z(n9825) );
  NAND U10030 ( .A(a[116]), .B(b[15]), .Z(n9824) );
  XOR U10031 ( .A(n9825), .B(n9824), .Z(n9843) );
  NAND U10032 ( .A(n19722), .B(n9778), .Z(n9780) );
  XNOR U10033 ( .A(b[5]), .B(n10525), .Z(n9834) );
  NANDN U10034 ( .A(n19640), .B(n9834), .Z(n9779) );
  NAND U10035 ( .A(n9780), .B(n9779), .Z(n9868) );
  XNOR U10036 ( .A(n19714), .B(n10369), .Z(n9837) );
  NANDN U10037 ( .A(n9837), .B(n19766), .Z(n9783) );
  NANDN U10038 ( .A(n9781), .B(n19767), .Z(n9782) );
  NAND U10039 ( .A(n9783), .B(n9782), .Z(n9865) );
  NAND U10040 ( .A(n19554), .B(n9784), .Z(n9786) );
  IV U10041 ( .A(a[130]), .Z(n10708) );
  XNOR U10042 ( .A(b[3]), .B(n10708), .Z(n9840) );
  NANDN U10043 ( .A(n19521), .B(n9840), .Z(n9785) );
  AND U10044 ( .A(n9786), .B(n9785), .Z(n9866) );
  XNOR U10045 ( .A(n9865), .B(n9866), .Z(n9867) );
  XOR U10046 ( .A(n9868), .B(n9867), .Z(n9844) );
  XOR U10047 ( .A(n9843), .B(n9844), .Z(n9845) );
  XNOR U10048 ( .A(n9846), .B(n9845), .Z(n9816) );
  NAND U10049 ( .A(n9788), .B(n9787), .Z(n9792) );
  NAND U10050 ( .A(n9790), .B(n9789), .Z(n9791) );
  NAND U10051 ( .A(n9792), .B(n9791), .Z(n9817) );
  XOR U10052 ( .A(n9816), .B(n9817), .Z(n9819) );
  XNOR U10053 ( .A(n9818), .B(n9819), .Z(n9877) );
  NANDN U10054 ( .A(n9794), .B(n9793), .Z(n9798) );
  NAND U10055 ( .A(n9796), .B(n9795), .Z(n9797) );
  NAND U10056 ( .A(n9798), .B(n9797), .Z(n9878) );
  XNOR U10057 ( .A(n9877), .B(n9878), .Z(n9879) );
  XOR U10058 ( .A(n9880), .B(n9879), .Z(n9810) );
  NANDN U10059 ( .A(n9800), .B(n9799), .Z(n9804) );
  NANDN U10060 ( .A(n9802), .B(n9801), .Z(n9803) );
  NAND U10061 ( .A(n9804), .B(n9803), .Z(n9811) );
  XNOR U10062 ( .A(n9810), .B(n9811), .Z(n9812) );
  XNOR U10063 ( .A(n9813), .B(n9812), .Z(n9883) );
  XNOR U10064 ( .A(n9883), .B(sreg[372]), .Z(n9885) );
  NAND U10065 ( .A(n9805), .B(sreg[371]), .Z(n9809) );
  OR U10066 ( .A(n9807), .B(n9806), .Z(n9808) );
  AND U10067 ( .A(n9809), .B(n9808), .Z(n9884) );
  XOR U10068 ( .A(n9885), .B(n9884), .Z(c[372]) );
  NANDN U10069 ( .A(n9811), .B(n9810), .Z(n9815) );
  NAND U10070 ( .A(n9813), .B(n9812), .Z(n9814) );
  NAND U10071 ( .A(n9815), .B(n9814), .Z(n9891) );
  NANDN U10072 ( .A(n9817), .B(n9816), .Z(n9821) );
  OR U10073 ( .A(n9819), .B(n9818), .Z(n9820) );
  NAND U10074 ( .A(n9821), .B(n9820), .Z(n9956) );
  NANDN U10075 ( .A(n9823), .B(n9822), .Z(n9827) );
  OR U10076 ( .A(n9825), .B(n9824), .Z(n9826) );
  NAND U10077 ( .A(n9827), .B(n9826), .Z(n9946) );
  XNOR U10078 ( .A(n20154), .B(n10006), .Z(n9931) );
  OR U10079 ( .A(n9931), .B(n20057), .Z(n9830) );
  NANDN U10080 ( .A(n9828), .B(n20098), .Z(n9829) );
  NAND U10081 ( .A(n9830), .B(n9829), .Z(n9922) );
  AND U10082 ( .A(a[133]), .B(b[0]), .Z(n9831) );
  XOR U10083 ( .A(b[1]), .B(n9831), .Z(n9833) );
  NAND U10084 ( .A(a[132]), .B(n98), .Z(n9832) );
  NAND U10085 ( .A(n9833), .B(n9832), .Z(n9923) );
  XNOR U10086 ( .A(n9922), .B(n9923), .Z(n9924) );
  NAND U10087 ( .A(a[117]), .B(b[15]), .Z(n9925) );
  XOR U10088 ( .A(n9924), .B(n9925), .Z(n9943) );
  NAND U10089 ( .A(n19722), .B(n9834), .Z(n9836) );
  XNOR U10090 ( .A(b[5]), .B(n10630), .Z(n9934) );
  NANDN U10091 ( .A(n19640), .B(n9934), .Z(n9835) );
  NAND U10092 ( .A(n9836), .B(n9835), .Z(n9919) );
  XNOR U10093 ( .A(n19714), .B(n10474), .Z(n9937) );
  NANDN U10094 ( .A(n9937), .B(n19766), .Z(n9839) );
  NANDN U10095 ( .A(n9837), .B(n19767), .Z(n9838) );
  NAND U10096 ( .A(n9839), .B(n9838), .Z(n9916) );
  NAND U10097 ( .A(n19554), .B(n9840), .Z(n9842) );
  IV U10098 ( .A(a[131]), .Z(n10786) );
  XNOR U10099 ( .A(b[3]), .B(n10786), .Z(n9940) );
  NANDN U10100 ( .A(n19521), .B(n9940), .Z(n9841) );
  AND U10101 ( .A(n9842), .B(n9841), .Z(n9917) );
  XNOR U10102 ( .A(n9916), .B(n9917), .Z(n9918) );
  XOR U10103 ( .A(n9919), .B(n9918), .Z(n9944) );
  XNOR U10104 ( .A(n9943), .B(n9944), .Z(n9945) );
  XNOR U10105 ( .A(n9946), .B(n9945), .Z(n9894) );
  NAND U10106 ( .A(n9844), .B(n9843), .Z(n9848) );
  NAND U10107 ( .A(n9846), .B(n9845), .Z(n9847) );
  NAND U10108 ( .A(n9848), .B(n9847), .Z(n9895) );
  XOR U10109 ( .A(n9894), .B(n9895), .Z(n9897) );
  XNOR U10110 ( .A(n20052), .B(n10135), .Z(n9900) );
  OR U10111 ( .A(n9900), .B(n20020), .Z(n9851) );
  NANDN U10112 ( .A(n9849), .B(n19960), .Z(n9850) );
  NAND U10113 ( .A(n9851), .B(n9850), .Z(n9913) );
  XNOR U10114 ( .A(n102), .B(n9852), .Z(n9904) );
  OR U10115 ( .A(n9904), .B(n20121), .Z(n9855) );
  NANDN U10116 ( .A(n9853), .B(n20122), .Z(n9854) );
  NAND U10117 ( .A(n9855), .B(n9854), .Z(n9910) );
  XNOR U10118 ( .A(n19975), .B(n10291), .Z(n9907) );
  NANDN U10119 ( .A(n9907), .B(n19883), .Z(n9858) );
  NANDN U10120 ( .A(n9856), .B(n19937), .Z(n9857) );
  AND U10121 ( .A(n9858), .B(n9857), .Z(n9911) );
  XNOR U10122 ( .A(n9910), .B(n9911), .Z(n9912) );
  XNOR U10123 ( .A(n9913), .B(n9912), .Z(n9947) );
  NANDN U10124 ( .A(n9860), .B(n9859), .Z(n9864) );
  NAND U10125 ( .A(n9862), .B(n9861), .Z(n9863) );
  NAND U10126 ( .A(n9864), .B(n9863), .Z(n9948) );
  XNOR U10127 ( .A(n9947), .B(n9948), .Z(n9949) );
  NANDN U10128 ( .A(n9866), .B(n9865), .Z(n9870) );
  NAND U10129 ( .A(n9868), .B(n9867), .Z(n9869) );
  AND U10130 ( .A(n9870), .B(n9869), .Z(n9950) );
  XNOR U10131 ( .A(n9949), .B(n9950), .Z(n9896) );
  XNOR U10132 ( .A(n9897), .B(n9896), .Z(n9953) );
  NANDN U10133 ( .A(n9872), .B(n9871), .Z(n9876) );
  NAND U10134 ( .A(n9874), .B(n9873), .Z(n9875) );
  NAND U10135 ( .A(n9876), .B(n9875), .Z(n9954) );
  XNOR U10136 ( .A(n9953), .B(n9954), .Z(n9955) );
  XOR U10137 ( .A(n9956), .B(n9955), .Z(n9888) );
  NANDN U10138 ( .A(n9878), .B(n9877), .Z(n9882) );
  NANDN U10139 ( .A(n9880), .B(n9879), .Z(n9881) );
  NAND U10140 ( .A(n9882), .B(n9881), .Z(n9889) );
  XNOR U10141 ( .A(n9888), .B(n9889), .Z(n9890) );
  XNOR U10142 ( .A(n9891), .B(n9890), .Z(n9959) );
  XNOR U10143 ( .A(n9959), .B(sreg[373]), .Z(n9961) );
  NAND U10144 ( .A(n9883), .B(sreg[372]), .Z(n9887) );
  OR U10145 ( .A(n9885), .B(n9884), .Z(n9886) );
  AND U10146 ( .A(n9887), .B(n9886), .Z(n9960) );
  XOR U10147 ( .A(n9961), .B(n9960), .Z(c[373]) );
  NANDN U10148 ( .A(n9889), .B(n9888), .Z(n9893) );
  NAND U10149 ( .A(n9891), .B(n9890), .Z(n9892) );
  NAND U10150 ( .A(n9893), .B(n9892), .Z(n9967) );
  NANDN U10151 ( .A(n9895), .B(n9894), .Z(n9899) );
  OR U10152 ( .A(n9897), .B(n9896), .Z(n9898) );
  NAND U10153 ( .A(n9899), .B(n9898), .Z(n10034) );
  XNOR U10154 ( .A(n20052), .B(n10213), .Z(n10003) );
  OR U10155 ( .A(n10003), .B(n20020), .Z(n9902) );
  NANDN U10156 ( .A(n9900), .B(n19960), .Z(n9901) );
  NAND U10157 ( .A(n9902), .B(n9901), .Z(n10016) );
  XNOR U10158 ( .A(n102), .B(n9903), .Z(n10007) );
  OR U10159 ( .A(n10007), .B(n20121), .Z(n9906) );
  NANDN U10160 ( .A(n9904), .B(n20122), .Z(n9905) );
  NAND U10161 ( .A(n9906), .B(n9905), .Z(n10013) );
  XNOR U10162 ( .A(n19975), .B(n10369), .Z(n10010) );
  NANDN U10163 ( .A(n10010), .B(n19883), .Z(n9909) );
  NANDN U10164 ( .A(n9907), .B(n19937), .Z(n9908) );
  AND U10165 ( .A(n9909), .B(n9908), .Z(n10014) );
  XNOR U10166 ( .A(n10013), .B(n10014), .Z(n10015) );
  XNOR U10167 ( .A(n10016), .B(n10015), .Z(n10025) );
  NANDN U10168 ( .A(n9911), .B(n9910), .Z(n9915) );
  NAND U10169 ( .A(n9913), .B(n9912), .Z(n9914) );
  NAND U10170 ( .A(n9915), .B(n9914), .Z(n10026) );
  XNOR U10171 ( .A(n10025), .B(n10026), .Z(n10027) );
  NANDN U10172 ( .A(n9917), .B(n9916), .Z(n9921) );
  NAND U10173 ( .A(n9919), .B(n9918), .Z(n9920) );
  AND U10174 ( .A(n9921), .B(n9920), .Z(n10028) );
  XNOR U10175 ( .A(n10027), .B(n10028), .Z(n9972) );
  NANDN U10176 ( .A(n9923), .B(n9922), .Z(n9927) );
  NANDN U10177 ( .A(n9925), .B(n9924), .Z(n9926) );
  NAND U10178 ( .A(n9927), .B(n9926), .Z(n10000) );
  NAND U10179 ( .A(b[0]), .B(a[134]), .Z(n9928) );
  XNOR U10180 ( .A(b[1]), .B(n9928), .Z(n9930) );
  NAND U10181 ( .A(a[133]), .B(n98), .Z(n9929) );
  AND U10182 ( .A(n9930), .B(n9929), .Z(n9976) );
  XNOR U10183 ( .A(n20154), .B(n10084), .Z(n9982) );
  OR U10184 ( .A(n9982), .B(n20057), .Z(n9933) );
  NANDN U10185 ( .A(n9931), .B(n20098), .Z(n9932) );
  AND U10186 ( .A(n9933), .B(n9932), .Z(n9977) );
  XOR U10187 ( .A(n9976), .B(n9977), .Z(n9979) );
  NAND U10188 ( .A(a[118]), .B(b[15]), .Z(n9978) );
  XOR U10189 ( .A(n9979), .B(n9978), .Z(n9997) );
  NAND U10190 ( .A(n19722), .B(n9934), .Z(n9936) );
  XNOR U10191 ( .A(b[5]), .B(n10708), .Z(n9988) );
  NANDN U10192 ( .A(n19640), .B(n9988), .Z(n9935) );
  NAND U10193 ( .A(n9936), .B(n9935), .Z(n10022) );
  XNOR U10194 ( .A(n19714), .B(n10525), .Z(n9991) );
  NANDN U10195 ( .A(n9991), .B(n19766), .Z(n9939) );
  NANDN U10196 ( .A(n9937), .B(n19767), .Z(n9938) );
  NAND U10197 ( .A(n9939), .B(n9938), .Z(n10019) );
  NAND U10198 ( .A(n19554), .B(n9940), .Z(n9942) );
  IV U10199 ( .A(a[132]), .Z(n10837) );
  XNOR U10200 ( .A(b[3]), .B(n10837), .Z(n9994) );
  NANDN U10201 ( .A(n19521), .B(n9994), .Z(n9941) );
  AND U10202 ( .A(n9942), .B(n9941), .Z(n10020) );
  XNOR U10203 ( .A(n10019), .B(n10020), .Z(n10021) );
  XOR U10204 ( .A(n10022), .B(n10021), .Z(n9998) );
  XOR U10205 ( .A(n9997), .B(n9998), .Z(n9999) );
  XNOR U10206 ( .A(n10000), .B(n9999), .Z(n9970) );
  XOR U10207 ( .A(n9970), .B(n9971), .Z(n9973) );
  XNOR U10208 ( .A(n9972), .B(n9973), .Z(n10031) );
  NANDN U10209 ( .A(n9948), .B(n9947), .Z(n9952) );
  NAND U10210 ( .A(n9950), .B(n9949), .Z(n9951) );
  NAND U10211 ( .A(n9952), .B(n9951), .Z(n10032) );
  XNOR U10212 ( .A(n10031), .B(n10032), .Z(n10033) );
  XOR U10213 ( .A(n10034), .B(n10033), .Z(n9964) );
  NANDN U10214 ( .A(n9954), .B(n9953), .Z(n9958) );
  NANDN U10215 ( .A(n9956), .B(n9955), .Z(n9957) );
  NAND U10216 ( .A(n9958), .B(n9957), .Z(n9965) );
  XNOR U10217 ( .A(n9964), .B(n9965), .Z(n9966) );
  XNOR U10218 ( .A(n9967), .B(n9966), .Z(n10037) );
  XNOR U10219 ( .A(n10037), .B(sreg[374]), .Z(n10039) );
  NAND U10220 ( .A(n9959), .B(sreg[373]), .Z(n9963) );
  OR U10221 ( .A(n9961), .B(n9960), .Z(n9962) );
  AND U10222 ( .A(n9963), .B(n9962), .Z(n10038) );
  XOR U10223 ( .A(n10039), .B(n10038), .Z(c[374]) );
  NANDN U10224 ( .A(n9965), .B(n9964), .Z(n9969) );
  NAND U10225 ( .A(n9967), .B(n9966), .Z(n9968) );
  NAND U10226 ( .A(n9969), .B(n9968), .Z(n10045) );
  NANDN U10227 ( .A(n9971), .B(n9970), .Z(n9975) );
  OR U10228 ( .A(n9973), .B(n9972), .Z(n9974) );
  NAND U10229 ( .A(n9975), .B(n9974), .Z(n10112) );
  NANDN U10230 ( .A(n9977), .B(n9976), .Z(n9981) );
  OR U10231 ( .A(n9979), .B(n9978), .Z(n9980) );
  NAND U10232 ( .A(n9981), .B(n9980), .Z(n10078) );
  XNOR U10233 ( .A(n20154), .B(n10135), .Z(n10063) );
  OR U10234 ( .A(n10063), .B(n20057), .Z(n9984) );
  NANDN U10235 ( .A(n9982), .B(n20098), .Z(n9983) );
  AND U10236 ( .A(n9984), .B(n9983), .Z(n10055) );
  NAND U10237 ( .A(b[0]), .B(a[135]), .Z(n9985) );
  XNOR U10238 ( .A(b[1]), .B(n9985), .Z(n9987) );
  NAND U10239 ( .A(a[134]), .B(n98), .Z(n9986) );
  AND U10240 ( .A(n9987), .B(n9986), .Z(n10054) );
  XOR U10241 ( .A(n10055), .B(n10054), .Z(n10057) );
  NAND U10242 ( .A(a[119]), .B(b[15]), .Z(n10056) );
  XOR U10243 ( .A(n10057), .B(n10056), .Z(n10075) );
  NAND U10244 ( .A(n19722), .B(n9988), .Z(n9990) );
  XNOR U10245 ( .A(b[5]), .B(n10786), .Z(n10066) );
  NANDN U10246 ( .A(n19640), .B(n10066), .Z(n9989) );
  NAND U10247 ( .A(n9990), .B(n9989), .Z(n10100) );
  XNOR U10248 ( .A(n19714), .B(n10630), .Z(n10069) );
  NANDN U10249 ( .A(n10069), .B(n19766), .Z(n9993) );
  NANDN U10250 ( .A(n9991), .B(n19767), .Z(n9992) );
  NAND U10251 ( .A(n9993), .B(n9992), .Z(n10097) );
  NAND U10252 ( .A(n19554), .B(n9994), .Z(n9996) );
  IV U10253 ( .A(a[133]), .Z(n10942) );
  XNOR U10254 ( .A(b[3]), .B(n10942), .Z(n10072) );
  NANDN U10255 ( .A(n19521), .B(n10072), .Z(n9995) );
  AND U10256 ( .A(n9996), .B(n9995), .Z(n10098) );
  XNOR U10257 ( .A(n10097), .B(n10098), .Z(n10099) );
  XOR U10258 ( .A(n10100), .B(n10099), .Z(n10076) );
  XOR U10259 ( .A(n10075), .B(n10076), .Z(n10077) );
  XNOR U10260 ( .A(n10078), .B(n10077), .Z(n10048) );
  NAND U10261 ( .A(n9998), .B(n9997), .Z(n10002) );
  NAND U10262 ( .A(n10000), .B(n9999), .Z(n10001) );
  NAND U10263 ( .A(n10002), .B(n10001), .Z(n10049) );
  XOR U10264 ( .A(n10048), .B(n10049), .Z(n10051) );
  XNOR U10265 ( .A(n20052), .B(n10291), .Z(n10081) );
  OR U10266 ( .A(n10081), .B(n20020), .Z(n10005) );
  NANDN U10267 ( .A(n10003), .B(n19960), .Z(n10004) );
  NAND U10268 ( .A(n10005), .B(n10004), .Z(n10094) );
  XNOR U10269 ( .A(n102), .B(n10006), .Z(n10085) );
  OR U10270 ( .A(n10085), .B(n20121), .Z(n10009) );
  NANDN U10271 ( .A(n10007), .B(n20122), .Z(n10008) );
  NAND U10272 ( .A(n10009), .B(n10008), .Z(n10091) );
  XNOR U10273 ( .A(n19975), .B(n10474), .Z(n10088) );
  NANDN U10274 ( .A(n10088), .B(n19883), .Z(n10012) );
  NANDN U10275 ( .A(n10010), .B(n19937), .Z(n10011) );
  AND U10276 ( .A(n10012), .B(n10011), .Z(n10092) );
  XNOR U10277 ( .A(n10091), .B(n10092), .Z(n10093) );
  XNOR U10278 ( .A(n10094), .B(n10093), .Z(n10103) );
  NANDN U10279 ( .A(n10014), .B(n10013), .Z(n10018) );
  NAND U10280 ( .A(n10016), .B(n10015), .Z(n10017) );
  NAND U10281 ( .A(n10018), .B(n10017), .Z(n10104) );
  XNOR U10282 ( .A(n10103), .B(n10104), .Z(n10105) );
  NANDN U10283 ( .A(n10020), .B(n10019), .Z(n10024) );
  NAND U10284 ( .A(n10022), .B(n10021), .Z(n10023) );
  AND U10285 ( .A(n10024), .B(n10023), .Z(n10106) );
  XNOR U10286 ( .A(n10105), .B(n10106), .Z(n10050) );
  XNOR U10287 ( .A(n10051), .B(n10050), .Z(n10109) );
  NANDN U10288 ( .A(n10026), .B(n10025), .Z(n10030) );
  NAND U10289 ( .A(n10028), .B(n10027), .Z(n10029) );
  NAND U10290 ( .A(n10030), .B(n10029), .Z(n10110) );
  XNOR U10291 ( .A(n10109), .B(n10110), .Z(n10111) );
  XOR U10292 ( .A(n10112), .B(n10111), .Z(n10042) );
  NANDN U10293 ( .A(n10032), .B(n10031), .Z(n10036) );
  NANDN U10294 ( .A(n10034), .B(n10033), .Z(n10035) );
  NAND U10295 ( .A(n10036), .B(n10035), .Z(n10043) );
  XNOR U10296 ( .A(n10042), .B(n10043), .Z(n10044) );
  XNOR U10297 ( .A(n10045), .B(n10044), .Z(n10115) );
  XNOR U10298 ( .A(n10115), .B(sreg[375]), .Z(n10117) );
  NAND U10299 ( .A(n10037), .B(sreg[374]), .Z(n10041) );
  OR U10300 ( .A(n10039), .B(n10038), .Z(n10040) );
  AND U10301 ( .A(n10041), .B(n10040), .Z(n10116) );
  XOR U10302 ( .A(n10117), .B(n10116), .Z(c[375]) );
  NANDN U10303 ( .A(n10043), .B(n10042), .Z(n10047) );
  NAND U10304 ( .A(n10045), .B(n10044), .Z(n10046) );
  NAND U10305 ( .A(n10047), .B(n10046), .Z(n10123) );
  NANDN U10306 ( .A(n10049), .B(n10048), .Z(n10053) );
  OR U10307 ( .A(n10051), .B(n10050), .Z(n10052) );
  NAND U10308 ( .A(n10053), .B(n10052), .Z(n10190) );
  NANDN U10309 ( .A(n10055), .B(n10054), .Z(n10059) );
  OR U10310 ( .A(n10057), .B(n10056), .Z(n10058) );
  NAND U10311 ( .A(n10059), .B(n10058), .Z(n10178) );
  NAND U10312 ( .A(b[0]), .B(a[136]), .Z(n10060) );
  XNOR U10313 ( .A(b[1]), .B(n10060), .Z(n10062) );
  NAND U10314 ( .A(a[135]), .B(n98), .Z(n10061) );
  AND U10315 ( .A(n10062), .B(n10061), .Z(n10154) );
  XNOR U10316 ( .A(n20154), .B(n10213), .Z(n10160) );
  OR U10317 ( .A(n10160), .B(n20057), .Z(n10065) );
  NANDN U10318 ( .A(n10063), .B(n20098), .Z(n10064) );
  AND U10319 ( .A(n10065), .B(n10064), .Z(n10155) );
  XOR U10320 ( .A(n10154), .B(n10155), .Z(n10157) );
  NAND U10321 ( .A(a[120]), .B(b[15]), .Z(n10156) );
  XOR U10322 ( .A(n10157), .B(n10156), .Z(n10175) );
  NAND U10323 ( .A(n19722), .B(n10066), .Z(n10068) );
  XNOR U10324 ( .A(b[5]), .B(n10837), .Z(n10166) );
  NANDN U10325 ( .A(n19640), .B(n10166), .Z(n10067) );
  NAND U10326 ( .A(n10068), .B(n10067), .Z(n10151) );
  XNOR U10327 ( .A(n19714), .B(n10708), .Z(n10169) );
  NANDN U10328 ( .A(n10169), .B(n19766), .Z(n10071) );
  NANDN U10329 ( .A(n10069), .B(n19767), .Z(n10070) );
  NAND U10330 ( .A(n10071), .B(n10070), .Z(n10148) );
  NAND U10331 ( .A(n19554), .B(n10072), .Z(n10074) );
  IV U10332 ( .A(a[134]), .Z(n11020) );
  XNOR U10333 ( .A(b[3]), .B(n11020), .Z(n10172) );
  NANDN U10334 ( .A(n19521), .B(n10172), .Z(n10073) );
  AND U10335 ( .A(n10074), .B(n10073), .Z(n10149) );
  XNOR U10336 ( .A(n10148), .B(n10149), .Z(n10150) );
  XOR U10337 ( .A(n10151), .B(n10150), .Z(n10176) );
  XOR U10338 ( .A(n10175), .B(n10176), .Z(n10177) );
  XNOR U10339 ( .A(n10178), .B(n10177), .Z(n10126) );
  NAND U10340 ( .A(n10076), .B(n10075), .Z(n10080) );
  NAND U10341 ( .A(n10078), .B(n10077), .Z(n10079) );
  NAND U10342 ( .A(n10080), .B(n10079), .Z(n10127) );
  XOR U10343 ( .A(n10126), .B(n10127), .Z(n10129) );
  XNOR U10344 ( .A(n20052), .B(n10369), .Z(n10132) );
  OR U10345 ( .A(n10132), .B(n20020), .Z(n10083) );
  NANDN U10346 ( .A(n10081), .B(n19960), .Z(n10082) );
  NAND U10347 ( .A(n10083), .B(n10082), .Z(n10145) );
  XNOR U10348 ( .A(n102), .B(n10084), .Z(n10136) );
  OR U10349 ( .A(n10136), .B(n20121), .Z(n10087) );
  NANDN U10350 ( .A(n10085), .B(n20122), .Z(n10086) );
  NAND U10351 ( .A(n10087), .B(n10086), .Z(n10142) );
  XNOR U10352 ( .A(n19975), .B(n10525), .Z(n10139) );
  NANDN U10353 ( .A(n10139), .B(n19883), .Z(n10090) );
  NANDN U10354 ( .A(n10088), .B(n19937), .Z(n10089) );
  AND U10355 ( .A(n10090), .B(n10089), .Z(n10143) );
  XNOR U10356 ( .A(n10142), .B(n10143), .Z(n10144) );
  XNOR U10357 ( .A(n10145), .B(n10144), .Z(n10181) );
  NANDN U10358 ( .A(n10092), .B(n10091), .Z(n10096) );
  NAND U10359 ( .A(n10094), .B(n10093), .Z(n10095) );
  NAND U10360 ( .A(n10096), .B(n10095), .Z(n10182) );
  XNOR U10361 ( .A(n10181), .B(n10182), .Z(n10183) );
  NANDN U10362 ( .A(n10098), .B(n10097), .Z(n10102) );
  NAND U10363 ( .A(n10100), .B(n10099), .Z(n10101) );
  AND U10364 ( .A(n10102), .B(n10101), .Z(n10184) );
  XNOR U10365 ( .A(n10183), .B(n10184), .Z(n10128) );
  XNOR U10366 ( .A(n10129), .B(n10128), .Z(n10187) );
  NANDN U10367 ( .A(n10104), .B(n10103), .Z(n10108) );
  NAND U10368 ( .A(n10106), .B(n10105), .Z(n10107) );
  NAND U10369 ( .A(n10108), .B(n10107), .Z(n10188) );
  XNOR U10370 ( .A(n10187), .B(n10188), .Z(n10189) );
  XOR U10371 ( .A(n10190), .B(n10189), .Z(n10120) );
  NANDN U10372 ( .A(n10110), .B(n10109), .Z(n10114) );
  NANDN U10373 ( .A(n10112), .B(n10111), .Z(n10113) );
  NAND U10374 ( .A(n10114), .B(n10113), .Z(n10121) );
  XNOR U10375 ( .A(n10120), .B(n10121), .Z(n10122) );
  XNOR U10376 ( .A(n10123), .B(n10122), .Z(n10193) );
  XNOR U10377 ( .A(n10193), .B(sreg[376]), .Z(n10195) );
  NAND U10378 ( .A(n10115), .B(sreg[375]), .Z(n10119) );
  OR U10379 ( .A(n10117), .B(n10116), .Z(n10118) );
  AND U10380 ( .A(n10119), .B(n10118), .Z(n10194) );
  XOR U10381 ( .A(n10195), .B(n10194), .Z(c[376]) );
  NANDN U10382 ( .A(n10121), .B(n10120), .Z(n10125) );
  NAND U10383 ( .A(n10123), .B(n10122), .Z(n10124) );
  NAND U10384 ( .A(n10125), .B(n10124), .Z(n10201) );
  NANDN U10385 ( .A(n10127), .B(n10126), .Z(n10131) );
  OR U10386 ( .A(n10129), .B(n10128), .Z(n10130) );
  NAND U10387 ( .A(n10131), .B(n10130), .Z(n10268) );
  XNOR U10388 ( .A(n20052), .B(n10474), .Z(n10210) );
  OR U10389 ( .A(n10210), .B(n20020), .Z(n10134) );
  NANDN U10390 ( .A(n10132), .B(n19960), .Z(n10133) );
  NAND U10391 ( .A(n10134), .B(n10133), .Z(n10223) );
  XNOR U10392 ( .A(n102), .B(n10135), .Z(n10214) );
  OR U10393 ( .A(n10214), .B(n20121), .Z(n10138) );
  NANDN U10394 ( .A(n10136), .B(n20122), .Z(n10137) );
  NAND U10395 ( .A(n10138), .B(n10137), .Z(n10220) );
  XNOR U10396 ( .A(n19975), .B(n10630), .Z(n10217) );
  NANDN U10397 ( .A(n10217), .B(n19883), .Z(n10141) );
  NANDN U10398 ( .A(n10139), .B(n19937), .Z(n10140) );
  AND U10399 ( .A(n10141), .B(n10140), .Z(n10221) );
  XNOR U10400 ( .A(n10220), .B(n10221), .Z(n10222) );
  XNOR U10401 ( .A(n10223), .B(n10222), .Z(n10259) );
  NANDN U10402 ( .A(n10143), .B(n10142), .Z(n10147) );
  NAND U10403 ( .A(n10145), .B(n10144), .Z(n10146) );
  NAND U10404 ( .A(n10147), .B(n10146), .Z(n10260) );
  XNOR U10405 ( .A(n10259), .B(n10260), .Z(n10261) );
  NANDN U10406 ( .A(n10149), .B(n10148), .Z(n10153) );
  NAND U10407 ( .A(n10151), .B(n10150), .Z(n10152) );
  AND U10408 ( .A(n10153), .B(n10152), .Z(n10262) );
  XNOR U10409 ( .A(n10261), .B(n10262), .Z(n10206) );
  NANDN U10410 ( .A(n10155), .B(n10154), .Z(n10159) );
  OR U10411 ( .A(n10157), .B(n10156), .Z(n10158) );
  NAND U10412 ( .A(n10159), .B(n10158), .Z(n10256) );
  XNOR U10413 ( .A(n20154), .B(n10291), .Z(n10241) );
  OR U10414 ( .A(n10241), .B(n20057), .Z(n10162) );
  NANDN U10415 ( .A(n10160), .B(n20098), .Z(n10161) );
  AND U10416 ( .A(n10162), .B(n10161), .Z(n10233) );
  NAND U10417 ( .A(b[0]), .B(a[137]), .Z(n10163) );
  XNOR U10418 ( .A(b[1]), .B(n10163), .Z(n10165) );
  NAND U10419 ( .A(a[136]), .B(n98), .Z(n10164) );
  AND U10420 ( .A(n10165), .B(n10164), .Z(n10232) );
  XOR U10421 ( .A(n10233), .B(n10232), .Z(n10235) );
  NAND U10422 ( .A(a[121]), .B(b[15]), .Z(n10234) );
  XOR U10423 ( .A(n10235), .B(n10234), .Z(n10253) );
  NAND U10424 ( .A(n19722), .B(n10166), .Z(n10168) );
  XNOR U10425 ( .A(b[5]), .B(n10942), .Z(n10244) );
  NANDN U10426 ( .A(n19640), .B(n10244), .Z(n10167) );
  NAND U10427 ( .A(n10168), .B(n10167), .Z(n10229) );
  XNOR U10428 ( .A(n19714), .B(n10786), .Z(n10247) );
  NANDN U10429 ( .A(n10247), .B(n19766), .Z(n10171) );
  NANDN U10430 ( .A(n10169), .B(n19767), .Z(n10170) );
  NAND U10431 ( .A(n10171), .B(n10170), .Z(n10226) );
  NAND U10432 ( .A(n19554), .B(n10172), .Z(n10174) );
  IV U10433 ( .A(a[135]), .Z(n11098) );
  XNOR U10434 ( .A(b[3]), .B(n11098), .Z(n10250) );
  NANDN U10435 ( .A(n19521), .B(n10250), .Z(n10173) );
  AND U10436 ( .A(n10174), .B(n10173), .Z(n10227) );
  XNOR U10437 ( .A(n10226), .B(n10227), .Z(n10228) );
  XOR U10438 ( .A(n10229), .B(n10228), .Z(n10254) );
  XOR U10439 ( .A(n10253), .B(n10254), .Z(n10255) );
  XNOR U10440 ( .A(n10256), .B(n10255), .Z(n10204) );
  NAND U10441 ( .A(n10176), .B(n10175), .Z(n10180) );
  NAND U10442 ( .A(n10178), .B(n10177), .Z(n10179) );
  NAND U10443 ( .A(n10180), .B(n10179), .Z(n10205) );
  XOR U10444 ( .A(n10204), .B(n10205), .Z(n10207) );
  XNOR U10445 ( .A(n10206), .B(n10207), .Z(n10265) );
  NANDN U10446 ( .A(n10182), .B(n10181), .Z(n10186) );
  NAND U10447 ( .A(n10184), .B(n10183), .Z(n10185) );
  NAND U10448 ( .A(n10186), .B(n10185), .Z(n10266) );
  XNOR U10449 ( .A(n10265), .B(n10266), .Z(n10267) );
  XOR U10450 ( .A(n10268), .B(n10267), .Z(n10198) );
  NANDN U10451 ( .A(n10188), .B(n10187), .Z(n10192) );
  NANDN U10452 ( .A(n10190), .B(n10189), .Z(n10191) );
  NAND U10453 ( .A(n10192), .B(n10191), .Z(n10199) );
  XNOR U10454 ( .A(n10198), .B(n10199), .Z(n10200) );
  XNOR U10455 ( .A(n10201), .B(n10200), .Z(n10271) );
  XNOR U10456 ( .A(n10271), .B(sreg[377]), .Z(n10273) );
  NAND U10457 ( .A(n10193), .B(sreg[376]), .Z(n10197) );
  OR U10458 ( .A(n10195), .B(n10194), .Z(n10196) );
  AND U10459 ( .A(n10197), .B(n10196), .Z(n10272) );
  XOR U10460 ( .A(n10273), .B(n10272), .Z(c[377]) );
  NANDN U10461 ( .A(n10199), .B(n10198), .Z(n10203) );
  NAND U10462 ( .A(n10201), .B(n10200), .Z(n10202) );
  NAND U10463 ( .A(n10203), .B(n10202), .Z(n10279) );
  NANDN U10464 ( .A(n10205), .B(n10204), .Z(n10209) );
  OR U10465 ( .A(n10207), .B(n10206), .Z(n10208) );
  NAND U10466 ( .A(n10209), .B(n10208), .Z(n10346) );
  XNOR U10467 ( .A(n20052), .B(n10525), .Z(n10288) );
  OR U10468 ( .A(n10288), .B(n20020), .Z(n10212) );
  NANDN U10469 ( .A(n10210), .B(n19960), .Z(n10211) );
  NAND U10470 ( .A(n10212), .B(n10211), .Z(n10301) );
  XNOR U10471 ( .A(n102), .B(n10213), .Z(n10292) );
  OR U10472 ( .A(n10292), .B(n20121), .Z(n10216) );
  NANDN U10473 ( .A(n10214), .B(n20122), .Z(n10215) );
  NAND U10474 ( .A(n10216), .B(n10215), .Z(n10298) );
  XNOR U10475 ( .A(n19975), .B(n10708), .Z(n10295) );
  NANDN U10476 ( .A(n10295), .B(n19883), .Z(n10219) );
  NANDN U10477 ( .A(n10217), .B(n19937), .Z(n10218) );
  AND U10478 ( .A(n10219), .B(n10218), .Z(n10299) );
  XNOR U10479 ( .A(n10298), .B(n10299), .Z(n10300) );
  XNOR U10480 ( .A(n10301), .B(n10300), .Z(n10337) );
  NANDN U10481 ( .A(n10221), .B(n10220), .Z(n10225) );
  NAND U10482 ( .A(n10223), .B(n10222), .Z(n10224) );
  NAND U10483 ( .A(n10225), .B(n10224), .Z(n10338) );
  XNOR U10484 ( .A(n10337), .B(n10338), .Z(n10339) );
  NANDN U10485 ( .A(n10227), .B(n10226), .Z(n10231) );
  NAND U10486 ( .A(n10229), .B(n10228), .Z(n10230) );
  AND U10487 ( .A(n10231), .B(n10230), .Z(n10340) );
  XNOR U10488 ( .A(n10339), .B(n10340), .Z(n10284) );
  NANDN U10489 ( .A(n10233), .B(n10232), .Z(n10237) );
  OR U10490 ( .A(n10235), .B(n10234), .Z(n10236) );
  NAND U10491 ( .A(n10237), .B(n10236), .Z(n10334) );
  NAND U10492 ( .A(b[0]), .B(a[138]), .Z(n10238) );
  XNOR U10493 ( .A(b[1]), .B(n10238), .Z(n10240) );
  NAND U10494 ( .A(a[137]), .B(n98), .Z(n10239) );
  AND U10495 ( .A(n10240), .B(n10239), .Z(n10310) );
  XNOR U10496 ( .A(n20154), .B(n10369), .Z(n10319) );
  OR U10497 ( .A(n10319), .B(n20057), .Z(n10243) );
  NANDN U10498 ( .A(n10241), .B(n20098), .Z(n10242) );
  AND U10499 ( .A(n10243), .B(n10242), .Z(n10311) );
  XOR U10500 ( .A(n10310), .B(n10311), .Z(n10313) );
  NAND U10501 ( .A(a[122]), .B(b[15]), .Z(n10312) );
  XOR U10502 ( .A(n10313), .B(n10312), .Z(n10331) );
  NAND U10503 ( .A(n19722), .B(n10244), .Z(n10246) );
  XNOR U10504 ( .A(b[5]), .B(n11020), .Z(n10322) );
  NANDN U10505 ( .A(n19640), .B(n10322), .Z(n10245) );
  NAND U10506 ( .A(n10246), .B(n10245), .Z(n10307) );
  XNOR U10507 ( .A(n19714), .B(n10837), .Z(n10325) );
  NANDN U10508 ( .A(n10325), .B(n19766), .Z(n10249) );
  NANDN U10509 ( .A(n10247), .B(n19767), .Z(n10248) );
  NAND U10510 ( .A(n10249), .B(n10248), .Z(n10304) );
  NAND U10511 ( .A(n19554), .B(n10250), .Z(n10252) );
  IV U10512 ( .A(a[136]), .Z(n11149) );
  XNOR U10513 ( .A(b[3]), .B(n11149), .Z(n10328) );
  NANDN U10514 ( .A(n19521), .B(n10328), .Z(n10251) );
  AND U10515 ( .A(n10252), .B(n10251), .Z(n10305) );
  XNOR U10516 ( .A(n10304), .B(n10305), .Z(n10306) );
  XOR U10517 ( .A(n10307), .B(n10306), .Z(n10332) );
  XOR U10518 ( .A(n10331), .B(n10332), .Z(n10333) );
  XNOR U10519 ( .A(n10334), .B(n10333), .Z(n10282) );
  NAND U10520 ( .A(n10254), .B(n10253), .Z(n10258) );
  NAND U10521 ( .A(n10256), .B(n10255), .Z(n10257) );
  NAND U10522 ( .A(n10258), .B(n10257), .Z(n10283) );
  XOR U10523 ( .A(n10282), .B(n10283), .Z(n10285) );
  XNOR U10524 ( .A(n10284), .B(n10285), .Z(n10343) );
  NANDN U10525 ( .A(n10260), .B(n10259), .Z(n10264) );
  NAND U10526 ( .A(n10262), .B(n10261), .Z(n10263) );
  NAND U10527 ( .A(n10264), .B(n10263), .Z(n10344) );
  XNOR U10528 ( .A(n10343), .B(n10344), .Z(n10345) );
  XOR U10529 ( .A(n10346), .B(n10345), .Z(n10276) );
  NANDN U10530 ( .A(n10266), .B(n10265), .Z(n10270) );
  NANDN U10531 ( .A(n10268), .B(n10267), .Z(n10269) );
  NAND U10532 ( .A(n10270), .B(n10269), .Z(n10277) );
  XNOR U10533 ( .A(n10276), .B(n10277), .Z(n10278) );
  XNOR U10534 ( .A(n10279), .B(n10278), .Z(n10349) );
  XNOR U10535 ( .A(n10349), .B(sreg[378]), .Z(n10351) );
  NAND U10536 ( .A(n10271), .B(sreg[377]), .Z(n10275) );
  OR U10537 ( .A(n10273), .B(n10272), .Z(n10274) );
  AND U10538 ( .A(n10275), .B(n10274), .Z(n10350) );
  XOR U10539 ( .A(n10351), .B(n10350), .Z(c[378]) );
  NANDN U10540 ( .A(n10277), .B(n10276), .Z(n10281) );
  NAND U10541 ( .A(n10279), .B(n10278), .Z(n10280) );
  NAND U10542 ( .A(n10281), .B(n10280), .Z(n10357) );
  NANDN U10543 ( .A(n10283), .B(n10282), .Z(n10287) );
  OR U10544 ( .A(n10285), .B(n10284), .Z(n10286) );
  NAND U10545 ( .A(n10287), .B(n10286), .Z(n10424) );
  XNOR U10546 ( .A(n20052), .B(n10630), .Z(n10366) );
  OR U10547 ( .A(n10366), .B(n20020), .Z(n10290) );
  NANDN U10548 ( .A(n10288), .B(n19960), .Z(n10289) );
  NAND U10549 ( .A(n10290), .B(n10289), .Z(n10379) );
  XNOR U10550 ( .A(n102), .B(n10291), .Z(n10370) );
  OR U10551 ( .A(n10370), .B(n20121), .Z(n10294) );
  NANDN U10552 ( .A(n10292), .B(n20122), .Z(n10293) );
  NAND U10553 ( .A(n10294), .B(n10293), .Z(n10376) );
  XNOR U10554 ( .A(n19975), .B(n10786), .Z(n10373) );
  NANDN U10555 ( .A(n10373), .B(n19883), .Z(n10297) );
  NANDN U10556 ( .A(n10295), .B(n19937), .Z(n10296) );
  AND U10557 ( .A(n10297), .B(n10296), .Z(n10377) );
  XNOR U10558 ( .A(n10376), .B(n10377), .Z(n10378) );
  XNOR U10559 ( .A(n10379), .B(n10378), .Z(n10415) );
  NANDN U10560 ( .A(n10299), .B(n10298), .Z(n10303) );
  NAND U10561 ( .A(n10301), .B(n10300), .Z(n10302) );
  NAND U10562 ( .A(n10303), .B(n10302), .Z(n10416) );
  XNOR U10563 ( .A(n10415), .B(n10416), .Z(n10417) );
  NANDN U10564 ( .A(n10305), .B(n10304), .Z(n10309) );
  NAND U10565 ( .A(n10307), .B(n10306), .Z(n10308) );
  AND U10566 ( .A(n10309), .B(n10308), .Z(n10418) );
  XNOR U10567 ( .A(n10417), .B(n10418), .Z(n10362) );
  NANDN U10568 ( .A(n10311), .B(n10310), .Z(n10315) );
  OR U10569 ( .A(n10313), .B(n10312), .Z(n10314) );
  NAND U10570 ( .A(n10315), .B(n10314), .Z(n10412) );
  NAND U10571 ( .A(b[0]), .B(a[139]), .Z(n10316) );
  XNOR U10572 ( .A(b[1]), .B(n10316), .Z(n10318) );
  NAND U10573 ( .A(a[138]), .B(n98), .Z(n10317) );
  AND U10574 ( .A(n10318), .B(n10317), .Z(n10388) );
  XNOR U10575 ( .A(n20154), .B(n10474), .Z(n10397) );
  OR U10576 ( .A(n10397), .B(n20057), .Z(n10321) );
  NANDN U10577 ( .A(n10319), .B(n20098), .Z(n10320) );
  AND U10578 ( .A(n10321), .B(n10320), .Z(n10389) );
  XOR U10579 ( .A(n10388), .B(n10389), .Z(n10391) );
  NAND U10580 ( .A(a[123]), .B(b[15]), .Z(n10390) );
  XOR U10581 ( .A(n10391), .B(n10390), .Z(n10409) );
  NAND U10582 ( .A(n19722), .B(n10322), .Z(n10324) );
  XNOR U10583 ( .A(b[5]), .B(n11098), .Z(n10400) );
  NANDN U10584 ( .A(n19640), .B(n10400), .Z(n10323) );
  NAND U10585 ( .A(n10324), .B(n10323), .Z(n10385) );
  XNOR U10586 ( .A(n19714), .B(n10942), .Z(n10403) );
  NANDN U10587 ( .A(n10403), .B(n19766), .Z(n10327) );
  NANDN U10588 ( .A(n10325), .B(n19767), .Z(n10326) );
  NAND U10589 ( .A(n10327), .B(n10326), .Z(n10382) );
  NAND U10590 ( .A(n19554), .B(n10328), .Z(n10330) );
  IV U10591 ( .A(a[137]), .Z(n11254) );
  XNOR U10592 ( .A(b[3]), .B(n11254), .Z(n10406) );
  NANDN U10593 ( .A(n19521), .B(n10406), .Z(n10329) );
  AND U10594 ( .A(n10330), .B(n10329), .Z(n10383) );
  XNOR U10595 ( .A(n10382), .B(n10383), .Z(n10384) );
  XOR U10596 ( .A(n10385), .B(n10384), .Z(n10410) );
  XOR U10597 ( .A(n10409), .B(n10410), .Z(n10411) );
  XNOR U10598 ( .A(n10412), .B(n10411), .Z(n10360) );
  NAND U10599 ( .A(n10332), .B(n10331), .Z(n10336) );
  NAND U10600 ( .A(n10334), .B(n10333), .Z(n10335) );
  NAND U10601 ( .A(n10336), .B(n10335), .Z(n10361) );
  XOR U10602 ( .A(n10360), .B(n10361), .Z(n10363) );
  XNOR U10603 ( .A(n10362), .B(n10363), .Z(n10421) );
  NANDN U10604 ( .A(n10338), .B(n10337), .Z(n10342) );
  NAND U10605 ( .A(n10340), .B(n10339), .Z(n10341) );
  NAND U10606 ( .A(n10342), .B(n10341), .Z(n10422) );
  XNOR U10607 ( .A(n10421), .B(n10422), .Z(n10423) );
  XOR U10608 ( .A(n10424), .B(n10423), .Z(n10354) );
  NANDN U10609 ( .A(n10344), .B(n10343), .Z(n10348) );
  NANDN U10610 ( .A(n10346), .B(n10345), .Z(n10347) );
  NAND U10611 ( .A(n10348), .B(n10347), .Z(n10355) );
  XNOR U10612 ( .A(n10354), .B(n10355), .Z(n10356) );
  XNOR U10613 ( .A(n10357), .B(n10356), .Z(n10427) );
  XNOR U10614 ( .A(n10427), .B(sreg[379]), .Z(n10429) );
  NAND U10615 ( .A(n10349), .B(sreg[378]), .Z(n10353) );
  OR U10616 ( .A(n10351), .B(n10350), .Z(n10352) );
  AND U10617 ( .A(n10353), .B(n10352), .Z(n10428) );
  XOR U10618 ( .A(n10429), .B(n10428), .Z(c[379]) );
  NANDN U10619 ( .A(n10355), .B(n10354), .Z(n10359) );
  NAND U10620 ( .A(n10357), .B(n10356), .Z(n10358) );
  NAND U10621 ( .A(n10359), .B(n10358), .Z(n10435) );
  NANDN U10622 ( .A(n10361), .B(n10360), .Z(n10365) );
  OR U10623 ( .A(n10363), .B(n10362), .Z(n10364) );
  NAND U10624 ( .A(n10365), .B(n10364), .Z(n10502) );
  XNOR U10625 ( .A(n20052), .B(n10708), .Z(n10471) );
  OR U10626 ( .A(n10471), .B(n20020), .Z(n10368) );
  NANDN U10627 ( .A(n10366), .B(n19960), .Z(n10367) );
  NAND U10628 ( .A(n10368), .B(n10367), .Z(n10484) );
  XNOR U10629 ( .A(n102), .B(n10369), .Z(n10475) );
  OR U10630 ( .A(n10475), .B(n20121), .Z(n10372) );
  NANDN U10631 ( .A(n10370), .B(n20122), .Z(n10371) );
  NAND U10632 ( .A(n10372), .B(n10371), .Z(n10481) );
  XNOR U10633 ( .A(n19975), .B(n10837), .Z(n10478) );
  NANDN U10634 ( .A(n10478), .B(n19883), .Z(n10375) );
  NANDN U10635 ( .A(n10373), .B(n19937), .Z(n10374) );
  AND U10636 ( .A(n10375), .B(n10374), .Z(n10482) );
  XNOR U10637 ( .A(n10481), .B(n10482), .Z(n10483) );
  XNOR U10638 ( .A(n10484), .B(n10483), .Z(n10493) );
  NANDN U10639 ( .A(n10377), .B(n10376), .Z(n10381) );
  NAND U10640 ( .A(n10379), .B(n10378), .Z(n10380) );
  NAND U10641 ( .A(n10381), .B(n10380), .Z(n10494) );
  XNOR U10642 ( .A(n10493), .B(n10494), .Z(n10495) );
  NANDN U10643 ( .A(n10383), .B(n10382), .Z(n10387) );
  NAND U10644 ( .A(n10385), .B(n10384), .Z(n10386) );
  AND U10645 ( .A(n10387), .B(n10386), .Z(n10496) );
  XNOR U10646 ( .A(n10495), .B(n10496), .Z(n10440) );
  NANDN U10647 ( .A(n10389), .B(n10388), .Z(n10393) );
  OR U10648 ( .A(n10391), .B(n10390), .Z(n10392) );
  NAND U10649 ( .A(n10393), .B(n10392), .Z(n10468) );
  NAND U10650 ( .A(b[0]), .B(a[140]), .Z(n10394) );
  XNOR U10651 ( .A(b[1]), .B(n10394), .Z(n10396) );
  NAND U10652 ( .A(a[139]), .B(n98), .Z(n10395) );
  AND U10653 ( .A(n10396), .B(n10395), .Z(n10444) );
  XNOR U10654 ( .A(n20154), .B(n10525), .Z(n10453) );
  OR U10655 ( .A(n10453), .B(n20057), .Z(n10399) );
  NANDN U10656 ( .A(n10397), .B(n20098), .Z(n10398) );
  AND U10657 ( .A(n10399), .B(n10398), .Z(n10445) );
  XOR U10658 ( .A(n10444), .B(n10445), .Z(n10447) );
  NAND U10659 ( .A(a[124]), .B(b[15]), .Z(n10446) );
  XOR U10660 ( .A(n10447), .B(n10446), .Z(n10465) );
  NAND U10661 ( .A(n19722), .B(n10400), .Z(n10402) );
  XNOR U10662 ( .A(b[5]), .B(n11149), .Z(n10456) );
  NANDN U10663 ( .A(n19640), .B(n10456), .Z(n10401) );
  NAND U10664 ( .A(n10402), .B(n10401), .Z(n10490) );
  XNOR U10665 ( .A(n19714), .B(n11020), .Z(n10459) );
  NANDN U10666 ( .A(n10459), .B(n19766), .Z(n10405) );
  NANDN U10667 ( .A(n10403), .B(n19767), .Z(n10404) );
  NAND U10668 ( .A(n10405), .B(n10404), .Z(n10487) );
  NAND U10669 ( .A(n19554), .B(n10406), .Z(n10408) );
  IV U10670 ( .A(a[138]), .Z(n11305) );
  XNOR U10671 ( .A(b[3]), .B(n11305), .Z(n10462) );
  NANDN U10672 ( .A(n19521), .B(n10462), .Z(n10407) );
  AND U10673 ( .A(n10408), .B(n10407), .Z(n10488) );
  XNOR U10674 ( .A(n10487), .B(n10488), .Z(n10489) );
  XOR U10675 ( .A(n10490), .B(n10489), .Z(n10466) );
  XOR U10676 ( .A(n10465), .B(n10466), .Z(n10467) );
  XNOR U10677 ( .A(n10468), .B(n10467), .Z(n10438) );
  NAND U10678 ( .A(n10410), .B(n10409), .Z(n10414) );
  NAND U10679 ( .A(n10412), .B(n10411), .Z(n10413) );
  NAND U10680 ( .A(n10414), .B(n10413), .Z(n10439) );
  XOR U10681 ( .A(n10438), .B(n10439), .Z(n10441) );
  XNOR U10682 ( .A(n10440), .B(n10441), .Z(n10499) );
  NANDN U10683 ( .A(n10416), .B(n10415), .Z(n10420) );
  NAND U10684 ( .A(n10418), .B(n10417), .Z(n10419) );
  NAND U10685 ( .A(n10420), .B(n10419), .Z(n10500) );
  XNOR U10686 ( .A(n10499), .B(n10500), .Z(n10501) );
  XOR U10687 ( .A(n10502), .B(n10501), .Z(n10432) );
  NANDN U10688 ( .A(n10422), .B(n10421), .Z(n10426) );
  NANDN U10689 ( .A(n10424), .B(n10423), .Z(n10425) );
  NAND U10690 ( .A(n10426), .B(n10425), .Z(n10433) );
  XNOR U10691 ( .A(n10432), .B(n10433), .Z(n10434) );
  XNOR U10692 ( .A(n10435), .B(n10434), .Z(n10505) );
  XNOR U10693 ( .A(n10505), .B(sreg[380]), .Z(n10507) );
  NAND U10694 ( .A(n10427), .B(sreg[379]), .Z(n10431) );
  OR U10695 ( .A(n10429), .B(n10428), .Z(n10430) );
  AND U10696 ( .A(n10431), .B(n10430), .Z(n10506) );
  XOR U10697 ( .A(n10507), .B(n10506), .Z(c[380]) );
  NANDN U10698 ( .A(n10433), .B(n10432), .Z(n10437) );
  NAND U10699 ( .A(n10435), .B(n10434), .Z(n10436) );
  NAND U10700 ( .A(n10437), .B(n10436), .Z(n10513) );
  NANDN U10701 ( .A(n10439), .B(n10438), .Z(n10443) );
  OR U10702 ( .A(n10441), .B(n10440), .Z(n10442) );
  NAND U10703 ( .A(n10443), .B(n10442), .Z(n10580) );
  NANDN U10704 ( .A(n10445), .B(n10444), .Z(n10449) );
  OR U10705 ( .A(n10447), .B(n10446), .Z(n10448) );
  NAND U10706 ( .A(n10449), .B(n10448), .Z(n10568) );
  NAND U10707 ( .A(b[0]), .B(a[141]), .Z(n10450) );
  XNOR U10708 ( .A(b[1]), .B(n10450), .Z(n10452) );
  NAND U10709 ( .A(a[140]), .B(n98), .Z(n10451) );
  AND U10710 ( .A(n10452), .B(n10451), .Z(n10544) );
  XNOR U10711 ( .A(n20154), .B(n10630), .Z(n10553) );
  OR U10712 ( .A(n10553), .B(n20057), .Z(n10455) );
  NANDN U10713 ( .A(n10453), .B(n20098), .Z(n10454) );
  AND U10714 ( .A(n10455), .B(n10454), .Z(n10545) );
  XOR U10715 ( .A(n10544), .B(n10545), .Z(n10547) );
  NAND U10716 ( .A(a[125]), .B(b[15]), .Z(n10546) );
  XOR U10717 ( .A(n10547), .B(n10546), .Z(n10565) );
  NAND U10718 ( .A(n19722), .B(n10456), .Z(n10458) );
  XNOR U10719 ( .A(b[5]), .B(n11254), .Z(n10556) );
  NANDN U10720 ( .A(n19640), .B(n10556), .Z(n10457) );
  NAND U10721 ( .A(n10458), .B(n10457), .Z(n10541) );
  XNOR U10722 ( .A(n19714), .B(n11098), .Z(n10559) );
  NANDN U10723 ( .A(n10559), .B(n19766), .Z(n10461) );
  NANDN U10724 ( .A(n10459), .B(n19767), .Z(n10460) );
  NAND U10725 ( .A(n10461), .B(n10460), .Z(n10538) );
  NAND U10726 ( .A(n19554), .B(n10462), .Z(n10464) );
  IV U10727 ( .A(a[139]), .Z(n11410) );
  XNOR U10728 ( .A(b[3]), .B(n11410), .Z(n10562) );
  NANDN U10729 ( .A(n19521), .B(n10562), .Z(n10463) );
  AND U10730 ( .A(n10464), .B(n10463), .Z(n10539) );
  XNOR U10731 ( .A(n10538), .B(n10539), .Z(n10540) );
  XOR U10732 ( .A(n10541), .B(n10540), .Z(n10566) );
  XOR U10733 ( .A(n10565), .B(n10566), .Z(n10567) );
  XNOR U10734 ( .A(n10568), .B(n10567), .Z(n10516) );
  NAND U10735 ( .A(n10466), .B(n10465), .Z(n10470) );
  NAND U10736 ( .A(n10468), .B(n10467), .Z(n10469) );
  NAND U10737 ( .A(n10470), .B(n10469), .Z(n10517) );
  XOR U10738 ( .A(n10516), .B(n10517), .Z(n10519) );
  XNOR U10739 ( .A(n20052), .B(n10786), .Z(n10522) );
  OR U10740 ( .A(n10522), .B(n20020), .Z(n10473) );
  NANDN U10741 ( .A(n10471), .B(n19960), .Z(n10472) );
  NAND U10742 ( .A(n10473), .B(n10472), .Z(n10535) );
  XNOR U10743 ( .A(n102), .B(n10474), .Z(n10526) );
  OR U10744 ( .A(n10526), .B(n20121), .Z(n10477) );
  NANDN U10745 ( .A(n10475), .B(n20122), .Z(n10476) );
  NAND U10746 ( .A(n10477), .B(n10476), .Z(n10532) );
  XNOR U10747 ( .A(n19975), .B(n10942), .Z(n10529) );
  NANDN U10748 ( .A(n10529), .B(n19883), .Z(n10480) );
  NANDN U10749 ( .A(n10478), .B(n19937), .Z(n10479) );
  AND U10750 ( .A(n10480), .B(n10479), .Z(n10533) );
  XNOR U10751 ( .A(n10532), .B(n10533), .Z(n10534) );
  XNOR U10752 ( .A(n10535), .B(n10534), .Z(n10571) );
  NANDN U10753 ( .A(n10482), .B(n10481), .Z(n10486) );
  NAND U10754 ( .A(n10484), .B(n10483), .Z(n10485) );
  NAND U10755 ( .A(n10486), .B(n10485), .Z(n10572) );
  XNOR U10756 ( .A(n10571), .B(n10572), .Z(n10573) );
  NANDN U10757 ( .A(n10488), .B(n10487), .Z(n10492) );
  NAND U10758 ( .A(n10490), .B(n10489), .Z(n10491) );
  AND U10759 ( .A(n10492), .B(n10491), .Z(n10574) );
  XNOR U10760 ( .A(n10573), .B(n10574), .Z(n10518) );
  XNOR U10761 ( .A(n10519), .B(n10518), .Z(n10577) );
  NANDN U10762 ( .A(n10494), .B(n10493), .Z(n10498) );
  NAND U10763 ( .A(n10496), .B(n10495), .Z(n10497) );
  NAND U10764 ( .A(n10498), .B(n10497), .Z(n10578) );
  XNOR U10765 ( .A(n10577), .B(n10578), .Z(n10579) );
  XOR U10766 ( .A(n10580), .B(n10579), .Z(n10510) );
  NANDN U10767 ( .A(n10500), .B(n10499), .Z(n10504) );
  NANDN U10768 ( .A(n10502), .B(n10501), .Z(n10503) );
  NAND U10769 ( .A(n10504), .B(n10503), .Z(n10511) );
  XNOR U10770 ( .A(n10510), .B(n10511), .Z(n10512) );
  XNOR U10771 ( .A(n10513), .B(n10512), .Z(n10583) );
  XNOR U10772 ( .A(n10583), .B(sreg[381]), .Z(n10585) );
  NAND U10773 ( .A(n10505), .B(sreg[380]), .Z(n10509) );
  OR U10774 ( .A(n10507), .B(n10506), .Z(n10508) );
  AND U10775 ( .A(n10509), .B(n10508), .Z(n10584) );
  XOR U10776 ( .A(n10585), .B(n10584), .Z(c[381]) );
  NANDN U10777 ( .A(n10511), .B(n10510), .Z(n10515) );
  NAND U10778 ( .A(n10513), .B(n10512), .Z(n10514) );
  NAND U10779 ( .A(n10515), .B(n10514), .Z(n10591) );
  NANDN U10780 ( .A(n10517), .B(n10516), .Z(n10521) );
  OR U10781 ( .A(n10519), .B(n10518), .Z(n10520) );
  NAND U10782 ( .A(n10521), .B(n10520), .Z(n10658) );
  XNOR U10783 ( .A(n20052), .B(n10837), .Z(n10627) );
  OR U10784 ( .A(n10627), .B(n20020), .Z(n10524) );
  NANDN U10785 ( .A(n10522), .B(n19960), .Z(n10523) );
  NAND U10786 ( .A(n10524), .B(n10523), .Z(n10640) );
  XNOR U10787 ( .A(n102), .B(n10525), .Z(n10631) );
  OR U10788 ( .A(n10631), .B(n20121), .Z(n10528) );
  NANDN U10789 ( .A(n10526), .B(n20122), .Z(n10527) );
  NAND U10790 ( .A(n10528), .B(n10527), .Z(n10637) );
  XNOR U10791 ( .A(n19975), .B(n11020), .Z(n10634) );
  NANDN U10792 ( .A(n10634), .B(n19883), .Z(n10531) );
  NANDN U10793 ( .A(n10529), .B(n19937), .Z(n10530) );
  AND U10794 ( .A(n10531), .B(n10530), .Z(n10638) );
  XNOR U10795 ( .A(n10637), .B(n10638), .Z(n10639) );
  XNOR U10796 ( .A(n10640), .B(n10639), .Z(n10649) );
  NANDN U10797 ( .A(n10533), .B(n10532), .Z(n10537) );
  NAND U10798 ( .A(n10535), .B(n10534), .Z(n10536) );
  NAND U10799 ( .A(n10537), .B(n10536), .Z(n10650) );
  XNOR U10800 ( .A(n10649), .B(n10650), .Z(n10651) );
  NANDN U10801 ( .A(n10539), .B(n10538), .Z(n10543) );
  NAND U10802 ( .A(n10541), .B(n10540), .Z(n10542) );
  AND U10803 ( .A(n10543), .B(n10542), .Z(n10652) );
  XNOR U10804 ( .A(n10651), .B(n10652), .Z(n10596) );
  NANDN U10805 ( .A(n10545), .B(n10544), .Z(n10549) );
  OR U10806 ( .A(n10547), .B(n10546), .Z(n10548) );
  NAND U10807 ( .A(n10549), .B(n10548), .Z(n10624) );
  NAND U10808 ( .A(b[0]), .B(a[142]), .Z(n10550) );
  XNOR U10809 ( .A(b[1]), .B(n10550), .Z(n10552) );
  NAND U10810 ( .A(a[141]), .B(n98), .Z(n10551) );
  AND U10811 ( .A(n10552), .B(n10551), .Z(n10600) );
  XNOR U10812 ( .A(n20154), .B(n10708), .Z(n10609) );
  OR U10813 ( .A(n10609), .B(n20057), .Z(n10555) );
  NANDN U10814 ( .A(n10553), .B(n20098), .Z(n10554) );
  AND U10815 ( .A(n10555), .B(n10554), .Z(n10601) );
  XOR U10816 ( .A(n10600), .B(n10601), .Z(n10603) );
  NAND U10817 ( .A(a[126]), .B(b[15]), .Z(n10602) );
  XOR U10818 ( .A(n10603), .B(n10602), .Z(n10621) );
  NAND U10819 ( .A(n19722), .B(n10556), .Z(n10558) );
  XNOR U10820 ( .A(b[5]), .B(n11305), .Z(n10612) );
  NANDN U10821 ( .A(n19640), .B(n10612), .Z(n10557) );
  NAND U10822 ( .A(n10558), .B(n10557), .Z(n10646) );
  XNOR U10823 ( .A(n19714), .B(n11149), .Z(n10615) );
  NANDN U10824 ( .A(n10615), .B(n19766), .Z(n10561) );
  NANDN U10825 ( .A(n10559), .B(n19767), .Z(n10560) );
  NAND U10826 ( .A(n10561), .B(n10560), .Z(n10643) );
  NAND U10827 ( .A(n19554), .B(n10562), .Z(n10564) );
  IV U10828 ( .A(a[140]), .Z(n11461) );
  XNOR U10829 ( .A(b[3]), .B(n11461), .Z(n10618) );
  NANDN U10830 ( .A(n19521), .B(n10618), .Z(n10563) );
  AND U10831 ( .A(n10564), .B(n10563), .Z(n10644) );
  XNOR U10832 ( .A(n10643), .B(n10644), .Z(n10645) );
  XOR U10833 ( .A(n10646), .B(n10645), .Z(n10622) );
  XOR U10834 ( .A(n10621), .B(n10622), .Z(n10623) );
  XNOR U10835 ( .A(n10624), .B(n10623), .Z(n10594) );
  NAND U10836 ( .A(n10566), .B(n10565), .Z(n10570) );
  NAND U10837 ( .A(n10568), .B(n10567), .Z(n10569) );
  NAND U10838 ( .A(n10570), .B(n10569), .Z(n10595) );
  XOR U10839 ( .A(n10594), .B(n10595), .Z(n10597) );
  XNOR U10840 ( .A(n10596), .B(n10597), .Z(n10655) );
  NANDN U10841 ( .A(n10572), .B(n10571), .Z(n10576) );
  NAND U10842 ( .A(n10574), .B(n10573), .Z(n10575) );
  NAND U10843 ( .A(n10576), .B(n10575), .Z(n10656) );
  XNOR U10844 ( .A(n10655), .B(n10656), .Z(n10657) );
  XOR U10845 ( .A(n10658), .B(n10657), .Z(n10588) );
  NANDN U10846 ( .A(n10578), .B(n10577), .Z(n10582) );
  NANDN U10847 ( .A(n10580), .B(n10579), .Z(n10581) );
  NAND U10848 ( .A(n10582), .B(n10581), .Z(n10589) );
  XNOR U10849 ( .A(n10588), .B(n10589), .Z(n10590) );
  XNOR U10850 ( .A(n10591), .B(n10590), .Z(n10661) );
  XNOR U10851 ( .A(n10661), .B(sreg[382]), .Z(n10663) );
  NAND U10852 ( .A(n10583), .B(sreg[381]), .Z(n10587) );
  OR U10853 ( .A(n10585), .B(n10584), .Z(n10586) );
  AND U10854 ( .A(n10587), .B(n10586), .Z(n10662) );
  XOR U10855 ( .A(n10663), .B(n10662), .Z(c[382]) );
  NANDN U10856 ( .A(n10589), .B(n10588), .Z(n10593) );
  NAND U10857 ( .A(n10591), .B(n10590), .Z(n10592) );
  NAND U10858 ( .A(n10593), .B(n10592), .Z(n10669) );
  NANDN U10859 ( .A(n10595), .B(n10594), .Z(n10599) );
  OR U10860 ( .A(n10597), .B(n10596), .Z(n10598) );
  NAND U10861 ( .A(n10599), .B(n10598), .Z(n10736) );
  NANDN U10862 ( .A(n10601), .B(n10600), .Z(n10605) );
  OR U10863 ( .A(n10603), .B(n10602), .Z(n10604) );
  NAND U10864 ( .A(n10605), .B(n10604), .Z(n10702) );
  NAND U10865 ( .A(b[0]), .B(a[143]), .Z(n10606) );
  XNOR U10866 ( .A(b[1]), .B(n10606), .Z(n10608) );
  NAND U10867 ( .A(a[142]), .B(n98), .Z(n10607) );
  AND U10868 ( .A(n10608), .B(n10607), .Z(n10678) );
  XNOR U10869 ( .A(n20154), .B(n10786), .Z(n10687) );
  OR U10870 ( .A(n10687), .B(n20057), .Z(n10611) );
  NANDN U10871 ( .A(n10609), .B(n20098), .Z(n10610) );
  AND U10872 ( .A(n10611), .B(n10610), .Z(n10679) );
  XOR U10873 ( .A(n10678), .B(n10679), .Z(n10681) );
  NAND U10874 ( .A(a[127]), .B(b[15]), .Z(n10680) );
  XOR U10875 ( .A(n10681), .B(n10680), .Z(n10699) );
  NAND U10876 ( .A(n19722), .B(n10612), .Z(n10614) );
  XNOR U10877 ( .A(b[5]), .B(n11410), .Z(n10690) );
  NANDN U10878 ( .A(n19640), .B(n10690), .Z(n10613) );
  NAND U10879 ( .A(n10614), .B(n10613), .Z(n10724) );
  XNOR U10880 ( .A(n19714), .B(n11254), .Z(n10693) );
  NANDN U10881 ( .A(n10693), .B(n19766), .Z(n10617) );
  NANDN U10882 ( .A(n10615), .B(n19767), .Z(n10616) );
  NAND U10883 ( .A(n10617), .B(n10616), .Z(n10721) );
  NAND U10884 ( .A(n19554), .B(n10618), .Z(n10620) );
  IV U10885 ( .A(a[141]), .Z(n11539) );
  XNOR U10886 ( .A(b[3]), .B(n11539), .Z(n10696) );
  NANDN U10887 ( .A(n19521), .B(n10696), .Z(n10619) );
  AND U10888 ( .A(n10620), .B(n10619), .Z(n10722) );
  XNOR U10889 ( .A(n10721), .B(n10722), .Z(n10723) );
  XOR U10890 ( .A(n10724), .B(n10723), .Z(n10700) );
  XOR U10891 ( .A(n10699), .B(n10700), .Z(n10701) );
  XNOR U10892 ( .A(n10702), .B(n10701), .Z(n10672) );
  NAND U10893 ( .A(n10622), .B(n10621), .Z(n10626) );
  NAND U10894 ( .A(n10624), .B(n10623), .Z(n10625) );
  NAND U10895 ( .A(n10626), .B(n10625), .Z(n10673) );
  XOR U10896 ( .A(n10672), .B(n10673), .Z(n10675) );
  XNOR U10897 ( .A(n20052), .B(n10942), .Z(n10705) );
  OR U10898 ( .A(n10705), .B(n20020), .Z(n10629) );
  NANDN U10899 ( .A(n10627), .B(n19960), .Z(n10628) );
  NAND U10900 ( .A(n10629), .B(n10628), .Z(n10718) );
  XNOR U10901 ( .A(n102), .B(n10630), .Z(n10709) );
  OR U10902 ( .A(n10709), .B(n20121), .Z(n10633) );
  NANDN U10903 ( .A(n10631), .B(n20122), .Z(n10632) );
  NAND U10904 ( .A(n10633), .B(n10632), .Z(n10715) );
  XNOR U10905 ( .A(n19975), .B(n11098), .Z(n10712) );
  NANDN U10906 ( .A(n10712), .B(n19883), .Z(n10636) );
  NANDN U10907 ( .A(n10634), .B(n19937), .Z(n10635) );
  AND U10908 ( .A(n10636), .B(n10635), .Z(n10716) );
  XNOR U10909 ( .A(n10715), .B(n10716), .Z(n10717) );
  XNOR U10910 ( .A(n10718), .B(n10717), .Z(n10727) );
  NANDN U10911 ( .A(n10638), .B(n10637), .Z(n10642) );
  NAND U10912 ( .A(n10640), .B(n10639), .Z(n10641) );
  NAND U10913 ( .A(n10642), .B(n10641), .Z(n10728) );
  XNOR U10914 ( .A(n10727), .B(n10728), .Z(n10729) );
  NANDN U10915 ( .A(n10644), .B(n10643), .Z(n10648) );
  NAND U10916 ( .A(n10646), .B(n10645), .Z(n10647) );
  AND U10917 ( .A(n10648), .B(n10647), .Z(n10730) );
  XNOR U10918 ( .A(n10729), .B(n10730), .Z(n10674) );
  XNOR U10919 ( .A(n10675), .B(n10674), .Z(n10733) );
  NANDN U10920 ( .A(n10650), .B(n10649), .Z(n10654) );
  NAND U10921 ( .A(n10652), .B(n10651), .Z(n10653) );
  NAND U10922 ( .A(n10654), .B(n10653), .Z(n10734) );
  XNOR U10923 ( .A(n10733), .B(n10734), .Z(n10735) );
  XOR U10924 ( .A(n10736), .B(n10735), .Z(n10666) );
  NANDN U10925 ( .A(n10656), .B(n10655), .Z(n10660) );
  NANDN U10926 ( .A(n10658), .B(n10657), .Z(n10659) );
  NAND U10927 ( .A(n10660), .B(n10659), .Z(n10667) );
  XNOR U10928 ( .A(n10666), .B(n10667), .Z(n10668) );
  XNOR U10929 ( .A(n10669), .B(n10668), .Z(n10739) );
  XNOR U10930 ( .A(n10739), .B(sreg[383]), .Z(n10741) );
  NAND U10931 ( .A(n10661), .B(sreg[382]), .Z(n10665) );
  OR U10932 ( .A(n10663), .B(n10662), .Z(n10664) );
  AND U10933 ( .A(n10665), .B(n10664), .Z(n10740) );
  XOR U10934 ( .A(n10741), .B(n10740), .Z(c[383]) );
  NANDN U10935 ( .A(n10667), .B(n10666), .Z(n10671) );
  NAND U10936 ( .A(n10669), .B(n10668), .Z(n10670) );
  NAND U10937 ( .A(n10671), .B(n10670), .Z(n10747) );
  NANDN U10938 ( .A(n10673), .B(n10672), .Z(n10677) );
  OR U10939 ( .A(n10675), .B(n10674), .Z(n10676) );
  NAND U10940 ( .A(n10677), .B(n10676), .Z(n10814) );
  NANDN U10941 ( .A(n10679), .B(n10678), .Z(n10683) );
  OR U10942 ( .A(n10681), .B(n10680), .Z(n10682) );
  NAND U10943 ( .A(n10683), .B(n10682), .Z(n10780) );
  NAND U10944 ( .A(b[0]), .B(a[144]), .Z(n10684) );
  XNOR U10945 ( .A(b[1]), .B(n10684), .Z(n10686) );
  NAND U10946 ( .A(a[143]), .B(n98), .Z(n10685) );
  AND U10947 ( .A(n10686), .B(n10685), .Z(n10756) );
  XNOR U10948 ( .A(n20154), .B(n10837), .Z(n10765) );
  OR U10949 ( .A(n10765), .B(n20057), .Z(n10689) );
  NANDN U10950 ( .A(n10687), .B(n20098), .Z(n10688) );
  AND U10951 ( .A(n10689), .B(n10688), .Z(n10757) );
  XOR U10952 ( .A(n10756), .B(n10757), .Z(n10759) );
  NAND U10953 ( .A(a[128]), .B(b[15]), .Z(n10758) );
  XOR U10954 ( .A(n10759), .B(n10758), .Z(n10777) );
  NAND U10955 ( .A(n19722), .B(n10690), .Z(n10692) );
  XNOR U10956 ( .A(b[5]), .B(n11461), .Z(n10768) );
  NANDN U10957 ( .A(n19640), .B(n10768), .Z(n10691) );
  NAND U10958 ( .A(n10692), .B(n10691), .Z(n10802) );
  XNOR U10959 ( .A(n19714), .B(n11305), .Z(n10771) );
  NANDN U10960 ( .A(n10771), .B(n19766), .Z(n10695) );
  NANDN U10961 ( .A(n10693), .B(n19767), .Z(n10694) );
  NAND U10962 ( .A(n10695), .B(n10694), .Z(n10799) );
  NAND U10963 ( .A(n19554), .B(n10696), .Z(n10698) );
  IV U10964 ( .A(a[142]), .Z(n11644) );
  XNOR U10965 ( .A(b[3]), .B(n11644), .Z(n10774) );
  NANDN U10966 ( .A(n19521), .B(n10774), .Z(n10697) );
  AND U10967 ( .A(n10698), .B(n10697), .Z(n10800) );
  XNOR U10968 ( .A(n10799), .B(n10800), .Z(n10801) );
  XOR U10969 ( .A(n10802), .B(n10801), .Z(n10778) );
  XOR U10970 ( .A(n10777), .B(n10778), .Z(n10779) );
  XNOR U10971 ( .A(n10780), .B(n10779), .Z(n10750) );
  NAND U10972 ( .A(n10700), .B(n10699), .Z(n10704) );
  NAND U10973 ( .A(n10702), .B(n10701), .Z(n10703) );
  NAND U10974 ( .A(n10704), .B(n10703), .Z(n10751) );
  XOR U10975 ( .A(n10750), .B(n10751), .Z(n10753) );
  XNOR U10976 ( .A(n20052), .B(n11020), .Z(n10783) );
  OR U10977 ( .A(n10783), .B(n20020), .Z(n10707) );
  NANDN U10978 ( .A(n10705), .B(n19960), .Z(n10706) );
  NAND U10979 ( .A(n10707), .B(n10706), .Z(n10796) );
  XNOR U10980 ( .A(n102), .B(n10708), .Z(n10787) );
  OR U10981 ( .A(n10787), .B(n20121), .Z(n10711) );
  NANDN U10982 ( .A(n10709), .B(n20122), .Z(n10710) );
  NAND U10983 ( .A(n10711), .B(n10710), .Z(n10793) );
  XNOR U10984 ( .A(n19975), .B(n11149), .Z(n10790) );
  NANDN U10985 ( .A(n10790), .B(n19883), .Z(n10714) );
  NANDN U10986 ( .A(n10712), .B(n19937), .Z(n10713) );
  AND U10987 ( .A(n10714), .B(n10713), .Z(n10794) );
  XNOR U10988 ( .A(n10793), .B(n10794), .Z(n10795) );
  XNOR U10989 ( .A(n10796), .B(n10795), .Z(n10805) );
  NANDN U10990 ( .A(n10716), .B(n10715), .Z(n10720) );
  NAND U10991 ( .A(n10718), .B(n10717), .Z(n10719) );
  NAND U10992 ( .A(n10720), .B(n10719), .Z(n10806) );
  XNOR U10993 ( .A(n10805), .B(n10806), .Z(n10807) );
  NANDN U10994 ( .A(n10722), .B(n10721), .Z(n10726) );
  NAND U10995 ( .A(n10724), .B(n10723), .Z(n10725) );
  AND U10996 ( .A(n10726), .B(n10725), .Z(n10808) );
  XNOR U10997 ( .A(n10807), .B(n10808), .Z(n10752) );
  XNOR U10998 ( .A(n10753), .B(n10752), .Z(n10811) );
  NANDN U10999 ( .A(n10728), .B(n10727), .Z(n10732) );
  NAND U11000 ( .A(n10730), .B(n10729), .Z(n10731) );
  NAND U11001 ( .A(n10732), .B(n10731), .Z(n10812) );
  XNOR U11002 ( .A(n10811), .B(n10812), .Z(n10813) );
  XOR U11003 ( .A(n10814), .B(n10813), .Z(n10744) );
  NANDN U11004 ( .A(n10734), .B(n10733), .Z(n10738) );
  NANDN U11005 ( .A(n10736), .B(n10735), .Z(n10737) );
  NAND U11006 ( .A(n10738), .B(n10737), .Z(n10745) );
  XNOR U11007 ( .A(n10744), .B(n10745), .Z(n10746) );
  XNOR U11008 ( .A(n10747), .B(n10746), .Z(n10817) );
  XNOR U11009 ( .A(n10817), .B(sreg[384]), .Z(n10819) );
  NAND U11010 ( .A(n10739), .B(sreg[383]), .Z(n10743) );
  OR U11011 ( .A(n10741), .B(n10740), .Z(n10742) );
  AND U11012 ( .A(n10743), .B(n10742), .Z(n10818) );
  XOR U11013 ( .A(n10819), .B(n10818), .Z(c[384]) );
  NANDN U11014 ( .A(n10745), .B(n10744), .Z(n10749) );
  NAND U11015 ( .A(n10747), .B(n10746), .Z(n10748) );
  NAND U11016 ( .A(n10749), .B(n10748), .Z(n10825) );
  NANDN U11017 ( .A(n10751), .B(n10750), .Z(n10755) );
  OR U11018 ( .A(n10753), .B(n10752), .Z(n10754) );
  NAND U11019 ( .A(n10755), .B(n10754), .Z(n10892) );
  NANDN U11020 ( .A(n10757), .B(n10756), .Z(n10761) );
  OR U11021 ( .A(n10759), .B(n10758), .Z(n10760) );
  NAND U11022 ( .A(n10761), .B(n10760), .Z(n10880) );
  NAND U11023 ( .A(b[0]), .B(a[145]), .Z(n10762) );
  XNOR U11024 ( .A(b[1]), .B(n10762), .Z(n10764) );
  NAND U11025 ( .A(a[144]), .B(n98), .Z(n10763) );
  AND U11026 ( .A(n10764), .B(n10763), .Z(n10856) );
  XNOR U11027 ( .A(n20154), .B(n10942), .Z(n10865) );
  OR U11028 ( .A(n10865), .B(n20057), .Z(n10767) );
  NANDN U11029 ( .A(n10765), .B(n20098), .Z(n10766) );
  AND U11030 ( .A(n10767), .B(n10766), .Z(n10857) );
  XOR U11031 ( .A(n10856), .B(n10857), .Z(n10859) );
  NAND U11032 ( .A(a[129]), .B(b[15]), .Z(n10858) );
  XOR U11033 ( .A(n10859), .B(n10858), .Z(n10877) );
  NAND U11034 ( .A(n19722), .B(n10768), .Z(n10770) );
  XNOR U11035 ( .A(b[5]), .B(n11539), .Z(n10868) );
  NANDN U11036 ( .A(n19640), .B(n10868), .Z(n10769) );
  NAND U11037 ( .A(n10770), .B(n10769), .Z(n10853) );
  XNOR U11038 ( .A(n19714), .B(n11410), .Z(n10871) );
  NANDN U11039 ( .A(n10871), .B(n19766), .Z(n10773) );
  NANDN U11040 ( .A(n10771), .B(n19767), .Z(n10772) );
  NAND U11041 ( .A(n10773), .B(n10772), .Z(n10850) );
  NAND U11042 ( .A(n19554), .B(n10774), .Z(n10776) );
  IV U11043 ( .A(a[143]), .Z(n11722) );
  XNOR U11044 ( .A(b[3]), .B(n11722), .Z(n10874) );
  NANDN U11045 ( .A(n19521), .B(n10874), .Z(n10775) );
  AND U11046 ( .A(n10776), .B(n10775), .Z(n10851) );
  XNOR U11047 ( .A(n10850), .B(n10851), .Z(n10852) );
  XOR U11048 ( .A(n10853), .B(n10852), .Z(n10878) );
  XOR U11049 ( .A(n10877), .B(n10878), .Z(n10879) );
  XNOR U11050 ( .A(n10880), .B(n10879), .Z(n10828) );
  NAND U11051 ( .A(n10778), .B(n10777), .Z(n10782) );
  NAND U11052 ( .A(n10780), .B(n10779), .Z(n10781) );
  NAND U11053 ( .A(n10782), .B(n10781), .Z(n10829) );
  XOR U11054 ( .A(n10828), .B(n10829), .Z(n10831) );
  XNOR U11055 ( .A(n20052), .B(n11098), .Z(n10834) );
  OR U11056 ( .A(n10834), .B(n20020), .Z(n10785) );
  NANDN U11057 ( .A(n10783), .B(n19960), .Z(n10784) );
  NAND U11058 ( .A(n10785), .B(n10784), .Z(n10847) );
  XNOR U11059 ( .A(n102), .B(n10786), .Z(n10838) );
  OR U11060 ( .A(n10838), .B(n20121), .Z(n10789) );
  NANDN U11061 ( .A(n10787), .B(n20122), .Z(n10788) );
  NAND U11062 ( .A(n10789), .B(n10788), .Z(n10844) );
  XNOR U11063 ( .A(n19975), .B(n11254), .Z(n10841) );
  NANDN U11064 ( .A(n10841), .B(n19883), .Z(n10792) );
  NANDN U11065 ( .A(n10790), .B(n19937), .Z(n10791) );
  AND U11066 ( .A(n10792), .B(n10791), .Z(n10845) );
  XNOR U11067 ( .A(n10844), .B(n10845), .Z(n10846) );
  XNOR U11068 ( .A(n10847), .B(n10846), .Z(n10883) );
  NANDN U11069 ( .A(n10794), .B(n10793), .Z(n10798) );
  NAND U11070 ( .A(n10796), .B(n10795), .Z(n10797) );
  NAND U11071 ( .A(n10798), .B(n10797), .Z(n10884) );
  XNOR U11072 ( .A(n10883), .B(n10884), .Z(n10885) );
  NANDN U11073 ( .A(n10800), .B(n10799), .Z(n10804) );
  NAND U11074 ( .A(n10802), .B(n10801), .Z(n10803) );
  AND U11075 ( .A(n10804), .B(n10803), .Z(n10886) );
  XNOR U11076 ( .A(n10885), .B(n10886), .Z(n10830) );
  XNOR U11077 ( .A(n10831), .B(n10830), .Z(n10889) );
  NANDN U11078 ( .A(n10806), .B(n10805), .Z(n10810) );
  NAND U11079 ( .A(n10808), .B(n10807), .Z(n10809) );
  NAND U11080 ( .A(n10810), .B(n10809), .Z(n10890) );
  XNOR U11081 ( .A(n10889), .B(n10890), .Z(n10891) );
  XOR U11082 ( .A(n10892), .B(n10891), .Z(n10822) );
  NANDN U11083 ( .A(n10812), .B(n10811), .Z(n10816) );
  NANDN U11084 ( .A(n10814), .B(n10813), .Z(n10815) );
  NAND U11085 ( .A(n10816), .B(n10815), .Z(n10823) );
  XNOR U11086 ( .A(n10822), .B(n10823), .Z(n10824) );
  XNOR U11087 ( .A(n10825), .B(n10824), .Z(n10895) );
  XNOR U11088 ( .A(n10895), .B(sreg[385]), .Z(n10897) );
  NAND U11089 ( .A(n10817), .B(sreg[384]), .Z(n10821) );
  OR U11090 ( .A(n10819), .B(n10818), .Z(n10820) );
  AND U11091 ( .A(n10821), .B(n10820), .Z(n10896) );
  XOR U11092 ( .A(n10897), .B(n10896), .Z(c[385]) );
  NANDN U11093 ( .A(n10823), .B(n10822), .Z(n10827) );
  NAND U11094 ( .A(n10825), .B(n10824), .Z(n10826) );
  NAND U11095 ( .A(n10827), .B(n10826), .Z(n10903) );
  NANDN U11096 ( .A(n10829), .B(n10828), .Z(n10833) );
  OR U11097 ( .A(n10831), .B(n10830), .Z(n10832) );
  NAND U11098 ( .A(n10833), .B(n10832), .Z(n10970) );
  XNOR U11099 ( .A(n20052), .B(n11149), .Z(n10939) );
  OR U11100 ( .A(n10939), .B(n20020), .Z(n10836) );
  NANDN U11101 ( .A(n10834), .B(n19960), .Z(n10835) );
  NAND U11102 ( .A(n10836), .B(n10835), .Z(n10952) );
  XNOR U11103 ( .A(n102), .B(n10837), .Z(n10943) );
  OR U11104 ( .A(n10943), .B(n20121), .Z(n10840) );
  NANDN U11105 ( .A(n10838), .B(n20122), .Z(n10839) );
  NAND U11106 ( .A(n10840), .B(n10839), .Z(n10949) );
  XNOR U11107 ( .A(n19975), .B(n11305), .Z(n10946) );
  NANDN U11108 ( .A(n10946), .B(n19883), .Z(n10843) );
  NANDN U11109 ( .A(n10841), .B(n19937), .Z(n10842) );
  AND U11110 ( .A(n10843), .B(n10842), .Z(n10950) );
  XNOR U11111 ( .A(n10949), .B(n10950), .Z(n10951) );
  XNOR U11112 ( .A(n10952), .B(n10951), .Z(n10961) );
  NANDN U11113 ( .A(n10845), .B(n10844), .Z(n10849) );
  NAND U11114 ( .A(n10847), .B(n10846), .Z(n10848) );
  NAND U11115 ( .A(n10849), .B(n10848), .Z(n10962) );
  XNOR U11116 ( .A(n10961), .B(n10962), .Z(n10963) );
  NANDN U11117 ( .A(n10851), .B(n10850), .Z(n10855) );
  NAND U11118 ( .A(n10853), .B(n10852), .Z(n10854) );
  AND U11119 ( .A(n10855), .B(n10854), .Z(n10964) );
  XNOR U11120 ( .A(n10963), .B(n10964), .Z(n10908) );
  NANDN U11121 ( .A(n10857), .B(n10856), .Z(n10861) );
  OR U11122 ( .A(n10859), .B(n10858), .Z(n10860) );
  NAND U11123 ( .A(n10861), .B(n10860), .Z(n10936) );
  NAND U11124 ( .A(b[0]), .B(a[146]), .Z(n10862) );
  XNOR U11125 ( .A(b[1]), .B(n10862), .Z(n10864) );
  NAND U11126 ( .A(a[145]), .B(n98), .Z(n10863) );
  AND U11127 ( .A(n10864), .B(n10863), .Z(n10912) );
  XNOR U11128 ( .A(n20154), .B(n11020), .Z(n10921) );
  OR U11129 ( .A(n10921), .B(n20057), .Z(n10867) );
  NANDN U11130 ( .A(n10865), .B(n20098), .Z(n10866) );
  AND U11131 ( .A(n10867), .B(n10866), .Z(n10913) );
  XOR U11132 ( .A(n10912), .B(n10913), .Z(n10915) );
  NAND U11133 ( .A(a[130]), .B(b[15]), .Z(n10914) );
  XOR U11134 ( .A(n10915), .B(n10914), .Z(n10933) );
  NAND U11135 ( .A(n19722), .B(n10868), .Z(n10870) );
  XNOR U11136 ( .A(b[5]), .B(n11644), .Z(n10924) );
  NANDN U11137 ( .A(n19640), .B(n10924), .Z(n10869) );
  NAND U11138 ( .A(n10870), .B(n10869), .Z(n10958) );
  XNOR U11139 ( .A(n19714), .B(n11461), .Z(n10927) );
  NANDN U11140 ( .A(n10927), .B(n19766), .Z(n10873) );
  NANDN U11141 ( .A(n10871), .B(n19767), .Z(n10872) );
  NAND U11142 ( .A(n10873), .B(n10872), .Z(n10955) );
  NAND U11143 ( .A(n19554), .B(n10874), .Z(n10876) );
  IV U11144 ( .A(a[144]), .Z(n11773) );
  XNOR U11145 ( .A(b[3]), .B(n11773), .Z(n10930) );
  NANDN U11146 ( .A(n19521), .B(n10930), .Z(n10875) );
  AND U11147 ( .A(n10876), .B(n10875), .Z(n10956) );
  XNOR U11148 ( .A(n10955), .B(n10956), .Z(n10957) );
  XOR U11149 ( .A(n10958), .B(n10957), .Z(n10934) );
  XOR U11150 ( .A(n10933), .B(n10934), .Z(n10935) );
  XNOR U11151 ( .A(n10936), .B(n10935), .Z(n10906) );
  NAND U11152 ( .A(n10878), .B(n10877), .Z(n10882) );
  NAND U11153 ( .A(n10880), .B(n10879), .Z(n10881) );
  NAND U11154 ( .A(n10882), .B(n10881), .Z(n10907) );
  XOR U11155 ( .A(n10906), .B(n10907), .Z(n10909) );
  XNOR U11156 ( .A(n10908), .B(n10909), .Z(n10967) );
  NANDN U11157 ( .A(n10884), .B(n10883), .Z(n10888) );
  NAND U11158 ( .A(n10886), .B(n10885), .Z(n10887) );
  NAND U11159 ( .A(n10888), .B(n10887), .Z(n10968) );
  XNOR U11160 ( .A(n10967), .B(n10968), .Z(n10969) );
  XOR U11161 ( .A(n10970), .B(n10969), .Z(n10900) );
  NANDN U11162 ( .A(n10890), .B(n10889), .Z(n10894) );
  NANDN U11163 ( .A(n10892), .B(n10891), .Z(n10893) );
  NAND U11164 ( .A(n10894), .B(n10893), .Z(n10901) );
  XNOR U11165 ( .A(n10900), .B(n10901), .Z(n10902) );
  XNOR U11166 ( .A(n10903), .B(n10902), .Z(n10973) );
  XNOR U11167 ( .A(n10973), .B(sreg[386]), .Z(n10975) );
  NAND U11168 ( .A(n10895), .B(sreg[385]), .Z(n10899) );
  OR U11169 ( .A(n10897), .B(n10896), .Z(n10898) );
  AND U11170 ( .A(n10899), .B(n10898), .Z(n10974) );
  XOR U11171 ( .A(n10975), .B(n10974), .Z(c[386]) );
  NANDN U11172 ( .A(n10901), .B(n10900), .Z(n10905) );
  NAND U11173 ( .A(n10903), .B(n10902), .Z(n10904) );
  NAND U11174 ( .A(n10905), .B(n10904), .Z(n10981) );
  NANDN U11175 ( .A(n10907), .B(n10906), .Z(n10911) );
  OR U11176 ( .A(n10909), .B(n10908), .Z(n10910) );
  NAND U11177 ( .A(n10911), .B(n10910), .Z(n11048) );
  NANDN U11178 ( .A(n10913), .B(n10912), .Z(n10917) );
  OR U11179 ( .A(n10915), .B(n10914), .Z(n10916) );
  NAND U11180 ( .A(n10917), .B(n10916), .Z(n11014) );
  NAND U11181 ( .A(b[0]), .B(a[147]), .Z(n10918) );
  XNOR U11182 ( .A(b[1]), .B(n10918), .Z(n10920) );
  NAND U11183 ( .A(a[146]), .B(n98), .Z(n10919) );
  AND U11184 ( .A(n10920), .B(n10919), .Z(n10990) );
  XNOR U11185 ( .A(n20154), .B(n11098), .Z(n10999) );
  OR U11186 ( .A(n10999), .B(n20057), .Z(n10923) );
  NANDN U11187 ( .A(n10921), .B(n20098), .Z(n10922) );
  AND U11188 ( .A(n10923), .B(n10922), .Z(n10991) );
  XOR U11189 ( .A(n10990), .B(n10991), .Z(n10993) );
  NAND U11190 ( .A(a[131]), .B(b[15]), .Z(n10992) );
  XOR U11191 ( .A(n10993), .B(n10992), .Z(n11011) );
  NAND U11192 ( .A(n19722), .B(n10924), .Z(n10926) );
  XNOR U11193 ( .A(b[5]), .B(n11722), .Z(n11002) );
  NANDN U11194 ( .A(n19640), .B(n11002), .Z(n10925) );
  NAND U11195 ( .A(n10926), .B(n10925), .Z(n11036) );
  XNOR U11196 ( .A(n19714), .B(n11539), .Z(n11005) );
  NANDN U11197 ( .A(n11005), .B(n19766), .Z(n10929) );
  NANDN U11198 ( .A(n10927), .B(n19767), .Z(n10928) );
  NAND U11199 ( .A(n10929), .B(n10928), .Z(n11033) );
  NAND U11200 ( .A(n19554), .B(n10930), .Z(n10932) );
  IV U11201 ( .A(a[145]), .Z(n11851) );
  XNOR U11202 ( .A(b[3]), .B(n11851), .Z(n11008) );
  NANDN U11203 ( .A(n19521), .B(n11008), .Z(n10931) );
  AND U11204 ( .A(n10932), .B(n10931), .Z(n11034) );
  XNOR U11205 ( .A(n11033), .B(n11034), .Z(n11035) );
  XOR U11206 ( .A(n11036), .B(n11035), .Z(n11012) );
  XOR U11207 ( .A(n11011), .B(n11012), .Z(n11013) );
  XNOR U11208 ( .A(n11014), .B(n11013), .Z(n10984) );
  NAND U11209 ( .A(n10934), .B(n10933), .Z(n10938) );
  NAND U11210 ( .A(n10936), .B(n10935), .Z(n10937) );
  NAND U11211 ( .A(n10938), .B(n10937), .Z(n10985) );
  XOR U11212 ( .A(n10984), .B(n10985), .Z(n10987) );
  XNOR U11213 ( .A(n20052), .B(n11254), .Z(n11017) );
  OR U11214 ( .A(n11017), .B(n20020), .Z(n10941) );
  NANDN U11215 ( .A(n10939), .B(n19960), .Z(n10940) );
  NAND U11216 ( .A(n10941), .B(n10940), .Z(n11030) );
  XNOR U11217 ( .A(n102), .B(n10942), .Z(n11021) );
  OR U11218 ( .A(n11021), .B(n20121), .Z(n10945) );
  NANDN U11219 ( .A(n10943), .B(n20122), .Z(n10944) );
  NAND U11220 ( .A(n10945), .B(n10944), .Z(n11027) );
  XNOR U11221 ( .A(n19975), .B(n11410), .Z(n11024) );
  NANDN U11222 ( .A(n11024), .B(n19883), .Z(n10948) );
  NANDN U11223 ( .A(n10946), .B(n19937), .Z(n10947) );
  AND U11224 ( .A(n10948), .B(n10947), .Z(n11028) );
  XNOR U11225 ( .A(n11027), .B(n11028), .Z(n11029) );
  XNOR U11226 ( .A(n11030), .B(n11029), .Z(n11039) );
  NANDN U11227 ( .A(n10950), .B(n10949), .Z(n10954) );
  NAND U11228 ( .A(n10952), .B(n10951), .Z(n10953) );
  NAND U11229 ( .A(n10954), .B(n10953), .Z(n11040) );
  XNOR U11230 ( .A(n11039), .B(n11040), .Z(n11041) );
  NANDN U11231 ( .A(n10956), .B(n10955), .Z(n10960) );
  NAND U11232 ( .A(n10958), .B(n10957), .Z(n10959) );
  AND U11233 ( .A(n10960), .B(n10959), .Z(n11042) );
  XNOR U11234 ( .A(n11041), .B(n11042), .Z(n10986) );
  XNOR U11235 ( .A(n10987), .B(n10986), .Z(n11045) );
  NANDN U11236 ( .A(n10962), .B(n10961), .Z(n10966) );
  NAND U11237 ( .A(n10964), .B(n10963), .Z(n10965) );
  NAND U11238 ( .A(n10966), .B(n10965), .Z(n11046) );
  XNOR U11239 ( .A(n11045), .B(n11046), .Z(n11047) );
  XOR U11240 ( .A(n11048), .B(n11047), .Z(n10978) );
  NANDN U11241 ( .A(n10968), .B(n10967), .Z(n10972) );
  NANDN U11242 ( .A(n10970), .B(n10969), .Z(n10971) );
  NAND U11243 ( .A(n10972), .B(n10971), .Z(n10979) );
  XNOR U11244 ( .A(n10978), .B(n10979), .Z(n10980) );
  XNOR U11245 ( .A(n10981), .B(n10980), .Z(n11051) );
  XNOR U11246 ( .A(n11051), .B(sreg[387]), .Z(n11053) );
  NAND U11247 ( .A(n10973), .B(sreg[386]), .Z(n10977) );
  OR U11248 ( .A(n10975), .B(n10974), .Z(n10976) );
  AND U11249 ( .A(n10977), .B(n10976), .Z(n11052) );
  XOR U11250 ( .A(n11053), .B(n11052), .Z(c[387]) );
  NANDN U11251 ( .A(n10979), .B(n10978), .Z(n10983) );
  NAND U11252 ( .A(n10981), .B(n10980), .Z(n10982) );
  NAND U11253 ( .A(n10983), .B(n10982), .Z(n11059) );
  NANDN U11254 ( .A(n10985), .B(n10984), .Z(n10989) );
  OR U11255 ( .A(n10987), .B(n10986), .Z(n10988) );
  NAND U11256 ( .A(n10989), .B(n10988), .Z(n11126) );
  NANDN U11257 ( .A(n10991), .B(n10990), .Z(n10995) );
  OR U11258 ( .A(n10993), .B(n10992), .Z(n10994) );
  NAND U11259 ( .A(n10995), .B(n10994), .Z(n11092) );
  NAND U11260 ( .A(b[0]), .B(a[148]), .Z(n10996) );
  XNOR U11261 ( .A(b[1]), .B(n10996), .Z(n10998) );
  NAND U11262 ( .A(a[147]), .B(n98), .Z(n10997) );
  AND U11263 ( .A(n10998), .B(n10997), .Z(n11068) );
  XNOR U11264 ( .A(n20154), .B(n11149), .Z(n11077) );
  OR U11265 ( .A(n11077), .B(n20057), .Z(n11001) );
  NANDN U11266 ( .A(n10999), .B(n20098), .Z(n11000) );
  AND U11267 ( .A(n11001), .B(n11000), .Z(n11069) );
  XOR U11268 ( .A(n11068), .B(n11069), .Z(n11071) );
  NAND U11269 ( .A(a[132]), .B(b[15]), .Z(n11070) );
  XOR U11270 ( .A(n11071), .B(n11070), .Z(n11089) );
  NAND U11271 ( .A(n19722), .B(n11002), .Z(n11004) );
  XNOR U11272 ( .A(b[5]), .B(n11773), .Z(n11080) );
  NANDN U11273 ( .A(n19640), .B(n11080), .Z(n11003) );
  NAND U11274 ( .A(n11004), .B(n11003), .Z(n11114) );
  XNOR U11275 ( .A(n19714), .B(n11644), .Z(n11083) );
  NANDN U11276 ( .A(n11083), .B(n19766), .Z(n11007) );
  NANDN U11277 ( .A(n11005), .B(n19767), .Z(n11006) );
  NAND U11278 ( .A(n11007), .B(n11006), .Z(n11111) );
  NAND U11279 ( .A(n19554), .B(n11008), .Z(n11010) );
  IV U11280 ( .A(a[146]), .Z(n11929) );
  XNOR U11281 ( .A(b[3]), .B(n11929), .Z(n11086) );
  NANDN U11282 ( .A(n19521), .B(n11086), .Z(n11009) );
  AND U11283 ( .A(n11010), .B(n11009), .Z(n11112) );
  XNOR U11284 ( .A(n11111), .B(n11112), .Z(n11113) );
  XOR U11285 ( .A(n11114), .B(n11113), .Z(n11090) );
  XOR U11286 ( .A(n11089), .B(n11090), .Z(n11091) );
  XNOR U11287 ( .A(n11092), .B(n11091), .Z(n11062) );
  NAND U11288 ( .A(n11012), .B(n11011), .Z(n11016) );
  NAND U11289 ( .A(n11014), .B(n11013), .Z(n11015) );
  NAND U11290 ( .A(n11016), .B(n11015), .Z(n11063) );
  XOR U11291 ( .A(n11062), .B(n11063), .Z(n11065) );
  XNOR U11292 ( .A(n20052), .B(n11305), .Z(n11095) );
  OR U11293 ( .A(n11095), .B(n20020), .Z(n11019) );
  NANDN U11294 ( .A(n11017), .B(n19960), .Z(n11018) );
  NAND U11295 ( .A(n11019), .B(n11018), .Z(n11108) );
  XNOR U11296 ( .A(n102), .B(n11020), .Z(n11099) );
  OR U11297 ( .A(n11099), .B(n20121), .Z(n11023) );
  NANDN U11298 ( .A(n11021), .B(n20122), .Z(n11022) );
  NAND U11299 ( .A(n11023), .B(n11022), .Z(n11105) );
  XNOR U11300 ( .A(n19975), .B(n11461), .Z(n11102) );
  NANDN U11301 ( .A(n11102), .B(n19883), .Z(n11026) );
  NANDN U11302 ( .A(n11024), .B(n19937), .Z(n11025) );
  AND U11303 ( .A(n11026), .B(n11025), .Z(n11106) );
  XNOR U11304 ( .A(n11105), .B(n11106), .Z(n11107) );
  XNOR U11305 ( .A(n11108), .B(n11107), .Z(n11117) );
  NANDN U11306 ( .A(n11028), .B(n11027), .Z(n11032) );
  NAND U11307 ( .A(n11030), .B(n11029), .Z(n11031) );
  NAND U11308 ( .A(n11032), .B(n11031), .Z(n11118) );
  XNOR U11309 ( .A(n11117), .B(n11118), .Z(n11119) );
  NANDN U11310 ( .A(n11034), .B(n11033), .Z(n11038) );
  NAND U11311 ( .A(n11036), .B(n11035), .Z(n11037) );
  AND U11312 ( .A(n11038), .B(n11037), .Z(n11120) );
  XNOR U11313 ( .A(n11119), .B(n11120), .Z(n11064) );
  XNOR U11314 ( .A(n11065), .B(n11064), .Z(n11123) );
  NANDN U11315 ( .A(n11040), .B(n11039), .Z(n11044) );
  NAND U11316 ( .A(n11042), .B(n11041), .Z(n11043) );
  NAND U11317 ( .A(n11044), .B(n11043), .Z(n11124) );
  XNOR U11318 ( .A(n11123), .B(n11124), .Z(n11125) );
  XOR U11319 ( .A(n11126), .B(n11125), .Z(n11056) );
  NANDN U11320 ( .A(n11046), .B(n11045), .Z(n11050) );
  NANDN U11321 ( .A(n11048), .B(n11047), .Z(n11049) );
  NAND U11322 ( .A(n11050), .B(n11049), .Z(n11057) );
  XNOR U11323 ( .A(n11056), .B(n11057), .Z(n11058) );
  XNOR U11324 ( .A(n11059), .B(n11058), .Z(n11129) );
  XNOR U11325 ( .A(n11129), .B(sreg[388]), .Z(n11131) );
  NAND U11326 ( .A(n11051), .B(sreg[387]), .Z(n11055) );
  OR U11327 ( .A(n11053), .B(n11052), .Z(n11054) );
  AND U11328 ( .A(n11055), .B(n11054), .Z(n11130) );
  XOR U11329 ( .A(n11131), .B(n11130), .Z(c[388]) );
  NANDN U11330 ( .A(n11057), .B(n11056), .Z(n11061) );
  NAND U11331 ( .A(n11059), .B(n11058), .Z(n11060) );
  NAND U11332 ( .A(n11061), .B(n11060), .Z(n11137) );
  NANDN U11333 ( .A(n11063), .B(n11062), .Z(n11067) );
  OR U11334 ( .A(n11065), .B(n11064), .Z(n11066) );
  NAND U11335 ( .A(n11067), .B(n11066), .Z(n11204) );
  NANDN U11336 ( .A(n11069), .B(n11068), .Z(n11073) );
  OR U11337 ( .A(n11071), .B(n11070), .Z(n11072) );
  NAND U11338 ( .A(n11073), .B(n11072), .Z(n11192) );
  NAND U11339 ( .A(b[0]), .B(a[149]), .Z(n11074) );
  XNOR U11340 ( .A(b[1]), .B(n11074), .Z(n11076) );
  NAND U11341 ( .A(a[148]), .B(n98), .Z(n11075) );
  AND U11342 ( .A(n11076), .B(n11075), .Z(n11168) );
  XNOR U11343 ( .A(n20154), .B(n11254), .Z(n11177) );
  OR U11344 ( .A(n11177), .B(n20057), .Z(n11079) );
  NANDN U11345 ( .A(n11077), .B(n20098), .Z(n11078) );
  AND U11346 ( .A(n11079), .B(n11078), .Z(n11169) );
  XOR U11347 ( .A(n11168), .B(n11169), .Z(n11171) );
  NAND U11348 ( .A(a[133]), .B(b[15]), .Z(n11170) );
  XOR U11349 ( .A(n11171), .B(n11170), .Z(n11189) );
  NAND U11350 ( .A(n19722), .B(n11080), .Z(n11082) );
  XNOR U11351 ( .A(b[5]), .B(n11851), .Z(n11180) );
  NANDN U11352 ( .A(n19640), .B(n11180), .Z(n11081) );
  NAND U11353 ( .A(n11082), .B(n11081), .Z(n11165) );
  XNOR U11354 ( .A(n19714), .B(n11722), .Z(n11183) );
  NANDN U11355 ( .A(n11183), .B(n19766), .Z(n11085) );
  NANDN U11356 ( .A(n11083), .B(n19767), .Z(n11084) );
  NAND U11357 ( .A(n11085), .B(n11084), .Z(n11162) );
  NAND U11358 ( .A(n19554), .B(n11086), .Z(n11088) );
  IV U11359 ( .A(a[147]), .Z(n12007) );
  XNOR U11360 ( .A(b[3]), .B(n12007), .Z(n11186) );
  NANDN U11361 ( .A(n19521), .B(n11186), .Z(n11087) );
  AND U11362 ( .A(n11088), .B(n11087), .Z(n11163) );
  XNOR U11363 ( .A(n11162), .B(n11163), .Z(n11164) );
  XOR U11364 ( .A(n11165), .B(n11164), .Z(n11190) );
  XOR U11365 ( .A(n11189), .B(n11190), .Z(n11191) );
  XNOR U11366 ( .A(n11192), .B(n11191), .Z(n11140) );
  NAND U11367 ( .A(n11090), .B(n11089), .Z(n11094) );
  NAND U11368 ( .A(n11092), .B(n11091), .Z(n11093) );
  NAND U11369 ( .A(n11094), .B(n11093), .Z(n11141) );
  XOR U11370 ( .A(n11140), .B(n11141), .Z(n11143) );
  XNOR U11371 ( .A(n20052), .B(n11410), .Z(n11146) );
  OR U11372 ( .A(n11146), .B(n20020), .Z(n11097) );
  NANDN U11373 ( .A(n11095), .B(n19960), .Z(n11096) );
  NAND U11374 ( .A(n11097), .B(n11096), .Z(n11159) );
  XNOR U11375 ( .A(n102), .B(n11098), .Z(n11150) );
  OR U11376 ( .A(n11150), .B(n20121), .Z(n11101) );
  NANDN U11377 ( .A(n11099), .B(n20122), .Z(n11100) );
  NAND U11378 ( .A(n11101), .B(n11100), .Z(n11156) );
  XNOR U11379 ( .A(n19975), .B(n11539), .Z(n11153) );
  NANDN U11380 ( .A(n11153), .B(n19883), .Z(n11104) );
  NANDN U11381 ( .A(n11102), .B(n19937), .Z(n11103) );
  AND U11382 ( .A(n11104), .B(n11103), .Z(n11157) );
  XNOR U11383 ( .A(n11156), .B(n11157), .Z(n11158) );
  XNOR U11384 ( .A(n11159), .B(n11158), .Z(n11195) );
  NANDN U11385 ( .A(n11106), .B(n11105), .Z(n11110) );
  NAND U11386 ( .A(n11108), .B(n11107), .Z(n11109) );
  NAND U11387 ( .A(n11110), .B(n11109), .Z(n11196) );
  XNOR U11388 ( .A(n11195), .B(n11196), .Z(n11197) );
  NANDN U11389 ( .A(n11112), .B(n11111), .Z(n11116) );
  NAND U11390 ( .A(n11114), .B(n11113), .Z(n11115) );
  AND U11391 ( .A(n11116), .B(n11115), .Z(n11198) );
  XNOR U11392 ( .A(n11197), .B(n11198), .Z(n11142) );
  XNOR U11393 ( .A(n11143), .B(n11142), .Z(n11201) );
  NANDN U11394 ( .A(n11118), .B(n11117), .Z(n11122) );
  NAND U11395 ( .A(n11120), .B(n11119), .Z(n11121) );
  NAND U11396 ( .A(n11122), .B(n11121), .Z(n11202) );
  XNOR U11397 ( .A(n11201), .B(n11202), .Z(n11203) );
  XOR U11398 ( .A(n11204), .B(n11203), .Z(n11134) );
  NANDN U11399 ( .A(n11124), .B(n11123), .Z(n11128) );
  NANDN U11400 ( .A(n11126), .B(n11125), .Z(n11127) );
  NAND U11401 ( .A(n11128), .B(n11127), .Z(n11135) );
  XNOR U11402 ( .A(n11134), .B(n11135), .Z(n11136) );
  XNOR U11403 ( .A(n11137), .B(n11136), .Z(n11207) );
  XNOR U11404 ( .A(n11207), .B(sreg[389]), .Z(n11209) );
  NAND U11405 ( .A(n11129), .B(sreg[388]), .Z(n11133) );
  OR U11406 ( .A(n11131), .B(n11130), .Z(n11132) );
  AND U11407 ( .A(n11133), .B(n11132), .Z(n11208) );
  XOR U11408 ( .A(n11209), .B(n11208), .Z(c[389]) );
  NANDN U11409 ( .A(n11135), .B(n11134), .Z(n11139) );
  NAND U11410 ( .A(n11137), .B(n11136), .Z(n11138) );
  NAND U11411 ( .A(n11139), .B(n11138), .Z(n11215) );
  NANDN U11412 ( .A(n11141), .B(n11140), .Z(n11145) );
  OR U11413 ( .A(n11143), .B(n11142), .Z(n11144) );
  NAND U11414 ( .A(n11145), .B(n11144), .Z(n11282) );
  XNOR U11415 ( .A(n20052), .B(n11461), .Z(n11251) );
  OR U11416 ( .A(n11251), .B(n20020), .Z(n11148) );
  NANDN U11417 ( .A(n11146), .B(n19960), .Z(n11147) );
  NAND U11418 ( .A(n11148), .B(n11147), .Z(n11264) );
  XNOR U11419 ( .A(n102), .B(n11149), .Z(n11255) );
  OR U11420 ( .A(n11255), .B(n20121), .Z(n11152) );
  NANDN U11421 ( .A(n11150), .B(n20122), .Z(n11151) );
  NAND U11422 ( .A(n11152), .B(n11151), .Z(n11261) );
  XNOR U11423 ( .A(n19975), .B(n11644), .Z(n11258) );
  NANDN U11424 ( .A(n11258), .B(n19883), .Z(n11155) );
  NANDN U11425 ( .A(n11153), .B(n19937), .Z(n11154) );
  AND U11426 ( .A(n11155), .B(n11154), .Z(n11262) );
  XNOR U11427 ( .A(n11261), .B(n11262), .Z(n11263) );
  XNOR U11428 ( .A(n11264), .B(n11263), .Z(n11273) );
  NANDN U11429 ( .A(n11157), .B(n11156), .Z(n11161) );
  NAND U11430 ( .A(n11159), .B(n11158), .Z(n11160) );
  NAND U11431 ( .A(n11161), .B(n11160), .Z(n11274) );
  XNOR U11432 ( .A(n11273), .B(n11274), .Z(n11275) );
  NANDN U11433 ( .A(n11163), .B(n11162), .Z(n11167) );
  NAND U11434 ( .A(n11165), .B(n11164), .Z(n11166) );
  AND U11435 ( .A(n11167), .B(n11166), .Z(n11276) );
  XNOR U11436 ( .A(n11275), .B(n11276), .Z(n11220) );
  NANDN U11437 ( .A(n11169), .B(n11168), .Z(n11173) );
  OR U11438 ( .A(n11171), .B(n11170), .Z(n11172) );
  NAND U11439 ( .A(n11173), .B(n11172), .Z(n11248) );
  NAND U11440 ( .A(b[0]), .B(a[150]), .Z(n11174) );
  XNOR U11441 ( .A(b[1]), .B(n11174), .Z(n11176) );
  NAND U11442 ( .A(a[149]), .B(n98), .Z(n11175) );
  AND U11443 ( .A(n11176), .B(n11175), .Z(n11224) );
  XNOR U11444 ( .A(n20154), .B(n11305), .Z(n11230) );
  OR U11445 ( .A(n11230), .B(n20057), .Z(n11179) );
  NANDN U11446 ( .A(n11177), .B(n20098), .Z(n11178) );
  AND U11447 ( .A(n11179), .B(n11178), .Z(n11225) );
  XOR U11448 ( .A(n11224), .B(n11225), .Z(n11227) );
  NAND U11449 ( .A(a[134]), .B(b[15]), .Z(n11226) );
  XOR U11450 ( .A(n11227), .B(n11226), .Z(n11245) );
  NAND U11451 ( .A(n19722), .B(n11180), .Z(n11182) );
  XNOR U11452 ( .A(b[5]), .B(n11929), .Z(n11236) );
  NANDN U11453 ( .A(n19640), .B(n11236), .Z(n11181) );
  NAND U11454 ( .A(n11182), .B(n11181), .Z(n11270) );
  XNOR U11455 ( .A(n19714), .B(n11773), .Z(n11239) );
  NANDN U11456 ( .A(n11239), .B(n19766), .Z(n11185) );
  NANDN U11457 ( .A(n11183), .B(n19767), .Z(n11184) );
  NAND U11458 ( .A(n11185), .B(n11184), .Z(n11267) );
  NAND U11459 ( .A(n19554), .B(n11186), .Z(n11188) );
  IV U11460 ( .A(a[148]), .Z(n12112) );
  XNOR U11461 ( .A(b[3]), .B(n12112), .Z(n11242) );
  NANDN U11462 ( .A(n19521), .B(n11242), .Z(n11187) );
  AND U11463 ( .A(n11188), .B(n11187), .Z(n11268) );
  XNOR U11464 ( .A(n11267), .B(n11268), .Z(n11269) );
  XOR U11465 ( .A(n11270), .B(n11269), .Z(n11246) );
  XOR U11466 ( .A(n11245), .B(n11246), .Z(n11247) );
  XNOR U11467 ( .A(n11248), .B(n11247), .Z(n11218) );
  NAND U11468 ( .A(n11190), .B(n11189), .Z(n11194) );
  NAND U11469 ( .A(n11192), .B(n11191), .Z(n11193) );
  NAND U11470 ( .A(n11194), .B(n11193), .Z(n11219) );
  XOR U11471 ( .A(n11218), .B(n11219), .Z(n11221) );
  XNOR U11472 ( .A(n11220), .B(n11221), .Z(n11279) );
  NANDN U11473 ( .A(n11196), .B(n11195), .Z(n11200) );
  NAND U11474 ( .A(n11198), .B(n11197), .Z(n11199) );
  NAND U11475 ( .A(n11200), .B(n11199), .Z(n11280) );
  XNOR U11476 ( .A(n11279), .B(n11280), .Z(n11281) );
  XOR U11477 ( .A(n11282), .B(n11281), .Z(n11212) );
  NANDN U11478 ( .A(n11202), .B(n11201), .Z(n11206) );
  NANDN U11479 ( .A(n11204), .B(n11203), .Z(n11205) );
  NAND U11480 ( .A(n11206), .B(n11205), .Z(n11213) );
  XNOR U11481 ( .A(n11212), .B(n11213), .Z(n11214) );
  XNOR U11482 ( .A(n11215), .B(n11214), .Z(n11285) );
  XNOR U11483 ( .A(n11285), .B(sreg[390]), .Z(n11287) );
  NAND U11484 ( .A(n11207), .B(sreg[389]), .Z(n11211) );
  OR U11485 ( .A(n11209), .B(n11208), .Z(n11210) );
  AND U11486 ( .A(n11211), .B(n11210), .Z(n11286) );
  XOR U11487 ( .A(n11287), .B(n11286), .Z(c[390]) );
  NANDN U11488 ( .A(n11213), .B(n11212), .Z(n11217) );
  NAND U11489 ( .A(n11215), .B(n11214), .Z(n11216) );
  NAND U11490 ( .A(n11217), .B(n11216), .Z(n11293) );
  NANDN U11491 ( .A(n11219), .B(n11218), .Z(n11223) );
  OR U11492 ( .A(n11221), .B(n11220), .Z(n11222) );
  NAND U11493 ( .A(n11223), .B(n11222), .Z(n11360) );
  NANDN U11494 ( .A(n11225), .B(n11224), .Z(n11229) );
  OR U11495 ( .A(n11227), .B(n11226), .Z(n11228) );
  NAND U11496 ( .A(n11229), .B(n11228), .Z(n11348) );
  XNOR U11497 ( .A(n20154), .B(n11410), .Z(n11333) );
  OR U11498 ( .A(n11333), .B(n20057), .Z(n11232) );
  NANDN U11499 ( .A(n11230), .B(n20098), .Z(n11231) );
  AND U11500 ( .A(n11232), .B(n11231), .Z(n11325) );
  NAND U11501 ( .A(b[0]), .B(a[151]), .Z(n11233) );
  XNOR U11502 ( .A(b[1]), .B(n11233), .Z(n11235) );
  NAND U11503 ( .A(a[150]), .B(n98), .Z(n11234) );
  AND U11504 ( .A(n11235), .B(n11234), .Z(n11324) );
  XOR U11505 ( .A(n11325), .B(n11324), .Z(n11327) );
  NAND U11506 ( .A(a[135]), .B(b[15]), .Z(n11326) );
  XOR U11507 ( .A(n11327), .B(n11326), .Z(n11345) );
  NAND U11508 ( .A(n19722), .B(n11236), .Z(n11238) );
  XNOR U11509 ( .A(b[5]), .B(n12007), .Z(n11336) );
  NANDN U11510 ( .A(n19640), .B(n11336), .Z(n11237) );
  NAND U11511 ( .A(n11238), .B(n11237), .Z(n11321) );
  XNOR U11512 ( .A(n19714), .B(n11851), .Z(n11339) );
  NANDN U11513 ( .A(n11339), .B(n19766), .Z(n11241) );
  NANDN U11514 ( .A(n11239), .B(n19767), .Z(n11240) );
  NAND U11515 ( .A(n11241), .B(n11240), .Z(n11318) );
  NAND U11516 ( .A(n19554), .B(n11242), .Z(n11244) );
  IV U11517 ( .A(a[149]), .Z(n12163) );
  XNOR U11518 ( .A(b[3]), .B(n12163), .Z(n11342) );
  NANDN U11519 ( .A(n19521), .B(n11342), .Z(n11243) );
  AND U11520 ( .A(n11244), .B(n11243), .Z(n11319) );
  XNOR U11521 ( .A(n11318), .B(n11319), .Z(n11320) );
  XOR U11522 ( .A(n11321), .B(n11320), .Z(n11346) );
  XOR U11523 ( .A(n11345), .B(n11346), .Z(n11347) );
  XNOR U11524 ( .A(n11348), .B(n11347), .Z(n11296) );
  NAND U11525 ( .A(n11246), .B(n11245), .Z(n11250) );
  NAND U11526 ( .A(n11248), .B(n11247), .Z(n11249) );
  NAND U11527 ( .A(n11250), .B(n11249), .Z(n11297) );
  XOR U11528 ( .A(n11296), .B(n11297), .Z(n11299) );
  XNOR U11529 ( .A(n20052), .B(n11539), .Z(n11302) );
  OR U11530 ( .A(n11302), .B(n20020), .Z(n11253) );
  NANDN U11531 ( .A(n11251), .B(n19960), .Z(n11252) );
  NAND U11532 ( .A(n11253), .B(n11252), .Z(n11315) );
  XNOR U11533 ( .A(n102), .B(n11254), .Z(n11306) );
  OR U11534 ( .A(n11306), .B(n20121), .Z(n11257) );
  NANDN U11535 ( .A(n11255), .B(n20122), .Z(n11256) );
  NAND U11536 ( .A(n11257), .B(n11256), .Z(n11312) );
  XNOR U11537 ( .A(n19975), .B(n11722), .Z(n11309) );
  NANDN U11538 ( .A(n11309), .B(n19883), .Z(n11260) );
  NANDN U11539 ( .A(n11258), .B(n19937), .Z(n11259) );
  AND U11540 ( .A(n11260), .B(n11259), .Z(n11313) );
  XNOR U11541 ( .A(n11312), .B(n11313), .Z(n11314) );
  XNOR U11542 ( .A(n11315), .B(n11314), .Z(n11351) );
  NANDN U11543 ( .A(n11262), .B(n11261), .Z(n11266) );
  NAND U11544 ( .A(n11264), .B(n11263), .Z(n11265) );
  NAND U11545 ( .A(n11266), .B(n11265), .Z(n11352) );
  XNOR U11546 ( .A(n11351), .B(n11352), .Z(n11353) );
  NANDN U11547 ( .A(n11268), .B(n11267), .Z(n11272) );
  NAND U11548 ( .A(n11270), .B(n11269), .Z(n11271) );
  AND U11549 ( .A(n11272), .B(n11271), .Z(n11354) );
  XNOR U11550 ( .A(n11353), .B(n11354), .Z(n11298) );
  XNOR U11551 ( .A(n11299), .B(n11298), .Z(n11357) );
  NANDN U11552 ( .A(n11274), .B(n11273), .Z(n11278) );
  NAND U11553 ( .A(n11276), .B(n11275), .Z(n11277) );
  NAND U11554 ( .A(n11278), .B(n11277), .Z(n11358) );
  XNOR U11555 ( .A(n11357), .B(n11358), .Z(n11359) );
  XOR U11556 ( .A(n11360), .B(n11359), .Z(n11290) );
  NANDN U11557 ( .A(n11280), .B(n11279), .Z(n11284) );
  NANDN U11558 ( .A(n11282), .B(n11281), .Z(n11283) );
  NAND U11559 ( .A(n11284), .B(n11283), .Z(n11291) );
  XNOR U11560 ( .A(n11290), .B(n11291), .Z(n11292) );
  XNOR U11561 ( .A(n11293), .B(n11292), .Z(n11363) );
  XNOR U11562 ( .A(n11363), .B(sreg[391]), .Z(n11365) );
  NAND U11563 ( .A(n11285), .B(sreg[390]), .Z(n11289) );
  OR U11564 ( .A(n11287), .B(n11286), .Z(n11288) );
  AND U11565 ( .A(n11289), .B(n11288), .Z(n11364) );
  XOR U11566 ( .A(n11365), .B(n11364), .Z(c[391]) );
  NANDN U11567 ( .A(n11291), .B(n11290), .Z(n11295) );
  NAND U11568 ( .A(n11293), .B(n11292), .Z(n11294) );
  NAND U11569 ( .A(n11295), .B(n11294), .Z(n11371) );
  NANDN U11570 ( .A(n11297), .B(n11296), .Z(n11301) );
  OR U11571 ( .A(n11299), .B(n11298), .Z(n11300) );
  NAND U11572 ( .A(n11301), .B(n11300), .Z(n11438) );
  XNOR U11573 ( .A(n20052), .B(n11644), .Z(n11407) );
  OR U11574 ( .A(n11407), .B(n20020), .Z(n11304) );
  NANDN U11575 ( .A(n11302), .B(n19960), .Z(n11303) );
  NAND U11576 ( .A(n11304), .B(n11303), .Z(n11420) );
  XNOR U11577 ( .A(n102), .B(n11305), .Z(n11411) );
  OR U11578 ( .A(n11411), .B(n20121), .Z(n11308) );
  NANDN U11579 ( .A(n11306), .B(n20122), .Z(n11307) );
  NAND U11580 ( .A(n11308), .B(n11307), .Z(n11417) );
  XNOR U11581 ( .A(n19975), .B(n11773), .Z(n11414) );
  NANDN U11582 ( .A(n11414), .B(n19883), .Z(n11311) );
  NANDN U11583 ( .A(n11309), .B(n19937), .Z(n11310) );
  AND U11584 ( .A(n11311), .B(n11310), .Z(n11418) );
  XNOR U11585 ( .A(n11417), .B(n11418), .Z(n11419) );
  XNOR U11586 ( .A(n11420), .B(n11419), .Z(n11429) );
  NANDN U11587 ( .A(n11313), .B(n11312), .Z(n11317) );
  NAND U11588 ( .A(n11315), .B(n11314), .Z(n11316) );
  NAND U11589 ( .A(n11317), .B(n11316), .Z(n11430) );
  XNOR U11590 ( .A(n11429), .B(n11430), .Z(n11431) );
  NANDN U11591 ( .A(n11319), .B(n11318), .Z(n11323) );
  NAND U11592 ( .A(n11321), .B(n11320), .Z(n11322) );
  AND U11593 ( .A(n11323), .B(n11322), .Z(n11432) );
  XNOR U11594 ( .A(n11431), .B(n11432), .Z(n11376) );
  NANDN U11595 ( .A(n11325), .B(n11324), .Z(n11329) );
  OR U11596 ( .A(n11327), .B(n11326), .Z(n11328) );
  NAND U11597 ( .A(n11329), .B(n11328), .Z(n11404) );
  NAND U11598 ( .A(b[0]), .B(a[152]), .Z(n11330) );
  XNOR U11599 ( .A(b[1]), .B(n11330), .Z(n11332) );
  NAND U11600 ( .A(a[151]), .B(n98), .Z(n11331) );
  AND U11601 ( .A(n11332), .B(n11331), .Z(n11380) );
  XNOR U11602 ( .A(n20154), .B(n11461), .Z(n11389) );
  OR U11603 ( .A(n11389), .B(n20057), .Z(n11335) );
  NANDN U11604 ( .A(n11333), .B(n20098), .Z(n11334) );
  AND U11605 ( .A(n11335), .B(n11334), .Z(n11381) );
  XOR U11606 ( .A(n11380), .B(n11381), .Z(n11383) );
  NAND U11607 ( .A(a[136]), .B(b[15]), .Z(n11382) );
  XOR U11608 ( .A(n11383), .B(n11382), .Z(n11401) );
  NAND U11609 ( .A(n19722), .B(n11336), .Z(n11338) );
  XNOR U11610 ( .A(b[5]), .B(n12112), .Z(n11392) );
  NANDN U11611 ( .A(n19640), .B(n11392), .Z(n11337) );
  NAND U11612 ( .A(n11338), .B(n11337), .Z(n11426) );
  XNOR U11613 ( .A(n19714), .B(n11929), .Z(n11395) );
  NANDN U11614 ( .A(n11395), .B(n19766), .Z(n11341) );
  NANDN U11615 ( .A(n11339), .B(n19767), .Z(n11340) );
  NAND U11616 ( .A(n11341), .B(n11340), .Z(n11423) );
  NAND U11617 ( .A(n19554), .B(n11342), .Z(n11344) );
  IV U11618 ( .A(a[150]), .Z(n12241) );
  XNOR U11619 ( .A(b[3]), .B(n12241), .Z(n11398) );
  NANDN U11620 ( .A(n19521), .B(n11398), .Z(n11343) );
  AND U11621 ( .A(n11344), .B(n11343), .Z(n11424) );
  XNOR U11622 ( .A(n11423), .B(n11424), .Z(n11425) );
  XOR U11623 ( .A(n11426), .B(n11425), .Z(n11402) );
  XOR U11624 ( .A(n11401), .B(n11402), .Z(n11403) );
  XNOR U11625 ( .A(n11404), .B(n11403), .Z(n11374) );
  NAND U11626 ( .A(n11346), .B(n11345), .Z(n11350) );
  NAND U11627 ( .A(n11348), .B(n11347), .Z(n11349) );
  NAND U11628 ( .A(n11350), .B(n11349), .Z(n11375) );
  XOR U11629 ( .A(n11374), .B(n11375), .Z(n11377) );
  XNOR U11630 ( .A(n11376), .B(n11377), .Z(n11435) );
  NANDN U11631 ( .A(n11352), .B(n11351), .Z(n11356) );
  NAND U11632 ( .A(n11354), .B(n11353), .Z(n11355) );
  NAND U11633 ( .A(n11356), .B(n11355), .Z(n11436) );
  XNOR U11634 ( .A(n11435), .B(n11436), .Z(n11437) );
  XOR U11635 ( .A(n11438), .B(n11437), .Z(n11368) );
  NANDN U11636 ( .A(n11358), .B(n11357), .Z(n11362) );
  NANDN U11637 ( .A(n11360), .B(n11359), .Z(n11361) );
  NAND U11638 ( .A(n11362), .B(n11361), .Z(n11369) );
  XNOR U11639 ( .A(n11368), .B(n11369), .Z(n11370) );
  XNOR U11640 ( .A(n11371), .B(n11370), .Z(n11441) );
  XNOR U11641 ( .A(n11441), .B(sreg[392]), .Z(n11443) );
  NAND U11642 ( .A(n11363), .B(sreg[391]), .Z(n11367) );
  OR U11643 ( .A(n11365), .B(n11364), .Z(n11366) );
  AND U11644 ( .A(n11367), .B(n11366), .Z(n11442) );
  XOR U11645 ( .A(n11443), .B(n11442), .Z(c[392]) );
  NANDN U11646 ( .A(n11369), .B(n11368), .Z(n11373) );
  NAND U11647 ( .A(n11371), .B(n11370), .Z(n11372) );
  NAND U11648 ( .A(n11373), .B(n11372), .Z(n11449) );
  NANDN U11649 ( .A(n11375), .B(n11374), .Z(n11379) );
  OR U11650 ( .A(n11377), .B(n11376), .Z(n11378) );
  NAND U11651 ( .A(n11379), .B(n11378), .Z(n11516) );
  NANDN U11652 ( .A(n11381), .B(n11380), .Z(n11385) );
  OR U11653 ( .A(n11383), .B(n11382), .Z(n11384) );
  NAND U11654 ( .A(n11385), .B(n11384), .Z(n11504) );
  NAND U11655 ( .A(b[0]), .B(a[153]), .Z(n11386) );
  XNOR U11656 ( .A(b[1]), .B(n11386), .Z(n11388) );
  NAND U11657 ( .A(a[152]), .B(n98), .Z(n11387) );
  AND U11658 ( .A(n11388), .B(n11387), .Z(n11480) );
  XNOR U11659 ( .A(n20154), .B(n11539), .Z(n11486) );
  OR U11660 ( .A(n11486), .B(n20057), .Z(n11391) );
  NANDN U11661 ( .A(n11389), .B(n20098), .Z(n11390) );
  AND U11662 ( .A(n11391), .B(n11390), .Z(n11481) );
  XOR U11663 ( .A(n11480), .B(n11481), .Z(n11483) );
  NAND U11664 ( .A(a[137]), .B(b[15]), .Z(n11482) );
  XOR U11665 ( .A(n11483), .B(n11482), .Z(n11501) );
  NAND U11666 ( .A(n19722), .B(n11392), .Z(n11394) );
  XNOR U11667 ( .A(b[5]), .B(n12163), .Z(n11492) );
  NANDN U11668 ( .A(n19640), .B(n11492), .Z(n11393) );
  NAND U11669 ( .A(n11394), .B(n11393), .Z(n11477) );
  XNOR U11670 ( .A(n19714), .B(n12007), .Z(n11495) );
  NANDN U11671 ( .A(n11495), .B(n19766), .Z(n11397) );
  NANDN U11672 ( .A(n11395), .B(n19767), .Z(n11396) );
  NAND U11673 ( .A(n11397), .B(n11396), .Z(n11474) );
  NAND U11674 ( .A(n19554), .B(n11398), .Z(n11400) );
  IV U11675 ( .A(a[151]), .Z(n12346) );
  XNOR U11676 ( .A(b[3]), .B(n12346), .Z(n11498) );
  NANDN U11677 ( .A(n19521), .B(n11498), .Z(n11399) );
  AND U11678 ( .A(n11400), .B(n11399), .Z(n11475) );
  XNOR U11679 ( .A(n11474), .B(n11475), .Z(n11476) );
  XOR U11680 ( .A(n11477), .B(n11476), .Z(n11502) );
  XOR U11681 ( .A(n11501), .B(n11502), .Z(n11503) );
  XNOR U11682 ( .A(n11504), .B(n11503), .Z(n11452) );
  NAND U11683 ( .A(n11402), .B(n11401), .Z(n11406) );
  NAND U11684 ( .A(n11404), .B(n11403), .Z(n11405) );
  NAND U11685 ( .A(n11406), .B(n11405), .Z(n11453) );
  XOR U11686 ( .A(n11452), .B(n11453), .Z(n11455) );
  XNOR U11687 ( .A(n20052), .B(n11722), .Z(n11458) );
  OR U11688 ( .A(n11458), .B(n20020), .Z(n11409) );
  NANDN U11689 ( .A(n11407), .B(n19960), .Z(n11408) );
  NAND U11690 ( .A(n11409), .B(n11408), .Z(n11471) );
  XNOR U11691 ( .A(n102), .B(n11410), .Z(n11462) );
  OR U11692 ( .A(n11462), .B(n20121), .Z(n11413) );
  NANDN U11693 ( .A(n11411), .B(n20122), .Z(n11412) );
  NAND U11694 ( .A(n11413), .B(n11412), .Z(n11468) );
  XNOR U11695 ( .A(n19975), .B(n11851), .Z(n11465) );
  NANDN U11696 ( .A(n11465), .B(n19883), .Z(n11416) );
  NANDN U11697 ( .A(n11414), .B(n19937), .Z(n11415) );
  AND U11698 ( .A(n11416), .B(n11415), .Z(n11469) );
  XNOR U11699 ( .A(n11468), .B(n11469), .Z(n11470) );
  XNOR U11700 ( .A(n11471), .B(n11470), .Z(n11507) );
  NANDN U11701 ( .A(n11418), .B(n11417), .Z(n11422) );
  NAND U11702 ( .A(n11420), .B(n11419), .Z(n11421) );
  NAND U11703 ( .A(n11422), .B(n11421), .Z(n11508) );
  XNOR U11704 ( .A(n11507), .B(n11508), .Z(n11509) );
  NANDN U11705 ( .A(n11424), .B(n11423), .Z(n11428) );
  NAND U11706 ( .A(n11426), .B(n11425), .Z(n11427) );
  AND U11707 ( .A(n11428), .B(n11427), .Z(n11510) );
  XNOR U11708 ( .A(n11509), .B(n11510), .Z(n11454) );
  XNOR U11709 ( .A(n11455), .B(n11454), .Z(n11513) );
  NANDN U11710 ( .A(n11430), .B(n11429), .Z(n11434) );
  NAND U11711 ( .A(n11432), .B(n11431), .Z(n11433) );
  NAND U11712 ( .A(n11434), .B(n11433), .Z(n11514) );
  XNOR U11713 ( .A(n11513), .B(n11514), .Z(n11515) );
  XOR U11714 ( .A(n11516), .B(n11515), .Z(n11446) );
  NANDN U11715 ( .A(n11436), .B(n11435), .Z(n11440) );
  NANDN U11716 ( .A(n11438), .B(n11437), .Z(n11439) );
  NAND U11717 ( .A(n11440), .B(n11439), .Z(n11447) );
  XNOR U11718 ( .A(n11446), .B(n11447), .Z(n11448) );
  XNOR U11719 ( .A(n11449), .B(n11448), .Z(n11519) );
  XNOR U11720 ( .A(n11519), .B(sreg[393]), .Z(n11521) );
  NAND U11721 ( .A(n11441), .B(sreg[392]), .Z(n11445) );
  OR U11722 ( .A(n11443), .B(n11442), .Z(n11444) );
  AND U11723 ( .A(n11445), .B(n11444), .Z(n11520) );
  XOR U11724 ( .A(n11521), .B(n11520), .Z(c[393]) );
  NANDN U11725 ( .A(n11447), .B(n11446), .Z(n11451) );
  NAND U11726 ( .A(n11449), .B(n11448), .Z(n11450) );
  NAND U11727 ( .A(n11451), .B(n11450), .Z(n11527) );
  NANDN U11728 ( .A(n11453), .B(n11452), .Z(n11457) );
  OR U11729 ( .A(n11455), .B(n11454), .Z(n11456) );
  NAND U11730 ( .A(n11457), .B(n11456), .Z(n11594) );
  XNOR U11731 ( .A(n20052), .B(n11773), .Z(n11536) );
  OR U11732 ( .A(n11536), .B(n20020), .Z(n11460) );
  NANDN U11733 ( .A(n11458), .B(n19960), .Z(n11459) );
  NAND U11734 ( .A(n11460), .B(n11459), .Z(n11549) );
  XNOR U11735 ( .A(n102), .B(n11461), .Z(n11540) );
  OR U11736 ( .A(n11540), .B(n20121), .Z(n11464) );
  NANDN U11737 ( .A(n11462), .B(n20122), .Z(n11463) );
  NAND U11738 ( .A(n11464), .B(n11463), .Z(n11546) );
  XNOR U11739 ( .A(n19975), .B(n11929), .Z(n11543) );
  NANDN U11740 ( .A(n11543), .B(n19883), .Z(n11467) );
  NANDN U11741 ( .A(n11465), .B(n19937), .Z(n11466) );
  AND U11742 ( .A(n11467), .B(n11466), .Z(n11547) );
  XNOR U11743 ( .A(n11546), .B(n11547), .Z(n11548) );
  XNOR U11744 ( .A(n11549), .B(n11548), .Z(n11585) );
  NANDN U11745 ( .A(n11469), .B(n11468), .Z(n11473) );
  NAND U11746 ( .A(n11471), .B(n11470), .Z(n11472) );
  NAND U11747 ( .A(n11473), .B(n11472), .Z(n11586) );
  XNOR U11748 ( .A(n11585), .B(n11586), .Z(n11587) );
  NANDN U11749 ( .A(n11475), .B(n11474), .Z(n11479) );
  NAND U11750 ( .A(n11477), .B(n11476), .Z(n11478) );
  AND U11751 ( .A(n11479), .B(n11478), .Z(n11588) );
  XNOR U11752 ( .A(n11587), .B(n11588), .Z(n11532) );
  NANDN U11753 ( .A(n11481), .B(n11480), .Z(n11485) );
  OR U11754 ( .A(n11483), .B(n11482), .Z(n11484) );
  NAND U11755 ( .A(n11485), .B(n11484), .Z(n11582) );
  XNOR U11756 ( .A(n20154), .B(n11644), .Z(n11567) );
  OR U11757 ( .A(n11567), .B(n20057), .Z(n11488) );
  NANDN U11758 ( .A(n11486), .B(n20098), .Z(n11487) );
  AND U11759 ( .A(n11488), .B(n11487), .Z(n11559) );
  NAND U11760 ( .A(b[0]), .B(a[154]), .Z(n11489) );
  XNOR U11761 ( .A(b[1]), .B(n11489), .Z(n11491) );
  NAND U11762 ( .A(a[153]), .B(n98), .Z(n11490) );
  AND U11763 ( .A(n11491), .B(n11490), .Z(n11558) );
  XOR U11764 ( .A(n11559), .B(n11558), .Z(n11561) );
  NAND U11765 ( .A(a[138]), .B(b[15]), .Z(n11560) );
  XOR U11766 ( .A(n11561), .B(n11560), .Z(n11579) );
  NAND U11767 ( .A(n19722), .B(n11492), .Z(n11494) );
  XNOR U11768 ( .A(b[5]), .B(n12241), .Z(n11570) );
  NANDN U11769 ( .A(n19640), .B(n11570), .Z(n11493) );
  NAND U11770 ( .A(n11494), .B(n11493), .Z(n11555) );
  XNOR U11771 ( .A(n19714), .B(n12112), .Z(n11573) );
  NANDN U11772 ( .A(n11573), .B(n19766), .Z(n11497) );
  NANDN U11773 ( .A(n11495), .B(n19767), .Z(n11496) );
  NAND U11774 ( .A(n11497), .B(n11496), .Z(n11552) );
  NAND U11775 ( .A(n19554), .B(n11498), .Z(n11500) );
  IV U11776 ( .A(a[152]), .Z(n12397) );
  XNOR U11777 ( .A(b[3]), .B(n12397), .Z(n11576) );
  NANDN U11778 ( .A(n19521), .B(n11576), .Z(n11499) );
  AND U11779 ( .A(n11500), .B(n11499), .Z(n11553) );
  XNOR U11780 ( .A(n11552), .B(n11553), .Z(n11554) );
  XOR U11781 ( .A(n11555), .B(n11554), .Z(n11580) );
  XOR U11782 ( .A(n11579), .B(n11580), .Z(n11581) );
  XNOR U11783 ( .A(n11582), .B(n11581), .Z(n11530) );
  NAND U11784 ( .A(n11502), .B(n11501), .Z(n11506) );
  NAND U11785 ( .A(n11504), .B(n11503), .Z(n11505) );
  NAND U11786 ( .A(n11506), .B(n11505), .Z(n11531) );
  XOR U11787 ( .A(n11530), .B(n11531), .Z(n11533) );
  XNOR U11788 ( .A(n11532), .B(n11533), .Z(n11591) );
  NANDN U11789 ( .A(n11508), .B(n11507), .Z(n11512) );
  NAND U11790 ( .A(n11510), .B(n11509), .Z(n11511) );
  NAND U11791 ( .A(n11512), .B(n11511), .Z(n11592) );
  XNOR U11792 ( .A(n11591), .B(n11592), .Z(n11593) );
  XOR U11793 ( .A(n11594), .B(n11593), .Z(n11524) );
  NANDN U11794 ( .A(n11514), .B(n11513), .Z(n11518) );
  NANDN U11795 ( .A(n11516), .B(n11515), .Z(n11517) );
  NAND U11796 ( .A(n11518), .B(n11517), .Z(n11525) );
  XNOR U11797 ( .A(n11524), .B(n11525), .Z(n11526) );
  XNOR U11798 ( .A(n11527), .B(n11526), .Z(n11597) );
  XNOR U11799 ( .A(n11597), .B(sreg[394]), .Z(n11599) );
  NAND U11800 ( .A(n11519), .B(sreg[393]), .Z(n11523) );
  OR U11801 ( .A(n11521), .B(n11520), .Z(n11522) );
  AND U11802 ( .A(n11523), .B(n11522), .Z(n11598) );
  XOR U11803 ( .A(n11599), .B(n11598), .Z(c[394]) );
  NANDN U11804 ( .A(n11525), .B(n11524), .Z(n11529) );
  NAND U11805 ( .A(n11527), .B(n11526), .Z(n11528) );
  NAND U11806 ( .A(n11529), .B(n11528), .Z(n11605) );
  NANDN U11807 ( .A(n11531), .B(n11530), .Z(n11535) );
  OR U11808 ( .A(n11533), .B(n11532), .Z(n11534) );
  NAND U11809 ( .A(n11535), .B(n11534), .Z(n11672) );
  XNOR U11810 ( .A(n20052), .B(n11851), .Z(n11641) );
  OR U11811 ( .A(n11641), .B(n20020), .Z(n11538) );
  NANDN U11812 ( .A(n11536), .B(n19960), .Z(n11537) );
  NAND U11813 ( .A(n11538), .B(n11537), .Z(n11654) );
  XNOR U11814 ( .A(n102), .B(n11539), .Z(n11645) );
  OR U11815 ( .A(n11645), .B(n20121), .Z(n11542) );
  NANDN U11816 ( .A(n11540), .B(n20122), .Z(n11541) );
  NAND U11817 ( .A(n11542), .B(n11541), .Z(n11651) );
  XNOR U11818 ( .A(n19975), .B(n12007), .Z(n11648) );
  NANDN U11819 ( .A(n11648), .B(n19883), .Z(n11545) );
  NANDN U11820 ( .A(n11543), .B(n19937), .Z(n11544) );
  AND U11821 ( .A(n11545), .B(n11544), .Z(n11652) );
  XNOR U11822 ( .A(n11651), .B(n11652), .Z(n11653) );
  XNOR U11823 ( .A(n11654), .B(n11653), .Z(n11663) );
  NANDN U11824 ( .A(n11547), .B(n11546), .Z(n11551) );
  NAND U11825 ( .A(n11549), .B(n11548), .Z(n11550) );
  NAND U11826 ( .A(n11551), .B(n11550), .Z(n11664) );
  XNOR U11827 ( .A(n11663), .B(n11664), .Z(n11665) );
  NANDN U11828 ( .A(n11553), .B(n11552), .Z(n11557) );
  NAND U11829 ( .A(n11555), .B(n11554), .Z(n11556) );
  AND U11830 ( .A(n11557), .B(n11556), .Z(n11666) );
  XNOR U11831 ( .A(n11665), .B(n11666), .Z(n11610) );
  NANDN U11832 ( .A(n11559), .B(n11558), .Z(n11563) );
  OR U11833 ( .A(n11561), .B(n11560), .Z(n11562) );
  NAND U11834 ( .A(n11563), .B(n11562), .Z(n11638) );
  NAND U11835 ( .A(b[0]), .B(a[155]), .Z(n11564) );
  XNOR U11836 ( .A(b[1]), .B(n11564), .Z(n11566) );
  NAND U11837 ( .A(a[154]), .B(n98), .Z(n11565) );
  AND U11838 ( .A(n11566), .B(n11565), .Z(n11614) );
  XNOR U11839 ( .A(n20154), .B(n11722), .Z(n11620) );
  OR U11840 ( .A(n11620), .B(n20057), .Z(n11569) );
  NANDN U11841 ( .A(n11567), .B(n20098), .Z(n11568) );
  AND U11842 ( .A(n11569), .B(n11568), .Z(n11615) );
  XOR U11843 ( .A(n11614), .B(n11615), .Z(n11617) );
  NAND U11844 ( .A(a[139]), .B(b[15]), .Z(n11616) );
  XOR U11845 ( .A(n11617), .B(n11616), .Z(n11635) );
  NAND U11846 ( .A(n19722), .B(n11570), .Z(n11572) );
  XNOR U11847 ( .A(b[5]), .B(n12346), .Z(n11626) );
  NANDN U11848 ( .A(n19640), .B(n11626), .Z(n11571) );
  NAND U11849 ( .A(n11572), .B(n11571), .Z(n11660) );
  XNOR U11850 ( .A(n19714), .B(n12163), .Z(n11629) );
  NANDN U11851 ( .A(n11629), .B(n19766), .Z(n11575) );
  NANDN U11852 ( .A(n11573), .B(n19767), .Z(n11574) );
  NAND U11853 ( .A(n11575), .B(n11574), .Z(n11657) );
  NAND U11854 ( .A(n19554), .B(n11576), .Z(n11578) );
  IV U11855 ( .A(a[153]), .Z(n12475) );
  XNOR U11856 ( .A(b[3]), .B(n12475), .Z(n11632) );
  NANDN U11857 ( .A(n19521), .B(n11632), .Z(n11577) );
  AND U11858 ( .A(n11578), .B(n11577), .Z(n11658) );
  XNOR U11859 ( .A(n11657), .B(n11658), .Z(n11659) );
  XOR U11860 ( .A(n11660), .B(n11659), .Z(n11636) );
  XOR U11861 ( .A(n11635), .B(n11636), .Z(n11637) );
  XNOR U11862 ( .A(n11638), .B(n11637), .Z(n11608) );
  NAND U11863 ( .A(n11580), .B(n11579), .Z(n11584) );
  NAND U11864 ( .A(n11582), .B(n11581), .Z(n11583) );
  NAND U11865 ( .A(n11584), .B(n11583), .Z(n11609) );
  XOR U11866 ( .A(n11608), .B(n11609), .Z(n11611) );
  XNOR U11867 ( .A(n11610), .B(n11611), .Z(n11669) );
  NANDN U11868 ( .A(n11586), .B(n11585), .Z(n11590) );
  NAND U11869 ( .A(n11588), .B(n11587), .Z(n11589) );
  NAND U11870 ( .A(n11590), .B(n11589), .Z(n11670) );
  XNOR U11871 ( .A(n11669), .B(n11670), .Z(n11671) );
  XOR U11872 ( .A(n11672), .B(n11671), .Z(n11602) );
  NANDN U11873 ( .A(n11592), .B(n11591), .Z(n11596) );
  NANDN U11874 ( .A(n11594), .B(n11593), .Z(n11595) );
  NAND U11875 ( .A(n11596), .B(n11595), .Z(n11603) );
  XNOR U11876 ( .A(n11602), .B(n11603), .Z(n11604) );
  XNOR U11877 ( .A(n11605), .B(n11604), .Z(n11675) );
  XNOR U11878 ( .A(n11675), .B(sreg[395]), .Z(n11677) );
  NAND U11879 ( .A(n11597), .B(sreg[394]), .Z(n11601) );
  OR U11880 ( .A(n11599), .B(n11598), .Z(n11600) );
  AND U11881 ( .A(n11601), .B(n11600), .Z(n11676) );
  XOR U11882 ( .A(n11677), .B(n11676), .Z(c[395]) );
  NANDN U11883 ( .A(n11603), .B(n11602), .Z(n11607) );
  NAND U11884 ( .A(n11605), .B(n11604), .Z(n11606) );
  NAND U11885 ( .A(n11607), .B(n11606), .Z(n11683) );
  NANDN U11886 ( .A(n11609), .B(n11608), .Z(n11613) );
  OR U11887 ( .A(n11611), .B(n11610), .Z(n11612) );
  NAND U11888 ( .A(n11613), .B(n11612), .Z(n11750) );
  NANDN U11889 ( .A(n11615), .B(n11614), .Z(n11619) );
  OR U11890 ( .A(n11617), .B(n11616), .Z(n11618) );
  NAND U11891 ( .A(n11619), .B(n11618), .Z(n11716) );
  XNOR U11892 ( .A(n20154), .B(n11773), .Z(n11701) );
  OR U11893 ( .A(n11701), .B(n20057), .Z(n11622) );
  NANDN U11894 ( .A(n11620), .B(n20098), .Z(n11621) );
  AND U11895 ( .A(n11622), .B(n11621), .Z(n11693) );
  NAND U11896 ( .A(b[0]), .B(a[156]), .Z(n11623) );
  XNOR U11897 ( .A(b[1]), .B(n11623), .Z(n11625) );
  NAND U11898 ( .A(a[155]), .B(n98), .Z(n11624) );
  AND U11899 ( .A(n11625), .B(n11624), .Z(n11692) );
  XOR U11900 ( .A(n11693), .B(n11692), .Z(n11695) );
  NAND U11901 ( .A(a[140]), .B(b[15]), .Z(n11694) );
  XOR U11902 ( .A(n11695), .B(n11694), .Z(n11713) );
  NAND U11903 ( .A(n19722), .B(n11626), .Z(n11628) );
  XNOR U11904 ( .A(b[5]), .B(n12397), .Z(n11704) );
  NANDN U11905 ( .A(n19640), .B(n11704), .Z(n11627) );
  NAND U11906 ( .A(n11628), .B(n11627), .Z(n11738) );
  XNOR U11907 ( .A(n19714), .B(n12241), .Z(n11707) );
  NANDN U11908 ( .A(n11707), .B(n19766), .Z(n11631) );
  NANDN U11909 ( .A(n11629), .B(n19767), .Z(n11630) );
  NAND U11910 ( .A(n11631), .B(n11630), .Z(n11735) );
  NAND U11911 ( .A(n19554), .B(n11632), .Z(n11634) );
  IV U11912 ( .A(a[154]), .Z(n12580) );
  XNOR U11913 ( .A(b[3]), .B(n12580), .Z(n11710) );
  NANDN U11914 ( .A(n19521), .B(n11710), .Z(n11633) );
  AND U11915 ( .A(n11634), .B(n11633), .Z(n11736) );
  XNOR U11916 ( .A(n11735), .B(n11736), .Z(n11737) );
  XOR U11917 ( .A(n11738), .B(n11737), .Z(n11714) );
  XOR U11918 ( .A(n11713), .B(n11714), .Z(n11715) );
  XNOR U11919 ( .A(n11716), .B(n11715), .Z(n11686) );
  NAND U11920 ( .A(n11636), .B(n11635), .Z(n11640) );
  NAND U11921 ( .A(n11638), .B(n11637), .Z(n11639) );
  NAND U11922 ( .A(n11640), .B(n11639), .Z(n11687) );
  XOR U11923 ( .A(n11686), .B(n11687), .Z(n11689) );
  XNOR U11924 ( .A(n20052), .B(n11929), .Z(n11719) );
  OR U11925 ( .A(n11719), .B(n20020), .Z(n11643) );
  NANDN U11926 ( .A(n11641), .B(n19960), .Z(n11642) );
  NAND U11927 ( .A(n11643), .B(n11642), .Z(n11732) );
  XNOR U11928 ( .A(n102), .B(n11644), .Z(n11723) );
  OR U11929 ( .A(n11723), .B(n20121), .Z(n11647) );
  NANDN U11930 ( .A(n11645), .B(n20122), .Z(n11646) );
  NAND U11931 ( .A(n11647), .B(n11646), .Z(n11729) );
  XNOR U11932 ( .A(n19975), .B(n12112), .Z(n11726) );
  NANDN U11933 ( .A(n11726), .B(n19883), .Z(n11650) );
  NANDN U11934 ( .A(n11648), .B(n19937), .Z(n11649) );
  AND U11935 ( .A(n11650), .B(n11649), .Z(n11730) );
  XNOR U11936 ( .A(n11729), .B(n11730), .Z(n11731) );
  XNOR U11937 ( .A(n11732), .B(n11731), .Z(n11741) );
  NANDN U11938 ( .A(n11652), .B(n11651), .Z(n11656) );
  NAND U11939 ( .A(n11654), .B(n11653), .Z(n11655) );
  NAND U11940 ( .A(n11656), .B(n11655), .Z(n11742) );
  XNOR U11941 ( .A(n11741), .B(n11742), .Z(n11743) );
  NANDN U11942 ( .A(n11658), .B(n11657), .Z(n11662) );
  NAND U11943 ( .A(n11660), .B(n11659), .Z(n11661) );
  AND U11944 ( .A(n11662), .B(n11661), .Z(n11744) );
  XNOR U11945 ( .A(n11743), .B(n11744), .Z(n11688) );
  XNOR U11946 ( .A(n11689), .B(n11688), .Z(n11747) );
  NANDN U11947 ( .A(n11664), .B(n11663), .Z(n11668) );
  NAND U11948 ( .A(n11666), .B(n11665), .Z(n11667) );
  NAND U11949 ( .A(n11668), .B(n11667), .Z(n11748) );
  XNOR U11950 ( .A(n11747), .B(n11748), .Z(n11749) );
  XOR U11951 ( .A(n11750), .B(n11749), .Z(n11680) );
  NANDN U11952 ( .A(n11670), .B(n11669), .Z(n11674) );
  NANDN U11953 ( .A(n11672), .B(n11671), .Z(n11673) );
  NAND U11954 ( .A(n11674), .B(n11673), .Z(n11681) );
  XNOR U11955 ( .A(n11680), .B(n11681), .Z(n11682) );
  XNOR U11956 ( .A(n11683), .B(n11682), .Z(n11753) );
  XNOR U11957 ( .A(n11753), .B(sreg[396]), .Z(n11755) );
  NAND U11958 ( .A(n11675), .B(sreg[395]), .Z(n11679) );
  OR U11959 ( .A(n11677), .B(n11676), .Z(n11678) );
  AND U11960 ( .A(n11679), .B(n11678), .Z(n11754) );
  XOR U11961 ( .A(n11755), .B(n11754), .Z(c[396]) );
  NANDN U11962 ( .A(n11681), .B(n11680), .Z(n11685) );
  NAND U11963 ( .A(n11683), .B(n11682), .Z(n11684) );
  NAND U11964 ( .A(n11685), .B(n11684), .Z(n11761) );
  NANDN U11965 ( .A(n11687), .B(n11686), .Z(n11691) );
  OR U11966 ( .A(n11689), .B(n11688), .Z(n11690) );
  NAND U11967 ( .A(n11691), .B(n11690), .Z(n11828) );
  NANDN U11968 ( .A(n11693), .B(n11692), .Z(n11697) );
  OR U11969 ( .A(n11695), .B(n11694), .Z(n11696) );
  NAND U11970 ( .A(n11697), .B(n11696), .Z(n11816) );
  NAND U11971 ( .A(b[0]), .B(a[157]), .Z(n11698) );
  XNOR U11972 ( .A(b[1]), .B(n11698), .Z(n11700) );
  NAND U11973 ( .A(a[156]), .B(n98), .Z(n11699) );
  AND U11974 ( .A(n11700), .B(n11699), .Z(n11792) );
  XNOR U11975 ( .A(n20154), .B(n11851), .Z(n11801) );
  OR U11976 ( .A(n11801), .B(n20057), .Z(n11703) );
  NANDN U11977 ( .A(n11701), .B(n20098), .Z(n11702) );
  AND U11978 ( .A(n11703), .B(n11702), .Z(n11793) );
  XOR U11979 ( .A(n11792), .B(n11793), .Z(n11795) );
  NAND U11980 ( .A(a[141]), .B(b[15]), .Z(n11794) );
  XOR U11981 ( .A(n11795), .B(n11794), .Z(n11813) );
  NAND U11982 ( .A(n19722), .B(n11704), .Z(n11706) );
  XNOR U11983 ( .A(b[5]), .B(n12475), .Z(n11804) );
  NANDN U11984 ( .A(n19640), .B(n11804), .Z(n11705) );
  NAND U11985 ( .A(n11706), .B(n11705), .Z(n11789) );
  XNOR U11986 ( .A(n19714), .B(n12346), .Z(n11807) );
  NANDN U11987 ( .A(n11807), .B(n19766), .Z(n11709) );
  NANDN U11988 ( .A(n11707), .B(n19767), .Z(n11708) );
  NAND U11989 ( .A(n11709), .B(n11708), .Z(n11786) );
  NAND U11990 ( .A(n19554), .B(n11710), .Z(n11712) );
  IV U11991 ( .A(a[155]), .Z(n12631) );
  XNOR U11992 ( .A(b[3]), .B(n12631), .Z(n11810) );
  NANDN U11993 ( .A(n19521), .B(n11810), .Z(n11711) );
  AND U11994 ( .A(n11712), .B(n11711), .Z(n11787) );
  XNOR U11995 ( .A(n11786), .B(n11787), .Z(n11788) );
  XOR U11996 ( .A(n11789), .B(n11788), .Z(n11814) );
  XOR U11997 ( .A(n11813), .B(n11814), .Z(n11815) );
  XNOR U11998 ( .A(n11816), .B(n11815), .Z(n11764) );
  NAND U11999 ( .A(n11714), .B(n11713), .Z(n11718) );
  NAND U12000 ( .A(n11716), .B(n11715), .Z(n11717) );
  NAND U12001 ( .A(n11718), .B(n11717), .Z(n11765) );
  XOR U12002 ( .A(n11764), .B(n11765), .Z(n11767) );
  XNOR U12003 ( .A(n20052), .B(n12007), .Z(n11770) );
  OR U12004 ( .A(n11770), .B(n20020), .Z(n11721) );
  NANDN U12005 ( .A(n11719), .B(n19960), .Z(n11720) );
  NAND U12006 ( .A(n11721), .B(n11720), .Z(n11783) );
  XNOR U12007 ( .A(n102), .B(n11722), .Z(n11774) );
  OR U12008 ( .A(n11774), .B(n20121), .Z(n11725) );
  NANDN U12009 ( .A(n11723), .B(n20122), .Z(n11724) );
  NAND U12010 ( .A(n11725), .B(n11724), .Z(n11780) );
  XNOR U12011 ( .A(n19975), .B(n12163), .Z(n11777) );
  NANDN U12012 ( .A(n11777), .B(n19883), .Z(n11728) );
  NANDN U12013 ( .A(n11726), .B(n19937), .Z(n11727) );
  AND U12014 ( .A(n11728), .B(n11727), .Z(n11781) );
  XNOR U12015 ( .A(n11780), .B(n11781), .Z(n11782) );
  XNOR U12016 ( .A(n11783), .B(n11782), .Z(n11819) );
  NANDN U12017 ( .A(n11730), .B(n11729), .Z(n11734) );
  NAND U12018 ( .A(n11732), .B(n11731), .Z(n11733) );
  NAND U12019 ( .A(n11734), .B(n11733), .Z(n11820) );
  XNOR U12020 ( .A(n11819), .B(n11820), .Z(n11821) );
  NANDN U12021 ( .A(n11736), .B(n11735), .Z(n11740) );
  NAND U12022 ( .A(n11738), .B(n11737), .Z(n11739) );
  AND U12023 ( .A(n11740), .B(n11739), .Z(n11822) );
  XNOR U12024 ( .A(n11821), .B(n11822), .Z(n11766) );
  XNOR U12025 ( .A(n11767), .B(n11766), .Z(n11825) );
  NANDN U12026 ( .A(n11742), .B(n11741), .Z(n11746) );
  NAND U12027 ( .A(n11744), .B(n11743), .Z(n11745) );
  NAND U12028 ( .A(n11746), .B(n11745), .Z(n11826) );
  XNOR U12029 ( .A(n11825), .B(n11826), .Z(n11827) );
  XOR U12030 ( .A(n11828), .B(n11827), .Z(n11758) );
  NANDN U12031 ( .A(n11748), .B(n11747), .Z(n11752) );
  NANDN U12032 ( .A(n11750), .B(n11749), .Z(n11751) );
  NAND U12033 ( .A(n11752), .B(n11751), .Z(n11759) );
  XNOR U12034 ( .A(n11758), .B(n11759), .Z(n11760) );
  XNOR U12035 ( .A(n11761), .B(n11760), .Z(n11831) );
  XNOR U12036 ( .A(n11831), .B(sreg[397]), .Z(n11833) );
  NAND U12037 ( .A(n11753), .B(sreg[396]), .Z(n11757) );
  OR U12038 ( .A(n11755), .B(n11754), .Z(n11756) );
  AND U12039 ( .A(n11757), .B(n11756), .Z(n11832) );
  XOR U12040 ( .A(n11833), .B(n11832), .Z(c[397]) );
  NANDN U12041 ( .A(n11759), .B(n11758), .Z(n11763) );
  NAND U12042 ( .A(n11761), .B(n11760), .Z(n11762) );
  NAND U12043 ( .A(n11763), .B(n11762), .Z(n11839) );
  NANDN U12044 ( .A(n11765), .B(n11764), .Z(n11769) );
  OR U12045 ( .A(n11767), .B(n11766), .Z(n11768) );
  NAND U12046 ( .A(n11769), .B(n11768), .Z(n11906) );
  XNOR U12047 ( .A(n20052), .B(n12112), .Z(n11848) );
  OR U12048 ( .A(n11848), .B(n20020), .Z(n11772) );
  NANDN U12049 ( .A(n11770), .B(n19960), .Z(n11771) );
  NAND U12050 ( .A(n11772), .B(n11771), .Z(n11861) );
  XNOR U12051 ( .A(n102), .B(n11773), .Z(n11852) );
  OR U12052 ( .A(n11852), .B(n20121), .Z(n11776) );
  NANDN U12053 ( .A(n11774), .B(n20122), .Z(n11775) );
  NAND U12054 ( .A(n11776), .B(n11775), .Z(n11858) );
  XNOR U12055 ( .A(n19975), .B(n12241), .Z(n11855) );
  NANDN U12056 ( .A(n11855), .B(n19883), .Z(n11779) );
  NANDN U12057 ( .A(n11777), .B(n19937), .Z(n11778) );
  AND U12058 ( .A(n11779), .B(n11778), .Z(n11859) );
  XNOR U12059 ( .A(n11858), .B(n11859), .Z(n11860) );
  XNOR U12060 ( .A(n11861), .B(n11860), .Z(n11897) );
  NANDN U12061 ( .A(n11781), .B(n11780), .Z(n11785) );
  NAND U12062 ( .A(n11783), .B(n11782), .Z(n11784) );
  NAND U12063 ( .A(n11785), .B(n11784), .Z(n11898) );
  XNOR U12064 ( .A(n11897), .B(n11898), .Z(n11899) );
  NANDN U12065 ( .A(n11787), .B(n11786), .Z(n11791) );
  NAND U12066 ( .A(n11789), .B(n11788), .Z(n11790) );
  AND U12067 ( .A(n11791), .B(n11790), .Z(n11900) );
  XNOR U12068 ( .A(n11899), .B(n11900), .Z(n11844) );
  NANDN U12069 ( .A(n11793), .B(n11792), .Z(n11797) );
  OR U12070 ( .A(n11795), .B(n11794), .Z(n11796) );
  NAND U12071 ( .A(n11797), .B(n11796), .Z(n11894) );
  NAND U12072 ( .A(b[0]), .B(a[158]), .Z(n11798) );
  XNOR U12073 ( .A(b[1]), .B(n11798), .Z(n11800) );
  NAND U12074 ( .A(a[157]), .B(n98), .Z(n11799) );
  AND U12075 ( .A(n11800), .B(n11799), .Z(n11870) );
  XNOR U12076 ( .A(n20154), .B(n11929), .Z(n11876) );
  OR U12077 ( .A(n11876), .B(n20057), .Z(n11803) );
  NANDN U12078 ( .A(n11801), .B(n20098), .Z(n11802) );
  AND U12079 ( .A(n11803), .B(n11802), .Z(n11871) );
  XOR U12080 ( .A(n11870), .B(n11871), .Z(n11873) );
  NAND U12081 ( .A(a[142]), .B(b[15]), .Z(n11872) );
  XOR U12082 ( .A(n11873), .B(n11872), .Z(n11891) );
  NAND U12083 ( .A(n19722), .B(n11804), .Z(n11806) );
  XNOR U12084 ( .A(b[5]), .B(n12580), .Z(n11882) );
  NANDN U12085 ( .A(n19640), .B(n11882), .Z(n11805) );
  NAND U12086 ( .A(n11806), .B(n11805), .Z(n11867) );
  XNOR U12087 ( .A(n19714), .B(n12397), .Z(n11885) );
  NANDN U12088 ( .A(n11885), .B(n19766), .Z(n11809) );
  NANDN U12089 ( .A(n11807), .B(n19767), .Z(n11808) );
  NAND U12090 ( .A(n11809), .B(n11808), .Z(n11864) );
  NAND U12091 ( .A(n19554), .B(n11810), .Z(n11812) );
  IV U12092 ( .A(a[156]), .Z(n12736) );
  XNOR U12093 ( .A(b[3]), .B(n12736), .Z(n11888) );
  NANDN U12094 ( .A(n19521), .B(n11888), .Z(n11811) );
  AND U12095 ( .A(n11812), .B(n11811), .Z(n11865) );
  XNOR U12096 ( .A(n11864), .B(n11865), .Z(n11866) );
  XOR U12097 ( .A(n11867), .B(n11866), .Z(n11892) );
  XOR U12098 ( .A(n11891), .B(n11892), .Z(n11893) );
  XNOR U12099 ( .A(n11894), .B(n11893), .Z(n11842) );
  NAND U12100 ( .A(n11814), .B(n11813), .Z(n11818) );
  NAND U12101 ( .A(n11816), .B(n11815), .Z(n11817) );
  NAND U12102 ( .A(n11818), .B(n11817), .Z(n11843) );
  XOR U12103 ( .A(n11842), .B(n11843), .Z(n11845) );
  XNOR U12104 ( .A(n11844), .B(n11845), .Z(n11903) );
  NANDN U12105 ( .A(n11820), .B(n11819), .Z(n11824) );
  NAND U12106 ( .A(n11822), .B(n11821), .Z(n11823) );
  NAND U12107 ( .A(n11824), .B(n11823), .Z(n11904) );
  XNOR U12108 ( .A(n11903), .B(n11904), .Z(n11905) );
  XOR U12109 ( .A(n11906), .B(n11905), .Z(n11836) );
  NANDN U12110 ( .A(n11826), .B(n11825), .Z(n11830) );
  NANDN U12111 ( .A(n11828), .B(n11827), .Z(n11829) );
  NAND U12112 ( .A(n11830), .B(n11829), .Z(n11837) );
  XNOR U12113 ( .A(n11836), .B(n11837), .Z(n11838) );
  XNOR U12114 ( .A(n11839), .B(n11838), .Z(n11909) );
  XNOR U12115 ( .A(n11909), .B(sreg[398]), .Z(n11911) );
  NAND U12116 ( .A(n11831), .B(sreg[397]), .Z(n11835) );
  OR U12117 ( .A(n11833), .B(n11832), .Z(n11834) );
  AND U12118 ( .A(n11835), .B(n11834), .Z(n11910) );
  XOR U12119 ( .A(n11911), .B(n11910), .Z(c[398]) );
  NANDN U12120 ( .A(n11837), .B(n11836), .Z(n11841) );
  NAND U12121 ( .A(n11839), .B(n11838), .Z(n11840) );
  NAND U12122 ( .A(n11841), .B(n11840), .Z(n11917) );
  NANDN U12123 ( .A(n11843), .B(n11842), .Z(n11847) );
  OR U12124 ( .A(n11845), .B(n11844), .Z(n11846) );
  NAND U12125 ( .A(n11847), .B(n11846), .Z(n11984) );
  XNOR U12126 ( .A(n20052), .B(n12163), .Z(n11926) );
  OR U12127 ( .A(n11926), .B(n20020), .Z(n11850) );
  NANDN U12128 ( .A(n11848), .B(n19960), .Z(n11849) );
  NAND U12129 ( .A(n11850), .B(n11849), .Z(n11939) );
  XNOR U12130 ( .A(n102), .B(n11851), .Z(n11930) );
  OR U12131 ( .A(n11930), .B(n20121), .Z(n11854) );
  NANDN U12132 ( .A(n11852), .B(n20122), .Z(n11853) );
  NAND U12133 ( .A(n11854), .B(n11853), .Z(n11936) );
  XNOR U12134 ( .A(n19975), .B(n12346), .Z(n11933) );
  NANDN U12135 ( .A(n11933), .B(n19883), .Z(n11857) );
  NANDN U12136 ( .A(n11855), .B(n19937), .Z(n11856) );
  AND U12137 ( .A(n11857), .B(n11856), .Z(n11937) );
  XNOR U12138 ( .A(n11936), .B(n11937), .Z(n11938) );
  XNOR U12139 ( .A(n11939), .B(n11938), .Z(n11975) );
  NANDN U12140 ( .A(n11859), .B(n11858), .Z(n11863) );
  NAND U12141 ( .A(n11861), .B(n11860), .Z(n11862) );
  NAND U12142 ( .A(n11863), .B(n11862), .Z(n11976) );
  XNOR U12143 ( .A(n11975), .B(n11976), .Z(n11977) );
  NANDN U12144 ( .A(n11865), .B(n11864), .Z(n11869) );
  NAND U12145 ( .A(n11867), .B(n11866), .Z(n11868) );
  AND U12146 ( .A(n11869), .B(n11868), .Z(n11978) );
  XNOR U12147 ( .A(n11977), .B(n11978), .Z(n11922) );
  NANDN U12148 ( .A(n11871), .B(n11870), .Z(n11875) );
  OR U12149 ( .A(n11873), .B(n11872), .Z(n11874) );
  NAND U12150 ( .A(n11875), .B(n11874), .Z(n11972) );
  XNOR U12151 ( .A(n20154), .B(n12007), .Z(n11957) );
  OR U12152 ( .A(n11957), .B(n20057), .Z(n11878) );
  NANDN U12153 ( .A(n11876), .B(n20098), .Z(n11877) );
  AND U12154 ( .A(n11878), .B(n11877), .Z(n11949) );
  NAND U12155 ( .A(b[0]), .B(a[159]), .Z(n11879) );
  XNOR U12156 ( .A(b[1]), .B(n11879), .Z(n11881) );
  NAND U12157 ( .A(a[158]), .B(n98), .Z(n11880) );
  AND U12158 ( .A(n11881), .B(n11880), .Z(n11948) );
  XOR U12159 ( .A(n11949), .B(n11948), .Z(n11951) );
  NAND U12160 ( .A(a[143]), .B(b[15]), .Z(n11950) );
  XOR U12161 ( .A(n11951), .B(n11950), .Z(n11969) );
  NAND U12162 ( .A(n19722), .B(n11882), .Z(n11884) );
  XNOR U12163 ( .A(b[5]), .B(n12631), .Z(n11960) );
  NANDN U12164 ( .A(n19640), .B(n11960), .Z(n11883) );
  NAND U12165 ( .A(n11884), .B(n11883), .Z(n11945) );
  XNOR U12166 ( .A(n19714), .B(n12475), .Z(n11963) );
  NANDN U12167 ( .A(n11963), .B(n19766), .Z(n11887) );
  NANDN U12168 ( .A(n11885), .B(n19767), .Z(n11886) );
  NAND U12169 ( .A(n11887), .B(n11886), .Z(n11942) );
  NAND U12170 ( .A(n19554), .B(n11888), .Z(n11890) );
  IV U12171 ( .A(a[157]), .Z(n12787) );
  XNOR U12172 ( .A(b[3]), .B(n12787), .Z(n11966) );
  NANDN U12173 ( .A(n19521), .B(n11966), .Z(n11889) );
  AND U12174 ( .A(n11890), .B(n11889), .Z(n11943) );
  XNOR U12175 ( .A(n11942), .B(n11943), .Z(n11944) );
  XOR U12176 ( .A(n11945), .B(n11944), .Z(n11970) );
  XOR U12177 ( .A(n11969), .B(n11970), .Z(n11971) );
  XNOR U12178 ( .A(n11972), .B(n11971), .Z(n11920) );
  NAND U12179 ( .A(n11892), .B(n11891), .Z(n11896) );
  NAND U12180 ( .A(n11894), .B(n11893), .Z(n11895) );
  NAND U12181 ( .A(n11896), .B(n11895), .Z(n11921) );
  XOR U12182 ( .A(n11920), .B(n11921), .Z(n11923) );
  XNOR U12183 ( .A(n11922), .B(n11923), .Z(n11981) );
  NANDN U12184 ( .A(n11898), .B(n11897), .Z(n11902) );
  NAND U12185 ( .A(n11900), .B(n11899), .Z(n11901) );
  NAND U12186 ( .A(n11902), .B(n11901), .Z(n11982) );
  XNOR U12187 ( .A(n11981), .B(n11982), .Z(n11983) );
  XOR U12188 ( .A(n11984), .B(n11983), .Z(n11914) );
  NANDN U12189 ( .A(n11904), .B(n11903), .Z(n11908) );
  NANDN U12190 ( .A(n11906), .B(n11905), .Z(n11907) );
  NAND U12191 ( .A(n11908), .B(n11907), .Z(n11915) );
  XNOR U12192 ( .A(n11914), .B(n11915), .Z(n11916) );
  XNOR U12193 ( .A(n11917), .B(n11916), .Z(n11987) );
  XNOR U12194 ( .A(n11987), .B(sreg[399]), .Z(n11989) );
  NAND U12195 ( .A(n11909), .B(sreg[398]), .Z(n11913) );
  OR U12196 ( .A(n11911), .B(n11910), .Z(n11912) );
  AND U12197 ( .A(n11913), .B(n11912), .Z(n11988) );
  XOR U12198 ( .A(n11989), .B(n11988), .Z(c[399]) );
  NANDN U12199 ( .A(n11915), .B(n11914), .Z(n11919) );
  NAND U12200 ( .A(n11917), .B(n11916), .Z(n11918) );
  NAND U12201 ( .A(n11919), .B(n11918), .Z(n11995) );
  NANDN U12202 ( .A(n11921), .B(n11920), .Z(n11925) );
  OR U12203 ( .A(n11923), .B(n11922), .Z(n11924) );
  NAND U12204 ( .A(n11925), .B(n11924), .Z(n12062) );
  XNOR U12205 ( .A(n20052), .B(n12241), .Z(n12004) );
  OR U12206 ( .A(n12004), .B(n20020), .Z(n11928) );
  NANDN U12207 ( .A(n11926), .B(n19960), .Z(n11927) );
  NAND U12208 ( .A(n11928), .B(n11927), .Z(n12017) );
  XNOR U12209 ( .A(n102), .B(n11929), .Z(n12008) );
  OR U12210 ( .A(n12008), .B(n20121), .Z(n11932) );
  NANDN U12211 ( .A(n11930), .B(n20122), .Z(n11931) );
  NAND U12212 ( .A(n11932), .B(n11931), .Z(n12014) );
  XNOR U12213 ( .A(n19975), .B(n12397), .Z(n12011) );
  NANDN U12214 ( .A(n12011), .B(n19883), .Z(n11935) );
  NANDN U12215 ( .A(n11933), .B(n19937), .Z(n11934) );
  AND U12216 ( .A(n11935), .B(n11934), .Z(n12015) );
  XNOR U12217 ( .A(n12014), .B(n12015), .Z(n12016) );
  XNOR U12218 ( .A(n12017), .B(n12016), .Z(n12053) );
  NANDN U12219 ( .A(n11937), .B(n11936), .Z(n11941) );
  NAND U12220 ( .A(n11939), .B(n11938), .Z(n11940) );
  NAND U12221 ( .A(n11941), .B(n11940), .Z(n12054) );
  XNOR U12222 ( .A(n12053), .B(n12054), .Z(n12055) );
  NANDN U12223 ( .A(n11943), .B(n11942), .Z(n11947) );
  NAND U12224 ( .A(n11945), .B(n11944), .Z(n11946) );
  AND U12225 ( .A(n11947), .B(n11946), .Z(n12056) );
  XNOR U12226 ( .A(n12055), .B(n12056), .Z(n12000) );
  NANDN U12227 ( .A(n11949), .B(n11948), .Z(n11953) );
  OR U12228 ( .A(n11951), .B(n11950), .Z(n11952) );
  NAND U12229 ( .A(n11953), .B(n11952), .Z(n12050) );
  NAND U12230 ( .A(b[0]), .B(a[160]), .Z(n11954) );
  XNOR U12231 ( .A(b[1]), .B(n11954), .Z(n11956) );
  NAND U12232 ( .A(a[159]), .B(n98), .Z(n11955) );
  AND U12233 ( .A(n11956), .B(n11955), .Z(n12026) );
  XNOR U12234 ( .A(n20154), .B(n12112), .Z(n12035) );
  OR U12235 ( .A(n12035), .B(n20057), .Z(n11959) );
  NANDN U12236 ( .A(n11957), .B(n20098), .Z(n11958) );
  AND U12237 ( .A(n11959), .B(n11958), .Z(n12027) );
  XOR U12238 ( .A(n12026), .B(n12027), .Z(n12029) );
  NAND U12239 ( .A(a[144]), .B(b[15]), .Z(n12028) );
  XOR U12240 ( .A(n12029), .B(n12028), .Z(n12047) );
  NAND U12241 ( .A(n19722), .B(n11960), .Z(n11962) );
  XNOR U12242 ( .A(b[5]), .B(n12736), .Z(n12038) );
  NANDN U12243 ( .A(n19640), .B(n12038), .Z(n11961) );
  NAND U12244 ( .A(n11962), .B(n11961), .Z(n12023) );
  XNOR U12245 ( .A(n19714), .B(n12580), .Z(n12041) );
  NANDN U12246 ( .A(n12041), .B(n19766), .Z(n11965) );
  NANDN U12247 ( .A(n11963), .B(n19767), .Z(n11964) );
  NAND U12248 ( .A(n11965), .B(n11964), .Z(n12020) );
  NAND U12249 ( .A(n19554), .B(n11966), .Z(n11968) );
  IV U12250 ( .A(a[158]), .Z(n12865) );
  XNOR U12251 ( .A(b[3]), .B(n12865), .Z(n12044) );
  NANDN U12252 ( .A(n19521), .B(n12044), .Z(n11967) );
  AND U12253 ( .A(n11968), .B(n11967), .Z(n12021) );
  XNOR U12254 ( .A(n12020), .B(n12021), .Z(n12022) );
  XOR U12255 ( .A(n12023), .B(n12022), .Z(n12048) );
  XOR U12256 ( .A(n12047), .B(n12048), .Z(n12049) );
  XNOR U12257 ( .A(n12050), .B(n12049), .Z(n11998) );
  NAND U12258 ( .A(n11970), .B(n11969), .Z(n11974) );
  NAND U12259 ( .A(n11972), .B(n11971), .Z(n11973) );
  NAND U12260 ( .A(n11974), .B(n11973), .Z(n11999) );
  XOR U12261 ( .A(n11998), .B(n11999), .Z(n12001) );
  XNOR U12262 ( .A(n12000), .B(n12001), .Z(n12059) );
  NANDN U12263 ( .A(n11976), .B(n11975), .Z(n11980) );
  NAND U12264 ( .A(n11978), .B(n11977), .Z(n11979) );
  NAND U12265 ( .A(n11980), .B(n11979), .Z(n12060) );
  XNOR U12266 ( .A(n12059), .B(n12060), .Z(n12061) );
  XOR U12267 ( .A(n12062), .B(n12061), .Z(n11992) );
  NANDN U12268 ( .A(n11982), .B(n11981), .Z(n11986) );
  NANDN U12269 ( .A(n11984), .B(n11983), .Z(n11985) );
  NAND U12270 ( .A(n11986), .B(n11985), .Z(n11993) );
  XNOR U12271 ( .A(n11992), .B(n11993), .Z(n11994) );
  XNOR U12272 ( .A(n11995), .B(n11994), .Z(n12065) );
  XNOR U12273 ( .A(n12065), .B(sreg[400]), .Z(n12067) );
  NAND U12274 ( .A(n11987), .B(sreg[399]), .Z(n11991) );
  OR U12275 ( .A(n11989), .B(n11988), .Z(n11990) );
  AND U12276 ( .A(n11991), .B(n11990), .Z(n12066) );
  XOR U12277 ( .A(n12067), .B(n12066), .Z(c[400]) );
  NANDN U12278 ( .A(n11993), .B(n11992), .Z(n11997) );
  NAND U12279 ( .A(n11995), .B(n11994), .Z(n11996) );
  NAND U12280 ( .A(n11997), .B(n11996), .Z(n12073) );
  NANDN U12281 ( .A(n11999), .B(n11998), .Z(n12003) );
  OR U12282 ( .A(n12001), .B(n12000), .Z(n12002) );
  NAND U12283 ( .A(n12003), .B(n12002), .Z(n12140) );
  XNOR U12284 ( .A(n20052), .B(n12346), .Z(n12109) );
  OR U12285 ( .A(n12109), .B(n20020), .Z(n12006) );
  NANDN U12286 ( .A(n12004), .B(n19960), .Z(n12005) );
  NAND U12287 ( .A(n12006), .B(n12005), .Z(n12122) );
  XNOR U12288 ( .A(n102), .B(n12007), .Z(n12113) );
  OR U12289 ( .A(n12113), .B(n20121), .Z(n12010) );
  NANDN U12290 ( .A(n12008), .B(n20122), .Z(n12009) );
  NAND U12291 ( .A(n12010), .B(n12009), .Z(n12119) );
  XNOR U12292 ( .A(n19975), .B(n12475), .Z(n12116) );
  NANDN U12293 ( .A(n12116), .B(n19883), .Z(n12013) );
  NANDN U12294 ( .A(n12011), .B(n19937), .Z(n12012) );
  AND U12295 ( .A(n12013), .B(n12012), .Z(n12120) );
  XNOR U12296 ( .A(n12119), .B(n12120), .Z(n12121) );
  XNOR U12297 ( .A(n12122), .B(n12121), .Z(n12131) );
  NANDN U12298 ( .A(n12015), .B(n12014), .Z(n12019) );
  NAND U12299 ( .A(n12017), .B(n12016), .Z(n12018) );
  NAND U12300 ( .A(n12019), .B(n12018), .Z(n12132) );
  XNOR U12301 ( .A(n12131), .B(n12132), .Z(n12133) );
  NANDN U12302 ( .A(n12021), .B(n12020), .Z(n12025) );
  NAND U12303 ( .A(n12023), .B(n12022), .Z(n12024) );
  AND U12304 ( .A(n12025), .B(n12024), .Z(n12134) );
  XNOR U12305 ( .A(n12133), .B(n12134), .Z(n12078) );
  NANDN U12306 ( .A(n12027), .B(n12026), .Z(n12031) );
  OR U12307 ( .A(n12029), .B(n12028), .Z(n12030) );
  NAND U12308 ( .A(n12031), .B(n12030), .Z(n12106) );
  NAND U12309 ( .A(b[0]), .B(a[161]), .Z(n12032) );
  XNOR U12310 ( .A(b[1]), .B(n12032), .Z(n12034) );
  NAND U12311 ( .A(a[160]), .B(n98), .Z(n12033) );
  AND U12312 ( .A(n12034), .B(n12033), .Z(n12082) );
  XNOR U12313 ( .A(n20154), .B(n12163), .Z(n12091) );
  OR U12314 ( .A(n12091), .B(n20057), .Z(n12037) );
  NANDN U12315 ( .A(n12035), .B(n20098), .Z(n12036) );
  AND U12316 ( .A(n12037), .B(n12036), .Z(n12083) );
  XOR U12317 ( .A(n12082), .B(n12083), .Z(n12085) );
  NAND U12318 ( .A(a[145]), .B(b[15]), .Z(n12084) );
  XOR U12319 ( .A(n12085), .B(n12084), .Z(n12103) );
  NAND U12320 ( .A(n19722), .B(n12038), .Z(n12040) );
  XNOR U12321 ( .A(b[5]), .B(n12787), .Z(n12094) );
  NANDN U12322 ( .A(n19640), .B(n12094), .Z(n12039) );
  NAND U12323 ( .A(n12040), .B(n12039), .Z(n12128) );
  XNOR U12324 ( .A(n19714), .B(n12631), .Z(n12097) );
  NANDN U12325 ( .A(n12097), .B(n19766), .Z(n12043) );
  NANDN U12326 ( .A(n12041), .B(n19767), .Z(n12042) );
  NAND U12327 ( .A(n12043), .B(n12042), .Z(n12125) );
  NAND U12328 ( .A(n19554), .B(n12044), .Z(n12046) );
  IV U12329 ( .A(a[159]), .Z(n12943) );
  XNOR U12330 ( .A(b[3]), .B(n12943), .Z(n12100) );
  NANDN U12331 ( .A(n19521), .B(n12100), .Z(n12045) );
  AND U12332 ( .A(n12046), .B(n12045), .Z(n12126) );
  XNOR U12333 ( .A(n12125), .B(n12126), .Z(n12127) );
  XOR U12334 ( .A(n12128), .B(n12127), .Z(n12104) );
  XOR U12335 ( .A(n12103), .B(n12104), .Z(n12105) );
  XNOR U12336 ( .A(n12106), .B(n12105), .Z(n12076) );
  NAND U12337 ( .A(n12048), .B(n12047), .Z(n12052) );
  NAND U12338 ( .A(n12050), .B(n12049), .Z(n12051) );
  NAND U12339 ( .A(n12052), .B(n12051), .Z(n12077) );
  XOR U12340 ( .A(n12076), .B(n12077), .Z(n12079) );
  XNOR U12341 ( .A(n12078), .B(n12079), .Z(n12137) );
  NANDN U12342 ( .A(n12054), .B(n12053), .Z(n12058) );
  NAND U12343 ( .A(n12056), .B(n12055), .Z(n12057) );
  NAND U12344 ( .A(n12058), .B(n12057), .Z(n12138) );
  XNOR U12345 ( .A(n12137), .B(n12138), .Z(n12139) );
  XOR U12346 ( .A(n12140), .B(n12139), .Z(n12070) );
  NANDN U12347 ( .A(n12060), .B(n12059), .Z(n12064) );
  NANDN U12348 ( .A(n12062), .B(n12061), .Z(n12063) );
  NAND U12349 ( .A(n12064), .B(n12063), .Z(n12071) );
  XNOR U12350 ( .A(n12070), .B(n12071), .Z(n12072) );
  XNOR U12351 ( .A(n12073), .B(n12072), .Z(n12143) );
  XNOR U12352 ( .A(n12143), .B(sreg[401]), .Z(n12145) );
  NAND U12353 ( .A(n12065), .B(sreg[400]), .Z(n12069) );
  OR U12354 ( .A(n12067), .B(n12066), .Z(n12068) );
  AND U12355 ( .A(n12069), .B(n12068), .Z(n12144) );
  XOR U12356 ( .A(n12145), .B(n12144), .Z(c[401]) );
  NANDN U12357 ( .A(n12071), .B(n12070), .Z(n12075) );
  NAND U12358 ( .A(n12073), .B(n12072), .Z(n12074) );
  NAND U12359 ( .A(n12075), .B(n12074), .Z(n12151) );
  NANDN U12360 ( .A(n12077), .B(n12076), .Z(n12081) );
  OR U12361 ( .A(n12079), .B(n12078), .Z(n12080) );
  NAND U12362 ( .A(n12081), .B(n12080), .Z(n12218) );
  NANDN U12363 ( .A(n12083), .B(n12082), .Z(n12087) );
  OR U12364 ( .A(n12085), .B(n12084), .Z(n12086) );
  NAND U12365 ( .A(n12087), .B(n12086), .Z(n12206) );
  NAND U12366 ( .A(b[0]), .B(a[162]), .Z(n12088) );
  XNOR U12367 ( .A(b[1]), .B(n12088), .Z(n12090) );
  NAND U12368 ( .A(a[161]), .B(n98), .Z(n12089) );
  AND U12369 ( .A(n12090), .B(n12089), .Z(n12182) );
  XNOR U12370 ( .A(n20154), .B(n12241), .Z(n12191) );
  OR U12371 ( .A(n12191), .B(n20057), .Z(n12093) );
  NANDN U12372 ( .A(n12091), .B(n20098), .Z(n12092) );
  AND U12373 ( .A(n12093), .B(n12092), .Z(n12183) );
  XOR U12374 ( .A(n12182), .B(n12183), .Z(n12185) );
  NAND U12375 ( .A(a[146]), .B(b[15]), .Z(n12184) );
  XOR U12376 ( .A(n12185), .B(n12184), .Z(n12203) );
  NAND U12377 ( .A(n19722), .B(n12094), .Z(n12096) );
  XNOR U12378 ( .A(b[5]), .B(n12865), .Z(n12194) );
  NANDN U12379 ( .A(n19640), .B(n12194), .Z(n12095) );
  NAND U12380 ( .A(n12096), .B(n12095), .Z(n12179) );
  XNOR U12381 ( .A(n19714), .B(n12736), .Z(n12197) );
  NANDN U12382 ( .A(n12197), .B(n19766), .Z(n12099) );
  NANDN U12383 ( .A(n12097), .B(n19767), .Z(n12098) );
  NAND U12384 ( .A(n12099), .B(n12098), .Z(n12176) );
  NAND U12385 ( .A(n19554), .B(n12100), .Z(n12102) );
  IV U12386 ( .A(a[160]), .Z(n13021) );
  XNOR U12387 ( .A(b[3]), .B(n13021), .Z(n12200) );
  NANDN U12388 ( .A(n19521), .B(n12200), .Z(n12101) );
  AND U12389 ( .A(n12102), .B(n12101), .Z(n12177) );
  XNOR U12390 ( .A(n12176), .B(n12177), .Z(n12178) );
  XOR U12391 ( .A(n12179), .B(n12178), .Z(n12204) );
  XOR U12392 ( .A(n12203), .B(n12204), .Z(n12205) );
  XNOR U12393 ( .A(n12206), .B(n12205), .Z(n12154) );
  NAND U12394 ( .A(n12104), .B(n12103), .Z(n12108) );
  NAND U12395 ( .A(n12106), .B(n12105), .Z(n12107) );
  NAND U12396 ( .A(n12108), .B(n12107), .Z(n12155) );
  XOR U12397 ( .A(n12154), .B(n12155), .Z(n12157) );
  XNOR U12398 ( .A(n20052), .B(n12397), .Z(n12160) );
  OR U12399 ( .A(n12160), .B(n20020), .Z(n12111) );
  NANDN U12400 ( .A(n12109), .B(n19960), .Z(n12110) );
  NAND U12401 ( .A(n12111), .B(n12110), .Z(n12173) );
  XNOR U12402 ( .A(n102), .B(n12112), .Z(n12164) );
  OR U12403 ( .A(n12164), .B(n20121), .Z(n12115) );
  NANDN U12404 ( .A(n12113), .B(n20122), .Z(n12114) );
  NAND U12405 ( .A(n12115), .B(n12114), .Z(n12170) );
  XNOR U12406 ( .A(n19975), .B(n12580), .Z(n12167) );
  NANDN U12407 ( .A(n12167), .B(n19883), .Z(n12118) );
  NANDN U12408 ( .A(n12116), .B(n19937), .Z(n12117) );
  AND U12409 ( .A(n12118), .B(n12117), .Z(n12171) );
  XNOR U12410 ( .A(n12170), .B(n12171), .Z(n12172) );
  XNOR U12411 ( .A(n12173), .B(n12172), .Z(n12209) );
  NANDN U12412 ( .A(n12120), .B(n12119), .Z(n12124) );
  NAND U12413 ( .A(n12122), .B(n12121), .Z(n12123) );
  NAND U12414 ( .A(n12124), .B(n12123), .Z(n12210) );
  XNOR U12415 ( .A(n12209), .B(n12210), .Z(n12211) );
  NANDN U12416 ( .A(n12126), .B(n12125), .Z(n12130) );
  NAND U12417 ( .A(n12128), .B(n12127), .Z(n12129) );
  AND U12418 ( .A(n12130), .B(n12129), .Z(n12212) );
  XNOR U12419 ( .A(n12211), .B(n12212), .Z(n12156) );
  XNOR U12420 ( .A(n12157), .B(n12156), .Z(n12215) );
  NANDN U12421 ( .A(n12132), .B(n12131), .Z(n12136) );
  NAND U12422 ( .A(n12134), .B(n12133), .Z(n12135) );
  NAND U12423 ( .A(n12136), .B(n12135), .Z(n12216) );
  XNOR U12424 ( .A(n12215), .B(n12216), .Z(n12217) );
  XOR U12425 ( .A(n12218), .B(n12217), .Z(n12148) );
  NANDN U12426 ( .A(n12138), .B(n12137), .Z(n12142) );
  NANDN U12427 ( .A(n12140), .B(n12139), .Z(n12141) );
  NAND U12428 ( .A(n12142), .B(n12141), .Z(n12149) );
  XNOR U12429 ( .A(n12148), .B(n12149), .Z(n12150) );
  XNOR U12430 ( .A(n12151), .B(n12150), .Z(n12221) );
  XNOR U12431 ( .A(n12221), .B(sreg[402]), .Z(n12223) );
  NAND U12432 ( .A(n12143), .B(sreg[401]), .Z(n12147) );
  OR U12433 ( .A(n12145), .B(n12144), .Z(n12146) );
  AND U12434 ( .A(n12147), .B(n12146), .Z(n12222) );
  XOR U12435 ( .A(n12223), .B(n12222), .Z(c[402]) );
  NANDN U12436 ( .A(n12149), .B(n12148), .Z(n12153) );
  NAND U12437 ( .A(n12151), .B(n12150), .Z(n12152) );
  NAND U12438 ( .A(n12153), .B(n12152), .Z(n12229) );
  NANDN U12439 ( .A(n12155), .B(n12154), .Z(n12159) );
  OR U12440 ( .A(n12157), .B(n12156), .Z(n12158) );
  NAND U12441 ( .A(n12159), .B(n12158), .Z(n12296) );
  XNOR U12442 ( .A(n20052), .B(n12475), .Z(n12238) );
  OR U12443 ( .A(n12238), .B(n20020), .Z(n12162) );
  NANDN U12444 ( .A(n12160), .B(n19960), .Z(n12161) );
  NAND U12445 ( .A(n12162), .B(n12161), .Z(n12251) );
  XNOR U12446 ( .A(n102), .B(n12163), .Z(n12242) );
  OR U12447 ( .A(n12242), .B(n20121), .Z(n12166) );
  NANDN U12448 ( .A(n12164), .B(n20122), .Z(n12165) );
  NAND U12449 ( .A(n12166), .B(n12165), .Z(n12248) );
  XNOR U12450 ( .A(n19975), .B(n12631), .Z(n12245) );
  NANDN U12451 ( .A(n12245), .B(n19883), .Z(n12169) );
  NANDN U12452 ( .A(n12167), .B(n19937), .Z(n12168) );
  AND U12453 ( .A(n12169), .B(n12168), .Z(n12249) );
  XNOR U12454 ( .A(n12248), .B(n12249), .Z(n12250) );
  XNOR U12455 ( .A(n12251), .B(n12250), .Z(n12287) );
  NANDN U12456 ( .A(n12171), .B(n12170), .Z(n12175) );
  NAND U12457 ( .A(n12173), .B(n12172), .Z(n12174) );
  NAND U12458 ( .A(n12175), .B(n12174), .Z(n12288) );
  XNOR U12459 ( .A(n12287), .B(n12288), .Z(n12289) );
  NANDN U12460 ( .A(n12177), .B(n12176), .Z(n12181) );
  NAND U12461 ( .A(n12179), .B(n12178), .Z(n12180) );
  AND U12462 ( .A(n12181), .B(n12180), .Z(n12290) );
  XNOR U12463 ( .A(n12289), .B(n12290), .Z(n12234) );
  NANDN U12464 ( .A(n12183), .B(n12182), .Z(n12187) );
  OR U12465 ( .A(n12185), .B(n12184), .Z(n12186) );
  NAND U12466 ( .A(n12187), .B(n12186), .Z(n12284) );
  NAND U12467 ( .A(b[0]), .B(a[163]), .Z(n12188) );
  XNOR U12468 ( .A(b[1]), .B(n12188), .Z(n12190) );
  NAND U12469 ( .A(a[162]), .B(n98), .Z(n12189) );
  AND U12470 ( .A(n12190), .B(n12189), .Z(n12260) );
  XNOR U12471 ( .A(n20154), .B(n12346), .Z(n12269) );
  OR U12472 ( .A(n12269), .B(n20057), .Z(n12193) );
  NANDN U12473 ( .A(n12191), .B(n20098), .Z(n12192) );
  AND U12474 ( .A(n12193), .B(n12192), .Z(n12261) );
  XOR U12475 ( .A(n12260), .B(n12261), .Z(n12263) );
  NAND U12476 ( .A(a[147]), .B(b[15]), .Z(n12262) );
  XOR U12477 ( .A(n12263), .B(n12262), .Z(n12281) );
  NAND U12478 ( .A(n19722), .B(n12194), .Z(n12196) );
  XNOR U12479 ( .A(b[5]), .B(n12943), .Z(n12272) );
  NANDN U12480 ( .A(n19640), .B(n12272), .Z(n12195) );
  NAND U12481 ( .A(n12196), .B(n12195), .Z(n12257) );
  XNOR U12482 ( .A(n19714), .B(n12787), .Z(n12275) );
  NANDN U12483 ( .A(n12275), .B(n19766), .Z(n12199) );
  NANDN U12484 ( .A(n12197), .B(n19767), .Z(n12198) );
  NAND U12485 ( .A(n12199), .B(n12198), .Z(n12254) );
  NAND U12486 ( .A(n19554), .B(n12200), .Z(n12202) );
  IV U12487 ( .A(a[161]), .Z(n13126) );
  XNOR U12488 ( .A(b[3]), .B(n13126), .Z(n12278) );
  NANDN U12489 ( .A(n19521), .B(n12278), .Z(n12201) );
  AND U12490 ( .A(n12202), .B(n12201), .Z(n12255) );
  XNOR U12491 ( .A(n12254), .B(n12255), .Z(n12256) );
  XOR U12492 ( .A(n12257), .B(n12256), .Z(n12282) );
  XOR U12493 ( .A(n12281), .B(n12282), .Z(n12283) );
  XNOR U12494 ( .A(n12284), .B(n12283), .Z(n12232) );
  NAND U12495 ( .A(n12204), .B(n12203), .Z(n12208) );
  NAND U12496 ( .A(n12206), .B(n12205), .Z(n12207) );
  NAND U12497 ( .A(n12208), .B(n12207), .Z(n12233) );
  XOR U12498 ( .A(n12232), .B(n12233), .Z(n12235) );
  XNOR U12499 ( .A(n12234), .B(n12235), .Z(n12293) );
  NANDN U12500 ( .A(n12210), .B(n12209), .Z(n12214) );
  NAND U12501 ( .A(n12212), .B(n12211), .Z(n12213) );
  NAND U12502 ( .A(n12214), .B(n12213), .Z(n12294) );
  XNOR U12503 ( .A(n12293), .B(n12294), .Z(n12295) );
  XOR U12504 ( .A(n12296), .B(n12295), .Z(n12226) );
  NANDN U12505 ( .A(n12216), .B(n12215), .Z(n12220) );
  NANDN U12506 ( .A(n12218), .B(n12217), .Z(n12219) );
  NAND U12507 ( .A(n12220), .B(n12219), .Z(n12227) );
  XNOR U12508 ( .A(n12226), .B(n12227), .Z(n12228) );
  XNOR U12509 ( .A(n12229), .B(n12228), .Z(n12299) );
  XNOR U12510 ( .A(n12299), .B(sreg[403]), .Z(n12301) );
  NAND U12511 ( .A(n12221), .B(sreg[402]), .Z(n12225) );
  OR U12512 ( .A(n12223), .B(n12222), .Z(n12224) );
  AND U12513 ( .A(n12225), .B(n12224), .Z(n12300) );
  XOR U12514 ( .A(n12301), .B(n12300), .Z(c[403]) );
  NANDN U12515 ( .A(n12227), .B(n12226), .Z(n12231) );
  NAND U12516 ( .A(n12229), .B(n12228), .Z(n12230) );
  NAND U12517 ( .A(n12231), .B(n12230), .Z(n12307) );
  NANDN U12518 ( .A(n12233), .B(n12232), .Z(n12237) );
  OR U12519 ( .A(n12235), .B(n12234), .Z(n12236) );
  NAND U12520 ( .A(n12237), .B(n12236), .Z(n12374) );
  XNOR U12521 ( .A(n20052), .B(n12580), .Z(n12343) );
  OR U12522 ( .A(n12343), .B(n20020), .Z(n12240) );
  NANDN U12523 ( .A(n12238), .B(n19960), .Z(n12239) );
  NAND U12524 ( .A(n12240), .B(n12239), .Z(n12356) );
  XNOR U12525 ( .A(n102), .B(n12241), .Z(n12347) );
  OR U12526 ( .A(n12347), .B(n20121), .Z(n12244) );
  NANDN U12527 ( .A(n12242), .B(n20122), .Z(n12243) );
  NAND U12528 ( .A(n12244), .B(n12243), .Z(n12353) );
  XNOR U12529 ( .A(n19975), .B(n12736), .Z(n12350) );
  NANDN U12530 ( .A(n12350), .B(n19883), .Z(n12247) );
  NANDN U12531 ( .A(n12245), .B(n19937), .Z(n12246) );
  AND U12532 ( .A(n12247), .B(n12246), .Z(n12354) );
  XNOR U12533 ( .A(n12353), .B(n12354), .Z(n12355) );
  XNOR U12534 ( .A(n12356), .B(n12355), .Z(n12365) );
  NANDN U12535 ( .A(n12249), .B(n12248), .Z(n12253) );
  NAND U12536 ( .A(n12251), .B(n12250), .Z(n12252) );
  NAND U12537 ( .A(n12253), .B(n12252), .Z(n12366) );
  XNOR U12538 ( .A(n12365), .B(n12366), .Z(n12367) );
  NANDN U12539 ( .A(n12255), .B(n12254), .Z(n12259) );
  NAND U12540 ( .A(n12257), .B(n12256), .Z(n12258) );
  AND U12541 ( .A(n12259), .B(n12258), .Z(n12368) );
  XNOR U12542 ( .A(n12367), .B(n12368), .Z(n12312) );
  NANDN U12543 ( .A(n12261), .B(n12260), .Z(n12265) );
  OR U12544 ( .A(n12263), .B(n12262), .Z(n12264) );
  NAND U12545 ( .A(n12265), .B(n12264), .Z(n12340) );
  NAND U12546 ( .A(b[0]), .B(a[164]), .Z(n12266) );
  XNOR U12547 ( .A(b[1]), .B(n12266), .Z(n12268) );
  NAND U12548 ( .A(a[163]), .B(n98), .Z(n12267) );
  AND U12549 ( .A(n12268), .B(n12267), .Z(n12316) );
  XNOR U12550 ( .A(n20154), .B(n12397), .Z(n12325) );
  OR U12551 ( .A(n12325), .B(n20057), .Z(n12271) );
  NANDN U12552 ( .A(n12269), .B(n20098), .Z(n12270) );
  AND U12553 ( .A(n12271), .B(n12270), .Z(n12317) );
  XOR U12554 ( .A(n12316), .B(n12317), .Z(n12319) );
  NAND U12555 ( .A(a[148]), .B(b[15]), .Z(n12318) );
  XOR U12556 ( .A(n12319), .B(n12318), .Z(n12337) );
  NAND U12557 ( .A(n19722), .B(n12272), .Z(n12274) );
  XNOR U12558 ( .A(b[5]), .B(n13021), .Z(n12328) );
  NANDN U12559 ( .A(n19640), .B(n12328), .Z(n12273) );
  NAND U12560 ( .A(n12274), .B(n12273), .Z(n12362) );
  XNOR U12561 ( .A(n19714), .B(n12865), .Z(n12331) );
  NANDN U12562 ( .A(n12331), .B(n19766), .Z(n12277) );
  NANDN U12563 ( .A(n12275), .B(n19767), .Z(n12276) );
  NAND U12564 ( .A(n12277), .B(n12276), .Z(n12359) );
  NAND U12565 ( .A(n19554), .B(n12278), .Z(n12280) );
  IV U12566 ( .A(a[162]), .Z(n13204) );
  XNOR U12567 ( .A(b[3]), .B(n13204), .Z(n12334) );
  NANDN U12568 ( .A(n19521), .B(n12334), .Z(n12279) );
  AND U12569 ( .A(n12280), .B(n12279), .Z(n12360) );
  XNOR U12570 ( .A(n12359), .B(n12360), .Z(n12361) );
  XOR U12571 ( .A(n12362), .B(n12361), .Z(n12338) );
  XOR U12572 ( .A(n12337), .B(n12338), .Z(n12339) );
  XNOR U12573 ( .A(n12340), .B(n12339), .Z(n12310) );
  NAND U12574 ( .A(n12282), .B(n12281), .Z(n12286) );
  NAND U12575 ( .A(n12284), .B(n12283), .Z(n12285) );
  NAND U12576 ( .A(n12286), .B(n12285), .Z(n12311) );
  XOR U12577 ( .A(n12310), .B(n12311), .Z(n12313) );
  XNOR U12578 ( .A(n12312), .B(n12313), .Z(n12371) );
  NANDN U12579 ( .A(n12288), .B(n12287), .Z(n12292) );
  NAND U12580 ( .A(n12290), .B(n12289), .Z(n12291) );
  NAND U12581 ( .A(n12292), .B(n12291), .Z(n12372) );
  XNOR U12582 ( .A(n12371), .B(n12372), .Z(n12373) );
  XOR U12583 ( .A(n12374), .B(n12373), .Z(n12304) );
  NANDN U12584 ( .A(n12294), .B(n12293), .Z(n12298) );
  NANDN U12585 ( .A(n12296), .B(n12295), .Z(n12297) );
  NAND U12586 ( .A(n12298), .B(n12297), .Z(n12305) );
  XNOR U12587 ( .A(n12304), .B(n12305), .Z(n12306) );
  XNOR U12588 ( .A(n12307), .B(n12306), .Z(n12377) );
  XNOR U12589 ( .A(n12377), .B(sreg[404]), .Z(n12379) );
  NAND U12590 ( .A(n12299), .B(sreg[403]), .Z(n12303) );
  OR U12591 ( .A(n12301), .B(n12300), .Z(n12302) );
  AND U12592 ( .A(n12303), .B(n12302), .Z(n12378) );
  XOR U12593 ( .A(n12379), .B(n12378), .Z(c[404]) );
  NANDN U12594 ( .A(n12305), .B(n12304), .Z(n12309) );
  NAND U12595 ( .A(n12307), .B(n12306), .Z(n12308) );
  NAND U12596 ( .A(n12309), .B(n12308), .Z(n12385) );
  NANDN U12597 ( .A(n12311), .B(n12310), .Z(n12315) );
  OR U12598 ( .A(n12313), .B(n12312), .Z(n12314) );
  NAND U12599 ( .A(n12315), .B(n12314), .Z(n12452) );
  NANDN U12600 ( .A(n12317), .B(n12316), .Z(n12321) );
  OR U12601 ( .A(n12319), .B(n12318), .Z(n12320) );
  NAND U12602 ( .A(n12321), .B(n12320), .Z(n12440) );
  NAND U12603 ( .A(b[0]), .B(a[165]), .Z(n12322) );
  XNOR U12604 ( .A(b[1]), .B(n12322), .Z(n12324) );
  NAND U12605 ( .A(a[164]), .B(n98), .Z(n12323) );
  AND U12606 ( .A(n12324), .B(n12323), .Z(n12416) );
  XNOR U12607 ( .A(n20154), .B(n12475), .Z(n12425) );
  OR U12608 ( .A(n12425), .B(n20057), .Z(n12327) );
  NANDN U12609 ( .A(n12325), .B(n20098), .Z(n12326) );
  AND U12610 ( .A(n12327), .B(n12326), .Z(n12417) );
  XOR U12611 ( .A(n12416), .B(n12417), .Z(n12419) );
  NAND U12612 ( .A(a[149]), .B(b[15]), .Z(n12418) );
  XOR U12613 ( .A(n12419), .B(n12418), .Z(n12437) );
  NAND U12614 ( .A(n19722), .B(n12328), .Z(n12330) );
  XNOR U12615 ( .A(b[5]), .B(n13126), .Z(n12428) );
  NANDN U12616 ( .A(n19640), .B(n12428), .Z(n12329) );
  NAND U12617 ( .A(n12330), .B(n12329), .Z(n12413) );
  XNOR U12618 ( .A(n19714), .B(n12943), .Z(n12431) );
  NANDN U12619 ( .A(n12431), .B(n19766), .Z(n12333) );
  NANDN U12620 ( .A(n12331), .B(n19767), .Z(n12332) );
  NAND U12621 ( .A(n12333), .B(n12332), .Z(n12410) );
  NAND U12622 ( .A(n19554), .B(n12334), .Z(n12336) );
  IV U12623 ( .A(a[163]), .Z(n13282) );
  XNOR U12624 ( .A(b[3]), .B(n13282), .Z(n12434) );
  NANDN U12625 ( .A(n19521), .B(n12434), .Z(n12335) );
  AND U12626 ( .A(n12336), .B(n12335), .Z(n12411) );
  XNOR U12627 ( .A(n12410), .B(n12411), .Z(n12412) );
  XOR U12628 ( .A(n12413), .B(n12412), .Z(n12438) );
  XOR U12629 ( .A(n12437), .B(n12438), .Z(n12439) );
  XNOR U12630 ( .A(n12440), .B(n12439), .Z(n12388) );
  NAND U12631 ( .A(n12338), .B(n12337), .Z(n12342) );
  NAND U12632 ( .A(n12340), .B(n12339), .Z(n12341) );
  NAND U12633 ( .A(n12342), .B(n12341), .Z(n12389) );
  XOR U12634 ( .A(n12388), .B(n12389), .Z(n12391) );
  XNOR U12635 ( .A(n20052), .B(n12631), .Z(n12394) );
  OR U12636 ( .A(n12394), .B(n20020), .Z(n12345) );
  NANDN U12637 ( .A(n12343), .B(n19960), .Z(n12344) );
  NAND U12638 ( .A(n12345), .B(n12344), .Z(n12407) );
  XNOR U12639 ( .A(n102), .B(n12346), .Z(n12398) );
  OR U12640 ( .A(n12398), .B(n20121), .Z(n12349) );
  NANDN U12641 ( .A(n12347), .B(n20122), .Z(n12348) );
  NAND U12642 ( .A(n12349), .B(n12348), .Z(n12404) );
  XNOR U12643 ( .A(n19975), .B(n12787), .Z(n12401) );
  NANDN U12644 ( .A(n12401), .B(n19883), .Z(n12352) );
  NANDN U12645 ( .A(n12350), .B(n19937), .Z(n12351) );
  AND U12646 ( .A(n12352), .B(n12351), .Z(n12405) );
  XNOR U12647 ( .A(n12404), .B(n12405), .Z(n12406) );
  XNOR U12648 ( .A(n12407), .B(n12406), .Z(n12443) );
  NANDN U12649 ( .A(n12354), .B(n12353), .Z(n12358) );
  NAND U12650 ( .A(n12356), .B(n12355), .Z(n12357) );
  NAND U12651 ( .A(n12358), .B(n12357), .Z(n12444) );
  XNOR U12652 ( .A(n12443), .B(n12444), .Z(n12445) );
  NANDN U12653 ( .A(n12360), .B(n12359), .Z(n12364) );
  NAND U12654 ( .A(n12362), .B(n12361), .Z(n12363) );
  AND U12655 ( .A(n12364), .B(n12363), .Z(n12446) );
  XNOR U12656 ( .A(n12445), .B(n12446), .Z(n12390) );
  XNOR U12657 ( .A(n12391), .B(n12390), .Z(n12449) );
  NANDN U12658 ( .A(n12366), .B(n12365), .Z(n12370) );
  NAND U12659 ( .A(n12368), .B(n12367), .Z(n12369) );
  NAND U12660 ( .A(n12370), .B(n12369), .Z(n12450) );
  XNOR U12661 ( .A(n12449), .B(n12450), .Z(n12451) );
  XOR U12662 ( .A(n12452), .B(n12451), .Z(n12382) );
  NANDN U12663 ( .A(n12372), .B(n12371), .Z(n12376) );
  NANDN U12664 ( .A(n12374), .B(n12373), .Z(n12375) );
  NAND U12665 ( .A(n12376), .B(n12375), .Z(n12383) );
  XNOR U12666 ( .A(n12382), .B(n12383), .Z(n12384) );
  XNOR U12667 ( .A(n12385), .B(n12384), .Z(n12455) );
  XNOR U12668 ( .A(n12455), .B(sreg[405]), .Z(n12457) );
  NAND U12669 ( .A(n12377), .B(sreg[404]), .Z(n12381) );
  OR U12670 ( .A(n12379), .B(n12378), .Z(n12380) );
  AND U12671 ( .A(n12381), .B(n12380), .Z(n12456) );
  XOR U12672 ( .A(n12457), .B(n12456), .Z(c[405]) );
  NANDN U12673 ( .A(n12383), .B(n12382), .Z(n12387) );
  NAND U12674 ( .A(n12385), .B(n12384), .Z(n12386) );
  NAND U12675 ( .A(n12387), .B(n12386), .Z(n12463) );
  NANDN U12676 ( .A(n12389), .B(n12388), .Z(n12393) );
  OR U12677 ( .A(n12391), .B(n12390), .Z(n12392) );
  NAND U12678 ( .A(n12393), .B(n12392), .Z(n12530) );
  XNOR U12679 ( .A(n20052), .B(n12736), .Z(n12472) );
  OR U12680 ( .A(n12472), .B(n20020), .Z(n12396) );
  NANDN U12681 ( .A(n12394), .B(n19960), .Z(n12395) );
  NAND U12682 ( .A(n12396), .B(n12395), .Z(n12485) );
  XNOR U12683 ( .A(n102), .B(n12397), .Z(n12476) );
  OR U12684 ( .A(n12476), .B(n20121), .Z(n12400) );
  NANDN U12685 ( .A(n12398), .B(n20122), .Z(n12399) );
  NAND U12686 ( .A(n12400), .B(n12399), .Z(n12482) );
  XNOR U12687 ( .A(n19975), .B(n12865), .Z(n12479) );
  NANDN U12688 ( .A(n12479), .B(n19883), .Z(n12403) );
  NANDN U12689 ( .A(n12401), .B(n19937), .Z(n12402) );
  AND U12690 ( .A(n12403), .B(n12402), .Z(n12483) );
  XNOR U12691 ( .A(n12482), .B(n12483), .Z(n12484) );
  XNOR U12692 ( .A(n12485), .B(n12484), .Z(n12521) );
  NANDN U12693 ( .A(n12405), .B(n12404), .Z(n12409) );
  NAND U12694 ( .A(n12407), .B(n12406), .Z(n12408) );
  NAND U12695 ( .A(n12409), .B(n12408), .Z(n12522) );
  XNOR U12696 ( .A(n12521), .B(n12522), .Z(n12523) );
  NANDN U12697 ( .A(n12411), .B(n12410), .Z(n12415) );
  NAND U12698 ( .A(n12413), .B(n12412), .Z(n12414) );
  AND U12699 ( .A(n12415), .B(n12414), .Z(n12524) );
  XNOR U12700 ( .A(n12523), .B(n12524), .Z(n12468) );
  NANDN U12701 ( .A(n12417), .B(n12416), .Z(n12421) );
  OR U12702 ( .A(n12419), .B(n12418), .Z(n12420) );
  NAND U12703 ( .A(n12421), .B(n12420), .Z(n12518) );
  NAND U12704 ( .A(b[0]), .B(a[166]), .Z(n12422) );
  XNOR U12705 ( .A(b[1]), .B(n12422), .Z(n12424) );
  NAND U12706 ( .A(a[165]), .B(n98), .Z(n12423) );
  AND U12707 ( .A(n12424), .B(n12423), .Z(n12494) );
  XNOR U12708 ( .A(n20154), .B(n12580), .Z(n12500) );
  OR U12709 ( .A(n12500), .B(n20057), .Z(n12427) );
  NANDN U12710 ( .A(n12425), .B(n20098), .Z(n12426) );
  AND U12711 ( .A(n12427), .B(n12426), .Z(n12495) );
  XOR U12712 ( .A(n12494), .B(n12495), .Z(n12497) );
  NAND U12713 ( .A(a[150]), .B(b[15]), .Z(n12496) );
  XOR U12714 ( .A(n12497), .B(n12496), .Z(n12515) );
  NAND U12715 ( .A(n19722), .B(n12428), .Z(n12430) );
  XNOR U12716 ( .A(b[5]), .B(n13204), .Z(n12506) );
  NANDN U12717 ( .A(n19640), .B(n12506), .Z(n12429) );
  NAND U12718 ( .A(n12430), .B(n12429), .Z(n12491) );
  XNOR U12719 ( .A(n19714), .B(n13021), .Z(n12509) );
  NANDN U12720 ( .A(n12509), .B(n19766), .Z(n12433) );
  NANDN U12721 ( .A(n12431), .B(n19767), .Z(n12432) );
  NAND U12722 ( .A(n12433), .B(n12432), .Z(n12488) );
  NAND U12723 ( .A(n19554), .B(n12434), .Z(n12436) );
  IV U12724 ( .A(a[164]), .Z(n13333) );
  XNOR U12725 ( .A(b[3]), .B(n13333), .Z(n12512) );
  NANDN U12726 ( .A(n19521), .B(n12512), .Z(n12435) );
  AND U12727 ( .A(n12436), .B(n12435), .Z(n12489) );
  XNOR U12728 ( .A(n12488), .B(n12489), .Z(n12490) );
  XOR U12729 ( .A(n12491), .B(n12490), .Z(n12516) );
  XOR U12730 ( .A(n12515), .B(n12516), .Z(n12517) );
  XNOR U12731 ( .A(n12518), .B(n12517), .Z(n12466) );
  NAND U12732 ( .A(n12438), .B(n12437), .Z(n12442) );
  NAND U12733 ( .A(n12440), .B(n12439), .Z(n12441) );
  NAND U12734 ( .A(n12442), .B(n12441), .Z(n12467) );
  XOR U12735 ( .A(n12466), .B(n12467), .Z(n12469) );
  XNOR U12736 ( .A(n12468), .B(n12469), .Z(n12527) );
  NANDN U12737 ( .A(n12444), .B(n12443), .Z(n12448) );
  NAND U12738 ( .A(n12446), .B(n12445), .Z(n12447) );
  NAND U12739 ( .A(n12448), .B(n12447), .Z(n12528) );
  XNOR U12740 ( .A(n12527), .B(n12528), .Z(n12529) );
  XOR U12741 ( .A(n12530), .B(n12529), .Z(n12460) );
  NANDN U12742 ( .A(n12450), .B(n12449), .Z(n12454) );
  NANDN U12743 ( .A(n12452), .B(n12451), .Z(n12453) );
  NAND U12744 ( .A(n12454), .B(n12453), .Z(n12461) );
  XNOR U12745 ( .A(n12460), .B(n12461), .Z(n12462) );
  XNOR U12746 ( .A(n12463), .B(n12462), .Z(n12533) );
  XNOR U12747 ( .A(n12533), .B(sreg[406]), .Z(n12535) );
  NAND U12748 ( .A(n12455), .B(sreg[405]), .Z(n12459) );
  OR U12749 ( .A(n12457), .B(n12456), .Z(n12458) );
  AND U12750 ( .A(n12459), .B(n12458), .Z(n12534) );
  XOR U12751 ( .A(n12535), .B(n12534), .Z(c[406]) );
  NANDN U12752 ( .A(n12461), .B(n12460), .Z(n12465) );
  NAND U12753 ( .A(n12463), .B(n12462), .Z(n12464) );
  NAND U12754 ( .A(n12465), .B(n12464), .Z(n12541) );
  NANDN U12755 ( .A(n12467), .B(n12466), .Z(n12471) );
  OR U12756 ( .A(n12469), .B(n12468), .Z(n12470) );
  NAND U12757 ( .A(n12471), .B(n12470), .Z(n12608) );
  XNOR U12758 ( .A(n20052), .B(n12787), .Z(n12577) );
  OR U12759 ( .A(n12577), .B(n20020), .Z(n12474) );
  NANDN U12760 ( .A(n12472), .B(n19960), .Z(n12473) );
  NAND U12761 ( .A(n12474), .B(n12473), .Z(n12590) );
  XNOR U12762 ( .A(n102), .B(n12475), .Z(n12581) );
  OR U12763 ( .A(n12581), .B(n20121), .Z(n12478) );
  NANDN U12764 ( .A(n12476), .B(n20122), .Z(n12477) );
  NAND U12765 ( .A(n12478), .B(n12477), .Z(n12587) );
  XNOR U12766 ( .A(n19975), .B(n12943), .Z(n12584) );
  NANDN U12767 ( .A(n12584), .B(n19883), .Z(n12481) );
  NANDN U12768 ( .A(n12479), .B(n19937), .Z(n12480) );
  AND U12769 ( .A(n12481), .B(n12480), .Z(n12588) );
  XNOR U12770 ( .A(n12587), .B(n12588), .Z(n12589) );
  XNOR U12771 ( .A(n12590), .B(n12589), .Z(n12599) );
  NANDN U12772 ( .A(n12483), .B(n12482), .Z(n12487) );
  NAND U12773 ( .A(n12485), .B(n12484), .Z(n12486) );
  NAND U12774 ( .A(n12487), .B(n12486), .Z(n12600) );
  XNOR U12775 ( .A(n12599), .B(n12600), .Z(n12601) );
  NANDN U12776 ( .A(n12489), .B(n12488), .Z(n12493) );
  NAND U12777 ( .A(n12491), .B(n12490), .Z(n12492) );
  AND U12778 ( .A(n12493), .B(n12492), .Z(n12602) );
  XNOR U12779 ( .A(n12601), .B(n12602), .Z(n12546) );
  NANDN U12780 ( .A(n12495), .B(n12494), .Z(n12499) );
  OR U12781 ( .A(n12497), .B(n12496), .Z(n12498) );
  NAND U12782 ( .A(n12499), .B(n12498), .Z(n12574) );
  XNOR U12783 ( .A(n20154), .B(n12631), .Z(n12556) );
  OR U12784 ( .A(n12556), .B(n20057), .Z(n12502) );
  NANDN U12785 ( .A(n12500), .B(n20098), .Z(n12501) );
  AND U12786 ( .A(n12502), .B(n12501), .Z(n12551) );
  NAND U12787 ( .A(b[0]), .B(a[167]), .Z(n12503) );
  XNOR U12788 ( .A(b[1]), .B(n12503), .Z(n12505) );
  NAND U12789 ( .A(a[166]), .B(n98), .Z(n12504) );
  AND U12790 ( .A(n12505), .B(n12504), .Z(n12550) );
  XOR U12791 ( .A(n12551), .B(n12550), .Z(n12553) );
  NAND U12792 ( .A(a[151]), .B(b[15]), .Z(n12552) );
  XOR U12793 ( .A(n12553), .B(n12552), .Z(n12571) );
  NAND U12794 ( .A(n19722), .B(n12506), .Z(n12508) );
  XNOR U12795 ( .A(b[5]), .B(n13282), .Z(n12562) );
  NANDN U12796 ( .A(n19640), .B(n12562), .Z(n12507) );
  NAND U12797 ( .A(n12508), .B(n12507), .Z(n12596) );
  XNOR U12798 ( .A(n19714), .B(n13126), .Z(n12565) );
  NANDN U12799 ( .A(n12565), .B(n19766), .Z(n12511) );
  NANDN U12800 ( .A(n12509), .B(n19767), .Z(n12510) );
  NAND U12801 ( .A(n12511), .B(n12510), .Z(n12593) );
  NAND U12802 ( .A(n19554), .B(n12512), .Z(n12514) );
  IV U12803 ( .A(a[165]), .Z(n13438) );
  XNOR U12804 ( .A(b[3]), .B(n13438), .Z(n12568) );
  NANDN U12805 ( .A(n19521), .B(n12568), .Z(n12513) );
  AND U12806 ( .A(n12514), .B(n12513), .Z(n12594) );
  XNOR U12807 ( .A(n12593), .B(n12594), .Z(n12595) );
  XOR U12808 ( .A(n12596), .B(n12595), .Z(n12572) );
  XOR U12809 ( .A(n12571), .B(n12572), .Z(n12573) );
  XNOR U12810 ( .A(n12574), .B(n12573), .Z(n12544) );
  NAND U12811 ( .A(n12516), .B(n12515), .Z(n12520) );
  NAND U12812 ( .A(n12518), .B(n12517), .Z(n12519) );
  NAND U12813 ( .A(n12520), .B(n12519), .Z(n12545) );
  XOR U12814 ( .A(n12544), .B(n12545), .Z(n12547) );
  XNOR U12815 ( .A(n12546), .B(n12547), .Z(n12605) );
  NANDN U12816 ( .A(n12522), .B(n12521), .Z(n12526) );
  NAND U12817 ( .A(n12524), .B(n12523), .Z(n12525) );
  NAND U12818 ( .A(n12526), .B(n12525), .Z(n12606) );
  XNOR U12819 ( .A(n12605), .B(n12606), .Z(n12607) );
  XOR U12820 ( .A(n12608), .B(n12607), .Z(n12538) );
  NANDN U12821 ( .A(n12528), .B(n12527), .Z(n12532) );
  NANDN U12822 ( .A(n12530), .B(n12529), .Z(n12531) );
  NAND U12823 ( .A(n12532), .B(n12531), .Z(n12539) );
  XNOR U12824 ( .A(n12538), .B(n12539), .Z(n12540) );
  XNOR U12825 ( .A(n12541), .B(n12540), .Z(n12611) );
  XNOR U12826 ( .A(n12611), .B(sreg[407]), .Z(n12613) );
  NAND U12827 ( .A(n12533), .B(sreg[406]), .Z(n12537) );
  OR U12828 ( .A(n12535), .B(n12534), .Z(n12536) );
  AND U12829 ( .A(n12537), .B(n12536), .Z(n12612) );
  XOR U12830 ( .A(n12613), .B(n12612), .Z(c[407]) );
  NANDN U12831 ( .A(n12539), .B(n12538), .Z(n12543) );
  NAND U12832 ( .A(n12541), .B(n12540), .Z(n12542) );
  NAND U12833 ( .A(n12543), .B(n12542), .Z(n12619) );
  NANDN U12834 ( .A(n12545), .B(n12544), .Z(n12549) );
  OR U12835 ( .A(n12547), .B(n12546), .Z(n12548) );
  NAND U12836 ( .A(n12549), .B(n12548), .Z(n12686) );
  NANDN U12837 ( .A(n12551), .B(n12550), .Z(n12555) );
  OR U12838 ( .A(n12553), .B(n12552), .Z(n12554) );
  NAND U12839 ( .A(n12555), .B(n12554), .Z(n12674) );
  XNOR U12840 ( .A(n20154), .B(n12736), .Z(n12659) );
  OR U12841 ( .A(n12659), .B(n20057), .Z(n12558) );
  NANDN U12842 ( .A(n12556), .B(n20098), .Z(n12557) );
  AND U12843 ( .A(n12558), .B(n12557), .Z(n12651) );
  NAND U12844 ( .A(b[0]), .B(a[168]), .Z(n12559) );
  XNOR U12845 ( .A(b[1]), .B(n12559), .Z(n12561) );
  NAND U12846 ( .A(a[167]), .B(n98), .Z(n12560) );
  AND U12847 ( .A(n12561), .B(n12560), .Z(n12650) );
  XOR U12848 ( .A(n12651), .B(n12650), .Z(n12653) );
  NAND U12849 ( .A(a[152]), .B(b[15]), .Z(n12652) );
  XOR U12850 ( .A(n12653), .B(n12652), .Z(n12671) );
  NAND U12851 ( .A(n19722), .B(n12562), .Z(n12564) );
  XNOR U12852 ( .A(b[5]), .B(n13333), .Z(n12662) );
  NANDN U12853 ( .A(n19640), .B(n12662), .Z(n12563) );
  NAND U12854 ( .A(n12564), .B(n12563), .Z(n12647) );
  XNOR U12855 ( .A(n19714), .B(n13204), .Z(n12665) );
  NANDN U12856 ( .A(n12665), .B(n19766), .Z(n12567) );
  NANDN U12857 ( .A(n12565), .B(n19767), .Z(n12566) );
  NAND U12858 ( .A(n12567), .B(n12566), .Z(n12644) );
  NAND U12859 ( .A(n19554), .B(n12568), .Z(n12570) );
  IV U12860 ( .A(a[166]), .Z(n13516) );
  XNOR U12861 ( .A(b[3]), .B(n13516), .Z(n12668) );
  NANDN U12862 ( .A(n19521), .B(n12668), .Z(n12569) );
  AND U12863 ( .A(n12570), .B(n12569), .Z(n12645) );
  XNOR U12864 ( .A(n12644), .B(n12645), .Z(n12646) );
  XOR U12865 ( .A(n12647), .B(n12646), .Z(n12672) );
  XOR U12866 ( .A(n12671), .B(n12672), .Z(n12673) );
  XNOR U12867 ( .A(n12674), .B(n12673), .Z(n12622) );
  NAND U12868 ( .A(n12572), .B(n12571), .Z(n12576) );
  NAND U12869 ( .A(n12574), .B(n12573), .Z(n12575) );
  NAND U12870 ( .A(n12576), .B(n12575), .Z(n12623) );
  XOR U12871 ( .A(n12622), .B(n12623), .Z(n12625) );
  XNOR U12872 ( .A(n20052), .B(n12865), .Z(n12628) );
  OR U12873 ( .A(n12628), .B(n20020), .Z(n12579) );
  NANDN U12874 ( .A(n12577), .B(n19960), .Z(n12578) );
  NAND U12875 ( .A(n12579), .B(n12578), .Z(n12641) );
  XNOR U12876 ( .A(n102), .B(n12580), .Z(n12632) );
  OR U12877 ( .A(n12632), .B(n20121), .Z(n12583) );
  NANDN U12878 ( .A(n12581), .B(n20122), .Z(n12582) );
  NAND U12879 ( .A(n12583), .B(n12582), .Z(n12638) );
  XNOR U12880 ( .A(n19975), .B(n13021), .Z(n12635) );
  NANDN U12881 ( .A(n12635), .B(n19883), .Z(n12586) );
  NANDN U12882 ( .A(n12584), .B(n19937), .Z(n12585) );
  AND U12883 ( .A(n12586), .B(n12585), .Z(n12639) );
  XNOR U12884 ( .A(n12638), .B(n12639), .Z(n12640) );
  XNOR U12885 ( .A(n12641), .B(n12640), .Z(n12677) );
  NANDN U12886 ( .A(n12588), .B(n12587), .Z(n12592) );
  NAND U12887 ( .A(n12590), .B(n12589), .Z(n12591) );
  NAND U12888 ( .A(n12592), .B(n12591), .Z(n12678) );
  XNOR U12889 ( .A(n12677), .B(n12678), .Z(n12679) );
  NANDN U12890 ( .A(n12594), .B(n12593), .Z(n12598) );
  NAND U12891 ( .A(n12596), .B(n12595), .Z(n12597) );
  AND U12892 ( .A(n12598), .B(n12597), .Z(n12680) );
  XNOR U12893 ( .A(n12679), .B(n12680), .Z(n12624) );
  XNOR U12894 ( .A(n12625), .B(n12624), .Z(n12683) );
  NANDN U12895 ( .A(n12600), .B(n12599), .Z(n12604) );
  NAND U12896 ( .A(n12602), .B(n12601), .Z(n12603) );
  NAND U12897 ( .A(n12604), .B(n12603), .Z(n12684) );
  XNOR U12898 ( .A(n12683), .B(n12684), .Z(n12685) );
  XOR U12899 ( .A(n12686), .B(n12685), .Z(n12616) );
  NANDN U12900 ( .A(n12606), .B(n12605), .Z(n12610) );
  NANDN U12901 ( .A(n12608), .B(n12607), .Z(n12609) );
  NAND U12902 ( .A(n12610), .B(n12609), .Z(n12617) );
  XNOR U12903 ( .A(n12616), .B(n12617), .Z(n12618) );
  XNOR U12904 ( .A(n12619), .B(n12618), .Z(n12689) );
  XNOR U12905 ( .A(n12689), .B(sreg[408]), .Z(n12691) );
  NAND U12906 ( .A(n12611), .B(sreg[407]), .Z(n12615) );
  OR U12907 ( .A(n12613), .B(n12612), .Z(n12614) );
  AND U12908 ( .A(n12615), .B(n12614), .Z(n12690) );
  XOR U12909 ( .A(n12691), .B(n12690), .Z(c[408]) );
  NANDN U12910 ( .A(n12617), .B(n12616), .Z(n12621) );
  NAND U12911 ( .A(n12619), .B(n12618), .Z(n12620) );
  NAND U12912 ( .A(n12621), .B(n12620), .Z(n12697) );
  NANDN U12913 ( .A(n12623), .B(n12622), .Z(n12627) );
  OR U12914 ( .A(n12625), .B(n12624), .Z(n12626) );
  NAND U12915 ( .A(n12627), .B(n12626), .Z(n12764) );
  XNOR U12916 ( .A(n20052), .B(n12943), .Z(n12733) );
  OR U12917 ( .A(n12733), .B(n20020), .Z(n12630) );
  NANDN U12918 ( .A(n12628), .B(n19960), .Z(n12629) );
  NAND U12919 ( .A(n12630), .B(n12629), .Z(n12746) );
  XNOR U12920 ( .A(n102), .B(n12631), .Z(n12737) );
  OR U12921 ( .A(n12737), .B(n20121), .Z(n12634) );
  NANDN U12922 ( .A(n12632), .B(n20122), .Z(n12633) );
  NAND U12923 ( .A(n12634), .B(n12633), .Z(n12743) );
  XNOR U12924 ( .A(n19975), .B(n13126), .Z(n12740) );
  NANDN U12925 ( .A(n12740), .B(n19883), .Z(n12637) );
  NANDN U12926 ( .A(n12635), .B(n19937), .Z(n12636) );
  AND U12927 ( .A(n12637), .B(n12636), .Z(n12744) );
  XNOR U12928 ( .A(n12743), .B(n12744), .Z(n12745) );
  XNOR U12929 ( .A(n12746), .B(n12745), .Z(n12755) );
  NANDN U12930 ( .A(n12639), .B(n12638), .Z(n12643) );
  NAND U12931 ( .A(n12641), .B(n12640), .Z(n12642) );
  NAND U12932 ( .A(n12643), .B(n12642), .Z(n12756) );
  XNOR U12933 ( .A(n12755), .B(n12756), .Z(n12757) );
  NANDN U12934 ( .A(n12645), .B(n12644), .Z(n12649) );
  NAND U12935 ( .A(n12647), .B(n12646), .Z(n12648) );
  AND U12936 ( .A(n12649), .B(n12648), .Z(n12758) );
  XNOR U12937 ( .A(n12757), .B(n12758), .Z(n12702) );
  NANDN U12938 ( .A(n12651), .B(n12650), .Z(n12655) );
  OR U12939 ( .A(n12653), .B(n12652), .Z(n12654) );
  NAND U12940 ( .A(n12655), .B(n12654), .Z(n12730) );
  NAND U12941 ( .A(b[0]), .B(a[169]), .Z(n12656) );
  XNOR U12942 ( .A(b[1]), .B(n12656), .Z(n12658) );
  NAND U12943 ( .A(a[168]), .B(n98), .Z(n12657) );
  AND U12944 ( .A(n12658), .B(n12657), .Z(n12706) );
  XNOR U12945 ( .A(n20154), .B(n12787), .Z(n12715) );
  OR U12946 ( .A(n12715), .B(n20057), .Z(n12661) );
  NANDN U12947 ( .A(n12659), .B(n20098), .Z(n12660) );
  AND U12948 ( .A(n12661), .B(n12660), .Z(n12707) );
  XOR U12949 ( .A(n12706), .B(n12707), .Z(n12709) );
  NAND U12950 ( .A(a[153]), .B(b[15]), .Z(n12708) );
  XOR U12951 ( .A(n12709), .B(n12708), .Z(n12727) );
  NAND U12952 ( .A(n19722), .B(n12662), .Z(n12664) );
  XNOR U12953 ( .A(b[5]), .B(n13438), .Z(n12718) );
  NANDN U12954 ( .A(n19640), .B(n12718), .Z(n12663) );
  NAND U12955 ( .A(n12664), .B(n12663), .Z(n12752) );
  XNOR U12956 ( .A(n19714), .B(n13282), .Z(n12721) );
  NANDN U12957 ( .A(n12721), .B(n19766), .Z(n12667) );
  NANDN U12958 ( .A(n12665), .B(n19767), .Z(n12666) );
  NAND U12959 ( .A(n12667), .B(n12666), .Z(n12749) );
  NAND U12960 ( .A(n19554), .B(n12668), .Z(n12670) );
  IV U12961 ( .A(a[167]), .Z(n13567) );
  XNOR U12962 ( .A(b[3]), .B(n13567), .Z(n12724) );
  NANDN U12963 ( .A(n19521), .B(n12724), .Z(n12669) );
  AND U12964 ( .A(n12670), .B(n12669), .Z(n12750) );
  XNOR U12965 ( .A(n12749), .B(n12750), .Z(n12751) );
  XOR U12966 ( .A(n12752), .B(n12751), .Z(n12728) );
  XOR U12967 ( .A(n12727), .B(n12728), .Z(n12729) );
  XNOR U12968 ( .A(n12730), .B(n12729), .Z(n12700) );
  NAND U12969 ( .A(n12672), .B(n12671), .Z(n12676) );
  NAND U12970 ( .A(n12674), .B(n12673), .Z(n12675) );
  NAND U12971 ( .A(n12676), .B(n12675), .Z(n12701) );
  XOR U12972 ( .A(n12700), .B(n12701), .Z(n12703) );
  XNOR U12973 ( .A(n12702), .B(n12703), .Z(n12761) );
  NANDN U12974 ( .A(n12678), .B(n12677), .Z(n12682) );
  NAND U12975 ( .A(n12680), .B(n12679), .Z(n12681) );
  NAND U12976 ( .A(n12682), .B(n12681), .Z(n12762) );
  XNOR U12977 ( .A(n12761), .B(n12762), .Z(n12763) );
  XOR U12978 ( .A(n12764), .B(n12763), .Z(n12694) );
  NANDN U12979 ( .A(n12684), .B(n12683), .Z(n12688) );
  NANDN U12980 ( .A(n12686), .B(n12685), .Z(n12687) );
  NAND U12981 ( .A(n12688), .B(n12687), .Z(n12695) );
  XNOR U12982 ( .A(n12694), .B(n12695), .Z(n12696) );
  XNOR U12983 ( .A(n12697), .B(n12696), .Z(n12767) );
  XNOR U12984 ( .A(n12767), .B(sreg[409]), .Z(n12769) );
  NAND U12985 ( .A(n12689), .B(sreg[408]), .Z(n12693) );
  OR U12986 ( .A(n12691), .B(n12690), .Z(n12692) );
  AND U12987 ( .A(n12693), .B(n12692), .Z(n12768) );
  XOR U12988 ( .A(n12769), .B(n12768), .Z(c[409]) );
  NANDN U12989 ( .A(n12695), .B(n12694), .Z(n12699) );
  NAND U12990 ( .A(n12697), .B(n12696), .Z(n12698) );
  NAND U12991 ( .A(n12699), .B(n12698), .Z(n12775) );
  NANDN U12992 ( .A(n12701), .B(n12700), .Z(n12705) );
  OR U12993 ( .A(n12703), .B(n12702), .Z(n12704) );
  NAND U12994 ( .A(n12705), .B(n12704), .Z(n12842) );
  NANDN U12995 ( .A(n12707), .B(n12706), .Z(n12711) );
  OR U12996 ( .A(n12709), .B(n12708), .Z(n12710) );
  NAND U12997 ( .A(n12711), .B(n12710), .Z(n12830) );
  NAND U12998 ( .A(b[0]), .B(a[170]), .Z(n12712) );
  XNOR U12999 ( .A(b[1]), .B(n12712), .Z(n12714) );
  NAND U13000 ( .A(a[169]), .B(n98), .Z(n12713) );
  AND U13001 ( .A(n12714), .B(n12713), .Z(n12806) );
  XNOR U13002 ( .A(n20154), .B(n12865), .Z(n12815) );
  OR U13003 ( .A(n12815), .B(n20057), .Z(n12717) );
  NANDN U13004 ( .A(n12715), .B(n20098), .Z(n12716) );
  AND U13005 ( .A(n12717), .B(n12716), .Z(n12807) );
  XOR U13006 ( .A(n12806), .B(n12807), .Z(n12809) );
  NAND U13007 ( .A(a[154]), .B(b[15]), .Z(n12808) );
  XOR U13008 ( .A(n12809), .B(n12808), .Z(n12827) );
  NAND U13009 ( .A(n19722), .B(n12718), .Z(n12720) );
  XNOR U13010 ( .A(b[5]), .B(n13516), .Z(n12818) );
  NANDN U13011 ( .A(n19640), .B(n12818), .Z(n12719) );
  NAND U13012 ( .A(n12720), .B(n12719), .Z(n12803) );
  XNOR U13013 ( .A(n19714), .B(n13333), .Z(n12821) );
  NANDN U13014 ( .A(n12821), .B(n19766), .Z(n12723) );
  NANDN U13015 ( .A(n12721), .B(n19767), .Z(n12722) );
  NAND U13016 ( .A(n12723), .B(n12722), .Z(n12800) );
  NAND U13017 ( .A(n19554), .B(n12724), .Z(n12726) );
  IV U13018 ( .A(a[168]), .Z(n13672) );
  XNOR U13019 ( .A(b[3]), .B(n13672), .Z(n12824) );
  NANDN U13020 ( .A(n19521), .B(n12824), .Z(n12725) );
  AND U13021 ( .A(n12726), .B(n12725), .Z(n12801) );
  XNOR U13022 ( .A(n12800), .B(n12801), .Z(n12802) );
  XOR U13023 ( .A(n12803), .B(n12802), .Z(n12828) );
  XOR U13024 ( .A(n12827), .B(n12828), .Z(n12829) );
  XNOR U13025 ( .A(n12830), .B(n12829), .Z(n12778) );
  NAND U13026 ( .A(n12728), .B(n12727), .Z(n12732) );
  NAND U13027 ( .A(n12730), .B(n12729), .Z(n12731) );
  NAND U13028 ( .A(n12732), .B(n12731), .Z(n12779) );
  XOR U13029 ( .A(n12778), .B(n12779), .Z(n12781) );
  XNOR U13030 ( .A(n20052), .B(n13021), .Z(n12784) );
  OR U13031 ( .A(n12784), .B(n20020), .Z(n12735) );
  NANDN U13032 ( .A(n12733), .B(n19960), .Z(n12734) );
  NAND U13033 ( .A(n12735), .B(n12734), .Z(n12797) );
  XNOR U13034 ( .A(n102), .B(n12736), .Z(n12788) );
  OR U13035 ( .A(n12788), .B(n20121), .Z(n12739) );
  NANDN U13036 ( .A(n12737), .B(n20122), .Z(n12738) );
  NAND U13037 ( .A(n12739), .B(n12738), .Z(n12794) );
  XNOR U13038 ( .A(n19975), .B(n13204), .Z(n12791) );
  NANDN U13039 ( .A(n12791), .B(n19883), .Z(n12742) );
  NANDN U13040 ( .A(n12740), .B(n19937), .Z(n12741) );
  AND U13041 ( .A(n12742), .B(n12741), .Z(n12795) );
  XNOR U13042 ( .A(n12794), .B(n12795), .Z(n12796) );
  XNOR U13043 ( .A(n12797), .B(n12796), .Z(n12833) );
  NANDN U13044 ( .A(n12744), .B(n12743), .Z(n12748) );
  NAND U13045 ( .A(n12746), .B(n12745), .Z(n12747) );
  NAND U13046 ( .A(n12748), .B(n12747), .Z(n12834) );
  XNOR U13047 ( .A(n12833), .B(n12834), .Z(n12835) );
  NANDN U13048 ( .A(n12750), .B(n12749), .Z(n12754) );
  NAND U13049 ( .A(n12752), .B(n12751), .Z(n12753) );
  AND U13050 ( .A(n12754), .B(n12753), .Z(n12836) );
  XNOR U13051 ( .A(n12835), .B(n12836), .Z(n12780) );
  XNOR U13052 ( .A(n12781), .B(n12780), .Z(n12839) );
  NANDN U13053 ( .A(n12756), .B(n12755), .Z(n12760) );
  NAND U13054 ( .A(n12758), .B(n12757), .Z(n12759) );
  NAND U13055 ( .A(n12760), .B(n12759), .Z(n12840) );
  XNOR U13056 ( .A(n12839), .B(n12840), .Z(n12841) );
  XOR U13057 ( .A(n12842), .B(n12841), .Z(n12772) );
  NANDN U13058 ( .A(n12762), .B(n12761), .Z(n12766) );
  NANDN U13059 ( .A(n12764), .B(n12763), .Z(n12765) );
  NAND U13060 ( .A(n12766), .B(n12765), .Z(n12773) );
  XNOR U13061 ( .A(n12772), .B(n12773), .Z(n12774) );
  XNOR U13062 ( .A(n12775), .B(n12774), .Z(n12845) );
  XNOR U13063 ( .A(n12845), .B(sreg[410]), .Z(n12847) );
  NAND U13064 ( .A(n12767), .B(sreg[409]), .Z(n12771) );
  OR U13065 ( .A(n12769), .B(n12768), .Z(n12770) );
  AND U13066 ( .A(n12771), .B(n12770), .Z(n12846) );
  XOR U13067 ( .A(n12847), .B(n12846), .Z(c[410]) );
  NANDN U13068 ( .A(n12773), .B(n12772), .Z(n12777) );
  NAND U13069 ( .A(n12775), .B(n12774), .Z(n12776) );
  NAND U13070 ( .A(n12777), .B(n12776), .Z(n12853) );
  NANDN U13071 ( .A(n12779), .B(n12778), .Z(n12783) );
  OR U13072 ( .A(n12781), .B(n12780), .Z(n12782) );
  NAND U13073 ( .A(n12783), .B(n12782), .Z(n12920) );
  XNOR U13074 ( .A(n20052), .B(n13126), .Z(n12862) );
  OR U13075 ( .A(n12862), .B(n20020), .Z(n12786) );
  NANDN U13076 ( .A(n12784), .B(n19960), .Z(n12785) );
  NAND U13077 ( .A(n12786), .B(n12785), .Z(n12875) );
  XNOR U13078 ( .A(n102), .B(n12787), .Z(n12866) );
  OR U13079 ( .A(n12866), .B(n20121), .Z(n12790) );
  NANDN U13080 ( .A(n12788), .B(n20122), .Z(n12789) );
  NAND U13081 ( .A(n12790), .B(n12789), .Z(n12872) );
  XNOR U13082 ( .A(n19975), .B(n13282), .Z(n12869) );
  NANDN U13083 ( .A(n12869), .B(n19883), .Z(n12793) );
  NANDN U13084 ( .A(n12791), .B(n19937), .Z(n12792) );
  AND U13085 ( .A(n12793), .B(n12792), .Z(n12873) );
  XNOR U13086 ( .A(n12872), .B(n12873), .Z(n12874) );
  XNOR U13087 ( .A(n12875), .B(n12874), .Z(n12911) );
  NANDN U13088 ( .A(n12795), .B(n12794), .Z(n12799) );
  NAND U13089 ( .A(n12797), .B(n12796), .Z(n12798) );
  NAND U13090 ( .A(n12799), .B(n12798), .Z(n12912) );
  XNOR U13091 ( .A(n12911), .B(n12912), .Z(n12913) );
  NANDN U13092 ( .A(n12801), .B(n12800), .Z(n12805) );
  NAND U13093 ( .A(n12803), .B(n12802), .Z(n12804) );
  AND U13094 ( .A(n12805), .B(n12804), .Z(n12914) );
  XNOR U13095 ( .A(n12913), .B(n12914), .Z(n12858) );
  NANDN U13096 ( .A(n12807), .B(n12806), .Z(n12811) );
  OR U13097 ( .A(n12809), .B(n12808), .Z(n12810) );
  NAND U13098 ( .A(n12811), .B(n12810), .Z(n12908) );
  NAND U13099 ( .A(b[0]), .B(a[171]), .Z(n12812) );
  XNOR U13100 ( .A(b[1]), .B(n12812), .Z(n12814) );
  NAND U13101 ( .A(a[170]), .B(n98), .Z(n12813) );
  AND U13102 ( .A(n12814), .B(n12813), .Z(n12884) );
  XNOR U13103 ( .A(n20154), .B(n12943), .Z(n12893) );
  OR U13104 ( .A(n12893), .B(n20057), .Z(n12817) );
  NANDN U13105 ( .A(n12815), .B(n20098), .Z(n12816) );
  AND U13106 ( .A(n12817), .B(n12816), .Z(n12885) );
  XOR U13107 ( .A(n12884), .B(n12885), .Z(n12887) );
  NAND U13108 ( .A(a[155]), .B(b[15]), .Z(n12886) );
  XOR U13109 ( .A(n12887), .B(n12886), .Z(n12905) );
  NAND U13110 ( .A(n19722), .B(n12818), .Z(n12820) );
  XNOR U13111 ( .A(b[5]), .B(n13567), .Z(n12896) );
  NANDN U13112 ( .A(n19640), .B(n12896), .Z(n12819) );
  NAND U13113 ( .A(n12820), .B(n12819), .Z(n12881) );
  XNOR U13114 ( .A(n19714), .B(n13438), .Z(n12899) );
  NANDN U13115 ( .A(n12899), .B(n19766), .Z(n12823) );
  NANDN U13116 ( .A(n12821), .B(n19767), .Z(n12822) );
  NAND U13117 ( .A(n12823), .B(n12822), .Z(n12878) );
  NAND U13118 ( .A(n19554), .B(n12824), .Z(n12826) );
  IV U13119 ( .A(a[169]), .Z(n13750) );
  XNOR U13120 ( .A(b[3]), .B(n13750), .Z(n12902) );
  NANDN U13121 ( .A(n19521), .B(n12902), .Z(n12825) );
  AND U13122 ( .A(n12826), .B(n12825), .Z(n12879) );
  XNOR U13123 ( .A(n12878), .B(n12879), .Z(n12880) );
  XOR U13124 ( .A(n12881), .B(n12880), .Z(n12906) );
  XOR U13125 ( .A(n12905), .B(n12906), .Z(n12907) );
  XNOR U13126 ( .A(n12908), .B(n12907), .Z(n12856) );
  NAND U13127 ( .A(n12828), .B(n12827), .Z(n12832) );
  NAND U13128 ( .A(n12830), .B(n12829), .Z(n12831) );
  NAND U13129 ( .A(n12832), .B(n12831), .Z(n12857) );
  XOR U13130 ( .A(n12856), .B(n12857), .Z(n12859) );
  XNOR U13131 ( .A(n12858), .B(n12859), .Z(n12917) );
  NANDN U13132 ( .A(n12834), .B(n12833), .Z(n12838) );
  NAND U13133 ( .A(n12836), .B(n12835), .Z(n12837) );
  NAND U13134 ( .A(n12838), .B(n12837), .Z(n12918) );
  XNOR U13135 ( .A(n12917), .B(n12918), .Z(n12919) );
  XOR U13136 ( .A(n12920), .B(n12919), .Z(n12850) );
  NANDN U13137 ( .A(n12840), .B(n12839), .Z(n12844) );
  NANDN U13138 ( .A(n12842), .B(n12841), .Z(n12843) );
  NAND U13139 ( .A(n12844), .B(n12843), .Z(n12851) );
  XNOR U13140 ( .A(n12850), .B(n12851), .Z(n12852) );
  XNOR U13141 ( .A(n12853), .B(n12852), .Z(n12923) );
  XNOR U13142 ( .A(n12923), .B(sreg[411]), .Z(n12925) );
  NAND U13143 ( .A(n12845), .B(sreg[410]), .Z(n12849) );
  OR U13144 ( .A(n12847), .B(n12846), .Z(n12848) );
  AND U13145 ( .A(n12849), .B(n12848), .Z(n12924) );
  XOR U13146 ( .A(n12925), .B(n12924), .Z(c[411]) );
  NANDN U13147 ( .A(n12851), .B(n12850), .Z(n12855) );
  NAND U13148 ( .A(n12853), .B(n12852), .Z(n12854) );
  NAND U13149 ( .A(n12855), .B(n12854), .Z(n12931) );
  NANDN U13150 ( .A(n12857), .B(n12856), .Z(n12861) );
  OR U13151 ( .A(n12859), .B(n12858), .Z(n12860) );
  NAND U13152 ( .A(n12861), .B(n12860), .Z(n12998) );
  XNOR U13153 ( .A(n20052), .B(n13204), .Z(n12940) );
  OR U13154 ( .A(n12940), .B(n20020), .Z(n12864) );
  NANDN U13155 ( .A(n12862), .B(n19960), .Z(n12863) );
  NAND U13156 ( .A(n12864), .B(n12863), .Z(n12953) );
  XNOR U13157 ( .A(n102), .B(n12865), .Z(n12944) );
  OR U13158 ( .A(n12944), .B(n20121), .Z(n12868) );
  NANDN U13159 ( .A(n12866), .B(n20122), .Z(n12867) );
  NAND U13160 ( .A(n12868), .B(n12867), .Z(n12950) );
  XNOR U13161 ( .A(n19975), .B(n13333), .Z(n12947) );
  NANDN U13162 ( .A(n12947), .B(n19883), .Z(n12871) );
  NANDN U13163 ( .A(n12869), .B(n19937), .Z(n12870) );
  AND U13164 ( .A(n12871), .B(n12870), .Z(n12951) );
  XNOR U13165 ( .A(n12950), .B(n12951), .Z(n12952) );
  XNOR U13166 ( .A(n12953), .B(n12952), .Z(n12989) );
  NANDN U13167 ( .A(n12873), .B(n12872), .Z(n12877) );
  NAND U13168 ( .A(n12875), .B(n12874), .Z(n12876) );
  NAND U13169 ( .A(n12877), .B(n12876), .Z(n12990) );
  XNOR U13170 ( .A(n12989), .B(n12990), .Z(n12991) );
  NANDN U13171 ( .A(n12879), .B(n12878), .Z(n12883) );
  NAND U13172 ( .A(n12881), .B(n12880), .Z(n12882) );
  AND U13173 ( .A(n12883), .B(n12882), .Z(n12992) );
  XNOR U13174 ( .A(n12991), .B(n12992), .Z(n12936) );
  NANDN U13175 ( .A(n12885), .B(n12884), .Z(n12889) );
  OR U13176 ( .A(n12887), .B(n12886), .Z(n12888) );
  NAND U13177 ( .A(n12889), .B(n12888), .Z(n12986) );
  NAND U13178 ( .A(b[0]), .B(a[172]), .Z(n12890) );
  XNOR U13179 ( .A(b[1]), .B(n12890), .Z(n12892) );
  NAND U13180 ( .A(a[171]), .B(n98), .Z(n12891) );
  AND U13181 ( .A(n12892), .B(n12891), .Z(n12962) );
  XNOR U13182 ( .A(n20154), .B(n13021), .Z(n12968) );
  OR U13183 ( .A(n12968), .B(n20057), .Z(n12895) );
  NANDN U13184 ( .A(n12893), .B(n20098), .Z(n12894) );
  AND U13185 ( .A(n12895), .B(n12894), .Z(n12963) );
  XOR U13186 ( .A(n12962), .B(n12963), .Z(n12965) );
  NAND U13187 ( .A(a[156]), .B(b[15]), .Z(n12964) );
  XOR U13188 ( .A(n12965), .B(n12964), .Z(n12983) );
  NAND U13189 ( .A(n19722), .B(n12896), .Z(n12898) );
  XNOR U13190 ( .A(b[5]), .B(n13672), .Z(n12974) );
  NANDN U13191 ( .A(n19640), .B(n12974), .Z(n12897) );
  NAND U13192 ( .A(n12898), .B(n12897), .Z(n12959) );
  XNOR U13193 ( .A(n19714), .B(n13516), .Z(n12977) );
  NANDN U13194 ( .A(n12977), .B(n19766), .Z(n12901) );
  NANDN U13195 ( .A(n12899), .B(n19767), .Z(n12900) );
  NAND U13196 ( .A(n12901), .B(n12900), .Z(n12956) );
  NAND U13197 ( .A(n19554), .B(n12902), .Z(n12904) );
  IV U13198 ( .A(a[170]), .Z(n13801) );
  XNOR U13199 ( .A(b[3]), .B(n13801), .Z(n12980) );
  NANDN U13200 ( .A(n19521), .B(n12980), .Z(n12903) );
  AND U13201 ( .A(n12904), .B(n12903), .Z(n12957) );
  XNOR U13202 ( .A(n12956), .B(n12957), .Z(n12958) );
  XOR U13203 ( .A(n12959), .B(n12958), .Z(n12984) );
  XOR U13204 ( .A(n12983), .B(n12984), .Z(n12985) );
  XNOR U13205 ( .A(n12986), .B(n12985), .Z(n12934) );
  NAND U13206 ( .A(n12906), .B(n12905), .Z(n12910) );
  NAND U13207 ( .A(n12908), .B(n12907), .Z(n12909) );
  NAND U13208 ( .A(n12910), .B(n12909), .Z(n12935) );
  XOR U13209 ( .A(n12934), .B(n12935), .Z(n12937) );
  XNOR U13210 ( .A(n12936), .B(n12937), .Z(n12995) );
  NANDN U13211 ( .A(n12912), .B(n12911), .Z(n12916) );
  NAND U13212 ( .A(n12914), .B(n12913), .Z(n12915) );
  NAND U13213 ( .A(n12916), .B(n12915), .Z(n12996) );
  XNOR U13214 ( .A(n12995), .B(n12996), .Z(n12997) );
  XOR U13215 ( .A(n12998), .B(n12997), .Z(n12928) );
  NANDN U13216 ( .A(n12918), .B(n12917), .Z(n12922) );
  NANDN U13217 ( .A(n12920), .B(n12919), .Z(n12921) );
  NAND U13218 ( .A(n12922), .B(n12921), .Z(n12929) );
  XNOR U13219 ( .A(n12928), .B(n12929), .Z(n12930) );
  XNOR U13220 ( .A(n12931), .B(n12930), .Z(n13001) );
  XNOR U13221 ( .A(n13001), .B(sreg[412]), .Z(n13003) );
  NAND U13222 ( .A(n12923), .B(sreg[411]), .Z(n12927) );
  OR U13223 ( .A(n12925), .B(n12924), .Z(n12926) );
  AND U13224 ( .A(n12927), .B(n12926), .Z(n13002) );
  XOR U13225 ( .A(n13003), .B(n13002), .Z(c[412]) );
  NANDN U13226 ( .A(n12929), .B(n12928), .Z(n12933) );
  NAND U13227 ( .A(n12931), .B(n12930), .Z(n12932) );
  NAND U13228 ( .A(n12933), .B(n12932), .Z(n13009) );
  NANDN U13229 ( .A(n12935), .B(n12934), .Z(n12939) );
  OR U13230 ( .A(n12937), .B(n12936), .Z(n12938) );
  NAND U13231 ( .A(n12939), .B(n12938), .Z(n13076) );
  XNOR U13232 ( .A(n20052), .B(n13282), .Z(n13018) );
  OR U13233 ( .A(n13018), .B(n20020), .Z(n12942) );
  NANDN U13234 ( .A(n12940), .B(n19960), .Z(n12941) );
  NAND U13235 ( .A(n12942), .B(n12941), .Z(n13031) );
  XNOR U13236 ( .A(n102), .B(n12943), .Z(n13022) );
  OR U13237 ( .A(n13022), .B(n20121), .Z(n12946) );
  NANDN U13238 ( .A(n12944), .B(n20122), .Z(n12945) );
  NAND U13239 ( .A(n12946), .B(n12945), .Z(n13028) );
  XNOR U13240 ( .A(n19975), .B(n13438), .Z(n13025) );
  NANDN U13241 ( .A(n13025), .B(n19883), .Z(n12949) );
  NANDN U13242 ( .A(n12947), .B(n19937), .Z(n12948) );
  AND U13243 ( .A(n12949), .B(n12948), .Z(n13029) );
  XNOR U13244 ( .A(n13028), .B(n13029), .Z(n13030) );
  XNOR U13245 ( .A(n13031), .B(n13030), .Z(n13067) );
  NANDN U13246 ( .A(n12951), .B(n12950), .Z(n12955) );
  NAND U13247 ( .A(n12953), .B(n12952), .Z(n12954) );
  NAND U13248 ( .A(n12955), .B(n12954), .Z(n13068) );
  XNOR U13249 ( .A(n13067), .B(n13068), .Z(n13069) );
  NANDN U13250 ( .A(n12957), .B(n12956), .Z(n12961) );
  NAND U13251 ( .A(n12959), .B(n12958), .Z(n12960) );
  AND U13252 ( .A(n12961), .B(n12960), .Z(n13070) );
  XNOR U13253 ( .A(n13069), .B(n13070), .Z(n13014) );
  NANDN U13254 ( .A(n12963), .B(n12962), .Z(n12967) );
  OR U13255 ( .A(n12965), .B(n12964), .Z(n12966) );
  NAND U13256 ( .A(n12967), .B(n12966), .Z(n13064) );
  XNOR U13257 ( .A(n20154), .B(n13126), .Z(n13049) );
  OR U13258 ( .A(n13049), .B(n20057), .Z(n12970) );
  NANDN U13259 ( .A(n12968), .B(n20098), .Z(n12969) );
  AND U13260 ( .A(n12970), .B(n12969), .Z(n13041) );
  NAND U13261 ( .A(b[0]), .B(a[173]), .Z(n12971) );
  XNOR U13262 ( .A(b[1]), .B(n12971), .Z(n12973) );
  NAND U13263 ( .A(a[172]), .B(n98), .Z(n12972) );
  AND U13264 ( .A(n12973), .B(n12972), .Z(n13040) );
  XOR U13265 ( .A(n13041), .B(n13040), .Z(n13043) );
  NAND U13266 ( .A(a[157]), .B(b[15]), .Z(n13042) );
  XOR U13267 ( .A(n13043), .B(n13042), .Z(n13061) );
  NAND U13268 ( .A(n19722), .B(n12974), .Z(n12976) );
  XNOR U13269 ( .A(b[5]), .B(n13750), .Z(n13052) );
  NANDN U13270 ( .A(n19640), .B(n13052), .Z(n12975) );
  NAND U13271 ( .A(n12976), .B(n12975), .Z(n13037) );
  XNOR U13272 ( .A(n19714), .B(n13567), .Z(n13055) );
  NANDN U13273 ( .A(n13055), .B(n19766), .Z(n12979) );
  NANDN U13274 ( .A(n12977), .B(n19767), .Z(n12978) );
  NAND U13275 ( .A(n12979), .B(n12978), .Z(n13034) );
  NAND U13276 ( .A(n19554), .B(n12980), .Z(n12982) );
  IV U13277 ( .A(a[171]), .Z(n13906) );
  XNOR U13278 ( .A(b[3]), .B(n13906), .Z(n13058) );
  NANDN U13279 ( .A(n19521), .B(n13058), .Z(n12981) );
  AND U13280 ( .A(n12982), .B(n12981), .Z(n13035) );
  XNOR U13281 ( .A(n13034), .B(n13035), .Z(n13036) );
  XOR U13282 ( .A(n13037), .B(n13036), .Z(n13062) );
  XOR U13283 ( .A(n13061), .B(n13062), .Z(n13063) );
  XNOR U13284 ( .A(n13064), .B(n13063), .Z(n13012) );
  NAND U13285 ( .A(n12984), .B(n12983), .Z(n12988) );
  NAND U13286 ( .A(n12986), .B(n12985), .Z(n12987) );
  NAND U13287 ( .A(n12988), .B(n12987), .Z(n13013) );
  XOR U13288 ( .A(n13012), .B(n13013), .Z(n13015) );
  XNOR U13289 ( .A(n13014), .B(n13015), .Z(n13073) );
  NANDN U13290 ( .A(n12990), .B(n12989), .Z(n12994) );
  NAND U13291 ( .A(n12992), .B(n12991), .Z(n12993) );
  NAND U13292 ( .A(n12994), .B(n12993), .Z(n13074) );
  XNOR U13293 ( .A(n13073), .B(n13074), .Z(n13075) );
  XOR U13294 ( .A(n13076), .B(n13075), .Z(n13006) );
  NANDN U13295 ( .A(n12996), .B(n12995), .Z(n13000) );
  NANDN U13296 ( .A(n12998), .B(n12997), .Z(n12999) );
  NAND U13297 ( .A(n13000), .B(n12999), .Z(n13007) );
  XNOR U13298 ( .A(n13006), .B(n13007), .Z(n13008) );
  XNOR U13299 ( .A(n13009), .B(n13008), .Z(n13079) );
  XNOR U13300 ( .A(n13079), .B(sreg[413]), .Z(n13081) );
  NAND U13301 ( .A(n13001), .B(sreg[412]), .Z(n13005) );
  OR U13302 ( .A(n13003), .B(n13002), .Z(n13004) );
  AND U13303 ( .A(n13005), .B(n13004), .Z(n13080) );
  XOR U13304 ( .A(n13081), .B(n13080), .Z(c[413]) );
  NANDN U13305 ( .A(n13007), .B(n13006), .Z(n13011) );
  NAND U13306 ( .A(n13009), .B(n13008), .Z(n13010) );
  NAND U13307 ( .A(n13011), .B(n13010), .Z(n13087) );
  NANDN U13308 ( .A(n13013), .B(n13012), .Z(n13017) );
  OR U13309 ( .A(n13015), .B(n13014), .Z(n13016) );
  NAND U13310 ( .A(n13017), .B(n13016), .Z(n13154) );
  XNOR U13311 ( .A(n20052), .B(n13333), .Z(n13123) );
  OR U13312 ( .A(n13123), .B(n20020), .Z(n13020) );
  NANDN U13313 ( .A(n13018), .B(n19960), .Z(n13019) );
  NAND U13314 ( .A(n13020), .B(n13019), .Z(n13136) );
  XNOR U13315 ( .A(n102), .B(n13021), .Z(n13127) );
  OR U13316 ( .A(n13127), .B(n20121), .Z(n13024) );
  NANDN U13317 ( .A(n13022), .B(n20122), .Z(n13023) );
  NAND U13318 ( .A(n13024), .B(n13023), .Z(n13133) );
  XNOR U13319 ( .A(n19975), .B(n13516), .Z(n13130) );
  NANDN U13320 ( .A(n13130), .B(n19883), .Z(n13027) );
  NANDN U13321 ( .A(n13025), .B(n19937), .Z(n13026) );
  AND U13322 ( .A(n13027), .B(n13026), .Z(n13134) );
  XNOR U13323 ( .A(n13133), .B(n13134), .Z(n13135) );
  XNOR U13324 ( .A(n13136), .B(n13135), .Z(n13145) );
  NANDN U13325 ( .A(n13029), .B(n13028), .Z(n13033) );
  NAND U13326 ( .A(n13031), .B(n13030), .Z(n13032) );
  NAND U13327 ( .A(n13033), .B(n13032), .Z(n13146) );
  XNOR U13328 ( .A(n13145), .B(n13146), .Z(n13147) );
  NANDN U13329 ( .A(n13035), .B(n13034), .Z(n13039) );
  NAND U13330 ( .A(n13037), .B(n13036), .Z(n13038) );
  AND U13331 ( .A(n13039), .B(n13038), .Z(n13148) );
  XNOR U13332 ( .A(n13147), .B(n13148), .Z(n13092) );
  NANDN U13333 ( .A(n13041), .B(n13040), .Z(n13045) );
  OR U13334 ( .A(n13043), .B(n13042), .Z(n13044) );
  NAND U13335 ( .A(n13045), .B(n13044), .Z(n13120) );
  NAND U13336 ( .A(b[0]), .B(a[174]), .Z(n13046) );
  XNOR U13337 ( .A(b[1]), .B(n13046), .Z(n13048) );
  NAND U13338 ( .A(a[173]), .B(n98), .Z(n13047) );
  AND U13339 ( .A(n13048), .B(n13047), .Z(n13096) );
  XNOR U13340 ( .A(n20154), .B(n13204), .Z(n13102) );
  OR U13341 ( .A(n13102), .B(n20057), .Z(n13051) );
  NANDN U13342 ( .A(n13049), .B(n20098), .Z(n13050) );
  AND U13343 ( .A(n13051), .B(n13050), .Z(n13097) );
  XOR U13344 ( .A(n13096), .B(n13097), .Z(n13099) );
  NAND U13345 ( .A(a[158]), .B(b[15]), .Z(n13098) );
  XOR U13346 ( .A(n13099), .B(n13098), .Z(n13117) );
  NAND U13347 ( .A(n19722), .B(n13052), .Z(n13054) );
  XNOR U13348 ( .A(b[5]), .B(n13801), .Z(n13108) );
  NANDN U13349 ( .A(n19640), .B(n13108), .Z(n13053) );
  NAND U13350 ( .A(n13054), .B(n13053), .Z(n13142) );
  XNOR U13351 ( .A(n19714), .B(n13672), .Z(n13111) );
  NANDN U13352 ( .A(n13111), .B(n19766), .Z(n13057) );
  NANDN U13353 ( .A(n13055), .B(n19767), .Z(n13056) );
  NAND U13354 ( .A(n13057), .B(n13056), .Z(n13139) );
  NAND U13355 ( .A(n19554), .B(n13058), .Z(n13060) );
  IV U13356 ( .A(a[172]), .Z(n13984) );
  XNOR U13357 ( .A(b[3]), .B(n13984), .Z(n13114) );
  NANDN U13358 ( .A(n19521), .B(n13114), .Z(n13059) );
  AND U13359 ( .A(n13060), .B(n13059), .Z(n13140) );
  XNOR U13360 ( .A(n13139), .B(n13140), .Z(n13141) );
  XOR U13361 ( .A(n13142), .B(n13141), .Z(n13118) );
  XOR U13362 ( .A(n13117), .B(n13118), .Z(n13119) );
  XNOR U13363 ( .A(n13120), .B(n13119), .Z(n13090) );
  NAND U13364 ( .A(n13062), .B(n13061), .Z(n13066) );
  NAND U13365 ( .A(n13064), .B(n13063), .Z(n13065) );
  NAND U13366 ( .A(n13066), .B(n13065), .Z(n13091) );
  XOR U13367 ( .A(n13090), .B(n13091), .Z(n13093) );
  XNOR U13368 ( .A(n13092), .B(n13093), .Z(n13151) );
  NANDN U13369 ( .A(n13068), .B(n13067), .Z(n13072) );
  NAND U13370 ( .A(n13070), .B(n13069), .Z(n13071) );
  NAND U13371 ( .A(n13072), .B(n13071), .Z(n13152) );
  XNOR U13372 ( .A(n13151), .B(n13152), .Z(n13153) );
  XOR U13373 ( .A(n13154), .B(n13153), .Z(n13084) );
  NANDN U13374 ( .A(n13074), .B(n13073), .Z(n13078) );
  NANDN U13375 ( .A(n13076), .B(n13075), .Z(n13077) );
  NAND U13376 ( .A(n13078), .B(n13077), .Z(n13085) );
  XNOR U13377 ( .A(n13084), .B(n13085), .Z(n13086) );
  XNOR U13378 ( .A(n13087), .B(n13086), .Z(n13157) );
  XNOR U13379 ( .A(n13157), .B(sreg[414]), .Z(n13159) );
  NAND U13380 ( .A(n13079), .B(sreg[413]), .Z(n13083) );
  OR U13381 ( .A(n13081), .B(n13080), .Z(n13082) );
  AND U13382 ( .A(n13083), .B(n13082), .Z(n13158) );
  XOR U13383 ( .A(n13159), .B(n13158), .Z(c[414]) );
  NANDN U13384 ( .A(n13085), .B(n13084), .Z(n13089) );
  NAND U13385 ( .A(n13087), .B(n13086), .Z(n13088) );
  NAND U13386 ( .A(n13089), .B(n13088), .Z(n13165) );
  NANDN U13387 ( .A(n13091), .B(n13090), .Z(n13095) );
  OR U13388 ( .A(n13093), .B(n13092), .Z(n13094) );
  NAND U13389 ( .A(n13095), .B(n13094), .Z(n13232) );
  NANDN U13390 ( .A(n13097), .B(n13096), .Z(n13101) );
  OR U13391 ( .A(n13099), .B(n13098), .Z(n13100) );
  NAND U13392 ( .A(n13101), .B(n13100), .Z(n13198) );
  XNOR U13393 ( .A(n20154), .B(n13282), .Z(n13183) );
  OR U13394 ( .A(n13183), .B(n20057), .Z(n13104) );
  NANDN U13395 ( .A(n13102), .B(n20098), .Z(n13103) );
  AND U13396 ( .A(n13104), .B(n13103), .Z(n13175) );
  NAND U13397 ( .A(b[0]), .B(a[175]), .Z(n13105) );
  XNOR U13398 ( .A(b[1]), .B(n13105), .Z(n13107) );
  NAND U13399 ( .A(a[174]), .B(n98), .Z(n13106) );
  AND U13400 ( .A(n13107), .B(n13106), .Z(n13174) );
  XOR U13401 ( .A(n13175), .B(n13174), .Z(n13177) );
  NAND U13402 ( .A(a[159]), .B(b[15]), .Z(n13176) );
  XOR U13403 ( .A(n13177), .B(n13176), .Z(n13195) );
  NAND U13404 ( .A(n19722), .B(n13108), .Z(n13110) );
  XNOR U13405 ( .A(b[5]), .B(n13906), .Z(n13186) );
  NANDN U13406 ( .A(n19640), .B(n13186), .Z(n13109) );
  NAND U13407 ( .A(n13110), .B(n13109), .Z(n13220) );
  XNOR U13408 ( .A(n19714), .B(n13750), .Z(n13189) );
  NANDN U13409 ( .A(n13189), .B(n19766), .Z(n13113) );
  NANDN U13410 ( .A(n13111), .B(n19767), .Z(n13112) );
  NAND U13411 ( .A(n13113), .B(n13112), .Z(n13217) );
  NAND U13412 ( .A(n19554), .B(n13114), .Z(n13116) );
  IV U13413 ( .A(a[173]), .Z(n14062) );
  XNOR U13414 ( .A(b[3]), .B(n14062), .Z(n13192) );
  NANDN U13415 ( .A(n19521), .B(n13192), .Z(n13115) );
  AND U13416 ( .A(n13116), .B(n13115), .Z(n13218) );
  XNOR U13417 ( .A(n13217), .B(n13218), .Z(n13219) );
  XOR U13418 ( .A(n13220), .B(n13219), .Z(n13196) );
  XOR U13419 ( .A(n13195), .B(n13196), .Z(n13197) );
  XNOR U13420 ( .A(n13198), .B(n13197), .Z(n13168) );
  NAND U13421 ( .A(n13118), .B(n13117), .Z(n13122) );
  NAND U13422 ( .A(n13120), .B(n13119), .Z(n13121) );
  NAND U13423 ( .A(n13122), .B(n13121), .Z(n13169) );
  XOR U13424 ( .A(n13168), .B(n13169), .Z(n13171) );
  XNOR U13425 ( .A(n20052), .B(n13438), .Z(n13201) );
  OR U13426 ( .A(n13201), .B(n20020), .Z(n13125) );
  NANDN U13427 ( .A(n13123), .B(n19960), .Z(n13124) );
  NAND U13428 ( .A(n13125), .B(n13124), .Z(n13214) );
  XNOR U13429 ( .A(n102), .B(n13126), .Z(n13205) );
  OR U13430 ( .A(n13205), .B(n20121), .Z(n13129) );
  NANDN U13431 ( .A(n13127), .B(n20122), .Z(n13128) );
  NAND U13432 ( .A(n13129), .B(n13128), .Z(n13211) );
  XNOR U13433 ( .A(n19975), .B(n13567), .Z(n13208) );
  NANDN U13434 ( .A(n13208), .B(n19883), .Z(n13132) );
  NANDN U13435 ( .A(n13130), .B(n19937), .Z(n13131) );
  AND U13436 ( .A(n13132), .B(n13131), .Z(n13212) );
  XNOR U13437 ( .A(n13211), .B(n13212), .Z(n13213) );
  XNOR U13438 ( .A(n13214), .B(n13213), .Z(n13223) );
  NANDN U13439 ( .A(n13134), .B(n13133), .Z(n13138) );
  NAND U13440 ( .A(n13136), .B(n13135), .Z(n13137) );
  NAND U13441 ( .A(n13138), .B(n13137), .Z(n13224) );
  XNOR U13442 ( .A(n13223), .B(n13224), .Z(n13225) );
  NANDN U13443 ( .A(n13140), .B(n13139), .Z(n13144) );
  NAND U13444 ( .A(n13142), .B(n13141), .Z(n13143) );
  AND U13445 ( .A(n13144), .B(n13143), .Z(n13226) );
  XNOR U13446 ( .A(n13225), .B(n13226), .Z(n13170) );
  XNOR U13447 ( .A(n13171), .B(n13170), .Z(n13229) );
  NANDN U13448 ( .A(n13146), .B(n13145), .Z(n13150) );
  NAND U13449 ( .A(n13148), .B(n13147), .Z(n13149) );
  NAND U13450 ( .A(n13150), .B(n13149), .Z(n13230) );
  XNOR U13451 ( .A(n13229), .B(n13230), .Z(n13231) );
  XOR U13452 ( .A(n13232), .B(n13231), .Z(n13162) );
  NANDN U13453 ( .A(n13152), .B(n13151), .Z(n13156) );
  NANDN U13454 ( .A(n13154), .B(n13153), .Z(n13155) );
  NAND U13455 ( .A(n13156), .B(n13155), .Z(n13163) );
  XNOR U13456 ( .A(n13162), .B(n13163), .Z(n13164) );
  XNOR U13457 ( .A(n13165), .B(n13164), .Z(n13235) );
  XNOR U13458 ( .A(n13235), .B(sreg[415]), .Z(n13237) );
  NAND U13459 ( .A(n13157), .B(sreg[414]), .Z(n13161) );
  OR U13460 ( .A(n13159), .B(n13158), .Z(n13160) );
  AND U13461 ( .A(n13161), .B(n13160), .Z(n13236) );
  XOR U13462 ( .A(n13237), .B(n13236), .Z(c[415]) );
  NANDN U13463 ( .A(n13163), .B(n13162), .Z(n13167) );
  NAND U13464 ( .A(n13165), .B(n13164), .Z(n13166) );
  NAND U13465 ( .A(n13167), .B(n13166), .Z(n13243) );
  NANDN U13466 ( .A(n13169), .B(n13168), .Z(n13173) );
  OR U13467 ( .A(n13171), .B(n13170), .Z(n13172) );
  NAND U13468 ( .A(n13173), .B(n13172), .Z(n13310) );
  NANDN U13469 ( .A(n13175), .B(n13174), .Z(n13179) );
  OR U13470 ( .A(n13177), .B(n13176), .Z(n13178) );
  NAND U13471 ( .A(n13179), .B(n13178), .Z(n13276) );
  NAND U13472 ( .A(b[0]), .B(a[176]), .Z(n13180) );
  XNOR U13473 ( .A(b[1]), .B(n13180), .Z(n13182) );
  NAND U13474 ( .A(a[175]), .B(n98), .Z(n13181) );
  AND U13475 ( .A(n13182), .B(n13181), .Z(n13252) );
  XNOR U13476 ( .A(n20154), .B(n13333), .Z(n13261) );
  OR U13477 ( .A(n13261), .B(n20057), .Z(n13185) );
  NANDN U13478 ( .A(n13183), .B(n20098), .Z(n13184) );
  AND U13479 ( .A(n13185), .B(n13184), .Z(n13253) );
  XOR U13480 ( .A(n13252), .B(n13253), .Z(n13255) );
  NAND U13481 ( .A(a[160]), .B(b[15]), .Z(n13254) );
  XOR U13482 ( .A(n13255), .B(n13254), .Z(n13273) );
  NAND U13483 ( .A(n19722), .B(n13186), .Z(n13188) );
  XNOR U13484 ( .A(b[5]), .B(n13984), .Z(n13264) );
  NANDN U13485 ( .A(n19640), .B(n13264), .Z(n13187) );
  NAND U13486 ( .A(n13188), .B(n13187), .Z(n13298) );
  XNOR U13487 ( .A(n19714), .B(n13801), .Z(n13267) );
  NANDN U13488 ( .A(n13267), .B(n19766), .Z(n13191) );
  NANDN U13489 ( .A(n13189), .B(n19767), .Z(n13190) );
  NAND U13490 ( .A(n13191), .B(n13190), .Z(n13295) );
  NAND U13491 ( .A(n19554), .B(n13192), .Z(n13194) );
  IV U13492 ( .A(a[174]), .Z(n14113) );
  XNOR U13493 ( .A(b[3]), .B(n14113), .Z(n13270) );
  NANDN U13494 ( .A(n19521), .B(n13270), .Z(n13193) );
  AND U13495 ( .A(n13194), .B(n13193), .Z(n13296) );
  XNOR U13496 ( .A(n13295), .B(n13296), .Z(n13297) );
  XOR U13497 ( .A(n13298), .B(n13297), .Z(n13274) );
  XOR U13498 ( .A(n13273), .B(n13274), .Z(n13275) );
  XNOR U13499 ( .A(n13276), .B(n13275), .Z(n13246) );
  NAND U13500 ( .A(n13196), .B(n13195), .Z(n13200) );
  NAND U13501 ( .A(n13198), .B(n13197), .Z(n13199) );
  NAND U13502 ( .A(n13200), .B(n13199), .Z(n13247) );
  XOR U13503 ( .A(n13246), .B(n13247), .Z(n13249) );
  XNOR U13504 ( .A(n20052), .B(n13516), .Z(n13279) );
  OR U13505 ( .A(n13279), .B(n20020), .Z(n13203) );
  NANDN U13506 ( .A(n13201), .B(n19960), .Z(n13202) );
  NAND U13507 ( .A(n13203), .B(n13202), .Z(n13292) );
  XNOR U13508 ( .A(n102), .B(n13204), .Z(n13283) );
  OR U13509 ( .A(n13283), .B(n20121), .Z(n13207) );
  NANDN U13510 ( .A(n13205), .B(n20122), .Z(n13206) );
  NAND U13511 ( .A(n13207), .B(n13206), .Z(n13289) );
  XNOR U13512 ( .A(n19975), .B(n13672), .Z(n13286) );
  NANDN U13513 ( .A(n13286), .B(n19883), .Z(n13210) );
  NANDN U13514 ( .A(n13208), .B(n19937), .Z(n13209) );
  AND U13515 ( .A(n13210), .B(n13209), .Z(n13290) );
  XNOR U13516 ( .A(n13289), .B(n13290), .Z(n13291) );
  XNOR U13517 ( .A(n13292), .B(n13291), .Z(n13301) );
  NANDN U13518 ( .A(n13212), .B(n13211), .Z(n13216) );
  NAND U13519 ( .A(n13214), .B(n13213), .Z(n13215) );
  NAND U13520 ( .A(n13216), .B(n13215), .Z(n13302) );
  XNOR U13521 ( .A(n13301), .B(n13302), .Z(n13303) );
  NANDN U13522 ( .A(n13218), .B(n13217), .Z(n13222) );
  NAND U13523 ( .A(n13220), .B(n13219), .Z(n13221) );
  AND U13524 ( .A(n13222), .B(n13221), .Z(n13304) );
  XNOR U13525 ( .A(n13303), .B(n13304), .Z(n13248) );
  XNOR U13526 ( .A(n13249), .B(n13248), .Z(n13307) );
  NANDN U13527 ( .A(n13224), .B(n13223), .Z(n13228) );
  NAND U13528 ( .A(n13226), .B(n13225), .Z(n13227) );
  NAND U13529 ( .A(n13228), .B(n13227), .Z(n13308) );
  XNOR U13530 ( .A(n13307), .B(n13308), .Z(n13309) );
  XOR U13531 ( .A(n13310), .B(n13309), .Z(n13240) );
  NANDN U13532 ( .A(n13230), .B(n13229), .Z(n13234) );
  NANDN U13533 ( .A(n13232), .B(n13231), .Z(n13233) );
  NAND U13534 ( .A(n13234), .B(n13233), .Z(n13241) );
  XNOR U13535 ( .A(n13240), .B(n13241), .Z(n13242) );
  XNOR U13536 ( .A(n13243), .B(n13242), .Z(n13313) );
  XNOR U13537 ( .A(n13313), .B(sreg[416]), .Z(n13315) );
  NAND U13538 ( .A(n13235), .B(sreg[415]), .Z(n13239) );
  OR U13539 ( .A(n13237), .B(n13236), .Z(n13238) );
  AND U13540 ( .A(n13239), .B(n13238), .Z(n13314) );
  XOR U13541 ( .A(n13315), .B(n13314), .Z(c[416]) );
  NANDN U13542 ( .A(n13241), .B(n13240), .Z(n13245) );
  NAND U13543 ( .A(n13243), .B(n13242), .Z(n13244) );
  NAND U13544 ( .A(n13245), .B(n13244), .Z(n13321) );
  NANDN U13545 ( .A(n13247), .B(n13246), .Z(n13251) );
  OR U13546 ( .A(n13249), .B(n13248), .Z(n13250) );
  NAND U13547 ( .A(n13251), .B(n13250), .Z(n13388) );
  NANDN U13548 ( .A(n13253), .B(n13252), .Z(n13257) );
  OR U13549 ( .A(n13255), .B(n13254), .Z(n13256) );
  NAND U13550 ( .A(n13257), .B(n13256), .Z(n13376) );
  NAND U13551 ( .A(b[0]), .B(a[177]), .Z(n13258) );
  XNOR U13552 ( .A(b[1]), .B(n13258), .Z(n13260) );
  NAND U13553 ( .A(a[176]), .B(n98), .Z(n13259) );
  AND U13554 ( .A(n13260), .B(n13259), .Z(n13352) );
  XNOR U13555 ( .A(n20154), .B(n13438), .Z(n13361) );
  OR U13556 ( .A(n13361), .B(n20057), .Z(n13263) );
  NANDN U13557 ( .A(n13261), .B(n20098), .Z(n13262) );
  AND U13558 ( .A(n13263), .B(n13262), .Z(n13353) );
  XOR U13559 ( .A(n13352), .B(n13353), .Z(n13355) );
  NAND U13560 ( .A(a[161]), .B(b[15]), .Z(n13354) );
  XOR U13561 ( .A(n13355), .B(n13354), .Z(n13373) );
  NAND U13562 ( .A(n19722), .B(n13264), .Z(n13266) );
  XNOR U13563 ( .A(b[5]), .B(n14062), .Z(n13364) );
  NANDN U13564 ( .A(n19640), .B(n13364), .Z(n13265) );
  NAND U13565 ( .A(n13266), .B(n13265), .Z(n13349) );
  XNOR U13566 ( .A(n19714), .B(n13906), .Z(n13367) );
  NANDN U13567 ( .A(n13367), .B(n19766), .Z(n13269) );
  NANDN U13568 ( .A(n13267), .B(n19767), .Z(n13268) );
  NAND U13569 ( .A(n13269), .B(n13268), .Z(n13346) );
  NAND U13570 ( .A(n19554), .B(n13270), .Z(n13272) );
  IV U13571 ( .A(a[175]), .Z(n14218) );
  XNOR U13572 ( .A(b[3]), .B(n14218), .Z(n13370) );
  NANDN U13573 ( .A(n19521), .B(n13370), .Z(n13271) );
  AND U13574 ( .A(n13272), .B(n13271), .Z(n13347) );
  XNOR U13575 ( .A(n13346), .B(n13347), .Z(n13348) );
  XOR U13576 ( .A(n13349), .B(n13348), .Z(n13374) );
  XOR U13577 ( .A(n13373), .B(n13374), .Z(n13375) );
  XNOR U13578 ( .A(n13376), .B(n13375), .Z(n13324) );
  NAND U13579 ( .A(n13274), .B(n13273), .Z(n13278) );
  NAND U13580 ( .A(n13276), .B(n13275), .Z(n13277) );
  NAND U13581 ( .A(n13278), .B(n13277), .Z(n13325) );
  XOR U13582 ( .A(n13324), .B(n13325), .Z(n13327) );
  XNOR U13583 ( .A(n20052), .B(n13567), .Z(n13330) );
  OR U13584 ( .A(n13330), .B(n20020), .Z(n13281) );
  NANDN U13585 ( .A(n13279), .B(n19960), .Z(n13280) );
  NAND U13586 ( .A(n13281), .B(n13280), .Z(n13343) );
  XNOR U13587 ( .A(n102), .B(n13282), .Z(n13334) );
  OR U13588 ( .A(n13334), .B(n20121), .Z(n13285) );
  NANDN U13589 ( .A(n13283), .B(n20122), .Z(n13284) );
  NAND U13590 ( .A(n13285), .B(n13284), .Z(n13340) );
  XNOR U13591 ( .A(n19975), .B(n13750), .Z(n13337) );
  NANDN U13592 ( .A(n13337), .B(n19883), .Z(n13288) );
  NANDN U13593 ( .A(n13286), .B(n19937), .Z(n13287) );
  AND U13594 ( .A(n13288), .B(n13287), .Z(n13341) );
  XNOR U13595 ( .A(n13340), .B(n13341), .Z(n13342) );
  XNOR U13596 ( .A(n13343), .B(n13342), .Z(n13379) );
  NANDN U13597 ( .A(n13290), .B(n13289), .Z(n13294) );
  NAND U13598 ( .A(n13292), .B(n13291), .Z(n13293) );
  NAND U13599 ( .A(n13294), .B(n13293), .Z(n13380) );
  XNOR U13600 ( .A(n13379), .B(n13380), .Z(n13381) );
  NANDN U13601 ( .A(n13296), .B(n13295), .Z(n13300) );
  NAND U13602 ( .A(n13298), .B(n13297), .Z(n13299) );
  AND U13603 ( .A(n13300), .B(n13299), .Z(n13382) );
  XNOR U13604 ( .A(n13381), .B(n13382), .Z(n13326) );
  XNOR U13605 ( .A(n13327), .B(n13326), .Z(n13385) );
  NANDN U13606 ( .A(n13302), .B(n13301), .Z(n13306) );
  NAND U13607 ( .A(n13304), .B(n13303), .Z(n13305) );
  NAND U13608 ( .A(n13306), .B(n13305), .Z(n13386) );
  XNOR U13609 ( .A(n13385), .B(n13386), .Z(n13387) );
  XOR U13610 ( .A(n13388), .B(n13387), .Z(n13318) );
  NANDN U13611 ( .A(n13308), .B(n13307), .Z(n13312) );
  NANDN U13612 ( .A(n13310), .B(n13309), .Z(n13311) );
  NAND U13613 ( .A(n13312), .B(n13311), .Z(n13319) );
  XNOR U13614 ( .A(n13318), .B(n13319), .Z(n13320) );
  XNOR U13615 ( .A(n13321), .B(n13320), .Z(n13391) );
  XNOR U13616 ( .A(n13391), .B(sreg[417]), .Z(n13393) );
  NAND U13617 ( .A(n13313), .B(sreg[416]), .Z(n13317) );
  OR U13618 ( .A(n13315), .B(n13314), .Z(n13316) );
  AND U13619 ( .A(n13317), .B(n13316), .Z(n13392) );
  XOR U13620 ( .A(n13393), .B(n13392), .Z(c[417]) );
  NANDN U13621 ( .A(n13319), .B(n13318), .Z(n13323) );
  NAND U13622 ( .A(n13321), .B(n13320), .Z(n13322) );
  NAND U13623 ( .A(n13323), .B(n13322), .Z(n13399) );
  NANDN U13624 ( .A(n13325), .B(n13324), .Z(n13329) );
  OR U13625 ( .A(n13327), .B(n13326), .Z(n13328) );
  NAND U13626 ( .A(n13329), .B(n13328), .Z(n13466) );
  XNOR U13627 ( .A(n20052), .B(n13672), .Z(n13435) );
  OR U13628 ( .A(n13435), .B(n20020), .Z(n13332) );
  NANDN U13629 ( .A(n13330), .B(n19960), .Z(n13331) );
  NAND U13630 ( .A(n13332), .B(n13331), .Z(n13448) );
  XNOR U13631 ( .A(n102), .B(n13333), .Z(n13439) );
  OR U13632 ( .A(n13439), .B(n20121), .Z(n13336) );
  NANDN U13633 ( .A(n13334), .B(n20122), .Z(n13335) );
  NAND U13634 ( .A(n13336), .B(n13335), .Z(n13445) );
  XNOR U13635 ( .A(n19975), .B(n13801), .Z(n13442) );
  NANDN U13636 ( .A(n13442), .B(n19883), .Z(n13339) );
  NANDN U13637 ( .A(n13337), .B(n19937), .Z(n13338) );
  AND U13638 ( .A(n13339), .B(n13338), .Z(n13446) );
  XNOR U13639 ( .A(n13445), .B(n13446), .Z(n13447) );
  XNOR U13640 ( .A(n13448), .B(n13447), .Z(n13457) );
  NANDN U13641 ( .A(n13341), .B(n13340), .Z(n13345) );
  NAND U13642 ( .A(n13343), .B(n13342), .Z(n13344) );
  NAND U13643 ( .A(n13345), .B(n13344), .Z(n13458) );
  XNOR U13644 ( .A(n13457), .B(n13458), .Z(n13459) );
  NANDN U13645 ( .A(n13347), .B(n13346), .Z(n13351) );
  NAND U13646 ( .A(n13349), .B(n13348), .Z(n13350) );
  AND U13647 ( .A(n13351), .B(n13350), .Z(n13460) );
  XNOR U13648 ( .A(n13459), .B(n13460), .Z(n13404) );
  NANDN U13649 ( .A(n13353), .B(n13352), .Z(n13357) );
  OR U13650 ( .A(n13355), .B(n13354), .Z(n13356) );
  NAND U13651 ( .A(n13357), .B(n13356), .Z(n13432) );
  NAND U13652 ( .A(b[0]), .B(a[178]), .Z(n13358) );
  XNOR U13653 ( .A(b[1]), .B(n13358), .Z(n13360) );
  NAND U13654 ( .A(a[177]), .B(n98), .Z(n13359) );
  AND U13655 ( .A(n13360), .B(n13359), .Z(n13408) );
  XNOR U13656 ( .A(n20154), .B(n13516), .Z(n13417) );
  OR U13657 ( .A(n13417), .B(n20057), .Z(n13363) );
  NANDN U13658 ( .A(n13361), .B(n20098), .Z(n13362) );
  AND U13659 ( .A(n13363), .B(n13362), .Z(n13409) );
  XOR U13660 ( .A(n13408), .B(n13409), .Z(n13411) );
  NAND U13661 ( .A(a[162]), .B(b[15]), .Z(n13410) );
  XOR U13662 ( .A(n13411), .B(n13410), .Z(n13429) );
  NAND U13663 ( .A(n19722), .B(n13364), .Z(n13366) );
  XNOR U13664 ( .A(b[5]), .B(n14113), .Z(n13420) );
  NANDN U13665 ( .A(n19640), .B(n13420), .Z(n13365) );
  NAND U13666 ( .A(n13366), .B(n13365), .Z(n13454) );
  XNOR U13667 ( .A(n19714), .B(n13984), .Z(n13423) );
  NANDN U13668 ( .A(n13423), .B(n19766), .Z(n13369) );
  NANDN U13669 ( .A(n13367), .B(n19767), .Z(n13368) );
  NAND U13670 ( .A(n13369), .B(n13368), .Z(n13451) );
  NAND U13671 ( .A(n19554), .B(n13370), .Z(n13372) );
  IV U13672 ( .A(a[176]), .Z(n14269) );
  XNOR U13673 ( .A(b[3]), .B(n14269), .Z(n13426) );
  NANDN U13674 ( .A(n19521), .B(n13426), .Z(n13371) );
  AND U13675 ( .A(n13372), .B(n13371), .Z(n13452) );
  XNOR U13676 ( .A(n13451), .B(n13452), .Z(n13453) );
  XOR U13677 ( .A(n13454), .B(n13453), .Z(n13430) );
  XOR U13678 ( .A(n13429), .B(n13430), .Z(n13431) );
  XNOR U13679 ( .A(n13432), .B(n13431), .Z(n13402) );
  NAND U13680 ( .A(n13374), .B(n13373), .Z(n13378) );
  NAND U13681 ( .A(n13376), .B(n13375), .Z(n13377) );
  NAND U13682 ( .A(n13378), .B(n13377), .Z(n13403) );
  XOR U13683 ( .A(n13402), .B(n13403), .Z(n13405) );
  XNOR U13684 ( .A(n13404), .B(n13405), .Z(n13463) );
  NANDN U13685 ( .A(n13380), .B(n13379), .Z(n13384) );
  NAND U13686 ( .A(n13382), .B(n13381), .Z(n13383) );
  NAND U13687 ( .A(n13384), .B(n13383), .Z(n13464) );
  XNOR U13688 ( .A(n13463), .B(n13464), .Z(n13465) );
  XOR U13689 ( .A(n13466), .B(n13465), .Z(n13396) );
  NANDN U13690 ( .A(n13386), .B(n13385), .Z(n13390) );
  NANDN U13691 ( .A(n13388), .B(n13387), .Z(n13389) );
  NAND U13692 ( .A(n13390), .B(n13389), .Z(n13397) );
  XNOR U13693 ( .A(n13396), .B(n13397), .Z(n13398) );
  XNOR U13694 ( .A(n13399), .B(n13398), .Z(n13469) );
  XNOR U13695 ( .A(n13469), .B(sreg[418]), .Z(n13471) );
  NAND U13696 ( .A(n13391), .B(sreg[417]), .Z(n13395) );
  OR U13697 ( .A(n13393), .B(n13392), .Z(n13394) );
  AND U13698 ( .A(n13395), .B(n13394), .Z(n13470) );
  XOR U13699 ( .A(n13471), .B(n13470), .Z(c[418]) );
  NANDN U13700 ( .A(n13397), .B(n13396), .Z(n13401) );
  NAND U13701 ( .A(n13399), .B(n13398), .Z(n13400) );
  NAND U13702 ( .A(n13401), .B(n13400), .Z(n13477) );
  NANDN U13703 ( .A(n13403), .B(n13402), .Z(n13407) );
  OR U13704 ( .A(n13405), .B(n13404), .Z(n13406) );
  NAND U13705 ( .A(n13407), .B(n13406), .Z(n13544) );
  NANDN U13706 ( .A(n13409), .B(n13408), .Z(n13413) );
  OR U13707 ( .A(n13411), .B(n13410), .Z(n13412) );
  NAND U13708 ( .A(n13413), .B(n13412), .Z(n13510) );
  NAND U13709 ( .A(b[0]), .B(a[179]), .Z(n13414) );
  XNOR U13710 ( .A(b[1]), .B(n13414), .Z(n13416) );
  NAND U13711 ( .A(a[178]), .B(n98), .Z(n13415) );
  AND U13712 ( .A(n13416), .B(n13415), .Z(n13486) );
  XNOR U13713 ( .A(n20154), .B(n13567), .Z(n13492) );
  OR U13714 ( .A(n13492), .B(n20057), .Z(n13419) );
  NANDN U13715 ( .A(n13417), .B(n20098), .Z(n13418) );
  AND U13716 ( .A(n13419), .B(n13418), .Z(n13487) );
  XOR U13717 ( .A(n13486), .B(n13487), .Z(n13489) );
  NAND U13718 ( .A(a[163]), .B(b[15]), .Z(n13488) );
  XOR U13719 ( .A(n13489), .B(n13488), .Z(n13507) );
  NAND U13720 ( .A(n19722), .B(n13420), .Z(n13422) );
  XNOR U13721 ( .A(b[5]), .B(n14218), .Z(n13498) );
  NANDN U13722 ( .A(n19640), .B(n13498), .Z(n13421) );
  NAND U13723 ( .A(n13422), .B(n13421), .Z(n13532) );
  XNOR U13724 ( .A(n19714), .B(n14062), .Z(n13501) );
  NANDN U13725 ( .A(n13501), .B(n19766), .Z(n13425) );
  NANDN U13726 ( .A(n13423), .B(n19767), .Z(n13424) );
  NAND U13727 ( .A(n13425), .B(n13424), .Z(n13529) );
  NAND U13728 ( .A(n19554), .B(n13426), .Z(n13428) );
  IV U13729 ( .A(a[177]), .Z(n14347) );
  XNOR U13730 ( .A(b[3]), .B(n14347), .Z(n13504) );
  NANDN U13731 ( .A(n19521), .B(n13504), .Z(n13427) );
  AND U13732 ( .A(n13428), .B(n13427), .Z(n13530) );
  XNOR U13733 ( .A(n13529), .B(n13530), .Z(n13531) );
  XOR U13734 ( .A(n13532), .B(n13531), .Z(n13508) );
  XOR U13735 ( .A(n13507), .B(n13508), .Z(n13509) );
  XNOR U13736 ( .A(n13510), .B(n13509), .Z(n13480) );
  NAND U13737 ( .A(n13430), .B(n13429), .Z(n13434) );
  NAND U13738 ( .A(n13432), .B(n13431), .Z(n13433) );
  NAND U13739 ( .A(n13434), .B(n13433), .Z(n13481) );
  XOR U13740 ( .A(n13480), .B(n13481), .Z(n13483) );
  XNOR U13741 ( .A(n20052), .B(n13750), .Z(n13513) );
  OR U13742 ( .A(n13513), .B(n20020), .Z(n13437) );
  NANDN U13743 ( .A(n13435), .B(n19960), .Z(n13436) );
  NAND U13744 ( .A(n13437), .B(n13436), .Z(n13526) );
  XNOR U13745 ( .A(n102), .B(n13438), .Z(n13517) );
  OR U13746 ( .A(n13517), .B(n20121), .Z(n13441) );
  NANDN U13747 ( .A(n13439), .B(n20122), .Z(n13440) );
  NAND U13748 ( .A(n13441), .B(n13440), .Z(n13523) );
  XNOR U13749 ( .A(n19975), .B(n13906), .Z(n13520) );
  NANDN U13750 ( .A(n13520), .B(n19883), .Z(n13444) );
  NANDN U13751 ( .A(n13442), .B(n19937), .Z(n13443) );
  AND U13752 ( .A(n13444), .B(n13443), .Z(n13524) );
  XNOR U13753 ( .A(n13523), .B(n13524), .Z(n13525) );
  XNOR U13754 ( .A(n13526), .B(n13525), .Z(n13535) );
  NANDN U13755 ( .A(n13446), .B(n13445), .Z(n13450) );
  NAND U13756 ( .A(n13448), .B(n13447), .Z(n13449) );
  NAND U13757 ( .A(n13450), .B(n13449), .Z(n13536) );
  XNOR U13758 ( .A(n13535), .B(n13536), .Z(n13537) );
  NANDN U13759 ( .A(n13452), .B(n13451), .Z(n13456) );
  NAND U13760 ( .A(n13454), .B(n13453), .Z(n13455) );
  AND U13761 ( .A(n13456), .B(n13455), .Z(n13538) );
  XNOR U13762 ( .A(n13537), .B(n13538), .Z(n13482) );
  XNOR U13763 ( .A(n13483), .B(n13482), .Z(n13541) );
  NANDN U13764 ( .A(n13458), .B(n13457), .Z(n13462) );
  NAND U13765 ( .A(n13460), .B(n13459), .Z(n13461) );
  NAND U13766 ( .A(n13462), .B(n13461), .Z(n13542) );
  XNOR U13767 ( .A(n13541), .B(n13542), .Z(n13543) );
  XOR U13768 ( .A(n13544), .B(n13543), .Z(n13474) );
  NANDN U13769 ( .A(n13464), .B(n13463), .Z(n13468) );
  NANDN U13770 ( .A(n13466), .B(n13465), .Z(n13467) );
  NAND U13771 ( .A(n13468), .B(n13467), .Z(n13475) );
  XNOR U13772 ( .A(n13474), .B(n13475), .Z(n13476) );
  XNOR U13773 ( .A(n13477), .B(n13476), .Z(n13547) );
  XNOR U13774 ( .A(n13547), .B(sreg[419]), .Z(n13549) );
  NAND U13775 ( .A(n13469), .B(sreg[418]), .Z(n13473) );
  OR U13776 ( .A(n13471), .B(n13470), .Z(n13472) );
  AND U13777 ( .A(n13473), .B(n13472), .Z(n13548) );
  XOR U13778 ( .A(n13549), .B(n13548), .Z(c[419]) );
  NANDN U13779 ( .A(n13475), .B(n13474), .Z(n13479) );
  NAND U13780 ( .A(n13477), .B(n13476), .Z(n13478) );
  NAND U13781 ( .A(n13479), .B(n13478), .Z(n13555) );
  NANDN U13782 ( .A(n13481), .B(n13480), .Z(n13485) );
  OR U13783 ( .A(n13483), .B(n13482), .Z(n13484) );
  NAND U13784 ( .A(n13485), .B(n13484), .Z(n13622) );
  NANDN U13785 ( .A(n13487), .B(n13486), .Z(n13491) );
  OR U13786 ( .A(n13489), .B(n13488), .Z(n13490) );
  NAND U13787 ( .A(n13491), .B(n13490), .Z(n13610) );
  XNOR U13788 ( .A(n20154), .B(n13672), .Z(n13595) );
  OR U13789 ( .A(n13595), .B(n20057), .Z(n13494) );
  NANDN U13790 ( .A(n13492), .B(n20098), .Z(n13493) );
  AND U13791 ( .A(n13494), .B(n13493), .Z(n13587) );
  NAND U13792 ( .A(b[0]), .B(a[180]), .Z(n13495) );
  XNOR U13793 ( .A(b[1]), .B(n13495), .Z(n13497) );
  NAND U13794 ( .A(a[179]), .B(n98), .Z(n13496) );
  AND U13795 ( .A(n13497), .B(n13496), .Z(n13586) );
  XOR U13796 ( .A(n13587), .B(n13586), .Z(n13589) );
  NAND U13797 ( .A(a[164]), .B(b[15]), .Z(n13588) );
  XOR U13798 ( .A(n13589), .B(n13588), .Z(n13607) );
  NAND U13799 ( .A(n19722), .B(n13498), .Z(n13500) );
  XNOR U13800 ( .A(b[5]), .B(n14269), .Z(n13598) );
  NANDN U13801 ( .A(n19640), .B(n13598), .Z(n13499) );
  NAND U13802 ( .A(n13500), .B(n13499), .Z(n13583) );
  XNOR U13803 ( .A(n19714), .B(n14113), .Z(n13601) );
  NANDN U13804 ( .A(n13601), .B(n19766), .Z(n13503) );
  NANDN U13805 ( .A(n13501), .B(n19767), .Z(n13502) );
  NAND U13806 ( .A(n13503), .B(n13502), .Z(n13580) );
  NAND U13807 ( .A(n19554), .B(n13504), .Z(n13506) );
  IV U13808 ( .A(a[178]), .Z(n14425) );
  XNOR U13809 ( .A(b[3]), .B(n14425), .Z(n13604) );
  NANDN U13810 ( .A(n19521), .B(n13604), .Z(n13505) );
  AND U13811 ( .A(n13506), .B(n13505), .Z(n13581) );
  XNOR U13812 ( .A(n13580), .B(n13581), .Z(n13582) );
  XOR U13813 ( .A(n13583), .B(n13582), .Z(n13608) );
  XOR U13814 ( .A(n13607), .B(n13608), .Z(n13609) );
  XNOR U13815 ( .A(n13610), .B(n13609), .Z(n13558) );
  NAND U13816 ( .A(n13508), .B(n13507), .Z(n13512) );
  NAND U13817 ( .A(n13510), .B(n13509), .Z(n13511) );
  NAND U13818 ( .A(n13512), .B(n13511), .Z(n13559) );
  XOR U13819 ( .A(n13558), .B(n13559), .Z(n13561) );
  XNOR U13820 ( .A(n20052), .B(n13801), .Z(n13564) );
  OR U13821 ( .A(n13564), .B(n20020), .Z(n13515) );
  NANDN U13822 ( .A(n13513), .B(n19960), .Z(n13514) );
  NAND U13823 ( .A(n13515), .B(n13514), .Z(n13577) );
  XNOR U13824 ( .A(n102), .B(n13516), .Z(n13568) );
  OR U13825 ( .A(n13568), .B(n20121), .Z(n13519) );
  NANDN U13826 ( .A(n13517), .B(n20122), .Z(n13518) );
  NAND U13827 ( .A(n13519), .B(n13518), .Z(n13574) );
  XNOR U13828 ( .A(n19975), .B(n13984), .Z(n13571) );
  NANDN U13829 ( .A(n13571), .B(n19883), .Z(n13522) );
  NANDN U13830 ( .A(n13520), .B(n19937), .Z(n13521) );
  AND U13831 ( .A(n13522), .B(n13521), .Z(n13575) );
  XNOR U13832 ( .A(n13574), .B(n13575), .Z(n13576) );
  XNOR U13833 ( .A(n13577), .B(n13576), .Z(n13613) );
  NANDN U13834 ( .A(n13524), .B(n13523), .Z(n13528) );
  NAND U13835 ( .A(n13526), .B(n13525), .Z(n13527) );
  NAND U13836 ( .A(n13528), .B(n13527), .Z(n13614) );
  XNOR U13837 ( .A(n13613), .B(n13614), .Z(n13615) );
  NANDN U13838 ( .A(n13530), .B(n13529), .Z(n13534) );
  NAND U13839 ( .A(n13532), .B(n13531), .Z(n13533) );
  AND U13840 ( .A(n13534), .B(n13533), .Z(n13616) );
  XNOR U13841 ( .A(n13615), .B(n13616), .Z(n13560) );
  XNOR U13842 ( .A(n13561), .B(n13560), .Z(n13619) );
  NANDN U13843 ( .A(n13536), .B(n13535), .Z(n13540) );
  NAND U13844 ( .A(n13538), .B(n13537), .Z(n13539) );
  NAND U13845 ( .A(n13540), .B(n13539), .Z(n13620) );
  XNOR U13846 ( .A(n13619), .B(n13620), .Z(n13621) );
  XOR U13847 ( .A(n13622), .B(n13621), .Z(n13552) );
  NANDN U13848 ( .A(n13542), .B(n13541), .Z(n13546) );
  NANDN U13849 ( .A(n13544), .B(n13543), .Z(n13545) );
  NAND U13850 ( .A(n13546), .B(n13545), .Z(n13553) );
  XNOR U13851 ( .A(n13552), .B(n13553), .Z(n13554) );
  XNOR U13852 ( .A(n13555), .B(n13554), .Z(n13625) );
  XNOR U13853 ( .A(n13625), .B(sreg[420]), .Z(n13627) );
  NAND U13854 ( .A(n13547), .B(sreg[419]), .Z(n13551) );
  OR U13855 ( .A(n13549), .B(n13548), .Z(n13550) );
  AND U13856 ( .A(n13551), .B(n13550), .Z(n13626) );
  XOR U13857 ( .A(n13627), .B(n13626), .Z(c[420]) );
  NANDN U13858 ( .A(n13553), .B(n13552), .Z(n13557) );
  NAND U13859 ( .A(n13555), .B(n13554), .Z(n13556) );
  NAND U13860 ( .A(n13557), .B(n13556), .Z(n13633) );
  NANDN U13861 ( .A(n13559), .B(n13558), .Z(n13563) );
  OR U13862 ( .A(n13561), .B(n13560), .Z(n13562) );
  NAND U13863 ( .A(n13563), .B(n13562), .Z(n13700) );
  XNOR U13864 ( .A(n20052), .B(n13906), .Z(n13669) );
  OR U13865 ( .A(n13669), .B(n20020), .Z(n13566) );
  NANDN U13866 ( .A(n13564), .B(n19960), .Z(n13565) );
  NAND U13867 ( .A(n13566), .B(n13565), .Z(n13682) );
  XNOR U13868 ( .A(n102), .B(n13567), .Z(n13673) );
  OR U13869 ( .A(n13673), .B(n20121), .Z(n13570) );
  NANDN U13870 ( .A(n13568), .B(n20122), .Z(n13569) );
  NAND U13871 ( .A(n13570), .B(n13569), .Z(n13679) );
  XNOR U13872 ( .A(n19975), .B(n14062), .Z(n13676) );
  NANDN U13873 ( .A(n13676), .B(n19883), .Z(n13573) );
  NANDN U13874 ( .A(n13571), .B(n19937), .Z(n13572) );
  AND U13875 ( .A(n13573), .B(n13572), .Z(n13680) );
  XNOR U13876 ( .A(n13679), .B(n13680), .Z(n13681) );
  XNOR U13877 ( .A(n13682), .B(n13681), .Z(n13691) );
  NANDN U13878 ( .A(n13575), .B(n13574), .Z(n13579) );
  NAND U13879 ( .A(n13577), .B(n13576), .Z(n13578) );
  NAND U13880 ( .A(n13579), .B(n13578), .Z(n13692) );
  XNOR U13881 ( .A(n13691), .B(n13692), .Z(n13693) );
  NANDN U13882 ( .A(n13581), .B(n13580), .Z(n13585) );
  NAND U13883 ( .A(n13583), .B(n13582), .Z(n13584) );
  AND U13884 ( .A(n13585), .B(n13584), .Z(n13694) );
  XNOR U13885 ( .A(n13693), .B(n13694), .Z(n13638) );
  NANDN U13886 ( .A(n13587), .B(n13586), .Z(n13591) );
  OR U13887 ( .A(n13589), .B(n13588), .Z(n13590) );
  NAND U13888 ( .A(n13591), .B(n13590), .Z(n13666) );
  NAND U13889 ( .A(b[0]), .B(a[181]), .Z(n13592) );
  XNOR U13890 ( .A(b[1]), .B(n13592), .Z(n13594) );
  NAND U13891 ( .A(a[180]), .B(n98), .Z(n13593) );
  AND U13892 ( .A(n13594), .B(n13593), .Z(n13642) );
  XNOR U13893 ( .A(n20154), .B(n13750), .Z(n13648) );
  OR U13894 ( .A(n13648), .B(n20057), .Z(n13597) );
  NANDN U13895 ( .A(n13595), .B(n20098), .Z(n13596) );
  AND U13896 ( .A(n13597), .B(n13596), .Z(n13643) );
  XOR U13897 ( .A(n13642), .B(n13643), .Z(n13645) );
  NAND U13898 ( .A(a[165]), .B(b[15]), .Z(n13644) );
  XOR U13899 ( .A(n13645), .B(n13644), .Z(n13663) );
  NAND U13900 ( .A(n19722), .B(n13598), .Z(n13600) );
  XNOR U13901 ( .A(b[5]), .B(n14347), .Z(n13654) );
  NANDN U13902 ( .A(n19640), .B(n13654), .Z(n13599) );
  NAND U13903 ( .A(n13600), .B(n13599), .Z(n13688) );
  XNOR U13904 ( .A(n19714), .B(n14218), .Z(n13657) );
  NANDN U13905 ( .A(n13657), .B(n19766), .Z(n13603) );
  NANDN U13906 ( .A(n13601), .B(n19767), .Z(n13602) );
  NAND U13907 ( .A(n13603), .B(n13602), .Z(n13685) );
  NAND U13908 ( .A(n19554), .B(n13604), .Z(n13606) );
  IV U13909 ( .A(a[179]), .Z(n14503) );
  XNOR U13910 ( .A(b[3]), .B(n14503), .Z(n13660) );
  NANDN U13911 ( .A(n19521), .B(n13660), .Z(n13605) );
  AND U13912 ( .A(n13606), .B(n13605), .Z(n13686) );
  XNOR U13913 ( .A(n13685), .B(n13686), .Z(n13687) );
  XOR U13914 ( .A(n13688), .B(n13687), .Z(n13664) );
  XOR U13915 ( .A(n13663), .B(n13664), .Z(n13665) );
  XNOR U13916 ( .A(n13666), .B(n13665), .Z(n13636) );
  NAND U13917 ( .A(n13608), .B(n13607), .Z(n13612) );
  NAND U13918 ( .A(n13610), .B(n13609), .Z(n13611) );
  NAND U13919 ( .A(n13612), .B(n13611), .Z(n13637) );
  XOR U13920 ( .A(n13636), .B(n13637), .Z(n13639) );
  XNOR U13921 ( .A(n13638), .B(n13639), .Z(n13697) );
  NANDN U13922 ( .A(n13614), .B(n13613), .Z(n13618) );
  NAND U13923 ( .A(n13616), .B(n13615), .Z(n13617) );
  NAND U13924 ( .A(n13618), .B(n13617), .Z(n13698) );
  XNOR U13925 ( .A(n13697), .B(n13698), .Z(n13699) );
  XOR U13926 ( .A(n13700), .B(n13699), .Z(n13630) );
  NANDN U13927 ( .A(n13620), .B(n13619), .Z(n13624) );
  NANDN U13928 ( .A(n13622), .B(n13621), .Z(n13623) );
  NAND U13929 ( .A(n13624), .B(n13623), .Z(n13631) );
  XNOR U13930 ( .A(n13630), .B(n13631), .Z(n13632) );
  XNOR U13931 ( .A(n13633), .B(n13632), .Z(n13703) );
  XNOR U13932 ( .A(n13703), .B(sreg[421]), .Z(n13705) );
  NAND U13933 ( .A(n13625), .B(sreg[420]), .Z(n13629) );
  OR U13934 ( .A(n13627), .B(n13626), .Z(n13628) );
  AND U13935 ( .A(n13629), .B(n13628), .Z(n13704) );
  XOR U13936 ( .A(n13705), .B(n13704), .Z(c[421]) );
  NANDN U13937 ( .A(n13631), .B(n13630), .Z(n13635) );
  NAND U13938 ( .A(n13633), .B(n13632), .Z(n13634) );
  NAND U13939 ( .A(n13635), .B(n13634), .Z(n13711) );
  NANDN U13940 ( .A(n13637), .B(n13636), .Z(n13641) );
  OR U13941 ( .A(n13639), .B(n13638), .Z(n13640) );
  NAND U13942 ( .A(n13641), .B(n13640), .Z(n13778) );
  NANDN U13943 ( .A(n13643), .B(n13642), .Z(n13647) );
  OR U13944 ( .A(n13645), .B(n13644), .Z(n13646) );
  NAND U13945 ( .A(n13647), .B(n13646), .Z(n13744) );
  XNOR U13946 ( .A(n20154), .B(n13801), .Z(n13729) );
  OR U13947 ( .A(n13729), .B(n20057), .Z(n13650) );
  NANDN U13948 ( .A(n13648), .B(n20098), .Z(n13649) );
  AND U13949 ( .A(n13650), .B(n13649), .Z(n13721) );
  NAND U13950 ( .A(b[0]), .B(a[182]), .Z(n13651) );
  XNOR U13951 ( .A(b[1]), .B(n13651), .Z(n13653) );
  NAND U13952 ( .A(a[181]), .B(n98), .Z(n13652) );
  AND U13953 ( .A(n13653), .B(n13652), .Z(n13720) );
  XOR U13954 ( .A(n13721), .B(n13720), .Z(n13723) );
  NAND U13955 ( .A(a[166]), .B(b[15]), .Z(n13722) );
  XOR U13956 ( .A(n13723), .B(n13722), .Z(n13741) );
  NAND U13957 ( .A(n19722), .B(n13654), .Z(n13656) );
  XNOR U13958 ( .A(b[5]), .B(n14425), .Z(n13732) );
  NANDN U13959 ( .A(n19640), .B(n13732), .Z(n13655) );
  NAND U13960 ( .A(n13656), .B(n13655), .Z(n13766) );
  XNOR U13961 ( .A(n19714), .B(n14269), .Z(n13735) );
  NANDN U13962 ( .A(n13735), .B(n19766), .Z(n13659) );
  NANDN U13963 ( .A(n13657), .B(n19767), .Z(n13658) );
  NAND U13964 ( .A(n13659), .B(n13658), .Z(n13763) );
  NAND U13965 ( .A(n19554), .B(n13660), .Z(n13662) );
  IV U13966 ( .A(a[180]), .Z(n14581) );
  XNOR U13967 ( .A(b[3]), .B(n14581), .Z(n13738) );
  NANDN U13968 ( .A(n19521), .B(n13738), .Z(n13661) );
  AND U13969 ( .A(n13662), .B(n13661), .Z(n13764) );
  XNOR U13970 ( .A(n13763), .B(n13764), .Z(n13765) );
  XOR U13971 ( .A(n13766), .B(n13765), .Z(n13742) );
  XOR U13972 ( .A(n13741), .B(n13742), .Z(n13743) );
  XNOR U13973 ( .A(n13744), .B(n13743), .Z(n13714) );
  NAND U13974 ( .A(n13664), .B(n13663), .Z(n13668) );
  NAND U13975 ( .A(n13666), .B(n13665), .Z(n13667) );
  NAND U13976 ( .A(n13668), .B(n13667), .Z(n13715) );
  XOR U13977 ( .A(n13714), .B(n13715), .Z(n13717) );
  XNOR U13978 ( .A(n20052), .B(n13984), .Z(n13747) );
  OR U13979 ( .A(n13747), .B(n20020), .Z(n13671) );
  NANDN U13980 ( .A(n13669), .B(n19960), .Z(n13670) );
  NAND U13981 ( .A(n13671), .B(n13670), .Z(n13760) );
  XNOR U13982 ( .A(n102), .B(n13672), .Z(n13751) );
  OR U13983 ( .A(n13751), .B(n20121), .Z(n13675) );
  NANDN U13984 ( .A(n13673), .B(n20122), .Z(n13674) );
  NAND U13985 ( .A(n13675), .B(n13674), .Z(n13757) );
  XNOR U13986 ( .A(n19975), .B(n14113), .Z(n13754) );
  NANDN U13987 ( .A(n13754), .B(n19883), .Z(n13678) );
  NANDN U13988 ( .A(n13676), .B(n19937), .Z(n13677) );
  AND U13989 ( .A(n13678), .B(n13677), .Z(n13758) );
  XNOR U13990 ( .A(n13757), .B(n13758), .Z(n13759) );
  XNOR U13991 ( .A(n13760), .B(n13759), .Z(n13769) );
  NANDN U13992 ( .A(n13680), .B(n13679), .Z(n13684) );
  NAND U13993 ( .A(n13682), .B(n13681), .Z(n13683) );
  NAND U13994 ( .A(n13684), .B(n13683), .Z(n13770) );
  XNOR U13995 ( .A(n13769), .B(n13770), .Z(n13771) );
  NANDN U13996 ( .A(n13686), .B(n13685), .Z(n13690) );
  NAND U13997 ( .A(n13688), .B(n13687), .Z(n13689) );
  AND U13998 ( .A(n13690), .B(n13689), .Z(n13772) );
  XNOR U13999 ( .A(n13771), .B(n13772), .Z(n13716) );
  XNOR U14000 ( .A(n13717), .B(n13716), .Z(n13775) );
  NANDN U14001 ( .A(n13692), .B(n13691), .Z(n13696) );
  NAND U14002 ( .A(n13694), .B(n13693), .Z(n13695) );
  NAND U14003 ( .A(n13696), .B(n13695), .Z(n13776) );
  XNOR U14004 ( .A(n13775), .B(n13776), .Z(n13777) );
  XOR U14005 ( .A(n13778), .B(n13777), .Z(n13708) );
  NANDN U14006 ( .A(n13698), .B(n13697), .Z(n13702) );
  NANDN U14007 ( .A(n13700), .B(n13699), .Z(n13701) );
  NAND U14008 ( .A(n13702), .B(n13701), .Z(n13709) );
  XNOR U14009 ( .A(n13708), .B(n13709), .Z(n13710) );
  XNOR U14010 ( .A(n13711), .B(n13710), .Z(n13781) );
  XNOR U14011 ( .A(n13781), .B(sreg[422]), .Z(n13783) );
  NAND U14012 ( .A(n13703), .B(sreg[421]), .Z(n13707) );
  OR U14013 ( .A(n13705), .B(n13704), .Z(n13706) );
  AND U14014 ( .A(n13707), .B(n13706), .Z(n13782) );
  XOR U14015 ( .A(n13783), .B(n13782), .Z(c[422]) );
  NANDN U14016 ( .A(n13709), .B(n13708), .Z(n13713) );
  NAND U14017 ( .A(n13711), .B(n13710), .Z(n13712) );
  NAND U14018 ( .A(n13713), .B(n13712), .Z(n13789) );
  NANDN U14019 ( .A(n13715), .B(n13714), .Z(n13719) );
  OR U14020 ( .A(n13717), .B(n13716), .Z(n13718) );
  NAND U14021 ( .A(n13719), .B(n13718), .Z(n13856) );
  NANDN U14022 ( .A(n13721), .B(n13720), .Z(n13725) );
  OR U14023 ( .A(n13723), .B(n13722), .Z(n13724) );
  NAND U14024 ( .A(n13725), .B(n13724), .Z(n13844) );
  NAND U14025 ( .A(b[0]), .B(a[183]), .Z(n13726) );
  XNOR U14026 ( .A(b[1]), .B(n13726), .Z(n13728) );
  NAND U14027 ( .A(a[182]), .B(n98), .Z(n13727) );
  AND U14028 ( .A(n13728), .B(n13727), .Z(n13820) );
  XNOR U14029 ( .A(n20154), .B(n13906), .Z(n13829) );
  OR U14030 ( .A(n13829), .B(n20057), .Z(n13731) );
  NANDN U14031 ( .A(n13729), .B(n20098), .Z(n13730) );
  AND U14032 ( .A(n13731), .B(n13730), .Z(n13821) );
  XOR U14033 ( .A(n13820), .B(n13821), .Z(n13823) );
  NAND U14034 ( .A(a[167]), .B(b[15]), .Z(n13822) );
  XOR U14035 ( .A(n13823), .B(n13822), .Z(n13841) );
  NAND U14036 ( .A(n19722), .B(n13732), .Z(n13734) );
  XNOR U14037 ( .A(b[5]), .B(n14503), .Z(n13832) );
  NANDN U14038 ( .A(n19640), .B(n13832), .Z(n13733) );
  NAND U14039 ( .A(n13734), .B(n13733), .Z(n13817) );
  XNOR U14040 ( .A(n19714), .B(n14347), .Z(n13835) );
  NANDN U14041 ( .A(n13835), .B(n19766), .Z(n13737) );
  NANDN U14042 ( .A(n13735), .B(n19767), .Z(n13736) );
  NAND U14043 ( .A(n13737), .B(n13736), .Z(n13814) );
  NAND U14044 ( .A(n19554), .B(n13738), .Z(n13740) );
  IV U14045 ( .A(a[181]), .Z(n14659) );
  XNOR U14046 ( .A(b[3]), .B(n14659), .Z(n13838) );
  NANDN U14047 ( .A(n19521), .B(n13838), .Z(n13739) );
  AND U14048 ( .A(n13740), .B(n13739), .Z(n13815) );
  XNOR U14049 ( .A(n13814), .B(n13815), .Z(n13816) );
  XOR U14050 ( .A(n13817), .B(n13816), .Z(n13842) );
  XOR U14051 ( .A(n13841), .B(n13842), .Z(n13843) );
  XNOR U14052 ( .A(n13844), .B(n13843), .Z(n13792) );
  NAND U14053 ( .A(n13742), .B(n13741), .Z(n13746) );
  NAND U14054 ( .A(n13744), .B(n13743), .Z(n13745) );
  NAND U14055 ( .A(n13746), .B(n13745), .Z(n13793) );
  XOR U14056 ( .A(n13792), .B(n13793), .Z(n13795) );
  XNOR U14057 ( .A(n20052), .B(n14062), .Z(n13798) );
  OR U14058 ( .A(n13798), .B(n20020), .Z(n13749) );
  NANDN U14059 ( .A(n13747), .B(n19960), .Z(n13748) );
  NAND U14060 ( .A(n13749), .B(n13748), .Z(n13811) );
  XNOR U14061 ( .A(n102), .B(n13750), .Z(n13802) );
  OR U14062 ( .A(n13802), .B(n20121), .Z(n13753) );
  NANDN U14063 ( .A(n13751), .B(n20122), .Z(n13752) );
  NAND U14064 ( .A(n13753), .B(n13752), .Z(n13808) );
  XNOR U14065 ( .A(n19975), .B(n14218), .Z(n13805) );
  NANDN U14066 ( .A(n13805), .B(n19883), .Z(n13756) );
  NANDN U14067 ( .A(n13754), .B(n19937), .Z(n13755) );
  AND U14068 ( .A(n13756), .B(n13755), .Z(n13809) );
  XNOR U14069 ( .A(n13808), .B(n13809), .Z(n13810) );
  XNOR U14070 ( .A(n13811), .B(n13810), .Z(n13847) );
  NANDN U14071 ( .A(n13758), .B(n13757), .Z(n13762) );
  NAND U14072 ( .A(n13760), .B(n13759), .Z(n13761) );
  NAND U14073 ( .A(n13762), .B(n13761), .Z(n13848) );
  XNOR U14074 ( .A(n13847), .B(n13848), .Z(n13849) );
  NANDN U14075 ( .A(n13764), .B(n13763), .Z(n13768) );
  NAND U14076 ( .A(n13766), .B(n13765), .Z(n13767) );
  AND U14077 ( .A(n13768), .B(n13767), .Z(n13850) );
  XNOR U14078 ( .A(n13849), .B(n13850), .Z(n13794) );
  XNOR U14079 ( .A(n13795), .B(n13794), .Z(n13853) );
  NANDN U14080 ( .A(n13770), .B(n13769), .Z(n13774) );
  NAND U14081 ( .A(n13772), .B(n13771), .Z(n13773) );
  NAND U14082 ( .A(n13774), .B(n13773), .Z(n13854) );
  XNOR U14083 ( .A(n13853), .B(n13854), .Z(n13855) );
  XOR U14084 ( .A(n13856), .B(n13855), .Z(n13786) );
  NANDN U14085 ( .A(n13776), .B(n13775), .Z(n13780) );
  NANDN U14086 ( .A(n13778), .B(n13777), .Z(n13779) );
  NAND U14087 ( .A(n13780), .B(n13779), .Z(n13787) );
  XNOR U14088 ( .A(n13786), .B(n13787), .Z(n13788) );
  XNOR U14089 ( .A(n13789), .B(n13788), .Z(n13859) );
  XNOR U14090 ( .A(n13859), .B(sreg[423]), .Z(n13861) );
  NAND U14091 ( .A(n13781), .B(sreg[422]), .Z(n13785) );
  OR U14092 ( .A(n13783), .B(n13782), .Z(n13784) );
  AND U14093 ( .A(n13785), .B(n13784), .Z(n13860) );
  XOR U14094 ( .A(n13861), .B(n13860), .Z(c[423]) );
  NANDN U14095 ( .A(n13787), .B(n13786), .Z(n13791) );
  NAND U14096 ( .A(n13789), .B(n13788), .Z(n13790) );
  NAND U14097 ( .A(n13791), .B(n13790), .Z(n13867) );
  NANDN U14098 ( .A(n13793), .B(n13792), .Z(n13797) );
  OR U14099 ( .A(n13795), .B(n13794), .Z(n13796) );
  NAND U14100 ( .A(n13797), .B(n13796), .Z(n13934) );
  XNOR U14101 ( .A(n20052), .B(n14113), .Z(n13903) );
  OR U14102 ( .A(n13903), .B(n20020), .Z(n13800) );
  NANDN U14103 ( .A(n13798), .B(n19960), .Z(n13799) );
  NAND U14104 ( .A(n13800), .B(n13799), .Z(n13916) );
  XNOR U14105 ( .A(n102), .B(n13801), .Z(n13907) );
  OR U14106 ( .A(n13907), .B(n20121), .Z(n13804) );
  NANDN U14107 ( .A(n13802), .B(n20122), .Z(n13803) );
  NAND U14108 ( .A(n13804), .B(n13803), .Z(n13913) );
  XNOR U14109 ( .A(n19975), .B(n14269), .Z(n13910) );
  NANDN U14110 ( .A(n13910), .B(n19883), .Z(n13807) );
  NANDN U14111 ( .A(n13805), .B(n19937), .Z(n13806) );
  AND U14112 ( .A(n13807), .B(n13806), .Z(n13914) );
  XNOR U14113 ( .A(n13913), .B(n13914), .Z(n13915) );
  XNOR U14114 ( .A(n13916), .B(n13915), .Z(n13925) );
  NANDN U14115 ( .A(n13809), .B(n13808), .Z(n13813) );
  NAND U14116 ( .A(n13811), .B(n13810), .Z(n13812) );
  NAND U14117 ( .A(n13813), .B(n13812), .Z(n13926) );
  XNOR U14118 ( .A(n13925), .B(n13926), .Z(n13927) );
  NANDN U14119 ( .A(n13815), .B(n13814), .Z(n13819) );
  NAND U14120 ( .A(n13817), .B(n13816), .Z(n13818) );
  AND U14121 ( .A(n13819), .B(n13818), .Z(n13928) );
  XNOR U14122 ( .A(n13927), .B(n13928), .Z(n13872) );
  NANDN U14123 ( .A(n13821), .B(n13820), .Z(n13825) );
  OR U14124 ( .A(n13823), .B(n13822), .Z(n13824) );
  NAND U14125 ( .A(n13825), .B(n13824), .Z(n13900) );
  NAND U14126 ( .A(b[0]), .B(a[184]), .Z(n13826) );
  XNOR U14127 ( .A(b[1]), .B(n13826), .Z(n13828) );
  NAND U14128 ( .A(a[183]), .B(n98), .Z(n13827) );
  AND U14129 ( .A(n13828), .B(n13827), .Z(n13876) );
  XNOR U14130 ( .A(n20154), .B(n13984), .Z(n13885) );
  OR U14131 ( .A(n13885), .B(n20057), .Z(n13831) );
  NANDN U14132 ( .A(n13829), .B(n20098), .Z(n13830) );
  AND U14133 ( .A(n13831), .B(n13830), .Z(n13877) );
  XOR U14134 ( .A(n13876), .B(n13877), .Z(n13879) );
  NAND U14135 ( .A(a[168]), .B(b[15]), .Z(n13878) );
  XOR U14136 ( .A(n13879), .B(n13878), .Z(n13897) );
  NAND U14137 ( .A(n19722), .B(n13832), .Z(n13834) );
  XNOR U14138 ( .A(b[5]), .B(n14581), .Z(n13888) );
  NANDN U14139 ( .A(n19640), .B(n13888), .Z(n13833) );
  NAND U14140 ( .A(n13834), .B(n13833), .Z(n13922) );
  XNOR U14141 ( .A(n19714), .B(n14425), .Z(n13891) );
  NANDN U14142 ( .A(n13891), .B(n19766), .Z(n13837) );
  NANDN U14143 ( .A(n13835), .B(n19767), .Z(n13836) );
  NAND U14144 ( .A(n13837), .B(n13836), .Z(n13919) );
  NAND U14145 ( .A(n19554), .B(n13838), .Z(n13840) );
  IV U14146 ( .A(a[182]), .Z(n14737) );
  XNOR U14147 ( .A(b[3]), .B(n14737), .Z(n13894) );
  NANDN U14148 ( .A(n19521), .B(n13894), .Z(n13839) );
  AND U14149 ( .A(n13840), .B(n13839), .Z(n13920) );
  XNOR U14150 ( .A(n13919), .B(n13920), .Z(n13921) );
  XOR U14151 ( .A(n13922), .B(n13921), .Z(n13898) );
  XOR U14152 ( .A(n13897), .B(n13898), .Z(n13899) );
  XNOR U14153 ( .A(n13900), .B(n13899), .Z(n13870) );
  NAND U14154 ( .A(n13842), .B(n13841), .Z(n13846) );
  NAND U14155 ( .A(n13844), .B(n13843), .Z(n13845) );
  NAND U14156 ( .A(n13846), .B(n13845), .Z(n13871) );
  XOR U14157 ( .A(n13870), .B(n13871), .Z(n13873) );
  XNOR U14158 ( .A(n13872), .B(n13873), .Z(n13931) );
  NANDN U14159 ( .A(n13848), .B(n13847), .Z(n13852) );
  NAND U14160 ( .A(n13850), .B(n13849), .Z(n13851) );
  NAND U14161 ( .A(n13852), .B(n13851), .Z(n13932) );
  XNOR U14162 ( .A(n13931), .B(n13932), .Z(n13933) );
  XOR U14163 ( .A(n13934), .B(n13933), .Z(n13864) );
  NANDN U14164 ( .A(n13854), .B(n13853), .Z(n13858) );
  NANDN U14165 ( .A(n13856), .B(n13855), .Z(n13857) );
  NAND U14166 ( .A(n13858), .B(n13857), .Z(n13865) );
  XNOR U14167 ( .A(n13864), .B(n13865), .Z(n13866) );
  XNOR U14168 ( .A(n13867), .B(n13866), .Z(n13937) );
  XNOR U14169 ( .A(n13937), .B(sreg[424]), .Z(n13939) );
  NAND U14170 ( .A(n13859), .B(sreg[423]), .Z(n13863) );
  OR U14171 ( .A(n13861), .B(n13860), .Z(n13862) );
  AND U14172 ( .A(n13863), .B(n13862), .Z(n13938) );
  XOR U14173 ( .A(n13939), .B(n13938), .Z(c[424]) );
  NANDN U14174 ( .A(n13865), .B(n13864), .Z(n13869) );
  NAND U14175 ( .A(n13867), .B(n13866), .Z(n13868) );
  NAND U14176 ( .A(n13869), .B(n13868), .Z(n13945) );
  NANDN U14177 ( .A(n13871), .B(n13870), .Z(n13875) );
  OR U14178 ( .A(n13873), .B(n13872), .Z(n13874) );
  NAND U14179 ( .A(n13875), .B(n13874), .Z(n14012) );
  NANDN U14180 ( .A(n13877), .B(n13876), .Z(n13881) );
  OR U14181 ( .A(n13879), .B(n13878), .Z(n13880) );
  NAND U14182 ( .A(n13881), .B(n13880), .Z(n13978) );
  NAND U14183 ( .A(b[0]), .B(a[185]), .Z(n13882) );
  XNOR U14184 ( .A(b[1]), .B(n13882), .Z(n13884) );
  NAND U14185 ( .A(a[184]), .B(n98), .Z(n13883) );
  AND U14186 ( .A(n13884), .B(n13883), .Z(n13954) );
  XNOR U14187 ( .A(n20154), .B(n14062), .Z(n13963) );
  OR U14188 ( .A(n13963), .B(n20057), .Z(n13887) );
  NANDN U14189 ( .A(n13885), .B(n20098), .Z(n13886) );
  AND U14190 ( .A(n13887), .B(n13886), .Z(n13955) );
  XOR U14191 ( .A(n13954), .B(n13955), .Z(n13957) );
  NAND U14192 ( .A(a[169]), .B(b[15]), .Z(n13956) );
  XOR U14193 ( .A(n13957), .B(n13956), .Z(n13975) );
  NAND U14194 ( .A(n19722), .B(n13888), .Z(n13890) );
  XNOR U14195 ( .A(b[5]), .B(n14659), .Z(n13966) );
  NANDN U14196 ( .A(n19640), .B(n13966), .Z(n13889) );
  NAND U14197 ( .A(n13890), .B(n13889), .Z(n14000) );
  XNOR U14198 ( .A(n19714), .B(n14503), .Z(n13969) );
  NANDN U14199 ( .A(n13969), .B(n19766), .Z(n13893) );
  NANDN U14200 ( .A(n13891), .B(n19767), .Z(n13892) );
  NAND U14201 ( .A(n13893), .B(n13892), .Z(n13997) );
  NAND U14202 ( .A(n19554), .B(n13894), .Z(n13896) );
  IV U14203 ( .A(a[183]), .Z(n14815) );
  XNOR U14204 ( .A(b[3]), .B(n14815), .Z(n13972) );
  NANDN U14205 ( .A(n19521), .B(n13972), .Z(n13895) );
  AND U14206 ( .A(n13896), .B(n13895), .Z(n13998) );
  XNOR U14207 ( .A(n13997), .B(n13998), .Z(n13999) );
  XOR U14208 ( .A(n14000), .B(n13999), .Z(n13976) );
  XOR U14209 ( .A(n13975), .B(n13976), .Z(n13977) );
  XNOR U14210 ( .A(n13978), .B(n13977), .Z(n13948) );
  NAND U14211 ( .A(n13898), .B(n13897), .Z(n13902) );
  NAND U14212 ( .A(n13900), .B(n13899), .Z(n13901) );
  NAND U14213 ( .A(n13902), .B(n13901), .Z(n13949) );
  XOR U14214 ( .A(n13948), .B(n13949), .Z(n13951) );
  XNOR U14215 ( .A(n20052), .B(n14218), .Z(n13981) );
  OR U14216 ( .A(n13981), .B(n20020), .Z(n13905) );
  NANDN U14217 ( .A(n13903), .B(n19960), .Z(n13904) );
  NAND U14218 ( .A(n13905), .B(n13904), .Z(n13994) );
  XNOR U14219 ( .A(n102), .B(n13906), .Z(n13985) );
  OR U14220 ( .A(n13985), .B(n20121), .Z(n13909) );
  NANDN U14221 ( .A(n13907), .B(n20122), .Z(n13908) );
  NAND U14222 ( .A(n13909), .B(n13908), .Z(n13991) );
  XNOR U14223 ( .A(n19975), .B(n14347), .Z(n13988) );
  NANDN U14224 ( .A(n13988), .B(n19883), .Z(n13912) );
  NANDN U14225 ( .A(n13910), .B(n19937), .Z(n13911) );
  AND U14226 ( .A(n13912), .B(n13911), .Z(n13992) );
  XNOR U14227 ( .A(n13991), .B(n13992), .Z(n13993) );
  XNOR U14228 ( .A(n13994), .B(n13993), .Z(n14003) );
  NANDN U14229 ( .A(n13914), .B(n13913), .Z(n13918) );
  NAND U14230 ( .A(n13916), .B(n13915), .Z(n13917) );
  NAND U14231 ( .A(n13918), .B(n13917), .Z(n14004) );
  XNOR U14232 ( .A(n14003), .B(n14004), .Z(n14005) );
  NANDN U14233 ( .A(n13920), .B(n13919), .Z(n13924) );
  NAND U14234 ( .A(n13922), .B(n13921), .Z(n13923) );
  AND U14235 ( .A(n13924), .B(n13923), .Z(n14006) );
  XNOR U14236 ( .A(n14005), .B(n14006), .Z(n13950) );
  XNOR U14237 ( .A(n13951), .B(n13950), .Z(n14009) );
  NANDN U14238 ( .A(n13926), .B(n13925), .Z(n13930) );
  NAND U14239 ( .A(n13928), .B(n13927), .Z(n13929) );
  NAND U14240 ( .A(n13930), .B(n13929), .Z(n14010) );
  XNOR U14241 ( .A(n14009), .B(n14010), .Z(n14011) );
  XOR U14242 ( .A(n14012), .B(n14011), .Z(n13942) );
  NANDN U14243 ( .A(n13932), .B(n13931), .Z(n13936) );
  NANDN U14244 ( .A(n13934), .B(n13933), .Z(n13935) );
  NAND U14245 ( .A(n13936), .B(n13935), .Z(n13943) );
  XNOR U14246 ( .A(n13942), .B(n13943), .Z(n13944) );
  XNOR U14247 ( .A(n13945), .B(n13944), .Z(n14015) );
  XNOR U14248 ( .A(n14015), .B(sreg[425]), .Z(n14017) );
  NAND U14249 ( .A(n13937), .B(sreg[424]), .Z(n13941) );
  OR U14250 ( .A(n13939), .B(n13938), .Z(n13940) );
  AND U14251 ( .A(n13941), .B(n13940), .Z(n14016) );
  XOR U14252 ( .A(n14017), .B(n14016), .Z(c[425]) );
  NANDN U14253 ( .A(n13943), .B(n13942), .Z(n13947) );
  NAND U14254 ( .A(n13945), .B(n13944), .Z(n13946) );
  NAND U14255 ( .A(n13947), .B(n13946), .Z(n14023) );
  NANDN U14256 ( .A(n13949), .B(n13948), .Z(n13953) );
  OR U14257 ( .A(n13951), .B(n13950), .Z(n13952) );
  NAND U14258 ( .A(n13953), .B(n13952), .Z(n14090) );
  NANDN U14259 ( .A(n13955), .B(n13954), .Z(n13959) );
  OR U14260 ( .A(n13957), .B(n13956), .Z(n13958) );
  NAND U14261 ( .A(n13959), .B(n13958), .Z(n14056) );
  NAND U14262 ( .A(b[0]), .B(a[186]), .Z(n13960) );
  XNOR U14263 ( .A(b[1]), .B(n13960), .Z(n13962) );
  NAND U14264 ( .A(a[185]), .B(n98), .Z(n13961) );
  AND U14265 ( .A(n13962), .B(n13961), .Z(n14032) );
  XNOR U14266 ( .A(n20154), .B(n14113), .Z(n14041) );
  OR U14267 ( .A(n14041), .B(n20057), .Z(n13965) );
  NANDN U14268 ( .A(n13963), .B(n20098), .Z(n13964) );
  AND U14269 ( .A(n13965), .B(n13964), .Z(n14033) );
  XOR U14270 ( .A(n14032), .B(n14033), .Z(n14035) );
  NAND U14271 ( .A(a[170]), .B(b[15]), .Z(n14034) );
  XOR U14272 ( .A(n14035), .B(n14034), .Z(n14053) );
  NAND U14273 ( .A(n19722), .B(n13966), .Z(n13968) );
  XNOR U14274 ( .A(b[5]), .B(n14737), .Z(n14044) );
  NANDN U14275 ( .A(n19640), .B(n14044), .Z(n13967) );
  NAND U14276 ( .A(n13968), .B(n13967), .Z(n14078) );
  XNOR U14277 ( .A(n19714), .B(n14581), .Z(n14047) );
  NANDN U14278 ( .A(n14047), .B(n19766), .Z(n13971) );
  NANDN U14279 ( .A(n13969), .B(n19767), .Z(n13970) );
  NAND U14280 ( .A(n13971), .B(n13970), .Z(n14075) );
  NAND U14281 ( .A(n19554), .B(n13972), .Z(n13974) );
  IV U14282 ( .A(a[184]), .Z(n14893) );
  XNOR U14283 ( .A(b[3]), .B(n14893), .Z(n14050) );
  NANDN U14284 ( .A(n19521), .B(n14050), .Z(n13973) );
  AND U14285 ( .A(n13974), .B(n13973), .Z(n14076) );
  XNOR U14286 ( .A(n14075), .B(n14076), .Z(n14077) );
  XOR U14287 ( .A(n14078), .B(n14077), .Z(n14054) );
  XOR U14288 ( .A(n14053), .B(n14054), .Z(n14055) );
  XNOR U14289 ( .A(n14056), .B(n14055), .Z(n14026) );
  NAND U14290 ( .A(n13976), .B(n13975), .Z(n13980) );
  NAND U14291 ( .A(n13978), .B(n13977), .Z(n13979) );
  NAND U14292 ( .A(n13980), .B(n13979), .Z(n14027) );
  XOR U14293 ( .A(n14026), .B(n14027), .Z(n14029) );
  XNOR U14294 ( .A(n20052), .B(n14269), .Z(n14059) );
  OR U14295 ( .A(n14059), .B(n20020), .Z(n13983) );
  NANDN U14296 ( .A(n13981), .B(n19960), .Z(n13982) );
  NAND U14297 ( .A(n13983), .B(n13982), .Z(n14072) );
  XNOR U14298 ( .A(n102), .B(n13984), .Z(n14063) );
  OR U14299 ( .A(n14063), .B(n20121), .Z(n13987) );
  NANDN U14300 ( .A(n13985), .B(n20122), .Z(n13986) );
  NAND U14301 ( .A(n13987), .B(n13986), .Z(n14069) );
  XNOR U14302 ( .A(n19975), .B(n14425), .Z(n14066) );
  NANDN U14303 ( .A(n14066), .B(n19883), .Z(n13990) );
  NANDN U14304 ( .A(n13988), .B(n19937), .Z(n13989) );
  AND U14305 ( .A(n13990), .B(n13989), .Z(n14070) );
  XNOR U14306 ( .A(n14069), .B(n14070), .Z(n14071) );
  XNOR U14307 ( .A(n14072), .B(n14071), .Z(n14081) );
  NANDN U14308 ( .A(n13992), .B(n13991), .Z(n13996) );
  NAND U14309 ( .A(n13994), .B(n13993), .Z(n13995) );
  NAND U14310 ( .A(n13996), .B(n13995), .Z(n14082) );
  XNOR U14311 ( .A(n14081), .B(n14082), .Z(n14083) );
  NANDN U14312 ( .A(n13998), .B(n13997), .Z(n14002) );
  NAND U14313 ( .A(n14000), .B(n13999), .Z(n14001) );
  AND U14314 ( .A(n14002), .B(n14001), .Z(n14084) );
  XNOR U14315 ( .A(n14083), .B(n14084), .Z(n14028) );
  XNOR U14316 ( .A(n14029), .B(n14028), .Z(n14087) );
  NANDN U14317 ( .A(n14004), .B(n14003), .Z(n14008) );
  NAND U14318 ( .A(n14006), .B(n14005), .Z(n14007) );
  NAND U14319 ( .A(n14008), .B(n14007), .Z(n14088) );
  XNOR U14320 ( .A(n14087), .B(n14088), .Z(n14089) );
  XOR U14321 ( .A(n14090), .B(n14089), .Z(n14020) );
  NANDN U14322 ( .A(n14010), .B(n14009), .Z(n14014) );
  NANDN U14323 ( .A(n14012), .B(n14011), .Z(n14013) );
  NAND U14324 ( .A(n14014), .B(n14013), .Z(n14021) );
  XNOR U14325 ( .A(n14020), .B(n14021), .Z(n14022) );
  XNOR U14326 ( .A(n14023), .B(n14022), .Z(n14093) );
  XNOR U14327 ( .A(n14093), .B(sreg[426]), .Z(n14095) );
  NAND U14328 ( .A(n14015), .B(sreg[425]), .Z(n14019) );
  OR U14329 ( .A(n14017), .B(n14016), .Z(n14018) );
  AND U14330 ( .A(n14019), .B(n14018), .Z(n14094) );
  XOR U14331 ( .A(n14095), .B(n14094), .Z(c[426]) );
  NANDN U14332 ( .A(n14021), .B(n14020), .Z(n14025) );
  NAND U14333 ( .A(n14023), .B(n14022), .Z(n14024) );
  NAND U14334 ( .A(n14025), .B(n14024), .Z(n14101) );
  NANDN U14335 ( .A(n14027), .B(n14026), .Z(n14031) );
  OR U14336 ( .A(n14029), .B(n14028), .Z(n14030) );
  NAND U14337 ( .A(n14031), .B(n14030), .Z(n14168) );
  NANDN U14338 ( .A(n14033), .B(n14032), .Z(n14037) );
  OR U14339 ( .A(n14035), .B(n14034), .Z(n14036) );
  NAND U14340 ( .A(n14037), .B(n14036), .Z(n14156) );
  NAND U14341 ( .A(b[0]), .B(a[187]), .Z(n14038) );
  XNOR U14342 ( .A(b[1]), .B(n14038), .Z(n14040) );
  NAND U14343 ( .A(a[186]), .B(n98), .Z(n14039) );
  AND U14344 ( .A(n14040), .B(n14039), .Z(n14132) );
  XNOR U14345 ( .A(n20154), .B(n14218), .Z(n14141) );
  OR U14346 ( .A(n14141), .B(n20057), .Z(n14043) );
  NANDN U14347 ( .A(n14041), .B(n20098), .Z(n14042) );
  AND U14348 ( .A(n14043), .B(n14042), .Z(n14133) );
  XOR U14349 ( .A(n14132), .B(n14133), .Z(n14135) );
  NAND U14350 ( .A(a[171]), .B(b[15]), .Z(n14134) );
  XOR U14351 ( .A(n14135), .B(n14134), .Z(n14153) );
  NAND U14352 ( .A(n19722), .B(n14044), .Z(n14046) );
  XNOR U14353 ( .A(b[5]), .B(n14815), .Z(n14144) );
  NANDN U14354 ( .A(n19640), .B(n14144), .Z(n14045) );
  NAND U14355 ( .A(n14046), .B(n14045), .Z(n14129) );
  XNOR U14356 ( .A(n19714), .B(n14659), .Z(n14147) );
  NANDN U14357 ( .A(n14147), .B(n19766), .Z(n14049) );
  NANDN U14358 ( .A(n14047), .B(n19767), .Z(n14048) );
  NAND U14359 ( .A(n14049), .B(n14048), .Z(n14126) );
  NAND U14360 ( .A(n19554), .B(n14050), .Z(n14052) );
  IV U14361 ( .A(a[185]), .Z(n14971) );
  XNOR U14362 ( .A(b[3]), .B(n14971), .Z(n14150) );
  NANDN U14363 ( .A(n19521), .B(n14150), .Z(n14051) );
  AND U14364 ( .A(n14052), .B(n14051), .Z(n14127) );
  XNOR U14365 ( .A(n14126), .B(n14127), .Z(n14128) );
  XOR U14366 ( .A(n14129), .B(n14128), .Z(n14154) );
  XOR U14367 ( .A(n14153), .B(n14154), .Z(n14155) );
  XNOR U14368 ( .A(n14156), .B(n14155), .Z(n14104) );
  NAND U14369 ( .A(n14054), .B(n14053), .Z(n14058) );
  NAND U14370 ( .A(n14056), .B(n14055), .Z(n14057) );
  NAND U14371 ( .A(n14058), .B(n14057), .Z(n14105) );
  XOR U14372 ( .A(n14104), .B(n14105), .Z(n14107) );
  XNOR U14373 ( .A(n20052), .B(n14347), .Z(n14110) );
  OR U14374 ( .A(n14110), .B(n20020), .Z(n14061) );
  NANDN U14375 ( .A(n14059), .B(n19960), .Z(n14060) );
  NAND U14376 ( .A(n14061), .B(n14060), .Z(n14123) );
  XNOR U14377 ( .A(n102), .B(n14062), .Z(n14114) );
  OR U14378 ( .A(n14114), .B(n20121), .Z(n14065) );
  NANDN U14379 ( .A(n14063), .B(n20122), .Z(n14064) );
  NAND U14380 ( .A(n14065), .B(n14064), .Z(n14120) );
  XNOR U14381 ( .A(n19975), .B(n14503), .Z(n14117) );
  NANDN U14382 ( .A(n14117), .B(n19883), .Z(n14068) );
  NANDN U14383 ( .A(n14066), .B(n19937), .Z(n14067) );
  AND U14384 ( .A(n14068), .B(n14067), .Z(n14121) );
  XNOR U14385 ( .A(n14120), .B(n14121), .Z(n14122) );
  XNOR U14386 ( .A(n14123), .B(n14122), .Z(n14159) );
  NANDN U14387 ( .A(n14070), .B(n14069), .Z(n14074) );
  NAND U14388 ( .A(n14072), .B(n14071), .Z(n14073) );
  NAND U14389 ( .A(n14074), .B(n14073), .Z(n14160) );
  XNOR U14390 ( .A(n14159), .B(n14160), .Z(n14161) );
  NANDN U14391 ( .A(n14076), .B(n14075), .Z(n14080) );
  NAND U14392 ( .A(n14078), .B(n14077), .Z(n14079) );
  AND U14393 ( .A(n14080), .B(n14079), .Z(n14162) );
  XNOR U14394 ( .A(n14161), .B(n14162), .Z(n14106) );
  XNOR U14395 ( .A(n14107), .B(n14106), .Z(n14165) );
  NANDN U14396 ( .A(n14082), .B(n14081), .Z(n14086) );
  NAND U14397 ( .A(n14084), .B(n14083), .Z(n14085) );
  NAND U14398 ( .A(n14086), .B(n14085), .Z(n14166) );
  XNOR U14399 ( .A(n14165), .B(n14166), .Z(n14167) );
  XOR U14400 ( .A(n14168), .B(n14167), .Z(n14098) );
  NANDN U14401 ( .A(n14088), .B(n14087), .Z(n14092) );
  NANDN U14402 ( .A(n14090), .B(n14089), .Z(n14091) );
  NAND U14403 ( .A(n14092), .B(n14091), .Z(n14099) );
  XNOR U14404 ( .A(n14098), .B(n14099), .Z(n14100) );
  XNOR U14405 ( .A(n14101), .B(n14100), .Z(n14171) );
  XNOR U14406 ( .A(n14171), .B(sreg[427]), .Z(n14173) );
  NAND U14407 ( .A(n14093), .B(sreg[426]), .Z(n14097) );
  OR U14408 ( .A(n14095), .B(n14094), .Z(n14096) );
  AND U14409 ( .A(n14097), .B(n14096), .Z(n14172) );
  XOR U14410 ( .A(n14173), .B(n14172), .Z(c[427]) );
  NANDN U14411 ( .A(n14099), .B(n14098), .Z(n14103) );
  NAND U14412 ( .A(n14101), .B(n14100), .Z(n14102) );
  NAND U14413 ( .A(n14103), .B(n14102), .Z(n14179) );
  NANDN U14414 ( .A(n14105), .B(n14104), .Z(n14109) );
  OR U14415 ( .A(n14107), .B(n14106), .Z(n14108) );
  NAND U14416 ( .A(n14109), .B(n14108), .Z(n14246) );
  XNOR U14417 ( .A(n20052), .B(n14425), .Z(n14215) );
  OR U14418 ( .A(n14215), .B(n20020), .Z(n14112) );
  NANDN U14419 ( .A(n14110), .B(n19960), .Z(n14111) );
  NAND U14420 ( .A(n14112), .B(n14111), .Z(n14228) );
  XNOR U14421 ( .A(n102), .B(n14113), .Z(n14219) );
  OR U14422 ( .A(n14219), .B(n20121), .Z(n14116) );
  NANDN U14423 ( .A(n14114), .B(n20122), .Z(n14115) );
  NAND U14424 ( .A(n14116), .B(n14115), .Z(n14225) );
  XNOR U14425 ( .A(n19975), .B(n14581), .Z(n14222) );
  NANDN U14426 ( .A(n14222), .B(n19883), .Z(n14119) );
  NANDN U14427 ( .A(n14117), .B(n19937), .Z(n14118) );
  AND U14428 ( .A(n14119), .B(n14118), .Z(n14226) );
  XNOR U14429 ( .A(n14225), .B(n14226), .Z(n14227) );
  XNOR U14430 ( .A(n14228), .B(n14227), .Z(n14237) );
  NANDN U14431 ( .A(n14121), .B(n14120), .Z(n14125) );
  NAND U14432 ( .A(n14123), .B(n14122), .Z(n14124) );
  NAND U14433 ( .A(n14125), .B(n14124), .Z(n14238) );
  XNOR U14434 ( .A(n14237), .B(n14238), .Z(n14239) );
  NANDN U14435 ( .A(n14127), .B(n14126), .Z(n14131) );
  NAND U14436 ( .A(n14129), .B(n14128), .Z(n14130) );
  AND U14437 ( .A(n14131), .B(n14130), .Z(n14240) );
  XNOR U14438 ( .A(n14239), .B(n14240), .Z(n14184) );
  NANDN U14439 ( .A(n14133), .B(n14132), .Z(n14137) );
  OR U14440 ( .A(n14135), .B(n14134), .Z(n14136) );
  NAND U14441 ( .A(n14137), .B(n14136), .Z(n14212) );
  NAND U14442 ( .A(b[0]), .B(a[188]), .Z(n14138) );
  XNOR U14443 ( .A(b[1]), .B(n14138), .Z(n14140) );
  NAND U14444 ( .A(a[187]), .B(n98), .Z(n14139) );
  AND U14445 ( .A(n14140), .B(n14139), .Z(n14188) );
  XNOR U14446 ( .A(n20154), .B(n14269), .Z(n14197) );
  OR U14447 ( .A(n14197), .B(n20057), .Z(n14143) );
  NANDN U14448 ( .A(n14141), .B(n20098), .Z(n14142) );
  AND U14449 ( .A(n14143), .B(n14142), .Z(n14189) );
  XOR U14450 ( .A(n14188), .B(n14189), .Z(n14191) );
  NAND U14451 ( .A(a[172]), .B(b[15]), .Z(n14190) );
  XOR U14452 ( .A(n14191), .B(n14190), .Z(n14209) );
  NAND U14453 ( .A(n19722), .B(n14144), .Z(n14146) );
  XNOR U14454 ( .A(b[5]), .B(n14893), .Z(n14200) );
  NANDN U14455 ( .A(n19640), .B(n14200), .Z(n14145) );
  NAND U14456 ( .A(n14146), .B(n14145), .Z(n14234) );
  XNOR U14457 ( .A(n19714), .B(n14737), .Z(n14203) );
  NANDN U14458 ( .A(n14203), .B(n19766), .Z(n14149) );
  NANDN U14459 ( .A(n14147), .B(n19767), .Z(n14148) );
  NAND U14460 ( .A(n14149), .B(n14148), .Z(n14231) );
  NAND U14461 ( .A(n19554), .B(n14150), .Z(n14152) );
  IV U14462 ( .A(a[186]), .Z(n15049) );
  XNOR U14463 ( .A(b[3]), .B(n15049), .Z(n14206) );
  NANDN U14464 ( .A(n19521), .B(n14206), .Z(n14151) );
  AND U14465 ( .A(n14152), .B(n14151), .Z(n14232) );
  XNOR U14466 ( .A(n14231), .B(n14232), .Z(n14233) );
  XOR U14467 ( .A(n14234), .B(n14233), .Z(n14210) );
  XOR U14468 ( .A(n14209), .B(n14210), .Z(n14211) );
  XNOR U14469 ( .A(n14212), .B(n14211), .Z(n14182) );
  NAND U14470 ( .A(n14154), .B(n14153), .Z(n14158) );
  NAND U14471 ( .A(n14156), .B(n14155), .Z(n14157) );
  NAND U14472 ( .A(n14158), .B(n14157), .Z(n14183) );
  XOR U14473 ( .A(n14182), .B(n14183), .Z(n14185) );
  XNOR U14474 ( .A(n14184), .B(n14185), .Z(n14243) );
  NANDN U14475 ( .A(n14160), .B(n14159), .Z(n14164) );
  NAND U14476 ( .A(n14162), .B(n14161), .Z(n14163) );
  NAND U14477 ( .A(n14164), .B(n14163), .Z(n14244) );
  XNOR U14478 ( .A(n14243), .B(n14244), .Z(n14245) );
  XOR U14479 ( .A(n14246), .B(n14245), .Z(n14176) );
  NANDN U14480 ( .A(n14166), .B(n14165), .Z(n14170) );
  NANDN U14481 ( .A(n14168), .B(n14167), .Z(n14169) );
  NAND U14482 ( .A(n14170), .B(n14169), .Z(n14177) );
  XNOR U14483 ( .A(n14176), .B(n14177), .Z(n14178) );
  XNOR U14484 ( .A(n14179), .B(n14178), .Z(n14249) );
  XNOR U14485 ( .A(n14249), .B(sreg[428]), .Z(n14251) );
  NAND U14486 ( .A(n14171), .B(sreg[427]), .Z(n14175) );
  OR U14487 ( .A(n14173), .B(n14172), .Z(n14174) );
  AND U14488 ( .A(n14175), .B(n14174), .Z(n14250) );
  XOR U14489 ( .A(n14251), .B(n14250), .Z(c[428]) );
  NANDN U14490 ( .A(n14177), .B(n14176), .Z(n14181) );
  NAND U14491 ( .A(n14179), .B(n14178), .Z(n14180) );
  NAND U14492 ( .A(n14181), .B(n14180), .Z(n14257) );
  NANDN U14493 ( .A(n14183), .B(n14182), .Z(n14187) );
  OR U14494 ( .A(n14185), .B(n14184), .Z(n14186) );
  NAND U14495 ( .A(n14187), .B(n14186), .Z(n14324) );
  NANDN U14496 ( .A(n14189), .B(n14188), .Z(n14193) );
  OR U14497 ( .A(n14191), .B(n14190), .Z(n14192) );
  NAND U14498 ( .A(n14193), .B(n14192), .Z(n14312) );
  NAND U14499 ( .A(b[0]), .B(a[189]), .Z(n14194) );
  XNOR U14500 ( .A(b[1]), .B(n14194), .Z(n14196) );
  NAND U14501 ( .A(a[188]), .B(n98), .Z(n14195) );
  AND U14502 ( .A(n14196), .B(n14195), .Z(n14288) );
  XNOR U14503 ( .A(n20154), .B(n14347), .Z(n14297) );
  OR U14504 ( .A(n14297), .B(n20057), .Z(n14199) );
  NANDN U14505 ( .A(n14197), .B(n20098), .Z(n14198) );
  AND U14506 ( .A(n14199), .B(n14198), .Z(n14289) );
  XOR U14507 ( .A(n14288), .B(n14289), .Z(n14291) );
  NAND U14508 ( .A(a[173]), .B(b[15]), .Z(n14290) );
  XOR U14509 ( .A(n14291), .B(n14290), .Z(n14309) );
  NAND U14510 ( .A(n19722), .B(n14200), .Z(n14202) );
  XNOR U14511 ( .A(b[5]), .B(n14971), .Z(n14300) );
  NANDN U14512 ( .A(n19640), .B(n14300), .Z(n14201) );
  NAND U14513 ( .A(n14202), .B(n14201), .Z(n14285) );
  XNOR U14514 ( .A(n19714), .B(n14815), .Z(n14303) );
  NANDN U14515 ( .A(n14303), .B(n19766), .Z(n14205) );
  NANDN U14516 ( .A(n14203), .B(n19767), .Z(n14204) );
  NAND U14517 ( .A(n14205), .B(n14204), .Z(n14282) );
  NAND U14518 ( .A(n19554), .B(n14206), .Z(n14208) );
  IV U14519 ( .A(a[187]), .Z(n15127) );
  XNOR U14520 ( .A(b[3]), .B(n15127), .Z(n14306) );
  NANDN U14521 ( .A(n19521), .B(n14306), .Z(n14207) );
  AND U14522 ( .A(n14208), .B(n14207), .Z(n14283) );
  XNOR U14523 ( .A(n14282), .B(n14283), .Z(n14284) );
  XOR U14524 ( .A(n14285), .B(n14284), .Z(n14310) );
  XOR U14525 ( .A(n14309), .B(n14310), .Z(n14311) );
  XNOR U14526 ( .A(n14312), .B(n14311), .Z(n14260) );
  NAND U14527 ( .A(n14210), .B(n14209), .Z(n14214) );
  NAND U14528 ( .A(n14212), .B(n14211), .Z(n14213) );
  NAND U14529 ( .A(n14214), .B(n14213), .Z(n14261) );
  XOR U14530 ( .A(n14260), .B(n14261), .Z(n14263) );
  XNOR U14531 ( .A(n20052), .B(n14503), .Z(n14266) );
  OR U14532 ( .A(n14266), .B(n20020), .Z(n14217) );
  NANDN U14533 ( .A(n14215), .B(n19960), .Z(n14216) );
  NAND U14534 ( .A(n14217), .B(n14216), .Z(n14279) );
  XNOR U14535 ( .A(n102), .B(n14218), .Z(n14270) );
  OR U14536 ( .A(n14270), .B(n20121), .Z(n14221) );
  NANDN U14537 ( .A(n14219), .B(n20122), .Z(n14220) );
  NAND U14538 ( .A(n14221), .B(n14220), .Z(n14276) );
  XNOR U14539 ( .A(n19975), .B(n14659), .Z(n14273) );
  NANDN U14540 ( .A(n14273), .B(n19883), .Z(n14224) );
  NANDN U14541 ( .A(n14222), .B(n19937), .Z(n14223) );
  AND U14542 ( .A(n14224), .B(n14223), .Z(n14277) );
  XNOR U14543 ( .A(n14276), .B(n14277), .Z(n14278) );
  XNOR U14544 ( .A(n14279), .B(n14278), .Z(n14315) );
  NANDN U14545 ( .A(n14226), .B(n14225), .Z(n14230) );
  NAND U14546 ( .A(n14228), .B(n14227), .Z(n14229) );
  NAND U14547 ( .A(n14230), .B(n14229), .Z(n14316) );
  XNOR U14548 ( .A(n14315), .B(n14316), .Z(n14317) );
  NANDN U14549 ( .A(n14232), .B(n14231), .Z(n14236) );
  NAND U14550 ( .A(n14234), .B(n14233), .Z(n14235) );
  AND U14551 ( .A(n14236), .B(n14235), .Z(n14318) );
  XNOR U14552 ( .A(n14317), .B(n14318), .Z(n14262) );
  XNOR U14553 ( .A(n14263), .B(n14262), .Z(n14321) );
  NANDN U14554 ( .A(n14238), .B(n14237), .Z(n14242) );
  NAND U14555 ( .A(n14240), .B(n14239), .Z(n14241) );
  NAND U14556 ( .A(n14242), .B(n14241), .Z(n14322) );
  XNOR U14557 ( .A(n14321), .B(n14322), .Z(n14323) );
  XOR U14558 ( .A(n14324), .B(n14323), .Z(n14254) );
  NANDN U14559 ( .A(n14244), .B(n14243), .Z(n14248) );
  NANDN U14560 ( .A(n14246), .B(n14245), .Z(n14247) );
  NAND U14561 ( .A(n14248), .B(n14247), .Z(n14255) );
  XNOR U14562 ( .A(n14254), .B(n14255), .Z(n14256) );
  XNOR U14563 ( .A(n14257), .B(n14256), .Z(n14327) );
  XNOR U14564 ( .A(n14327), .B(sreg[429]), .Z(n14329) );
  NAND U14565 ( .A(n14249), .B(sreg[428]), .Z(n14253) );
  OR U14566 ( .A(n14251), .B(n14250), .Z(n14252) );
  AND U14567 ( .A(n14253), .B(n14252), .Z(n14328) );
  XOR U14568 ( .A(n14329), .B(n14328), .Z(c[429]) );
  NANDN U14569 ( .A(n14255), .B(n14254), .Z(n14259) );
  NAND U14570 ( .A(n14257), .B(n14256), .Z(n14258) );
  NAND U14571 ( .A(n14259), .B(n14258), .Z(n14335) );
  NANDN U14572 ( .A(n14261), .B(n14260), .Z(n14265) );
  OR U14573 ( .A(n14263), .B(n14262), .Z(n14264) );
  NAND U14574 ( .A(n14265), .B(n14264), .Z(n14402) );
  XNOR U14575 ( .A(n20052), .B(n14581), .Z(n14344) );
  OR U14576 ( .A(n14344), .B(n20020), .Z(n14268) );
  NANDN U14577 ( .A(n14266), .B(n19960), .Z(n14267) );
  NAND U14578 ( .A(n14268), .B(n14267), .Z(n14357) );
  XNOR U14579 ( .A(n102), .B(n14269), .Z(n14348) );
  OR U14580 ( .A(n14348), .B(n20121), .Z(n14272) );
  NANDN U14581 ( .A(n14270), .B(n20122), .Z(n14271) );
  NAND U14582 ( .A(n14272), .B(n14271), .Z(n14354) );
  XNOR U14583 ( .A(n19975), .B(n14737), .Z(n14351) );
  NANDN U14584 ( .A(n14351), .B(n19883), .Z(n14275) );
  NANDN U14585 ( .A(n14273), .B(n19937), .Z(n14274) );
  AND U14586 ( .A(n14275), .B(n14274), .Z(n14355) );
  XNOR U14587 ( .A(n14354), .B(n14355), .Z(n14356) );
  XNOR U14588 ( .A(n14357), .B(n14356), .Z(n14393) );
  NANDN U14589 ( .A(n14277), .B(n14276), .Z(n14281) );
  NAND U14590 ( .A(n14279), .B(n14278), .Z(n14280) );
  NAND U14591 ( .A(n14281), .B(n14280), .Z(n14394) );
  XNOR U14592 ( .A(n14393), .B(n14394), .Z(n14395) );
  NANDN U14593 ( .A(n14283), .B(n14282), .Z(n14287) );
  NAND U14594 ( .A(n14285), .B(n14284), .Z(n14286) );
  AND U14595 ( .A(n14287), .B(n14286), .Z(n14396) );
  XNOR U14596 ( .A(n14395), .B(n14396), .Z(n14340) );
  NANDN U14597 ( .A(n14289), .B(n14288), .Z(n14293) );
  OR U14598 ( .A(n14291), .B(n14290), .Z(n14292) );
  NAND U14599 ( .A(n14293), .B(n14292), .Z(n14390) );
  NAND U14600 ( .A(b[0]), .B(a[190]), .Z(n14294) );
  XNOR U14601 ( .A(b[1]), .B(n14294), .Z(n14296) );
  NAND U14602 ( .A(a[189]), .B(n98), .Z(n14295) );
  AND U14603 ( .A(n14296), .B(n14295), .Z(n14366) );
  XNOR U14604 ( .A(n20154), .B(n14425), .Z(n14375) );
  OR U14605 ( .A(n14375), .B(n20057), .Z(n14299) );
  NANDN U14606 ( .A(n14297), .B(n20098), .Z(n14298) );
  AND U14607 ( .A(n14299), .B(n14298), .Z(n14367) );
  XOR U14608 ( .A(n14366), .B(n14367), .Z(n14369) );
  NAND U14609 ( .A(a[174]), .B(b[15]), .Z(n14368) );
  XOR U14610 ( .A(n14369), .B(n14368), .Z(n14387) );
  NAND U14611 ( .A(n19722), .B(n14300), .Z(n14302) );
  XNOR U14612 ( .A(b[5]), .B(n15049), .Z(n14378) );
  NANDN U14613 ( .A(n19640), .B(n14378), .Z(n14301) );
  NAND U14614 ( .A(n14302), .B(n14301), .Z(n14363) );
  XNOR U14615 ( .A(n19714), .B(n14893), .Z(n14381) );
  NANDN U14616 ( .A(n14381), .B(n19766), .Z(n14305) );
  NANDN U14617 ( .A(n14303), .B(n19767), .Z(n14304) );
  NAND U14618 ( .A(n14305), .B(n14304), .Z(n14360) );
  NAND U14619 ( .A(n19554), .B(n14306), .Z(n14308) );
  IV U14620 ( .A(a[188]), .Z(n15204) );
  XNOR U14621 ( .A(b[3]), .B(n15204), .Z(n14384) );
  NANDN U14622 ( .A(n19521), .B(n14384), .Z(n14307) );
  AND U14623 ( .A(n14308), .B(n14307), .Z(n14361) );
  XNOR U14624 ( .A(n14360), .B(n14361), .Z(n14362) );
  XOR U14625 ( .A(n14363), .B(n14362), .Z(n14388) );
  XOR U14626 ( .A(n14387), .B(n14388), .Z(n14389) );
  XNOR U14627 ( .A(n14390), .B(n14389), .Z(n14338) );
  NAND U14628 ( .A(n14310), .B(n14309), .Z(n14314) );
  NAND U14629 ( .A(n14312), .B(n14311), .Z(n14313) );
  NAND U14630 ( .A(n14314), .B(n14313), .Z(n14339) );
  XOR U14631 ( .A(n14338), .B(n14339), .Z(n14341) );
  XNOR U14632 ( .A(n14340), .B(n14341), .Z(n14399) );
  NANDN U14633 ( .A(n14316), .B(n14315), .Z(n14320) );
  NAND U14634 ( .A(n14318), .B(n14317), .Z(n14319) );
  NAND U14635 ( .A(n14320), .B(n14319), .Z(n14400) );
  XNOR U14636 ( .A(n14399), .B(n14400), .Z(n14401) );
  XOR U14637 ( .A(n14402), .B(n14401), .Z(n14332) );
  NANDN U14638 ( .A(n14322), .B(n14321), .Z(n14326) );
  NANDN U14639 ( .A(n14324), .B(n14323), .Z(n14325) );
  NAND U14640 ( .A(n14326), .B(n14325), .Z(n14333) );
  XNOR U14641 ( .A(n14332), .B(n14333), .Z(n14334) );
  XNOR U14642 ( .A(n14335), .B(n14334), .Z(n14405) );
  XNOR U14643 ( .A(n14405), .B(sreg[430]), .Z(n14407) );
  NAND U14644 ( .A(n14327), .B(sreg[429]), .Z(n14331) );
  OR U14645 ( .A(n14329), .B(n14328), .Z(n14330) );
  AND U14646 ( .A(n14331), .B(n14330), .Z(n14406) );
  XOR U14647 ( .A(n14407), .B(n14406), .Z(c[430]) );
  NANDN U14648 ( .A(n14333), .B(n14332), .Z(n14337) );
  NAND U14649 ( .A(n14335), .B(n14334), .Z(n14336) );
  NAND U14650 ( .A(n14337), .B(n14336), .Z(n14413) );
  NANDN U14651 ( .A(n14339), .B(n14338), .Z(n14343) );
  OR U14652 ( .A(n14341), .B(n14340), .Z(n14342) );
  NAND U14653 ( .A(n14343), .B(n14342), .Z(n14480) );
  XNOR U14654 ( .A(n20052), .B(n14659), .Z(n14422) );
  OR U14655 ( .A(n14422), .B(n20020), .Z(n14346) );
  NANDN U14656 ( .A(n14344), .B(n19960), .Z(n14345) );
  NAND U14657 ( .A(n14346), .B(n14345), .Z(n14435) );
  XNOR U14658 ( .A(n102), .B(n14347), .Z(n14426) );
  OR U14659 ( .A(n14426), .B(n20121), .Z(n14350) );
  NANDN U14660 ( .A(n14348), .B(n20122), .Z(n14349) );
  NAND U14661 ( .A(n14350), .B(n14349), .Z(n14432) );
  XNOR U14662 ( .A(n19975), .B(n14815), .Z(n14429) );
  NANDN U14663 ( .A(n14429), .B(n19883), .Z(n14353) );
  NANDN U14664 ( .A(n14351), .B(n19937), .Z(n14352) );
  AND U14665 ( .A(n14353), .B(n14352), .Z(n14433) );
  XNOR U14666 ( .A(n14432), .B(n14433), .Z(n14434) );
  XNOR U14667 ( .A(n14435), .B(n14434), .Z(n14471) );
  NANDN U14668 ( .A(n14355), .B(n14354), .Z(n14359) );
  NAND U14669 ( .A(n14357), .B(n14356), .Z(n14358) );
  NAND U14670 ( .A(n14359), .B(n14358), .Z(n14472) );
  XNOR U14671 ( .A(n14471), .B(n14472), .Z(n14473) );
  NANDN U14672 ( .A(n14361), .B(n14360), .Z(n14365) );
  NAND U14673 ( .A(n14363), .B(n14362), .Z(n14364) );
  AND U14674 ( .A(n14365), .B(n14364), .Z(n14474) );
  XNOR U14675 ( .A(n14473), .B(n14474), .Z(n14418) );
  NANDN U14676 ( .A(n14367), .B(n14366), .Z(n14371) );
  OR U14677 ( .A(n14369), .B(n14368), .Z(n14370) );
  NAND U14678 ( .A(n14371), .B(n14370), .Z(n14468) );
  NAND U14679 ( .A(b[0]), .B(a[191]), .Z(n14372) );
  XNOR U14680 ( .A(b[1]), .B(n14372), .Z(n14374) );
  NAND U14681 ( .A(a[190]), .B(n98), .Z(n14373) );
  AND U14682 ( .A(n14374), .B(n14373), .Z(n14444) );
  XNOR U14683 ( .A(n20154), .B(n14503), .Z(n14453) );
  OR U14684 ( .A(n14453), .B(n20057), .Z(n14377) );
  NANDN U14685 ( .A(n14375), .B(n20098), .Z(n14376) );
  AND U14686 ( .A(n14377), .B(n14376), .Z(n14445) );
  XOR U14687 ( .A(n14444), .B(n14445), .Z(n14447) );
  NAND U14688 ( .A(a[175]), .B(b[15]), .Z(n14446) );
  XOR U14689 ( .A(n14447), .B(n14446), .Z(n14465) );
  NAND U14690 ( .A(n19722), .B(n14378), .Z(n14380) );
  XNOR U14691 ( .A(b[5]), .B(n15127), .Z(n14456) );
  NANDN U14692 ( .A(n19640), .B(n14456), .Z(n14379) );
  NAND U14693 ( .A(n14380), .B(n14379), .Z(n14441) );
  XNOR U14694 ( .A(n19714), .B(n14971), .Z(n14459) );
  NANDN U14695 ( .A(n14459), .B(n19766), .Z(n14383) );
  NANDN U14696 ( .A(n14381), .B(n19767), .Z(n14382) );
  NAND U14697 ( .A(n14383), .B(n14382), .Z(n14438) );
  NAND U14698 ( .A(n19554), .B(n14384), .Z(n14386) );
  IV U14699 ( .A(a[189]), .Z(n15280) );
  XNOR U14700 ( .A(b[3]), .B(n15280), .Z(n14462) );
  NANDN U14701 ( .A(n19521), .B(n14462), .Z(n14385) );
  AND U14702 ( .A(n14386), .B(n14385), .Z(n14439) );
  XNOR U14703 ( .A(n14438), .B(n14439), .Z(n14440) );
  XOR U14704 ( .A(n14441), .B(n14440), .Z(n14466) );
  XOR U14705 ( .A(n14465), .B(n14466), .Z(n14467) );
  XNOR U14706 ( .A(n14468), .B(n14467), .Z(n14416) );
  NAND U14707 ( .A(n14388), .B(n14387), .Z(n14392) );
  NAND U14708 ( .A(n14390), .B(n14389), .Z(n14391) );
  NAND U14709 ( .A(n14392), .B(n14391), .Z(n14417) );
  XOR U14710 ( .A(n14416), .B(n14417), .Z(n14419) );
  XNOR U14711 ( .A(n14418), .B(n14419), .Z(n14477) );
  NANDN U14712 ( .A(n14394), .B(n14393), .Z(n14398) );
  NAND U14713 ( .A(n14396), .B(n14395), .Z(n14397) );
  NAND U14714 ( .A(n14398), .B(n14397), .Z(n14478) );
  XNOR U14715 ( .A(n14477), .B(n14478), .Z(n14479) );
  XOR U14716 ( .A(n14480), .B(n14479), .Z(n14410) );
  NANDN U14717 ( .A(n14400), .B(n14399), .Z(n14404) );
  NANDN U14718 ( .A(n14402), .B(n14401), .Z(n14403) );
  NAND U14719 ( .A(n14404), .B(n14403), .Z(n14411) );
  XNOR U14720 ( .A(n14410), .B(n14411), .Z(n14412) );
  XNOR U14721 ( .A(n14413), .B(n14412), .Z(n14483) );
  XNOR U14722 ( .A(n14483), .B(sreg[431]), .Z(n14485) );
  NAND U14723 ( .A(n14405), .B(sreg[430]), .Z(n14409) );
  OR U14724 ( .A(n14407), .B(n14406), .Z(n14408) );
  AND U14725 ( .A(n14409), .B(n14408), .Z(n14484) );
  XOR U14726 ( .A(n14485), .B(n14484), .Z(c[431]) );
  NANDN U14727 ( .A(n14411), .B(n14410), .Z(n14415) );
  NAND U14728 ( .A(n14413), .B(n14412), .Z(n14414) );
  NAND U14729 ( .A(n14415), .B(n14414), .Z(n14491) );
  NANDN U14730 ( .A(n14417), .B(n14416), .Z(n14421) );
  OR U14731 ( .A(n14419), .B(n14418), .Z(n14420) );
  NAND U14732 ( .A(n14421), .B(n14420), .Z(n14558) );
  XNOR U14733 ( .A(n20052), .B(n14737), .Z(n14500) );
  OR U14734 ( .A(n14500), .B(n20020), .Z(n14424) );
  NANDN U14735 ( .A(n14422), .B(n19960), .Z(n14423) );
  NAND U14736 ( .A(n14424), .B(n14423), .Z(n14513) );
  XNOR U14737 ( .A(n102), .B(n14425), .Z(n14504) );
  OR U14738 ( .A(n14504), .B(n20121), .Z(n14428) );
  NANDN U14739 ( .A(n14426), .B(n20122), .Z(n14427) );
  NAND U14740 ( .A(n14428), .B(n14427), .Z(n14510) );
  XNOR U14741 ( .A(n19975), .B(n14893), .Z(n14507) );
  NANDN U14742 ( .A(n14507), .B(n19883), .Z(n14431) );
  NANDN U14743 ( .A(n14429), .B(n19937), .Z(n14430) );
  AND U14744 ( .A(n14431), .B(n14430), .Z(n14511) );
  XNOR U14745 ( .A(n14510), .B(n14511), .Z(n14512) );
  XNOR U14746 ( .A(n14513), .B(n14512), .Z(n14549) );
  NANDN U14747 ( .A(n14433), .B(n14432), .Z(n14437) );
  NAND U14748 ( .A(n14435), .B(n14434), .Z(n14436) );
  NAND U14749 ( .A(n14437), .B(n14436), .Z(n14550) );
  XNOR U14750 ( .A(n14549), .B(n14550), .Z(n14551) );
  NANDN U14751 ( .A(n14439), .B(n14438), .Z(n14443) );
  NAND U14752 ( .A(n14441), .B(n14440), .Z(n14442) );
  AND U14753 ( .A(n14443), .B(n14442), .Z(n14552) );
  XNOR U14754 ( .A(n14551), .B(n14552), .Z(n14496) );
  NANDN U14755 ( .A(n14445), .B(n14444), .Z(n14449) );
  OR U14756 ( .A(n14447), .B(n14446), .Z(n14448) );
  NAND U14757 ( .A(n14449), .B(n14448), .Z(n14546) );
  NAND U14758 ( .A(b[0]), .B(a[192]), .Z(n14450) );
  XNOR U14759 ( .A(b[1]), .B(n14450), .Z(n14452) );
  NAND U14760 ( .A(a[191]), .B(n98), .Z(n14451) );
  AND U14761 ( .A(n14452), .B(n14451), .Z(n14522) );
  XNOR U14762 ( .A(n20154), .B(n14581), .Z(n14531) );
  OR U14763 ( .A(n14531), .B(n20057), .Z(n14455) );
  NANDN U14764 ( .A(n14453), .B(n20098), .Z(n14454) );
  AND U14765 ( .A(n14455), .B(n14454), .Z(n14523) );
  XOR U14766 ( .A(n14522), .B(n14523), .Z(n14525) );
  NAND U14767 ( .A(a[176]), .B(b[15]), .Z(n14524) );
  XOR U14768 ( .A(n14525), .B(n14524), .Z(n14543) );
  NAND U14769 ( .A(n19722), .B(n14456), .Z(n14458) );
  XNOR U14770 ( .A(b[5]), .B(n15204), .Z(n14534) );
  NANDN U14771 ( .A(n19640), .B(n14534), .Z(n14457) );
  NAND U14772 ( .A(n14458), .B(n14457), .Z(n14519) );
  XNOR U14773 ( .A(n19714), .B(n15049), .Z(n14537) );
  NANDN U14774 ( .A(n14537), .B(n19766), .Z(n14461) );
  NANDN U14775 ( .A(n14459), .B(n19767), .Z(n14460) );
  NAND U14776 ( .A(n14461), .B(n14460), .Z(n14516) );
  NAND U14777 ( .A(n19554), .B(n14462), .Z(n14464) );
  IV U14778 ( .A(a[190]), .Z(n15385) );
  XNOR U14779 ( .A(b[3]), .B(n15385), .Z(n14540) );
  NANDN U14780 ( .A(n19521), .B(n14540), .Z(n14463) );
  AND U14781 ( .A(n14464), .B(n14463), .Z(n14517) );
  XNOR U14782 ( .A(n14516), .B(n14517), .Z(n14518) );
  XOR U14783 ( .A(n14519), .B(n14518), .Z(n14544) );
  XOR U14784 ( .A(n14543), .B(n14544), .Z(n14545) );
  XNOR U14785 ( .A(n14546), .B(n14545), .Z(n14494) );
  NAND U14786 ( .A(n14466), .B(n14465), .Z(n14470) );
  NAND U14787 ( .A(n14468), .B(n14467), .Z(n14469) );
  NAND U14788 ( .A(n14470), .B(n14469), .Z(n14495) );
  XOR U14789 ( .A(n14494), .B(n14495), .Z(n14497) );
  XNOR U14790 ( .A(n14496), .B(n14497), .Z(n14555) );
  NANDN U14791 ( .A(n14472), .B(n14471), .Z(n14476) );
  NAND U14792 ( .A(n14474), .B(n14473), .Z(n14475) );
  NAND U14793 ( .A(n14476), .B(n14475), .Z(n14556) );
  XNOR U14794 ( .A(n14555), .B(n14556), .Z(n14557) );
  XOR U14795 ( .A(n14558), .B(n14557), .Z(n14488) );
  NANDN U14796 ( .A(n14478), .B(n14477), .Z(n14482) );
  NANDN U14797 ( .A(n14480), .B(n14479), .Z(n14481) );
  NAND U14798 ( .A(n14482), .B(n14481), .Z(n14489) );
  XNOR U14799 ( .A(n14488), .B(n14489), .Z(n14490) );
  XNOR U14800 ( .A(n14491), .B(n14490), .Z(n14561) );
  XNOR U14801 ( .A(n14561), .B(sreg[432]), .Z(n14563) );
  NAND U14802 ( .A(n14483), .B(sreg[431]), .Z(n14487) );
  OR U14803 ( .A(n14485), .B(n14484), .Z(n14486) );
  AND U14804 ( .A(n14487), .B(n14486), .Z(n14562) );
  XOR U14805 ( .A(n14563), .B(n14562), .Z(c[432]) );
  NANDN U14806 ( .A(n14489), .B(n14488), .Z(n14493) );
  NAND U14807 ( .A(n14491), .B(n14490), .Z(n14492) );
  NAND U14808 ( .A(n14493), .B(n14492), .Z(n14569) );
  NANDN U14809 ( .A(n14495), .B(n14494), .Z(n14499) );
  OR U14810 ( .A(n14497), .B(n14496), .Z(n14498) );
  NAND U14811 ( .A(n14499), .B(n14498), .Z(n14636) );
  XNOR U14812 ( .A(n20052), .B(n14815), .Z(n14578) );
  OR U14813 ( .A(n14578), .B(n20020), .Z(n14502) );
  NANDN U14814 ( .A(n14500), .B(n19960), .Z(n14501) );
  NAND U14815 ( .A(n14502), .B(n14501), .Z(n14591) );
  XNOR U14816 ( .A(n102), .B(n14503), .Z(n14582) );
  OR U14817 ( .A(n14582), .B(n20121), .Z(n14506) );
  NANDN U14818 ( .A(n14504), .B(n20122), .Z(n14505) );
  NAND U14819 ( .A(n14506), .B(n14505), .Z(n14588) );
  XNOR U14820 ( .A(n19975), .B(n14971), .Z(n14585) );
  NANDN U14821 ( .A(n14585), .B(n19883), .Z(n14509) );
  NANDN U14822 ( .A(n14507), .B(n19937), .Z(n14508) );
  AND U14823 ( .A(n14509), .B(n14508), .Z(n14589) );
  XNOR U14824 ( .A(n14588), .B(n14589), .Z(n14590) );
  XNOR U14825 ( .A(n14591), .B(n14590), .Z(n14627) );
  NANDN U14826 ( .A(n14511), .B(n14510), .Z(n14515) );
  NAND U14827 ( .A(n14513), .B(n14512), .Z(n14514) );
  NAND U14828 ( .A(n14515), .B(n14514), .Z(n14628) );
  XNOR U14829 ( .A(n14627), .B(n14628), .Z(n14629) );
  NANDN U14830 ( .A(n14517), .B(n14516), .Z(n14521) );
  NAND U14831 ( .A(n14519), .B(n14518), .Z(n14520) );
  AND U14832 ( .A(n14521), .B(n14520), .Z(n14630) );
  XNOR U14833 ( .A(n14629), .B(n14630), .Z(n14574) );
  NANDN U14834 ( .A(n14523), .B(n14522), .Z(n14527) );
  OR U14835 ( .A(n14525), .B(n14524), .Z(n14526) );
  NAND U14836 ( .A(n14527), .B(n14526), .Z(n14624) );
  NAND U14837 ( .A(b[0]), .B(a[193]), .Z(n14528) );
  XNOR U14838 ( .A(b[1]), .B(n14528), .Z(n14530) );
  NAND U14839 ( .A(a[192]), .B(n98), .Z(n14529) );
  AND U14840 ( .A(n14530), .B(n14529), .Z(n14600) );
  XNOR U14841 ( .A(n20154), .B(n14659), .Z(n14609) );
  OR U14842 ( .A(n14609), .B(n20057), .Z(n14533) );
  NANDN U14843 ( .A(n14531), .B(n20098), .Z(n14532) );
  AND U14844 ( .A(n14533), .B(n14532), .Z(n14601) );
  XOR U14845 ( .A(n14600), .B(n14601), .Z(n14603) );
  NAND U14846 ( .A(a[177]), .B(b[15]), .Z(n14602) );
  XOR U14847 ( .A(n14603), .B(n14602), .Z(n14621) );
  NAND U14848 ( .A(n19722), .B(n14534), .Z(n14536) );
  XNOR U14849 ( .A(b[5]), .B(n15280), .Z(n14612) );
  NANDN U14850 ( .A(n19640), .B(n14612), .Z(n14535) );
  NAND U14851 ( .A(n14536), .B(n14535), .Z(n14597) );
  XNOR U14852 ( .A(n19714), .B(n15127), .Z(n14615) );
  NANDN U14853 ( .A(n14615), .B(n19766), .Z(n14539) );
  NANDN U14854 ( .A(n14537), .B(n19767), .Z(n14538) );
  NAND U14855 ( .A(n14539), .B(n14538), .Z(n14594) );
  NAND U14856 ( .A(n19554), .B(n14540), .Z(n14542) );
  IV U14857 ( .A(a[191]), .Z(n15436) );
  XNOR U14858 ( .A(b[3]), .B(n15436), .Z(n14618) );
  NANDN U14859 ( .A(n19521), .B(n14618), .Z(n14541) );
  AND U14860 ( .A(n14542), .B(n14541), .Z(n14595) );
  XNOR U14861 ( .A(n14594), .B(n14595), .Z(n14596) );
  XOR U14862 ( .A(n14597), .B(n14596), .Z(n14622) );
  XOR U14863 ( .A(n14621), .B(n14622), .Z(n14623) );
  XNOR U14864 ( .A(n14624), .B(n14623), .Z(n14572) );
  NAND U14865 ( .A(n14544), .B(n14543), .Z(n14548) );
  NAND U14866 ( .A(n14546), .B(n14545), .Z(n14547) );
  NAND U14867 ( .A(n14548), .B(n14547), .Z(n14573) );
  XOR U14868 ( .A(n14572), .B(n14573), .Z(n14575) );
  XNOR U14869 ( .A(n14574), .B(n14575), .Z(n14633) );
  NANDN U14870 ( .A(n14550), .B(n14549), .Z(n14554) );
  NAND U14871 ( .A(n14552), .B(n14551), .Z(n14553) );
  NAND U14872 ( .A(n14554), .B(n14553), .Z(n14634) );
  XNOR U14873 ( .A(n14633), .B(n14634), .Z(n14635) );
  XOR U14874 ( .A(n14636), .B(n14635), .Z(n14566) );
  NANDN U14875 ( .A(n14556), .B(n14555), .Z(n14560) );
  NANDN U14876 ( .A(n14558), .B(n14557), .Z(n14559) );
  NAND U14877 ( .A(n14560), .B(n14559), .Z(n14567) );
  XNOR U14878 ( .A(n14566), .B(n14567), .Z(n14568) );
  XNOR U14879 ( .A(n14569), .B(n14568), .Z(n14639) );
  XNOR U14880 ( .A(n14639), .B(sreg[433]), .Z(n14641) );
  NAND U14881 ( .A(n14561), .B(sreg[432]), .Z(n14565) );
  OR U14882 ( .A(n14563), .B(n14562), .Z(n14564) );
  AND U14883 ( .A(n14565), .B(n14564), .Z(n14640) );
  XOR U14884 ( .A(n14641), .B(n14640), .Z(c[433]) );
  NANDN U14885 ( .A(n14567), .B(n14566), .Z(n14571) );
  NAND U14886 ( .A(n14569), .B(n14568), .Z(n14570) );
  NAND U14887 ( .A(n14571), .B(n14570), .Z(n14647) );
  NANDN U14888 ( .A(n14573), .B(n14572), .Z(n14577) );
  OR U14889 ( .A(n14575), .B(n14574), .Z(n14576) );
  NAND U14890 ( .A(n14577), .B(n14576), .Z(n14714) );
  XNOR U14891 ( .A(n20052), .B(n14893), .Z(n14656) );
  OR U14892 ( .A(n14656), .B(n20020), .Z(n14580) );
  NANDN U14893 ( .A(n14578), .B(n19960), .Z(n14579) );
  NAND U14894 ( .A(n14580), .B(n14579), .Z(n14669) );
  XNOR U14895 ( .A(n102), .B(n14581), .Z(n14660) );
  OR U14896 ( .A(n14660), .B(n20121), .Z(n14584) );
  NANDN U14897 ( .A(n14582), .B(n20122), .Z(n14583) );
  NAND U14898 ( .A(n14584), .B(n14583), .Z(n14666) );
  XNOR U14899 ( .A(n19975), .B(n15049), .Z(n14663) );
  NANDN U14900 ( .A(n14663), .B(n19883), .Z(n14587) );
  NANDN U14901 ( .A(n14585), .B(n19937), .Z(n14586) );
  AND U14902 ( .A(n14587), .B(n14586), .Z(n14667) );
  XNOR U14903 ( .A(n14666), .B(n14667), .Z(n14668) );
  XNOR U14904 ( .A(n14669), .B(n14668), .Z(n14705) );
  NANDN U14905 ( .A(n14589), .B(n14588), .Z(n14593) );
  NAND U14906 ( .A(n14591), .B(n14590), .Z(n14592) );
  NAND U14907 ( .A(n14593), .B(n14592), .Z(n14706) );
  XNOR U14908 ( .A(n14705), .B(n14706), .Z(n14707) );
  NANDN U14909 ( .A(n14595), .B(n14594), .Z(n14599) );
  NAND U14910 ( .A(n14597), .B(n14596), .Z(n14598) );
  AND U14911 ( .A(n14599), .B(n14598), .Z(n14708) );
  XNOR U14912 ( .A(n14707), .B(n14708), .Z(n14652) );
  NANDN U14913 ( .A(n14601), .B(n14600), .Z(n14605) );
  OR U14914 ( .A(n14603), .B(n14602), .Z(n14604) );
  NAND U14915 ( .A(n14605), .B(n14604), .Z(n14702) );
  NAND U14916 ( .A(b[0]), .B(a[194]), .Z(n14606) );
  XNOR U14917 ( .A(b[1]), .B(n14606), .Z(n14608) );
  NAND U14918 ( .A(a[193]), .B(n98), .Z(n14607) );
  AND U14919 ( .A(n14608), .B(n14607), .Z(n14678) );
  XNOR U14920 ( .A(n20154), .B(n14737), .Z(n14684) );
  OR U14921 ( .A(n14684), .B(n20057), .Z(n14611) );
  NANDN U14922 ( .A(n14609), .B(n20098), .Z(n14610) );
  AND U14923 ( .A(n14611), .B(n14610), .Z(n14679) );
  XOR U14924 ( .A(n14678), .B(n14679), .Z(n14681) );
  NAND U14925 ( .A(a[178]), .B(b[15]), .Z(n14680) );
  XOR U14926 ( .A(n14681), .B(n14680), .Z(n14699) );
  NAND U14927 ( .A(n19722), .B(n14612), .Z(n14614) );
  XNOR U14928 ( .A(b[5]), .B(n15385), .Z(n14690) );
  NANDN U14929 ( .A(n19640), .B(n14690), .Z(n14613) );
  NAND U14930 ( .A(n14614), .B(n14613), .Z(n14675) );
  XNOR U14931 ( .A(n19714), .B(n15204), .Z(n14693) );
  NANDN U14932 ( .A(n14693), .B(n19766), .Z(n14617) );
  NANDN U14933 ( .A(n14615), .B(n19767), .Z(n14616) );
  NAND U14934 ( .A(n14617), .B(n14616), .Z(n14672) );
  NAND U14935 ( .A(n19554), .B(n14618), .Z(n14620) );
  IV U14936 ( .A(a[192]), .Z(n15514) );
  XNOR U14937 ( .A(b[3]), .B(n15514), .Z(n14696) );
  NANDN U14938 ( .A(n19521), .B(n14696), .Z(n14619) );
  AND U14939 ( .A(n14620), .B(n14619), .Z(n14673) );
  XNOR U14940 ( .A(n14672), .B(n14673), .Z(n14674) );
  XOR U14941 ( .A(n14675), .B(n14674), .Z(n14700) );
  XOR U14942 ( .A(n14699), .B(n14700), .Z(n14701) );
  XNOR U14943 ( .A(n14702), .B(n14701), .Z(n14650) );
  NAND U14944 ( .A(n14622), .B(n14621), .Z(n14626) );
  NAND U14945 ( .A(n14624), .B(n14623), .Z(n14625) );
  NAND U14946 ( .A(n14626), .B(n14625), .Z(n14651) );
  XOR U14947 ( .A(n14650), .B(n14651), .Z(n14653) );
  XNOR U14948 ( .A(n14652), .B(n14653), .Z(n14711) );
  NANDN U14949 ( .A(n14628), .B(n14627), .Z(n14632) );
  NAND U14950 ( .A(n14630), .B(n14629), .Z(n14631) );
  NAND U14951 ( .A(n14632), .B(n14631), .Z(n14712) );
  XNOR U14952 ( .A(n14711), .B(n14712), .Z(n14713) );
  XOR U14953 ( .A(n14714), .B(n14713), .Z(n14644) );
  NANDN U14954 ( .A(n14634), .B(n14633), .Z(n14638) );
  NANDN U14955 ( .A(n14636), .B(n14635), .Z(n14637) );
  NAND U14956 ( .A(n14638), .B(n14637), .Z(n14645) );
  XNOR U14957 ( .A(n14644), .B(n14645), .Z(n14646) );
  XNOR U14958 ( .A(n14647), .B(n14646), .Z(n14717) );
  XNOR U14959 ( .A(n14717), .B(sreg[434]), .Z(n14719) );
  NAND U14960 ( .A(n14639), .B(sreg[433]), .Z(n14643) );
  OR U14961 ( .A(n14641), .B(n14640), .Z(n14642) );
  AND U14962 ( .A(n14643), .B(n14642), .Z(n14718) );
  XOR U14963 ( .A(n14719), .B(n14718), .Z(c[434]) );
  NANDN U14964 ( .A(n14645), .B(n14644), .Z(n14649) );
  NAND U14965 ( .A(n14647), .B(n14646), .Z(n14648) );
  NAND U14966 ( .A(n14649), .B(n14648), .Z(n14725) );
  NANDN U14967 ( .A(n14651), .B(n14650), .Z(n14655) );
  OR U14968 ( .A(n14653), .B(n14652), .Z(n14654) );
  NAND U14969 ( .A(n14655), .B(n14654), .Z(n14792) );
  XNOR U14970 ( .A(n20052), .B(n14971), .Z(n14734) );
  OR U14971 ( .A(n14734), .B(n20020), .Z(n14658) );
  NANDN U14972 ( .A(n14656), .B(n19960), .Z(n14657) );
  NAND U14973 ( .A(n14658), .B(n14657), .Z(n14747) );
  XNOR U14974 ( .A(n102), .B(n14659), .Z(n14738) );
  OR U14975 ( .A(n14738), .B(n20121), .Z(n14662) );
  NANDN U14976 ( .A(n14660), .B(n20122), .Z(n14661) );
  NAND U14977 ( .A(n14662), .B(n14661), .Z(n14744) );
  XNOR U14978 ( .A(n19975), .B(n15127), .Z(n14741) );
  NANDN U14979 ( .A(n14741), .B(n19883), .Z(n14665) );
  NANDN U14980 ( .A(n14663), .B(n19937), .Z(n14664) );
  AND U14981 ( .A(n14665), .B(n14664), .Z(n14745) );
  XNOR U14982 ( .A(n14744), .B(n14745), .Z(n14746) );
  XNOR U14983 ( .A(n14747), .B(n14746), .Z(n14783) );
  NANDN U14984 ( .A(n14667), .B(n14666), .Z(n14671) );
  NAND U14985 ( .A(n14669), .B(n14668), .Z(n14670) );
  NAND U14986 ( .A(n14671), .B(n14670), .Z(n14784) );
  XNOR U14987 ( .A(n14783), .B(n14784), .Z(n14785) );
  NANDN U14988 ( .A(n14673), .B(n14672), .Z(n14677) );
  NAND U14989 ( .A(n14675), .B(n14674), .Z(n14676) );
  AND U14990 ( .A(n14677), .B(n14676), .Z(n14786) );
  XNOR U14991 ( .A(n14785), .B(n14786), .Z(n14730) );
  NANDN U14992 ( .A(n14679), .B(n14678), .Z(n14683) );
  OR U14993 ( .A(n14681), .B(n14680), .Z(n14682) );
  NAND U14994 ( .A(n14683), .B(n14682), .Z(n14780) );
  XNOR U14995 ( .A(n20154), .B(n14815), .Z(n14765) );
  OR U14996 ( .A(n14765), .B(n20057), .Z(n14686) );
  NANDN U14997 ( .A(n14684), .B(n20098), .Z(n14685) );
  AND U14998 ( .A(n14686), .B(n14685), .Z(n14757) );
  NAND U14999 ( .A(b[0]), .B(a[195]), .Z(n14687) );
  XNOR U15000 ( .A(b[1]), .B(n14687), .Z(n14689) );
  NAND U15001 ( .A(a[194]), .B(n98), .Z(n14688) );
  AND U15002 ( .A(n14689), .B(n14688), .Z(n14756) );
  XOR U15003 ( .A(n14757), .B(n14756), .Z(n14759) );
  NAND U15004 ( .A(a[179]), .B(b[15]), .Z(n14758) );
  XOR U15005 ( .A(n14759), .B(n14758), .Z(n14777) );
  NAND U15006 ( .A(n19722), .B(n14690), .Z(n14692) );
  XNOR U15007 ( .A(b[5]), .B(n15436), .Z(n14768) );
  NANDN U15008 ( .A(n19640), .B(n14768), .Z(n14691) );
  NAND U15009 ( .A(n14692), .B(n14691), .Z(n14753) );
  XNOR U15010 ( .A(n19714), .B(n15280), .Z(n14771) );
  NANDN U15011 ( .A(n14771), .B(n19766), .Z(n14695) );
  NANDN U15012 ( .A(n14693), .B(n19767), .Z(n14694) );
  NAND U15013 ( .A(n14695), .B(n14694), .Z(n14750) );
  NAND U15014 ( .A(n19554), .B(n14696), .Z(n14698) );
  IV U15015 ( .A(a[193]), .Z(n15619) );
  XNOR U15016 ( .A(b[3]), .B(n15619), .Z(n14774) );
  NANDN U15017 ( .A(n19521), .B(n14774), .Z(n14697) );
  AND U15018 ( .A(n14698), .B(n14697), .Z(n14751) );
  XNOR U15019 ( .A(n14750), .B(n14751), .Z(n14752) );
  XOR U15020 ( .A(n14753), .B(n14752), .Z(n14778) );
  XOR U15021 ( .A(n14777), .B(n14778), .Z(n14779) );
  XNOR U15022 ( .A(n14780), .B(n14779), .Z(n14728) );
  NAND U15023 ( .A(n14700), .B(n14699), .Z(n14704) );
  NAND U15024 ( .A(n14702), .B(n14701), .Z(n14703) );
  NAND U15025 ( .A(n14704), .B(n14703), .Z(n14729) );
  XOR U15026 ( .A(n14728), .B(n14729), .Z(n14731) );
  XNOR U15027 ( .A(n14730), .B(n14731), .Z(n14789) );
  NANDN U15028 ( .A(n14706), .B(n14705), .Z(n14710) );
  NAND U15029 ( .A(n14708), .B(n14707), .Z(n14709) );
  NAND U15030 ( .A(n14710), .B(n14709), .Z(n14790) );
  XNOR U15031 ( .A(n14789), .B(n14790), .Z(n14791) );
  XOR U15032 ( .A(n14792), .B(n14791), .Z(n14722) );
  NANDN U15033 ( .A(n14712), .B(n14711), .Z(n14716) );
  NANDN U15034 ( .A(n14714), .B(n14713), .Z(n14715) );
  NAND U15035 ( .A(n14716), .B(n14715), .Z(n14723) );
  XNOR U15036 ( .A(n14722), .B(n14723), .Z(n14724) );
  XNOR U15037 ( .A(n14725), .B(n14724), .Z(n14795) );
  XNOR U15038 ( .A(n14795), .B(sreg[435]), .Z(n14797) );
  NAND U15039 ( .A(n14717), .B(sreg[434]), .Z(n14721) );
  OR U15040 ( .A(n14719), .B(n14718), .Z(n14720) );
  AND U15041 ( .A(n14721), .B(n14720), .Z(n14796) );
  XOR U15042 ( .A(n14797), .B(n14796), .Z(c[435]) );
  NANDN U15043 ( .A(n14723), .B(n14722), .Z(n14727) );
  NAND U15044 ( .A(n14725), .B(n14724), .Z(n14726) );
  NAND U15045 ( .A(n14727), .B(n14726), .Z(n14803) );
  NANDN U15046 ( .A(n14729), .B(n14728), .Z(n14733) );
  OR U15047 ( .A(n14731), .B(n14730), .Z(n14732) );
  NAND U15048 ( .A(n14733), .B(n14732), .Z(n14870) );
  XNOR U15049 ( .A(n20052), .B(n15049), .Z(n14812) );
  OR U15050 ( .A(n14812), .B(n20020), .Z(n14736) );
  NANDN U15051 ( .A(n14734), .B(n19960), .Z(n14735) );
  NAND U15052 ( .A(n14736), .B(n14735), .Z(n14825) );
  XNOR U15053 ( .A(n102), .B(n14737), .Z(n14816) );
  OR U15054 ( .A(n14816), .B(n20121), .Z(n14740) );
  NANDN U15055 ( .A(n14738), .B(n20122), .Z(n14739) );
  NAND U15056 ( .A(n14740), .B(n14739), .Z(n14822) );
  XNOR U15057 ( .A(n19975), .B(n15204), .Z(n14819) );
  NANDN U15058 ( .A(n14819), .B(n19883), .Z(n14743) );
  NANDN U15059 ( .A(n14741), .B(n19937), .Z(n14742) );
  AND U15060 ( .A(n14743), .B(n14742), .Z(n14823) );
  XNOR U15061 ( .A(n14822), .B(n14823), .Z(n14824) );
  XNOR U15062 ( .A(n14825), .B(n14824), .Z(n14861) );
  NANDN U15063 ( .A(n14745), .B(n14744), .Z(n14749) );
  NAND U15064 ( .A(n14747), .B(n14746), .Z(n14748) );
  NAND U15065 ( .A(n14749), .B(n14748), .Z(n14862) );
  XNOR U15066 ( .A(n14861), .B(n14862), .Z(n14863) );
  NANDN U15067 ( .A(n14751), .B(n14750), .Z(n14755) );
  NAND U15068 ( .A(n14753), .B(n14752), .Z(n14754) );
  AND U15069 ( .A(n14755), .B(n14754), .Z(n14864) );
  XNOR U15070 ( .A(n14863), .B(n14864), .Z(n14808) );
  NANDN U15071 ( .A(n14757), .B(n14756), .Z(n14761) );
  OR U15072 ( .A(n14759), .B(n14758), .Z(n14760) );
  NAND U15073 ( .A(n14761), .B(n14760), .Z(n14858) );
  NAND U15074 ( .A(b[0]), .B(a[196]), .Z(n14762) );
  XNOR U15075 ( .A(b[1]), .B(n14762), .Z(n14764) );
  NAND U15076 ( .A(a[195]), .B(n98), .Z(n14763) );
  AND U15077 ( .A(n14764), .B(n14763), .Z(n14834) );
  XNOR U15078 ( .A(n20154), .B(n14893), .Z(n14840) );
  OR U15079 ( .A(n14840), .B(n20057), .Z(n14767) );
  NANDN U15080 ( .A(n14765), .B(n20098), .Z(n14766) );
  AND U15081 ( .A(n14767), .B(n14766), .Z(n14835) );
  XOR U15082 ( .A(n14834), .B(n14835), .Z(n14837) );
  NAND U15083 ( .A(a[180]), .B(b[15]), .Z(n14836) );
  XOR U15084 ( .A(n14837), .B(n14836), .Z(n14855) );
  NAND U15085 ( .A(n19722), .B(n14768), .Z(n14770) );
  XNOR U15086 ( .A(b[5]), .B(n15514), .Z(n14846) );
  NANDN U15087 ( .A(n19640), .B(n14846), .Z(n14769) );
  NAND U15088 ( .A(n14770), .B(n14769), .Z(n14831) );
  XNOR U15089 ( .A(n19714), .B(n15385), .Z(n14849) );
  NANDN U15090 ( .A(n14849), .B(n19766), .Z(n14773) );
  NANDN U15091 ( .A(n14771), .B(n19767), .Z(n14772) );
  NAND U15092 ( .A(n14773), .B(n14772), .Z(n14828) );
  NAND U15093 ( .A(n19554), .B(n14774), .Z(n14776) );
  IV U15094 ( .A(a[194]), .Z(n15697) );
  XNOR U15095 ( .A(b[3]), .B(n15697), .Z(n14852) );
  NANDN U15096 ( .A(n19521), .B(n14852), .Z(n14775) );
  AND U15097 ( .A(n14776), .B(n14775), .Z(n14829) );
  XNOR U15098 ( .A(n14828), .B(n14829), .Z(n14830) );
  XOR U15099 ( .A(n14831), .B(n14830), .Z(n14856) );
  XOR U15100 ( .A(n14855), .B(n14856), .Z(n14857) );
  XNOR U15101 ( .A(n14858), .B(n14857), .Z(n14806) );
  NAND U15102 ( .A(n14778), .B(n14777), .Z(n14782) );
  NAND U15103 ( .A(n14780), .B(n14779), .Z(n14781) );
  NAND U15104 ( .A(n14782), .B(n14781), .Z(n14807) );
  XOR U15105 ( .A(n14806), .B(n14807), .Z(n14809) );
  XNOR U15106 ( .A(n14808), .B(n14809), .Z(n14867) );
  NANDN U15107 ( .A(n14784), .B(n14783), .Z(n14788) );
  NAND U15108 ( .A(n14786), .B(n14785), .Z(n14787) );
  NAND U15109 ( .A(n14788), .B(n14787), .Z(n14868) );
  XNOR U15110 ( .A(n14867), .B(n14868), .Z(n14869) );
  XOR U15111 ( .A(n14870), .B(n14869), .Z(n14800) );
  NANDN U15112 ( .A(n14790), .B(n14789), .Z(n14794) );
  NANDN U15113 ( .A(n14792), .B(n14791), .Z(n14793) );
  NAND U15114 ( .A(n14794), .B(n14793), .Z(n14801) );
  XNOR U15115 ( .A(n14800), .B(n14801), .Z(n14802) );
  XNOR U15116 ( .A(n14803), .B(n14802), .Z(n14873) );
  XNOR U15117 ( .A(n14873), .B(sreg[436]), .Z(n14875) );
  NAND U15118 ( .A(n14795), .B(sreg[435]), .Z(n14799) );
  OR U15119 ( .A(n14797), .B(n14796), .Z(n14798) );
  AND U15120 ( .A(n14799), .B(n14798), .Z(n14874) );
  XOR U15121 ( .A(n14875), .B(n14874), .Z(c[436]) );
  NANDN U15122 ( .A(n14801), .B(n14800), .Z(n14805) );
  NAND U15123 ( .A(n14803), .B(n14802), .Z(n14804) );
  NAND U15124 ( .A(n14805), .B(n14804), .Z(n14881) );
  NANDN U15125 ( .A(n14807), .B(n14806), .Z(n14811) );
  OR U15126 ( .A(n14809), .B(n14808), .Z(n14810) );
  NAND U15127 ( .A(n14811), .B(n14810), .Z(n14948) );
  XNOR U15128 ( .A(n20052), .B(n15127), .Z(n14890) );
  OR U15129 ( .A(n14890), .B(n20020), .Z(n14814) );
  NANDN U15130 ( .A(n14812), .B(n19960), .Z(n14813) );
  NAND U15131 ( .A(n14814), .B(n14813), .Z(n14903) );
  XNOR U15132 ( .A(n102), .B(n14815), .Z(n14894) );
  OR U15133 ( .A(n14894), .B(n20121), .Z(n14818) );
  NANDN U15134 ( .A(n14816), .B(n20122), .Z(n14817) );
  NAND U15135 ( .A(n14818), .B(n14817), .Z(n14900) );
  XNOR U15136 ( .A(n19975), .B(n15280), .Z(n14897) );
  NANDN U15137 ( .A(n14897), .B(n19883), .Z(n14821) );
  NANDN U15138 ( .A(n14819), .B(n19937), .Z(n14820) );
  AND U15139 ( .A(n14821), .B(n14820), .Z(n14901) );
  XNOR U15140 ( .A(n14900), .B(n14901), .Z(n14902) );
  XNOR U15141 ( .A(n14903), .B(n14902), .Z(n14939) );
  NANDN U15142 ( .A(n14823), .B(n14822), .Z(n14827) );
  NAND U15143 ( .A(n14825), .B(n14824), .Z(n14826) );
  NAND U15144 ( .A(n14827), .B(n14826), .Z(n14940) );
  XNOR U15145 ( .A(n14939), .B(n14940), .Z(n14941) );
  NANDN U15146 ( .A(n14829), .B(n14828), .Z(n14833) );
  NAND U15147 ( .A(n14831), .B(n14830), .Z(n14832) );
  AND U15148 ( .A(n14833), .B(n14832), .Z(n14942) );
  XNOR U15149 ( .A(n14941), .B(n14942), .Z(n14886) );
  NANDN U15150 ( .A(n14835), .B(n14834), .Z(n14839) );
  OR U15151 ( .A(n14837), .B(n14836), .Z(n14838) );
  NAND U15152 ( .A(n14839), .B(n14838), .Z(n14936) );
  XNOR U15153 ( .A(n20154), .B(n14971), .Z(n14921) );
  OR U15154 ( .A(n14921), .B(n20057), .Z(n14842) );
  NANDN U15155 ( .A(n14840), .B(n20098), .Z(n14841) );
  AND U15156 ( .A(n14842), .B(n14841), .Z(n14913) );
  NAND U15157 ( .A(b[0]), .B(a[197]), .Z(n14843) );
  XNOR U15158 ( .A(b[1]), .B(n14843), .Z(n14845) );
  NAND U15159 ( .A(a[196]), .B(n98), .Z(n14844) );
  AND U15160 ( .A(n14845), .B(n14844), .Z(n14912) );
  XOR U15161 ( .A(n14913), .B(n14912), .Z(n14915) );
  NAND U15162 ( .A(a[181]), .B(b[15]), .Z(n14914) );
  XOR U15163 ( .A(n14915), .B(n14914), .Z(n14933) );
  NAND U15164 ( .A(n19722), .B(n14846), .Z(n14848) );
  XNOR U15165 ( .A(b[5]), .B(n15619), .Z(n14924) );
  NANDN U15166 ( .A(n19640), .B(n14924), .Z(n14847) );
  NAND U15167 ( .A(n14848), .B(n14847), .Z(n14909) );
  XNOR U15168 ( .A(n19714), .B(n15436), .Z(n14927) );
  NANDN U15169 ( .A(n14927), .B(n19766), .Z(n14851) );
  NANDN U15170 ( .A(n14849), .B(n19767), .Z(n14850) );
  NAND U15171 ( .A(n14851), .B(n14850), .Z(n14906) );
  NAND U15172 ( .A(n19554), .B(n14852), .Z(n14854) );
  IV U15173 ( .A(a[195]), .Z(n15775) );
  XNOR U15174 ( .A(b[3]), .B(n15775), .Z(n14930) );
  NANDN U15175 ( .A(n19521), .B(n14930), .Z(n14853) );
  AND U15176 ( .A(n14854), .B(n14853), .Z(n14907) );
  XNOR U15177 ( .A(n14906), .B(n14907), .Z(n14908) );
  XOR U15178 ( .A(n14909), .B(n14908), .Z(n14934) );
  XOR U15179 ( .A(n14933), .B(n14934), .Z(n14935) );
  XNOR U15180 ( .A(n14936), .B(n14935), .Z(n14884) );
  NAND U15181 ( .A(n14856), .B(n14855), .Z(n14860) );
  NAND U15182 ( .A(n14858), .B(n14857), .Z(n14859) );
  NAND U15183 ( .A(n14860), .B(n14859), .Z(n14885) );
  XOR U15184 ( .A(n14884), .B(n14885), .Z(n14887) );
  XNOR U15185 ( .A(n14886), .B(n14887), .Z(n14945) );
  NANDN U15186 ( .A(n14862), .B(n14861), .Z(n14866) );
  NAND U15187 ( .A(n14864), .B(n14863), .Z(n14865) );
  NAND U15188 ( .A(n14866), .B(n14865), .Z(n14946) );
  XNOR U15189 ( .A(n14945), .B(n14946), .Z(n14947) );
  XOR U15190 ( .A(n14948), .B(n14947), .Z(n14878) );
  NANDN U15191 ( .A(n14868), .B(n14867), .Z(n14872) );
  NANDN U15192 ( .A(n14870), .B(n14869), .Z(n14871) );
  NAND U15193 ( .A(n14872), .B(n14871), .Z(n14879) );
  XNOR U15194 ( .A(n14878), .B(n14879), .Z(n14880) );
  XNOR U15195 ( .A(n14881), .B(n14880), .Z(n14951) );
  XNOR U15196 ( .A(n14951), .B(sreg[437]), .Z(n14953) );
  NAND U15197 ( .A(n14873), .B(sreg[436]), .Z(n14877) );
  OR U15198 ( .A(n14875), .B(n14874), .Z(n14876) );
  AND U15199 ( .A(n14877), .B(n14876), .Z(n14952) );
  XOR U15200 ( .A(n14953), .B(n14952), .Z(c[437]) );
  NANDN U15201 ( .A(n14879), .B(n14878), .Z(n14883) );
  NAND U15202 ( .A(n14881), .B(n14880), .Z(n14882) );
  NAND U15203 ( .A(n14883), .B(n14882), .Z(n14959) );
  NANDN U15204 ( .A(n14885), .B(n14884), .Z(n14889) );
  OR U15205 ( .A(n14887), .B(n14886), .Z(n14888) );
  NAND U15206 ( .A(n14889), .B(n14888), .Z(n15026) );
  XNOR U15207 ( .A(n20052), .B(n15204), .Z(n14968) );
  OR U15208 ( .A(n14968), .B(n20020), .Z(n14892) );
  NANDN U15209 ( .A(n14890), .B(n19960), .Z(n14891) );
  NAND U15210 ( .A(n14892), .B(n14891), .Z(n14981) );
  XNOR U15211 ( .A(n102), .B(n14893), .Z(n14972) );
  OR U15212 ( .A(n14972), .B(n20121), .Z(n14896) );
  NANDN U15213 ( .A(n14894), .B(n20122), .Z(n14895) );
  NAND U15214 ( .A(n14896), .B(n14895), .Z(n14978) );
  XNOR U15215 ( .A(n19975), .B(n15385), .Z(n14975) );
  NANDN U15216 ( .A(n14975), .B(n19883), .Z(n14899) );
  NANDN U15217 ( .A(n14897), .B(n19937), .Z(n14898) );
  AND U15218 ( .A(n14899), .B(n14898), .Z(n14979) );
  XNOR U15219 ( .A(n14978), .B(n14979), .Z(n14980) );
  XNOR U15220 ( .A(n14981), .B(n14980), .Z(n15017) );
  NANDN U15221 ( .A(n14901), .B(n14900), .Z(n14905) );
  NAND U15222 ( .A(n14903), .B(n14902), .Z(n14904) );
  NAND U15223 ( .A(n14905), .B(n14904), .Z(n15018) );
  XNOR U15224 ( .A(n15017), .B(n15018), .Z(n15019) );
  NANDN U15225 ( .A(n14907), .B(n14906), .Z(n14911) );
  NAND U15226 ( .A(n14909), .B(n14908), .Z(n14910) );
  AND U15227 ( .A(n14911), .B(n14910), .Z(n15020) );
  XNOR U15228 ( .A(n15019), .B(n15020), .Z(n14964) );
  NANDN U15229 ( .A(n14913), .B(n14912), .Z(n14917) );
  OR U15230 ( .A(n14915), .B(n14914), .Z(n14916) );
  NAND U15231 ( .A(n14917), .B(n14916), .Z(n15014) );
  NAND U15232 ( .A(b[0]), .B(a[198]), .Z(n14918) );
  XNOR U15233 ( .A(b[1]), .B(n14918), .Z(n14920) );
  NAND U15234 ( .A(a[197]), .B(n98), .Z(n14919) );
  AND U15235 ( .A(n14920), .B(n14919), .Z(n14990) );
  XNOR U15236 ( .A(n20154), .B(n15049), .Z(n14999) );
  OR U15237 ( .A(n14999), .B(n20057), .Z(n14923) );
  NANDN U15238 ( .A(n14921), .B(n20098), .Z(n14922) );
  AND U15239 ( .A(n14923), .B(n14922), .Z(n14991) );
  XOR U15240 ( .A(n14990), .B(n14991), .Z(n14993) );
  NAND U15241 ( .A(a[182]), .B(b[15]), .Z(n14992) );
  XOR U15242 ( .A(n14993), .B(n14992), .Z(n15011) );
  NAND U15243 ( .A(n19722), .B(n14924), .Z(n14926) );
  XNOR U15244 ( .A(b[5]), .B(n15697), .Z(n15002) );
  NANDN U15245 ( .A(n19640), .B(n15002), .Z(n14925) );
  NAND U15246 ( .A(n14926), .B(n14925), .Z(n14987) );
  XNOR U15247 ( .A(n19714), .B(n15514), .Z(n15005) );
  NANDN U15248 ( .A(n15005), .B(n19766), .Z(n14929) );
  NANDN U15249 ( .A(n14927), .B(n19767), .Z(n14928) );
  NAND U15250 ( .A(n14929), .B(n14928), .Z(n14984) );
  NAND U15251 ( .A(n19554), .B(n14930), .Z(n14932) );
  IV U15252 ( .A(a[196]), .Z(n15826) );
  XNOR U15253 ( .A(b[3]), .B(n15826), .Z(n15008) );
  NANDN U15254 ( .A(n19521), .B(n15008), .Z(n14931) );
  AND U15255 ( .A(n14932), .B(n14931), .Z(n14985) );
  XNOR U15256 ( .A(n14984), .B(n14985), .Z(n14986) );
  XOR U15257 ( .A(n14987), .B(n14986), .Z(n15012) );
  XOR U15258 ( .A(n15011), .B(n15012), .Z(n15013) );
  XNOR U15259 ( .A(n15014), .B(n15013), .Z(n14962) );
  NAND U15260 ( .A(n14934), .B(n14933), .Z(n14938) );
  NAND U15261 ( .A(n14936), .B(n14935), .Z(n14937) );
  NAND U15262 ( .A(n14938), .B(n14937), .Z(n14963) );
  XOR U15263 ( .A(n14962), .B(n14963), .Z(n14965) );
  XNOR U15264 ( .A(n14964), .B(n14965), .Z(n15023) );
  NANDN U15265 ( .A(n14940), .B(n14939), .Z(n14944) );
  NAND U15266 ( .A(n14942), .B(n14941), .Z(n14943) );
  NAND U15267 ( .A(n14944), .B(n14943), .Z(n15024) );
  XNOR U15268 ( .A(n15023), .B(n15024), .Z(n15025) );
  XOR U15269 ( .A(n15026), .B(n15025), .Z(n14956) );
  NANDN U15270 ( .A(n14946), .B(n14945), .Z(n14950) );
  NANDN U15271 ( .A(n14948), .B(n14947), .Z(n14949) );
  NAND U15272 ( .A(n14950), .B(n14949), .Z(n14957) );
  XNOR U15273 ( .A(n14956), .B(n14957), .Z(n14958) );
  XNOR U15274 ( .A(n14959), .B(n14958), .Z(n15029) );
  XNOR U15275 ( .A(n15029), .B(sreg[438]), .Z(n15031) );
  NAND U15276 ( .A(n14951), .B(sreg[437]), .Z(n14955) );
  OR U15277 ( .A(n14953), .B(n14952), .Z(n14954) );
  AND U15278 ( .A(n14955), .B(n14954), .Z(n15030) );
  XOR U15279 ( .A(n15031), .B(n15030), .Z(c[438]) );
  NANDN U15280 ( .A(n14957), .B(n14956), .Z(n14961) );
  NAND U15281 ( .A(n14959), .B(n14958), .Z(n14960) );
  NAND U15282 ( .A(n14961), .B(n14960), .Z(n15037) );
  NANDN U15283 ( .A(n14963), .B(n14962), .Z(n14967) );
  OR U15284 ( .A(n14965), .B(n14964), .Z(n14966) );
  NAND U15285 ( .A(n14967), .B(n14966), .Z(n15104) );
  XNOR U15286 ( .A(n20052), .B(n15280), .Z(n15046) );
  OR U15287 ( .A(n15046), .B(n20020), .Z(n14970) );
  NANDN U15288 ( .A(n14968), .B(n19960), .Z(n14969) );
  NAND U15289 ( .A(n14970), .B(n14969), .Z(n15059) );
  XNOR U15290 ( .A(n102), .B(n14971), .Z(n15050) );
  OR U15291 ( .A(n15050), .B(n20121), .Z(n14974) );
  NANDN U15292 ( .A(n14972), .B(n20122), .Z(n14973) );
  NAND U15293 ( .A(n14974), .B(n14973), .Z(n15056) );
  XNOR U15294 ( .A(n19975), .B(n15436), .Z(n15053) );
  NANDN U15295 ( .A(n15053), .B(n19883), .Z(n14977) );
  NANDN U15296 ( .A(n14975), .B(n19937), .Z(n14976) );
  AND U15297 ( .A(n14977), .B(n14976), .Z(n15057) );
  XNOR U15298 ( .A(n15056), .B(n15057), .Z(n15058) );
  XNOR U15299 ( .A(n15059), .B(n15058), .Z(n15095) );
  NANDN U15300 ( .A(n14979), .B(n14978), .Z(n14983) );
  NAND U15301 ( .A(n14981), .B(n14980), .Z(n14982) );
  NAND U15302 ( .A(n14983), .B(n14982), .Z(n15096) );
  XNOR U15303 ( .A(n15095), .B(n15096), .Z(n15097) );
  NANDN U15304 ( .A(n14985), .B(n14984), .Z(n14989) );
  NAND U15305 ( .A(n14987), .B(n14986), .Z(n14988) );
  AND U15306 ( .A(n14989), .B(n14988), .Z(n15098) );
  XNOR U15307 ( .A(n15097), .B(n15098), .Z(n15042) );
  NANDN U15308 ( .A(n14991), .B(n14990), .Z(n14995) );
  OR U15309 ( .A(n14993), .B(n14992), .Z(n14994) );
  NAND U15310 ( .A(n14995), .B(n14994), .Z(n15092) );
  NAND U15311 ( .A(b[0]), .B(a[199]), .Z(n14996) );
  XNOR U15312 ( .A(b[1]), .B(n14996), .Z(n14998) );
  NAND U15313 ( .A(a[198]), .B(n98), .Z(n14997) );
  AND U15314 ( .A(n14998), .B(n14997), .Z(n15068) );
  XNOR U15315 ( .A(n20154), .B(n15127), .Z(n15074) );
  OR U15316 ( .A(n15074), .B(n20057), .Z(n15001) );
  NANDN U15317 ( .A(n14999), .B(n20098), .Z(n15000) );
  AND U15318 ( .A(n15001), .B(n15000), .Z(n15069) );
  XOR U15319 ( .A(n15068), .B(n15069), .Z(n15071) );
  NAND U15320 ( .A(a[183]), .B(b[15]), .Z(n15070) );
  XOR U15321 ( .A(n15071), .B(n15070), .Z(n15089) );
  NAND U15322 ( .A(n19722), .B(n15002), .Z(n15004) );
  XNOR U15323 ( .A(b[5]), .B(n15775), .Z(n15080) );
  NANDN U15324 ( .A(n19640), .B(n15080), .Z(n15003) );
  NAND U15325 ( .A(n15004), .B(n15003), .Z(n15065) );
  XNOR U15326 ( .A(n19714), .B(n15619), .Z(n15083) );
  NANDN U15327 ( .A(n15083), .B(n19766), .Z(n15007) );
  NANDN U15328 ( .A(n15005), .B(n19767), .Z(n15006) );
  NAND U15329 ( .A(n15007), .B(n15006), .Z(n15062) );
  NAND U15330 ( .A(n19554), .B(n15008), .Z(n15010) );
  IV U15331 ( .A(a[197]), .Z(n15931) );
  XNOR U15332 ( .A(b[3]), .B(n15931), .Z(n15086) );
  NANDN U15333 ( .A(n19521), .B(n15086), .Z(n15009) );
  AND U15334 ( .A(n15010), .B(n15009), .Z(n15063) );
  XNOR U15335 ( .A(n15062), .B(n15063), .Z(n15064) );
  XOR U15336 ( .A(n15065), .B(n15064), .Z(n15090) );
  XOR U15337 ( .A(n15089), .B(n15090), .Z(n15091) );
  XNOR U15338 ( .A(n15092), .B(n15091), .Z(n15040) );
  NAND U15339 ( .A(n15012), .B(n15011), .Z(n15016) );
  NAND U15340 ( .A(n15014), .B(n15013), .Z(n15015) );
  NAND U15341 ( .A(n15016), .B(n15015), .Z(n15041) );
  XOR U15342 ( .A(n15040), .B(n15041), .Z(n15043) );
  XNOR U15343 ( .A(n15042), .B(n15043), .Z(n15101) );
  NANDN U15344 ( .A(n15018), .B(n15017), .Z(n15022) );
  NAND U15345 ( .A(n15020), .B(n15019), .Z(n15021) );
  NAND U15346 ( .A(n15022), .B(n15021), .Z(n15102) );
  XNOR U15347 ( .A(n15101), .B(n15102), .Z(n15103) );
  XOR U15348 ( .A(n15104), .B(n15103), .Z(n15034) );
  NANDN U15349 ( .A(n15024), .B(n15023), .Z(n15028) );
  NANDN U15350 ( .A(n15026), .B(n15025), .Z(n15027) );
  NAND U15351 ( .A(n15028), .B(n15027), .Z(n15035) );
  XNOR U15352 ( .A(n15034), .B(n15035), .Z(n15036) );
  XNOR U15353 ( .A(n15037), .B(n15036), .Z(n15107) );
  XNOR U15354 ( .A(n15107), .B(sreg[439]), .Z(n15109) );
  NAND U15355 ( .A(n15029), .B(sreg[438]), .Z(n15033) );
  OR U15356 ( .A(n15031), .B(n15030), .Z(n15032) );
  AND U15357 ( .A(n15033), .B(n15032), .Z(n15108) );
  XOR U15358 ( .A(n15109), .B(n15108), .Z(c[439]) );
  NANDN U15359 ( .A(n15035), .B(n15034), .Z(n15039) );
  NAND U15360 ( .A(n15037), .B(n15036), .Z(n15038) );
  NAND U15361 ( .A(n15039), .B(n15038), .Z(n15115) );
  NANDN U15362 ( .A(n15041), .B(n15040), .Z(n15045) );
  OR U15363 ( .A(n15043), .B(n15042), .Z(n15044) );
  NAND U15364 ( .A(n15045), .B(n15044), .Z(n15181) );
  XNOR U15365 ( .A(n20052), .B(n15385), .Z(n15124) );
  OR U15366 ( .A(n15124), .B(n20020), .Z(n15048) );
  NANDN U15367 ( .A(n15046), .B(n19960), .Z(n15047) );
  NAND U15368 ( .A(n15048), .B(n15047), .Z(n15137) );
  XNOR U15369 ( .A(n102), .B(n15049), .Z(n15128) );
  OR U15370 ( .A(n15128), .B(n20121), .Z(n15052) );
  NANDN U15371 ( .A(n15050), .B(n20122), .Z(n15051) );
  NAND U15372 ( .A(n15052), .B(n15051), .Z(n15134) );
  XNOR U15373 ( .A(n19975), .B(n15514), .Z(n15131) );
  NANDN U15374 ( .A(n15131), .B(n19883), .Z(n15055) );
  NANDN U15375 ( .A(n15053), .B(n19937), .Z(n15054) );
  AND U15376 ( .A(n15055), .B(n15054), .Z(n15135) );
  XNOR U15377 ( .A(n15134), .B(n15135), .Z(n15136) );
  XNOR U15378 ( .A(n15137), .B(n15136), .Z(n15172) );
  NANDN U15379 ( .A(n15057), .B(n15056), .Z(n15061) );
  NAND U15380 ( .A(n15059), .B(n15058), .Z(n15060) );
  NAND U15381 ( .A(n15061), .B(n15060), .Z(n15173) );
  XNOR U15382 ( .A(n15172), .B(n15173), .Z(n15174) );
  NANDN U15383 ( .A(n15063), .B(n15062), .Z(n15067) );
  NAND U15384 ( .A(n15065), .B(n15064), .Z(n15066) );
  AND U15385 ( .A(n15067), .B(n15066), .Z(n15175) );
  XNOR U15386 ( .A(n15174), .B(n15175), .Z(n15120) );
  NANDN U15387 ( .A(n15069), .B(n15068), .Z(n15073) );
  OR U15388 ( .A(n15071), .B(n15070), .Z(n15072) );
  NAND U15389 ( .A(n15073), .B(n15072), .Z(n15171) );
  XNOR U15390 ( .A(n20154), .B(n15204), .Z(n15152) );
  OR U15391 ( .A(n15152), .B(n20057), .Z(n15076) );
  NANDN U15392 ( .A(n15074), .B(n20098), .Z(n15075) );
  NAND U15393 ( .A(n15076), .B(n15075), .Z(n15146) );
  AND U15394 ( .A(a[200]), .B(b[0]), .Z(n15077) );
  XOR U15395 ( .A(b[1]), .B(n15077), .Z(n15079) );
  NAND U15396 ( .A(a[199]), .B(n98), .Z(n15078) );
  NAND U15397 ( .A(n15079), .B(n15078), .Z(n15147) );
  XNOR U15398 ( .A(n15146), .B(n15147), .Z(n15148) );
  NAND U15399 ( .A(a[184]), .B(b[15]), .Z(n15149) );
  XOR U15400 ( .A(n15148), .B(n15149), .Z(n15168) );
  NAND U15401 ( .A(n19722), .B(n15080), .Z(n15082) );
  XNOR U15402 ( .A(b[5]), .B(n15826), .Z(n15159) );
  NANDN U15403 ( .A(n19640), .B(n15159), .Z(n15081) );
  NAND U15404 ( .A(n15082), .B(n15081), .Z(n15143) );
  XNOR U15405 ( .A(n19714), .B(n15697), .Z(n15162) );
  NANDN U15406 ( .A(n15162), .B(n19766), .Z(n15085) );
  NANDN U15407 ( .A(n15083), .B(n19767), .Z(n15084) );
  NAND U15408 ( .A(n15085), .B(n15084), .Z(n15140) );
  NAND U15409 ( .A(n19554), .B(n15086), .Z(n15088) );
  IV U15410 ( .A(a[198]), .Z(n16009) );
  XNOR U15411 ( .A(b[3]), .B(n16009), .Z(n15165) );
  NANDN U15412 ( .A(n19521), .B(n15165), .Z(n15087) );
  AND U15413 ( .A(n15088), .B(n15087), .Z(n15141) );
  XNOR U15414 ( .A(n15140), .B(n15141), .Z(n15142) );
  XOR U15415 ( .A(n15143), .B(n15142), .Z(n15169) );
  XNOR U15416 ( .A(n15168), .B(n15169), .Z(n15170) );
  XNOR U15417 ( .A(n15171), .B(n15170), .Z(n15118) );
  NAND U15418 ( .A(n15090), .B(n15089), .Z(n15094) );
  NAND U15419 ( .A(n15092), .B(n15091), .Z(n15093) );
  NAND U15420 ( .A(n15094), .B(n15093), .Z(n15119) );
  XOR U15421 ( .A(n15118), .B(n15119), .Z(n15121) );
  XNOR U15422 ( .A(n15120), .B(n15121), .Z(n15178) );
  NANDN U15423 ( .A(n15096), .B(n15095), .Z(n15100) );
  NAND U15424 ( .A(n15098), .B(n15097), .Z(n15099) );
  NAND U15425 ( .A(n15100), .B(n15099), .Z(n15179) );
  XNOR U15426 ( .A(n15178), .B(n15179), .Z(n15180) );
  XOR U15427 ( .A(n15181), .B(n15180), .Z(n15112) );
  NANDN U15428 ( .A(n15102), .B(n15101), .Z(n15106) );
  NANDN U15429 ( .A(n15104), .B(n15103), .Z(n15105) );
  NAND U15430 ( .A(n15106), .B(n15105), .Z(n15113) );
  XNOR U15431 ( .A(n15112), .B(n15113), .Z(n15114) );
  XNOR U15432 ( .A(n15115), .B(n15114), .Z(n15184) );
  XNOR U15433 ( .A(n15184), .B(sreg[440]), .Z(n15186) );
  NAND U15434 ( .A(n15107), .B(sreg[439]), .Z(n15111) );
  OR U15435 ( .A(n15109), .B(n15108), .Z(n15110) );
  AND U15436 ( .A(n15111), .B(n15110), .Z(n15185) );
  XOR U15437 ( .A(n15186), .B(n15185), .Z(c[440]) );
  NANDN U15438 ( .A(n15113), .B(n15112), .Z(n15117) );
  NAND U15439 ( .A(n15115), .B(n15114), .Z(n15116) );
  NAND U15440 ( .A(n15117), .B(n15116), .Z(n15192) );
  NANDN U15441 ( .A(n15119), .B(n15118), .Z(n15123) );
  OR U15442 ( .A(n15121), .B(n15120), .Z(n15122) );
  NAND U15443 ( .A(n15123), .B(n15122), .Z(n15257) );
  XNOR U15444 ( .A(n20052), .B(n15436), .Z(n15201) );
  OR U15445 ( .A(n15201), .B(n20020), .Z(n15126) );
  NANDN U15446 ( .A(n15124), .B(n19960), .Z(n15125) );
  NAND U15447 ( .A(n15126), .B(n15125), .Z(n15214) );
  XNOR U15448 ( .A(n102), .B(n15127), .Z(n15205) );
  OR U15449 ( .A(n15205), .B(n20121), .Z(n15130) );
  NANDN U15450 ( .A(n15128), .B(n20122), .Z(n15129) );
  NAND U15451 ( .A(n15130), .B(n15129), .Z(n15211) );
  XNOR U15452 ( .A(n19975), .B(n15619), .Z(n15208) );
  NANDN U15453 ( .A(n15208), .B(n19883), .Z(n15133) );
  NANDN U15454 ( .A(n15131), .B(n19937), .Z(n15132) );
  AND U15455 ( .A(n15133), .B(n15132), .Z(n15212) );
  XNOR U15456 ( .A(n15211), .B(n15212), .Z(n15213) );
  XNOR U15457 ( .A(n15214), .B(n15213), .Z(n15248) );
  NANDN U15458 ( .A(n15135), .B(n15134), .Z(n15139) );
  NAND U15459 ( .A(n15137), .B(n15136), .Z(n15138) );
  NAND U15460 ( .A(n15139), .B(n15138), .Z(n15249) );
  XNOR U15461 ( .A(n15248), .B(n15249), .Z(n15250) );
  NANDN U15462 ( .A(n15141), .B(n15140), .Z(n15145) );
  NAND U15463 ( .A(n15143), .B(n15142), .Z(n15144) );
  AND U15464 ( .A(n15145), .B(n15144), .Z(n15251) );
  XNOR U15465 ( .A(n15250), .B(n15251), .Z(n15197) );
  NANDN U15466 ( .A(n15147), .B(n15146), .Z(n15151) );
  NANDN U15467 ( .A(n15149), .B(n15148), .Z(n15150) );
  NAND U15468 ( .A(n15151), .B(n15150), .Z(n15247) );
  XNOR U15469 ( .A(n20154), .B(n15280), .Z(n15232) );
  OR U15470 ( .A(n15232), .B(n20057), .Z(n15154) );
  NANDN U15471 ( .A(n15152), .B(n20098), .Z(n15153) );
  NAND U15472 ( .A(n15154), .B(n15153), .Z(n15223) );
  AND U15473 ( .A(a[201]), .B(b[0]), .Z(n15155) );
  XOR U15474 ( .A(b[1]), .B(n15155), .Z(n15158) );
  NANDN U15475 ( .A(n15156), .B(a[200]), .Z(n15157) );
  NAND U15476 ( .A(n15158), .B(n15157), .Z(n15224) );
  XNOR U15477 ( .A(n15223), .B(n15224), .Z(n15225) );
  NAND U15478 ( .A(a[185]), .B(b[15]), .Z(n15226) );
  XOR U15479 ( .A(n15225), .B(n15226), .Z(n15244) );
  NAND U15480 ( .A(n19722), .B(n15159), .Z(n15161) );
  XNOR U15481 ( .A(b[5]), .B(n15931), .Z(n15235) );
  NANDN U15482 ( .A(n19640), .B(n15235), .Z(n15160) );
  NAND U15483 ( .A(n15161), .B(n15160), .Z(n15220) );
  XNOR U15484 ( .A(n19714), .B(n15775), .Z(n15238) );
  NANDN U15485 ( .A(n15238), .B(n19766), .Z(n15164) );
  NANDN U15486 ( .A(n15162), .B(n19767), .Z(n15163) );
  NAND U15487 ( .A(n15164), .B(n15163), .Z(n15217) );
  NAND U15488 ( .A(n19554), .B(n15165), .Z(n15167) );
  IV U15489 ( .A(a[199]), .Z(n16060) );
  XNOR U15490 ( .A(b[3]), .B(n16060), .Z(n15241) );
  NANDN U15491 ( .A(n19521), .B(n15241), .Z(n15166) );
  AND U15492 ( .A(n15167), .B(n15166), .Z(n15218) );
  XNOR U15493 ( .A(n15217), .B(n15218), .Z(n15219) );
  XOR U15494 ( .A(n15220), .B(n15219), .Z(n15245) );
  XNOR U15495 ( .A(n15244), .B(n15245), .Z(n15246) );
  XNOR U15496 ( .A(n15247), .B(n15246), .Z(n15195) );
  XOR U15497 ( .A(n15195), .B(n15196), .Z(n15198) );
  XNOR U15498 ( .A(n15197), .B(n15198), .Z(n15254) );
  NANDN U15499 ( .A(n15173), .B(n15172), .Z(n15177) );
  NAND U15500 ( .A(n15175), .B(n15174), .Z(n15176) );
  NAND U15501 ( .A(n15177), .B(n15176), .Z(n15255) );
  XNOR U15502 ( .A(n15254), .B(n15255), .Z(n15256) );
  XOR U15503 ( .A(n15257), .B(n15256), .Z(n15189) );
  NANDN U15504 ( .A(n15179), .B(n15178), .Z(n15183) );
  NANDN U15505 ( .A(n15181), .B(n15180), .Z(n15182) );
  NAND U15506 ( .A(n15183), .B(n15182), .Z(n15190) );
  XNOR U15507 ( .A(n15189), .B(n15190), .Z(n15191) );
  XNOR U15508 ( .A(n15192), .B(n15191), .Z(n15260) );
  XNOR U15509 ( .A(n15260), .B(sreg[441]), .Z(n15262) );
  NAND U15510 ( .A(n15184), .B(sreg[440]), .Z(n15188) );
  OR U15511 ( .A(n15186), .B(n15185), .Z(n15187) );
  AND U15512 ( .A(n15188), .B(n15187), .Z(n15261) );
  XOR U15513 ( .A(n15262), .B(n15261), .Z(c[441]) );
  NANDN U15514 ( .A(n15190), .B(n15189), .Z(n15194) );
  NAND U15515 ( .A(n15192), .B(n15191), .Z(n15193) );
  NAND U15516 ( .A(n15194), .B(n15193), .Z(n15268) );
  NANDN U15517 ( .A(n15196), .B(n15195), .Z(n15200) );
  OR U15518 ( .A(n15198), .B(n15197), .Z(n15199) );
  NAND U15519 ( .A(n15200), .B(n15199), .Z(n15335) );
  XNOR U15520 ( .A(n20052), .B(n15514), .Z(n15277) );
  OR U15521 ( .A(n15277), .B(n20020), .Z(n15203) );
  NANDN U15522 ( .A(n15201), .B(n19960), .Z(n15202) );
  NAND U15523 ( .A(n15203), .B(n15202), .Z(n15290) );
  XNOR U15524 ( .A(n102), .B(n15204), .Z(n15281) );
  OR U15525 ( .A(n15281), .B(n20121), .Z(n15207) );
  NANDN U15526 ( .A(n15205), .B(n20122), .Z(n15206) );
  NAND U15527 ( .A(n15207), .B(n15206), .Z(n15287) );
  XNOR U15528 ( .A(n19975), .B(n15697), .Z(n15284) );
  NANDN U15529 ( .A(n15284), .B(n19883), .Z(n15210) );
  NANDN U15530 ( .A(n15208), .B(n19937), .Z(n15209) );
  AND U15531 ( .A(n15210), .B(n15209), .Z(n15288) );
  XNOR U15532 ( .A(n15287), .B(n15288), .Z(n15289) );
  XNOR U15533 ( .A(n15290), .B(n15289), .Z(n15326) );
  NANDN U15534 ( .A(n15212), .B(n15211), .Z(n15216) );
  NAND U15535 ( .A(n15214), .B(n15213), .Z(n15215) );
  NAND U15536 ( .A(n15216), .B(n15215), .Z(n15327) );
  XNOR U15537 ( .A(n15326), .B(n15327), .Z(n15328) );
  NANDN U15538 ( .A(n15218), .B(n15217), .Z(n15222) );
  NAND U15539 ( .A(n15220), .B(n15219), .Z(n15221) );
  AND U15540 ( .A(n15222), .B(n15221), .Z(n15329) );
  XNOR U15541 ( .A(n15328), .B(n15329), .Z(n15273) );
  NANDN U15542 ( .A(n15224), .B(n15223), .Z(n15228) );
  NANDN U15543 ( .A(n15226), .B(n15225), .Z(n15227) );
  NAND U15544 ( .A(n15228), .B(n15227), .Z(n15323) );
  NAND U15545 ( .A(b[0]), .B(a[202]), .Z(n15229) );
  XNOR U15546 ( .A(b[1]), .B(n15229), .Z(n15231) );
  NAND U15547 ( .A(a[201]), .B(n98), .Z(n15230) );
  AND U15548 ( .A(n15231), .B(n15230), .Z(n15299) );
  XNOR U15549 ( .A(n20154), .B(n15385), .Z(n15308) );
  OR U15550 ( .A(n15308), .B(n20057), .Z(n15234) );
  NANDN U15551 ( .A(n15232), .B(n20098), .Z(n15233) );
  AND U15552 ( .A(n15234), .B(n15233), .Z(n15300) );
  XOR U15553 ( .A(n15299), .B(n15300), .Z(n15302) );
  NAND U15554 ( .A(a[186]), .B(b[15]), .Z(n15301) );
  XOR U15555 ( .A(n15302), .B(n15301), .Z(n15320) );
  NAND U15556 ( .A(n19722), .B(n15235), .Z(n15237) );
  XNOR U15557 ( .A(b[5]), .B(n16009), .Z(n15311) );
  NANDN U15558 ( .A(n19640), .B(n15311), .Z(n15236) );
  NAND U15559 ( .A(n15237), .B(n15236), .Z(n15296) );
  XNOR U15560 ( .A(n19714), .B(n15826), .Z(n15314) );
  NANDN U15561 ( .A(n15314), .B(n19766), .Z(n15240) );
  NANDN U15562 ( .A(n15238), .B(n19767), .Z(n15239) );
  NAND U15563 ( .A(n15240), .B(n15239), .Z(n15293) );
  NAND U15564 ( .A(n19554), .B(n15241), .Z(n15243) );
  IV U15565 ( .A(a[200]), .Z(n16165) );
  XNOR U15566 ( .A(b[3]), .B(n16165), .Z(n15317) );
  NANDN U15567 ( .A(n19521), .B(n15317), .Z(n15242) );
  AND U15568 ( .A(n15243), .B(n15242), .Z(n15294) );
  XNOR U15569 ( .A(n15293), .B(n15294), .Z(n15295) );
  XOR U15570 ( .A(n15296), .B(n15295), .Z(n15321) );
  XOR U15571 ( .A(n15320), .B(n15321), .Z(n15322) );
  XNOR U15572 ( .A(n15323), .B(n15322), .Z(n15271) );
  XOR U15573 ( .A(n15271), .B(n15272), .Z(n15274) );
  XNOR U15574 ( .A(n15273), .B(n15274), .Z(n15332) );
  NANDN U15575 ( .A(n15249), .B(n15248), .Z(n15253) );
  NAND U15576 ( .A(n15251), .B(n15250), .Z(n15252) );
  NAND U15577 ( .A(n15253), .B(n15252), .Z(n15333) );
  XNOR U15578 ( .A(n15332), .B(n15333), .Z(n15334) );
  XOR U15579 ( .A(n15335), .B(n15334), .Z(n15265) );
  NANDN U15580 ( .A(n15255), .B(n15254), .Z(n15259) );
  NANDN U15581 ( .A(n15257), .B(n15256), .Z(n15258) );
  NAND U15582 ( .A(n15259), .B(n15258), .Z(n15266) );
  XNOR U15583 ( .A(n15265), .B(n15266), .Z(n15267) );
  XNOR U15584 ( .A(n15268), .B(n15267), .Z(n15338) );
  XNOR U15585 ( .A(n15338), .B(sreg[442]), .Z(n15340) );
  NAND U15586 ( .A(n15260), .B(sreg[441]), .Z(n15264) );
  OR U15587 ( .A(n15262), .B(n15261), .Z(n15263) );
  AND U15588 ( .A(n15264), .B(n15263), .Z(n15339) );
  XOR U15589 ( .A(n15340), .B(n15339), .Z(c[442]) );
  NANDN U15590 ( .A(n15266), .B(n15265), .Z(n15270) );
  NAND U15591 ( .A(n15268), .B(n15267), .Z(n15269) );
  NAND U15592 ( .A(n15270), .B(n15269), .Z(n15346) );
  NANDN U15593 ( .A(n15272), .B(n15271), .Z(n15276) );
  OR U15594 ( .A(n15274), .B(n15273), .Z(n15275) );
  NAND U15595 ( .A(n15276), .B(n15275), .Z(n15413) );
  XNOR U15596 ( .A(n20052), .B(n15619), .Z(n15382) );
  OR U15597 ( .A(n15382), .B(n20020), .Z(n15279) );
  NANDN U15598 ( .A(n15277), .B(n19960), .Z(n15278) );
  NAND U15599 ( .A(n15279), .B(n15278), .Z(n15395) );
  XNOR U15600 ( .A(n102), .B(n15280), .Z(n15386) );
  OR U15601 ( .A(n15386), .B(n20121), .Z(n15283) );
  NANDN U15602 ( .A(n15281), .B(n20122), .Z(n15282) );
  NAND U15603 ( .A(n15283), .B(n15282), .Z(n15392) );
  XNOR U15604 ( .A(n19975), .B(n15775), .Z(n15389) );
  NANDN U15605 ( .A(n15389), .B(n19883), .Z(n15286) );
  NANDN U15606 ( .A(n15284), .B(n19937), .Z(n15285) );
  AND U15607 ( .A(n15286), .B(n15285), .Z(n15393) );
  XNOR U15608 ( .A(n15392), .B(n15393), .Z(n15394) );
  XNOR U15609 ( .A(n15395), .B(n15394), .Z(n15404) );
  NANDN U15610 ( .A(n15288), .B(n15287), .Z(n15292) );
  NAND U15611 ( .A(n15290), .B(n15289), .Z(n15291) );
  NAND U15612 ( .A(n15292), .B(n15291), .Z(n15405) );
  XNOR U15613 ( .A(n15404), .B(n15405), .Z(n15406) );
  NANDN U15614 ( .A(n15294), .B(n15293), .Z(n15298) );
  NAND U15615 ( .A(n15296), .B(n15295), .Z(n15297) );
  AND U15616 ( .A(n15298), .B(n15297), .Z(n15407) );
  XNOR U15617 ( .A(n15406), .B(n15407), .Z(n15351) );
  NANDN U15618 ( .A(n15300), .B(n15299), .Z(n15304) );
  OR U15619 ( .A(n15302), .B(n15301), .Z(n15303) );
  NAND U15620 ( .A(n15304), .B(n15303), .Z(n15379) );
  NAND U15621 ( .A(b[0]), .B(a[203]), .Z(n15305) );
  XNOR U15622 ( .A(b[1]), .B(n15305), .Z(n15307) );
  NAND U15623 ( .A(a[202]), .B(n98), .Z(n15306) );
  AND U15624 ( .A(n15307), .B(n15306), .Z(n15355) );
  XNOR U15625 ( .A(n20154), .B(n15436), .Z(n15364) );
  OR U15626 ( .A(n15364), .B(n20057), .Z(n15310) );
  NANDN U15627 ( .A(n15308), .B(n20098), .Z(n15309) );
  AND U15628 ( .A(n15310), .B(n15309), .Z(n15356) );
  XOR U15629 ( .A(n15355), .B(n15356), .Z(n15358) );
  NAND U15630 ( .A(a[187]), .B(b[15]), .Z(n15357) );
  XOR U15631 ( .A(n15358), .B(n15357), .Z(n15376) );
  NAND U15632 ( .A(n19722), .B(n15311), .Z(n15313) );
  XNOR U15633 ( .A(b[5]), .B(n16060), .Z(n15367) );
  NANDN U15634 ( .A(n19640), .B(n15367), .Z(n15312) );
  NAND U15635 ( .A(n15313), .B(n15312), .Z(n15401) );
  XNOR U15636 ( .A(n19714), .B(n15931), .Z(n15370) );
  NANDN U15637 ( .A(n15370), .B(n19766), .Z(n15316) );
  NANDN U15638 ( .A(n15314), .B(n19767), .Z(n15315) );
  NAND U15639 ( .A(n15316), .B(n15315), .Z(n15398) );
  NAND U15640 ( .A(n19554), .B(n15317), .Z(n15319) );
  IV U15641 ( .A(a[201]), .Z(n16216) );
  XNOR U15642 ( .A(b[3]), .B(n16216), .Z(n15373) );
  NANDN U15643 ( .A(n19521), .B(n15373), .Z(n15318) );
  AND U15644 ( .A(n15319), .B(n15318), .Z(n15399) );
  XNOR U15645 ( .A(n15398), .B(n15399), .Z(n15400) );
  XOR U15646 ( .A(n15401), .B(n15400), .Z(n15377) );
  XOR U15647 ( .A(n15376), .B(n15377), .Z(n15378) );
  XNOR U15648 ( .A(n15379), .B(n15378), .Z(n15349) );
  NAND U15649 ( .A(n15321), .B(n15320), .Z(n15325) );
  NAND U15650 ( .A(n15323), .B(n15322), .Z(n15324) );
  NAND U15651 ( .A(n15325), .B(n15324), .Z(n15350) );
  XOR U15652 ( .A(n15349), .B(n15350), .Z(n15352) );
  XNOR U15653 ( .A(n15351), .B(n15352), .Z(n15410) );
  NANDN U15654 ( .A(n15327), .B(n15326), .Z(n15331) );
  NAND U15655 ( .A(n15329), .B(n15328), .Z(n15330) );
  NAND U15656 ( .A(n15331), .B(n15330), .Z(n15411) );
  XNOR U15657 ( .A(n15410), .B(n15411), .Z(n15412) );
  XOR U15658 ( .A(n15413), .B(n15412), .Z(n15343) );
  NANDN U15659 ( .A(n15333), .B(n15332), .Z(n15337) );
  NANDN U15660 ( .A(n15335), .B(n15334), .Z(n15336) );
  NAND U15661 ( .A(n15337), .B(n15336), .Z(n15344) );
  XNOR U15662 ( .A(n15343), .B(n15344), .Z(n15345) );
  XNOR U15663 ( .A(n15346), .B(n15345), .Z(n15416) );
  XNOR U15664 ( .A(n15416), .B(sreg[443]), .Z(n15418) );
  NAND U15665 ( .A(n15338), .B(sreg[442]), .Z(n15342) );
  OR U15666 ( .A(n15340), .B(n15339), .Z(n15341) );
  AND U15667 ( .A(n15342), .B(n15341), .Z(n15417) );
  XOR U15668 ( .A(n15418), .B(n15417), .Z(c[443]) );
  NANDN U15669 ( .A(n15344), .B(n15343), .Z(n15348) );
  NAND U15670 ( .A(n15346), .B(n15345), .Z(n15347) );
  NAND U15671 ( .A(n15348), .B(n15347), .Z(n15424) );
  NANDN U15672 ( .A(n15350), .B(n15349), .Z(n15354) );
  OR U15673 ( .A(n15352), .B(n15351), .Z(n15353) );
  NAND U15674 ( .A(n15354), .B(n15353), .Z(n15491) );
  NANDN U15675 ( .A(n15356), .B(n15355), .Z(n15360) );
  OR U15676 ( .A(n15358), .B(n15357), .Z(n15359) );
  NAND U15677 ( .A(n15360), .B(n15359), .Z(n15479) );
  NAND U15678 ( .A(b[0]), .B(a[204]), .Z(n15361) );
  XNOR U15679 ( .A(b[1]), .B(n15361), .Z(n15363) );
  NAND U15680 ( .A(a[203]), .B(n98), .Z(n15362) );
  AND U15681 ( .A(n15363), .B(n15362), .Z(n15455) );
  XNOR U15682 ( .A(n20154), .B(n15514), .Z(n15461) );
  OR U15683 ( .A(n15461), .B(n20057), .Z(n15366) );
  NANDN U15684 ( .A(n15364), .B(n20098), .Z(n15365) );
  AND U15685 ( .A(n15366), .B(n15365), .Z(n15456) );
  XOR U15686 ( .A(n15455), .B(n15456), .Z(n15458) );
  NAND U15687 ( .A(a[188]), .B(b[15]), .Z(n15457) );
  XOR U15688 ( .A(n15458), .B(n15457), .Z(n15476) );
  NAND U15689 ( .A(n19722), .B(n15367), .Z(n15369) );
  XNOR U15690 ( .A(b[5]), .B(n16165), .Z(n15467) );
  NANDN U15691 ( .A(n19640), .B(n15467), .Z(n15368) );
  NAND U15692 ( .A(n15369), .B(n15368), .Z(n15452) );
  XNOR U15693 ( .A(n19714), .B(n16009), .Z(n15470) );
  NANDN U15694 ( .A(n15470), .B(n19766), .Z(n15372) );
  NANDN U15695 ( .A(n15370), .B(n19767), .Z(n15371) );
  NAND U15696 ( .A(n15372), .B(n15371), .Z(n15449) );
  NAND U15697 ( .A(n19554), .B(n15373), .Z(n15375) );
  IV U15698 ( .A(a[202]), .Z(n16294) );
  XNOR U15699 ( .A(b[3]), .B(n16294), .Z(n15473) );
  NANDN U15700 ( .A(n19521), .B(n15473), .Z(n15374) );
  AND U15701 ( .A(n15375), .B(n15374), .Z(n15450) );
  XNOR U15702 ( .A(n15449), .B(n15450), .Z(n15451) );
  XOR U15703 ( .A(n15452), .B(n15451), .Z(n15477) );
  XOR U15704 ( .A(n15476), .B(n15477), .Z(n15478) );
  XNOR U15705 ( .A(n15479), .B(n15478), .Z(n15427) );
  NAND U15706 ( .A(n15377), .B(n15376), .Z(n15381) );
  NAND U15707 ( .A(n15379), .B(n15378), .Z(n15380) );
  NAND U15708 ( .A(n15381), .B(n15380), .Z(n15428) );
  XOR U15709 ( .A(n15427), .B(n15428), .Z(n15430) );
  XNOR U15710 ( .A(n20052), .B(n15697), .Z(n15433) );
  OR U15711 ( .A(n15433), .B(n20020), .Z(n15384) );
  NANDN U15712 ( .A(n15382), .B(n19960), .Z(n15383) );
  NAND U15713 ( .A(n15384), .B(n15383), .Z(n15446) );
  XNOR U15714 ( .A(n102), .B(n15385), .Z(n15437) );
  OR U15715 ( .A(n15437), .B(n20121), .Z(n15388) );
  NANDN U15716 ( .A(n15386), .B(n20122), .Z(n15387) );
  NAND U15717 ( .A(n15388), .B(n15387), .Z(n15443) );
  XNOR U15718 ( .A(n19975), .B(n15826), .Z(n15440) );
  NANDN U15719 ( .A(n15440), .B(n19883), .Z(n15391) );
  NANDN U15720 ( .A(n15389), .B(n19937), .Z(n15390) );
  AND U15721 ( .A(n15391), .B(n15390), .Z(n15444) );
  XNOR U15722 ( .A(n15443), .B(n15444), .Z(n15445) );
  XNOR U15723 ( .A(n15446), .B(n15445), .Z(n15482) );
  NANDN U15724 ( .A(n15393), .B(n15392), .Z(n15397) );
  NAND U15725 ( .A(n15395), .B(n15394), .Z(n15396) );
  NAND U15726 ( .A(n15397), .B(n15396), .Z(n15483) );
  XNOR U15727 ( .A(n15482), .B(n15483), .Z(n15484) );
  NANDN U15728 ( .A(n15399), .B(n15398), .Z(n15403) );
  NAND U15729 ( .A(n15401), .B(n15400), .Z(n15402) );
  AND U15730 ( .A(n15403), .B(n15402), .Z(n15485) );
  XNOR U15731 ( .A(n15484), .B(n15485), .Z(n15429) );
  XNOR U15732 ( .A(n15430), .B(n15429), .Z(n15488) );
  NANDN U15733 ( .A(n15405), .B(n15404), .Z(n15409) );
  NAND U15734 ( .A(n15407), .B(n15406), .Z(n15408) );
  NAND U15735 ( .A(n15409), .B(n15408), .Z(n15489) );
  XNOR U15736 ( .A(n15488), .B(n15489), .Z(n15490) );
  XOR U15737 ( .A(n15491), .B(n15490), .Z(n15421) );
  NANDN U15738 ( .A(n15411), .B(n15410), .Z(n15415) );
  NANDN U15739 ( .A(n15413), .B(n15412), .Z(n15414) );
  NAND U15740 ( .A(n15415), .B(n15414), .Z(n15422) );
  XNOR U15741 ( .A(n15421), .B(n15422), .Z(n15423) );
  XNOR U15742 ( .A(n15424), .B(n15423), .Z(n15494) );
  XNOR U15743 ( .A(n15494), .B(sreg[444]), .Z(n15496) );
  NAND U15744 ( .A(n15416), .B(sreg[443]), .Z(n15420) );
  OR U15745 ( .A(n15418), .B(n15417), .Z(n15419) );
  AND U15746 ( .A(n15420), .B(n15419), .Z(n15495) );
  XOR U15747 ( .A(n15496), .B(n15495), .Z(c[444]) );
  NANDN U15748 ( .A(n15422), .B(n15421), .Z(n15426) );
  NAND U15749 ( .A(n15424), .B(n15423), .Z(n15425) );
  NAND U15750 ( .A(n15426), .B(n15425), .Z(n15502) );
  NANDN U15751 ( .A(n15428), .B(n15427), .Z(n15432) );
  OR U15752 ( .A(n15430), .B(n15429), .Z(n15431) );
  NAND U15753 ( .A(n15432), .B(n15431), .Z(n15569) );
  XNOR U15754 ( .A(n20052), .B(n15775), .Z(n15511) );
  OR U15755 ( .A(n15511), .B(n20020), .Z(n15435) );
  NANDN U15756 ( .A(n15433), .B(n19960), .Z(n15434) );
  NAND U15757 ( .A(n15435), .B(n15434), .Z(n15524) );
  XNOR U15758 ( .A(n102), .B(n15436), .Z(n15515) );
  OR U15759 ( .A(n15515), .B(n20121), .Z(n15439) );
  NANDN U15760 ( .A(n15437), .B(n20122), .Z(n15438) );
  NAND U15761 ( .A(n15439), .B(n15438), .Z(n15521) );
  XNOR U15762 ( .A(n19975), .B(n15931), .Z(n15518) );
  NANDN U15763 ( .A(n15518), .B(n19883), .Z(n15442) );
  NANDN U15764 ( .A(n15440), .B(n19937), .Z(n15441) );
  AND U15765 ( .A(n15442), .B(n15441), .Z(n15522) );
  XNOR U15766 ( .A(n15521), .B(n15522), .Z(n15523) );
  XNOR U15767 ( .A(n15524), .B(n15523), .Z(n15560) );
  NANDN U15768 ( .A(n15444), .B(n15443), .Z(n15448) );
  NAND U15769 ( .A(n15446), .B(n15445), .Z(n15447) );
  NAND U15770 ( .A(n15448), .B(n15447), .Z(n15561) );
  XNOR U15771 ( .A(n15560), .B(n15561), .Z(n15562) );
  NANDN U15772 ( .A(n15450), .B(n15449), .Z(n15454) );
  NAND U15773 ( .A(n15452), .B(n15451), .Z(n15453) );
  AND U15774 ( .A(n15454), .B(n15453), .Z(n15563) );
  XNOR U15775 ( .A(n15562), .B(n15563), .Z(n15507) );
  NANDN U15776 ( .A(n15456), .B(n15455), .Z(n15460) );
  OR U15777 ( .A(n15458), .B(n15457), .Z(n15459) );
  NAND U15778 ( .A(n15460), .B(n15459), .Z(n15557) );
  XNOR U15779 ( .A(n20154), .B(n15619), .Z(n15542) );
  OR U15780 ( .A(n15542), .B(n20057), .Z(n15463) );
  NANDN U15781 ( .A(n15461), .B(n20098), .Z(n15462) );
  AND U15782 ( .A(n15463), .B(n15462), .Z(n15534) );
  NAND U15783 ( .A(b[0]), .B(a[205]), .Z(n15464) );
  XNOR U15784 ( .A(b[1]), .B(n15464), .Z(n15466) );
  NAND U15785 ( .A(a[204]), .B(n98), .Z(n15465) );
  AND U15786 ( .A(n15466), .B(n15465), .Z(n15533) );
  XOR U15787 ( .A(n15534), .B(n15533), .Z(n15536) );
  NAND U15788 ( .A(a[189]), .B(b[15]), .Z(n15535) );
  XOR U15789 ( .A(n15536), .B(n15535), .Z(n15554) );
  NAND U15790 ( .A(n19722), .B(n15467), .Z(n15469) );
  XNOR U15791 ( .A(b[5]), .B(n16216), .Z(n15545) );
  NANDN U15792 ( .A(n19640), .B(n15545), .Z(n15468) );
  NAND U15793 ( .A(n15469), .B(n15468), .Z(n15530) );
  XNOR U15794 ( .A(n19714), .B(n16060), .Z(n15548) );
  NANDN U15795 ( .A(n15548), .B(n19766), .Z(n15472) );
  NANDN U15796 ( .A(n15470), .B(n19767), .Z(n15471) );
  NAND U15797 ( .A(n15472), .B(n15471), .Z(n15527) );
  NAND U15798 ( .A(n19554), .B(n15473), .Z(n15475) );
  IV U15799 ( .A(a[203]), .Z(n16399) );
  XNOR U15800 ( .A(b[3]), .B(n16399), .Z(n15551) );
  NANDN U15801 ( .A(n19521), .B(n15551), .Z(n15474) );
  AND U15802 ( .A(n15475), .B(n15474), .Z(n15528) );
  XNOR U15803 ( .A(n15527), .B(n15528), .Z(n15529) );
  XOR U15804 ( .A(n15530), .B(n15529), .Z(n15555) );
  XOR U15805 ( .A(n15554), .B(n15555), .Z(n15556) );
  XNOR U15806 ( .A(n15557), .B(n15556), .Z(n15505) );
  NAND U15807 ( .A(n15477), .B(n15476), .Z(n15481) );
  NAND U15808 ( .A(n15479), .B(n15478), .Z(n15480) );
  NAND U15809 ( .A(n15481), .B(n15480), .Z(n15506) );
  XOR U15810 ( .A(n15505), .B(n15506), .Z(n15508) );
  XNOR U15811 ( .A(n15507), .B(n15508), .Z(n15566) );
  NANDN U15812 ( .A(n15483), .B(n15482), .Z(n15487) );
  NAND U15813 ( .A(n15485), .B(n15484), .Z(n15486) );
  NAND U15814 ( .A(n15487), .B(n15486), .Z(n15567) );
  XNOR U15815 ( .A(n15566), .B(n15567), .Z(n15568) );
  XOR U15816 ( .A(n15569), .B(n15568), .Z(n15499) );
  NANDN U15817 ( .A(n15489), .B(n15488), .Z(n15493) );
  NANDN U15818 ( .A(n15491), .B(n15490), .Z(n15492) );
  NAND U15819 ( .A(n15493), .B(n15492), .Z(n15500) );
  XNOR U15820 ( .A(n15499), .B(n15500), .Z(n15501) );
  XNOR U15821 ( .A(n15502), .B(n15501), .Z(n15572) );
  XNOR U15822 ( .A(n15572), .B(sreg[445]), .Z(n15574) );
  NAND U15823 ( .A(n15494), .B(sreg[444]), .Z(n15498) );
  OR U15824 ( .A(n15496), .B(n15495), .Z(n15497) );
  AND U15825 ( .A(n15498), .B(n15497), .Z(n15573) );
  XOR U15826 ( .A(n15574), .B(n15573), .Z(c[445]) );
  NANDN U15827 ( .A(n15500), .B(n15499), .Z(n15504) );
  NAND U15828 ( .A(n15502), .B(n15501), .Z(n15503) );
  NAND U15829 ( .A(n15504), .B(n15503), .Z(n15580) );
  NANDN U15830 ( .A(n15506), .B(n15505), .Z(n15510) );
  OR U15831 ( .A(n15508), .B(n15507), .Z(n15509) );
  NAND U15832 ( .A(n15510), .B(n15509), .Z(n15647) );
  XNOR U15833 ( .A(n20052), .B(n15826), .Z(n15616) );
  OR U15834 ( .A(n15616), .B(n20020), .Z(n15513) );
  NANDN U15835 ( .A(n15511), .B(n19960), .Z(n15512) );
  NAND U15836 ( .A(n15513), .B(n15512), .Z(n15629) );
  XNOR U15837 ( .A(n102), .B(n15514), .Z(n15620) );
  OR U15838 ( .A(n15620), .B(n20121), .Z(n15517) );
  NANDN U15839 ( .A(n15515), .B(n20122), .Z(n15516) );
  NAND U15840 ( .A(n15517), .B(n15516), .Z(n15626) );
  XNOR U15841 ( .A(n19975), .B(n16009), .Z(n15623) );
  NANDN U15842 ( .A(n15623), .B(n19883), .Z(n15520) );
  NANDN U15843 ( .A(n15518), .B(n19937), .Z(n15519) );
  AND U15844 ( .A(n15520), .B(n15519), .Z(n15627) );
  XNOR U15845 ( .A(n15626), .B(n15627), .Z(n15628) );
  XNOR U15846 ( .A(n15629), .B(n15628), .Z(n15638) );
  NANDN U15847 ( .A(n15522), .B(n15521), .Z(n15526) );
  NAND U15848 ( .A(n15524), .B(n15523), .Z(n15525) );
  NAND U15849 ( .A(n15526), .B(n15525), .Z(n15639) );
  XNOR U15850 ( .A(n15638), .B(n15639), .Z(n15640) );
  NANDN U15851 ( .A(n15528), .B(n15527), .Z(n15532) );
  NAND U15852 ( .A(n15530), .B(n15529), .Z(n15531) );
  AND U15853 ( .A(n15532), .B(n15531), .Z(n15641) );
  XNOR U15854 ( .A(n15640), .B(n15641), .Z(n15585) );
  NANDN U15855 ( .A(n15534), .B(n15533), .Z(n15538) );
  OR U15856 ( .A(n15536), .B(n15535), .Z(n15537) );
  NAND U15857 ( .A(n15538), .B(n15537), .Z(n15613) );
  NAND U15858 ( .A(b[0]), .B(a[206]), .Z(n15539) );
  XNOR U15859 ( .A(b[1]), .B(n15539), .Z(n15541) );
  NAND U15860 ( .A(a[205]), .B(n98), .Z(n15540) );
  AND U15861 ( .A(n15541), .B(n15540), .Z(n15589) );
  XNOR U15862 ( .A(n20154), .B(n15697), .Z(n15598) );
  OR U15863 ( .A(n15598), .B(n20057), .Z(n15544) );
  NANDN U15864 ( .A(n15542), .B(n20098), .Z(n15543) );
  AND U15865 ( .A(n15544), .B(n15543), .Z(n15590) );
  XOR U15866 ( .A(n15589), .B(n15590), .Z(n15592) );
  NAND U15867 ( .A(a[190]), .B(b[15]), .Z(n15591) );
  XOR U15868 ( .A(n15592), .B(n15591), .Z(n15610) );
  NAND U15869 ( .A(n19722), .B(n15545), .Z(n15547) );
  XNOR U15870 ( .A(b[5]), .B(n16294), .Z(n15601) );
  NANDN U15871 ( .A(n19640), .B(n15601), .Z(n15546) );
  NAND U15872 ( .A(n15547), .B(n15546), .Z(n15635) );
  XNOR U15873 ( .A(n19714), .B(n16165), .Z(n15604) );
  NANDN U15874 ( .A(n15604), .B(n19766), .Z(n15550) );
  NANDN U15875 ( .A(n15548), .B(n19767), .Z(n15549) );
  NAND U15876 ( .A(n15550), .B(n15549), .Z(n15632) );
  NAND U15877 ( .A(n19554), .B(n15551), .Z(n15553) );
  IV U15878 ( .A(a[204]), .Z(n16477) );
  XNOR U15879 ( .A(b[3]), .B(n16477), .Z(n15607) );
  NANDN U15880 ( .A(n19521), .B(n15607), .Z(n15552) );
  AND U15881 ( .A(n15553), .B(n15552), .Z(n15633) );
  XNOR U15882 ( .A(n15632), .B(n15633), .Z(n15634) );
  XOR U15883 ( .A(n15635), .B(n15634), .Z(n15611) );
  XOR U15884 ( .A(n15610), .B(n15611), .Z(n15612) );
  XNOR U15885 ( .A(n15613), .B(n15612), .Z(n15583) );
  NAND U15886 ( .A(n15555), .B(n15554), .Z(n15559) );
  NAND U15887 ( .A(n15557), .B(n15556), .Z(n15558) );
  NAND U15888 ( .A(n15559), .B(n15558), .Z(n15584) );
  XOR U15889 ( .A(n15583), .B(n15584), .Z(n15586) );
  XNOR U15890 ( .A(n15585), .B(n15586), .Z(n15644) );
  NANDN U15891 ( .A(n15561), .B(n15560), .Z(n15565) );
  NAND U15892 ( .A(n15563), .B(n15562), .Z(n15564) );
  NAND U15893 ( .A(n15565), .B(n15564), .Z(n15645) );
  XNOR U15894 ( .A(n15644), .B(n15645), .Z(n15646) );
  XOR U15895 ( .A(n15647), .B(n15646), .Z(n15577) );
  NANDN U15896 ( .A(n15567), .B(n15566), .Z(n15571) );
  NANDN U15897 ( .A(n15569), .B(n15568), .Z(n15570) );
  NAND U15898 ( .A(n15571), .B(n15570), .Z(n15578) );
  XNOR U15899 ( .A(n15577), .B(n15578), .Z(n15579) );
  XNOR U15900 ( .A(n15580), .B(n15579), .Z(n15650) );
  XNOR U15901 ( .A(n15650), .B(sreg[446]), .Z(n15652) );
  NAND U15902 ( .A(n15572), .B(sreg[445]), .Z(n15576) );
  OR U15903 ( .A(n15574), .B(n15573), .Z(n15575) );
  AND U15904 ( .A(n15576), .B(n15575), .Z(n15651) );
  XOR U15905 ( .A(n15652), .B(n15651), .Z(c[446]) );
  NANDN U15906 ( .A(n15578), .B(n15577), .Z(n15582) );
  NAND U15907 ( .A(n15580), .B(n15579), .Z(n15581) );
  NAND U15908 ( .A(n15582), .B(n15581), .Z(n15658) );
  NANDN U15909 ( .A(n15584), .B(n15583), .Z(n15588) );
  OR U15910 ( .A(n15586), .B(n15585), .Z(n15587) );
  NAND U15911 ( .A(n15588), .B(n15587), .Z(n15725) );
  NANDN U15912 ( .A(n15590), .B(n15589), .Z(n15594) );
  OR U15913 ( .A(n15592), .B(n15591), .Z(n15593) );
  NAND U15914 ( .A(n15594), .B(n15593), .Z(n15691) );
  NAND U15915 ( .A(b[0]), .B(a[207]), .Z(n15595) );
  XNOR U15916 ( .A(b[1]), .B(n15595), .Z(n15597) );
  NAND U15917 ( .A(a[206]), .B(n98), .Z(n15596) );
  AND U15918 ( .A(n15597), .B(n15596), .Z(n15667) );
  XNOR U15919 ( .A(n20154), .B(n15775), .Z(n15673) );
  OR U15920 ( .A(n15673), .B(n20057), .Z(n15600) );
  NANDN U15921 ( .A(n15598), .B(n20098), .Z(n15599) );
  AND U15922 ( .A(n15600), .B(n15599), .Z(n15668) );
  XOR U15923 ( .A(n15667), .B(n15668), .Z(n15670) );
  NAND U15924 ( .A(a[191]), .B(b[15]), .Z(n15669) );
  XOR U15925 ( .A(n15670), .B(n15669), .Z(n15688) );
  NAND U15926 ( .A(n19722), .B(n15601), .Z(n15603) );
  XNOR U15927 ( .A(b[5]), .B(n16399), .Z(n15679) );
  NANDN U15928 ( .A(n19640), .B(n15679), .Z(n15602) );
  NAND U15929 ( .A(n15603), .B(n15602), .Z(n15713) );
  XNOR U15930 ( .A(n19714), .B(n16216), .Z(n15682) );
  NANDN U15931 ( .A(n15682), .B(n19766), .Z(n15606) );
  NANDN U15932 ( .A(n15604), .B(n19767), .Z(n15605) );
  NAND U15933 ( .A(n15606), .B(n15605), .Z(n15710) );
  NAND U15934 ( .A(n19554), .B(n15607), .Z(n15609) );
  IV U15935 ( .A(a[205]), .Z(n16555) );
  XNOR U15936 ( .A(b[3]), .B(n16555), .Z(n15685) );
  NANDN U15937 ( .A(n19521), .B(n15685), .Z(n15608) );
  AND U15938 ( .A(n15609), .B(n15608), .Z(n15711) );
  XNOR U15939 ( .A(n15710), .B(n15711), .Z(n15712) );
  XOR U15940 ( .A(n15713), .B(n15712), .Z(n15689) );
  XOR U15941 ( .A(n15688), .B(n15689), .Z(n15690) );
  XNOR U15942 ( .A(n15691), .B(n15690), .Z(n15661) );
  NAND U15943 ( .A(n15611), .B(n15610), .Z(n15615) );
  NAND U15944 ( .A(n15613), .B(n15612), .Z(n15614) );
  NAND U15945 ( .A(n15615), .B(n15614), .Z(n15662) );
  XOR U15946 ( .A(n15661), .B(n15662), .Z(n15664) );
  XNOR U15947 ( .A(n20052), .B(n15931), .Z(n15694) );
  OR U15948 ( .A(n15694), .B(n20020), .Z(n15618) );
  NANDN U15949 ( .A(n15616), .B(n19960), .Z(n15617) );
  NAND U15950 ( .A(n15618), .B(n15617), .Z(n15707) );
  XNOR U15951 ( .A(n102), .B(n15619), .Z(n15698) );
  OR U15952 ( .A(n15698), .B(n20121), .Z(n15622) );
  NANDN U15953 ( .A(n15620), .B(n20122), .Z(n15621) );
  NAND U15954 ( .A(n15622), .B(n15621), .Z(n15704) );
  XNOR U15955 ( .A(n19975), .B(n16060), .Z(n15701) );
  NANDN U15956 ( .A(n15701), .B(n19883), .Z(n15625) );
  NANDN U15957 ( .A(n15623), .B(n19937), .Z(n15624) );
  AND U15958 ( .A(n15625), .B(n15624), .Z(n15705) );
  XNOR U15959 ( .A(n15704), .B(n15705), .Z(n15706) );
  XNOR U15960 ( .A(n15707), .B(n15706), .Z(n15716) );
  NANDN U15961 ( .A(n15627), .B(n15626), .Z(n15631) );
  NAND U15962 ( .A(n15629), .B(n15628), .Z(n15630) );
  NAND U15963 ( .A(n15631), .B(n15630), .Z(n15717) );
  XNOR U15964 ( .A(n15716), .B(n15717), .Z(n15718) );
  NANDN U15965 ( .A(n15633), .B(n15632), .Z(n15637) );
  NAND U15966 ( .A(n15635), .B(n15634), .Z(n15636) );
  AND U15967 ( .A(n15637), .B(n15636), .Z(n15719) );
  XNOR U15968 ( .A(n15718), .B(n15719), .Z(n15663) );
  XNOR U15969 ( .A(n15664), .B(n15663), .Z(n15722) );
  NANDN U15970 ( .A(n15639), .B(n15638), .Z(n15643) );
  NAND U15971 ( .A(n15641), .B(n15640), .Z(n15642) );
  NAND U15972 ( .A(n15643), .B(n15642), .Z(n15723) );
  XNOR U15973 ( .A(n15722), .B(n15723), .Z(n15724) );
  XOR U15974 ( .A(n15725), .B(n15724), .Z(n15655) );
  NANDN U15975 ( .A(n15645), .B(n15644), .Z(n15649) );
  NANDN U15976 ( .A(n15647), .B(n15646), .Z(n15648) );
  NAND U15977 ( .A(n15649), .B(n15648), .Z(n15656) );
  XNOR U15978 ( .A(n15655), .B(n15656), .Z(n15657) );
  XNOR U15979 ( .A(n15658), .B(n15657), .Z(n15728) );
  XNOR U15980 ( .A(n15728), .B(sreg[447]), .Z(n15730) );
  NAND U15981 ( .A(n15650), .B(sreg[446]), .Z(n15654) );
  OR U15982 ( .A(n15652), .B(n15651), .Z(n15653) );
  AND U15983 ( .A(n15654), .B(n15653), .Z(n15729) );
  XOR U15984 ( .A(n15730), .B(n15729), .Z(c[447]) );
  NANDN U15985 ( .A(n15656), .B(n15655), .Z(n15660) );
  NAND U15986 ( .A(n15658), .B(n15657), .Z(n15659) );
  NAND U15987 ( .A(n15660), .B(n15659), .Z(n15736) );
  NANDN U15988 ( .A(n15662), .B(n15661), .Z(n15666) );
  OR U15989 ( .A(n15664), .B(n15663), .Z(n15665) );
  NAND U15990 ( .A(n15666), .B(n15665), .Z(n15803) );
  NANDN U15991 ( .A(n15668), .B(n15667), .Z(n15672) );
  OR U15992 ( .A(n15670), .B(n15669), .Z(n15671) );
  NAND U15993 ( .A(n15672), .B(n15671), .Z(n15769) );
  XNOR U15994 ( .A(n20154), .B(n15826), .Z(n15751) );
  OR U15995 ( .A(n15751), .B(n20057), .Z(n15675) );
  NANDN U15996 ( .A(n15673), .B(n20098), .Z(n15674) );
  AND U15997 ( .A(n15675), .B(n15674), .Z(n15746) );
  NAND U15998 ( .A(b[0]), .B(a[208]), .Z(n15676) );
  XNOR U15999 ( .A(b[1]), .B(n15676), .Z(n15678) );
  NAND U16000 ( .A(a[207]), .B(n98), .Z(n15677) );
  AND U16001 ( .A(n15678), .B(n15677), .Z(n15745) );
  XOR U16002 ( .A(n15746), .B(n15745), .Z(n15748) );
  NAND U16003 ( .A(a[192]), .B(b[15]), .Z(n15747) );
  XOR U16004 ( .A(n15748), .B(n15747), .Z(n15766) );
  NAND U16005 ( .A(n19722), .B(n15679), .Z(n15681) );
  XNOR U16006 ( .A(b[5]), .B(n16477), .Z(n15757) );
  NANDN U16007 ( .A(n19640), .B(n15757), .Z(n15680) );
  NAND U16008 ( .A(n15681), .B(n15680), .Z(n15791) );
  XNOR U16009 ( .A(n19714), .B(n16294), .Z(n15760) );
  NANDN U16010 ( .A(n15760), .B(n19766), .Z(n15684) );
  NANDN U16011 ( .A(n15682), .B(n19767), .Z(n15683) );
  NAND U16012 ( .A(n15684), .B(n15683), .Z(n15788) );
  NAND U16013 ( .A(n19554), .B(n15685), .Z(n15687) );
  IV U16014 ( .A(a[206]), .Z(n16606) );
  XNOR U16015 ( .A(b[3]), .B(n16606), .Z(n15763) );
  NANDN U16016 ( .A(n19521), .B(n15763), .Z(n15686) );
  AND U16017 ( .A(n15687), .B(n15686), .Z(n15789) );
  XNOR U16018 ( .A(n15788), .B(n15789), .Z(n15790) );
  XOR U16019 ( .A(n15791), .B(n15790), .Z(n15767) );
  XOR U16020 ( .A(n15766), .B(n15767), .Z(n15768) );
  XNOR U16021 ( .A(n15769), .B(n15768), .Z(n15739) );
  NAND U16022 ( .A(n15689), .B(n15688), .Z(n15693) );
  NAND U16023 ( .A(n15691), .B(n15690), .Z(n15692) );
  NAND U16024 ( .A(n15693), .B(n15692), .Z(n15740) );
  XOR U16025 ( .A(n15739), .B(n15740), .Z(n15742) );
  XNOR U16026 ( .A(n20052), .B(n16009), .Z(n15772) );
  OR U16027 ( .A(n15772), .B(n20020), .Z(n15696) );
  NANDN U16028 ( .A(n15694), .B(n19960), .Z(n15695) );
  NAND U16029 ( .A(n15696), .B(n15695), .Z(n15785) );
  XNOR U16030 ( .A(n102), .B(n15697), .Z(n15776) );
  OR U16031 ( .A(n15776), .B(n20121), .Z(n15700) );
  NANDN U16032 ( .A(n15698), .B(n20122), .Z(n15699) );
  NAND U16033 ( .A(n15700), .B(n15699), .Z(n15782) );
  XNOR U16034 ( .A(n19975), .B(n16165), .Z(n15779) );
  NANDN U16035 ( .A(n15779), .B(n19883), .Z(n15703) );
  NANDN U16036 ( .A(n15701), .B(n19937), .Z(n15702) );
  AND U16037 ( .A(n15703), .B(n15702), .Z(n15783) );
  XNOR U16038 ( .A(n15782), .B(n15783), .Z(n15784) );
  XNOR U16039 ( .A(n15785), .B(n15784), .Z(n15794) );
  NANDN U16040 ( .A(n15705), .B(n15704), .Z(n15709) );
  NAND U16041 ( .A(n15707), .B(n15706), .Z(n15708) );
  NAND U16042 ( .A(n15709), .B(n15708), .Z(n15795) );
  XNOR U16043 ( .A(n15794), .B(n15795), .Z(n15796) );
  NANDN U16044 ( .A(n15711), .B(n15710), .Z(n15715) );
  NAND U16045 ( .A(n15713), .B(n15712), .Z(n15714) );
  AND U16046 ( .A(n15715), .B(n15714), .Z(n15797) );
  XNOR U16047 ( .A(n15796), .B(n15797), .Z(n15741) );
  XNOR U16048 ( .A(n15742), .B(n15741), .Z(n15800) );
  NANDN U16049 ( .A(n15717), .B(n15716), .Z(n15721) );
  NAND U16050 ( .A(n15719), .B(n15718), .Z(n15720) );
  NAND U16051 ( .A(n15721), .B(n15720), .Z(n15801) );
  XNOR U16052 ( .A(n15800), .B(n15801), .Z(n15802) );
  XOR U16053 ( .A(n15803), .B(n15802), .Z(n15733) );
  NANDN U16054 ( .A(n15723), .B(n15722), .Z(n15727) );
  NANDN U16055 ( .A(n15725), .B(n15724), .Z(n15726) );
  NAND U16056 ( .A(n15727), .B(n15726), .Z(n15734) );
  XNOR U16057 ( .A(n15733), .B(n15734), .Z(n15735) );
  XNOR U16058 ( .A(n15736), .B(n15735), .Z(n15806) );
  XNOR U16059 ( .A(n15806), .B(sreg[448]), .Z(n15808) );
  NAND U16060 ( .A(n15728), .B(sreg[447]), .Z(n15732) );
  OR U16061 ( .A(n15730), .B(n15729), .Z(n15731) );
  AND U16062 ( .A(n15732), .B(n15731), .Z(n15807) );
  XOR U16063 ( .A(n15808), .B(n15807), .Z(c[448]) );
  NANDN U16064 ( .A(n15734), .B(n15733), .Z(n15738) );
  NAND U16065 ( .A(n15736), .B(n15735), .Z(n15737) );
  NAND U16066 ( .A(n15738), .B(n15737), .Z(n15814) );
  NANDN U16067 ( .A(n15740), .B(n15739), .Z(n15744) );
  OR U16068 ( .A(n15742), .B(n15741), .Z(n15743) );
  NAND U16069 ( .A(n15744), .B(n15743), .Z(n15881) );
  NANDN U16070 ( .A(n15746), .B(n15745), .Z(n15750) );
  OR U16071 ( .A(n15748), .B(n15747), .Z(n15749) );
  NAND U16072 ( .A(n15750), .B(n15749), .Z(n15869) );
  XNOR U16073 ( .A(n20154), .B(n15931), .Z(n15854) );
  OR U16074 ( .A(n15854), .B(n20057), .Z(n15753) );
  NANDN U16075 ( .A(n15751), .B(n20098), .Z(n15752) );
  AND U16076 ( .A(n15753), .B(n15752), .Z(n15846) );
  NAND U16077 ( .A(b[0]), .B(a[209]), .Z(n15754) );
  XNOR U16078 ( .A(b[1]), .B(n15754), .Z(n15756) );
  NAND U16079 ( .A(a[208]), .B(n98), .Z(n15755) );
  AND U16080 ( .A(n15756), .B(n15755), .Z(n15845) );
  XOR U16081 ( .A(n15846), .B(n15845), .Z(n15848) );
  NAND U16082 ( .A(a[193]), .B(b[15]), .Z(n15847) );
  XOR U16083 ( .A(n15848), .B(n15847), .Z(n15866) );
  NAND U16084 ( .A(n19722), .B(n15757), .Z(n15759) );
  XNOR U16085 ( .A(b[5]), .B(n16555), .Z(n15857) );
  NANDN U16086 ( .A(n19640), .B(n15857), .Z(n15758) );
  NAND U16087 ( .A(n15759), .B(n15758), .Z(n15842) );
  XNOR U16088 ( .A(n19714), .B(n16399), .Z(n15860) );
  NANDN U16089 ( .A(n15860), .B(n19766), .Z(n15762) );
  NANDN U16090 ( .A(n15760), .B(n19767), .Z(n15761) );
  NAND U16091 ( .A(n15762), .B(n15761), .Z(n15839) );
  NAND U16092 ( .A(n19554), .B(n15763), .Z(n15765) );
  IV U16093 ( .A(a[207]), .Z(n16684) );
  XNOR U16094 ( .A(b[3]), .B(n16684), .Z(n15863) );
  NANDN U16095 ( .A(n19521), .B(n15863), .Z(n15764) );
  AND U16096 ( .A(n15765), .B(n15764), .Z(n15840) );
  XNOR U16097 ( .A(n15839), .B(n15840), .Z(n15841) );
  XOR U16098 ( .A(n15842), .B(n15841), .Z(n15867) );
  XOR U16099 ( .A(n15866), .B(n15867), .Z(n15868) );
  XNOR U16100 ( .A(n15869), .B(n15868), .Z(n15817) );
  NAND U16101 ( .A(n15767), .B(n15766), .Z(n15771) );
  NAND U16102 ( .A(n15769), .B(n15768), .Z(n15770) );
  NAND U16103 ( .A(n15771), .B(n15770), .Z(n15818) );
  XOR U16104 ( .A(n15817), .B(n15818), .Z(n15820) );
  XNOR U16105 ( .A(n20052), .B(n16060), .Z(n15823) );
  OR U16106 ( .A(n15823), .B(n20020), .Z(n15774) );
  NANDN U16107 ( .A(n15772), .B(n19960), .Z(n15773) );
  NAND U16108 ( .A(n15774), .B(n15773), .Z(n15836) );
  XNOR U16109 ( .A(n102), .B(n15775), .Z(n15827) );
  OR U16110 ( .A(n15827), .B(n20121), .Z(n15778) );
  NANDN U16111 ( .A(n15776), .B(n20122), .Z(n15777) );
  NAND U16112 ( .A(n15778), .B(n15777), .Z(n15833) );
  XNOR U16113 ( .A(n19975), .B(n16216), .Z(n15830) );
  NANDN U16114 ( .A(n15830), .B(n19883), .Z(n15781) );
  NANDN U16115 ( .A(n15779), .B(n19937), .Z(n15780) );
  AND U16116 ( .A(n15781), .B(n15780), .Z(n15834) );
  XNOR U16117 ( .A(n15833), .B(n15834), .Z(n15835) );
  XNOR U16118 ( .A(n15836), .B(n15835), .Z(n15872) );
  NANDN U16119 ( .A(n15783), .B(n15782), .Z(n15787) );
  NAND U16120 ( .A(n15785), .B(n15784), .Z(n15786) );
  NAND U16121 ( .A(n15787), .B(n15786), .Z(n15873) );
  XNOR U16122 ( .A(n15872), .B(n15873), .Z(n15874) );
  NANDN U16123 ( .A(n15789), .B(n15788), .Z(n15793) );
  NAND U16124 ( .A(n15791), .B(n15790), .Z(n15792) );
  AND U16125 ( .A(n15793), .B(n15792), .Z(n15875) );
  XNOR U16126 ( .A(n15874), .B(n15875), .Z(n15819) );
  XNOR U16127 ( .A(n15820), .B(n15819), .Z(n15878) );
  NANDN U16128 ( .A(n15795), .B(n15794), .Z(n15799) );
  NAND U16129 ( .A(n15797), .B(n15796), .Z(n15798) );
  NAND U16130 ( .A(n15799), .B(n15798), .Z(n15879) );
  XNOR U16131 ( .A(n15878), .B(n15879), .Z(n15880) );
  XOR U16132 ( .A(n15881), .B(n15880), .Z(n15811) );
  NANDN U16133 ( .A(n15801), .B(n15800), .Z(n15805) );
  NANDN U16134 ( .A(n15803), .B(n15802), .Z(n15804) );
  NAND U16135 ( .A(n15805), .B(n15804), .Z(n15812) );
  XNOR U16136 ( .A(n15811), .B(n15812), .Z(n15813) );
  XNOR U16137 ( .A(n15814), .B(n15813), .Z(n15884) );
  XNOR U16138 ( .A(n15884), .B(sreg[449]), .Z(n15886) );
  NAND U16139 ( .A(n15806), .B(sreg[448]), .Z(n15810) );
  OR U16140 ( .A(n15808), .B(n15807), .Z(n15809) );
  AND U16141 ( .A(n15810), .B(n15809), .Z(n15885) );
  XOR U16142 ( .A(n15886), .B(n15885), .Z(c[449]) );
  NANDN U16143 ( .A(n15812), .B(n15811), .Z(n15816) );
  NAND U16144 ( .A(n15814), .B(n15813), .Z(n15815) );
  NAND U16145 ( .A(n15816), .B(n15815), .Z(n15892) );
  NANDN U16146 ( .A(n15818), .B(n15817), .Z(n15822) );
  OR U16147 ( .A(n15820), .B(n15819), .Z(n15821) );
  NAND U16148 ( .A(n15822), .B(n15821), .Z(n15959) );
  XNOR U16149 ( .A(n20052), .B(n16165), .Z(n15928) );
  OR U16150 ( .A(n15928), .B(n20020), .Z(n15825) );
  NANDN U16151 ( .A(n15823), .B(n19960), .Z(n15824) );
  NAND U16152 ( .A(n15825), .B(n15824), .Z(n15941) );
  XNOR U16153 ( .A(n102), .B(n15826), .Z(n15932) );
  OR U16154 ( .A(n15932), .B(n20121), .Z(n15829) );
  NANDN U16155 ( .A(n15827), .B(n20122), .Z(n15828) );
  NAND U16156 ( .A(n15829), .B(n15828), .Z(n15938) );
  XNOR U16157 ( .A(n19975), .B(n16294), .Z(n15935) );
  NANDN U16158 ( .A(n15935), .B(n19883), .Z(n15832) );
  NANDN U16159 ( .A(n15830), .B(n19937), .Z(n15831) );
  AND U16160 ( .A(n15832), .B(n15831), .Z(n15939) );
  XNOR U16161 ( .A(n15938), .B(n15939), .Z(n15940) );
  XNOR U16162 ( .A(n15941), .B(n15940), .Z(n15950) );
  NANDN U16163 ( .A(n15834), .B(n15833), .Z(n15838) );
  NAND U16164 ( .A(n15836), .B(n15835), .Z(n15837) );
  NAND U16165 ( .A(n15838), .B(n15837), .Z(n15951) );
  XNOR U16166 ( .A(n15950), .B(n15951), .Z(n15952) );
  NANDN U16167 ( .A(n15840), .B(n15839), .Z(n15844) );
  NAND U16168 ( .A(n15842), .B(n15841), .Z(n15843) );
  AND U16169 ( .A(n15844), .B(n15843), .Z(n15953) );
  XNOR U16170 ( .A(n15952), .B(n15953), .Z(n15897) );
  NANDN U16171 ( .A(n15846), .B(n15845), .Z(n15850) );
  OR U16172 ( .A(n15848), .B(n15847), .Z(n15849) );
  NAND U16173 ( .A(n15850), .B(n15849), .Z(n15925) );
  NAND U16174 ( .A(b[0]), .B(a[210]), .Z(n15851) );
  XNOR U16175 ( .A(b[1]), .B(n15851), .Z(n15853) );
  NAND U16176 ( .A(a[209]), .B(n98), .Z(n15852) );
  AND U16177 ( .A(n15853), .B(n15852), .Z(n15901) );
  XNOR U16178 ( .A(n20154), .B(n16009), .Z(n15907) );
  OR U16179 ( .A(n15907), .B(n20057), .Z(n15856) );
  NANDN U16180 ( .A(n15854), .B(n20098), .Z(n15855) );
  AND U16181 ( .A(n15856), .B(n15855), .Z(n15902) );
  XOR U16182 ( .A(n15901), .B(n15902), .Z(n15904) );
  NAND U16183 ( .A(a[194]), .B(b[15]), .Z(n15903) );
  XOR U16184 ( .A(n15904), .B(n15903), .Z(n15922) );
  NAND U16185 ( .A(n19722), .B(n15857), .Z(n15859) );
  XNOR U16186 ( .A(b[5]), .B(n16606), .Z(n15913) );
  NANDN U16187 ( .A(n19640), .B(n15913), .Z(n15858) );
  NAND U16188 ( .A(n15859), .B(n15858), .Z(n15947) );
  XNOR U16189 ( .A(n19714), .B(n16477), .Z(n15916) );
  NANDN U16190 ( .A(n15916), .B(n19766), .Z(n15862) );
  NANDN U16191 ( .A(n15860), .B(n19767), .Z(n15861) );
  NAND U16192 ( .A(n15862), .B(n15861), .Z(n15944) );
  NAND U16193 ( .A(n19554), .B(n15863), .Z(n15865) );
  IV U16194 ( .A(a[208]), .Z(n16762) );
  XNOR U16195 ( .A(b[3]), .B(n16762), .Z(n15919) );
  NANDN U16196 ( .A(n19521), .B(n15919), .Z(n15864) );
  AND U16197 ( .A(n15865), .B(n15864), .Z(n15945) );
  XNOR U16198 ( .A(n15944), .B(n15945), .Z(n15946) );
  XOR U16199 ( .A(n15947), .B(n15946), .Z(n15923) );
  XOR U16200 ( .A(n15922), .B(n15923), .Z(n15924) );
  XNOR U16201 ( .A(n15925), .B(n15924), .Z(n15895) );
  NAND U16202 ( .A(n15867), .B(n15866), .Z(n15871) );
  NAND U16203 ( .A(n15869), .B(n15868), .Z(n15870) );
  NAND U16204 ( .A(n15871), .B(n15870), .Z(n15896) );
  XOR U16205 ( .A(n15895), .B(n15896), .Z(n15898) );
  XNOR U16206 ( .A(n15897), .B(n15898), .Z(n15956) );
  NANDN U16207 ( .A(n15873), .B(n15872), .Z(n15877) );
  NAND U16208 ( .A(n15875), .B(n15874), .Z(n15876) );
  NAND U16209 ( .A(n15877), .B(n15876), .Z(n15957) );
  XNOR U16210 ( .A(n15956), .B(n15957), .Z(n15958) );
  XOR U16211 ( .A(n15959), .B(n15958), .Z(n15889) );
  NANDN U16212 ( .A(n15879), .B(n15878), .Z(n15883) );
  NANDN U16213 ( .A(n15881), .B(n15880), .Z(n15882) );
  NAND U16214 ( .A(n15883), .B(n15882), .Z(n15890) );
  XNOR U16215 ( .A(n15889), .B(n15890), .Z(n15891) );
  XNOR U16216 ( .A(n15892), .B(n15891), .Z(n15962) );
  XNOR U16217 ( .A(n15962), .B(sreg[450]), .Z(n15964) );
  NAND U16218 ( .A(n15884), .B(sreg[449]), .Z(n15888) );
  OR U16219 ( .A(n15886), .B(n15885), .Z(n15887) );
  AND U16220 ( .A(n15888), .B(n15887), .Z(n15963) );
  XOR U16221 ( .A(n15964), .B(n15963), .Z(c[450]) );
  NANDN U16222 ( .A(n15890), .B(n15889), .Z(n15894) );
  NAND U16223 ( .A(n15892), .B(n15891), .Z(n15893) );
  NAND U16224 ( .A(n15894), .B(n15893), .Z(n15970) );
  NANDN U16225 ( .A(n15896), .B(n15895), .Z(n15900) );
  OR U16226 ( .A(n15898), .B(n15897), .Z(n15899) );
  NAND U16227 ( .A(n15900), .B(n15899), .Z(n16037) );
  NANDN U16228 ( .A(n15902), .B(n15901), .Z(n15906) );
  OR U16229 ( .A(n15904), .B(n15903), .Z(n15905) );
  NAND U16230 ( .A(n15906), .B(n15905), .Z(n16003) );
  XNOR U16231 ( .A(n20154), .B(n16060), .Z(n15988) );
  OR U16232 ( .A(n15988), .B(n20057), .Z(n15909) );
  NANDN U16233 ( .A(n15907), .B(n20098), .Z(n15908) );
  AND U16234 ( .A(n15909), .B(n15908), .Z(n15980) );
  NAND U16235 ( .A(b[0]), .B(a[211]), .Z(n15910) );
  XNOR U16236 ( .A(b[1]), .B(n15910), .Z(n15912) );
  NAND U16237 ( .A(a[210]), .B(n98), .Z(n15911) );
  AND U16238 ( .A(n15912), .B(n15911), .Z(n15979) );
  XOR U16239 ( .A(n15980), .B(n15979), .Z(n15982) );
  NAND U16240 ( .A(a[195]), .B(b[15]), .Z(n15981) );
  XOR U16241 ( .A(n15982), .B(n15981), .Z(n16000) );
  NAND U16242 ( .A(n19722), .B(n15913), .Z(n15915) );
  XNOR U16243 ( .A(b[5]), .B(n16684), .Z(n15991) );
  NANDN U16244 ( .A(n19640), .B(n15991), .Z(n15914) );
  NAND U16245 ( .A(n15915), .B(n15914), .Z(n16025) );
  XNOR U16246 ( .A(n19714), .B(n16555), .Z(n15994) );
  NANDN U16247 ( .A(n15994), .B(n19766), .Z(n15918) );
  NANDN U16248 ( .A(n15916), .B(n19767), .Z(n15917) );
  NAND U16249 ( .A(n15918), .B(n15917), .Z(n16022) );
  NAND U16250 ( .A(n19554), .B(n15919), .Z(n15921) );
  IV U16251 ( .A(a[209]), .Z(n16867) );
  XNOR U16252 ( .A(b[3]), .B(n16867), .Z(n15997) );
  NANDN U16253 ( .A(n19521), .B(n15997), .Z(n15920) );
  AND U16254 ( .A(n15921), .B(n15920), .Z(n16023) );
  XNOR U16255 ( .A(n16022), .B(n16023), .Z(n16024) );
  XOR U16256 ( .A(n16025), .B(n16024), .Z(n16001) );
  XOR U16257 ( .A(n16000), .B(n16001), .Z(n16002) );
  XNOR U16258 ( .A(n16003), .B(n16002), .Z(n15973) );
  NAND U16259 ( .A(n15923), .B(n15922), .Z(n15927) );
  NAND U16260 ( .A(n15925), .B(n15924), .Z(n15926) );
  NAND U16261 ( .A(n15927), .B(n15926), .Z(n15974) );
  XOR U16262 ( .A(n15973), .B(n15974), .Z(n15976) );
  XNOR U16263 ( .A(n20052), .B(n16216), .Z(n16006) );
  OR U16264 ( .A(n16006), .B(n20020), .Z(n15930) );
  NANDN U16265 ( .A(n15928), .B(n19960), .Z(n15929) );
  NAND U16266 ( .A(n15930), .B(n15929), .Z(n16019) );
  XNOR U16267 ( .A(n102), .B(n15931), .Z(n16010) );
  OR U16268 ( .A(n16010), .B(n20121), .Z(n15934) );
  NANDN U16269 ( .A(n15932), .B(n20122), .Z(n15933) );
  NAND U16270 ( .A(n15934), .B(n15933), .Z(n16016) );
  XNOR U16271 ( .A(n19975), .B(n16399), .Z(n16013) );
  NANDN U16272 ( .A(n16013), .B(n19883), .Z(n15937) );
  NANDN U16273 ( .A(n15935), .B(n19937), .Z(n15936) );
  AND U16274 ( .A(n15937), .B(n15936), .Z(n16017) );
  XNOR U16275 ( .A(n16016), .B(n16017), .Z(n16018) );
  XNOR U16276 ( .A(n16019), .B(n16018), .Z(n16028) );
  NANDN U16277 ( .A(n15939), .B(n15938), .Z(n15943) );
  NAND U16278 ( .A(n15941), .B(n15940), .Z(n15942) );
  NAND U16279 ( .A(n15943), .B(n15942), .Z(n16029) );
  XNOR U16280 ( .A(n16028), .B(n16029), .Z(n16030) );
  NANDN U16281 ( .A(n15945), .B(n15944), .Z(n15949) );
  NAND U16282 ( .A(n15947), .B(n15946), .Z(n15948) );
  AND U16283 ( .A(n15949), .B(n15948), .Z(n16031) );
  XNOR U16284 ( .A(n16030), .B(n16031), .Z(n15975) );
  XNOR U16285 ( .A(n15976), .B(n15975), .Z(n16034) );
  NANDN U16286 ( .A(n15951), .B(n15950), .Z(n15955) );
  NAND U16287 ( .A(n15953), .B(n15952), .Z(n15954) );
  NAND U16288 ( .A(n15955), .B(n15954), .Z(n16035) );
  XNOR U16289 ( .A(n16034), .B(n16035), .Z(n16036) );
  XOR U16290 ( .A(n16037), .B(n16036), .Z(n15967) );
  NANDN U16291 ( .A(n15957), .B(n15956), .Z(n15961) );
  NANDN U16292 ( .A(n15959), .B(n15958), .Z(n15960) );
  NAND U16293 ( .A(n15961), .B(n15960), .Z(n15968) );
  XNOR U16294 ( .A(n15967), .B(n15968), .Z(n15969) );
  XNOR U16295 ( .A(n15970), .B(n15969), .Z(n16040) );
  XNOR U16296 ( .A(n16040), .B(sreg[451]), .Z(n16042) );
  NAND U16297 ( .A(n15962), .B(sreg[450]), .Z(n15966) );
  OR U16298 ( .A(n15964), .B(n15963), .Z(n15965) );
  AND U16299 ( .A(n15966), .B(n15965), .Z(n16041) );
  XOR U16300 ( .A(n16042), .B(n16041), .Z(c[451]) );
  NANDN U16301 ( .A(n15968), .B(n15967), .Z(n15972) );
  NAND U16302 ( .A(n15970), .B(n15969), .Z(n15971) );
  NAND U16303 ( .A(n15972), .B(n15971), .Z(n16048) );
  NANDN U16304 ( .A(n15974), .B(n15973), .Z(n15978) );
  OR U16305 ( .A(n15976), .B(n15975), .Z(n15977) );
  NAND U16306 ( .A(n15978), .B(n15977), .Z(n16115) );
  NANDN U16307 ( .A(n15980), .B(n15979), .Z(n15984) );
  OR U16308 ( .A(n15982), .B(n15981), .Z(n15983) );
  NAND U16309 ( .A(n15984), .B(n15983), .Z(n16103) );
  NAND U16310 ( .A(b[0]), .B(a[212]), .Z(n15985) );
  XNOR U16311 ( .A(b[1]), .B(n15985), .Z(n15987) );
  NAND U16312 ( .A(a[211]), .B(n98), .Z(n15986) );
  AND U16313 ( .A(n15987), .B(n15986), .Z(n16079) );
  XNOR U16314 ( .A(n20154), .B(n16165), .Z(n16088) );
  OR U16315 ( .A(n16088), .B(n20057), .Z(n15990) );
  NANDN U16316 ( .A(n15988), .B(n20098), .Z(n15989) );
  AND U16317 ( .A(n15990), .B(n15989), .Z(n16080) );
  XOR U16318 ( .A(n16079), .B(n16080), .Z(n16082) );
  NAND U16319 ( .A(a[196]), .B(b[15]), .Z(n16081) );
  XOR U16320 ( .A(n16082), .B(n16081), .Z(n16100) );
  NAND U16321 ( .A(n19722), .B(n15991), .Z(n15993) );
  XNOR U16322 ( .A(b[5]), .B(n16762), .Z(n16091) );
  NANDN U16323 ( .A(n19640), .B(n16091), .Z(n15992) );
  NAND U16324 ( .A(n15993), .B(n15992), .Z(n16076) );
  XNOR U16325 ( .A(n19714), .B(n16606), .Z(n16094) );
  NANDN U16326 ( .A(n16094), .B(n19766), .Z(n15996) );
  NANDN U16327 ( .A(n15994), .B(n19767), .Z(n15995) );
  NAND U16328 ( .A(n15996), .B(n15995), .Z(n16073) );
  NAND U16329 ( .A(n19554), .B(n15997), .Z(n15999) );
  IV U16330 ( .A(a[210]), .Z(n16918) );
  XNOR U16331 ( .A(b[3]), .B(n16918), .Z(n16097) );
  NANDN U16332 ( .A(n19521), .B(n16097), .Z(n15998) );
  AND U16333 ( .A(n15999), .B(n15998), .Z(n16074) );
  XNOR U16334 ( .A(n16073), .B(n16074), .Z(n16075) );
  XOR U16335 ( .A(n16076), .B(n16075), .Z(n16101) );
  XOR U16336 ( .A(n16100), .B(n16101), .Z(n16102) );
  XNOR U16337 ( .A(n16103), .B(n16102), .Z(n16051) );
  NAND U16338 ( .A(n16001), .B(n16000), .Z(n16005) );
  NAND U16339 ( .A(n16003), .B(n16002), .Z(n16004) );
  NAND U16340 ( .A(n16005), .B(n16004), .Z(n16052) );
  XOR U16341 ( .A(n16051), .B(n16052), .Z(n16054) );
  XNOR U16342 ( .A(n20052), .B(n16294), .Z(n16057) );
  OR U16343 ( .A(n16057), .B(n20020), .Z(n16008) );
  NANDN U16344 ( .A(n16006), .B(n19960), .Z(n16007) );
  NAND U16345 ( .A(n16008), .B(n16007), .Z(n16070) );
  XNOR U16346 ( .A(n102), .B(n16009), .Z(n16061) );
  OR U16347 ( .A(n16061), .B(n20121), .Z(n16012) );
  NANDN U16348 ( .A(n16010), .B(n20122), .Z(n16011) );
  NAND U16349 ( .A(n16012), .B(n16011), .Z(n16067) );
  XNOR U16350 ( .A(n19975), .B(n16477), .Z(n16064) );
  NANDN U16351 ( .A(n16064), .B(n19883), .Z(n16015) );
  NANDN U16352 ( .A(n16013), .B(n19937), .Z(n16014) );
  AND U16353 ( .A(n16015), .B(n16014), .Z(n16068) );
  XNOR U16354 ( .A(n16067), .B(n16068), .Z(n16069) );
  XNOR U16355 ( .A(n16070), .B(n16069), .Z(n16106) );
  NANDN U16356 ( .A(n16017), .B(n16016), .Z(n16021) );
  NAND U16357 ( .A(n16019), .B(n16018), .Z(n16020) );
  NAND U16358 ( .A(n16021), .B(n16020), .Z(n16107) );
  XNOR U16359 ( .A(n16106), .B(n16107), .Z(n16108) );
  NANDN U16360 ( .A(n16023), .B(n16022), .Z(n16027) );
  NAND U16361 ( .A(n16025), .B(n16024), .Z(n16026) );
  AND U16362 ( .A(n16027), .B(n16026), .Z(n16109) );
  XNOR U16363 ( .A(n16108), .B(n16109), .Z(n16053) );
  XNOR U16364 ( .A(n16054), .B(n16053), .Z(n16112) );
  NANDN U16365 ( .A(n16029), .B(n16028), .Z(n16033) );
  NAND U16366 ( .A(n16031), .B(n16030), .Z(n16032) );
  NAND U16367 ( .A(n16033), .B(n16032), .Z(n16113) );
  XNOR U16368 ( .A(n16112), .B(n16113), .Z(n16114) );
  XOR U16369 ( .A(n16115), .B(n16114), .Z(n16045) );
  NANDN U16370 ( .A(n16035), .B(n16034), .Z(n16039) );
  NANDN U16371 ( .A(n16037), .B(n16036), .Z(n16038) );
  NAND U16372 ( .A(n16039), .B(n16038), .Z(n16046) );
  XNOR U16373 ( .A(n16045), .B(n16046), .Z(n16047) );
  XNOR U16374 ( .A(n16048), .B(n16047), .Z(n16118) );
  XNOR U16375 ( .A(n16118), .B(sreg[452]), .Z(n16120) );
  NAND U16376 ( .A(n16040), .B(sreg[451]), .Z(n16044) );
  OR U16377 ( .A(n16042), .B(n16041), .Z(n16043) );
  AND U16378 ( .A(n16044), .B(n16043), .Z(n16119) );
  XOR U16379 ( .A(n16120), .B(n16119), .Z(c[452]) );
  NANDN U16380 ( .A(n16046), .B(n16045), .Z(n16050) );
  NAND U16381 ( .A(n16048), .B(n16047), .Z(n16049) );
  NAND U16382 ( .A(n16050), .B(n16049), .Z(n16126) );
  NANDN U16383 ( .A(n16052), .B(n16051), .Z(n16056) );
  OR U16384 ( .A(n16054), .B(n16053), .Z(n16055) );
  NAND U16385 ( .A(n16056), .B(n16055), .Z(n16193) );
  XNOR U16386 ( .A(n20052), .B(n16399), .Z(n16162) );
  OR U16387 ( .A(n16162), .B(n20020), .Z(n16059) );
  NANDN U16388 ( .A(n16057), .B(n19960), .Z(n16058) );
  NAND U16389 ( .A(n16059), .B(n16058), .Z(n16175) );
  XNOR U16390 ( .A(n102), .B(n16060), .Z(n16166) );
  OR U16391 ( .A(n16166), .B(n20121), .Z(n16063) );
  NANDN U16392 ( .A(n16061), .B(n20122), .Z(n16062) );
  NAND U16393 ( .A(n16063), .B(n16062), .Z(n16172) );
  XNOR U16394 ( .A(n19975), .B(n16555), .Z(n16169) );
  NANDN U16395 ( .A(n16169), .B(n19883), .Z(n16066) );
  NANDN U16396 ( .A(n16064), .B(n19937), .Z(n16065) );
  AND U16397 ( .A(n16066), .B(n16065), .Z(n16173) );
  XNOR U16398 ( .A(n16172), .B(n16173), .Z(n16174) );
  XNOR U16399 ( .A(n16175), .B(n16174), .Z(n16184) );
  NANDN U16400 ( .A(n16068), .B(n16067), .Z(n16072) );
  NAND U16401 ( .A(n16070), .B(n16069), .Z(n16071) );
  NAND U16402 ( .A(n16072), .B(n16071), .Z(n16185) );
  XNOR U16403 ( .A(n16184), .B(n16185), .Z(n16186) );
  NANDN U16404 ( .A(n16074), .B(n16073), .Z(n16078) );
  NAND U16405 ( .A(n16076), .B(n16075), .Z(n16077) );
  AND U16406 ( .A(n16078), .B(n16077), .Z(n16187) );
  XNOR U16407 ( .A(n16186), .B(n16187), .Z(n16131) );
  NANDN U16408 ( .A(n16080), .B(n16079), .Z(n16084) );
  OR U16409 ( .A(n16082), .B(n16081), .Z(n16083) );
  NAND U16410 ( .A(n16084), .B(n16083), .Z(n16159) );
  NAND U16411 ( .A(b[0]), .B(a[213]), .Z(n16085) );
  XNOR U16412 ( .A(b[1]), .B(n16085), .Z(n16087) );
  NAND U16413 ( .A(a[212]), .B(n98), .Z(n16086) );
  AND U16414 ( .A(n16087), .B(n16086), .Z(n16135) );
  XNOR U16415 ( .A(n20154), .B(n16216), .Z(n16144) );
  OR U16416 ( .A(n16144), .B(n20057), .Z(n16090) );
  NANDN U16417 ( .A(n16088), .B(n20098), .Z(n16089) );
  AND U16418 ( .A(n16090), .B(n16089), .Z(n16136) );
  XOR U16419 ( .A(n16135), .B(n16136), .Z(n16138) );
  NAND U16420 ( .A(a[197]), .B(b[15]), .Z(n16137) );
  XOR U16421 ( .A(n16138), .B(n16137), .Z(n16156) );
  NAND U16422 ( .A(n19722), .B(n16091), .Z(n16093) );
  XNOR U16423 ( .A(b[5]), .B(n16867), .Z(n16147) );
  NANDN U16424 ( .A(n19640), .B(n16147), .Z(n16092) );
  NAND U16425 ( .A(n16093), .B(n16092), .Z(n16181) );
  XNOR U16426 ( .A(n19714), .B(n16684), .Z(n16150) );
  NANDN U16427 ( .A(n16150), .B(n19766), .Z(n16096) );
  NANDN U16428 ( .A(n16094), .B(n19767), .Z(n16095) );
  NAND U16429 ( .A(n16096), .B(n16095), .Z(n16178) );
  NAND U16430 ( .A(n19554), .B(n16097), .Z(n16099) );
  IV U16431 ( .A(a[211]), .Z(n17008) );
  XNOR U16432 ( .A(b[3]), .B(n17008), .Z(n16153) );
  NANDN U16433 ( .A(n19521), .B(n16153), .Z(n16098) );
  AND U16434 ( .A(n16099), .B(n16098), .Z(n16179) );
  XNOR U16435 ( .A(n16178), .B(n16179), .Z(n16180) );
  XOR U16436 ( .A(n16181), .B(n16180), .Z(n16157) );
  XOR U16437 ( .A(n16156), .B(n16157), .Z(n16158) );
  XNOR U16438 ( .A(n16159), .B(n16158), .Z(n16129) );
  NAND U16439 ( .A(n16101), .B(n16100), .Z(n16105) );
  NAND U16440 ( .A(n16103), .B(n16102), .Z(n16104) );
  NAND U16441 ( .A(n16105), .B(n16104), .Z(n16130) );
  XOR U16442 ( .A(n16129), .B(n16130), .Z(n16132) );
  XNOR U16443 ( .A(n16131), .B(n16132), .Z(n16190) );
  NANDN U16444 ( .A(n16107), .B(n16106), .Z(n16111) );
  NAND U16445 ( .A(n16109), .B(n16108), .Z(n16110) );
  NAND U16446 ( .A(n16111), .B(n16110), .Z(n16191) );
  XNOR U16447 ( .A(n16190), .B(n16191), .Z(n16192) );
  XOR U16448 ( .A(n16193), .B(n16192), .Z(n16123) );
  NANDN U16449 ( .A(n16113), .B(n16112), .Z(n16117) );
  NANDN U16450 ( .A(n16115), .B(n16114), .Z(n16116) );
  NAND U16451 ( .A(n16117), .B(n16116), .Z(n16124) );
  XNOR U16452 ( .A(n16123), .B(n16124), .Z(n16125) );
  XNOR U16453 ( .A(n16126), .B(n16125), .Z(n16196) );
  XNOR U16454 ( .A(n16196), .B(sreg[453]), .Z(n16198) );
  NAND U16455 ( .A(n16118), .B(sreg[452]), .Z(n16122) );
  OR U16456 ( .A(n16120), .B(n16119), .Z(n16121) );
  AND U16457 ( .A(n16122), .B(n16121), .Z(n16197) );
  XOR U16458 ( .A(n16198), .B(n16197), .Z(c[453]) );
  NANDN U16459 ( .A(n16124), .B(n16123), .Z(n16128) );
  NAND U16460 ( .A(n16126), .B(n16125), .Z(n16127) );
  NAND U16461 ( .A(n16128), .B(n16127), .Z(n16204) );
  NANDN U16462 ( .A(n16130), .B(n16129), .Z(n16134) );
  OR U16463 ( .A(n16132), .B(n16131), .Z(n16133) );
  NAND U16464 ( .A(n16134), .B(n16133), .Z(n16271) );
  NANDN U16465 ( .A(n16136), .B(n16135), .Z(n16140) );
  OR U16466 ( .A(n16138), .B(n16137), .Z(n16139) );
  NAND U16467 ( .A(n16140), .B(n16139), .Z(n16259) );
  NAND U16468 ( .A(b[0]), .B(a[214]), .Z(n16141) );
  XNOR U16469 ( .A(b[1]), .B(n16141), .Z(n16143) );
  NAND U16470 ( .A(a[213]), .B(n98), .Z(n16142) );
  AND U16471 ( .A(n16143), .B(n16142), .Z(n16235) );
  XNOR U16472 ( .A(n20154), .B(n16294), .Z(n16244) );
  OR U16473 ( .A(n16244), .B(n20057), .Z(n16146) );
  NANDN U16474 ( .A(n16144), .B(n20098), .Z(n16145) );
  AND U16475 ( .A(n16146), .B(n16145), .Z(n16236) );
  XOR U16476 ( .A(n16235), .B(n16236), .Z(n16238) );
  NAND U16477 ( .A(a[198]), .B(b[15]), .Z(n16237) );
  XOR U16478 ( .A(n16238), .B(n16237), .Z(n16256) );
  NAND U16479 ( .A(n19722), .B(n16147), .Z(n16149) );
  XNOR U16480 ( .A(b[5]), .B(n16918), .Z(n16247) );
  NANDN U16481 ( .A(n19640), .B(n16247), .Z(n16148) );
  NAND U16482 ( .A(n16149), .B(n16148), .Z(n16232) );
  XNOR U16483 ( .A(n19714), .B(n16762), .Z(n16250) );
  NANDN U16484 ( .A(n16250), .B(n19766), .Z(n16152) );
  NANDN U16485 ( .A(n16150), .B(n19767), .Z(n16151) );
  NAND U16486 ( .A(n16152), .B(n16151), .Z(n16229) );
  NAND U16487 ( .A(n19554), .B(n16153), .Z(n16155) );
  IV U16488 ( .A(a[212]), .Z(n17074) );
  XNOR U16489 ( .A(b[3]), .B(n17074), .Z(n16253) );
  NANDN U16490 ( .A(n19521), .B(n16253), .Z(n16154) );
  AND U16491 ( .A(n16155), .B(n16154), .Z(n16230) );
  XNOR U16492 ( .A(n16229), .B(n16230), .Z(n16231) );
  XOR U16493 ( .A(n16232), .B(n16231), .Z(n16257) );
  XOR U16494 ( .A(n16256), .B(n16257), .Z(n16258) );
  XNOR U16495 ( .A(n16259), .B(n16258), .Z(n16207) );
  NAND U16496 ( .A(n16157), .B(n16156), .Z(n16161) );
  NAND U16497 ( .A(n16159), .B(n16158), .Z(n16160) );
  NAND U16498 ( .A(n16161), .B(n16160), .Z(n16208) );
  XOR U16499 ( .A(n16207), .B(n16208), .Z(n16210) );
  XNOR U16500 ( .A(n20052), .B(n16477), .Z(n16213) );
  OR U16501 ( .A(n16213), .B(n20020), .Z(n16164) );
  NANDN U16502 ( .A(n16162), .B(n19960), .Z(n16163) );
  NAND U16503 ( .A(n16164), .B(n16163), .Z(n16226) );
  XNOR U16504 ( .A(n102), .B(n16165), .Z(n16217) );
  OR U16505 ( .A(n16217), .B(n20121), .Z(n16168) );
  NANDN U16506 ( .A(n16166), .B(n20122), .Z(n16167) );
  NAND U16507 ( .A(n16168), .B(n16167), .Z(n16223) );
  XNOR U16508 ( .A(n19975), .B(n16606), .Z(n16220) );
  NANDN U16509 ( .A(n16220), .B(n19883), .Z(n16171) );
  NANDN U16510 ( .A(n16169), .B(n19937), .Z(n16170) );
  AND U16511 ( .A(n16171), .B(n16170), .Z(n16224) );
  XNOR U16512 ( .A(n16223), .B(n16224), .Z(n16225) );
  XNOR U16513 ( .A(n16226), .B(n16225), .Z(n16262) );
  NANDN U16514 ( .A(n16173), .B(n16172), .Z(n16177) );
  NAND U16515 ( .A(n16175), .B(n16174), .Z(n16176) );
  NAND U16516 ( .A(n16177), .B(n16176), .Z(n16263) );
  XNOR U16517 ( .A(n16262), .B(n16263), .Z(n16264) );
  NANDN U16518 ( .A(n16179), .B(n16178), .Z(n16183) );
  NAND U16519 ( .A(n16181), .B(n16180), .Z(n16182) );
  AND U16520 ( .A(n16183), .B(n16182), .Z(n16265) );
  XNOR U16521 ( .A(n16264), .B(n16265), .Z(n16209) );
  XNOR U16522 ( .A(n16210), .B(n16209), .Z(n16268) );
  NANDN U16523 ( .A(n16185), .B(n16184), .Z(n16189) );
  NAND U16524 ( .A(n16187), .B(n16186), .Z(n16188) );
  NAND U16525 ( .A(n16189), .B(n16188), .Z(n16269) );
  XNOR U16526 ( .A(n16268), .B(n16269), .Z(n16270) );
  XOR U16527 ( .A(n16271), .B(n16270), .Z(n16201) );
  NANDN U16528 ( .A(n16191), .B(n16190), .Z(n16195) );
  NANDN U16529 ( .A(n16193), .B(n16192), .Z(n16194) );
  NAND U16530 ( .A(n16195), .B(n16194), .Z(n16202) );
  XNOR U16531 ( .A(n16201), .B(n16202), .Z(n16203) );
  XNOR U16532 ( .A(n16204), .B(n16203), .Z(n16274) );
  XNOR U16533 ( .A(n16274), .B(sreg[454]), .Z(n16276) );
  NAND U16534 ( .A(n16196), .B(sreg[453]), .Z(n16200) );
  OR U16535 ( .A(n16198), .B(n16197), .Z(n16199) );
  AND U16536 ( .A(n16200), .B(n16199), .Z(n16275) );
  XOR U16537 ( .A(n16276), .B(n16275), .Z(c[454]) );
  NANDN U16538 ( .A(n16202), .B(n16201), .Z(n16206) );
  NAND U16539 ( .A(n16204), .B(n16203), .Z(n16205) );
  NAND U16540 ( .A(n16206), .B(n16205), .Z(n16282) );
  NANDN U16541 ( .A(n16208), .B(n16207), .Z(n16212) );
  OR U16542 ( .A(n16210), .B(n16209), .Z(n16211) );
  NAND U16543 ( .A(n16212), .B(n16211), .Z(n16349) );
  XNOR U16544 ( .A(n20052), .B(n16555), .Z(n16291) );
  OR U16545 ( .A(n16291), .B(n20020), .Z(n16215) );
  NANDN U16546 ( .A(n16213), .B(n19960), .Z(n16214) );
  NAND U16547 ( .A(n16215), .B(n16214), .Z(n16304) );
  XNOR U16548 ( .A(n102), .B(n16216), .Z(n16295) );
  OR U16549 ( .A(n16295), .B(n20121), .Z(n16219) );
  NANDN U16550 ( .A(n16217), .B(n20122), .Z(n16218) );
  NAND U16551 ( .A(n16219), .B(n16218), .Z(n16301) );
  XNOR U16552 ( .A(n19975), .B(n16684), .Z(n16298) );
  NANDN U16553 ( .A(n16298), .B(n19883), .Z(n16222) );
  NANDN U16554 ( .A(n16220), .B(n19937), .Z(n16221) );
  AND U16555 ( .A(n16222), .B(n16221), .Z(n16302) );
  XNOR U16556 ( .A(n16301), .B(n16302), .Z(n16303) );
  XNOR U16557 ( .A(n16304), .B(n16303), .Z(n16340) );
  NANDN U16558 ( .A(n16224), .B(n16223), .Z(n16228) );
  NAND U16559 ( .A(n16226), .B(n16225), .Z(n16227) );
  NAND U16560 ( .A(n16228), .B(n16227), .Z(n16341) );
  XNOR U16561 ( .A(n16340), .B(n16341), .Z(n16342) );
  NANDN U16562 ( .A(n16230), .B(n16229), .Z(n16234) );
  NAND U16563 ( .A(n16232), .B(n16231), .Z(n16233) );
  AND U16564 ( .A(n16234), .B(n16233), .Z(n16343) );
  XNOR U16565 ( .A(n16342), .B(n16343), .Z(n16287) );
  NANDN U16566 ( .A(n16236), .B(n16235), .Z(n16240) );
  OR U16567 ( .A(n16238), .B(n16237), .Z(n16239) );
  NAND U16568 ( .A(n16240), .B(n16239), .Z(n16337) );
  NAND U16569 ( .A(b[0]), .B(a[215]), .Z(n16241) );
  XNOR U16570 ( .A(b[1]), .B(n16241), .Z(n16243) );
  NAND U16571 ( .A(a[214]), .B(n98), .Z(n16242) );
  AND U16572 ( .A(n16243), .B(n16242), .Z(n16313) );
  XNOR U16573 ( .A(n20154), .B(n16399), .Z(n16322) );
  OR U16574 ( .A(n16322), .B(n20057), .Z(n16246) );
  NANDN U16575 ( .A(n16244), .B(n20098), .Z(n16245) );
  AND U16576 ( .A(n16246), .B(n16245), .Z(n16314) );
  XOR U16577 ( .A(n16313), .B(n16314), .Z(n16316) );
  NAND U16578 ( .A(a[199]), .B(b[15]), .Z(n16315) );
  XOR U16579 ( .A(n16316), .B(n16315), .Z(n16334) );
  NAND U16580 ( .A(n19722), .B(n16247), .Z(n16249) );
  XNOR U16581 ( .A(b[5]), .B(n17008), .Z(n16325) );
  NANDN U16582 ( .A(n19640), .B(n16325), .Z(n16248) );
  NAND U16583 ( .A(n16249), .B(n16248), .Z(n16310) );
  XNOR U16584 ( .A(n19714), .B(n16867), .Z(n16328) );
  NANDN U16585 ( .A(n16328), .B(n19766), .Z(n16252) );
  NANDN U16586 ( .A(n16250), .B(n19767), .Z(n16251) );
  NAND U16587 ( .A(n16252), .B(n16251), .Z(n16307) );
  NAND U16588 ( .A(n19554), .B(n16253), .Z(n16255) );
  IV U16589 ( .A(a[213]), .Z(n17152) );
  XNOR U16590 ( .A(b[3]), .B(n17152), .Z(n16331) );
  NANDN U16591 ( .A(n19521), .B(n16331), .Z(n16254) );
  AND U16592 ( .A(n16255), .B(n16254), .Z(n16308) );
  XNOR U16593 ( .A(n16307), .B(n16308), .Z(n16309) );
  XOR U16594 ( .A(n16310), .B(n16309), .Z(n16335) );
  XOR U16595 ( .A(n16334), .B(n16335), .Z(n16336) );
  XNOR U16596 ( .A(n16337), .B(n16336), .Z(n16285) );
  NAND U16597 ( .A(n16257), .B(n16256), .Z(n16261) );
  NAND U16598 ( .A(n16259), .B(n16258), .Z(n16260) );
  NAND U16599 ( .A(n16261), .B(n16260), .Z(n16286) );
  XOR U16600 ( .A(n16285), .B(n16286), .Z(n16288) );
  XNOR U16601 ( .A(n16287), .B(n16288), .Z(n16346) );
  NANDN U16602 ( .A(n16263), .B(n16262), .Z(n16267) );
  NAND U16603 ( .A(n16265), .B(n16264), .Z(n16266) );
  NAND U16604 ( .A(n16267), .B(n16266), .Z(n16347) );
  XNOR U16605 ( .A(n16346), .B(n16347), .Z(n16348) );
  XOR U16606 ( .A(n16349), .B(n16348), .Z(n16279) );
  NANDN U16607 ( .A(n16269), .B(n16268), .Z(n16273) );
  NANDN U16608 ( .A(n16271), .B(n16270), .Z(n16272) );
  NAND U16609 ( .A(n16273), .B(n16272), .Z(n16280) );
  XNOR U16610 ( .A(n16279), .B(n16280), .Z(n16281) );
  XNOR U16611 ( .A(n16282), .B(n16281), .Z(n16352) );
  XNOR U16612 ( .A(n16352), .B(sreg[455]), .Z(n16354) );
  NAND U16613 ( .A(n16274), .B(sreg[454]), .Z(n16278) );
  OR U16614 ( .A(n16276), .B(n16275), .Z(n16277) );
  AND U16615 ( .A(n16278), .B(n16277), .Z(n16353) );
  XOR U16616 ( .A(n16354), .B(n16353), .Z(c[455]) );
  NANDN U16617 ( .A(n16280), .B(n16279), .Z(n16284) );
  NAND U16618 ( .A(n16282), .B(n16281), .Z(n16283) );
  NAND U16619 ( .A(n16284), .B(n16283), .Z(n16360) );
  NANDN U16620 ( .A(n16286), .B(n16285), .Z(n16290) );
  OR U16621 ( .A(n16288), .B(n16287), .Z(n16289) );
  NAND U16622 ( .A(n16290), .B(n16289), .Z(n16427) );
  XNOR U16623 ( .A(n20052), .B(n16606), .Z(n16396) );
  OR U16624 ( .A(n16396), .B(n20020), .Z(n16293) );
  NANDN U16625 ( .A(n16291), .B(n19960), .Z(n16292) );
  NAND U16626 ( .A(n16293), .B(n16292), .Z(n16409) );
  XNOR U16627 ( .A(n102), .B(n16294), .Z(n16400) );
  OR U16628 ( .A(n16400), .B(n20121), .Z(n16297) );
  NANDN U16629 ( .A(n16295), .B(n20122), .Z(n16296) );
  NAND U16630 ( .A(n16297), .B(n16296), .Z(n16406) );
  XNOR U16631 ( .A(n19975), .B(n16762), .Z(n16403) );
  NANDN U16632 ( .A(n16403), .B(n19883), .Z(n16300) );
  NANDN U16633 ( .A(n16298), .B(n19937), .Z(n16299) );
  AND U16634 ( .A(n16300), .B(n16299), .Z(n16407) );
  XNOR U16635 ( .A(n16406), .B(n16407), .Z(n16408) );
  XNOR U16636 ( .A(n16409), .B(n16408), .Z(n16418) );
  NANDN U16637 ( .A(n16302), .B(n16301), .Z(n16306) );
  NAND U16638 ( .A(n16304), .B(n16303), .Z(n16305) );
  NAND U16639 ( .A(n16306), .B(n16305), .Z(n16419) );
  XNOR U16640 ( .A(n16418), .B(n16419), .Z(n16420) );
  NANDN U16641 ( .A(n16308), .B(n16307), .Z(n16312) );
  NAND U16642 ( .A(n16310), .B(n16309), .Z(n16311) );
  AND U16643 ( .A(n16312), .B(n16311), .Z(n16421) );
  XNOR U16644 ( .A(n16420), .B(n16421), .Z(n16365) );
  NANDN U16645 ( .A(n16314), .B(n16313), .Z(n16318) );
  OR U16646 ( .A(n16316), .B(n16315), .Z(n16317) );
  NAND U16647 ( .A(n16318), .B(n16317), .Z(n16393) );
  NAND U16648 ( .A(b[0]), .B(a[216]), .Z(n16319) );
  XNOR U16649 ( .A(b[1]), .B(n16319), .Z(n16321) );
  NAND U16650 ( .A(a[215]), .B(n98), .Z(n16320) );
  AND U16651 ( .A(n16321), .B(n16320), .Z(n16369) );
  XNOR U16652 ( .A(n20154), .B(n16477), .Z(n16378) );
  OR U16653 ( .A(n16378), .B(n20057), .Z(n16324) );
  NANDN U16654 ( .A(n16322), .B(n20098), .Z(n16323) );
  AND U16655 ( .A(n16324), .B(n16323), .Z(n16370) );
  XOR U16656 ( .A(n16369), .B(n16370), .Z(n16372) );
  NAND U16657 ( .A(a[200]), .B(b[15]), .Z(n16371) );
  XOR U16658 ( .A(n16372), .B(n16371), .Z(n16390) );
  NAND U16659 ( .A(n19722), .B(n16325), .Z(n16327) );
  XNOR U16660 ( .A(b[5]), .B(n17074), .Z(n16381) );
  NANDN U16661 ( .A(n19640), .B(n16381), .Z(n16326) );
  NAND U16662 ( .A(n16327), .B(n16326), .Z(n16415) );
  XNOR U16663 ( .A(n19714), .B(n16918), .Z(n16384) );
  NANDN U16664 ( .A(n16384), .B(n19766), .Z(n16330) );
  NANDN U16665 ( .A(n16328), .B(n19767), .Z(n16329) );
  NAND U16666 ( .A(n16330), .B(n16329), .Z(n16412) );
  NAND U16667 ( .A(n19554), .B(n16331), .Z(n16333) );
  IV U16668 ( .A(a[214]), .Z(n17257) );
  XNOR U16669 ( .A(b[3]), .B(n17257), .Z(n16387) );
  NANDN U16670 ( .A(n19521), .B(n16387), .Z(n16332) );
  AND U16671 ( .A(n16333), .B(n16332), .Z(n16413) );
  XNOR U16672 ( .A(n16412), .B(n16413), .Z(n16414) );
  XOR U16673 ( .A(n16415), .B(n16414), .Z(n16391) );
  XOR U16674 ( .A(n16390), .B(n16391), .Z(n16392) );
  XNOR U16675 ( .A(n16393), .B(n16392), .Z(n16363) );
  NAND U16676 ( .A(n16335), .B(n16334), .Z(n16339) );
  NAND U16677 ( .A(n16337), .B(n16336), .Z(n16338) );
  NAND U16678 ( .A(n16339), .B(n16338), .Z(n16364) );
  XOR U16679 ( .A(n16363), .B(n16364), .Z(n16366) );
  XNOR U16680 ( .A(n16365), .B(n16366), .Z(n16424) );
  NANDN U16681 ( .A(n16341), .B(n16340), .Z(n16345) );
  NAND U16682 ( .A(n16343), .B(n16342), .Z(n16344) );
  NAND U16683 ( .A(n16345), .B(n16344), .Z(n16425) );
  XNOR U16684 ( .A(n16424), .B(n16425), .Z(n16426) );
  XOR U16685 ( .A(n16427), .B(n16426), .Z(n16357) );
  NANDN U16686 ( .A(n16347), .B(n16346), .Z(n16351) );
  NANDN U16687 ( .A(n16349), .B(n16348), .Z(n16350) );
  NAND U16688 ( .A(n16351), .B(n16350), .Z(n16358) );
  XNOR U16689 ( .A(n16357), .B(n16358), .Z(n16359) );
  XNOR U16690 ( .A(n16360), .B(n16359), .Z(n16430) );
  XNOR U16691 ( .A(n16430), .B(sreg[456]), .Z(n16432) );
  NAND U16692 ( .A(n16352), .B(sreg[455]), .Z(n16356) );
  OR U16693 ( .A(n16354), .B(n16353), .Z(n16355) );
  AND U16694 ( .A(n16356), .B(n16355), .Z(n16431) );
  XOR U16695 ( .A(n16432), .B(n16431), .Z(c[456]) );
  NANDN U16696 ( .A(n16358), .B(n16357), .Z(n16362) );
  NAND U16697 ( .A(n16360), .B(n16359), .Z(n16361) );
  NAND U16698 ( .A(n16362), .B(n16361), .Z(n16438) );
  NANDN U16699 ( .A(n16364), .B(n16363), .Z(n16368) );
  OR U16700 ( .A(n16366), .B(n16365), .Z(n16367) );
  NAND U16701 ( .A(n16368), .B(n16367), .Z(n16505) );
  NANDN U16702 ( .A(n16370), .B(n16369), .Z(n16374) );
  OR U16703 ( .A(n16372), .B(n16371), .Z(n16373) );
  NAND U16704 ( .A(n16374), .B(n16373), .Z(n16471) );
  NAND U16705 ( .A(b[0]), .B(a[217]), .Z(n16375) );
  XNOR U16706 ( .A(b[1]), .B(n16375), .Z(n16377) );
  NAND U16707 ( .A(a[216]), .B(n98), .Z(n16376) );
  AND U16708 ( .A(n16377), .B(n16376), .Z(n16447) );
  XNOR U16709 ( .A(n20154), .B(n16555), .Z(n16453) );
  OR U16710 ( .A(n16453), .B(n20057), .Z(n16380) );
  NANDN U16711 ( .A(n16378), .B(n20098), .Z(n16379) );
  AND U16712 ( .A(n16380), .B(n16379), .Z(n16448) );
  XOR U16713 ( .A(n16447), .B(n16448), .Z(n16450) );
  NAND U16714 ( .A(a[201]), .B(b[15]), .Z(n16449) );
  XOR U16715 ( .A(n16450), .B(n16449), .Z(n16468) );
  NAND U16716 ( .A(n19722), .B(n16381), .Z(n16383) );
  XNOR U16717 ( .A(b[5]), .B(n17152), .Z(n16459) );
  NANDN U16718 ( .A(n19640), .B(n16459), .Z(n16382) );
  NAND U16719 ( .A(n16383), .B(n16382), .Z(n16493) );
  XNOR U16720 ( .A(n19714), .B(n17008), .Z(n16462) );
  NANDN U16721 ( .A(n16462), .B(n19766), .Z(n16386) );
  NANDN U16722 ( .A(n16384), .B(n19767), .Z(n16385) );
  NAND U16723 ( .A(n16386), .B(n16385), .Z(n16490) );
  NAND U16724 ( .A(n19554), .B(n16387), .Z(n16389) );
  IV U16725 ( .A(a[215]), .Z(n17308) );
  XNOR U16726 ( .A(b[3]), .B(n17308), .Z(n16465) );
  NANDN U16727 ( .A(n19521), .B(n16465), .Z(n16388) );
  AND U16728 ( .A(n16389), .B(n16388), .Z(n16491) );
  XNOR U16729 ( .A(n16490), .B(n16491), .Z(n16492) );
  XOR U16730 ( .A(n16493), .B(n16492), .Z(n16469) );
  XOR U16731 ( .A(n16468), .B(n16469), .Z(n16470) );
  XNOR U16732 ( .A(n16471), .B(n16470), .Z(n16441) );
  NAND U16733 ( .A(n16391), .B(n16390), .Z(n16395) );
  NAND U16734 ( .A(n16393), .B(n16392), .Z(n16394) );
  NAND U16735 ( .A(n16395), .B(n16394), .Z(n16442) );
  XOR U16736 ( .A(n16441), .B(n16442), .Z(n16444) );
  XNOR U16737 ( .A(n20052), .B(n16684), .Z(n16474) );
  OR U16738 ( .A(n16474), .B(n20020), .Z(n16398) );
  NANDN U16739 ( .A(n16396), .B(n19960), .Z(n16397) );
  NAND U16740 ( .A(n16398), .B(n16397), .Z(n16487) );
  XNOR U16741 ( .A(n102), .B(n16399), .Z(n16478) );
  OR U16742 ( .A(n16478), .B(n20121), .Z(n16402) );
  NANDN U16743 ( .A(n16400), .B(n20122), .Z(n16401) );
  NAND U16744 ( .A(n16402), .B(n16401), .Z(n16484) );
  XNOR U16745 ( .A(n19975), .B(n16867), .Z(n16481) );
  NANDN U16746 ( .A(n16481), .B(n19883), .Z(n16405) );
  NANDN U16747 ( .A(n16403), .B(n19937), .Z(n16404) );
  AND U16748 ( .A(n16405), .B(n16404), .Z(n16485) );
  XNOR U16749 ( .A(n16484), .B(n16485), .Z(n16486) );
  XNOR U16750 ( .A(n16487), .B(n16486), .Z(n16496) );
  NANDN U16751 ( .A(n16407), .B(n16406), .Z(n16411) );
  NAND U16752 ( .A(n16409), .B(n16408), .Z(n16410) );
  NAND U16753 ( .A(n16411), .B(n16410), .Z(n16497) );
  XNOR U16754 ( .A(n16496), .B(n16497), .Z(n16498) );
  NANDN U16755 ( .A(n16413), .B(n16412), .Z(n16417) );
  NAND U16756 ( .A(n16415), .B(n16414), .Z(n16416) );
  AND U16757 ( .A(n16417), .B(n16416), .Z(n16499) );
  XNOR U16758 ( .A(n16498), .B(n16499), .Z(n16443) );
  XNOR U16759 ( .A(n16444), .B(n16443), .Z(n16502) );
  NANDN U16760 ( .A(n16419), .B(n16418), .Z(n16423) );
  NAND U16761 ( .A(n16421), .B(n16420), .Z(n16422) );
  NAND U16762 ( .A(n16423), .B(n16422), .Z(n16503) );
  XNOR U16763 ( .A(n16502), .B(n16503), .Z(n16504) );
  XOR U16764 ( .A(n16505), .B(n16504), .Z(n16435) );
  NANDN U16765 ( .A(n16425), .B(n16424), .Z(n16429) );
  NANDN U16766 ( .A(n16427), .B(n16426), .Z(n16428) );
  NAND U16767 ( .A(n16429), .B(n16428), .Z(n16436) );
  XNOR U16768 ( .A(n16435), .B(n16436), .Z(n16437) );
  XNOR U16769 ( .A(n16438), .B(n16437), .Z(n16508) );
  XNOR U16770 ( .A(n16508), .B(sreg[457]), .Z(n16510) );
  NAND U16771 ( .A(n16430), .B(sreg[456]), .Z(n16434) );
  OR U16772 ( .A(n16432), .B(n16431), .Z(n16433) );
  AND U16773 ( .A(n16434), .B(n16433), .Z(n16509) );
  XOR U16774 ( .A(n16510), .B(n16509), .Z(c[457]) );
  NANDN U16775 ( .A(n16436), .B(n16435), .Z(n16440) );
  NAND U16776 ( .A(n16438), .B(n16437), .Z(n16439) );
  NAND U16777 ( .A(n16440), .B(n16439), .Z(n16516) );
  NANDN U16778 ( .A(n16442), .B(n16441), .Z(n16446) );
  OR U16779 ( .A(n16444), .B(n16443), .Z(n16445) );
  NAND U16780 ( .A(n16446), .B(n16445), .Z(n16583) );
  NANDN U16781 ( .A(n16448), .B(n16447), .Z(n16452) );
  OR U16782 ( .A(n16450), .B(n16449), .Z(n16451) );
  NAND U16783 ( .A(n16452), .B(n16451), .Z(n16549) );
  XNOR U16784 ( .A(n20154), .B(n16606), .Z(n16534) );
  OR U16785 ( .A(n16534), .B(n20057), .Z(n16455) );
  NANDN U16786 ( .A(n16453), .B(n20098), .Z(n16454) );
  AND U16787 ( .A(n16455), .B(n16454), .Z(n16526) );
  NAND U16788 ( .A(b[0]), .B(a[218]), .Z(n16456) );
  XNOR U16789 ( .A(b[1]), .B(n16456), .Z(n16458) );
  NAND U16790 ( .A(a[217]), .B(n98), .Z(n16457) );
  AND U16791 ( .A(n16458), .B(n16457), .Z(n16525) );
  XOR U16792 ( .A(n16526), .B(n16525), .Z(n16528) );
  NAND U16793 ( .A(a[202]), .B(b[15]), .Z(n16527) );
  XOR U16794 ( .A(n16528), .B(n16527), .Z(n16546) );
  NAND U16795 ( .A(n19722), .B(n16459), .Z(n16461) );
  XNOR U16796 ( .A(b[5]), .B(n17257), .Z(n16537) );
  NANDN U16797 ( .A(n19640), .B(n16537), .Z(n16460) );
  NAND U16798 ( .A(n16461), .B(n16460), .Z(n16571) );
  XNOR U16799 ( .A(n19714), .B(n17074), .Z(n16540) );
  NANDN U16800 ( .A(n16540), .B(n19766), .Z(n16464) );
  NANDN U16801 ( .A(n16462), .B(n19767), .Z(n16463) );
  NAND U16802 ( .A(n16464), .B(n16463), .Z(n16568) );
  NAND U16803 ( .A(n19554), .B(n16465), .Z(n16467) );
  IV U16804 ( .A(a[216]), .Z(n17413) );
  XNOR U16805 ( .A(b[3]), .B(n17413), .Z(n16543) );
  NANDN U16806 ( .A(n19521), .B(n16543), .Z(n16466) );
  AND U16807 ( .A(n16467), .B(n16466), .Z(n16569) );
  XNOR U16808 ( .A(n16568), .B(n16569), .Z(n16570) );
  XOR U16809 ( .A(n16571), .B(n16570), .Z(n16547) );
  XOR U16810 ( .A(n16546), .B(n16547), .Z(n16548) );
  XNOR U16811 ( .A(n16549), .B(n16548), .Z(n16519) );
  NAND U16812 ( .A(n16469), .B(n16468), .Z(n16473) );
  NAND U16813 ( .A(n16471), .B(n16470), .Z(n16472) );
  NAND U16814 ( .A(n16473), .B(n16472), .Z(n16520) );
  XOR U16815 ( .A(n16519), .B(n16520), .Z(n16522) );
  XNOR U16816 ( .A(n20052), .B(n16762), .Z(n16552) );
  OR U16817 ( .A(n16552), .B(n20020), .Z(n16476) );
  NANDN U16818 ( .A(n16474), .B(n19960), .Z(n16475) );
  NAND U16819 ( .A(n16476), .B(n16475), .Z(n16565) );
  XNOR U16820 ( .A(n102), .B(n16477), .Z(n16556) );
  OR U16821 ( .A(n16556), .B(n20121), .Z(n16480) );
  NANDN U16822 ( .A(n16478), .B(n20122), .Z(n16479) );
  NAND U16823 ( .A(n16480), .B(n16479), .Z(n16562) );
  XNOR U16824 ( .A(n19975), .B(n16918), .Z(n16559) );
  NANDN U16825 ( .A(n16559), .B(n19883), .Z(n16483) );
  NANDN U16826 ( .A(n16481), .B(n19937), .Z(n16482) );
  AND U16827 ( .A(n16483), .B(n16482), .Z(n16563) );
  XNOR U16828 ( .A(n16562), .B(n16563), .Z(n16564) );
  XNOR U16829 ( .A(n16565), .B(n16564), .Z(n16574) );
  NANDN U16830 ( .A(n16485), .B(n16484), .Z(n16489) );
  NAND U16831 ( .A(n16487), .B(n16486), .Z(n16488) );
  NAND U16832 ( .A(n16489), .B(n16488), .Z(n16575) );
  XNOR U16833 ( .A(n16574), .B(n16575), .Z(n16576) );
  NANDN U16834 ( .A(n16491), .B(n16490), .Z(n16495) );
  NAND U16835 ( .A(n16493), .B(n16492), .Z(n16494) );
  AND U16836 ( .A(n16495), .B(n16494), .Z(n16577) );
  XNOR U16837 ( .A(n16576), .B(n16577), .Z(n16521) );
  XNOR U16838 ( .A(n16522), .B(n16521), .Z(n16580) );
  NANDN U16839 ( .A(n16497), .B(n16496), .Z(n16501) );
  NAND U16840 ( .A(n16499), .B(n16498), .Z(n16500) );
  NAND U16841 ( .A(n16501), .B(n16500), .Z(n16581) );
  XNOR U16842 ( .A(n16580), .B(n16581), .Z(n16582) );
  XOR U16843 ( .A(n16583), .B(n16582), .Z(n16513) );
  NANDN U16844 ( .A(n16503), .B(n16502), .Z(n16507) );
  NANDN U16845 ( .A(n16505), .B(n16504), .Z(n16506) );
  NAND U16846 ( .A(n16507), .B(n16506), .Z(n16514) );
  XNOR U16847 ( .A(n16513), .B(n16514), .Z(n16515) );
  XNOR U16848 ( .A(n16516), .B(n16515), .Z(n16586) );
  XNOR U16849 ( .A(n16586), .B(sreg[458]), .Z(n16588) );
  NAND U16850 ( .A(n16508), .B(sreg[457]), .Z(n16512) );
  OR U16851 ( .A(n16510), .B(n16509), .Z(n16511) );
  AND U16852 ( .A(n16512), .B(n16511), .Z(n16587) );
  XOR U16853 ( .A(n16588), .B(n16587), .Z(c[458]) );
  NANDN U16854 ( .A(n16514), .B(n16513), .Z(n16518) );
  NAND U16855 ( .A(n16516), .B(n16515), .Z(n16517) );
  NAND U16856 ( .A(n16518), .B(n16517), .Z(n16594) );
  NANDN U16857 ( .A(n16520), .B(n16519), .Z(n16524) );
  OR U16858 ( .A(n16522), .B(n16521), .Z(n16523) );
  NAND U16859 ( .A(n16524), .B(n16523), .Z(n16661) );
  NANDN U16860 ( .A(n16526), .B(n16525), .Z(n16530) );
  OR U16861 ( .A(n16528), .B(n16527), .Z(n16529) );
  NAND U16862 ( .A(n16530), .B(n16529), .Z(n16649) );
  NAND U16863 ( .A(b[0]), .B(a[219]), .Z(n16531) );
  XNOR U16864 ( .A(b[1]), .B(n16531), .Z(n16533) );
  NAND U16865 ( .A(a[218]), .B(n98), .Z(n16532) );
  AND U16866 ( .A(n16533), .B(n16532), .Z(n16625) );
  XNOR U16867 ( .A(n20154), .B(n16684), .Z(n16631) );
  OR U16868 ( .A(n16631), .B(n20057), .Z(n16536) );
  NANDN U16869 ( .A(n16534), .B(n20098), .Z(n16535) );
  AND U16870 ( .A(n16536), .B(n16535), .Z(n16626) );
  XOR U16871 ( .A(n16625), .B(n16626), .Z(n16628) );
  NAND U16872 ( .A(a[203]), .B(b[15]), .Z(n16627) );
  XOR U16873 ( .A(n16628), .B(n16627), .Z(n16646) );
  NAND U16874 ( .A(n19722), .B(n16537), .Z(n16539) );
  XNOR U16875 ( .A(b[5]), .B(n17308), .Z(n16637) );
  NANDN U16876 ( .A(n19640), .B(n16637), .Z(n16538) );
  NAND U16877 ( .A(n16539), .B(n16538), .Z(n16622) );
  XNOR U16878 ( .A(n19714), .B(n17152), .Z(n16640) );
  NANDN U16879 ( .A(n16640), .B(n19766), .Z(n16542) );
  NANDN U16880 ( .A(n16540), .B(n19767), .Z(n16541) );
  NAND U16881 ( .A(n16542), .B(n16541), .Z(n16619) );
  NAND U16882 ( .A(n19554), .B(n16543), .Z(n16545) );
  IV U16883 ( .A(a[217]), .Z(n17464) );
  XNOR U16884 ( .A(b[3]), .B(n17464), .Z(n16643) );
  NANDN U16885 ( .A(n19521), .B(n16643), .Z(n16544) );
  AND U16886 ( .A(n16545), .B(n16544), .Z(n16620) );
  XNOR U16887 ( .A(n16619), .B(n16620), .Z(n16621) );
  XOR U16888 ( .A(n16622), .B(n16621), .Z(n16647) );
  XOR U16889 ( .A(n16646), .B(n16647), .Z(n16648) );
  XNOR U16890 ( .A(n16649), .B(n16648), .Z(n16597) );
  NAND U16891 ( .A(n16547), .B(n16546), .Z(n16551) );
  NAND U16892 ( .A(n16549), .B(n16548), .Z(n16550) );
  NAND U16893 ( .A(n16551), .B(n16550), .Z(n16598) );
  XOR U16894 ( .A(n16597), .B(n16598), .Z(n16600) );
  XNOR U16895 ( .A(n20052), .B(n16867), .Z(n16603) );
  OR U16896 ( .A(n16603), .B(n20020), .Z(n16554) );
  NANDN U16897 ( .A(n16552), .B(n19960), .Z(n16553) );
  NAND U16898 ( .A(n16554), .B(n16553), .Z(n16616) );
  XNOR U16899 ( .A(n102), .B(n16555), .Z(n16607) );
  OR U16900 ( .A(n16607), .B(n20121), .Z(n16558) );
  NANDN U16901 ( .A(n16556), .B(n20122), .Z(n16557) );
  NAND U16902 ( .A(n16558), .B(n16557), .Z(n16613) );
  XNOR U16903 ( .A(n19975), .B(n17008), .Z(n16610) );
  NANDN U16904 ( .A(n16610), .B(n19883), .Z(n16561) );
  NANDN U16905 ( .A(n16559), .B(n19937), .Z(n16560) );
  AND U16906 ( .A(n16561), .B(n16560), .Z(n16614) );
  XNOR U16907 ( .A(n16613), .B(n16614), .Z(n16615) );
  XNOR U16908 ( .A(n16616), .B(n16615), .Z(n16652) );
  NANDN U16909 ( .A(n16563), .B(n16562), .Z(n16567) );
  NAND U16910 ( .A(n16565), .B(n16564), .Z(n16566) );
  NAND U16911 ( .A(n16567), .B(n16566), .Z(n16653) );
  XNOR U16912 ( .A(n16652), .B(n16653), .Z(n16654) );
  NANDN U16913 ( .A(n16569), .B(n16568), .Z(n16573) );
  NAND U16914 ( .A(n16571), .B(n16570), .Z(n16572) );
  AND U16915 ( .A(n16573), .B(n16572), .Z(n16655) );
  XNOR U16916 ( .A(n16654), .B(n16655), .Z(n16599) );
  XNOR U16917 ( .A(n16600), .B(n16599), .Z(n16658) );
  NANDN U16918 ( .A(n16575), .B(n16574), .Z(n16579) );
  NAND U16919 ( .A(n16577), .B(n16576), .Z(n16578) );
  NAND U16920 ( .A(n16579), .B(n16578), .Z(n16659) );
  XNOR U16921 ( .A(n16658), .B(n16659), .Z(n16660) );
  XOR U16922 ( .A(n16661), .B(n16660), .Z(n16591) );
  NANDN U16923 ( .A(n16581), .B(n16580), .Z(n16585) );
  NANDN U16924 ( .A(n16583), .B(n16582), .Z(n16584) );
  NAND U16925 ( .A(n16585), .B(n16584), .Z(n16592) );
  XNOR U16926 ( .A(n16591), .B(n16592), .Z(n16593) );
  XNOR U16927 ( .A(n16594), .B(n16593), .Z(n16664) );
  XNOR U16928 ( .A(n16664), .B(sreg[459]), .Z(n16666) );
  NAND U16929 ( .A(n16586), .B(sreg[458]), .Z(n16590) );
  OR U16930 ( .A(n16588), .B(n16587), .Z(n16589) );
  AND U16931 ( .A(n16590), .B(n16589), .Z(n16665) );
  XOR U16932 ( .A(n16666), .B(n16665), .Z(c[459]) );
  NANDN U16933 ( .A(n16592), .B(n16591), .Z(n16596) );
  NAND U16934 ( .A(n16594), .B(n16593), .Z(n16595) );
  NAND U16935 ( .A(n16596), .B(n16595), .Z(n16672) );
  NANDN U16936 ( .A(n16598), .B(n16597), .Z(n16602) );
  OR U16937 ( .A(n16600), .B(n16599), .Z(n16601) );
  NAND U16938 ( .A(n16602), .B(n16601), .Z(n16739) );
  XNOR U16939 ( .A(n20052), .B(n16918), .Z(n16681) );
  OR U16940 ( .A(n16681), .B(n20020), .Z(n16605) );
  NANDN U16941 ( .A(n16603), .B(n19960), .Z(n16604) );
  NAND U16942 ( .A(n16605), .B(n16604), .Z(n16694) );
  XNOR U16943 ( .A(n102), .B(n16606), .Z(n16685) );
  OR U16944 ( .A(n16685), .B(n20121), .Z(n16609) );
  NANDN U16945 ( .A(n16607), .B(n20122), .Z(n16608) );
  NAND U16946 ( .A(n16609), .B(n16608), .Z(n16691) );
  XNOR U16947 ( .A(n19975), .B(n17074), .Z(n16688) );
  NANDN U16948 ( .A(n16688), .B(n19883), .Z(n16612) );
  NANDN U16949 ( .A(n16610), .B(n19937), .Z(n16611) );
  AND U16950 ( .A(n16612), .B(n16611), .Z(n16692) );
  XNOR U16951 ( .A(n16691), .B(n16692), .Z(n16693) );
  XNOR U16952 ( .A(n16694), .B(n16693), .Z(n16730) );
  NANDN U16953 ( .A(n16614), .B(n16613), .Z(n16618) );
  NAND U16954 ( .A(n16616), .B(n16615), .Z(n16617) );
  NAND U16955 ( .A(n16618), .B(n16617), .Z(n16731) );
  XNOR U16956 ( .A(n16730), .B(n16731), .Z(n16732) );
  NANDN U16957 ( .A(n16620), .B(n16619), .Z(n16624) );
  NAND U16958 ( .A(n16622), .B(n16621), .Z(n16623) );
  AND U16959 ( .A(n16624), .B(n16623), .Z(n16733) );
  XNOR U16960 ( .A(n16732), .B(n16733), .Z(n16677) );
  NANDN U16961 ( .A(n16626), .B(n16625), .Z(n16630) );
  OR U16962 ( .A(n16628), .B(n16627), .Z(n16629) );
  NAND U16963 ( .A(n16630), .B(n16629), .Z(n16727) );
  XNOR U16964 ( .A(n20154), .B(n16762), .Z(n16712) );
  OR U16965 ( .A(n16712), .B(n20057), .Z(n16633) );
  NANDN U16966 ( .A(n16631), .B(n20098), .Z(n16632) );
  AND U16967 ( .A(n16633), .B(n16632), .Z(n16704) );
  NAND U16968 ( .A(b[0]), .B(a[220]), .Z(n16634) );
  XNOR U16969 ( .A(b[1]), .B(n16634), .Z(n16636) );
  NAND U16970 ( .A(a[219]), .B(n98), .Z(n16635) );
  AND U16971 ( .A(n16636), .B(n16635), .Z(n16703) );
  XOR U16972 ( .A(n16704), .B(n16703), .Z(n16706) );
  NAND U16973 ( .A(a[204]), .B(b[15]), .Z(n16705) );
  XOR U16974 ( .A(n16706), .B(n16705), .Z(n16724) );
  NAND U16975 ( .A(n19722), .B(n16637), .Z(n16639) );
  XNOR U16976 ( .A(b[5]), .B(n17413), .Z(n16715) );
  NANDN U16977 ( .A(n19640), .B(n16715), .Z(n16638) );
  NAND U16978 ( .A(n16639), .B(n16638), .Z(n16700) );
  XNOR U16979 ( .A(n19714), .B(n17257), .Z(n16718) );
  NANDN U16980 ( .A(n16718), .B(n19766), .Z(n16642) );
  NANDN U16981 ( .A(n16640), .B(n19767), .Z(n16641) );
  NAND U16982 ( .A(n16642), .B(n16641), .Z(n16697) );
  NAND U16983 ( .A(n19554), .B(n16643), .Z(n16645) );
  IV U16984 ( .A(a[218]), .Z(n17542) );
  XNOR U16985 ( .A(b[3]), .B(n17542), .Z(n16721) );
  NANDN U16986 ( .A(n19521), .B(n16721), .Z(n16644) );
  AND U16987 ( .A(n16645), .B(n16644), .Z(n16698) );
  XNOR U16988 ( .A(n16697), .B(n16698), .Z(n16699) );
  XOR U16989 ( .A(n16700), .B(n16699), .Z(n16725) );
  XOR U16990 ( .A(n16724), .B(n16725), .Z(n16726) );
  XNOR U16991 ( .A(n16727), .B(n16726), .Z(n16675) );
  NAND U16992 ( .A(n16647), .B(n16646), .Z(n16651) );
  NAND U16993 ( .A(n16649), .B(n16648), .Z(n16650) );
  NAND U16994 ( .A(n16651), .B(n16650), .Z(n16676) );
  XOR U16995 ( .A(n16675), .B(n16676), .Z(n16678) );
  XNOR U16996 ( .A(n16677), .B(n16678), .Z(n16736) );
  NANDN U16997 ( .A(n16653), .B(n16652), .Z(n16657) );
  NAND U16998 ( .A(n16655), .B(n16654), .Z(n16656) );
  NAND U16999 ( .A(n16657), .B(n16656), .Z(n16737) );
  XNOR U17000 ( .A(n16736), .B(n16737), .Z(n16738) );
  XOR U17001 ( .A(n16739), .B(n16738), .Z(n16669) );
  NANDN U17002 ( .A(n16659), .B(n16658), .Z(n16663) );
  NANDN U17003 ( .A(n16661), .B(n16660), .Z(n16662) );
  NAND U17004 ( .A(n16663), .B(n16662), .Z(n16670) );
  XNOR U17005 ( .A(n16669), .B(n16670), .Z(n16671) );
  XNOR U17006 ( .A(n16672), .B(n16671), .Z(n16742) );
  XNOR U17007 ( .A(n16742), .B(sreg[460]), .Z(n16744) );
  NAND U17008 ( .A(n16664), .B(sreg[459]), .Z(n16668) );
  OR U17009 ( .A(n16666), .B(n16665), .Z(n16667) );
  AND U17010 ( .A(n16668), .B(n16667), .Z(n16743) );
  XOR U17011 ( .A(n16744), .B(n16743), .Z(c[460]) );
  NANDN U17012 ( .A(n16670), .B(n16669), .Z(n16674) );
  NAND U17013 ( .A(n16672), .B(n16671), .Z(n16673) );
  NAND U17014 ( .A(n16674), .B(n16673), .Z(n16750) );
  NANDN U17015 ( .A(n16676), .B(n16675), .Z(n16680) );
  OR U17016 ( .A(n16678), .B(n16677), .Z(n16679) );
  NAND U17017 ( .A(n16680), .B(n16679), .Z(n16817) );
  XNOR U17018 ( .A(n20052), .B(n17008), .Z(n16759) );
  OR U17019 ( .A(n16759), .B(n20020), .Z(n16683) );
  NANDN U17020 ( .A(n16681), .B(n19960), .Z(n16682) );
  NAND U17021 ( .A(n16683), .B(n16682), .Z(n16772) );
  XNOR U17022 ( .A(n102), .B(n16684), .Z(n16763) );
  OR U17023 ( .A(n16763), .B(n20121), .Z(n16687) );
  NANDN U17024 ( .A(n16685), .B(n20122), .Z(n16686) );
  NAND U17025 ( .A(n16687), .B(n16686), .Z(n16769) );
  XNOR U17026 ( .A(n19975), .B(n17152), .Z(n16766) );
  NANDN U17027 ( .A(n16766), .B(n19883), .Z(n16690) );
  NANDN U17028 ( .A(n16688), .B(n19937), .Z(n16689) );
  AND U17029 ( .A(n16690), .B(n16689), .Z(n16770) );
  XNOR U17030 ( .A(n16769), .B(n16770), .Z(n16771) );
  XNOR U17031 ( .A(n16772), .B(n16771), .Z(n16808) );
  NANDN U17032 ( .A(n16692), .B(n16691), .Z(n16696) );
  NAND U17033 ( .A(n16694), .B(n16693), .Z(n16695) );
  NAND U17034 ( .A(n16696), .B(n16695), .Z(n16809) );
  XNOR U17035 ( .A(n16808), .B(n16809), .Z(n16810) );
  NANDN U17036 ( .A(n16698), .B(n16697), .Z(n16702) );
  NAND U17037 ( .A(n16700), .B(n16699), .Z(n16701) );
  AND U17038 ( .A(n16702), .B(n16701), .Z(n16811) );
  XNOR U17039 ( .A(n16810), .B(n16811), .Z(n16755) );
  NANDN U17040 ( .A(n16704), .B(n16703), .Z(n16708) );
  OR U17041 ( .A(n16706), .B(n16705), .Z(n16707) );
  NAND U17042 ( .A(n16708), .B(n16707), .Z(n16805) );
  NAND U17043 ( .A(b[0]), .B(a[221]), .Z(n16709) );
  XNOR U17044 ( .A(b[1]), .B(n16709), .Z(n16711) );
  NAND U17045 ( .A(a[220]), .B(n98), .Z(n16710) );
  AND U17046 ( .A(n16711), .B(n16710), .Z(n16781) );
  XNOR U17047 ( .A(n20154), .B(n16867), .Z(n16790) );
  OR U17048 ( .A(n16790), .B(n20057), .Z(n16714) );
  NANDN U17049 ( .A(n16712), .B(n20098), .Z(n16713) );
  AND U17050 ( .A(n16714), .B(n16713), .Z(n16782) );
  XOR U17051 ( .A(n16781), .B(n16782), .Z(n16784) );
  NAND U17052 ( .A(a[205]), .B(b[15]), .Z(n16783) );
  XOR U17053 ( .A(n16784), .B(n16783), .Z(n16802) );
  NAND U17054 ( .A(n19722), .B(n16715), .Z(n16717) );
  XNOR U17055 ( .A(b[5]), .B(n17464), .Z(n16793) );
  NANDN U17056 ( .A(n19640), .B(n16793), .Z(n16716) );
  NAND U17057 ( .A(n16717), .B(n16716), .Z(n16778) );
  XNOR U17058 ( .A(n19714), .B(n17308), .Z(n16796) );
  NANDN U17059 ( .A(n16796), .B(n19766), .Z(n16720) );
  NANDN U17060 ( .A(n16718), .B(n19767), .Z(n16719) );
  NAND U17061 ( .A(n16720), .B(n16719), .Z(n16775) );
  NAND U17062 ( .A(n19554), .B(n16721), .Z(n16723) );
  IV U17063 ( .A(a[219]), .Z(n17620) );
  XNOR U17064 ( .A(b[3]), .B(n17620), .Z(n16799) );
  NANDN U17065 ( .A(n19521), .B(n16799), .Z(n16722) );
  AND U17066 ( .A(n16723), .B(n16722), .Z(n16776) );
  XNOR U17067 ( .A(n16775), .B(n16776), .Z(n16777) );
  XOR U17068 ( .A(n16778), .B(n16777), .Z(n16803) );
  XOR U17069 ( .A(n16802), .B(n16803), .Z(n16804) );
  XNOR U17070 ( .A(n16805), .B(n16804), .Z(n16753) );
  NAND U17071 ( .A(n16725), .B(n16724), .Z(n16729) );
  NAND U17072 ( .A(n16727), .B(n16726), .Z(n16728) );
  NAND U17073 ( .A(n16729), .B(n16728), .Z(n16754) );
  XOR U17074 ( .A(n16753), .B(n16754), .Z(n16756) );
  XNOR U17075 ( .A(n16755), .B(n16756), .Z(n16814) );
  NANDN U17076 ( .A(n16731), .B(n16730), .Z(n16735) );
  NAND U17077 ( .A(n16733), .B(n16732), .Z(n16734) );
  NAND U17078 ( .A(n16735), .B(n16734), .Z(n16815) );
  XNOR U17079 ( .A(n16814), .B(n16815), .Z(n16816) );
  XOR U17080 ( .A(n16817), .B(n16816), .Z(n16747) );
  NANDN U17081 ( .A(n16737), .B(n16736), .Z(n16741) );
  NANDN U17082 ( .A(n16739), .B(n16738), .Z(n16740) );
  NAND U17083 ( .A(n16741), .B(n16740), .Z(n16748) );
  XNOR U17084 ( .A(n16747), .B(n16748), .Z(n16749) );
  XNOR U17085 ( .A(n16750), .B(n16749), .Z(n16820) );
  XNOR U17086 ( .A(n16820), .B(sreg[461]), .Z(n16822) );
  NAND U17087 ( .A(n16742), .B(sreg[460]), .Z(n16746) );
  OR U17088 ( .A(n16744), .B(n16743), .Z(n16745) );
  AND U17089 ( .A(n16746), .B(n16745), .Z(n16821) );
  XOR U17090 ( .A(n16822), .B(n16821), .Z(c[461]) );
  NANDN U17091 ( .A(n16748), .B(n16747), .Z(n16752) );
  NAND U17092 ( .A(n16750), .B(n16749), .Z(n16751) );
  NAND U17093 ( .A(n16752), .B(n16751), .Z(n16828) );
  NANDN U17094 ( .A(n16754), .B(n16753), .Z(n16758) );
  OR U17095 ( .A(n16756), .B(n16755), .Z(n16757) );
  NAND U17096 ( .A(n16758), .B(n16757), .Z(n16895) );
  XNOR U17097 ( .A(n20052), .B(n17074), .Z(n16864) );
  OR U17098 ( .A(n16864), .B(n20020), .Z(n16761) );
  NANDN U17099 ( .A(n16759), .B(n19960), .Z(n16760) );
  NAND U17100 ( .A(n16761), .B(n16760), .Z(n16877) );
  XNOR U17101 ( .A(n102), .B(n16762), .Z(n16868) );
  OR U17102 ( .A(n16868), .B(n20121), .Z(n16765) );
  NANDN U17103 ( .A(n16763), .B(n20122), .Z(n16764) );
  NAND U17104 ( .A(n16765), .B(n16764), .Z(n16874) );
  XNOR U17105 ( .A(n19975), .B(n17257), .Z(n16871) );
  NANDN U17106 ( .A(n16871), .B(n19883), .Z(n16768) );
  NANDN U17107 ( .A(n16766), .B(n19937), .Z(n16767) );
  AND U17108 ( .A(n16768), .B(n16767), .Z(n16875) );
  XNOR U17109 ( .A(n16874), .B(n16875), .Z(n16876) );
  XNOR U17110 ( .A(n16877), .B(n16876), .Z(n16886) );
  NANDN U17111 ( .A(n16770), .B(n16769), .Z(n16774) );
  NAND U17112 ( .A(n16772), .B(n16771), .Z(n16773) );
  NAND U17113 ( .A(n16774), .B(n16773), .Z(n16887) );
  XNOR U17114 ( .A(n16886), .B(n16887), .Z(n16888) );
  NANDN U17115 ( .A(n16776), .B(n16775), .Z(n16780) );
  NAND U17116 ( .A(n16778), .B(n16777), .Z(n16779) );
  AND U17117 ( .A(n16780), .B(n16779), .Z(n16889) );
  XNOR U17118 ( .A(n16888), .B(n16889), .Z(n16833) );
  NANDN U17119 ( .A(n16782), .B(n16781), .Z(n16786) );
  OR U17120 ( .A(n16784), .B(n16783), .Z(n16785) );
  NAND U17121 ( .A(n16786), .B(n16785), .Z(n16861) );
  NAND U17122 ( .A(b[0]), .B(a[222]), .Z(n16787) );
  XNOR U17123 ( .A(b[1]), .B(n16787), .Z(n16789) );
  NAND U17124 ( .A(a[221]), .B(n98), .Z(n16788) );
  AND U17125 ( .A(n16789), .B(n16788), .Z(n16837) );
  XNOR U17126 ( .A(n20154), .B(n16918), .Z(n16846) );
  OR U17127 ( .A(n16846), .B(n20057), .Z(n16792) );
  NANDN U17128 ( .A(n16790), .B(n20098), .Z(n16791) );
  AND U17129 ( .A(n16792), .B(n16791), .Z(n16838) );
  XOR U17130 ( .A(n16837), .B(n16838), .Z(n16840) );
  NAND U17131 ( .A(a[206]), .B(b[15]), .Z(n16839) );
  XOR U17132 ( .A(n16840), .B(n16839), .Z(n16858) );
  NAND U17133 ( .A(n19722), .B(n16793), .Z(n16795) );
  XNOR U17134 ( .A(b[5]), .B(n17542), .Z(n16849) );
  NANDN U17135 ( .A(n19640), .B(n16849), .Z(n16794) );
  NAND U17136 ( .A(n16795), .B(n16794), .Z(n16883) );
  XNOR U17137 ( .A(n19714), .B(n17413), .Z(n16852) );
  NANDN U17138 ( .A(n16852), .B(n19766), .Z(n16798) );
  NANDN U17139 ( .A(n16796), .B(n19767), .Z(n16797) );
  NAND U17140 ( .A(n16798), .B(n16797), .Z(n16880) );
  NAND U17141 ( .A(n19554), .B(n16799), .Z(n16801) );
  IV U17142 ( .A(a[220]), .Z(n17725) );
  XNOR U17143 ( .A(b[3]), .B(n17725), .Z(n16855) );
  NANDN U17144 ( .A(n19521), .B(n16855), .Z(n16800) );
  AND U17145 ( .A(n16801), .B(n16800), .Z(n16881) );
  XNOR U17146 ( .A(n16880), .B(n16881), .Z(n16882) );
  XOR U17147 ( .A(n16883), .B(n16882), .Z(n16859) );
  XOR U17148 ( .A(n16858), .B(n16859), .Z(n16860) );
  XNOR U17149 ( .A(n16861), .B(n16860), .Z(n16831) );
  NAND U17150 ( .A(n16803), .B(n16802), .Z(n16807) );
  NAND U17151 ( .A(n16805), .B(n16804), .Z(n16806) );
  NAND U17152 ( .A(n16807), .B(n16806), .Z(n16832) );
  XOR U17153 ( .A(n16831), .B(n16832), .Z(n16834) );
  XNOR U17154 ( .A(n16833), .B(n16834), .Z(n16892) );
  NANDN U17155 ( .A(n16809), .B(n16808), .Z(n16813) );
  NAND U17156 ( .A(n16811), .B(n16810), .Z(n16812) );
  NAND U17157 ( .A(n16813), .B(n16812), .Z(n16893) );
  XNOR U17158 ( .A(n16892), .B(n16893), .Z(n16894) );
  XOR U17159 ( .A(n16895), .B(n16894), .Z(n16825) );
  NANDN U17160 ( .A(n16815), .B(n16814), .Z(n16819) );
  NANDN U17161 ( .A(n16817), .B(n16816), .Z(n16818) );
  NAND U17162 ( .A(n16819), .B(n16818), .Z(n16826) );
  XNOR U17163 ( .A(n16825), .B(n16826), .Z(n16827) );
  XNOR U17164 ( .A(n16828), .B(n16827), .Z(n16898) );
  XNOR U17165 ( .A(n16898), .B(sreg[462]), .Z(n16900) );
  NAND U17166 ( .A(n16820), .B(sreg[461]), .Z(n16824) );
  OR U17167 ( .A(n16822), .B(n16821), .Z(n16823) );
  AND U17168 ( .A(n16824), .B(n16823), .Z(n16899) );
  XOR U17169 ( .A(n16900), .B(n16899), .Z(c[462]) );
  NANDN U17170 ( .A(n16826), .B(n16825), .Z(n16830) );
  NAND U17171 ( .A(n16828), .B(n16827), .Z(n16829) );
  NAND U17172 ( .A(n16830), .B(n16829), .Z(n16906) );
  NANDN U17173 ( .A(n16832), .B(n16831), .Z(n16836) );
  OR U17174 ( .A(n16834), .B(n16833), .Z(n16835) );
  NAND U17175 ( .A(n16836), .B(n16835), .Z(n16973) );
  NANDN U17176 ( .A(n16838), .B(n16837), .Z(n16842) );
  OR U17177 ( .A(n16840), .B(n16839), .Z(n16841) );
  NAND U17178 ( .A(n16842), .B(n16841), .Z(n16961) );
  NAND U17179 ( .A(b[0]), .B(a[223]), .Z(n16843) );
  XNOR U17180 ( .A(b[1]), .B(n16843), .Z(n16845) );
  NAND U17181 ( .A(a[222]), .B(n98), .Z(n16844) );
  AND U17182 ( .A(n16845), .B(n16844), .Z(n16937) );
  XNOR U17183 ( .A(n20154), .B(n17008), .Z(n16946) );
  OR U17184 ( .A(n16946), .B(n20057), .Z(n16848) );
  NANDN U17185 ( .A(n16846), .B(n20098), .Z(n16847) );
  AND U17186 ( .A(n16848), .B(n16847), .Z(n16938) );
  XOR U17187 ( .A(n16937), .B(n16938), .Z(n16940) );
  NAND U17188 ( .A(a[207]), .B(b[15]), .Z(n16939) );
  XOR U17189 ( .A(n16940), .B(n16939), .Z(n16958) );
  NAND U17190 ( .A(n19722), .B(n16849), .Z(n16851) );
  XNOR U17191 ( .A(b[5]), .B(n17620), .Z(n16949) );
  NANDN U17192 ( .A(n19640), .B(n16949), .Z(n16850) );
  NAND U17193 ( .A(n16851), .B(n16850), .Z(n16934) );
  XNOR U17194 ( .A(n19714), .B(n17464), .Z(n16952) );
  NANDN U17195 ( .A(n16952), .B(n19766), .Z(n16854) );
  NANDN U17196 ( .A(n16852), .B(n19767), .Z(n16853) );
  NAND U17197 ( .A(n16854), .B(n16853), .Z(n16931) );
  NAND U17198 ( .A(n19554), .B(n16855), .Z(n16857) );
  IV U17199 ( .A(a[221]), .Z(n17776) );
  XNOR U17200 ( .A(b[3]), .B(n17776), .Z(n16955) );
  NANDN U17201 ( .A(n19521), .B(n16955), .Z(n16856) );
  AND U17202 ( .A(n16857), .B(n16856), .Z(n16932) );
  XNOR U17203 ( .A(n16931), .B(n16932), .Z(n16933) );
  XOR U17204 ( .A(n16934), .B(n16933), .Z(n16959) );
  XOR U17205 ( .A(n16958), .B(n16959), .Z(n16960) );
  XNOR U17206 ( .A(n16961), .B(n16960), .Z(n16909) );
  NAND U17207 ( .A(n16859), .B(n16858), .Z(n16863) );
  NAND U17208 ( .A(n16861), .B(n16860), .Z(n16862) );
  NAND U17209 ( .A(n16863), .B(n16862), .Z(n16910) );
  XOR U17210 ( .A(n16909), .B(n16910), .Z(n16912) );
  XNOR U17211 ( .A(n20052), .B(n17152), .Z(n16915) );
  OR U17212 ( .A(n16915), .B(n20020), .Z(n16866) );
  NANDN U17213 ( .A(n16864), .B(n19960), .Z(n16865) );
  NAND U17214 ( .A(n16866), .B(n16865), .Z(n16928) );
  XNOR U17215 ( .A(n102), .B(n16867), .Z(n16919) );
  OR U17216 ( .A(n16919), .B(n20121), .Z(n16870) );
  NANDN U17217 ( .A(n16868), .B(n20122), .Z(n16869) );
  NAND U17218 ( .A(n16870), .B(n16869), .Z(n16925) );
  XNOR U17219 ( .A(n19975), .B(n17308), .Z(n16922) );
  NANDN U17220 ( .A(n16922), .B(n19883), .Z(n16873) );
  NANDN U17221 ( .A(n16871), .B(n19937), .Z(n16872) );
  AND U17222 ( .A(n16873), .B(n16872), .Z(n16926) );
  XNOR U17223 ( .A(n16925), .B(n16926), .Z(n16927) );
  XNOR U17224 ( .A(n16928), .B(n16927), .Z(n16964) );
  NANDN U17225 ( .A(n16875), .B(n16874), .Z(n16879) );
  NAND U17226 ( .A(n16877), .B(n16876), .Z(n16878) );
  NAND U17227 ( .A(n16879), .B(n16878), .Z(n16965) );
  XNOR U17228 ( .A(n16964), .B(n16965), .Z(n16966) );
  NANDN U17229 ( .A(n16881), .B(n16880), .Z(n16885) );
  NAND U17230 ( .A(n16883), .B(n16882), .Z(n16884) );
  AND U17231 ( .A(n16885), .B(n16884), .Z(n16967) );
  XNOR U17232 ( .A(n16966), .B(n16967), .Z(n16911) );
  XNOR U17233 ( .A(n16912), .B(n16911), .Z(n16970) );
  NANDN U17234 ( .A(n16887), .B(n16886), .Z(n16891) );
  NAND U17235 ( .A(n16889), .B(n16888), .Z(n16890) );
  NAND U17236 ( .A(n16891), .B(n16890), .Z(n16971) );
  XNOR U17237 ( .A(n16970), .B(n16971), .Z(n16972) );
  XOR U17238 ( .A(n16973), .B(n16972), .Z(n16903) );
  NANDN U17239 ( .A(n16893), .B(n16892), .Z(n16897) );
  NANDN U17240 ( .A(n16895), .B(n16894), .Z(n16896) );
  NAND U17241 ( .A(n16897), .B(n16896), .Z(n16904) );
  XNOR U17242 ( .A(n16903), .B(n16904), .Z(n16905) );
  XNOR U17243 ( .A(n16906), .B(n16905), .Z(n16976) );
  XNOR U17244 ( .A(n16976), .B(sreg[463]), .Z(n16978) );
  NAND U17245 ( .A(n16898), .B(sreg[462]), .Z(n16902) );
  OR U17246 ( .A(n16900), .B(n16899), .Z(n16901) );
  AND U17247 ( .A(n16902), .B(n16901), .Z(n16977) );
  XOR U17248 ( .A(n16978), .B(n16977), .Z(c[463]) );
  NANDN U17249 ( .A(n16904), .B(n16903), .Z(n16908) );
  NAND U17250 ( .A(n16906), .B(n16905), .Z(n16907) );
  NAND U17251 ( .A(n16908), .B(n16907), .Z(n16984) );
  NANDN U17252 ( .A(n16910), .B(n16909), .Z(n16914) );
  OR U17253 ( .A(n16912), .B(n16911), .Z(n16913) );
  NAND U17254 ( .A(n16914), .B(n16913), .Z(n17051) );
  XNOR U17255 ( .A(n20052), .B(n17257), .Z(n17005) );
  OR U17256 ( .A(n17005), .B(n20020), .Z(n16917) );
  NANDN U17257 ( .A(n16915), .B(n19960), .Z(n16916) );
  NAND U17258 ( .A(n16917), .B(n16916), .Z(n17002) );
  XNOR U17259 ( .A(n102), .B(n16918), .Z(n17009) );
  OR U17260 ( .A(n17009), .B(n20121), .Z(n16921) );
  NANDN U17261 ( .A(n16919), .B(n20122), .Z(n16920) );
  NAND U17262 ( .A(n16921), .B(n16920), .Z(n16999) );
  XNOR U17263 ( .A(n19975), .B(n17413), .Z(n17012) );
  NANDN U17264 ( .A(n17012), .B(n19883), .Z(n16924) );
  NANDN U17265 ( .A(n16922), .B(n19937), .Z(n16923) );
  AND U17266 ( .A(n16924), .B(n16923), .Z(n17000) );
  XNOR U17267 ( .A(n16999), .B(n17000), .Z(n17001) );
  XNOR U17268 ( .A(n17002), .B(n17001), .Z(n17042) );
  NANDN U17269 ( .A(n16926), .B(n16925), .Z(n16930) );
  NAND U17270 ( .A(n16928), .B(n16927), .Z(n16929) );
  NAND U17271 ( .A(n16930), .B(n16929), .Z(n17043) );
  XNOR U17272 ( .A(n17042), .B(n17043), .Z(n17044) );
  NANDN U17273 ( .A(n16932), .B(n16931), .Z(n16936) );
  NAND U17274 ( .A(n16934), .B(n16933), .Z(n16935) );
  AND U17275 ( .A(n16936), .B(n16935), .Z(n17045) );
  XNOR U17276 ( .A(n17044), .B(n17045), .Z(n16989) );
  NANDN U17277 ( .A(n16938), .B(n16937), .Z(n16942) );
  OR U17278 ( .A(n16940), .B(n16939), .Z(n16941) );
  NAND U17279 ( .A(n16942), .B(n16941), .Z(n17039) );
  NAND U17280 ( .A(b[0]), .B(a[224]), .Z(n16943) );
  XNOR U17281 ( .A(b[1]), .B(n16943), .Z(n16945) );
  NAND U17282 ( .A(a[223]), .B(n98), .Z(n16944) );
  AND U17283 ( .A(n16945), .B(n16944), .Z(n17015) );
  XNOR U17284 ( .A(n20154), .B(n17074), .Z(n17024) );
  OR U17285 ( .A(n17024), .B(n20057), .Z(n16948) );
  NANDN U17286 ( .A(n16946), .B(n20098), .Z(n16947) );
  AND U17287 ( .A(n16948), .B(n16947), .Z(n17016) );
  XOR U17288 ( .A(n17015), .B(n17016), .Z(n17018) );
  NAND U17289 ( .A(a[208]), .B(b[15]), .Z(n17017) );
  XOR U17290 ( .A(n17018), .B(n17017), .Z(n17036) );
  NAND U17291 ( .A(n19722), .B(n16949), .Z(n16951) );
  XNOR U17292 ( .A(b[5]), .B(n17725), .Z(n17027) );
  NANDN U17293 ( .A(n19640), .B(n17027), .Z(n16950) );
  NAND U17294 ( .A(n16951), .B(n16950), .Z(n16996) );
  XNOR U17295 ( .A(n19714), .B(n17542), .Z(n17030) );
  NANDN U17296 ( .A(n17030), .B(n19766), .Z(n16954) );
  NANDN U17297 ( .A(n16952), .B(n19767), .Z(n16953) );
  NAND U17298 ( .A(n16954), .B(n16953), .Z(n16993) );
  NAND U17299 ( .A(n19554), .B(n16955), .Z(n16957) );
  IV U17300 ( .A(a[222]), .Z(n17854) );
  XNOR U17301 ( .A(b[3]), .B(n17854), .Z(n17033) );
  NANDN U17302 ( .A(n19521), .B(n17033), .Z(n16956) );
  AND U17303 ( .A(n16957), .B(n16956), .Z(n16994) );
  XNOR U17304 ( .A(n16993), .B(n16994), .Z(n16995) );
  XOR U17305 ( .A(n16996), .B(n16995), .Z(n17037) );
  XOR U17306 ( .A(n17036), .B(n17037), .Z(n17038) );
  XNOR U17307 ( .A(n17039), .B(n17038), .Z(n16987) );
  NAND U17308 ( .A(n16959), .B(n16958), .Z(n16963) );
  NAND U17309 ( .A(n16961), .B(n16960), .Z(n16962) );
  NAND U17310 ( .A(n16963), .B(n16962), .Z(n16988) );
  XOR U17311 ( .A(n16987), .B(n16988), .Z(n16990) );
  XNOR U17312 ( .A(n16989), .B(n16990), .Z(n17048) );
  NANDN U17313 ( .A(n16965), .B(n16964), .Z(n16969) );
  NAND U17314 ( .A(n16967), .B(n16966), .Z(n16968) );
  NAND U17315 ( .A(n16969), .B(n16968), .Z(n17049) );
  XNOR U17316 ( .A(n17048), .B(n17049), .Z(n17050) );
  XOR U17317 ( .A(n17051), .B(n17050), .Z(n16981) );
  NANDN U17318 ( .A(n16971), .B(n16970), .Z(n16975) );
  NANDN U17319 ( .A(n16973), .B(n16972), .Z(n16974) );
  NAND U17320 ( .A(n16975), .B(n16974), .Z(n16982) );
  XNOR U17321 ( .A(n16981), .B(n16982), .Z(n16983) );
  XNOR U17322 ( .A(n16984), .B(n16983), .Z(n17054) );
  XNOR U17323 ( .A(n17054), .B(sreg[464]), .Z(n17056) );
  NAND U17324 ( .A(n16976), .B(sreg[463]), .Z(n16980) );
  OR U17325 ( .A(n16978), .B(n16977), .Z(n16979) );
  AND U17326 ( .A(n16980), .B(n16979), .Z(n17055) );
  XOR U17327 ( .A(n17056), .B(n17055), .Z(c[464]) );
  NANDN U17328 ( .A(n16982), .B(n16981), .Z(n16986) );
  NAND U17329 ( .A(n16984), .B(n16983), .Z(n16985) );
  NAND U17330 ( .A(n16986), .B(n16985), .Z(n17062) );
  NANDN U17331 ( .A(n16988), .B(n16987), .Z(n16992) );
  OR U17332 ( .A(n16990), .B(n16989), .Z(n16991) );
  NAND U17333 ( .A(n16992), .B(n16991), .Z(n17129) );
  NANDN U17334 ( .A(n16994), .B(n16993), .Z(n16998) );
  NAND U17335 ( .A(n16996), .B(n16995), .Z(n16997) );
  NAND U17336 ( .A(n16998), .B(n16997), .Z(n17123) );
  NANDN U17337 ( .A(n17000), .B(n16999), .Z(n17004) );
  NAND U17338 ( .A(n17002), .B(n17001), .Z(n17003) );
  NAND U17339 ( .A(n17004), .B(n17003), .Z(n17120) );
  XNOR U17340 ( .A(n20052), .B(n17308), .Z(n17071) );
  OR U17341 ( .A(n17071), .B(n20020), .Z(n17007) );
  NANDN U17342 ( .A(n17005), .B(n19960), .Z(n17006) );
  NAND U17343 ( .A(n17007), .B(n17006), .Z(n17084) );
  XNOR U17344 ( .A(n102), .B(n17008), .Z(n17075) );
  OR U17345 ( .A(n17075), .B(n20121), .Z(n17011) );
  NANDN U17346 ( .A(n17009), .B(n20122), .Z(n17010) );
  NAND U17347 ( .A(n17011), .B(n17010), .Z(n17081) );
  XNOR U17348 ( .A(n19975), .B(n17464), .Z(n17078) );
  NANDN U17349 ( .A(n17078), .B(n19883), .Z(n17014) );
  NANDN U17350 ( .A(n17012), .B(n19937), .Z(n17013) );
  AND U17351 ( .A(n17014), .B(n17013), .Z(n17082) );
  XNOR U17352 ( .A(n17081), .B(n17082), .Z(n17083) );
  XNOR U17353 ( .A(n17084), .B(n17083), .Z(n17121) );
  XNOR U17354 ( .A(n17120), .B(n17121), .Z(n17122) );
  XNOR U17355 ( .A(n17123), .B(n17122), .Z(n17068) );
  NANDN U17356 ( .A(n17016), .B(n17015), .Z(n17020) );
  OR U17357 ( .A(n17018), .B(n17017), .Z(n17019) );
  NAND U17358 ( .A(n17020), .B(n17019), .Z(n17117) );
  NAND U17359 ( .A(b[0]), .B(a[225]), .Z(n17021) );
  XNOR U17360 ( .A(b[1]), .B(n17021), .Z(n17023) );
  NAND U17361 ( .A(a[224]), .B(n98), .Z(n17022) );
  AND U17362 ( .A(n17023), .B(n17022), .Z(n17093) );
  XNOR U17363 ( .A(n20154), .B(n17152), .Z(n17099) );
  OR U17364 ( .A(n17099), .B(n20057), .Z(n17026) );
  NANDN U17365 ( .A(n17024), .B(n20098), .Z(n17025) );
  AND U17366 ( .A(n17026), .B(n17025), .Z(n17094) );
  XOR U17367 ( .A(n17093), .B(n17094), .Z(n17096) );
  NAND U17368 ( .A(a[209]), .B(b[15]), .Z(n17095) );
  XOR U17369 ( .A(n17096), .B(n17095), .Z(n17114) );
  NAND U17370 ( .A(n19722), .B(n17027), .Z(n17029) );
  XNOR U17371 ( .A(b[5]), .B(n17776), .Z(n17105) );
  NANDN U17372 ( .A(n19640), .B(n17105), .Z(n17028) );
  NAND U17373 ( .A(n17029), .B(n17028), .Z(n17090) );
  XNOR U17374 ( .A(n19714), .B(n17620), .Z(n17108) );
  NANDN U17375 ( .A(n17108), .B(n19766), .Z(n17032) );
  NANDN U17376 ( .A(n17030), .B(n19767), .Z(n17031) );
  NAND U17377 ( .A(n17032), .B(n17031), .Z(n17087) );
  NAND U17378 ( .A(n19554), .B(n17033), .Z(n17035) );
  IV U17379 ( .A(a[223]), .Z(n17932) );
  XNOR U17380 ( .A(b[3]), .B(n17932), .Z(n17111) );
  NANDN U17381 ( .A(n19521), .B(n17111), .Z(n17034) );
  AND U17382 ( .A(n17035), .B(n17034), .Z(n17088) );
  XNOR U17383 ( .A(n17087), .B(n17088), .Z(n17089) );
  XOR U17384 ( .A(n17090), .B(n17089), .Z(n17115) );
  XOR U17385 ( .A(n17114), .B(n17115), .Z(n17116) );
  XNOR U17386 ( .A(n17117), .B(n17116), .Z(n17065) );
  NAND U17387 ( .A(n17037), .B(n17036), .Z(n17041) );
  NAND U17388 ( .A(n17039), .B(n17038), .Z(n17040) );
  NAND U17389 ( .A(n17041), .B(n17040), .Z(n17066) );
  XNOR U17390 ( .A(n17065), .B(n17066), .Z(n17067) );
  XOR U17391 ( .A(n17068), .B(n17067), .Z(n17126) );
  NANDN U17392 ( .A(n17043), .B(n17042), .Z(n17047) );
  NAND U17393 ( .A(n17045), .B(n17044), .Z(n17046) );
  NAND U17394 ( .A(n17047), .B(n17046), .Z(n17127) );
  XOR U17395 ( .A(n17126), .B(n17127), .Z(n17128) );
  XOR U17396 ( .A(n17129), .B(n17128), .Z(n17059) );
  NANDN U17397 ( .A(n17049), .B(n17048), .Z(n17053) );
  NANDN U17398 ( .A(n17051), .B(n17050), .Z(n17052) );
  NAND U17399 ( .A(n17053), .B(n17052), .Z(n17060) );
  XNOR U17400 ( .A(n17059), .B(n17060), .Z(n17061) );
  XNOR U17401 ( .A(n17062), .B(n17061), .Z(n17132) );
  XNOR U17402 ( .A(n17132), .B(sreg[465]), .Z(n17134) );
  NAND U17403 ( .A(n17054), .B(sreg[464]), .Z(n17058) );
  OR U17404 ( .A(n17056), .B(n17055), .Z(n17057) );
  AND U17405 ( .A(n17058), .B(n17057), .Z(n17133) );
  XOR U17406 ( .A(n17134), .B(n17133), .Z(c[465]) );
  NANDN U17407 ( .A(n17060), .B(n17059), .Z(n17064) );
  NAND U17408 ( .A(n17062), .B(n17061), .Z(n17063) );
  NAND U17409 ( .A(n17064), .B(n17063), .Z(n17140) );
  NANDN U17410 ( .A(n17066), .B(n17065), .Z(n17070) );
  NAND U17411 ( .A(n17068), .B(n17067), .Z(n17069) );
  NAND U17412 ( .A(n17070), .B(n17069), .Z(n17207) );
  XNOR U17413 ( .A(n20052), .B(n17413), .Z(n17149) );
  OR U17414 ( .A(n17149), .B(n20020), .Z(n17073) );
  NANDN U17415 ( .A(n17071), .B(n19960), .Z(n17072) );
  NAND U17416 ( .A(n17073), .B(n17072), .Z(n17162) );
  XNOR U17417 ( .A(n102), .B(n17074), .Z(n17153) );
  OR U17418 ( .A(n17153), .B(n20121), .Z(n17077) );
  NANDN U17419 ( .A(n17075), .B(n20122), .Z(n17076) );
  NAND U17420 ( .A(n17077), .B(n17076), .Z(n17159) );
  XNOR U17421 ( .A(n19975), .B(n17542), .Z(n17156) );
  NANDN U17422 ( .A(n17156), .B(n19883), .Z(n17080) );
  NANDN U17423 ( .A(n17078), .B(n19937), .Z(n17079) );
  AND U17424 ( .A(n17080), .B(n17079), .Z(n17160) );
  XNOR U17425 ( .A(n17159), .B(n17160), .Z(n17161) );
  XNOR U17426 ( .A(n17162), .B(n17161), .Z(n17198) );
  NANDN U17427 ( .A(n17082), .B(n17081), .Z(n17086) );
  NAND U17428 ( .A(n17084), .B(n17083), .Z(n17085) );
  NAND U17429 ( .A(n17086), .B(n17085), .Z(n17199) );
  XNOR U17430 ( .A(n17198), .B(n17199), .Z(n17200) );
  NANDN U17431 ( .A(n17088), .B(n17087), .Z(n17092) );
  NAND U17432 ( .A(n17090), .B(n17089), .Z(n17091) );
  AND U17433 ( .A(n17092), .B(n17091), .Z(n17201) );
  XNOR U17434 ( .A(n17200), .B(n17201), .Z(n17145) );
  NANDN U17435 ( .A(n17094), .B(n17093), .Z(n17098) );
  OR U17436 ( .A(n17096), .B(n17095), .Z(n17097) );
  NAND U17437 ( .A(n17098), .B(n17097), .Z(n17195) );
  XNOR U17438 ( .A(n20154), .B(n17257), .Z(n17180) );
  OR U17439 ( .A(n17180), .B(n20057), .Z(n17101) );
  NANDN U17440 ( .A(n17099), .B(n20098), .Z(n17100) );
  AND U17441 ( .A(n17101), .B(n17100), .Z(n17172) );
  NAND U17442 ( .A(b[0]), .B(a[226]), .Z(n17102) );
  XNOR U17443 ( .A(b[1]), .B(n17102), .Z(n17104) );
  NAND U17444 ( .A(a[225]), .B(n98), .Z(n17103) );
  AND U17445 ( .A(n17104), .B(n17103), .Z(n17171) );
  XOR U17446 ( .A(n17172), .B(n17171), .Z(n17174) );
  NAND U17447 ( .A(a[210]), .B(b[15]), .Z(n17173) );
  XOR U17448 ( .A(n17174), .B(n17173), .Z(n17192) );
  NAND U17449 ( .A(n19722), .B(n17105), .Z(n17107) );
  XNOR U17450 ( .A(b[5]), .B(n17854), .Z(n17183) );
  NANDN U17451 ( .A(n19640), .B(n17183), .Z(n17106) );
  NAND U17452 ( .A(n17107), .B(n17106), .Z(n17168) );
  XNOR U17453 ( .A(n19714), .B(n17725), .Z(n17186) );
  NANDN U17454 ( .A(n17186), .B(n19766), .Z(n17110) );
  NANDN U17455 ( .A(n17108), .B(n19767), .Z(n17109) );
  NAND U17456 ( .A(n17110), .B(n17109), .Z(n17165) );
  NAND U17457 ( .A(n19554), .B(n17111), .Z(n17113) );
  IV U17458 ( .A(a[224]), .Z(n18037) );
  XNOR U17459 ( .A(b[3]), .B(n18037), .Z(n17189) );
  NANDN U17460 ( .A(n19521), .B(n17189), .Z(n17112) );
  AND U17461 ( .A(n17113), .B(n17112), .Z(n17166) );
  XNOR U17462 ( .A(n17165), .B(n17166), .Z(n17167) );
  XOR U17463 ( .A(n17168), .B(n17167), .Z(n17193) );
  XOR U17464 ( .A(n17192), .B(n17193), .Z(n17194) );
  XNOR U17465 ( .A(n17195), .B(n17194), .Z(n17143) );
  NAND U17466 ( .A(n17115), .B(n17114), .Z(n17119) );
  NAND U17467 ( .A(n17117), .B(n17116), .Z(n17118) );
  NAND U17468 ( .A(n17119), .B(n17118), .Z(n17144) );
  XOR U17469 ( .A(n17143), .B(n17144), .Z(n17146) );
  XNOR U17470 ( .A(n17145), .B(n17146), .Z(n17204) );
  NANDN U17471 ( .A(n17121), .B(n17120), .Z(n17125) );
  NAND U17472 ( .A(n17123), .B(n17122), .Z(n17124) );
  AND U17473 ( .A(n17125), .B(n17124), .Z(n17205) );
  XNOR U17474 ( .A(n17204), .B(n17205), .Z(n17206) );
  XOR U17475 ( .A(n17207), .B(n17206), .Z(n17137) );
  OR U17476 ( .A(n17127), .B(n17126), .Z(n17131) );
  NANDN U17477 ( .A(n17129), .B(n17128), .Z(n17130) );
  NAND U17478 ( .A(n17131), .B(n17130), .Z(n17138) );
  XNOR U17479 ( .A(n17137), .B(n17138), .Z(n17139) );
  XNOR U17480 ( .A(n17140), .B(n17139), .Z(n17210) );
  XNOR U17481 ( .A(n17210), .B(sreg[466]), .Z(n17212) );
  NAND U17482 ( .A(n17132), .B(sreg[465]), .Z(n17136) );
  OR U17483 ( .A(n17134), .B(n17133), .Z(n17135) );
  AND U17484 ( .A(n17136), .B(n17135), .Z(n17211) );
  XOR U17485 ( .A(n17212), .B(n17211), .Z(c[466]) );
  NANDN U17486 ( .A(n17138), .B(n17137), .Z(n17142) );
  NAND U17487 ( .A(n17140), .B(n17139), .Z(n17141) );
  NAND U17488 ( .A(n17142), .B(n17141), .Z(n17218) );
  NANDN U17489 ( .A(n17144), .B(n17143), .Z(n17148) );
  OR U17490 ( .A(n17146), .B(n17145), .Z(n17147) );
  NAND U17491 ( .A(n17148), .B(n17147), .Z(n17285) );
  XNOR U17492 ( .A(n20052), .B(n17464), .Z(n17254) );
  OR U17493 ( .A(n17254), .B(n20020), .Z(n17151) );
  NANDN U17494 ( .A(n17149), .B(n19960), .Z(n17150) );
  NAND U17495 ( .A(n17151), .B(n17150), .Z(n17267) );
  XNOR U17496 ( .A(n102), .B(n17152), .Z(n17258) );
  OR U17497 ( .A(n17258), .B(n20121), .Z(n17155) );
  NANDN U17498 ( .A(n17153), .B(n20122), .Z(n17154) );
  NAND U17499 ( .A(n17155), .B(n17154), .Z(n17264) );
  XNOR U17500 ( .A(n19975), .B(n17620), .Z(n17261) );
  NANDN U17501 ( .A(n17261), .B(n19883), .Z(n17158) );
  NANDN U17502 ( .A(n17156), .B(n19937), .Z(n17157) );
  AND U17503 ( .A(n17158), .B(n17157), .Z(n17265) );
  XNOR U17504 ( .A(n17264), .B(n17265), .Z(n17266) );
  XNOR U17505 ( .A(n17267), .B(n17266), .Z(n17276) );
  NANDN U17506 ( .A(n17160), .B(n17159), .Z(n17164) );
  NAND U17507 ( .A(n17162), .B(n17161), .Z(n17163) );
  NAND U17508 ( .A(n17164), .B(n17163), .Z(n17277) );
  XNOR U17509 ( .A(n17276), .B(n17277), .Z(n17278) );
  NANDN U17510 ( .A(n17166), .B(n17165), .Z(n17170) );
  NAND U17511 ( .A(n17168), .B(n17167), .Z(n17169) );
  AND U17512 ( .A(n17170), .B(n17169), .Z(n17279) );
  XNOR U17513 ( .A(n17278), .B(n17279), .Z(n17223) );
  NANDN U17514 ( .A(n17172), .B(n17171), .Z(n17176) );
  OR U17515 ( .A(n17174), .B(n17173), .Z(n17175) );
  NAND U17516 ( .A(n17176), .B(n17175), .Z(n17251) );
  NAND U17517 ( .A(b[0]), .B(a[227]), .Z(n17177) );
  XNOR U17518 ( .A(b[1]), .B(n17177), .Z(n17179) );
  NAND U17519 ( .A(a[226]), .B(n98), .Z(n17178) );
  AND U17520 ( .A(n17179), .B(n17178), .Z(n17227) );
  XNOR U17521 ( .A(n20154), .B(n17308), .Z(n17236) );
  OR U17522 ( .A(n17236), .B(n20057), .Z(n17182) );
  NANDN U17523 ( .A(n17180), .B(n20098), .Z(n17181) );
  AND U17524 ( .A(n17182), .B(n17181), .Z(n17228) );
  XOR U17525 ( .A(n17227), .B(n17228), .Z(n17230) );
  NAND U17526 ( .A(a[211]), .B(b[15]), .Z(n17229) );
  XOR U17527 ( .A(n17230), .B(n17229), .Z(n17248) );
  NAND U17528 ( .A(n19722), .B(n17183), .Z(n17185) );
  XNOR U17529 ( .A(b[5]), .B(n17932), .Z(n17239) );
  NANDN U17530 ( .A(n19640), .B(n17239), .Z(n17184) );
  NAND U17531 ( .A(n17185), .B(n17184), .Z(n17273) );
  XNOR U17532 ( .A(n19714), .B(n17776), .Z(n17242) );
  NANDN U17533 ( .A(n17242), .B(n19766), .Z(n17188) );
  NANDN U17534 ( .A(n17186), .B(n19767), .Z(n17187) );
  NAND U17535 ( .A(n17188), .B(n17187), .Z(n17270) );
  NAND U17536 ( .A(n19554), .B(n17189), .Z(n17191) );
  IV U17537 ( .A(a[225]), .Z(n18115) );
  XNOR U17538 ( .A(b[3]), .B(n18115), .Z(n17245) );
  NANDN U17539 ( .A(n19521), .B(n17245), .Z(n17190) );
  AND U17540 ( .A(n17191), .B(n17190), .Z(n17271) );
  XNOR U17541 ( .A(n17270), .B(n17271), .Z(n17272) );
  XOR U17542 ( .A(n17273), .B(n17272), .Z(n17249) );
  XOR U17543 ( .A(n17248), .B(n17249), .Z(n17250) );
  XNOR U17544 ( .A(n17251), .B(n17250), .Z(n17221) );
  NAND U17545 ( .A(n17193), .B(n17192), .Z(n17197) );
  NAND U17546 ( .A(n17195), .B(n17194), .Z(n17196) );
  NAND U17547 ( .A(n17197), .B(n17196), .Z(n17222) );
  XOR U17548 ( .A(n17221), .B(n17222), .Z(n17224) );
  XNOR U17549 ( .A(n17223), .B(n17224), .Z(n17282) );
  NANDN U17550 ( .A(n17199), .B(n17198), .Z(n17203) );
  NAND U17551 ( .A(n17201), .B(n17200), .Z(n17202) );
  NAND U17552 ( .A(n17203), .B(n17202), .Z(n17283) );
  XNOR U17553 ( .A(n17282), .B(n17283), .Z(n17284) );
  XOR U17554 ( .A(n17285), .B(n17284), .Z(n17215) );
  NANDN U17555 ( .A(n17205), .B(n17204), .Z(n17209) );
  NANDN U17556 ( .A(n17207), .B(n17206), .Z(n17208) );
  NAND U17557 ( .A(n17209), .B(n17208), .Z(n17216) );
  XNOR U17558 ( .A(n17215), .B(n17216), .Z(n17217) );
  XNOR U17559 ( .A(n17218), .B(n17217), .Z(n17288) );
  XNOR U17560 ( .A(n17288), .B(sreg[467]), .Z(n17290) );
  NAND U17561 ( .A(n17210), .B(sreg[466]), .Z(n17214) );
  OR U17562 ( .A(n17212), .B(n17211), .Z(n17213) );
  AND U17563 ( .A(n17214), .B(n17213), .Z(n17289) );
  XOR U17564 ( .A(n17290), .B(n17289), .Z(c[467]) );
  NANDN U17565 ( .A(n17216), .B(n17215), .Z(n17220) );
  NAND U17566 ( .A(n17218), .B(n17217), .Z(n17219) );
  NAND U17567 ( .A(n17220), .B(n17219), .Z(n17296) );
  NANDN U17568 ( .A(n17222), .B(n17221), .Z(n17226) );
  OR U17569 ( .A(n17224), .B(n17223), .Z(n17225) );
  NAND U17570 ( .A(n17226), .B(n17225), .Z(n17363) );
  NANDN U17571 ( .A(n17228), .B(n17227), .Z(n17232) );
  OR U17572 ( .A(n17230), .B(n17229), .Z(n17231) );
  NAND U17573 ( .A(n17232), .B(n17231), .Z(n17351) );
  NAND U17574 ( .A(b[0]), .B(a[228]), .Z(n17233) );
  XNOR U17575 ( .A(b[1]), .B(n17233), .Z(n17235) );
  NAND U17576 ( .A(a[227]), .B(n98), .Z(n17234) );
  AND U17577 ( .A(n17235), .B(n17234), .Z(n17327) );
  XNOR U17578 ( .A(n20154), .B(n17413), .Z(n17333) );
  OR U17579 ( .A(n17333), .B(n20057), .Z(n17238) );
  NANDN U17580 ( .A(n17236), .B(n20098), .Z(n17237) );
  AND U17581 ( .A(n17238), .B(n17237), .Z(n17328) );
  XOR U17582 ( .A(n17327), .B(n17328), .Z(n17330) );
  NAND U17583 ( .A(a[212]), .B(b[15]), .Z(n17329) );
  XOR U17584 ( .A(n17330), .B(n17329), .Z(n17348) );
  NAND U17585 ( .A(n19722), .B(n17239), .Z(n17241) );
  XNOR U17586 ( .A(b[5]), .B(n18037), .Z(n17339) );
  NANDN U17587 ( .A(n19640), .B(n17339), .Z(n17240) );
  NAND U17588 ( .A(n17241), .B(n17240), .Z(n17324) );
  XNOR U17589 ( .A(n19714), .B(n17854), .Z(n17342) );
  NANDN U17590 ( .A(n17342), .B(n19766), .Z(n17244) );
  NANDN U17591 ( .A(n17242), .B(n19767), .Z(n17243) );
  NAND U17592 ( .A(n17244), .B(n17243), .Z(n17321) );
  NAND U17593 ( .A(n19554), .B(n17245), .Z(n17247) );
  IV U17594 ( .A(a[226]), .Z(n18193) );
  XNOR U17595 ( .A(b[3]), .B(n18193), .Z(n17345) );
  NANDN U17596 ( .A(n19521), .B(n17345), .Z(n17246) );
  AND U17597 ( .A(n17247), .B(n17246), .Z(n17322) );
  XNOR U17598 ( .A(n17321), .B(n17322), .Z(n17323) );
  XOR U17599 ( .A(n17324), .B(n17323), .Z(n17349) );
  XOR U17600 ( .A(n17348), .B(n17349), .Z(n17350) );
  XNOR U17601 ( .A(n17351), .B(n17350), .Z(n17299) );
  NAND U17602 ( .A(n17249), .B(n17248), .Z(n17253) );
  NAND U17603 ( .A(n17251), .B(n17250), .Z(n17252) );
  NAND U17604 ( .A(n17253), .B(n17252), .Z(n17300) );
  XOR U17605 ( .A(n17299), .B(n17300), .Z(n17302) );
  XNOR U17606 ( .A(n20052), .B(n17542), .Z(n17305) );
  OR U17607 ( .A(n17305), .B(n20020), .Z(n17256) );
  NANDN U17608 ( .A(n17254), .B(n19960), .Z(n17255) );
  NAND U17609 ( .A(n17256), .B(n17255), .Z(n17318) );
  XNOR U17610 ( .A(n102), .B(n17257), .Z(n17309) );
  OR U17611 ( .A(n17309), .B(n20121), .Z(n17260) );
  NANDN U17612 ( .A(n17258), .B(n20122), .Z(n17259) );
  NAND U17613 ( .A(n17260), .B(n17259), .Z(n17315) );
  XNOR U17614 ( .A(n19975), .B(n17725), .Z(n17312) );
  NANDN U17615 ( .A(n17312), .B(n19883), .Z(n17263) );
  NANDN U17616 ( .A(n17261), .B(n19937), .Z(n17262) );
  AND U17617 ( .A(n17263), .B(n17262), .Z(n17316) );
  XNOR U17618 ( .A(n17315), .B(n17316), .Z(n17317) );
  XNOR U17619 ( .A(n17318), .B(n17317), .Z(n17354) );
  NANDN U17620 ( .A(n17265), .B(n17264), .Z(n17269) );
  NAND U17621 ( .A(n17267), .B(n17266), .Z(n17268) );
  NAND U17622 ( .A(n17269), .B(n17268), .Z(n17355) );
  XNOR U17623 ( .A(n17354), .B(n17355), .Z(n17356) );
  NANDN U17624 ( .A(n17271), .B(n17270), .Z(n17275) );
  NAND U17625 ( .A(n17273), .B(n17272), .Z(n17274) );
  AND U17626 ( .A(n17275), .B(n17274), .Z(n17357) );
  XNOR U17627 ( .A(n17356), .B(n17357), .Z(n17301) );
  XNOR U17628 ( .A(n17302), .B(n17301), .Z(n17360) );
  NANDN U17629 ( .A(n17277), .B(n17276), .Z(n17281) );
  NAND U17630 ( .A(n17279), .B(n17278), .Z(n17280) );
  NAND U17631 ( .A(n17281), .B(n17280), .Z(n17361) );
  XNOR U17632 ( .A(n17360), .B(n17361), .Z(n17362) );
  XOR U17633 ( .A(n17363), .B(n17362), .Z(n17293) );
  NANDN U17634 ( .A(n17283), .B(n17282), .Z(n17287) );
  NANDN U17635 ( .A(n17285), .B(n17284), .Z(n17286) );
  NAND U17636 ( .A(n17287), .B(n17286), .Z(n17294) );
  XNOR U17637 ( .A(n17293), .B(n17294), .Z(n17295) );
  XNOR U17638 ( .A(n17296), .B(n17295), .Z(n17366) );
  XNOR U17639 ( .A(n17366), .B(sreg[468]), .Z(n17368) );
  NAND U17640 ( .A(n17288), .B(sreg[467]), .Z(n17292) );
  OR U17641 ( .A(n17290), .B(n17289), .Z(n17291) );
  AND U17642 ( .A(n17292), .B(n17291), .Z(n17367) );
  XOR U17643 ( .A(n17368), .B(n17367), .Z(c[468]) );
  NANDN U17644 ( .A(n17294), .B(n17293), .Z(n17298) );
  NAND U17645 ( .A(n17296), .B(n17295), .Z(n17297) );
  NAND U17646 ( .A(n17298), .B(n17297), .Z(n17374) );
  NANDN U17647 ( .A(n17300), .B(n17299), .Z(n17304) );
  OR U17648 ( .A(n17302), .B(n17301), .Z(n17303) );
  NAND U17649 ( .A(n17304), .B(n17303), .Z(n17441) );
  XNOR U17650 ( .A(n20052), .B(n17620), .Z(n17410) );
  OR U17651 ( .A(n17410), .B(n20020), .Z(n17307) );
  NANDN U17652 ( .A(n17305), .B(n19960), .Z(n17306) );
  NAND U17653 ( .A(n17307), .B(n17306), .Z(n17423) );
  XNOR U17654 ( .A(n102), .B(n17308), .Z(n17414) );
  OR U17655 ( .A(n17414), .B(n20121), .Z(n17311) );
  NANDN U17656 ( .A(n17309), .B(n20122), .Z(n17310) );
  NAND U17657 ( .A(n17311), .B(n17310), .Z(n17420) );
  XNOR U17658 ( .A(n19975), .B(n17776), .Z(n17417) );
  NANDN U17659 ( .A(n17417), .B(n19883), .Z(n17314) );
  NANDN U17660 ( .A(n17312), .B(n19937), .Z(n17313) );
  AND U17661 ( .A(n17314), .B(n17313), .Z(n17421) );
  XNOR U17662 ( .A(n17420), .B(n17421), .Z(n17422) );
  XNOR U17663 ( .A(n17423), .B(n17422), .Z(n17432) );
  NANDN U17664 ( .A(n17316), .B(n17315), .Z(n17320) );
  NAND U17665 ( .A(n17318), .B(n17317), .Z(n17319) );
  NAND U17666 ( .A(n17320), .B(n17319), .Z(n17433) );
  XNOR U17667 ( .A(n17432), .B(n17433), .Z(n17434) );
  NANDN U17668 ( .A(n17322), .B(n17321), .Z(n17326) );
  NAND U17669 ( .A(n17324), .B(n17323), .Z(n17325) );
  AND U17670 ( .A(n17326), .B(n17325), .Z(n17435) );
  XNOR U17671 ( .A(n17434), .B(n17435), .Z(n17379) );
  NANDN U17672 ( .A(n17328), .B(n17327), .Z(n17332) );
  OR U17673 ( .A(n17330), .B(n17329), .Z(n17331) );
  NAND U17674 ( .A(n17332), .B(n17331), .Z(n17407) );
  XNOR U17675 ( .A(n20154), .B(n17464), .Z(n17392) );
  OR U17676 ( .A(n17392), .B(n20057), .Z(n17335) );
  NANDN U17677 ( .A(n17333), .B(n20098), .Z(n17334) );
  AND U17678 ( .A(n17335), .B(n17334), .Z(n17384) );
  NAND U17679 ( .A(b[0]), .B(a[229]), .Z(n17336) );
  XNOR U17680 ( .A(b[1]), .B(n17336), .Z(n17338) );
  NAND U17681 ( .A(a[228]), .B(n98), .Z(n17337) );
  AND U17682 ( .A(n17338), .B(n17337), .Z(n17383) );
  XOR U17683 ( .A(n17384), .B(n17383), .Z(n17386) );
  NAND U17684 ( .A(a[213]), .B(b[15]), .Z(n17385) );
  XOR U17685 ( .A(n17386), .B(n17385), .Z(n17404) );
  NAND U17686 ( .A(n19722), .B(n17339), .Z(n17341) );
  XNOR U17687 ( .A(b[5]), .B(n18115), .Z(n17395) );
  NANDN U17688 ( .A(n19640), .B(n17395), .Z(n17340) );
  NAND U17689 ( .A(n17341), .B(n17340), .Z(n17429) );
  XNOR U17690 ( .A(n19714), .B(n17932), .Z(n17398) );
  NANDN U17691 ( .A(n17398), .B(n19766), .Z(n17344) );
  NANDN U17692 ( .A(n17342), .B(n19767), .Z(n17343) );
  NAND U17693 ( .A(n17344), .B(n17343), .Z(n17426) );
  NAND U17694 ( .A(n19554), .B(n17345), .Z(n17347) );
  IV U17695 ( .A(a[227]), .Z(n18244) );
  XNOR U17696 ( .A(b[3]), .B(n18244), .Z(n17401) );
  NANDN U17697 ( .A(n19521), .B(n17401), .Z(n17346) );
  AND U17698 ( .A(n17347), .B(n17346), .Z(n17427) );
  XNOR U17699 ( .A(n17426), .B(n17427), .Z(n17428) );
  XOR U17700 ( .A(n17429), .B(n17428), .Z(n17405) );
  XOR U17701 ( .A(n17404), .B(n17405), .Z(n17406) );
  XNOR U17702 ( .A(n17407), .B(n17406), .Z(n17377) );
  NAND U17703 ( .A(n17349), .B(n17348), .Z(n17353) );
  NAND U17704 ( .A(n17351), .B(n17350), .Z(n17352) );
  NAND U17705 ( .A(n17353), .B(n17352), .Z(n17378) );
  XOR U17706 ( .A(n17377), .B(n17378), .Z(n17380) );
  XNOR U17707 ( .A(n17379), .B(n17380), .Z(n17438) );
  NANDN U17708 ( .A(n17355), .B(n17354), .Z(n17359) );
  NAND U17709 ( .A(n17357), .B(n17356), .Z(n17358) );
  NAND U17710 ( .A(n17359), .B(n17358), .Z(n17439) );
  XNOR U17711 ( .A(n17438), .B(n17439), .Z(n17440) );
  XOR U17712 ( .A(n17441), .B(n17440), .Z(n17371) );
  NANDN U17713 ( .A(n17361), .B(n17360), .Z(n17365) );
  NANDN U17714 ( .A(n17363), .B(n17362), .Z(n17364) );
  NAND U17715 ( .A(n17365), .B(n17364), .Z(n17372) );
  XNOR U17716 ( .A(n17371), .B(n17372), .Z(n17373) );
  XNOR U17717 ( .A(n17374), .B(n17373), .Z(n17444) );
  XNOR U17718 ( .A(n17444), .B(sreg[469]), .Z(n17446) );
  NAND U17719 ( .A(n17366), .B(sreg[468]), .Z(n17370) );
  OR U17720 ( .A(n17368), .B(n17367), .Z(n17369) );
  AND U17721 ( .A(n17370), .B(n17369), .Z(n17445) );
  XOR U17722 ( .A(n17446), .B(n17445), .Z(c[469]) );
  NANDN U17723 ( .A(n17372), .B(n17371), .Z(n17376) );
  NAND U17724 ( .A(n17374), .B(n17373), .Z(n17375) );
  NAND U17725 ( .A(n17376), .B(n17375), .Z(n17452) );
  NANDN U17726 ( .A(n17378), .B(n17377), .Z(n17382) );
  OR U17727 ( .A(n17380), .B(n17379), .Z(n17381) );
  NAND U17728 ( .A(n17382), .B(n17381), .Z(n17519) );
  NANDN U17729 ( .A(n17384), .B(n17383), .Z(n17388) );
  OR U17730 ( .A(n17386), .B(n17385), .Z(n17387) );
  NAND U17731 ( .A(n17388), .B(n17387), .Z(n17507) );
  NAND U17732 ( .A(b[0]), .B(a[230]), .Z(n17389) );
  XNOR U17733 ( .A(b[1]), .B(n17389), .Z(n17391) );
  NAND U17734 ( .A(a[229]), .B(n98), .Z(n17390) );
  AND U17735 ( .A(n17391), .B(n17390), .Z(n17483) );
  XNOR U17736 ( .A(n20154), .B(n17542), .Z(n17492) );
  OR U17737 ( .A(n17492), .B(n20057), .Z(n17394) );
  NANDN U17738 ( .A(n17392), .B(n20098), .Z(n17393) );
  AND U17739 ( .A(n17394), .B(n17393), .Z(n17484) );
  XOR U17740 ( .A(n17483), .B(n17484), .Z(n17486) );
  NAND U17741 ( .A(a[214]), .B(b[15]), .Z(n17485) );
  XOR U17742 ( .A(n17486), .B(n17485), .Z(n17504) );
  NAND U17743 ( .A(n19722), .B(n17395), .Z(n17397) );
  XNOR U17744 ( .A(b[5]), .B(n18193), .Z(n17495) );
  NANDN U17745 ( .A(n19640), .B(n17495), .Z(n17396) );
  NAND U17746 ( .A(n17397), .B(n17396), .Z(n17480) );
  XNOR U17747 ( .A(n19714), .B(n18037), .Z(n17498) );
  NANDN U17748 ( .A(n17498), .B(n19766), .Z(n17400) );
  NANDN U17749 ( .A(n17398), .B(n19767), .Z(n17399) );
  NAND U17750 ( .A(n17400), .B(n17399), .Z(n17477) );
  NAND U17751 ( .A(n19554), .B(n17401), .Z(n17403) );
  IV U17752 ( .A(a[228]), .Z(n18322) );
  XNOR U17753 ( .A(b[3]), .B(n18322), .Z(n17501) );
  NANDN U17754 ( .A(n19521), .B(n17501), .Z(n17402) );
  AND U17755 ( .A(n17403), .B(n17402), .Z(n17478) );
  XNOR U17756 ( .A(n17477), .B(n17478), .Z(n17479) );
  XOR U17757 ( .A(n17480), .B(n17479), .Z(n17505) );
  XOR U17758 ( .A(n17504), .B(n17505), .Z(n17506) );
  XNOR U17759 ( .A(n17507), .B(n17506), .Z(n17455) );
  NAND U17760 ( .A(n17405), .B(n17404), .Z(n17409) );
  NAND U17761 ( .A(n17407), .B(n17406), .Z(n17408) );
  NAND U17762 ( .A(n17409), .B(n17408), .Z(n17456) );
  XOR U17763 ( .A(n17455), .B(n17456), .Z(n17458) );
  XNOR U17764 ( .A(n20052), .B(n17725), .Z(n17461) );
  OR U17765 ( .A(n17461), .B(n20020), .Z(n17412) );
  NANDN U17766 ( .A(n17410), .B(n19960), .Z(n17411) );
  NAND U17767 ( .A(n17412), .B(n17411), .Z(n17474) );
  XNOR U17768 ( .A(n102), .B(n17413), .Z(n17465) );
  OR U17769 ( .A(n17465), .B(n20121), .Z(n17416) );
  NANDN U17770 ( .A(n17414), .B(n20122), .Z(n17415) );
  NAND U17771 ( .A(n17416), .B(n17415), .Z(n17471) );
  XNOR U17772 ( .A(n19975), .B(n17854), .Z(n17468) );
  NANDN U17773 ( .A(n17468), .B(n19883), .Z(n17419) );
  NANDN U17774 ( .A(n17417), .B(n19937), .Z(n17418) );
  AND U17775 ( .A(n17419), .B(n17418), .Z(n17472) );
  XNOR U17776 ( .A(n17471), .B(n17472), .Z(n17473) );
  XNOR U17777 ( .A(n17474), .B(n17473), .Z(n17510) );
  NANDN U17778 ( .A(n17421), .B(n17420), .Z(n17425) );
  NAND U17779 ( .A(n17423), .B(n17422), .Z(n17424) );
  NAND U17780 ( .A(n17425), .B(n17424), .Z(n17511) );
  XNOR U17781 ( .A(n17510), .B(n17511), .Z(n17512) );
  NANDN U17782 ( .A(n17427), .B(n17426), .Z(n17431) );
  NAND U17783 ( .A(n17429), .B(n17428), .Z(n17430) );
  AND U17784 ( .A(n17431), .B(n17430), .Z(n17513) );
  XNOR U17785 ( .A(n17512), .B(n17513), .Z(n17457) );
  XNOR U17786 ( .A(n17458), .B(n17457), .Z(n17516) );
  NANDN U17787 ( .A(n17433), .B(n17432), .Z(n17437) );
  NAND U17788 ( .A(n17435), .B(n17434), .Z(n17436) );
  NAND U17789 ( .A(n17437), .B(n17436), .Z(n17517) );
  XNOR U17790 ( .A(n17516), .B(n17517), .Z(n17518) );
  XOR U17791 ( .A(n17519), .B(n17518), .Z(n17449) );
  NANDN U17792 ( .A(n17439), .B(n17438), .Z(n17443) );
  NANDN U17793 ( .A(n17441), .B(n17440), .Z(n17442) );
  NAND U17794 ( .A(n17443), .B(n17442), .Z(n17450) );
  XNOR U17795 ( .A(n17449), .B(n17450), .Z(n17451) );
  XNOR U17796 ( .A(n17452), .B(n17451), .Z(n17522) );
  XNOR U17797 ( .A(n17522), .B(sreg[470]), .Z(n17524) );
  NAND U17798 ( .A(n17444), .B(sreg[469]), .Z(n17448) );
  OR U17799 ( .A(n17446), .B(n17445), .Z(n17447) );
  AND U17800 ( .A(n17448), .B(n17447), .Z(n17523) );
  XOR U17801 ( .A(n17524), .B(n17523), .Z(c[470]) );
  NANDN U17802 ( .A(n17450), .B(n17449), .Z(n17454) );
  NAND U17803 ( .A(n17452), .B(n17451), .Z(n17453) );
  NAND U17804 ( .A(n17454), .B(n17453), .Z(n17530) );
  NANDN U17805 ( .A(n17456), .B(n17455), .Z(n17460) );
  OR U17806 ( .A(n17458), .B(n17457), .Z(n17459) );
  NAND U17807 ( .A(n17460), .B(n17459), .Z(n17597) );
  XNOR U17808 ( .A(n20052), .B(n17776), .Z(n17539) );
  OR U17809 ( .A(n17539), .B(n20020), .Z(n17463) );
  NANDN U17810 ( .A(n17461), .B(n19960), .Z(n17462) );
  NAND U17811 ( .A(n17463), .B(n17462), .Z(n17552) );
  XNOR U17812 ( .A(n102), .B(n17464), .Z(n17543) );
  OR U17813 ( .A(n17543), .B(n20121), .Z(n17467) );
  NANDN U17814 ( .A(n17465), .B(n20122), .Z(n17466) );
  NAND U17815 ( .A(n17467), .B(n17466), .Z(n17549) );
  XNOR U17816 ( .A(n19975), .B(n17932), .Z(n17546) );
  NANDN U17817 ( .A(n17546), .B(n19883), .Z(n17470) );
  NANDN U17818 ( .A(n17468), .B(n19937), .Z(n17469) );
  AND U17819 ( .A(n17470), .B(n17469), .Z(n17550) );
  XNOR U17820 ( .A(n17549), .B(n17550), .Z(n17551) );
  XNOR U17821 ( .A(n17552), .B(n17551), .Z(n17588) );
  NANDN U17822 ( .A(n17472), .B(n17471), .Z(n17476) );
  NAND U17823 ( .A(n17474), .B(n17473), .Z(n17475) );
  NAND U17824 ( .A(n17476), .B(n17475), .Z(n17589) );
  XNOR U17825 ( .A(n17588), .B(n17589), .Z(n17590) );
  NANDN U17826 ( .A(n17478), .B(n17477), .Z(n17482) );
  NAND U17827 ( .A(n17480), .B(n17479), .Z(n17481) );
  AND U17828 ( .A(n17482), .B(n17481), .Z(n17591) );
  XNOR U17829 ( .A(n17590), .B(n17591), .Z(n17535) );
  NANDN U17830 ( .A(n17484), .B(n17483), .Z(n17488) );
  OR U17831 ( .A(n17486), .B(n17485), .Z(n17487) );
  NAND U17832 ( .A(n17488), .B(n17487), .Z(n17585) );
  NAND U17833 ( .A(b[0]), .B(a[231]), .Z(n17489) );
  XNOR U17834 ( .A(b[1]), .B(n17489), .Z(n17491) );
  NAND U17835 ( .A(a[230]), .B(n98), .Z(n17490) );
  AND U17836 ( .A(n17491), .B(n17490), .Z(n17561) );
  XNOR U17837 ( .A(n20154), .B(n17620), .Z(n17570) );
  OR U17838 ( .A(n17570), .B(n20057), .Z(n17494) );
  NANDN U17839 ( .A(n17492), .B(n20098), .Z(n17493) );
  AND U17840 ( .A(n17494), .B(n17493), .Z(n17562) );
  XOR U17841 ( .A(n17561), .B(n17562), .Z(n17564) );
  NAND U17842 ( .A(a[215]), .B(b[15]), .Z(n17563) );
  XOR U17843 ( .A(n17564), .B(n17563), .Z(n17582) );
  NAND U17844 ( .A(n19722), .B(n17495), .Z(n17497) );
  XNOR U17845 ( .A(b[5]), .B(n18244), .Z(n17573) );
  NANDN U17846 ( .A(n19640), .B(n17573), .Z(n17496) );
  NAND U17847 ( .A(n17497), .B(n17496), .Z(n17558) );
  XNOR U17848 ( .A(n19714), .B(n18115), .Z(n17576) );
  NANDN U17849 ( .A(n17576), .B(n19766), .Z(n17500) );
  NANDN U17850 ( .A(n17498), .B(n19767), .Z(n17499) );
  NAND U17851 ( .A(n17500), .B(n17499), .Z(n17555) );
  NAND U17852 ( .A(n19554), .B(n17501), .Z(n17503) );
  IV U17853 ( .A(a[229]), .Z(n18427) );
  XNOR U17854 ( .A(b[3]), .B(n18427), .Z(n17579) );
  NANDN U17855 ( .A(n19521), .B(n17579), .Z(n17502) );
  AND U17856 ( .A(n17503), .B(n17502), .Z(n17556) );
  XNOR U17857 ( .A(n17555), .B(n17556), .Z(n17557) );
  XOR U17858 ( .A(n17558), .B(n17557), .Z(n17583) );
  XOR U17859 ( .A(n17582), .B(n17583), .Z(n17584) );
  XNOR U17860 ( .A(n17585), .B(n17584), .Z(n17533) );
  NAND U17861 ( .A(n17505), .B(n17504), .Z(n17509) );
  NAND U17862 ( .A(n17507), .B(n17506), .Z(n17508) );
  NAND U17863 ( .A(n17509), .B(n17508), .Z(n17534) );
  XOR U17864 ( .A(n17533), .B(n17534), .Z(n17536) );
  XNOR U17865 ( .A(n17535), .B(n17536), .Z(n17594) );
  NANDN U17866 ( .A(n17511), .B(n17510), .Z(n17515) );
  NAND U17867 ( .A(n17513), .B(n17512), .Z(n17514) );
  NAND U17868 ( .A(n17515), .B(n17514), .Z(n17595) );
  XNOR U17869 ( .A(n17594), .B(n17595), .Z(n17596) );
  XOR U17870 ( .A(n17597), .B(n17596), .Z(n17527) );
  NANDN U17871 ( .A(n17517), .B(n17516), .Z(n17521) );
  NANDN U17872 ( .A(n17519), .B(n17518), .Z(n17520) );
  NAND U17873 ( .A(n17521), .B(n17520), .Z(n17528) );
  XNOR U17874 ( .A(n17527), .B(n17528), .Z(n17529) );
  XNOR U17875 ( .A(n17530), .B(n17529), .Z(n17600) );
  XNOR U17876 ( .A(n17600), .B(sreg[471]), .Z(n17602) );
  NAND U17877 ( .A(n17522), .B(sreg[470]), .Z(n17526) );
  OR U17878 ( .A(n17524), .B(n17523), .Z(n17525) );
  AND U17879 ( .A(n17526), .B(n17525), .Z(n17601) );
  XOR U17880 ( .A(n17602), .B(n17601), .Z(c[471]) );
  NANDN U17881 ( .A(n17528), .B(n17527), .Z(n17532) );
  NAND U17882 ( .A(n17530), .B(n17529), .Z(n17531) );
  NAND U17883 ( .A(n17532), .B(n17531), .Z(n17608) );
  NANDN U17884 ( .A(n17534), .B(n17533), .Z(n17538) );
  OR U17885 ( .A(n17536), .B(n17535), .Z(n17537) );
  NAND U17886 ( .A(n17538), .B(n17537), .Z(n17675) );
  XNOR U17887 ( .A(n20052), .B(n17854), .Z(n17617) );
  OR U17888 ( .A(n17617), .B(n20020), .Z(n17541) );
  NANDN U17889 ( .A(n17539), .B(n19960), .Z(n17540) );
  NAND U17890 ( .A(n17541), .B(n17540), .Z(n17630) );
  XNOR U17891 ( .A(n102), .B(n17542), .Z(n17621) );
  OR U17892 ( .A(n17621), .B(n20121), .Z(n17545) );
  NANDN U17893 ( .A(n17543), .B(n20122), .Z(n17544) );
  NAND U17894 ( .A(n17545), .B(n17544), .Z(n17627) );
  XNOR U17895 ( .A(n19975), .B(n18037), .Z(n17624) );
  NANDN U17896 ( .A(n17624), .B(n19883), .Z(n17548) );
  NANDN U17897 ( .A(n17546), .B(n19937), .Z(n17547) );
  AND U17898 ( .A(n17548), .B(n17547), .Z(n17628) );
  XNOR U17899 ( .A(n17627), .B(n17628), .Z(n17629) );
  XNOR U17900 ( .A(n17630), .B(n17629), .Z(n17666) );
  NANDN U17901 ( .A(n17550), .B(n17549), .Z(n17554) );
  NAND U17902 ( .A(n17552), .B(n17551), .Z(n17553) );
  NAND U17903 ( .A(n17554), .B(n17553), .Z(n17667) );
  XNOR U17904 ( .A(n17666), .B(n17667), .Z(n17668) );
  NANDN U17905 ( .A(n17556), .B(n17555), .Z(n17560) );
  NAND U17906 ( .A(n17558), .B(n17557), .Z(n17559) );
  AND U17907 ( .A(n17560), .B(n17559), .Z(n17669) );
  XNOR U17908 ( .A(n17668), .B(n17669), .Z(n17613) );
  NANDN U17909 ( .A(n17562), .B(n17561), .Z(n17566) );
  OR U17910 ( .A(n17564), .B(n17563), .Z(n17565) );
  NAND U17911 ( .A(n17566), .B(n17565), .Z(n17663) );
  NAND U17912 ( .A(b[0]), .B(a[232]), .Z(n17567) );
  XNOR U17913 ( .A(b[1]), .B(n17567), .Z(n17569) );
  NAND U17914 ( .A(a[231]), .B(n98), .Z(n17568) );
  AND U17915 ( .A(n17569), .B(n17568), .Z(n17639) );
  XNOR U17916 ( .A(n20154), .B(n17725), .Z(n17648) );
  OR U17917 ( .A(n17648), .B(n20057), .Z(n17572) );
  NANDN U17918 ( .A(n17570), .B(n20098), .Z(n17571) );
  AND U17919 ( .A(n17572), .B(n17571), .Z(n17640) );
  XOR U17920 ( .A(n17639), .B(n17640), .Z(n17642) );
  NAND U17921 ( .A(a[216]), .B(b[15]), .Z(n17641) );
  XOR U17922 ( .A(n17642), .B(n17641), .Z(n17660) );
  NAND U17923 ( .A(n19722), .B(n17573), .Z(n17575) );
  XNOR U17924 ( .A(b[5]), .B(n18322), .Z(n17651) );
  NANDN U17925 ( .A(n19640), .B(n17651), .Z(n17574) );
  NAND U17926 ( .A(n17575), .B(n17574), .Z(n17636) );
  XNOR U17927 ( .A(n19714), .B(n18193), .Z(n17654) );
  NANDN U17928 ( .A(n17654), .B(n19766), .Z(n17578) );
  NANDN U17929 ( .A(n17576), .B(n19767), .Z(n17577) );
  NAND U17930 ( .A(n17578), .B(n17577), .Z(n17633) );
  NAND U17931 ( .A(n19554), .B(n17579), .Z(n17581) );
  IV U17932 ( .A(a[230]), .Z(n18505) );
  XNOR U17933 ( .A(b[3]), .B(n18505), .Z(n17657) );
  NANDN U17934 ( .A(n19521), .B(n17657), .Z(n17580) );
  AND U17935 ( .A(n17581), .B(n17580), .Z(n17634) );
  XNOR U17936 ( .A(n17633), .B(n17634), .Z(n17635) );
  XOR U17937 ( .A(n17636), .B(n17635), .Z(n17661) );
  XOR U17938 ( .A(n17660), .B(n17661), .Z(n17662) );
  XNOR U17939 ( .A(n17663), .B(n17662), .Z(n17611) );
  NAND U17940 ( .A(n17583), .B(n17582), .Z(n17587) );
  NAND U17941 ( .A(n17585), .B(n17584), .Z(n17586) );
  NAND U17942 ( .A(n17587), .B(n17586), .Z(n17612) );
  XOR U17943 ( .A(n17611), .B(n17612), .Z(n17614) );
  XNOR U17944 ( .A(n17613), .B(n17614), .Z(n17672) );
  NANDN U17945 ( .A(n17589), .B(n17588), .Z(n17593) );
  NAND U17946 ( .A(n17591), .B(n17590), .Z(n17592) );
  NAND U17947 ( .A(n17593), .B(n17592), .Z(n17673) );
  XNOR U17948 ( .A(n17672), .B(n17673), .Z(n17674) );
  XOR U17949 ( .A(n17675), .B(n17674), .Z(n17605) );
  NANDN U17950 ( .A(n17595), .B(n17594), .Z(n17599) );
  NANDN U17951 ( .A(n17597), .B(n17596), .Z(n17598) );
  NAND U17952 ( .A(n17599), .B(n17598), .Z(n17606) );
  XNOR U17953 ( .A(n17605), .B(n17606), .Z(n17607) );
  XNOR U17954 ( .A(n17608), .B(n17607), .Z(n17678) );
  XNOR U17955 ( .A(n17678), .B(sreg[472]), .Z(n17680) );
  NAND U17956 ( .A(n17600), .B(sreg[471]), .Z(n17604) );
  OR U17957 ( .A(n17602), .B(n17601), .Z(n17603) );
  AND U17958 ( .A(n17604), .B(n17603), .Z(n17679) );
  XOR U17959 ( .A(n17680), .B(n17679), .Z(c[472]) );
  NANDN U17960 ( .A(n17606), .B(n17605), .Z(n17610) );
  NAND U17961 ( .A(n17608), .B(n17607), .Z(n17609) );
  NAND U17962 ( .A(n17610), .B(n17609), .Z(n17686) );
  NANDN U17963 ( .A(n17612), .B(n17611), .Z(n17616) );
  OR U17964 ( .A(n17614), .B(n17613), .Z(n17615) );
  NAND U17965 ( .A(n17616), .B(n17615), .Z(n17753) );
  XNOR U17966 ( .A(n20052), .B(n17932), .Z(n17722) );
  OR U17967 ( .A(n17722), .B(n20020), .Z(n17619) );
  NANDN U17968 ( .A(n17617), .B(n19960), .Z(n17618) );
  NAND U17969 ( .A(n17619), .B(n17618), .Z(n17735) );
  XNOR U17970 ( .A(n102), .B(n17620), .Z(n17726) );
  OR U17971 ( .A(n17726), .B(n20121), .Z(n17623) );
  NANDN U17972 ( .A(n17621), .B(n20122), .Z(n17622) );
  NAND U17973 ( .A(n17623), .B(n17622), .Z(n17732) );
  XNOR U17974 ( .A(n19975), .B(n18115), .Z(n17729) );
  NANDN U17975 ( .A(n17729), .B(n19883), .Z(n17626) );
  NANDN U17976 ( .A(n17624), .B(n19937), .Z(n17625) );
  AND U17977 ( .A(n17626), .B(n17625), .Z(n17733) );
  XNOR U17978 ( .A(n17732), .B(n17733), .Z(n17734) );
  XNOR U17979 ( .A(n17735), .B(n17734), .Z(n17744) );
  NANDN U17980 ( .A(n17628), .B(n17627), .Z(n17632) );
  NAND U17981 ( .A(n17630), .B(n17629), .Z(n17631) );
  NAND U17982 ( .A(n17632), .B(n17631), .Z(n17745) );
  XNOR U17983 ( .A(n17744), .B(n17745), .Z(n17746) );
  NANDN U17984 ( .A(n17634), .B(n17633), .Z(n17638) );
  NAND U17985 ( .A(n17636), .B(n17635), .Z(n17637) );
  AND U17986 ( .A(n17638), .B(n17637), .Z(n17747) );
  XNOR U17987 ( .A(n17746), .B(n17747), .Z(n17691) );
  NANDN U17988 ( .A(n17640), .B(n17639), .Z(n17644) );
  OR U17989 ( .A(n17642), .B(n17641), .Z(n17643) );
  NAND U17990 ( .A(n17644), .B(n17643), .Z(n17719) );
  NAND U17991 ( .A(b[0]), .B(a[233]), .Z(n17645) );
  XNOR U17992 ( .A(b[1]), .B(n17645), .Z(n17647) );
  NAND U17993 ( .A(a[232]), .B(n98), .Z(n17646) );
  AND U17994 ( .A(n17647), .B(n17646), .Z(n17695) );
  XNOR U17995 ( .A(n20154), .B(n17776), .Z(n17701) );
  OR U17996 ( .A(n17701), .B(n20057), .Z(n17650) );
  NANDN U17997 ( .A(n17648), .B(n20098), .Z(n17649) );
  AND U17998 ( .A(n17650), .B(n17649), .Z(n17696) );
  XOR U17999 ( .A(n17695), .B(n17696), .Z(n17698) );
  NAND U18000 ( .A(a[217]), .B(b[15]), .Z(n17697) );
  XOR U18001 ( .A(n17698), .B(n17697), .Z(n17716) );
  NAND U18002 ( .A(n19722), .B(n17651), .Z(n17653) );
  XNOR U18003 ( .A(b[5]), .B(n18427), .Z(n17707) );
  NANDN U18004 ( .A(n19640), .B(n17707), .Z(n17652) );
  NAND U18005 ( .A(n17653), .B(n17652), .Z(n17741) );
  XNOR U18006 ( .A(n19714), .B(n18244), .Z(n17710) );
  NANDN U18007 ( .A(n17710), .B(n19766), .Z(n17656) );
  NANDN U18008 ( .A(n17654), .B(n19767), .Z(n17655) );
  NAND U18009 ( .A(n17656), .B(n17655), .Z(n17738) );
  NAND U18010 ( .A(n19554), .B(n17657), .Z(n17659) );
  IV U18011 ( .A(a[231]), .Z(n18556) );
  XNOR U18012 ( .A(b[3]), .B(n18556), .Z(n17713) );
  NANDN U18013 ( .A(n19521), .B(n17713), .Z(n17658) );
  AND U18014 ( .A(n17659), .B(n17658), .Z(n17739) );
  XNOR U18015 ( .A(n17738), .B(n17739), .Z(n17740) );
  XOR U18016 ( .A(n17741), .B(n17740), .Z(n17717) );
  XOR U18017 ( .A(n17716), .B(n17717), .Z(n17718) );
  XNOR U18018 ( .A(n17719), .B(n17718), .Z(n17689) );
  NAND U18019 ( .A(n17661), .B(n17660), .Z(n17665) );
  NAND U18020 ( .A(n17663), .B(n17662), .Z(n17664) );
  NAND U18021 ( .A(n17665), .B(n17664), .Z(n17690) );
  XOR U18022 ( .A(n17689), .B(n17690), .Z(n17692) );
  XNOR U18023 ( .A(n17691), .B(n17692), .Z(n17750) );
  NANDN U18024 ( .A(n17667), .B(n17666), .Z(n17671) );
  NAND U18025 ( .A(n17669), .B(n17668), .Z(n17670) );
  NAND U18026 ( .A(n17671), .B(n17670), .Z(n17751) );
  XNOR U18027 ( .A(n17750), .B(n17751), .Z(n17752) );
  XOR U18028 ( .A(n17753), .B(n17752), .Z(n17683) );
  NANDN U18029 ( .A(n17673), .B(n17672), .Z(n17677) );
  NANDN U18030 ( .A(n17675), .B(n17674), .Z(n17676) );
  NAND U18031 ( .A(n17677), .B(n17676), .Z(n17684) );
  XNOR U18032 ( .A(n17683), .B(n17684), .Z(n17685) );
  XNOR U18033 ( .A(n17686), .B(n17685), .Z(n17756) );
  XNOR U18034 ( .A(n17756), .B(sreg[473]), .Z(n17758) );
  NAND U18035 ( .A(n17678), .B(sreg[472]), .Z(n17682) );
  OR U18036 ( .A(n17680), .B(n17679), .Z(n17681) );
  AND U18037 ( .A(n17682), .B(n17681), .Z(n17757) );
  XOR U18038 ( .A(n17758), .B(n17757), .Z(c[473]) );
  NANDN U18039 ( .A(n17684), .B(n17683), .Z(n17688) );
  NAND U18040 ( .A(n17686), .B(n17685), .Z(n17687) );
  NAND U18041 ( .A(n17688), .B(n17687), .Z(n17764) );
  NANDN U18042 ( .A(n17690), .B(n17689), .Z(n17694) );
  OR U18043 ( .A(n17692), .B(n17691), .Z(n17693) );
  NAND U18044 ( .A(n17694), .B(n17693), .Z(n17831) );
  NANDN U18045 ( .A(n17696), .B(n17695), .Z(n17700) );
  OR U18046 ( .A(n17698), .B(n17697), .Z(n17699) );
  NAND U18047 ( .A(n17700), .B(n17699), .Z(n17819) );
  XNOR U18048 ( .A(n20154), .B(n17854), .Z(n17804) );
  OR U18049 ( .A(n17804), .B(n20057), .Z(n17703) );
  NANDN U18050 ( .A(n17701), .B(n20098), .Z(n17702) );
  AND U18051 ( .A(n17703), .B(n17702), .Z(n17796) );
  NAND U18052 ( .A(b[0]), .B(a[234]), .Z(n17704) );
  XNOR U18053 ( .A(b[1]), .B(n17704), .Z(n17706) );
  NAND U18054 ( .A(a[233]), .B(n98), .Z(n17705) );
  AND U18055 ( .A(n17706), .B(n17705), .Z(n17795) );
  XOR U18056 ( .A(n17796), .B(n17795), .Z(n17798) );
  NAND U18057 ( .A(a[218]), .B(b[15]), .Z(n17797) );
  XOR U18058 ( .A(n17798), .B(n17797), .Z(n17816) );
  NAND U18059 ( .A(n19722), .B(n17707), .Z(n17709) );
  XNOR U18060 ( .A(b[5]), .B(n18505), .Z(n17807) );
  NANDN U18061 ( .A(n19640), .B(n17807), .Z(n17708) );
  NAND U18062 ( .A(n17709), .B(n17708), .Z(n17792) );
  XNOR U18063 ( .A(n19714), .B(n18322), .Z(n17810) );
  NANDN U18064 ( .A(n17810), .B(n19766), .Z(n17712) );
  NANDN U18065 ( .A(n17710), .B(n19767), .Z(n17711) );
  NAND U18066 ( .A(n17712), .B(n17711), .Z(n17789) );
  NAND U18067 ( .A(n19554), .B(n17713), .Z(n17715) );
  IV U18068 ( .A(a[232]), .Z(n18661) );
  XNOR U18069 ( .A(b[3]), .B(n18661), .Z(n17813) );
  NANDN U18070 ( .A(n19521), .B(n17813), .Z(n17714) );
  AND U18071 ( .A(n17715), .B(n17714), .Z(n17790) );
  XNOR U18072 ( .A(n17789), .B(n17790), .Z(n17791) );
  XOR U18073 ( .A(n17792), .B(n17791), .Z(n17817) );
  XOR U18074 ( .A(n17816), .B(n17817), .Z(n17818) );
  XNOR U18075 ( .A(n17819), .B(n17818), .Z(n17767) );
  NAND U18076 ( .A(n17717), .B(n17716), .Z(n17721) );
  NAND U18077 ( .A(n17719), .B(n17718), .Z(n17720) );
  NAND U18078 ( .A(n17721), .B(n17720), .Z(n17768) );
  XOR U18079 ( .A(n17767), .B(n17768), .Z(n17770) );
  XNOR U18080 ( .A(n20052), .B(n18037), .Z(n17773) );
  OR U18081 ( .A(n17773), .B(n20020), .Z(n17724) );
  NANDN U18082 ( .A(n17722), .B(n19960), .Z(n17723) );
  NAND U18083 ( .A(n17724), .B(n17723), .Z(n17786) );
  XNOR U18084 ( .A(n102), .B(n17725), .Z(n17777) );
  OR U18085 ( .A(n17777), .B(n20121), .Z(n17728) );
  NANDN U18086 ( .A(n17726), .B(n20122), .Z(n17727) );
  NAND U18087 ( .A(n17728), .B(n17727), .Z(n17783) );
  XNOR U18088 ( .A(n19975), .B(n18193), .Z(n17780) );
  NANDN U18089 ( .A(n17780), .B(n19883), .Z(n17731) );
  NANDN U18090 ( .A(n17729), .B(n19937), .Z(n17730) );
  AND U18091 ( .A(n17731), .B(n17730), .Z(n17784) );
  XNOR U18092 ( .A(n17783), .B(n17784), .Z(n17785) );
  XNOR U18093 ( .A(n17786), .B(n17785), .Z(n17822) );
  NANDN U18094 ( .A(n17733), .B(n17732), .Z(n17737) );
  NAND U18095 ( .A(n17735), .B(n17734), .Z(n17736) );
  NAND U18096 ( .A(n17737), .B(n17736), .Z(n17823) );
  XNOR U18097 ( .A(n17822), .B(n17823), .Z(n17824) );
  NANDN U18098 ( .A(n17739), .B(n17738), .Z(n17743) );
  NAND U18099 ( .A(n17741), .B(n17740), .Z(n17742) );
  AND U18100 ( .A(n17743), .B(n17742), .Z(n17825) );
  XNOR U18101 ( .A(n17824), .B(n17825), .Z(n17769) );
  XNOR U18102 ( .A(n17770), .B(n17769), .Z(n17828) );
  NANDN U18103 ( .A(n17745), .B(n17744), .Z(n17749) );
  NAND U18104 ( .A(n17747), .B(n17746), .Z(n17748) );
  NAND U18105 ( .A(n17749), .B(n17748), .Z(n17829) );
  XNOR U18106 ( .A(n17828), .B(n17829), .Z(n17830) );
  XOR U18107 ( .A(n17831), .B(n17830), .Z(n17761) );
  NANDN U18108 ( .A(n17751), .B(n17750), .Z(n17755) );
  NANDN U18109 ( .A(n17753), .B(n17752), .Z(n17754) );
  NAND U18110 ( .A(n17755), .B(n17754), .Z(n17762) );
  XNOR U18111 ( .A(n17761), .B(n17762), .Z(n17763) );
  XNOR U18112 ( .A(n17764), .B(n17763), .Z(n17834) );
  XNOR U18113 ( .A(n17834), .B(sreg[474]), .Z(n17836) );
  NAND U18114 ( .A(n17756), .B(sreg[473]), .Z(n17760) );
  OR U18115 ( .A(n17758), .B(n17757), .Z(n17759) );
  AND U18116 ( .A(n17760), .B(n17759), .Z(n17835) );
  XOR U18117 ( .A(n17836), .B(n17835), .Z(c[474]) );
  NANDN U18118 ( .A(n17762), .B(n17761), .Z(n17766) );
  NAND U18119 ( .A(n17764), .B(n17763), .Z(n17765) );
  NAND U18120 ( .A(n17766), .B(n17765), .Z(n17842) );
  NANDN U18121 ( .A(n17768), .B(n17767), .Z(n17772) );
  OR U18122 ( .A(n17770), .B(n17769), .Z(n17771) );
  NAND U18123 ( .A(n17772), .B(n17771), .Z(n17909) );
  XNOR U18124 ( .A(n20052), .B(n18115), .Z(n17851) );
  OR U18125 ( .A(n17851), .B(n20020), .Z(n17775) );
  NANDN U18126 ( .A(n17773), .B(n19960), .Z(n17774) );
  NAND U18127 ( .A(n17775), .B(n17774), .Z(n17864) );
  XNOR U18128 ( .A(n102), .B(n17776), .Z(n17855) );
  OR U18129 ( .A(n17855), .B(n20121), .Z(n17779) );
  NANDN U18130 ( .A(n17777), .B(n20122), .Z(n17778) );
  NAND U18131 ( .A(n17779), .B(n17778), .Z(n17861) );
  XNOR U18132 ( .A(n19975), .B(n18244), .Z(n17858) );
  NANDN U18133 ( .A(n17858), .B(n19883), .Z(n17782) );
  NANDN U18134 ( .A(n17780), .B(n19937), .Z(n17781) );
  AND U18135 ( .A(n17782), .B(n17781), .Z(n17862) );
  XNOR U18136 ( .A(n17861), .B(n17862), .Z(n17863) );
  XNOR U18137 ( .A(n17864), .B(n17863), .Z(n17900) );
  NANDN U18138 ( .A(n17784), .B(n17783), .Z(n17788) );
  NAND U18139 ( .A(n17786), .B(n17785), .Z(n17787) );
  NAND U18140 ( .A(n17788), .B(n17787), .Z(n17901) );
  XNOR U18141 ( .A(n17900), .B(n17901), .Z(n17902) );
  NANDN U18142 ( .A(n17790), .B(n17789), .Z(n17794) );
  NAND U18143 ( .A(n17792), .B(n17791), .Z(n17793) );
  AND U18144 ( .A(n17794), .B(n17793), .Z(n17903) );
  XNOR U18145 ( .A(n17902), .B(n17903), .Z(n17847) );
  NANDN U18146 ( .A(n17796), .B(n17795), .Z(n17800) );
  OR U18147 ( .A(n17798), .B(n17797), .Z(n17799) );
  NAND U18148 ( .A(n17800), .B(n17799), .Z(n17897) );
  NAND U18149 ( .A(b[0]), .B(a[235]), .Z(n17801) );
  XNOR U18150 ( .A(b[1]), .B(n17801), .Z(n17803) );
  NAND U18151 ( .A(a[234]), .B(n98), .Z(n17802) );
  AND U18152 ( .A(n17803), .B(n17802), .Z(n17873) );
  XNOR U18153 ( .A(n20154), .B(n17932), .Z(n17879) );
  OR U18154 ( .A(n17879), .B(n20057), .Z(n17806) );
  NANDN U18155 ( .A(n17804), .B(n20098), .Z(n17805) );
  AND U18156 ( .A(n17806), .B(n17805), .Z(n17874) );
  XOR U18157 ( .A(n17873), .B(n17874), .Z(n17876) );
  NAND U18158 ( .A(a[219]), .B(b[15]), .Z(n17875) );
  XOR U18159 ( .A(n17876), .B(n17875), .Z(n17894) );
  NAND U18160 ( .A(n19722), .B(n17807), .Z(n17809) );
  XNOR U18161 ( .A(b[5]), .B(n18556), .Z(n17885) );
  NANDN U18162 ( .A(n19640), .B(n17885), .Z(n17808) );
  NAND U18163 ( .A(n17809), .B(n17808), .Z(n17870) );
  XNOR U18164 ( .A(n19714), .B(n18427), .Z(n17888) );
  NANDN U18165 ( .A(n17888), .B(n19766), .Z(n17812) );
  NANDN U18166 ( .A(n17810), .B(n19767), .Z(n17811) );
  NAND U18167 ( .A(n17812), .B(n17811), .Z(n17867) );
  NAND U18168 ( .A(n19554), .B(n17813), .Z(n17815) );
  IV U18169 ( .A(a[233]), .Z(n18712) );
  XNOR U18170 ( .A(b[3]), .B(n18712), .Z(n17891) );
  NANDN U18171 ( .A(n19521), .B(n17891), .Z(n17814) );
  AND U18172 ( .A(n17815), .B(n17814), .Z(n17868) );
  XNOR U18173 ( .A(n17867), .B(n17868), .Z(n17869) );
  XOR U18174 ( .A(n17870), .B(n17869), .Z(n17895) );
  XOR U18175 ( .A(n17894), .B(n17895), .Z(n17896) );
  XNOR U18176 ( .A(n17897), .B(n17896), .Z(n17845) );
  NAND U18177 ( .A(n17817), .B(n17816), .Z(n17821) );
  NAND U18178 ( .A(n17819), .B(n17818), .Z(n17820) );
  NAND U18179 ( .A(n17821), .B(n17820), .Z(n17846) );
  XOR U18180 ( .A(n17845), .B(n17846), .Z(n17848) );
  XNOR U18181 ( .A(n17847), .B(n17848), .Z(n17906) );
  NANDN U18182 ( .A(n17823), .B(n17822), .Z(n17827) );
  NAND U18183 ( .A(n17825), .B(n17824), .Z(n17826) );
  NAND U18184 ( .A(n17827), .B(n17826), .Z(n17907) );
  XNOR U18185 ( .A(n17906), .B(n17907), .Z(n17908) );
  XOR U18186 ( .A(n17909), .B(n17908), .Z(n17839) );
  NANDN U18187 ( .A(n17829), .B(n17828), .Z(n17833) );
  NANDN U18188 ( .A(n17831), .B(n17830), .Z(n17832) );
  NAND U18189 ( .A(n17833), .B(n17832), .Z(n17840) );
  XNOR U18190 ( .A(n17839), .B(n17840), .Z(n17841) );
  XNOR U18191 ( .A(n17842), .B(n17841), .Z(n17912) );
  XNOR U18192 ( .A(n17912), .B(sreg[475]), .Z(n17914) );
  NAND U18193 ( .A(n17834), .B(sreg[474]), .Z(n17838) );
  OR U18194 ( .A(n17836), .B(n17835), .Z(n17837) );
  AND U18195 ( .A(n17838), .B(n17837), .Z(n17913) );
  XOR U18196 ( .A(n17914), .B(n17913), .Z(c[475]) );
  NANDN U18197 ( .A(n17840), .B(n17839), .Z(n17844) );
  NAND U18198 ( .A(n17842), .B(n17841), .Z(n17843) );
  NAND U18199 ( .A(n17844), .B(n17843), .Z(n17920) );
  NANDN U18200 ( .A(n17846), .B(n17845), .Z(n17850) );
  OR U18201 ( .A(n17848), .B(n17847), .Z(n17849) );
  NAND U18202 ( .A(n17850), .B(n17849), .Z(n17987) );
  XNOR U18203 ( .A(n20052), .B(n18193), .Z(n17929) );
  OR U18204 ( .A(n17929), .B(n20020), .Z(n17853) );
  NANDN U18205 ( .A(n17851), .B(n19960), .Z(n17852) );
  NAND U18206 ( .A(n17853), .B(n17852), .Z(n17942) );
  XNOR U18207 ( .A(n102), .B(n17854), .Z(n17933) );
  OR U18208 ( .A(n17933), .B(n20121), .Z(n17857) );
  NANDN U18209 ( .A(n17855), .B(n20122), .Z(n17856) );
  NAND U18210 ( .A(n17857), .B(n17856), .Z(n17939) );
  XNOR U18211 ( .A(n19975), .B(n18322), .Z(n17936) );
  NANDN U18212 ( .A(n17936), .B(n19883), .Z(n17860) );
  NANDN U18213 ( .A(n17858), .B(n19937), .Z(n17859) );
  AND U18214 ( .A(n17860), .B(n17859), .Z(n17940) );
  XNOR U18215 ( .A(n17939), .B(n17940), .Z(n17941) );
  XNOR U18216 ( .A(n17942), .B(n17941), .Z(n17978) );
  NANDN U18217 ( .A(n17862), .B(n17861), .Z(n17866) );
  NAND U18218 ( .A(n17864), .B(n17863), .Z(n17865) );
  NAND U18219 ( .A(n17866), .B(n17865), .Z(n17979) );
  XNOR U18220 ( .A(n17978), .B(n17979), .Z(n17980) );
  NANDN U18221 ( .A(n17868), .B(n17867), .Z(n17872) );
  NAND U18222 ( .A(n17870), .B(n17869), .Z(n17871) );
  AND U18223 ( .A(n17872), .B(n17871), .Z(n17981) );
  XNOR U18224 ( .A(n17980), .B(n17981), .Z(n17925) );
  NANDN U18225 ( .A(n17874), .B(n17873), .Z(n17878) );
  OR U18226 ( .A(n17876), .B(n17875), .Z(n17877) );
  NAND U18227 ( .A(n17878), .B(n17877), .Z(n17975) );
  XNOR U18228 ( .A(n20154), .B(n18037), .Z(n17960) );
  OR U18229 ( .A(n17960), .B(n20057), .Z(n17881) );
  NANDN U18230 ( .A(n17879), .B(n20098), .Z(n17880) );
  AND U18231 ( .A(n17881), .B(n17880), .Z(n17952) );
  NAND U18232 ( .A(b[0]), .B(a[236]), .Z(n17882) );
  XNOR U18233 ( .A(b[1]), .B(n17882), .Z(n17884) );
  NAND U18234 ( .A(a[235]), .B(n98), .Z(n17883) );
  AND U18235 ( .A(n17884), .B(n17883), .Z(n17951) );
  XOR U18236 ( .A(n17952), .B(n17951), .Z(n17954) );
  NAND U18237 ( .A(a[220]), .B(b[15]), .Z(n17953) );
  XOR U18238 ( .A(n17954), .B(n17953), .Z(n17972) );
  NAND U18239 ( .A(n19722), .B(n17885), .Z(n17887) );
  XNOR U18240 ( .A(b[5]), .B(n18661), .Z(n17963) );
  NANDN U18241 ( .A(n19640), .B(n17963), .Z(n17886) );
  NAND U18242 ( .A(n17887), .B(n17886), .Z(n17948) );
  XNOR U18243 ( .A(n19714), .B(n18505), .Z(n17966) );
  NANDN U18244 ( .A(n17966), .B(n19766), .Z(n17890) );
  NANDN U18245 ( .A(n17888), .B(n19767), .Z(n17889) );
  NAND U18246 ( .A(n17890), .B(n17889), .Z(n17945) );
  NAND U18247 ( .A(n19554), .B(n17891), .Z(n17893) );
  IV U18248 ( .A(a[234]), .Z(n18790) );
  XNOR U18249 ( .A(b[3]), .B(n18790), .Z(n17969) );
  NANDN U18250 ( .A(n19521), .B(n17969), .Z(n17892) );
  AND U18251 ( .A(n17893), .B(n17892), .Z(n17946) );
  XNOR U18252 ( .A(n17945), .B(n17946), .Z(n17947) );
  XOR U18253 ( .A(n17948), .B(n17947), .Z(n17973) );
  XOR U18254 ( .A(n17972), .B(n17973), .Z(n17974) );
  XNOR U18255 ( .A(n17975), .B(n17974), .Z(n17923) );
  NAND U18256 ( .A(n17895), .B(n17894), .Z(n17899) );
  NAND U18257 ( .A(n17897), .B(n17896), .Z(n17898) );
  NAND U18258 ( .A(n17899), .B(n17898), .Z(n17924) );
  XOR U18259 ( .A(n17923), .B(n17924), .Z(n17926) );
  XNOR U18260 ( .A(n17925), .B(n17926), .Z(n17984) );
  NANDN U18261 ( .A(n17901), .B(n17900), .Z(n17905) );
  NAND U18262 ( .A(n17903), .B(n17902), .Z(n17904) );
  NAND U18263 ( .A(n17905), .B(n17904), .Z(n17985) );
  XNOR U18264 ( .A(n17984), .B(n17985), .Z(n17986) );
  XOR U18265 ( .A(n17987), .B(n17986), .Z(n17917) );
  NANDN U18266 ( .A(n17907), .B(n17906), .Z(n17911) );
  NANDN U18267 ( .A(n17909), .B(n17908), .Z(n17910) );
  NAND U18268 ( .A(n17911), .B(n17910), .Z(n17918) );
  XNOR U18269 ( .A(n17917), .B(n17918), .Z(n17919) );
  XNOR U18270 ( .A(n17920), .B(n17919), .Z(n17990) );
  XNOR U18271 ( .A(n17990), .B(sreg[476]), .Z(n17992) );
  NAND U18272 ( .A(n17912), .B(sreg[475]), .Z(n17916) );
  OR U18273 ( .A(n17914), .B(n17913), .Z(n17915) );
  AND U18274 ( .A(n17916), .B(n17915), .Z(n17991) );
  XOR U18275 ( .A(n17992), .B(n17991), .Z(c[476]) );
  NANDN U18276 ( .A(n17918), .B(n17917), .Z(n17922) );
  NAND U18277 ( .A(n17920), .B(n17919), .Z(n17921) );
  NAND U18278 ( .A(n17922), .B(n17921), .Z(n17998) );
  NANDN U18279 ( .A(n17924), .B(n17923), .Z(n17928) );
  OR U18280 ( .A(n17926), .B(n17925), .Z(n17927) );
  NAND U18281 ( .A(n17928), .B(n17927), .Z(n18065) );
  XNOR U18282 ( .A(n20052), .B(n18244), .Z(n18034) );
  OR U18283 ( .A(n18034), .B(n20020), .Z(n17931) );
  NANDN U18284 ( .A(n17929), .B(n19960), .Z(n17930) );
  NAND U18285 ( .A(n17931), .B(n17930), .Z(n18047) );
  XNOR U18286 ( .A(n102), .B(n17932), .Z(n18038) );
  OR U18287 ( .A(n18038), .B(n20121), .Z(n17935) );
  NANDN U18288 ( .A(n17933), .B(n20122), .Z(n17934) );
  NAND U18289 ( .A(n17935), .B(n17934), .Z(n18044) );
  XNOR U18290 ( .A(n19975), .B(n18427), .Z(n18041) );
  NANDN U18291 ( .A(n18041), .B(n19883), .Z(n17938) );
  NANDN U18292 ( .A(n17936), .B(n19937), .Z(n17937) );
  AND U18293 ( .A(n17938), .B(n17937), .Z(n18045) );
  XNOR U18294 ( .A(n18044), .B(n18045), .Z(n18046) );
  XNOR U18295 ( .A(n18047), .B(n18046), .Z(n18056) );
  NANDN U18296 ( .A(n17940), .B(n17939), .Z(n17944) );
  NAND U18297 ( .A(n17942), .B(n17941), .Z(n17943) );
  NAND U18298 ( .A(n17944), .B(n17943), .Z(n18057) );
  XNOR U18299 ( .A(n18056), .B(n18057), .Z(n18058) );
  NANDN U18300 ( .A(n17946), .B(n17945), .Z(n17950) );
  NAND U18301 ( .A(n17948), .B(n17947), .Z(n17949) );
  AND U18302 ( .A(n17950), .B(n17949), .Z(n18059) );
  XNOR U18303 ( .A(n18058), .B(n18059), .Z(n18003) );
  NANDN U18304 ( .A(n17952), .B(n17951), .Z(n17956) );
  OR U18305 ( .A(n17954), .B(n17953), .Z(n17955) );
  NAND U18306 ( .A(n17956), .B(n17955), .Z(n18031) );
  NAND U18307 ( .A(b[0]), .B(a[237]), .Z(n17957) );
  XNOR U18308 ( .A(b[1]), .B(n17957), .Z(n17959) );
  NAND U18309 ( .A(a[236]), .B(n98), .Z(n17958) );
  AND U18310 ( .A(n17959), .B(n17958), .Z(n18007) );
  XNOR U18311 ( .A(n20154), .B(n18115), .Z(n18016) );
  OR U18312 ( .A(n18016), .B(n20057), .Z(n17962) );
  NANDN U18313 ( .A(n17960), .B(n20098), .Z(n17961) );
  AND U18314 ( .A(n17962), .B(n17961), .Z(n18008) );
  XOR U18315 ( .A(n18007), .B(n18008), .Z(n18010) );
  NAND U18316 ( .A(a[221]), .B(b[15]), .Z(n18009) );
  XOR U18317 ( .A(n18010), .B(n18009), .Z(n18028) );
  NAND U18318 ( .A(n19722), .B(n17963), .Z(n17965) );
  XNOR U18319 ( .A(b[5]), .B(n18712), .Z(n18019) );
  NANDN U18320 ( .A(n19640), .B(n18019), .Z(n17964) );
  NAND U18321 ( .A(n17965), .B(n17964), .Z(n18053) );
  XNOR U18322 ( .A(n19714), .B(n18556), .Z(n18022) );
  NANDN U18323 ( .A(n18022), .B(n19766), .Z(n17968) );
  NANDN U18324 ( .A(n17966), .B(n19767), .Z(n17967) );
  NAND U18325 ( .A(n17968), .B(n17967), .Z(n18050) );
  NAND U18326 ( .A(n19554), .B(n17969), .Z(n17971) );
  IV U18327 ( .A(a[235]), .Z(n18868) );
  XNOR U18328 ( .A(b[3]), .B(n18868), .Z(n18025) );
  NANDN U18329 ( .A(n19521), .B(n18025), .Z(n17970) );
  AND U18330 ( .A(n17971), .B(n17970), .Z(n18051) );
  XNOR U18331 ( .A(n18050), .B(n18051), .Z(n18052) );
  XOR U18332 ( .A(n18053), .B(n18052), .Z(n18029) );
  XOR U18333 ( .A(n18028), .B(n18029), .Z(n18030) );
  XNOR U18334 ( .A(n18031), .B(n18030), .Z(n18001) );
  NAND U18335 ( .A(n17973), .B(n17972), .Z(n17977) );
  NAND U18336 ( .A(n17975), .B(n17974), .Z(n17976) );
  NAND U18337 ( .A(n17977), .B(n17976), .Z(n18002) );
  XOR U18338 ( .A(n18001), .B(n18002), .Z(n18004) );
  XNOR U18339 ( .A(n18003), .B(n18004), .Z(n18062) );
  NANDN U18340 ( .A(n17979), .B(n17978), .Z(n17983) );
  NAND U18341 ( .A(n17981), .B(n17980), .Z(n17982) );
  NAND U18342 ( .A(n17983), .B(n17982), .Z(n18063) );
  XNOR U18343 ( .A(n18062), .B(n18063), .Z(n18064) );
  XOR U18344 ( .A(n18065), .B(n18064), .Z(n17995) );
  NANDN U18345 ( .A(n17985), .B(n17984), .Z(n17989) );
  NANDN U18346 ( .A(n17987), .B(n17986), .Z(n17988) );
  NAND U18347 ( .A(n17989), .B(n17988), .Z(n17996) );
  XNOR U18348 ( .A(n17995), .B(n17996), .Z(n17997) );
  XNOR U18349 ( .A(n17998), .B(n17997), .Z(n18068) );
  XNOR U18350 ( .A(n18068), .B(sreg[477]), .Z(n18070) );
  NAND U18351 ( .A(n17990), .B(sreg[476]), .Z(n17994) );
  OR U18352 ( .A(n17992), .B(n17991), .Z(n17993) );
  AND U18353 ( .A(n17994), .B(n17993), .Z(n18069) );
  XOR U18354 ( .A(n18070), .B(n18069), .Z(c[477]) );
  NANDN U18355 ( .A(n17996), .B(n17995), .Z(n18000) );
  NAND U18356 ( .A(n17998), .B(n17997), .Z(n17999) );
  NAND U18357 ( .A(n18000), .B(n17999), .Z(n18076) );
  NANDN U18358 ( .A(n18002), .B(n18001), .Z(n18006) );
  OR U18359 ( .A(n18004), .B(n18003), .Z(n18005) );
  NAND U18360 ( .A(n18006), .B(n18005), .Z(n18143) );
  NANDN U18361 ( .A(n18008), .B(n18007), .Z(n18012) );
  OR U18362 ( .A(n18010), .B(n18009), .Z(n18011) );
  NAND U18363 ( .A(n18012), .B(n18011), .Z(n18109) );
  NAND U18364 ( .A(b[0]), .B(a[238]), .Z(n18013) );
  XNOR U18365 ( .A(b[1]), .B(n18013), .Z(n18015) );
  NAND U18366 ( .A(n98), .B(a[237]), .Z(n18014) );
  AND U18367 ( .A(n18015), .B(n18014), .Z(n18085) );
  XNOR U18368 ( .A(n20154), .B(n18193), .Z(n18094) );
  OR U18369 ( .A(n18094), .B(n20057), .Z(n18018) );
  NANDN U18370 ( .A(n18016), .B(n20098), .Z(n18017) );
  AND U18371 ( .A(n18018), .B(n18017), .Z(n18086) );
  XOR U18372 ( .A(n18085), .B(n18086), .Z(n18088) );
  NAND U18373 ( .A(a[222]), .B(b[15]), .Z(n18087) );
  XOR U18374 ( .A(n18088), .B(n18087), .Z(n18106) );
  NAND U18375 ( .A(n19722), .B(n18019), .Z(n18021) );
  XNOR U18376 ( .A(b[5]), .B(n18790), .Z(n18097) );
  NANDN U18377 ( .A(n19640), .B(n18097), .Z(n18020) );
  NAND U18378 ( .A(n18021), .B(n18020), .Z(n18131) );
  XNOR U18379 ( .A(n19714), .B(n18661), .Z(n18100) );
  NANDN U18380 ( .A(n18100), .B(n19766), .Z(n18024) );
  NANDN U18381 ( .A(n18022), .B(n19767), .Z(n18023) );
  NAND U18382 ( .A(n18024), .B(n18023), .Z(n18128) );
  NAND U18383 ( .A(n19554), .B(n18025), .Z(n18027) );
  IV U18384 ( .A(a[236]), .Z(n18946) );
  XNOR U18385 ( .A(b[3]), .B(n18946), .Z(n18103) );
  NANDN U18386 ( .A(n19521), .B(n18103), .Z(n18026) );
  AND U18387 ( .A(n18027), .B(n18026), .Z(n18129) );
  XNOR U18388 ( .A(n18128), .B(n18129), .Z(n18130) );
  XOR U18389 ( .A(n18131), .B(n18130), .Z(n18107) );
  XOR U18390 ( .A(n18106), .B(n18107), .Z(n18108) );
  XNOR U18391 ( .A(n18109), .B(n18108), .Z(n18079) );
  NAND U18392 ( .A(n18029), .B(n18028), .Z(n18033) );
  NAND U18393 ( .A(n18031), .B(n18030), .Z(n18032) );
  NAND U18394 ( .A(n18033), .B(n18032), .Z(n18080) );
  XOR U18395 ( .A(n18079), .B(n18080), .Z(n18082) );
  XNOR U18396 ( .A(n20052), .B(n18322), .Z(n18112) );
  OR U18397 ( .A(n18112), .B(n20020), .Z(n18036) );
  NANDN U18398 ( .A(n18034), .B(n19960), .Z(n18035) );
  NAND U18399 ( .A(n18036), .B(n18035), .Z(n18125) );
  XNOR U18400 ( .A(n102), .B(n18037), .Z(n18116) );
  OR U18401 ( .A(n18116), .B(n20121), .Z(n18040) );
  NANDN U18402 ( .A(n18038), .B(n20122), .Z(n18039) );
  NAND U18403 ( .A(n18040), .B(n18039), .Z(n18122) );
  XNOR U18404 ( .A(n19975), .B(n18505), .Z(n18119) );
  NANDN U18405 ( .A(n18119), .B(n19883), .Z(n18043) );
  NANDN U18406 ( .A(n18041), .B(n19937), .Z(n18042) );
  AND U18407 ( .A(n18043), .B(n18042), .Z(n18123) );
  XNOR U18408 ( .A(n18122), .B(n18123), .Z(n18124) );
  XNOR U18409 ( .A(n18125), .B(n18124), .Z(n18134) );
  NANDN U18410 ( .A(n18045), .B(n18044), .Z(n18049) );
  NAND U18411 ( .A(n18047), .B(n18046), .Z(n18048) );
  NAND U18412 ( .A(n18049), .B(n18048), .Z(n18135) );
  XNOR U18413 ( .A(n18134), .B(n18135), .Z(n18136) );
  NANDN U18414 ( .A(n18051), .B(n18050), .Z(n18055) );
  NAND U18415 ( .A(n18053), .B(n18052), .Z(n18054) );
  AND U18416 ( .A(n18055), .B(n18054), .Z(n18137) );
  XNOR U18417 ( .A(n18136), .B(n18137), .Z(n18081) );
  XNOR U18418 ( .A(n18082), .B(n18081), .Z(n18140) );
  NANDN U18419 ( .A(n18057), .B(n18056), .Z(n18061) );
  NAND U18420 ( .A(n18059), .B(n18058), .Z(n18060) );
  NAND U18421 ( .A(n18061), .B(n18060), .Z(n18141) );
  XNOR U18422 ( .A(n18140), .B(n18141), .Z(n18142) );
  XOR U18423 ( .A(n18143), .B(n18142), .Z(n18073) );
  NANDN U18424 ( .A(n18063), .B(n18062), .Z(n18067) );
  NANDN U18425 ( .A(n18065), .B(n18064), .Z(n18066) );
  NAND U18426 ( .A(n18067), .B(n18066), .Z(n18074) );
  XNOR U18427 ( .A(n18073), .B(n18074), .Z(n18075) );
  XNOR U18428 ( .A(n18076), .B(n18075), .Z(n18146) );
  XNOR U18429 ( .A(n18146), .B(sreg[478]), .Z(n18148) );
  NAND U18430 ( .A(n18068), .B(sreg[477]), .Z(n18072) );
  OR U18431 ( .A(n18070), .B(n18069), .Z(n18071) );
  AND U18432 ( .A(n18072), .B(n18071), .Z(n18147) );
  XOR U18433 ( .A(n18148), .B(n18147), .Z(c[478]) );
  NANDN U18434 ( .A(n18074), .B(n18073), .Z(n18078) );
  NAND U18435 ( .A(n18076), .B(n18075), .Z(n18077) );
  NAND U18436 ( .A(n18078), .B(n18077), .Z(n18154) );
  NANDN U18437 ( .A(n18080), .B(n18079), .Z(n18084) );
  OR U18438 ( .A(n18082), .B(n18081), .Z(n18083) );
  NAND U18439 ( .A(n18084), .B(n18083), .Z(n18221) );
  NANDN U18440 ( .A(n18086), .B(n18085), .Z(n18090) );
  OR U18441 ( .A(n18088), .B(n18087), .Z(n18089) );
  NAND U18442 ( .A(n18090), .B(n18089), .Z(n18187) );
  NAND U18443 ( .A(b[0]), .B(a[239]), .Z(n18091) );
  XNOR U18444 ( .A(b[1]), .B(n18091), .Z(n18093) );
  NAND U18445 ( .A(a[238]), .B(n98), .Z(n18092) );
  AND U18446 ( .A(n18093), .B(n18092), .Z(n18163) );
  XNOR U18447 ( .A(n20154), .B(n18244), .Z(n18172) );
  OR U18448 ( .A(n18172), .B(n20057), .Z(n18096) );
  NANDN U18449 ( .A(n18094), .B(n20098), .Z(n18095) );
  AND U18450 ( .A(n18096), .B(n18095), .Z(n18164) );
  XOR U18451 ( .A(n18163), .B(n18164), .Z(n18166) );
  NAND U18452 ( .A(a[223]), .B(b[15]), .Z(n18165) );
  XOR U18453 ( .A(n18166), .B(n18165), .Z(n18184) );
  NAND U18454 ( .A(n19722), .B(n18097), .Z(n18099) );
  XNOR U18455 ( .A(b[5]), .B(n18868), .Z(n18175) );
  NANDN U18456 ( .A(n19640), .B(n18175), .Z(n18098) );
  NAND U18457 ( .A(n18099), .B(n18098), .Z(n18209) );
  XNOR U18458 ( .A(n19714), .B(n18712), .Z(n18178) );
  NANDN U18459 ( .A(n18178), .B(n19766), .Z(n18102) );
  NANDN U18460 ( .A(n18100), .B(n19767), .Z(n18101) );
  NAND U18461 ( .A(n18102), .B(n18101), .Z(n18206) );
  NAND U18462 ( .A(n19554), .B(n18103), .Z(n18105) );
  XOR U18463 ( .A(b[3]), .B(a[237]), .Z(n18181) );
  NANDN U18464 ( .A(n19521), .B(n18181), .Z(n18104) );
  AND U18465 ( .A(n18105), .B(n18104), .Z(n18207) );
  XNOR U18466 ( .A(n18206), .B(n18207), .Z(n18208) );
  XOR U18467 ( .A(n18209), .B(n18208), .Z(n18185) );
  XOR U18468 ( .A(n18184), .B(n18185), .Z(n18186) );
  XNOR U18469 ( .A(n18187), .B(n18186), .Z(n18157) );
  NAND U18470 ( .A(n18107), .B(n18106), .Z(n18111) );
  NAND U18471 ( .A(n18109), .B(n18108), .Z(n18110) );
  NAND U18472 ( .A(n18111), .B(n18110), .Z(n18158) );
  XOR U18473 ( .A(n18157), .B(n18158), .Z(n18160) );
  XNOR U18474 ( .A(n20052), .B(n18427), .Z(n18190) );
  OR U18475 ( .A(n18190), .B(n20020), .Z(n18114) );
  NANDN U18476 ( .A(n18112), .B(n19960), .Z(n18113) );
  NAND U18477 ( .A(n18114), .B(n18113), .Z(n18203) );
  XNOR U18478 ( .A(n102), .B(n18115), .Z(n18194) );
  OR U18479 ( .A(n18194), .B(n20121), .Z(n18118) );
  NANDN U18480 ( .A(n18116), .B(n20122), .Z(n18117) );
  NAND U18481 ( .A(n18118), .B(n18117), .Z(n18200) );
  XNOR U18482 ( .A(n19975), .B(n18556), .Z(n18197) );
  NANDN U18483 ( .A(n18197), .B(n19883), .Z(n18121) );
  NANDN U18484 ( .A(n18119), .B(n19937), .Z(n18120) );
  AND U18485 ( .A(n18121), .B(n18120), .Z(n18201) );
  XNOR U18486 ( .A(n18200), .B(n18201), .Z(n18202) );
  XNOR U18487 ( .A(n18203), .B(n18202), .Z(n18212) );
  NANDN U18488 ( .A(n18123), .B(n18122), .Z(n18127) );
  NAND U18489 ( .A(n18125), .B(n18124), .Z(n18126) );
  NAND U18490 ( .A(n18127), .B(n18126), .Z(n18213) );
  XNOR U18491 ( .A(n18212), .B(n18213), .Z(n18214) );
  NANDN U18492 ( .A(n18129), .B(n18128), .Z(n18133) );
  NAND U18493 ( .A(n18131), .B(n18130), .Z(n18132) );
  AND U18494 ( .A(n18133), .B(n18132), .Z(n18215) );
  XNOR U18495 ( .A(n18214), .B(n18215), .Z(n18159) );
  XNOR U18496 ( .A(n18160), .B(n18159), .Z(n18218) );
  NANDN U18497 ( .A(n18135), .B(n18134), .Z(n18139) );
  NAND U18498 ( .A(n18137), .B(n18136), .Z(n18138) );
  NAND U18499 ( .A(n18139), .B(n18138), .Z(n18219) );
  XNOR U18500 ( .A(n18218), .B(n18219), .Z(n18220) );
  XOR U18501 ( .A(n18221), .B(n18220), .Z(n18151) );
  NANDN U18502 ( .A(n18141), .B(n18140), .Z(n18145) );
  NANDN U18503 ( .A(n18143), .B(n18142), .Z(n18144) );
  NAND U18504 ( .A(n18145), .B(n18144), .Z(n18152) );
  XNOR U18505 ( .A(n18151), .B(n18152), .Z(n18153) );
  XNOR U18506 ( .A(n18154), .B(n18153), .Z(n18224) );
  XNOR U18507 ( .A(n18224), .B(sreg[479]), .Z(n18226) );
  NAND U18508 ( .A(n18146), .B(sreg[478]), .Z(n18150) );
  OR U18509 ( .A(n18148), .B(n18147), .Z(n18149) );
  AND U18510 ( .A(n18150), .B(n18149), .Z(n18225) );
  XOR U18511 ( .A(n18226), .B(n18225), .Z(c[479]) );
  NANDN U18512 ( .A(n18152), .B(n18151), .Z(n18156) );
  NAND U18513 ( .A(n18154), .B(n18153), .Z(n18155) );
  NAND U18514 ( .A(n18156), .B(n18155), .Z(n18232) );
  NANDN U18515 ( .A(n18158), .B(n18157), .Z(n18162) );
  OR U18516 ( .A(n18160), .B(n18159), .Z(n18161) );
  NAND U18517 ( .A(n18162), .B(n18161), .Z(n18299) );
  NANDN U18518 ( .A(n18164), .B(n18163), .Z(n18168) );
  OR U18519 ( .A(n18166), .B(n18165), .Z(n18167) );
  NAND U18520 ( .A(n18168), .B(n18167), .Z(n18287) );
  NAND U18521 ( .A(b[0]), .B(a[240]), .Z(n18169) );
  XNOR U18522 ( .A(b[1]), .B(n18169), .Z(n18171) );
  NAND U18523 ( .A(n98), .B(a[239]), .Z(n18170) );
  AND U18524 ( .A(n18171), .B(n18170), .Z(n18263) );
  XNOR U18525 ( .A(n20154), .B(n18322), .Z(n18272) );
  OR U18526 ( .A(n18272), .B(n20057), .Z(n18174) );
  NANDN U18527 ( .A(n18172), .B(n20098), .Z(n18173) );
  AND U18528 ( .A(n18174), .B(n18173), .Z(n18264) );
  XOR U18529 ( .A(n18263), .B(n18264), .Z(n18266) );
  NAND U18530 ( .A(a[224]), .B(b[15]), .Z(n18265) );
  XOR U18531 ( .A(n18266), .B(n18265), .Z(n18284) );
  NAND U18532 ( .A(n19722), .B(n18175), .Z(n18177) );
  XNOR U18533 ( .A(b[5]), .B(n18946), .Z(n18275) );
  NANDN U18534 ( .A(n19640), .B(n18275), .Z(n18176) );
  NAND U18535 ( .A(n18177), .B(n18176), .Z(n18260) );
  XNOR U18536 ( .A(n19714), .B(n18790), .Z(n18278) );
  NANDN U18537 ( .A(n18278), .B(n19766), .Z(n18180) );
  NANDN U18538 ( .A(n18178), .B(n19767), .Z(n18179) );
  NAND U18539 ( .A(n18180), .B(n18179), .Z(n18257) );
  NAND U18540 ( .A(n19554), .B(n18181), .Z(n18183) );
  IV U18541 ( .A(a[238]), .Z(n19128) );
  XNOR U18542 ( .A(b[3]), .B(n19128), .Z(n18281) );
  NANDN U18543 ( .A(n19521), .B(n18281), .Z(n18182) );
  AND U18544 ( .A(n18183), .B(n18182), .Z(n18258) );
  XNOR U18545 ( .A(n18257), .B(n18258), .Z(n18259) );
  XOR U18546 ( .A(n18260), .B(n18259), .Z(n18285) );
  XOR U18547 ( .A(n18284), .B(n18285), .Z(n18286) );
  XNOR U18548 ( .A(n18287), .B(n18286), .Z(n18235) );
  NAND U18549 ( .A(n18185), .B(n18184), .Z(n18189) );
  NAND U18550 ( .A(n18187), .B(n18186), .Z(n18188) );
  NAND U18551 ( .A(n18189), .B(n18188), .Z(n18236) );
  XOR U18552 ( .A(n18235), .B(n18236), .Z(n18238) );
  XNOR U18553 ( .A(n20052), .B(n18505), .Z(n18241) );
  OR U18554 ( .A(n18241), .B(n20020), .Z(n18192) );
  NANDN U18555 ( .A(n18190), .B(n19960), .Z(n18191) );
  NAND U18556 ( .A(n18192), .B(n18191), .Z(n18254) );
  XNOR U18557 ( .A(n102), .B(n18193), .Z(n18245) );
  OR U18558 ( .A(n18245), .B(n20121), .Z(n18196) );
  NANDN U18559 ( .A(n18194), .B(n20122), .Z(n18195) );
  NAND U18560 ( .A(n18196), .B(n18195), .Z(n18251) );
  XNOR U18561 ( .A(n19975), .B(n18661), .Z(n18248) );
  NANDN U18562 ( .A(n18248), .B(n19883), .Z(n18199) );
  NANDN U18563 ( .A(n18197), .B(n19937), .Z(n18198) );
  AND U18564 ( .A(n18199), .B(n18198), .Z(n18252) );
  XNOR U18565 ( .A(n18251), .B(n18252), .Z(n18253) );
  XNOR U18566 ( .A(n18254), .B(n18253), .Z(n18290) );
  NANDN U18567 ( .A(n18201), .B(n18200), .Z(n18205) );
  NAND U18568 ( .A(n18203), .B(n18202), .Z(n18204) );
  NAND U18569 ( .A(n18205), .B(n18204), .Z(n18291) );
  XNOR U18570 ( .A(n18290), .B(n18291), .Z(n18292) );
  NANDN U18571 ( .A(n18207), .B(n18206), .Z(n18211) );
  NAND U18572 ( .A(n18209), .B(n18208), .Z(n18210) );
  AND U18573 ( .A(n18211), .B(n18210), .Z(n18293) );
  XNOR U18574 ( .A(n18292), .B(n18293), .Z(n18237) );
  XNOR U18575 ( .A(n18238), .B(n18237), .Z(n18296) );
  NANDN U18576 ( .A(n18213), .B(n18212), .Z(n18217) );
  NAND U18577 ( .A(n18215), .B(n18214), .Z(n18216) );
  NAND U18578 ( .A(n18217), .B(n18216), .Z(n18297) );
  XNOR U18579 ( .A(n18296), .B(n18297), .Z(n18298) );
  XOR U18580 ( .A(n18299), .B(n18298), .Z(n18229) );
  NANDN U18581 ( .A(n18219), .B(n18218), .Z(n18223) );
  NANDN U18582 ( .A(n18221), .B(n18220), .Z(n18222) );
  NAND U18583 ( .A(n18223), .B(n18222), .Z(n18230) );
  XNOR U18584 ( .A(n18229), .B(n18230), .Z(n18231) );
  XNOR U18585 ( .A(n18232), .B(n18231), .Z(n18302) );
  XNOR U18586 ( .A(n18302), .B(sreg[480]), .Z(n18304) );
  NAND U18587 ( .A(n18224), .B(sreg[479]), .Z(n18228) );
  OR U18588 ( .A(n18226), .B(n18225), .Z(n18227) );
  AND U18589 ( .A(n18228), .B(n18227), .Z(n18303) );
  XOR U18590 ( .A(n18304), .B(n18303), .Z(c[480]) );
  NANDN U18591 ( .A(n18230), .B(n18229), .Z(n18234) );
  NAND U18592 ( .A(n18232), .B(n18231), .Z(n18233) );
  NAND U18593 ( .A(n18234), .B(n18233), .Z(n18310) );
  NANDN U18594 ( .A(n18236), .B(n18235), .Z(n18240) );
  OR U18595 ( .A(n18238), .B(n18237), .Z(n18239) );
  NAND U18596 ( .A(n18240), .B(n18239), .Z(n18377) );
  XNOR U18597 ( .A(n20052), .B(n18556), .Z(n18319) );
  OR U18598 ( .A(n18319), .B(n20020), .Z(n18243) );
  NANDN U18599 ( .A(n18241), .B(n19960), .Z(n18242) );
  NAND U18600 ( .A(n18243), .B(n18242), .Z(n18332) );
  XNOR U18601 ( .A(n102), .B(n18244), .Z(n18323) );
  OR U18602 ( .A(n18323), .B(n20121), .Z(n18247) );
  NANDN U18603 ( .A(n18245), .B(n20122), .Z(n18246) );
  NAND U18604 ( .A(n18247), .B(n18246), .Z(n18329) );
  XNOR U18605 ( .A(n19975), .B(n18712), .Z(n18326) );
  NANDN U18606 ( .A(n18326), .B(n19883), .Z(n18250) );
  NANDN U18607 ( .A(n18248), .B(n19937), .Z(n18249) );
  AND U18608 ( .A(n18250), .B(n18249), .Z(n18330) );
  XNOR U18609 ( .A(n18329), .B(n18330), .Z(n18331) );
  XNOR U18610 ( .A(n18332), .B(n18331), .Z(n18368) );
  NANDN U18611 ( .A(n18252), .B(n18251), .Z(n18256) );
  NAND U18612 ( .A(n18254), .B(n18253), .Z(n18255) );
  NAND U18613 ( .A(n18256), .B(n18255), .Z(n18369) );
  XNOR U18614 ( .A(n18368), .B(n18369), .Z(n18370) );
  NANDN U18615 ( .A(n18258), .B(n18257), .Z(n18262) );
  NAND U18616 ( .A(n18260), .B(n18259), .Z(n18261) );
  AND U18617 ( .A(n18262), .B(n18261), .Z(n18371) );
  XNOR U18618 ( .A(n18370), .B(n18371), .Z(n18315) );
  NANDN U18619 ( .A(n18264), .B(n18263), .Z(n18268) );
  OR U18620 ( .A(n18266), .B(n18265), .Z(n18267) );
  NAND U18621 ( .A(n18268), .B(n18267), .Z(n18365) );
  NAND U18622 ( .A(b[0]), .B(a[241]), .Z(n18269) );
  XNOR U18623 ( .A(b[1]), .B(n18269), .Z(n18271) );
  NAND U18624 ( .A(n98), .B(a[240]), .Z(n18270) );
  AND U18625 ( .A(n18271), .B(n18270), .Z(n18341) );
  XNOR U18626 ( .A(n20154), .B(n18427), .Z(n18350) );
  OR U18627 ( .A(n18350), .B(n20057), .Z(n18274) );
  NANDN U18628 ( .A(n18272), .B(n20098), .Z(n18273) );
  AND U18629 ( .A(n18274), .B(n18273), .Z(n18342) );
  XOR U18630 ( .A(n18341), .B(n18342), .Z(n18344) );
  NAND U18631 ( .A(a[225]), .B(b[15]), .Z(n18343) );
  XOR U18632 ( .A(n18344), .B(n18343), .Z(n18362) );
  NAND U18633 ( .A(n19722), .B(n18275), .Z(n18277) );
  XOR U18634 ( .A(b[5]), .B(a[237]), .Z(n18353) );
  NANDN U18635 ( .A(n19640), .B(n18353), .Z(n18276) );
  NAND U18636 ( .A(n18277), .B(n18276), .Z(n18338) );
  XNOR U18637 ( .A(n19714), .B(n18868), .Z(n18356) );
  NANDN U18638 ( .A(n18356), .B(n19766), .Z(n18280) );
  NANDN U18639 ( .A(n18278), .B(n19767), .Z(n18279) );
  NAND U18640 ( .A(n18280), .B(n18279), .Z(n18335) );
  NAND U18641 ( .A(n19554), .B(n18281), .Z(n18283) );
  XOR U18642 ( .A(b[3]), .B(a[239]), .Z(n18359) );
  NANDN U18643 ( .A(n19521), .B(n18359), .Z(n18282) );
  AND U18644 ( .A(n18283), .B(n18282), .Z(n18336) );
  XNOR U18645 ( .A(n18335), .B(n18336), .Z(n18337) );
  XOR U18646 ( .A(n18338), .B(n18337), .Z(n18363) );
  XOR U18647 ( .A(n18362), .B(n18363), .Z(n18364) );
  XNOR U18648 ( .A(n18365), .B(n18364), .Z(n18313) );
  NAND U18649 ( .A(n18285), .B(n18284), .Z(n18289) );
  NAND U18650 ( .A(n18287), .B(n18286), .Z(n18288) );
  NAND U18651 ( .A(n18289), .B(n18288), .Z(n18314) );
  XOR U18652 ( .A(n18313), .B(n18314), .Z(n18316) );
  XNOR U18653 ( .A(n18315), .B(n18316), .Z(n18374) );
  NANDN U18654 ( .A(n18291), .B(n18290), .Z(n18295) );
  NAND U18655 ( .A(n18293), .B(n18292), .Z(n18294) );
  NAND U18656 ( .A(n18295), .B(n18294), .Z(n18375) );
  XNOR U18657 ( .A(n18374), .B(n18375), .Z(n18376) );
  XOR U18658 ( .A(n18377), .B(n18376), .Z(n18307) );
  NANDN U18659 ( .A(n18297), .B(n18296), .Z(n18301) );
  NANDN U18660 ( .A(n18299), .B(n18298), .Z(n18300) );
  NAND U18661 ( .A(n18301), .B(n18300), .Z(n18308) );
  XNOR U18662 ( .A(n18307), .B(n18308), .Z(n18309) );
  XNOR U18663 ( .A(n18310), .B(n18309), .Z(n18380) );
  XNOR U18664 ( .A(n18380), .B(sreg[481]), .Z(n18382) );
  NAND U18665 ( .A(n18302), .B(sreg[480]), .Z(n18306) );
  OR U18666 ( .A(n18304), .B(n18303), .Z(n18305) );
  AND U18667 ( .A(n18306), .B(n18305), .Z(n18381) );
  XOR U18668 ( .A(n18382), .B(n18381), .Z(c[481]) );
  NANDN U18669 ( .A(n18308), .B(n18307), .Z(n18312) );
  NAND U18670 ( .A(n18310), .B(n18309), .Z(n18311) );
  NAND U18671 ( .A(n18312), .B(n18311), .Z(n18388) );
  NANDN U18672 ( .A(n18314), .B(n18313), .Z(n18318) );
  OR U18673 ( .A(n18316), .B(n18315), .Z(n18317) );
  NAND U18674 ( .A(n18318), .B(n18317), .Z(n18455) );
  XNOR U18675 ( .A(n20052), .B(n18661), .Z(n18424) );
  OR U18676 ( .A(n18424), .B(n20020), .Z(n18321) );
  NANDN U18677 ( .A(n18319), .B(n19960), .Z(n18320) );
  NAND U18678 ( .A(n18321), .B(n18320), .Z(n18437) );
  XNOR U18679 ( .A(n102), .B(n18322), .Z(n18428) );
  OR U18680 ( .A(n18428), .B(n20121), .Z(n18325) );
  NANDN U18681 ( .A(n18323), .B(n20122), .Z(n18324) );
  NAND U18682 ( .A(n18325), .B(n18324), .Z(n18434) );
  XNOR U18683 ( .A(n19975), .B(n18790), .Z(n18431) );
  NANDN U18684 ( .A(n18431), .B(n19883), .Z(n18328) );
  NANDN U18685 ( .A(n18326), .B(n19937), .Z(n18327) );
  AND U18686 ( .A(n18328), .B(n18327), .Z(n18435) );
  XNOR U18687 ( .A(n18434), .B(n18435), .Z(n18436) );
  XNOR U18688 ( .A(n18437), .B(n18436), .Z(n18446) );
  NANDN U18689 ( .A(n18330), .B(n18329), .Z(n18334) );
  NAND U18690 ( .A(n18332), .B(n18331), .Z(n18333) );
  NAND U18691 ( .A(n18334), .B(n18333), .Z(n18447) );
  XNOR U18692 ( .A(n18446), .B(n18447), .Z(n18448) );
  NANDN U18693 ( .A(n18336), .B(n18335), .Z(n18340) );
  NAND U18694 ( .A(n18338), .B(n18337), .Z(n18339) );
  AND U18695 ( .A(n18340), .B(n18339), .Z(n18449) );
  XNOR U18696 ( .A(n18448), .B(n18449), .Z(n18393) );
  NANDN U18697 ( .A(n18342), .B(n18341), .Z(n18346) );
  OR U18698 ( .A(n18344), .B(n18343), .Z(n18345) );
  NAND U18699 ( .A(n18346), .B(n18345), .Z(n18421) );
  NAND U18700 ( .A(b[0]), .B(a[242]), .Z(n18347) );
  XNOR U18701 ( .A(b[1]), .B(n18347), .Z(n18349) );
  NAND U18702 ( .A(n98), .B(a[241]), .Z(n18348) );
  AND U18703 ( .A(n18349), .B(n18348), .Z(n18397) );
  XNOR U18704 ( .A(n20154), .B(n18505), .Z(n18406) );
  OR U18705 ( .A(n18406), .B(n20057), .Z(n18352) );
  NANDN U18706 ( .A(n18350), .B(n20098), .Z(n18351) );
  AND U18707 ( .A(n18352), .B(n18351), .Z(n18398) );
  XOR U18708 ( .A(n18397), .B(n18398), .Z(n18400) );
  NAND U18709 ( .A(a[226]), .B(b[15]), .Z(n18399) );
  XOR U18710 ( .A(n18400), .B(n18399), .Z(n18418) );
  NAND U18711 ( .A(n19722), .B(n18353), .Z(n18355) );
  XNOR U18712 ( .A(b[5]), .B(n19128), .Z(n18409) );
  NANDN U18713 ( .A(n19640), .B(n18409), .Z(n18354) );
  NAND U18714 ( .A(n18355), .B(n18354), .Z(n18443) );
  XNOR U18715 ( .A(n19714), .B(n18946), .Z(n18412) );
  NANDN U18716 ( .A(n18412), .B(n19766), .Z(n18358) );
  NANDN U18717 ( .A(n18356), .B(n19767), .Z(n18357) );
  NAND U18718 ( .A(n18358), .B(n18357), .Z(n18440) );
  NAND U18719 ( .A(n19554), .B(n18359), .Z(n18361) );
  XOR U18720 ( .A(b[3]), .B(a[240]), .Z(n18415) );
  NANDN U18721 ( .A(n19521), .B(n18415), .Z(n18360) );
  AND U18722 ( .A(n18361), .B(n18360), .Z(n18441) );
  XNOR U18723 ( .A(n18440), .B(n18441), .Z(n18442) );
  XOR U18724 ( .A(n18443), .B(n18442), .Z(n18419) );
  XOR U18725 ( .A(n18418), .B(n18419), .Z(n18420) );
  XNOR U18726 ( .A(n18421), .B(n18420), .Z(n18391) );
  NAND U18727 ( .A(n18363), .B(n18362), .Z(n18367) );
  NAND U18728 ( .A(n18365), .B(n18364), .Z(n18366) );
  NAND U18729 ( .A(n18367), .B(n18366), .Z(n18392) );
  XOR U18730 ( .A(n18391), .B(n18392), .Z(n18394) );
  XNOR U18731 ( .A(n18393), .B(n18394), .Z(n18452) );
  NANDN U18732 ( .A(n18369), .B(n18368), .Z(n18373) );
  NAND U18733 ( .A(n18371), .B(n18370), .Z(n18372) );
  NAND U18734 ( .A(n18373), .B(n18372), .Z(n18453) );
  XNOR U18735 ( .A(n18452), .B(n18453), .Z(n18454) );
  XOR U18736 ( .A(n18455), .B(n18454), .Z(n18385) );
  NANDN U18737 ( .A(n18375), .B(n18374), .Z(n18379) );
  NANDN U18738 ( .A(n18377), .B(n18376), .Z(n18378) );
  NAND U18739 ( .A(n18379), .B(n18378), .Z(n18386) );
  XNOR U18740 ( .A(n18385), .B(n18386), .Z(n18387) );
  XNOR U18741 ( .A(n18388), .B(n18387), .Z(n18458) );
  XNOR U18742 ( .A(n18458), .B(sreg[482]), .Z(n18460) );
  NAND U18743 ( .A(n18380), .B(sreg[481]), .Z(n18384) );
  OR U18744 ( .A(n18382), .B(n18381), .Z(n18383) );
  AND U18745 ( .A(n18384), .B(n18383), .Z(n18459) );
  XOR U18746 ( .A(n18460), .B(n18459), .Z(c[482]) );
  NANDN U18747 ( .A(n18386), .B(n18385), .Z(n18390) );
  NAND U18748 ( .A(n18388), .B(n18387), .Z(n18389) );
  NAND U18749 ( .A(n18390), .B(n18389), .Z(n18466) );
  NANDN U18750 ( .A(n18392), .B(n18391), .Z(n18396) );
  OR U18751 ( .A(n18394), .B(n18393), .Z(n18395) );
  NAND U18752 ( .A(n18396), .B(n18395), .Z(n18533) );
  NANDN U18753 ( .A(n18398), .B(n18397), .Z(n18402) );
  OR U18754 ( .A(n18400), .B(n18399), .Z(n18401) );
  NAND U18755 ( .A(n18402), .B(n18401), .Z(n18499) );
  NAND U18756 ( .A(b[0]), .B(a[243]), .Z(n18403) );
  XNOR U18757 ( .A(b[1]), .B(n18403), .Z(n18405) );
  NAND U18758 ( .A(a[242]), .B(n98), .Z(n18404) );
  AND U18759 ( .A(n18405), .B(n18404), .Z(n18475) );
  XNOR U18760 ( .A(n20154), .B(n18556), .Z(n18481) );
  OR U18761 ( .A(n18481), .B(n20057), .Z(n18408) );
  NANDN U18762 ( .A(n18406), .B(n20098), .Z(n18407) );
  AND U18763 ( .A(n18408), .B(n18407), .Z(n18476) );
  XOR U18764 ( .A(n18475), .B(n18476), .Z(n18478) );
  NAND U18765 ( .A(a[227]), .B(b[15]), .Z(n18477) );
  XOR U18766 ( .A(n18478), .B(n18477), .Z(n18496) );
  NAND U18767 ( .A(n19722), .B(n18409), .Z(n18411) );
  XOR U18768 ( .A(b[5]), .B(a[239]), .Z(n18487) );
  NANDN U18769 ( .A(n19640), .B(n18487), .Z(n18410) );
  NAND U18770 ( .A(n18411), .B(n18410), .Z(n18521) );
  XOR U18771 ( .A(n19714), .B(a[237]), .Z(n18490) );
  NANDN U18772 ( .A(n18490), .B(n19766), .Z(n18414) );
  NANDN U18773 ( .A(n18412), .B(n19767), .Z(n18413) );
  NAND U18774 ( .A(n18414), .B(n18413), .Z(n18518) );
  NAND U18775 ( .A(n19554), .B(n18415), .Z(n18417) );
  XOR U18776 ( .A(b[3]), .B(a[241]), .Z(n18493) );
  NANDN U18777 ( .A(n19521), .B(n18493), .Z(n18416) );
  AND U18778 ( .A(n18417), .B(n18416), .Z(n18519) );
  XNOR U18779 ( .A(n18518), .B(n18519), .Z(n18520) );
  XOR U18780 ( .A(n18521), .B(n18520), .Z(n18497) );
  XOR U18781 ( .A(n18496), .B(n18497), .Z(n18498) );
  XNOR U18782 ( .A(n18499), .B(n18498), .Z(n18469) );
  NAND U18783 ( .A(n18419), .B(n18418), .Z(n18423) );
  NAND U18784 ( .A(n18421), .B(n18420), .Z(n18422) );
  NAND U18785 ( .A(n18423), .B(n18422), .Z(n18470) );
  XOR U18786 ( .A(n18469), .B(n18470), .Z(n18472) );
  XNOR U18787 ( .A(n20052), .B(n18712), .Z(n18502) );
  OR U18788 ( .A(n18502), .B(n20020), .Z(n18426) );
  NANDN U18789 ( .A(n18424), .B(n19960), .Z(n18425) );
  NAND U18790 ( .A(n18426), .B(n18425), .Z(n18515) );
  XNOR U18791 ( .A(n102), .B(n18427), .Z(n18506) );
  OR U18792 ( .A(n18506), .B(n20121), .Z(n18430) );
  NANDN U18793 ( .A(n18428), .B(n20122), .Z(n18429) );
  NAND U18794 ( .A(n18430), .B(n18429), .Z(n18512) );
  XNOR U18795 ( .A(n19975), .B(n18868), .Z(n18509) );
  NANDN U18796 ( .A(n18509), .B(n19883), .Z(n18433) );
  NANDN U18797 ( .A(n18431), .B(n19937), .Z(n18432) );
  AND U18798 ( .A(n18433), .B(n18432), .Z(n18513) );
  XNOR U18799 ( .A(n18512), .B(n18513), .Z(n18514) );
  XNOR U18800 ( .A(n18515), .B(n18514), .Z(n18524) );
  NANDN U18801 ( .A(n18435), .B(n18434), .Z(n18439) );
  NAND U18802 ( .A(n18437), .B(n18436), .Z(n18438) );
  NAND U18803 ( .A(n18439), .B(n18438), .Z(n18525) );
  XNOR U18804 ( .A(n18524), .B(n18525), .Z(n18526) );
  NANDN U18805 ( .A(n18441), .B(n18440), .Z(n18445) );
  NAND U18806 ( .A(n18443), .B(n18442), .Z(n18444) );
  AND U18807 ( .A(n18445), .B(n18444), .Z(n18527) );
  XNOR U18808 ( .A(n18526), .B(n18527), .Z(n18471) );
  XNOR U18809 ( .A(n18472), .B(n18471), .Z(n18530) );
  NANDN U18810 ( .A(n18447), .B(n18446), .Z(n18451) );
  NAND U18811 ( .A(n18449), .B(n18448), .Z(n18450) );
  NAND U18812 ( .A(n18451), .B(n18450), .Z(n18531) );
  XNOR U18813 ( .A(n18530), .B(n18531), .Z(n18532) );
  XOR U18814 ( .A(n18533), .B(n18532), .Z(n18463) );
  NANDN U18815 ( .A(n18453), .B(n18452), .Z(n18457) );
  NANDN U18816 ( .A(n18455), .B(n18454), .Z(n18456) );
  NAND U18817 ( .A(n18457), .B(n18456), .Z(n18464) );
  XNOR U18818 ( .A(n18463), .B(n18464), .Z(n18465) );
  XNOR U18819 ( .A(n18466), .B(n18465), .Z(n18536) );
  XNOR U18820 ( .A(n18536), .B(sreg[483]), .Z(n18538) );
  NAND U18821 ( .A(n18458), .B(sreg[482]), .Z(n18462) );
  OR U18822 ( .A(n18460), .B(n18459), .Z(n18461) );
  AND U18823 ( .A(n18462), .B(n18461), .Z(n18537) );
  XOR U18824 ( .A(n18538), .B(n18537), .Z(c[483]) );
  NANDN U18825 ( .A(n18464), .B(n18463), .Z(n18468) );
  NAND U18826 ( .A(n18466), .B(n18465), .Z(n18467) );
  NAND U18827 ( .A(n18468), .B(n18467), .Z(n18544) );
  NANDN U18828 ( .A(n18470), .B(n18469), .Z(n18474) );
  OR U18829 ( .A(n18472), .B(n18471), .Z(n18473) );
  NAND U18830 ( .A(n18474), .B(n18473), .Z(n18611) );
  NANDN U18831 ( .A(n18476), .B(n18475), .Z(n18480) );
  OR U18832 ( .A(n18478), .B(n18477), .Z(n18479) );
  NAND U18833 ( .A(n18480), .B(n18479), .Z(n18599) );
  XNOR U18834 ( .A(n20154), .B(n18661), .Z(n18584) );
  OR U18835 ( .A(n18584), .B(n20057), .Z(n18483) );
  NANDN U18836 ( .A(n18481), .B(n20098), .Z(n18482) );
  AND U18837 ( .A(n18483), .B(n18482), .Z(n18576) );
  NAND U18838 ( .A(b[0]), .B(a[244]), .Z(n18484) );
  XNOR U18839 ( .A(b[1]), .B(n18484), .Z(n18486) );
  NAND U18840 ( .A(n98), .B(a[243]), .Z(n18485) );
  AND U18841 ( .A(n18486), .B(n18485), .Z(n18575) );
  XOR U18842 ( .A(n18576), .B(n18575), .Z(n18578) );
  NAND U18843 ( .A(a[228]), .B(b[15]), .Z(n18577) );
  XOR U18844 ( .A(n18578), .B(n18577), .Z(n18596) );
  NAND U18845 ( .A(n19722), .B(n18487), .Z(n18489) );
  XOR U18846 ( .A(b[5]), .B(a[240]), .Z(n18587) );
  NANDN U18847 ( .A(n19640), .B(n18587), .Z(n18488) );
  NAND U18848 ( .A(n18489), .B(n18488), .Z(n18572) );
  XNOR U18849 ( .A(n19714), .B(n19128), .Z(n18590) );
  NANDN U18850 ( .A(n18590), .B(n19766), .Z(n18492) );
  NANDN U18851 ( .A(n18490), .B(n19767), .Z(n18491) );
  NAND U18852 ( .A(n18492), .B(n18491), .Z(n18569) );
  NAND U18853 ( .A(n19554), .B(n18493), .Z(n18495) );
  IV U18854 ( .A(a[242]), .Z(n19433) );
  XNOR U18855 ( .A(b[3]), .B(n19433), .Z(n18593) );
  NANDN U18856 ( .A(n19521), .B(n18593), .Z(n18494) );
  AND U18857 ( .A(n18495), .B(n18494), .Z(n18570) );
  XNOR U18858 ( .A(n18569), .B(n18570), .Z(n18571) );
  XOR U18859 ( .A(n18572), .B(n18571), .Z(n18597) );
  XOR U18860 ( .A(n18596), .B(n18597), .Z(n18598) );
  XNOR U18861 ( .A(n18599), .B(n18598), .Z(n18547) );
  NAND U18862 ( .A(n18497), .B(n18496), .Z(n18501) );
  NAND U18863 ( .A(n18499), .B(n18498), .Z(n18500) );
  NAND U18864 ( .A(n18501), .B(n18500), .Z(n18548) );
  XOR U18865 ( .A(n18547), .B(n18548), .Z(n18550) );
  XNOR U18866 ( .A(n20052), .B(n18790), .Z(n18553) );
  OR U18867 ( .A(n18553), .B(n20020), .Z(n18504) );
  NANDN U18868 ( .A(n18502), .B(n19960), .Z(n18503) );
  NAND U18869 ( .A(n18504), .B(n18503), .Z(n18566) );
  XNOR U18870 ( .A(n102), .B(n18505), .Z(n18557) );
  OR U18871 ( .A(n18557), .B(n20121), .Z(n18508) );
  NANDN U18872 ( .A(n18506), .B(n20122), .Z(n18507) );
  NAND U18873 ( .A(n18508), .B(n18507), .Z(n18563) );
  XNOR U18874 ( .A(n19975), .B(n18946), .Z(n18560) );
  NANDN U18875 ( .A(n18560), .B(n19883), .Z(n18511) );
  NANDN U18876 ( .A(n18509), .B(n19937), .Z(n18510) );
  AND U18877 ( .A(n18511), .B(n18510), .Z(n18564) );
  XNOR U18878 ( .A(n18563), .B(n18564), .Z(n18565) );
  XNOR U18879 ( .A(n18566), .B(n18565), .Z(n18602) );
  NANDN U18880 ( .A(n18513), .B(n18512), .Z(n18517) );
  NAND U18881 ( .A(n18515), .B(n18514), .Z(n18516) );
  NAND U18882 ( .A(n18517), .B(n18516), .Z(n18603) );
  XNOR U18883 ( .A(n18602), .B(n18603), .Z(n18604) );
  NANDN U18884 ( .A(n18519), .B(n18518), .Z(n18523) );
  NAND U18885 ( .A(n18521), .B(n18520), .Z(n18522) );
  AND U18886 ( .A(n18523), .B(n18522), .Z(n18605) );
  XNOR U18887 ( .A(n18604), .B(n18605), .Z(n18549) );
  XNOR U18888 ( .A(n18550), .B(n18549), .Z(n18608) );
  NANDN U18889 ( .A(n18525), .B(n18524), .Z(n18529) );
  NAND U18890 ( .A(n18527), .B(n18526), .Z(n18528) );
  NAND U18891 ( .A(n18529), .B(n18528), .Z(n18609) );
  XNOR U18892 ( .A(n18608), .B(n18609), .Z(n18610) );
  XOR U18893 ( .A(n18611), .B(n18610), .Z(n18541) );
  NANDN U18894 ( .A(n18531), .B(n18530), .Z(n18535) );
  NANDN U18895 ( .A(n18533), .B(n18532), .Z(n18534) );
  NAND U18896 ( .A(n18535), .B(n18534), .Z(n18542) );
  XNOR U18897 ( .A(n18541), .B(n18542), .Z(n18543) );
  XNOR U18898 ( .A(n18544), .B(n18543), .Z(n18614) );
  XNOR U18899 ( .A(n18614), .B(sreg[484]), .Z(n18616) );
  NAND U18900 ( .A(n18536), .B(sreg[483]), .Z(n18540) );
  OR U18901 ( .A(n18538), .B(n18537), .Z(n18539) );
  AND U18902 ( .A(n18540), .B(n18539), .Z(n18615) );
  XOR U18903 ( .A(n18616), .B(n18615), .Z(c[484]) );
  NANDN U18904 ( .A(n18542), .B(n18541), .Z(n18546) );
  NAND U18905 ( .A(n18544), .B(n18543), .Z(n18545) );
  NAND U18906 ( .A(n18546), .B(n18545), .Z(n18622) );
  NANDN U18907 ( .A(n18548), .B(n18547), .Z(n18552) );
  OR U18908 ( .A(n18550), .B(n18549), .Z(n18551) );
  NAND U18909 ( .A(n18552), .B(n18551), .Z(n18689) );
  XNOR U18910 ( .A(n20052), .B(n18868), .Z(n18658) );
  OR U18911 ( .A(n18658), .B(n20020), .Z(n18555) );
  NANDN U18912 ( .A(n18553), .B(n19960), .Z(n18554) );
  NAND U18913 ( .A(n18555), .B(n18554), .Z(n18671) );
  XNOR U18914 ( .A(n102), .B(n18556), .Z(n18662) );
  OR U18915 ( .A(n18662), .B(n20121), .Z(n18559) );
  NANDN U18916 ( .A(n18557), .B(n20122), .Z(n18558) );
  NAND U18917 ( .A(n18559), .B(n18558), .Z(n18668) );
  XOR U18918 ( .A(n19975), .B(a[237]), .Z(n18665) );
  NANDN U18919 ( .A(n18665), .B(n19883), .Z(n18562) );
  NANDN U18920 ( .A(n18560), .B(n19937), .Z(n18561) );
  AND U18921 ( .A(n18562), .B(n18561), .Z(n18669) );
  XNOR U18922 ( .A(n18668), .B(n18669), .Z(n18670) );
  XNOR U18923 ( .A(n18671), .B(n18670), .Z(n18680) );
  NANDN U18924 ( .A(n18564), .B(n18563), .Z(n18568) );
  NAND U18925 ( .A(n18566), .B(n18565), .Z(n18567) );
  NAND U18926 ( .A(n18568), .B(n18567), .Z(n18681) );
  XNOR U18927 ( .A(n18680), .B(n18681), .Z(n18682) );
  NANDN U18928 ( .A(n18570), .B(n18569), .Z(n18574) );
  NAND U18929 ( .A(n18572), .B(n18571), .Z(n18573) );
  AND U18930 ( .A(n18574), .B(n18573), .Z(n18683) );
  XNOR U18931 ( .A(n18682), .B(n18683), .Z(n18627) );
  NANDN U18932 ( .A(n18576), .B(n18575), .Z(n18580) );
  OR U18933 ( .A(n18578), .B(n18577), .Z(n18579) );
  NAND U18934 ( .A(n18580), .B(n18579), .Z(n18655) );
  NAND U18935 ( .A(b[0]), .B(a[245]), .Z(n18581) );
  XNOR U18936 ( .A(b[1]), .B(n18581), .Z(n18583) );
  NAND U18937 ( .A(a[244]), .B(n98), .Z(n18582) );
  AND U18938 ( .A(n18583), .B(n18582), .Z(n18631) );
  XNOR U18939 ( .A(n20154), .B(n18712), .Z(n18637) );
  OR U18940 ( .A(n18637), .B(n20057), .Z(n18586) );
  NANDN U18941 ( .A(n18584), .B(n20098), .Z(n18585) );
  AND U18942 ( .A(n18586), .B(n18585), .Z(n18632) );
  XOR U18943 ( .A(n18631), .B(n18632), .Z(n18634) );
  NAND U18944 ( .A(a[229]), .B(b[15]), .Z(n18633) );
  XOR U18945 ( .A(n18634), .B(n18633), .Z(n18652) );
  NAND U18946 ( .A(n19722), .B(n18587), .Z(n18589) );
  XOR U18947 ( .A(b[5]), .B(a[241]), .Z(n18643) );
  NANDN U18948 ( .A(n19640), .B(n18643), .Z(n18588) );
  NAND U18949 ( .A(n18589), .B(n18588), .Z(n18677) );
  XOR U18950 ( .A(n19714), .B(a[239]), .Z(n18646) );
  NANDN U18951 ( .A(n18646), .B(n19766), .Z(n18592) );
  NANDN U18952 ( .A(n18590), .B(n19767), .Z(n18591) );
  NAND U18953 ( .A(n18592), .B(n18591), .Z(n18674) );
  NAND U18954 ( .A(n19554), .B(n18593), .Z(n18595) );
  XOR U18955 ( .A(b[3]), .B(a[243]), .Z(n18649) );
  NANDN U18956 ( .A(n19521), .B(n18649), .Z(n18594) );
  AND U18957 ( .A(n18595), .B(n18594), .Z(n18675) );
  XNOR U18958 ( .A(n18674), .B(n18675), .Z(n18676) );
  XOR U18959 ( .A(n18677), .B(n18676), .Z(n18653) );
  XOR U18960 ( .A(n18652), .B(n18653), .Z(n18654) );
  XNOR U18961 ( .A(n18655), .B(n18654), .Z(n18625) );
  NAND U18962 ( .A(n18597), .B(n18596), .Z(n18601) );
  NAND U18963 ( .A(n18599), .B(n18598), .Z(n18600) );
  NAND U18964 ( .A(n18601), .B(n18600), .Z(n18626) );
  XOR U18965 ( .A(n18625), .B(n18626), .Z(n18628) );
  XNOR U18966 ( .A(n18627), .B(n18628), .Z(n18686) );
  NANDN U18967 ( .A(n18603), .B(n18602), .Z(n18607) );
  NAND U18968 ( .A(n18605), .B(n18604), .Z(n18606) );
  NAND U18969 ( .A(n18607), .B(n18606), .Z(n18687) );
  XNOR U18970 ( .A(n18686), .B(n18687), .Z(n18688) );
  XOR U18971 ( .A(n18689), .B(n18688), .Z(n18619) );
  NANDN U18972 ( .A(n18609), .B(n18608), .Z(n18613) );
  NANDN U18973 ( .A(n18611), .B(n18610), .Z(n18612) );
  NAND U18974 ( .A(n18613), .B(n18612), .Z(n18620) );
  XNOR U18975 ( .A(n18619), .B(n18620), .Z(n18621) );
  XNOR U18976 ( .A(n18622), .B(n18621), .Z(n18692) );
  XNOR U18977 ( .A(n18692), .B(sreg[485]), .Z(n18694) );
  NAND U18978 ( .A(n18614), .B(sreg[484]), .Z(n18618) );
  OR U18979 ( .A(n18616), .B(n18615), .Z(n18617) );
  AND U18980 ( .A(n18618), .B(n18617), .Z(n18693) );
  XOR U18981 ( .A(n18694), .B(n18693), .Z(c[485]) );
  NANDN U18982 ( .A(n18620), .B(n18619), .Z(n18624) );
  NAND U18983 ( .A(n18622), .B(n18621), .Z(n18623) );
  NAND U18984 ( .A(n18624), .B(n18623), .Z(n18700) );
  NANDN U18985 ( .A(n18626), .B(n18625), .Z(n18630) );
  OR U18986 ( .A(n18628), .B(n18627), .Z(n18629) );
  NAND U18987 ( .A(n18630), .B(n18629), .Z(n18767) );
  NANDN U18988 ( .A(n18632), .B(n18631), .Z(n18636) );
  OR U18989 ( .A(n18634), .B(n18633), .Z(n18635) );
  NAND U18990 ( .A(n18636), .B(n18635), .Z(n18755) );
  XNOR U18991 ( .A(n20154), .B(n18790), .Z(n18740) );
  OR U18992 ( .A(n18740), .B(n20057), .Z(n18639) );
  NANDN U18993 ( .A(n18637), .B(n20098), .Z(n18638) );
  AND U18994 ( .A(n18639), .B(n18638), .Z(n18732) );
  NAND U18995 ( .A(b[0]), .B(a[246]), .Z(n18640) );
  XNOR U18996 ( .A(b[1]), .B(n18640), .Z(n18642) );
  NAND U18997 ( .A(a[245]), .B(n98), .Z(n18641) );
  AND U18998 ( .A(n18642), .B(n18641), .Z(n18731) );
  XOR U18999 ( .A(n18732), .B(n18731), .Z(n18734) );
  NAND U19000 ( .A(a[230]), .B(b[15]), .Z(n18733) );
  XOR U19001 ( .A(n18734), .B(n18733), .Z(n18752) );
  NAND U19002 ( .A(n19722), .B(n18643), .Z(n18645) );
  XNOR U19003 ( .A(b[5]), .B(n19433), .Z(n18743) );
  NANDN U19004 ( .A(n19640), .B(n18743), .Z(n18644) );
  NAND U19005 ( .A(n18645), .B(n18644), .Z(n18728) );
  XOR U19006 ( .A(n19714), .B(a[240]), .Z(n18746) );
  NANDN U19007 ( .A(n18746), .B(n19766), .Z(n18648) );
  NANDN U19008 ( .A(n18646), .B(n19767), .Z(n18647) );
  NAND U19009 ( .A(n18648), .B(n18647), .Z(n18725) );
  NAND U19010 ( .A(n19554), .B(n18649), .Z(n18651) );
  XNOR U19011 ( .A(a[244]), .B(n100), .Z(n18749) );
  NANDN U19012 ( .A(n19521), .B(n18749), .Z(n18650) );
  AND U19013 ( .A(n18651), .B(n18650), .Z(n18726) );
  XNOR U19014 ( .A(n18725), .B(n18726), .Z(n18727) );
  XOR U19015 ( .A(n18728), .B(n18727), .Z(n18753) );
  XOR U19016 ( .A(n18752), .B(n18753), .Z(n18754) );
  XNOR U19017 ( .A(n18755), .B(n18754), .Z(n18703) );
  NAND U19018 ( .A(n18653), .B(n18652), .Z(n18657) );
  NAND U19019 ( .A(n18655), .B(n18654), .Z(n18656) );
  NAND U19020 ( .A(n18657), .B(n18656), .Z(n18704) );
  XOR U19021 ( .A(n18703), .B(n18704), .Z(n18706) );
  XNOR U19022 ( .A(n20052), .B(n18946), .Z(n18709) );
  OR U19023 ( .A(n18709), .B(n20020), .Z(n18660) );
  NANDN U19024 ( .A(n18658), .B(n19960), .Z(n18659) );
  NAND U19025 ( .A(n18660), .B(n18659), .Z(n18722) );
  XNOR U19026 ( .A(n102), .B(n18661), .Z(n18713) );
  OR U19027 ( .A(n18713), .B(n20121), .Z(n18664) );
  NANDN U19028 ( .A(n18662), .B(n20122), .Z(n18663) );
  NAND U19029 ( .A(n18664), .B(n18663), .Z(n18719) );
  XNOR U19030 ( .A(n19975), .B(n19128), .Z(n18716) );
  NANDN U19031 ( .A(n18716), .B(n19883), .Z(n18667) );
  NANDN U19032 ( .A(n18665), .B(n19937), .Z(n18666) );
  AND U19033 ( .A(n18667), .B(n18666), .Z(n18720) );
  XNOR U19034 ( .A(n18719), .B(n18720), .Z(n18721) );
  XNOR U19035 ( .A(n18722), .B(n18721), .Z(n18758) );
  NANDN U19036 ( .A(n18669), .B(n18668), .Z(n18673) );
  NAND U19037 ( .A(n18671), .B(n18670), .Z(n18672) );
  NAND U19038 ( .A(n18673), .B(n18672), .Z(n18759) );
  XNOR U19039 ( .A(n18758), .B(n18759), .Z(n18760) );
  NANDN U19040 ( .A(n18675), .B(n18674), .Z(n18679) );
  NAND U19041 ( .A(n18677), .B(n18676), .Z(n18678) );
  AND U19042 ( .A(n18679), .B(n18678), .Z(n18761) );
  XNOR U19043 ( .A(n18760), .B(n18761), .Z(n18705) );
  XNOR U19044 ( .A(n18706), .B(n18705), .Z(n18764) );
  NANDN U19045 ( .A(n18681), .B(n18680), .Z(n18685) );
  NAND U19046 ( .A(n18683), .B(n18682), .Z(n18684) );
  NAND U19047 ( .A(n18685), .B(n18684), .Z(n18765) );
  XNOR U19048 ( .A(n18764), .B(n18765), .Z(n18766) );
  XOR U19049 ( .A(n18767), .B(n18766), .Z(n18697) );
  NANDN U19050 ( .A(n18687), .B(n18686), .Z(n18691) );
  NANDN U19051 ( .A(n18689), .B(n18688), .Z(n18690) );
  NAND U19052 ( .A(n18691), .B(n18690), .Z(n18698) );
  XNOR U19053 ( .A(n18697), .B(n18698), .Z(n18699) );
  XNOR U19054 ( .A(n18700), .B(n18699), .Z(n18770) );
  XNOR U19055 ( .A(n18770), .B(sreg[486]), .Z(n18772) );
  NAND U19056 ( .A(n18692), .B(sreg[485]), .Z(n18696) );
  OR U19057 ( .A(n18694), .B(n18693), .Z(n18695) );
  AND U19058 ( .A(n18696), .B(n18695), .Z(n18771) );
  XOR U19059 ( .A(n18772), .B(n18771), .Z(c[486]) );
  NANDN U19060 ( .A(n18698), .B(n18697), .Z(n18702) );
  NAND U19061 ( .A(n18700), .B(n18699), .Z(n18701) );
  NAND U19062 ( .A(n18702), .B(n18701), .Z(n18778) );
  NANDN U19063 ( .A(n18704), .B(n18703), .Z(n18708) );
  OR U19064 ( .A(n18706), .B(n18705), .Z(n18707) );
  NAND U19065 ( .A(n18708), .B(n18707), .Z(n18845) );
  XOR U19066 ( .A(n20052), .B(a[237]), .Z(n18787) );
  OR U19067 ( .A(n18787), .B(n20020), .Z(n18711) );
  NANDN U19068 ( .A(n18709), .B(n19960), .Z(n18710) );
  NAND U19069 ( .A(n18711), .B(n18710), .Z(n18800) );
  XNOR U19070 ( .A(n102), .B(n18712), .Z(n18791) );
  OR U19071 ( .A(n18791), .B(n20121), .Z(n18715) );
  NANDN U19072 ( .A(n18713), .B(n20122), .Z(n18714) );
  NAND U19073 ( .A(n18715), .B(n18714), .Z(n18797) );
  XOR U19074 ( .A(n19975), .B(a[239]), .Z(n18794) );
  NANDN U19075 ( .A(n18794), .B(n19883), .Z(n18718) );
  NANDN U19076 ( .A(n18716), .B(n19937), .Z(n18717) );
  AND U19077 ( .A(n18718), .B(n18717), .Z(n18798) );
  XNOR U19078 ( .A(n18797), .B(n18798), .Z(n18799) );
  XNOR U19079 ( .A(n18800), .B(n18799), .Z(n18836) );
  NANDN U19080 ( .A(n18720), .B(n18719), .Z(n18724) );
  NAND U19081 ( .A(n18722), .B(n18721), .Z(n18723) );
  NAND U19082 ( .A(n18724), .B(n18723), .Z(n18837) );
  XNOR U19083 ( .A(n18836), .B(n18837), .Z(n18838) );
  NANDN U19084 ( .A(n18726), .B(n18725), .Z(n18730) );
  NAND U19085 ( .A(n18728), .B(n18727), .Z(n18729) );
  AND U19086 ( .A(n18730), .B(n18729), .Z(n18839) );
  XNOR U19087 ( .A(n18838), .B(n18839), .Z(n18783) );
  NANDN U19088 ( .A(n18732), .B(n18731), .Z(n18736) );
  OR U19089 ( .A(n18734), .B(n18733), .Z(n18735) );
  NAND U19090 ( .A(n18736), .B(n18735), .Z(n18833) );
  NAND U19091 ( .A(b[0]), .B(a[247]), .Z(n18737) );
  XNOR U19092 ( .A(b[1]), .B(n18737), .Z(n18739) );
  NAND U19093 ( .A(a[246]), .B(n98), .Z(n18738) );
  AND U19094 ( .A(n18739), .B(n18738), .Z(n18809) );
  XNOR U19095 ( .A(n20154), .B(n18868), .Z(n18818) );
  OR U19096 ( .A(n18818), .B(n20057), .Z(n18742) );
  NANDN U19097 ( .A(n18740), .B(n20098), .Z(n18741) );
  AND U19098 ( .A(n18742), .B(n18741), .Z(n18810) );
  XOR U19099 ( .A(n18809), .B(n18810), .Z(n18812) );
  NAND U19100 ( .A(a[231]), .B(b[15]), .Z(n18811) );
  XOR U19101 ( .A(n18812), .B(n18811), .Z(n18830) );
  NAND U19102 ( .A(n19722), .B(n18743), .Z(n18745) );
  XOR U19103 ( .A(b[5]), .B(a[243]), .Z(n18821) );
  NANDN U19104 ( .A(n19640), .B(n18821), .Z(n18744) );
  NAND U19105 ( .A(n18745), .B(n18744), .Z(n18806) );
  XOR U19106 ( .A(n19714), .B(a[241]), .Z(n18824) );
  NANDN U19107 ( .A(n18824), .B(n19766), .Z(n18748) );
  NANDN U19108 ( .A(n18746), .B(n19767), .Z(n18747) );
  NAND U19109 ( .A(n18748), .B(n18747), .Z(n18803) );
  NAND U19110 ( .A(n19554), .B(n18749), .Z(n18751) );
  IV U19111 ( .A(a[245]), .Z(n19647) );
  XNOR U19112 ( .A(b[3]), .B(n19647), .Z(n18827) );
  NANDN U19113 ( .A(n19521), .B(n18827), .Z(n18750) );
  AND U19114 ( .A(n18751), .B(n18750), .Z(n18804) );
  XNOR U19115 ( .A(n18803), .B(n18804), .Z(n18805) );
  XOR U19116 ( .A(n18806), .B(n18805), .Z(n18831) );
  XOR U19117 ( .A(n18830), .B(n18831), .Z(n18832) );
  XNOR U19118 ( .A(n18833), .B(n18832), .Z(n18781) );
  NAND U19119 ( .A(n18753), .B(n18752), .Z(n18757) );
  NAND U19120 ( .A(n18755), .B(n18754), .Z(n18756) );
  NAND U19121 ( .A(n18757), .B(n18756), .Z(n18782) );
  XOR U19122 ( .A(n18781), .B(n18782), .Z(n18784) );
  XNOR U19123 ( .A(n18783), .B(n18784), .Z(n18842) );
  NANDN U19124 ( .A(n18759), .B(n18758), .Z(n18763) );
  NAND U19125 ( .A(n18761), .B(n18760), .Z(n18762) );
  NAND U19126 ( .A(n18763), .B(n18762), .Z(n18843) );
  XNOR U19127 ( .A(n18842), .B(n18843), .Z(n18844) );
  XOR U19128 ( .A(n18845), .B(n18844), .Z(n18775) );
  NANDN U19129 ( .A(n18765), .B(n18764), .Z(n18769) );
  NANDN U19130 ( .A(n18767), .B(n18766), .Z(n18768) );
  NAND U19131 ( .A(n18769), .B(n18768), .Z(n18776) );
  XNOR U19132 ( .A(n18775), .B(n18776), .Z(n18777) );
  XNOR U19133 ( .A(n18778), .B(n18777), .Z(n18848) );
  XNOR U19134 ( .A(n18848), .B(sreg[487]), .Z(n18850) );
  NAND U19135 ( .A(n18770), .B(sreg[486]), .Z(n18774) );
  OR U19136 ( .A(n18772), .B(n18771), .Z(n18773) );
  AND U19137 ( .A(n18774), .B(n18773), .Z(n18849) );
  XOR U19138 ( .A(n18850), .B(n18849), .Z(c[487]) );
  NANDN U19139 ( .A(n18776), .B(n18775), .Z(n18780) );
  NAND U19140 ( .A(n18778), .B(n18777), .Z(n18779) );
  NAND U19141 ( .A(n18780), .B(n18779), .Z(n18856) );
  NANDN U19142 ( .A(n18782), .B(n18781), .Z(n18786) );
  OR U19143 ( .A(n18784), .B(n18783), .Z(n18785) );
  NAND U19144 ( .A(n18786), .B(n18785), .Z(n18923) );
  XNOR U19145 ( .A(n20052), .B(n19128), .Z(n18865) );
  OR U19146 ( .A(n18865), .B(n20020), .Z(n18789) );
  NANDN U19147 ( .A(n18787), .B(n19960), .Z(n18788) );
  NAND U19148 ( .A(n18789), .B(n18788), .Z(n18878) );
  XNOR U19149 ( .A(n102), .B(n18790), .Z(n18869) );
  OR U19150 ( .A(n18869), .B(n20121), .Z(n18793) );
  NANDN U19151 ( .A(n18791), .B(n20122), .Z(n18792) );
  NAND U19152 ( .A(n18793), .B(n18792), .Z(n18875) );
  XOR U19153 ( .A(n19975), .B(a[240]), .Z(n18872) );
  NANDN U19154 ( .A(n18872), .B(n19883), .Z(n18796) );
  NANDN U19155 ( .A(n18794), .B(n19937), .Z(n18795) );
  AND U19156 ( .A(n18796), .B(n18795), .Z(n18876) );
  XNOR U19157 ( .A(n18875), .B(n18876), .Z(n18877) );
  XNOR U19158 ( .A(n18878), .B(n18877), .Z(n18914) );
  NANDN U19159 ( .A(n18798), .B(n18797), .Z(n18802) );
  NAND U19160 ( .A(n18800), .B(n18799), .Z(n18801) );
  NAND U19161 ( .A(n18802), .B(n18801), .Z(n18915) );
  XNOR U19162 ( .A(n18914), .B(n18915), .Z(n18916) );
  NANDN U19163 ( .A(n18804), .B(n18803), .Z(n18808) );
  NAND U19164 ( .A(n18806), .B(n18805), .Z(n18807) );
  AND U19165 ( .A(n18808), .B(n18807), .Z(n18917) );
  XNOR U19166 ( .A(n18916), .B(n18917), .Z(n18861) );
  NANDN U19167 ( .A(n18810), .B(n18809), .Z(n18814) );
  OR U19168 ( .A(n18812), .B(n18811), .Z(n18813) );
  NAND U19169 ( .A(n18814), .B(n18813), .Z(n18911) );
  NAND U19170 ( .A(b[0]), .B(a[248]), .Z(n18815) );
  XNOR U19171 ( .A(b[1]), .B(n18815), .Z(n18817) );
  NAND U19172 ( .A(a[247]), .B(n98), .Z(n18816) );
  AND U19173 ( .A(n18817), .B(n18816), .Z(n18887) );
  XNOR U19174 ( .A(n20154), .B(n18946), .Z(n18896) );
  OR U19175 ( .A(n18896), .B(n20057), .Z(n18820) );
  NANDN U19176 ( .A(n18818), .B(n20098), .Z(n18819) );
  AND U19177 ( .A(n18820), .B(n18819), .Z(n18888) );
  XOR U19178 ( .A(n18887), .B(n18888), .Z(n18890) );
  NAND U19179 ( .A(a[232]), .B(b[15]), .Z(n18889) );
  XOR U19180 ( .A(n18890), .B(n18889), .Z(n18908) );
  NAND U19181 ( .A(n19722), .B(n18821), .Z(n18823) );
  IV U19182 ( .A(a[244]), .Z(n19558) );
  XNOR U19183 ( .A(b[5]), .B(n19558), .Z(n18899) );
  NANDN U19184 ( .A(n19640), .B(n18899), .Z(n18822) );
  NAND U19185 ( .A(n18823), .B(n18822), .Z(n18884) );
  XNOR U19186 ( .A(n19714), .B(n19433), .Z(n18902) );
  NANDN U19187 ( .A(n18902), .B(n19766), .Z(n18826) );
  NANDN U19188 ( .A(n18824), .B(n19767), .Z(n18825) );
  NAND U19189 ( .A(n18826), .B(n18825), .Z(n18881) );
  NAND U19190 ( .A(n19554), .B(n18827), .Z(n18829) );
  XNOR U19191 ( .A(a[246]), .B(n100), .Z(n18905) );
  NANDN U19192 ( .A(n19521), .B(n18905), .Z(n18828) );
  AND U19193 ( .A(n18829), .B(n18828), .Z(n18882) );
  XNOR U19194 ( .A(n18881), .B(n18882), .Z(n18883) );
  XOR U19195 ( .A(n18884), .B(n18883), .Z(n18909) );
  XOR U19196 ( .A(n18908), .B(n18909), .Z(n18910) );
  XNOR U19197 ( .A(n18911), .B(n18910), .Z(n18859) );
  NAND U19198 ( .A(n18831), .B(n18830), .Z(n18835) );
  NAND U19199 ( .A(n18833), .B(n18832), .Z(n18834) );
  NAND U19200 ( .A(n18835), .B(n18834), .Z(n18860) );
  XOR U19201 ( .A(n18859), .B(n18860), .Z(n18862) );
  XNOR U19202 ( .A(n18861), .B(n18862), .Z(n18920) );
  NANDN U19203 ( .A(n18837), .B(n18836), .Z(n18841) );
  NAND U19204 ( .A(n18839), .B(n18838), .Z(n18840) );
  NAND U19205 ( .A(n18841), .B(n18840), .Z(n18921) );
  XNOR U19206 ( .A(n18920), .B(n18921), .Z(n18922) );
  XOR U19207 ( .A(n18923), .B(n18922), .Z(n18853) );
  NANDN U19208 ( .A(n18843), .B(n18842), .Z(n18847) );
  NANDN U19209 ( .A(n18845), .B(n18844), .Z(n18846) );
  NAND U19210 ( .A(n18847), .B(n18846), .Z(n18854) );
  XNOR U19211 ( .A(n18853), .B(n18854), .Z(n18855) );
  XNOR U19212 ( .A(n18856), .B(n18855), .Z(n18926) );
  XNOR U19213 ( .A(n18926), .B(sreg[488]), .Z(n18928) );
  NAND U19214 ( .A(n18848), .B(sreg[487]), .Z(n18852) );
  OR U19215 ( .A(n18850), .B(n18849), .Z(n18851) );
  AND U19216 ( .A(n18852), .B(n18851), .Z(n18927) );
  XOR U19217 ( .A(n18928), .B(n18927), .Z(c[488]) );
  NANDN U19218 ( .A(n18854), .B(n18853), .Z(n18858) );
  NAND U19219 ( .A(n18856), .B(n18855), .Z(n18857) );
  NAND U19220 ( .A(n18858), .B(n18857), .Z(n18934) );
  NANDN U19221 ( .A(n18860), .B(n18859), .Z(n18864) );
  OR U19222 ( .A(n18862), .B(n18861), .Z(n18863) );
  NAND U19223 ( .A(n18864), .B(n18863), .Z(n19001) );
  XOR U19224 ( .A(n20052), .B(a[239]), .Z(n18943) );
  OR U19225 ( .A(n18943), .B(n20020), .Z(n18867) );
  NANDN U19226 ( .A(n18865), .B(n19960), .Z(n18866) );
  NAND U19227 ( .A(n18867), .B(n18866), .Z(n18956) );
  XNOR U19228 ( .A(n102), .B(n18868), .Z(n18947) );
  OR U19229 ( .A(n18947), .B(n20121), .Z(n18871) );
  NANDN U19230 ( .A(n18869), .B(n20122), .Z(n18870) );
  NAND U19231 ( .A(n18871), .B(n18870), .Z(n18953) );
  XOR U19232 ( .A(n19975), .B(a[241]), .Z(n18950) );
  NANDN U19233 ( .A(n18950), .B(n19883), .Z(n18874) );
  NANDN U19234 ( .A(n18872), .B(n19937), .Z(n18873) );
  AND U19235 ( .A(n18874), .B(n18873), .Z(n18954) );
  XNOR U19236 ( .A(n18953), .B(n18954), .Z(n18955) );
  XNOR U19237 ( .A(n18956), .B(n18955), .Z(n18992) );
  NANDN U19238 ( .A(n18876), .B(n18875), .Z(n18880) );
  NAND U19239 ( .A(n18878), .B(n18877), .Z(n18879) );
  NAND U19240 ( .A(n18880), .B(n18879), .Z(n18993) );
  XNOR U19241 ( .A(n18992), .B(n18993), .Z(n18994) );
  NANDN U19242 ( .A(n18882), .B(n18881), .Z(n18886) );
  NAND U19243 ( .A(n18884), .B(n18883), .Z(n18885) );
  AND U19244 ( .A(n18886), .B(n18885), .Z(n18995) );
  XNOR U19245 ( .A(n18994), .B(n18995), .Z(n18939) );
  NANDN U19246 ( .A(n18888), .B(n18887), .Z(n18892) );
  OR U19247 ( .A(n18890), .B(n18889), .Z(n18891) );
  NAND U19248 ( .A(n18892), .B(n18891), .Z(n18989) );
  NAND U19249 ( .A(b[0]), .B(a[249]), .Z(n18893) );
  XNOR U19250 ( .A(b[1]), .B(n18893), .Z(n18895) );
  NAND U19251 ( .A(a[248]), .B(n98), .Z(n18894) );
  AND U19252 ( .A(n18895), .B(n18894), .Z(n18965) );
  XOR U19253 ( .A(n20154), .B(a[237]), .Z(n18974) );
  OR U19254 ( .A(n18974), .B(n20057), .Z(n18898) );
  NANDN U19255 ( .A(n18896), .B(n20098), .Z(n18897) );
  AND U19256 ( .A(n18898), .B(n18897), .Z(n18966) );
  XOR U19257 ( .A(n18965), .B(n18966), .Z(n18968) );
  NAND U19258 ( .A(a[233]), .B(b[15]), .Z(n18967) );
  XOR U19259 ( .A(n18968), .B(n18967), .Z(n18986) );
  NAND U19260 ( .A(n19722), .B(n18899), .Z(n18901) );
  XNOR U19261 ( .A(b[5]), .B(n19647), .Z(n18977) );
  NANDN U19262 ( .A(n19640), .B(n18977), .Z(n18900) );
  NAND U19263 ( .A(n18901), .B(n18900), .Z(n18962) );
  XOR U19264 ( .A(n19714), .B(a[243]), .Z(n18980) );
  NANDN U19265 ( .A(n18980), .B(n19766), .Z(n18904) );
  NANDN U19266 ( .A(n18902), .B(n19767), .Z(n18903) );
  NAND U19267 ( .A(n18904), .B(n18903), .Z(n18959) );
  NAND U19268 ( .A(n19554), .B(n18905), .Z(n18907) );
  XNOR U19269 ( .A(a[247]), .B(n100), .Z(n18983) );
  NANDN U19270 ( .A(n19521), .B(n18983), .Z(n18906) );
  AND U19271 ( .A(n18907), .B(n18906), .Z(n18960) );
  XNOR U19272 ( .A(n18959), .B(n18960), .Z(n18961) );
  XOR U19273 ( .A(n18962), .B(n18961), .Z(n18987) );
  XOR U19274 ( .A(n18986), .B(n18987), .Z(n18988) );
  XNOR U19275 ( .A(n18989), .B(n18988), .Z(n18937) );
  NAND U19276 ( .A(n18909), .B(n18908), .Z(n18913) );
  NAND U19277 ( .A(n18911), .B(n18910), .Z(n18912) );
  NAND U19278 ( .A(n18913), .B(n18912), .Z(n18938) );
  XOR U19279 ( .A(n18937), .B(n18938), .Z(n18940) );
  XNOR U19280 ( .A(n18939), .B(n18940), .Z(n18998) );
  NANDN U19281 ( .A(n18915), .B(n18914), .Z(n18919) );
  NAND U19282 ( .A(n18917), .B(n18916), .Z(n18918) );
  NAND U19283 ( .A(n18919), .B(n18918), .Z(n18999) );
  XNOR U19284 ( .A(n18998), .B(n18999), .Z(n19000) );
  XOR U19285 ( .A(n19001), .B(n19000), .Z(n18931) );
  NANDN U19286 ( .A(n18921), .B(n18920), .Z(n18925) );
  NANDN U19287 ( .A(n18923), .B(n18922), .Z(n18924) );
  NAND U19288 ( .A(n18925), .B(n18924), .Z(n18932) );
  XNOR U19289 ( .A(n18931), .B(n18932), .Z(n18933) );
  XNOR U19290 ( .A(n18934), .B(n18933), .Z(n19004) );
  XNOR U19291 ( .A(n19004), .B(sreg[489]), .Z(n19006) );
  NAND U19292 ( .A(n18926), .B(sreg[488]), .Z(n18930) );
  OR U19293 ( .A(n18928), .B(n18927), .Z(n18929) );
  AND U19294 ( .A(n18930), .B(n18929), .Z(n19005) );
  XOR U19295 ( .A(n19006), .B(n19005), .Z(c[489]) );
  NANDN U19296 ( .A(n18932), .B(n18931), .Z(n18936) );
  NAND U19297 ( .A(n18934), .B(n18933), .Z(n18935) );
  NAND U19298 ( .A(n18936), .B(n18935), .Z(n19012) );
  NANDN U19299 ( .A(n18938), .B(n18937), .Z(n18942) );
  OR U19300 ( .A(n18940), .B(n18939), .Z(n18941) );
  NAND U19301 ( .A(n18942), .B(n18941), .Z(n19078) );
  XOR U19302 ( .A(n20052), .B(a[240]), .Z(n19021) );
  OR U19303 ( .A(n19021), .B(n20020), .Z(n18945) );
  NANDN U19304 ( .A(n18943), .B(n19960), .Z(n18944) );
  NAND U19305 ( .A(n18945), .B(n18944), .Z(n19033) );
  XNOR U19306 ( .A(n102), .B(n18946), .Z(n19024) );
  OR U19307 ( .A(n19024), .B(n20121), .Z(n18949) );
  NANDN U19308 ( .A(n18947), .B(n20122), .Z(n18948) );
  NAND U19309 ( .A(n18949), .B(n18948), .Z(n19030) );
  XNOR U19310 ( .A(n19975), .B(n19433), .Z(n19027) );
  NANDN U19311 ( .A(n19027), .B(n19883), .Z(n18952) );
  NANDN U19312 ( .A(n18950), .B(n19937), .Z(n18951) );
  AND U19313 ( .A(n18952), .B(n18951), .Z(n19031) );
  XNOR U19314 ( .A(n19030), .B(n19031), .Z(n19032) );
  XNOR U19315 ( .A(n19033), .B(n19032), .Z(n19069) );
  NANDN U19316 ( .A(n18954), .B(n18953), .Z(n18958) );
  NAND U19317 ( .A(n18956), .B(n18955), .Z(n18957) );
  NAND U19318 ( .A(n18958), .B(n18957), .Z(n19070) );
  XNOR U19319 ( .A(n19069), .B(n19070), .Z(n19071) );
  NANDN U19320 ( .A(n18960), .B(n18959), .Z(n18964) );
  NAND U19321 ( .A(n18962), .B(n18961), .Z(n18963) );
  AND U19322 ( .A(n18964), .B(n18963), .Z(n19072) );
  XNOR U19323 ( .A(n19071), .B(n19072), .Z(n19017) );
  NANDN U19324 ( .A(n18966), .B(n18965), .Z(n18970) );
  OR U19325 ( .A(n18968), .B(n18967), .Z(n18969) );
  NAND U19326 ( .A(n18970), .B(n18969), .Z(n19066) );
  NAND U19327 ( .A(b[0]), .B(a[250]), .Z(n18971) );
  XNOR U19328 ( .A(b[1]), .B(n18971), .Z(n18973) );
  NAND U19329 ( .A(n98), .B(a[249]), .Z(n18972) );
  AND U19330 ( .A(n18973), .B(n18972), .Z(n19042) );
  XNOR U19331 ( .A(n20154), .B(n19128), .Z(n19051) );
  OR U19332 ( .A(n19051), .B(n20057), .Z(n18976) );
  NANDN U19333 ( .A(n18974), .B(n20098), .Z(n18975) );
  AND U19334 ( .A(n18976), .B(n18975), .Z(n19043) );
  XOR U19335 ( .A(n19042), .B(n19043), .Z(n19045) );
  NAND U19336 ( .A(a[234]), .B(b[15]), .Z(n19044) );
  XOR U19337 ( .A(n19045), .B(n19044), .Z(n19063) );
  NAND U19338 ( .A(n19722), .B(n18977), .Z(n18979) );
  IV U19339 ( .A(a[246]), .Z(n19576) );
  XNOR U19340 ( .A(b[5]), .B(n19576), .Z(n19054) );
  NANDN U19341 ( .A(n19640), .B(n19054), .Z(n18978) );
  NAND U19342 ( .A(n18979), .B(n18978), .Z(n19039) );
  XNOR U19343 ( .A(n19714), .B(n19558), .Z(n19057) );
  NANDN U19344 ( .A(n19057), .B(n19766), .Z(n18982) );
  NANDN U19345 ( .A(n18980), .B(n19767), .Z(n18981) );
  NAND U19346 ( .A(n18982), .B(n18981), .Z(n19036) );
  NAND U19347 ( .A(n19554), .B(n18983), .Z(n18985) );
  XNOR U19348 ( .A(a[248]), .B(n100), .Z(n19060) );
  NANDN U19349 ( .A(n19521), .B(n19060), .Z(n18984) );
  AND U19350 ( .A(n18985), .B(n18984), .Z(n19037) );
  XNOR U19351 ( .A(n19036), .B(n19037), .Z(n19038) );
  XOR U19352 ( .A(n19039), .B(n19038), .Z(n19064) );
  XOR U19353 ( .A(n19063), .B(n19064), .Z(n19065) );
  XNOR U19354 ( .A(n19066), .B(n19065), .Z(n19015) );
  NAND U19355 ( .A(n18987), .B(n18986), .Z(n18991) );
  NAND U19356 ( .A(n18989), .B(n18988), .Z(n18990) );
  NAND U19357 ( .A(n18991), .B(n18990), .Z(n19016) );
  XOR U19358 ( .A(n19015), .B(n19016), .Z(n19018) );
  XNOR U19359 ( .A(n19017), .B(n19018), .Z(n19075) );
  NANDN U19360 ( .A(n18993), .B(n18992), .Z(n18997) );
  NAND U19361 ( .A(n18995), .B(n18994), .Z(n18996) );
  NAND U19362 ( .A(n18997), .B(n18996), .Z(n19076) );
  XNOR U19363 ( .A(n19075), .B(n19076), .Z(n19077) );
  XOR U19364 ( .A(n19078), .B(n19077), .Z(n19009) );
  NANDN U19365 ( .A(n18999), .B(n18998), .Z(n19003) );
  NANDN U19366 ( .A(n19001), .B(n19000), .Z(n19002) );
  NAND U19367 ( .A(n19003), .B(n19002), .Z(n19010) );
  XNOR U19368 ( .A(n19009), .B(n19010), .Z(n19011) );
  XNOR U19369 ( .A(n19012), .B(n19011), .Z(n19081) );
  XNOR U19370 ( .A(n19081), .B(sreg[490]), .Z(n19083) );
  NAND U19371 ( .A(n19004), .B(sreg[489]), .Z(n19008) );
  OR U19372 ( .A(n19006), .B(n19005), .Z(n19007) );
  AND U19373 ( .A(n19008), .B(n19007), .Z(n19082) );
  XOR U19374 ( .A(n19083), .B(n19082), .Z(c[490]) );
  NANDN U19375 ( .A(n19010), .B(n19009), .Z(n19014) );
  NAND U19376 ( .A(n19012), .B(n19011), .Z(n19013) );
  NAND U19377 ( .A(n19014), .B(n19013), .Z(n19089) );
  NANDN U19378 ( .A(n19016), .B(n19015), .Z(n19020) );
  OR U19379 ( .A(n19018), .B(n19017), .Z(n19019) );
  NAND U19380 ( .A(n19020), .B(n19019), .Z(n19156) );
  XOR U19381 ( .A(n20052), .B(a[241]), .Z(n19125) );
  OR U19382 ( .A(n19125), .B(n20020), .Z(n19023) );
  NANDN U19383 ( .A(n19021), .B(n19960), .Z(n19022) );
  NAND U19384 ( .A(n19023), .B(n19022), .Z(n19138) );
  XOR U19385 ( .A(n102), .B(a[237]), .Z(n19129) );
  OR U19386 ( .A(n19129), .B(n20121), .Z(n19026) );
  NANDN U19387 ( .A(n19024), .B(n20122), .Z(n19025) );
  NAND U19388 ( .A(n19026), .B(n19025), .Z(n19135) );
  XOR U19389 ( .A(n19975), .B(a[243]), .Z(n19132) );
  NANDN U19390 ( .A(n19132), .B(n19883), .Z(n19029) );
  NANDN U19391 ( .A(n19027), .B(n19937), .Z(n19028) );
  AND U19392 ( .A(n19029), .B(n19028), .Z(n19136) );
  XNOR U19393 ( .A(n19135), .B(n19136), .Z(n19137) );
  XNOR U19394 ( .A(n19138), .B(n19137), .Z(n19147) );
  NANDN U19395 ( .A(n19031), .B(n19030), .Z(n19035) );
  NAND U19396 ( .A(n19033), .B(n19032), .Z(n19034) );
  NAND U19397 ( .A(n19035), .B(n19034), .Z(n19148) );
  XNOR U19398 ( .A(n19147), .B(n19148), .Z(n19149) );
  NANDN U19399 ( .A(n19037), .B(n19036), .Z(n19041) );
  NAND U19400 ( .A(n19039), .B(n19038), .Z(n19040) );
  AND U19401 ( .A(n19041), .B(n19040), .Z(n19150) );
  XNOR U19402 ( .A(n19149), .B(n19150), .Z(n19094) );
  NANDN U19403 ( .A(n19043), .B(n19042), .Z(n19047) );
  OR U19404 ( .A(n19045), .B(n19044), .Z(n19046) );
  NAND U19405 ( .A(n19047), .B(n19046), .Z(n19122) );
  NAND U19406 ( .A(b[0]), .B(a[251]), .Z(n19048) );
  XNOR U19407 ( .A(b[1]), .B(n19048), .Z(n19050) );
  NAND U19408 ( .A(a[250]), .B(n98), .Z(n19049) );
  AND U19409 ( .A(n19050), .B(n19049), .Z(n19098) );
  XOR U19410 ( .A(n20154), .B(a[239]), .Z(n19104) );
  OR U19411 ( .A(n19104), .B(n20057), .Z(n19053) );
  NANDN U19412 ( .A(n19051), .B(n20098), .Z(n19052) );
  AND U19413 ( .A(n19053), .B(n19052), .Z(n19099) );
  XOR U19414 ( .A(n19098), .B(n19099), .Z(n19101) );
  NAND U19415 ( .A(a[235]), .B(b[15]), .Z(n19100) );
  XOR U19416 ( .A(n19101), .B(n19100), .Z(n19119) );
  NAND U19417 ( .A(n19722), .B(n19054), .Z(n19056) );
  IV U19418 ( .A(a[247]), .Z(n19775) );
  XNOR U19419 ( .A(b[5]), .B(n19775), .Z(n19110) );
  NANDN U19420 ( .A(n19640), .B(n19110), .Z(n19055) );
  NAND U19421 ( .A(n19056), .B(n19055), .Z(n19144) );
  XNOR U19422 ( .A(n19714), .B(n19647), .Z(n19113) );
  NANDN U19423 ( .A(n19113), .B(n19766), .Z(n19059) );
  NANDN U19424 ( .A(n19057), .B(n19767), .Z(n19058) );
  NAND U19425 ( .A(n19059), .B(n19058), .Z(n19141) );
  NAND U19426 ( .A(n19554), .B(n19060), .Z(n19062) );
  XOR U19427 ( .A(a[249]), .B(b[3]), .Z(n19116) );
  NANDN U19428 ( .A(n19521), .B(n19116), .Z(n19061) );
  AND U19429 ( .A(n19062), .B(n19061), .Z(n19142) );
  XNOR U19430 ( .A(n19141), .B(n19142), .Z(n19143) );
  XOR U19431 ( .A(n19144), .B(n19143), .Z(n19120) );
  XOR U19432 ( .A(n19119), .B(n19120), .Z(n19121) );
  XNOR U19433 ( .A(n19122), .B(n19121), .Z(n19092) );
  NAND U19434 ( .A(n19064), .B(n19063), .Z(n19068) );
  NAND U19435 ( .A(n19066), .B(n19065), .Z(n19067) );
  NAND U19436 ( .A(n19068), .B(n19067), .Z(n19093) );
  XOR U19437 ( .A(n19092), .B(n19093), .Z(n19095) );
  XNOR U19438 ( .A(n19094), .B(n19095), .Z(n19153) );
  NANDN U19439 ( .A(n19070), .B(n19069), .Z(n19074) );
  NAND U19440 ( .A(n19072), .B(n19071), .Z(n19073) );
  NAND U19441 ( .A(n19074), .B(n19073), .Z(n19154) );
  XNOR U19442 ( .A(n19153), .B(n19154), .Z(n19155) );
  XOR U19443 ( .A(n19156), .B(n19155), .Z(n19086) );
  NANDN U19444 ( .A(n19076), .B(n19075), .Z(n19080) );
  NANDN U19445 ( .A(n19078), .B(n19077), .Z(n19079) );
  NAND U19446 ( .A(n19080), .B(n19079), .Z(n19087) );
  XNOR U19447 ( .A(n19086), .B(n19087), .Z(n19088) );
  XNOR U19448 ( .A(n19089), .B(n19088), .Z(n19159) );
  XNOR U19449 ( .A(n19159), .B(sreg[491]), .Z(n19161) );
  NAND U19450 ( .A(n19081), .B(sreg[490]), .Z(n19085) );
  OR U19451 ( .A(n19083), .B(n19082), .Z(n19084) );
  AND U19452 ( .A(n19085), .B(n19084), .Z(n19160) );
  XOR U19453 ( .A(n19161), .B(n19160), .Z(c[491]) );
  NANDN U19454 ( .A(n19087), .B(n19086), .Z(n19091) );
  NAND U19455 ( .A(n19089), .B(n19088), .Z(n19090) );
  NAND U19456 ( .A(n19091), .B(n19090), .Z(n19167) );
  NANDN U19457 ( .A(n19093), .B(n19092), .Z(n19097) );
  OR U19458 ( .A(n19095), .B(n19094), .Z(n19096) );
  NAND U19459 ( .A(n19097), .B(n19096), .Z(n19233) );
  NANDN U19460 ( .A(n19099), .B(n19098), .Z(n19103) );
  OR U19461 ( .A(n19101), .B(n19100), .Z(n19102) );
  NAND U19462 ( .A(n19103), .B(n19102), .Z(n19221) );
  XOR U19463 ( .A(n20154), .B(a[240]), .Z(n19206) );
  OR U19464 ( .A(n19206), .B(n20057), .Z(n19106) );
  NANDN U19465 ( .A(n19104), .B(n20098), .Z(n19105) );
  AND U19466 ( .A(n19106), .B(n19105), .Z(n19198) );
  NAND U19467 ( .A(b[0]), .B(a[252]), .Z(n19107) );
  XNOR U19468 ( .A(b[1]), .B(n19107), .Z(n19109) );
  NAND U19469 ( .A(n98), .B(a[251]), .Z(n19108) );
  AND U19470 ( .A(n19109), .B(n19108), .Z(n19197) );
  XOR U19471 ( .A(n19198), .B(n19197), .Z(n19200) );
  NAND U19472 ( .A(a[236]), .B(b[15]), .Z(n19199) );
  XOR U19473 ( .A(n19200), .B(n19199), .Z(n19218) );
  NAND U19474 ( .A(n19722), .B(n19110), .Z(n19112) );
  XNOR U19475 ( .A(a[248]), .B(n101), .Z(n19212) );
  NANDN U19476 ( .A(n19640), .B(n19212), .Z(n19111) );
  NAND U19477 ( .A(n19112), .B(n19111), .Z(n19194) );
  XNOR U19478 ( .A(n19714), .B(n19576), .Z(n19215) );
  NANDN U19479 ( .A(n19215), .B(n19766), .Z(n19115) );
  NANDN U19480 ( .A(n19113), .B(n19767), .Z(n19114) );
  NAND U19481 ( .A(n19115), .B(n19114), .Z(n19191) );
  NAND U19482 ( .A(n19554), .B(n19116), .Z(n19118) );
  XNOR U19483 ( .A(a[250]), .B(n100), .Z(n19209) );
  NANDN U19484 ( .A(n19521), .B(n19209), .Z(n19117) );
  AND U19485 ( .A(n19118), .B(n19117), .Z(n19192) );
  XNOR U19486 ( .A(n19191), .B(n19192), .Z(n19193) );
  XOR U19487 ( .A(n19194), .B(n19193), .Z(n19219) );
  XOR U19488 ( .A(n19218), .B(n19219), .Z(n19220) );
  XNOR U19489 ( .A(n19221), .B(n19220), .Z(n19170) );
  NAND U19490 ( .A(n19120), .B(n19119), .Z(n19124) );
  NAND U19491 ( .A(n19122), .B(n19121), .Z(n19123) );
  NAND U19492 ( .A(n19124), .B(n19123), .Z(n19171) );
  XOR U19493 ( .A(n19170), .B(n19171), .Z(n19173) );
  XNOR U19494 ( .A(n20052), .B(n19433), .Z(n19179) );
  OR U19495 ( .A(n19179), .B(n20020), .Z(n19127) );
  NANDN U19496 ( .A(n19125), .B(n19960), .Z(n19126) );
  NAND U19497 ( .A(n19127), .B(n19126), .Z(n19188) );
  XNOR U19498 ( .A(n102), .B(n19128), .Z(n19182) );
  OR U19499 ( .A(n19182), .B(n20121), .Z(n19131) );
  NANDN U19500 ( .A(n19129), .B(n20122), .Z(n19130) );
  NAND U19501 ( .A(n19131), .B(n19130), .Z(n19185) );
  XNOR U19502 ( .A(n19975), .B(n19558), .Z(n19176) );
  NANDN U19503 ( .A(n19176), .B(n19883), .Z(n19134) );
  NANDN U19504 ( .A(n19132), .B(n19937), .Z(n19133) );
  AND U19505 ( .A(n19134), .B(n19133), .Z(n19186) );
  XNOR U19506 ( .A(n19185), .B(n19186), .Z(n19187) );
  XNOR U19507 ( .A(n19188), .B(n19187), .Z(n19224) );
  NANDN U19508 ( .A(n19136), .B(n19135), .Z(n19140) );
  NAND U19509 ( .A(n19138), .B(n19137), .Z(n19139) );
  NAND U19510 ( .A(n19140), .B(n19139), .Z(n19225) );
  XNOR U19511 ( .A(n19224), .B(n19225), .Z(n19226) );
  NANDN U19512 ( .A(n19142), .B(n19141), .Z(n19146) );
  NAND U19513 ( .A(n19144), .B(n19143), .Z(n19145) );
  AND U19514 ( .A(n19146), .B(n19145), .Z(n19227) );
  XNOR U19515 ( .A(n19226), .B(n19227), .Z(n19172) );
  XNOR U19516 ( .A(n19173), .B(n19172), .Z(n19230) );
  NANDN U19517 ( .A(n19148), .B(n19147), .Z(n19152) );
  NAND U19518 ( .A(n19150), .B(n19149), .Z(n19151) );
  NAND U19519 ( .A(n19152), .B(n19151), .Z(n19231) );
  XNOR U19520 ( .A(n19230), .B(n19231), .Z(n19232) );
  XOR U19521 ( .A(n19233), .B(n19232), .Z(n19164) );
  NANDN U19522 ( .A(n19154), .B(n19153), .Z(n19158) );
  NANDN U19523 ( .A(n19156), .B(n19155), .Z(n19157) );
  NAND U19524 ( .A(n19158), .B(n19157), .Z(n19165) );
  XNOR U19525 ( .A(n19164), .B(n19165), .Z(n19166) );
  XNOR U19526 ( .A(n19167), .B(n19166), .Z(n19236) );
  XNOR U19527 ( .A(n19236), .B(sreg[492]), .Z(n19238) );
  NAND U19528 ( .A(n19159), .B(sreg[491]), .Z(n19163) );
  OR U19529 ( .A(n19161), .B(n19160), .Z(n19162) );
  AND U19530 ( .A(n19163), .B(n19162), .Z(n19237) );
  XOR U19531 ( .A(n19238), .B(n19237), .Z(c[492]) );
  NANDN U19532 ( .A(n19165), .B(n19164), .Z(n19169) );
  NAND U19533 ( .A(n19167), .B(n19166), .Z(n19168) );
  NAND U19534 ( .A(n19169), .B(n19168), .Z(n19244) );
  NANDN U19535 ( .A(n19171), .B(n19170), .Z(n19175) );
  OR U19536 ( .A(n19173), .B(n19172), .Z(n19174) );
  NAND U19537 ( .A(n19175), .B(n19174), .Z(n19310) );
  XNOR U19538 ( .A(n19975), .B(n19647), .Z(n19280) );
  NANDN U19539 ( .A(n19280), .B(n19883), .Z(n19178) );
  NANDN U19540 ( .A(n19176), .B(n19937), .Z(n19177) );
  NAND U19541 ( .A(n19178), .B(n19177), .Z(n19277) );
  XOR U19542 ( .A(n20052), .B(a[243]), .Z(n19283) );
  OR U19543 ( .A(n19283), .B(n20020), .Z(n19181) );
  NANDN U19544 ( .A(n19179), .B(n19960), .Z(n19180) );
  NAND U19545 ( .A(n19181), .B(n19180), .Z(n19274) );
  XOR U19546 ( .A(n102), .B(a[239]), .Z(n19286) );
  OR U19547 ( .A(n19286), .B(n20121), .Z(n19184) );
  NANDN U19548 ( .A(n19182), .B(n20122), .Z(n19183) );
  AND U19549 ( .A(n19184), .B(n19183), .Z(n19275) );
  XNOR U19550 ( .A(n19274), .B(n19275), .Z(n19276) );
  XNOR U19551 ( .A(n19277), .B(n19276), .Z(n19301) );
  NANDN U19552 ( .A(n19186), .B(n19185), .Z(n19190) );
  NAND U19553 ( .A(n19188), .B(n19187), .Z(n19189) );
  NAND U19554 ( .A(n19190), .B(n19189), .Z(n19302) );
  XNOR U19555 ( .A(n19301), .B(n19302), .Z(n19303) );
  NANDN U19556 ( .A(n19192), .B(n19191), .Z(n19196) );
  NAND U19557 ( .A(n19194), .B(n19193), .Z(n19195) );
  AND U19558 ( .A(n19196), .B(n19195), .Z(n19304) );
  XNOR U19559 ( .A(n19303), .B(n19304), .Z(n19249) );
  NANDN U19560 ( .A(n19198), .B(n19197), .Z(n19202) );
  OR U19561 ( .A(n19200), .B(n19199), .Z(n19201) );
  NAND U19562 ( .A(n19202), .B(n19201), .Z(n19298) );
  NAND U19563 ( .A(b[0]), .B(a[253]), .Z(n19203) );
  XNOR U19564 ( .A(b[1]), .B(n19203), .Z(n19205) );
  NAND U19565 ( .A(a[252]), .B(n98), .Z(n19204) );
  AND U19566 ( .A(n19205), .B(n19204), .Z(n19255) );
  XOR U19567 ( .A(b[13]), .B(a[241]), .Z(n19262) );
  NANDN U19568 ( .A(n20057), .B(n19262), .Z(n19208) );
  NANDN U19569 ( .A(n19206), .B(n20098), .Z(n19207) );
  NAND U19570 ( .A(n19208), .B(n19207), .Z(n19253) );
  NAND U19571 ( .A(b[15]), .B(a[237]), .Z(n19254) );
  XNOR U19572 ( .A(n19253), .B(n19254), .Z(n19256) );
  XOR U19573 ( .A(n19255), .B(n19256), .Z(n19295) );
  NAND U19574 ( .A(n19554), .B(n19209), .Z(n19211) );
  XOR U19575 ( .A(a[251]), .B(b[3]), .Z(n19265) );
  NANDN U19576 ( .A(n19521), .B(n19265), .Z(n19210) );
  NAND U19577 ( .A(n19211), .B(n19210), .Z(n19291) );
  NAND U19578 ( .A(n19722), .B(n19212), .Z(n19214) );
  XOR U19579 ( .A(a[249]), .B(b[5]), .Z(n19268) );
  NANDN U19580 ( .A(n19640), .B(n19268), .Z(n19213) );
  NAND U19581 ( .A(n19214), .B(n19213), .Z(n19289) );
  XNOR U19582 ( .A(n19714), .B(n19775), .Z(n19271) );
  NANDN U19583 ( .A(n19271), .B(n19766), .Z(n19217) );
  NANDN U19584 ( .A(n19215), .B(n19767), .Z(n19216) );
  AND U19585 ( .A(n19217), .B(n19216), .Z(n19290) );
  XOR U19586 ( .A(n19291), .B(n19292), .Z(n19296) );
  XNOR U19587 ( .A(n19295), .B(n19296), .Z(n19297) );
  XNOR U19588 ( .A(n19298), .B(n19297), .Z(n19247) );
  NAND U19589 ( .A(n19219), .B(n19218), .Z(n19223) );
  NAND U19590 ( .A(n19221), .B(n19220), .Z(n19222) );
  NAND U19591 ( .A(n19223), .B(n19222), .Z(n19248) );
  XOR U19592 ( .A(n19247), .B(n19248), .Z(n19250) );
  XNOR U19593 ( .A(n19249), .B(n19250), .Z(n19307) );
  NANDN U19594 ( .A(n19225), .B(n19224), .Z(n19229) );
  NAND U19595 ( .A(n19227), .B(n19226), .Z(n19228) );
  NAND U19596 ( .A(n19229), .B(n19228), .Z(n19308) );
  XNOR U19597 ( .A(n19307), .B(n19308), .Z(n19309) );
  XOR U19598 ( .A(n19310), .B(n19309), .Z(n19241) );
  NANDN U19599 ( .A(n19231), .B(n19230), .Z(n19235) );
  NANDN U19600 ( .A(n19233), .B(n19232), .Z(n19234) );
  NAND U19601 ( .A(n19235), .B(n19234), .Z(n19242) );
  XNOR U19602 ( .A(n19241), .B(n19242), .Z(n19243) );
  XNOR U19603 ( .A(n19244), .B(n19243), .Z(n19313) );
  XNOR U19604 ( .A(n19313), .B(sreg[493]), .Z(n19315) );
  NAND U19605 ( .A(n19236), .B(sreg[492]), .Z(n19240) );
  OR U19606 ( .A(n19238), .B(n19237), .Z(n19239) );
  AND U19607 ( .A(n19240), .B(n19239), .Z(n19314) );
  XOR U19608 ( .A(n19315), .B(n19314), .Z(c[493]) );
  NANDN U19609 ( .A(n19242), .B(n19241), .Z(n19246) );
  NAND U19610 ( .A(n19244), .B(n19243), .Z(n19245) );
  NAND U19611 ( .A(n19246), .B(n19245), .Z(n19321) );
  NANDN U19612 ( .A(n19248), .B(n19247), .Z(n19252) );
  OR U19613 ( .A(n19250), .B(n19249), .Z(n19251) );
  NAND U19614 ( .A(n19252), .B(n19251), .Z(n19327) );
  NANDN U19615 ( .A(n19254), .B(n19253), .Z(n19258) );
  NAND U19616 ( .A(n19256), .B(n19255), .Z(n19257) );
  NAND U19617 ( .A(n19258), .B(n19257), .Z(n19375) );
  AND U19618 ( .A(b[15]), .B(a[238]), .Z(n19369) );
  NAND U19619 ( .A(b[0]), .B(a[254]), .Z(n19259) );
  XNOR U19620 ( .A(b[1]), .B(n19259), .Z(n19261) );
  NAND U19621 ( .A(n98), .B(a[253]), .Z(n19260) );
  AND U19622 ( .A(n19261), .B(n19260), .Z(n19367) );
  NAND U19623 ( .A(n20098), .B(n19262), .Z(n19264) );
  XOR U19624 ( .A(b[13]), .B(a[242]), .Z(n19354) );
  NANDN U19625 ( .A(n20057), .B(n19354), .Z(n19263) );
  AND U19626 ( .A(n19264), .B(n19263), .Z(n19366) );
  XNOR U19627 ( .A(n19367), .B(n19366), .Z(n19368) );
  XOR U19628 ( .A(n19369), .B(n19368), .Z(n19372) );
  NAND U19629 ( .A(n19554), .B(n19265), .Z(n19267) );
  XNOR U19630 ( .A(a[252]), .B(n100), .Z(n19357) );
  NANDN U19631 ( .A(n19521), .B(n19357), .Z(n19266) );
  NAND U19632 ( .A(n19267), .B(n19266), .Z(n19348) );
  NAND U19633 ( .A(n19722), .B(n19268), .Z(n19270) );
  XNOR U19634 ( .A(a[250]), .B(n101), .Z(n19360) );
  NANDN U19635 ( .A(n19640), .B(n19360), .Z(n19269) );
  NAND U19636 ( .A(n19270), .B(n19269), .Z(n19345) );
  IV U19637 ( .A(a[248]), .Z(n19562) );
  XNOR U19638 ( .A(n19714), .B(n19562), .Z(n19363) );
  NANDN U19639 ( .A(n19363), .B(n19766), .Z(n19273) );
  NANDN U19640 ( .A(n19271), .B(n19767), .Z(n19272) );
  AND U19641 ( .A(n19273), .B(n19272), .Z(n19346) );
  XNOR U19642 ( .A(n19345), .B(n19346), .Z(n19347) );
  XNOR U19643 ( .A(n19348), .B(n19347), .Z(n19373) );
  XOR U19644 ( .A(n19372), .B(n19373), .Z(n19374) );
  XOR U19645 ( .A(n19375), .B(n19374), .Z(n19379) );
  NANDN U19646 ( .A(n19275), .B(n19274), .Z(n19279) );
  NAND U19647 ( .A(n19277), .B(n19276), .Z(n19278) );
  NAND U19648 ( .A(n19279), .B(n19278), .Z(n19383) );
  XNOR U19649 ( .A(n19975), .B(n19576), .Z(n19330) );
  NANDN U19650 ( .A(n19330), .B(n19883), .Z(n19282) );
  NANDN U19651 ( .A(n19280), .B(n19937), .Z(n19281) );
  NAND U19652 ( .A(n19282), .B(n19281), .Z(n19342) );
  XNOR U19653 ( .A(n20052), .B(n19558), .Z(n19333) );
  OR U19654 ( .A(n19333), .B(n20020), .Z(n19285) );
  NANDN U19655 ( .A(n19283), .B(n19960), .Z(n19284) );
  NAND U19656 ( .A(n19285), .B(n19284), .Z(n19339) );
  XOR U19657 ( .A(n102), .B(a[240]), .Z(n19336) );
  OR U19658 ( .A(n19336), .B(n20121), .Z(n19288) );
  NANDN U19659 ( .A(n19286), .B(n20122), .Z(n19287) );
  AND U19660 ( .A(n19288), .B(n19287), .Z(n19340) );
  XNOR U19661 ( .A(n19339), .B(n19340), .Z(n19341) );
  XOR U19662 ( .A(n19342), .B(n19341), .Z(n19382) );
  XNOR U19663 ( .A(n19383), .B(n19382), .Z(n19385) );
  NANDN U19664 ( .A(n19290), .B(n19289), .Z(n19294) );
  NANDN U19665 ( .A(n19292), .B(n19291), .Z(n19293) );
  NAND U19666 ( .A(n19294), .B(n19293), .Z(n19384) );
  XOR U19667 ( .A(n19385), .B(n19384), .Z(n19376) );
  NANDN U19668 ( .A(n19296), .B(n19295), .Z(n19300) );
  NAND U19669 ( .A(n19298), .B(n19297), .Z(n19299) );
  AND U19670 ( .A(n19300), .B(n19299), .Z(n19377) );
  XOR U19671 ( .A(n19376), .B(n19377), .Z(n19378) );
  XOR U19672 ( .A(n19379), .B(n19378), .Z(n19324) );
  NANDN U19673 ( .A(n19302), .B(n19301), .Z(n19306) );
  NAND U19674 ( .A(n19304), .B(n19303), .Z(n19305) );
  NAND U19675 ( .A(n19306), .B(n19305), .Z(n19325) );
  XOR U19676 ( .A(n19324), .B(n19325), .Z(n19326) );
  XOR U19677 ( .A(n19327), .B(n19326), .Z(n19318) );
  NANDN U19678 ( .A(n19308), .B(n19307), .Z(n19312) );
  NANDN U19679 ( .A(n19310), .B(n19309), .Z(n19311) );
  NAND U19680 ( .A(n19312), .B(n19311), .Z(n19319) );
  XNOR U19681 ( .A(n19318), .B(n19319), .Z(n19320) );
  XNOR U19682 ( .A(n19321), .B(n19320), .Z(n19388) );
  XNOR U19683 ( .A(n19388), .B(sreg[494]), .Z(n19390) );
  NAND U19684 ( .A(n19313), .B(sreg[493]), .Z(n19317) );
  OR U19685 ( .A(n19315), .B(n19314), .Z(n19316) );
  AND U19686 ( .A(n19317), .B(n19316), .Z(n19389) );
  XOR U19687 ( .A(n19390), .B(n19389), .Z(c[494]) );
  NANDN U19688 ( .A(n19319), .B(n19318), .Z(n19323) );
  NAND U19689 ( .A(n19321), .B(n19320), .Z(n19322) );
  NAND U19690 ( .A(n19323), .B(n19322), .Z(n19396) );
  OR U19691 ( .A(n19325), .B(n19324), .Z(n19329) );
  NANDN U19692 ( .A(n19327), .B(n19326), .Z(n19328) );
  NAND U19693 ( .A(n19329), .B(n19328), .Z(n19394) );
  XNOR U19694 ( .A(n19975), .B(n19775), .Z(n19427) );
  NANDN U19695 ( .A(n19427), .B(n19883), .Z(n19332) );
  NANDN U19696 ( .A(n19330), .B(n19937), .Z(n19331) );
  NAND U19697 ( .A(n19332), .B(n19331), .Z(n19424) );
  XNOR U19698 ( .A(n20052), .B(n19647), .Z(n19430) );
  OR U19699 ( .A(n19430), .B(n20020), .Z(n19335) );
  NANDN U19700 ( .A(n19333), .B(n19960), .Z(n19334) );
  NAND U19701 ( .A(n19335), .B(n19334), .Z(n19421) );
  XOR U19702 ( .A(n102), .B(a[241]), .Z(n19434) );
  OR U19703 ( .A(n19434), .B(n20121), .Z(n19338) );
  NANDN U19704 ( .A(n19336), .B(n20122), .Z(n19337) );
  AND U19705 ( .A(n19338), .B(n19337), .Z(n19422) );
  XNOR U19706 ( .A(n19421), .B(n19422), .Z(n19423) );
  XNOR U19707 ( .A(n19424), .B(n19423), .Z(n19412) );
  NANDN U19708 ( .A(n19340), .B(n19339), .Z(n19344) );
  NAND U19709 ( .A(n19342), .B(n19341), .Z(n19343) );
  NAND U19710 ( .A(n19344), .B(n19343), .Z(n19410) );
  NANDN U19711 ( .A(n19346), .B(n19345), .Z(n19350) );
  NAND U19712 ( .A(n19348), .B(n19347), .Z(n19349) );
  AND U19713 ( .A(n19350), .B(n19349), .Z(n19409) );
  XNOR U19714 ( .A(n19410), .B(n19409), .Z(n19411) );
  XOR U19715 ( .A(n19412), .B(n19411), .Z(n19405) );
  NAND U19716 ( .A(a[255]), .B(b[0]), .Z(n19351) );
  XNOR U19717 ( .A(b[1]), .B(n19351), .Z(n19353) );
  NAND U19718 ( .A(n98), .B(a[254]), .Z(n19352) );
  AND U19719 ( .A(n19353), .B(n19352), .Z(n19445) );
  XOR U19720 ( .A(n20154), .B(a[243]), .Z(n19458) );
  OR U19721 ( .A(n19458), .B(n20057), .Z(n19356) );
  NAND U19722 ( .A(n19354), .B(n20098), .Z(n19355) );
  NAND U19723 ( .A(n19356), .B(n19355), .Z(n19443) );
  NAND U19724 ( .A(b[15]), .B(a[239]), .Z(n19444) );
  XNOR U19725 ( .A(n19443), .B(n19444), .Z(n19446) );
  XOR U19726 ( .A(n19445), .B(n19446), .Z(n19437) );
  NAND U19727 ( .A(n19554), .B(n19357), .Z(n19359) );
  XOR U19728 ( .A(a[253]), .B(b[3]), .Z(n19455) );
  NANDN U19729 ( .A(n19521), .B(n19455), .Z(n19358) );
  NAND U19730 ( .A(n19359), .B(n19358), .Z(n19417) );
  NAND U19731 ( .A(n19722), .B(n19360), .Z(n19362) );
  XOR U19732 ( .A(a[251]), .B(b[5]), .Z(n19452) );
  NANDN U19733 ( .A(n19640), .B(n19452), .Z(n19361) );
  NAND U19734 ( .A(n19362), .B(n19361), .Z(n19415) );
  XOR U19735 ( .A(b[7]), .B(a[249]), .Z(n19449) );
  NAND U19736 ( .A(n19449), .B(n19766), .Z(n19365) );
  NANDN U19737 ( .A(n19363), .B(n19767), .Z(n19364) );
  AND U19738 ( .A(n19365), .B(n19364), .Z(n19416) );
  XOR U19739 ( .A(n19417), .B(n19418), .Z(n19438) );
  XNOR U19740 ( .A(n19437), .B(n19438), .Z(n19439) );
  NANDN U19741 ( .A(n19367), .B(n19366), .Z(n19371) );
  NANDN U19742 ( .A(n19369), .B(n19368), .Z(n19370) );
  NAND U19743 ( .A(n19371), .B(n19370), .Z(n19440) );
  XOR U19744 ( .A(n19439), .B(n19440), .Z(n19403) );
  XNOR U19745 ( .A(n19403), .B(n19404), .Z(n19406) );
  XOR U19746 ( .A(n19405), .B(n19406), .Z(n19399) );
  NAND U19747 ( .A(n19377), .B(n19376), .Z(n19381) );
  NAND U19748 ( .A(n19379), .B(n19378), .Z(n19380) );
  NAND U19749 ( .A(n19381), .B(n19380), .Z(n19397) );
  OR U19750 ( .A(n19383), .B(n19382), .Z(n19387) );
  OR U19751 ( .A(n19385), .B(n19384), .Z(n19386) );
  AND U19752 ( .A(n19387), .B(n19386), .Z(n19398) );
  XNOR U19753 ( .A(n19397), .B(n19398), .Z(n19400) );
  XOR U19754 ( .A(n19399), .B(n19400), .Z(n19393) );
  XOR U19755 ( .A(n19394), .B(n19393), .Z(n19395) );
  XOR U19756 ( .A(n19396), .B(n19395), .Z(n19461) );
  XNOR U19757 ( .A(n19461), .B(sreg[495]), .Z(n19463) );
  NAND U19758 ( .A(n19388), .B(sreg[494]), .Z(n19392) );
  OR U19759 ( .A(n19390), .B(n19389), .Z(n19391) );
  AND U19760 ( .A(n19392), .B(n19391), .Z(n19462) );
  XOR U19761 ( .A(n19463), .B(n19462), .Z(c[495]) );
  NANDN U19762 ( .A(n19398), .B(n19397), .Z(n19402) );
  NAND U19763 ( .A(n19400), .B(n19399), .Z(n19401) );
  NAND U19764 ( .A(n19402), .B(n19401), .Z(n19469) );
  NANDN U19765 ( .A(n19404), .B(n19403), .Z(n19408) );
  NAND U19766 ( .A(n19406), .B(n19405), .Z(n19407) );
  NAND U19767 ( .A(n19408), .B(n19407), .Z(n19476) );
  NANDN U19768 ( .A(n19410), .B(n19409), .Z(n19414) );
  NAND U19769 ( .A(n19412), .B(n19411), .Z(n19413) );
  NAND U19770 ( .A(n19414), .B(n19413), .Z(n19475) );
  NANDN U19771 ( .A(n19416), .B(n19415), .Z(n19420) );
  NANDN U19772 ( .A(n19418), .B(n19417), .Z(n19419) );
  NAND U19773 ( .A(n19420), .B(n19419), .Z(n19489) );
  NANDN U19774 ( .A(n19422), .B(n19421), .Z(n19426) );
  NAND U19775 ( .A(n19424), .B(n19423), .Z(n19425) );
  NAND U19776 ( .A(n19426), .B(n19425), .Z(n19487) );
  XNOR U19777 ( .A(n19975), .B(n19562), .Z(n19495) );
  NANDN U19778 ( .A(n19495), .B(n19883), .Z(n19429) );
  NANDN U19779 ( .A(n19427), .B(n19937), .Z(n19428) );
  NAND U19780 ( .A(n19429), .B(n19428), .Z(n19504) );
  XNOR U19781 ( .A(n20052), .B(n19576), .Z(n19498) );
  OR U19782 ( .A(n19498), .B(n20020), .Z(n19432) );
  NANDN U19783 ( .A(n19430), .B(n19960), .Z(n19431) );
  NAND U19784 ( .A(n19432), .B(n19431), .Z(n19501) );
  XNOR U19785 ( .A(n102), .B(n19433), .Z(n19530) );
  OR U19786 ( .A(n19530), .B(n20121), .Z(n19436) );
  NANDN U19787 ( .A(n19434), .B(n20122), .Z(n19435) );
  AND U19788 ( .A(n19436), .B(n19435), .Z(n19502) );
  XNOR U19789 ( .A(n19501), .B(n19502), .Z(n19503) );
  XOR U19790 ( .A(n19504), .B(n19503), .Z(n19486) );
  XNOR U19791 ( .A(n19487), .B(n19486), .Z(n19488) );
  XNOR U19792 ( .A(n19489), .B(n19488), .Z(n19481) );
  NANDN U19793 ( .A(n19438), .B(n19437), .Z(n19442) );
  NANDN U19794 ( .A(n19440), .B(n19439), .Z(n19441) );
  AND U19795 ( .A(n19442), .B(n19441), .Z(n19480) );
  XNOR U19796 ( .A(n19481), .B(n19480), .Z(n19482) );
  NANDN U19797 ( .A(n19444), .B(n19443), .Z(n19448) );
  NAND U19798 ( .A(n19446), .B(n19445), .Z(n19447) );
  NAND U19799 ( .A(n19448), .B(n19447), .Z(n19514) );
  NAND U19800 ( .A(n19767), .B(n19449), .Z(n19451) );
  IV U19801 ( .A(a[250]), .Z(n19941) );
  XNOR U19802 ( .A(n19941), .B(n19714), .Z(n19492) );
  NANDN U19803 ( .A(n19492), .B(n19766), .Z(n19450) );
  AND U19804 ( .A(n19451), .B(n19450), .Z(n19507) );
  NAND U19805 ( .A(n19722), .B(n19452), .Z(n19454) );
  XNOR U19806 ( .A(a[252]), .B(n101), .Z(n19517) );
  NANDN U19807 ( .A(n19640), .B(n19517), .Z(n19453) );
  AND U19808 ( .A(n19454), .B(n19453), .Z(n19508) );
  XOR U19809 ( .A(n19507), .B(n19508), .Z(n19509) );
  NAND U19810 ( .A(n19554), .B(n19455), .Z(n19457) );
  XOR U19811 ( .A(a[254]), .B(b[3]), .Z(n19520) );
  NANDN U19812 ( .A(n19521), .B(n19520), .Z(n19456) );
  AND U19813 ( .A(n19457), .B(n19456), .Z(n19510) );
  XNOR U19814 ( .A(n19509), .B(n19510), .Z(n19512) );
  IV U19815 ( .A(a[255]), .Z(n20120) );
  XNOR U19816 ( .A(n20154), .B(n19558), .Z(n19533) );
  OR U19817 ( .A(n19533), .B(n20057), .Z(n19460) );
  NANDN U19818 ( .A(n19458), .B(n20098), .Z(n19459) );
  NAND U19819 ( .A(n19460), .B(n19459), .Z(n19524) );
  NAND U19820 ( .A(b[15]), .B(a[240]), .Z(n19525) );
  XNOR U19821 ( .A(n19524), .B(n19525), .Z(n19526) );
  XOR U19822 ( .A(n19527), .B(n19526), .Z(n19511) );
  XOR U19823 ( .A(n19512), .B(n19511), .Z(n19513) );
  XOR U19824 ( .A(n19514), .B(n19513), .Z(n19483) );
  XNOR U19825 ( .A(n19482), .B(n19483), .Z(n19474) );
  XNOR U19826 ( .A(n19475), .B(n19474), .Z(n19477) );
  XNOR U19827 ( .A(n19476), .B(n19477), .Z(n19468) );
  XOR U19828 ( .A(n19469), .B(n19468), .Z(n19470) );
  XOR U19829 ( .A(n19471), .B(n19470), .Z(n19467) );
  NAND U19830 ( .A(n19461), .B(sreg[495]), .Z(n19465) );
  OR U19831 ( .A(n19463), .B(n19462), .Z(n19464) );
  AND U19832 ( .A(n19465), .B(n19464), .Z(n19466) );
  XOR U19833 ( .A(n19467), .B(n19466), .Z(c[496]) );
  OR U19834 ( .A(n19467), .B(n19466), .Z(n19606) );
  NAND U19835 ( .A(n19469), .B(n19468), .Z(n19473) );
  NAND U19836 ( .A(n19471), .B(n19470), .Z(n19472) );
  NAND U19837 ( .A(n19473), .B(n19472), .Z(n19539) );
  NAND U19838 ( .A(n19475), .B(n19474), .Z(n19479) );
  NANDN U19839 ( .A(n19477), .B(n19476), .Z(n19478) );
  NAND U19840 ( .A(n19479), .B(n19478), .Z(n19537) );
  NANDN U19841 ( .A(n19481), .B(n19480), .Z(n19485) );
  NANDN U19842 ( .A(n19483), .B(n19482), .Z(n19484) );
  NAND U19843 ( .A(n19485), .B(n19484), .Z(n19598) );
  OR U19844 ( .A(n19487), .B(n19486), .Z(n19491) );
  OR U19845 ( .A(n19489), .B(n19488), .Z(n19490) );
  AND U19846 ( .A(n19491), .B(n19490), .Z(n19599) );
  XNOR U19847 ( .A(n19598), .B(n19599), .Z(n19600) );
  XOR U19848 ( .A(a[251]), .B(n19714), .Z(n19569) );
  NANDN U19849 ( .A(n19569), .B(n19766), .Z(n19494) );
  NANDN U19850 ( .A(n19492), .B(n19767), .Z(n19493) );
  NAND U19851 ( .A(n19494), .B(n19493), .Z(n19587) );
  XOR U19852 ( .A(n19975), .B(a[249]), .Z(n19566) );
  NANDN U19853 ( .A(n19566), .B(n19883), .Z(n19497) );
  NANDN U19854 ( .A(n19495), .B(n19937), .Z(n19496) );
  NAND U19855 ( .A(n19497), .B(n19496), .Z(n19584) );
  XNOR U19856 ( .A(n20052), .B(n19775), .Z(n19563) );
  OR U19857 ( .A(n19563), .B(n20020), .Z(n19500) );
  NANDN U19858 ( .A(n19498), .B(n19960), .Z(n19499) );
  AND U19859 ( .A(n19500), .B(n19499), .Z(n19585) );
  XNOR U19860 ( .A(n19584), .B(n19585), .Z(n19586) );
  XOR U19861 ( .A(n19587), .B(n19586), .Z(n19597) );
  NANDN U19862 ( .A(n19502), .B(n19501), .Z(n19506) );
  NAND U19863 ( .A(n19504), .B(n19503), .Z(n19505) );
  NAND U19864 ( .A(n19506), .B(n19505), .Z(n19595) );
  XOR U19865 ( .A(n19595), .B(n19594), .Z(n19596) );
  XOR U19866 ( .A(n19597), .B(n19596), .Z(n19592) );
  OR U19867 ( .A(n19512), .B(n19511), .Z(n19516) );
  NANDN U19868 ( .A(n19514), .B(n19513), .Z(n19515) );
  NAND U19869 ( .A(n19516), .B(n19515), .Z(n19591) );
  NAND U19870 ( .A(n19722), .B(n19517), .Z(n19519) );
  XOR U19871 ( .A(a[253]), .B(b[5]), .Z(n19572) );
  NANDN U19872 ( .A(n19640), .B(n19572), .Z(n19518) );
  NAND U19873 ( .A(n19519), .B(n19518), .Z(n19579) );
  XNOR U19874 ( .A(n99), .B(n19579), .Z(n19581) );
  NAND U19875 ( .A(n19554), .B(n19520), .Z(n19523) );
  XNOR U19876 ( .A(a[255]), .B(n100), .Z(n19553) );
  NANDN U19877 ( .A(n19521), .B(n19553), .Z(n19522) );
  NAND U19878 ( .A(n19523), .B(n19522), .Z(n19580) );
  XOR U19879 ( .A(n19581), .B(n19580), .Z(n19542) );
  NANDN U19880 ( .A(n19525), .B(n19524), .Z(n19529) );
  NAND U19881 ( .A(n19527), .B(n19526), .Z(n19528) );
  AND U19882 ( .A(n19529), .B(n19528), .Z(n19543) );
  XNOR U19883 ( .A(n19542), .B(n19543), .Z(n19545) );
  NANDN U19884 ( .A(n19530), .B(n20122), .Z(n19532) );
  XOR U19885 ( .A(b[15]), .B(a[243]), .Z(n19559) );
  NANDN U19886 ( .A(n20121), .B(n19559), .Z(n19531) );
  NAND U19887 ( .A(n19532), .B(n19531), .Z(n19550) );
  ANDN U19888 ( .B(a[241]), .A(n102), .Z(n19698) );
  IV U19889 ( .A(n19698), .Z(n19557) );
  NANDN U19890 ( .A(n19533), .B(n20098), .Z(n19535) );
  XNOR U19891 ( .A(b[13]), .B(n19647), .Z(n19575) );
  NANDN U19892 ( .A(n20057), .B(n19575), .Z(n19534) );
  NAND U19893 ( .A(n19535), .B(n19534), .Z(n19548) );
  XOR U19894 ( .A(n19557), .B(n19548), .Z(n19549) );
  XOR U19895 ( .A(n19545), .B(n19544), .Z(n19590) );
  XOR U19896 ( .A(n19591), .B(n19590), .Z(n19593) );
  XOR U19897 ( .A(n19592), .B(n19593), .Z(n19601) );
  XOR U19898 ( .A(n19600), .B(n19601), .Z(n19536) );
  XOR U19899 ( .A(n19537), .B(n19536), .Z(n19538) );
  XOR U19900 ( .A(n19539), .B(n19538), .Z(n19605) );
  XOR U19901 ( .A(n19606), .B(n19605), .Z(c[497]) );
  NAND U19902 ( .A(n19537), .B(n19536), .Z(n19541) );
  NAND U19903 ( .A(n19539), .B(n19538), .Z(n19540) );
  NAND U19904 ( .A(n19541), .B(n19540), .Z(n19613) );
  NAND U19905 ( .A(n19543), .B(n19542), .Z(n19547) );
  NANDN U19906 ( .A(n19545), .B(n19544), .Z(n19546) );
  NAND U19907 ( .A(n19547), .B(n19546), .Z(n19660) );
  NANDN U19908 ( .A(n19548), .B(n19698), .Z(n19552) );
  NANDN U19909 ( .A(n19550), .B(n19549), .Z(n19551) );
  AND U19910 ( .A(n19552), .B(n19551), .Z(n19661) );
  XNOR U19911 ( .A(n19660), .B(n19661), .Z(n19662) );
  NAND U19912 ( .A(a[242]), .B(b[15]), .Z(n19624) );
  NAND U19913 ( .A(n19554), .B(n19553), .Z(n19555) );
  NANDN U19914 ( .A(n19556), .B(n19555), .Z(n19622) );
  XOR U19915 ( .A(n19557), .B(n19622), .Z(n19623) );
  XNOR U19916 ( .A(n19624), .B(n19623), .Z(n19630) );
  XNOR U19917 ( .A(n102), .B(n19558), .Z(n19648) );
  OR U19918 ( .A(n19648), .B(n20121), .Z(n19561) );
  NAND U19919 ( .A(n19559), .B(n20122), .Z(n19560) );
  NAND U19920 ( .A(n19561), .B(n19560), .Z(n19627) );
  XNOR U19921 ( .A(n20052), .B(n19562), .Z(n19643) );
  OR U19922 ( .A(n19643), .B(n20020), .Z(n19565) );
  NANDN U19923 ( .A(n19563), .B(n19960), .Z(n19564) );
  AND U19924 ( .A(n19565), .B(n19564), .Z(n19628) );
  XNOR U19925 ( .A(n19627), .B(n19628), .Z(n19629) );
  XOR U19926 ( .A(n19630), .B(n19629), .Z(n19635) );
  XNOR U19927 ( .A(b[9]), .B(n19941), .Z(n19654) );
  NAND U19928 ( .A(n19883), .B(n19654), .Z(n19568) );
  NANDN U19929 ( .A(n19566), .B(n19937), .Z(n19567) );
  NAND U19930 ( .A(n19568), .B(n19567), .Z(n19619) );
  IV U19931 ( .A(a[252]), .Z(n20094) );
  XNOR U19932 ( .A(n20094), .B(n19714), .Z(n19657) );
  NANDN U19933 ( .A(n19657), .B(n19766), .Z(n19571) );
  NANDN U19934 ( .A(n19569), .B(n19767), .Z(n19570) );
  NAND U19935 ( .A(n19571), .B(n19570), .Z(n19616) );
  NAND U19936 ( .A(n19722), .B(n19572), .Z(n19574) );
  XOR U19937 ( .A(a[254]), .B(n101), .Z(n19639) );
  OR U19938 ( .A(n19639), .B(n19640), .Z(n19573) );
  AND U19939 ( .A(n19574), .B(n19573), .Z(n19617) );
  XNOR U19940 ( .A(n19616), .B(n19617), .Z(n19618) );
  XNOR U19941 ( .A(n19619), .B(n19618), .Z(n19633) );
  NAND U19942 ( .A(n20098), .B(n19575), .Z(n19578) );
  XNOR U19943 ( .A(b[13]), .B(n19576), .Z(n19651) );
  NANDN U19944 ( .A(n20057), .B(n19651), .Z(n19577) );
  NAND U19945 ( .A(n19578), .B(n19577), .Z(n19634) );
  XOR U19946 ( .A(n19633), .B(n19634), .Z(n19636) );
  XOR U19947 ( .A(n19635), .B(n19636), .Z(n19668) );
  NANDN U19948 ( .A(n19579), .B(b[1]), .Z(n19583) );
  OR U19949 ( .A(n19581), .B(n19580), .Z(n19582) );
  AND U19950 ( .A(n19583), .B(n19582), .Z(n19666) );
  NANDN U19951 ( .A(n19585), .B(n19584), .Z(n19589) );
  NAND U19952 ( .A(n19587), .B(n19586), .Z(n19588) );
  NAND U19953 ( .A(n19589), .B(n19588), .Z(n19667) );
  XNOR U19954 ( .A(n19666), .B(n19667), .Z(n19669) );
  XOR U19955 ( .A(n19662), .B(n19663), .Z(n19675) );
  XNOR U19956 ( .A(n19673), .B(n19672), .Z(n19674) );
  XNOR U19957 ( .A(n19675), .B(n19674), .Z(n19611) );
  IV U19958 ( .A(n19611), .Z(n19609) );
  NANDN U19959 ( .A(n19599), .B(n19598), .Z(n19603) );
  NAND U19960 ( .A(n19601), .B(n19600), .Z(n19602) );
  AND U19961 ( .A(n19603), .B(n19602), .Z(n19610) );
  XNOR U19962 ( .A(n19609), .B(n19610), .Z(n19604) );
  XNOR U19963 ( .A(n19613), .B(n19604), .Z(n19608) );
  OR U19964 ( .A(n19606), .B(n19605), .Z(n19607) );
  XOR U19965 ( .A(n19608), .B(n19607), .Z(c[498]) );
  OR U19966 ( .A(n19608), .B(n19607), .Z(n19742) );
  NAND U19967 ( .A(n19609), .B(n19610), .Z(n19615) );
  ANDN U19968 ( .B(n19611), .A(n19610), .Z(n19612) );
  OR U19969 ( .A(n19613), .B(n19612), .Z(n19614) );
  NAND U19970 ( .A(n19615), .B(n19614), .Z(n19681) );
  NANDN U19971 ( .A(n19617), .B(n19616), .Z(n19621) );
  NAND U19972 ( .A(n19619), .B(n19618), .Z(n19620) );
  NAND U19973 ( .A(n19621), .B(n19620), .Z(n19731) );
  NANDN U19974 ( .A(n19622), .B(n19698), .Z(n19626) );
  NAND U19975 ( .A(n19624), .B(n19623), .Z(n19625) );
  NAND U19976 ( .A(n19626), .B(n19625), .Z(n19728) );
  NANDN U19977 ( .A(n19628), .B(n19627), .Z(n19632) );
  NAND U19978 ( .A(n19630), .B(n19629), .Z(n19631) );
  NAND U19979 ( .A(n19632), .B(n19631), .Z(n19729) );
  XNOR U19980 ( .A(n19728), .B(n19729), .Z(n19730) );
  XOR U19981 ( .A(n19731), .B(n19730), .Z(n19684) );
  NANDN U19982 ( .A(n19634), .B(n19633), .Z(n19638) );
  OR U19983 ( .A(n19636), .B(n19635), .Z(n19637) );
  NAND U19984 ( .A(n19638), .B(n19637), .Z(n19685) );
  XNOR U19985 ( .A(n19684), .B(n19685), .Z(n19686) );
  NANDN U19986 ( .A(n19639), .B(n19722), .Z(n19642) );
  XNOR U19987 ( .A(a[255]), .B(n101), .Z(n19721) );
  NANDN U19988 ( .A(n19640), .B(n19721), .Z(n19641) );
  AND U19989 ( .A(n19642), .B(n19641), .Z(n19694) );
  XOR U19990 ( .A(n20052), .B(a[249]), .Z(n19708) );
  OR U19991 ( .A(n19708), .B(n20020), .Z(n19645) );
  NANDN U19992 ( .A(n19643), .B(n19960), .Z(n19644) );
  AND U19993 ( .A(n19645), .B(n19644), .Z(n19695) );
  XOR U19994 ( .A(n19694), .B(n19695), .Z(n19696) );
  NAND U19995 ( .A(b[15]), .B(a[243]), .Z(n19701) );
  NAND U19996 ( .A(b[1]), .B(b[2]), .Z(n19646) );
  AND U19997 ( .A(n19646), .B(b[3]), .Z(n19699) );
  XOR U19998 ( .A(n19698), .B(n19699), .Z(n19700) );
  XNOR U19999 ( .A(n19701), .B(n19700), .Z(n19697) );
  XOR U20000 ( .A(n19696), .B(n19697), .Z(n19706) );
  XNOR U20001 ( .A(n102), .B(n19647), .Z(n19725) );
  OR U20002 ( .A(n19725), .B(n20121), .Z(n19650) );
  NANDN U20003 ( .A(n19648), .B(n20122), .Z(n19649) );
  NAND U20004 ( .A(n19650), .B(n19649), .Z(n19705) );
  NAND U20005 ( .A(n20098), .B(n19651), .Z(n19653) );
  XNOR U20006 ( .A(b[13]), .B(n19775), .Z(n19718) );
  NANDN U20007 ( .A(n20057), .B(n19718), .Z(n19652) );
  AND U20008 ( .A(n19653), .B(n19652), .Z(n19692) );
  NAND U20009 ( .A(n19937), .B(n19654), .Z(n19656) );
  XOR U20010 ( .A(b[9]), .B(a[251]), .Z(n19711) );
  NAND U20011 ( .A(n19883), .B(n19711), .Z(n19655) );
  AND U20012 ( .A(n19656), .B(n19655), .Z(n19690) );
  XOR U20013 ( .A(a[253]), .B(n19714), .Z(n19715) );
  NANDN U20014 ( .A(n19715), .B(n19766), .Z(n19659) );
  NANDN U20015 ( .A(n19657), .B(n19767), .Z(n19658) );
  AND U20016 ( .A(n19659), .B(n19658), .Z(n19691) );
  XOR U20017 ( .A(n19690), .B(n19691), .Z(n19693) );
  XOR U20018 ( .A(n19692), .B(n19693), .Z(n19704) );
  XOR U20019 ( .A(n19705), .B(n19704), .Z(n19707) );
  XOR U20020 ( .A(n19706), .B(n19707), .Z(n19687) );
  XNOR U20021 ( .A(n19686), .B(n19687), .Z(n19737) );
  NANDN U20022 ( .A(n19661), .B(n19660), .Z(n19665) );
  NANDN U20023 ( .A(n19663), .B(n19662), .Z(n19664) );
  NAND U20024 ( .A(n19665), .B(n19664), .Z(n19734) );
  OR U20025 ( .A(n19667), .B(n19666), .Z(n19671) );
  NANDN U20026 ( .A(n19669), .B(n19668), .Z(n19670) );
  AND U20027 ( .A(n19671), .B(n19670), .Z(n19735) );
  XNOR U20028 ( .A(n19734), .B(n19735), .Z(n19736) );
  XNOR U20029 ( .A(n19737), .B(n19736), .Z(n19679) );
  NANDN U20030 ( .A(n19673), .B(n19672), .Z(n19677) );
  NAND U20031 ( .A(n19675), .B(n19674), .Z(n19676) );
  AND U20032 ( .A(n19677), .B(n19676), .Z(n19678) );
  XNOR U20033 ( .A(n19679), .B(n19678), .Z(n19680) );
  XNOR U20034 ( .A(n19681), .B(n19680), .Z(n19741) );
  XOR U20035 ( .A(n19742), .B(n19741), .Z(c[499]) );
  NANDN U20036 ( .A(n19679), .B(n19678), .Z(n19683) );
  NANDN U20037 ( .A(n19681), .B(n19680), .Z(n19682) );
  NAND U20038 ( .A(n19683), .B(n19682), .Z(n19747) );
  NANDN U20039 ( .A(n19685), .B(n19684), .Z(n19689) );
  NAND U20040 ( .A(n19687), .B(n19686), .Z(n19688) );
  NAND U20041 ( .A(n19689), .B(n19688), .Z(n19750) );
  NANDN U20042 ( .A(n19699), .B(n19698), .Z(n19703) );
  OR U20043 ( .A(n19701), .B(n19700), .Z(n19702) );
  NAND U20044 ( .A(n19703), .B(n19702), .Z(n19788) );
  XOR U20045 ( .A(n19789), .B(n19788), .Z(n19790) );
  XNOR U20046 ( .A(n19791), .B(n19790), .Z(n19795) );
  XNOR U20047 ( .A(n20052), .B(n19941), .Z(n19771) );
  OR U20048 ( .A(n19771), .B(n20020), .Z(n19710) );
  NANDN U20049 ( .A(n19708), .B(n19960), .Z(n19709) );
  NAND U20050 ( .A(n19710), .B(n19709), .Z(n19763) );
  XNOR U20051 ( .A(n20094), .B(n19975), .Z(n19779) );
  NANDN U20052 ( .A(n19779), .B(n19883), .Z(n19713) );
  NAND U20053 ( .A(n19711), .B(n19937), .Z(n19712) );
  NAND U20054 ( .A(n19713), .B(n19712), .Z(n19760) );
  XOR U20055 ( .A(a[254]), .B(n19714), .Z(n19768) );
  NANDN U20056 ( .A(n19768), .B(n19766), .Z(n19717) );
  NANDN U20057 ( .A(n19715), .B(n19767), .Z(n19716) );
  AND U20058 ( .A(n19717), .B(n19716), .Z(n19761) );
  XNOR U20059 ( .A(n19760), .B(n19761), .Z(n19762) );
  XNOR U20060 ( .A(n19763), .B(n19762), .Z(n19757) );
  NAND U20061 ( .A(n20098), .B(n19718), .Z(n19720) );
  XOR U20062 ( .A(b[13]), .B(a[248]), .Z(n19782) );
  NANDN U20063 ( .A(n20057), .B(n19782), .Z(n19719) );
  NAND U20064 ( .A(n19720), .B(n19719), .Z(n19754) );
  NAND U20065 ( .A(n19722), .B(n19721), .Z(n19723) );
  NANDN U20066 ( .A(n19724), .B(n19723), .Z(n19785) );
  ANDN U20067 ( .B(a[244]), .A(n102), .Z(n19810) );
  XOR U20068 ( .A(n19785), .B(n19810), .Z(n19786) );
  NANDN U20069 ( .A(n19725), .B(n20122), .Z(n19727) );
  XOR U20070 ( .A(b[15]), .B(a[246]), .Z(n19776) );
  NANDN U20071 ( .A(n20121), .B(n19776), .Z(n19726) );
  AND U20072 ( .A(n19727), .B(n19726), .Z(n19787) );
  XOR U20073 ( .A(n19786), .B(n19787), .Z(n19755) );
  XOR U20074 ( .A(n19754), .B(n19755), .Z(n19756) );
  XOR U20075 ( .A(n19757), .B(n19756), .Z(n19793) );
  XNOR U20076 ( .A(n19792), .B(n19793), .Z(n19794) );
  XNOR U20077 ( .A(n19795), .B(n19794), .Z(n19748) );
  NANDN U20078 ( .A(n19729), .B(n19728), .Z(n19733) );
  NANDN U20079 ( .A(n19731), .B(n19730), .Z(n19732) );
  AND U20080 ( .A(n19733), .B(n19732), .Z(n19749) );
  XNOR U20081 ( .A(n19748), .B(n19749), .Z(n19751) );
  XOR U20082 ( .A(n19750), .B(n19751), .Z(n19745) );
  NANDN U20083 ( .A(n19735), .B(n19734), .Z(n19739) );
  NAND U20084 ( .A(n19737), .B(n19736), .Z(n19738) );
  AND U20085 ( .A(n19739), .B(n19738), .Z(n19746) );
  XOR U20086 ( .A(n19745), .B(n19746), .Z(n19740) );
  XOR U20087 ( .A(n19747), .B(n19740), .Z(n19743) );
  OR U20088 ( .A(n19742), .B(n19741), .Z(n19744) );
  XNOR U20089 ( .A(n19743), .B(n19744), .Z(c[500]) );
  NANDN U20090 ( .A(n19744), .B(n19743), .Z(n19856) );
  NAND U20091 ( .A(n19749), .B(n19748), .Z(n19753) );
  NANDN U20092 ( .A(n19751), .B(n19750), .Z(n19752) );
  NAND U20093 ( .A(n19753), .B(n19752), .Z(n19849) );
  OR U20094 ( .A(n19755), .B(n19754), .Z(n19759) );
  NAND U20095 ( .A(n19757), .B(n19756), .Z(n19758) );
  NAND U20096 ( .A(n19759), .B(n19758), .Z(n19805) );
  NANDN U20097 ( .A(n19761), .B(n19760), .Z(n19765) );
  NAND U20098 ( .A(n19763), .B(n19762), .Z(n19764) );
  AND U20099 ( .A(n19765), .B(n19764), .Z(n19801) );
  XOR U20100 ( .A(a[255]), .B(b[7]), .Z(n19831) );
  NAND U20101 ( .A(n19831), .B(n19766), .Z(n19770) );
  NANDN U20102 ( .A(n19768), .B(n19767), .Z(n19769) );
  NAND U20103 ( .A(n19770), .B(n19769), .Z(n19837) );
  XOR U20104 ( .A(n20052), .B(a[251]), .Z(n19823) );
  OR U20105 ( .A(n19823), .B(n20020), .Z(n19773) );
  NANDN U20106 ( .A(n19771), .B(n19960), .Z(n19772) );
  AND U20107 ( .A(n19773), .B(n19772), .Z(n19838) );
  XNOR U20108 ( .A(n19837), .B(n19838), .Z(n19839) );
  NAND U20109 ( .A(b[4]), .B(b[3]), .Z(n19774) );
  NAND U20110 ( .A(b[5]), .B(n19774), .Z(n19809) );
  AND U20111 ( .A(b[15]), .B(a[245]), .Z(n19808) );
  XNOR U20112 ( .A(n19809), .B(n19808), .Z(n19811) );
  XOR U20113 ( .A(n19810), .B(n19811), .Z(n19840) );
  XOR U20114 ( .A(n19839), .B(n19840), .Z(n19798) );
  XNOR U20115 ( .A(n102), .B(n19775), .Z(n19834) );
  OR U20116 ( .A(n19834), .B(n20121), .Z(n19778) );
  NAND U20117 ( .A(n19776), .B(n20122), .Z(n19777) );
  NAND U20118 ( .A(n19778), .B(n19777), .Z(n19817) );
  XOR U20119 ( .A(a[253]), .B(n19975), .Z(n19826) );
  NANDN U20120 ( .A(n19826), .B(n19883), .Z(n19781) );
  NANDN U20121 ( .A(n19779), .B(n19937), .Z(n19780) );
  NAND U20122 ( .A(n19781), .B(n19780), .Z(n19814) );
  XOR U20123 ( .A(n20154), .B(a[249]), .Z(n19820) );
  OR U20124 ( .A(n19820), .B(n20057), .Z(n19784) );
  NAND U20125 ( .A(n19782), .B(n20098), .Z(n19783) );
  AND U20126 ( .A(n19784), .B(n19783), .Z(n19815) );
  XNOR U20127 ( .A(n19814), .B(n19815), .Z(n19816) );
  XOR U20128 ( .A(n19817), .B(n19816), .Z(n19799) );
  XOR U20129 ( .A(n19798), .B(n19799), .Z(n19800) );
  XOR U20130 ( .A(n19801), .B(n19800), .Z(n19803) );
  XOR U20131 ( .A(n19803), .B(n19802), .Z(n19804) );
  XNOR U20132 ( .A(n19805), .B(n19804), .Z(n19846) );
  NANDN U20133 ( .A(n19793), .B(n19792), .Z(n19797) );
  NANDN U20134 ( .A(n19795), .B(n19794), .Z(n19796) );
  NAND U20135 ( .A(n19797), .B(n19796), .Z(n19844) );
  XNOR U20136 ( .A(n19843), .B(n19844), .Z(n19845) );
  XOR U20137 ( .A(n19846), .B(n19845), .Z(n19850) );
  XOR U20138 ( .A(n19849), .B(n19850), .Z(n19852) );
  XOR U20139 ( .A(n19851), .B(n19852), .Z(n19855) );
  XOR U20140 ( .A(n19856), .B(n19855), .Z(c[501]) );
  OR U20141 ( .A(n19803), .B(n19802), .Z(n19807) );
  NAND U20142 ( .A(n19805), .B(n19804), .Z(n19806) );
  NAND U20143 ( .A(n19807), .B(n19806), .Z(n19902) );
  XNOR U20144 ( .A(n19901), .B(n19902), .Z(n19903) );
  NAND U20145 ( .A(n19809), .B(n19808), .Z(n19813) );
  NANDN U20146 ( .A(n19811), .B(n19810), .Z(n19812) );
  NAND U20147 ( .A(n19813), .B(n19812), .Z(n19873) );
  NANDN U20148 ( .A(n19815), .B(n19814), .Z(n19819) );
  NAND U20149 ( .A(n19817), .B(n19816), .Z(n19818) );
  NAND U20150 ( .A(n19819), .B(n19818), .Z(n19868) );
  XNOR U20151 ( .A(n20154), .B(n19941), .Z(n19887) );
  OR U20152 ( .A(n19887), .B(n20057), .Z(n19822) );
  NANDN U20153 ( .A(n19820), .B(n20098), .Z(n19821) );
  NAND U20154 ( .A(n19822), .B(n19821), .Z(n19898) );
  XNOR U20155 ( .A(n20052), .B(n20094), .Z(n19880) );
  OR U20156 ( .A(n19880), .B(n20020), .Z(n19825) );
  NANDN U20157 ( .A(n19823), .B(n19960), .Z(n19824) );
  NAND U20158 ( .A(n19825), .B(n19824), .Z(n19895) );
  XOR U20159 ( .A(a[254]), .B(n19975), .Z(n19884) );
  NANDN U20160 ( .A(n19884), .B(n19883), .Z(n19828) );
  NANDN U20161 ( .A(n19826), .B(n19937), .Z(n19827) );
  AND U20162 ( .A(n19828), .B(n19827), .Z(n19896) );
  XNOR U20163 ( .A(n19895), .B(n19896), .Z(n19897) );
  XOR U20164 ( .A(n19898), .B(n19897), .Z(n19865) );
  XNOR U20165 ( .A(b[7]), .B(n19829), .Z(n19833) );
  XNOR U20166 ( .A(b[6]), .B(b[5]), .Z(n19830) );
  NANDN U20167 ( .A(n19831), .B(n19830), .Z(n19832) );
  AND U20168 ( .A(n19833), .B(n19832), .Z(n19890) );
  ANDN U20169 ( .B(a[246]), .A(n102), .Z(n19925) );
  XNOR U20170 ( .A(n19890), .B(n19925), .Z(n19891) );
  NANDN U20171 ( .A(n19834), .B(n20122), .Z(n19836) );
  XOR U20172 ( .A(b[15]), .B(a[248]), .Z(n19877) );
  NANDN U20173 ( .A(n20121), .B(n19877), .Z(n19835) );
  AND U20174 ( .A(n19836), .B(n19835), .Z(n19892) );
  XNOR U20175 ( .A(n19891), .B(n19892), .Z(n19866) );
  XNOR U20176 ( .A(n19865), .B(n19866), .Z(n19867) );
  XNOR U20177 ( .A(n19868), .B(n19867), .Z(n19871) );
  NANDN U20178 ( .A(n19838), .B(n19837), .Z(n19842) );
  NANDN U20179 ( .A(n19840), .B(n19839), .Z(n19841) );
  AND U20180 ( .A(n19842), .B(n19841), .Z(n19872) );
  XOR U20181 ( .A(n19871), .B(n19872), .Z(n19874) );
  XNOR U20182 ( .A(n19873), .B(n19874), .Z(n19904) );
  XNOR U20183 ( .A(n19903), .B(n19904), .Z(n19860) );
  NANDN U20184 ( .A(n19844), .B(n19843), .Z(n19848) );
  NANDN U20185 ( .A(n19846), .B(n19845), .Z(n19847) );
  AND U20186 ( .A(n19848), .B(n19847), .Z(n19859) );
  XNOR U20187 ( .A(n19860), .B(n19859), .Z(n19861) );
  OR U20188 ( .A(n19850), .B(n19849), .Z(n19854) );
  NAND U20189 ( .A(n19852), .B(n19851), .Z(n19853) );
  AND U20190 ( .A(n19854), .B(n19853), .Z(n19862) );
  XNOR U20191 ( .A(n19861), .B(n19862), .Z(n19858) );
  OR U20192 ( .A(n19856), .B(n19855), .Z(n19857) );
  XOR U20193 ( .A(n19858), .B(n19857), .Z(c[502]) );
  OR U20194 ( .A(n19858), .B(n19857), .Z(n19909) );
  NANDN U20195 ( .A(n19860), .B(n19859), .Z(n19864) );
  NAND U20196 ( .A(n19862), .B(n19861), .Z(n19863) );
  AND U20197 ( .A(n19864), .B(n19863), .Z(n19912) );
  OR U20198 ( .A(n19866), .B(n19865), .Z(n19870) );
  OR U20199 ( .A(n19868), .B(n19867), .Z(n19869) );
  NAND U20200 ( .A(n19870), .B(n19869), .Z(n19951) );
  NANDN U20201 ( .A(n19872), .B(n19871), .Z(n19876) );
  NANDN U20202 ( .A(n19874), .B(n19873), .Z(n19875) );
  NAND U20203 ( .A(n19876), .B(n19875), .Z(n19952) );
  XNOR U20204 ( .A(n19951), .B(n19952), .Z(n19953) );
  XOR U20205 ( .A(n102), .B(a[249]), .Z(n19942) );
  OR U20206 ( .A(n19942), .B(n20121), .Z(n19879) );
  NAND U20207 ( .A(n19877), .B(n20122), .Z(n19878) );
  NAND U20208 ( .A(n19879), .B(n19878), .Z(n19948) );
  XOR U20209 ( .A(n20052), .B(a[253]), .Z(n19934) );
  OR U20210 ( .A(n19934), .B(n20020), .Z(n19882) );
  NANDN U20211 ( .A(n19880), .B(n19960), .Z(n19881) );
  NAND U20212 ( .A(n19882), .B(n19881), .Z(n19946) );
  XOR U20213 ( .A(n19926), .B(n19925), .Z(n19928) );
  NAND U20214 ( .A(a[247]), .B(b[15]), .Z(n19927) );
  XOR U20215 ( .A(n19928), .B(n19927), .Z(n19921) );
  XNOR U20216 ( .A(n20120), .B(n19975), .Z(n19938) );
  NANDN U20217 ( .A(n19938), .B(n19883), .Z(n19886) );
  NANDN U20218 ( .A(n19884), .B(n19937), .Z(n19885) );
  NAND U20219 ( .A(n19886), .B(n19885), .Z(n19919) );
  XOR U20220 ( .A(n20154), .B(a[251]), .Z(n19931) );
  OR U20221 ( .A(n19931), .B(n20057), .Z(n19889) );
  NANDN U20222 ( .A(n19887), .B(n20098), .Z(n19888) );
  AND U20223 ( .A(n19889), .B(n19888), .Z(n19920) );
  XNOR U20224 ( .A(n19919), .B(n19920), .Z(n19922) );
  XOR U20225 ( .A(n19921), .B(n19922), .Z(n19945) );
  XOR U20226 ( .A(n19946), .B(n19945), .Z(n19947) );
  XNOR U20227 ( .A(n19948), .B(n19947), .Z(n19916) );
  NANDN U20228 ( .A(n19890), .B(n19925), .Z(n19894) );
  NAND U20229 ( .A(n19892), .B(n19891), .Z(n19893) );
  NAND U20230 ( .A(n19894), .B(n19893), .Z(n19913) );
  NANDN U20231 ( .A(n19896), .B(n19895), .Z(n19900) );
  NAND U20232 ( .A(n19898), .B(n19897), .Z(n19899) );
  NAND U20233 ( .A(n19900), .B(n19899), .Z(n19914) );
  XNOR U20234 ( .A(n19913), .B(n19914), .Z(n19915) );
  XOR U20235 ( .A(n19916), .B(n19915), .Z(n19954) );
  XNOR U20236 ( .A(n19953), .B(n19954), .Z(n19910) );
  NANDN U20237 ( .A(n19902), .B(n19901), .Z(n19906) );
  NAND U20238 ( .A(n19904), .B(n19903), .Z(n19905) );
  AND U20239 ( .A(n19906), .B(n19905), .Z(n19911) );
  XOR U20240 ( .A(n19910), .B(n19911), .Z(n19907) );
  XNOR U20241 ( .A(n19912), .B(n19907), .Z(n19908) );
  XOR U20242 ( .A(n19909), .B(n19908), .Z(c[503]) );
  OR U20243 ( .A(n19909), .B(n19908), .Z(n19959) );
  NANDN U20244 ( .A(n19914), .B(n19913), .Z(n19918) );
  NAND U20245 ( .A(n19916), .B(n19915), .Z(n19917) );
  NAND U20246 ( .A(n19918), .B(n19917), .Z(n19992) );
  NANDN U20247 ( .A(n19920), .B(n19919), .Z(n19924) );
  NAND U20248 ( .A(n19922), .B(n19921), .Z(n19923) );
  NAND U20249 ( .A(n19924), .B(n19923), .Z(n19983) );
  NANDN U20250 ( .A(n19926), .B(n19925), .Z(n19930) );
  OR U20251 ( .A(n19928), .B(n19927), .Z(n19929) );
  NAND U20252 ( .A(n19930), .B(n19929), .Z(n19980) );
  XNOR U20253 ( .A(n20154), .B(n20094), .Z(n19969) );
  OR U20254 ( .A(n19969), .B(n20057), .Z(n19933) );
  NANDN U20255 ( .A(n19931), .B(n20098), .Z(n19932) );
  NAND U20256 ( .A(n19933), .B(n19932), .Z(n19977) );
  XOR U20257 ( .A(n20052), .B(a[254]), .Z(n19961) );
  OR U20258 ( .A(n19961), .B(n20020), .Z(n19936) );
  NANDN U20259 ( .A(n19934), .B(n19960), .Z(n19935) );
  AND U20260 ( .A(n19936), .B(n19935), .Z(n19978) );
  XNOR U20261 ( .A(n19977), .B(n19978), .Z(n19979) );
  XNOR U20262 ( .A(n19980), .B(n19979), .Z(n19984) );
  XNOR U20263 ( .A(n19983), .B(n19984), .Z(n19985) );
  NANDN U20264 ( .A(n19938), .B(n19937), .Z(n19940) );
  ANDN U20265 ( .B(n19940), .A(n19939), .Z(n19966) );
  ANDN U20266 ( .B(a[248]), .A(n102), .Z(n20016) );
  XNOR U20267 ( .A(n102), .B(n19941), .Z(n19972) );
  OR U20268 ( .A(n19972), .B(n20121), .Z(n19944) );
  NANDN U20269 ( .A(n19942), .B(n20122), .Z(n19943) );
  AND U20270 ( .A(n19944), .B(n19943), .Z(n19964) );
  XOR U20271 ( .A(n20016), .B(n19964), .Z(n19965) );
  XNOR U20272 ( .A(n19966), .B(n19965), .Z(n19986) );
  XOR U20273 ( .A(n19985), .B(n19986), .Z(n19989) );
  NAND U20274 ( .A(n19946), .B(n19945), .Z(n19950) );
  NAND U20275 ( .A(n19948), .B(n19947), .Z(n19949) );
  NAND U20276 ( .A(n19950), .B(n19949), .Z(n19990) );
  XOR U20277 ( .A(n19989), .B(n19990), .Z(n19991) );
  XNOR U20278 ( .A(n19992), .B(n19991), .Z(n19993) );
  NANDN U20279 ( .A(n19952), .B(n19951), .Z(n19956) );
  NAND U20280 ( .A(n19954), .B(n19953), .Z(n19955) );
  AND U20281 ( .A(n19956), .B(n19955), .Z(n19994) );
  XOR U20282 ( .A(n19993), .B(n19994), .Z(n19957) );
  XOR U20283 ( .A(n19995), .B(n19957), .Z(n19958) );
  XNOR U20284 ( .A(n19959), .B(n19958), .Z(c[504]) );
  NANDN U20285 ( .A(n19959), .B(n19958), .Z(n19998) );
  XOR U20286 ( .A(a[255]), .B(b[11]), .Z(n20021) );
  NANDN U20287 ( .A(n20020), .B(n20021), .Z(n19963) );
  NANDN U20288 ( .A(n19961), .B(n19960), .Z(n19962) );
  NAND U20289 ( .A(n19963), .B(n19962), .Z(n20008) );
  OR U20290 ( .A(n20016), .B(n19964), .Z(n19968) );
  NANDN U20291 ( .A(n19966), .B(n19965), .Z(n19967) );
  AND U20292 ( .A(n19968), .B(n19967), .Z(n20009) );
  XNOR U20293 ( .A(n20008), .B(n20009), .Z(n20010) );
  XOR U20294 ( .A(b[13]), .B(a[253]), .Z(n20027) );
  NANDN U20295 ( .A(n20057), .B(n20027), .Z(n19971) );
  NANDN U20296 ( .A(n19969), .B(n20098), .Z(n19970) );
  NAND U20297 ( .A(n19971), .B(n19970), .Z(n20030) );
  XOR U20298 ( .A(n102), .B(a[251]), .Z(n20024) );
  OR U20299 ( .A(n20024), .B(n20121), .Z(n19974) );
  NANDN U20300 ( .A(n19972), .B(n20122), .Z(n19973) );
  AND U20301 ( .A(n19974), .B(n19973), .Z(n20031) );
  XNOR U20302 ( .A(n20030), .B(n20031), .Z(n20032) );
  NAND U20303 ( .A(b[7]), .B(b[8]), .Z(n19976) );
  ANDN U20304 ( .B(n19976), .A(n19975), .Z(n20014) );
  NAND U20305 ( .A(b[15]), .B(a[249]), .Z(n20015) );
  XOR U20306 ( .A(n20014), .B(n20015), .Z(n20017) );
  XNOR U20307 ( .A(n20016), .B(n20017), .Z(n20033) );
  XOR U20308 ( .A(n20032), .B(n20033), .Z(n20011) );
  XOR U20309 ( .A(n20010), .B(n20011), .Z(n20002) );
  NANDN U20310 ( .A(n19978), .B(n19977), .Z(n19982) );
  NAND U20311 ( .A(n19980), .B(n19979), .Z(n19981) );
  NAND U20312 ( .A(n19982), .B(n19981), .Z(n20003) );
  XNOR U20313 ( .A(n20002), .B(n20003), .Z(n20004) );
  NANDN U20314 ( .A(n19984), .B(n19983), .Z(n19988) );
  NAND U20315 ( .A(n19986), .B(n19985), .Z(n19987) );
  AND U20316 ( .A(n19988), .B(n19987), .Z(n20005) );
  XOR U20317 ( .A(n20004), .B(n20005), .Z(n20000) );
  XNOR U20318 ( .A(n19999), .B(n20001), .Z(n19996) );
  XOR U20319 ( .A(n20000), .B(n19996), .Z(n19997) );
  XNOR U20320 ( .A(n19998), .B(n19997), .Z(c[505]) );
  NANDN U20321 ( .A(n19998), .B(n19997), .Z(n20067) );
  NANDN U20322 ( .A(n20003), .B(n20002), .Z(n20007) );
  NAND U20323 ( .A(n20005), .B(n20004), .Z(n20006) );
  NAND U20324 ( .A(n20007), .B(n20006), .Z(n20036) );
  NANDN U20325 ( .A(n20009), .B(n20008), .Z(n20013) );
  NANDN U20326 ( .A(n20011), .B(n20010), .Z(n20012) );
  NAND U20327 ( .A(n20013), .B(n20012), .Z(n20063) );
  OR U20328 ( .A(n20015), .B(n20014), .Z(n20019) );
  NAND U20329 ( .A(n20017), .B(n20016), .Z(n20018) );
  NAND U20330 ( .A(n20019), .B(n20018), .Z(n20042) );
  NAND U20331 ( .A(b[9]), .B(b[10]), .Z(n20051) );
  XNOR U20332 ( .A(b[11]), .B(n20051), .Z(n20023) );
  NANDN U20333 ( .A(n20021), .B(n20020), .Z(n20022) );
  AND U20334 ( .A(n20023), .B(n20022), .Z(n20048) );
  ANDN U20335 ( .B(a[250]), .A(n102), .Z(n20084) );
  XOR U20336 ( .A(n20048), .B(n20084), .Z(n20049) );
  NANDN U20337 ( .A(n20024), .B(n20122), .Z(n20026) );
  XNOR U20338 ( .A(n102), .B(n20094), .Z(n20053) );
  OR U20339 ( .A(n20053), .B(n20121), .Z(n20025) );
  AND U20340 ( .A(n20026), .B(n20025), .Z(n20050) );
  XOR U20341 ( .A(n20049), .B(n20050), .Z(n20043) );
  XOR U20342 ( .A(n20042), .B(n20043), .Z(n20044) );
  NAND U20343 ( .A(n20098), .B(n20027), .Z(n20029) );
  XOR U20344 ( .A(b[13]), .B(a[254]), .Z(n20056) );
  NANDN U20345 ( .A(n20057), .B(n20056), .Z(n20028) );
  NAND U20346 ( .A(n20029), .B(n20028), .Z(n20045) );
  XOR U20347 ( .A(n20044), .B(n20045), .Z(n20060) );
  NANDN U20348 ( .A(n20031), .B(n20030), .Z(n20035) );
  NANDN U20349 ( .A(n20033), .B(n20032), .Z(n20034) );
  AND U20350 ( .A(n20035), .B(n20034), .Z(n20061) );
  XNOR U20351 ( .A(n20060), .B(n20061), .Z(n20062) );
  XOR U20352 ( .A(n20063), .B(n20062), .Z(n20037) );
  XNOR U20353 ( .A(n20036), .B(n20037), .Z(n20038) );
  XNOR U20354 ( .A(n20039), .B(n20038), .Z(n20066) );
  XOR U20355 ( .A(n20067), .B(n20066), .Z(c[506]) );
  NANDN U20356 ( .A(n20037), .B(n20036), .Z(n20041) );
  NANDN U20357 ( .A(n20039), .B(n20038), .Z(n20040) );
  NAND U20358 ( .A(n20041), .B(n20040), .Z(n20072) );
  OR U20359 ( .A(n20043), .B(n20042), .Z(n20047) );
  NANDN U20360 ( .A(n20045), .B(n20044), .Z(n20046) );
  NAND U20361 ( .A(n20047), .B(n20046), .Z(n20079) );
  NANDN U20362 ( .A(n20052), .B(n20051), .Z(n20082) );
  NAND U20363 ( .A(b[15]), .B(a[251]), .Z(n20083) );
  XOR U20364 ( .A(n20082), .B(n20083), .Z(n20085) );
  XNOR U20365 ( .A(n20084), .B(n20085), .Z(n20088) );
  NANDN U20366 ( .A(n20053), .B(n20122), .Z(n20055) );
  XOR U20367 ( .A(b[15]), .B(a[253]), .Z(n20095) );
  NANDN U20368 ( .A(n20121), .B(n20095), .Z(n20054) );
  NAND U20369 ( .A(n20055), .B(n20054), .Z(n20089) );
  XOR U20370 ( .A(n20088), .B(n20089), .Z(n20090) );
  NAND U20371 ( .A(n20098), .B(n20056), .Z(n20059) );
  XNOR U20372 ( .A(b[13]), .B(n20120), .Z(n20099) );
  NANDN U20373 ( .A(n20057), .B(n20099), .Z(n20058) );
  AND U20374 ( .A(n20059), .B(n20058), .Z(n20091) );
  XNOR U20375 ( .A(n20090), .B(n20091), .Z(n20077) );
  XNOR U20376 ( .A(n20076), .B(n20077), .Z(n20078) );
  XNOR U20377 ( .A(n20079), .B(n20078), .Z(n20070) );
  NANDN U20378 ( .A(n20061), .B(n20060), .Z(n20065) );
  NAND U20379 ( .A(n20063), .B(n20062), .Z(n20064) );
  AND U20380 ( .A(n20065), .B(n20064), .Z(n20071) );
  XOR U20381 ( .A(n20070), .B(n20071), .Z(n20073) );
  XOR U20382 ( .A(n20072), .B(n20073), .Z(n20068) );
  OR U20383 ( .A(n20067), .B(n20066), .Z(n20069) );
  XNOR U20384 ( .A(n20068), .B(n20069), .Z(c[507]) );
  NANDN U20385 ( .A(n20069), .B(n20068), .Z(n20104) );
  NANDN U20386 ( .A(n20071), .B(n20070), .Z(n20075) );
  OR U20387 ( .A(n20073), .B(n20072), .Z(n20074) );
  NAND U20388 ( .A(n20075), .B(n20074), .Z(n20107) );
  NANDN U20389 ( .A(n20077), .B(n20076), .Z(n20081) );
  NAND U20390 ( .A(n20079), .B(n20078), .Z(n20080) );
  AND U20391 ( .A(n20081), .B(n20080), .Z(n20105) );
  NANDN U20392 ( .A(n20083), .B(n20082), .Z(n20087) );
  NANDN U20393 ( .A(n20085), .B(n20084), .Z(n20086) );
  NAND U20394 ( .A(n20087), .B(n20086), .Z(n20108) );
  OR U20395 ( .A(n20089), .B(n20088), .Z(n20093) );
  NAND U20396 ( .A(n20091), .B(n20090), .Z(n20092) );
  NAND U20397 ( .A(n20093), .B(n20092), .Z(n20109) );
  XNOR U20398 ( .A(n20108), .B(n20109), .Z(n20110) );
  ANDN U20399 ( .B(b[15]), .A(n20094), .Z(n20135) );
  XOR U20400 ( .A(n102), .B(a[254]), .Z(n20123) );
  OR U20401 ( .A(n20123), .B(n20121), .Z(n20097) );
  NAND U20402 ( .A(n20095), .B(n20122), .Z(n20096) );
  AND U20403 ( .A(n20097), .B(n20096), .Z(n20115) );
  XOR U20404 ( .A(n20135), .B(n20115), .Z(n20116) );
  NAND U20405 ( .A(n20099), .B(n20098), .Z(n20101) );
  ANDN U20406 ( .B(n20101), .A(n20100), .Z(n20117) );
  XNOR U20407 ( .A(n20116), .B(n20117), .Z(n20111) );
  XNOR U20408 ( .A(n20110), .B(n20111), .Z(n20106) );
  XNOR U20409 ( .A(n20105), .B(n20106), .Z(n20102) );
  XOR U20410 ( .A(n20107), .B(n20102), .Z(n20103) );
  XNOR U20411 ( .A(n20104), .B(n20103), .Z(c[508]) );
  NANDN U20412 ( .A(n20104), .B(n20103), .Z(n20150) );
  NANDN U20413 ( .A(n20109), .B(n20108), .Z(n20113) );
  NAND U20414 ( .A(n20111), .B(n20110), .Z(n20112) );
  AND U20415 ( .A(n20113), .B(n20112), .Z(n20140) );
  NAND U20416 ( .A(b[11]), .B(b[12]), .Z(n20114) );
  ANDN U20417 ( .B(n20114), .A(n20154), .Z(n20132) );
  NAND U20418 ( .A(b[15]), .B(a[253]), .Z(n20133) );
  XOR U20419 ( .A(n20132), .B(n20133), .Z(n20134) );
  XNOR U20420 ( .A(n20135), .B(n20134), .Z(n20145) );
  OR U20421 ( .A(n20115), .B(n20135), .Z(n20119) );
  NANDN U20422 ( .A(n20117), .B(n20116), .Z(n20118) );
  AND U20423 ( .A(n20119), .B(n20118), .Z(n20142) );
  XNOR U20424 ( .A(n102), .B(n20120), .Z(n20128) );
  OR U20425 ( .A(n20128), .B(n20121), .Z(n20125) );
  NANDN U20426 ( .A(n20123), .B(n20122), .Z(n20124) );
  AND U20427 ( .A(n20125), .B(n20124), .Z(n20143) );
  XOR U20428 ( .A(n20142), .B(n20143), .Z(n20144) );
  XNOR U20429 ( .A(n20140), .B(n20139), .Z(n20126) );
  XOR U20430 ( .A(n20141), .B(n20126), .Z(n20149) );
  XNOR U20431 ( .A(n20150), .B(n20149), .Z(c[509]) );
  AND U20432 ( .A(b[14]), .B(b[13]), .Z(n20127) );
  XNOR U20433 ( .A(n102), .B(n20127), .Z(n20131) );
  XNOR U20434 ( .A(b[13]), .B(b[14]), .Z(n20129) );
  NAND U20435 ( .A(n20129), .B(n20128), .Z(n20130) );
  NAND U20436 ( .A(n20131), .B(n20130), .Z(n20156) );
  OR U20437 ( .A(n20133), .B(n20132), .Z(n20137) );
  NAND U20438 ( .A(n20135), .B(n20134), .Z(n20136) );
  NAND U20439 ( .A(n20137), .B(n20136), .Z(n20157) );
  ANDN U20440 ( .B(a[254]), .A(n102), .Z(n20155) );
  XNOR U20441 ( .A(n20157), .B(n20155), .Z(n20138) );
  XOR U20442 ( .A(n20156), .B(n20138), .Z(n20151) );
  OR U20443 ( .A(n20143), .B(n20142), .Z(n20147) );
  NANDN U20444 ( .A(n20145), .B(n20144), .Z(n20146) );
  AND U20445 ( .A(n20147), .B(n20146), .Z(n20153) );
  XNOR U20446 ( .A(n20152), .B(n20153), .Z(n20148) );
  XNOR U20447 ( .A(n20151), .B(n20148), .Z(n20158) );
  NANDN U20448 ( .A(n20150), .B(n20149), .Z(n20159) );
  XNOR U20449 ( .A(n20158), .B(n20159), .Z(c[510]) );
endmodule

