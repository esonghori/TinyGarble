
module k_nns_seq_W31_K8 ( clk, rst, q, DB, min_val_out );
  input [30:0] q;
  input [30:0] DB;
  output [247:0] min_val_out;
  input clk, rst;
  wire   \min_dist_reg[7][4] , \min_dist_reg[7][3] , \min_dist_reg[7][2] ,
         \min_dist_reg[7][1] , \min_dist_reg[7][0] , \min_dist_reg[6][4] ,
         \min_dist_reg[6][3] , \min_dist_reg[6][2] , \min_dist_reg[6][1] ,
         \min_dist_reg[6][0] , \min_dist_reg[5][4] , \min_dist_reg[5][3] ,
         \min_dist_reg[5][2] , \min_dist_reg[5][1] , \min_dist_reg[5][0] ,
         \min_dist_reg[4][4] , \min_dist_reg[4][3] , \min_dist_reg[4][2] ,
         \min_dist_reg[4][1] , \min_dist_reg[4][0] , \min_dist_reg[3][4] ,
         \min_dist_reg[3][3] , \min_dist_reg[3][2] , \min_dist_reg[3][1] ,
         \min_dist_reg[3][0] , \min_dist_reg[2][4] , \min_dist_reg[2][3] ,
         \min_dist_reg[2][2] , \min_dist_reg[2][1] , \min_dist_reg[2][0] ,
         \min_dist_reg[1][4] , \min_dist_reg[1][3] , \min_dist_reg[1][2] ,
         \min_dist_reg[1][1] , \min_dist_reg[1][0] , \min_dist_reg[0][4] ,
         \min_dist_reg[0][3] , \min_dist_reg[0][2] , \min_dist_reg[0][1] ,
         \min_dist_reg[0][0] , \local_min_dist[0][4] , \local_min_dist[0][3] ,
         \local_min_dist[0][2] , \local_min_dist[0][1] ,
         \local_min_dist[0][0] , \min_dist[7][4] , \min_dist[7][3] ,
         \min_dist[7][2] , \min_dist[7][1] , \min_dist[7][0] ,
         \min_dist[6][4] , \min_dist[6][3] , \min_dist[6][2] ,
         \min_dist[6][1] , \min_dist[6][0] , \min_dist[5][4] ,
         \min_dist[5][3] , \min_dist[5][2] , \min_dist[5][1] ,
         \min_dist[5][0] , \min_dist[4][4] , \min_dist[4][3] ,
         \min_dist[4][2] , \min_dist[4][1] , \min_dist[4][0] ,
         \min_dist[3][4] , \min_dist[3][3] , \min_dist[3][2] ,
         \min_dist[3][1] , \min_dist[3][0] , \min_dist[2][4] ,
         \min_dist[2][3] , \min_dist[2][2] , \min_dist[2][1] ,
         \min_dist[2][0] , \min_dist[1][4] , \min_dist[1][3] ,
         \min_dist[1][2] , \min_dist[1][1] , \min_dist[1][0] ,
         \min_val_reg[7][30] , \min_val_reg[7][29] , \min_val_reg[7][28] ,
         \min_val_reg[7][27] , \min_val_reg[7][26] , \min_val_reg[7][25] ,
         \min_val_reg[7][24] , \min_val_reg[7][23] , \min_val_reg[7][22] ,
         \min_val_reg[7][21] , \min_val_reg[7][20] , \min_val_reg[7][19] ,
         \min_val_reg[7][18] , \min_val_reg[7][17] , \min_val_reg[7][16] ,
         \min_val_reg[7][15] , \min_val_reg[7][14] , \min_val_reg[7][13] ,
         \min_val_reg[7][12] , \min_val_reg[7][11] , \min_val_reg[7][10] ,
         \min_val_reg[7][9] , \min_val_reg[7][8] , \min_val_reg[7][7] ,
         \min_val_reg[7][6] , \min_val_reg[7][5] , \min_val_reg[7][4] ,
         \min_val_reg[7][3] , \min_val_reg[7][2] , \min_val_reg[7][1] ,
         \min_val_reg[7][0] , \min_val_reg[6][30] , \min_val_reg[6][29] ,
         \min_val_reg[6][28] , \min_val_reg[6][27] , \min_val_reg[6][26] ,
         \min_val_reg[6][25] , \min_val_reg[6][24] , \min_val_reg[6][23] ,
         \min_val_reg[6][22] , \min_val_reg[6][21] , \min_val_reg[6][20] ,
         \min_val_reg[6][19] , \min_val_reg[6][18] , \min_val_reg[6][17] ,
         \min_val_reg[6][16] , \min_val_reg[6][15] , \min_val_reg[6][14] ,
         \min_val_reg[6][13] , \min_val_reg[6][12] , \min_val_reg[6][11] ,
         \min_val_reg[6][10] , \min_val_reg[6][9] , \min_val_reg[6][8] ,
         \min_val_reg[6][7] , \min_val_reg[6][6] , \min_val_reg[6][5] ,
         \min_val_reg[6][4] , \min_val_reg[6][3] , \min_val_reg[6][2] ,
         \min_val_reg[6][1] , \min_val_reg[6][0] , \min_val_reg[5][30] ,
         \min_val_reg[5][29] , \min_val_reg[5][28] , \min_val_reg[5][27] ,
         \min_val_reg[5][26] , \min_val_reg[5][25] , \min_val_reg[5][24] ,
         \min_val_reg[5][23] , \min_val_reg[5][22] , \min_val_reg[5][21] ,
         \min_val_reg[5][20] , \min_val_reg[5][19] , \min_val_reg[5][18] ,
         \min_val_reg[5][17] , \min_val_reg[5][16] , \min_val_reg[5][15] ,
         \min_val_reg[5][14] , \min_val_reg[5][13] , \min_val_reg[5][12] ,
         \min_val_reg[5][11] , \min_val_reg[5][10] , \min_val_reg[5][9] ,
         \min_val_reg[5][8] , \min_val_reg[5][7] , \min_val_reg[5][6] ,
         \min_val_reg[5][5] , \min_val_reg[5][4] , \min_val_reg[5][3] ,
         \min_val_reg[5][2] , \min_val_reg[5][1] , \min_val_reg[5][0] ,
         \min_val_reg[4][30] , \min_val_reg[4][29] , \min_val_reg[4][28] ,
         \min_val_reg[4][27] , \min_val_reg[4][26] , \min_val_reg[4][25] ,
         \min_val_reg[4][24] , \min_val_reg[4][23] , \min_val_reg[4][22] ,
         \min_val_reg[4][21] , \min_val_reg[4][20] , \min_val_reg[4][19] ,
         \min_val_reg[4][18] , \min_val_reg[4][17] , \min_val_reg[4][16] ,
         \min_val_reg[4][15] , \min_val_reg[4][14] , \min_val_reg[4][13] ,
         \min_val_reg[4][12] , \min_val_reg[4][11] , \min_val_reg[4][10] ,
         \min_val_reg[4][9] , \min_val_reg[4][8] , \min_val_reg[4][7] ,
         \min_val_reg[4][6] , \min_val_reg[4][5] , \min_val_reg[4][4] ,
         \min_val_reg[4][3] , \min_val_reg[4][2] , \min_val_reg[4][1] ,
         \min_val_reg[4][0] , \min_val_reg[3][30] , \min_val_reg[3][29] ,
         \min_val_reg[3][28] , \min_val_reg[3][27] , \min_val_reg[3][26] ,
         \min_val_reg[3][25] , \min_val_reg[3][24] , \min_val_reg[3][23] ,
         \min_val_reg[3][22] , \min_val_reg[3][21] , \min_val_reg[3][20] ,
         \min_val_reg[3][19] , \min_val_reg[3][18] , \min_val_reg[3][17] ,
         \min_val_reg[3][16] , \min_val_reg[3][15] , \min_val_reg[3][14] ,
         \min_val_reg[3][13] , \min_val_reg[3][12] , \min_val_reg[3][11] ,
         \min_val_reg[3][10] , \min_val_reg[3][9] , \min_val_reg[3][8] ,
         \min_val_reg[3][7] , \min_val_reg[3][6] , \min_val_reg[3][5] ,
         \min_val_reg[3][4] , \min_val_reg[3][3] , \min_val_reg[3][2] ,
         \min_val_reg[3][1] , \min_val_reg[3][0] , \min_val_reg[2][30] ,
         \min_val_reg[2][29] , \min_val_reg[2][28] , \min_val_reg[2][27] ,
         \min_val_reg[2][26] , \min_val_reg[2][25] , \min_val_reg[2][24] ,
         \min_val_reg[2][23] , \min_val_reg[2][22] , \min_val_reg[2][21] ,
         \min_val_reg[2][20] , \min_val_reg[2][19] , \min_val_reg[2][18] ,
         \min_val_reg[2][17] , \min_val_reg[2][16] , \min_val_reg[2][15] ,
         \min_val_reg[2][14] , \min_val_reg[2][13] , \min_val_reg[2][12] ,
         \min_val_reg[2][11] , \min_val_reg[2][10] , \min_val_reg[2][9] ,
         \min_val_reg[2][8] , \min_val_reg[2][7] , \min_val_reg[2][6] ,
         \min_val_reg[2][5] , \min_val_reg[2][4] , \min_val_reg[2][3] ,
         \min_val_reg[2][2] , \min_val_reg[2][1] , \min_val_reg[2][0] ,
         \min_val_reg[1][30] , \min_val_reg[1][29] , \min_val_reg[1][28] ,
         \min_val_reg[1][27] , \min_val_reg[1][26] , \min_val_reg[1][25] ,
         \min_val_reg[1][24] , \min_val_reg[1][23] , \min_val_reg[1][22] ,
         \min_val_reg[1][21] , \min_val_reg[1][20] , \min_val_reg[1][19] ,
         \min_val_reg[1][18] , \min_val_reg[1][17] , \min_val_reg[1][16] ,
         \min_val_reg[1][15] , \min_val_reg[1][14] , \min_val_reg[1][13] ,
         \min_val_reg[1][12] , \min_val_reg[1][11] , \min_val_reg[1][10] ,
         \min_val_reg[1][9] , \min_val_reg[1][8] , \min_val_reg[1][7] ,
         \min_val_reg[1][6] , \min_val_reg[1][5] , \min_val_reg[1][4] ,
         \min_val_reg[1][3] , \min_val_reg[1][2] , \min_val_reg[1][1] ,
         \min_val_reg[1][0] , \min_val_reg[0][30] , \min_val_reg[0][29] ,
         \min_val_reg[0][28] , \min_val_reg[0][27] , \min_val_reg[0][26] ,
         \min_val_reg[0][25] , \min_val_reg[0][24] , \min_val_reg[0][23] ,
         \min_val_reg[0][22] , \min_val_reg[0][21] , \min_val_reg[0][20] ,
         \min_val_reg[0][19] , \min_val_reg[0][18] , \min_val_reg[0][17] ,
         \min_val_reg[0][16] , \min_val_reg[0][15] , \min_val_reg[0][14] ,
         \min_val_reg[0][13] , \min_val_reg[0][12] , \min_val_reg[0][11] ,
         \min_val_reg[0][10] , \min_val_reg[0][9] , \min_val_reg[0][8] ,
         \min_val_reg[0][7] , \min_val_reg[0][6] , \min_val_reg[0][5] ,
         \min_val_reg[0][4] , \min_val_reg[0][3] , \min_val_reg[0][2] ,
         \min_val_reg[0][1] , \min_val_reg[0][0] , n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784;

  DFF \min_dist_reg_reg[0][0]  ( .D(\local_min_dist[0][0] ), .CLK(clk), .RST(
        rst), .I(1'b1), .Q(\min_dist_reg[0][0] ) );
  DFF \min_dist_reg_reg[0][1]  ( .D(\local_min_dist[0][1] ), .CLK(clk), .RST(
        rst), .I(1'b1), .Q(\min_dist_reg[0][1] ) );
  DFF \min_dist_reg_reg[0][2]  ( .D(\local_min_dist[0][2] ), .CLK(clk), .RST(
        rst), .I(1'b1), .Q(\min_dist_reg[0][2] ) );
  DFF \min_dist_reg_reg[0][3]  ( .D(\local_min_dist[0][3] ), .CLK(clk), .RST(
        rst), .I(1'b1), .Q(\min_dist_reg[0][3] ) );
  DFF \min_dist_reg_reg[0][4]  ( .D(\local_min_dist[0][4] ), .CLK(clk), .RST(
        rst), .I(1'b1), .Q(\min_dist_reg[0][4] ) );
  DFF \min_dist_reg_reg[1][0]  ( .D(\min_dist[1][0] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][0] ) );
  DFF \min_dist_reg_reg[1][1]  ( .D(\min_dist[1][1] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][1] ) );
  DFF \min_dist_reg_reg[1][2]  ( .D(\min_dist[1][2] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][2] ) );
  DFF \min_dist_reg_reg[1][3]  ( .D(\min_dist[1][3] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][3] ) );
  DFF \min_dist_reg_reg[1][4]  ( .D(\min_dist[1][4] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][4] ) );
  DFF \min_dist_reg_reg[2][0]  ( .D(\min_dist[2][0] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][0] ) );
  DFF \min_dist_reg_reg[2][1]  ( .D(\min_dist[2][1] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][1] ) );
  DFF \min_dist_reg_reg[2][2]  ( .D(\min_dist[2][2] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][2] ) );
  DFF \min_dist_reg_reg[2][3]  ( .D(\min_dist[2][3] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][3] ) );
  DFF \min_dist_reg_reg[2][4]  ( .D(\min_dist[2][4] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][4] ) );
  DFF \min_dist_reg_reg[3][0]  ( .D(\min_dist[3][0] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][0] ) );
  DFF \min_dist_reg_reg[3][1]  ( .D(\min_dist[3][1] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][1] ) );
  DFF \min_dist_reg_reg[3][2]  ( .D(\min_dist[3][2] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][2] ) );
  DFF \min_dist_reg_reg[3][3]  ( .D(\min_dist[3][3] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][3] ) );
  DFF \min_dist_reg_reg[3][4]  ( .D(\min_dist[3][4] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][4] ) );
  DFF \min_dist_reg_reg[4][0]  ( .D(\min_dist[4][0] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[4][0] ) );
  DFF \min_dist_reg_reg[4][1]  ( .D(\min_dist[4][1] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[4][1] ) );
  DFF \min_dist_reg_reg[4][2]  ( .D(\min_dist[4][2] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[4][2] ) );
  DFF \min_dist_reg_reg[4][3]  ( .D(\min_dist[4][3] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[4][3] ) );
  DFF \min_dist_reg_reg[4][4]  ( .D(\min_dist[4][4] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[4][4] ) );
  DFF \min_dist_reg_reg[5][0]  ( .D(\min_dist[5][0] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[5][0] ) );
  DFF \min_dist_reg_reg[5][1]  ( .D(\min_dist[5][1] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[5][1] ) );
  DFF \min_dist_reg_reg[5][2]  ( .D(\min_dist[5][2] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[5][2] ) );
  DFF \min_dist_reg_reg[5][3]  ( .D(\min_dist[5][3] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[5][3] ) );
  DFF \min_dist_reg_reg[5][4]  ( .D(\min_dist[5][4] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[5][4] ) );
  DFF \min_dist_reg_reg[6][0]  ( .D(\min_dist[6][0] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[6][0] ) );
  DFF \min_dist_reg_reg[6][1]  ( .D(\min_dist[6][1] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[6][1] ) );
  DFF \min_dist_reg_reg[6][2]  ( .D(\min_dist[6][2] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[6][2] ) );
  DFF \min_dist_reg_reg[6][3]  ( .D(\min_dist[6][3] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[6][3] ) );
  DFF \min_dist_reg_reg[6][4]  ( .D(\min_dist[6][4] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[6][4] ) );
  DFF \min_dist_reg_reg[7][0]  ( .D(\min_dist[7][0] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[7][0] ) );
  DFF \min_dist_reg_reg[7][1]  ( .D(\min_dist[7][1] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[7][1] ) );
  DFF \min_dist_reg_reg[7][2]  ( .D(\min_dist[7][2] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[7][2] ) );
  DFF \min_dist_reg_reg[7][3]  ( .D(\min_dist[7][3] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[7][3] ) );
  DFF \min_dist_reg_reg[7][4]  ( .D(\min_dist[7][4] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[7][4] ) );
  DFF \min_val_reg_reg[0][0]  ( .D(min_val_out[0]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[0][0] ) );
  DFF \min_val_reg_reg[0][1]  ( .D(min_val_out[1]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[0][1] ) );
  DFF \min_val_reg_reg[0][2]  ( .D(min_val_out[2]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[0][2] ) );
  DFF \min_val_reg_reg[0][3]  ( .D(min_val_out[3]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[0][3] ) );
  DFF \min_val_reg_reg[0][4]  ( .D(min_val_out[4]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[0][4] ) );
  DFF \min_val_reg_reg[0][5]  ( .D(min_val_out[5]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[0][5] ) );
  DFF \min_val_reg_reg[0][6]  ( .D(min_val_out[6]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[0][6] ) );
  DFF \min_val_reg_reg[0][7]  ( .D(min_val_out[7]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[0][7] ) );
  DFF \min_val_reg_reg[0][8]  ( .D(min_val_out[8]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[0][8] ) );
  DFF \min_val_reg_reg[0][9]  ( .D(min_val_out[9]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[0][9] ) );
  DFF \min_val_reg_reg[0][10]  ( .D(min_val_out[10]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][10] ) );
  DFF \min_val_reg_reg[0][11]  ( .D(min_val_out[11]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][11] ) );
  DFF \min_val_reg_reg[0][12]  ( .D(min_val_out[12]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][12] ) );
  DFF \min_val_reg_reg[0][13]  ( .D(min_val_out[13]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][13] ) );
  DFF \min_val_reg_reg[0][14]  ( .D(min_val_out[14]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][14] ) );
  DFF \min_val_reg_reg[0][15]  ( .D(min_val_out[15]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][15] ) );
  DFF \min_val_reg_reg[0][16]  ( .D(min_val_out[16]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][16] ) );
  DFF \min_val_reg_reg[0][17]  ( .D(min_val_out[17]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][17] ) );
  DFF \min_val_reg_reg[0][18]  ( .D(min_val_out[18]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][18] ) );
  DFF \min_val_reg_reg[0][19]  ( .D(min_val_out[19]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][19] ) );
  DFF \min_val_reg_reg[0][20]  ( .D(min_val_out[20]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][20] ) );
  DFF \min_val_reg_reg[0][21]  ( .D(min_val_out[21]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][21] ) );
  DFF \min_val_reg_reg[0][22]  ( .D(min_val_out[22]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][22] ) );
  DFF \min_val_reg_reg[0][23]  ( .D(min_val_out[23]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][23] ) );
  DFF \min_val_reg_reg[0][24]  ( .D(min_val_out[24]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][24] ) );
  DFF \min_val_reg_reg[0][25]  ( .D(min_val_out[25]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][25] ) );
  DFF \min_val_reg_reg[0][26]  ( .D(min_val_out[26]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][26] ) );
  DFF \min_val_reg_reg[0][27]  ( .D(min_val_out[27]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][27] ) );
  DFF \min_val_reg_reg[0][28]  ( .D(min_val_out[28]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][28] ) );
  DFF \min_val_reg_reg[0][29]  ( .D(min_val_out[29]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][29] ) );
  DFF \min_val_reg_reg[0][30]  ( .D(min_val_out[30]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][30] ) );
  DFF \min_val_reg_reg[1][0]  ( .D(min_val_out[31]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[1][0] ) );
  DFF \min_val_reg_reg[1][1]  ( .D(min_val_out[32]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[1][1] ) );
  DFF \min_val_reg_reg[1][2]  ( .D(min_val_out[33]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[1][2] ) );
  DFF \min_val_reg_reg[1][3]  ( .D(min_val_out[34]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[1][3] ) );
  DFF \min_val_reg_reg[1][4]  ( .D(min_val_out[35]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[1][4] ) );
  DFF \min_val_reg_reg[1][5]  ( .D(min_val_out[36]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[1][5] ) );
  DFF \min_val_reg_reg[1][6]  ( .D(min_val_out[37]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[1][6] ) );
  DFF \min_val_reg_reg[1][7]  ( .D(min_val_out[38]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[1][7] ) );
  DFF \min_val_reg_reg[1][8]  ( .D(min_val_out[39]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[1][8] ) );
  DFF \min_val_reg_reg[1][9]  ( .D(min_val_out[40]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[1][9] ) );
  DFF \min_val_reg_reg[1][10]  ( .D(min_val_out[41]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][10] ) );
  DFF \min_val_reg_reg[1][11]  ( .D(min_val_out[42]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][11] ) );
  DFF \min_val_reg_reg[1][12]  ( .D(min_val_out[43]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][12] ) );
  DFF \min_val_reg_reg[1][13]  ( .D(min_val_out[44]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][13] ) );
  DFF \min_val_reg_reg[1][14]  ( .D(min_val_out[45]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][14] ) );
  DFF \min_val_reg_reg[1][15]  ( .D(min_val_out[46]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][15] ) );
  DFF \min_val_reg_reg[1][16]  ( .D(min_val_out[47]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][16] ) );
  DFF \min_val_reg_reg[1][17]  ( .D(min_val_out[48]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][17] ) );
  DFF \min_val_reg_reg[1][18]  ( .D(min_val_out[49]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][18] ) );
  DFF \min_val_reg_reg[1][19]  ( .D(min_val_out[50]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][19] ) );
  DFF \min_val_reg_reg[1][20]  ( .D(min_val_out[51]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][20] ) );
  DFF \min_val_reg_reg[1][21]  ( .D(min_val_out[52]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][21] ) );
  DFF \min_val_reg_reg[1][22]  ( .D(min_val_out[53]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][22] ) );
  DFF \min_val_reg_reg[1][23]  ( .D(min_val_out[54]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][23] ) );
  DFF \min_val_reg_reg[1][24]  ( .D(min_val_out[55]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][24] ) );
  DFF \min_val_reg_reg[1][25]  ( .D(min_val_out[56]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][25] ) );
  DFF \min_val_reg_reg[1][26]  ( .D(min_val_out[57]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][26] ) );
  DFF \min_val_reg_reg[1][27]  ( .D(min_val_out[58]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][27] ) );
  DFF \min_val_reg_reg[1][28]  ( .D(min_val_out[59]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][28] ) );
  DFF \min_val_reg_reg[1][29]  ( .D(min_val_out[60]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][29] ) );
  DFF \min_val_reg_reg[1][30]  ( .D(min_val_out[61]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][30] ) );
  DFF \min_val_reg_reg[2][0]  ( .D(min_val_out[62]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[2][0] ) );
  DFF \min_val_reg_reg[2][1]  ( .D(min_val_out[63]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[2][1] ) );
  DFF \min_val_reg_reg[2][2]  ( .D(min_val_out[64]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[2][2] ) );
  DFF \min_val_reg_reg[2][3]  ( .D(min_val_out[65]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[2][3] ) );
  DFF \min_val_reg_reg[2][4]  ( .D(min_val_out[66]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[2][4] ) );
  DFF \min_val_reg_reg[2][5]  ( .D(min_val_out[67]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[2][5] ) );
  DFF \min_val_reg_reg[2][6]  ( .D(min_val_out[68]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[2][6] ) );
  DFF \min_val_reg_reg[2][7]  ( .D(min_val_out[69]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[2][7] ) );
  DFF \min_val_reg_reg[2][8]  ( .D(min_val_out[70]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[2][8] ) );
  DFF \min_val_reg_reg[2][9]  ( .D(min_val_out[71]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[2][9] ) );
  DFF \min_val_reg_reg[2][10]  ( .D(min_val_out[72]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][10] ) );
  DFF \min_val_reg_reg[2][11]  ( .D(min_val_out[73]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][11] ) );
  DFF \min_val_reg_reg[2][12]  ( .D(min_val_out[74]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][12] ) );
  DFF \min_val_reg_reg[2][13]  ( .D(min_val_out[75]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][13] ) );
  DFF \min_val_reg_reg[2][14]  ( .D(min_val_out[76]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][14] ) );
  DFF \min_val_reg_reg[2][15]  ( .D(min_val_out[77]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][15] ) );
  DFF \min_val_reg_reg[2][16]  ( .D(min_val_out[78]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][16] ) );
  DFF \min_val_reg_reg[2][17]  ( .D(min_val_out[79]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][17] ) );
  DFF \min_val_reg_reg[2][18]  ( .D(min_val_out[80]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][18] ) );
  DFF \min_val_reg_reg[2][19]  ( .D(min_val_out[81]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][19] ) );
  DFF \min_val_reg_reg[2][20]  ( .D(min_val_out[82]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][20] ) );
  DFF \min_val_reg_reg[2][21]  ( .D(min_val_out[83]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][21] ) );
  DFF \min_val_reg_reg[2][22]  ( .D(min_val_out[84]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][22] ) );
  DFF \min_val_reg_reg[2][23]  ( .D(min_val_out[85]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][23] ) );
  DFF \min_val_reg_reg[2][24]  ( .D(min_val_out[86]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][24] ) );
  DFF \min_val_reg_reg[2][25]  ( .D(min_val_out[87]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][25] ) );
  DFF \min_val_reg_reg[2][26]  ( .D(min_val_out[88]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][26] ) );
  DFF \min_val_reg_reg[2][27]  ( .D(min_val_out[89]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][27] ) );
  DFF \min_val_reg_reg[2][28]  ( .D(min_val_out[90]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][28] ) );
  DFF \min_val_reg_reg[2][29]  ( .D(min_val_out[91]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][29] ) );
  DFF \min_val_reg_reg[2][30]  ( .D(min_val_out[92]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][30] ) );
  DFF \min_val_reg_reg[3][0]  ( .D(min_val_out[93]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[3][0] ) );
  DFF \min_val_reg_reg[3][1]  ( .D(min_val_out[94]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[3][1] ) );
  DFF \min_val_reg_reg[3][2]  ( .D(min_val_out[95]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[3][2] ) );
  DFF \min_val_reg_reg[3][3]  ( .D(min_val_out[96]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[3][3] ) );
  DFF \min_val_reg_reg[3][4]  ( .D(min_val_out[97]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[3][4] ) );
  DFF \min_val_reg_reg[3][5]  ( .D(min_val_out[98]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[3][5] ) );
  DFF \min_val_reg_reg[3][6]  ( .D(min_val_out[99]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[3][6] ) );
  DFF \min_val_reg_reg[3][7]  ( .D(min_val_out[100]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][7] ) );
  DFF \min_val_reg_reg[3][8]  ( .D(min_val_out[101]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][8] ) );
  DFF \min_val_reg_reg[3][9]  ( .D(min_val_out[102]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][9] ) );
  DFF \min_val_reg_reg[3][10]  ( .D(min_val_out[103]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][10] ) );
  DFF \min_val_reg_reg[3][11]  ( .D(min_val_out[104]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][11] ) );
  DFF \min_val_reg_reg[3][12]  ( .D(min_val_out[105]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][12] ) );
  DFF \min_val_reg_reg[3][13]  ( .D(min_val_out[106]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][13] ) );
  DFF \min_val_reg_reg[3][14]  ( .D(min_val_out[107]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][14] ) );
  DFF \min_val_reg_reg[3][15]  ( .D(min_val_out[108]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][15] ) );
  DFF \min_val_reg_reg[3][16]  ( .D(min_val_out[109]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][16] ) );
  DFF \min_val_reg_reg[3][17]  ( .D(min_val_out[110]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][17] ) );
  DFF \min_val_reg_reg[3][18]  ( .D(min_val_out[111]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][18] ) );
  DFF \min_val_reg_reg[3][19]  ( .D(min_val_out[112]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][19] ) );
  DFF \min_val_reg_reg[3][20]  ( .D(min_val_out[113]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][20] ) );
  DFF \min_val_reg_reg[3][21]  ( .D(min_val_out[114]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][21] ) );
  DFF \min_val_reg_reg[3][22]  ( .D(min_val_out[115]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][22] ) );
  DFF \min_val_reg_reg[3][23]  ( .D(min_val_out[116]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][23] ) );
  DFF \min_val_reg_reg[3][24]  ( .D(min_val_out[117]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][24] ) );
  DFF \min_val_reg_reg[3][25]  ( .D(min_val_out[118]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][25] ) );
  DFF \min_val_reg_reg[3][26]  ( .D(min_val_out[119]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][26] ) );
  DFF \min_val_reg_reg[3][27]  ( .D(min_val_out[120]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][27] ) );
  DFF \min_val_reg_reg[3][28]  ( .D(min_val_out[121]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][28] ) );
  DFF \min_val_reg_reg[3][29]  ( .D(min_val_out[122]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][29] ) );
  DFF \min_val_reg_reg[3][30]  ( .D(min_val_out[123]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][30] ) );
  DFF \min_val_reg_reg[4][0]  ( .D(min_val_out[124]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][0] ) );
  DFF \min_val_reg_reg[4][1]  ( .D(min_val_out[125]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][1] ) );
  DFF \min_val_reg_reg[4][2]  ( .D(min_val_out[126]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][2] ) );
  DFF \min_val_reg_reg[4][3]  ( .D(min_val_out[127]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][3] ) );
  DFF \min_val_reg_reg[4][4]  ( .D(min_val_out[128]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][4] ) );
  DFF \min_val_reg_reg[4][5]  ( .D(min_val_out[129]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][5] ) );
  DFF \min_val_reg_reg[4][6]  ( .D(min_val_out[130]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][6] ) );
  DFF \min_val_reg_reg[4][7]  ( .D(min_val_out[131]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][7] ) );
  DFF \min_val_reg_reg[4][8]  ( .D(min_val_out[132]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][8] ) );
  DFF \min_val_reg_reg[4][9]  ( .D(min_val_out[133]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][9] ) );
  DFF \min_val_reg_reg[4][10]  ( .D(min_val_out[134]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][10] ) );
  DFF \min_val_reg_reg[4][11]  ( .D(min_val_out[135]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][11] ) );
  DFF \min_val_reg_reg[4][12]  ( .D(min_val_out[136]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][12] ) );
  DFF \min_val_reg_reg[4][13]  ( .D(min_val_out[137]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][13] ) );
  DFF \min_val_reg_reg[4][14]  ( .D(min_val_out[138]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][14] ) );
  DFF \min_val_reg_reg[4][15]  ( .D(min_val_out[139]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][15] ) );
  DFF \min_val_reg_reg[4][16]  ( .D(min_val_out[140]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][16] ) );
  DFF \min_val_reg_reg[4][17]  ( .D(min_val_out[141]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][17] ) );
  DFF \min_val_reg_reg[4][18]  ( .D(min_val_out[142]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][18] ) );
  DFF \min_val_reg_reg[4][19]  ( .D(min_val_out[143]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][19] ) );
  DFF \min_val_reg_reg[4][20]  ( .D(min_val_out[144]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][20] ) );
  DFF \min_val_reg_reg[4][21]  ( .D(min_val_out[145]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][21] ) );
  DFF \min_val_reg_reg[4][22]  ( .D(min_val_out[146]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][22] ) );
  DFF \min_val_reg_reg[4][23]  ( .D(min_val_out[147]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][23] ) );
  DFF \min_val_reg_reg[4][24]  ( .D(min_val_out[148]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][24] ) );
  DFF \min_val_reg_reg[4][25]  ( .D(min_val_out[149]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][25] ) );
  DFF \min_val_reg_reg[4][26]  ( .D(min_val_out[150]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][26] ) );
  DFF \min_val_reg_reg[4][27]  ( .D(min_val_out[151]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][27] ) );
  DFF \min_val_reg_reg[4][28]  ( .D(min_val_out[152]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][28] ) );
  DFF \min_val_reg_reg[4][29]  ( .D(min_val_out[153]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][29] ) );
  DFF \min_val_reg_reg[4][30]  ( .D(min_val_out[154]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][30] ) );
  DFF \min_val_reg_reg[5][0]  ( .D(min_val_out[155]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][0] ) );
  DFF \min_val_reg_reg[5][1]  ( .D(min_val_out[156]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][1] ) );
  DFF \min_val_reg_reg[5][2]  ( .D(min_val_out[157]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][2] ) );
  DFF \min_val_reg_reg[5][3]  ( .D(min_val_out[158]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][3] ) );
  DFF \min_val_reg_reg[5][4]  ( .D(min_val_out[159]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][4] ) );
  DFF \min_val_reg_reg[5][5]  ( .D(min_val_out[160]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][5] ) );
  DFF \min_val_reg_reg[5][6]  ( .D(min_val_out[161]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][6] ) );
  DFF \min_val_reg_reg[5][7]  ( .D(min_val_out[162]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][7] ) );
  DFF \min_val_reg_reg[5][8]  ( .D(min_val_out[163]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][8] ) );
  DFF \min_val_reg_reg[5][9]  ( .D(min_val_out[164]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][9] ) );
  DFF \min_val_reg_reg[5][10]  ( .D(min_val_out[165]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][10] ) );
  DFF \min_val_reg_reg[5][11]  ( .D(min_val_out[166]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][11] ) );
  DFF \min_val_reg_reg[5][12]  ( .D(min_val_out[167]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][12] ) );
  DFF \min_val_reg_reg[5][13]  ( .D(min_val_out[168]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][13] ) );
  DFF \min_val_reg_reg[5][14]  ( .D(min_val_out[169]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][14] ) );
  DFF \min_val_reg_reg[5][15]  ( .D(min_val_out[170]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][15] ) );
  DFF \min_val_reg_reg[5][16]  ( .D(min_val_out[171]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][16] ) );
  DFF \min_val_reg_reg[5][17]  ( .D(min_val_out[172]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][17] ) );
  DFF \min_val_reg_reg[5][18]  ( .D(min_val_out[173]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][18] ) );
  DFF \min_val_reg_reg[5][19]  ( .D(min_val_out[174]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][19] ) );
  DFF \min_val_reg_reg[5][20]  ( .D(min_val_out[175]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][20] ) );
  DFF \min_val_reg_reg[5][21]  ( .D(min_val_out[176]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][21] ) );
  DFF \min_val_reg_reg[5][22]  ( .D(min_val_out[177]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][22] ) );
  DFF \min_val_reg_reg[5][23]  ( .D(min_val_out[178]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][23] ) );
  DFF \min_val_reg_reg[5][24]  ( .D(min_val_out[179]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][24] ) );
  DFF \min_val_reg_reg[5][25]  ( .D(min_val_out[180]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][25] ) );
  DFF \min_val_reg_reg[5][26]  ( .D(min_val_out[181]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][26] ) );
  DFF \min_val_reg_reg[5][27]  ( .D(min_val_out[182]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][27] ) );
  DFF \min_val_reg_reg[5][28]  ( .D(min_val_out[183]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][28] ) );
  DFF \min_val_reg_reg[5][29]  ( .D(min_val_out[184]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][29] ) );
  DFF \min_val_reg_reg[5][30]  ( .D(min_val_out[185]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][30] ) );
  DFF \min_val_reg_reg[6][0]  ( .D(min_val_out[186]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][0] ) );
  DFF \min_val_reg_reg[6][1]  ( .D(min_val_out[187]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][1] ) );
  DFF \min_val_reg_reg[6][2]  ( .D(min_val_out[188]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][2] ) );
  DFF \min_val_reg_reg[6][3]  ( .D(min_val_out[189]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][3] ) );
  DFF \min_val_reg_reg[6][4]  ( .D(min_val_out[190]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][4] ) );
  DFF \min_val_reg_reg[6][5]  ( .D(min_val_out[191]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][5] ) );
  DFF \min_val_reg_reg[6][6]  ( .D(min_val_out[192]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][6] ) );
  DFF \min_val_reg_reg[6][7]  ( .D(min_val_out[193]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][7] ) );
  DFF \min_val_reg_reg[6][8]  ( .D(min_val_out[194]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][8] ) );
  DFF \min_val_reg_reg[6][9]  ( .D(min_val_out[195]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][9] ) );
  DFF \min_val_reg_reg[6][10]  ( .D(min_val_out[196]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][10] ) );
  DFF \min_val_reg_reg[6][11]  ( .D(min_val_out[197]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][11] ) );
  DFF \min_val_reg_reg[6][12]  ( .D(min_val_out[198]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][12] ) );
  DFF \min_val_reg_reg[6][13]  ( .D(min_val_out[199]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][13] ) );
  DFF \min_val_reg_reg[6][14]  ( .D(min_val_out[200]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][14] ) );
  DFF \min_val_reg_reg[6][15]  ( .D(min_val_out[201]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][15] ) );
  DFF \min_val_reg_reg[6][16]  ( .D(min_val_out[202]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][16] ) );
  DFF \min_val_reg_reg[6][17]  ( .D(min_val_out[203]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][17] ) );
  DFF \min_val_reg_reg[6][18]  ( .D(min_val_out[204]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][18] ) );
  DFF \min_val_reg_reg[6][19]  ( .D(min_val_out[205]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][19] ) );
  DFF \min_val_reg_reg[6][20]  ( .D(min_val_out[206]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][20] ) );
  DFF \min_val_reg_reg[6][21]  ( .D(min_val_out[207]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][21] ) );
  DFF \min_val_reg_reg[6][22]  ( .D(min_val_out[208]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][22] ) );
  DFF \min_val_reg_reg[6][23]  ( .D(min_val_out[209]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][23] ) );
  DFF \min_val_reg_reg[6][24]  ( .D(min_val_out[210]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][24] ) );
  DFF \min_val_reg_reg[6][25]  ( .D(min_val_out[211]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][25] ) );
  DFF \min_val_reg_reg[6][26]  ( .D(min_val_out[212]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][26] ) );
  DFF \min_val_reg_reg[6][27]  ( .D(min_val_out[213]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][27] ) );
  DFF \min_val_reg_reg[6][28]  ( .D(min_val_out[214]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][28] ) );
  DFF \min_val_reg_reg[6][29]  ( .D(min_val_out[215]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][29] ) );
  DFF \min_val_reg_reg[6][30]  ( .D(min_val_out[216]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][30] ) );
  DFF \min_val_reg_reg[7][0]  ( .D(min_val_out[217]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][0] ) );
  DFF \min_val_reg_reg[7][1]  ( .D(min_val_out[218]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][1] ) );
  DFF \min_val_reg_reg[7][2]  ( .D(min_val_out[219]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][2] ) );
  DFF \min_val_reg_reg[7][3]  ( .D(min_val_out[220]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][3] ) );
  DFF \min_val_reg_reg[7][4]  ( .D(min_val_out[221]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][4] ) );
  DFF \min_val_reg_reg[7][5]  ( .D(min_val_out[222]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][5] ) );
  DFF \min_val_reg_reg[7][6]  ( .D(min_val_out[223]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][6] ) );
  DFF \min_val_reg_reg[7][7]  ( .D(min_val_out[224]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][7] ) );
  DFF \min_val_reg_reg[7][8]  ( .D(min_val_out[225]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][8] ) );
  DFF \min_val_reg_reg[7][9]  ( .D(min_val_out[226]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][9] ) );
  DFF \min_val_reg_reg[7][10]  ( .D(min_val_out[227]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][10] ) );
  DFF \min_val_reg_reg[7][11]  ( .D(min_val_out[228]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][11] ) );
  DFF \min_val_reg_reg[7][12]  ( .D(min_val_out[229]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][12] ) );
  DFF \min_val_reg_reg[7][13]  ( .D(min_val_out[230]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][13] ) );
  DFF \min_val_reg_reg[7][14]  ( .D(min_val_out[231]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][14] ) );
  DFF \min_val_reg_reg[7][15]  ( .D(min_val_out[232]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][15] ) );
  DFF \min_val_reg_reg[7][16]  ( .D(min_val_out[233]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][16] ) );
  DFF \min_val_reg_reg[7][17]  ( .D(min_val_out[234]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][17] ) );
  DFF \min_val_reg_reg[7][18]  ( .D(min_val_out[235]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][18] ) );
  DFF \min_val_reg_reg[7][19]  ( .D(min_val_out[236]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][19] ) );
  DFF \min_val_reg_reg[7][20]  ( .D(min_val_out[237]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][20] ) );
  DFF \min_val_reg_reg[7][21]  ( .D(min_val_out[238]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][21] ) );
  DFF \min_val_reg_reg[7][22]  ( .D(min_val_out[239]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][22] ) );
  DFF \min_val_reg_reg[7][23]  ( .D(min_val_out[240]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][23] ) );
  DFF \min_val_reg_reg[7][24]  ( .D(min_val_out[241]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][24] ) );
  DFF \min_val_reg_reg[7][25]  ( .D(min_val_out[242]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][25] ) );
  DFF \min_val_reg_reg[7][26]  ( .D(min_val_out[243]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][26] ) );
  DFF \min_val_reg_reg[7][27]  ( .D(min_val_out[244]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][27] ) );
  DFF \min_val_reg_reg[7][28]  ( .D(min_val_out[245]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][28] ) );
  DFF \min_val_reg_reg[7][29]  ( .D(min_val_out[246]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][29] ) );
  DFF \min_val_reg_reg[7][30]  ( .D(min_val_out[247]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][30] ) );
  XOR U322 ( .A(\min_val_reg[0][9] ), .B(n289), .Z(min_val_out[9]) );
  AND U323 ( .A(n290), .B(n291), .Z(n289) );
  XOR U324 ( .A(n292), .B(n293), .Z(min_val_out[99]) );
  AND U325 ( .A(n294), .B(n295), .Z(n292) );
  XOR U326 ( .A(n296), .B(n297), .Z(min_val_out[98]) );
  AND U327 ( .A(n294), .B(n298), .Z(n296) );
  XOR U328 ( .A(n299), .B(n300), .Z(min_val_out[97]) );
  AND U329 ( .A(n294), .B(n301), .Z(n299) );
  XOR U330 ( .A(n302), .B(n303), .Z(min_val_out[96]) );
  AND U331 ( .A(n294), .B(n304), .Z(n302) );
  XOR U332 ( .A(n305), .B(n306), .Z(min_val_out[95]) );
  AND U333 ( .A(n294), .B(n307), .Z(n305) );
  XOR U334 ( .A(n308), .B(n309), .Z(min_val_out[94]) );
  AND U335 ( .A(n294), .B(n310), .Z(n308) );
  XOR U336 ( .A(n311), .B(n312), .Z(min_val_out[93]) );
  AND U337 ( .A(n294), .B(n313), .Z(n311) );
  XOR U338 ( .A(n314), .B(n315), .Z(min_val_out[92]) );
  AND U339 ( .A(n316), .B(n317), .Z(n314) );
  XOR U340 ( .A(n318), .B(n319), .Z(min_val_out[91]) );
  AND U341 ( .A(n316), .B(n320), .Z(n318) );
  XOR U342 ( .A(n321), .B(n322), .Z(min_val_out[90]) );
  AND U343 ( .A(n316), .B(n323), .Z(n321) );
  XOR U344 ( .A(\min_val_reg[0][8] ), .B(n324), .Z(min_val_out[8]) );
  AND U345 ( .A(n290), .B(n325), .Z(n324) );
  XOR U346 ( .A(n326), .B(n327), .Z(min_val_out[89]) );
  AND U347 ( .A(n316), .B(n328), .Z(n326) );
  XOR U348 ( .A(n329), .B(n330), .Z(min_val_out[88]) );
  AND U349 ( .A(n316), .B(n331), .Z(n329) );
  XOR U350 ( .A(n332), .B(n333), .Z(min_val_out[87]) );
  AND U351 ( .A(n316), .B(n334), .Z(n332) );
  XOR U352 ( .A(n335), .B(n336), .Z(min_val_out[86]) );
  AND U353 ( .A(n316), .B(n337), .Z(n335) );
  XOR U354 ( .A(n338), .B(n339), .Z(min_val_out[85]) );
  AND U355 ( .A(n316), .B(n340), .Z(n338) );
  XOR U356 ( .A(n341), .B(n342), .Z(min_val_out[84]) );
  AND U357 ( .A(n316), .B(n343), .Z(n341) );
  XOR U358 ( .A(n344), .B(n345), .Z(min_val_out[83]) );
  AND U359 ( .A(n316), .B(n346), .Z(n344) );
  XOR U360 ( .A(n347), .B(n348), .Z(min_val_out[82]) );
  AND U361 ( .A(n316), .B(n349), .Z(n347) );
  XOR U362 ( .A(n350), .B(n351), .Z(min_val_out[81]) );
  AND U363 ( .A(n316), .B(n352), .Z(n350) );
  XOR U364 ( .A(n353), .B(n354), .Z(min_val_out[80]) );
  AND U365 ( .A(n316), .B(n355), .Z(n353) );
  XOR U366 ( .A(\min_val_reg[0][7] ), .B(n356), .Z(min_val_out[7]) );
  AND U367 ( .A(n290), .B(n357), .Z(n356) );
  XOR U368 ( .A(n358), .B(n359), .Z(min_val_out[79]) );
  AND U369 ( .A(n316), .B(n360), .Z(n358) );
  XOR U370 ( .A(n361), .B(n362), .Z(min_val_out[78]) );
  AND U371 ( .A(n316), .B(n363), .Z(n361) );
  XOR U372 ( .A(n364), .B(n365), .Z(min_val_out[77]) );
  AND U373 ( .A(n316), .B(n366), .Z(n364) );
  XOR U374 ( .A(n367), .B(n368), .Z(min_val_out[76]) );
  AND U375 ( .A(n316), .B(n369), .Z(n367) );
  XOR U376 ( .A(n370), .B(n371), .Z(min_val_out[75]) );
  AND U377 ( .A(n316), .B(n372), .Z(n370) );
  XOR U378 ( .A(n373), .B(n374), .Z(min_val_out[74]) );
  AND U379 ( .A(n316), .B(n375), .Z(n373) );
  XOR U380 ( .A(n376), .B(n377), .Z(min_val_out[73]) );
  AND U381 ( .A(n316), .B(n378), .Z(n376) );
  XOR U382 ( .A(n379), .B(n380), .Z(min_val_out[72]) );
  AND U383 ( .A(n316), .B(n381), .Z(n379) );
  XOR U384 ( .A(n382), .B(n383), .Z(min_val_out[71]) );
  AND U385 ( .A(n316), .B(n384), .Z(n382) );
  XOR U386 ( .A(n385), .B(n386), .Z(min_val_out[70]) );
  AND U387 ( .A(n316), .B(n387), .Z(n385) );
  XOR U388 ( .A(\min_val_reg[0][6] ), .B(n388), .Z(min_val_out[6]) );
  AND U389 ( .A(n290), .B(n389), .Z(n388) );
  XOR U390 ( .A(n390), .B(n391), .Z(min_val_out[69]) );
  AND U391 ( .A(n316), .B(n392), .Z(n390) );
  XNOR U392 ( .A(n393), .B(n394), .Z(min_val_out[68]) );
  AND U393 ( .A(n316), .B(n395), .Z(n393) );
  XNOR U394 ( .A(n396), .B(n397), .Z(min_val_out[67]) );
  AND U395 ( .A(n316), .B(n398), .Z(n396) );
  XNOR U396 ( .A(n399), .B(n400), .Z(min_val_out[66]) );
  AND U397 ( .A(n316), .B(n401), .Z(n399) );
  XNOR U398 ( .A(n402), .B(n403), .Z(min_val_out[65]) );
  AND U399 ( .A(n316), .B(n404), .Z(n402) );
  XNOR U400 ( .A(n405), .B(n406), .Z(min_val_out[64]) );
  AND U401 ( .A(n316), .B(n407), .Z(n405) );
  XNOR U402 ( .A(n408), .B(n409), .Z(min_val_out[63]) );
  AND U403 ( .A(n316), .B(n410), .Z(n408) );
  XNOR U404 ( .A(n411), .B(n412), .Z(min_val_out[62]) );
  AND U405 ( .A(n316), .B(n413), .Z(n411) );
  XNOR U406 ( .A(n414), .B(n415), .Z(min_val_out[61]) );
  AND U407 ( .A(n416), .B(n417), .Z(n414) );
  XNOR U408 ( .A(n418), .B(n419), .Z(min_val_out[60]) );
  AND U409 ( .A(n416), .B(n420), .Z(n418) );
  XOR U410 ( .A(\min_val_reg[0][5] ), .B(n421), .Z(min_val_out[5]) );
  AND U411 ( .A(n290), .B(n422), .Z(n421) );
  XNOR U412 ( .A(n423), .B(n424), .Z(min_val_out[59]) );
  AND U413 ( .A(n416), .B(n425), .Z(n423) );
  XNOR U414 ( .A(n426), .B(n427), .Z(min_val_out[58]) );
  AND U415 ( .A(n416), .B(n428), .Z(n426) );
  XNOR U416 ( .A(n429), .B(n430), .Z(min_val_out[57]) );
  AND U417 ( .A(n416), .B(n431), .Z(n429) );
  XNOR U418 ( .A(n432), .B(n433), .Z(min_val_out[56]) );
  AND U419 ( .A(n416), .B(n434), .Z(n432) );
  XNOR U420 ( .A(n435), .B(n436), .Z(min_val_out[55]) );
  AND U421 ( .A(n416), .B(n437), .Z(n435) );
  XNOR U422 ( .A(n438), .B(n439), .Z(min_val_out[54]) );
  AND U423 ( .A(n416), .B(n440), .Z(n438) );
  XNOR U424 ( .A(n441), .B(n442), .Z(min_val_out[53]) );
  AND U425 ( .A(n416), .B(n443), .Z(n441) );
  XNOR U426 ( .A(n444), .B(n445), .Z(min_val_out[52]) );
  AND U427 ( .A(n416), .B(n446), .Z(n444) );
  XNOR U428 ( .A(n447), .B(n448), .Z(min_val_out[51]) );
  AND U429 ( .A(n416), .B(n449), .Z(n447) );
  XNOR U430 ( .A(n450), .B(n451), .Z(min_val_out[50]) );
  AND U431 ( .A(n416), .B(n452), .Z(n450) );
  XOR U432 ( .A(\min_val_reg[0][4] ), .B(n453), .Z(min_val_out[4]) );
  AND U433 ( .A(n290), .B(n454), .Z(n453) );
  XNOR U434 ( .A(n455), .B(n456), .Z(min_val_out[49]) );
  AND U435 ( .A(n416), .B(n457), .Z(n455) );
  XNOR U436 ( .A(n458), .B(n459), .Z(min_val_out[48]) );
  AND U437 ( .A(n416), .B(n460), .Z(n458) );
  XNOR U438 ( .A(n461), .B(n462), .Z(min_val_out[47]) );
  AND U439 ( .A(n416), .B(n463), .Z(n461) );
  XNOR U440 ( .A(n464), .B(n465), .Z(min_val_out[46]) );
  AND U441 ( .A(n416), .B(n466), .Z(n464) );
  XNOR U442 ( .A(n467), .B(n468), .Z(min_val_out[45]) );
  AND U443 ( .A(n416), .B(n469), .Z(n467) );
  XNOR U444 ( .A(n470), .B(n471), .Z(min_val_out[44]) );
  AND U445 ( .A(n416), .B(n472), .Z(n470) );
  XNOR U446 ( .A(n473), .B(n474), .Z(min_val_out[43]) );
  AND U447 ( .A(n416), .B(n475), .Z(n473) );
  XNOR U448 ( .A(n476), .B(n477), .Z(min_val_out[42]) );
  AND U449 ( .A(n416), .B(n478), .Z(n476) );
  XNOR U450 ( .A(n479), .B(n480), .Z(min_val_out[41]) );
  AND U451 ( .A(n416), .B(n481), .Z(n479) );
  XOR U452 ( .A(n482), .B(n483), .Z(min_val_out[40]) );
  AND U453 ( .A(n416), .B(n291), .Z(n482) );
  XOR U454 ( .A(\min_val_reg[0][9] ), .B(n483), .Z(n291) );
  XNOR U455 ( .A(\min_val_reg[1][9] ), .B(n484), .Z(n483) );
  NAND U456 ( .A(n384), .B(n316), .Z(n484) );
  XOR U457 ( .A(\min_val_reg[1][9] ), .B(n383), .Z(n384) );
  XNOR U458 ( .A(\min_val_reg[2][9] ), .B(n485), .Z(n383) );
  NAND U459 ( .A(n486), .B(n294), .Z(n485) );
  XOR U460 ( .A(\min_val_reg[0][3] ), .B(n487), .Z(min_val_out[3]) );
  AND U461 ( .A(n290), .B(n488), .Z(n487) );
  XOR U462 ( .A(n489), .B(n490), .Z(min_val_out[39]) );
  AND U463 ( .A(n416), .B(n325), .Z(n489) );
  XOR U464 ( .A(\min_val_reg[0][8] ), .B(n490), .Z(n325) );
  XNOR U465 ( .A(\min_val_reg[1][8] ), .B(n491), .Z(n490) );
  NAND U466 ( .A(n387), .B(n316), .Z(n491) );
  XOR U467 ( .A(\min_val_reg[1][8] ), .B(n386), .Z(n387) );
  XNOR U468 ( .A(\min_val_reg[2][8] ), .B(n492), .Z(n386) );
  NAND U469 ( .A(n493), .B(n294), .Z(n492) );
  XOR U470 ( .A(n494), .B(n495), .Z(min_val_out[38]) );
  AND U471 ( .A(n416), .B(n357), .Z(n494) );
  XOR U472 ( .A(\min_val_reg[0][7] ), .B(n495), .Z(n357) );
  XNOR U473 ( .A(\min_val_reg[1][7] ), .B(n496), .Z(n495) );
  NAND U474 ( .A(n392), .B(n316), .Z(n496) );
  XOR U475 ( .A(\min_val_reg[1][7] ), .B(n391), .Z(n392) );
  XNOR U476 ( .A(\min_val_reg[2][7] ), .B(n497), .Z(n391) );
  NAND U477 ( .A(n498), .B(n294), .Z(n497) );
  XOR U478 ( .A(n499), .B(n500), .Z(min_val_out[37]) );
  AND U479 ( .A(n416), .B(n389), .Z(n499) );
  XOR U480 ( .A(\min_val_reg[0][6] ), .B(n500), .Z(n389) );
  XNOR U481 ( .A(\min_val_reg[1][6] ), .B(n501), .Z(n500) );
  NAND U482 ( .A(n395), .B(n316), .Z(n501) );
  XNOR U483 ( .A(\min_val_reg[1][6] ), .B(n394), .Z(n395) );
  XOR U484 ( .A(\min_val_reg[2][6] ), .B(n502), .Z(n394) );
  NAND U485 ( .A(n295), .B(n294), .Z(n502) );
  XOR U486 ( .A(\min_val_reg[2][6] ), .B(n293), .Z(n295) );
  XNOR U487 ( .A(\min_val_reg[3][6] ), .B(n503), .Z(n293) );
  NAND U488 ( .A(n504), .B(n505), .Z(n503) );
  XNOR U489 ( .A(n506), .B(n507), .Z(min_val_out[36]) );
  AND U490 ( .A(n416), .B(n422), .Z(n506) );
  XNOR U491 ( .A(\min_val_reg[0][5] ), .B(n507), .Z(n422) );
  XOR U492 ( .A(\min_val_reg[1][5] ), .B(n508), .Z(n507) );
  NAND U493 ( .A(n398), .B(n316), .Z(n508) );
  XNOR U494 ( .A(\min_val_reg[1][5] ), .B(n397), .Z(n398) );
  XOR U495 ( .A(\min_val_reg[2][5] ), .B(n509), .Z(n397) );
  NAND U496 ( .A(n298), .B(n294), .Z(n509) );
  XOR U497 ( .A(\min_val_reg[2][5] ), .B(n297), .Z(n298) );
  XNOR U498 ( .A(\min_val_reg[3][5] ), .B(n510), .Z(n297) );
  NAND U499 ( .A(n511), .B(n505), .Z(n510) );
  XNOR U500 ( .A(n512), .B(n513), .Z(min_val_out[35]) );
  AND U501 ( .A(n416), .B(n454), .Z(n512) );
  XNOR U502 ( .A(\min_val_reg[0][4] ), .B(n513), .Z(n454) );
  XOR U503 ( .A(\min_val_reg[1][4] ), .B(n514), .Z(n513) );
  NAND U504 ( .A(n401), .B(n316), .Z(n514) );
  XNOR U505 ( .A(\min_val_reg[1][4] ), .B(n400), .Z(n401) );
  XOR U506 ( .A(\min_val_reg[2][4] ), .B(n515), .Z(n400) );
  NAND U507 ( .A(n301), .B(n294), .Z(n515) );
  XOR U508 ( .A(\min_val_reg[2][4] ), .B(n300), .Z(n301) );
  XNOR U509 ( .A(\min_val_reg[3][4] ), .B(n516), .Z(n300) );
  NAND U510 ( .A(n517), .B(n505), .Z(n516) );
  XNOR U511 ( .A(n518), .B(n519), .Z(min_val_out[34]) );
  AND U512 ( .A(n416), .B(n488), .Z(n518) );
  XNOR U513 ( .A(\min_val_reg[0][3] ), .B(n519), .Z(n488) );
  XOR U514 ( .A(\min_val_reg[1][3] ), .B(n520), .Z(n519) );
  NAND U515 ( .A(n404), .B(n316), .Z(n520) );
  XNOR U516 ( .A(\min_val_reg[1][3] ), .B(n403), .Z(n404) );
  XOR U517 ( .A(\min_val_reg[2][3] ), .B(n521), .Z(n403) );
  NAND U518 ( .A(n304), .B(n294), .Z(n521) );
  XOR U519 ( .A(\min_val_reg[2][3] ), .B(n303), .Z(n304) );
  XNOR U520 ( .A(\min_val_reg[3][3] ), .B(n522), .Z(n303) );
  NAND U521 ( .A(n523), .B(n505), .Z(n522) );
  XNOR U522 ( .A(n524), .B(n525), .Z(min_val_out[33]) );
  AND U523 ( .A(n416), .B(n526), .Z(n524) );
  XNOR U524 ( .A(n527), .B(n528), .Z(min_val_out[32]) );
  AND U525 ( .A(n416), .B(n529), .Z(n527) );
  XNOR U526 ( .A(n530), .B(n531), .Z(min_val_out[31]) );
  AND U527 ( .A(n416), .B(n532), .Z(n530) );
  XOR U528 ( .A(\min_val_reg[0][30] ), .B(n533), .Z(min_val_out[30]) );
  AND U529 ( .A(n290), .B(n417), .Z(n533) );
  XNOR U530 ( .A(\min_val_reg[0][30] ), .B(n415), .Z(n417) );
  XOR U531 ( .A(\min_val_reg[1][30] ), .B(n534), .Z(n415) );
  NAND U532 ( .A(n317), .B(n316), .Z(n534) );
  XOR U533 ( .A(\min_val_reg[1][30] ), .B(n315), .Z(n317) );
  XNOR U534 ( .A(\min_val_reg[2][30] ), .B(n535), .Z(n315) );
  NAND U535 ( .A(n536), .B(n294), .Z(n535) );
  XOR U536 ( .A(\min_val_reg[0][2] ), .B(n537), .Z(min_val_out[2]) );
  AND U537 ( .A(n290), .B(n526), .Z(n537) );
  XNOR U538 ( .A(\min_val_reg[0][2] ), .B(n525), .Z(n526) );
  XOR U539 ( .A(\min_val_reg[1][2] ), .B(n538), .Z(n525) );
  NAND U540 ( .A(n407), .B(n316), .Z(n538) );
  XNOR U541 ( .A(\min_val_reg[1][2] ), .B(n406), .Z(n407) );
  XOR U542 ( .A(\min_val_reg[2][2] ), .B(n539), .Z(n406) );
  NAND U543 ( .A(n307), .B(n294), .Z(n539) );
  XOR U544 ( .A(\min_val_reg[2][2] ), .B(n306), .Z(n307) );
  XNOR U545 ( .A(\min_val_reg[3][2] ), .B(n540), .Z(n306) );
  NAND U546 ( .A(n541), .B(n505), .Z(n540) );
  XOR U547 ( .A(\min_val_reg[0][29] ), .B(n542), .Z(min_val_out[29]) );
  AND U548 ( .A(n290), .B(n420), .Z(n542) );
  XNOR U549 ( .A(\min_val_reg[0][29] ), .B(n419), .Z(n420) );
  XOR U550 ( .A(\min_val_reg[1][29] ), .B(n543), .Z(n419) );
  NAND U551 ( .A(n320), .B(n316), .Z(n543) );
  XOR U552 ( .A(\min_val_reg[1][29] ), .B(n319), .Z(n320) );
  XNOR U553 ( .A(\min_val_reg[2][29] ), .B(n544), .Z(n319) );
  NAND U554 ( .A(n545), .B(n294), .Z(n544) );
  XOR U555 ( .A(\min_val_reg[0][28] ), .B(n546), .Z(min_val_out[28]) );
  AND U556 ( .A(n290), .B(n425), .Z(n546) );
  XNOR U557 ( .A(\min_val_reg[0][28] ), .B(n424), .Z(n425) );
  XOR U558 ( .A(\min_val_reg[1][28] ), .B(n547), .Z(n424) );
  NAND U559 ( .A(n323), .B(n316), .Z(n547) );
  XOR U560 ( .A(\min_val_reg[1][28] ), .B(n322), .Z(n323) );
  XNOR U561 ( .A(\min_val_reg[2][28] ), .B(n548), .Z(n322) );
  NAND U562 ( .A(n549), .B(n294), .Z(n548) );
  XOR U563 ( .A(\min_val_reg[0][27] ), .B(n550), .Z(min_val_out[27]) );
  AND U564 ( .A(n290), .B(n428), .Z(n550) );
  XNOR U565 ( .A(\min_val_reg[0][27] ), .B(n427), .Z(n428) );
  XOR U566 ( .A(\min_val_reg[1][27] ), .B(n551), .Z(n427) );
  NAND U567 ( .A(n328), .B(n316), .Z(n551) );
  XOR U568 ( .A(\min_val_reg[1][27] ), .B(n327), .Z(n328) );
  XNOR U569 ( .A(\min_val_reg[2][27] ), .B(n552), .Z(n327) );
  NAND U570 ( .A(n553), .B(n294), .Z(n552) );
  XOR U571 ( .A(\min_val_reg[0][26] ), .B(n554), .Z(min_val_out[26]) );
  AND U572 ( .A(n290), .B(n431), .Z(n554) );
  XNOR U573 ( .A(\min_val_reg[0][26] ), .B(n430), .Z(n431) );
  XOR U574 ( .A(\min_val_reg[1][26] ), .B(n555), .Z(n430) );
  NAND U575 ( .A(n331), .B(n316), .Z(n555) );
  XOR U576 ( .A(\min_val_reg[1][26] ), .B(n330), .Z(n331) );
  XNOR U577 ( .A(\min_val_reg[2][26] ), .B(n556), .Z(n330) );
  NAND U578 ( .A(n557), .B(n294), .Z(n556) );
  XOR U579 ( .A(\min_val_reg[0][25] ), .B(n558), .Z(min_val_out[25]) );
  AND U580 ( .A(n290), .B(n434), .Z(n558) );
  XNOR U581 ( .A(\min_val_reg[0][25] ), .B(n433), .Z(n434) );
  XOR U582 ( .A(\min_val_reg[1][25] ), .B(n559), .Z(n433) );
  NAND U583 ( .A(n334), .B(n316), .Z(n559) );
  XOR U584 ( .A(\min_val_reg[1][25] ), .B(n333), .Z(n334) );
  XNOR U585 ( .A(\min_val_reg[2][25] ), .B(n560), .Z(n333) );
  NAND U586 ( .A(n561), .B(n294), .Z(n560) );
  XOR U587 ( .A(\min_val_reg[0][24] ), .B(n562), .Z(min_val_out[24]) );
  AND U588 ( .A(n290), .B(n437), .Z(n562) );
  XNOR U589 ( .A(\min_val_reg[0][24] ), .B(n436), .Z(n437) );
  XOR U590 ( .A(\min_val_reg[1][24] ), .B(n563), .Z(n436) );
  NAND U591 ( .A(n337), .B(n316), .Z(n563) );
  XOR U592 ( .A(\min_val_reg[1][24] ), .B(n336), .Z(n337) );
  XNOR U593 ( .A(\min_val_reg[2][24] ), .B(n564), .Z(n336) );
  NAND U594 ( .A(n565), .B(n294), .Z(n564) );
  XNOR U595 ( .A(n566), .B(n567), .Z(min_val_out[247]) );
  AND U596 ( .A(n568), .B(n569), .Z(n566) );
  XNOR U597 ( .A(n570), .B(n571), .Z(min_val_out[246]) );
  AND U598 ( .A(n568), .B(n572), .Z(n570) );
  XNOR U599 ( .A(n573), .B(n574), .Z(min_val_out[245]) );
  AND U600 ( .A(n568), .B(n575), .Z(n573) );
  XNOR U601 ( .A(n576), .B(n577), .Z(min_val_out[244]) );
  AND U602 ( .A(n568), .B(n578), .Z(n576) );
  XNOR U603 ( .A(n579), .B(n580), .Z(min_val_out[243]) );
  AND U604 ( .A(n568), .B(n581), .Z(n579) );
  XNOR U605 ( .A(n582), .B(n583), .Z(min_val_out[242]) );
  AND U606 ( .A(n568), .B(n584), .Z(n582) );
  XNOR U607 ( .A(n585), .B(n586), .Z(min_val_out[241]) );
  AND U608 ( .A(n568), .B(n587), .Z(n585) );
  XNOR U609 ( .A(n588), .B(n589), .Z(min_val_out[240]) );
  AND U610 ( .A(n568), .B(n590), .Z(n588) );
  XOR U611 ( .A(\min_val_reg[0][23] ), .B(n591), .Z(min_val_out[23]) );
  AND U612 ( .A(n290), .B(n440), .Z(n591) );
  XNOR U613 ( .A(\min_val_reg[0][23] ), .B(n439), .Z(n440) );
  XOR U614 ( .A(\min_val_reg[1][23] ), .B(n592), .Z(n439) );
  NAND U615 ( .A(n340), .B(n316), .Z(n592) );
  XOR U616 ( .A(\min_val_reg[1][23] ), .B(n339), .Z(n340) );
  XNOR U617 ( .A(\min_val_reg[2][23] ), .B(n593), .Z(n339) );
  NAND U618 ( .A(n594), .B(n294), .Z(n593) );
  XNOR U619 ( .A(n595), .B(n596), .Z(min_val_out[239]) );
  AND U620 ( .A(n568), .B(n597), .Z(n595) );
  XNOR U621 ( .A(n598), .B(n599), .Z(min_val_out[238]) );
  AND U622 ( .A(n568), .B(n600), .Z(n598) );
  XNOR U623 ( .A(n601), .B(n602), .Z(min_val_out[237]) );
  AND U624 ( .A(n568), .B(n603), .Z(n601) );
  XNOR U625 ( .A(n604), .B(n605), .Z(min_val_out[236]) );
  AND U626 ( .A(n568), .B(n606), .Z(n604) );
  XNOR U627 ( .A(n607), .B(n608), .Z(min_val_out[235]) );
  AND U628 ( .A(n568), .B(n609), .Z(n607) );
  XNOR U629 ( .A(n610), .B(n611), .Z(min_val_out[234]) );
  AND U630 ( .A(n568), .B(n612), .Z(n610) );
  XNOR U631 ( .A(n613), .B(n614), .Z(min_val_out[233]) );
  AND U632 ( .A(n568), .B(n615), .Z(n613) );
  XNOR U633 ( .A(n616), .B(n617), .Z(min_val_out[232]) );
  AND U634 ( .A(n568), .B(n618), .Z(n616) );
  XNOR U635 ( .A(n619), .B(n620), .Z(min_val_out[231]) );
  AND U636 ( .A(n568), .B(n621), .Z(n619) );
  XNOR U637 ( .A(n622), .B(n623), .Z(min_val_out[230]) );
  AND U638 ( .A(n568), .B(n624), .Z(n622) );
  XOR U639 ( .A(\min_val_reg[0][22] ), .B(n625), .Z(min_val_out[22]) );
  AND U640 ( .A(n290), .B(n443), .Z(n625) );
  XNOR U641 ( .A(\min_val_reg[0][22] ), .B(n442), .Z(n443) );
  XOR U642 ( .A(\min_val_reg[1][22] ), .B(n626), .Z(n442) );
  NAND U643 ( .A(n343), .B(n316), .Z(n626) );
  XOR U644 ( .A(\min_val_reg[1][22] ), .B(n342), .Z(n343) );
  XNOR U645 ( .A(\min_val_reg[2][22] ), .B(n627), .Z(n342) );
  NAND U646 ( .A(n628), .B(n294), .Z(n627) );
  XNOR U647 ( .A(n629), .B(n630), .Z(min_val_out[229]) );
  AND U648 ( .A(n568), .B(n631), .Z(n629) );
  XNOR U649 ( .A(n632), .B(n633), .Z(min_val_out[228]) );
  AND U650 ( .A(n568), .B(n634), .Z(n632) );
  XNOR U651 ( .A(n635), .B(n636), .Z(min_val_out[227]) );
  AND U652 ( .A(n568), .B(n637), .Z(n635) );
  XNOR U653 ( .A(n638), .B(n639), .Z(min_val_out[226]) );
  AND U654 ( .A(n568), .B(n640), .Z(n638) );
  XNOR U655 ( .A(n641), .B(n642), .Z(min_val_out[225]) );
  AND U656 ( .A(n568), .B(n643), .Z(n641) );
  XNOR U657 ( .A(n644), .B(n645), .Z(min_val_out[224]) );
  AND U658 ( .A(n568), .B(n646), .Z(n644) );
  XNOR U659 ( .A(n647), .B(n648), .Z(min_val_out[223]) );
  AND U660 ( .A(n568), .B(n649), .Z(n647) );
  XNOR U661 ( .A(n650), .B(n651), .Z(min_val_out[222]) );
  AND U662 ( .A(n568), .B(n652), .Z(n650) );
  XNOR U663 ( .A(n653), .B(n654), .Z(min_val_out[221]) );
  AND U664 ( .A(n568), .B(n655), .Z(n653) );
  XNOR U665 ( .A(n656), .B(n657), .Z(min_val_out[220]) );
  AND U666 ( .A(n568), .B(n658), .Z(n656) );
  XOR U667 ( .A(\min_val_reg[0][21] ), .B(n659), .Z(min_val_out[21]) );
  AND U668 ( .A(n290), .B(n446), .Z(n659) );
  XNOR U669 ( .A(\min_val_reg[0][21] ), .B(n445), .Z(n446) );
  XOR U670 ( .A(\min_val_reg[1][21] ), .B(n660), .Z(n445) );
  NAND U671 ( .A(n346), .B(n316), .Z(n660) );
  XOR U672 ( .A(\min_val_reg[1][21] ), .B(n345), .Z(n346) );
  XNOR U673 ( .A(\min_val_reg[2][21] ), .B(n661), .Z(n345) );
  NAND U674 ( .A(n662), .B(n294), .Z(n661) );
  XNOR U675 ( .A(n663), .B(n664), .Z(min_val_out[219]) );
  AND U676 ( .A(n568), .B(n665), .Z(n663) );
  XNOR U677 ( .A(n666), .B(n667), .Z(min_val_out[218]) );
  AND U678 ( .A(n568), .B(n668), .Z(n666) );
  XNOR U679 ( .A(n669), .B(n670), .Z(min_val_out[217]) );
  AND U680 ( .A(n568), .B(n671), .Z(n669) );
  XOR U681 ( .A(n672), .B(n673), .Z(min_val_out[216]) );
  AND U682 ( .A(n674), .B(n675), .Z(n672) );
  XOR U683 ( .A(n676), .B(n677), .Z(min_val_out[215]) );
  AND U684 ( .A(n674), .B(n678), .Z(n676) );
  XOR U685 ( .A(n679), .B(n680), .Z(min_val_out[214]) );
  AND U686 ( .A(n674), .B(n681), .Z(n679) );
  XOR U687 ( .A(n682), .B(n683), .Z(min_val_out[213]) );
  AND U688 ( .A(n674), .B(n684), .Z(n682) );
  XOR U689 ( .A(n685), .B(n686), .Z(min_val_out[212]) );
  AND U690 ( .A(n674), .B(n687), .Z(n685) );
  XOR U691 ( .A(n688), .B(n689), .Z(min_val_out[211]) );
  AND U692 ( .A(n674), .B(n690), .Z(n688) );
  XOR U693 ( .A(n691), .B(n692), .Z(min_val_out[210]) );
  AND U694 ( .A(n674), .B(n693), .Z(n691) );
  XOR U695 ( .A(\min_val_reg[0][20] ), .B(n694), .Z(min_val_out[20]) );
  AND U696 ( .A(n290), .B(n449), .Z(n694) );
  XNOR U697 ( .A(\min_val_reg[0][20] ), .B(n448), .Z(n449) );
  XOR U698 ( .A(\min_val_reg[1][20] ), .B(n695), .Z(n448) );
  NAND U699 ( .A(n349), .B(n316), .Z(n695) );
  XOR U700 ( .A(\min_val_reg[1][20] ), .B(n348), .Z(n349) );
  XNOR U701 ( .A(\min_val_reg[2][20] ), .B(n696), .Z(n348) );
  NAND U702 ( .A(n697), .B(n294), .Z(n696) );
  XOR U703 ( .A(n698), .B(n699), .Z(min_val_out[209]) );
  AND U704 ( .A(n674), .B(n700), .Z(n698) );
  XOR U705 ( .A(n701), .B(n702), .Z(min_val_out[208]) );
  AND U706 ( .A(n674), .B(n703), .Z(n701) );
  XOR U707 ( .A(n704), .B(n705), .Z(min_val_out[207]) );
  AND U708 ( .A(n674), .B(n706), .Z(n704) );
  XOR U709 ( .A(n707), .B(n708), .Z(min_val_out[206]) );
  AND U710 ( .A(n674), .B(n709), .Z(n707) );
  XOR U711 ( .A(n710), .B(n711), .Z(min_val_out[205]) );
  AND U712 ( .A(n674), .B(n712), .Z(n710) );
  XOR U713 ( .A(n713), .B(n714), .Z(min_val_out[204]) );
  AND U714 ( .A(n674), .B(n715), .Z(n713) );
  XOR U715 ( .A(n716), .B(n717), .Z(min_val_out[203]) );
  AND U716 ( .A(n674), .B(n718), .Z(n716) );
  XOR U717 ( .A(n719), .B(n720), .Z(min_val_out[202]) );
  AND U718 ( .A(n674), .B(n721), .Z(n719) );
  XOR U719 ( .A(n722), .B(n723), .Z(min_val_out[201]) );
  AND U720 ( .A(n674), .B(n724), .Z(n722) );
  XOR U721 ( .A(n725), .B(n726), .Z(min_val_out[200]) );
  AND U722 ( .A(n674), .B(n727), .Z(n725) );
  XOR U723 ( .A(\min_val_reg[0][1] ), .B(n728), .Z(min_val_out[1]) );
  AND U724 ( .A(n290), .B(n529), .Z(n728) );
  XNOR U725 ( .A(\min_val_reg[0][1] ), .B(n528), .Z(n529) );
  XOR U726 ( .A(\min_val_reg[1][1] ), .B(n729), .Z(n528) );
  NAND U727 ( .A(n410), .B(n316), .Z(n729) );
  XNOR U728 ( .A(\min_val_reg[1][1] ), .B(n409), .Z(n410) );
  XOR U729 ( .A(\min_val_reg[2][1] ), .B(n730), .Z(n409) );
  NAND U730 ( .A(n310), .B(n294), .Z(n730) );
  XOR U731 ( .A(\min_val_reg[2][1] ), .B(n309), .Z(n310) );
  XNOR U732 ( .A(\min_val_reg[3][1] ), .B(n731), .Z(n309) );
  NAND U733 ( .A(n732), .B(n505), .Z(n731) );
  XOR U734 ( .A(\min_val_reg[0][19] ), .B(n733), .Z(min_val_out[19]) );
  AND U735 ( .A(n290), .B(n452), .Z(n733) );
  XNOR U736 ( .A(\min_val_reg[0][19] ), .B(n451), .Z(n452) );
  XOR U737 ( .A(\min_val_reg[1][19] ), .B(n734), .Z(n451) );
  NAND U738 ( .A(n352), .B(n316), .Z(n734) );
  XOR U739 ( .A(\min_val_reg[1][19] ), .B(n351), .Z(n352) );
  XNOR U740 ( .A(\min_val_reg[2][19] ), .B(n735), .Z(n351) );
  NAND U741 ( .A(n736), .B(n294), .Z(n735) );
  XOR U742 ( .A(n737), .B(n738), .Z(min_val_out[199]) );
  AND U743 ( .A(n674), .B(n739), .Z(n737) );
  XOR U744 ( .A(n740), .B(n741), .Z(min_val_out[198]) );
  AND U745 ( .A(n674), .B(n742), .Z(n740) );
  XOR U746 ( .A(n743), .B(n744), .Z(min_val_out[197]) );
  AND U747 ( .A(n674), .B(n745), .Z(n743) );
  XOR U748 ( .A(n746), .B(n747), .Z(min_val_out[196]) );
  AND U749 ( .A(n674), .B(n748), .Z(n746) );
  XOR U750 ( .A(n749), .B(n750), .Z(min_val_out[195]) );
  AND U751 ( .A(n674), .B(n751), .Z(n749) );
  XOR U752 ( .A(n752), .B(n753), .Z(min_val_out[194]) );
  AND U753 ( .A(n674), .B(n754), .Z(n752) );
  XOR U754 ( .A(n755), .B(n756), .Z(min_val_out[193]) );
  AND U755 ( .A(n674), .B(n757), .Z(n755) );
  XOR U756 ( .A(n758), .B(n759), .Z(min_val_out[192]) );
  AND U757 ( .A(n674), .B(n760), .Z(n758) );
  XOR U758 ( .A(n761), .B(n762), .Z(min_val_out[191]) );
  AND U759 ( .A(n674), .B(n763), .Z(n761) );
  XOR U760 ( .A(n764), .B(n765), .Z(min_val_out[190]) );
  AND U761 ( .A(n674), .B(n766), .Z(n764) );
  XOR U762 ( .A(\min_val_reg[0][18] ), .B(n767), .Z(min_val_out[18]) );
  AND U763 ( .A(n290), .B(n457), .Z(n767) );
  XNOR U764 ( .A(\min_val_reg[0][18] ), .B(n456), .Z(n457) );
  XOR U765 ( .A(\min_val_reg[1][18] ), .B(n768), .Z(n456) );
  NAND U766 ( .A(n355), .B(n316), .Z(n768) );
  XOR U767 ( .A(\min_val_reg[1][18] ), .B(n354), .Z(n355) );
  XNOR U768 ( .A(\min_val_reg[2][18] ), .B(n769), .Z(n354) );
  NAND U769 ( .A(n770), .B(n294), .Z(n769) );
  XOR U770 ( .A(n771), .B(n772), .Z(min_val_out[189]) );
  AND U771 ( .A(n674), .B(n773), .Z(n771) );
  XOR U772 ( .A(n774), .B(n775), .Z(min_val_out[188]) );
  AND U773 ( .A(n674), .B(n776), .Z(n774) );
  XOR U774 ( .A(n777), .B(n778), .Z(min_val_out[187]) );
  AND U775 ( .A(n674), .B(n779), .Z(n777) );
  XOR U776 ( .A(n780), .B(n781), .Z(min_val_out[186]) );
  AND U777 ( .A(n674), .B(n782), .Z(n780) );
  XOR U778 ( .A(n783), .B(n784), .Z(min_val_out[185]) );
  AND U779 ( .A(n785), .B(n786), .Z(n783) );
  XOR U780 ( .A(n787), .B(n788), .Z(min_val_out[184]) );
  AND U781 ( .A(n785), .B(n789), .Z(n787) );
  XOR U782 ( .A(n790), .B(n791), .Z(min_val_out[183]) );
  AND U783 ( .A(n785), .B(n792), .Z(n790) );
  XOR U784 ( .A(n793), .B(n794), .Z(min_val_out[182]) );
  AND U785 ( .A(n785), .B(n795), .Z(n793) );
  XOR U786 ( .A(n796), .B(n797), .Z(min_val_out[181]) );
  AND U787 ( .A(n785), .B(n798), .Z(n796) );
  XOR U788 ( .A(n799), .B(n800), .Z(min_val_out[180]) );
  AND U789 ( .A(n785), .B(n801), .Z(n799) );
  XOR U790 ( .A(\min_val_reg[0][17] ), .B(n802), .Z(min_val_out[17]) );
  AND U791 ( .A(n290), .B(n460), .Z(n802) );
  XNOR U792 ( .A(\min_val_reg[0][17] ), .B(n459), .Z(n460) );
  XOR U793 ( .A(\min_val_reg[1][17] ), .B(n803), .Z(n459) );
  NAND U794 ( .A(n360), .B(n316), .Z(n803) );
  XOR U795 ( .A(\min_val_reg[1][17] ), .B(n359), .Z(n360) );
  XNOR U796 ( .A(\min_val_reg[2][17] ), .B(n804), .Z(n359) );
  NAND U797 ( .A(n805), .B(n294), .Z(n804) );
  XOR U798 ( .A(n806), .B(n807), .Z(min_val_out[179]) );
  AND U799 ( .A(n785), .B(n808), .Z(n806) );
  XOR U800 ( .A(n809), .B(n810), .Z(min_val_out[178]) );
  AND U801 ( .A(n785), .B(n811), .Z(n809) );
  XOR U802 ( .A(n812), .B(n813), .Z(min_val_out[177]) );
  AND U803 ( .A(n785), .B(n814), .Z(n812) );
  XOR U804 ( .A(n815), .B(n816), .Z(min_val_out[176]) );
  AND U805 ( .A(n785), .B(n817), .Z(n815) );
  XOR U806 ( .A(n818), .B(n819), .Z(min_val_out[175]) );
  AND U807 ( .A(n785), .B(n820), .Z(n818) );
  XOR U808 ( .A(n821), .B(n822), .Z(min_val_out[174]) );
  AND U809 ( .A(n785), .B(n823), .Z(n821) );
  XOR U810 ( .A(n824), .B(n825), .Z(min_val_out[173]) );
  AND U811 ( .A(n785), .B(n826), .Z(n824) );
  XOR U812 ( .A(n827), .B(n828), .Z(min_val_out[172]) );
  AND U813 ( .A(n785), .B(n829), .Z(n827) );
  XOR U814 ( .A(n830), .B(n831), .Z(min_val_out[171]) );
  AND U815 ( .A(n785), .B(n832), .Z(n830) );
  XOR U816 ( .A(n833), .B(n834), .Z(min_val_out[170]) );
  AND U817 ( .A(n785), .B(n835), .Z(n833) );
  XOR U818 ( .A(\min_val_reg[0][16] ), .B(n836), .Z(min_val_out[16]) );
  AND U819 ( .A(n290), .B(n463), .Z(n836) );
  XNOR U820 ( .A(\min_val_reg[0][16] ), .B(n462), .Z(n463) );
  XOR U821 ( .A(\min_val_reg[1][16] ), .B(n837), .Z(n462) );
  NAND U822 ( .A(n363), .B(n316), .Z(n837) );
  XOR U823 ( .A(\min_val_reg[1][16] ), .B(n362), .Z(n363) );
  XNOR U824 ( .A(\min_val_reg[2][16] ), .B(n838), .Z(n362) );
  NAND U825 ( .A(n839), .B(n294), .Z(n838) );
  XOR U826 ( .A(n840), .B(n841), .Z(min_val_out[169]) );
  AND U827 ( .A(n785), .B(n842), .Z(n840) );
  XOR U828 ( .A(n843), .B(n844), .Z(min_val_out[168]) );
  AND U829 ( .A(n785), .B(n845), .Z(n843) );
  XOR U830 ( .A(n846), .B(n847), .Z(min_val_out[167]) );
  AND U831 ( .A(n785), .B(n848), .Z(n846) );
  XOR U832 ( .A(n849), .B(n850), .Z(min_val_out[166]) );
  AND U833 ( .A(n785), .B(n851), .Z(n849) );
  XOR U834 ( .A(n852), .B(n853), .Z(min_val_out[165]) );
  AND U835 ( .A(n785), .B(n854), .Z(n852) );
  XOR U836 ( .A(n855), .B(n856), .Z(min_val_out[164]) );
  AND U837 ( .A(n785), .B(n857), .Z(n855) );
  XOR U838 ( .A(n858), .B(n859), .Z(min_val_out[163]) );
  AND U839 ( .A(n785), .B(n860), .Z(n858) );
  XOR U840 ( .A(n861), .B(n862), .Z(min_val_out[162]) );
  AND U841 ( .A(n785), .B(n863), .Z(n861) );
  XOR U842 ( .A(n864), .B(n865), .Z(min_val_out[161]) );
  AND U843 ( .A(n785), .B(n866), .Z(n864) );
  XOR U844 ( .A(n867), .B(n868), .Z(min_val_out[160]) );
  AND U845 ( .A(n785), .B(n869), .Z(n867) );
  XOR U846 ( .A(\min_val_reg[0][15] ), .B(n870), .Z(min_val_out[15]) );
  AND U847 ( .A(n290), .B(n466), .Z(n870) );
  XNOR U848 ( .A(\min_val_reg[0][15] ), .B(n465), .Z(n466) );
  XOR U849 ( .A(\min_val_reg[1][15] ), .B(n871), .Z(n465) );
  NAND U850 ( .A(n366), .B(n316), .Z(n871) );
  XOR U851 ( .A(\min_val_reg[1][15] ), .B(n365), .Z(n366) );
  XNOR U852 ( .A(\min_val_reg[2][15] ), .B(n872), .Z(n365) );
  NAND U853 ( .A(n873), .B(n294), .Z(n872) );
  XOR U854 ( .A(n874), .B(n875), .Z(min_val_out[159]) );
  AND U855 ( .A(n785), .B(n876), .Z(n874) );
  XOR U856 ( .A(n877), .B(n878), .Z(min_val_out[158]) );
  AND U857 ( .A(n785), .B(n879), .Z(n877) );
  XOR U858 ( .A(n880), .B(n881), .Z(min_val_out[157]) );
  AND U859 ( .A(n785), .B(n882), .Z(n880) );
  XOR U860 ( .A(n883), .B(n884), .Z(min_val_out[156]) );
  AND U861 ( .A(n785), .B(n885), .Z(n883) );
  XOR U862 ( .A(n886), .B(n887), .Z(min_val_out[155]) );
  AND U863 ( .A(n785), .B(n888), .Z(n886) );
  XOR U864 ( .A(n889), .B(n890), .Z(min_val_out[154]) );
  AND U865 ( .A(n505), .B(n891), .Z(n889) );
  XOR U866 ( .A(n892), .B(n893), .Z(min_val_out[153]) );
  AND U867 ( .A(n505), .B(n894), .Z(n892) );
  XOR U868 ( .A(n895), .B(n896), .Z(min_val_out[152]) );
  AND U869 ( .A(n505), .B(n897), .Z(n895) );
  XOR U870 ( .A(n898), .B(n899), .Z(min_val_out[151]) );
  AND U871 ( .A(n505), .B(n900), .Z(n898) );
  XOR U872 ( .A(n901), .B(n902), .Z(min_val_out[150]) );
  AND U873 ( .A(n505), .B(n903), .Z(n901) );
  XOR U874 ( .A(\min_val_reg[0][14] ), .B(n904), .Z(min_val_out[14]) );
  AND U875 ( .A(n290), .B(n469), .Z(n904) );
  XNOR U876 ( .A(\min_val_reg[0][14] ), .B(n468), .Z(n469) );
  XOR U877 ( .A(\min_val_reg[1][14] ), .B(n905), .Z(n468) );
  NAND U878 ( .A(n369), .B(n316), .Z(n905) );
  XOR U879 ( .A(\min_val_reg[1][14] ), .B(n368), .Z(n369) );
  XNOR U880 ( .A(\min_val_reg[2][14] ), .B(n906), .Z(n368) );
  NAND U881 ( .A(n907), .B(n294), .Z(n906) );
  XOR U882 ( .A(n908), .B(n909), .Z(min_val_out[149]) );
  AND U883 ( .A(n505), .B(n910), .Z(n908) );
  XOR U884 ( .A(n911), .B(n912), .Z(min_val_out[148]) );
  AND U885 ( .A(n505), .B(n913), .Z(n911) );
  XOR U886 ( .A(n914), .B(n915), .Z(min_val_out[147]) );
  AND U887 ( .A(n505), .B(n916), .Z(n914) );
  XOR U888 ( .A(n917), .B(n918), .Z(min_val_out[146]) );
  AND U889 ( .A(n505), .B(n919), .Z(n917) );
  XOR U890 ( .A(n920), .B(n921), .Z(min_val_out[145]) );
  AND U891 ( .A(n505), .B(n922), .Z(n920) );
  XOR U892 ( .A(n923), .B(n924), .Z(min_val_out[144]) );
  AND U893 ( .A(n505), .B(n925), .Z(n923) );
  XOR U894 ( .A(n926), .B(n927), .Z(min_val_out[143]) );
  AND U895 ( .A(n505), .B(n928), .Z(n926) );
  XOR U896 ( .A(n929), .B(n930), .Z(min_val_out[142]) );
  AND U897 ( .A(n505), .B(n931), .Z(n929) );
  XOR U898 ( .A(n932), .B(n933), .Z(min_val_out[141]) );
  AND U899 ( .A(n505), .B(n934), .Z(n932) );
  XOR U900 ( .A(n935), .B(n936), .Z(min_val_out[140]) );
  AND U901 ( .A(n505), .B(n937), .Z(n935) );
  XOR U902 ( .A(\min_val_reg[0][13] ), .B(n938), .Z(min_val_out[13]) );
  AND U903 ( .A(n290), .B(n472), .Z(n938) );
  XNOR U904 ( .A(\min_val_reg[0][13] ), .B(n471), .Z(n472) );
  XOR U905 ( .A(\min_val_reg[1][13] ), .B(n939), .Z(n471) );
  NAND U906 ( .A(n372), .B(n316), .Z(n939) );
  XOR U907 ( .A(\min_val_reg[1][13] ), .B(n371), .Z(n372) );
  XNOR U908 ( .A(\min_val_reg[2][13] ), .B(n940), .Z(n371) );
  NAND U909 ( .A(n941), .B(n294), .Z(n940) );
  XOR U910 ( .A(n942), .B(n943), .Z(min_val_out[139]) );
  AND U911 ( .A(n505), .B(n944), .Z(n942) );
  XOR U912 ( .A(n945), .B(n946), .Z(min_val_out[138]) );
  AND U913 ( .A(n505), .B(n947), .Z(n945) );
  XOR U914 ( .A(n948), .B(n949), .Z(min_val_out[137]) );
  AND U915 ( .A(n505), .B(n950), .Z(n948) );
  XOR U916 ( .A(n951), .B(n952), .Z(min_val_out[136]) );
  AND U917 ( .A(n505), .B(n953), .Z(n951) );
  XOR U918 ( .A(n954), .B(n955), .Z(min_val_out[135]) );
  AND U919 ( .A(n505), .B(n956), .Z(n954) );
  XOR U920 ( .A(n957), .B(n958), .Z(min_val_out[134]) );
  AND U921 ( .A(n505), .B(n959), .Z(n957) );
  XOR U922 ( .A(n960), .B(n961), .Z(min_val_out[133]) );
  AND U923 ( .A(n505), .B(n962), .Z(n960) );
  XOR U924 ( .A(n963), .B(n964), .Z(min_val_out[132]) );
  AND U925 ( .A(n505), .B(n965), .Z(n963) );
  XOR U926 ( .A(n966), .B(n967), .Z(min_val_out[131]) );
  AND U927 ( .A(n505), .B(n968), .Z(n966) );
  XOR U928 ( .A(n969), .B(n970), .Z(min_val_out[130]) );
  AND U929 ( .A(n505), .B(n504), .Z(n969) );
  XOR U930 ( .A(\min_val_reg[3][6] ), .B(n970), .Z(n504) );
  XNOR U931 ( .A(\min_val_reg[4][6] ), .B(n971), .Z(n970) );
  NAND U932 ( .A(n866), .B(n785), .Z(n971) );
  XOR U933 ( .A(\min_val_reg[4][6] ), .B(n865), .Z(n866) );
  XNOR U934 ( .A(\min_val_reg[5][6] ), .B(n972), .Z(n865) );
  NAND U935 ( .A(n760), .B(n674), .Z(n972) );
  XOR U936 ( .A(\min_val_reg[5][6] ), .B(n759), .Z(n760) );
  XNOR U937 ( .A(\min_val_reg[6][6] ), .B(n973), .Z(n759) );
  NAND U938 ( .A(n649), .B(n974), .Z(n973) );
  XNOR U939 ( .A(\min_val_reg[6][6] ), .B(n648), .Z(n649) );
  XOR U940 ( .A(\min_val_reg[7][6] ), .B(n975), .Z(n648) );
  NAND U941 ( .A(n976), .B(n977), .Z(n975) );
  XOR U942 ( .A(\min_val_reg[7][6] ), .B(DB[6]), .Z(n976) );
  XOR U943 ( .A(\min_val_reg[0][12] ), .B(n978), .Z(min_val_out[12]) );
  AND U944 ( .A(n290), .B(n475), .Z(n978) );
  XNOR U945 ( .A(\min_val_reg[0][12] ), .B(n474), .Z(n475) );
  XOR U946 ( .A(\min_val_reg[1][12] ), .B(n979), .Z(n474) );
  NAND U947 ( .A(n375), .B(n316), .Z(n979) );
  XOR U948 ( .A(\min_val_reg[1][12] ), .B(n374), .Z(n375) );
  XNOR U949 ( .A(\min_val_reg[2][12] ), .B(n980), .Z(n374) );
  NAND U950 ( .A(n981), .B(n294), .Z(n980) );
  XOR U951 ( .A(n982), .B(n983), .Z(min_val_out[129]) );
  AND U952 ( .A(n505), .B(n511), .Z(n982) );
  XOR U953 ( .A(\min_val_reg[3][5] ), .B(n983), .Z(n511) );
  XNOR U954 ( .A(\min_val_reg[4][5] ), .B(n984), .Z(n983) );
  NAND U955 ( .A(n869), .B(n785), .Z(n984) );
  XOR U956 ( .A(\min_val_reg[4][5] ), .B(n868), .Z(n869) );
  XNOR U957 ( .A(\min_val_reg[5][5] ), .B(n985), .Z(n868) );
  NAND U958 ( .A(n763), .B(n674), .Z(n985) );
  XOR U959 ( .A(\min_val_reg[5][5] ), .B(n762), .Z(n763) );
  XNOR U960 ( .A(\min_val_reg[6][5] ), .B(n986), .Z(n762) );
  NAND U961 ( .A(n652), .B(n974), .Z(n986) );
  XNOR U962 ( .A(\min_val_reg[6][5] ), .B(n651), .Z(n652) );
  XOR U963 ( .A(\min_val_reg[7][5] ), .B(n987), .Z(n651) );
  NAND U964 ( .A(n988), .B(n977), .Z(n987) );
  XOR U965 ( .A(\min_val_reg[7][5] ), .B(DB[5]), .Z(n988) );
  XOR U966 ( .A(n989), .B(n990), .Z(min_val_out[128]) );
  AND U967 ( .A(n505), .B(n517), .Z(n989) );
  XOR U968 ( .A(\min_val_reg[3][4] ), .B(n990), .Z(n517) );
  XNOR U969 ( .A(\min_val_reg[4][4] ), .B(n991), .Z(n990) );
  NAND U970 ( .A(n876), .B(n785), .Z(n991) );
  XOR U971 ( .A(\min_val_reg[4][4] ), .B(n875), .Z(n876) );
  XNOR U972 ( .A(\min_val_reg[5][4] ), .B(n992), .Z(n875) );
  NAND U973 ( .A(n766), .B(n674), .Z(n992) );
  XOR U974 ( .A(\min_val_reg[5][4] ), .B(n765), .Z(n766) );
  XNOR U975 ( .A(\min_val_reg[6][4] ), .B(n993), .Z(n765) );
  NAND U976 ( .A(n655), .B(n974), .Z(n993) );
  XNOR U977 ( .A(\min_val_reg[6][4] ), .B(n654), .Z(n655) );
  XOR U978 ( .A(\min_val_reg[7][4] ), .B(n994), .Z(n654) );
  NAND U979 ( .A(n995), .B(n977), .Z(n994) );
  XOR U980 ( .A(\min_val_reg[7][4] ), .B(DB[4]), .Z(n995) );
  XOR U981 ( .A(n996), .B(n997), .Z(min_val_out[127]) );
  AND U982 ( .A(n505), .B(n523), .Z(n996) );
  XOR U983 ( .A(\min_val_reg[3][3] ), .B(n997), .Z(n523) );
  XNOR U984 ( .A(\min_val_reg[4][3] ), .B(n998), .Z(n997) );
  NAND U985 ( .A(n879), .B(n785), .Z(n998) );
  XOR U986 ( .A(\min_val_reg[4][3] ), .B(n878), .Z(n879) );
  XNOR U987 ( .A(\min_val_reg[5][3] ), .B(n999), .Z(n878) );
  NAND U988 ( .A(n773), .B(n674), .Z(n999) );
  XOR U989 ( .A(\min_val_reg[5][3] ), .B(n772), .Z(n773) );
  XNOR U990 ( .A(\min_val_reg[6][3] ), .B(n1000), .Z(n772) );
  NAND U991 ( .A(n658), .B(n974), .Z(n1000) );
  XNOR U992 ( .A(\min_val_reg[6][3] ), .B(n657), .Z(n658) );
  XOR U993 ( .A(\min_val_reg[7][3] ), .B(n1001), .Z(n657) );
  NAND U994 ( .A(n1002), .B(n977), .Z(n1001) );
  XOR U995 ( .A(\min_val_reg[7][3] ), .B(DB[3]), .Z(n1002) );
  XOR U996 ( .A(n1003), .B(n1004), .Z(min_val_out[126]) );
  AND U997 ( .A(n505), .B(n541), .Z(n1003) );
  XOR U998 ( .A(\min_val_reg[3][2] ), .B(n1004), .Z(n541) );
  XNOR U999 ( .A(\min_val_reg[4][2] ), .B(n1005), .Z(n1004) );
  NAND U1000 ( .A(n882), .B(n785), .Z(n1005) );
  XOR U1001 ( .A(\min_val_reg[4][2] ), .B(n881), .Z(n882) );
  XNOR U1002 ( .A(\min_val_reg[5][2] ), .B(n1006), .Z(n881) );
  NAND U1003 ( .A(n776), .B(n674), .Z(n1006) );
  XOR U1004 ( .A(\min_val_reg[5][2] ), .B(n775), .Z(n776) );
  XNOR U1005 ( .A(\min_val_reg[6][2] ), .B(n1007), .Z(n775) );
  NAND U1006 ( .A(n665), .B(n974), .Z(n1007) );
  XNOR U1007 ( .A(\min_val_reg[6][2] ), .B(n664), .Z(n665) );
  XOR U1008 ( .A(\min_val_reg[7][2] ), .B(n1008), .Z(n664) );
  NAND U1009 ( .A(n1009), .B(n977), .Z(n1008) );
  XOR U1010 ( .A(\min_val_reg[7][2] ), .B(DB[2]), .Z(n1009) );
  XOR U1011 ( .A(n1010), .B(n1011), .Z(min_val_out[125]) );
  AND U1012 ( .A(n505), .B(n732), .Z(n1010) );
  XOR U1013 ( .A(\min_val_reg[3][1] ), .B(n1011), .Z(n732) );
  XNOR U1014 ( .A(\min_val_reg[4][1] ), .B(n1012), .Z(n1011) );
  NAND U1015 ( .A(n885), .B(n785), .Z(n1012) );
  XOR U1016 ( .A(\min_val_reg[4][1] ), .B(n884), .Z(n885) );
  XNOR U1017 ( .A(\min_val_reg[5][1] ), .B(n1013), .Z(n884) );
  NAND U1018 ( .A(n779), .B(n674), .Z(n1013) );
  XOR U1019 ( .A(\min_val_reg[5][1] ), .B(n778), .Z(n779) );
  XNOR U1020 ( .A(\min_val_reg[6][1] ), .B(n1014), .Z(n778) );
  NAND U1021 ( .A(n668), .B(n974), .Z(n1014) );
  XNOR U1022 ( .A(\min_val_reg[6][1] ), .B(n667), .Z(n668) );
  XOR U1023 ( .A(\min_val_reg[7][1] ), .B(n1015), .Z(n667) );
  NAND U1024 ( .A(n1016), .B(n977), .Z(n1015) );
  XOR U1025 ( .A(\min_val_reg[7][1] ), .B(DB[1]), .Z(n1016) );
  XOR U1026 ( .A(n1017), .B(n1018), .Z(min_val_out[124]) );
  AND U1027 ( .A(n505), .B(n1019), .Z(n1017) );
  XOR U1028 ( .A(n1020), .B(n1021), .Z(min_val_out[123]) );
  AND U1029 ( .A(n294), .B(n536), .Z(n1020) );
  XOR U1030 ( .A(\min_val_reg[2][30] ), .B(n1021), .Z(n536) );
  XNOR U1031 ( .A(\min_val_reg[3][30] ), .B(n1022), .Z(n1021) );
  NAND U1032 ( .A(n891), .B(n505), .Z(n1022) );
  XOR U1033 ( .A(\min_val_reg[3][30] ), .B(n890), .Z(n891) );
  XNOR U1034 ( .A(\min_val_reg[4][30] ), .B(n1023), .Z(n890) );
  NAND U1035 ( .A(n786), .B(n785), .Z(n1023) );
  XOR U1036 ( .A(\min_val_reg[4][30] ), .B(n784), .Z(n786) );
  XNOR U1037 ( .A(\min_val_reg[5][30] ), .B(n1024), .Z(n784) );
  NAND U1038 ( .A(n675), .B(n674), .Z(n1024) );
  XOR U1039 ( .A(\min_val_reg[5][30] ), .B(n673), .Z(n675) );
  XNOR U1040 ( .A(\min_val_reg[6][30] ), .B(n1025), .Z(n673) );
  NAND U1041 ( .A(n569), .B(n974), .Z(n1025) );
  XNOR U1042 ( .A(\min_val_reg[6][30] ), .B(n567), .Z(n569) );
  XOR U1043 ( .A(\min_val_reg[7][30] ), .B(n1026), .Z(n567) );
  NAND U1044 ( .A(n1027), .B(n977), .Z(n1026) );
  XOR U1045 ( .A(\min_val_reg[7][30] ), .B(DB[30]), .Z(n1027) );
  XOR U1046 ( .A(n1028), .B(n1029), .Z(min_val_out[122]) );
  AND U1047 ( .A(n294), .B(n545), .Z(n1028) );
  XOR U1048 ( .A(\min_val_reg[2][29] ), .B(n1029), .Z(n545) );
  XNOR U1049 ( .A(\min_val_reg[3][29] ), .B(n1030), .Z(n1029) );
  NAND U1050 ( .A(n894), .B(n505), .Z(n1030) );
  XOR U1051 ( .A(\min_val_reg[3][29] ), .B(n893), .Z(n894) );
  XNOR U1052 ( .A(\min_val_reg[4][29] ), .B(n1031), .Z(n893) );
  NAND U1053 ( .A(n789), .B(n785), .Z(n1031) );
  XOR U1054 ( .A(\min_val_reg[4][29] ), .B(n788), .Z(n789) );
  XNOR U1055 ( .A(\min_val_reg[5][29] ), .B(n1032), .Z(n788) );
  NAND U1056 ( .A(n678), .B(n674), .Z(n1032) );
  XOR U1057 ( .A(\min_val_reg[5][29] ), .B(n677), .Z(n678) );
  XNOR U1058 ( .A(\min_val_reg[6][29] ), .B(n1033), .Z(n677) );
  NAND U1059 ( .A(n572), .B(n974), .Z(n1033) );
  XNOR U1060 ( .A(\min_val_reg[6][29] ), .B(n571), .Z(n572) );
  XOR U1061 ( .A(\min_val_reg[7][29] ), .B(n1034), .Z(n571) );
  NAND U1062 ( .A(n1035), .B(n977), .Z(n1034) );
  XOR U1063 ( .A(\min_val_reg[7][29] ), .B(DB[29]), .Z(n1035) );
  XOR U1064 ( .A(n1036), .B(n1037), .Z(min_val_out[121]) );
  AND U1065 ( .A(n294), .B(n549), .Z(n1036) );
  XOR U1066 ( .A(\min_val_reg[2][28] ), .B(n1037), .Z(n549) );
  XNOR U1067 ( .A(\min_val_reg[3][28] ), .B(n1038), .Z(n1037) );
  NAND U1068 ( .A(n897), .B(n505), .Z(n1038) );
  XOR U1069 ( .A(\min_val_reg[3][28] ), .B(n896), .Z(n897) );
  XNOR U1070 ( .A(\min_val_reg[4][28] ), .B(n1039), .Z(n896) );
  NAND U1071 ( .A(n792), .B(n785), .Z(n1039) );
  XOR U1072 ( .A(\min_val_reg[4][28] ), .B(n791), .Z(n792) );
  XNOR U1073 ( .A(\min_val_reg[5][28] ), .B(n1040), .Z(n791) );
  NAND U1074 ( .A(n681), .B(n674), .Z(n1040) );
  XOR U1075 ( .A(\min_val_reg[5][28] ), .B(n680), .Z(n681) );
  XNOR U1076 ( .A(\min_val_reg[6][28] ), .B(n1041), .Z(n680) );
  NAND U1077 ( .A(n575), .B(n974), .Z(n1041) );
  XNOR U1078 ( .A(\min_val_reg[6][28] ), .B(n574), .Z(n575) );
  XOR U1079 ( .A(\min_val_reg[7][28] ), .B(n1042), .Z(n574) );
  NAND U1080 ( .A(n1043), .B(n977), .Z(n1042) );
  XOR U1081 ( .A(\min_val_reg[7][28] ), .B(DB[28]), .Z(n1043) );
  XOR U1082 ( .A(n1044), .B(n1045), .Z(min_val_out[120]) );
  AND U1083 ( .A(n294), .B(n553), .Z(n1044) );
  XOR U1084 ( .A(\min_val_reg[2][27] ), .B(n1045), .Z(n553) );
  XNOR U1085 ( .A(\min_val_reg[3][27] ), .B(n1046), .Z(n1045) );
  NAND U1086 ( .A(n900), .B(n505), .Z(n1046) );
  XOR U1087 ( .A(\min_val_reg[3][27] ), .B(n899), .Z(n900) );
  XNOR U1088 ( .A(\min_val_reg[4][27] ), .B(n1047), .Z(n899) );
  NAND U1089 ( .A(n795), .B(n785), .Z(n1047) );
  XOR U1090 ( .A(\min_val_reg[4][27] ), .B(n794), .Z(n795) );
  XNOR U1091 ( .A(\min_val_reg[5][27] ), .B(n1048), .Z(n794) );
  NAND U1092 ( .A(n684), .B(n674), .Z(n1048) );
  XOR U1093 ( .A(\min_val_reg[5][27] ), .B(n683), .Z(n684) );
  XNOR U1094 ( .A(\min_val_reg[6][27] ), .B(n1049), .Z(n683) );
  NAND U1095 ( .A(n578), .B(n974), .Z(n1049) );
  XNOR U1096 ( .A(\min_val_reg[6][27] ), .B(n577), .Z(n578) );
  XOR U1097 ( .A(\min_val_reg[7][27] ), .B(n1050), .Z(n577) );
  NAND U1098 ( .A(n1051), .B(n977), .Z(n1050) );
  XOR U1099 ( .A(\min_val_reg[7][27] ), .B(DB[27]), .Z(n1051) );
  XOR U1100 ( .A(\min_val_reg[0][11] ), .B(n1052), .Z(min_val_out[11]) );
  AND U1101 ( .A(n290), .B(n478), .Z(n1052) );
  XNOR U1102 ( .A(\min_val_reg[0][11] ), .B(n477), .Z(n478) );
  XOR U1103 ( .A(\min_val_reg[1][11] ), .B(n1053), .Z(n477) );
  NAND U1104 ( .A(n378), .B(n316), .Z(n1053) );
  XOR U1105 ( .A(\min_val_reg[1][11] ), .B(n377), .Z(n378) );
  XNOR U1106 ( .A(\min_val_reg[2][11] ), .B(n1054), .Z(n377) );
  NAND U1107 ( .A(n1055), .B(n294), .Z(n1054) );
  XOR U1108 ( .A(n1056), .B(n1057), .Z(min_val_out[119]) );
  AND U1109 ( .A(n294), .B(n557), .Z(n1056) );
  XOR U1110 ( .A(\min_val_reg[2][26] ), .B(n1057), .Z(n557) );
  XNOR U1111 ( .A(\min_val_reg[3][26] ), .B(n1058), .Z(n1057) );
  NAND U1112 ( .A(n903), .B(n505), .Z(n1058) );
  XOR U1113 ( .A(\min_val_reg[3][26] ), .B(n902), .Z(n903) );
  XNOR U1114 ( .A(\min_val_reg[4][26] ), .B(n1059), .Z(n902) );
  NAND U1115 ( .A(n798), .B(n785), .Z(n1059) );
  XOR U1116 ( .A(\min_val_reg[4][26] ), .B(n797), .Z(n798) );
  XNOR U1117 ( .A(\min_val_reg[5][26] ), .B(n1060), .Z(n797) );
  NAND U1118 ( .A(n687), .B(n674), .Z(n1060) );
  XOR U1119 ( .A(\min_val_reg[5][26] ), .B(n686), .Z(n687) );
  XNOR U1120 ( .A(\min_val_reg[6][26] ), .B(n1061), .Z(n686) );
  NAND U1121 ( .A(n581), .B(n974), .Z(n1061) );
  XNOR U1122 ( .A(\min_val_reg[6][26] ), .B(n580), .Z(n581) );
  XOR U1123 ( .A(\min_val_reg[7][26] ), .B(n1062), .Z(n580) );
  NAND U1124 ( .A(n1063), .B(n977), .Z(n1062) );
  XOR U1125 ( .A(\min_val_reg[7][26] ), .B(DB[26]), .Z(n1063) );
  XOR U1126 ( .A(n1064), .B(n1065), .Z(min_val_out[118]) );
  AND U1127 ( .A(n294), .B(n561), .Z(n1064) );
  XOR U1128 ( .A(\min_val_reg[2][25] ), .B(n1065), .Z(n561) );
  XNOR U1129 ( .A(\min_val_reg[3][25] ), .B(n1066), .Z(n1065) );
  NAND U1130 ( .A(n910), .B(n505), .Z(n1066) );
  XOR U1131 ( .A(\min_val_reg[3][25] ), .B(n909), .Z(n910) );
  XNOR U1132 ( .A(\min_val_reg[4][25] ), .B(n1067), .Z(n909) );
  NAND U1133 ( .A(n801), .B(n785), .Z(n1067) );
  XOR U1134 ( .A(\min_val_reg[4][25] ), .B(n800), .Z(n801) );
  XNOR U1135 ( .A(\min_val_reg[5][25] ), .B(n1068), .Z(n800) );
  NAND U1136 ( .A(n690), .B(n674), .Z(n1068) );
  XOR U1137 ( .A(\min_val_reg[5][25] ), .B(n689), .Z(n690) );
  XNOR U1138 ( .A(\min_val_reg[6][25] ), .B(n1069), .Z(n689) );
  NAND U1139 ( .A(n584), .B(n974), .Z(n1069) );
  XNOR U1140 ( .A(\min_val_reg[6][25] ), .B(n583), .Z(n584) );
  XOR U1141 ( .A(\min_val_reg[7][25] ), .B(n1070), .Z(n583) );
  NAND U1142 ( .A(n1071), .B(n977), .Z(n1070) );
  XOR U1143 ( .A(\min_val_reg[7][25] ), .B(DB[25]), .Z(n1071) );
  XOR U1144 ( .A(n1072), .B(n1073), .Z(min_val_out[117]) );
  AND U1145 ( .A(n294), .B(n565), .Z(n1072) );
  XOR U1146 ( .A(\min_val_reg[2][24] ), .B(n1073), .Z(n565) );
  XNOR U1147 ( .A(\min_val_reg[3][24] ), .B(n1074), .Z(n1073) );
  NAND U1148 ( .A(n913), .B(n505), .Z(n1074) );
  XOR U1149 ( .A(\min_val_reg[3][24] ), .B(n912), .Z(n913) );
  XNOR U1150 ( .A(\min_val_reg[4][24] ), .B(n1075), .Z(n912) );
  NAND U1151 ( .A(n808), .B(n785), .Z(n1075) );
  XOR U1152 ( .A(\min_val_reg[4][24] ), .B(n807), .Z(n808) );
  XNOR U1153 ( .A(\min_val_reg[5][24] ), .B(n1076), .Z(n807) );
  NAND U1154 ( .A(n693), .B(n674), .Z(n1076) );
  XOR U1155 ( .A(\min_val_reg[5][24] ), .B(n692), .Z(n693) );
  XNOR U1156 ( .A(\min_val_reg[6][24] ), .B(n1077), .Z(n692) );
  NAND U1157 ( .A(n587), .B(n974), .Z(n1077) );
  XNOR U1158 ( .A(\min_val_reg[6][24] ), .B(n586), .Z(n587) );
  XOR U1159 ( .A(\min_val_reg[7][24] ), .B(n1078), .Z(n586) );
  NAND U1160 ( .A(n1079), .B(n977), .Z(n1078) );
  XOR U1161 ( .A(\min_val_reg[7][24] ), .B(DB[24]), .Z(n1079) );
  XOR U1162 ( .A(n1080), .B(n1081), .Z(min_val_out[116]) );
  AND U1163 ( .A(n294), .B(n594), .Z(n1080) );
  XOR U1164 ( .A(\min_val_reg[2][23] ), .B(n1081), .Z(n594) );
  XNOR U1165 ( .A(\min_val_reg[3][23] ), .B(n1082), .Z(n1081) );
  NAND U1166 ( .A(n916), .B(n505), .Z(n1082) );
  XOR U1167 ( .A(\min_val_reg[3][23] ), .B(n915), .Z(n916) );
  XNOR U1168 ( .A(\min_val_reg[4][23] ), .B(n1083), .Z(n915) );
  NAND U1169 ( .A(n811), .B(n785), .Z(n1083) );
  XOR U1170 ( .A(\min_val_reg[4][23] ), .B(n810), .Z(n811) );
  XNOR U1171 ( .A(\min_val_reg[5][23] ), .B(n1084), .Z(n810) );
  NAND U1172 ( .A(n700), .B(n674), .Z(n1084) );
  XOR U1173 ( .A(\min_val_reg[5][23] ), .B(n699), .Z(n700) );
  XNOR U1174 ( .A(\min_val_reg[6][23] ), .B(n1085), .Z(n699) );
  NAND U1175 ( .A(n590), .B(n974), .Z(n1085) );
  XNOR U1176 ( .A(\min_val_reg[6][23] ), .B(n589), .Z(n590) );
  XOR U1177 ( .A(\min_val_reg[7][23] ), .B(n1086), .Z(n589) );
  NAND U1178 ( .A(n1087), .B(n977), .Z(n1086) );
  XOR U1179 ( .A(\min_val_reg[7][23] ), .B(DB[23]), .Z(n1087) );
  XOR U1180 ( .A(n1088), .B(n1089), .Z(min_val_out[115]) );
  AND U1181 ( .A(n294), .B(n628), .Z(n1088) );
  XOR U1182 ( .A(\min_val_reg[2][22] ), .B(n1089), .Z(n628) );
  XNOR U1183 ( .A(\min_val_reg[3][22] ), .B(n1090), .Z(n1089) );
  NAND U1184 ( .A(n919), .B(n505), .Z(n1090) );
  XOR U1185 ( .A(\min_val_reg[3][22] ), .B(n918), .Z(n919) );
  XNOR U1186 ( .A(\min_val_reg[4][22] ), .B(n1091), .Z(n918) );
  NAND U1187 ( .A(n814), .B(n785), .Z(n1091) );
  XOR U1188 ( .A(\min_val_reg[4][22] ), .B(n813), .Z(n814) );
  XNOR U1189 ( .A(\min_val_reg[5][22] ), .B(n1092), .Z(n813) );
  NAND U1190 ( .A(n703), .B(n674), .Z(n1092) );
  XOR U1191 ( .A(\min_val_reg[5][22] ), .B(n702), .Z(n703) );
  XNOR U1192 ( .A(\min_val_reg[6][22] ), .B(n1093), .Z(n702) );
  NAND U1193 ( .A(n597), .B(n974), .Z(n1093) );
  XNOR U1194 ( .A(\min_val_reg[6][22] ), .B(n596), .Z(n597) );
  XOR U1195 ( .A(\min_val_reg[7][22] ), .B(n1094), .Z(n596) );
  NAND U1196 ( .A(n1095), .B(n977), .Z(n1094) );
  XOR U1197 ( .A(\min_val_reg[7][22] ), .B(DB[22]), .Z(n1095) );
  XOR U1198 ( .A(n1096), .B(n1097), .Z(min_val_out[114]) );
  AND U1199 ( .A(n294), .B(n662), .Z(n1096) );
  XOR U1200 ( .A(\min_val_reg[2][21] ), .B(n1097), .Z(n662) );
  XNOR U1201 ( .A(\min_val_reg[3][21] ), .B(n1098), .Z(n1097) );
  NAND U1202 ( .A(n922), .B(n505), .Z(n1098) );
  XOR U1203 ( .A(\min_val_reg[3][21] ), .B(n921), .Z(n922) );
  XNOR U1204 ( .A(\min_val_reg[4][21] ), .B(n1099), .Z(n921) );
  NAND U1205 ( .A(n817), .B(n785), .Z(n1099) );
  XOR U1206 ( .A(\min_val_reg[4][21] ), .B(n816), .Z(n817) );
  XNOR U1207 ( .A(\min_val_reg[5][21] ), .B(n1100), .Z(n816) );
  NAND U1208 ( .A(n706), .B(n674), .Z(n1100) );
  XOR U1209 ( .A(\min_val_reg[5][21] ), .B(n705), .Z(n706) );
  XNOR U1210 ( .A(\min_val_reg[6][21] ), .B(n1101), .Z(n705) );
  NAND U1211 ( .A(n600), .B(n974), .Z(n1101) );
  XNOR U1212 ( .A(\min_val_reg[6][21] ), .B(n599), .Z(n600) );
  XOR U1213 ( .A(\min_val_reg[7][21] ), .B(n1102), .Z(n599) );
  NAND U1214 ( .A(n1103), .B(n977), .Z(n1102) );
  XOR U1215 ( .A(\min_val_reg[7][21] ), .B(DB[21]), .Z(n1103) );
  XOR U1216 ( .A(n1104), .B(n1105), .Z(min_val_out[113]) );
  AND U1217 ( .A(n294), .B(n697), .Z(n1104) );
  XOR U1218 ( .A(\min_val_reg[2][20] ), .B(n1105), .Z(n697) );
  XNOR U1219 ( .A(\min_val_reg[3][20] ), .B(n1106), .Z(n1105) );
  NAND U1220 ( .A(n925), .B(n505), .Z(n1106) );
  XOR U1221 ( .A(\min_val_reg[3][20] ), .B(n924), .Z(n925) );
  XNOR U1222 ( .A(\min_val_reg[4][20] ), .B(n1107), .Z(n924) );
  NAND U1223 ( .A(n820), .B(n785), .Z(n1107) );
  XOR U1224 ( .A(\min_val_reg[4][20] ), .B(n819), .Z(n820) );
  XNOR U1225 ( .A(\min_val_reg[5][20] ), .B(n1108), .Z(n819) );
  NAND U1226 ( .A(n709), .B(n674), .Z(n1108) );
  XOR U1227 ( .A(\min_val_reg[5][20] ), .B(n708), .Z(n709) );
  XNOR U1228 ( .A(\min_val_reg[6][20] ), .B(n1109), .Z(n708) );
  NAND U1229 ( .A(n603), .B(n974), .Z(n1109) );
  XNOR U1230 ( .A(\min_val_reg[6][20] ), .B(n602), .Z(n603) );
  XOR U1231 ( .A(\min_val_reg[7][20] ), .B(n1110), .Z(n602) );
  NAND U1232 ( .A(n1111), .B(n977), .Z(n1110) );
  XOR U1233 ( .A(\min_val_reg[7][20] ), .B(DB[20]), .Z(n1111) );
  XOR U1234 ( .A(n1112), .B(n1113), .Z(min_val_out[112]) );
  AND U1235 ( .A(n294), .B(n736), .Z(n1112) );
  XOR U1236 ( .A(\min_val_reg[2][19] ), .B(n1113), .Z(n736) );
  XNOR U1237 ( .A(\min_val_reg[3][19] ), .B(n1114), .Z(n1113) );
  NAND U1238 ( .A(n928), .B(n505), .Z(n1114) );
  XOR U1239 ( .A(\min_val_reg[3][19] ), .B(n927), .Z(n928) );
  XNOR U1240 ( .A(\min_val_reg[4][19] ), .B(n1115), .Z(n927) );
  NAND U1241 ( .A(n823), .B(n785), .Z(n1115) );
  XOR U1242 ( .A(\min_val_reg[4][19] ), .B(n822), .Z(n823) );
  XNOR U1243 ( .A(\min_val_reg[5][19] ), .B(n1116), .Z(n822) );
  NAND U1244 ( .A(n712), .B(n674), .Z(n1116) );
  XOR U1245 ( .A(\min_val_reg[5][19] ), .B(n711), .Z(n712) );
  XNOR U1246 ( .A(\min_val_reg[6][19] ), .B(n1117), .Z(n711) );
  NAND U1247 ( .A(n606), .B(n974), .Z(n1117) );
  XNOR U1248 ( .A(\min_val_reg[6][19] ), .B(n605), .Z(n606) );
  XOR U1249 ( .A(\min_val_reg[7][19] ), .B(n1118), .Z(n605) );
  NAND U1250 ( .A(n1119), .B(n977), .Z(n1118) );
  XOR U1251 ( .A(\min_val_reg[7][19] ), .B(DB[19]), .Z(n1119) );
  XOR U1252 ( .A(n1120), .B(n1121), .Z(min_val_out[111]) );
  AND U1253 ( .A(n294), .B(n770), .Z(n1120) );
  XOR U1254 ( .A(\min_val_reg[2][18] ), .B(n1121), .Z(n770) );
  XNOR U1255 ( .A(\min_val_reg[3][18] ), .B(n1122), .Z(n1121) );
  NAND U1256 ( .A(n931), .B(n505), .Z(n1122) );
  XOR U1257 ( .A(\min_val_reg[3][18] ), .B(n930), .Z(n931) );
  XNOR U1258 ( .A(\min_val_reg[4][18] ), .B(n1123), .Z(n930) );
  NAND U1259 ( .A(n826), .B(n785), .Z(n1123) );
  XOR U1260 ( .A(\min_val_reg[4][18] ), .B(n825), .Z(n826) );
  XNOR U1261 ( .A(\min_val_reg[5][18] ), .B(n1124), .Z(n825) );
  NAND U1262 ( .A(n715), .B(n674), .Z(n1124) );
  XOR U1263 ( .A(\min_val_reg[5][18] ), .B(n714), .Z(n715) );
  XNOR U1264 ( .A(\min_val_reg[6][18] ), .B(n1125), .Z(n714) );
  NAND U1265 ( .A(n609), .B(n974), .Z(n1125) );
  XNOR U1266 ( .A(\min_val_reg[6][18] ), .B(n608), .Z(n609) );
  XOR U1267 ( .A(\min_val_reg[7][18] ), .B(n1126), .Z(n608) );
  NAND U1268 ( .A(n1127), .B(n977), .Z(n1126) );
  XOR U1269 ( .A(\min_val_reg[7][18] ), .B(DB[18]), .Z(n1127) );
  XOR U1270 ( .A(n1128), .B(n1129), .Z(min_val_out[110]) );
  AND U1271 ( .A(n294), .B(n805), .Z(n1128) );
  XOR U1272 ( .A(\min_val_reg[2][17] ), .B(n1129), .Z(n805) );
  XNOR U1273 ( .A(\min_val_reg[3][17] ), .B(n1130), .Z(n1129) );
  NAND U1274 ( .A(n934), .B(n505), .Z(n1130) );
  XOR U1275 ( .A(\min_val_reg[3][17] ), .B(n933), .Z(n934) );
  XNOR U1276 ( .A(\min_val_reg[4][17] ), .B(n1131), .Z(n933) );
  NAND U1277 ( .A(n829), .B(n785), .Z(n1131) );
  XOR U1278 ( .A(\min_val_reg[4][17] ), .B(n828), .Z(n829) );
  XNOR U1279 ( .A(\min_val_reg[5][17] ), .B(n1132), .Z(n828) );
  NAND U1280 ( .A(n718), .B(n674), .Z(n1132) );
  XOR U1281 ( .A(\min_val_reg[5][17] ), .B(n717), .Z(n718) );
  XNOR U1282 ( .A(\min_val_reg[6][17] ), .B(n1133), .Z(n717) );
  NAND U1283 ( .A(n612), .B(n974), .Z(n1133) );
  XNOR U1284 ( .A(\min_val_reg[6][17] ), .B(n611), .Z(n612) );
  XOR U1285 ( .A(\min_val_reg[7][17] ), .B(n1134), .Z(n611) );
  NAND U1286 ( .A(n1135), .B(n977), .Z(n1134) );
  XOR U1287 ( .A(\min_val_reg[7][17] ), .B(DB[17]), .Z(n1135) );
  XOR U1288 ( .A(\min_val_reg[0][10] ), .B(n1136), .Z(min_val_out[10]) );
  AND U1289 ( .A(n290), .B(n481), .Z(n1136) );
  XNOR U1290 ( .A(\min_val_reg[0][10] ), .B(n480), .Z(n481) );
  XOR U1291 ( .A(\min_val_reg[1][10] ), .B(n1137), .Z(n480) );
  NAND U1292 ( .A(n381), .B(n316), .Z(n1137) );
  XOR U1293 ( .A(\min_val_reg[1][10] ), .B(n380), .Z(n381) );
  XNOR U1294 ( .A(\min_val_reg[2][10] ), .B(n1138), .Z(n380) );
  NAND U1295 ( .A(n1139), .B(n294), .Z(n1138) );
  XOR U1296 ( .A(n1140), .B(n1141), .Z(min_val_out[109]) );
  AND U1297 ( .A(n294), .B(n839), .Z(n1140) );
  XOR U1298 ( .A(\min_val_reg[2][16] ), .B(n1141), .Z(n839) );
  XNOR U1299 ( .A(\min_val_reg[3][16] ), .B(n1142), .Z(n1141) );
  NAND U1300 ( .A(n937), .B(n505), .Z(n1142) );
  XOR U1301 ( .A(\min_val_reg[3][16] ), .B(n936), .Z(n937) );
  XNOR U1302 ( .A(\min_val_reg[4][16] ), .B(n1143), .Z(n936) );
  NAND U1303 ( .A(n832), .B(n785), .Z(n1143) );
  XOR U1304 ( .A(\min_val_reg[4][16] ), .B(n831), .Z(n832) );
  XNOR U1305 ( .A(\min_val_reg[5][16] ), .B(n1144), .Z(n831) );
  NAND U1306 ( .A(n721), .B(n674), .Z(n1144) );
  XOR U1307 ( .A(\min_val_reg[5][16] ), .B(n720), .Z(n721) );
  XNOR U1308 ( .A(\min_val_reg[6][16] ), .B(n1145), .Z(n720) );
  NAND U1309 ( .A(n615), .B(n974), .Z(n1145) );
  XNOR U1310 ( .A(\min_val_reg[6][16] ), .B(n614), .Z(n615) );
  XOR U1311 ( .A(\min_val_reg[7][16] ), .B(n1146), .Z(n614) );
  NAND U1312 ( .A(n1147), .B(n977), .Z(n1146) );
  XOR U1313 ( .A(\min_val_reg[7][16] ), .B(DB[16]), .Z(n1147) );
  XOR U1314 ( .A(n1148), .B(n1149), .Z(min_val_out[108]) );
  AND U1315 ( .A(n294), .B(n873), .Z(n1148) );
  XOR U1316 ( .A(\min_val_reg[2][15] ), .B(n1149), .Z(n873) );
  XNOR U1317 ( .A(\min_val_reg[3][15] ), .B(n1150), .Z(n1149) );
  NAND U1318 ( .A(n944), .B(n505), .Z(n1150) );
  XOR U1319 ( .A(\min_val_reg[3][15] ), .B(n943), .Z(n944) );
  XNOR U1320 ( .A(\min_val_reg[4][15] ), .B(n1151), .Z(n943) );
  NAND U1321 ( .A(n835), .B(n785), .Z(n1151) );
  XOR U1322 ( .A(\min_val_reg[4][15] ), .B(n834), .Z(n835) );
  XNOR U1323 ( .A(\min_val_reg[5][15] ), .B(n1152), .Z(n834) );
  NAND U1324 ( .A(n724), .B(n674), .Z(n1152) );
  XOR U1325 ( .A(\min_val_reg[5][15] ), .B(n723), .Z(n724) );
  XNOR U1326 ( .A(\min_val_reg[6][15] ), .B(n1153), .Z(n723) );
  NAND U1327 ( .A(n618), .B(n974), .Z(n1153) );
  XNOR U1328 ( .A(\min_val_reg[6][15] ), .B(n617), .Z(n618) );
  XOR U1329 ( .A(\min_val_reg[7][15] ), .B(n1154), .Z(n617) );
  NAND U1330 ( .A(n1155), .B(n977), .Z(n1154) );
  XOR U1331 ( .A(\min_val_reg[7][15] ), .B(DB[15]), .Z(n1155) );
  XOR U1332 ( .A(n1156), .B(n1157), .Z(min_val_out[107]) );
  AND U1333 ( .A(n294), .B(n907), .Z(n1156) );
  XOR U1334 ( .A(\min_val_reg[2][14] ), .B(n1157), .Z(n907) );
  XNOR U1335 ( .A(\min_val_reg[3][14] ), .B(n1158), .Z(n1157) );
  NAND U1336 ( .A(n947), .B(n505), .Z(n1158) );
  XOR U1337 ( .A(\min_val_reg[3][14] ), .B(n946), .Z(n947) );
  XNOR U1338 ( .A(\min_val_reg[4][14] ), .B(n1159), .Z(n946) );
  NAND U1339 ( .A(n842), .B(n785), .Z(n1159) );
  XOR U1340 ( .A(\min_val_reg[4][14] ), .B(n841), .Z(n842) );
  XNOR U1341 ( .A(\min_val_reg[5][14] ), .B(n1160), .Z(n841) );
  NAND U1342 ( .A(n727), .B(n674), .Z(n1160) );
  XOR U1343 ( .A(\min_val_reg[5][14] ), .B(n726), .Z(n727) );
  XNOR U1344 ( .A(\min_val_reg[6][14] ), .B(n1161), .Z(n726) );
  NAND U1345 ( .A(n621), .B(n974), .Z(n1161) );
  XNOR U1346 ( .A(\min_val_reg[6][14] ), .B(n620), .Z(n621) );
  XOR U1347 ( .A(\min_val_reg[7][14] ), .B(n1162), .Z(n620) );
  NAND U1348 ( .A(n1163), .B(n977), .Z(n1162) );
  XOR U1349 ( .A(\min_val_reg[7][14] ), .B(DB[14]), .Z(n1163) );
  XOR U1350 ( .A(n1164), .B(n1165), .Z(min_val_out[106]) );
  AND U1351 ( .A(n294), .B(n941), .Z(n1164) );
  XOR U1352 ( .A(\min_val_reg[2][13] ), .B(n1165), .Z(n941) );
  XNOR U1353 ( .A(\min_val_reg[3][13] ), .B(n1166), .Z(n1165) );
  NAND U1354 ( .A(n950), .B(n505), .Z(n1166) );
  XOR U1355 ( .A(\min_val_reg[3][13] ), .B(n949), .Z(n950) );
  XNOR U1356 ( .A(\min_val_reg[4][13] ), .B(n1167), .Z(n949) );
  NAND U1357 ( .A(n845), .B(n785), .Z(n1167) );
  XOR U1358 ( .A(\min_val_reg[4][13] ), .B(n844), .Z(n845) );
  XNOR U1359 ( .A(\min_val_reg[5][13] ), .B(n1168), .Z(n844) );
  NAND U1360 ( .A(n739), .B(n674), .Z(n1168) );
  XOR U1361 ( .A(\min_val_reg[5][13] ), .B(n738), .Z(n739) );
  XNOR U1362 ( .A(\min_val_reg[6][13] ), .B(n1169), .Z(n738) );
  NAND U1363 ( .A(n624), .B(n974), .Z(n1169) );
  XNOR U1364 ( .A(\min_val_reg[6][13] ), .B(n623), .Z(n624) );
  XOR U1365 ( .A(\min_val_reg[7][13] ), .B(n1170), .Z(n623) );
  NAND U1366 ( .A(n1171), .B(n977), .Z(n1170) );
  XOR U1367 ( .A(\min_val_reg[7][13] ), .B(DB[13]), .Z(n1171) );
  XOR U1368 ( .A(n1172), .B(n1173), .Z(min_val_out[105]) );
  AND U1369 ( .A(n294), .B(n981), .Z(n1172) );
  XOR U1370 ( .A(\min_val_reg[2][12] ), .B(n1173), .Z(n981) );
  XNOR U1371 ( .A(\min_val_reg[3][12] ), .B(n1174), .Z(n1173) );
  NAND U1372 ( .A(n953), .B(n505), .Z(n1174) );
  XOR U1373 ( .A(\min_val_reg[3][12] ), .B(n952), .Z(n953) );
  XNOR U1374 ( .A(\min_val_reg[4][12] ), .B(n1175), .Z(n952) );
  NAND U1375 ( .A(n848), .B(n785), .Z(n1175) );
  XOR U1376 ( .A(\min_val_reg[4][12] ), .B(n847), .Z(n848) );
  XNOR U1377 ( .A(\min_val_reg[5][12] ), .B(n1176), .Z(n847) );
  NAND U1378 ( .A(n742), .B(n674), .Z(n1176) );
  XOR U1379 ( .A(\min_val_reg[5][12] ), .B(n741), .Z(n742) );
  XNOR U1380 ( .A(\min_val_reg[6][12] ), .B(n1177), .Z(n741) );
  NAND U1381 ( .A(n631), .B(n974), .Z(n1177) );
  XNOR U1382 ( .A(\min_val_reg[6][12] ), .B(n630), .Z(n631) );
  XOR U1383 ( .A(\min_val_reg[7][12] ), .B(n1178), .Z(n630) );
  NAND U1384 ( .A(n1179), .B(n977), .Z(n1178) );
  XOR U1385 ( .A(\min_val_reg[7][12] ), .B(DB[12]), .Z(n1179) );
  XOR U1386 ( .A(n1180), .B(n1181), .Z(min_val_out[104]) );
  AND U1387 ( .A(n294), .B(n1055), .Z(n1180) );
  XOR U1388 ( .A(\min_val_reg[2][11] ), .B(n1181), .Z(n1055) );
  XNOR U1389 ( .A(\min_val_reg[3][11] ), .B(n1182), .Z(n1181) );
  NAND U1390 ( .A(n956), .B(n505), .Z(n1182) );
  XOR U1391 ( .A(\min_val_reg[3][11] ), .B(n955), .Z(n956) );
  XNOR U1392 ( .A(\min_val_reg[4][11] ), .B(n1183), .Z(n955) );
  NAND U1393 ( .A(n851), .B(n785), .Z(n1183) );
  XOR U1394 ( .A(\min_val_reg[4][11] ), .B(n850), .Z(n851) );
  XNOR U1395 ( .A(\min_val_reg[5][11] ), .B(n1184), .Z(n850) );
  NAND U1396 ( .A(n745), .B(n674), .Z(n1184) );
  XOR U1397 ( .A(\min_val_reg[5][11] ), .B(n744), .Z(n745) );
  XNOR U1398 ( .A(\min_val_reg[6][11] ), .B(n1185), .Z(n744) );
  NAND U1399 ( .A(n634), .B(n974), .Z(n1185) );
  XNOR U1400 ( .A(\min_val_reg[6][11] ), .B(n633), .Z(n634) );
  XOR U1401 ( .A(\min_val_reg[7][11] ), .B(n1186), .Z(n633) );
  NAND U1402 ( .A(n1187), .B(n977), .Z(n1186) );
  XOR U1403 ( .A(\min_val_reg[7][11] ), .B(DB[11]), .Z(n1187) );
  XOR U1404 ( .A(n1188), .B(n1189), .Z(min_val_out[103]) );
  AND U1405 ( .A(n294), .B(n1139), .Z(n1188) );
  XOR U1406 ( .A(\min_val_reg[2][10] ), .B(n1189), .Z(n1139) );
  XNOR U1407 ( .A(\min_val_reg[3][10] ), .B(n1190), .Z(n1189) );
  NAND U1408 ( .A(n959), .B(n505), .Z(n1190) );
  XOR U1409 ( .A(\min_val_reg[3][10] ), .B(n958), .Z(n959) );
  XNOR U1410 ( .A(\min_val_reg[4][10] ), .B(n1191), .Z(n958) );
  NAND U1411 ( .A(n854), .B(n785), .Z(n1191) );
  XOR U1412 ( .A(\min_val_reg[4][10] ), .B(n853), .Z(n854) );
  XNOR U1413 ( .A(\min_val_reg[5][10] ), .B(n1192), .Z(n853) );
  NAND U1414 ( .A(n748), .B(n674), .Z(n1192) );
  XOR U1415 ( .A(\min_val_reg[5][10] ), .B(n747), .Z(n748) );
  XNOR U1416 ( .A(\min_val_reg[6][10] ), .B(n1193), .Z(n747) );
  NAND U1417 ( .A(n637), .B(n974), .Z(n1193) );
  XNOR U1418 ( .A(\min_val_reg[6][10] ), .B(n636), .Z(n637) );
  XOR U1419 ( .A(\min_val_reg[7][10] ), .B(n1194), .Z(n636) );
  NAND U1420 ( .A(n1195), .B(n977), .Z(n1194) );
  XOR U1421 ( .A(\min_val_reg[7][10] ), .B(DB[10]), .Z(n1195) );
  XOR U1422 ( .A(n1196), .B(n1197), .Z(min_val_out[102]) );
  AND U1423 ( .A(n294), .B(n486), .Z(n1196) );
  XOR U1424 ( .A(\min_val_reg[2][9] ), .B(n1197), .Z(n486) );
  XNOR U1425 ( .A(\min_val_reg[3][9] ), .B(n1198), .Z(n1197) );
  NAND U1426 ( .A(n962), .B(n505), .Z(n1198) );
  XOR U1427 ( .A(\min_val_reg[3][9] ), .B(n961), .Z(n962) );
  XNOR U1428 ( .A(\min_val_reg[4][9] ), .B(n1199), .Z(n961) );
  NAND U1429 ( .A(n857), .B(n785), .Z(n1199) );
  XOR U1430 ( .A(\min_val_reg[4][9] ), .B(n856), .Z(n857) );
  XNOR U1431 ( .A(\min_val_reg[5][9] ), .B(n1200), .Z(n856) );
  NAND U1432 ( .A(n751), .B(n674), .Z(n1200) );
  XOR U1433 ( .A(\min_val_reg[5][9] ), .B(n750), .Z(n751) );
  XNOR U1434 ( .A(\min_val_reg[6][9] ), .B(n1201), .Z(n750) );
  NAND U1435 ( .A(n640), .B(n974), .Z(n1201) );
  XNOR U1436 ( .A(\min_val_reg[6][9] ), .B(n639), .Z(n640) );
  XOR U1437 ( .A(\min_val_reg[7][9] ), .B(n1202), .Z(n639) );
  NAND U1438 ( .A(n1203), .B(n977), .Z(n1202) );
  XOR U1439 ( .A(\min_val_reg[7][9] ), .B(DB[9]), .Z(n1203) );
  XOR U1440 ( .A(n1204), .B(n1205), .Z(min_val_out[101]) );
  AND U1441 ( .A(n294), .B(n493), .Z(n1204) );
  XOR U1442 ( .A(\min_val_reg[2][8] ), .B(n1205), .Z(n493) );
  XNOR U1443 ( .A(\min_val_reg[3][8] ), .B(n1206), .Z(n1205) );
  NAND U1444 ( .A(n965), .B(n505), .Z(n1206) );
  XOR U1445 ( .A(\min_val_reg[3][8] ), .B(n964), .Z(n965) );
  XNOR U1446 ( .A(\min_val_reg[4][8] ), .B(n1207), .Z(n964) );
  NAND U1447 ( .A(n860), .B(n785), .Z(n1207) );
  XOR U1448 ( .A(\min_val_reg[4][8] ), .B(n859), .Z(n860) );
  XNOR U1449 ( .A(\min_val_reg[5][8] ), .B(n1208), .Z(n859) );
  NAND U1450 ( .A(n754), .B(n674), .Z(n1208) );
  XOR U1451 ( .A(\min_val_reg[5][8] ), .B(n753), .Z(n754) );
  XNOR U1452 ( .A(\min_val_reg[6][8] ), .B(n1209), .Z(n753) );
  NAND U1453 ( .A(n643), .B(n974), .Z(n1209) );
  XNOR U1454 ( .A(\min_val_reg[6][8] ), .B(n642), .Z(n643) );
  XOR U1455 ( .A(\min_val_reg[7][8] ), .B(n1210), .Z(n642) );
  NAND U1456 ( .A(n1211), .B(n977), .Z(n1210) );
  XOR U1457 ( .A(\min_val_reg[7][8] ), .B(DB[8]), .Z(n1211) );
  XOR U1458 ( .A(n1212), .B(n1213), .Z(min_val_out[100]) );
  AND U1459 ( .A(n294), .B(n498), .Z(n1212) );
  XOR U1460 ( .A(\min_val_reg[2][7] ), .B(n1213), .Z(n498) );
  XNOR U1461 ( .A(\min_val_reg[3][7] ), .B(n1214), .Z(n1213) );
  NAND U1462 ( .A(n968), .B(n505), .Z(n1214) );
  XOR U1463 ( .A(\min_val_reg[3][7] ), .B(n967), .Z(n968) );
  XNOR U1464 ( .A(\min_val_reg[4][7] ), .B(n1215), .Z(n967) );
  NAND U1465 ( .A(n863), .B(n785), .Z(n1215) );
  XOR U1466 ( .A(\min_val_reg[4][7] ), .B(n862), .Z(n863) );
  XNOR U1467 ( .A(\min_val_reg[5][7] ), .B(n1216), .Z(n862) );
  NAND U1468 ( .A(n757), .B(n674), .Z(n1216) );
  XOR U1469 ( .A(\min_val_reg[5][7] ), .B(n756), .Z(n757) );
  XNOR U1470 ( .A(\min_val_reg[6][7] ), .B(n1217), .Z(n756) );
  NAND U1471 ( .A(n646), .B(n974), .Z(n1217) );
  XNOR U1472 ( .A(\min_val_reg[6][7] ), .B(n645), .Z(n646) );
  XOR U1473 ( .A(\min_val_reg[7][7] ), .B(n1218), .Z(n645) );
  NAND U1474 ( .A(n1219), .B(n977), .Z(n1218) );
  XOR U1475 ( .A(\min_val_reg[7][7] ), .B(DB[7]), .Z(n1219) );
  XOR U1476 ( .A(\min_val_reg[0][0] ), .B(n1220), .Z(min_val_out[0]) );
  AND U1477 ( .A(n290), .B(n532), .Z(n1220) );
  XNOR U1478 ( .A(\min_val_reg[0][0] ), .B(n531), .Z(n532) );
  XOR U1479 ( .A(\min_val_reg[1][0] ), .B(n1221), .Z(n531) );
  NAND U1480 ( .A(n413), .B(n316), .Z(n1221) );
  XNOR U1481 ( .A(\min_val_reg[1][0] ), .B(n412), .Z(n413) );
  XOR U1482 ( .A(\min_val_reg[2][0] ), .B(n1222), .Z(n412) );
  NAND U1483 ( .A(n313), .B(n294), .Z(n1222) );
  XOR U1484 ( .A(\min_val_reg[2][0] ), .B(n312), .Z(n313) );
  XNOR U1485 ( .A(\min_val_reg[3][0] ), .B(n1223), .Z(n312) );
  NAND U1486 ( .A(n1019), .B(n505), .Z(n1223) );
  XOR U1487 ( .A(\min_val_reg[3][0] ), .B(n1018), .Z(n1019) );
  XNOR U1488 ( .A(\min_val_reg[4][0] ), .B(n1224), .Z(n1018) );
  NAND U1489 ( .A(n888), .B(n785), .Z(n1224) );
  XOR U1490 ( .A(\min_val_reg[4][0] ), .B(n887), .Z(n888) );
  XNOR U1491 ( .A(\min_val_reg[5][0] ), .B(n1225), .Z(n887) );
  NAND U1492 ( .A(n782), .B(n674), .Z(n1225) );
  XOR U1493 ( .A(\min_val_reg[5][0] ), .B(n781), .Z(n782) );
  XNOR U1494 ( .A(\min_val_reg[6][0] ), .B(n1226), .Z(n781) );
  NAND U1495 ( .A(n671), .B(n974), .Z(n1226) );
  XNOR U1496 ( .A(\min_val_reg[6][0] ), .B(n670), .Z(n671) );
  XOR U1497 ( .A(\min_val_reg[7][0] ), .B(n1227), .Z(n670) );
  NAND U1498 ( .A(n1228), .B(n977), .Z(n1227) );
  XOR U1499 ( .A(\min_val_reg[7][0] ), .B(DB[0]), .Z(n1228) );
  XOR U1500 ( .A(n1229), .B(n1230), .Z(\min_dist[7][4] ) );
  AND U1501 ( .A(n568), .B(n1231), .Z(n1229) );
  XOR U1502 ( .A(\min_dist_reg[6][4] ), .B(n1230), .Z(n1231) );
  XOR U1503 ( .A(n1232), .B(n1233), .Z(\min_dist[7][3] ) );
  AND U1504 ( .A(n568), .B(n1234), .Z(n1232) );
  XNOR U1505 ( .A(\min_dist_reg[6][3] ), .B(n1235), .Z(n1234) );
  XOR U1506 ( .A(n1236), .B(n1237), .Z(\min_dist[7][2] ) );
  AND U1507 ( .A(n568), .B(n1238), .Z(n1236) );
  XNOR U1508 ( .A(\min_dist_reg[6][2] ), .B(n1239), .Z(n1238) );
  XOR U1509 ( .A(n1240), .B(n1241), .Z(\min_dist[7][1] ) );
  AND U1510 ( .A(n568), .B(n1242), .Z(n1240) );
  XNOR U1511 ( .A(\min_dist_reg[6][1] ), .B(n1243), .Z(n1242) );
  XOR U1512 ( .A(n1244), .B(n1245), .Z(\min_dist[7][0] ) );
  AND U1513 ( .A(n568), .B(n1246), .Z(n1244) );
  XOR U1514 ( .A(n1247), .B(n1248), .Z(n568) );
  AND U1515 ( .A(n1249), .B(n1250), .Z(n1247) );
  XNOR U1516 ( .A(n1230), .B(n1248), .Z(n1250) );
  XNOR U1517 ( .A(n1251), .B(n1248), .Z(n1249) );
  XOR U1518 ( .A(n1252), .B(n1253), .Z(n1248) );
  AND U1519 ( .A(n1254), .B(n1255), .Z(n1252) );
  XNOR U1520 ( .A(n1235), .B(n1256), .Z(n1255) );
  IV U1521 ( .A(n1253), .Z(n1256) );
  IV U1522 ( .A(n1233), .Z(n1235) );
  XOR U1523 ( .A(n1257), .B(n1258), .Z(\min_dist[6][4] ) );
  AND U1524 ( .A(n674), .B(n1259), .Z(n1257) );
  XOR U1525 ( .A(\min_dist_reg[5][4] ), .B(n1258), .Z(n1259) );
  XOR U1526 ( .A(n1260), .B(n1261), .Z(\min_dist[6][3] ) );
  AND U1527 ( .A(n674), .B(n1262), .Z(n1260) );
  XOR U1528 ( .A(\min_dist_reg[5][3] ), .B(n1261), .Z(n1262) );
  XOR U1529 ( .A(n1263), .B(n1264), .Z(\min_dist[6][2] ) );
  AND U1530 ( .A(n674), .B(n1265), .Z(n1263) );
  XOR U1531 ( .A(\min_dist_reg[5][2] ), .B(n1264), .Z(n1265) );
  XOR U1532 ( .A(n1266), .B(n1267), .Z(\min_dist[6][1] ) );
  AND U1533 ( .A(n674), .B(n1268), .Z(n1266) );
  XOR U1534 ( .A(\min_dist_reg[5][1] ), .B(n1267), .Z(n1268) );
  XOR U1535 ( .A(n1269), .B(n1270), .Z(\min_dist[6][0] ) );
  AND U1536 ( .A(n674), .B(n1271), .Z(n1269) );
  XOR U1537 ( .A(n1272), .B(n1273), .Z(\min_dist[5][4] ) );
  AND U1538 ( .A(n785), .B(n1274), .Z(n1272) );
  XOR U1539 ( .A(\min_dist_reg[4][4] ), .B(n1273), .Z(n1274) );
  XOR U1540 ( .A(n1275), .B(n1276), .Z(\min_dist[5][3] ) );
  AND U1541 ( .A(n785), .B(n1277), .Z(n1275) );
  XOR U1542 ( .A(\min_dist_reg[4][3] ), .B(n1276), .Z(n1277) );
  XOR U1543 ( .A(n1278), .B(n1279), .Z(\min_dist[5][2] ) );
  AND U1544 ( .A(n785), .B(n1280), .Z(n1278) );
  XOR U1545 ( .A(\min_dist_reg[4][2] ), .B(n1279), .Z(n1280) );
  XOR U1546 ( .A(n1281), .B(n1282), .Z(\min_dist[5][1] ) );
  AND U1547 ( .A(n785), .B(n1283), .Z(n1281) );
  XOR U1548 ( .A(\min_dist_reg[4][1] ), .B(n1282), .Z(n1283) );
  XOR U1549 ( .A(n1284), .B(n1285), .Z(\min_dist[5][0] ) );
  AND U1550 ( .A(n785), .B(n1286), .Z(n1284) );
  XOR U1551 ( .A(n1287), .B(n1288), .Z(\min_dist[4][4] ) );
  AND U1552 ( .A(n505), .B(n1289), .Z(n1287) );
  XOR U1553 ( .A(\min_dist_reg[3][4] ), .B(n1288), .Z(n1289) );
  XOR U1554 ( .A(n1290), .B(n1291), .Z(\min_dist[4][3] ) );
  AND U1555 ( .A(n505), .B(n1292), .Z(n1290) );
  XOR U1556 ( .A(\min_dist_reg[3][3] ), .B(n1291), .Z(n1292) );
  XOR U1557 ( .A(n1293), .B(n1294), .Z(\min_dist[4][2] ) );
  AND U1558 ( .A(n505), .B(n1295), .Z(n1293) );
  XOR U1559 ( .A(\min_dist_reg[3][2] ), .B(n1294), .Z(n1295) );
  XOR U1560 ( .A(n1296), .B(n1297), .Z(\min_dist[4][1] ) );
  AND U1561 ( .A(n505), .B(n1298), .Z(n1296) );
  XOR U1562 ( .A(\min_dist_reg[3][1] ), .B(n1297), .Z(n1298) );
  XOR U1563 ( .A(n1299), .B(n1300), .Z(\min_dist[4][0] ) );
  AND U1564 ( .A(n505), .B(n1301), .Z(n1299) );
  XOR U1565 ( .A(n1302), .B(n1303), .Z(\min_dist[3][4] ) );
  AND U1566 ( .A(n294), .B(n1304), .Z(n1302) );
  XOR U1567 ( .A(\min_dist_reg[2][4] ), .B(n1303), .Z(n1304) );
  XOR U1568 ( .A(n1305), .B(n1306), .Z(\min_dist[3][3] ) );
  AND U1569 ( .A(n294), .B(n1307), .Z(n1305) );
  XOR U1570 ( .A(\min_dist_reg[2][3] ), .B(n1306), .Z(n1307) );
  XOR U1571 ( .A(n1308), .B(n1309), .Z(\min_dist[3][2] ) );
  AND U1572 ( .A(n294), .B(n1310), .Z(n1308) );
  XOR U1573 ( .A(\min_dist_reg[2][2] ), .B(n1309), .Z(n1310) );
  XOR U1574 ( .A(n1311), .B(n1312), .Z(\min_dist[3][1] ) );
  AND U1575 ( .A(n294), .B(n1313), .Z(n1311) );
  XOR U1576 ( .A(\min_dist_reg[2][1] ), .B(n1312), .Z(n1313) );
  XOR U1577 ( .A(n1314), .B(n1315), .Z(\min_dist[3][0] ) );
  AND U1578 ( .A(n294), .B(n1316), .Z(n1314) );
  XOR U1579 ( .A(n1317), .B(n1318), .Z(\min_dist[2][4] ) );
  AND U1580 ( .A(n316), .B(n1319), .Z(n1317) );
  XOR U1581 ( .A(\min_dist_reg[1][4] ), .B(n1318), .Z(n1319) );
  XOR U1582 ( .A(n1320), .B(n1321), .Z(\min_dist[2][3] ) );
  AND U1583 ( .A(n316), .B(n1322), .Z(n1320) );
  XOR U1584 ( .A(\min_dist_reg[1][3] ), .B(n1321), .Z(n1322) );
  XOR U1585 ( .A(n1323), .B(n1324), .Z(\min_dist[2][2] ) );
  AND U1586 ( .A(n316), .B(n1325), .Z(n1323) );
  XOR U1587 ( .A(\min_dist_reg[1][2] ), .B(n1324), .Z(n1325) );
  XOR U1588 ( .A(n1326), .B(n1327), .Z(\min_dist[2][1] ) );
  AND U1589 ( .A(n316), .B(n1328), .Z(n1326) );
  XOR U1590 ( .A(\min_dist_reg[1][1] ), .B(n1327), .Z(n1328) );
  XOR U1591 ( .A(n1329), .B(n1330), .Z(\min_dist[2][0] ) );
  AND U1592 ( .A(n316), .B(n1331), .Z(n1329) );
  XOR U1593 ( .A(n1332), .B(n1333), .Z(\min_dist[1][4] ) );
  AND U1594 ( .A(n416), .B(n1334), .Z(n1332) );
  XOR U1595 ( .A(\min_dist_reg[0][4] ), .B(n1333), .Z(n1334) );
  XOR U1596 ( .A(n1335), .B(n1336), .Z(\min_dist[1][3] ) );
  AND U1597 ( .A(n416), .B(n1337), .Z(n1335) );
  XOR U1598 ( .A(n1338), .B(n1339), .Z(\min_dist[1][2] ) );
  AND U1599 ( .A(n416), .B(n1340), .Z(n1338) );
  XOR U1600 ( .A(n1341), .B(n1342), .Z(\min_dist[1][1] ) );
  AND U1601 ( .A(n416), .B(n1343), .Z(n1341) );
  XNOR U1602 ( .A(n1344), .B(n1345), .Z(\min_dist[1][0] ) );
  AND U1603 ( .A(n416), .B(n1346), .Z(n1344) );
  XNOR U1604 ( .A(\min_dist_reg[0][0] ), .B(n1345), .Z(n1346) );
  XNOR U1605 ( .A(n1347), .B(n1348), .Z(n416) );
  AND U1606 ( .A(n1349), .B(n1350), .Z(n1347) );
  XOR U1607 ( .A(n1333), .B(n1348), .Z(n1350) );
  XNOR U1608 ( .A(\min_dist_reg[0][4] ), .B(n1348), .Z(n1349) );
  XOR U1609 ( .A(n1351), .B(n1352), .Z(n1348) );
  AND U1610 ( .A(n1353), .B(n1354), .Z(n1351) );
  XNOR U1611 ( .A(n1336), .B(n1355), .Z(n1354) );
  XNOR U1612 ( .A(\min_dist_reg[0][3] ), .B(n1352), .Z(n1353) );
  IV U1613 ( .A(n1355), .Z(n1352) );
  XOR U1614 ( .A(n1356), .B(n1357), .Z(n1355) );
  AND U1615 ( .A(n1358), .B(n1359), .Z(n1356) );
  XNOR U1616 ( .A(n1339), .B(n1357), .Z(n1359) );
  XOR U1617 ( .A(\min_dist_reg[0][2] ), .B(n1357), .Z(n1358) );
  XOR U1618 ( .A(n1360), .B(n1361), .Z(n1357) );
  NAND U1619 ( .A(n1362), .B(n1363), .Z(n1361) );
  XOR U1620 ( .A(n1360), .B(n1342), .Z(n1363) );
  XNOR U1621 ( .A(\min_dist_reg[0][1] ), .B(n1360), .Z(n1362) );
  NOR U1622 ( .A(n1345), .B(\min_dist_reg[0][0] ), .Z(n1360) );
  AND U1623 ( .A(\min_dist_reg[0][4] ), .B(n1364), .Z(\local_min_dist[0][4] )
         );
  NANDN U1624 ( .A(n1333), .B(n290), .Z(n1364) );
  XOR U1625 ( .A(\min_dist_reg[0][3] ), .B(n1365), .Z(\local_min_dist[0][3] )
         );
  AND U1626 ( .A(n290), .B(n1337), .Z(n1365) );
  XOR U1627 ( .A(\min_dist_reg[0][3] ), .B(n1336), .Z(n1337) );
  XOR U1628 ( .A(\min_dist_reg[0][2] ), .B(n1366), .Z(\local_min_dist[0][2] )
         );
  AND U1629 ( .A(n290), .B(n1340), .Z(n1366) );
  XOR U1630 ( .A(\min_dist_reg[0][2] ), .B(n1339), .Z(n1340) );
  XOR U1631 ( .A(\min_dist_reg[0][1] ), .B(n1367), .Z(\local_min_dist[0][1] )
         );
  AND U1632 ( .A(n290), .B(n1343), .Z(n1367) );
  XOR U1633 ( .A(\min_dist_reg[0][1] ), .B(n1342), .Z(n1343) );
  XOR U1634 ( .A(\min_dist_reg[0][0] ), .B(n1368), .Z(\local_min_dist[0][0] )
         );
  AND U1635 ( .A(n290), .B(n1369), .Z(n1368) );
  XOR U1636 ( .A(\min_dist_reg[0][0] ), .B(n1370), .Z(n1369) );
  XNOR U1637 ( .A(n1371), .B(n1372), .Z(n290) );
  AND U1638 ( .A(n1373), .B(n1374), .Z(n1371) );
  XOR U1639 ( .A(n1333), .B(n1372), .Z(n1374) );
  AND U1640 ( .A(n1375), .B(\min_dist_reg[1][4] ), .Z(n1333) );
  NANDN U1641 ( .A(n1318), .B(n316), .Z(n1375) );
  XNOR U1642 ( .A(\min_dist_reg[0][4] ), .B(n1372), .Z(n1373) );
  XOR U1643 ( .A(n1376), .B(n1377), .Z(n1372) );
  AND U1644 ( .A(n1378), .B(n1379), .Z(n1376) );
  XNOR U1645 ( .A(n1380), .B(n1336), .Z(n1379) );
  XNOR U1646 ( .A(\min_dist_reg[1][3] ), .B(n1381), .Z(n1336) );
  NAND U1647 ( .A(n1382), .B(n316), .Z(n1381) );
  XNOR U1648 ( .A(n1383), .B(n1321), .Z(n1382) );
  XNOR U1649 ( .A(\min_dist_reg[0][3] ), .B(n1377), .Z(n1378) );
  IV U1650 ( .A(n1380), .Z(n1377) );
  XOR U1651 ( .A(n1384), .B(n1385), .Z(n1380) );
  AND U1652 ( .A(n1386), .B(n1387), .Z(n1384) );
  XNOR U1653 ( .A(n1385), .B(n1339), .Z(n1387) );
  XNOR U1654 ( .A(\min_dist_reg[1][2] ), .B(n1388), .Z(n1339) );
  NAND U1655 ( .A(n1389), .B(n316), .Z(n1388) );
  XNOR U1656 ( .A(n1390), .B(n1324), .Z(n1389) );
  XOR U1657 ( .A(\min_dist_reg[0][2] ), .B(n1385), .Z(n1386) );
  XOR U1658 ( .A(n1391), .B(n1392), .Z(n1385) );
  NAND U1659 ( .A(n1393), .B(n1394), .Z(n1392) );
  XOR U1660 ( .A(n1391), .B(n1342), .Z(n1394) );
  XNOR U1661 ( .A(\min_dist_reg[1][1] ), .B(n1395), .Z(n1342) );
  NAND U1662 ( .A(n1396), .B(n316), .Z(n1395) );
  XNOR U1663 ( .A(n1397), .B(n1327), .Z(n1396) );
  XNOR U1664 ( .A(\min_dist_reg[0][1] ), .B(n1391), .Z(n1393) );
  ANDN U1665 ( .B(n1370), .A(\min_dist_reg[0][0] ), .Z(n1391) );
  IV U1666 ( .A(n1345), .Z(n1370) );
  XOR U1667 ( .A(\min_dist_reg[1][0] ), .B(n1398), .Z(n1345) );
  NAND U1668 ( .A(n1331), .B(n316), .Z(n1398) );
  XOR U1669 ( .A(n1399), .B(n1400), .Z(n316) );
  AND U1670 ( .A(n1401), .B(n1402), .Z(n1399) );
  XNOR U1671 ( .A(n1318), .B(n1400), .Z(n1402) );
  AND U1672 ( .A(n1403), .B(\min_dist_reg[2][4] ), .Z(n1318) );
  NANDN U1673 ( .A(n1303), .B(n294), .Z(n1403) );
  XNOR U1674 ( .A(n1404), .B(n1400), .Z(n1401) );
  XOR U1675 ( .A(n1405), .B(n1406), .Z(n1400) );
  AND U1676 ( .A(n1407), .B(n1408), .Z(n1405) );
  XNOR U1677 ( .A(n1321), .B(n1406), .Z(n1408) );
  XNOR U1678 ( .A(\min_dist_reg[2][3] ), .B(n1409), .Z(n1321) );
  NAND U1679 ( .A(n1410), .B(n294), .Z(n1409) );
  XNOR U1680 ( .A(n1411), .B(n1306), .Z(n1410) );
  XNOR U1681 ( .A(n1383), .B(n1406), .Z(n1407) );
  XOR U1682 ( .A(n1412), .B(n1413), .Z(n1406) );
  AND U1683 ( .A(n1414), .B(n1415), .Z(n1412) );
  XNOR U1684 ( .A(n1324), .B(n1413), .Z(n1415) );
  XNOR U1685 ( .A(\min_dist_reg[2][2] ), .B(n1416), .Z(n1324) );
  NAND U1686 ( .A(n1417), .B(n294), .Z(n1416) );
  XNOR U1687 ( .A(n1418), .B(n1309), .Z(n1417) );
  XNOR U1688 ( .A(n1390), .B(n1413), .Z(n1414) );
  XOR U1689 ( .A(n1419), .B(n1420), .Z(n1413) );
  NAND U1690 ( .A(n1421), .B(n1422), .Z(n1420) );
  XOR U1691 ( .A(n1419), .B(n1327), .Z(n1422) );
  XNOR U1692 ( .A(\min_dist_reg[2][1] ), .B(n1423), .Z(n1327) );
  NAND U1693 ( .A(n1424), .B(n294), .Z(n1423) );
  XNOR U1694 ( .A(n1425), .B(n1312), .Z(n1424) );
  XOR U1695 ( .A(n1397), .B(n1419), .Z(n1421) );
  IV U1696 ( .A(\min_dist_reg[1][1] ), .Z(n1397) );
  AND U1697 ( .A(n1330), .B(n1426), .Z(n1419) );
  IV U1698 ( .A(\min_dist_reg[1][2] ), .Z(n1390) );
  IV U1699 ( .A(\min_dist_reg[1][3] ), .Z(n1383) );
  IV U1700 ( .A(\min_dist_reg[1][4] ), .Z(n1404) );
  XNOR U1701 ( .A(n1426), .B(n1330), .Z(n1331) );
  XNOR U1702 ( .A(\min_dist_reg[2][0] ), .B(n1427), .Z(n1330) );
  NAND U1703 ( .A(n1316), .B(n294), .Z(n1427) );
  XOR U1704 ( .A(n1428), .B(n1429), .Z(n294) );
  AND U1705 ( .A(n1430), .B(n1431), .Z(n1428) );
  XNOR U1706 ( .A(n1303), .B(n1429), .Z(n1431) );
  AND U1707 ( .A(n1432), .B(\min_dist_reg[3][4] ), .Z(n1303) );
  NANDN U1708 ( .A(n1288), .B(n505), .Z(n1432) );
  XNOR U1709 ( .A(n1433), .B(n1429), .Z(n1430) );
  XOR U1710 ( .A(n1434), .B(n1435), .Z(n1429) );
  AND U1711 ( .A(n1436), .B(n1437), .Z(n1434) );
  XNOR U1712 ( .A(n1306), .B(n1435), .Z(n1437) );
  XNOR U1713 ( .A(\min_dist_reg[3][3] ), .B(n1438), .Z(n1306) );
  NAND U1714 ( .A(n1439), .B(n505), .Z(n1438) );
  XNOR U1715 ( .A(n1440), .B(n1291), .Z(n1439) );
  XNOR U1716 ( .A(n1411), .B(n1435), .Z(n1436) );
  XOR U1717 ( .A(n1441), .B(n1442), .Z(n1435) );
  AND U1718 ( .A(n1443), .B(n1444), .Z(n1441) );
  XNOR U1719 ( .A(n1309), .B(n1442), .Z(n1444) );
  XNOR U1720 ( .A(\min_dist_reg[3][2] ), .B(n1445), .Z(n1309) );
  NAND U1721 ( .A(n1446), .B(n505), .Z(n1445) );
  XNOR U1722 ( .A(n1447), .B(n1294), .Z(n1446) );
  XNOR U1723 ( .A(n1418), .B(n1442), .Z(n1443) );
  XOR U1724 ( .A(n1448), .B(n1449), .Z(n1442) );
  NAND U1725 ( .A(n1450), .B(n1451), .Z(n1449) );
  XOR U1726 ( .A(n1448), .B(n1312), .Z(n1451) );
  XNOR U1727 ( .A(\min_dist_reg[3][1] ), .B(n1452), .Z(n1312) );
  NAND U1728 ( .A(n1453), .B(n505), .Z(n1452) );
  XNOR U1729 ( .A(n1454), .B(n1297), .Z(n1453) );
  XOR U1730 ( .A(n1425), .B(n1448), .Z(n1450) );
  IV U1731 ( .A(\min_dist_reg[2][1] ), .Z(n1425) );
  ANDN U1732 ( .B(n1315), .A(\min_dist_reg[2][0] ), .Z(n1448) );
  IV U1733 ( .A(\min_dist_reg[2][2] ), .Z(n1418) );
  IV U1734 ( .A(\min_dist_reg[2][3] ), .Z(n1411) );
  IV U1735 ( .A(\min_dist_reg[2][4] ), .Z(n1433) );
  XOR U1736 ( .A(\min_dist_reg[2][0] ), .B(n1315), .Z(n1316) );
  XNOR U1737 ( .A(\min_dist_reg[3][0] ), .B(n1455), .Z(n1315) );
  NAND U1738 ( .A(n1301), .B(n505), .Z(n1455) );
  XOR U1739 ( .A(n1456), .B(n1457), .Z(n505) );
  AND U1740 ( .A(n1458), .B(n1459), .Z(n1456) );
  XNOR U1741 ( .A(n1288), .B(n1457), .Z(n1459) );
  AND U1742 ( .A(n1460), .B(\min_dist_reg[4][4] ), .Z(n1288) );
  NANDN U1743 ( .A(n1273), .B(n785), .Z(n1460) );
  XNOR U1744 ( .A(n1461), .B(n1457), .Z(n1458) );
  XOR U1745 ( .A(n1462), .B(n1463), .Z(n1457) );
  AND U1746 ( .A(n1464), .B(n1465), .Z(n1462) );
  XNOR U1747 ( .A(n1291), .B(n1463), .Z(n1465) );
  XNOR U1748 ( .A(\min_dist_reg[4][3] ), .B(n1466), .Z(n1291) );
  NAND U1749 ( .A(n1467), .B(n785), .Z(n1466) );
  XNOR U1750 ( .A(n1468), .B(n1276), .Z(n1467) );
  XNOR U1751 ( .A(n1440), .B(n1463), .Z(n1464) );
  XOR U1752 ( .A(n1469), .B(n1470), .Z(n1463) );
  AND U1753 ( .A(n1471), .B(n1472), .Z(n1469) );
  XNOR U1754 ( .A(n1294), .B(n1470), .Z(n1472) );
  XNOR U1755 ( .A(\min_dist_reg[4][2] ), .B(n1473), .Z(n1294) );
  NAND U1756 ( .A(n1474), .B(n785), .Z(n1473) );
  XNOR U1757 ( .A(n1475), .B(n1279), .Z(n1474) );
  XNOR U1758 ( .A(n1447), .B(n1470), .Z(n1471) );
  XOR U1759 ( .A(n1476), .B(n1477), .Z(n1470) );
  NAND U1760 ( .A(n1478), .B(n1479), .Z(n1477) );
  XOR U1761 ( .A(n1476), .B(n1297), .Z(n1479) );
  XNOR U1762 ( .A(\min_dist_reg[4][1] ), .B(n1480), .Z(n1297) );
  NAND U1763 ( .A(n1481), .B(n785), .Z(n1480) );
  XNOR U1764 ( .A(n1482), .B(n1282), .Z(n1481) );
  XOR U1765 ( .A(n1454), .B(n1476), .Z(n1478) );
  IV U1766 ( .A(\min_dist_reg[3][1] ), .Z(n1454) );
  ANDN U1767 ( .B(n1300), .A(\min_dist_reg[3][0] ), .Z(n1476) );
  IV U1768 ( .A(\min_dist_reg[3][2] ), .Z(n1447) );
  IV U1769 ( .A(\min_dist_reg[3][3] ), .Z(n1440) );
  IV U1770 ( .A(\min_dist_reg[3][4] ), .Z(n1461) );
  XOR U1771 ( .A(\min_dist_reg[3][0] ), .B(n1300), .Z(n1301) );
  XNOR U1772 ( .A(\min_dist_reg[4][0] ), .B(n1483), .Z(n1300) );
  NAND U1773 ( .A(n1286), .B(n785), .Z(n1483) );
  XOR U1774 ( .A(n1484), .B(n1485), .Z(n785) );
  AND U1775 ( .A(n1486), .B(n1487), .Z(n1484) );
  XNOR U1776 ( .A(n1273), .B(n1485), .Z(n1487) );
  AND U1777 ( .A(n1488), .B(\min_dist_reg[5][4] ), .Z(n1273) );
  NANDN U1778 ( .A(n1258), .B(n674), .Z(n1488) );
  XNOR U1779 ( .A(n1489), .B(n1485), .Z(n1486) );
  XOR U1780 ( .A(n1490), .B(n1491), .Z(n1485) );
  AND U1781 ( .A(n1492), .B(n1493), .Z(n1490) );
  XNOR U1782 ( .A(n1276), .B(n1491), .Z(n1493) );
  XNOR U1783 ( .A(\min_dist_reg[5][3] ), .B(n1494), .Z(n1276) );
  NAND U1784 ( .A(n1495), .B(n674), .Z(n1494) );
  XNOR U1785 ( .A(n1496), .B(n1261), .Z(n1495) );
  XNOR U1786 ( .A(n1468), .B(n1491), .Z(n1492) );
  XOR U1787 ( .A(n1497), .B(n1498), .Z(n1491) );
  AND U1788 ( .A(n1499), .B(n1500), .Z(n1497) );
  XNOR U1789 ( .A(n1279), .B(n1498), .Z(n1500) );
  XNOR U1790 ( .A(\min_dist_reg[5][2] ), .B(n1501), .Z(n1279) );
  NAND U1791 ( .A(n1502), .B(n674), .Z(n1501) );
  XNOR U1792 ( .A(n1503), .B(n1264), .Z(n1502) );
  XNOR U1793 ( .A(n1475), .B(n1498), .Z(n1499) );
  XOR U1794 ( .A(n1504), .B(n1505), .Z(n1498) );
  NAND U1795 ( .A(n1506), .B(n1507), .Z(n1505) );
  XOR U1796 ( .A(n1504), .B(n1282), .Z(n1507) );
  XNOR U1797 ( .A(\min_dist_reg[5][1] ), .B(n1508), .Z(n1282) );
  NAND U1798 ( .A(n1509), .B(n674), .Z(n1508) );
  XNOR U1799 ( .A(n1510), .B(n1267), .Z(n1509) );
  XOR U1800 ( .A(n1482), .B(n1504), .Z(n1506) );
  IV U1801 ( .A(\min_dist_reg[4][1] ), .Z(n1482) );
  ANDN U1802 ( .B(n1285), .A(\min_dist_reg[4][0] ), .Z(n1504) );
  IV U1803 ( .A(\min_dist_reg[4][2] ), .Z(n1475) );
  IV U1804 ( .A(\min_dist_reg[4][3] ), .Z(n1468) );
  IV U1805 ( .A(\min_dist_reg[4][4] ), .Z(n1489) );
  XOR U1806 ( .A(\min_dist_reg[4][0] ), .B(n1285), .Z(n1286) );
  XNOR U1807 ( .A(\min_dist_reg[5][0] ), .B(n1511), .Z(n1285) );
  NAND U1808 ( .A(n1271), .B(n674), .Z(n1511) );
  XOR U1809 ( .A(n1512), .B(n1513), .Z(n674) );
  AND U1810 ( .A(n1514), .B(n1515), .Z(n1512) );
  XNOR U1811 ( .A(n1258), .B(n1513), .Z(n1515) );
  AND U1812 ( .A(n1516), .B(\min_dist_reg[6][4] ), .Z(n1258) );
  NANDN U1813 ( .A(n1230), .B(n974), .Z(n1516) );
  XNOR U1814 ( .A(n1517), .B(n1513), .Z(n1514) );
  XOR U1815 ( .A(n1518), .B(n1519), .Z(n1513) );
  AND U1816 ( .A(n1520), .B(n1521), .Z(n1518) );
  XNOR U1817 ( .A(n1261), .B(n1519), .Z(n1521) );
  XNOR U1818 ( .A(\min_dist_reg[6][3] ), .B(n1522), .Z(n1261) );
  NAND U1819 ( .A(n1523), .B(n974), .Z(n1522) );
  XNOR U1820 ( .A(n1524), .B(n1233), .Z(n1523) );
  XNOR U1821 ( .A(n1496), .B(n1519), .Z(n1520) );
  XOR U1822 ( .A(n1525), .B(n1526), .Z(n1519) );
  AND U1823 ( .A(n1527), .B(n1528), .Z(n1525) );
  XNOR U1824 ( .A(n1264), .B(n1526), .Z(n1528) );
  XNOR U1825 ( .A(\min_dist_reg[6][2] ), .B(n1529), .Z(n1264) );
  NAND U1826 ( .A(n1530), .B(n974), .Z(n1529) );
  XNOR U1827 ( .A(n1531), .B(n1237), .Z(n1530) );
  XNOR U1828 ( .A(n1503), .B(n1526), .Z(n1527) );
  XOR U1829 ( .A(n1532), .B(n1533), .Z(n1526) );
  NAND U1830 ( .A(n1534), .B(n1535), .Z(n1533) );
  XOR U1831 ( .A(n1532), .B(n1267), .Z(n1535) );
  XNOR U1832 ( .A(\min_dist_reg[6][1] ), .B(n1536), .Z(n1267) );
  NAND U1833 ( .A(n1537), .B(n974), .Z(n1536) );
  XNOR U1834 ( .A(n1538), .B(n1241), .Z(n1537) );
  XOR U1835 ( .A(n1510), .B(n1532), .Z(n1534) );
  IV U1836 ( .A(\min_dist_reg[5][1] ), .Z(n1510) );
  ANDN U1837 ( .B(n1270), .A(\min_dist_reg[5][0] ), .Z(n1532) );
  IV U1838 ( .A(\min_dist_reg[5][2] ), .Z(n1503) );
  IV U1839 ( .A(\min_dist_reg[5][3] ), .Z(n1496) );
  IV U1840 ( .A(\min_dist_reg[5][4] ), .Z(n1517) );
  XOR U1841 ( .A(\min_dist_reg[5][0] ), .B(n1270), .Z(n1271) );
  XNOR U1842 ( .A(\min_dist_reg[6][0] ), .B(n1539), .Z(n1270) );
  NAND U1843 ( .A(n1246), .B(n974), .Z(n1539) );
  XOR U1844 ( .A(n1540), .B(n1541), .Z(n974) );
  AND U1845 ( .A(n1542), .B(n1543), .Z(n1540) );
  XNOR U1846 ( .A(n1541), .B(n1230), .Z(n1543) );
  XNOR U1847 ( .A(\min_dist_reg[7][4] ), .B(n1544), .Z(n1230) );
  NAND U1848 ( .A(n1545), .B(n977), .Z(n1544) );
  XOR U1849 ( .A(\min_dist_reg[7][4] ), .B(n1546), .Z(n1545) );
  XNOR U1850 ( .A(n1251), .B(n1541), .Z(n1542) );
  XOR U1851 ( .A(n1547), .B(n1253), .Z(n1541) );
  AND U1852 ( .A(n1254), .B(n1548), .Z(n1547) );
  XNOR U1853 ( .A(n1253), .B(n1233), .Z(n1548) );
  XNOR U1854 ( .A(\min_dist_reg[7][3] ), .B(n1549), .Z(n1233) );
  NAND U1855 ( .A(n1550), .B(n977), .Z(n1549) );
  XNOR U1856 ( .A(\min_dist_reg[7][3] ), .B(n1551), .Z(n1550) );
  XNOR U1857 ( .A(n1524), .B(n1253), .Z(n1254) );
  XOR U1858 ( .A(n1552), .B(n1553), .Z(n1253) );
  AND U1859 ( .A(n1554), .B(n1555), .Z(n1552) );
  XOR U1860 ( .A(n1239), .B(n1553), .Z(n1555) );
  IV U1861 ( .A(n1237), .Z(n1239) );
  XNOR U1862 ( .A(\min_dist_reg[7][2] ), .B(n1556), .Z(n1237) );
  NAND U1863 ( .A(n1557), .B(n977), .Z(n1556) );
  XNOR U1864 ( .A(\min_dist_reg[7][2] ), .B(n1558), .Z(n1557) );
  XNOR U1865 ( .A(n1531), .B(n1553), .Z(n1554) );
  XOR U1866 ( .A(n1559), .B(n1560), .Z(n1553) );
  NAND U1867 ( .A(n1561), .B(n1562), .Z(n1560) );
  XNOR U1868 ( .A(n1559), .B(n1243), .Z(n1562) );
  IV U1869 ( .A(n1241), .Z(n1243) );
  XNOR U1870 ( .A(\min_dist_reg[7][1] ), .B(n1563), .Z(n1241) );
  NAND U1871 ( .A(n1564), .B(n977), .Z(n1563) );
  XNOR U1872 ( .A(\min_dist_reg[7][1] ), .B(n1565), .Z(n1564) );
  XOR U1873 ( .A(n1538), .B(n1559), .Z(n1561) );
  IV U1874 ( .A(\min_dist_reg[6][1] ), .Z(n1538) );
  ANDN U1875 ( .B(n1245), .A(\min_dist_reg[6][0] ), .Z(n1559) );
  IV U1876 ( .A(\min_dist_reg[6][2] ), .Z(n1531) );
  IV U1877 ( .A(\min_dist_reg[6][3] ), .Z(n1524) );
  IV U1878 ( .A(\min_dist_reg[6][4] ), .Z(n1251) );
  XOR U1879 ( .A(\min_dist_reg[6][0] ), .B(n1245), .Z(n1246) );
  XOR U1880 ( .A(n1566), .B(n1567), .Z(n1245) );
  NAND U1881 ( .A(n1568), .B(n977), .Z(n1567) );
  XNOR U1882 ( .A(n1569), .B(n1570), .Z(n977) );
  AND U1883 ( .A(n1571), .B(n1572), .Z(n1569) );
  XNOR U1884 ( .A(n1573), .B(n1546), .Z(n1572) );
  XNOR U1885 ( .A(n1574), .B(n1575), .Z(n1546) );
  ANDN U1886 ( .B(n1576), .A(n1577), .Z(n1574) );
  XOR U1887 ( .A(n1575), .B(n1578), .Z(n1576) );
  XNOR U1888 ( .A(\min_dist_reg[7][4] ), .B(n1570), .Z(n1571) );
  IV U1889 ( .A(n1573), .Z(n1570) );
  XOR U1890 ( .A(n1579), .B(n1580), .Z(n1573) );
  AND U1891 ( .A(n1581), .B(n1582), .Z(n1579) );
  XOR U1892 ( .A(n1580), .B(n1551), .Z(n1582) );
  XOR U1893 ( .A(n1583), .B(n1578), .Z(n1551) );
  XNOR U1894 ( .A(n1584), .B(n1585), .Z(n1578) );
  ANDN U1895 ( .B(n1586), .A(n1587), .Z(n1584) );
  XOR U1896 ( .A(n1588), .B(n1589), .Z(n1586) );
  IV U1897 ( .A(n1577), .Z(n1583) );
  XOR U1898 ( .A(n1590), .B(n1591), .Z(n1577) );
  XNOR U1899 ( .A(n1592), .B(n1593), .Z(n1591) );
  ANDN U1900 ( .B(n1594), .A(n1595), .Z(n1592) );
  XNOR U1901 ( .A(n1596), .B(n1597), .Z(n1594) );
  IV U1902 ( .A(n1575), .Z(n1590) );
  XOR U1903 ( .A(n1598), .B(n1599), .Z(n1575) );
  ANDN U1904 ( .B(n1600), .A(n1601), .Z(n1598) );
  XOR U1905 ( .A(n1599), .B(n1602), .Z(n1600) );
  XNOR U1906 ( .A(\min_dist_reg[7][3] ), .B(n1603), .Z(n1581) );
  IV U1907 ( .A(n1580), .Z(n1603) );
  XOR U1908 ( .A(n1604), .B(n1605), .Z(n1580) );
  AND U1909 ( .A(n1606), .B(n1607), .Z(n1604) );
  XOR U1910 ( .A(n1605), .B(n1558), .Z(n1607) );
  XOR U1911 ( .A(n1608), .B(n1602), .Z(n1558) );
  XOR U1912 ( .A(n1609), .B(n1589), .Z(n1602) );
  XNOR U1913 ( .A(n1610), .B(n1611), .Z(n1589) );
  ANDN U1914 ( .B(n1612), .A(n1613), .Z(n1610) );
  XOR U1915 ( .A(n1614), .B(n1615), .Z(n1612) );
  IV U1916 ( .A(n1587), .Z(n1609) );
  XOR U1917 ( .A(n1585), .B(n1616), .Z(n1587) );
  XNOR U1918 ( .A(n1617), .B(n1618), .Z(n1616) );
  ANDN U1919 ( .B(n1619), .A(n1620), .Z(n1617) );
  XNOR U1920 ( .A(n1621), .B(n1622), .Z(n1619) );
  IV U1921 ( .A(n1588), .Z(n1585) );
  XOR U1922 ( .A(n1623), .B(n1624), .Z(n1588) );
  ANDN U1923 ( .B(n1625), .A(n1626), .Z(n1623) );
  XOR U1924 ( .A(n1624), .B(n1627), .Z(n1625) );
  IV U1925 ( .A(n1601), .Z(n1608) );
  XOR U1926 ( .A(n1628), .B(n1629), .Z(n1601) );
  XNOR U1927 ( .A(n1596), .B(n1630), .Z(n1629) );
  IV U1928 ( .A(n1599), .Z(n1630) );
  XOR U1929 ( .A(n1631), .B(n1632), .Z(n1599) );
  ANDN U1930 ( .B(n1633), .A(n1634), .Z(n1631) );
  XOR U1931 ( .A(n1632), .B(n1635), .Z(n1633) );
  XNOR U1932 ( .A(n1636), .B(n1637), .Z(n1596) );
  ANDN U1933 ( .B(n1638), .A(n1639), .Z(n1636) );
  XOR U1934 ( .A(n1637), .B(n1640), .Z(n1638) );
  IV U1935 ( .A(n1595), .Z(n1628) );
  XOR U1936 ( .A(n1593), .B(n1641), .Z(n1595) );
  XNOR U1937 ( .A(n1642), .B(n1643), .Z(n1641) );
  ANDN U1938 ( .B(n1644), .A(n1645), .Z(n1642) );
  XNOR U1939 ( .A(n1646), .B(n1647), .Z(n1644) );
  IV U1940 ( .A(n1597), .Z(n1593) );
  XOR U1941 ( .A(n1648), .B(n1649), .Z(n1597) );
  ANDN U1942 ( .B(n1650), .A(n1651), .Z(n1648) );
  XOR U1943 ( .A(n1652), .B(n1649), .Z(n1650) );
  XOR U1944 ( .A(\min_dist_reg[7][2] ), .B(n1605), .Z(n1606) );
  XOR U1945 ( .A(n1653), .B(n1654), .Z(n1605) );
  NAND U1946 ( .A(n1655), .B(n1656), .Z(n1654) );
  XNOR U1947 ( .A(n1653), .B(n1565), .Z(n1656) );
  XOR U1948 ( .A(n1657), .B(n1635), .Z(n1565) );
  XOR U1949 ( .A(n1658), .B(n1627), .Z(n1635) );
  XOR U1950 ( .A(n1659), .B(n1615), .Z(n1627) );
  XNOR U1951 ( .A(n1660), .B(n1661), .Z(n1615) );
  ANDN U1952 ( .B(n1662), .A(n1663), .Z(n1660) );
  XNOR U1953 ( .A(n1661), .B(n1664), .Z(n1662) );
  IV U1954 ( .A(n1613), .Z(n1659) );
  XOR U1955 ( .A(n1611), .B(n1665), .Z(n1613) );
  XNOR U1956 ( .A(n1666), .B(n1667), .Z(n1665) );
  ANDN U1957 ( .B(n1668), .A(n1669), .Z(n1666) );
  XNOR U1958 ( .A(n1670), .B(n1671), .Z(n1668) );
  IV U1959 ( .A(n1667), .Z(n1671) );
  IV U1960 ( .A(n1614), .Z(n1611) );
  XNOR U1961 ( .A(n1672), .B(n1673), .Z(n1614) );
  ANDN U1962 ( .B(n1674), .A(n1675), .Z(n1672) );
  XNOR U1963 ( .A(n1673), .B(n1676), .Z(n1674) );
  IV U1964 ( .A(n1626), .Z(n1658) );
  XOR U1965 ( .A(n1677), .B(n1678), .Z(n1626) );
  XNOR U1966 ( .A(n1621), .B(n1679), .Z(n1678) );
  IV U1967 ( .A(n1624), .Z(n1679) );
  XNOR U1968 ( .A(n1680), .B(n1681), .Z(n1624) );
  ANDN U1969 ( .B(n1682), .A(n1683), .Z(n1680) );
  XNOR U1970 ( .A(n1681), .B(n1684), .Z(n1682) );
  XOR U1971 ( .A(n1685), .B(n1686), .Z(n1621) );
  ANDN U1972 ( .B(n1687), .A(n1688), .Z(n1685) );
  XNOR U1973 ( .A(n1686), .B(n1689), .Z(n1687) );
  IV U1974 ( .A(n1620), .Z(n1677) );
  XOR U1975 ( .A(n1618), .B(n1690), .Z(n1620) );
  XNOR U1976 ( .A(n1691), .B(n1692), .Z(n1690) );
  ANDN U1977 ( .B(n1693), .A(n1694), .Z(n1691) );
  XNOR U1978 ( .A(n1695), .B(n1696), .Z(n1693) );
  IV U1979 ( .A(n1692), .Z(n1696) );
  IV U1980 ( .A(n1622), .Z(n1618) );
  XNOR U1981 ( .A(n1697), .B(n1698), .Z(n1622) );
  ANDN U1982 ( .B(n1699), .A(n1700), .Z(n1697) );
  XNOR U1983 ( .A(n1701), .B(n1698), .Z(n1699) );
  IV U1984 ( .A(n1634), .Z(n1657) );
  XOR U1985 ( .A(n1702), .B(n1703), .Z(n1634) );
  XOR U1986 ( .A(n1652), .B(n1704), .Z(n1703) );
  IV U1987 ( .A(n1632), .Z(n1704) );
  XNOR U1988 ( .A(n1705), .B(n1706), .Z(n1632) );
  ANDN U1989 ( .B(n1707), .A(n1708), .Z(n1705) );
  XNOR U1990 ( .A(n1706), .B(n1709), .Z(n1707) );
  XOR U1991 ( .A(n1710), .B(n1640), .Z(n1652) );
  XNOR U1992 ( .A(n1711), .B(n1712), .Z(n1640) );
  ANDN U1993 ( .B(n1713), .A(n1714), .Z(n1711) );
  XNOR U1994 ( .A(n1712), .B(n1715), .Z(n1713) );
  IV U1995 ( .A(n1639), .Z(n1710) );
  XOR U1996 ( .A(n1716), .B(n1717), .Z(n1639) );
  XNOR U1997 ( .A(n1718), .B(n1719), .Z(n1717) );
  ANDN U1998 ( .B(n1720), .A(n1721), .Z(n1718) );
  XNOR U1999 ( .A(n1722), .B(n1723), .Z(n1720) );
  IV U2000 ( .A(n1719), .Z(n1723) );
  IV U2001 ( .A(n1637), .Z(n1716) );
  XNOR U2002 ( .A(n1724), .B(n1725), .Z(n1637) );
  ANDN U2003 ( .B(n1726), .A(n1727), .Z(n1724) );
  XNOR U2004 ( .A(n1725), .B(n1728), .Z(n1726) );
  IV U2005 ( .A(n1651), .Z(n1702) );
  XOR U2006 ( .A(n1729), .B(n1730), .Z(n1651) );
  XNOR U2007 ( .A(n1646), .B(n1731), .Z(n1730) );
  IV U2008 ( .A(n1649), .Z(n1731) );
  XNOR U2009 ( .A(n1732), .B(n1733), .Z(n1649) );
  ANDN U2010 ( .B(n1734), .A(n1735), .Z(n1732) );
  XNOR U2011 ( .A(n1736), .B(n1733), .Z(n1734) );
  XOR U2012 ( .A(n1737), .B(n1738), .Z(n1646) );
  ANDN U2013 ( .B(n1739), .A(n1740), .Z(n1737) );
  XNOR U2014 ( .A(n1738), .B(n1741), .Z(n1739) );
  IV U2015 ( .A(n1645), .Z(n1729) );
  XOR U2016 ( .A(n1643), .B(n1742), .Z(n1645) );
  XNOR U2017 ( .A(n1743), .B(n1744), .Z(n1742) );
  ANDN U2018 ( .B(n1745), .A(n1746), .Z(n1743) );
  XNOR U2019 ( .A(n1747), .B(n1748), .Z(n1745) );
  IV U2020 ( .A(n1744), .Z(n1748) );
  IV U2021 ( .A(n1647), .Z(n1643) );
  XNOR U2022 ( .A(n1749), .B(n1750), .Z(n1647) );
  ANDN U2023 ( .B(n1751), .A(n1752), .Z(n1749) );
  XNOR U2024 ( .A(n1753), .B(n1750), .Z(n1751) );
  XNOR U2025 ( .A(\min_dist_reg[7][1] ), .B(n1653), .Z(n1655) );
  NOR U2026 ( .A(\min_dist_reg[7][0] ), .B(n1754), .Z(n1653) );
  XOR U2027 ( .A(n1566), .B(n1754), .Z(n1568) );
  XOR U2028 ( .A(n1755), .B(n1709), .Z(n1754) );
  XOR U2029 ( .A(n1756), .B(n1684), .Z(n1709) );
  XOR U2030 ( .A(n1757), .B(n1676), .Z(n1684) );
  XOR U2031 ( .A(n1758), .B(n1664), .Z(n1676) );
  XNOR U2032 ( .A(q[30]), .B(DB[30]), .Z(n1664) );
  IV U2033 ( .A(n1663), .Z(n1758) );
  XOR U2034 ( .A(n1661), .B(n1759), .Z(n1663) );
  XNOR U2035 ( .A(q[29]), .B(DB[29]), .Z(n1759) );
  XOR U2036 ( .A(q[28]), .B(DB[28]), .Z(n1661) );
  IV U2037 ( .A(n1675), .Z(n1757) );
  XOR U2038 ( .A(n1760), .B(n1761), .Z(n1675) );
  XNOR U2039 ( .A(n1670), .B(n1673), .Z(n1761) );
  XOR U2040 ( .A(q[24]), .B(DB[24]), .Z(n1673) );
  XOR U2041 ( .A(q[27]), .B(DB[27]), .Z(n1670) );
  IV U2042 ( .A(n1669), .Z(n1760) );
  XOR U2043 ( .A(n1667), .B(n1762), .Z(n1669) );
  XNOR U2044 ( .A(q[26]), .B(DB[26]), .Z(n1762) );
  XOR U2045 ( .A(q[25]), .B(DB[25]), .Z(n1667) );
  IV U2046 ( .A(n1683), .Z(n1756) );
  XOR U2047 ( .A(n1763), .B(n1764), .Z(n1683) );
  XOR U2048 ( .A(n1701), .B(n1681), .Z(n1764) );
  XOR U2049 ( .A(q[16]), .B(DB[16]), .Z(n1681) );
  XOR U2050 ( .A(n1765), .B(n1689), .Z(n1701) );
  XNOR U2051 ( .A(q[23]), .B(DB[23]), .Z(n1689) );
  IV U2052 ( .A(n1688), .Z(n1765) );
  XOR U2053 ( .A(n1686), .B(n1766), .Z(n1688) );
  XNOR U2054 ( .A(q[22]), .B(DB[22]), .Z(n1766) );
  XOR U2055 ( .A(q[21]), .B(DB[21]), .Z(n1686) );
  IV U2056 ( .A(n1700), .Z(n1763) );
  XOR U2057 ( .A(n1767), .B(n1768), .Z(n1700) );
  XNOR U2058 ( .A(n1695), .B(n1698), .Z(n1768) );
  XOR U2059 ( .A(q[17]), .B(DB[17]), .Z(n1698) );
  XOR U2060 ( .A(q[20]), .B(DB[20]), .Z(n1695) );
  IV U2061 ( .A(n1694), .Z(n1767) );
  XOR U2062 ( .A(n1692), .B(n1769), .Z(n1694) );
  XNOR U2063 ( .A(q[19]), .B(DB[19]), .Z(n1769) );
  XOR U2064 ( .A(q[18]), .B(DB[18]), .Z(n1692) );
  IV U2065 ( .A(n1708), .Z(n1755) );
  XOR U2066 ( .A(n1770), .B(n1771), .Z(n1708) );
  XOR U2067 ( .A(n1736), .B(n1706), .Z(n1771) );
  XOR U2068 ( .A(q[0]), .B(DB[0]), .Z(n1706) );
  XOR U2069 ( .A(n1772), .B(n1728), .Z(n1736) );
  XOR U2070 ( .A(n1773), .B(n1715), .Z(n1728) );
  XNOR U2071 ( .A(q[15]), .B(DB[15]), .Z(n1715) );
  IV U2072 ( .A(n1714), .Z(n1773) );
  XOR U2073 ( .A(n1712), .B(n1774), .Z(n1714) );
  XNOR U2074 ( .A(q[14]), .B(DB[14]), .Z(n1774) );
  XOR U2075 ( .A(q[13]), .B(DB[13]), .Z(n1712) );
  IV U2076 ( .A(n1727), .Z(n1772) );
  XOR U2077 ( .A(n1775), .B(n1776), .Z(n1727) );
  XNOR U2078 ( .A(n1722), .B(n1725), .Z(n1776) );
  XOR U2079 ( .A(q[9]), .B(DB[9]), .Z(n1725) );
  XOR U2080 ( .A(q[12]), .B(DB[12]), .Z(n1722) );
  IV U2081 ( .A(n1721), .Z(n1775) );
  XOR U2082 ( .A(n1719), .B(n1777), .Z(n1721) );
  XNOR U2083 ( .A(q[11]), .B(DB[11]), .Z(n1777) );
  XOR U2084 ( .A(q[10]), .B(DB[10]), .Z(n1719) );
  IV U2085 ( .A(n1735), .Z(n1770) );
  XOR U2086 ( .A(n1778), .B(n1779), .Z(n1735) );
  XOR U2087 ( .A(n1753), .B(n1733), .Z(n1779) );
  XOR U2088 ( .A(q[1]), .B(DB[1]), .Z(n1733) );
  XOR U2089 ( .A(n1780), .B(n1741), .Z(n1753) );
  XNOR U2090 ( .A(q[8]), .B(DB[8]), .Z(n1741) );
  IV U2091 ( .A(n1740), .Z(n1780) );
  XOR U2092 ( .A(n1738), .B(n1781), .Z(n1740) );
  XNOR U2093 ( .A(q[7]), .B(DB[7]), .Z(n1781) );
  XOR U2094 ( .A(q[6]), .B(DB[6]), .Z(n1738) );
  IV U2095 ( .A(n1752), .Z(n1778) );
  XOR U2096 ( .A(n1782), .B(n1783), .Z(n1752) );
  XNOR U2097 ( .A(n1747), .B(n1750), .Z(n1783) );
  XOR U2098 ( .A(q[2]), .B(DB[2]), .Z(n1750) );
  XOR U2099 ( .A(q[5]), .B(DB[5]), .Z(n1747) );
  IV U2100 ( .A(n1746), .Z(n1782) );
  XOR U2101 ( .A(n1744), .B(n1784), .Z(n1746) );
  XNOR U2102 ( .A(q[4]), .B(DB[4]), .Z(n1784) );
  XOR U2103 ( .A(q[3]), .B(DB[3]), .Z(n1744) );
  IV U2104 ( .A(\min_dist_reg[7][0] ), .Z(n1566) );
  IV U2105 ( .A(\min_dist_reg[1][0] ), .Z(n1426) );
endmodule

