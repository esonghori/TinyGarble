
module sum_N256_CC1 ( clk, rst, a, b, c );
  input [255:0] a;
  input [255:0] b;
  output [255:0] c;
  input clk, rst;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020;

  NANDN U2 ( .A(n854), .B(b[254]), .Z(n2) );
  XNOR U3 ( .A(n854), .B(b[254]), .Z(n3) );
  NAND U4 ( .A(n3), .B(a[254]), .Z(n4) );
  NAND U5 ( .A(n2), .B(n4), .Z(n5) );
  XNOR U6 ( .A(a[255]), .B(n5), .Z(n6) );
  XNOR U7 ( .A(b[255]), .B(n6), .Z(c[255]) );
  XOR U8 ( .A(a[0]), .B(b[0]), .Z(c[0]) );
  XOR U9 ( .A(a[100]), .B(b[100]), .Z(n205) );
  NAND U10 ( .A(b[99]), .B(a[99]), .Z(n204) );
  XNOR U11 ( .A(b[99]), .B(a[99]), .Z(n1018) );
  NAND U12 ( .A(b[98]), .B(a[98]), .Z(n202) );
  NAND U13 ( .A(b[97]), .B(a[97]), .Z(n200) );
  NAND U14 ( .A(b[96]), .B(a[96]), .Z(n198) );
  NAND U15 ( .A(b[95]), .B(a[95]), .Z(n196) );
  NAND U16 ( .A(b[94]), .B(a[94]), .Z(n194) );
  NAND U17 ( .A(b[93]), .B(a[93]), .Z(n192) );
  NAND U18 ( .A(b[92]), .B(a[92]), .Z(n190) );
  NAND U19 ( .A(b[91]), .B(a[91]), .Z(n188) );
  NAND U20 ( .A(b[90]), .B(a[90]), .Z(n186) );
  NAND U21 ( .A(b[89]), .B(a[89]), .Z(n184) );
  NAND U22 ( .A(b[88]), .B(a[88]), .Z(n182) );
  NAND U23 ( .A(b[87]), .B(a[87]), .Z(n180) );
  NAND U24 ( .A(b[86]), .B(a[86]), .Z(n178) );
  NAND U25 ( .A(b[85]), .B(a[85]), .Z(n176) );
  NAND U26 ( .A(b[84]), .B(a[84]), .Z(n174) );
  NAND U27 ( .A(b[83]), .B(a[83]), .Z(n172) );
  NAND U28 ( .A(b[82]), .B(a[82]), .Z(n170) );
  NAND U29 ( .A(b[81]), .B(a[81]), .Z(n168) );
  NAND U30 ( .A(b[80]), .B(a[80]), .Z(n166) );
  NAND U31 ( .A(b[79]), .B(a[79]), .Z(n164) );
  NAND U32 ( .A(b[78]), .B(a[78]), .Z(n162) );
  NAND U33 ( .A(b[77]), .B(a[77]), .Z(n160) );
  NAND U34 ( .A(b[76]), .B(a[76]), .Z(n158) );
  NAND U35 ( .A(b[75]), .B(a[75]), .Z(n156) );
  NAND U36 ( .A(b[74]), .B(a[74]), .Z(n154) );
  NAND U37 ( .A(b[73]), .B(a[73]), .Z(n152) );
  NAND U38 ( .A(b[72]), .B(a[72]), .Z(n150) );
  NAND U39 ( .A(b[71]), .B(a[71]), .Z(n148) );
  NAND U40 ( .A(b[70]), .B(a[70]), .Z(n146) );
  NAND U41 ( .A(b[69]), .B(a[69]), .Z(n144) );
  NAND U42 ( .A(b[68]), .B(a[68]), .Z(n142) );
  NAND U43 ( .A(b[67]), .B(a[67]), .Z(n140) );
  NAND U44 ( .A(b[66]), .B(a[66]), .Z(n138) );
  NAND U45 ( .A(b[65]), .B(a[65]), .Z(n136) );
  NAND U46 ( .A(b[64]), .B(a[64]), .Z(n134) );
  NAND U47 ( .A(b[63]), .B(a[63]), .Z(n132) );
  NAND U48 ( .A(b[62]), .B(a[62]), .Z(n130) );
  NAND U49 ( .A(b[61]), .B(a[61]), .Z(n128) );
  NAND U50 ( .A(b[60]), .B(a[60]), .Z(n126) );
  NAND U51 ( .A(b[59]), .B(a[59]), .Z(n124) );
  NAND U52 ( .A(b[58]), .B(a[58]), .Z(n122) );
  NAND U53 ( .A(b[57]), .B(a[57]), .Z(n120) );
  NAND U54 ( .A(b[56]), .B(a[56]), .Z(n118) );
  NAND U55 ( .A(b[55]), .B(a[55]), .Z(n116) );
  NAND U56 ( .A(b[54]), .B(a[54]), .Z(n114) );
  NAND U57 ( .A(b[53]), .B(a[53]), .Z(n112) );
  NAND U58 ( .A(b[52]), .B(a[52]), .Z(n110) );
  NAND U59 ( .A(b[51]), .B(a[51]), .Z(n108) );
  NAND U60 ( .A(b[50]), .B(a[50]), .Z(n106) );
  NAND U61 ( .A(b[49]), .B(a[49]), .Z(n104) );
  NAND U62 ( .A(b[48]), .B(a[48]), .Z(n102) );
  NAND U63 ( .A(b[47]), .B(a[47]), .Z(n100) );
  NAND U64 ( .A(b[46]), .B(a[46]), .Z(n98) );
  NAND U65 ( .A(b[45]), .B(a[45]), .Z(n96) );
  NAND U66 ( .A(b[44]), .B(a[44]), .Z(n94) );
  NAND U67 ( .A(b[43]), .B(a[43]), .Z(n92) );
  NAND U68 ( .A(b[42]), .B(a[42]), .Z(n90) );
  NAND U69 ( .A(b[41]), .B(a[41]), .Z(n88) );
  NAND U70 ( .A(b[40]), .B(a[40]), .Z(n86) );
  NAND U71 ( .A(b[39]), .B(a[39]), .Z(n84) );
  NAND U72 ( .A(b[38]), .B(a[38]), .Z(n82) );
  NAND U73 ( .A(b[37]), .B(a[37]), .Z(n80) );
  NAND U74 ( .A(b[36]), .B(a[36]), .Z(n78) );
  NAND U75 ( .A(b[35]), .B(a[35]), .Z(n76) );
  NAND U76 ( .A(b[34]), .B(a[34]), .Z(n74) );
  NAND U77 ( .A(b[33]), .B(a[33]), .Z(n72) );
  NAND U78 ( .A(b[32]), .B(a[32]), .Z(n70) );
  NAND U79 ( .A(b[31]), .B(a[31]), .Z(n68) );
  NAND U80 ( .A(b[30]), .B(a[30]), .Z(n66) );
  NAND U81 ( .A(b[29]), .B(a[29]), .Z(n64) );
  NAND U82 ( .A(b[28]), .B(a[28]), .Z(n62) );
  NAND U83 ( .A(b[27]), .B(a[27]), .Z(n60) );
  NAND U84 ( .A(b[26]), .B(a[26]), .Z(n58) );
  NAND U85 ( .A(b[25]), .B(a[25]), .Z(n56) );
  NAND U86 ( .A(b[24]), .B(a[24]), .Z(n54) );
  NAND U87 ( .A(b[23]), .B(a[23]), .Z(n52) );
  NAND U88 ( .A(b[22]), .B(a[22]), .Z(n50) );
  NAND U89 ( .A(b[21]), .B(a[21]), .Z(n48) );
  NAND U90 ( .A(b[20]), .B(a[20]), .Z(n46) );
  NAND U91 ( .A(b[19]), .B(a[19]), .Z(n44) );
  NAND U92 ( .A(b[18]), .B(a[18]), .Z(n42) );
  NAND U93 ( .A(b[17]), .B(a[17]), .Z(n40) );
  NAND U94 ( .A(b[16]), .B(a[16]), .Z(n38) );
  NAND U95 ( .A(b[15]), .B(a[15]), .Z(n36) );
  NAND U96 ( .A(b[14]), .B(a[14]), .Z(n34) );
  NAND U97 ( .A(b[13]), .B(a[13]), .Z(n32) );
  NAND U98 ( .A(b[12]), .B(a[12]), .Z(n30) );
  NAND U99 ( .A(b[11]), .B(a[11]), .Z(n28) );
  NAND U100 ( .A(b[10]), .B(a[10]), .Z(n26) );
  NAND U101 ( .A(b[9]), .B(a[9]), .Z(n24) );
  XNOR U102 ( .A(b[9]), .B(a[9]), .Z(n1020) );
  NAND U103 ( .A(b[8]), .B(a[8]), .Z(n22) );
  NAND U104 ( .A(b[7]), .B(a[7]), .Z(n20) );
  NAND U105 ( .A(b[6]), .B(a[6]), .Z(n18) );
  NAND U106 ( .A(b[5]), .B(a[5]), .Z(n16) );
  NAND U107 ( .A(b[4]), .B(a[4]), .Z(n14) );
  NAND U108 ( .A(b[3]), .B(a[3]), .Z(n12) );
  NAND U109 ( .A(b[2]), .B(a[2]), .Z(n10) );
  NAND U110 ( .A(b[1]), .B(a[1]), .Z(n8) );
  NAND U111 ( .A(a[0]), .B(b[0]), .Z(n621) );
  XOR U112 ( .A(a[1]), .B(b[1]), .Z(n622) );
  NANDN U113 ( .A(n621), .B(n622), .Z(n7) );
  AND U114 ( .A(n8), .B(n7), .Z(n865) );
  XOR U115 ( .A(a[2]), .B(b[2]), .Z(n866) );
  NANDN U116 ( .A(n865), .B(n866), .Z(n9) );
  AND U117 ( .A(n10), .B(n9), .Z(n887) );
  XOR U118 ( .A(a[3]), .B(b[3]), .Z(n888) );
  NANDN U119 ( .A(n887), .B(n888), .Z(n11) );
  AND U120 ( .A(n12), .B(n11), .Z(n909) );
  XOR U121 ( .A(a[4]), .B(b[4]), .Z(n910) );
  NANDN U122 ( .A(n909), .B(n910), .Z(n13) );
  AND U123 ( .A(n14), .B(n13), .Z(n931) );
  XOR U124 ( .A(a[5]), .B(b[5]), .Z(n932) );
  NANDN U125 ( .A(n931), .B(n932), .Z(n15) );
  AND U126 ( .A(n16), .B(n15), .Z(n953) );
  XOR U127 ( .A(a[6]), .B(b[6]), .Z(n954) );
  NANDN U128 ( .A(n953), .B(n954), .Z(n17) );
  AND U129 ( .A(n18), .B(n17), .Z(n975) );
  XOR U130 ( .A(a[7]), .B(b[7]), .Z(n976) );
  NANDN U131 ( .A(n975), .B(n976), .Z(n19) );
  AND U132 ( .A(n20), .B(n19), .Z(n997) );
  XOR U133 ( .A(a[8]), .B(b[8]), .Z(n998) );
  NANDN U134 ( .A(n997), .B(n998), .Z(n21) );
  AND U135 ( .A(n22), .B(n21), .Z(n1019) );
  OR U136 ( .A(n1020), .B(n1019), .Z(n23) );
  AND U137 ( .A(n24), .B(n23), .Z(n241) );
  XOR U138 ( .A(a[10]), .B(b[10]), .Z(n242) );
  NANDN U139 ( .A(n241), .B(n242), .Z(n25) );
  AND U140 ( .A(n26), .B(n25), .Z(n283) );
  XOR U141 ( .A(a[11]), .B(b[11]), .Z(n284) );
  NANDN U142 ( .A(n283), .B(n284), .Z(n27) );
  AND U143 ( .A(n28), .B(n27), .Z(n325) );
  XOR U144 ( .A(a[12]), .B(b[12]), .Z(n326) );
  NANDN U145 ( .A(n325), .B(n326), .Z(n29) );
  AND U146 ( .A(n30), .B(n29), .Z(n367) );
  XOR U147 ( .A(a[13]), .B(b[13]), .Z(n368) );
  NANDN U148 ( .A(n367), .B(n368), .Z(n31) );
  AND U149 ( .A(n32), .B(n31), .Z(n409) );
  XOR U150 ( .A(a[14]), .B(b[14]), .Z(n410) );
  NANDN U151 ( .A(n409), .B(n410), .Z(n33) );
  AND U152 ( .A(n34), .B(n33), .Z(n451) );
  XOR U153 ( .A(a[15]), .B(b[15]), .Z(n452) );
  NANDN U154 ( .A(n451), .B(n452), .Z(n35) );
  AND U155 ( .A(n36), .B(n35), .Z(n493) );
  XOR U156 ( .A(a[16]), .B(b[16]), .Z(n494) );
  NANDN U157 ( .A(n493), .B(n494), .Z(n37) );
  AND U158 ( .A(n38), .B(n37), .Z(n535) );
  XOR U159 ( .A(a[17]), .B(b[17]), .Z(n536) );
  NANDN U160 ( .A(n535), .B(n536), .Z(n39) );
  AND U161 ( .A(n40), .B(n39), .Z(n577) );
  XOR U162 ( .A(a[18]), .B(b[18]), .Z(n578) );
  NANDN U163 ( .A(n577), .B(n578), .Z(n41) );
  AND U164 ( .A(n42), .B(n41), .Z(n619) );
  XOR U165 ( .A(a[19]), .B(b[19]), .Z(n620) );
  NANDN U166 ( .A(n619), .B(n620), .Z(n43) );
  AND U167 ( .A(n44), .B(n43), .Z(n663) );
  XOR U168 ( .A(a[20]), .B(b[20]), .Z(n664) );
  NANDN U169 ( .A(n663), .B(n664), .Z(n45) );
  AND U170 ( .A(n46), .B(n45), .Z(n705) );
  XOR U171 ( .A(a[21]), .B(b[21]), .Z(n706) );
  NANDN U172 ( .A(n705), .B(n706), .Z(n47) );
  AND U173 ( .A(n48), .B(n47), .Z(n747) );
  XOR U174 ( .A(a[22]), .B(b[22]), .Z(n748) );
  NANDN U175 ( .A(n747), .B(n748), .Z(n49) );
  AND U176 ( .A(n50), .B(n49), .Z(n789) );
  XOR U177 ( .A(a[23]), .B(b[23]), .Z(n790) );
  NANDN U178 ( .A(n789), .B(n790), .Z(n51) );
  AND U179 ( .A(n52), .B(n51), .Z(n831) );
  XOR U180 ( .A(a[24]), .B(b[24]), .Z(n832) );
  NANDN U181 ( .A(n831), .B(n832), .Z(n53) );
  AND U182 ( .A(n54), .B(n53), .Z(n855) );
  XOR U183 ( .A(a[25]), .B(b[25]), .Z(n856) );
  NANDN U184 ( .A(n855), .B(n856), .Z(n55) );
  AND U185 ( .A(n56), .B(n55), .Z(n857) );
  XOR U186 ( .A(a[26]), .B(b[26]), .Z(n858) );
  NANDN U187 ( .A(n857), .B(n858), .Z(n57) );
  AND U188 ( .A(n58), .B(n57), .Z(n859) );
  XOR U189 ( .A(a[27]), .B(b[27]), .Z(n860) );
  NANDN U190 ( .A(n859), .B(n860), .Z(n59) );
  AND U191 ( .A(n60), .B(n59), .Z(n861) );
  XOR U192 ( .A(a[28]), .B(b[28]), .Z(n862) );
  NANDN U193 ( .A(n861), .B(n862), .Z(n61) );
  AND U194 ( .A(n62), .B(n61), .Z(n863) );
  XOR U195 ( .A(a[29]), .B(b[29]), .Z(n864) );
  NANDN U196 ( .A(n863), .B(n864), .Z(n63) );
  AND U197 ( .A(n64), .B(n63), .Z(n867) );
  XOR U198 ( .A(a[30]), .B(b[30]), .Z(n868) );
  NANDN U199 ( .A(n867), .B(n868), .Z(n65) );
  AND U200 ( .A(n66), .B(n65), .Z(n869) );
  XOR U201 ( .A(a[31]), .B(b[31]), .Z(n870) );
  NANDN U202 ( .A(n869), .B(n870), .Z(n67) );
  AND U203 ( .A(n68), .B(n67), .Z(n871) );
  XOR U204 ( .A(a[32]), .B(b[32]), .Z(n872) );
  NANDN U205 ( .A(n871), .B(n872), .Z(n69) );
  AND U206 ( .A(n70), .B(n69), .Z(n873) );
  XOR U207 ( .A(a[33]), .B(b[33]), .Z(n874) );
  NANDN U208 ( .A(n873), .B(n874), .Z(n71) );
  AND U209 ( .A(n72), .B(n71), .Z(n875) );
  XOR U210 ( .A(a[34]), .B(b[34]), .Z(n876) );
  NANDN U211 ( .A(n875), .B(n876), .Z(n73) );
  AND U212 ( .A(n74), .B(n73), .Z(n877) );
  XOR U213 ( .A(a[35]), .B(b[35]), .Z(n878) );
  NANDN U214 ( .A(n877), .B(n878), .Z(n75) );
  AND U215 ( .A(n76), .B(n75), .Z(n879) );
  XOR U216 ( .A(a[36]), .B(b[36]), .Z(n880) );
  NANDN U217 ( .A(n879), .B(n880), .Z(n77) );
  AND U218 ( .A(n78), .B(n77), .Z(n881) );
  XOR U219 ( .A(a[37]), .B(b[37]), .Z(n882) );
  NANDN U220 ( .A(n881), .B(n882), .Z(n79) );
  AND U221 ( .A(n80), .B(n79), .Z(n883) );
  XOR U222 ( .A(a[38]), .B(b[38]), .Z(n884) );
  NANDN U223 ( .A(n883), .B(n884), .Z(n81) );
  AND U224 ( .A(n82), .B(n81), .Z(n885) );
  XOR U225 ( .A(a[39]), .B(b[39]), .Z(n886) );
  NANDN U226 ( .A(n885), .B(n886), .Z(n83) );
  AND U227 ( .A(n84), .B(n83), .Z(n889) );
  XOR U228 ( .A(a[40]), .B(b[40]), .Z(n890) );
  NANDN U229 ( .A(n889), .B(n890), .Z(n85) );
  AND U230 ( .A(n86), .B(n85), .Z(n891) );
  XOR U231 ( .A(a[41]), .B(b[41]), .Z(n892) );
  NANDN U232 ( .A(n891), .B(n892), .Z(n87) );
  AND U233 ( .A(n88), .B(n87), .Z(n893) );
  XOR U234 ( .A(a[42]), .B(b[42]), .Z(n894) );
  NANDN U235 ( .A(n893), .B(n894), .Z(n89) );
  AND U236 ( .A(n90), .B(n89), .Z(n895) );
  XOR U237 ( .A(a[43]), .B(b[43]), .Z(n896) );
  NANDN U238 ( .A(n895), .B(n896), .Z(n91) );
  AND U239 ( .A(n92), .B(n91), .Z(n897) );
  XOR U240 ( .A(a[44]), .B(b[44]), .Z(n898) );
  NANDN U241 ( .A(n897), .B(n898), .Z(n93) );
  AND U242 ( .A(n94), .B(n93), .Z(n899) );
  XOR U243 ( .A(a[45]), .B(b[45]), .Z(n900) );
  NANDN U244 ( .A(n899), .B(n900), .Z(n95) );
  AND U245 ( .A(n96), .B(n95), .Z(n901) );
  XOR U246 ( .A(a[46]), .B(b[46]), .Z(n902) );
  NANDN U247 ( .A(n901), .B(n902), .Z(n97) );
  AND U248 ( .A(n98), .B(n97), .Z(n903) );
  XOR U249 ( .A(a[47]), .B(b[47]), .Z(n904) );
  NANDN U250 ( .A(n903), .B(n904), .Z(n99) );
  AND U251 ( .A(n100), .B(n99), .Z(n905) );
  XOR U252 ( .A(a[48]), .B(b[48]), .Z(n906) );
  NANDN U253 ( .A(n905), .B(n906), .Z(n101) );
  AND U254 ( .A(n102), .B(n101), .Z(n907) );
  XOR U255 ( .A(a[49]), .B(b[49]), .Z(n908) );
  NANDN U256 ( .A(n907), .B(n908), .Z(n103) );
  AND U257 ( .A(n104), .B(n103), .Z(n911) );
  XOR U258 ( .A(a[50]), .B(b[50]), .Z(n912) );
  NANDN U259 ( .A(n911), .B(n912), .Z(n105) );
  AND U260 ( .A(n106), .B(n105), .Z(n913) );
  XOR U261 ( .A(a[51]), .B(b[51]), .Z(n914) );
  NANDN U262 ( .A(n913), .B(n914), .Z(n107) );
  AND U263 ( .A(n108), .B(n107), .Z(n915) );
  XOR U264 ( .A(a[52]), .B(b[52]), .Z(n916) );
  NANDN U265 ( .A(n915), .B(n916), .Z(n109) );
  AND U266 ( .A(n110), .B(n109), .Z(n917) );
  XOR U267 ( .A(a[53]), .B(b[53]), .Z(n918) );
  NANDN U268 ( .A(n917), .B(n918), .Z(n111) );
  AND U269 ( .A(n112), .B(n111), .Z(n919) );
  XOR U270 ( .A(a[54]), .B(b[54]), .Z(n920) );
  NANDN U271 ( .A(n919), .B(n920), .Z(n113) );
  AND U272 ( .A(n114), .B(n113), .Z(n921) );
  XOR U273 ( .A(a[55]), .B(b[55]), .Z(n922) );
  NANDN U274 ( .A(n921), .B(n922), .Z(n115) );
  AND U275 ( .A(n116), .B(n115), .Z(n923) );
  XOR U276 ( .A(a[56]), .B(b[56]), .Z(n924) );
  NANDN U277 ( .A(n923), .B(n924), .Z(n117) );
  AND U278 ( .A(n118), .B(n117), .Z(n925) );
  XOR U279 ( .A(a[57]), .B(b[57]), .Z(n926) );
  NANDN U280 ( .A(n925), .B(n926), .Z(n119) );
  AND U281 ( .A(n120), .B(n119), .Z(n927) );
  XOR U282 ( .A(a[58]), .B(b[58]), .Z(n928) );
  NANDN U283 ( .A(n927), .B(n928), .Z(n121) );
  AND U284 ( .A(n122), .B(n121), .Z(n929) );
  XOR U285 ( .A(a[59]), .B(b[59]), .Z(n930) );
  NANDN U286 ( .A(n929), .B(n930), .Z(n123) );
  AND U287 ( .A(n124), .B(n123), .Z(n933) );
  XOR U288 ( .A(a[60]), .B(b[60]), .Z(n934) );
  NANDN U289 ( .A(n933), .B(n934), .Z(n125) );
  AND U290 ( .A(n126), .B(n125), .Z(n935) );
  XOR U291 ( .A(a[61]), .B(b[61]), .Z(n936) );
  NANDN U292 ( .A(n935), .B(n936), .Z(n127) );
  AND U293 ( .A(n128), .B(n127), .Z(n937) );
  XOR U294 ( .A(a[62]), .B(b[62]), .Z(n938) );
  NANDN U295 ( .A(n937), .B(n938), .Z(n129) );
  AND U296 ( .A(n130), .B(n129), .Z(n939) );
  XOR U297 ( .A(a[63]), .B(b[63]), .Z(n940) );
  NANDN U298 ( .A(n939), .B(n940), .Z(n131) );
  AND U299 ( .A(n132), .B(n131), .Z(n941) );
  XOR U300 ( .A(a[64]), .B(b[64]), .Z(n942) );
  NANDN U301 ( .A(n941), .B(n942), .Z(n133) );
  AND U302 ( .A(n134), .B(n133), .Z(n943) );
  XOR U303 ( .A(a[65]), .B(b[65]), .Z(n944) );
  NANDN U304 ( .A(n943), .B(n944), .Z(n135) );
  AND U305 ( .A(n136), .B(n135), .Z(n945) );
  XOR U306 ( .A(a[66]), .B(b[66]), .Z(n946) );
  NANDN U307 ( .A(n945), .B(n946), .Z(n137) );
  AND U308 ( .A(n138), .B(n137), .Z(n947) );
  XOR U309 ( .A(a[67]), .B(b[67]), .Z(n948) );
  NANDN U310 ( .A(n947), .B(n948), .Z(n139) );
  AND U311 ( .A(n140), .B(n139), .Z(n949) );
  XOR U312 ( .A(a[68]), .B(b[68]), .Z(n950) );
  NANDN U313 ( .A(n949), .B(n950), .Z(n141) );
  AND U314 ( .A(n142), .B(n141), .Z(n951) );
  XOR U315 ( .A(a[69]), .B(b[69]), .Z(n952) );
  NANDN U316 ( .A(n951), .B(n952), .Z(n143) );
  AND U317 ( .A(n144), .B(n143), .Z(n955) );
  XOR U318 ( .A(a[70]), .B(b[70]), .Z(n956) );
  NANDN U319 ( .A(n955), .B(n956), .Z(n145) );
  AND U320 ( .A(n146), .B(n145), .Z(n957) );
  XOR U321 ( .A(a[71]), .B(b[71]), .Z(n958) );
  NANDN U322 ( .A(n957), .B(n958), .Z(n147) );
  AND U323 ( .A(n148), .B(n147), .Z(n959) );
  XOR U324 ( .A(a[72]), .B(b[72]), .Z(n960) );
  NANDN U325 ( .A(n959), .B(n960), .Z(n149) );
  AND U326 ( .A(n150), .B(n149), .Z(n961) );
  XOR U327 ( .A(a[73]), .B(b[73]), .Z(n962) );
  NANDN U328 ( .A(n961), .B(n962), .Z(n151) );
  AND U329 ( .A(n152), .B(n151), .Z(n963) );
  XOR U330 ( .A(a[74]), .B(b[74]), .Z(n964) );
  NANDN U331 ( .A(n963), .B(n964), .Z(n153) );
  AND U332 ( .A(n154), .B(n153), .Z(n965) );
  XOR U333 ( .A(a[75]), .B(b[75]), .Z(n966) );
  NANDN U334 ( .A(n965), .B(n966), .Z(n155) );
  AND U335 ( .A(n156), .B(n155), .Z(n967) );
  XOR U336 ( .A(a[76]), .B(b[76]), .Z(n968) );
  NANDN U337 ( .A(n967), .B(n968), .Z(n157) );
  AND U338 ( .A(n158), .B(n157), .Z(n969) );
  XOR U339 ( .A(a[77]), .B(b[77]), .Z(n970) );
  NANDN U340 ( .A(n969), .B(n970), .Z(n159) );
  AND U341 ( .A(n160), .B(n159), .Z(n971) );
  XOR U342 ( .A(a[78]), .B(b[78]), .Z(n972) );
  NANDN U343 ( .A(n971), .B(n972), .Z(n161) );
  AND U344 ( .A(n162), .B(n161), .Z(n973) );
  XOR U345 ( .A(a[79]), .B(b[79]), .Z(n974) );
  NANDN U346 ( .A(n973), .B(n974), .Z(n163) );
  AND U347 ( .A(n164), .B(n163), .Z(n977) );
  XOR U348 ( .A(a[80]), .B(b[80]), .Z(n978) );
  NANDN U349 ( .A(n977), .B(n978), .Z(n165) );
  AND U350 ( .A(n166), .B(n165), .Z(n979) );
  XOR U351 ( .A(a[81]), .B(b[81]), .Z(n980) );
  NANDN U352 ( .A(n979), .B(n980), .Z(n167) );
  AND U353 ( .A(n168), .B(n167), .Z(n981) );
  XOR U354 ( .A(a[82]), .B(b[82]), .Z(n982) );
  NANDN U355 ( .A(n981), .B(n982), .Z(n169) );
  AND U356 ( .A(n170), .B(n169), .Z(n983) );
  XOR U357 ( .A(a[83]), .B(b[83]), .Z(n984) );
  NANDN U358 ( .A(n983), .B(n984), .Z(n171) );
  AND U359 ( .A(n172), .B(n171), .Z(n985) );
  XOR U360 ( .A(a[84]), .B(b[84]), .Z(n986) );
  NANDN U361 ( .A(n985), .B(n986), .Z(n173) );
  AND U362 ( .A(n174), .B(n173), .Z(n987) );
  XOR U363 ( .A(a[85]), .B(b[85]), .Z(n988) );
  NANDN U364 ( .A(n987), .B(n988), .Z(n175) );
  AND U365 ( .A(n176), .B(n175), .Z(n989) );
  XOR U366 ( .A(a[86]), .B(b[86]), .Z(n990) );
  NANDN U367 ( .A(n989), .B(n990), .Z(n177) );
  AND U368 ( .A(n178), .B(n177), .Z(n991) );
  XOR U369 ( .A(a[87]), .B(b[87]), .Z(n992) );
  NANDN U370 ( .A(n991), .B(n992), .Z(n179) );
  AND U371 ( .A(n180), .B(n179), .Z(n993) );
  XOR U372 ( .A(a[88]), .B(b[88]), .Z(n994) );
  NANDN U373 ( .A(n993), .B(n994), .Z(n181) );
  AND U374 ( .A(n182), .B(n181), .Z(n995) );
  XOR U375 ( .A(a[89]), .B(b[89]), .Z(n996) );
  NANDN U376 ( .A(n995), .B(n996), .Z(n183) );
  AND U377 ( .A(n184), .B(n183), .Z(n999) );
  XOR U378 ( .A(a[90]), .B(b[90]), .Z(n1000) );
  NANDN U379 ( .A(n999), .B(n1000), .Z(n185) );
  AND U380 ( .A(n186), .B(n185), .Z(n1001) );
  XOR U381 ( .A(a[91]), .B(b[91]), .Z(n1002) );
  NANDN U382 ( .A(n1001), .B(n1002), .Z(n187) );
  AND U383 ( .A(n188), .B(n187), .Z(n1003) );
  XOR U384 ( .A(a[92]), .B(b[92]), .Z(n1004) );
  NANDN U385 ( .A(n1003), .B(n1004), .Z(n189) );
  AND U386 ( .A(n190), .B(n189), .Z(n1005) );
  XOR U387 ( .A(a[93]), .B(b[93]), .Z(n1006) );
  NANDN U388 ( .A(n1005), .B(n1006), .Z(n191) );
  AND U389 ( .A(n192), .B(n191), .Z(n1007) );
  XOR U390 ( .A(a[94]), .B(b[94]), .Z(n1008) );
  NANDN U391 ( .A(n1007), .B(n1008), .Z(n193) );
  AND U392 ( .A(n194), .B(n193), .Z(n1009) );
  XOR U393 ( .A(a[95]), .B(b[95]), .Z(n1010) );
  NANDN U394 ( .A(n1009), .B(n1010), .Z(n195) );
  AND U395 ( .A(n196), .B(n195), .Z(n1011) );
  XOR U396 ( .A(a[96]), .B(b[96]), .Z(n1012) );
  NANDN U397 ( .A(n1011), .B(n1012), .Z(n197) );
  AND U398 ( .A(n198), .B(n197), .Z(n1013) );
  XOR U399 ( .A(a[97]), .B(b[97]), .Z(n1014) );
  NANDN U400 ( .A(n1013), .B(n1014), .Z(n199) );
  AND U401 ( .A(n200), .B(n199), .Z(n1015) );
  XOR U402 ( .A(a[98]), .B(b[98]), .Z(n1016) );
  NANDN U403 ( .A(n1015), .B(n1016), .Z(n201) );
  AND U404 ( .A(n202), .B(n201), .Z(n1017) );
  OR U405 ( .A(n1018), .B(n1017), .Z(n203) );
  AND U406 ( .A(n204), .B(n203), .Z(n206) );
  XNOR U407 ( .A(n205), .B(n206), .Z(c[100]) );
  XOR U408 ( .A(a[101]), .B(b[101]), .Z(n209) );
  NAND U409 ( .A(b[100]), .B(a[100]), .Z(n208) );
  NANDN U410 ( .A(n206), .B(n205), .Z(n207) );
  AND U411 ( .A(n208), .B(n207), .Z(n210) );
  XNOR U412 ( .A(n209), .B(n210), .Z(c[101]) );
  XOR U413 ( .A(a[102]), .B(b[102]), .Z(n213) );
  NAND U414 ( .A(b[101]), .B(a[101]), .Z(n212) );
  NANDN U415 ( .A(n210), .B(n209), .Z(n211) );
  AND U416 ( .A(n212), .B(n211), .Z(n214) );
  XNOR U417 ( .A(n213), .B(n214), .Z(c[102]) );
  XOR U418 ( .A(a[103]), .B(b[103]), .Z(n217) );
  NAND U419 ( .A(b[102]), .B(a[102]), .Z(n216) );
  NANDN U420 ( .A(n214), .B(n213), .Z(n215) );
  AND U421 ( .A(n216), .B(n215), .Z(n218) );
  XNOR U422 ( .A(n217), .B(n218), .Z(c[103]) );
  XOR U423 ( .A(a[104]), .B(b[104]), .Z(n221) );
  NAND U424 ( .A(b[103]), .B(a[103]), .Z(n220) );
  NANDN U425 ( .A(n218), .B(n217), .Z(n219) );
  AND U426 ( .A(n220), .B(n219), .Z(n222) );
  XNOR U427 ( .A(n221), .B(n222), .Z(c[104]) );
  XOR U428 ( .A(a[105]), .B(b[105]), .Z(n225) );
  NAND U429 ( .A(b[104]), .B(a[104]), .Z(n224) );
  NANDN U430 ( .A(n222), .B(n221), .Z(n223) );
  AND U431 ( .A(n224), .B(n223), .Z(n226) );
  XNOR U432 ( .A(n225), .B(n226), .Z(c[105]) );
  XOR U433 ( .A(a[106]), .B(b[106]), .Z(n229) );
  NAND U434 ( .A(b[105]), .B(a[105]), .Z(n228) );
  NANDN U435 ( .A(n226), .B(n225), .Z(n227) );
  AND U436 ( .A(n228), .B(n227), .Z(n230) );
  XNOR U437 ( .A(n229), .B(n230), .Z(c[106]) );
  XOR U438 ( .A(a[107]), .B(b[107]), .Z(n233) );
  NAND U439 ( .A(b[106]), .B(a[106]), .Z(n232) );
  NANDN U440 ( .A(n230), .B(n229), .Z(n231) );
  AND U441 ( .A(n232), .B(n231), .Z(n234) );
  XNOR U442 ( .A(n233), .B(n234), .Z(c[107]) );
  XOR U443 ( .A(a[108]), .B(b[108]), .Z(n237) );
  NAND U444 ( .A(b[107]), .B(a[107]), .Z(n236) );
  NANDN U445 ( .A(n234), .B(n233), .Z(n235) );
  AND U446 ( .A(n236), .B(n235), .Z(n238) );
  XNOR U447 ( .A(n237), .B(n238), .Z(c[108]) );
  XOR U448 ( .A(a[109]), .B(b[109]), .Z(n243) );
  NAND U449 ( .A(b[108]), .B(a[108]), .Z(n240) );
  NANDN U450 ( .A(n238), .B(n237), .Z(n239) );
  AND U451 ( .A(n240), .B(n239), .Z(n244) );
  XNOR U452 ( .A(n243), .B(n244), .Z(c[109]) );
  XNOR U453 ( .A(n242), .B(n241), .Z(c[10]) );
  XOR U454 ( .A(a[110]), .B(b[110]), .Z(n247) );
  NAND U455 ( .A(b[109]), .B(a[109]), .Z(n246) );
  NANDN U456 ( .A(n244), .B(n243), .Z(n245) );
  AND U457 ( .A(n246), .B(n245), .Z(n248) );
  XNOR U458 ( .A(n247), .B(n248), .Z(c[110]) );
  XOR U459 ( .A(a[111]), .B(b[111]), .Z(n251) );
  NAND U460 ( .A(b[110]), .B(a[110]), .Z(n250) );
  NANDN U461 ( .A(n248), .B(n247), .Z(n249) );
  AND U462 ( .A(n250), .B(n249), .Z(n252) );
  XNOR U463 ( .A(n251), .B(n252), .Z(c[111]) );
  XOR U464 ( .A(a[112]), .B(b[112]), .Z(n255) );
  NAND U465 ( .A(b[111]), .B(a[111]), .Z(n254) );
  NANDN U466 ( .A(n252), .B(n251), .Z(n253) );
  AND U467 ( .A(n254), .B(n253), .Z(n256) );
  XNOR U468 ( .A(n255), .B(n256), .Z(c[112]) );
  XOR U469 ( .A(a[113]), .B(b[113]), .Z(n259) );
  NAND U470 ( .A(b[112]), .B(a[112]), .Z(n258) );
  NANDN U471 ( .A(n256), .B(n255), .Z(n257) );
  AND U472 ( .A(n258), .B(n257), .Z(n260) );
  XNOR U473 ( .A(n259), .B(n260), .Z(c[113]) );
  XOR U474 ( .A(a[114]), .B(b[114]), .Z(n263) );
  NAND U475 ( .A(b[113]), .B(a[113]), .Z(n262) );
  NANDN U476 ( .A(n260), .B(n259), .Z(n261) );
  AND U477 ( .A(n262), .B(n261), .Z(n264) );
  XNOR U478 ( .A(n263), .B(n264), .Z(c[114]) );
  XOR U479 ( .A(a[115]), .B(b[115]), .Z(n267) );
  NAND U480 ( .A(b[114]), .B(a[114]), .Z(n266) );
  NANDN U481 ( .A(n264), .B(n263), .Z(n265) );
  AND U482 ( .A(n266), .B(n265), .Z(n268) );
  XNOR U483 ( .A(n267), .B(n268), .Z(c[115]) );
  XOR U484 ( .A(a[116]), .B(b[116]), .Z(n271) );
  NAND U485 ( .A(b[115]), .B(a[115]), .Z(n270) );
  NANDN U486 ( .A(n268), .B(n267), .Z(n269) );
  AND U487 ( .A(n270), .B(n269), .Z(n272) );
  XNOR U488 ( .A(n271), .B(n272), .Z(c[116]) );
  XOR U489 ( .A(a[117]), .B(b[117]), .Z(n275) );
  NAND U490 ( .A(b[116]), .B(a[116]), .Z(n274) );
  NANDN U491 ( .A(n272), .B(n271), .Z(n273) );
  AND U492 ( .A(n274), .B(n273), .Z(n276) );
  XNOR U493 ( .A(n275), .B(n276), .Z(c[117]) );
  XOR U494 ( .A(a[118]), .B(b[118]), .Z(n279) );
  NAND U495 ( .A(b[117]), .B(a[117]), .Z(n278) );
  NANDN U496 ( .A(n276), .B(n275), .Z(n277) );
  AND U497 ( .A(n278), .B(n277), .Z(n280) );
  XNOR U498 ( .A(n279), .B(n280), .Z(c[118]) );
  XOR U499 ( .A(a[119]), .B(b[119]), .Z(n285) );
  NAND U500 ( .A(b[118]), .B(a[118]), .Z(n282) );
  NANDN U501 ( .A(n280), .B(n279), .Z(n281) );
  AND U502 ( .A(n282), .B(n281), .Z(n286) );
  XNOR U503 ( .A(n285), .B(n286), .Z(c[119]) );
  XNOR U504 ( .A(n284), .B(n283), .Z(c[11]) );
  XOR U505 ( .A(a[120]), .B(b[120]), .Z(n289) );
  NAND U506 ( .A(b[119]), .B(a[119]), .Z(n288) );
  NANDN U507 ( .A(n286), .B(n285), .Z(n287) );
  AND U508 ( .A(n288), .B(n287), .Z(n290) );
  XNOR U509 ( .A(n289), .B(n290), .Z(c[120]) );
  XOR U510 ( .A(a[121]), .B(b[121]), .Z(n293) );
  NAND U511 ( .A(b[120]), .B(a[120]), .Z(n292) );
  NANDN U512 ( .A(n290), .B(n289), .Z(n291) );
  AND U513 ( .A(n292), .B(n291), .Z(n294) );
  XNOR U514 ( .A(n293), .B(n294), .Z(c[121]) );
  XOR U515 ( .A(a[122]), .B(b[122]), .Z(n297) );
  NAND U516 ( .A(b[121]), .B(a[121]), .Z(n296) );
  NANDN U517 ( .A(n294), .B(n293), .Z(n295) );
  AND U518 ( .A(n296), .B(n295), .Z(n298) );
  XNOR U519 ( .A(n297), .B(n298), .Z(c[122]) );
  XOR U520 ( .A(a[123]), .B(b[123]), .Z(n301) );
  NAND U521 ( .A(b[122]), .B(a[122]), .Z(n300) );
  NANDN U522 ( .A(n298), .B(n297), .Z(n299) );
  AND U523 ( .A(n300), .B(n299), .Z(n302) );
  XNOR U524 ( .A(n301), .B(n302), .Z(c[123]) );
  XOR U525 ( .A(a[124]), .B(b[124]), .Z(n305) );
  NAND U526 ( .A(b[123]), .B(a[123]), .Z(n304) );
  NANDN U527 ( .A(n302), .B(n301), .Z(n303) );
  AND U528 ( .A(n304), .B(n303), .Z(n306) );
  XNOR U529 ( .A(n305), .B(n306), .Z(c[124]) );
  XOR U530 ( .A(a[125]), .B(b[125]), .Z(n309) );
  NAND U531 ( .A(b[124]), .B(a[124]), .Z(n308) );
  NANDN U532 ( .A(n306), .B(n305), .Z(n307) );
  AND U533 ( .A(n308), .B(n307), .Z(n310) );
  XNOR U534 ( .A(n309), .B(n310), .Z(c[125]) );
  XOR U535 ( .A(a[126]), .B(b[126]), .Z(n313) );
  NAND U536 ( .A(b[125]), .B(a[125]), .Z(n312) );
  NANDN U537 ( .A(n310), .B(n309), .Z(n311) );
  AND U538 ( .A(n312), .B(n311), .Z(n314) );
  XNOR U539 ( .A(n313), .B(n314), .Z(c[126]) );
  XOR U540 ( .A(a[127]), .B(b[127]), .Z(n317) );
  NAND U541 ( .A(b[126]), .B(a[126]), .Z(n316) );
  NANDN U542 ( .A(n314), .B(n313), .Z(n315) );
  AND U543 ( .A(n316), .B(n315), .Z(n318) );
  XNOR U544 ( .A(n317), .B(n318), .Z(c[127]) );
  XOR U545 ( .A(a[128]), .B(b[128]), .Z(n321) );
  NAND U546 ( .A(b[127]), .B(a[127]), .Z(n320) );
  NANDN U547 ( .A(n318), .B(n317), .Z(n319) );
  AND U548 ( .A(n320), .B(n319), .Z(n322) );
  XNOR U549 ( .A(n321), .B(n322), .Z(c[128]) );
  XOR U550 ( .A(a[129]), .B(b[129]), .Z(n327) );
  NAND U551 ( .A(b[128]), .B(a[128]), .Z(n324) );
  NANDN U552 ( .A(n322), .B(n321), .Z(n323) );
  AND U553 ( .A(n324), .B(n323), .Z(n328) );
  XNOR U554 ( .A(n327), .B(n328), .Z(c[129]) );
  XNOR U555 ( .A(n326), .B(n325), .Z(c[12]) );
  XOR U556 ( .A(a[130]), .B(b[130]), .Z(n331) );
  NAND U557 ( .A(b[129]), .B(a[129]), .Z(n330) );
  NANDN U558 ( .A(n328), .B(n327), .Z(n329) );
  AND U559 ( .A(n330), .B(n329), .Z(n332) );
  XNOR U560 ( .A(n331), .B(n332), .Z(c[130]) );
  XOR U561 ( .A(a[131]), .B(b[131]), .Z(n335) );
  NAND U562 ( .A(b[130]), .B(a[130]), .Z(n334) );
  NANDN U563 ( .A(n332), .B(n331), .Z(n333) );
  AND U564 ( .A(n334), .B(n333), .Z(n336) );
  XNOR U565 ( .A(n335), .B(n336), .Z(c[131]) );
  XOR U566 ( .A(a[132]), .B(b[132]), .Z(n339) );
  NAND U567 ( .A(b[131]), .B(a[131]), .Z(n338) );
  NANDN U568 ( .A(n336), .B(n335), .Z(n337) );
  AND U569 ( .A(n338), .B(n337), .Z(n340) );
  XNOR U570 ( .A(n339), .B(n340), .Z(c[132]) );
  XOR U571 ( .A(a[133]), .B(b[133]), .Z(n343) );
  NAND U572 ( .A(b[132]), .B(a[132]), .Z(n342) );
  NANDN U573 ( .A(n340), .B(n339), .Z(n341) );
  AND U574 ( .A(n342), .B(n341), .Z(n344) );
  XNOR U575 ( .A(n343), .B(n344), .Z(c[133]) );
  XOR U576 ( .A(a[134]), .B(b[134]), .Z(n347) );
  NAND U577 ( .A(b[133]), .B(a[133]), .Z(n346) );
  NANDN U578 ( .A(n344), .B(n343), .Z(n345) );
  AND U579 ( .A(n346), .B(n345), .Z(n348) );
  XNOR U580 ( .A(n347), .B(n348), .Z(c[134]) );
  XOR U581 ( .A(a[135]), .B(b[135]), .Z(n351) );
  NAND U582 ( .A(b[134]), .B(a[134]), .Z(n350) );
  NANDN U583 ( .A(n348), .B(n347), .Z(n349) );
  AND U584 ( .A(n350), .B(n349), .Z(n352) );
  XNOR U585 ( .A(n351), .B(n352), .Z(c[135]) );
  XOR U586 ( .A(a[136]), .B(b[136]), .Z(n355) );
  NAND U587 ( .A(b[135]), .B(a[135]), .Z(n354) );
  NANDN U588 ( .A(n352), .B(n351), .Z(n353) );
  AND U589 ( .A(n354), .B(n353), .Z(n356) );
  XNOR U590 ( .A(n355), .B(n356), .Z(c[136]) );
  XOR U591 ( .A(a[137]), .B(b[137]), .Z(n359) );
  NAND U592 ( .A(b[136]), .B(a[136]), .Z(n358) );
  NANDN U593 ( .A(n356), .B(n355), .Z(n357) );
  AND U594 ( .A(n358), .B(n357), .Z(n360) );
  XNOR U595 ( .A(n359), .B(n360), .Z(c[137]) );
  XOR U596 ( .A(a[138]), .B(b[138]), .Z(n363) );
  NAND U597 ( .A(b[137]), .B(a[137]), .Z(n362) );
  NANDN U598 ( .A(n360), .B(n359), .Z(n361) );
  AND U599 ( .A(n362), .B(n361), .Z(n364) );
  XNOR U600 ( .A(n363), .B(n364), .Z(c[138]) );
  XOR U601 ( .A(a[139]), .B(b[139]), .Z(n369) );
  NAND U602 ( .A(b[138]), .B(a[138]), .Z(n366) );
  NANDN U603 ( .A(n364), .B(n363), .Z(n365) );
  AND U604 ( .A(n366), .B(n365), .Z(n370) );
  XNOR U605 ( .A(n369), .B(n370), .Z(c[139]) );
  XNOR U606 ( .A(n368), .B(n367), .Z(c[13]) );
  XOR U607 ( .A(a[140]), .B(b[140]), .Z(n373) );
  NAND U608 ( .A(b[139]), .B(a[139]), .Z(n372) );
  NANDN U609 ( .A(n370), .B(n369), .Z(n371) );
  AND U610 ( .A(n372), .B(n371), .Z(n374) );
  XNOR U611 ( .A(n373), .B(n374), .Z(c[140]) );
  XOR U612 ( .A(a[141]), .B(b[141]), .Z(n377) );
  NAND U613 ( .A(b[140]), .B(a[140]), .Z(n376) );
  NANDN U614 ( .A(n374), .B(n373), .Z(n375) );
  AND U615 ( .A(n376), .B(n375), .Z(n378) );
  XNOR U616 ( .A(n377), .B(n378), .Z(c[141]) );
  XOR U617 ( .A(a[142]), .B(b[142]), .Z(n381) );
  NAND U618 ( .A(b[141]), .B(a[141]), .Z(n380) );
  NANDN U619 ( .A(n378), .B(n377), .Z(n379) );
  AND U620 ( .A(n380), .B(n379), .Z(n382) );
  XNOR U621 ( .A(n381), .B(n382), .Z(c[142]) );
  XOR U622 ( .A(a[143]), .B(b[143]), .Z(n385) );
  NAND U623 ( .A(b[142]), .B(a[142]), .Z(n384) );
  NANDN U624 ( .A(n382), .B(n381), .Z(n383) );
  AND U625 ( .A(n384), .B(n383), .Z(n386) );
  XNOR U626 ( .A(n385), .B(n386), .Z(c[143]) );
  XOR U627 ( .A(a[144]), .B(b[144]), .Z(n389) );
  NAND U628 ( .A(b[143]), .B(a[143]), .Z(n388) );
  NANDN U629 ( .A(n386), .B(n385), .Z(n387) );
  AND U630 ( .A(n388), .B(n387), .Z(n390) );
  XNOR U631 ( .A(n389), .B(n390), .Z(c[144]) );
  XOR U632 ( .A(a[145]), .B(b[145]), .Z(n393) );
  NAND U633 ( .A(b[144]), .B(a[144]), .Z(n392) );
  NANDN U634 ( .A(n390), .B(n389), .Z(n391) );
  AND U635 ( .A(n392), .B(n391), .Z(n394) );
  XNOR U636 ( .A(n393), .B(n394), .Z(c[145]) );
  XOR U637 ( .A(a[146]), .B(b[146]), .Z(n397) );
  NAND U638 ( .A(b[145]), .B(a[145]), .Z(n396) );
  NANDN U639 ( .A(n394), .B(n393), .Z(n395) );
  AND U640 ( .A(n396), .B(n395), .Z(n398) );
  XNOR U641 ( .A(n397), .B(n398), .Z(c[146]) );
  XOR U642 ( .A(a[147]), .B(b[147]), .Z(n401) );
  NAND U643 ( .A(b[146]), .B(a[146]), .Z(n400) );
  NANDN U644 ( .A(n398), .B(n397), .Z(n399) );
  AND U645 ( .A(n400), .B(n399), .Z(n402) );
  XNOR U646 ( .A(n401), .B(n402), .Z(c[147]) );
  XOR U647 ( .A(a[148]), .B(b[148]), .Z(n405) );
  NAND U648 ( .A(b[147]), .B(a[147]), .Z(n404) );
  NANDN U649 ( .A(n402), .B(n401), .Z(n403) );
  AND U650 ( .A(n404), .B(n403), .Z(n406) );
  XNOR U651 ( .A(n405), .B(n406), .Z(c[148]) );
  XOR U652 ( .A(a[149]), .B(b[149]), .Z(n411) );
  NAND U653 ( .A(b[148]), .B(a[148]), .Z(n408) );
  NANDN U654 ( .A(n406), .B(n405), .Z(n407) );
  AND U655 ( .A(n408), .B(n407), .Z(n412) );
  XNOR U656 ( .A(n411), .B(n412), .Z(c[149]) );
  XNOR U657 ( .A(n410), .B(n409), .Z(c[14]) );
  XOR U658 ( .A(a[150]), .B(b[150]), .Z(n415) );
  NAND U659 ( .A(b[149]), .B(a[149]), .Z(n414) );
  NANDN U660 ( .A(n412), .B(n411), .Z(n413) );
  AND U661 ( .A(n414), .B(n413), .Z(n416) );
  XNOR U662 ( .A(n415), .B(n416), .Z(c[150]) );
  XOR U663 ( .A(a[151]), .B(b[151]), .Z(n419) );
  NAND U664 ( .A(b[150]), .B(a[150]), .Z(n418) );
  NANDN U665 ( .A(n416), .B(n415), .Z(n417) );
  AND U666 ( .A(n418), .B(n417), .Z(n420) );
  XNOR U667 ( .A(n419), .B(n420), .Z(c[151]) );
  XOR U668 ( .A(a[152]), .B(b[152]), .Z(n423) );
  NAND U669 ( .A(b[151]), .B(a[151]), .Z(n422) );
  NANDN U670 ( .A(n420), .B(n419), .Z(n421) );
  AND U671 ( .A(n422), .B(n421), .Z(n424) );
  XNOR U672 ( .A(n423), .B(n424), .Z(c[152]) );
  XOR U673 ( .A(a[153]), .B(b[153]), .Z(n427) );
  NAND U674 ( .A(b[152]), .B(a[152]), .Z(n426) );
  NANDN U675 ( .A(n424), .B(n423), .Z(n425) );
  AND U676 ( .A(n426), .B(n425), .Z(n428) );
  XNOR U677 ( .A(n427), .B(n428), .Z(c[153]) );
  XOR U678 ( .A(a[154]), .B(b[154]), .Z(n431) );
  NAND U679 ( .A(b[153]), .B(a[153]), .Z(n430) );
  NANDN U680 ( .A(n428), .B(n427), .Z(n429) );
  AND U681 ( .A(n430), .B(n429), .Z(n432) );
  XNOR U682 ( .A(n431), .B(n432), .Z(c[154]) );
  XOR U683 ( .A(a[155]), .B(b[155]), .Z(n435) );
  NAND U684 ( .A(b[154]), .B(a[154]), .Z(n434) );
  NANDN U685 ( .A(n432), .B(n431), .Z(n433) );
  AND U686 ( .A(n434), .B(n433), .Z(n436) );
  XNOR U687 ( .A(n435), .B(n436), .Z(c[155]) );
  XOR U688 ( .A(a[156]), .B(b[156]), .Z(n439) );
  NAND U689 ( .A(b[155]), .B(a[155]), .Z(n438) );
  NANDN U690 ( .A(n436), .B(n435), .Z(n437) );
  AND U691 ( .A(n438), .B(n437), .Z(n440) );
  XNOR U692 ( .A(n439), .B(n440), .Z(c[156]) );
  XOR U693 ( .A(a[157]), .B(b[157]), .Z(n443) );
  NAND U694 ( .A(b[156]), .B(a[156]), .Z(n442) );
  NANDN U695 ( .A(n440), .B(n439), .Z(n441) );
  AND U696 ( .A(n442), .B(n441), .Z(n444) );
  XNOR U697 ( .A(n443), .B(n444), .Z(c[157]) );
  XOR U698 ( .A(a[158]), .B(b[158]), .Z(n447) );
  NAND U699 ( .A(b[157]), .B(a[157]), .Z(n446) );
  NANDN U700 ( .A(n444), .B(n443), .Z(n445) );
  AND U701 ( .A(n446), .B(n445), .Z(n448) );
  XNOR U702 ( .A(n447), .B(n448), .Z(c[158]) );
  XOR U703 ( .A(a[159]), .B(b[159]), .Z(n453) );
  NAND U704 ( .A(b[158]), .B(a[158]), .Z(n450) );
  NANDN U705 ( .A(n448), .B(n447), .Z(n449) );
  AND U706 ( .A(n450), .B(n449), .Z(n454) );
  XNOR U707 ( .A(n453), .B(n454), .Z(c[159]) );
  XNOR U708 ( .A(n452), .B(n451), .Z(c[15]) );
  XOR U709 ( .A(a[160]), .B(b[160]), .Z(n457) );
  NAND U710 ( .A(b[159]), .B(a[159]), .Z(n456) );
  NANDN U711 ( .A(n454), .B(n453), .Z(n455) );
  AND U712 ( .A(n456), .B(n455), .Z(n458) );
  XNOR U713 ( .A(n457), .B(n458), .Z(c[160]) );
  XOR U714 ( .A(a[161]), .B(b[161]), .Z(n461) );
  NAND U715 ( .A(b[160]), .B(a[160]), .Z(n460) );
  NANDN U716 ( .A(n458), .B(n457), .Z(n459) );
  AND U717 ( .A(n460), .B(n459), .Z(n462) );
  XNOR U718 ( .A(n461), .B(n462), .Z(c[161]) );
  XOR U719 ( .A(a[162]), .B(b[162]), .Z(n465) );
  NAND U720 ( .A(b[161]), .B(a[161]), .Z(n464) );
  NANDN U721 ( .A(n462), .B(n461), .Z(n463) );
  AND U722 ( .A(n464), .B(n463), .Z(n466) );
  XNOR U723 ( .A(n465), .B(n466), .Z(c[162]) );
  XOR U724 ( .A(a[163]), .B(b[163]), .Z(n469) );
  NAND U725 ( .A(b[162]), .B(a[162]), .Z(n468) );
  NANDN U726 ( .A(n466), .B(n465), .Z(n467) );
  AND U727 ( .A(n468), .B(n467), .Z(n470) );
  XNOR U728 ( .A(n469), .B(n470), .Z(c[163]) );
  XOR U729 ( .A(a[164]), .B(b[164]), .Z(n473) );
  NAND U730 ( .A(b[163]), .B(a[163]), .Z(n472) );
  NANDN U731 ( .A(n470), .B(n469), .Z(n471) );
  AND U732 ( .A(n472), .B(n471), .Z(n474) );
  XNOR U733 ( .A(n473), .B(n474), .Z(c[164]) );
  XOR U734 ( .A(a[165]), .B(b[165]), .Z(n477) );
  NAND U735 ( .A(b[164]), .B(a[164]), .Z(n476) );
  NANDN U736 ( .A(n474), .B(n473), .Z(n475) );
  AND U737 ( .A(n476), .B(n475), .Z(n478) );
  XNOR U738 ( .A(n477), .B(n478), .Z(c[165]) );
  XOR U739 ( .A(a[166]), .B(b[166]), .Z(n481) );
  NAND U740 ( .A(b[165]), .B(a[165]), .Z(n480) );
  NANDN U741 ( .A(n478), .B(n477), .Z(n479) );
  AND U742 ( .A(n480), .B(n479), .Z(n482) );
  XNOR U743 ( .A(n481), .B(n482), .Z(c[166]) );
  XOR U744 ( .A(a[167]), .B(b[167]), .Z(n485) );
  NAND U745 ( .A(b[166]), .B(a[166]), .Z(n484) );
  NANDN U746 ( .A(n482), .B(n481), .Z(n483) );
  AND U747 ( .A(n484), .B(n483), .Z(n486) );
  XNOR U748 ( .A(n485), .B(n486), .Z(c[167]) );
  XOR U749 ( .A(a[168]), .B(b[168]), .Z(n489) );
  NAND U750 ( .A(b[167]), .B(a[167]), .Z(n488) );
  NANDN U751 ( .A(n486), .B(n485), .Z(n487) );
  AND U752 ( .A(n488), .B(n487), .Z(n490) );
  XNOR U753 ( .A(n489), .B(n490), .Z(c[168]) );
  XOR U754 ( .A(a[169]), .B(b[169]), .Z(n495) );
  NAND U755 ( .A(b[168]), .B(a[168]), .Z(n492) );
  NANDN U756 ( .A(n490), .B(n489), .Z(n491) );
  AND U757 ( .A(n492), .B(n491), .Z(n496) );
  XNOR U758 ( .A(n495), .B(n496), .Z(c[169]) );
  XNOR U759 ( .A(n494), .B(n493), .Z(c[16]) );
  XOR U760 ( .A(a[170]), .B(b[170]), .Z(n499) );
  NAND U761 ( .A(b[169]), .B(a[169]), .Z(n498) );
  NANDN U762 ( .A(n496), .B(n495), .Z(n497) );
  AND U763 ( .A(n498), .B(n497), .Z(n500) );
  XNOR U764 ( .A(n499), .B(n500), .Z(c[170]) );
  XOR U765 ( .A(a[171]), .B(b[171]), .Z(n503) );
  NAND U766 ( .A(b[170]), .B(a[170]), .Z(n502) );
  NANDN U767 ( .A(n500), .B(n499), .Z(n501) );
  AND U768 ( .A(n502), .B(n501), .Z(n504) );
  XNOR U769 ( .A(n503), .B(n504), .Z(c[171]) );
  XOR U770 ( .A(a[172]), .B(b[172]), .Z(n507) );
  NAND U771 ( .A(b[171]), .B(a[171]), .Z(n506) );
  NANDN U772 ( .A(n504), .B(n503), .Z(n505) );
  AND U773 ( .A(n506), .B(n505), .Z(n508) );
  XNOR U774 ( .A(n507), .B(n508), .Z(c[172]) );
  XOR U775 ( .A(a[173]), .B(b[173]), .Z(n511) );
  NAND U776 ( .A(b[172]), .B(a[172]), .Z(n510) );
  NANDN U777 ( .A(n508), .B(n507), .Z(n509) );
  AND U778 ( .A(n510), .B(n509), .Z(n512) );
  XNOR U779 ( .A(n511), .B(n512), .Z(c[173]) );
  XOR U780 ( .A(a[174]), .B(b[174]), .Z(n515) );
  NAND U781 ( .A(b[173]), .B(a[173]), .Z(n514) );
  NANDN U782 ( .A(n512), .B(n511), .Z(n513) );
  AND U783 ( .A(n514), .B(n513), .Z(n516) );
  XNOR U784 ( .A(n515), .B(n516), .Z(c[174]) );
  XOR U785 ( .A(a[175]), .B(b[175]), .Z(n519) );
  NAND U786 ( .A(b[174]), .B(a[174]), .Z(n518) );
  NANDN U787 ( .A(n516), .B(n515), .Z(n517) );
  AND U788 ( .A(n518), .B(n517), .Z(n520) );
  XNOR U789 ( .A(n519), .B(n520), .Z(c[175]) );
  XOR U790 ( .A(a[176]), .B(b[176]), .Z(n523) );
  NAND U791 ( .A(b[175]), .B(a[175]), .Z(n522) );
  NANDN U792 ( .A(n520), .B(n519), .Z(n521) );
  AND U793 ( .A(n522), .B(n521), .Z(n524) );
  XNOR U794 ( .A(n523), .B(n524), .Z(c[176]) );
  XOR U795 ( .A(a[177]), .B(b[177]), .Z(n527) );
  NAND U796 ( .A(b[176]), .B(a[176]), .Z(n526) );
  NANDN U797 ( .A(n524), .B(n523), .Z(n525) );
  AND U798 ( .A(n526), .B(n525), .Z(n528) );
  XNOR U799 ( .A(n527), .B(n528), .Z(c[177]) );
  XOR U800 ( .A(a[178]), .B(b[178]), .Z(n531) );
  NAND U801 ( .A(b[177]), .B(a[177]), .Z(n530) );
  NANDN U802 ( .A(n528), .B(n527), .Z(n529) );
  AND U803 ( .A(n530), .B(n529), .Z(n532) );
  XNOR U804 ( .A(n531), .B(n532), .Z(c[178]) );
  XOR U805 ( .A(a[179]), .B(b[179]), .Z(n537) );
  NAND U806 ( .A(b[178]), .B(a[178]), .Z(n534) );
  NANDN U807 ( .A(n532), .B(n531), .Z(n533) );
  AND U808 ( .A(n534), .B(n533), .Z(n538) );
  XNOR U809 ( .A(n537), .B(n538), .Z(c[179]) );
  XNOR U810 ( .A(n536), .B(n535), .Z(c[17]) );
  XOR U811 ( .A(a[180]), .B(b[180]), .Z(n541) );
  NAND U812 ( .A(b[179]), .B(a[179]), .Z(n540) );
  NANDN U813 ( .A(n538), .B(n537), .Z(n539) );
  AND U814 ( .A(n540), .B(n539), .Z(n542) );
  XNOR U815 ( .A(n541), .B(n542), .Z(c[180]) );
  XOR U816 ( .A(a[181]), .B(b[181]), .Z(n545) );
  NAND U817 ( .A(b[180]), .B(a[180]), .Z(n544) );
  NANDN U818 ( .A(n542), .B(n541), .Z(n543) );
  AND U819 ( .A(n544), .B(n543), .Z(n546) );
  XNOR U820 ( .A(n545), .B(n546), .Z(c[181]) );
  XOR U821 ( .A(a[182]), .B(b[182]), .Z(n549) );
  NAND U822 ( .A(b[181]), .B(a[181]), .Z(n548) );
  NANDN U823 ( .A(n546), .B(n545), .Z(n547) );
  AND U824 ( .A(n548), .B(n547), .Z(n550) );
  XNOR U825 ( .A(n549), .B(n550), .Z(c[182]) );
  XOR U826 ( .A(a[183]), .B(b[183]), .Z(n553) );
  NAND U827 ( .A(b[182]), .B(a[182]), .Z(n552) );
  NANDN U828 ( .A(n550), .B(n549), .Z(n551) );
  AND U829 ( .A(n552), .B(n551), .Z(n554) );
  XNOR U830 ( .A(n553), .B(n554), .Z(c[183]) );
  XOR U831 ( .A(a[184]), .B(b[184]), .Z(n557) );
  NAND U832 ( .A(b[183]), .B(a[183]), .Z(n556) );
  NANDN U833 ( .A(n554), .B(n553), .Z(n555) );
  AND U834 ( .A(n556), .B(n555), .Z(n558) );
  XNOR U835 ( .A(n557), .B(n558), .Z(c[184]) );
  XOR U836 ( .A(a[185]), .B(b[185]), .Z(n561) );
  NAND U837 ( .A(b[184]), .B(a[184]), .Z(n560) );
  NANDN U838 ( .A(n558), .B(n557), .Z(n559) );
  AND U839 ( .A(n560), .B(n559), .Z(n562) );
  XNOR U840 ( .A(n561), .B(n562), .Z(c[185]) );
  XOR U841 ( .A(a[186]), .B(b[186]), .Z(n565) );
  NAND U842 ( .A(b[185]), .B(a[185]), .Z(n564) );
  NANDN U843 ( .A(n562), .B(n561), .Z(n563) );
  AND U844 ( .A(n564), .B(n563), .Z(n566) );
  XNOR U845 ( .A(n565), .B(n566), .Z(c[186]) );
  XOR U846 ( .A(a[187]), .B(b[187]), .Z(n569) );
  NAND U847 ( .A(b[186]), .B(a[186]), .Z(n568) );
  NANDN U848 ( .A(n566), .B(n565), .Z(n567) );
  AND U849 ( .A(n568), .B(n567), .Z(n570) );
  XNOR U850 ( .A(n569), .B(n570), .Z(c[187]) );
  XOR U851 ( .A(a[188]), .B(b[188]), .Z(n573) );
  NAND U852 ( .A(b[187]), .B(a[187]), .Z(n572) );
  NANDN U853 ( .A(n570), .B(n569), .Z(n571) );
  AND U854 ( .A(n572), .B(n571), .Z(n574) );
  XNOR U855 ( .A(n573), .B(n574), .Z(c[188]) );
  XOR U856 ( .A(a[189]), .B(b[189]), .Z(n579) );
  NAND U857 ( .A(b[188]), .B(a[188]), .Z(n576) );
  NANDN U858 ( .A(n574), .B(n573), .Z(n575) );
  AND U859 ( .A(n576), .B(n575), .Z(n580) );
  XNOR U860 ( .A(n579), .B(n580), .Z(c[189]) );
  XNOR U861 ( .A(n578), .B(n577), .Z(c[18]) );
  XOR U862 ( .A(a[190]), .B(b[190]), .Z(n583) );
  NAND U863 ( .A(b[189]), .B(a[189]), .Z(n582) );
  NANDN U864 ( .A(n580), .B(n579), .Z(n581) );
  AND U865 ( .A(n582), .B(n581), .Z(n584) );
  XNOR U866 ( .A(n583), .B(n584), .Z(c[190]) );
  XOR U867 ( .A(a[191]), .B(b[191]), .Z(n587) );
  NAND U868 ( .A(b[190]), .B(a[190]), .Z(n586) );
  NANDN U869 ( .A(n584), .B(n583), .Z(n585) );
  AND U870 ( .A(n586), .B(n585), .Z(n588) );
  XNOR U871 ( .A(n587), .B(n588), .Z(c[191]) );
  XOR U872 ( .A(a[192]), .B(b[192]), .Z(n591) );
  NAND U873 ( .A(b[191]), .B(a[191]), .Z(n590) );
  NANDN U874 ( .A(n588), .B(n587), .Z(n589) );
  AND U875 ( .A(n590), .B(n589), .Z(n592) );
  XNOR U876 ( .A(n591), .B(n592), .Z(c[192]) );
  XOR U877 ( .A(a[193]), .B(b[193]), .Z(n595) );
  NAND U878 ( .A(b[192]), .B(a[192]), .Z(n594) );
  NANDN U879 ( .A(n592), .B(n591), .Z(n593) );
  AND U880 ( .A(n594), .B(n593), .Z(n596) );
  XNOR U881 ( .A(n595), .B(n596), .Z(c[193]) );
  XOR U882 ( .A(a[194]), .B(b[194]), .Z(n599) );
  NAND U883 ( .A(b[193]), .B(a[193]), .Z(n598) );
  NANDN U884 ( .A(n596), .B(n595), .Z(n597) );
  AND U885 ( .A(n598), .B(n597), .Z(n600) );
  XNOR U886 ( .A(n599), .B(n600), .Z(c[194]) );
  XOR U887 ( .A(a[195]), .B(b[195]), .Z(n603) );
  NAND U888 ( .A(b[194]), .B(a[194]), .Z(n602) );
  NANDN U889 ( .A(n600), .B(n599), .Z(n601) );
  AND U890 ( .A(n602), .B(n601), .Z(n604) );
  XNOR U891 ( .A(n603), .B(n604), .Z(c[195]) );
  XOR U892 ( .A(a[196]), .B(b[196]), .Z(n607) );
  NAND U893 ( .A(b[195]), .B(a[195]), .Z(n606) );
  NANDN U894 ( .A(n604), .B(n603), .Z(n605) );
  AND U895 ( .A(n606), .B(n605), .Z(n608) );
  XNOR U896 ( .A(n607), .B(n608), .Z(c[196]) );
  XOR U897 ( .A(a[197]), .B(b[197]), .Z(n611) );
  NAND U898 ( .A(b[196]), .B(a[196]), .Z(n610) );
  NANDN U899 ( .A(n608), .B(n607), .Z(n609) );
  AND U900 ( .A(n610), .B(n609), .Z(n612) );
  XNOR U901 ( .A(n611), .B(n612), .Z(c[197]) );
  XOR U902 ( .A(a[198]), .B(b[198]), .Z(n615) );
  NAND U903 ( .A(b[197]), .B(a[197]), .Z(n614) );
  NANDN U904 ( .A(n612), .B(n611), .Z(n613) );
  AND U905 ( .A(n614), .B(n613), .Z(n616) );
  XNOR U906 ( .A(n615), .B(n616), .Z(c[198]) );
  XOR U907 ( .A(a[199]), .B(b[199]), .Z(n623) );
  NAND U908 ( .A(b[198]), .B(a[198]), .Z(n618) );
  NANDN U909 ( .A(n616), .B(n615), .Z(n617) );
  AND U910 ( .A(n618), .B(n617), .Z(n624) );
  XNOR U911 ( .A(n623), .B(n624), .Z(c[199]) );
  XNOR U912 ( .A(n620), .B(n619), .Z(c[19]) );
  XNOR U913 ( .A(n622), .B(n621), .Z(c[1]) );
  XOR U914 ( .A(a[200]), .B(b[200]), .Z(n627) );
  NAND U915 ( .A(b[199]), .B(a[199]), .Z(n626) );
  NANDN U916 ( .A(n624), .B(n623), .Z(n625) );
  AND U917 ( .A(n626), .B(n625), .Z(n628) );
  XNOR U918 ( .A(n627), .B(n628), .Z(c[200]) );
  XOR U919 ( .A(a[201]), .B(b[201]), .Z(n631) );
  NAND U920 ( .A(b[200]), .B(a[200]), .Z(n630) );
  NANDN U921 ( .A(n628), .B(n627), .Z(n629) );
  AND U922 ( .A(n630), .B(n629), .Z(n632) );
  XNOR U923 ( .A(n631), .B(n632), .Z(c[201]) );
  XOR U924 ( .A(a[202]), .B(b[202]), .Z(n635) );
  NAND U925 ( .A(b[201]), .B(a[201]), .Z(n634) );
  NANDN U926 ( .A(n632), .B(n631), .Z(n633) );
  AND U927 ( .A(n634), .B(n633), .Z(n636) );
  XNOR U928 ( .A(n635), .B(n636), .Z(c[202]) );
  XOR U929 ( .A(a[203]), .B(b[203]), .Z(n639) );
  NAND U930 ( .A(b[202]), .B(a[202]), .Z(n638) );
  NANDN U931 ( .A(n636), .B(n635), .Z(n637) );
  AND U932 ( .A(n638), .B(n637), .Z(n640) );
  XNOR U933 ( .A(n639), .B(n640), .Z(c[203]) );
  XOR U934 ( .A(a[204]), .B(b[204]), .Z(n643) );
  NAND U935 ( .A(b[203]), .B(a[203]), .Z(n642) );
  NANDN U936 ( .A(n640), .B(n639), .Z(n641) );
  AND U937 ( .A(n642), .B(n641), .Z(n644) );
  XNOR U938 ( .A(n643), .B(n644), .Z(c[204]) );
  XOR U939 ( .A(a[205]), .B(b[205]), .Z(n647) );
  NAND U940 ( .A(b[204]), .B(a[204]), .Z(n646) );
  NANDN U941 ( .A(n644), .B(n643), .Z(n645) );
  AND U942 ( .A(n646), .B(n645), .Z(n648) );
  XNOR U943 ( .A(n647), .B(n648), .Z(c[205]) );
  XOR U944 ( .A(a[206]), .B(b[206]), .Z(n651) );
  NAND U945 ( .A(b[205]), .B(a[205]), .Z(n650) );
  NANDN U946 ( .A(n648), .B(n647), .Z(n649) );
  AND U947 ( .A(n650), .B(n649), .Z(n652) );
  XNOR U948 ( .A(n651), .B(n652), .Z(c[206]) );
  XOR U949 ( .A(a[207]), .B(b[207]), .Z(n655) );
  NAND U950 ( .A(b[206]), .B(a[206]), .Z(n654) );
  NANDN U951 ( .A(n652), .B(n651), .Z(n653) );
  AND U952 ( .A(n654), .B(n653), .Z(n656) );
  XNOR U953 ( .A(n655), .B(n656), .Z(c[207]) );
  XOR U954 ( .A(a[208]), .B(b[208]), .Z(n659) );
  NAND U955 ( .A(b[207]), .B(a[207]), .Z(n658) );
  NANDN U956 ( .A(n656), .B(n655), .Z(n657) );
  AND U957 ( .A(n658), .B(n657), .Z(n660) );
  XNOR U958 ( .A(n659), .B(n660), .Z(c[208]) );
  XOR U959 ( .A(a[209]), .B(b[209]), .Z(n665) );
  NAND U960 ( .A(b[208]), .B(a[208]), .Z(n662) );
  NANDN U961 ( .A(n660), .B(n659), .Z(n661) );
  AND U962 ( .A(n662), .B(n661), .Z(n666) );
  XNOR U963 ( .A(n665), .B(n666), .Z(c[209]) );
  XNOR U964 ( .A(n664), .B(n663), .Z(c[20]) );
  XOR U965 ( .A(a[210]), .B(b[210]), .Z(n669) );
  NAND U966 ( .A(b[209]), .B(a[209]), .Z(n668) );
  NANDN U967 ( .A(n666), .B(n665), .Z(n667) );
  AND U968 ( .A(n668), .B(n667), .Z(n670) );
  XNOR U969 ( .A(n669), .B(n670), .Z(c[210]) );
  XOR U970 ( .A(a[211]), .B(b[211]), .Z(n673) );
  NAND U971 ( .A(b[210]), .B(a[210]), .Z(n672) );
  NANDN U972 ( .A(n670), .B(n669), .Z(n671) );
  AND U973 ( .A(n672), .B(n671), .Z(n674) );
  XNOR U974 ( .A(n673), .B(n674), .Z(c[211]) );
  XOR U975 ( .A(a[212]), .B(b[212]), .Z(n677) );
  NAND U976 ( .A(b[211]), .B(a[211]), .Z(n676) );
  NANDN U977 ( .A(n674), .B(n673), .Z(n675) );
  AND U978 ( .A(n676), .B(n675), .Z(n678) );
  XNOR U979 ( .A(n677), .B(n678), .Z(c[212]) );
  XOR U980 ( .A(a[213]), .B(b[213]), .Z(n681) );
  NAND U981 ( .A(b[212]), .B(a[212]), .Z(n680) );
  NANDN U982 ( .A(n678), .B(n677), .Z(n679) );
  AND U983 ( .A(n680), .B(n679), .Z(n682) );
  XNOR U984 ( .A(n681), .B(n682), .Z(c[213]) );
  XOR U985 ( .A(a[214]), .B(b[214]), .Z(n685) );
  NAND U986 ( .A(b[213]), .B(a[213]), .Z(n684) );
  NANDN U987 ( .A(n682), .B(n681), .Z(n683) );
  AND U988 ( .A(n684), .B(n683), .Z(n686) );
  XNOR U989 ( .A(n685), .B(n686), .Z(c[214]) );
  XOR U990 ( .A(a[215]), .B(b[215]), .Z(n689) );
  NAND U991 ( .A(b[214]), .B(a[214]), .Z(n688) );
  NANDN U992 ( .A(n686), .B(n685), .Z(n687) );
  AND U993 ( .A(n688), .B(n687), .Z(n690) );
  XNOR U994 ( .A(n689), .B(n690), .Z(c[215]) );
  XOR U995 ( .A(a[216]), .B(b[216]), .Z(n693) );
  NAND U996 ( .A(b[215]), .B(a[215]), .Z(n692) );
  NANDN U997 ( .A(n690), .B(n689), .Z(n691) );
  AND U998 ( .A(n692), .B(n691), .Z(n694) );
  XNOR U999 ( .A(n693), .B(n694), .Z(c[216]) );
  XOR U1000 ( .A(a[217]), .B(b[217]), .Z(n697) );
  NAND U1001 ( .A(b[216]), .B(a[216]), .Z(n696) );
  NANDN U1002 ( .A(n694), .B(n693), .Z(n695) );
  AND U1003 ( .A(n696), .B(n695), .Z(n698) );
  XNOR U1004 ( .A(n697), .B(n698), .Z(c[217]) );
  XOR U1005 ( .A(a[218]), .B(b[218]), .Z(n701) );
  NAND U1006 ( .A(b[217]), .B(a[217]), .Z(n700) );
  NANDN U1007 ( .A(n698), .B(n697), .Z(n699) );
  AND U1008 ( .A(n700), .B(n699), .Z(n702) );
  XNOR U1009 ( .A(n701), .B(n702), .Z(c[218]) );
  XOR U1010 ( .A(a[219]), .B(b[219]), .Z(n707) );
  NAND U1011 ( .A(b[218]), .B(a[218]), .Z(n704) );
  NANDN U1012 ( .A(n702), .B(n701), .Z(n703) );
  AND U1013 ( .A(n704), .B(n703), .Z(n708) );
  XNOR U1014 ( .A(n707), .B(n708), .Z(c[219]) );
  XNOR U1015 ( .A(n706), .B(n705), .Z(c[21]) );
  XOR U1016 ( .A(a[220]), .B(b[220]), .Z(n711) );
  NAND U1017 ( .A(b[219]), .B(a[219]), .Z(n710) );
  NANDN U1018 ( .A(n708), .B(n707), .Z(n709) );
  AND U1019 ( .A(n710), .B(n709), .Z(n712) );
  XNOR U1020 ( .A(n711), .B(n712), .Z(c[220]) );
  XOR U1021 ( .A(a[221]), .B(b[221]), .Z(n715) );
  NAND U1022 ( .A(b[220]), .B(a[220]), .Z(n714) );
  NANDN U1023 ( .A(n712), .B(n711), .Z(n713) );
  AND U1024 ( .A(n714), .B(n713), .Z(n716) );
  XNOR U1025 ( .A(n715), .B(n716), .Z(c[221]) );
  XOR U1026 ( .A(a[222]), .B(b[222]), .Z(n719) );
  NAND U1027 ( .A(b[221]), .B(a[221]), .Z(n718) );
  NANDN U1028 ( .A(n716), .B(n715), .Z(n717) );
  AND U1029 ( .A(n718), .B(n717), .Z(n720) );
  XNOR U1030 ( .A(n719), .B(n720), .Z(c[222]) );
  XOR U1031 ( .A(a[223]), .B(b[223]), .Z(n723) );
  NAND U1032 ( .A(b[222]), .B(a[222]), .Z(n722) );
  NANDN U1033 ( .A(n720), .B(n719), .Z(n721) );
  AND U1034 ( .A(n722), .B(n721), .Z(n724) );
  XNOR U1035 ( .A(n723), .B(n724), .Z(c[223]) );
  XOR U1036 ( .A(a[224]), .B(b[224]), .Z(n727) );
  NAND U1037 ( .A(b[223]), .B(a[223]), .Z(n726) );
  NANDN U1038 ( .A(n724), .B(n723), .Z(n725) );
  AND U1039 ( .A(n726), .B(n725), .Z(n728) );
  XNOR U1040 ( .A(n727), .B(n728), .Z(c[224]) );
  XOR U1041 ( .A(a[225]), .B(b[225]), .Z(n731) );
  NAND U1042 ( .A(b[224]), .B(a[224]), .Z(n730) );
  NANDN U1043 ( .A(n728), .B(n727), .Z(n729) );
  AND U1044 ( .A(n730), .B(n729), .Z(n732) );
  XNOR U1045 ( .A(n731), .B(n732), .Z(c[225]) );
  XOR U1046 ( .A(a[226]), .B(b[226]), .Z(n735) );
  NAND U1047 ( .A(b[225]), .B(a[225]), .Z(n734) );
  NANDN U1048 ( .A(n732), .B(n731), .Z(n733) );
  AND U1049 ( .A(n734), .B(n733), .Z(n736) );
  XNOR U1050 ( .A(n735), .B(n736), .Z(c[226]) );
  XOR U1051 ( .A(a[227]), .B(b[227]), .Z(n739) );
  NAND U1052 ( .A(b[226]), .B(a[226]), .Z(n738) );
  NANDN U1053 ( .A(n736), .B(n735), .Z(n737) );
  AND U1054 ( .A(n738), .B(n737), .Z(n740) );
  XNOR U1055 ( .A(n739), .B(n740), .Z(c[227]) );
  XOR U1056 ( .A(a[228]), .B(b[228]), .Z(n743) );
  NAND U1057 ( .A(b[227]), .B(a[227]), .Z(n742) );
  NANDN U1058 ( .A(n740), .B(n739), .Z(n741) );
  AND U1059 ( .A(n742), .B(n741), .Z(n744) );
  XNOR U1060 ( .A(n743), .B(n744), .Z(c[228]) );
  XOR U1061 ( .A(a[229]), .B(b[229]), .Z(n749) );
  NAND U1062 ( .A(b[228]), .B(a[228]), .Z(n746) );
  NANDN U1063 ( .A(n744), .B(n743), .Z(n745) );
  AND U1064 ( .A(n746), .B(n745), .Z(n750) );
  XNOR U1065 ( .A(n749), .B(n750), .Z(c[229]) );
  XNOR U1066 ( .A(n748), .B(n747), .Z(c[22]) );
  XOR U1067 ( .A(a[230]), .B(b[230]), .Z(n753) );
  NAND U1068 ( .A(b[229]), .B(a[229]), .Z(n752) );
  NANDN U1069 ( .A(n750), .B(n749), .Z(n751) );
  AND U1070 ( .A(n752), .B(n751), .Z(n754) );
  XNOR U1071 ( .A(n753), .B(n754), .Z(c[230]) );
  XOR U1072 ( .A(a[231]), .B(b[231]), .Z(n757) );
  NAND U1073 ( .A(b[230]), .B(a[230]), .Z(n756) );
  NANDN U1074 ( .A(n754), .B(n753), .Z(n755) );
  AND U1075 ( .A(n756), .B(n755), .Z(n758) );
  XNOR U1076 ( .A(n757), .B(n758), .Z(c[231]) );
  XOR U1077 ( .A(a[232]), .B(b[232]), .Z(n761) );
  NAND U1078 ( .A(b[231]), .B(a[231]), .Z(n760) );
  NANDN U1079 ( .A(n758), .B(n757), .Z(n759) );
  AND U1080 ( .A(n760), .B(n759), .Z(n762) );
  XNOR U1081 ( .A(n761), .B(n762), .Z(c[232]) );
  XOR U1082 ( .A(a[233]), .B(b[233]), .Z(n765) );
  NAND U1083 ( .A(b[232]), .B(a[232]), .Z(n764) );
  NANDN U1084 ( .A(n762), .B(n761), .Z(n763) );
  AND U1085 ( .A(n764), .B(n763), .Z(n766) );
  XNOR U1086 ( .A(n765), .B(n766), .Z(c[233]) );
  XOR U1087 ( .A(a[234]), .B(b[234]), .Z(n769) );
  NAND U1088 ( .A(b[233]), .B(a[233]), .Z(n768) );
  NANDN U1089 ( .A(n766), .B(n765), .Z(n767) );
  AND U1090 ( .A(n768), .B(n767), .Z(n770) );
  XNOR U1091 ( .A(n769), .B(n770), .Z(c[234]) );
  XOR U1092 ( .A(a[235]), .B(b[235]), .Z(n773) );
  NAND U1093 ( .A(b[234]), .B(a[234]), .Z(n772) );
  NANDN U1094 ( .A(n770), .B(n769), .Z(n771) );
  AND U1095 ( .A(n772), .B(n771), .Z(n774) );
  XNOR U1096 ( .A(n773), .B(n774), .Z(c[235]) );
  XOR U1097 ( .A(a[236]), .B(b[236]), .Z(n777) );
  NAND U1098 ( .A(b[235]), .B(a[235]), .Z(n776) );
  NANDN U1099 ( .A(n774), .B(n773), .Z(n775) );
  AND U1100 ( .A(n776), .B(n775), .Z(n778) );
  XNOR U1101 ( .A(n777), .B(n778), .Z(c[236]) );
  XOR U1102 ( .A(a[237]), .B(b[237]), .Z(n781) );
  NAND U1103 ( .A(b[236]), .B(a[236]), .Z(n780) );
  NANDN U1104 ( .A(n778), .B(n777), .Z(n779) );
  AND U1105 ( .A(n780), .B(n779), .Z(n782) );
  XNOR U1106 ( .A(n781), .B(n782), .Z(c[237]) );
  XOR U1107 ( .A(a[238]), .B(b[238]), .Z(n785) );
  NAND U1108 ( .A(b[237]), .B(a[237]), .Z(n784) );
  NANDN U1109 ( .A(n782), .B(n781), .Z(n783) );
  AND U1110 ( .A(n784), .B(n783), .Z(n786) );
  XNOR U1111 ( .A(n785), .B(n786), .Z(c[238]) );
  XOR U1112 ( .A(a[239]), .B(b[239]), .Z(n791) );
  NAND U1113 ( .A(b[238]), .B(a[238]), .Z(n788) );
  NANDN U1114 ( .A(n786), .B(n785), .Z(n787) );
  AND U1115 ( .A(n788), .B(n787), .Z(n792) );
  XNOR U1116 ( .A(n791), .B(n792), .Z(c[239]) );
  XNOR U1117 ( .A(n790), .B(n789), .Z(c[23]) );
  XOR U1118 ( .A(a[240]), .B(b[240]), .Z(n795) );
  NAND U1119 ( .A(b[239]), .B(a[239]), .Z(n794) );
  NANDN U1120 ( .A(n792), .B(n791), .Z(n793) );
  AND U1121 ( .A(n794), .B(n793), .Z(n796) );
  XNOR U1122 ( .A(n795), .B(n796), .Z(c[240]) );
  XOR U1123 ( .A(a[241]), .B(b[241]), .Z(n799) );
  NAND U1124 ( .A(b[240]), .B(a[240]), .Z(n798) );
  NANDN U1125 ( .A(n796), .B(n795), .Z(n797) );
  AND U1126 ( .A(n798), .B(n797), .Z(n800) );
  XNOR U1127 ( .A(n799), .B(n800), .Z(c[241]) );
  XOR U1128 ( .A(a[242]), .B(b[242]), .Z(n803) );
  NAND U1129 ( .A(b[241]), .B(a[241]), .Z(n802) );
  NANDN U1130 ( .A(n800), .B(n799), .Z(n801) );
  AND U1131 ( .A(n802), .B(n801), .Z(n804) );
  XNOR U1132 ( .A(n803), .B(n804), .Z(c[242]) );
  XOR U1133 ( .A(a[243]), .B(b[243]), .Z(n807) );
  NAND U1134 ( .A(b[242]), .B(a[242]), .Z(n806) );
  NANDN U1135 ( .A(n804), .B(n803), .Z(n805) );
  AND U1136 ( .A(n806), .B(n805), .Z(n808) );
  XNOR U1137 ( .A(n807), .B(n808), .Z(c[243]) );
  XOR U1138 ( .A(a[244]), .B(b[244]), .Z(n811) );
  NAND U1139 ( .A(b[243]), .B(a[243]), .Z(n810) );
  NANDN U1140 ( .A(n808), .B(n807), .Z(n809) );
  AND U1141 ( .A(n810), .B(n809), .Z(n812) );
  XNOR U1142 ( .A(n811), .B(n812), .Z(c[244]) );
  XOR U1143 ( .A(a[245]), .B(b[245]), .Z(n815) );
  NAND U1144 ( .A(b[244]), .B(a[244]), .Z(n814) );
  NANDN U1145 ( .A(n812), .B(n811), .Z(n813) );
  AND U1146 ( .A(n814), .B(n813), .Z(n816) );
  XNOR U1147 ( .A(n815), .B(n816), .Z(c[245]) );
  XOR U1148 ( .A(a[246]), .B(b[246]), .Z(n819) );
  NAND U1149 ( .A(b[245]), .B(a[245]), .Z(n818) );
  NANDN U1150 ( .A(n816), .B(n815), .Z(n817) );
  AND U1151 ( .A(n818), .B(n817), .Z(n820) );
  XNOR U1152 ( .A(n819), .B(n820), .Z(c[246]) );
  XOR U1153 ( .A(a[247]), .B(b[247]), .Z(n823) );
  NAND U1154 ( .A(b[246]), .B(a[246]), .Z(n822) );
  NANDN U1155 ( .A(n820), .B(n819), .Z(n821) );
  AND U1156 ( .A(n822), .B(n821), .Z(n824) );
  XNOR U1157 ( .A(n823), .B(n824), .Z(c[247]) );
  XOR U1158 ( .A(a[248]), .B(b[248]), .Z(n827) );
  NAND U1159 ( .A(b[247]), .B(a[247]), .Z(n826) );
  NANDN U1160 ( .A(n824), .B(n823), .Z(n825) );
  AND U1161 ( .A(n826), .B(n825), .Z(n828) );
  XNOR U1162 ( .A(n827), .B(n828), .Z(c[248]) );
  XOR U1163 ( .A(a[249]), .B(b[249]), .Z(n833) );
  NAND U1164 ( .A(b[248]), .B(a[248]), .Z(n830) );
  NANDN U1165 ( .A(n828), .B(n827), .Z(n829) );
  AND U1166 ( .A(n830), .B(n829), .Z(n834) );
  XNOR U1167 ( .A(n833), .B(n834), .Z(c[249]) );
  XNOR U1168 ( .A(n832), .B(n831), .Z(c[24]) );
  XOR U1169 ( .A(a[250]), .B(b[250]), .Z(n837) );
  NAND U1170 ( .A(b[249]), .B(a[249]), .Z(n836) );
  NANDN U1171 ( .A(n834), .B(n833), .Z(n835) );
  AND U1172 ( .A(n836), .B(n835), .Z(n838) );
  XNOR U1173 ( .A(n837), .B(n838), .Z(c[250]) );
  XOR U1174 ( .A(a[251]), .B(b[251]), .Z(n841) );
  NAND U1175 ( .A(b[250]), .B(a[250]), .Z(n840) );
  NANDN U1176 ( .A(n838), .B(n837), .Z(n839) );
  AND U1177 ( .A(n840), .B(n839), .Z(n842) );
  XNOR U1178 ( .A(n841), .B(n842), .Z(c[251]) );
  XOR U1179 ( .A(a[252]), .B(b[252]), .Z(n845) );
  NAND U1180 ( .A(b[251]), .B(a[251]), .Z(n844) );
  NANDN U1181 ( .A(n842), .B(n841), .Z(n843) );
  AND U1182 ( .A(n844), .B(n843), .Z(n846) );
  XNOR U1183 ( .A(n845), .B(n846), .Z(c[252]) );
  XOR U1184 ( .A(a[253]), .B(b[253]), .Z(n849) );
  NAND U1185 ( .A(b[252]), .B(a[252]), .Z(n848) );
  NANDN U1186 ( .A(n846), .B(n845), .Z(n847) );
  AND U1187 ( .A(n848), .B(n847), .Z(n850) );
  XNOR U1188 ( .A(n849), .B(n850), .Z(c[253]) );
  NAND U1189 ( .A(b[253]), .B(a[253]), .Z(n852) );
  NANDN U1190 ( .A(n850), .B(n849), .Z(n851) );
  AND U1191 ( .A(n852), .B(n851), .Z(n854) );
  XOR U1192 ( .A(a[254]), .B(n854), .Z(n853) );
  XNOR U1193 ( .A(b[254]), .B(n853), .Z(c[254]) );
  XNOR U1194 ( .A(n856), .B(n855), .Z(c[25]) );
  XNOR U1195 ( .A(n858), .B(n857), .Z(c[26]) );
  XNOR U1196 ( .A(n860), .B(n859), .Z(c[27]) );
  XNOR U1197 ( .A(n862), .B(n861), .Z(c[28]) );
  XNOR U1198 ( .A(n864), .B(n863), .Z(c[29]) );
  XNOR U1199 ( .A(n866), .B(n865), .Z(c[2]) );
  XNOR U1200 ( .A(n868), .B(n867), .Z(c[30]) );
  XNOR U1201 ( .A(n870), .B(n869), .Z(c[31]) );
  XNOR U1202 ( .A(n872), .B(n871), .Z(c[32]) );
  XNOR U1203 ( .A(n874), .B(n873), .Z(c[33]) );
  XNOR U1204 ( .A(n876), .B(n875), .Z(c[34]) );
  XNOR U1205 ( .A(n878), .B(n877), .Z(c[35]) );
  XNOR U1206 ( .A(n880), .B(n879), .Z(c[36]) );
  XNOR U1207 ( .A(n882), .B(n881), .Z(c[37]) );
  XNOR U1208 ( .A(n884), .B(n883), .Z(c[38]) );
  XNOR U1209 ( .A(n886), .B(n885), .Z(c[39]) );
  XNOR U1210 ( .A(n888), .B(n887), .Z(c[3]) );
  XNOR U1211 ( .A(n890), .B(n889), .Z(c[40]) );
  XNOR U1212 ( .A(n892), .B(n891), .Z(c[41]) );
  XNOR U1213 ( .A(n894), .B(n893), .Z(c[42]) );
  XNOR U1214 ( .A(n896), .B(n895), .Z(c[43]) );
  XNOR U1215 ( .A(n898), .B(n897), .Z(c[44]) );
  XNOR U1216 ( .A(n900), .B(n899), .Z(c[45]) );
  XNOR U1217 ( .A(n902), .B(n901), .Z(c[46]) );
  XNOR U1218 ( .A(n904), .B(n903), .Z(c[47]) );
  XNOR U1219 ( .A(n906), .B(n905), .Z(c[48]) );
  XNOR U1220 ( .A(n908), .B(n907), .Z(c[49]) );
  XNOR U1221 ( .A(n910), .B(n909), .Z(c[4]) );
  XNOR U1222 ( .A(n912), .B(n911), .Z(c[50]) );
  XNOR U1223 ( .A(n914), .B(n913), .Z(c[51]) );
  XNOR U1224 ( .A(n916), .B(n915), .Z(c[52]) );
  XNOR U1225 ( .A(n918), .B(n917), .Z(c[53]) );
  XNOR U1226 ( .A(n920), .B(n919), .Z(c[54]) );
  XNOR U1227 ( .A(n922), .B(n921), .Z(c[55]) );
  XNOR U1228 ( .A(n924), .B(n923), .Z(c[56]) );
  XNOR U1229 ( .A(n926), .B(n925), .Z(c[57]) );
  XNOR U1230 ( .A(n928), .B(n927), .Z(c[58]) );
  XNOR U1231 ( .A(n930), .B(n929), .Z(c[59]) );
  XNOR U1232 ( .A(n932), .B(n931), .Z(c[5]) );
  XNOR U1233 ( .A(n934), .B(n933), .Z(c[60]) );
  XNOR U1234 ( .A(n936), .B(n935), .Z(c[61]) );
  XNOR U1235 ( .A(n938), .B(n937), .Z(c[62]) );
  XNOR U1236 ( .A(n940), .B(n939), .Z(c[63]) );
  XNOR U1237 ( .A(n942), .B(n941), .Z(c[64]) );
  XNOR U1238 ( .A(n944), .B(n943), .Z(c[65]) );
  XNOR U1239 ( .A(n946), .B(n945), .Z(c[66]) );
  XNOR U1240 ( .A(n948), .B(n947), .Z(c[67]) );
  XNOR U1241 ( .A(n950), .B(n949), .Z(c[68]) );
  XNOR U1242 ( .A(n952), .B(n951), .Z(c[69]) );
  XNOR U1243 ( .A(n954), .B(n953), .Z(c[6]) );
  XNOR U1244 ( .A(n956), .B(n955), .Z(c[70]) );
  XNOR U1245 ( .A(n958), .B(n957), .Z(c[71]) );
  XNOR U1246 ( .A(n960), .B(n959), .Z(c[72]) );
  XNOR U1247 ( .A(n962), .B(n961), .Z(c[73]) );
  XNOR U1248 ( .A(n964), .B(n963), .Z(c[74]) );
  XNOR U1249 ( .A(n966), .B(n965), .Z(c[75]) );
  XNOR U1250 ( .A(n968), .B(n967), .Z(c[76]) );
  XNOR U1251 ( .A(n970), .B(n969), .Z(c[77]) );
  XNOR U1252 ( .A(n972), .B(n971), .Z(c[78]) );
  XNOR U1253 ( .A(n974), .B(n973), .Z(c[79]) );
  XNOR U1254 ( .A(n976), .B(n975), .Z(c[7]) );
  XNOR U1255 ( .A(n978), .B(n977), .Z(c[80]) );
  XNOR U1256 ( .A(n980), .B(n979), .Z(c[81]) );
  XNOR U1257 ( .A(n982), .B(n981), .Z(c[82]) );
  XNOR U1258 ( .A(n984), .B(n983), .Z(c[83]) );
  XNOR U1259 ( .A(n986), .B(n985), .Z(c[84]) );
  XNOR U1260 ( .A(n988), .B(n987), .Z(c[85]) );
  XNOR U1261 ( .A(n990), .B(n989), .Z(c[86]) );
  XNOR U1262 ( .A(n992), .B(n991), .Z(c[87]) );
  XNOR U1263 ( .A(n994), .B(n993), .Z(c[88]) );
  XNOR U1264 ( .A(n996), .B(n995), .Z(c[89]) );
  XNOR U1265 ( .A(n998), .B(n997), .Z(c[8]) );
  XNOR U1266 ( .A(n1000), .B(n999), .Z(c[90]) );
  XNOR U1267 ( .A(n1002), .B(n1001), .Z(c[91]) );
  XNOR U1268 ( .A(n1004), .B(n1003), .Z(c[92]) );
  XNOR U1269 ( .A(n1006), .B(n1005), .Z(c[93]) );
  XNOR U1270 ( .A(n1008), .B(n1007), .Z(c[94]) );
  XNOR U1271 ( .A(n1010), .B(n1009), .Z(c[95]) );
  XNOR U1272 ( .A(n1012), .B(n1011), .Z(c[96]) );
  XNOR U1273 ( .A(n1014), .B(n1013), .Z(c[97]) );
  XNOR U1274 ( .A(n1016), .B(n1015), .Z(c[98]) );
  XOR U1275 ( .A(n1018), .B(n1017), .Z(c[99]) );
  XOR U1276 ( .A(n1020), .B(n1019), .Z(c[9]) );
endmodule

