
module hamming_N160_CC1 ( clk, rst, x, y, o );
  input [159:0] x;
  input [159:0] y;
  output [7:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795;

  XOR U161 ( .A(n267), .B(n265), .Z(n257) );
  MUX U162 ( .IN0(n604), .IN1(n606), .SEL(n605), .F(n1) );
  IV U163 ( .A(n1), .Z(n333) );
  MUX U164 ( .IN0(n699), .IN1(n701), .SEL(n700), .F(n2) );
  IV U165 ( .A(n2), .Z(n389) );
  MUX U166 ( .IN0(n420), .IN1(n418), .SEL(n419), .F(n3) );
  IV U167 ( .A(n3), .Z(n230) );
  MUX U168 ( .IN0(n695), .IN1(n693), .SEL(n694), .F(n687) );
  MUX U169 ( .IN0(n526), .IN1(n524), .SEL(n525), .F(n520) );
  MUX U170 ( .IN0(n506), .IN1(n504), .SEL(n505), .F(n498) );
  MUX U171 ( .IN0(n4), .IN1(n538), .SEL(n539), .F(n294) );
  IV U172 ( .A(n540), .Z(n4) );
  MUX U173 ( .IN0(n586), .IN1(n584), .SEL(n585), .F(n580) );
  MUX U174 ( .IN0(n451), .IN1(n449), .SEL(n450), .F(n5) );
  IV U175 ( .A(n5), .Z(n245) );
  MUX U176 ( .IN0(n438), .IN1(n436), .SEL(n437), .F(n432) );
  MUX U177 ( .IN0(n360), .IN1(n363), .SEL(n361), .F(n196) );
  XNOR U178 ( .A(n310), .B(n311), .Z(n177) );
  MUX U179 ( .IN0(n221), .IN1(n6), .SEL(n222), .F(n133) );
  IV U180 ( .A(n223), .Z(n6) );
  MUX U181 ( .IN0(n201), .IN1(n204), .SEL(n202), .F(n131) );
  MUX U182 ( .IN0(n15), .IN1(n192), .SEL(n190), .F(n183) );
  XNOR U183 ( .A(n168), .B(n169), .Z(n109) );
  MUX U184 ( .IN0(n105), .IN1(n108), .SEL(n106), .F(n99) );
  MUX U185 ( .IN0(n715), .IN1(n713), .SEL(n714), .F(n709) );
  XOR U186 ( .A(n388), .B(n387), .Z(n395) );
  MUX U187 ( .IN0(n669), .IN1(n667), .SEL(n668), .F(n663) );
  MUX U188 ( .IN0(n7), .IN1(n680), .SEL(n681), .F(n381) );
  IV U189 ( .A(n682), .Z(n7) );
  MUX U190 ( .IN0(n597), .IN1(n595), .SEL(n596), .F(n8) );
  IV U191 ( .A(n8), .Z(n331) );
  MUX U192 ( .IN0(n9), .IN1(n507), .SEL(n508), .F(n277) );
  IV U193 ( .A(n509), .Z(n9) );
  MUX U194 ( .IN0(n464), .IN1(n462), .SEL(n463), .F(n263) );
  MUX U195 ( .IN0(n10), .IN1(n587), .SEL(n588), .F(n322) );
  IV U196 ( .A(n589), .Z(n10) );
  MUX U197 ( .IN0(n493), .IN1(n495), .SEL(n494), .F(n11) );
  IV U198 ( .A(n11), .Z(n268) );
  MUX U199 ( .IN0(n22), .IN1(n384), .SEL(n383), .F(n12) );
  IV U200 ( .A(n12), .Z(n205) );
  MUX U201 ( .IN0(n245), .IN1(n13), .SEL(n246), .F(n145) );
  IV U202 ( .A(n247), .Z(n13) );
  MUX U203 ( .IN0(n14), .IN1(n426), .SEL(n427), .F(n231) );
  IV U204 ( .A(n428), .Z(n14) );
  MUX U205 ( .IN0(n26), .IN1(n341), .SEL(n340), .F(n15) );
  IV U206 ( .A(n15), .Z(n191) );
  MUX U207 ( .IN0(n50), .IN1(n288), .SEL(n286), .F(n281) );
  MUX U208 ( .IN0(n21), .IN1(n267), .SEL(n265), .F(n153) );
  MUX U209 ( .IN0(n29), .IN1(n318), .SEL(n316), .F(n309) );
  MUX U210 ( .IN0(n31), .IN1(n199), .SEL(n198), .F(n16) );
  IV U211 ( .A(n16), .Z(n119) );
  MUX U212 ( .IN0(n45), .IN1(n227), .SEL(n225), .F(n219) );
  MUX U213 ( .IN0(n193), .IN1(n196), .SEL(n194), .F(n118) );
  MUX U214 ( .IN0(n173), .IN1(n176), .SEL(n174), .F(n167) );
  MUX U215 ( .IN0(n128), .IN1(n131), .SEL(n129), .F(n124) );
  XNOR U216 ( .A(n100), .B(n101), .Z(n73) );
  MUX U217 ( .IN0(n76), .IN1(n78), .SEL(n77), .F(n65) );
  MUX U218 ( .IN0(n583), .IN1(n581), .SEL(n582), .F(n17) );
  IV U219 ( .A(n17), .Z(n321) );
  MUX U220 ( .IN0(n435), .IN1(n433), .SEL(n434), .F(n18) );
  IV U221 ( .A(n18), .Z(n237) );
  MUX U222 ( .IN0(n455), .IN1(n453), .SEL(n454), .F(n19) );
  IV U223 ( .A(n19), .Z(n250) );
  MUX U224 ( .IN0(n20), .IN1(n696), .SEL(n697), .F(n388) );
  IV U225 ( .A(n698), .Z(n20) );
  MUX U226 ( .IN0(n657), .IN1(n655), .SEL(n656), .F(n377) );
  MUX U227 ( .IN0(n620), .IN1(n618), .SEL(n619), .F(n614) );
  MUX U228 ( .IN0(n600), .IN1(n598), .SEL(n599), .F(n594) );
  MUX U229 ( .IN0(n636), .IN1(n634), .SEL(n635), .F(n630) );
  MUX U230 ( .IN0(n646), .IN1(n644), .SEL(n645), .F(n638) );
  MUX U231 ( .IN0(n482), .IN1(n480), .SEL(n481), .F(n21) );
  IV U232 ( .A(n21), .Z(n266) );
  MUX U233 ( .IN0(n559), .IN1(n557), .SEL(n558), .F(n553) );
  XOR U234 ( .A(n257), .B(n256), .Z(n280) );
  MUX U235 ( .IN0(n683), .IN1(n685), .SEL(n684), .F(n22) );
  IV U236 ( .A(n22), .Z(n382) );
  MUX U237 ( .IN0(n416), .IN1(n414), .SEL(n415), .F(n410) );
  MUX U238 ( .IN0(n46), .IN1(n399), .SEL(n397), .F(n392) );
  MUX U239 ( .IN0(n24), .IN1(n381), .SEL(n379), .F(n204) );
  XOR U240 ( .A(n297), .B(n296), .Z(n272) );
  MUX U241 ( .IN0(n228), .IN1(n231), .SEL(n229), .F(n135) );
  MUX U242 ( .IN0(n163), .IN1(n166), .SEL(n164), .F(n159) );
  MUX U243 ( .IN0(n23), .IN1(n429), .SEL(n591), .F(n323) );
  IV U244 ( .A(n590), .Z(n23) );
  XOR U245 ( .A(n158), .B(n157), .Z(n199) );
  MUX U246 ( .IN0(n143), .IN1(n146), .SEL(n144), .F(n138) );
  MUX U247 ( .IN0(n109), .IN1(n111), .SEL(n110), .F(n75) );
  MUX U248 ( .IN0(n84), .IN1(n87), .SEL(n85), .F(n80) );
  MUX U249 ( .IN0(n705), .IN1(n703), .SEL(n704), .F(n399) );
  XOR U250 ( .A(n688), .B(n689), .Z(n386) );
  MUX U251 ( .IN0(n674), .IN1(n672), .SEL(n673), .F(n24) );
  IV U252 ( .A(n24), .Z(n380) );
  MUX U253 ( .IN0(n25), .IN1(n601), .SEL(n602), .F(n332) );
  IV U254 ( .A(n603), .Z(n25) );
  MUX U255 ( .IN0(n613), .IN1(n611), .SEL(n612), .F(n26) );
  IV U256 ( .A(n26), .Z(n339) );
  MUX U257 ( .IN0(n624), .IN1(n622), .SEL(n623), .F(n359) );
  MUX U258 ( .IN0(n27), .IN1(n647), .SEL(n648), .F(n363) );
  IV U259 ( .A(n649), .Z(n27) );
  MUX U260 ( .IN0(n516), .IN1(n514), .SEL(n515), .F(n288) );
  MUX U261 ( .IN0(n510), .IN1(n512), .SEL(n511), .F(n28) );
  IV U262 ( .A(n28), .Z(n278) );
  MUX U263 ( .IN0(n549), .IN1(n547), .SEL(n548), .F(n307) );
  MUX U264 ( .IN0(n573), .IN1(n571), .SEL(n572), .F(n29) );
  IV U265 ( .A(n29), .Z(n317) );
  MUX U266 ( .IN0(n458), .IN1(n456), .SEL(n457), .F(n452) );
  MUX U267 ( .IN0(n389), .IN1(n30), .SEL(n390), .F(n209) );
  IV U268 ( .A(n391), .Z(n30) );
  MUX U269 ( .IN0(n274), .IN1(n277), .SEL(n275), .F(n166) );
  XOR U270 ( .A(n153), .B(n151), .Z(n162) );
  MUX U271 ( .IN0(n53), .IN1(n294), .SEL(n292), .F(n176) );
  MUX U272 ( .IN0(n319), .IN1(n322), .SEL(n320), .F(n179) );
  XOR U273 ( .A(n545), .B(n544), .Z(n495) );
  XOR U274 ( .A(n231), .B(n229), .Z(n223) );
  XOR U275 ( .A(n238), .B(n236), .Z(n247) );
  MUX U276 ( .IN0(n40), .IN1(n366), .SEL(n365), .F(n31) );
  IV U277 ( .A(n31), .Z(n197) );
  MUX U278 ( .IN0(n205), .IN1(n32), .SEL(n206), .F(n125) );
  IV U279 ( .A(n207), .Z(n32) );
  MUX U280 ( .IN0(n112), .IN1(n96), .SEL(n113), .F(n76) );
  MUX U281 ( .IN0(n140), .IN1(n33), .SEL(n141), .F(n90) );
  IV U282 ( .A(n142), .Z(n33) );
  MUX U283 ( .IN0(n115), .IN1(n118), .SEL(n116), .F(n87) );
  MUX U284 ( .IN0(n73), .IN1(n75), .SEL(n74), .F(n71) );
  MUX U285 ( .IN0(n569), .IN1(n567), .SEL(n568), .F(n34) );
  IV U286 ( .A(n34), .Z(n310) );
  MUX U287 ( .IN0(n708), .IN1(n706), .SEL(n707), .F(n35) );
  IV U288 ( .A(n35), .Z(n393) );
  MUX U289 ( .IN0(n610), .IN1(n608), .SEL(n609), .F(n347) );
  XOR U290 ( .A(n332), .B(n330), .Z(n341) );
  MUX U291 ( .IN0(n519), .IN1(n517), .SEL(n518), .F(n36) );
  IV U292 ( .A(n36), .Z(n282) );
  MUX U293 ( .IN0(n552), .IN1(n550), .SEL(n551), .F(n37) );
  IV U294 ( .A(n37), .Z(n299) );
  XOR U295 ( .A(n353), .B(n352), .Z(n337) );
  XOR U296 ( .A(n371), .B(n370), .Z(n391) );
  MUX U297 ( .IN0(n404), .IN1(n402), .SEL(n403), .F(n227) );
  MUX U298 ( .IN0(n448), .IN1(n446), .SEL(n447), .F(n251) );
  MUX U299 ( .IN0(n386), .IN1(n388), .SEL(n387), .F(n217) );
  XOR U300 ( .A(n204), .B(n202), .Z(n211) );
  XOR U301 ( .A(n196), .B(n194), .Z(n188) );
  MUX U302 ( .IN0(n278), .IN1(n38), .SEL(n279), .F(n160) );
  IV U303 ( .A(n280), .Z(n38) );
  MUX U304 ( .IN0(n295), .IN1(n39), .SEL(n296), .F(n168) );
  IV U305 ( .A(n297), .Z(n39) );
  MUX U306 ( .IN0(n650), .IN1(n652), .SEL(n651), .F(n40) );
  IV U307 ( .A(n40), .Z(n364) );
  MUX U308 ( .IN0(n41), .IN1(n444), .SEL(n443), .F(n239) );
  IV U309 ( .A(n442), .Z(n41) );
  MUX U310 ( .IN0(n235), .IN1(n238), .SEL(n236), .F(n146) );
  XOR U311 ( .A(n111), .B(n110), .Z(n104) );
  MUX U312 ( .IN0(n150), .IN1(n153), .SEL(n151), .F(n108) );
  MUX U313 ( .IN0(n323), .IN1(n232), .SEL(n324), .F(n180) );
  XOR U314 ( .A(n135), .B(n134), .Z(n142) );
  MUX U315 ( .IN0(n81), .IN1(n42), .SEL(n82), .F(n70) );
  IV U316 ( .A(n83), .Z(n42) );
  MUX U317 ( .IN0(n125), .IN1(n43), .SEL(n126), .F(n86) );
  IV U318 ( .A(n127), .Z(n43) );
  MUX U319 ( .IN0(n65), .IN1(n44), .SEL(n66), .F(n63) );
  IV U320 ( .A(n67), .Z(n44) );
  MUX U321 ( .IN0(n413), .IN1(n411), .SEL(n412), .F(n45) );
  IV U322 ( .A(n45), .Z(n226) );
  MUX U323 ( .IN0(n712), .IN1(n710), .SEL(n711), .F(n46) );
  IV U324 ( .A(n46), .Z(n398) );
  MUX U325 ( .IN0(n666), .IN1(n664), .SEL(n665), .F(n47) );
  IV U326 ( .A(n47), .Z(n376) );
  MUX U327 ( .IN0(n617), .IN1(n615), .SEL(n616), .F(n48) );
  IV U328 ( .A(n48), .Z(n346) );
  MUX U329 ( .IN0(n633), .IN1(n631), .SEL(n632), .F(n49) );
  IV U330 ( .A(n49), .Z(n358) );
  MUX U331 ( .IN0(n523), .IN1(n521), .SEL(n522), .F(n50) );
  IV U332 ( .A(n50), .Z(n287) );
  MUX U333 ( .IN0(n473), .IN1(n471), .SEL(n472), .F(n51) );
  IV U334 ( .A(n51), .Z(n262) );
  MUX U335 ( .IN0(n556), .IN1(n554), .SEL(n555), .F(n52) );
  IV U336 ( .A(n52), .Z(n306) );
  MUX U337 ( .IN0(n532), .IN1(n530), .SEL(n531), .F(n53) );
  IV U338 ( .A(n53), .Z(n293) );
  MUX U339 ( .IN0(n54), .IN1(n439), .SEL(n440), .F(n238) );
  IV U340 ( .A(n441), .Z(n54) );
  MUX U341 ( .IN0(n393), .IN1(n55), .SEL(n394), .F(n216) );
  IV U342 ( .A(n395), .Z(n55) );
  MUX U343 ( .IN0(n369), .IN1(n56), .SEL(n370), .F(n203) );
  IV U344 ( .A(n371), .Z(n56) );
  MUX U345 ( .IN0(n282), .IN1(n57), .SEL(n283), .F(n165) );
  IV U346 ( .A(n284), .Z(n57) );
  MUX U347 ( .IN0(n255), .IN1(n58), .SEL(n256), .F(n152) );
  IV U348 ( .A(n257), .Z(n58) );
  MUX U349 ( .IN0(n299), .IN1(n59), .SEL(n300), .F(n175) );
  IV U350 ( .A(n301), .Z(n59) );
  XOR U351 ( .A(n606), .B(n605), .Z(n685) );
  XOR U352 ( .A(n337), .B(n336), .Z(n384) );
  XOR U353 ( .A(n188), .B(n187), .Z(n207) );
  MUX U354 ( .IN0(n248), .IN1(n251), .SEL(n249), .F(n244) );
  MUX U355 ( .IN0(n209), .IN1(n60), .SEL(n210), .F(n130) );
  IV U356 ( .A(n211), .Z(n60) );
  XOR U357 ( .A(n118), .B(n116), .Z(n127) );
  MUX U358 ( .IN0(n160), .IN1(n61), .SEL(n161), .F(n107) );
  IV U359 ( .A(n162), .Z(n61) );
  MUX U360 ( .IN0(n177), .IN1(n179), .SEL(n178), .F(n111) );
  XOR U361 ( .A(n495), .B(n494), .Z(n652) );
  XOR U362 ( .A(n272), .B(n271), .Z(n366) );
  XOR U363 ( .A(n223), .B(n222), .Z(n243) );
  MUX U364 ( .IN0(n180), .IN1(n136), .SEL(n181), .F(n112) );
  MUX U365 ( .IN0(n133), .IN1(n62), .SEL(n134), .F(n94) );
  IV U366 ( .A(n135), .Z(n62) );
  MUX U367 ( .IN0(n68), .IN1(n71), .SEL(n69), .F(n64) );
  ANDN U368 ( .B(n63), .A(o[6]), .Z(o[7]) );
  XNOR U369 ( .A(n64), .B(n63), .Z(o[6]) );
  XNOR U370 ( .A(n67), .B(n66), .Z(o[5]) );
  XOR U371 ( .A(n72), .B(n71), .Z(n66) );
  XNOR U372 ( .A(n69), .B(n65), .Z(n72) );
  IV U373 ( .A(n79), .Z(n78) );
  XOR U374 ( .A(n80), .B(n68), .Z(n69) );
  IV U375 ( .A(n70), .Z(n68) );
  NANDN U376 ( .A(n88), .B(n79), .Z(n67) );
  XNOR U377 ( .A(n77), .B(n79), .Z(o[4]) );
  XOR U378 ( .A(n89), .B(n90), .Z(n79) );
  XOR U379 ( .A(n88), .B(n91), .Z(n89) );
  AND U380 ( .A(n92), .B(n93), .Z(n91) );
  XOR U381 ( .A(n90), .B(n94), .Z(n93) );
  OR U382 ( .A(n95), .B(n96), .Z(n88) );
  XOR U383 ( .A(n97), .B(n83), .Z(n77) );
  XNOR U384 ( .A(n75), .B(n98), .Z(n83) );
  IV U385 ( .A(n74), .Z(n98) );
  XOR U386 ( .A(n99), .B(n73), .Z(n74) );
  AND U387 ( .A(n102), .B(n103), .Z(n101) );
  XNOR U388 ( .A(n100), .B(n104), .Z(n102) );
  XNOR U389 ( .A(n82), .B(n76), .Z(n97) );
  XOR U390 ( .A(n114), .B(n87), .Z(n82) );
  XNOR U391 ( .A(n85), .B(n81), .Z(n114) );
  XOR U392 ( .A(n119), .B(n120), .Z(n81) );
  AND U393 ( .A(n121), .B(n122), .Z(n120) );
  XNOR U394 ( .A(n119), .B(n123), .Z(n122) );
  XOR U395 ( .A(n124), .B(n84), .Z(n85) );
  IV U396 ( .A(n86), .Z(n84) );
  XOR U397 ( .A(n113), .B(n96), .Z(o[3]) );
  XNOR U398 ( .A(n132), .B(n94), .Z(n96) );
  XOR U399 ( .A(n92), .B(n95), .Z(n132) );
  OR U400 ( .A(n136), .B(n137), .Z(n95) );
  XOR U401 ( .A(n138), .B(n139), .Z(n92) );
  IV U402 ( .A(n90), .Z(n139) );
  XOR U403 ( .A(n147), .B(n123), .Z(n113) );
  XNOR U404 ( .A(n104), .B(n148), .Z(n123) );
  IV U405 ( .A(n103), .Z(n148) );
  XOR U406 ( .A(n149), .B(n108), .Z(n103) );
  XNOR U407 ( .A(n106), .B(n100), .Z(n149) );
  XOR U408 ( .A(n154), .B(n155), .Z(n100) );
  AND U409 ( .A(n156), .B(n157), .Z(n155) );
  XNOR U410 ( .A(n154), .B(n158), .Z(n156) );
  XOR U411 ( .A(n159), .B(n105), .Z(n106) );
  IV U412 ( .A(n107), .Z(n105) );
  XOR U413 ( .A(n167), .B(n109), .Z(n110) );
  AND U414 ( .A(n170), .B(n171), .Z(n169) );
  XNOR U415 ( .A(n168), .B(n172), .Z(n170) );
  XNOR U416 ( .A(n121), .B(n112), .Z(n147) );
  XOR U417 ( .A(n182), .B(n127), .Z(n121) );
  XOR U418 ( .A(n183), .B(n115), .Z(n116) );
  IV U419 ( .A(n117), .Z(n115) );
  XOR U420 ( .A(n184), .B(n185), .Z(n117) );
  AND U421 ( .A(n186), .B(n187), .Z(n185) );
  XNOR U422 ( .A(n184), .B(n188), .Z(n186) );
  XNOR U423 ( .A(n126), .B(n119), .Z(n182) );
  XOR U424 ( .A(n200), .B(n131), .Z(n126) );
  XNOR U425 ( .A(n129), .B(n125), .Z(n200) );
  XOR U426 ( .A(n208), .B(n128), .Z(n129) );
  IV U427 ( .A(n130), .Z(n128) );
  XOR U428 ( .A(n212), .B(n213), .Z(n208) );
  AND U429 ( .A(n214), .B(n215), .Z(n213) );
  XNOR U430 ( .A(n216), .B(n217), .Z(n215) );
  XOR U431 ( .A(n181), .B(n136), .Z(o[2]) );
  XOR U432 ( .A(n218), .B(n142), .Z(n136) );
  XOR U433 ( .A(n219), .B(n220), .Z(n134) );
  IV U434 ( .A(n133), .Z(n220) );
  XOR U435 ( .A(n141), .B(n137), .Z(n218) );
  OR U436 ( .A(n232), .B(n233), .Z(n137) );
  XOR U437 ( .A(n234), .B(n146), .Z(n141) );
  XNOR U438 ( .A(n144), .B(n140), .Z(n234) );
  XOR U439 ( .A(n239), .B(n240), .Z(n140) );
  AND U440 ( .A(n241), .B(n242), .Z(n240) );
  XNOR U441 ( .A(n239), .B(n243), .Z(n242) );
  XOR U442 ( .A(n244), .B(n143), .Z(n144) );
  IV U443 ( .A(n145), .Z(n143) );
  XOR U444 ( .A(n252), .B(n199), .Z(n181) );
  XOR U445 ( .A(n253), .B(n162), .Z(n157) );
  XOR U446 ( .A(n254), .B(n150), .Z(n151) );
  IV U447 ( .A(n152), .Z(n150) );
  XOR U448 ( .A(n258), .B(n259), .Z(n254) );
  AND U449 ( .A(n260), .B(n261), .Z(n259) );
  XNOR U450 ( .A(n262), .B(n263), .Z(n261) );
  XNOR U451 ( .A(n161), .B(n154), .Z(n253) );
  XOR U452 ( .A(n268), .B(n269), .Z(n154) );
  AND U453 ( .A(n270), .B(n271), .Z(n269) );
  XNOR U454 ( .A(n268), .B(n272), .Z(n270) );
  XOR U455 ( .A(n273), .B(n166), .Z(n161) );
  XNOR U456 ( .A(n164), .B(n160), .Z(n273) );
  XOR U457 ( .A(n281), .B(n163), .Z(n164) );
  IV U458 ( .A(n165), .Z(n163) );
  XNOR U459 ( .A(n172), .B(n289), .Z(n158) );
  IV U460 ( .A(n171), .Z(n289) );
  XOR U461 ( .A(n290), .B(n176), .Z(n171) );
  XNOR U462 ( .A(n174), .B(n168), .Z(n290) );
  XOR U463 ( .A(n298), .B(n173), .Z(n174) );
  IV U464 ( .A(n175), .Z(n173) );
  XOR U465 ( .A(n302), .B(n303), .Z(n298) );
  AND U466 ( .A(n304), .B(n305), .Z(n303) );
  XNOR U467 ( .A(n306), .B(n307), .Z(n305) );
  XNOR U468 ( .A(n179), .B(n308), .Z(n172) );
  IV U469 ( .A(n178), .Z(n308) );
  XOR U470 ( .A(n309), .B(n177), .Z(n178) );
  AND U471 ( .A(n312), .B(n313), .Z(n311) );
  XNOR U472 ( .A(n310), .B(n314), .Z(n312) );
  XNOR U473 ( .A(n198), .B(n180), .Z(n252) );
  XOR U474 ( .A(n325), .B(n207), .Z(n198) );
  XOR U475 ( .A(n326), .B(n192), .Z(n187) );
  XOR U476 ( .A(n327), .B(n328), .Z(n192) );
  AND U477 ( .A(n329), .B(n330), .Z(n328) );
  XNOR U478 ( .A(n331), .B(n332), .Z(n329) );
  XNOR U479 ( .A(n190), .B(n184), .Z(n326) );
  XOR U480 ( .A(n333), .B(n334), .Z(n184) );
  AND U481 ( .A(n335), .B(n336), .Z(n334) );
  XNOR U482 ( .A(n333), .B(n337), .Z(n335) );
  XOR U483 ( .A(n338), .B(n189), .Z(n190) );
  IV U484 ( .A(n191), .Z(n189) );
  XOR U485 ( .A(n342), .B(n343), .Z(n338) );
  AND U486 ( .A(n344), .B(n345), .Z(n343) );
  XNOR U487 ( .A(n346), .B(n347), .Z(n345) );
  XOR U488 ( .A(n348), .B(n193), .Z(n194) );
  IV U489 ( .A(n195), .Z(n193) );
  XOR U490 ( .A(n349), .B(n350), .Z(n195) );
  AND U491 ( .A(n351), .B(n352), .Z(n350) );
  XNOR U492 ( .A(n349), .B(n353), .Z(n351) );
  XOR U493 ( .A(n354), .B(n355), .Z(n348) );
  AND U494 ( .A(n356), .B(n357), .Z(n355) );
  XNOR U495 ( .A(n358), .B(n359), .Z(n357) );
  XNOR U496 ( .A(n206), .B(n197), .Z(n325) );
  XOR U497 ( .A(n367), .B(n211), .Z(n206) );
  XOR U498 ( .A(n368), .B(n201), .Z(n202) );
  IV U499 ( .A(n203), .Z(n201) );
  XOR U500 ( .A(n372), .B(n373), .Z(n368) );
  AND U501 ( .A(n374), .B(n375), .Z(n373) );
  XNOR U502 ( .A(n376), .B(n377), .Z(n375) );
  XNOR U503 ( .A(n210), .B(n205), .Z(n367) );
  XOR U504 ( .A(n385), .B(n217), .Z(n210) );
  XNOR U505 ( .A(n214), .B(n209), .Z(n385) );
  XOR U506 ( .A(n392), .B(n212), .Z(n214) );
  IV U507 ( .A(n216), .Z(n212) );
  XOR U508 ( .A(n324), .B(n232), .Z(o[1]) );
  XOR U509 ( .A(n400), .B(n243), .Z(n232) );
  XOR U510 ( .A(n401), .B(n227), .Z(n222) );
  XNOR U511 ( .A(n225), .B(n221), .Z(n401) );
  XNOR U512 ( .A(n405), .B(n406), .Z(n221) );
  ANDN U513 ( .B(n407), .A(n408), .Z(n406) );
  XOR U514 ( .A(n405), .B(n409), .Z(n407) );
  XOR U515 ( .A(n410), .B(n224), .Z(n225) );
  IV U516 ( .A(n226), .Z(n224) );
  XOR U517 ( .A(n417), .B(n228), .Z(n229) );
  IV U518 ( .A(n230), .Z(n228) );
  XOR U519 ( .A(n421), .B(n422), .Z(n417) );
  ANDN U520 ( .B(n423), .A(n424), .Z(n422) );
  XOR U521 ( .A(n421), .B(n425), .Z(n423) );
  XOR U522 ( .A(n241), .B(n233), .Z(n400) );
  OR U523 ( .A(n429), .B(n430), .Z(n233) );
  XOR U524 ( .A(n431), .B(n247), .Z(n241) );
  XOR U525 ( .A(n432), .B(n235), .Z(n236) );
  IV U526 ( .A(n237), .Z(n235) );
  XNOR U527 ( .A(n246), .B(n239), .Z(n431) );
  XOR U528 ( .A(n445), .B(n251), .Z(n246) );
  XNOR U529 ( .A(n249), .B(n245), .Z(n445) );
  XOR U530 ( .A(n452), .B(n248), .Z(n249) );
  IV U531 ( .A(n250), .Z(n248) );
  XOR U532 ( .A(n459), .B(n366), .Z(n324) );
  XOR U533 ( .A(n460), .B(n280), .Z(n271) );
  XOR U534 ( .A(n461), .B(n263), .Z(n256) );
  XNOR U535 ( .A(n260), .B(n255), .Z(n461) );
  XNOR U536 ( .A(n465), .B(n466), .Z(n255) );
  ANDN U537 ( .B(n467), .A(n468), .Z(n466) );
  XOR U538 ( .A(n465), .B(n469), .Z(n467) );
  XOR U539 ( .A(n470), .B(n258), .Z(n260) );
  IV U540 ( .A(n262), .Z(n258) );
  XOR U541 ( .A(n474), .B(n475), .Z(n470) );
  ANDN U542 ( .B(n476), .A(n477), .Z(n475) );
  XOR U543 ( .A(n474), .B(n478), .Z(n476) );
  XOR U544 ( .A(n479), .B(n264), .Z(n265) );
  IV U545 ( .A(n266), .Z(n264) );
  XOR U546 ( .A(n483), .B(n484), .Z(n479) );
  ANDN U547 ( .B(n485), .A(n486), .Z(n484) );
  XOR U548 ( .A(n483), .B(n487), .Z(n485) );
  XOR U549 ( .A(n488), .B(n489), .Z(n267) );
  ANDN U550 ( .B(n490), .A(n491), .Z(n489) );
  XNOR U551 ( .A(n488), .B(n492), .Z(n490) );
  XNOR U552 ( .A(n279), .B(n268), .Z(n460) );
  XOR U553 ( .A(n496), .B(n284), .Z(n279) );
  XNOR U554 ( .A(n277), .B(n497), .Z(n284) );
  IV U555 ( .A(n275), .Z(n497) );
  XOR U556 ( .A(n498), .B(n274), .Z(n275) );
  IV U557 ( .A(n276), .Z(n274) );
  XNOR U558 ( .A(n499), .B(n500), .Z(n276) );
  ANDN U559 ( .B(n501), .A(n502), .Z(n500) );
  XOR U560 ( .A(n499), .B(n503), .Z(n501) );
  XNOR U561 ( .A(n283), .B(n278), .Z(n496) );
  XOR U562 ( .A(n513), .B(n288), .Z(n283) );
  XNOR U563 ( .A(n286), .B(n282), .Z(n513) );
  XOR U564 ( .A(n520), .B(n285), .Z(n286) );
  IV U565 ( .A(n287), .Z(n285) );
  XOR U566 ( .A(n527), .B(n301), .Z(n296) );
  XNOR U567 ( .A(n294), .B(n528), .Z(n301) );
  IV U568 ( .A(n292), .Z(n528) );
  XOR U569 ( .A(n529), .B(n291), .Z(n292) );
  IV U570 ( .A(n293), .Z(n291) );
  XOR U571 ( .A(n533), .B(n534), .Z(n529) );
  ANDN U572 ( .B(n535), .A(n536), .Z(n534) );
  XOR U573 ( .A(n533), .B(n537), .Z(n535) );
  XNOR U574 ( .A(n300), .B(n295), .Z(n527) );
  XNOR U575 ( .A(n541), .B(n542), .Z(n295) );
  AND U576 ( .A(n543), .B(n544), .Z(n542) );
  XOR U577 ( .A(n541), .B(n545), .Z(n543) );
  XOR U578 ( .A(n546), .B(n307), .Z(n300) );
  XNOR U579 ( .A(n304), .B(n299), .Z(n546) );
  XOR U580 ( .A(n553), .B(n302), .Z(n304) );
  IV U581 ( .A(n306), .Z(n302) );
  XNOR U582 ( .A(n314), .B(n560), .Z(n297) );
  IV U583 ( .A(n313), .Z(n560) );
  XOR U584 ( .A(n561), .B(n318), .Z(n313) );
  XOR U585 ( .A(n562), .B(n563), .Z(n318) );
  ANDN U586 ( .B(n564), .A(n565), .Z(n563) );
  XOR U587 ( .A(n562), .B(n566), .Z(n564) );
  XNOR U588 ( .A(n316), .B(n310), .Z(n561) );
  XOR U589 ( .A(n570), .B(n315), .Z(n316) );
  IV U590 ( .A(n317), .Z(n315) );
  XOR U591 ( .A(n574), .B(n575), .Z(n570) );
  ANDN U592 ( .B(n576), .A(n577), .Z(n575) );
  XOR U593 ( .A(n574), .B(n578), .Z(n576) );
  XNOR U594 ( .A(n322), .B(n579), .Z(n314) );
  IV U595 ( .A(n320), .Z(n579) );
  XOR U596 ( .A(n580), .B(n319), .Z(n320) );
  IV U597 ( .A(n321), .Z(n319) );
  XNOR U598 ( .A(n365), .B(n323), .Z(n459) );
  XOR U599 ( .A(n592), .B(n384), .Z(n365) );
  XOR U600 ( .A(n593), .B(n341), .Z(n336) );
  XOR U601 ( .A(n594), .B(n327), .Z(n330) );
  IV U602 ( .A(n331), .Z(n327) );
  XNOR U603 ( .A(n340), .B(n333), .Z(n593) );
  XOR U604 ( .A(n607), .B(n347), .Z(n340) );
  XNOR U605 ( .A(n344), .B(n339), .Z(n607) );
  XOR U606 ( .A(n614), .B(n342), .Z(n344) );
  IV U607 ( .A(n346), .Z(n342) );
  XOR U608 ( .A(n621), .B(n359), .Z(n352) );
  XNOR U609 ( .A(n356), .B(n349), .Z(n621) );
  XNOR U610 ( .A(n625), .B(n626), .Z(n349) );
  ANDN U611 ( .B(n627), .A(n628), .Z(n626) );
  XOR U612 ( .A(n625), .B(n629), .Z(n627) );
  XOR U613 ( .A(n630), .B(n354), .Z(n356) );
  IV U614 ( .A(n358), .Z(n354) );
  XNOR U615 ( .A(n363), .B(n637), .Z(n353) );
  IV U616 ( .A(n361), .Z(n637) );
  XOR U617 ( .A(n638), .B(n360), .Z(n361) );
  IV U618 ( .A(n362), .Z(n360) );
  XNOR U619 ( .A(n639), .B(n640), .Z(n362) );
  ANDN U620 ( .B(n641), .A(n642), .Z(n640) );
  XOR U621 ( .A(n639), .B(n643), .Z(n641) );
  XNOR U622 ( .A(n383), .B(n364), .Z(n592) );
  XOR U623 ( .A(n653), .B(n391), .Z(n383) );
  XOR U624 ( .A(n654), .B(n377), .Z(n370) );
  XNOR U625 ( .A(n374), .B(n369), .Z(n654) );
  XNOR U626 ( .A(n658), .B(n659), .Z(n369) );
  ANDN U627 ( .B(n660), .A(n661), .Z(n659) );
  XOR U628 ( .A(n658), .B(n662), .Z(n660) );
  XOR U629 ( .A(n663), .B(n372), .Z(n374) );
  IV U630 ( .A(n376), .Z(n372) );
  XNOR U631 ( .A(n381), .B(n670), .Z(n371) );
  IV U632 ( .A(n379), .Z(n670) );
  XOR U633 ( .A(n671), .B(n378), .Z(n379) );
  IV U634 ( .A(n380), .Z(n378) );
  XOR U635 ( .A(n675), .B(n676), .Z(n671) );
  ANDN U636 ( .B(n677), .A(n678), .Z(n676) );
  XOR U637 ( .A(n675), .B(n679), .Z(n677) );
  XNOR U638 ( .A(n390), .B(n382), .Z(n653) );
  XOR U639 ( .A(n686), .B(n395), .Z(n390) );
  XOR U640 ( .A(n687), .B(n386), .Z(n387) );
  ANDN U641 ( .B(n690), .A(n691), .Z(n689) );
  XOR U642 ( .A(n688), .B(n692), .Z(n690) );
  XNOR U643 ( .A(n394), .B(n389), .Z(n686) );
  XOR U644 ( .A(n702), .B(n399), .Z(n394) );
  XNOR U645 ( .A(n397), .B(n393), .Z(n702) );
  XOR U646 ( .A(n709), .B(n396), .Z(n397) );
  IV U647 ( .A(n398), .Z(n396) );
  XOR U648 ( .A(n591), .B(n429), .Z(o[0]) );
  XNOR U649 ( .A(n716), .B(n444), .Z(n429) );
  XOR U650 ( .A(n409), .B(n408), .Z(n444) );
  XNOR U651 ( .A(n717), .B(n413), .Z(n408) );
  XNOR U652 ( .A(n404), .B(n403), .Z(n413) );
  XNOR U653 ( .A(n718), .B(n402), .Z(n403) );
  XNOR U654 ( .A(y[12]), .B(x[12]), .Z(n402) );
  XNOR U655 ( .A(y[13]), .B(x[13]), .Z(n718) );
  XNOR U656 ( .A(y[14]), .B(x[14]), .Z(n404) );
  XNOR U657 ( .A(n412), .B(n405), .Z(n717) );
  XNOR U658 ( .A(y[3]), .B(x[3]), .Z(n405) );
  XNOR U659 ( .A(n719), .B(n416), .Z(n412) );
  XNOR U660 ( .A(y[17]), .B(x[17]), .Z(n416) );
  XNOR U661 ( .A(n415), .B(n411), .Z(n719) );
  XNOR U662 ( .A(y[11]), .B(x[11]), .Z(n411) );
  XNOR U663 ( .A(n720), .B(n414), .Z(n415) );
  XNOR U664 ( .A(y[15]), .B(x[15]), .Z(n414) );
  XNOR U665 ( .A(y[16]), .B(x[16]), .Z(n720) );
  XNOR U666 ( .A(n420), .B(n419), .Z(n409) );
  XNOR U667 ( .A(n721), .B(n425), .Z(n419) );
  XNOR U668 ( .A(y[10]), .B(x[10]), .Z(n425) );
  XNOR U669 ( .A(n424), .B(n418), .Z(n721) );
  XNOR U670 ( .A(y[4]), .B(x[4]), .Z(n418) );
  XNOR U671 ( .A(n722), .B(n421), .Z(n424) );
  XNOR U672 ( .A(y[8]), .B(x[8]), .Z(n421) );
  XNOR U673 ( .A(y[9]), .B(x[9]), .Z(n722) );
  XOR U674 ( .A(n428), .B(n427), .Z(n420) );
  XNOR U675 ( .A(n723), .B(n426), .Z(n427) );
  XNOR U676 ( .A(y[5]), .B(x[5]), .Z(n426) );
  XNOR U677 ( .A(y[6]), .B(x[6]), .Z(n723) );
  XOR U678 ( .A(y[7]), .B(x[7]), .Z(n428) );
  XOR U679 ( .A(n443), .B(n430), .Z(n716) );
  XNOR U680 ( .A(y[1]), .B(x[1]), .Z(n430) );
  XOR U681 ( .A(n724), .B(n451), .Z(n443) );
  XNOR U682 ( .A(n435), .B(n434), .Z(n451) );
  XNOR U683 ( .A(n725), .B(n438), .Z(n434) );
  XNOR U684 ( .A(y[25]), .B(x[25]), .Z(n438) );
  XNOR U685 ( .A(n437), .B(n433), .Z(n725) );
  XNOR U686 ( .A(y[19]), .B(x[19]), .Z(n433) );
  XNOR U687 ( .A(n726), .B(n436), .Z(n437) );
  XNOR U688 ( .A(y[23]), .B(x[23]), .Z(n436) );
  XNOR U689 ( .A(y[24]), .B(x[24]), .Z(n726) );
  XOR U690 ( .A(n441), .B(n440), .Z(n435) );
  XNOR U691 ( .A(n727), .B(n439), .Z(n440) );
  XNOR U692 ( .A(y[20]), .B(x[20]), .Z(n439) );
  XNOR U693 ( .A(y[21]), .B(x[21]), .Z(n727) );
  XOR U694 ( .A(y[22]), .B(x[22]), .Z(n441) );
  XNOR U695 ( .A(n450), .B(n442), .Z(n724) );
  XNOR U696 ( .A(y[2]), .B(x[2]), .Z(n442) );
  XNOR U697 ( .A(n728), .B(n455), .Z(n450) );
  XNOR U698 ( .A(n448), .B(n447), .Z(n455) );
  XNOR U699 ( .A(n729), .B(n446), .Z(n447) );
  XNOR U700 ( .A(y[27]), .B(x[27]), .Z(n446) );
  XNOR U701 ( .A(y[28]), .B(x[28]), .Z(n729) );
  XNOR U702 ( .A(y[29]), .B(x[29]), .Z(n448) );
  XNOR U703 ( .A(n454), .B(n449), .Z(n728) );
  XNOR U704 ( .A(y[18]), .B(x[18]), .Z(n449) );
  XNOR U705 ( .A(n730), .B(n458), .Z(n454) );
  XNOR U706 ( .A(y[32]), .B(x[32]), .Z(n458) );
  XNOR U707 ( .A(n457), .B(n453), .Z(n730) );
  XNOR U708 ( .A(y[26]), .B(x[26]), .Z(n453) );
  XNOR U709 ( .A(n731), .B(n456), .Z(n457) );
  XNOR U710 ( .A(y[30]), .B(x[30]), .Z(n456) );
  XNOR U711 ( .A(y[31]), .B(x[31]), .Z(n731) );
  XOR U712 ( .A(n732), .B(n652), .Z(n591) );
  XOR U713 ( .A(n733), .B(n512), .Z(n494) );
  XNOR U714 ( .A(n469), .B(n468), .Z(n512) );
  XNOR U715 ( .A(n734), .B(n473), .Z(n468) );
  XNOR U716 ( .A(n464), .B(n463), .Z(n473) );
  XNOR U717 ( .A(n735), .B(n462), .Z(n463) );
  XNOR U718 ( .A(y[76]), .B(x[76]), .Z(n462) );
  XNOR U719 ( .A(y[77]), .B(x[77]), .Z(n735) );
  XNOR U720 ( .A(y[78]), .B(x[78]), .Z(n464) );
  XNOR U721 ( .A(n472), .B(n465), .Z(n734) );
  XNOR U722 ( .A(y[67]), .B(x[67]), .Z(n465) );
  XNOR U723 ( .A(n736), .B(n478), .Z(n472) );
  XNOR U724 ( .A(y[81]), .B(x[81]), .Z(n478) );
  XNOR U725 ( .A(n477), .B(n471), .Z(n736) );
  XNOR U726 ( .A(y[75]), .B(x[75]), .Z(n471) );
  XNOR U727 ( .A(n737), .B(n474), .Z(n477) );
  XNOR U728 ( .A(y[79]), .B(x[79]), .Z(n474) );
  XNOR U729 ( .A(y[80]), .B(x[80]), .Z(n737) );
  XNOR U730 ( .A(n482), .B(n481), .Z(n469) );
  XNOR U731 ( .A(n738), .B(n487), .Z(n481) );
  XNOR U732 ( .A(y[74]), .B(x[74]), .Z(n487) );
  XNOR U733 ( .A(n486), .B(n480), .Z(n738) );
  XNOR U734 ( .A(y[68]), .B(x[68]), .Z(n480) );
  XNOR U735 ( .A(n739), .B(n483), .Z(n486) );
  XNOR U736 ( .A(y[72]), .B(x[72]), .Z(n483) );
  XNOR U737 ( .A(y[73]), .B(x[73]), .Z(n739) );
  XOR U738 ( .A(n492), .B(n491), .Z(n482) );
  XNOR U739 ( .A(n740), .B(n488), .Z(n491) );
  XNOR U740 ( .A(y[69]), .B(x[69]), .Z(n488) );
  XNOR U741 ( .A(y[70]), .B(x[70]), .Z(n740) );
  XOR U742 ( .A(y[71]), .B(x[71]), .Z(n492) );
  XOR U743 ( .A(n511), .B(n493), .Z(n733) );
  XNOR U744 ( .A(y[34]), .B(x[34]), .Z(n493) );
  XOR U745 ( .A(n741), .B(n519), .Z(n511) );
  XNOR U746 ( .A(n503), .B(n502), .Z(n519) );
  XNOR U747 ( .A(n742), .B(n506), .Z(n502) );
  XNOR U748 ( .A(y[89]), .B(x[89]), .Z(n506) );
  XNOR U749 ( .A(n505), .B(n499), .Z(n742) );
  XNOR U750 ( .A(y[83]), .B(x[83]), .Z(n499) );
  XNOR U751 ( .A(n743), .B(n504), .Z(n505) );
  XNOR U752 ( .A(y[87]), .B(x[87]), .Z(n504) );
  XNOR U753 ( .A(y[88]), .B(x[88]), .Z(n743) );
  XOR U754 ( .A(n509), .B(n508), .Z(n503) );
  XNOR U755 ( .A(n744), .B(n507), .Z(n508) );
  XNOR U756 ( .A(y[84]), .B(x[84]), .Z(n507) );
  XNOR U757 ( .A(y[85]), .B(x[85]), .Z(n744) );
  XOR U758 ( .A(y[86]), .B(x[86]), .Z(n509) );
  XNOR U759 ( .A(n518), .B(n510), .Z(n741) );
  XNOR U760 ( .A(y[66]), .B(x[66]), .Z(n510) );
  XNOR U761 ( .A(n745), .B(n523), .Z(n518) );
  XNOR U762 ( .A(n516), .B(n515), .Z(n523) );
  XNOR U763 ( .A(n746), .B(n514), .Z(n515) );
  XNOR U764 ( .A(y[91]), .B(x[91]), .Z(n514) );
  XNOR U765 ( .A(y[92]), .B(x[92]), .Z(n746) );
  XNOR U766 ( .A(y[93]), .B(x[93]), .Z(n516) );
  XNOR U767 ( .A(n522), .B(n517), .Z(n745) );
  XNOR U768 ( .A(y[82]), .B(x[82]), .Z(n517) );
  XNOR U769 ( .A(n747), .B(n526), .Z(n522) );
  XNOR U770 ( .A(y[96]), .B(x[96]), .Z(n526) );
  XNOR U771 ( .A(n525), .B(n521), .Z(n747) );
  XNOR U772 ( .A(y[90]), .B(x[90]), .Z(n521) );
  XNOR U773 ( .A(n748), .B(n524), .Z(n525) );
  XNOR U774 ( .A(y[94]), .B(x[94]), .Z(n524) );
  XNOR U775 ( .A(y[95]), .B(x[95]), .Z(n748) );
  XOR U776 ( .A(n749), .B(n552), .Z(n544) );
  XNOR U777 ( .A(n532), .B(n531), .Z(n552) );
  XNOR U778 ( .A(n750), .B(n537), .Z(n531) );
  XNOR U779 ( .A(y[58]), .B(x[58]), .Z(n537) );
  XNOR U780 ( .A(n536), .B(n530), .Z(n750) );
  XNOR U781 ( .A(y[52]), .B(x[52]), .Z(n530) );
  XNOR U782 ( .A(n751), .B(n533), .Z(n536) );
  XNOR U783 ( .A(y[56]), .B(x[56]), .Z(n533) );
  XNOR U784 ( .A(y[57]), .B(x[57]), .Z(n751) );
  XOR U785 ( .A(n540), .B(n539), .Z(n532) );
  XNOR U786 ( .A(n752), .B(n538), .Z(n539) );
  XNOR U787 ( .A(y[53]), .B(x[53]), .Z(n538) );
  XNOR U788 ( .A(y[54]), .B(x[54]), .Z(n752) );
  XOR U789 ( .A(y[55]), .B(x[55]), .Z(n540) );
  XNOR U790 ( .A(n551), .B(n541), .Z(n749) );
  XNOR U791 ( .A(y[35]), .B(x[35]), .Z(n541) );
  XNOR U792 ( .A(n753), .B(n556), .Z(n551) );
  XNOR U793 ( .A(n549), .B(n548), .Z(n556) );
  XNOR U794 ( .A(n754), .B(n547), .Z(n548) );
  XNOR U795 ( .A(y[60]), .B(x[60]), .Z(n547) );
  XNOR U796 ( .A(y[61]), .B(x[61]), .Z(n754) );
  XNOR U797 ( .A(y[62]), .B(x[62]), .Z(n549) );
  XNOR U798 ( .A(n555), .B(n550), .Z(n753) );
  XNOR U799 ( .A(y[51]), .B(x[51]), .Z(n550) );
  XNOR U800 ( .A(n755), .B(n559), .Z(n555) );
  XNOR U801 ( .A(y[65]), .B(x[65]), .Z(n559) );
  XNOR U802 ( .A(n558), .B(n554), .Z(n755) );
  XNOR U803 ( .A(y[59]), .B(x[59]), .Z(n554) );
  XNOR U804 ( .A(n756), .B(n557), .Z(n558) );
  XNOR U805 ( .A(y[63]), .B(x[63]), .Z(n557) );
  XNOR U806 ( .A(y[64]), .B(x[64]), .Z(n756) );
  XNOR U807 ( .A(n569), .B(n568), .Z(n545) );
  XNOR U808 ( .A(n757), .B(n573), .Z(n568) );
  XNOR U809 ( .A(n566), .B(n565), .Z(n573) );
  XNOR U810 ( .A(n758), .B(n562), .Z(n565) );
  XNOR U811 ( .A(y[45]), .B(x[45]), .Z(n562) );
  XNOR U812 ( .A(y[46]), .B(x[46]), .Z(n758) );
  XNOR U813 ( .A(y[47]), .B(x[47]), .Z(n566) );
  XNOR U814 ( .A(n572), .B(n567), .Z(n757) );
  XNOR U815 ( .A(y[36]), .B(x[36]), .Z(n567) );
  XNOR U816 ( .A(n759), .B(n578), .Z(n572) );
  XNOR U817 ( .A(y[50]), .B(x[50]), .Z(n578) );
  XNOR U818 ( .A(n577), .B(n571), .Z(n759) );
  XNOR U819 ( .A(y[44]), .B(x[44]), .Z(n571) );
  XNOR U820 ( .A(n760), .B(n574), .Z(n577) );
  XNOR U821 ( .A(y[48]), .B(x[48]), .Z(n574) );
  XNOR U822 ( .A(y[49]), .B(x[49]), .Z(n760) );
  XNOR U823 ( .A(n583), .B(n582), .Z(n569) );
  XNOR U824 ( .A(n761), .B(n586), .Z(n582) );
  XNOR U825 ( .A(y[43]), .B(x[43]), .Z(n586) );
  XNOR U826 ( .A(n585), .B(n581), .Z(n761) );
  XNOR U827 ( .A(y[37]), .B(x[37]), .Z(n581) );
  XNOR U828 ( .A(n762), .B(n584), .Z(n585) );
  XNOR U829 ( .A(y[41]), .B(x[41]), .Z(n584) );
  XNOR U830 ( .A(y[42]), .B(x[42]), .Z(n762) );
  XOR U831 ( .A(n589), .B(n588), .Z(n583) );
  XNOR U832 ( .A(n763), .B(n587), .Z(n588) );
  XNOR U833 ( .A(y[38]), .B(x[38]), .Z(n587) );
  XNOR U834 ( .A(y[39]), .B(x[39]), .Z(n763) );
  XOR U835 ( .A(y[40]), .B(x[40]), .Z(n589) );
  XOR U836 ( .A(n651), .B(n590), .Z(n732) );
  XNOR U837 ( .A(y[0]), .B(x[0]), .Z(n590) );
  XOR U838 ( .A(n764), .B(n685), .Z(n651) );
  XOR U839 ( .A(n765), .B(n613), .Z(n605) );
  XNOR U840 ( .A(n597), .B(n596), .Z(n613) );
  XNOR U841 ( .A(n766), .B(n600), .Z(n596) );
  XNOR U842 ( .A(y[121]), .B(x[121]), .Z(n600) );
  XNOR U843 ( .A(n599), .B(n595), .Z(n766) );
  XNOR U844 ( .A(y[115]), .B(x[115]), .Z(n595) );
  XNOR U845 ( .A(n767), .B(n598), .Z(n599) );
  XNOR U846 ( .A(y[119]), .B(x[119]), .Z(n598) );
  XNOR U847 ( .A(y[120]), .B(x[120]), .Z(n767) );
  XOR U848 ( .A(n603), .B(n602), .Z(n597) );
  XNOR U849 ( .A(n768), .B(n601), .Z(n602) );
  XNOR U850 ( .A(y[116]), .B(x[116]), .Z(n601) );
  XNOR U851 ( .A(y[117]), .B(x[117]), .Z(n768) );
  XOR U852 ( .A(y[118]), .B(x[118]), .Z(n603) );
  XNOR U853 ( .A(n612), .B(n604), .Z(n765) );
  XNOR U854 ( .A(y[98]), .B(x[98]), .Z(n604) );
  XNOR U855 ( .A(n769), .B(n617), .Z(n612) );
  XNOR U856 ( .A(n610), .B(n609), .Z(n617) );
  XNOR U857 ( .A(n770), .B(n608), .Z(n609) );
  XNOR U858 ( .A(y[123]), .B(x[123]), .Z(n608) );
  XNOR U859 ( .A(y[124]), .B(x[124]), .Z(n770) );
  XNOR U860 ( .A(y[125]), .B(x[125]), .Z(n610) );
  XNOR U861 ( .A(n616), .B(n611), .Z(n769) );
  XNOR U862 ( .A(y[114]), .B(x[114]), .Z(n611) );
  XNOR U863 ( .A(n771), .B(n620), .Z(n616) );
  XNOR U864 ( .A(y[128]), .B(x[128]), .Z(n620) );
  XNOR U865 ( .A(n619), .B(n615), .Z(n771) );
  XNOR U866 ( .A(y[122]), .B(x[122]), .Z(n615) );
  XNOR U867 ( .A(n772), .B(n618), .Z(n619) );
  XNOR U868 ( .A(y[126]), .B(x[126]), .Z(n618) );
  XNOR U869 ( .A(y[127]), .B(x[127]), .Z(n772) );
  XNOR U870 ( .A(n629), .B(n628), .Z(n606) );
  XNOR U871 ( .A(n773), .B(n633), .Z(n628) );
  XNOR U872 ( .A(n624), .B(n623), .Z(n633) );
  XNOR U873 ( .A(n774), .B(n622), .Z(n623) );
  XNOR U874 ( .A(y[108]), .B(x[108]), .Z(n622) );
  XNOR U875 ( .A(y[109]), .B(x[109]), .Z(n774) );
  XNOR U876 ( .A(y[110]), .B(x[110]), .Z(n624) );
  XNOR U877 ( .A(n632), .B(n625), .Z(n773) );
  XNOR U878 ( .A(y[99]), .B(x[99]), .Z(n625) );
  XNOR U879 ( .A(n775), .B(n636), .Z(n632) );
  XNOR U880 ( .A(y[113]), .B(x[113]), .Z(n636) );
  XNOR U881 ( .A(n635), .B(n631), .Z(n775) );
  XNOR U882 ( .A(y[107]), .B(x[107]), .Z(n631) );
  XNOR U883 ( .A(n776), .B(n634), .Z(n635) );
  XNOR U884 ( .A(y[111]), .B(x[111]), .Z(n634) );
  XNOR U885 ( .A(y[112]), .B(x[112]), .Z(n776) );
  XNOR U886 ( .A(n643), .B(n642), .Z(n629) );
  XNOR U887 ( .A(n777), .B(n646), .Z(n642) );
  XNOR U888 ( .A(y[106]), .B(x[106]), .Z(n646) );
  XNOR U889 ( .A(n645), .B(n639), .Z(n777) );
  XNOR U890 ( .A(y[100]), .B(x[100]), .Z(n639) );
  XNOR U891 ( .A(n778), .B(n644), .Z(n645) );
  XNOR U892 ( .A(y[104]), .B(x[104]), .Z(n644) );
  XNOR U893 ( .A(y[105]), .B(x[105]), .Z(n778) );
  XOR U894 ( .A(n649), .B(n648), .Z(n643) );
  XNOR U895 ( .A(n779), .B(n647), .Z(n648) );
  XNOR U896 ( .A(y[101]), .B(x[101]), .Z(n647) );
  XNOR U897 ( .A(y[102]), .B(x[102]), .Z(n779) );
  XOR U898 ( .A(y[103]), .B(x[103]), .Z(n649) );
  XOR U899 ( .A(n684), .B(n650), .Z(n764) );
  XNOR U900 ( .A(y[33]), .B(x[33]), .Z(n650) );
  XOR U901 ( .A(n780), .B(n701), .Z(n684) );
  XNOR U902 ( .A(n662), .B(n661), .Z(n701) );
  XNOR U903 ( .A(n781), .B(n666), .Z(n661) );
  XNOR U904 ( .A(n657), .B(n656), .Z(n666) );
  XNOR U905 ( .A(n782), .B(n655), .Z(n656) );
  XNOR U906 ( .A(y[139]), .B(x[139]), .Z(n655) );
  XNOR U907 ( .A(y[140]), .B(x[140]), .Z(n782) );
  XNOR U908 ( .A(y[141]), .B(x[141]), .Z(n657) );
  XNOR U909 ( .A(n665), .B(n658), .Z(n781) );
  XNOR U910 ( .A(y[130]), .B(x[130]), .Z(n658) );
  XNOR U911 ( .A(n783), .B(n669), .Z(n665) );
  XNOR U912 ( .A(y[144]), .B(x[144]), .Z(n669) );
  XNOR U913 ( .A(n668), .B(n664), .Z(n783) );
  XNOR U914 ( .A(y[138]), .B(x[138]), .Z(n664) );
  XNOR U915 ( .A(n784), .B(n667), .Z(n668) );
  XNOR U916 ( .A(y[142]), .B(x[142]), .Z(n667) );
  XNOR U917 ( .A(y[143]), .B(x[143]), .Z(n784) );
  XNOR U918 ( .A(n674), .B(n673), .Z(n662) );
  XNOR U919 ( .A(n785), .B(n679), .Z(n673) );
  XNOR U920 ( .A(y[137]), .B(x[137]), .Z(n679) );
  XNOR U921 ( .A(n678), .B(n672), .Z(n785) );
  XNOR U922 ( .A(y[131]), .B(x[131]), .Z(n672) );
  XNOR U923 ( .A(n786), .B(n675), .Z(n678) );
  XNOR U924 ( .A(y[135]), .B(x[135]), .Z(n675) );
  XNOR U925 ( .A(y[136]), .B(x[136]), .Z(n786) );
  XOR U926 ( .A(n682), .B(n681), .Z(n674) );
  XNOR U927 ( .A(n787), .B(n680), .Z(n681) );
  XNOR U928 ( .A(y[132]), .B(x[132]), .Z(n680) );
  XNOR U929 ( .A(y[133]), .B(x[133]), .Z(n787) );
  XOR U930 ( .A(y[134]), .B(x[134]), .Z(n682) );
  XOR U931 ( .A(n700), .B(n683), .Z(n780) );
  XNOR U932 ( .A(y[97]), .B(x[97]), .Z(n683) );
  XOR U933 ( .A(n788), .B(n708), .Z(n700) );
  XNOR U934 ( .A(n692), .B(n691), .Z(n708) );
  XNOR U935 ( .A(n789), .B(n695), .Z(n691) );
  XNOR U936 ( .A(y[152]), .B(x[152]), .Z(n695) );
  XNOR U937 ( .A(n694), .B(n688), .Z(n789) );
  XNOR U938 ( .A(y[146]), .B(x[146]), .Z(n688) );
  XNOR U939 ( .A(n790), .B(n693), .Z(n694) );
  XNOR U940 ( .A(y[150]), .B(x[150]), .Z(n693) );
  XNOR U941 ( .A(y[151]), .B(x[151]), .Z(n790) );
  XOR U942 ( .A(n698), .B(n697), .Z(n692) );
  XNOR U943 ( .A(n791), .B(n696), .Z(n697) );
  XNOR U944 ( .A(y[147]), .B(x[147]), .Z(n696) );
  XNOR U945 ( .A(y[148]), .B(x[148]), .Z(n791) );
  XOR U946 ( .A(y[149]), .B(x[149]), .Z(n698) );
  XNOR U947 ( .A(n707), .B(n699), .Z(n788) );
  XNOR U948 ( .A(y[129]), .B(x[129]), .Z(n699) );
  XNOR U949 ( .A(n792), .B(n712), .Z(n707) );
  XNOR U950 ( .A(n705), .B(n704), .Z(n712) );
  XNOR U951 ( .A(n793), .B(n703), .Z(n704) );
  XNOR U952 ( .A(y[154]), .B(x[154]), .Z(n703) );
  XNOR U953 ( .A(y[155]), .B(x[155]), .Z(n793) );
  XNOR U954 ( .A(y[156]), .B(x[156]), .Z(n705) );
  XNOR U955 ( .A(n711), .B(n706), .Z(n792) );
  XNOR U956 ( .A(y[145]), .B(x[145]), .Z(n706) );
  XNOR U957 ( .A(n794), .B(n715), .Z(n711) );
  XNOR U958 ( .A(y[159]), .B(x[159]), .Z(n715) );
  XNOR U959 ( .A(n714), .B(n710), .Z(n794) );
  XNOR U960 ( .A(y[153]), .B(x[153]), .Z(n710) );
  XNOR U961 ( .A(n795), .B(n713), .Z(n714) );
  XNOR U962 ( .A(y[157]), .B(x[157]), .Z(n713) );
  XNOR U963 ( .A(y[158]), .B(x[158]), .Z(n795) );
endmodule

