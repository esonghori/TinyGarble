
module hamming_N16000_CC16 ( clk, rst, x, y, o );
  input [999:0] x;
  input [999:0] y;
  output [13:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095;
  wire   [13:0] oglobal;

  DFF \oglobal_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .Q(oglobal[13]) );
  DFF \oglobal_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .Q(oglobal[12]) );
  DFF \oglobal_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .Q(oglobal[11]) );
  DFF \oglobal_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .Q(oglobal[10]) );
  DFF \oglobal_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .Q(oglobal[9]) );
  DFF \oglobal_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .Q(oglobal[8]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(oglobal[7]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(oglobal[6]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(oglobal[5]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(oglobal[4]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(oglobal[3]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(oglobal[2]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(oglobal[1]) );
  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(oglobal[0]) );
  NANDN U1003 ( .A(n2018), .B(n2017), .Z(n1) );
  NANDN U1004 ( .A(n2019), .B(n2020), .Z(n2) );
  NAND U1005 ( .A(n1), .B(n2), .Z(n3651) );
  XOR U1006 ( .A(n4269), .B(n4268), .Z(n4640) );
  NAND U1007 ( .A(n4078), .B(n4080), .Z(n3) );
  XOR U1008 ( .A(n4078), .B(n4080), .Z(n4) );
  NAND U1009 ( .A(n4), .B(n4079), .Z(n5) );
  NAND U1010 ( .A(n3), .B(n5), .Z(n5252) );
  NAND U1011 ( .A(n1927), .B(n1928), .Z(n6) );
  NANDN U1012 ( .A(n1925), .B(n1926), .Z(n7) );
  NAND U1013 ( .A(n6), .B(n7), .Z(n3535) );
  NAND U1014 ( .A(n5007), .B(n5008), .Z(n8) );
  XOR U1015 ( .A(n5007), .B(n5008), .Z(n9) );
  NANDN U1016 ( .A(n5006), .B(n9), .Z(n10) );
  NAND U1017 ( .A(n8), .B(n10), .Z(n5547) );
  XOR U1018 ( .A(n5459), .B(n5458), .Z(n5546) );
  XOR U1019 ( .A(n5614), .B(n5613), .Z(n5540) );
  XOR U1020 ( .A(n5469), .B(n5468), .Z(n5470) );
  NAND U1021 ( .A(n4815), .B(n4816), .Z(n11) );
  XOR U1022 ( .A(n4815), .B(n4816), .Z(n12) );
  NANDN U1023 ( .A(n4814), .B(n12), .Z(n13) );
  NAND U1024 ( .A(n11), .B(n13), .Z(n5704) );
  XOR U1025 ( .A(n5857), .B(n5856), .Z(n5858) );
  XOR U1026 ( .A(n5839), .B(n5838), .Z(n5840) );
  XOR U1027 ( .A(n5760), .B(n5759), .Z(n5761) );
  XOR U1028 ( .A(n5796), .B(n5795), .Z(n5797) );
  XNOR U1029 ( .A(n5489), .B(n5488), .Z(n5402) );
  XOR U1030 ( .A(n3754), .B(n3753), .Z(n3755) );
  XOR U1031 ( .A(n4143), .B(n4142), .Z(n4144) );
  XOR U1032 ( .A(n4236), .B(n4235), .Z(n4237) );
  XOR U1033 ( .A(n4010), .B(n4009), .Z(n4012) );
  XOR U1034 ( .A(n4097), .B(n4096), .Z(n3737) );
  XNOR U1035 ( .A(n3732), .B(n3731), .Z(n3783) );
  XOR U1036 ( .A(n4471), .B(n4470), .Z(n4472) );
  NAND U1037 ( .A(n3690), .B(n3691), .Z(n14) );
  XOR U1038 ( .A(n3690), .B(n3691), .Z(n15) );
  NANDN U1039 ( .A(n3689), .B(n15), .Z(n16) );
  NAND U1040 ( .A(n14), .B(n16), .Z(n5003) );
  XOR U1041 ( .A(n5131), .B(n5130), .Z(n5132) );
  NAND U1042 ( .A(n3586), .B(n3588), .Z(n17) );
  XOR U1043 ( .A(n3586), .B(n3588), .Z(n18) );
  NAND U1044 ( .A(n18), .B(n3587), .Z(n19) );
  NAND U1045 ( .A(n17), .B(n19), .Z(n4802) );
  XOR U1046 ( .A(n5253), .B(n5252), .Z(n5254) );
  XOR U1047 ( .A(n4866), .B(n4865), .Z(n4867) );
  NAND U1048 ( .A(n4191), .B(n4192), .Z(n20) );
  XOR U1049 ( .A(n4191), .B(n4192), .Z(n21) );
  NANDN U1050 ( .A(n4190), .B(n21), .Z(n22) );
  NAND U1051 ( .A(n20), .B(n22), .Z(n5168) );
  XOR U1052 ( .A(n4071), .B(n4069), .Z(n23) );
  NANDN U1053 ( .A(n4070), .B(n23), .Z(n24) );
  NAND U1054 ( .A(n4071), .B(n4069), .Z(n25) );
  AND U1055 ( .A(n24), .B(n25), .Z(n4927) );
  NAND U1056 ( .A(n4629), .B(n4631), .Z(n26) );
  XOR U1057 ( .A(n4629), .B(n4631), .Z(n27) );
  NAND U1058 ( .A(n27), .B(n4630), .Z(n28) );
  NAND U1059 ( .A(n26), .B(n28), .Z(n4933) );
  NAND U1060 ( .A(n3703), .B(n3704), .Z(n29) );
  XOR U1061 ( .A(n3703), .B(n3704), .Z(n30) );
  NANDN U1062 ( .A(n3702), .B(n30), .Z(n31) );
  NAND U1063 ( .A(n29), .B(n31), .Z(n4796) );
  XNOR U1064 ( .A(n4856), .B(n4855), .Z(n4789) );
  NAND U1065 ( .A(n3472), .B(n3473), .Z(n32) );
  XOR U1066 ( .A(n3472), .B(n3473), .Z(n33) );
  NANDN U1067 ( .A(n3471), .B(n33), .Z(n34) );
  NAND U1068 ( .A(n32), .B(n34), .Z(n4786) );
  XOR U1069 ( .A(n4608), .B(n4606), .Z(n35) );
  NANDN U1070 ( .A(n4607), .B(n35), .Z(n36) );
  NAND U1071 ( .A(n4608), .B(n4606), .Z(n37) );
  AND U1072 ( .A(n36), .B(n37), .Z(n4775) );
  XOR U1073 ( .A(n4988), .B(n4987), .Z(n4716) );
  XOR U1074 ( .A(n1298), .B(n1297), .Z(n1299) );
  XOR U1075 ( .A(n2880), .B(n2879), .Z(n1847) );
  NANDN U1076 ( .A(n2014), .B(n2013), .Z(n38) );
  NANDN U1077 ( .A(n2015), .B(n2016), .Z(n39) );
  NAND U1078 ( .A(n38), .B(n39), .Z(n3653) );
  NANDN U1079 ( .A(n2135), .B(n2136), .Z(n40) );
  NANDN U1080 ( .A(n2138), .B(n2137), .Z(n41) );
  NAND U1081 ( .A(n40), .B(n41), .Z(n3647) );
  XOR U1082 ( .A(n3639), .B(n3638), .Z(n3640) );
  NAND U1083 ( .A(n4806), .B(n4805), .Z(n42) );
  XOR U1084 ( .A(n4806), .B(n4805), .Z(n43) );
  NANDN U1085 ( .A(n4807), .B(n43), .Z(n44) );
  NAND U1086 ( .A(n42), .B(n44), .Z(n5642) );
  XOR U1087 ( .A(n5612), .B(n5611), .Z(n5613) );
  XOR U1088 ( .A(n5451), .B(n5450), .Z(n5452) );
  XOR U1089 ( .A(n2004), .B(n2003), .Z(n1926) );
  XOR U1090 ( .A(n3408), .B(n3406), .Z(n45) );
  NANDN U1091 ( .A(n3407), .B(n45), .Z(n46) );
  NAND U1092 ( .A(n3408), .B(n3406), .Z(n47) );
  AND U1093 ( .A(n46), .B(n47), .Z(n4924) );
  NAND U1094 ( .A(n3394), .B(n3395), .Z(n48) );
  XOR U1095 ( .A(n3394), .B(n3395), .Z(n49) );
  NANDN U1096 ( .A(n3393), .B(n49), .Z(n50) );
  NAND U1097 ( .A(n48), .B(n50), .Z(n4829) );
  XOR U1098 ( .A(n4940), .B(n4941), .Z(n51) );
  XNOR U1099 ( .A(n4942), .B(n51), .Z(n4761) );
  NAND U1100 ( .A(n3779), .B(n3780), .Z(n52) );
  XOR U1101 ( .A(n3779), .B(n3780), .Z(n53) );
  NANDN U1102 ( .A(n3778), .B(n53), .Z(n54) );
  NAND U1103 ( .A(n52), .B(n54), .Z(n4970) );
  XNOR U1104 ( .A(n5477), .B(n5476), .Z(n5511) );
  XOR U1105 ( .A(n5678), .B(n5677), .Z(n5681) );
  XOR U1106 ( .A(n5447), .B(n5446), .Z(n5414) );
  NAND U1107 ( .A(n4832), .B(n4833), .Z(n55) );
  XOR U1108 ( .A(n4832), .B(n4833), .Z(n56) );
  NANDN U1109 ( .A(n4834), .B(n56), .Z(n57) );
  NAND U1110 ( .A(n55), .B(n57), .Z(n5432) );
  XOR U1111 ( .A(n5754), .B(n5753), .Z(n5755) );
  NAND U1112 ( .A(n5710), .B(n5712), .Z(n58) );
  XOR U1113 ( .A(n5710), .B(n5712), .Z(n59) );
  NAND U1114 ( .A(n59), .B(n5711), .Z(n60) );
  NAND U1115 ( .A(n58), .B(n60), .Z(n5807) );
  XOR U1116 ( .A(n5853), .B(n5852), .Z(n5777) );
  XOR U1117 ( .A(n5859), .B(n5858), .Z(n5783) );
  XOR U1118 ( .A(n5790), .B(n5789), .Z(n5792) );
  XOR U1119 ( .A(n5798), .B(n5797), .Z(n5874) );
  XNOR U1120 ( .A(n5974), .B(n5973), .Z(n5979) );
  NAND U1121 ( .A(n5719), .B(n5721), .Z(n61) );
  XOR U1122 ( .A(n5719), .B(n5721), .Z(n62) );
  NAND U1123 ( .A(n62), .B(n5720), .Z(n63) );
  NAND U1124 ( .A(n61), .B(n63), .Z(n5911) );
  XOR U1125 ( .A(n3205), .B(n3204), .Z(n3206) );
  XOR U1126 ( .A(n1942), .B(n1941), .Z(n1943) );
  XOR U1127 ( .A(n2028), .B(n2027), .Z(n2029) );
  XOR U1128 ( .A(n3187), .B(n3186), .Z(n3188) );
  XOR U1129 ( .A(n2497), .B(n2496), .Z(n2498) );
  XOR U1130 ( .A(n2232), .B(n2231), .Z(n2233) );
  XOR U1131 ( .A(n3235), .B(n3234), .Z(n3236) );
  XOR U1132 ( .A(n3053), .B(n3052), .Z(n3054) );
  XOR U1133 ( .A(n2569), .B(n2568), .Z(n2570) );
  XOR U1134 ( .A(n3326), .B(n3325), .Z(n3328) );
  XOR U1135 ( .A(n4162), .B(n4161), .Z(n4163) );
  XOR U1136 ( .A(n4119), .B(n4118), .Z(n4121) );
  XOR U1137 ( .A(n4125), .B(n4124), .Z(n4127) );
  XOR U1138 ( .A(n4113), .B(n4112), .Z(n4115) );
  XOR U1139 ( .A(n4393), .B(n4392), .Z(n4395) );
  XOR U1140 ( .A(n4052), .B(n4051), .Z(n4053) );
  XOR U1141 ( .A(n4212), .B(n4211), .Z(n4214) );
  XOR U1142 ( .A(n3819), .B(n3818), .Z(n3821) );
  XOR U1143 ( .A(n3813), .B(n3812), .Z(n3815) );
  XOR U1144 ( .A(n3825), .B(n3824), .Z(n3827) );
  XOR U1145 ( .A(n3609), .B(n3608), .Z(n3611) );
  XOR U1146 ( .A(n3878), .B(n3877), .Z(n3879) );
  XOR U1147 ( .A(n4417), .B(n4416), .Z(n4418) );
  XOR U1148 ( .A(n3597), .B(n3596), .Z(n3598) );
  XOR U1149 ( .A(n3603), .B(n3602), .Z(n3605) );
  XOR U1150 ( .A(n3591), .B(n3590), .Z(n3593) );
  XOR U1151 ( .A(n4107), .B(n4106), .Z(n4109) );
  XOR U1152 ( .A(n4435), .B(n4434), .Z(n4436) );
  XOR U1153 ( .A(n2317), .B(n2316), .Z(n2318) );
  XOR U1154 ( .A(n2577), .B(n2576), .Z(n1929) );
  XOR U1155 ( .A(n3583), .B(n3584), .Z(n64) );
  XNOR U1156 ( .A(n3585), .B(n64), .Z(n4634) );
  XOR U1157 ( .A(n4465), .B(n4464), .Z(n4466) );
  XOR U1158 ( .A(n3724), .B(n3723), .Z(n3725) );
  XOR U1159 ( .A(n4610), .B(n4612), .Z(n65) );
  XNOR U1160 ( .A(n4613), .B(n65), .Z(n3650) );
  NANDN U1161 ( .A(n1967), .B(n1966), .Z(n66) );
  NANDN U1162 ( .A(n1968), .B(n1969), .Z(n67) );
  NAND U1163 ( .A(n66), .B(n67), .Z(n3541) );
  XOR U1164 ( .A(n4238), .B(n4237), .Z(n4639) );
  XOR U1165 ( .A(n5279), .B(n5278), .Z(n5007) );
  XOR U1166 ( .A(n5137), .B(n5136), .Z(n5138) );
  XOR U1167 ( .A(n5125), .B(n5124), .Z(n5126) );
  XOR U1168 ( .A(n4879), .B(n4878), .Z(n4895) );
  NAND U1169 ( .A(n3308), .B(n3309), .Z(n68) );
  XOR U1170 ( .A(n3308), .B(n3309), .Z(n69) );
  NANDN U1171 ( .A(n3307), .B(n69), .Z(n70) );
  NAND U1172 ( .A(n68), .B(n70), .Z(n4805) );
  XOR U1173 ( .A(n5259), .B(n5258), .Z(n5260) );
  XOR U1174 ( .A(n5247), .B(n5246), .Z(n5248) );
  XOR U1175 ( .A(n4848), .B(n4847), .Z(n4849) );
  XOR U1176 ( .A(n4842), .B(n4841), .Z(n4843) );
  NAND U1177 ( .A(n3456), .B(n3455), .Z(n71) );
  XOR U1178 ( .A(n3456), .B(n3455), .Z(n72) );
  NANDN U1179 ( .A(n3457), .B(n72), .Z(n73) );
  NAND U1180 ( .A(n71), .B(n73), .Z(n4853) );
  XOR U1181 ( .A(n4860), .B(n4859), .Z(n4861) );
  XOR U1182 ( .A(n5094), .B(n5093), .Z(n5095) );
  XNOR U1183 ( .A(n4769), .B(n4770), .Z(n74) );
  XNOR U1184 ( .A(n4768), .B(n74), .Z(n4741) );
  NAND U1185 ( .A(n4642), .B(n4643), .Z(n75) );
  XOR U1186 ( .A(n4642), .B(n4643), .Z(n76) );
  NANDN U1187 ( .A(n4641), .B(n76), .Z(n77) );
  NAND U1188 ( .A(n75), .B(n77), .Z(n4985) );
  XNOR U1189 ( .A(n5042), .B(n5041), .Z(n4700) );
  XNOR U1190 ( .A(n5255), .B(n5254), .Z(n4928) );
  NAND U1191 ( .A(n4627), .B(n4628), .Z(n78) );
  XOR U1192 ( .A(n4627), .B(n4628), .Z(n79) );
  NANDN U1193 ( .A(n4626), .B(n79), .Z(n80) );
  NAND U1194 ( .A(n78), .B(n80), .Z(n4934) );
  NAND U1195 ( .A(n3700), .B(n3701), .Z(n81) );
  XOR U1196 ( .A(n3700), .B(n3701), .Z(n82) );
  NANDN U1197 ( .A(n3699), .B(n82), .Z(n83) );
  NAND U1198 ( .A(n81), .B(n83), .Z(n4797) );
  XOR U1199 ( .A(n3460), .B(n3458), .Z(n84) );
  NANDN U1200 ( .A(n3459), .B(n84), .Z(n85) );
  NAND U1201 ( .A(n3460), .B(n3458), .Z(n86) );
  AND U1202 ( .A(n85), .B(n86), .Z(n4790) );
  XOR U1203 ( .A(n3470), .B(n3468), .Z(n87) );
  NANDN U1204 ( .A(n3469), .B(n87), .Z(n88) );
  NAND U1205 ( .A(n3470), .B(n3468), .Z(n89) );
  AND U1206 ( .A(n88), .B(n89), .Z(n4787) );
  XOR U1207 ( .A(n5143), .B(n5142), .Z(n5145) );
  XOR U1208 ( .A(n5229), .B(n5228), .Z(n5231) );
  XOR U1209 ( .A(n5267), .B(n5266), .Z(n4964) );
  XNOR U1210 ( .A(n4777), .B(n4776), .Z(n4939) );
  XOR U1211 ( .A(n2935), .B(n2934), .Z(n2345) );
  XNOR U1212 ( .A(n3097), .B(n3096), .Z(n2589) );
  XOR U1213 ( .A(n4477), .B(n4476), .Z(n4478) );
  XOR U1214 ( .A(n3645), .B(n3644), .Z(n3646) );
  XOR U1215 ( .A(n4249), .B(n4248), .Z(n4250) );
  NAND U1216 ( .A(n1063), .B(n1064), .Z(n90) );
  NANDN U1217 ( .A(n1061), .B(n1062), .Z(n91) );
  NAND U1218 ( .A(n90), .B(n91), .Z(n3553) );
  XOR U1219 ( .A(n3801), .B(n3800), .Z(n3802) );
  XOR U1220 ( .A(n718), .B(n717), .Z(n247) );
  XOR U1221 ( .A(n5082), .B(n5081), .Z(n5083) );
  NANDN U1222 ( .A(n2342), .B(n2341), .Z(n92) );
  NANDN U1223 ( .A(n2343), .B(n2344), .Z(n93) );
  NAND U1224 ( .A(n92), .B(n93), .Z(n4281) );
  XNOR U1225 ( .A(n5133), .B(n5132), .Z(n5188) );
  XOR U1226 ( .A(n4961), .B(n4960), .Z(n4824) );
  NAND U1227 ( .A(n5004), .B(n5005), .Z(n94) );
  XOR U1228 ( .A(n5004), .B(n5005), .Z(n95) );
  NANDN U1229 ( .A(n5003), .B(n95), .Z(n96) );
  NAND U1230 ( .A(n94), .B(n96), .Z(n5548) );
  XOR U1231 ( .A(n5457), .B(n5456), .Z(n5458) );
  XOR U1232 ( .A(n4802), .B(n4803), .Z(n97) );
  NANDN U1233 ( .A(n4804), .B(n97), .Z(n98) );
  NAND U1234 ( .A(n4802), .B(n4803), .Z(n99) );
  AND U1235 ( .A(n98), .B(n99), .Z(n5641) );
  XOR U1236 ( .A(n4773), .B(n4771), .Z(n100) );
  NANDN U1237 ( .A(n4772), .B(n100), .Z(n101) );
  NAND U1238 ( .A(n4773), .B(n4771), .Z(n102) );
  AND U1239 ( .A(n101), .B(n102), .Z(n5653) );
  XOR U1240 ( .A(n5670), .B(n5669), .Z(n5671) );
  NAND U1241 ( .A(n4930), .B(n4932), .Z(n103) );
  XOR U1242 ( .A(n4930), .B(n4932), .Z(n104) );
  NAND U1243 ( .A(n104), .B(n4931), .Z(n105) );
  NAND U1244 ( .A(n103), .B(n105), .Z(n5623) );
  XOR U1245 ( .A(n5618), .B(n5617), .Z(n5620) );
  XOR U1246 ( .A(n5707), .B(n5706), .Z(n5578) );
  XOR U1247 ( .A(n3809), .B(n3808), .Z(n4664) );
  XOR U1248 ( .A(n3536), .B(n3535), .Z(n3537) );
  XNOR U1249 ( .A(n3532), .B(n3531), .Z(n3500) );
  XOR U1250 ( .A(n3566), .B(n3565), .Z(n3567) );
  XOR U1251 ( .A(n3633), .B(n3632), .Z(n3634) );
  NAND U1252 ( .A(n4028), .B(n4029), .Z(n106) );
  XOR U1253 ( .A(n4028), .B(n4029), .Z(n107) );
  NANDN U1254 ( .A(n4027), .B(n107), .Z(n108) );
  NAND U1255 ( .A(n106), .B(n108), .Z(n5332) );
  XOR U1256 ( .A(n5523), .B(n5522), .Z(n5524) );
  XNOR U1257 ( .A(n5556), .B(n5555), .Z(n5493) );
  NAND U1258 ( .A(n4971), .B(n4972), .Z(n109) );
  XOR U1259 ( .A(n4971), .B(n4972), .Z(n110) );
  NANDN U1260 ( .A(n4970), .B(n110), .Z(n111) );
  NAND U1261 ( .A(n109), .B(n111), .Z(n5682) );
  XOR U1262 ( .A(n4924), .B(n4925), .Z(n112) );
  NANDN U1263 ( .A(n4926), .B(n112), .Z(n113) );
  NAND U1264 ( .A(n4924), .B(n4925), .Z(n114) );
  AND U1265 ( .A(n113), .B(n114), .Z(n5415) );
  NAND U1266 ( .A(n4829), .B(n4830), .Z(n115) );
  XOR U1267 ( .A(n4829), .B(n4830), .Z(n116) );
  NANDN U1268 ( .A(n4831), .B(n116), .Z(n117) );
  NAND U1269 ( .A(n115), .B(n117), .Z(n5433) );
  NAND U1270 ( .A(n5659), .B(n5661), .Z(n118) );
  XOR U1271 ( .A(n5659), .B(n5661), .Z(n119) );
  NAND U1272 ( .A(n119), .B(n5660), .Z(n120) );
  NAND U1273 ( .A(n118), .B(n120), .Z(n5825) );
  XOR U1274 ( .A(n5841), .B(n5840), .Z(n5762) );
  XOR U1275 ( .A(n5834), .B(n5833), .Z(n5765) );
  XOR U1276 ( .A(n5810), .B(n5809), .Z(n5801) );
  NAND U1277 ( .A(n5584), .B(n5586), .Z(n121) );
  XOR U1278 ( .A(n5584), .B(n5586), .Z(n122) );
  NAND U1279 ( .A(n122), .B(n5585), .Z(n123) );
  NAND U1280 ( .A(n121), .B(n123), .Z(n5795) );
  NANDN U1281 ( .A(n5534), .B(n5537), .Z(n124) );
  OR U1282 ( .A(n5537), .B(n5536), .Z(n125) );
  NAND U1283 ( .A(n5535), .B(n125), .Z(n126) );
  NAND U1284 ( .A(n124), .B(n126), .Z(n5778) );
  XOR U1285 ( .A(n5784), .B(n5783), .Z(n5785) );
  XNOR U1286 ( .A(n5423), .B(n5422), .Z(n5388) );
  XNOR U1287 ( .A(n5441), .B(n5440), .Z(n5487) );
  XNOR U1288 ( .A(n5750), .B(n5749), .Z(n5865) );
  XOR U1289 ( .A(n5962), .B(n5961), .Z(n5967) );
  XOR U1290 ( .A(n4022), .B(n4021), .Z(n4023) );
  XOR U1291 ( .A(n5877), .B(n5876), .Z(n5899) );
  XNOR U1292 ( .A(n6041), .B(n6040), .Z(n6023) );
  XOR U1293 ( .A(n5400), .B(n5399), .Z(n5401) );
  XOR U1294 ( .A(n6067), .B(n6066), .Z(n6068) );
  NAND U1295 ( .A(n5350), .B(n5351), .Z(n127) );
  XOR U1296 ( .A(n5350), .B(n5351), .Z(n128) );
  NANDN U1297 ( .A(n5349), .B(n128), .Z(n129) );
  NAND U1298 ( .A(n127), .B(n129), .Z(n5720) );
  NAND U1299 ( .A(n6077), .B(n6079), .Z(n130) );
  XOR U1300 ( .A(n6077), .B(n6079), .Z(n131) );
  NAND U1301 ( .A(n131), .B(n6078), .Z(n132) );
  NAND U1302 ( .A(n130), .B(n132), .Z(n6086) );
  XOR U1303 ( .A(n1500), .B(n1499), .Z(n1501) );
  XOR U1304 ( .A(n3217), .B(n3216), .Z(n3218) );
  XOR U1305 ( .A(n2443), .B(n2442), .Z(n2444) );
  XOR U1306 ( .A(n2425), .B(n2424), .Z(n2426) );
  XOR U1307 ( .A(n2951), .B(n2950), .Z(n2952) );
  XOR U1308 ( .A(n1954), .B(n1953), .Z(n1955) );
  XOR U1309 ( .A(n2281), .B(n2280), .Z(n2282) );
  XOR U1310 ( .A(n2293), .B(n2292), .Z(n2294) );
  XOR U1311 ( .A(n1195), .B(n1194), .Z(n1196) );
  XOR U1312 ( .A(n2220), .B(n2219), .Z(n2221) );
  XOR U1313 ( .A(n2262), .B(n2261), .Z(n2263) );
  XOR U1314 ( .A(n910), .B(n909), .Z(n911) );
  XOR U1315 ( .A(n2981), .B(n2980), .Z(n2982) );
  XOR U1316 ( .A(n2975), .B(n2974), .Z(n2976) );
  XOR U1317 ( .A(n2503), .B(n2502), .Z(n2504) );
  XOR U1318 ( .A(n952), .B(n951), .Z(n953) );
  XOR U1319 ( .A(n1626), .B(n1625), .Z(n1627) );
  XOR U1320 ( .A(n851), .B(n850), .Z(n852) );
  XOR U1321 ( .A(n845), .B(n844), .Z(n846) );
  XOR U1322 ( .A(n2040), .B(n2039), .Z(n2041) );
  XOR U1323 ( .A(n2684), .B(n2683), .Z(n2685) );
  XOR U1324 ( .A(n1596), .B(n1595), .Z(n1597) );
  XOR U1325 ( .A(n3199), .B(n3198), .Z(n3200) );
  XOR U1326 ( .A(n2226), .B(n2225), .Z(n2227) );
  XOR U1327 ( .A(n2305), .B(n2304), .Z(n2306) );
  XOR U1328 ( .A(n2244), .B(n2243), .Z(n2245) );
  XOR U1329 ( .A(n2485), .B(n2484), .Z(n2486) );
  XOR U1330 ( .A(n3145), .B(n3144), .Z(n3146) );
  XOR U1331 ( .A(n2945), .B(n2944), .Z(n2946) );
  XOR U1332 ( .A(n2575), .B(n2574), .Z(n2576) );
  XOR U1333 ( .A(n1020), .B(n1019), .Z(n1021) );
  XOR U1334 ( .A(n1590), .B(n1589), .Z(n1591) );
  XNOR U1335 ( .A(n4164), .B(n4163), .Z(n3331) );
  XOR U1336 ( .A(n4447), .B(n4446), .Z(n4448) );
  XOR U1337 ( .A(n4453), .B(n4452), .Z(n4454) );
  XOR U1338 ( .A(n4261), .B(n4260), .Z(n4263) );
  XOR U1339 ( .A(n4531), .B(n4530), .Z(n4533) );
  XOR U1340 ( .A(n3980), .B(n3979), .Z(n3982) );
  XOR U1341 ( .A(n3986), .B(n3985), .Z(n3988) );
  XOR U1342 ( .A(n4156), .B(n4155), .Z(n4158) );
  XOR U1343 ( .A(n4381), .B(n4380), .Z(n4383) );
  XOR U1344 ( .A(n4131), .B(n4130), .Z(n4133) );
  XOR U1345 ( .A(n4137), .B(n4136), .Z(n4139) );
  XOR U1346 ( .A(n4315), .B(n4314), .Z(n4317) );
  XOR U1347 ( .A(n4573), .B(n4572), .Z(n4575) );
  XOR U1348 ( .A(n4297), .B(n4296), .Z(n4299) );
  XOR U1349 ( .A(n3615), .B(n3614), .Z(n3617) );
  XOR U1350 ( .A(n4363), .B(n4362), .Z(n4364) );
  XOR U1351 ( .A(n3962), .B(n3961), .Z(n3964) );
  XOR U1352 ( .A(n3956), .B(n3955), .Z(n3958) );
  XOR U1353 ( .A(n3950), .B(n3949), .Z(n3951) );
  XOR U1354 ( .A(n4095), .B(n4094), .Z(n4096) );
  XOR U1355 ( .A(n3932), .B(n3931), .Z(n3934) );
  XOR U1356 ( .A(n4016), .B(n4015), .Z(n4018) );
  XOR U1357 ( .A(n4004), .B(n4003), .Z(n4006) );
  XOR U1358 ( .A(n4459), .B(n4458), .Z(n4460) );
  NAND U1359 ( .A(n606), .B(n605), .Z(n133) );
  NANDN U1360 ( .A(n603), .B(n604), .Z(n134) );
  AND U1361 ( .A(n133), .B(n134), .Z(n4587) );
  XOR U1362 ( .A(n3083), .B(n3082), .Z(n3084) );
  XOR U1363 ( .A(n2678), .B(n2677), .Z(n2679) );
  XOR U1364 ( .A(n2196), .B(n2195), .Z(n2197) );
  XOR U1365 ( .A(n2268), .B(n2267), .Z(n2269) );
  XOR U1366 ( .A(n3055), .B(n3054), .Z(n2720) );
  XOR U1367 ( .A(n2545), .B(n2544), .Z(n2546) );
  XOR U1368 ( .A(n2571), .B(n2570), .Z(n1930) );
  XOR U1369 ( .A(n2592), .B(n2591), .Z(n2593) );
  XOR U1370 ( .A(n4208), .B(n4207), .Z(n3469) );
  XOR U1371 ( .A(n3712), .B(n3711), .Z(n3713) );
  XOR U1372 ( .A(n4501), .B(n4500), .Z(n4502) );
  XOR U1373 ( .A(n3739), .B(n3741), .Z(n135) );
  XNOR U1374 ( .A(n3742), .B(n135), .Z(n3529) );
  XNOR U1375 ( .A(n5285), .B(n5284), .Z(n4894) );
  XNOR U1376 ( .A(n5072), .B(n5071), .Z(n4889) );
  XOR U1377 ( .A(n4907), .B(n4906), .Z(n4908) );
  NAND U1378 ( .A(n3349), .B(n3350), .Z(n136) );
  XOR U1379 ( .A(n3349), .B(n3350), .Z(n137) );
  NANDN U1380 ( .A(n3348), .B(n137), .Z(n138) );
  NAND U1381 ( .A(n136), .B(n138), .Z(n5300) );
  XOR U1382 ( .A(n5289), .B(n5288), .Z(n5290) );
  XOR U1383 ( .A(n5076), .B(n5075), .Z(n5077) );
  XOR U1384 ( .A(n4809), .B(n4808), .Z(n4810) );
  XOR U1385 ( .A(n4872), .B(n4871), .Z(n4873) );
  XOR U1386 ( .A(n5048), .B(n5047), .Z(n4868) );
  XOR U1387 ( .A(n3294), .B(n3293), .Z(n139) );
  NANDN U1388 ( .A(n3292), .B(n139), .Z(n140) );
  NAND U1389 ( .A(n3294), .B(n3293), .Z(n141) );
  AND U1390 ( .A(n140), .B(n141), .Z(n5276) );
  XOR U1391 ( .A(n5157), .B(n5156), .Z(n5158) );
  NAND U1392 ( .A(n4188), .B(n4189), .Z(n142) );
  XOR U1393 ( .A(n4188), .B(n4189), .Z(n143) );
  NANDN U1394 ( .A(n4187), .B(n143), .Z(n144) );
  NAND U1395 ( .A(n142), .B(n144), .Z(n5169) );
  XOR U1396 ( .A(n5163), .B(n5162), .Z(n5164) );
  XOR U1397 ( .A(n5100), .B(n5099), .Z(n5101) );
  XNOR U1398 ( .A(n5096), .B(n5095), .Z(n4743) );
  NAND U1399 ( .A(n4639), .B(n4640), .Z(n145) );
  XOR U1400 ( .A(n4639), .B(n4640), .Z(n146) );
  NANDN U1401 ( .A(n4638), .B(n146), .Z(n147) );
  NAND U1402 ( .A(n145), .B(n147), .Z(n4986) );
  XOR U1403 ( .A(n4980), .B(n4979), .Z(n4982) );
  XOR U1404 ( .A(n5175), .B(n5174), .Z(n5176) );
  XOR U1405 ( .A(n5052), .B(n5051), .Z(n5053) );
  XOR U1406 ( .A(n4592), .B(n4590), .Z(n148) );
  NANDN U1407 ( .A(n4591), .B(n148), .Z(n149) );
  NAND U1408 ( .A(n4592), .B(n4590), .Z(n150) );
  AND U1409 ( .A(n149), .B(n150), .Z(n4815) );
  XOR U1410 ( .A(n5307), .B(n5306), .Z(n5309) );
  XNOR U1411 ( .A(n5273), .B(n5272), .Z(n4782) );
  NAND U1412 ( .A(n4152), .B(n4154), .Z(n151) );
  XOR U1413 ( .A(n4152), .B(n4154), .Z(n152) );
  NAND U1414 ( .A(n152), .B(n4153), .Z(n153) );
  NAND U1415 ( .A(n151), .B(n153), .Z(n5217) );
  XOR U1416 ( .A(n4936), .B(n4935), .Z(n4717) );
  XOR U1417 ( .A(n5315), .B(n5314), .Z(n4965) );
  XOR U1418 ( .A(n2256), .B(n2255), .Z(n2257) );
  XOR U1419 ( .A(n2146), .B(n2145), .Z(n2147) );
  XOR U1420 ( .A(n3011), .B(n3010), .Z(n3012) );
  XOR U1421 ( .A(n1108), .B(n1107), .Z(n1109) );
  XOR U1422 ( .A(n1104), .B(n1103), .Z(n1848) );
  XNOR U1423 ( .A(n4467), .B(n4466), .Z(n3784) );
  XOR U1424 ( .A(n3651), .B(n3650), .Z(n3652) );
  XNOR U1425 ( .A(n4000), .B(n3999), .Z(n3873) );
  XOR U1426 ( .A(n3675), .B(n3674), .Z(n3677) );
  XOR U1427 ( .A(n4089), .B(n4088), .Z(n4091) );
  XOR U1428 ( .A(n4883), .B(n4882), .Z(n4884) );
  XNOR U1429 ( .A(n5139), .B(n5138), .Z(n4946) );
  XOR U1430 ( .A(n5320), .B(n5319), .Z(n5322) );
  NANDN U1431 ( .A(n2589), .B(n2590), .Z(n154) );
  NANDN U1432 ( .A(n2588), .B(n2587), .Z(n155) );
  AND U1433 ( .A(n154), .B(n155), .Z(n3708) );
  XOR U1434 ( .A(n4617), .B(n4618), .Z(n156) );
  NANDN U1435 ( .A(n4619), .B(n156), .Z(n157) );
  NAND U1436 ( .A(n4617), .B(n4618), .Z(n158) );
  AND U1437 ( .A(n157), .B(n158), .Z(n4940) );
  XOR U1438 ( .A(n5193), .B(n5192), .Z(n5195) );
  XNOR U1439 ( .A(n4736), .B(n4735), .Z(n4738) );
  XOR U1440 ( .A(n5539), .B(n5538), .Z(n5541) );
  XOR U1441 ( .A(n5642), .B(n5641), .Z(n5644) );
  XOR U1442 ( .A(n5572), .B(n5571), .Z(n5573) );
  XOR U1443 ( .A(n5566), .B(n5565), .Z(n5567) );
  XOR U1444 ( .A(n5600), .B(n5599), .Z(n5601) );
  XOR U1445 ( .A(n5630), .B(n5629), .Z(n5631) );
  NAND U1446 ( .A(n4928), .B(n4929), .Z(n159) );
  XOR U1447 ( .A(n4928), .B(n4929), .Z(n160) );
  NANDN U1448 ( .A(n4927), .B(n160), .Z(n161) );
  NAND U1449 ( .A(n159), .B(n161), .Z(n5624) );
  XOR U1450 ( .A(n5699), .B(n5698), .Z(n5700) );
  XOR U1451 ( .A(n5714), .B(n5713), .Z(n5715) );
  XOR U1452 ( .A(n5596), .B(n5595), .Z(n5579) );
  XOR U1453 ( .A(n5588), .B(n5587), .Z(n5589) );
  XOR U1454 ( .A(n5550), .B(n5549), .Z(n5675) );
  XOR U1455 ( .A(n2909), .B(n2908), .Z(n2910) );
  XNOR U1456 ( .A(n2048), .B(n2047), .Z(n2015) );
  XOR U1457 ( .A(n4479), .B(n4478), .Z(n3769) );
  XNOR U1458 ( .A(n3647), .B(n3646), .Z(n3404) );
  XOR U1459 ( .A(n5235), .B(n5234), .Z(n5236) );
  XOR U1460 ( .A(n4281), .B(n4280), .Z(n3418) );
  NAND U1461 ( .A(n4663), .B(n4664), .Z(n162) );
  XOR U1462 ( .A(n4663), .B(n4664), .Z(n163) );
  NANDN U1463 ( .A(n4662), .B(n163), .Z(n164) );
  NAND U1464 ( .A(n162), .B(n164), .Z(n4759) );
  NAND U1465 ( .A(n3776), .B(n3777), .Z(n165) );
  XOR U1466 ( .A(n3776), .B(n3777), .Z(n166) );
  NANDN U1467 ( .A(n3775), .B(n166), .Z(n167) );
  NAND U1468 ( .A(n165), .B(n167), .Z(n4971) );
  XOR U1469 ( .A(n5121), .B(n5120), .Z(n5325) );
  XOR U1470 ( .A(n5493), .B(n5492), .Z(n5495) );
  XOR U1471 ( .A(n5453), .B(n5452), .Z(n5684) );
  XNOR U1472 ( .A(n5417), .B(n5416), .Z(n5409) );
  NAND U1473 ( .A(n5545), .B(n5546), .Z(n168) );
  XOR U1474 ( .A(n5545), .B(n5546), .Z(n169) );
  NANDN U1475 ( .A(n5544), .B(n169), .Z(n170) );
  NAND U1476 ( .A(n168), .B(n170), .Z(n5851) );
  XOR U1477 ( .A(n5845), .B(n5844), .Z(n5846) );
  XOR U1478 ( .A(n5837), .B(oglobal[4]), .Z(n5831) );
  XOR U1479 ( .A(n5820), .B(n5819), .Z(n5821) );
  XOR U1480 ( .A(n5826), .B(n5825), .Z(n5827) );
  XOR U1481 ( .A(n5808), .B(n5807), .Z(n5809) );
  NAND U1482 ( .A(n5696), .B(n5697), .Z(n171) );
  XOR U1483 ( .A(n5696), .B(n5697), .Z(n172) );
  NANDN U1484 ( .A(n5695), .B(n172), .Z(n173) );
  NAND U1485 ( .A(n171), .B(n173), .Z(n5802) );
  XOR U1486 ( .A(n3538), .B(n3537), .Z(n3501) );
  XNOR U1487 ( .A(n3568), .B(n3567), .Z(n3395) );
  XNOR U1488 ( .A(n4955), .B(n4954), .Z(n4689) );
  XOR U1489 ( .A(n5388), .B(n5387), .Z(n5389) );
  XOR U1490 ( .A(n5875), .B(n5874), .Z(n5876) );
  XNOR U1491 ( .A(n5334), .B(n5333), .Z(n5363) );
  XNOR U1492 ( .A(n5865), .B(n5864), .Z(n5901) );
  XOR U1493 ( .A(n5992), .B(n5991), .Z(n5937) );
  XOR U1494 ( .A(n5986), .B(n5985), .Z(n5931) );
  XNOR U1495 ( .A(n6030), .B(n6029), .Z(n6039) );
  XOR U1496 ( .A(n6022), .B(n6021), .Z(n6024) );
  XOR U1497 ( .A(n5402), .B(n5401), .Z(n5721) );
  NAND U1498 ( .A(n5354), .B(n5355), .Z(n174) );
  XOR U1499 ( .A(n5354), .B(n5355), .Z(n175) );
  NANDN U1500 ( .A(n5353), .B(n175), .Z(n176) );
  NAND U1501 ( .A(n174), .B(n176), .Z(n5405) );
  NAND U1502 ( .A(n6087), .B(n6088), .Z(n177) );
  XOR U1503 ( .A(n6087), .B(n6088), .Z(n178) );
  NAND U1504 ( .A(n178), .B(n6086), .Z(n179) );
  NAND U1505 ( .A(n177), .B(n179), .Z(n6090) );
  XOR U1506 ( .A(n3211), .B(n3210), .Z(n3212) );
  XOR U1507 ( .A(n3133), .B(n3132), .Z(n3134) );
  XOR U1508 ( .A(n2455), .B(n2454), .Z(n2456) );
  XOR U1509 ( .A(n2323), .B(n2322), .Z(n2324) );
  XOR U1510 ( .A(n324), .B(n323), .Z(n325) );
  XOR U1511 ( .A(n1360), .B(n1359), .Z(n1361) );
  XOR U1512 ( .A(n1354), .B(n1353), .Z(n1355) );
  XOR U1513 ( .A(n1470), .B(n1469), .Z(n1471) );
  XOR U1514 ( .A(n1482), .B(n1481), .Z(n1483) );
  XOR U1515 ( .A(n3041), .B(n3040), .Z(n3042) );
  XOR U1516 ( .A(n3035), .B(n3034), .Z(n3036) );
  XOR U1517 ( .A(n3047), .B(n3046), .Z(n3048) );
  XOR U1518 ( .A(n1753), .B(n1752), .Z(n1754) );
  XOR U1519 ( .A(n1759), .B(n1758), .Z(n1760) );
  XOR U1520 ( .A(n1914), .B(n1913), .Z(n1915) );
  XOR U1521 ( .A(n1828), .B(n1827), .Z(n1829) );
  XOR U1522 ( .A(n771), .B(n770), .Z(n772) );
  XOR U1523 ( .A(n3005), .B(n3004), .Z(n3006) );
  XOR U1524 ( .A(n2274), .B(n2273), .Z(n2275) );
  XOR U1525 ( .A(n904), .B(n903), .Z(n905) );
  XOR U1526 ( .A(n898), .B(n897), .Z(n899) );
  XOR U1527 ( .A(n2853), .B(n2852), .Z(n2854) );
  XOR U1528 ( .A(n2859), .B(n2858), .Z(n2860) );
  XOR U1529 ( .A(n2987), .B(n2986), .Z(n2988) );
  XOR U1530 ( .A(n2184), .B(n2183), .Z(n2185) );
  XOR U1531 ( .A(n1710), .B(n1709), .Z(n1711) );
  XOR U1532 ( .A(n1722), .B(n1721), .Z(n1723) );
  XOR U1533 ( .A(n2388), .B(n2387), .Z(n2389) );
  XOR U1534 ( .A(n2915), .B(n2914), .Z(n2916) );
  XOR U1535 ( .A(n857), .B(n856), .Z(n858) );
  XOR U1536 ( .A(n1638), .B(n1637), .Z(n1639) );
  XOR U1537 ( .A(n1644), .B(n1643), .Z(n1645) );
  XOR U1538 ( .A(n1662), .B(n1661), .Z(n1663) );
  XOR U1539 ( .A(n3175), .B(n3174), .Z(n3176) );
  XOR U1540 ( .A(n3181), .B(n3180), .Z(n3182) );
  XOR U1541 ( .A(n2757), .B(n2756), .Z(n2758) );
  XOR U1542 ( .A(n2751), .B(n2750), .Z(n2752) );
  XOR U1543 ( .A(n2696), .B(n2695), .Z(n2697) );
  XOR U1544 ( .A(n2805), .B(n2804), .Z(n2806) );
  XOR U1545 ( .A(n2811), .B(n2810), .Z(n2812) );
  XOR U1546 ( .A(n2158), .B(n2157), .Z(n2159) );
  XOR U1547 ( .A(n2672), .B(n2671), .Z(n2673) );
  XOR U1548 ( .A(n2733), .B(n2732), .Z(n2734) );
  XOR U1549 ( .A(n2745), .B(n2744), .Z(n2746) );
  XOR U1550 ( .A(n1316), .B(n1315), .Z(n1317) );
  XOR U1551 ( .A(n1310), .B(n1309), .Z(n1311) );
  XOR U1552 ( .A(n1304), .B(n1303), .Z(n1305) );
  XOR U1553 ( .A(n1995), .B(n1994), .Z(n1996) );
  XOR U1554 ( .A(n1983), .B(n1982), .Z(n1984) );
  XOR U1555 ( .A(n2666), .B(n2665), .Z(n2667) );
  XOR U1556 ( .A(n1280), .B(n1279), .Z(n1281) );
  XOR U1557 ( .A(n734), .B(n733), .Z(n735) );
  XOR U1558 ( .A(n1268), .B(n1267), .Z(n1269) );
  XOR U1559 ( .A(n2521), .B(n2520), .Z(n2522) );
  XOR U1560 ( .A(n2533), .B(n2532), .Z(n2534) );
  XOR U1561 ( .A(n1686), .B(n1685), .Z(n1687) );
  XOR U1562 ( .A(n1232), .B(n1231), .Z(n1233) );
  XOR U1563 ( .A(n1244), .B(n1243), .Z(n1245) );
  XOR U1564 ( .A(n1716), .B(n1715), .Z(n1717) );
  XOR U1565 ( .A(n1078), .B(n1077), .Z(n1079) );
  XOR U1566 ( .A(n3077), .B(n3076), .Z(n3078) );
  XOR U1567 ( .A(n3089), .B(n3088), .Z(n3090) );
  XOR U1568 ( .A(n2437), .B(n2436), .Z(n2438) );
  XOR U1569 ( .A(n2190), .B(n2189), .Z(n2191) );
  XOR U1570 ( .A(n2660), .B(n2659), .Z(n2661) );
  XOR U1571 ( .A(n2739), .B(n2738), .Z(n2740) );
  XOR U1572 ( .A(n2250), .B(n2249), .Z(n2251) );
  XOR U1573 ( .A(n2329), .B(n2328), .Z(n2330) );
  XOR U1574 ( .A(n2311), .B(n2310), .Z(n2312) );
  XOR U1575 ( .A(n2400), .B(n2399), .Z(n2401) );
  XOR U1576 ( .A(n524), .B(n523), .Z(n525) );
  XOR U1577 ( .A(n3163), .B(n3162), .Z(n3164) );
  XOR U1578 ( .A(n2208), .B(n2207), .Z(n2209) );
  XOR U1579 ( .A(n2034), .B(n2033), .Z(n2035) );
  XOR U1580 ( .A(n2467), .B(n2466), .Z(n2468) );
  XOR U1581 ( .A(n1201), .B(n1200), .Z(n1202) );
  XOR U1582 ( .A(n3017), .B(n3016), .Z(n3018) );
  XOR U1583 ( .A(n2999), .B(n2998), .Z(n3000) );
  XOR U1584 ( .A(n2461), .B(n2460), .Z(n2462) );
  XOR U1585 ( .A(n3223), .B(n3222), .Z(n3224) );
  XOR U1586 ( .A(n1422), .B(n1421), .Z(n1423) );
  XOR U1587 ( .A(n1834), .B(n1833), .Z(n1835) );
  XOR U1588 ( .A(n1747), .B(n1746), .Z(n1748) );
  XOR U1589 ( .A(n728), .B(n727), .Z(n729) );
  XOR U1590 ( .A(n2799), .B(n2798), .Z(n2800) );
  XOR U1591 ( .A(n2847), .B(n2846), .Z(n2848) );
  XOR U1592 ( .A(n1566), .B(n1565), .Z(n1567) );
  XOR U1593 ( .A(n3065), .B(n3064), .Z(n3066) );
  XOR U1594 ( .A(n2214), .B(n2213), .Z(n2215) );
  XOR U1595 ( .A(n2202), .B(n2201), .Z(n2203) );
  XOR U1596 ( .A(n2835), .B(n2834), .Z(n2836) );
  XOR U1597 ( .A(n1366), .B(n1365), .Z(n1367) );
  XOR U1598 ( .A(n4273), .B(n4272), .Z(n4275) );
  XOR U1599 ( .A(n4267), .B(n4266), .Z(n4268) );
  XOR U1600 ( .A(n4543), .B(n4542), .Z(n4545) );
  XOR U1601 ( .A(n4537), .B(n4536), .Z(n4539) );
  XOR U1602 ( .A(n3340), .B(n3339), .Z(n3342) );
  XOR U1603 ( .A(n3974), .B(n3973), .Z(n3976) );
  XOR U1604 ( .A(n4387), .B(n4386), .Z(n4389) );
  XOR U1605 ( .A(n3299), .B(n3298), .Z(n3301) );
  XOR U1606 ( .A(n4058), .B(n4057), .Z(n4060) );
  XOR U1607 ( .A(n4064), .B(n4063), .Z(n4066) );
  XOR U1608 ( .A(n4073), .B(n4072), .Z(n4075) );
  XOR U1609 ( .A(n4567), .B(n4566), .Z(n4569) );
  XOR U1610 ( .A(n4561), .B(n4560), .Z(n4563) );
  XOR U1611 ( .A(n4206), .B(n4205), .Z(n4207) );
  XOR U1612 ( .A(n3621), .B(n3620), .Z(n3623) );
  XOR U1613 ( .A(n3884), .B(n3883), .Z(n3886) );
  XOR U1614 ( .A(n4513), .B(n4512), .Z(n4515) );
  XOR U1615 ( .A(n4507), .B(n4506), .Z(n4509) );
  XOR U1616 ( .A(n4411), .B(n4410), .Z(n4413) );
  XOR U1617 ( .A(n4405), .B(n4404), .Z(n4407) );
  XOR U1618 ( .A(n3831), .B(n3830), .Z(n3833) );
  XOR U1619 ( .A(n3837), .B(n3836), .Z(n3839) );
  XOR U1620 ( .A(n3284), .B(n3283), .Z(n3286) );
  XOR U1621 ( .A(n3908), .B(n3907), .Z(n3910) );
  XOR U1622 ( .A(n4224), .B(n4223), .Z(n4226) );
  XOR U1623 ( .A(n4182), .B(n4181), .Z(n4184) );
  XOR U1624 ( .A(n4101), .B(n4100), .Z(n4103) );
  XOR U1625 ( .A(n3938), .B(n3937), .Z(n3940) );
  XOR U1626 ( .A(n4078), .B(n4079), .Z(n180) );
  XNOR U1627 ( .A(n4080), .B(n180), .Z(n3351) );
  XOR U1628 ( .A(n4489), .B(n4488), .Z(n4490) );
  XOR U1629 ( .A(n3730), .B(n3729), .Z(n3731) );
  XNOR U1630 ( .A(n4419), .B(n4418), .Z(n3738) );
  XOR U1631 ( .A(n4145), .B(n4144), .Z(n4464) );
  XOR U1632 ( .A(n3896), .B(n3895), .Z(n3898) );
  XOR U1633 ( .A(n3586), .B(n3587), .Z(n181) );
  XNOR U1634 ( .A(n3588), .B(n181), .Z(n4242) );
  XNOR U1635 ( .A(n4365), .B(n4364), .Z(n4609) );
  XOR U1636 ( .A(n4054), .B(n4053), .Z(n4607) );
  XOR U1637 ( .A(n2993), .B(n2992), .Z(n2994) );
  XOR U1638 ( .A(n1620), .B(n1619), .Z(n1621) );
  XOR U1639 ( .A(n1476), .B(n1475), .Z(n1477) );
  XOR U1640 ( .A(n3229), .B(n3228), .Z(n3230) );
  XOR U1641 ( .A(n2527), .B(n2526), .Z(n2528) );
  XOR U1642 ( .A(n2491), .B(n2490), .Z(n2492) );
  XOR U1643 ( .A(n2690), .B(n2689), .Z(n2691) );
  XOR U1644 ( .A(n976), .B(n975), .Z(n977) );
  XOR U1645 ( .A(n2933), .B(n2932), .Z(n2934) );
  XOR U1646 ( .A(n3029), .B(n3028), .Z(n3030) );
  XOR U1647 ( .A(n3095), .B(n3094), .Z(n3096) );
  XOR U1648 ( .A(n3169), .B(n3168), .Z(n3170) );
  XOR U1649 ( .A(n3718), .B(n3717), .Z(n3719) );
  XOR U1650 ( .A(n2878), .B(n2877), .Z(n2879) );
  XOR U1651 ( .A(n1102), .B(n1101), .Z(n1103) );
  XOR U1652 ( .A(n1840), .B(n1839), .Z(n1841) );
  XOR U1653 ( .A(n3998), .B(n3997), .Z(n3999) );
  XNOR U1654 ( .A(n3952), .B(n3951), .Z(n4173) );
  XOR U1655 ( .A(n3364), .B(n3363), .Z(n3365) );
  XOR U1656 ( .A(n716), .B(n715), .Z(n717) );
  NAND U1657 ( .A(n3296), .B(n3297), .Z(n182) );
  XOR U1658 ( .A(n3296), .B(n3297), .Z(n183) );
  NANDN U1659 ( .A(n3295), .B(n183), .Z(n184) );
  NAND U1660 ( .A(n182), .B(n184), .Z(n5006) );
  NAND U1661 ( .A(n3687), .B(n3688), .Z(n185) );
  XOR U1662 ( .A(n3687), .B(n3688), .Z(n186) );
  NANDN U1663 ( .A(n3686), .B(n186), .Z(n187) );
  NAND U1664 ( .A(n185), .B(n187), .Z(n5004) );
  XNOR U1665 ( .A(n4909), .B(n4908), .Z(n4999) );
  XOR U1666 ( .A(n5265), .B(n5264), .Z(n5266) );
  XNOR U1667 ( .A(n5165), .B(n5164), .Z(n4890) );
  NAND U1668 ( .A(n3346), .B(n3347), .Z(n188) );
  XOR U1669 ( .A(n3346), .B(n3347), .Z(n189) );
  NANDN U1670 ( .A(n3345), .B(n189), .Z(n190) );
  NAND U1671 ( .A(n188), .B(n190), .Z(n5301) );
  XOR U1672 ( .A(n5295), .B(n5294), .Z(n5296) );
  XOR U1673 ( .A(n5070), .B(n5069), .Z(n5071) );
  XOR U1674 ( .A(n5064), .B(n5063), .Z(n5066) );
  NAND U1675 ( .A(n3305), .B(n3306), .Z(n191) );
  XOR U1676 ( .A(n3305), .B(n3306), .Z(n192) );
  NANDN U1677 ( .A(n3304), .B(n192), .Z(n193) );
  NAND U1678 ( .A(n191), .B(n193), .Z(n4806) );
  NAND U1679 ( .A(n3583), .B(n3585), .Z(n194) );
  XOR U1680 ( .A(n3583), .B(n3585), .Z(n195) );
  NAND U1681 ( .A(n195), .B(n3584), .Z(n196) );
  NAND U1682 ( .A(n194), .B(n196), .Z(n4803) );
  XOR U1683 ( .A(n5271), .B(n5270), .Z(n5272) );
  XOR U1684 ( .A(n5046), .B(n5045), .Z(n5047) );
  XOR U1685 ( .A(n5040), .B(n5039), .Z(n5041) );
  NAND U1686 ( .A(n3290), .B(n3291), .Z(n197) );
  XOR U1687 ( .A(n3290), .B(n3291), .Z(n198) );
  NANDN U1688 ( .A(n3289), .B(n198), .Z(n199) );
  NAND U1689 ( .A(n197), .B(n199), .Z(n5277) );
  XOR U1690 ( .A(n5283), .B(n5282), .Z(n5284) );
  NAND U1691 ( .A(n3453), .B(n3452), .Z(n200) );
  XOR U1692 ( .A(n3453), .B(n3452), .Z(n201) );
  NANDN U1693 ( .A(n3454), .B(n201), .Z(n202) );
  NAND U1694 ( .A(n200), .B(n202), .Z(n4854) );
  XOR U1695 ( .A(n5088), .B(n5087), .Z(n5089) );
  XNOR U1696 ( .A(n5291), .B(n5290), .Z(n4975) );
  XNOR U1697 ( .A(n5159), .B(n5158), .Z(n5181) );
  NAND U1698 ( .A(n3736), .B(n3737), .Z(n203) );
  XOR U1699 ( .A(n3736), .B(n3737), .Z(n204) );
  NANDN U1700 ( .A(n3735), .B(n204), .Z(n205) );
  NAND U1701 ( .A(n203), .B(n205), .Z(n4931) );
  XOR U1702 ( .A(n4850), .B(n4849), .Z(n4792) );
  XOR U1703 ( .A(n5058), .B(n5057), .Z(n5060) );
  XNOR U1704 ( .A(n5078), .B(n5077), .Z(n4819) );
  XOR U1705 ( .A(n5313), .B(n5312), .Z(n5314) );
  XNOR U1706 ( .A(n4844), .B(n4843), .Z(n5308) );
  XOR U1707 ( .A(n2002), .B(n2001), .Z(n2003) );
  XOR U1708 ( .A(n3193), .B(n3192), .Z(n3194) );
  XOR U1709 ( .A(n2412), .B(n2411), .Z(n2413) );
  XOR U1710 ( .A(n2517), .B(n2516), .Z(n2007) );
  XOR U1711 ( .A(n2046), .B(n2045), .Z(n2047) );
  XOR U1712 ( .A(n3107), .B(n3106), .Z(n3109) );
  XNOR U1713 ( .A(n3714), .B(n3713), .Z(n3388) );
  XOR U1714 ( .A(n2547), .B(n2546), .Z(n1931) );
  XOR U1715 ( .A(n3807), .B(n3806), .Z(n3808) );
  XOR U1716 ( .A(n4503), .B(n4502), .Z(n3397) );
  XOR U1717 ( .A(n2594), .B(n2593), .Z(n1889) );
  XOR U1718 ( .A(n3530), .B(n3529), .Z(n3531) );
  XOR U1719 ( .A(n3332), .B(n3334), .Z(n206) );
  XNOR U1720 ( .A(n3335), .B(n206), .Z(n3511) );
  XOR U1721 ( .A(n3669), .B(n3668), .Z(n3671) );
  XOR U1722 ( .A(n4194), .B(n4193), .Z(n4196) );
  XOR U1723 ( .A(n3627), .B(n3626), .Z(n3628) );
  XOR U1724 ( .A(n4799), .B(n4798), .Z(n4692) );
  XOR U1725 ( .A(n4279), .B(n4278), .Z(n4280) );
  XOR U1726 ( .A(n5054), .B(n5053), .Z(n4966) );
  XOR U1727 ( .A(n5223), .B(n5222), .Z(n5225) );
  XOR U1728 ( .A(n5115), .B(n5114), .Z(n5010) );
  XNOR U1729 ( .A(n5177), .B(n5176), .Z(n5205) );
  XOR U1730 ( .A(n5199), .B(n5198), .Z(n5201) );
  XOR U1731 ( .A(n5481), .B(n5480), .Z(n5482) );
  XOR U1732 ( .A(n5463), .B(n5462), .Z(n5464) );
  XOR U1733 ( .A(n5636), .B(n5635), .Z(n5637) );
  XOR U1734 ( .A(n5606), .B(n5605), .Z(n5607) );
  NAND U1735 ( .A(n4769), .B(n4770), .Z(n207) );
  XOR U1736 ( .A(n4769), .B(n4770), .Z(n208) );
  NANDN U1737 ( .A(n4768), .B(n208), .Z(n209) );
  NAND U1738 ( .A(n207), .B(n209), .Z(n5654) );
  XOR U1739 ( .A(n5648), .B(n5647), .Z(n5649) );
  XOR U1740 ( .A(n5602), .B(n5601), .Z(n5672) );
  XOR U1741 ( .A(n5664), .B(n5663), .Z(n5666) );
  XOR U1742 ( .A(n5560), .B(n5559), .Z(n5561) );
  XOR U1743 ( .A(n5659), .B(n5660), .Z(n210) );
  XNOR U1744 ( .A(n5661), .B(n210), .Z(n5553) );
  XOR U1745 ( .A(n4786), .B(n4787), .Z(n211) );
  NANDN U1746 ( .A(n4788), .B(n211), .Z(n212) );
  NAND U1747 ( .A(n4786), .B(n4787), .Z(n213) );
  AND U1748 ( .A(n212), .B(n213), .Z(n5594) );
  XOR U1749 ( .A(n5705), .B(n5704), .Z(n5706) );
  XOR U1750 ( .A(n5701), .B(n5700), .Z(n5581) );
  XNOR U1751 ( .A(n5632), .B(n5631), .Z(n5534) );
  XOR U1752 ( .A(n5445), .B(n5444), .Z(n5446) );
  XOR U1753 ( .A(n5676), .B(n5675), .Z(n5677) );
  XNOR U1754 ( .A(n2258), .B(n2257), .Z(n1925) );
  XOR U1755 ( .A(n1961), .B(n1960), .Z(n1962) );
  XNOR U1756 ( .A(n2148), .B(n2147), .Z(n1968) );
  XNOR U1757 ( .A(n3013), .B(n3012), .Z(n2135) );
  XOR U1758 ( .A(n2727), .B(n2726), .Z(n2729) );
  XOR U1759 ( .A(n2723), .B(n2722), .Z(n2780) );
  XOR U1760 ( .A(n1300), .B(n1299), .Z(n1064) );
  XOR U1761 ( .A(n1110), .B(n1109), .Z(n1849) );
  XNOR U1762 ( .A(n4618), .B(n4617), .Z(n214) );
  XNOR U1763 ( .A(n4619), .B(n214), .Z(n3416) );
  NAND U1764 ( .A(n3404), .B(n3405), .Z(n215) );
  XOR U1765 ( .A(n3404), .B(n3405), .Z(n216) );
  NANDN U1766 ( .A(n3403), .B(n216), .Z(n217) );
  NAND U1767 ( .A(n215), .B(n217), .Z(n4925) );
  XOR U1768 ( .A(n3653), .B(n3652), .Z(n3477) );
  XOR U1769 ( .A(n3560), .B(n3559), .Z(n3562) );
  XOR U1770 ( .A(n3803), .B(n3802), .Z(n3520) );
  XOR U1771 ( .A(n3411), .B(n3410), .Z(n3412) );
  XOR U1772 ( .A(n5084), .B(n5083), .Z(n5029) );
  XNOR U1773 ( .A(n4885), .B(n4884), .Z(n4948) );
  XOR U1774 ( .A(n5241), .B(n5240), .Z(n5242) );
  XOR U1775 ( .A(n4953), .B(n4952), .Z(n4954) );
  NANDN U1776 ( .A(n4148), .B(n4151), .Z(n218) );
  OR U1777 ( .A(n4151), .B(n4150), .Z(n219) );
  NAND U1778 ( .A(n4149), .B(n219), .Z(n220) );
  NAND U1779 ( .A(n218), .B(n220), .Z(n5119) );
  XNOR U1780 ( .A(n5511), .B(n5510), .Z(n5513) );
  XNOR U1781 ( .A(n5519), .B(n5518), .Z(n5689) );
  NAND U1782 ( .A(n4760), .B(n4761), .Z(n221) );
  XOR U1783 ( .A(n4760), .B(n4761), .Z(n222) );
  NANDN U1784 ( .A(n4759), .B(n222), .Z(n223) );
  NAND U1785 ( .A(n221), .B(n223), .Z(n5421) );
  XNOR U1786 ( .A(n5584), .B(n5585), .Z(n224) );
  XNOR U1787 ( .A(n5586), .B(n224), .Z(n5439) );
  XOR U1788 ( .A(n5832), .B(n5831), .Z(n5833) );
  XNOR U1789 ( .A(n5756), .B(n5755), .Z(n5791) );
  XNOR U1790 ( .A(n2911), .B(n2910), .Z(n2343) );
  XOR U1791 ( .A(n2787), .B(n2786), .Z(n2789) );
  XOR U1792 ( .A(n3101), .B(n3100), .Z(n3103) );
  XNOR U1793 ( .A(n3635), .B(n3634), .Z(n3394) );
  XOR U1794 ( .A(n3665), .B(n3664), .Z(n3775) );
  NAND U1795 ( .A(n3766), .B(n3767), .Z(n225) );
  XOR U1796 ( .A(n3766), .B(n3767), .Z(n226) );
  NANDN U1797 ( .A(n3765), .B(n226), .Z(n227) );
  NAND U1798 ( .A(n225), .B(n227), .Z(n4832) );
  XOR U1799 ( .A(n5237), .B(n5236), .Z(n4681) );
  XOR U1800 ( .A(n5409), .B(n5408), .Z(n5411) );
  XOR U1801 ( .A(n5525), .B(n5524), .Z(n5486) );
  XOR U1802 ( .A(n5730), .B(n5729), .Z(n5732) );
  XOR U1803 ( .A(n5978), .B(n5977), .Z(n5980) );
  XOR U1804 ( .A(n5972), .B(n5971), .Z(n5973) );
  XOR U1805 ( .A(n5966), .B(n5965), .Z(n5968) );
  XOR U1806 ( .A(n5984), .B(n5983), .Z(n5985) );
  XOR U1807 ( .A(n5955), .B(n5954), .Z(n5957) );
  XOR U1808 ( .A(n5996), .B(n5995), .Z(n5998) );
  XOR U1809 ( .A(n5990), .B(n5989), .Z(n5991) );
  XOR U1810 ( .A(n5344), .B(n5343), .Z(n5346) );
  NAND U1811 ( .A(n2632), .B(n2631), .Z(n228) );
  NANDN U1812 ( .A(n2633), .B(n2634), .Z(n229) );
  AND U1813 ( .A(n228), .B(n229), .Z(n3494) );
  XOR U1814 ( .A(n5390), .B(n5389), .Z(n5723) );
  XOR U1815 ( .A(n5901), .B(n5900), .Z(n5887) );
  XNOR U1816 ( .A(n5925), .B(n5924), .Z(n5927) );
  XNOR U1817 ( .A(n4024), .B(n4023), .Z(n3488) );
  XOR U1818 ( .A(n5363), .B(n5362), .Z(n5364) );
  XNOR U1819 ( .A(n5951), .B(n5950), .Z(n5945) );
  XNOR U1820 ( .A(n5881), .B(n5880), .Z(n5883) );
  XOR U1821 ( .A(n6069), .B(n6068), .Z(n6061) );
  NAND U1822 ( .A(n5406), .B(n5407), .Z(n230) );
  XOR U1823 ( .A(n5406), .B(n5407), .Z(n231) );
  NANDN U1824 ( .A(n5405), .B(n231), .Z(n232) );
  NAND U1825 ( .A(n230), .B(n232), .Z(n5906) );
  NAND U1826 ( .A(n6050), .B(n6052), .Z(n233) );
  XOR U1827 ( .A(n6050), .B(n6052), .Z(n234) );
  NAND U1828 ( .A(n234), .B(n6051), .Z(n235) );
  NAND U1829 ( .A(n233), .B(n235), .Z(n6078) );
  NAND U1830 ( .A(n6090), .B(n6091), .Z(n236) );
  XOR U1831 ( .A(n6090), .B(n6091), .Z(n237) );
  NAND U1832 ( .A(n237), .B(oglobal[9]), .Z(n238) );
  NAND U1833 ( .A(n236), .B(n238), .Z(n6092) );
  XOR U1834 ( .A(x[266]), .B(y[266]), .Z(n2240) );
  XOR U1835 ( .A(x[177]), .B(y[177]), .Z(n2237) );
  XNOR U1836 ( .A(x[270]), .B(y[270]), .Z(n2238) );
  XNOR U1837 ( .A(n2237), .B(n2238), .Z(n2239) );
  XOR U1838 ( .A(n2240), .B(n2239), .Z(n1325) );
  XOR U1839 ( .A(x[256]), .B(y[256]), .Z(n2301) );
  XOR U1840 ( .A(x[258]), .B(y[258]), .Z(n2298) );
  XNOR U1841 ( .A(x[260]), .B(y[260]), .Z(n2299) );
  XNOR U1842 ( .A(n2298), .B(n2299), .Z(n2300) );
  XOR U1843 ( .A(n2301), .B(n2300), .Z(n1323) );
  XOR U1844 ( .A(x[230]), .B(y[230]), .Z(n2656) );
  XOR U1845 ( .A(x[195]), .B(y[195]), .Z(n2653) );
  XNOR U1846 ( .A(x[232]), .B(y[232]), .Z(n2654) );
  XNOR U1847 ( .A(n2653), .B(n2654), .Z(n2655) );
  XNOR U1848 ( .A(n2656), .B(n2655), .Z(n1322) );
  XNOR U1849 ( .A(n1323), .B(n1322), .Z(n1324) );
  XNOR U1850 ( .A(n1325), .B(n1324), .Z(n3100) );
  XOR U1851 ( .A(x[208]), .B(y[208]), .Z(n936) );
  XOR U1852 ( .A(x[210]), .B(y[210]), .Z(n933) );
  XNOR U1853 ( .A(x[216]), .B(y[216]), .Z(n934) );
  XNOR U1854 ( .A(n933), .B(n934), .Z(n935) );
  XOR U1855 ( .A(n936), .B(n935), .Z(n1818) );
  XOR U1856 ( .A(x[170]), .B(y[170]), .Z(n2463) );
  XOR U1857 ( .A(x[172]), .B(y[172]), .Z(n2460) );
  XOR U1858 ( .A(x[176]), .B(y[176]), .Z(n2461) );
  XOR U1859 ( .A(n2463), .B(n2462), .Z(n1816) );
  XOR U1860 ( .A(x[154]), .B(y[154]), .Z(n3147) );
  XOR U1861 ( .A(x[160]), .B(y[160]), .Z(n3144) );
  XOR U1862 ( .A(x[166]), .B(y[166]), .Z(n3145) );
  XNOR U1863 ( .A(n3147), .B(n3146), .Z(n1815) );
  XNOR U1864 ( .A(n1816), .B(n1815), .Z(n1817) );
  XNOR U1865 ( .A(n1818), .B(n1817), .Z(n3101) );
  XOR U1866 ( .A(x[148]), .B(y[148]), .Z(n368) );
  XOR U1867 ( .A(x[150]), .B(y[150]), .Z(n365) );
  XNOR U1868 ( .A(x[231]), .B(y[231]), .Z(n366) );
  XNOR U1869 ( .A(n365), .B(n366), .Z(n367) );
  XOR U1870 ( .A(n368), .B(n367), .Z(n1824) );
  XOR U1871 ( .A(x[142]), .B(y[142]), .Z(n3171) );
  XOR U1872 ( .A(x[144]), .B(y[144]), .Z(n3168) );
  XOR U1873 ( .A(x[235]), .B(y[235]), .Z(n3169) );
  XOR U1874 ( .A(n3171), .B(n3170), .Z(n1822) );
  XOR U1875 ( .A(x[126]), .B(y[126]), .Z(n308) );
  XOR U1876 ( .A(x[132]), .B(y[132]), .Z(n305) );
  XNOR U1877 ( .A(x[138]), .B(y[138]), .Z(n306) );
  XNOR U1878 ( .A(n305), .B(n306), .Z(n307) );
  XNOR U1879 ( .A(n308), .B(n307), .Z(n1821) );
  XNOR U1880 ( .A(n1822), .B(n1821), .Z(n1823) );
  XNOR U1881 ( .A(n1824), .B(n1823), .Z(n3102) );
  XOR U1882 ( .A(n3103), .B(n3102), .Z(n2717) );
  XOR U1883 ( .A(x[60]), .B(y[60]), .Z(n2825) );
  XOR U1884 ( .A(x[62]), .B(y[62]), .Z(n2822) );
  XNOR U1885 ( .A(x[271]), .B(y[271]), .Z(n2823) );
  XNOR U1886 ( .A(n2822), .B(n2823), .Z(n2824) );
  XNOR U1887 ( .A(n2825), .B(n2824), .Z(n1300) );
  XOR U1888 ( .A(x[52]), .B(y[52]), .Z(n2831) );
  XOR U1889 ( .A(x[56]), .B(y[56]), .Z(n2828) );
  XNOR U1890 ( .A(x[58]), .B(y[58]), .Z(n2829) );
  XNOR U1891 ( .A(n2828), .B(n2829), .Z(n2830) );
  XNOR U1892 ( .A(n2831), .B(n2830), .Z(n1298) );
  XOR U1893 ( .A(x[44]), .B(y[44]), .Z(n1172) );
  XOR U1894 ( .A(x[46]), .B(y[46]), .Z(n1169) );
  XNOR U1895 ( .A(x[48]), .B(y[48]), .Z(n1170) );
  XNOR U1896 ( .A(n1169), .B(n1170), .Z(n1171) );
  XNOR U1897 ( .A(n1172), .B(n1171), .Z(n1297) );
  XOR U1898 ( .A(x[88]), .B(y[88]), .Z(n502) );
  XOR U1899 ( .A(x[92]), .B(y[92]), .Z(n499) );
  XNOR U1900 ( .A(x[94]), .B(y[94]), .Z(n500) );
  XNOR U1901 ( .A(n499), .B(n500), .Z(n501) );
  XOR U1902 ( .A(n502), .B(n501), .Z(n724) );
  XOR U1903 ( .A(x[76]), .B(y[76]), .Z(n490) );
  XOR U1904 ( .A(x[82]), .B(y[82]), .Z(n487) );
  XNOR U1905 ( .A(x[84]), .B(y[84]), .Z(n488) );
  XNOR U1906 ( .A(n487), .B(n488), .Z(n489) );
  XOR U1907 ( .A(n490), .B(n489), .Z(n722) );
  XOR U1908 ( .A(x[66]), .B(y[66]), .Z(n272) );
  XOR U1909 ( .A(x[70]), .B(y[70]), .Z(n269) );
  XNOR U1910 ( .A(x[267]), .B(y[267]), .Z(n270) );
  XNOR U1911 ( .A(n269), .B(n270), .Z(n271) );
  XNOR U1912 ( .A(n272), .B(n271), .Z(n721) );
  XNOR U1913 ( .A(n722), .B(n721), .Z(n723) );
  XNOR U1914 ( .A(n724), .B(n723), .Z(n1062) );
  XOR U1915 ( .A(x[116]), .B(y[116]), .Z(n314) );
  XOR U1916 ( .A(x[120]), .B(y[120]), .Z(n311) );
  XNOR U1917 ( .A(x[122]), .B(y[122]), .Z(n312) );
  XNOR U1918 ( .A(n311), .B(n312), .Z(n313) );
  XOR U1919 ( .A(n314), .B(n313), .Z(n1430) );
  XOR U1920 ( .A(x[110]), .B(y[110]), .Z(n302) );
  XOR U1921 ( .A(x[114]), .B(y[114]), .Z(n299) );
  XNOR U1922 ( .A(x[249]), .B(y[249]), .Z(n300) );
  XNOR U1923 ( .A(n299), .B(n300), .Z(n301) );
  XOR U1924 ( .A(n302), .B(n301), .Z(n1428) );
  XOR U1925 ( .A(x[98]), .B(y[98]), .Z(n332) );
  XOR U1926 ( .A(x[104]), .B(y[104]), .Z(n329) );
  XNOR U1927 ( .A(x[253]), .B(y[253]), .Z(n330) );
  XNOR U1928 ( .A(n329), .B(n330), .Z(n331) );
  XNOR U1929 ( .A(n332), .B(n331), .Z(n1427) );
  XNOR U1930 ( .A(n1428), .B(n1427), .Z(n1429) );
  XOR U1931 ( .A(n1430), .B(n1429), .Z(n1061) );
  XNOR U1932 ( .A(n1062), .B(n1061), .Z(n1063) );
  XOR U1933 ( .A(n1064), .B(n1063), .Z(n2715) );
  XOR U1934 ( .A(x[13]), .B(y[13]), .Z(n2959) );
  XOR U1935 ( .A(x[11]), .B(y[11]), .Z(n2956) );
  XNOR U1936 ( .A(x[321]), .B(y[321]), .Z(n2957) );
  XNOR U1937 ( .A(n2956), .B(n2957), .Z(n2958) );
  XOR U1938 ( .A(n2959), .B(n2958), .Z(n631) );
  XOR U1939 ( .A(x[7]), .B(y[7]), .Z(n1122) );
  XOR U1940 ( .A(x[1]), .B(y[1]), .Z(n1119) );
  XNOR U1941 ( .A(x[5]), .B(y[5]), .Z(n1120) );
  XNOR U1942 ( .A(n1119), .B(n1120), .Z(n1121) );
  XOR U1943 ( .A(n1122), .B(n1121), .Z(n632) );
  XOR U1944 ( .A(n631), .B(n632), .Z(n634) );
  XOR U1945 ( .A(x[2]), .B(y[2]), .Z(n1116) );
  XOR U1946 ( .A(x[4]), .B(y[4]), .Z(n1113) );
  XNOR U1947 ( .A(x[6]), .B(y[6]), .Z(n1114) );
  XNOR U1948 ( .A(n1113), .B(n1114), .Z(n1115) );
  XOR U1949 ( .A(n1116), .B(n1115), .Z(n633) );
  XOR U1950 ( .A(n634), .B(n633), .Z(n1495) );
  XOR U1951 ( .A(x[8]), .B(y[8]), .Z(n1128) );
  XOR U1952 ( .A(x[10]), .B(y[10]), .Z(n1125) );
  XNOR U1953 ( .A(x[307]), .B(y[307]), .Z(n1126) );
  XNOR U1954 ( .A(n1125), .B(n1126), .Z(n1127) );
  XOR U1955 ( .A(n1128), .B(n1127), .Z(n604) );
  XOR U1956 ( .A(x[12]), .B(y[12]), .Z(n2898) );
  XOR U1957 ( .A(x[16]), .B(y[16]), .Z(n2895) );
  XNOR U1958 ( .A(x[303]), .B(y[303]), .Z(n2896) );
  XNOR U1959 ( .A(n2895), .B(n2896), .Z(n2897) );
  XNOR U1960 ( .A(n2898), .B(n2897), .Z(n603) );
  XNOR U1961 ( .A(n604), .B(n603), .Z(n606) );
  XOR U1962 ( .A(x[20]), .B(y[20]), .Z(n2892) );
  XOR U1963 ( .A(x[22]), .B(y[22]), .Z(n2889) );
  XNOR U1964 ( .A(x[24]), .B(y[24]), .Z(n2890) );
  XNOR U1965 ( .A(n2889), .B(n2890), .Z(n2891) );
  XOR U1966 ( .A(n2892), .B(n2891), .Z(n605) );
  XOR U1967 ( .A(n606), .B(n605), .Z(n1494) );
  XOR U1968 ( .A(x[40]), .B(y[40]), .Z(n1160) );
  XOR U1969 ( .A(x[42]), .B(y[42]), .Z(n1157) );
  XNOR U1970 ( .A(x[285]), .B(y[285]), .Z(n1158) );
  XNOR U1971 ( .A(n1157), .B(n1158), .Z(n1159) );
  XOR U1972 ( .A(n1160), .B(n1159), .Z(n748) );
  XOR U1973 ( .A(x[34]), .B(y[34]), .Z(n1166) );
  XOR U1974 ( .A(x[38]), .B(y[38]), .Z(n1163) );
  XNOR U1975 ( .A(x[289]), .B(y[289]), .Z(n1164) );
  XNOR U1976 ( .A(n1163), .B(n1164), .Z(n1165) );
  XOR U1977 ( .A(n1166), .B(n1165), .Z(n746) );
  XOR U1978 ( .A(x[26]), .B(y[26]), .Z(n2904) );
  XOR U1979 ( .A(x[28]), .B(y[28]), .Z(n2901) );
  XNOR U1980 ( .A(x[30]), .B(y[30]), .Z(n2902) );
  XNOR U1981 ( .A(n2901), .B(n2902), .Z(n2903) );
  XNOR U1982 ( .A(n2904), .B(n2903), .Z(n745) );
  XNOR U1983 ( .A(n746), .B(n745), .Z(n747) );
  XNOR U1984 ( .A(n748), .B(n747), .Z(n1493) );
  XOR U1985 ( .A(n1494), .B(n1493), .Z(n1496) );
  XNOR U1986 ( .A(n1495), .B(n1496), .Z(n2714) );
  XNOR U1987 ( .A(n2715), .B(n2714), .Z(n2716) );
  XNOR U1988 ( .A(n2717), .B(n2716), .Z(n3256) );
  XOR U1989 ( .A(x[742]), .B(y[742]), .Z(n1282) );
  XOR U1990 ( .A(x[74]), .B(y[74]), .Z(n1279) );
  XOR U1991 ( .A(x[744]), .B(y[744]), .Z(n1280) );
  XOR U1992 ( .A(n1282), .B(n1281), .Z(n1016) );
  XOR U1993 ( .A(x[890]), .B(y[890]), .Z(n2917) );
  XOR U1994 ( .A(x[174]), .B(y[174]), .Z(n2914) );
  XOR U1995 ( .A(x[892]), .B(y[892]), .Z(n2915) );
  XOR U1996 ( .A(n2917), .B(n2916), .Z(n1014) );
  XOR U1997 ( .A(x[738]), .B(y[738]), .Z(n1270) );
  XOR U1998 ( .A(x[740]), .B(y[740]), .Z(n1267) );
  XOR U1999 ( .A(x[965]), .B(y[965]), .Z(n1268) );
  XNOR U2000 ( .A(n1270), .B(n1269), .Z(n1013) );
  XNOR U2001 ( .A(n1014), .B(n1013), .Z(n1015) );
  XNOR U2002 ( .A(n1016), .B(n1015), .Z(n2587) );
  XOR U2003 ( .A(x[734]), .B(y[734]), .Z(n1264) );
  XOR U2004 ( .A(x[68]), .B(y[68]), .Z(n1261) );
  XNOR U2005 ( .A(x[736]), .B(y[736]), .Z(n1262) );
  XNOR U2006 ( .A(n1261), .B(n1262), .Z(n1263) );
  XOR U2007 ( .A(n1264), .B(n1263), .Z(n1706) );
  XOR U2008 ( .A(x[894]), .B(y[894]), .Z(n2120) );
  XOR U2009 ( .A(x[178]), .B(y[178]), .Z(n2117) );
  XNOR U2010 ( .A(x[896]), .B(y[896]), .Z(n2118) );
  XNOR U2011 ( .A(n2117), .B(n2118), .Z(n2119) );
  XOR U2012 ( .A(n2120), .B(n2119), .Z(n1704) );
  XOR U2013 ( .A(x[730]), .B(y[730]), .Z(n3007) );
  XOR U2014 ( .A(x[64]), .B(y[64]), .Z(n3004) );
  XOR U2015 ( .A(x[732]), .B(y[732]), .Z(n3005) );
  XNOR U2016 ( .A(n3007), .B(n3006), .Z(n1703) );
  XNOR U2017 ( .A(n1704), .B(n1703), .Z(n1705) );
  XOR U2018 ( .A(n1706), .B(n1705), .Z(n2588) );
  XNOR U2019 ( .A(n2587), .B(n2588), .Z(n2590) );
  XOR U2020 ( .A(x[726]), .B(y[726]), .Z(n3001) );
  XOR U2021 ( .A(x[169]), .B(y[169]), .Z(n2998) );
  XOR U2022 ( .A(x[728]), .B(y[728]), .Z(n2999) );
  XNOR U2023 ( .A(n3001), .B(n3000), .Z(n3097) );
  XOR U2024 ( .A(x[898]), .B(y[898]), .Z(n2078) );
  XOR U2025 ( .A(x[900]), .B(y[900]), .Z(n2075) );
  XNOR U2026 ( .A(x[985]), .B(y[985]), .Z(n2076) );
  XNOR U2027 ( .A(n2075), .B(n2076), .Z(n2077) );
  XNOR U2028 ( .A(n2078), .B(n2077), .Z(n3095) );
  XOR U2029 ( .A(x[722]), .B(y[722]), .Z(n1532) );
  XOR U2030 ( .A(x[326]), .B(y[326]), .Z(n1529) );
  XNOR U2031 ( .A(x[724]), .B(y[724]), .Z(n1530) );
  XNOR U2032 ( .A(n1529), .B(n1530), .Z(n1531) );
  XNOR U2033 ( .A(n1532), .B(n1531), .Z(n3094) );
  XNOR U2034 ( .A(n2590), .B(n2589), .Z(n2781) );
  XOR U2035 ( .A(x[794]), .B(y[794]), .Z(n2977) );
  XOR U2036 ( .A(x[108]), .B(y[108]), .Z(n2974) );
  XOR U2037 ( .A(x[796]), .B(y[796]), .Z(n2975) );
  XOR U2038 ( .A(n2977), .B(n2976), .Z(n2841) );
  XOR U2039 ( .A(x[862]), .B(y[862]), .Z(n2983) );
  XOR U2040 ( .A(x[156]), .B(y[156]), .Z(n2980) );
  XOR U2041 ( .A(x[864]), .B(y[864]), .Z(n2981) );
  XOR U2042 ( .A(n2983), .B(n2982), .Z(n2840) );
  XOR U2043 ( .A(n2841), .B(n2840), .Z(n2843) );
  XOR U2044 ( .A(x[798]), .B(y[798]), .Z(n1681) );
  XOR U2045 ( .A(x[112]), .B(y[112]), .Z(n1679) );
  XNOR U2046 ( .A(x[800]), .B(y[800]), .Z(n1680) );
  XOR U2047 ( .A(n1679), .B(n1680), .Z(n1682) );
  XNOR U2048 ( .A(n1681), .B(n1682), .Z(n2842) );
  XNOR U2049 ( .A(n2843), .B(n2842), .Z(n2723) );
  XOR U2050 ( .A(x[806]), .B(y[806]), .Z(n1628) );
  XOR U2051 ( .A(x[118]), .B(y[118]), .Z(n1625) );
  XOR U2052 ( .A(x[808]), .B(y[808]), .Z(n1626) );
  XOR U2053 ( .A(n1628), .B(n1627), .Z(n1610) );
  XOR U2054 ( .A(x[858]), .B(y[858]), .Z(n2989) );
  XOR U2055 ( .A(x[152]), .B(y[152]), .Z(n2986) );
  XOR U2056 ( .A(x[860]), .B(y[860]), .Z(n2987) );
  XOR U2057 ( .A(n2989), .B(n2988), .Z(n1608) );
  XOR U2058 ( .A(x[802]), .B(y[802]), .Z(n1664) );
  XOR U2059 ( .A(x[804]), .B(y[804]), .Z(n1661) );
  XOR U2060 ( .A(x[973]), .B(y[973]), .Z(n1662) );
  XNOR U2061 ( .A(n1664), .B(n1663), .Z(n1607) );
  XNOR U2062 ( .A(n1608), .B(n1607), .Z(n1609) );
  XNOR U2063 ( .A(n1610), .B(n1609), .Z(n2721) );
  XOR U2064 ( .A(x[830]), .B(y[830]), .Z(n3043) );
  XOR U2065 ( .A(x[134]), .B(y[134]), .Z(n3040) );
  XOR U2066 ( .A(x[832]), .B(y[832]), .Z(n3041) );
  XNOR U2067 ( .A(n3043), .B(n3042), .Z(n3055) );
  XOR U2068 ( .A(x[826]), .B(y[826]), .Z(n3049) );
  XOR U2069 ( .A(x[130]), .B(y[130]), .Z(n3046) );
  XOR U2070 ( .A(x[828]), .B(y[828]), .Z(n3047) );
  XNOR U2071 ( .A(n3049), .B(n3048), .Z(n3053) );
  XOR U2072 ( .A(x[838]), .B(y[838]), .Z(n1574) );
  XOR U2073 ( .A(x[140]), .B(y[140]), .Z(n1571) );
  XNOR U2074 ( .A(x[840]), .B(y[840]), .Z(n1572) );
  XNOR U2075 ( .A(n1571), .B(n1572), .Z(n1573) );
  XNOR U2076 ( .A(n1574), .B(n1573), .Z(n3052) );
  XOR U2077 ( .A(n2721), .B(n2720), .Z(n2722) );
  XOR U2078 ( .A(n2781), .B(n2780), .Z(n2783) );
  XOR U2079 ( .A(x[766]), .B(y[766]), .Z(n1670) );
  XOR U2080 ( .A(x[90]), .B(y[90]), .Z(n1667) );
  XNOR U2081 ( .A(x[768]), .B(y[768]), .Z(n1668) );
  XNOR U2082 ( .A(n1667), .B(n1668), .Z(n1669) );
  XNOR U2083 ( .A(n1670), .B(n1669), .Z(n2935) );
  XOR U2084 ( .A(x[878]), .B(y[878]), .Z(n1520) );
  XOR U2085 ( .A(x[75]), .B(y[75]), .Z(n1517) );
  XNOR U2086 ( .A(x[880]), .B(y[880]), .Z(n1518) );
  XNOR U2087 ( .A(n1517), .B(n1518), .Z(n1519) );
  XNOR U2088 ( .A(n1520), .B(n1519), .Z(n2933) );
  XOR U2089 ( .A(x[762]), .B(y[762]), .Z(n1562) );
  XOR U2090 ( .A(x[86]), .B(y[86]), .Z(n1559) );
  XNOR U2091 ( .A(x[764]), .B(y[764]), .Z(n1560) );
  XNOR U2092 ( .A(n1559), .B(n1560), .Z(n1561) );
  XNOR U2093 ( .A(n1562), .B(n1561), .Z(n2932) );
  XOR U2094 ( .A(x[758]), .B(y[758]), .Z(n3019) );
  XOR U2095 ( .A(x[149]), .B(y[149]), .Z(n3016) );
  XOR U2096 ( .A(x[760]), .B(y[760]), .Z(n3017) );
  XOR U2097 ( .A(n3019), .B(n3018), .Z(n1058) );
  XOR U2098 ( .A(x[882]), .B(y[882]), .Z(n1502) );
  XOR U2099 ( .A(x[168]), .B(y[168]), .Z(n1499) );
  XOR U2100 ( .A(x[884]), .B(y[884]), .Z(n1500) );
  XOR U2101 ( .A(n1502), .B(n1501), .Z(n1056) );
  XOR U2102 ( .A(x[754]), .B(y[754]), .Z(n3037) );
  XOR U2103 ( .A(x[80]), .B(y[80]), .Z(n3034) );
  XOR U2104 ( .A(x[756]), .B(y[756]), .Z(n3035) );
  XNOR U2105 ( .A(n3037), .B(n3036), .Z(n1055) );
  XNOR U2106 ( .A(n1056), .B(n1055), .Z(n1057) );
  XOR U2107 ( .A(n1058), .B(n1057), .Z(n2346) );
  XNOR U2108 ( .A(n2345), .B(n2346), .Z(n2347) );
  XOR U2109 ( .A(x[750]), .B(y[750]), .Z(n3031) );
  XOR U2110 ( .A(x[155]), .B(y[155]), .Z(n3028) );
  XOR U2111 ( .A(x[752]), .B(y[752]), .Z(n3029) );
  XOR U2112 ( .A(n3031), .B(n3030), .Z(n991) );
  XOR U2113 ( .A(x[886]), .B(y[886]), .Z(n1022) );
  XOR U2114 ( .A(x[69]), .B(y[69]), .Z(n1019) );
  XOR U2115 ( .A(x[888]), .B(y[888]), .Z(n1020) );
  XOR U2116 ( .A(n1022), .B(n1021), .Z(n989) );
  XOR U2117 ( .A(x[746]), .B(y[746]), .Z(n1568) );
  XOR U2118 ( .A(x[748]), .B(y[748]), .Z(n1565) );
  XOR U2119 ( .A(x[967]), .B(y[967]), .Z(n1566) );
  XNOR U2120 ( .A(n1568), .B(n1567), .Z(n988) );
  XNOR U2121 ( .A(n989), .B(n988), .Z(n990) );
  XOR U2122 ( .A(n991), .B(n990), .Z(n2348) );
  XNOR U2123 ( .A(n2347), .B(n2348), .Z(n2782) );
  XOR U2124 ( .A(n2783), .B(n2782), .Z(n3254) );
  XOR U2125 ( .A(x[502]), .B(y[502]), .Z(n1799) );
  XOR U2126 ( .A(x[54]), .B(y[54]), .Z(n1796) );
  XNOR U2127 ( .A(x[504]), .B(y[504]), .Z(n1797) );
  XNOR U2128 ( .A(n1796), .B(n1797), .Z(n1798) );
  XOR U2129 ( .A(n1799), .B(n1798), .Z(n2625) );
  XOR U2130 ( .A(x[498]), .B(y[498]), .Z(n1337) );
  XOR U2131 ( .A(x[50]), .B(y[50]), .Z(n1334) );
  XNOR U2132 ( .A(x[500]), .B(y[500]), .Z(n1335) );
  XNOR U2133 ( .A(n1334), .B(n1335), .Z(n1336) );
  XOR U2134 ( .A(n1337), .B(n1336), .Z(n2623) );
  XOR U2135 ( .A(x[492]), .B(y[492]), .Z(n1343) );
  XOR U2136 ( .A(x[494]), .B(y[494]), .Z(n1340) );
  XNOR U2137 ( .A(x[496]), .B(y[496]), .Z(n1341) );
  XNOR U2138 ( .A(n1340), .B(n1341), .Z(n1342) );
  XNOR U2139 ( .A(n1343), .B(n1342), .Z(n2622) );
  XNOR U2140 ( .A(n2623), .B(n2622), .Z(n2624) );
  XNOR U2141 ( .A(n2625), .B(n2624), .Z(n2726) );
  XOR U2142 ( .A(x[486]), .B(y[486]), .Z(n1349) );
  XOR U2143 ( .A(x[488]), .B(y[488]), .Z(n1346) );
  XNOR U2144 ( .A(x[490]), .B(y[490]), .Z(n1347) );
  XNOR U2145 ( .A(n1346), .B(n1347), .Z(n1348) );
  XOR U2146 ( .A(n1349), .B(n1348), .Z(n2354) );
  XOR U2147 ( .A(x[482]), .B(y[482]), .Z(n1454) );
  XOR U2148 ( .A(x[36]), .B(y[36]), .Z(n1451) );
  XNOR U2149 ( .A(x[484]), .B(y[484]), .Z(n1452) );
  XNOR U2150 ( .A(n1451), .B(n1452), .Z(n1453) );
  XOR U2151 ( .A(n1454), .B(n1453), .Z(n2352) );
  XOR U2152 ( .A(x[478]), .B(y[478]), .Z(n1442) );
  XOR U2153 ( .A(x[32]), .B(y[32]), .Z(n1439) );
  XNOR U2154 ( .A(x[480]), .B(y[480]), .Z(n1440) );
  XNOR U2155 ( .A(n1439), .B(n1440), .Z(n1441) );
  XNOR U2156 ( .A(n1442), .B(n1441), .Z(n2351) );
  XNOR U2157 ( .A(n2352), .B(n2351), .Z(n2353) );
  XNOR U2158 ( .A(n2354), .B(n2353), .Z(n2727) );
  XOR U2159 ( .A(x[472]), .B(y[472]), .Z(n2172) );
  XOR U2160 ( .A(x[474]), .B(y[474]), .Z(n2169) );
  XNOR U2161 ( .A(x[476]), .B(y[476]), .Z(n2170) );
  XNOR U2162 ( .A(n2169), .B(n2170), .Z(n2171) );
  XOR U2163 ( .A(n2172), .B(n2171), .Z(n2366) );
  XOR U2164 ( .A(x[466]), .B(y[466]), .Z(n2114) );
  XOR U2165 ( .A(x[468]), .B(y[468]), .Z(n2111) );
  XNOR U2166 ( .A(x[470]), .B(y[470]), .Z(n2112) );
  XNOR U2167 ( .A(n2111), .B(n2112), .Z(n2113) );
  XOR U2168 ( .A(n2114), .B(n2113), .Z(n2364) );
  XOR U2169 ( .A(x[462]), .B(y[462]), .Z(n1448) );
  XOR U2170 ( .A(x[18]), .B(y[18]), .Z(n1445) );
  XNOR U2171 ( .A(x[464]), .B(y[464]), .Z(n1446) );
  XNOR U2172 ( .A(n1445), .B(n1446), .Z(n1447) );
  XNOR U2173 ( .A(n1448), .B(n1447), .Z(n2363) );
  XNOR U2174 ( .A(n2364), .B(n2363), .Z(n2365) );
  XNOR U2175 ( .A(n2366), .B(n2365), .Z(n2728) );
  XOR U2176 ( .A(n2729), .B(n2728), .Z(n3243) );
  XOR U2177 ( .A(x[458]), .B(y[458]), .Z(n1368) );
  XOR U2178 ( .A(x[14]), .B(y[14]), .Z(n1365) );
  XOR U2179 ( .A(x[460]), .B(y[460]), .Z(n1366) );
  XOR U2180 ( .A(n1368), .B(n1367), .Z(n2559) );
  XOR U2181 ( .A(x[452]), .B(y[452]), .Z(n1356) );
  XOR U2182 ( .A(x[454]), .B(y[454]), .Z(n1353) );
  XOR U2183 ( .A(x[456]), .B(y[456]), .Z(n1354) );
  XOR U2184 ( .A(n1356), .B(n1355), .Z(n2557) );
  XOR U2185 ( .A(x[442]), .B(y[442]), .Z(n1362) );
  XOR U2186 ( .A(x[0]), .B(y[0]), .Z(n1359) );
  XOR U2187 ( .A(x[444]), .B(y[444]), .Z(n1360) );
  XNOR U2188 ( .A(n1362), .B(n1361), .Z(n2556) );
  XNOR U2189 ( .A(n2557), .B(n2556), .Z(n2558) );
  XNOR U2190 ( .A(n2559), .B(n2558), .Z(n245) );
  XOR U2191 ( .A(x[432]), .B(y[432]), .Z(n2837) );
  XOR U2192 ( .A(x[434]), .B(y[434]), .Z(n2834) );
  XOR U2193 ( .A(x[436]), .B(y[436]), .Z(n2835) );
  XOR U2194 ( .A(n2837), .B(n2836), .Z(n2600) );
  XOR U2195 ( .A(x[422]), .B(y[422]), .Z(n326) );
  XOR U2196 ( .A(x[21]), .B(y[21]), .Z(n323) );
  XOR U2197 ( .A(x[424]), .B(y[424]), .Z(n324) );
  XOR U2198 ( .A(n326), .B(n325), .Z(n2598) );
  XOR U2199 ( .A(x[412]), .B(y[412]), .Z(n3177) );
  XOR U2200 ( .A(x[414]), .B(y[414]), .Z(n3174) );
  XOR U2201 ( .A(x[416]), .B(y[416]), .Z(n3175) );
  XNOR U2202 ( .A(n3177), .B(n3176), .Z(n2597) );
  XNOR U2203 ( .A(n2598), .B(n2597), .Z(n2599) );
  XNOR U2204 ( .A(n2600), .B(n2599), .Z(n246) );
  XOR U2205 ( .A(n245), .B(n246), .Z(n248) );
  XOR U2206 ( .A(x[402]), .B(y[402]), .Z(n3141) );
  XOR U2207 ( .A(x[43]), .B(y[43]), .Z(n3138) );
  XNOR U2208 ( .A(x[404]), .B(y[404]), .Z(n3139) );
  XNOR U2209 ( .A(n3138), .B(n3139), .Z(n3140) );
  XNOR U2210 ( .A(n3141), .B(n3140), .Z(n718) );
  XOR U2211 ( .A(x[392]), .B(y[392]), .Z(n2396) );
  XOR U2212 ( .A(x[394]), .B(y[394]), .Z(n2393) );
  XNOR U2213 ( .A(x[396]), .B(y[396]), .Z(n2394) );
  XNOR U2214 ( .A(n2393), .B(n2394), .Z(n2395) );
  XNOR U2215 ( .A(n2396), .B(n2395), .Z(n716) );
  XOR U2216 ( .A(x[382]), .B(y[382]), .Z(n2765) );
  XOR U2217 ( .A(x[65]), .B(y[65]), .Z(n2762) );
  XNOR U2218 ( .A(x[384]), .B(y[384]), .Z(n2763) );
  XNOR U2219 ( .A(n2762), .B(n2763), .Z(n2764) );
  XNOR U2220 ( .A(n2765), .B(n2764), .Z(n715) );
  XOR U2221 ( .A(n248), .B(n247), .Z(n3241) );
  XOR U2222 ( .A(x[372]), .B(y[372]), .Z(n2704) );
  XOR U2223 ( .A(x[374]), .B(y[374]), .Z(n2701) );
  XNOR U2224 ( .A(x[376]), .B(y[376]), .Z(n2702) );
  XNOR U2225 ( .A(n2701), .B(n2702), .Z(n2703) );
  XOR U2226 ( .A(n2704), .B(n2703), .Z(n688) );
  XOR U2227 ( .A(x[362]), .B(y[362]), .Z(n3159) );
  XOR U2228 ( .A(x[87]), .B(y[87]), .Z(n3156) );
  XNOR U2229 ( .A(x[364]), .B(y[364]), .Z(n3157) );
  XNOR U2230 ( .A(n3156), .B(n3157), .Z(n3158) );
  XOR U2231 ( .A(n3159), .B(n3158), .Z(n686) );
  XOR U2232 ( .A(x[352]), .B(y[352]), .Z(n3153) );
  XOR U2233 ( .A(x[354]), .B(y[354]), .Z(n3150) );
  XNOR U2234 ( .A(x[356]), .B(y[356]), .Z(n3151) );
  XNOR U2235 ( .A(n3150), .B(n3151), .Z(n3152) );
  XNOR U2236 ( .A(n3153), .B(n3152), .Z(n685) );
  XNOR U2237 ( .A(n686), .B(n685), .Z(n687) );
  XNOR U2238 ( .A(n688), .B(n687), .Z(n3106) );
  XOR U2239 ( .A(x[342]), .B(y[342]), .Z(n3207) );
  XOR U2240 ( .A(x[111]), .B(y[111]), .Z(n3204) );
  XOR U2241 ( .A(x[344]), .B(y[344]), .Z(n3205) );
  XOR U2242 ( .A(n3207), .B(n3206), .Z(n755) );
  XOR U2243 ( .A(x[332]), .B(y[332]), .Z(n2372) );
  XOR U2244 ( .A(x[334]), .B(y[334]), .Z(n2369) );
  XNOR U2245 ( .A(x[336]), .B(y[336]), .Z(n2370) );
  XNOR U2246 ( .A(n2369), .B(n2370), .Z(n2371) );
  XOR U2247 ( .A(n2372), .B(n2371), .Z(n753) );
  XOR U2248 ( .A(x[318]), .B(y[318]), .Z(n2481) );
  XOR U2249 ( .A(x[133]), .B(y[133]), .Z(n2478) );
  XNOR U2250 ( .A(x[320]), .B(y[320]), .Z(n2479) );
  XNOR U2251 ( .A(n2478), .B(n2479), .Z(n2480) );
  XNOR U2252 ( .A(n2481), .B(n2480), .Z(n752) );
  XNOR U2253 ( .A(n753), .B(n752), .Z(n754) );
  XNOR U2254 ( .A(n755), .B(n754), .Z(n3107) );
  XOR U2255 ( .A(x[306]), .B(y[306]), .Z(n3225) );
  XOR U2256 ( .A(x[310]), .B(y[310]), .Z(n3222) );
  XOR U2257 ( .A(x[312]), .B(y[312]), .Z(n3223) );
  XOR U2258 ( .A(n3225), .B(n3224), .Z(n1406) );
  XOR U2259 ( .A(x[294]), .B(y[294]), .Z(n2186) );
  XOR U2260 ( .A(x[157]), .B(y[157]), .Z(n2183) );
  XOR U2261 ( .A(x[296]), .B(y[296]), .Z(n2184) );
  XOR U2262 ( .A(n2186), .B(n2185), .Z(n1404) );
  XOR U2263 ( .A(x[280]), .B(y[280]), .Z(n2222) );
  XOR U2264 ( .A(x[282]), .B(y[282]), .Z(n2219) );
  XOR U2265 ( .A(x[284]), .B(y[284]), .Z(n2220) );
  XNOR U2266 ( .A(n2222), .B(n2221), .Z(n1403) );
  XNOR U2267 ( .A(n1404), .B(n1403), .Z(n1405) );
  XNOR U2268 ( .A(n1406), .B(n1405), .Z(n3108) );
  XNOR U2269 ( .A(n3109), .B(n3108), .Z(n3240) );
  XNOR U2270 ( .A(n3241), .B(n3240), .Z(n3242) );
  XNOR U2271 ( .A(n3243), .B(n3242), .Z(n3253) );
  XNOR U2272 ( .A(n3254), .B(n3253), .Z(n3255) );
  XOR U2273 ( .A(n3256), .B(n3255), .Z(n240) );
  XOR U2274 ( .A(x[421]), .B(y[421]), .Z(n417) );
  XOR U2275 ( .A(x[419]), .B(y[419]), .Z(n414) );
  XNOR U2276 ( .A(x[689]), .B(y[689]), .Z(n415) );
  XNOR U2277 ( .A(n414), .B(n415), .Z(n416) );
  XOR U2278 ( .A(n417), .B(n416), .Z(n600) );
  XOR U2279 ( .A(x[406]), .B(y[406]), .Z(n3183) );
  XOR U2280 ( .A(x[408]), .B(y[408]), .Z(n3180) );
  XOR U2281 ( .A(x[410]), .B(y[410]), .Z(n3181) );
  XOR U2282 ( .A(n3183), .B(n3182), .Z(n598) );
  XOR U2283 ( .A(x[425]), .B(y[425]), .Z(n423) );
  XOR U2284 ( .A(x[423]), .B(y[423]), .Z(n420) );
  XNOR U2285 ( .A(x[901]), .B(y[901]), .Z(n421) );
  XNOR U2286 ( .A(n420), .B(n421), .Z(n422) );
  XNOR U2287 ( .A(n423), .B(n422), .Z(n597) );
  XNOR U2288 ( .A(n598), .B(n597), .Z(n599) );
  XNOR U2289 ( .A(n600), .B(n599), .Z(n2017) );
  XOR U2290 ( .A(x[429]), .B(y[429]), .Z(n1203) );
  XOR U2291 ( .A(x[427]), .B(y[427]), .Z(n1200) );
  XOR U2292 ( .A(x[693]), .B(y[693]), .Z(n1201) );
  XOR U2293 ( .A(n1203), .B(n1202), .Z(n435) );
  XOR U2294 ( .A(x[930]), .B(y[930]), .Z(n3135) );
  XOR U2295 ( .A(x[932]), .B(y[932]), .Z(n3132) );
  XOR U2296 ( .A(x[989]), .B(y[989]), .Z(n3133) );
  XOR U2297 ( .A(n3135), .B(n3134), .Z(n433) );
  XOR U2298 ( .A(x[433]), .B(y[433]), .Z(n1197) );
  XOR U2299 ( .A(x[431]), .B(y[431]), .Z(n1194) );
  XOR U2300 ( .A(x[899]), .B(y[899]), .Z(n1195) );
  XNOR U2301 ( .A(n1197), .B(n1196), .Z(n432) );
  XNOR U2302 ( .A(n433), .B(n432), .Z(n434) );
  XOR U2303 ( .A(n435), .B(n434), .Z(n2018) );
  XNOR U2304 ( .A(n2017), .B(n2018), .Z(n2020) );
  XOR U2305 ( .A(x[437]), .B(y[437]), .Z(n1191) );
  XOR U2306 ( .A(x[435]), .B(y[435]), .Z(n1188) );
  XNOR U2307 ( .A(x[697]), .B(y[697]), .Z(n1189) );
  XNOR U2308 ( .A(n1188), .B(n1189), .Z(n1190) );
  XOR U2309 ( .A(n1191), .B(n1190), .Z(n2126) );
  XOR U2310 ( .A(x[398]), .B(y[398]), .Z(n2469) );
  XOR U2311 ( .A(x[47]), .B(y[47]), .Z(n2466) );
  XOR U2312 ( .A(x[400]), .B(y[400]), .Z(n2467) );
  XOR U2313 ( .A(n2469), .B(n2468), .Z(n2124) );
  XOR U2314 ( .A(x[443]), .B(y[443]), .Z(n2108) );
  XOR U2315 ( .A(x[439]), .B(y[439]), .Z(n2105) );
  XNOR U2316 ( .A(x[441]), .B(y[441]), .Z(n2106) );
  XNOR U2317 ( .A(n2105), .B(n2106), .Z(n2107) );
  XNOR U2318 ( .A(n2108), .B(n2107), .Z(n2123) );
  XNOR U2319 ( .A(n2124), .B(n2123), .Z(n2125) );
  XOR U2320 ( .A(n2126), .B(n2125), .Z(n2019) );
  XNOR U2321 ( .A(n2020), .B(n2019), .Z(n2644) );
  XOR U2322 ( .A(x[449]), .B(y[449]), .Z(n2066) );
  XOR U2323 ( .A(x[445]), .B(y[445]), .Z(n2063) );
  XNOR U2324 ( .A(x[447]), .B(y[447]), .Z(n2064) );
  XNOR U2325 ( .A(n2063), .B(n2064), .Z(n2065) );
  XOR U2326 ( .A(n2066), .B(n2065), .Z(n2060) );
  XOR U2327 ( .A(x[934]), .B(y[934]), .Z(n2427) );
  XOR U2328 ( .A(x[206]), .B(y[206]), .Z(n2424) );
  XOR U2329 ( .A(x[936]), .B(y[936]), .Z(n2425) );
  XOR U2330 ( .A(n2427), .B(n2426), .Z(n2058) );
  XOR U2331 ( .A(x[455]), .B(y[455]), .Z(n2160) );
  XOR U2332 ( .A(x[451]), .B(y[451]), .Z(n2157) );
  XOR U2333 ( .A(x[453]), .B(y[453]), .Z(n2158) );
  XNOR U2334 ( .A(n2160), .B(n2159), .Z(n2057) );
  XNOR U2335 ( .A(n2058), .B(n2057), .Z(n2059) );
  XNOR U2336 ( .A(n2060), .B(n2059), .Z(n2051) );
  XOR U2337 ( .A(x[461]), .B(y[461]), .Z(n2042) );
  XOR U2338 ( .A(x[457]), .B(y[457]), .Z(n2039) );
  XOR U2339 ( .A(x[459]), .B(y[459]), .Z(n2040) );
  XOR U2340 ( .A(n2042), .B(n2041), .Z(n1898) );
  XOR U2341 ( .A(x[386]), .B(y[386]), .Z(n2505) );
  XOR U2342 ( .A(x[388]), .B(y[388]), .Z(n2502) );
  XOR U2343 ( .A(x[390]), .B(y[390]), .Z(n2503) );
  XOR U2344 ( .A(n2505), .B(n2504), .Z(n1896) );
  XOR U2345 ( .A(x[467]), .B(y[467]), .Z(n2030) );
  XOR U2346 ( .A(x[463]), .B(y[463]), .Z(n2027) );
  XOR U2347 ( .A(x[465]), .B(y[465]), .Z(n2028) );
  XNOR U2348 ( .A(n2030), .B(n2029), .Z(n1895) );
  XNOR U2349 ( .A(n1896), .B(n1895), .Z(n1897) );
  XOR U2350 ( .A(n1898), .B(n1897), .Z(n2052) );
  XNOR U2351 ( .A(n2051), .B(n2052), .Z(n2053) );
  XOR U2352 ( .A(x[473]), .B(y[473]), .Z(n2036) );
  XOR U2353 ( .A(x[469]), .B(y[469]), .Z(n2033) );
  XOR U2354 ( .A(x[471]), .B(y[471]), .Z(n2034) );
  XOR U2355 ( .A(n2036), .B(n2035), .Z(n1886) );
  XOR U2356 ( .A(x[938]), .B(y[938]), .Z(n2325) );
  XOR U2357 ( .A(x[940]), .B(y[940]), .Z(n2322) );
  XOR U2358 ( .A(x[991]), .B(y[991]), .Z(n2323) );
  XOR U2359 ( .A(n2325), .B(n2324), .Z(n1884) );
  XOR U2360 ( .A(x[479]), .B(y[479]), .Z(n1985) );
  XOR U2361 ( .A(x[475]), .B(y[475]), .Z(n1982) );
  XOR U2362 ( .A(x[477]), .B(y[477]), .Z(n1983) );
  XNOR U2363 ( .A(n1985), .B(n1984), .Z(n1883) );
  XNOR U2364 ( .A(n1884), .B(n1883), .Z(n1885) );
  XOR U2365 ( .A(n1886), .B(n1885), .Z(n2054) );
  XOR U2366 ( .A(n2053), .B(n2054), .Z(n2642) );
  XOR U2367 ( .A(x[485]), .B(y[485]), .Z(n1997) );
  XOR U2368 ( .A(x[481]), .B(y[481]), .Z(n1994) );
  XOR U2369 ( .A(x[483]), .B(y[483]), .Z(n1995) );
  XOR U2370 ( .A(n1997), .B(n1996), .Z(n1922) );
  XOR U2371 ( .A(x[378]), .B(y[378]), .Z(n2698) );
  XOR U2372 ( .A(x[71]), .B(y[71]), .Z(n2695) );
  XOR U2373 ( .A(x[380]), .B(y[380]), .Z(n2696) );
  XOR U2374 ( .A(n2698), .B(n2697), .Z(n1920) );
  XOR U2375 ( .A(x[491]), .B(y[491]), .Z(n1944) );
  XOR U2376 ( .A(x[487]), .B(y[487]), .Z(n1941) );
  XOR U2377 ( .A(x[489]), .B(y[489]), .Z(n1942) );
  XNOR U2378 ( .A(n1944), .B(n1943), .Z(n1919) );
  XNOR U2379 ( .A(n1920), .B(n1919), .Z(n1921) );
  XNOR U2380 ( .A(n1922), .B(n1921), .Z(n2087) );
  XOR U2381 ( .A(x[497]), .B(y[497]), .Z(n1956) );
  XOR U2382 ( .A(x[493]), .B(y[493]), .Z(n1953) );
  XOR U2383 ( .A(x[495]), .B(y[495]), .Z(n1954) );
  XOR U2384 ( .A(n1956), .B(n1955), .Z(n1862) );
  XOR U2385 ( .A(x[942]), .B(y[942]), .Z(n2753) );
  XOR U2386 ( .A(x[35]), .B(y[35]), .Z(n2750) );
  XOR U2387 ( .A(x[944]), .B(y[944]), .Z(n2751) );
  XOR U2388 ( .A(n2753), .B(n2752), .Z(n1860) );
  XOR U2389 ( .A(x[503]), .B(y[503]), .Z(n1916) );
  XOR U2390 ( .A(x[499]), .B(y[499]), .Z(n1913) );
  XOR U2391 ( .A(x[501]), .B(y[501]), .Z(n1914) );
  XNOR U2392 ( .A(n1916), .B(n1915), .Z(n1859) );
  XNOR U2393 ( .A(n1860), .B(n1859), .Z(n1861) );
  XOR U2394 ( .A(n1862), .B(n1861), .Z(n2088) );
  XNOR U2395 ( .A(n2087), .B(n2088), .Z(n2090) );
  XOR U2396 ( .A(x[509]), .B(y[509]), .Z(n1910) );
  XOR U2397 ( .A(x[505]), .B(y[505]), .Z(n1907) );
  XNOR U2398 ( .A(x[507]), .B(y[507]), .Z(n1908) );
  XNOR U2399 ( .A(n1907), .B(n1908), .Z(n1909) );
  XOR U2400 ( .A(n1910), .B(n1909), .Z(n1185) );
  XOR U2401 ( .A(x[366]), .B(y[366]), .Z(n960) );
  XOR U2402 ( .A(x[368]), .B(y[368]), .Z(n957) );
  XNOR U2403 ( .A(x[370]), .B(y[370]), .Z(n958) );
  XNOR U2404 ( .A(n957), .B(n958), .Z(n959) );
  XOR U2405 ( .A(n960), .B(n959), .Z(n1183) );
  XOR U2406 ( .A(x[515]), .B(y[515]), .Z(n1880) );
  XOR U2407 ( .A(x[511]), .B(y[511]), .Z(n1877) );
  XNOR U2408 ( .A(x[513]), .B(y[513]), .Z(n1878) );
  XNOR U2409 ( .A(n1877), .B(n1878), .Z(n1879) );
  XNOR U2410 ( .A(n1880), .B(n1879), .Z(n1182) );
  XNOR U2411 ( .A(n1183), .B(n1182), .Z(n1184) );
  XNOR U2412 ( .A(n1185), .B(n1184), .Z(n2089) );
  XNOR U2413 ( .A(n2090), .B(n2089), .Z(n2641) );
  XOR U2414 ( .A(n2642), .B(n2641), .Z(n2643) );
  XNOR U2415 ( .A(n2644), .B(n2643), .Z(n2872) );
  XOR U2416 ( .A(x[521]), .B(y[521]), .Z(n1874) );
  XOR U2417 ( .A(x[517]), .B(y[517]), .Z(n1871) );
  XNOR U2418 ( .A(x[519]), .B(y[519]), .Z(n1872) );
  XNOR U2419 ( .A(n1871), .B(n1872), .Z(n1873) );
  XOR U2420 ( .A(n1874), .B(n1873), .Z(n290) );
  XOR U2421 ( .A(x[946]), .B(y[946]), .Z(n954) );
  XOR U2422 ( .A(x[212]), .B(y[212]), .Z(n951) );
  XOR U2423 ( .A(x[948]), .B(y[948]), .Z(n952) );
  XOR U2424 ( .A(n954), .B(n953), .Z(n288) );
  XOR U2425 ( .A(x[527]), .B(y[527]), .Z(n284) );
  XOR U2426 ( .A(x[523]), .B(y[523]), .Z(n281) );
  XNOR U2427 ( .A(x[525]), .B(y[525]), .Z(n282) );
  XNOR U2428 ( .A(n281), .B(n282), .Z(n283) );
  XNOR U2429 ( .A(n284), .B(n283), .Z(n287) );
  XNOR U2430 ( .A(n288), .B(n287), .Z(n289) );
  XNOR U2431 ( .A(n290), .B(n289), .Z(n2129) );
  XOR U2432 ( .A(x[188]), .B(y[188]), .Z(n918) );
  XOR U2433 ( .A(x[194]), .B(y[194]), .Z(n915) );
  XNOR U2434 ( .A(x[213]), .B(y[213]), .Z(n916) );
  XNOR U2435 ( .A(n915), .B(n916), .Z(n917) );
  XOR U2436 ( .A(n918), .B(n917), .Z(n1634) );
  XOR U2437 ( .A(x[180]), .B(y[180]), .Z(n1640) );
  XOR U2438 ( .A(x[182]), .B(y[182]), .Z(n1637) );
  XOR U2439 ( .A(x[217]), .B(y[217]), .Z(n1638) );
  XOR U2440 ( .A(n1640), .B(n1639), .Z(n1632) );
  XOR U2441 ( .A(x[837]), .B(y[837]), .Z(n871) );
  XOR U2442 ( .A(x[849]), .B(y[849]), .Z(n868) );
  XNOR U2443 ( .A(x[855]), .B(y[855]), .Z(n869) );
  XNOR U2444 ( .A(n868), .B(n869), .Z(n870) );
  XNOR U2445 ( .A(n871), .B(n870), .Z(n1631) );
  XNOR U2446 ( .A(n1632), .B(n1631), .Z(n1633) );
  XOR U2447 ( .A(n1634), .B(n1633), .Z(n2130) );
  XNOR U2448 ( .A(n2129), .B(n2130), .Z(n2131) );
  XOR U2449 ( .A(x[533]), .B(y[533]), .Z(n278) );
  XOR U2450 ( .A(x[529]), .B(y[529]), .Z(n275) );
  XNOR U2451 ( .A(x[531]), .B(y[531]), .Z(n276) );
  XNOR U2452 ( .A(n275), .B(n276), .Z(n277) );
  XOR U2453 ( .A(n278), .B(n277), .Z(n484) );
  XOR U2454 ( .A(x[358]), .B(y[358]), .Z(n3165) );
  XOR U2455 ( .A(x[93]), .B(y[93]), .Z(n3162) );
  XOR U2456 ( .A(x[360]), .B(y[360]), .Z(n3163) );
  XOR U2457 ( .A(n3165), .B(n3164), .Z(n482) );
  XOR U2458 ( .A(x[539]), .B(y[539]), .Z(n526) );
  XOR U2459 ( .A(x[535]), .B(y[535]), .Z(n523) );
  XOR U2460 ( .A(x[537]), .B(y[537]), .Z(n524) );
  XNOR U2461 ( .A(n526), .B(n525), .Z(n481) );
  XNOR U2462 ( .A(n482), .B(n481), .Z(n483) );
  XOR U2463 ( .A(n484), .B(n483), .Z(n2132) );
  XOR U2464 ( .A(n2131), .B(n2132), .Z(n2776) );
  XOR U2465 ( .A(x[831]), .B(y[831]), .Z(n834) );
  XOR U2466 ( .A(x[829]), .B(y[829]), .Z(n832) );
  XNOR U2467 ( .A(x[857]), .B(y[857]), .Z(n833) );
  XOR U2468 ( .A(n832), .B(n833), .Z(n835) );
  XNOR U2469 ( .A(n834), .B(n835), .Z(n1697) );
  XOR U2470 ( .A(x[998]), .B(y[998]), .Z(n875) );
  XNOR U2471 ( .A(x[254]), .B(y[254]), .Z(n874) );
  XOR U2472 ( .A(oglobal[0]), .B(n874), .Z(n876) );
  XOR U2473 ( .A(n875), .B(n876), .Z(n1698) );
  XNOR U2474 ( .A(n1697), .B(n1698), .Z(n1700) );
  XOR U2475 ( .A(x[851]), .B(y[851]), .Z(n862) );
  XNOR U2476 ( .A(x[853]), .B(y[853]), .Z(n863) );
  XNOR U2477 ( .A(n862), .B(n863), .Z(n864) );
  XOR U2478 ( .A(x[250]), .B(y[250]), .Z(n1646) );
  XOR U2479 ( .A(x[252]), .B(y[252]), .Z(n1643) );
  XOR U2480 ( .A(x[999]), .B(y[999]), .Z(n1644) );
  XOR U2481 ( .A(n1646), .B(n1645), .Z(n865) );
  XOR U2482 ( .A(n864), .B(n865), .Z(n1699) );
  XOR U2483 ( .A(n1700), .B(n1699), .Z(n2094) );
  XOR U2484 ( .A(x[545]), .B(y[545]), .Z(n532) );
  XOR U2485 ( .A(x[541]), .B(y[541]), .Z(n529) );
  XNOR U2486 ( .A(x[543]), .B(y[543]), .Z(n530) );
  XNOR U2487 ( .A(n529), .B(n530), .Z(n531) );
  XOR U2488 ( .A(n532), .B(n531), .Z(n441) );
  XOR U2489 ( .A(x[950]), .B(y[950]), .Z(n2204) );
  XOR U2490 ( .A(x[29]), .B(y[29]), .Z(n2201) );
  XOR U2491 ( .A(x[952]), .B(y[952]), .Z(n2202) );
  XOR U2492 ( .A(n2204), .B(n2203), .Z(n439) );
  XOR U2493 ( .A(x[551]), .B(y[551]), .Z(n2216) );
  XOR U2494 ( .A(x[547]), .B(y[547]), .Z(n2213) );
  XOR U2495 ( .A(x[549]), .B(y[549]), .Z(n2214) );
  XNOR U2496 ( .A(n2216), .B(n2215), .Z(n438) );
  XNOR U2497 ( .A(n439), .B(n438), .Z(n440) );
  XNOR U2498 ( .A(n441), .B(n440), .Z(n2093) );
  XNOR U2499 ( .A(n2094), .B(n2093), .Z(n2095) );
  XOR U2500 ( .A(x[557]), .B(y[557]), .Z(n2210) );
  XOR U2501 ( .A(x[553]), .B(y[553]), .Z(n2207) );
  XOR U2502 ( .A(x[555]), .B(y[555]), .Z(n2208) );
  XOR U2503 ( .A(n2210), .B(n2209), .Z(n1209) );
  XOR U2504 ( .A(x[346]), .B(y[346]), .Z(n966) );
  XOR U2505 ( .A(x[348]), .B(y[348]), .Z(n963) );
  XNOR U2506 ( .A(x[350]), .B(y[350]), .Z(n964) );
  XNOR U2507 ( .A(n963), .B(n964), .Z(n965) );
  XOR U2508 ( .A(n966), .B(n965), .Z(n1207) );
  XOR U2509 ( .A(x[563]), .B(y[563]), .Z(n3219) );
  XOR U2510 ( .A(x[559]), .B(y[559]), .Z(n3216) );
  XOR U2511 ( .A(x[561]), .B(y[561]), .Z(n3217) );
  XNOR U2512 ( .A(n3219), .B(n3218), .Z(n1206) );
  XNOR U2513 ( .A(n1207), .B(n1206), .Z(n1208) );
  XOR U2514 ( .A(n1209), .B(n1208), .Z(n2096) );
  XOR U2515 ( .A(n2095), .B(n2096), .Z(n2775) );
  XOR U2516 ( .A(x[571]), .B(y[571]), .Z(n3213) );
  XOR U2517 ( .A(x[565]), .B(y[565]), .Z(n3210) );
  XOR U2518 ( .A(x[567]), .B(y[567]), .Z(n3211) );
  XOR U2519 ( .A(n3213), .B(n3212), .Z(n2102) );
  XOR U2520 ( .A(x[954]), .B(y[954]), .Z(n2445) );
  XOR U2521 ( .A(x[218]), .B(y[218]), .Z(n2442) );
  XOR U2522 ( .A(x[956]), .B(y[956]), .Z(n2443) );
  XOR U2523 ( .A(n2445), .B(n2444), .Z(n2100) );
  XOR U2524 ( .A(x[583]), .B(y[583]), .Z(n2457) );
  XOR U2525 ( .A(x[575]), .B(y[575]), .Z(n2454) );
  XOR U2526 ( .A(x[579]), .B(y[579]), .Z(n2455) );
  XNOR U2527 ( .A(n2457), .B(n2456), .Z(n2099) );
  XNOR U2528 ( .A(n2100), .B(n2099), .Z(n2101) );
  XNOR U2529 ( .A(n2102), .B(n2101), .Z(n2139) );
  XOR U2530 ( .A(x[825]), .B(y[825]), .Z(n924) );
  XOR U2531 ( .A(x[823]), .B(y[823]), .Z(n921) );
  XNOR U2532 ( .A(x[833]), .B(y[833]), .Z(n922) );
  XNOR U2533 ( .A(n921), .B(n922), .Z(n923) );
  XOR U2534 ( .A(n924), .B(n923), .Z(n1580) );
  XOR U2535 ( .A(x[994]), .B(y[994]), .Z(n829) );
  XOR U2536 ( .A(x[996]), .B(y[996]), .Z(n826) );
  XNOR U2537 ( .A(x[997]), .B(y[997]), .Z(n827) );
  XNOR U2538 ( .A(n826), .B(n827), .Z(n828) );
  XOR U2539 ( .A(n829), .B(n828), .Z(n1578) );
  XOR U2540 ( .A(x[859]), .B(y[859]), .Z(n841) );
  XOR U2541 ( .A(x[827]), .B(y[827]), .Z(n838) );
  XNOR U2542 ( .A(x[861]), .B(y[861]), .Z(n839) );
  XNOR U2543 ( .A(n838), .B(n839), .Z(n840) );
  XNOR U2544 ( .A(n841), .B(n840), .Z(n1577) );
  XNOR U2545 ( .A(n1578), .B(n1577), .Z(n1579) );
  XOR U2546 ( .A(n1580), .B(n1579), .Z(n2140) );
  XNOR U2547 ( .A(n2139), .B(n2140), .Z(n2142) );
  XOR U2548 ( .A(x[595]), .B(y[595]), .Z(n2451) );
  XOR U2549 ( .A(x[587]), .B(y[587]), .Z(n2448) );
  XNOR U2550 ( .A(x[591]), .B(y[591]), .Z(n2449) );
  XNOR U2551 ( .A(n2448), .B(n2449), .Z(n2450) );
  XOR U2552 ( .A(n2451), .B(n2450), .Z(n2154) );
  XOR U2553 ( .A(x[338]), .B(y[338]), .Z(n2759) );
  XOR U2554 ( .A(x[117]), .B(y[117]), .Z(n2756) );
  XOR U2555 ( .A(x[340]), .B(y[340]), .Z(n2757) );
  XOR U2556 ( .A(n2759), .B(n2758), .Z(n2152) );
  XOR U2557 ( .A(x[607]), .B(y[607]), .Z(n2384) );
  XOR U2558 ( .A(x[599]), .B(y[599]), .Z(n2381) );
  XNOR U2559 ( .A(x[603]), .B(y[603]), .Z(n2382) );
  XNOR U2560 ( .A(n2381), .B(n2382), .Z(n2383) );
  XNOR U2561 ( .A(n2384), .B(n2383), .Z(n2151) );
  XNOR U2562 ( .A(n2152), .B(n2151), .Z(n2153) );
  XNOR U2563 ( .A(n2154), .B(n2153), .Z(n2141) );
  XNOR U2564 ( .A(n2142), .B(n2141), .Z(n2774) );
  XOR U2565 ( .A(n2775), .B(n2774), .Z(n2777) );
  XOR U2566 ( .A(n2776), .B(n2777), .Z(n2871) );
  XOR U2567 ( .A(n2872), .B(n2871), .Z(n2874) );
  XOR U2568 ( .A(x[619]), .B(y[619]), .Z(n2378) );
  XOR U2569 ( .A(x[611]), .B(y[611]), .Z(n2375) );
  XNOR U2570 ( .A(x[615]), .B(y[615]), .Z(n2376) );
  XNOR U2571 ( .A(n2375), .B(n2376), .Z(n2377) );
  XOR U2572 ( .A(n2378), .B(n2377), .Z(n2024) );
  XOR U2573 ( .A(x[958]), .B(y[958]), .Z(n2408) );
  XOR U2574 ( .A(x[222]), .B(y[222]), .Z(n2405) );
  XNOR U2575 ( .A(x[960]), .B(y[960]), .Z(n2406) );
  XNOR U2576 ( .A(n2405), .B(n2406), .Z(n2407) );
  XOR U2577 ( .A(n2408), .B(n2407), .Z(n2022) );
  XOR U2578 ( .A(x[631]), .B(y[631]), .Z(n2420) );
  XOR U2579 ( .A(x[623]), .B(y[623]), .Z(n2417) );
  XNOR U2580 ( .A(x[627]), .B(y[627]), .Z(n2418) );
  XNOR U2581 ( .A(n2417), .B(n2418), .Z(n2419) );
  XNOR U2582 ( .A(n2420), .B(n2419), .Z(n2021) );
  XNOR U2583 ( .A(n2022), .B(n2021), .Z(n2023) );
  XNOR U2584 ( .A(n2024), .B(n2023), .Z(n2136) );
  XOR U2585 ( .A(x[821]), .B(y[821]), .Z(n888) );
  XOR U2586 ( .A(x[835]), .B(y[835]), .Z(n885) );
  XNOR U2587 ( .A(x[867]), .B(y[867]), .Z(n886) );
  XNOR U2588 ( .A(n885), .B(n886), .Z(n887) );
  XNOR U2589 ( .A(n888), .B(n887), .Z(n3013) );
  XOR U2590 ( .A(x[198]), .B(y[198]), .Z(n2475) );
  XOR U2591 ( .A(x[202]), .B(y[202]), .Z(n2472) );
  XNOR U2592 ( .A(x[204]), .B(y[204]), .Z(n2473) );
  XNOR U2593 ( .A(n2472), .B(n2473), .Z(n2474) );
  XNOR U2594 ( .A(n2475), .B(n2474), .Z(n3011) );
  XOR U2595 ( .A(x[863]), .B(y[863]), .Z(n930) );
  XOR U2596 ( .A(x[843]), .B(y[843]), .Z(n927) );
  XNOR U2597 ( .A(x[865]), .B(y[865]), .Z(n928) );
  XNOR U2598 ( .A(n927), .B(n928), .Z(n929) );
  XNOR U2599 ( .A(n930), .B(n929), .Z(n3010) );
  XNOR U2600 ( .A(n2136), .B(n2135), .Z(n2137) );
  XOR U2601 ( .A(x[643]), .B(y[643]), .Z(n2414) );
  XOR U2602 ( .A(x[635]), .B(y[635]), .Z(n2411) );
  XOR U2603 ( .A(x[639]), .B(y[639]), .Z(n2412) );
  XOR U2604 ( .A(n2414), .B(n2413), .Z(n1979) );
  XOR U2605 ( .A(x[324]), .B(y[324]), .Z(n2692) );
  XOR U2606 ( .A(x[328]), .B(y[328]), .Z(n2689) );
  XOR U2607 ( .A(x[330]), .B(y[330]), .Z(n2690) );
  XOR U2608 ( .A(n2692), .B(n2691), .Z(n1977) );
  XOR U2609 ( .A(x[655]), .B(y[655]), .Z(n2493) );
  XOR U2610 ( .A(x[647]), .B(y[647]), .Z(n2490) );
  XOR U2611 ( .A(x[651]), .B(y[651]), .Z(n2491) );
  XNOR U2612 ( .A(n2493), .B(n2492), .Z(n1976) );
  XNOR U2613 ( .A(n1977), .B(n1976), .Z(n1978) );
  XOR U2614 ( .A(n1979), .B(n1978), .Z(n2138) );
  XOR U2615 ( .A(n2137), .B(n2138), .Z(n3248) );
  XOR U2616 ( .A(x[667]), .B(y[667]), .Z(n2487) );
  XOR U2617 ( .A(x[659]), .B(y[659]), .Z(n2484) );
  XOR U2618 ( .A(x[663]), .B(y[663]), .Z(n2485) );
  XOR U2619 ( .A(n2487), .B(n2486), .Z(n2084) );
  XOR U2620 ( .A(x[962]), .B(y[962]), .Z(n2295) );
  XOR U2621 ( .A(x[964]), .B(y[964]), .Z(n2292) );
  XOR U2622 ( .A(x[993]), .B(y[993]), .Z(n2293) );
  XOR U2623 ( .A(n2295), .B(n2294), .Z(n2082) );
  XOR U2624 ( .A(x[679]), .B(y[679]), .Z(n2283) );
  XOR U2625 ( .A(x[671]), .B(y[671]), .Z(n2280) );
  XOR U2626 ( .A(x[675]), .B(y[675]), .Z(n2281) );
  XNOR U2627 ( .A(n2283), .B(n2282), .Z(n2081) );
  XNOR U2628 ( .A(n2082), .B(n2081), .Z(n2083) );
  XNOR U2629 ( .A(n2084), .B(n2083), .Z(n2013) );
  XOR U2630 ( .A(x[871]), .B(y[871]), .Z(n942) );
  XOR U2631 ( .A(x[817]), .B(y[817]), .Z(n939) );
  XNOR U2632 ( .A(x[841]), .B(y[841]), .Z(n940) );
  XNOR U2633 ( .A(n939), .B(n940), .Z(n941) );
  XOR U2634 ( .A(n942), .B(n941), .Z(n1538) );
  XOR U2635 ( .A(x[990]), .B(y[990]), .Z(n882) );
  XOR U2636 ( .A(x[244]), .B(y[244]), .Z(n879) );
  XNOR U2637 ( .A(x[992]), .B(y[992]), .Z(n880) );
  XNOR U2638 ( .A(n879), .B(n880), .Z(n881) );
  XOR U2639 ( .A(n882), .B(n881), .Z(n1536) );
  XOR U2640 ( .A(x[819]), .B(y[819]), .Z(n894) );
  XOR U2641 ( .A(x[839]), .B(y[839]), .Z(n891) );
  XNOR U2642 ( .A(x[869]), .B(y[869]), .Z(n892) );
  XNOR U2643 ( .A(n891), .B(n892), .Z(n893) );
  XNOR U2644 ( .A(n894), .B(n893), .Z(n1535) );
  XNOR U2645 ( .A(n1536), .B(n1535), .Z(n1537) );
  XOR U2646 ( .A(n1538), .B(n1537), .Z(n2014) );
  XNOR U2647 ( .A(n2013), .B(n2014), .Z(n2016) );
  XOR U2648 ( .A(x[691]), .B(y[691]), .Z(n2289) );
  XOR U2649 ( .A(x[683]), .B(y[683]), .Z(n2286) );
  XNOR U2650 ( .A(x[687]), .B(y[687]), .Z(n2287) );
  XNOR U2651 ( .A(n2286), .B(n2287), .Z(n2288) );
  XNOR U2652 ( .A(n2289), .B(n2288), .Z(n2048) );
  XOR U2653 ( .A(x[314]), .B(y[314]), .Z(n2511) );
  XOR U2654 ( .A(x[139]), .B(y[139]), .Z(n2508) );
  XNOR U2655 ( .A(x[316]), .B(y[316]), .Z(n2509) );
  XNOR U2656 ( .A(n2508), .B(n2509), .Z(n2510) );
  XNOR U2657 ( .A(n2511), .B(n2510), .Z(n2046) );
  XOR U2658 ( .A(x[701]), .B(y[701]), .Z(n3237) );
  XOR U2659 ( .A(x[695]), .B(y[695]), .Z(n3234) );
  XOR U2660 ( .A(x[699]), .B(y[699]), .Z(n3235) );
  XNOR U2661 ( .A(n3237), .B(n3236), .Z(n2045) );
  XNOR U2662 ( .A(n2016), .B(n2015), .Z(n3247) );
  XOR U2663 ( .A(x[779]), .B(y[779]), .Z(n2246) );
  XOR U2664 ( .A(x[775]), .B(y[775]), .Z(n2243) );
  XOR U2665 ( .A(x[777]), .B(y[777]), .Z(n2244) );
  XNOR U2666 ( .A(n2246), .B(n2245), .Z(n2517) );
  XOR U2667 ( .A(x[978]), .B(y[978]), .Z(n971) );
  XOR U2668 ( .A(x[234]), .B(y[234]), .Z(n969) );
  XNOR U2669 ( .A(x[980]), .B(y[980]), .Z(n970) );
  XOR U2670 ( .A(n969), .B(n970), .Z(n972) );
  XOR U2671 ( .A(n971), .B(n972), .Z(n2515) );
  XOR U2672 ( .A(x[783]), .B(y[783]), .Z(n984) );
  XOR U2673 ( .A(x[781]), .B(y[781]), .Z(n981) );
  XNOR U2674 ( .A(x[897]), .B(y[897]), .Z(n982) );
  XNOR U2675 ( .A(n981), .B(n982), .Z(n983) );
  XNOR U2676 ( .A(n984), .B(n983), .Z(n2514) );
  XOR U2677 ( .A(n2515), .B(n2514), .Z(n2516) );
  XOR U2678 ( .A(x[795]), .B(y[795]), .Z(n2307) );
  XOR U2679 ( .A(x[793]), .B(y[793]), .Z(n2304) );
  XOR U2680 ( .A(x[891]), .B(y[891]), .Z(n2305) );
  XOR U2681 ( .A(n2307), .B(n2306), .Z(n356) );
  XOR U2682 ( .A(x[982]), .B(y[982]), .Z(n2735) );
  XOR U2683 ( .A(x[9]), .B(y[9]), .Z(n2732) );
  XOR U2684 ( .A(x[984]), .B(y[984]), .Z(n2733) );
  XOR U2685 ( .A(n2735), .B(n2734), .Z(n354) );
  XOR U2686 ( .A(x[887]), .B(y[887]), .Z(n2747) );
  XOR U2687 ( .A(x[797]), .B(y[797]), .Z(n2744) );
  XOR U2688 ( .A(x[889]), .B(y[889]), .Z(n2745) );
  XNOR U2689 ( .A(n2747), .B(n2746), .Z(n353) );
  XNOR U2690 ( .A(n354), .B(n353), .Z(n355) );
  XOR U2691 ( .A(n356), .B(n355), .Z(n2008) );
  XNOR U2692 ( .A(n2007), .B(n2008), .Z(n2010) );
  XOR U2693 ( .A(x[787]), .B(y[787]), .Z(n978) );
  XOR U2694 ( .A(x[785]), .B(y[785]), .Z(n975) );
  XOR U2695 ( .A(x[895]), .B(y[895]), .Z(n976) );
  XOR U2696 ( .A(n978), .B(n977), .Z(n405) );
  XOR U2697 ( .A(x[262]), .B(y[262]), .Z(n2402) );
  XOR U2698 ( .A(x[181]), .B(y[181]), .Z(n2399) );
  XOR U2699 ( .A(x[264]), .B(y[264]), .Z(n2400) );
  XOR U2700 ( .A(n2402), .B(n2401), .Z(n403) );
  XOR U2701 ( .A(x[791]), .B(y[791]), .Z(n2313) );
  XOR U2702 ( .A(x[789]), .B(y[789]), .Z(n2310) );
  XOR U2703 ( .A(x[893]), .B(y[893]), .Z(n2311) );
  XNOR U2704 ( .A(n2313), .B(n2312), .Z(n402) );
  XNOR U2705 ( .A(n403), .B(n402), .Z(n404) );
  XNOR U2706 ( .A(n405), .B(n404), .Z(n2009) );
  XNOR U2707 ( .A(n2010), .B(n2009), .Z(n3246) );
  XNOR U2708 ( .A(n3247), .B(n3246), .Z(n3249) );
  XOR U2709 ( .A(n3248), .B(n3249), .Z(n2873) );
  XNOR U2710 ( .A(n2874), .B(n2873), .Z(n239) );
  XNOR U2711 ( .A(n240), .B(n239), .Z(n242) );
  XOR U2712 ( .A(x[707]), .B(y[707]), .Z(n3231) );
  XOR U2713 ( .A(x[703]), .B(y[703]), .Z(n3228) );
  XOR U2714 ( .A(x[705]), .B(y[705]), .Z(n3229) );
  XNOR U2715 ( .A(n3231), .B(n3230), .Z(n2004) );
  XOR U2716 ( .A(x[966]), .B(y[966]), .Z(n3189) );
  XOR U2717 ( .A(x[228]), .B(y[228]), .Z(n3186) );
  XOR U2718 ( .A(x[968]), .B(y[968]), .Z(n3187) );
  XNOR U2719 ( .A(n3189), .B(n3188), .Z(n2002) );
  XOR U2720 ( .A(x[713]), .B(y[713]), .Z(n3201) );
  XOR U2721 ( .A(x[709]), .B(y[709]), .Z(n3198) );
  XOR U2722 ( .A(x[711]), .B(y[711]), .Z(n3199) );
  XNOR U2723 ( .A(n3201), .B(n3200), .Z(n2001) );
  XOR U2724 ( .A(x[805]), .B(y[805]), .Z(n2680) );
  XOR U2725 ( .A(x[847]), .B(y[847]), .Z(n2677) );
  XOR U2726 ( .A(x[875]), .B(y[875]), .Z(n2678) );
  XNOR U2727 ( .A(n2680), .B(n2679), .Z(n2258) );
  XOR U2728 ( .A(x[224]), .B(y[224]), .Z(n2439) );
  XOR U2729 ( .A(x[199]), .B(y[199]), .Z(n2436) );
  XOR U2730 ( .A(x[226]), .B(y[226]), .Z(n2437) );
  XNOR U2731 ( .A(n2439), .B(n2438), .Z(n2256) );
  XOR U2732 ( .A(x[873]), .B(y[873]), .Z(n948) );
  XOR U2733 ( .A(x[815]), .B(y[815]), .Z(n945) );
  XNOR U2734 ( .A(x[845]), .B(y[845]), .Z(n946) );
  XNOR U2735 ( .A(n945), .B(n946), .Z(n947) );
  XNOR U2736 ( .A(n948), .B(n947), .Z(n2255) );
  XNOR U2737 ( .A(n1926), .B(n1925), .Z(n1927) );
  XOR U2738 ( .A(x[719]), .B(y[719]), .Z(n3195) );
  XOR U2739 ( .A(x[715]), .B(y[715]), .Z(n3192) );
  XOR U2740 ( .A(x[717]), .B(y[717]), .Z(n3193) );
  XOR U2741 ( .A(n3195), .B(n3194), .Z(n1963) );
  XOR U2742 ( .A(x[298]), .B(y[298]), .Z(n2319) );
  XOR U2743 ( .A(x[300]), .B(y[300]), .Z(n2316) );
  XOR U2744 ( .A(x[302]), .B(y[302]), .Z(n2317) );
  XNOR U2745 ( .A(n2319), .B(n2318), .Z(n1961) );
  XOR U2746 ( .A(x[725]), .B(y[725]), .Z(n2198) );
  XOR U2747 ( .A(x[721]), .B(y[721]), .Z(n2195) );
  XOR U2748 ( .A(x[723]), .B(y[723]), .Z(n2196) );
  XNOR U2749 ( .A(n2198), .B(n2197), .Z(n1960) );
  XNOR U2750 ( .A(n1963), .B(n1962), .Z(n1928) );
  XNOR U2751 ( .A(n1927), .B(n1928), .Z(n2866) );
  XOR U2752 ( .A(x[755]), .B(y[755]), .Z(n2228) );
  XOR U2753 ( .A(x[751]), .B(y[751]), .Z(n2225) );
  XOR U2754 ( .A(x[753]), .B(y[753]), .Z(n2226) );
  XOR U2755 ( .A(n2228), .B(n2227), .Z(n546) );
  XOR U2756 ( .A(x[974]), .B(y[974]), .Z(n2523) );
  XOR U2757 ( .A(x[15]), .B(y[15]), .Z(n2520) );
  XOR U2758 ( .A(x[976]), .B(y[976]), .Z(n2521) );
  XOR U2759 ( .A(n2523), .B(n2522), .Z(n544) );
  XOR U2760 ( .A(x[761]), .B(y[761]), .Z(n2535) );
  XOR U2761 ( .A(x[757]), .B(y[757]), .Z(n2532) );
  XOR U2762 ( .A(x[759]), .B(y[759]), .Z(n2533) );
  XNOR U2763 ( .A(n2535), .B(n2534), .Z(n543) );
  XNOR U2764 ( .A(n544), .B(n543), .Z(n545) );
  XNOR U2765 ( .A(n546), .B(n545), .Z(n1970) );
  XOR U2766 ( .A(x[801]), .B(y[801]), .Z(n2741) );
  XOR U2767 ( .A(x[799]), .B(y[799]), .Z(n2738) );
  XOR U2768 ( .A(x[811]), .B(y[811]), .Z(n2739) );
  XOR U2769 ( .A(n2741), .B(n2740), .Z(n381) );
  XOR U2770 ( .A(x[236]), .B(y[236]), .Z(n2390) );
  XOR U2771 ( .A(x[238]), .B(y[238]), .Z(n2387) );
  XOR U2772 ( .A(x[246]), .B(y[246]), .Z(n2388) );
  XOR U2773 ( .A(n2390), .B(n2389), .Z(n379) );
  XOR U2774 ( .A(x[883]), .B(y[883]), .Z(n2668) );
  XOR U2775 ( .A(x[813]), .B(y[813]), .Z(n2665) );
  XOR U2776 ( .A(x[885]), .B(y[885]), .Z(n2666) );
  XNOR U2777 ( .A(n2668), .B(n2667), .Z(n378) );
  XNOR U2778 ( .A(n379), .B(n378), .Z(n380) );
  XOR U2779 ( .A(n381), .B(n380), .Z(n1971) );
  XNOR U2780 ( .A(n1970), .B(n1971), .Z(n1972) );
  XOR U2781 ( .A(x[767]), .B(y[767]), .Z(n2529) );
  XOR U2782 ( .A(x[763]), .B(y[763]), .Z(n2526) );
  XOR U2783 ( .A(x[765]), .B(y[765]), .Z(n2527) );
  XOR U2784 ( .A(n2529), .B(n2528), .Z(n570) );
  XOR U2785 ( .A(x[274]), .B(y[274]), .Z(n2331) );
  XOR U2786 ( .A(x[276]), .B(y[276]), .Z(n2328) );
  XOR U2787 ( .A(x[278]), .B(y[278]), .Z(n2329) );
  XOR U2788 ( .A(n2331), .B(n2330), .Z(n568) );
  XOR U2789 ( .A(x[773]), .B(y[773]), .Z(n2252) );
  XOR U2790 ( .A(x[769]), .B(y[769]), .Z(n2249) );
  XOR U2791 ( .A(x[771]), .B(y[771]), .Z(n2250) );
  XNOR U2792 ( .A(n2252), .B(n2251), .Z(n567) );
  XNOR U2793 ( .A(n568), .B(n567), .Z(n569) );
  XOR U2794 ( .A(n570), .B(n569), .Z(n1973) );
  XOR U2795 ( .A(n1972), .B(n1973), .Z(n2864) );
  XOR U2796 ( .A(x[731]), .B(y[731]), .Z(n2192) );
  XOR U2797 ( .A(x[727]), .B(y[727]), .Z(n2189) );
  XOR U2798 ( .A(x[729]), .B(y[729]), .Z(n2190) );
  XOR U2799 ( .A(n2192), .B(n2191), .Z(n1938) );
  XOR U2800 ( .A(x[970]), .B(y[970]), .Z(n2264) );
  XOR U2801 ( .A(x[972]), .B(y[972]), .Z(n2261) );
  XOR U2802 ( .A(x[995]), .B(y[995]), .Z(n2262) );
  XOR U2803 ( .A(n2264), .B(n2263), .Z(n1936) );
  XOR U2804 ( .A(x[737]), .B(y[737]), .Z(n2276) );
  XOR U2805 ( .A(x[733]), .B(y[733]), .Z(n2273) );
  XOR U2806 ( .A(x[735]), .B(y[735]), .Z(n2274) );
  XNOR U2807 ( .A(n2276), .B(n2275), .Z(n1935) );
  XNOR U2808 ( .A(n1936), .B(n1935), .Z(n1937) );
  XNOR U2809 ( .A(n1938), .B(n1937), .Z(n1966) );
  XOR U2810 ( .A(x[881]), .B(y[881]), .Z(n2662) );
  XOR U2811 ( .A(x[803]), .B(y[803]), .Z(n2659) );
  XOR U2812 ( .A(x[807]), .B(y[807]), .Z(n2660) );
  XOR U2813 ( .A(n2662), .B(n2661), .Z(n411) );
  XOR U2814 ( .A(x[986]), .B(y[986]), .Z(n2674) );
  XOR U2815 ( .A(x[240]), .B(y[240]), .Z(n2671) );
  XOR U2816 ( .A(x[988]), .B(y[988]), .Z(n2672) );
  XOR U2817 ( .A(n2674), .B(n2673), .Z(n409) );
  XOR U2818 ( .A(x[877]), .B(y[877]), .Z(n2686) );
  XOR U2819 ( .A(x[809]), .B(y[809]), .Z(n2683) );
  XOR U2820 ( .A(x[879]), .B(y[879]), .Z(n2684) );
  XNOR U2821 ( .A(n2686), .B(n2685), .Z(n408) );
  XNOR U2822 ( .A(n409), .B(n408), .Z(n410) );
  XOR U2823 ( .A(n411), .B(n410), .Z(n1967) );
  XNOR U2824 ( .A(n1966), .B(n1967), .Z(n1969) );
  XOR U2825 ( .A(x[743]), .B(y[743]), .Z(n2270) );
  XOR U2826 ( .A(x[739]), .B(y[739]), .Z(n2267) );
  XOR U2827 ( .A(x[741]), .B(y[741]), .Z(n2268) );
  XNOR U2828 ( .A(n2270), .B(n2269), .Z(n2148) );
  XOR U2829 ( .A(x[288]), .B(y[288]), .Z(n2499) );
  XOR U2830 ( .A(x[161]), .B(y[161]), .Z(n2496) );
  XOR U2831 ( .A(x[292]), .B(y[292]), .Z(n2497) );
  XNOR U2832 ( .A(n2499), .B(n2498), .Z(n2146) );
  XOR U2833 ( .A(x[749]), .B(y[749]), .Z(n2234) );
  XOR U2834 ( .A(x[745]), .B(y[745]), .Z(n2231) );
  XOR U2835 ( .A(x[747]), .B(y[747]), .Z(n2232) );
  XNOR U2836 ( .A(n2234), .B(n2233), .Z(n2145) );
  XNOR U2837 ( .A(n1969), .B(n1968), .Z(n2865) );
  XOR U2838 ( .A(n2864), .B(n2865), .Z(n2867) );
  XOR U2839 ( .A(n2866), .B(n2867), .Z(n2632) );
  XOR U2840 ( .A(x[19]), .B(y[19]), .Z(n2947) );
  XOR U2841 ( .A(x[17]), .B(y[17]), .Z(n2944) );
  XOR U2842 ( .A(x[325]), .B(y[325]), .Z(n2945) );
  XOR U2843 ( .A(n2947), .B(n2946), .Z(n628) );
  XOR U2844 ( .A(x[31]), .B(y[31]), .Z(n2953) );
  XOR U2845 ( .A(x[23]), .B(y[23]), .Z(n2950) );
  XOR U2846 ( .A(x[27]), .B(y[27]), .Z(n2951) );
  XOR U2847 ( .A(n2953), .B(n2952), .Z(n626) );
  XOR U2848 ( .A(x[39]), .B(y[39]), .Z(n1761) );
  XOR U2849 ( .A(x[33]), .B(y[33]), .Z(n1758) );
  XOR U2850 ( .A(x[37]), .B(y[37]), .Z(n1759) );
  XNOR U2851 ( .A(n1761), .B(n1760), .Z(n625) );
  XNOR U2852 ( .A(n626), .B(n625), .Z(n627) );
  XNOR U2853 ( .A(n628), .B(n627), .Z(n1809) );
  XOR U2854 ( .A(x[45]), .B(y[45]), .Z(n1749) );
  XOR U2855 ( .A(x[41]), .B(y[41]), .Z(n1746) );
  XOR U2856 ( .A(x[339]), .B(y[339]), .Z(n1747) );
  XOR U2857 ( .A(n1749), .B(n1748), .Z(n809) );
  XOR U2858 ( .A(x[53]), .B(y[53]), .Z(n1755) );
  XOR U2859 ( .A(x[51]), .B(y[51]), .Z(n1752) );
  XOR U2860 ( .A(x[343]), .B(y[343]), .Z(n1753) );
  XOR U2861 ( .A(n1755), .B(n1754), .Z(n807) );
  XOR U2862 ( .A(x[61]), .B(y[61]), .Z(n1830) );
  XOR U2863 ( .A(x[57]), .B(y[57]), .Z(n1827) );
  XOR U2864 ( .A(x[59]), .B(y[59]), .Z(n1828) );
  XNOR U2865 ( .A(n1830), .B(n1829), .Z(n806) );
  XNOR U2866 ( .A(n807), .B(n806), .Z(n808) );
  XOR U2867 ( .A(n809), .B(n808), .Z(n1810) );
  XNOR U2868 ( .A(n1809), .B(n1810), .Z(n1812) );
  XOR U2869 ( .A(x[73]), .B(y[73]), .Z(n1842) );
  XOR U2870 ( .A(x[63]), .B(y[63]), .Z(n1839) );
  XOR U2871 ( .A(x[67]), .B(y[67]), .Z(n1840) );
  XOR U2872 ( .A(n1842), .B(n1841), .Z(n779) );
  XOR U2873 ( .A(x[79]), .B(y[79]), .Z(n1836) );
  XOR U2874 ( .A(x[77]), .B(y[77]), .Z(n1833) );
  XOR U2875 ( .A(x[357]), .B(y[357]), .Z(n1834) );
  XOR U2876 ( .A(n1836), .B(n1835), .Z(n777) );
  XOR U2877 ( .A(x[83]), .B(y[83]), .Z(n1424) );
  XOR U2878 ( .A(x[81]), .B(y[81]), .Z(n1421) );
  XOR U2879 ( .A(x[361]), .B(y[361]), .Z(n1422) );
  XNOR U2880 ( .A(n1424), .B(n1423), .Z(n776) );
  XNOR U2881 ( .A(n777), .B(n776), .Z(n778) );
  XNOR U2882 ( .A(n779), .B(n778), .Z(n1811) );
  XOR U2883 ( .A(n1812), .B(n1811), .Z(n2638) );
  XOR U2884 ( .A(x[97]), .B(y[97]), .Z(n1412) );
  XOR U2885 ( .A(x[85]), .B(y[85]), .Z(n1409) );
  XNOR U2886 ( .A(x[91]), .B(y[91]), .Z(n1410) );
  XNOR U2887 ( .A(n1409), .B(n1410), .Z(n1411) );
  XOR U2888 ( .A(n1412), .B(n1411), .Z(n785) );
  XOR U2889 ( .A(x[103]), .B(y[103]), .Z(n1418) );
  XOR U2890 ( .A(x[99]), .B(y[99]), .Z(n1415) );
  XNOR U2891 ( .A(x[101]), .B(y[101]), .Z(n1416) );
  XNOR U2892 ( .A(n1415), .B(n1416), .Z(n1417) );
  XOR U2893 ( .A(n1418), .B(n1417), .Z(n783) );
  XOR U2894 ( .A(x[107]), .B(y[107]), .Z(n1306) );
  XOR U2895 ( .A(x[105]), .B(y[105]), .Z(n1303) );
  XOR U2896 ( .A(x[963]), .B(y[963]), .Z(n1304) );
  XNOR U2897 ( .A(n1306), .B(n1305), .Z(n782) );
  XNOR U2898 ( .A(n783), .B(n782), .Z(n784) );
  XNOR U2899 ( .A(n785), .B(n784), .Z(n1853) );
  XOR U2900 ( .A(x[119]), .B(y[119]), .Z(n1312) );
  XOR U2901 ( .A(x[113]), .B(y[113]), .Z(n1309) );
  XOR U2902 ( .A(x[569]), .B(y[569]), .Z(n1310) );
  XOR U2903 ( .A(n1312), .B(n1311), .Z(n658) );
  XOR U2904 ( .A(x[123]), .B(y[123]), .Z(n1318) );
  XOR U2905 ( .A(x[121]), .B(y[121]), .Z(n1315) );
  XOR U2906 ( .A(x[961]), .B(y[961]), .Z(n1316) );
  XOR U2907 ( .A(n1318), .B(n1317), .Z(n656) );
  XOR U2908 ( .A(x[127]), .B(y[127]), .Z(n594) );
  XOR U2909 ( .A(x[125]), .B(y[125]), .Z(n591) );
  XNOR U2910 ( .A(x[573]), .B(y[573]), .Z(n592) );
  XNOR U2911 ( .A(n591), .B(n592), .Z(n593) );
  XNOR U2912 ( .A(n594), .B(n593), .Z(n655) );
  XNOR U2913 ( .A(n656), .B(n655), .Z(n657) );
  XOR U2914 ( .A(n658), .B(n657), .Z(n1854) );
  XNOR U2915 ( .A(n1853), .B(n1854), .Z(n1856) );
  XOR U2916 ( .A(x[137]), .B(y[137]), .Z(n582) );
  XOR U2917 ( .A(x[131]), .B(y[131]), .Z(n579) );
  XNOR U2918 ( .A(x[959]), .B(y[959]), .Z(n580) );
  XNOR U2919 ( .A(n579), .B(n580), .Z(n581) );
  XOR U2920 ( .A(n582), .B(n581), .Z(n664) );
  XOR U2921 ( .A(x[143]), .B(y[143]), .Z(n588) );
  XOR U2922 ( .A(x[141]), .B(y[141]), .Z(n585) );
  XNOR U2923 ( .A(x[577]), .B(y[577]), .Z(n586) );
  XNOR U2924 ( .A(n585), .B(n586), .Z(n587) );
  XOR U2925 ( .A(n588), .B(n587), .Z(n662) );
  XOR U2926 ( .A(x[147]), .B(y[147]), .Z(n622) );
  XOR U2927 ( .A(x[145]), .B(y[145]), .Z(n619) );
  XNOR U2928 ( .A(x[957]), .B(y[957]), .Z(n620) );
  XNOR U2929 ( .A(n619), .B(n620), .Z(n621) );
  XNOR U2930 ( .A(n622), .B(n621), .Z(n661) );
  XNOR U2931 ( .A(n662), .B(n661), .Z(n663) );
  XNOR U2932 ( .A(n664), .B(n663), .Z(n1855) );
  XOR U2933 ( .A(n1856), .B(n1855), .Z(n2636) );
  XOR U2934 ( .A(x[153]), .B(y[153]), .Z(n610) );
  XOR U2935 ( .A(x[151]), .B(y[151]), .Z(n607) );
  XNOR U2936 ( .A(x[581]), .B(y[581]), .Z(n608) );
  XNOR U2937 ( .A(n607), .B(n608), .Z(n609) );
  XNOR U2938 ( .A(n610), .B(n609), .Z(n2594) );
  XOR U2939 ( .A(x[163]), .B(y[163]), .Z(n616) );
  XOR U2940 ( .A(x[159]), .B(y[159]), .Z(n613) );
  XNOR U2941 ( .A(x[955]), .B(y[955]), .Z(n614) );
  XNOR U2942 ( .A(n613), .B(n614), .Z(n615) );
  XNOR U2943 ( .A(n616), .B(n615), .Z(n2592) );
  XOR U2944 ( .A(x[167]), .B(y[167]), .Z(n742) );
  XOR U2945 ( .A(x[165]), .B(y[165]), .Z(n739) );
  XNOR U2946 ( .A(x[585]), .B(y[585]), .Z(n740) );
  XNOR U2947 ( .A(n739), .B(n740), .Z(n741) );
  XNOR U2948 ( .A(n742), .B(n741), .Z(n2591) );
  XOR U2949 ( .A(x[173]), .B(y[173]), .Z(n730) );
  XOR U2950 ( .A(x[171]), .B(y[171]), .Z(n727) );
  XOR U2951 ( .A(x[953]), .B(y[953]), .Z(n728) );
  XOR U2952 ( .A(n730), .B(n729), .Z(n694) );
  XOR U2953 ( .A(x[179]), .B(y[179]), .Z(n736) );
  XOR U2954 ( .A(x[175]), .B(y[175]), .Z(n733) );
  XOR U2955 ( .A(x[589]), .B(y[589]), .Z(n734) );
  XOR U2956 ( .A(n736), .B(n735), .Z(n692) );
  XOR U2957 ( .A(x[185]), .B(y[185]), .Z(n773) );
  XOR U2958 ( .A(x[183]), .B(y[183]), .Z(n770) );
  XOR U2959 ( .A(x[951]), .B(y[951]), .Z(n771) );
  XNOR U2960 ( .A(n773), .B(n772), .Z(n691) );
  XNOR U2961 ( .A(n692), .B(n691), .Z(n693) );
  XOR U2962 ( .A(n694), .B(n693), .Z(n1890) );
  XNOR U2963 ( .A(n1889), .B(n1890), .Z(n1892) );
  XOR U2964 ( .A(x[189]), .B(y[189]), .Z(n761) );
  XOR U2965 ( .A(x[187]), .B(y[187]), .Z(n758) );
  XNOR U2966 ( .A(x[593]), .B(y[593]), .Z(n759) );
  XNOR U2967 ( .A(n758), .B(n759), .Z(n760) );
  XOR U2968 ( .A(n761), .B(n760), .Z(n1737) );
  XOR U2969 ( .A(x[193]), .B(y[193]), .Z(n767) );
  XOR U2970 ( .A(x[191]), .B(y[191]), .Z(n764) );
  XNOR U2971 ( .A(x[949]), .B(y[949]), .Z(n765) );
  XNOR U2972 ( .A(n764), .B(n765), .Z(n766) );
  XOR U2973 ( .A(n767), .B(n766), .Z(n1735) );
  XOR U2974 ( .A(x[201]), .B(y[201]), .Z(n803) );
  XOR U2975 ( .A(x[197]), .B(y[197]), .Z(n800) );
  XNOR U2976 ( .A(x[597]), .B(y[597]), .Z(n801) );
  XNOR U2977 ( .A(n800), .B(n801), .Z(n802) );
  XNOR U2978 ( .A(n803), .B(n802), .Z(n1734) );
  XNOR U2979 ( .A(n1735), .B(n1734), .Z(n1736) );
  XNOR U2980 ( .A(n1737), .B(n1736), .Z(n1891) );
  XNOR U2981 ( .A(n1892), .B(n1891), .Z(n2635) );
  XNOR U2982 ( .A(n2636), .B(n2635), .Z(n2637) );
  XNOR U2983 ( .A(n2638), .B(n2637), .Z(n3121) );
  XOR U2984 ( .A(x[297]), .B(y[297]), .Z(n847) );
  XOR U2985 ( .A(x[295]), .B(y[295]), .Z(n844) );
  XOR U2986 ( .A(x[929]), .B(y[929]), .Z(n845) );
  XOR U2987 ( .A(n847), .B(n846), .Z(n576) );
  XOR U2988 ( .A(x[301]), .B(y[301]), .Z(n853) );
  XOR U2989 ( .A(x[299]), .B(y[299]), .Z(n850) );
  XOR U2990 ( .A(x[637]), .B(y[637]), .Z(n851) );
  XOR U2991 ( .A(n853), .B(n852), .Z(n574) );
  XOR U2992 ( .A(x[309]), .B(y[309]), .Z(n912) );
  XOR U2993 ( .A(x[305]), .B(y[305]), .Z(n909) );
  XOR U2994 ( .A(x[927]), .B(y[927]), .Z(n910) );
  XNOR U2995 ( .A(n912), .B(n911), .Z(n573) );
  XNOR U2996 ( .A(n574), .B(n573), .Z(n575) );
  XNOR U2997 ( .A(n576), .B(n575), .Z(n1096) );
  XOR U2998 ( .A(x[313]), .B(y[313]), .Z(n900) );
  XOR U2999 ( .A(x[311]), .B(y[311]), .Z(n897) );
  XOR U3000 ( .A(x[641]), .B(y[641]), .Z(n898) );
  XOR U3001 ( .A(n900), .B(n899), .Z(n2819) );
  XOR U3002 ( .A(x[317]), .B(y[317]), .Z(n906) );
  XOR U3003 ( .A(x[315]), .B(y[315]), .Z(n903) );
  XOR U3004 ( .A(x[925]), .B(y[925]), .Z(n904) );
  XOR U3005 ( .A(n906), .B(n905), .Z(n2817) );
  XOR U3006 ( .A(x[323]), .B(y[323]), .Z(n564) );
  XOR U3007 ( .A(x[319]), .B(y[319]), .Z(n561) );
  XNOR U3008 ( .A(x[645]), .B(y[645]), .Z(n562) );
  XNOR U3009 ( .A(n561), .B(n562), .Z(n563) );
  XNOR U3010 ( .A(n564), .B(n563), .Z(n2816) );
  XNOR U3011 ( .A(n2817), .B(n2816), .Z(n2818) );
  XNOR U3012 ( .A(n2819), .B(n2818), .Z(n1095) );
  XOR U3013 ( .A(n1096), .B(n1095), .Z(n1098) );
  XOR U3014 ( .A(x[329]), .B(y[329]), .Z(n552) );
  XOR U3015 ( .A(x[327]), .B(y[327]), .Z(n549) );
  XNOR U3016 ( .A(x[923]), .B(y[923]), .Z(n550) );
  XNOR U3017 ( .A(n549), .B(n550), .Z(n551) );
  XOR U3018 ( .A(n552), .B(n551), .Z(n2606) );
  XOR U3019 ( .A(x[333]), .B(y[333]), .Z(n558) );
  XOR U3020 ( .A(x[331]), .B(y[331]), .Z(n555) );
  XNOR U3021 ( .A(x[649]), .B(y[649]), .Z(n556) );
  XNOR U3022 ( .A(n555), .B(n556), .Z(n557) );
  XOR U3023 ( .A(n558), .B(n557), .Z(n2604) );
  XOR U3024 ( .A(x[337]), .B(y[337]), .Z(n399) );
  XOR U3025 ( .A(x[335]), .B(y[335]), .Z(n396) );
  XNOR U3026 ( .A(x[921]), .B(y[921]), .Z(n397) );
  XNOR U3027 ( .A(n396), .B(n397), .Z(n398) );
  XNOR U3028 ( .A(n399), .B(n398), .Z(n2603) );
  XNOR U3029 ( .A(n2604), .B(n2603), .Z(n2605) );
  XNOR U3030 ( .A(n2606), .B(n2605), .Z(n1097) );
  XOR U3031 ( .A(n1098), .B(n1097), .Z(n814) );
  XOR U3032 ( .A(x[251]), .B(y[251]), .Z(n700) );
  XOR U3033 ( .A(x[247]), .B(y[247]), .Z(n697) );
  XNOR U3034 ( .A(x[617]), .B(y[617]), .Z(n698) );
  XNOR U3035 ( .A(n697), .B(n698), .Z(n699) );
  XOR U3036 ( .A(n700), .B(n699), .Z(n2965) );
  XOR U3037 ( .A(x[257]), .B(y[257]), .Z(n706) );
  XOR U3038 ( .A(x[255]), .B(y[255]), .Z(n703) );
  XNOR U3039 ( .A(x[937]), .B(y[937]), .Z(n704) );
  XNOR U3040 ( .A(n703), .B(n704), .Z(n705) );
  XOR U3041 ( .A(n706), .B(n705), .Z(n2963) );
  XOR U3042 ( .A(x[261]), .B(y[261]), .Z(n2813) );
  XOR U3043 ( .A(x[259]), .B(y[259]), .Z(n2810) );
  XOR U3044 ( .A(x[621]), .B(y[621]), .Z(n2811) );
  XNOR U3045 ( .A(n2813), .B(n2812), .Z(n2962) );
  XNOR U3046 ( .A(n2963), .B(n2962), .Z(n2964) );
  XNOR U3047 ( .A(n2965), .B(n2964), .Z(n1133) );
  XOR U3048 ( .A(x[265]), .B(y[265]), .Z(n2801) );
  XOR U3049 ( .A(x[263]), .B(y[263]), .Z(n2798) );
  XOR U3050 ( .A(x[935]), .B(y[935]), .Z(n2799) );
  XOR U3051 ( .A(n2801), .B(n2800), .Z(n2941) );
  XOR U3052 ( .A(x[273]), .B(y[273]), .Z(n2807) );
  XOR U3053 ( .A(x[269]), .B(y[269]), .Z(n2804) );
  XOR U3054 ( .A(x[625]), .B(y[625]), .Z(n2805) );
  XOR U3055 ( .A(n2807), .B(n2806), .Z(n2939) );
  XOR U3056 ( .A(x[277]), .B(y[277]), .Z(n2861) );
  XOR U3057 ( .A(x[275]), .B(y[275]), .Z(n2858) );
  XOR U3058 ( .A(x[933]), .B(y[933]), .Z(n2859) );
  XNOR U3059 ( .A(n2861), .B(n2860), .Z(n2938) );
  XNOR U3060 ( .A(n2939), .B(n2938), .Z(n2940) );
  XNOR U3061 ( .A(n2941), .B(n2940), .Z(n1132) );
  XOR U3062 ( .A(n1133), .B(n1132), .Z(n1135) );
  XOR U3063 ( .A(x[281]), .B(y[281]), .Z(n2849) );
  XOR U3064 ( .A(x[279]), .B(y[279]), .Z(n2846) );
  XOR U3065 ( .A(x[629]), .B(y[629]), .Z(n2847) );
  XOR U3066 ( .A(n2849), .B(n2848), .Z(n1743) );
  XOR U3067 ( .A(x[287]), .B(y[287]), .Z(n2855) );
  XOR U3068 ( .A(x[283]), .B(y[283]), .Z(n2852) );
  XOR U3069 ( .A(x[931]), .B(y[931]), .Z(n2853) );
  XOR U3070 ( .A(n2855), .B(n2854), .Z(n1741) );
  XOR U3071 ( .A(x[293]), .B(y[293]), .Z(n859) );
  XOR U3072 ( .A(x[291]), .B(y[291]), .Z(n856) );
  XOR U3073 ( .A(x[633]), .B(y[633]), .Z(n857) );
  XNOR U3074 ( .A(n859), .B(n858), .Z(n1740) );
  XNOR U3075 ( .A(n1741), .B(n1740), .Z(n1742) );
  XNOR U3076 ( .A(n1743), .B(n1742), .Z(n1134) );
  XOR U3077 ( .A(n1135), .B(n1134), .Z(n815) );
  XOR U3078 ( .A(n814), .B(n815), .Z(n816) );
  XOR U3079 ( .A(x[205]), .B(y[205]), .Z(n791) );
  XOR U3080 ( .A(x[203]), .B(y[203]), .Z(n788) );
  XNOR U3081 ( .A(x[947]), .B(y[947]), .Z(n789) );
  XNOR U3082 ( .A(n788), .B(n789), .Z(n790) );
  XNOR U3083 ( .A(n791), .B(n790), .Z(n1104) );
  XOR U3084 ( .A(x[209]), .B(y[209]), .Z(n797) );
  XOR U3085 ( .A(x[207]), .B(y[207]), .Z(n794) );
  XNOR U3086 ( .A(x[601]), .B(y[601]), .Z(n795) );
  XNOR U3087 ( .A(n794), .B(n795), .Z(n796) );
  XNOR U3088 ( .A(n797), .B(n796), .Z(n1102) );
  XOR U3089 ( .A(x[215]), .B(y[215]), .Z(n652) );
  XOR U3090 ( .A(x[211]), .B(y[211]), .Z(n649) );
  XNOR U3091 ( .A(x[945]), .B(y[945]), .Z(n650) );
  XNOR U3092 ( .A(n649), .B(n650), .Z(n651) );
  XNOR U3093 ( .A(n652), .B(n651), .Z(n1101) );
  XOR U3094 ( .A(x[221]), .B(y[221]), .Z(n640) );
  XOR U3095 ( .A(x[219]), .B(y[219]), .Z(n637) );
  XNOR U3096 ( .A(x[605]), .B(y[605]), .Z(n638) );
  XNOR U3097 ( .A(n637), .B(n638), .Z(n639) );
  XNOR U3098 ( .A(n640), .B(n639), .Z(n2880) );
  XOR U3099 ( .A(x[225]), .B(y[225]), .Z(n646) );
  XOR U3100 ( .A(x[223]), .B(y[223]), .Z(n643) );
  XNOR U3101 ( .A(x[943]), .B(y[943]), .Z(n644) );
  XNOR U3102 ( .A(n643), .B(n644), .Z(n645) );
  XNOR U3103 ( .A(n646), .B(n645), .Z(n2878) );
  XOR U3104 ( .A(x[229]), .B(y[229]), .Z(n682) );
  XOR U3105 ( .A(x[227]), .B(y[227]), .Z(n679) );
  XNOR U3106 ( .A(x[609]), .B(y[609]), .Z(n680) );
  XNOR U3107 ( .A(n679), .B(n680), .Z(n681) );
  XNOR U3108 ( .A(n682), .B(n681), .Z(n2877) );
  XOR U3109 ( .A(n1848), .B(n1847), .Z(n1850) );
  XOR U3110 ( .A(x[237]), .B(y[237]), .Z(n670) );
  XOR U3111 ( .A(x[233]), .B(y[233]), .Z(n667) );
  XNOR U3112 ( .A(x[941]), .B(y[941]), .Z(n668) );
  XNOR U3113 ( .A(n667), .B(n668), .Z(n669) );
  XNOR U3114 ( .A(n670), .B(n669), .Z(n1110) );
  XOR U3115 ( .A(x[241]), .B(y[241]), .Z(n676) );
  XOR U3116 ( .A(x[239]), .B(y[239]), .Z(n673) );
  XNOR U3117 ( .A(x[613]), .B(y[613]), .Z(n674) );
  XNOR U3118 ( .A(n673), .B(n674), .Z(n675) );
  XNOR U3119 ( .A(n676), .B(n675), .Z(n1108) );
  XOR U3120 ( .A(x[245]), .B(y[245]), .Z(n712) );
  XOR U3121 ( .A(x[243]), .B(y[243]), .Z(n709) );
  XNOR U3122 ( .A(x[939]), .B(y[939]), .Z(n710) );
  XNOR U3123 ( .A(n709), .B(n710), .Z(n711) );
  XNOR U3124 ( .A(n712), .B(n711), .Z(n1107) );
  XOR U3125 ( .A(n1850), .B(n1849), .Z(n817) );
  XOR U3126 ( .A(n816), .B(n817), .Z(n3120) );
  XNOR U3127 ( .A(n3121), .B(n3120), .Z(n3123) );
  XOR U3128 ( .A(x[373]), .B(y[373]), .Z(n520) );
  XOR U3129 ( .A(x[371]), .B(y[371]), .Z(n517) );
  XNOR U3130 ( .A(x[665]), .B(y[665]), .Z(n518) );
  XNOR U3131 ( .A(n517), .B(n518), .Z(n519) );
  XOR U3132 ( .A(n520), .B(n519), .Z(n1154) );
  XOR U3133 ( .A(x[438]), .B(y[438]), .Z(n1904) );
  XOR U3134 ( .A(x[3]), .B(y[3]), .Z(n1901) );
  XNOR U3135 ( .A(x[440]), .B(y[440]), .Z(n1902) );
  XNOR U3136 ( .A(n1901), .B(n1902), .Z(n1903) );
  XOR U3137 ( .A(n1904), .B(n1903), .Z(n1152) );
  XOR U3138 ( .A(x[377]), .B(y[377]), .Z(n514) );
  XOR U3139 ( .A(x[375]), .B(y[375]), .Z(n511) );
  XNOR U3140 ( .A(x[913]), .B(y[913]), .Z(n512) );
  XNOR U3141 ( .A(n511), .B(n512), .Z(n513) );
  XNOR U3142 ( .A(n514), .B(n513), .Z(n1151) );
  XNOR U3143 ( .A(n1152), .B(n1151), .Z(n1153) );
  XNOR U3144 ( .A(n1154), .B(n1153), .Z(n1145) );
  XOR U3145 ( .A(x[381]), .B(y[381]), .Z(n266) );
  XOR U3146 ( .A(x[379]), .B(y[379]), .Z(n263) );
  XNOR U3147 ( .A(x[669]), .B(y[669]), .Z(n264) );
  XNOR U3148 ( .A(n263), .B(n264), .Z(n265) );
  XOR U3149 ( .A(n266), .B(n265), .Z(n1178) );
  XOR U3150 ( .A(x[918]), .B(y[918]), .Z(n538) );
  XOR U3151 ( .A(x[49]), .B(y[49]), .Z(n535) );
  XNOR U3152 ( .A(x[920]), .B(y[920]), .Z(n536) );
  XNOR U3153 ( .A(n535), .B(n536), .Z(n537) );
  XOR U3154 ( .A(n538), .B(n537), .Z(n1176) );
  XOR U3155 ( .A(x[385]), .B(y[385]), .Z(n254) );
  XOR U3156 ( .A(x[383]), .B(y[383]), .Z(n251) );
  XNOR U3157 ( .A(x[911]), .B(y[911]), .Z(n252) );
  XNOR U3158 ( .A(n251), .B(n252), .Z(n253) );
  XNOR U3159 ( .A(n254), .B(n253), .Z(n1175) );
  XNOR U3160 ( .A(n1176), .B(n1175), .Z(n1177) );
  XNOR U3161 ( .A(n1178), .B(n1177), .Z(n1144) );
  XOR U3162 ( .A(n1145), .B(n1144), .Z(n1147) );
  XOR U3163 ( .A(x[389]), .B(y[389]), .Z(n260) );
  XOR U3164 ( .A(x[387]), .B(y[387]), .Z(n257) );
  XNOR U3165 ( .A(x[673]), .B(y[673]), .Z(n258) );
  XNOR U3166 ( .A(n257), .B(n258), .Z(n259) );
  XOR U3167 ( .A(n260), .B(n259), .Z(n2886) );
  XOR U3168 ( .A(x[426]), .B(y[426]), .Z(n496) );
  XOR U3169 ( .A(x[428]), .B(y[428]), .Z(n493) );
  XNOR U3170 ( .A(x[430]), .B(y[430]), .Z(n494) );
  XNOR U3171 ( .A(n493), .B(n494), .Z(n495) );
  XOR U3172 ( .A(n496), .B(n495), .Z(n2884) );
  XOR U3173 ( .A(x[393]), .B(y[393]), .Z(n447) );
  XOR U3174 ( .A(x[391]), .B(y[391]), .Z(n444) );
  XNOR U3175 ( .A(x[909]), .B(y[909]), .Z(n445) );
  XNOR U3176 ( .A(n444), .B(n445), .Z(n446) );
  XNOR U3177 ( .A(n447), .B(n446), .Z(n2883) );
  XNOR U3178 ( .A(n2884), .B(n2883), .Z(n2885) );
  XNOR U3179 ( .A(n2886), .B(n2885), .Z(n1146) );
  XOR U3180 ( .A(n1147), .B(n1146), .Z(n820) );
  XOR U3181 ( .A(x[397]), .B(y[397]), .Z(n459) );
  XOR U3182 ( .A(x[395]), .B(y[395]), .Z(n456) );
  XNOR U3183 ( .A(x[677]), .B(y[677]), .Z(n457) );
  XNOR U3184 ( .A(n456), .B(n457), .Z(n458) );
  XNOR U3185 ( .A(n459), .B(n458), .Z(n2571) );
  XOR U3186 ( .A(x[922]), .B(y[922]), .Z(n320) );
  XOR U3187 ( .A(x[196]), .B(y[196]), .Z(n317) );
  XNOR U3188 ( .A(x[924]), .B(y[924]), .Z(n318) );
  XNOR U3189 ( .A(n317), .B(n318), .Z(n319) );
  XNOR U3190 ( .A(n320), .B(n319), .Z(n2569) );
  XOR U3191 ( .A(x[401]), .B(y[401]), .Z(n453) );
  XOR U3192 ( .A(x[399]), .B(y[399]), .Z(n450) );
  XNOR U3193 ( .A(x[907]), .B(y[907]), .Z(n451) );
  XNOR U3194 ( .A(n450), .B(n451), .Z(n452) );
  XNOR U3195 ( .A(n453), .B(n452), .Z(n2568) );
  XOR U3196 ( .A(x[405]), .B(y[405]), .Z(n478) );
  XOR U3197 ( .A(x[403]), .B(y[403]), .Z(n475) );
  XNOR U3198 ( .A(x[681]), .B(y[681]), .Z(n476) );
  XNOR U3199 ( .A(n475), .B(n476), .Z(n477) );
  XNOR U3200 ( .A(n478), .B(n477), .Z(n2577) );
  XOR U3201 ( .A(x[418]), .B(y[418]), .Z(n362) );
  XOR U3202 ( .A(x[25]), .B(y[25]), .Z(n359) );
  XNOR U3203 ( .A(x[420]), .B(y[420]), .Z(n360) );
  XNOR U3204 ( .A(n359), .B(n360), .Z(n361) );
  XNOR U3205 ( .A(n362), .B(n361), .Z(n2575) );
  XOR U3206 ( .A(x[409]), .B(y[409]), .Z(n466) );
  XOR U3207 ( .A(x[407]), .B(y[407]), .Z(n463) );
  XNOR U3208 ( .A(x[905]), .B(y[905]), .Z(n464) );
  XNOR U3209 ( .A(n463), .B(n464), .Z(n465) );
  XNOR U3210 ( .A(n466), .B(n465), .Z(n2574) );
  XOR U3211 ( .A(n1930), .B(n1929), .Z(n1932) );
  XOR U3212 ( .A(x[413]), .B(y[413]), .Z(n472) );
  XOR U3213 ( .A(x[411]), .B(y[411]), .Z(n469) );
  XNOR U3214 ( .A(x[685]), .B(y[685]), .Z(n470) );
  XNOR U3215 ( .A(n469), .B(n470), .Z(n471) );
  XNOR U3216 ( .A(n472), .B(n471), .Z(n2547) );
  XOR U3217 ( .A(x[926]), .B(y[926]), .Z(n374) );
  XOR U3218 ( .A(x[200]), .B(y[200]), .Z(n371) );
  XNOR U3219 ( .A(x[928]), .B(y[928]), .Z(n372) );
  XNOR U3220 ( .A(n371), .B(n372), .Z(n373) );
  XNOR U3221 ( .A(n374), .B(n373), .Z(n2545) );
  XOR U3222 ( .A(x[417]), .B(y[417]), .Z(n429) );
  XOR U3223 ( .A(x[415]), .B(y[415]), .Z(n426) );
  XNOR U3224 ( .A(x[903]), .B(y[903]), .Z(n427) );
  XNOR U3225 ( .A(n426), .B(n427), .Z(n428) );
  XNOR U3226 ( .A(n429), .B(n428), .Z(n2544) );
  XOR U3227 ( .A(n1932), .B(n1931), .Z(n821) );
  XOR U3228 ( .A(n820), .B(n821), .Z(n823) );
  XOR U3229 ( .A(x[345]), .B(y[345]), .Z(n387) );
  XOR U3230 ( .A(x[341]), .B(y[341]), .Z(n384) );
  XNOR U3231 ( .A(x[653]), .B(y[653]), .Z(n385) );
  XNOR U3232 ( .A(n384), .B(n385), .Z(n386) );
  XOR U3233 ( .A(n387), .B(n386), .Z(n2360) );
  XOR U3234 ( .A(x[910]), .B(y[910]), .Z(n1950) );
  XOR U3235 ( .A(x[55]), .B(y[55]), .Z(n1947) );
  XNOR U3236 ( .A(x[912]), .B(y[912]), .Z(n1948) );
  XNOR U3237 ( .A(n1947), .B(n1948), .Z(n1949) );
  XOR U3238 ( .A(n1950), .B(n1949), .Z(n2358) );
  XOR U3239 ( .A(x[349]), .B(y[349]), .Z(n393) );
  XOR U3240 ( .A(x[347]), .B(y[347]), .Z(n390) );
  XNOR U3241 ( .A(x[919]), .B(y[919]), .Z(n391) );
  XNOR U3242 ( .A(n390), .B(n391), .Z(n392) );
  XNOR U3243 ( .A(n393), .B(n392), .Z(n2357) );
  XNOR U3244 ( .A(n2358), .B(n2357), .Z(n2359) );
  XNOR U3245 ( .A(n2360), .B(n2359), .Z(n1139) );
  XOR U3246 ( .A(x[353]), .B(y[353]), .Z(n350) );
  XOR U3247 ( .A(x[351]), .B(y[351]), .Z(n347) );
  XNOR U3248 ( .A(x[657]), .B(y[657]), .Z(n348) );
  XNOR U3249 ( .A(n347), .B(n348), .Z(n349) );
  XOR U3250 ( .A(n350), .B(n349), .Z(n2613) );
  XOR U3251 ( .A(x[446]), .B(y[446]), .Z(n1991) );
  XOR U3252 ( .A(x[448]), .B(y[448]), .Z(n1988) );
  XNOR U3253 ( .A(x[450]), .B(y[450]), .Z(n1989) );
  XNOR U3254 ( .A(n1988), .B(n1989), .Z(n1990) );
  XOR U3255 ( .A(n1991), .B(n1990), .Z(n2611) );
  XOR U3256 ( .A(x[359]), .B(y[359]), .Z(n338) );
  XOR U3257 ( .A(x[355]), .B(y[355]), .Z(n335) );
  XNOR U3258 ( .A(x[917]), .B(y[917]), .Z(n336) );
  XNOR U3259 ( .A(n335), .B(n336), .Z(n337) );
  XNOR U3260 ( .A(n338), .B(n337), .Z(n2610) );
  XNOR U3261 ( .A(n2611), .B(n2610), .Z(n2612) );
  XNOR U3262 ( .A(n2613), .B(n2612), .Z(n1138) );
  XOR U3263 ( .A(n1139), .B(n1138), .Z(n1141) );
  XOR U3264 ( .A(x[365]), .B(y[365]), .Z(n344) );
  XOR U3265 ( .A(x[363]), .B(y[363]), .Z(n341) );
  XNOR U3266 ( .A(x[661]), .B(y[661]), .Z(n342) );
  XNOR U3267 ( .A(n341), .B(n342), .Z(n343) );
  XOR U3268 ( .A(n344), .B(n343), .Z(n2619) );
  XOR U3269 ( .A(x[914]), .B(y[914]), .Z(n1868) );
  XOR U3270 ( .A(x[190]), .B(y[190]), .Z(n1865) );
  XNOR U3271 ( .A(x[916]), .B(y[916]), .Z(n1866) );
  XNOR U3272 ( .A(n1865), .B(n1866), .Z(n1867) );
  XOR U3273 ( .A(n1868), .B(n1867), .Z(n2617) );
  XOR U3274 ( .A(x[369]), .B(y[369]), .Z(n508) );
  XOR U3275 ( .A(x[367]), .B(y[367]), .Z(n505) );
  XNOR U3276 ( .A(x[915]), .B(y[915]), .Z(n506) );
  XNOR U3277 ( .A(n505), .B(n506), .Z(n507) );
  XNOR U3278 ( .A(n508), .B(n507), .Z(n2616) );
  XNOR U3279 ( .A(n2617), .B(n2616), .Z(n2618) );
  XNOR U3280 ( .A(n2619), .B(n2618), .Z(n1140) );
  XOR U3281 ( .A(n1141), .B(n1140), .Z(n822) );
  XOR U3282 ( .A(n823), .B(n822), .Z(n3122) );
  XOR U3283 ( .A(n3123), .B(n3122), .Z(n2631) );
  XOR U3284 ( .A(n2632), .B(n2631), .Z(n2634) );
  XOR U3285 ( .A(x[638]), .B(y[638]), .Z(n1009) );
  XOR U3286 ( .A(x[242]), .B(y[242]), .Z(n1006) );
  XNOR U3287 ( .A(x[640]), .B(y[640]), .Z(n1007) );
  XNOR U3288 ( .A(n1006), .B(n1007), .Z(n1008) );
  XOR U3289 ( .A(n1009), .B(n1008), .Z(n1399) );
  XOR U3290 ( .A(x[632]), .B(y[632]), .Z(n3091) );
  XOR U3291 ( .A(x[634]), .B(y[634]), .Z(n3088) );
  XOR U3292 ( .A(x[636]), .B(y[636]), .Z(n3089) );
  XOR U3293 ( .A(n3091), .B(n3090), .Z(n1397) );
  XOR U3294 ( .A(x[626]), .B(y[626]), .Z(n3079) );
  XOR U3295 ( .A(x[628]), .B(y[628]), .Z(n3076) );
  XOR U3296 ( .A(x[630]), .B(y[630]), .Z(n3077) );
  XNOR U3297 ( .A(n3079), .B(n3078), .Z(n1396) );
  XNOR U3298 ( .A(n1397), .B(n1396), .Z(n1398) );
  XNOR U3299 ( .A(n1399), .B(n1398), .Z(n2786) );
  XOR U3300 ( .A(x[622]), .B(y[622]), .Z(n3085) );
  XOR U3301 ( .A(x[220]), .B(y[220]), .Z(n3082) );
  XOR U3302 ( .A(x[624]), .B(y[624]), .Z(n3083) );
  XOR U3303 ( .A(n3085), .B(n3084), .Z(n1787) );
  XOR U3304 ( .A(x[618]), .B(y[618]), .Z(n1215) );
  XOR U3305 ( .A(x[214]), .B(y[214]), .Z(n1212) );
  XNOR U3306 ( .A(x[620]), .B(y[620]), .Z(n1213) );
  XNOR U3307 ( .A(n1212), .B(n1213), .Z(n1214) );
  XOR U3308 ( .A(n1215), .B(n1214), .Z(n1785) );
  XOR U3309 ( .A(x[612]), .B(y[612]), .Z(n1227) );
  XOR U3310 ( .A(x[614]), .B(y[614]), .Z(n1224) );
  XNOR U3311 ( .A(x[616]), .B(y[616]), .Z(n1225) );
  XNOR U3312 ( .A(n1224), .B(n1225), .Z(n1226) );
  XNOR U3313 ( .A(n1227), .B(n1226), .Z(n1784) );
  XNOR U3314 ( .A(n1785), .B(n1784), .Z(n1786) );
  XNOR U3315 ( .A(n1787), .B(n1786), .Z(n2787) );
  XOR U3316 ( .A(x[606]), .B(y[606]), .Z(n1221) );
  XOR U3317 ( .A(x[608]), .B(y[608]), .Z(n1218) );
  XNOR U3318 ( .A(x[610]), .B(y[610]), .Z(n1219) );
  XNOR U3319 ( .A(n1218), .B(n1219), .Z(n1220) );
  XOR U3320 ( .A(n1221), .B(n1220), .Z(n1436) );
  XOR U3321 ( .A(x[602]), .B(y[602]), .Z(n1086) );
  XOR U3322 ( .A(x[192]), .B(y[192]), .Z(n1083) );
  XNOR U3323 ( .A(x[604]), .B(y[604]), .Z(n1084) );
  XNOR U3324 ( .A(n1083), .B(n1084), .Z(n1085) );
  XOR U3325 ( .A(n1086), .B(n1085), .Z(n1434) );
  XOR U3326 ( .A(x[598]), .B(y[598]), .Z(n1074) );
  XOR U3327 ( .A(x[186]), .B(y[186]), .Z(n1071) );
  XNOR U3328 ( .A(x[600]), .B(y[600]), .Z(n1072) );
  XNOR U3329 ( .A(n1071), .B(n1072), .Z(n1073) );
  XNOR U3330 ( .A(n1074), .B(n1073), .Z(n1433) );
  XNOR U3331 ( .A(n1434), .B(n1433), .Z(n1435) );
  XNOR U3332 ( .A(n1436), .B(n1435), .Z(n2788) );
  XOR U3333 ( .A(n2789), .B(n2788), .Z(n2337) );
  XOR U3334 ( .A(x[592]), .B(y[592]), .Z(n1080) );
  XOR U3335 ( .A(x[594]), .B(y[594]), .Z(n1077) );
  XOR U3336 ( .A(x[596]), .B(y[596]), .Z(n1078) );
  XOR U3337 ( .A(n1080), .B(n1079), .Z(n1460) );
  XOR U3338 ( .A(x[586]), .B(y[586]), .Z(n1724) );
  XOR U3339 ( .A(x[588]), .B(y[588]), .Z(n1721) );
  XOR U3340 ( .A(x[590]), .B(y[590]), .Z(n1722) );
  XOR U3341 ( .A(n1724), .B(n1723), .Z(n1458) );
  XOR U3342 ( .A(x[582]), .B(y[582]), .Z(n1712) );
  XOR U3343 ( .A(x[164]), .B(y[164]), .Z(n1709) );
  XOR U3344 ( .A(x[584]), .B(y[584]), .Z(n1710) );
  XNOR U3345 ( .A(n1712), .B(n1711), .Z(n1457) );
  XNOR U3346 ( .A(n1458), .B(n1457), .Z(n1459) );
  XNOR U3347 ( .A(n1460), .B(n1459), .Z(n293) );
  XOR U3348 ( .A(x[578]), .B(y[578]), .Z(n1718) );
  XOR U3349 ( .A(x[158]), .B(y[158]), .Z(n1715) );
  XOR U3350 ( .A(x[580]), .B(y[580]), .Z(n1716) );
  XOR U3351 ( .A(n1718), .B(n1717), .Z(n2583) );
  XOR U3352 ( .A(x[572]), .B(y[572]), .Z(n1484) );
  XOR U3353 ( .A(x[574]), .B(y[574]), .Z(n1481) );
  XOR U3354 ( .A(x[576]), .B(y[576]), .Z(n1482) );
  XOR U3355 ( .A(n1484), .B(n1483), .Z(n2581) );
  XOR U3356 ( .A(x[566]), .B(y[566]), .Z(n1472) );
  XOR U3357 ( .A(x[568]), .B(y[568]), .Z(n1469) );
  XOR U3358 ( .A(x[570]), .B(y[570]), .Z(n1470) );
  XNOR U3359 ( .A(n1472), .B(n1471), .Z(n2580) );
  XNOR U3360 ( .A(n2581), .B(n2580), .Z(n2582) );
  XNOR U3361 ( .A(n2583), .B(n2582), .Z(n294) );
  XOR U3362 ( .A(n293), .B(n294), .Z(n296) );
  XOR U3363 ( .A(x[562]), .B(y[562]), .Z(n1478) );
  XOR U3364 ( .A(x[136]), .B(y[136]), .Z(n1475) );
  XOR U3365 ( .A(x[564]), .B(y[564]), .Z(n1476) );
  XOR U3366 ( .A(n1478), .B(n1477), .Z(n1331) );
  XOR U3367 ( .A(x[558]), .B(y[558]), .Z(n1246) );
  XOR U3368 ( .A(x[128]), .B(y[128]), .Z(n1243) );
  XOR U3369 ( .A(x[560]), .B(y[560]), .Z(n1244) );
  XOR U3370 ( .A(n1246), .B(n1245), .Z(n1329) );
  XOR U3371 ( .A(x[552]), .B(y[552]), .Z(n1234) );
  XOR U3372 ( .A(x[554]), .B(y[554]), .Z(n1231) );
  XOR U3373 ( .A(x[556]), .B(y[556]), .Z(n1232) );
  XNOR U3374 ( .A(n1234), .B(n1233), .Z(n1328) );
  XNOR U3375 ( .A(n1329), .B(n1328), .Z(n1330) );
  XNOR U3376 ( .A(n1331), .B(n1330), .Z(n295) );
  XOR U3377 ( .A(n296), .B(n295), .Z(n2336) );
  XOR U3378 ( .A(x[546]), .B(y[546]), .Z(n1240) );
  XOR U3379 ( .A(x[548]), .B(y[548]), .Z(n1237) );
  XNOR U3380 ( .A(x[550]), .B(y[550]), .Z(n1238) );
  XNOR U3381 ( .A(n1237), .B(n1238), .Z(n1239) );
  XOR U3382 ( .A(n1240), .B(n1239), .Z(n2541) );
  XOR U3383 ( .A(x[542]), .B(y[542]), .Z(n1781) );
  XOR U3384 ( .A(x[106]), .B(y[106]), .Z(n1778) );
  XNOR U3385 ( .A(x[544]), .B(y[544]), .Z(n1779) );
  XNOR U3386 ( .A(n1778), .B(n1779), .Z(n1780) );
  XOR U3387 ( .A(n1781), .B(n1780), .Z(n2539) );
  XOR U3388 ( .A(x[538]), .B(y[538]), .Z(n1769) );
  XOR U3389 ( .A(x[100]), .B(y[100]), .Z(n1766) );
  XNOR U3390 ( .A(x[540]), .B(y[540]), .Z(n1767) );
  XNOR U3391 ( .A(n1766), .B(n1767), .Z(n1768) );
  XNOR U3392 ( .A(n1769), .B(n1768), .Z(n2538) );
  XNOR U3393 ( .A(n2539), .B(n2538), .Z(n2540) );
  XNOR U3394 ( .A(n2541), .B(n2540), .Z(n3127) );
  XOR U3395 ( .A(x[532]), .B(y[532]), .Z(n1775) );
  XOR U3396 ( .A(x[534]), .B(y[534]), .Z(n1772) );
  XNOR U3397 ( .A(x[536]), .B(y[536]), .Z(n1773) );
  XNOR U3398 ( .A(n1772), .B(n1773), .Z(n1774) );
  XOR U3399 ( .A(n1775), .B(n1774), .Z(n2565) );
  XOR U3400 ( .A(x[526]), .B(y[526]), .Z(n1393) );
  XOR U3401 ( .A(x[528]), .B(y[528]), .Z(n1390) );
  XNOR U3402 ( .A(x[530]), .B(y[530]), .Z(n1391) );
  XNOR U3403 ( .A(n1390), .B(n1391), .Z(n1392) );
  XOR U3404 ( .A(n1393), .B(n1392), .Z(n2563) );
  XOR U3405 ( .A(x[522]), .B(y[522]), .Z(n1381) );
  XOR U3406 ( .A(x[78]), .B(y[78]), .Z(n1378) );
  XNOR U3407 ( .A(x[524]), .B(y[524]), .Z(n1379) );
  XNOR U3408 ( .A(n1378), .B(n1379), .Z(n1380) );
  XNOR U3409 ( .A(n1381), .B(n1380), .Z(n2562) );
  XNOR U3410 ( .A(n2563), .B(n2562), .Z(n2564) );
  XNOR U3411 ( .A(n2565), .B(n2564), .Z(n3126) );
  XOR U3412 ( .A(n3127), .B(n3126), .Z(n3129) );
  XOR U3413 ( .A(x[518]), .B(y[518]), .Z(n1387) );
  XOR U3414 ( .A(x[72]), .B(y[72]), .Z(n1384) );
  XNOR U3415 ( .A(x[520]), .B(y[520]), .Z(n1385) );
  XNOR U3416 ( .A(n1384), .B(n1385), .Z(n1386) );
  XOR U3417 ( .A(n1387), .B(n1386), .Z(n2553) );
  XOR U3418 ( .A(x[512]), .B(y[512]), .Z(n1805) );
  XOR U3419 ( .A(x[514]), .B(y[514]), .Z(n1802) );
  XNOR U3420 ( .A(x[516]), .B(y[516]), .Z(n1803) );
  XNOR U3421 ( .A(n1802), .B(n1803), .Z(n1804) );
  XOR U3422 ( .A(n1805), .B(n1804), .Z(n2551) );
  XOR U3423 ( .A(x[506]), .B(y[506]), .Z(n1793) );
  XOR U3424 ( .A(x[508]), .B(y[508]), .Z(n1790) );
  XNOR U3425 ( .A(x[510]), .B(y[510]), .Z(n1791) );
  XNOR U3426 ( .A(n1790), .B(n1791), .Z(n1792) );
  XNOR U3427 ( .A(n1793), .B(n1792), .Z(n2550) );
  XNOR U3428 ( .A(n2551), .B(n2550), .Z(n2552) );
  XNOR U3429 ( .A(n2553), .B(n2552), .Z(n3128) );
  XNOR U3430 ( .A(n3129), .B(n3128), .Z(n2335) );
  XOR U3431 ( .A(n2336), .B(n2335), .Z(n2338) );
  XOR U3432 ( .A(n2337), .B(n2338), .Z(n3117) );
  XOR U3433 ( .A(x[718]), .B(y[718]), .Z(n1526) );
  XOR U3434 ( .A(x[322]), .B(y[322]), .Z(n1523) );
  XNOR U3435 ( .A(x[720]), .B(y[720]), .Z(n1524) );
  XNOR U3436 ( .A(n1523), .B(n1524), .Z(n1525) );
  XOR U3437 ( .A(n1526), .B(n1525), .Z(n1068) );
  XOR U3438 ( .A(x[902]), .B(y[902]), .Z(n2072) );
  XOR U3439 ( .A(x[184]), .B(y[184]), .Z(n2069) );
  XNOR U3440 ( .A(x[904]), .B(y[904]), .Z(n2070) );
  XNOR U3441 ( .A(n2069), .B(n2070), .Z(n2071) );
  XOR U3442 ( .A(n2072), .B(n2071), .Z(n1066) );
  XOR U3443 ( .A(x[712]), .B(y[712]), .Z(n1514) );
  XOR U3444 ( .A(x[714]), .B(y[714]), .Z(n1511) );
  XNOR U3445 ( .A(x[716]), .B(y[716]), .Z(n1512) );
  XNOR U3446 ( .A(n1511), .B(n1512), .Z(n1513) );
  XNOR U3447 ( .A(n1514), .B(n1513), .Z(n1065) );
  XNOR U3448 ( .A(n1066), .B(n1065), .Z(n1067) );
  XNOR U3449 ( .A(n1068), .B(n1067), .Z(n2708) );
  XOR U3450 ( .A(x[706]), .B(y[706]), .Z(n1508) );
  XOR U3451 ( .A(x[708]), .B(y[708]), .Z(n1505) );
  XNOR U3452 ( .A(x[710]), .B(y[710]), .Z(n1506) );
  XNOR U3453 ( .A(n1505), .B(n1506), .Z(n1507) );
  XOR U3454 ( .A(n1508), .B(n1507), .Z(n1092) );
  XOR U3455 ( .A(x[906]), .B(y[906]), .Z(n2166) );
  XOR U3456 ( .A(x[908]), .B(y[908]), .Z(n2163) );
  XNOR U3457 ( .A(x[987]), .B(y[987]), .Z(n2164) );
  XNOR U3458 ( .A(n2163), .B(n2164), .Z(n2165) );
  XOR U3459 ( .A(n2166), .B(n2165), .Z(n1090) );
  XOR U3460 ( .A(x[702]), .B(y[702]), .Z(n1034) );
  XOR U3461 ( .A(x[308]), .B(y[308]), .Z(n1031) );
  XNOR U3462 ( .A(x[704]), .B(y[704]), .Z(n1032) );
  XNOR U3463 ( .A(n1031), .B(n1032), .Z(n1033) );
  XNOR U3464 ( .A(n1034), .B(n1033), .Z(n1089) );
  XNOR U3465 ( .A(n1090), .B(n1089), .Z(n1091) );
  XOR U3466 ( .A(n1092), .B(n1091), .Z(n2709) );
  XNOR U3467 ( .A(n2708), .B(n2709), .Z(n2711) );
  XOR U3468 ( .A(x[698]), .B(y[698]), .Z(n1028) );
  XOR U3469 ( .A(x[304]), .B(y[304]), .Z(n1025) );
  XNOR U3470 ( .A(x[700]), .B(y[700]), .Z(n1026) );
  XNOR U3471 ( .A(n1025), .B(n1026), .Z(n1027) );
  XOR U3472 ( .A(n1028), .B(n1027), .Z(n1730) );
  XOR U3473 ( .A(x[692]), .B(y[692]), .Z(n2929) );
  XOR U3474 ( .A(x[694]), .B(y[694]), .Z(n2926) );
  XNOR U3475 ( .A(x[696]), .B(y[696]), .Z(n2927) );
  XNOR U3476 ( .A(n2926), .B(n2927), .Z(n2928) );
  XOR U3477 ( .A(n2929), .B(n2928), .Z(n1728) );
  XOR U3478 ( .A(x[686]), .B(y[686]), .Z(n2433) );
  XOR U3479 ( .A(x[688]), .B(y[688]), .Z(n2430) );
  XNOR U3480 ( .A(x[690]), .B(y[690]), .Z(n2431) );
  XNOR U3481 ( .A(n2430), .B(n2431), .Z(n2432) );
  XNOR U3482 ( .A(n2433), .B(n2432), .Z(n1727) );
  XNOR U3483 ( .A(n1728), .B(n1727), .Z(n1729) );
  XNOR U3484 ( .A(n1730), .B(n1729), .Z(n2710) );
  XOR U3485 ( .A(n2711), .B(n2710), .Z(n2179) );
  XOR U3486 ( .A(x[814]), .B(y[814]), .Z(n1652) );
  XOR U3487 ( .A(x[115]), .B(y[115]), .Z(n1649) );
  XNOR U3488 ( .A(x[816]), .B(y[816]), .Z(n1650) );
  XNOR U3489 ( .A(n1649), .B(n1650), .Z(n1651) );
  XOR U3490 ( .A(n1652), .B(n1651), .Z(n1294) );
  XOR U3491 ( .A(x[850]), .B(y[850]), .Z(n1288) );
  XOR U3492 ( .A(x[146]), .B(y[146]), .Z(n1285) );
  XNOR U3493 ( .A(x[852]), .B(y[852]), .Z(n1286) );
  XNOR U3494 ( .A(n1285), .B(n1286), .Z(n1287) );
  XOR U3495 ( .A(n1288), .B(n1287), .Z(n1292) );
  XOR U3496 ( .A(x[846]), .B(y[846]), .Z(n1550) );
  XOR U3497 ( .A(x[95]), .B(y[95]), .Z(n1547) );
  XNOR U3498 ( .A(x[848]), .B(y[848]), .Z(n1548) );
  XNOR U3499 ( .A(n1547), .B(n1548), .Z(n1549) );
  XNOR U3500 ( .A(n1550), .B(n1549), .Z(n1291) );
  XNOR U3501 ( .A(n1292), .B(n1291), .Z(n1293) );
  XNOR U3502 ( .A(n1294), .B(n1293), .Z(n2969) );
  XOR U3503 ( .A(x[822]), .B(y[822]), .Z(n1694) );
  XOR U3504 ( .A(x[109]), .B(y[109]), .Z(n1691) );
  XNOR U3505 ( .A(x[824]), .B(y[824]), .Z(n1692) );
  XNOR U3506 ( .A(n1691), .B(n1692), .Z(n1693) );
  XOR U3507 ( .A(n1694), .B(n1693), .Z(n2795) );
  XOR U3508 ( .A(x[818]), .B(y[818]), .Z(n1616) );
  XOR U3509 ( .A(x[124]), .B(y[124]), .Z(n1613) );
  XNOR U3510 ( .A(x[820]), .B(y[820]), .Z(n1614) );
  XNOR U3511 ( .A(n1613), .B(n1614), .Z(n1615) );
  XOR U3512 ( .A(n1616), .B(n1615), .Z(n2793) );
  XOR U3513 ( .A(x[842]), .B(y[842]), .Z(n1556) );
  XOR U3514 ( .A(x[844]), .B(y[844]), .Z(n1553) );
  XNOR U3515 ( .A(x[979]), .B(y[979]), .Z(n1554) );
  XNOR U3516 ( .A(n1553), .B(n1554), .Z(n1555) );
  XNOR U3517 ( .A(n1556), .B(n1555), .Z(n2792) );
  XNOR U3518 ( .A(n2793), .B(n2792), .Z(n2794) );
  XNOR U3519 ( .A(n2795), .B(n2794), .Z(n2968) );
  XOR U3520 ( .A(n2969), .B(n2968), .Z(n2971) );
  XOR U3521 ( .A(x[810]), .B(y[810]), .Z(n1658) );
  XOR U3522 ( .A(x[812]), .B(y[812]), .Z(n1655) );
  XNOR U3523 ( .A(x[975]), .B(y[975]), .Z(n1656) );
  XNOR U3524 ( .A(n1655), .B(n1656), .Z(n1657) );
  XOR U3525 ( .A(n1658), .B(n1657), .Z(n2771) );
  XOR U3526 ( .A(x[834]), .B(y[834]), .Z(n3025) );
  XOR U3527 ( .A(x[836]), .B(y[836]), .Z(n3022) );
  XNOR U3528 ( .A(x[977]), .B(y[977]), .Z(n3023) );
  XNOR U3529 ( .A(n3022), .B(n3023), .Z(n3024) );
  XOR U3530 ( .A(n3025), .B(n3024), .Z(n2769) );
  XOR U3531 ( .A(x[854]), .B(y[854]), .Z(n1258) );
  XOR U3532 ( .A(x[89]), .B(y[89]), .Z(n1255) );
  XNOR U3533 ( .A(x[856]), .B(y[856]), .Z(n1256) );
  XNOR U3534 ( .A(n1255), .B(n1256), .Z(n1257) );
  XNOR U3535 ( .A(n1258), .B(n1257), .Z(n2768) );
  XNOR U3536 ( .A(n2769), .B(n2768), .Z(n2770) );
  XNOR U3537 ( .A(n2771), .B(n2770), .Z(n2970) );
  XOR U3538 ( .A(n2971), .B(n2970), .Z(n2178) );
  XOR U3539 ( .A(x[682]), .B(y[682]), .Z(n2923) );
  XOR U3540 ( .A(x[290]), .B(y[290]), .Z(n2920) );
  XNOR U3541 ( .A(x[684]), .B(y[684]), .Z(n2921) );
  XNOR U3542 ( .A(n2920), .B(n2921), .Z(n2922) );
  XOR U3543 ( .A(n2923), .B(n2922), .Z(n1490) );
  XOR U3544 ( .A(x[678]), .B(y[678]), .Z(n1052) );
  XOR U3545 ( .A(x[286]), .B(y[286]), .Z(n1049) );
  XNOR U3546 ( .A(x[680]), .B(y[680]), .Z(n1050) );
  XNOR U3547 ( .A(n1049), .B(n1050), .Z(n1051) );
  XOR U3548 ( .A(n1052), .B(n1051), .Z(n1488) );
  XOR U3549 ( .A(x[672]), .B(y[672]), .Z(n1040) );
  XOR U3550 ( .A(x[674]), .B(y[674]), .Z(n1037) );
  XNOR U3551 ( .A(x[676]), .B(y[676]), .Z(n1038) );
  XNOR U3552 ( .A(n1037), .B(n1038), .Z(n1039) );
  XNOR U3553 ( .A(n1040), .B(n1039), .Z(n1487) );
  XNOR U3554 ( .A(n1488), .B(n1487), .Z(n1489) );
  XNOR U3555 ( .A(n1490), .B(n1489), .Z(n2647) );
  XOR U3556 ( .A(x[666]), .B(y[666]), .Z(n1046) );
  XOR U3557 ( .A(x[668]), .B(y[668]), .Z(n1043) );
  XNOR U3558 ( .A(x[670]), .B(y[670]), .Z(n1044) );
  XNOR U3559 ( .A(n1043), .B(n1044), .Z(n1045) );
  XOR U3560 ( .A(n1046), .B(n1045), .Z(n1252) );
  XOR U3561 ( .A(x[662]), .B(y[662]), .Z(n3073) );
  XOR U3562 ( .A(x[272]), .B(y[272]), .Z(n3070) );
  XNOR U3563 ( .A(x[664]), .B(y[664]), .Z(n3071) );
  XNOR U3564 ( .A(n3070), .B(n3071), .Z(n3072) );
  XOR U3565 ( .A(n3073), .B(n3072), .Z(n1250) );
  XOR U3566 ( .A(x[658]), .B(y[658]), .Z(n3061) );
  XOR U3567 ( .A(x[268]), .B(y[268]), .Z(n3058) );
  XNOR U3568 ( .A(x[660]), .B(y[660]), .Z(n3059) );
  XNOR U3569 ( .A(n3058), .B(n3059), .Z(n3060) );
  XNOR U3570 ( .A(n3061), .B(n3060), .Z(n1249) );
  XNOR U3571 ( .A(n1250), .B(n1249), .Z(n1251) );
  XOR U3572 ( .A(n1252), .B(n1251), .Z(n2648) );
  XNOR U3573 ( .A(n2647), .B(n2648), .Z(n2650) );
  XOR U3574 ( .A(x[652]), .B(y[652]), .Z(n3067) );
  XOR U3575 ( .A(x[654]), .B(y[654]), .Z(n3064) );
  XOR U3576 ( .A(x[656]), .B(y[656]), .Z(n3065) );
  XOR U3577 ( .A(n3067), .B(n3066), .Z(n1375) );
  XOR U3578 ( .A(x[646]), .B(y[646]), .Z(n997) );
  XOR U3579 ( .A(x[648]), .B(y[648]), .Z(n994) );
  XNOR U3580 ( .A(x[650]), .B(y[650]), .Z(n995) );
  XNOR U3581 ( .A(n994), .B(n995), .Z(n996) );
  XOR U3582 ( .A(n997), .B(n996), .Z(n1373) );
  XOR U3583 ( .A(x[642]), .B(y[642]), .Z(n1003) );
  XOR U3584 ( .A(x[248]), .B(y[248]), .Z(n1000) );
  XNOR U3585 ( .A(x[644]), .B(y[644]), .Z(n1001) );
  XNOR U3586 ( .A(n1000), .B(n1001), .Z(n1002) );
  XNOR U3587 ( .A(n1003), .B(n1002), .Z(n1372) );
  XNOR U3588 ( .A(n1373), .B(n1372), .Z(n1374) );
  XNOR U3589 ( .A(n1375), .B(n1374), .Z(n2649) );
  XNOR U3590 ( .A(n2650), .B(n2649), .Z(n2177) );
  XOR U3591 ( .A(n2178), .B(n2177), .Z(n2180) );
  XOR U3592 ( .A(n2179), .B(n2180), .Z(n3115) );
  XOR U3593 ( .A(x[790]), .B(y[790]), .Z(n1622) );
  XOR U3594 ( .A(x[129]), .B(y[129]), .Z(n1619) );
  XOR U3595 ( .A(x[792]), .B(y[792]), .Z(n1620) );
  XOR U3596 ( .A(n1622), .B(n1621), .Z(n1466) );
  XOR U3597 ( .A(x[866]), .B(y[866]), .Z(n1592) );
  XOR U3598 ( .A(x[868]), .B(y[868]), .Z(n1589) );
  XOR U3599 ( .A(x[981]), .B(y[981]), .Z(n1590) );
  XOR U3600 ( .A(n1592), .B(n1591), .Z(n1464) );
  XOR U3601 ( .A(x[786]), .B(y[786]), .Z(n1276) );
  XOR U3602 ( .A(x[102]), .B(y[102]), .Z(n1273) );
  XNOR U3603 ( .A(x[788]), .B(y[788]), .Z(n1274) );
  XNOR U3604 ( .A(n1273), .B(n1274), .Z(n1275) );
  XNOR U3605 ( .A(n1276), .B(n1275), .Z(n1463) );
  XNOR U3606 ( .A(n1464), .B(n1463), .Z(n1465) );
  XNOR U3607 ( .A(n1466), .B(n1465), .Z(n2341) );
  XOR U3608 ( .A(x[782]), .B(y[782]), .Z(n2995) );
  XOR U3609 ( .A(x[135]), .B(y[135]), .Z(n2992) );
  XOR U3610 ( .A(x[784]), .B(y[784]), .Z(n2993) );
  XOR U3611 ( .A(n2995), .B(n2994), .Z(n1586) );
  XOR U3612 ( .A(x[870]), .B(y[870]), .Z(n1598) );
  XOR U3613 ( .A(x[162]), .B(y[162]), .Z(n1595) );
  XOR U3614 ( .A(x[872]), .B(y[872]), .Z(n1596) );
  XOR U3615 ( .A(n1598), .B(n1597), .Z(n1584) );
  XOR U3616 ( .A(x[778]), .B(y[778]), .Z(n1688) );
  XOR U3617 ( .A(x[780]), .B(y[780]), .Z(n1685) );
  XOR U3618 ( .A(x[971]), .B(y[971]), .Z(n1686) );
  XNOR U3619 ( .A(n1688), .B(n1687), .Z(n1583) );
  XNOR U3620 ( .A(n1584), .B(n1583), .Z(n1585) );
  XOR U3621 ( .A(n1586), .B(n1585), .Z(n2342) );
  XNOR U3622 ( .A(n2341), .B(n2342), .Z(n2344) );
  XOR U3623 ( .A(x[774]), .B(y[774]), .Z(n1544) );
  XOR U3624 ( .A(x[96]), .B(y[96]), .Z(n1541) );
  XNOR U3625 ( .A(x[776]), .B(y[776]), .Z(n1542) );
  XNOR U3626 ( .A(n1541), .B(n1542), .Z(n1543) );
  XNOR U3627 ( .A(n1544), .B(n1543), .Z(n2911) );
  XOR U3628 ( .A(x[874]), .B(y[874]), .Z(n1604) );
  XOR U3629 ( .A(x[876]), .B(y[876]), .Z(n1601) );
  XNOR U3630 ( .A(x[983]), .B(y[983]), .Z(n1602) );
  XNOR U3631 ( .A(n1601), .B(n1602), .Z(n1603) );
  XNOR U3632 ( .A(n1604), .B(n1603), .Z(n2909) );
  XOR U3633 ( .A(x[770]), .B(y[770]), .Z(n1676) );
  XOR U3634 ( .A(x[772]), .B(y[772]), .Z(n1673) );
  XNOR U3635 ( .A(x[969]), .B(y[969]), .Z(n1674) );
  XNOR U3636 ( .A(n1673), .B(n1674), .Z(n1675) );
  XNOR U3637 ( .A(n1676), .B(n1675), .Z(n2908) );
  XNOR U3638 ( .A(n2344), .B(n2343), .Z(n3114) );
  XNOR U3639 ( .A(n3115), .B(n3114), .Z(n3116) );
  XOR U3640 ( .A(n3117), .B(n3116), .Z(n2633) );
  XNOR U3641 ( .A(n2634), .B(n2633), .Z(n241) );
  XNOR U3642 ( .A(n242), .B(n241), .Z(o[0]) );
  NANDN U3643 ( .A(n240), .B(n239), .Z(n244) );
  NAND U3644 ( .A(n242), .B(n241), .Z(n243) );
  AND U3645 ( .A(n244), .B(n243), .Z(n3482) );
  NAND U3646 ( .A(n246), .B(n245), .Z(n250) );
  NAND U3647 ( .A(n248), .B(n247), .Z(n249) );
  NAND U3648 ( .A(n250), .B(n249), .Z(n3665) );
  NANDN U3649 ( .A(n252), .B(n251), .Z(n256) );
  NAND U3650 ( .A(n254), .B(n253), .Z(n255) );
  AND U3651 ( .A(n256), .B(n255), .Z(n4072) );
  NANDN U3652 ( .A(n258), .B(n257), .Z(n262) );
  NAND U3653 ( .A(n260), .B(n259), .Z(n261) );
  AND U3654 ( .A(n262), .B(n261), .Z(n4073) );
  NANDN U3655 ( .A(n264), .B(n263), .Z(n268) );
  NAND U3656 ( .A(n266), .B(n265), .Z(n267) );
  AND U3657 ( .A(n268), .B(n267), .Z(n4074) );
  XOR U3658 ( .A(n4075), .B(n4074), .Z(n4497) );
  NANDN U3659 ( .A(n270), .B(n269), .Z(n274) );
  NAND U3660 ( .A(n272), .B(n271), .Z(n273) );
  AND U3661 ( .A(n274), .B(n273), .Z(n3283) );
  NANDN U3662 ( .A(n276), .B(n275), .Z(n280) );
  NAND U3663 ( .A(n278), .B(n277), .Z(n279) );
  AND U3664 ( .A(n280), .B(n279), .Z(n3284) );
  NANDN U3665 ( .A(n282), .B(n281), .Z(n286) );
  NAND U3666 ( .A(n284), .B(n283), .Z(n285) );
  AND U3667 ( .A(n286), .B(n285), .Z(n3285) );
  XOR U3668 ( .A(n3286), .B(n3285), .Z(n4495) );
  NANDN U3669 ( .A(n288), .B(n287), .Z(n292) );
  NANDN U3670 ( .A(n290), .B(n289), .Z(n291) );
  AND U3671 ( .A(n292), .B(n291), .Z(n4494) );
  XNOR U3672 ( .A(n4495), .B(n4494), .Z(n4496) );
  XOR U3673 ( .A(n4497), .B(n4496), .Z(n3663) );
  NAND U3674 ( .A(n294), .B(n293), .Z(n298) );
  NAND U3675 ( .A(n296), .B(n295), .Z(n297) );
  NAND U3676 ( .A(n298), .B(n297), .Z(n3662) );
  XOR U3677 ( .A(n3663), .B(n3662), .Z(n3664) );
  NANDN U3678 ( .A(n300), .B(n299), .Z(n304) );
  NAND U3679 ( .A(n302), .B(n301), .Z(n303) );
  AND U3680 ( .A(n304), .B(n303), .Z(n3428) );
  NANDN U3681 ( .A(n306), .B(n305), .Z(n310) );
  NAND U3682 ( .A(n308), .B(n307), .Z(n309) );
  NAND U3683 ( .A(n310), .B(n309), .Z(n3429) );
  XNOR U3684 ( .A(n3428), .B(n3429), .Z(n3431) );
  NANDN U3685 ( .A(n312), .B(n311), .Z(n316) );
  NAND U3686 ( .A(n314), .B(n313), .Z(n315) );
  AND U3687 ( .A(n316), .B(n315), .Z(n3430) );
  XOR U3688 ( .A(n3431), .B(n3430), .Z(n3360) );
  NANDN U3689 ( .A(n318), .B(n317), .Z(n322) );
  NAND U3690 ( .A(n320), .B(n319), .Z(n321) );
  AND U3691 ( .A(n322), .B(n321), .Z(n3979) );
  NAND U3692 ( .A(n324), .B(n323), .Z(n328) );
  NAND U3693 ( .A(n326), .B(n325), .Z(n327) );
  AND U3694 ( .A(n328), .B(n327), .Z(n3980) );
  NANDN U3695 ( .A(n330), .B(n329), .Z(n334) );
  NAND U3696 ( .A(n332), .B(n331), .Z(n333) );
  AND U3697 ( .A(n334), .B(n333), .Z(n3981) );
  XOR U3698 ( .A(n3982), .B(n3981), .Z(n3358) );
  NANDN U3699 ( .A(n336), .B(n335), .Z(n340) );
  NAND U3700 ( .A(n338), .B(n337), .Z(n339) );
  AND U3701 ( .A(n340), .B(n339), .Z(n4302) );
  NANDN U3702 ( .A(n342), .B(n341), .Z(n346) );
  NAND U3703 ( .A(n344), .B(n343), .Z(n345) );
  NAND U3704 ( .A(n346), .B(n345), .Z(n4303) );
  XNOR U3705 ( .A(n4302), .B(n4303), .Z(n4305) );
  NANDN U3706 ( .A(n348), .B(n347), .Z(n352) );
  NAND U3707 ( .A(n350), .B(n349), .Z(n351) );
  AND U3708 ( .A(n352), .B(n351), .Z(n4304) );
  XNOR U3709 ( .A(n4305), .B(n4304), .Z(n3357) );
  XNOR U3710 ( .A(n3358), .B(n3357), .Z(n3359) );
  XOR U3711 ( .A(n3360), .B(n3359), .Z(n3561) );
  NANDN U3712 ( .A(n354), .B(n353), .Z(n358) );
  NANDN U3713 ( .A(n356), .B(n355), .Z(n357) );
  AND U3714 ( .A(n358), .B(n357), .Z(n3791) );
  NANDN U3715 ( .A(n360), .B(n359), .Z(n364) );
  NAND U3716 ( .A(n362), .B(n361), .Z(n363) );
  NAND U3717 ( .A(n364), .B(n363), .Z(n3457) );
  NANDN U3718 ( .A(n366), .B(n365), .Z(n370) );
  NAND U3719 ( .A(n368), .B(n367), .Z(n369) );
  AND U3720 ( .A(n370), .B(n369), .Z(n3456) );
  NANDN U3721 ( .A(n372), .B(n371), .Z(n376) );
  NAND U3722 ( .A(n374), .B(n373), .Z(n375) );
  AND U3723 ( .A(n376), .B(n375), .Z(n3455) );
  XNOR U3724 ( .A(n3456), .B(n3455), .Z(n377) );
  XNOR U3725 ( .A(n3457), .B(n377), .Z(n3788) );
  NANDN U3726 ( .A(n379), .B(n378), .Z(n383) );
  NANDN U3727 ( .A(n381), .B(n380), .Z(n382) );
  AND U3728 ( .A(n383), .B(n382), .Z(n3789) );
  XOR U3729 ( .A(n3788), .B(n3789), .Z(n3790) );
  XNOR U3730 ( .A(n3791), .B(n3790), .Z(n3560) );
  NANDN U3731 ( .A(n385), .B(n384), .Z(n389) );
  NAND U3732 ( .A(n387), .B(n386), .Z(n388) );
  AND U3733 ( .A(n389), .B(n388), .Z(n3830) );
  NANDN U3734 ( .A(n391), .B(n390), .Z(n395) );
  NAND U3735 ( .A(n393), .B(n392), .Z(n394) );
  AND U3736 ( .A(n395), .B(n394), .Z(n3831) );
  NANDN U3737 ( .A(n397), .B(n396), .Z(n401) );
  NAND U3738 ( .A(n399), .B(n398), .Z(n400) );
  AND U3739 ( .A(n401), .B(n400), .Z(n3832) );
  XOR U3740 ( .A(n3833), .B(n3832), .Z(n3382) );
  NANDN U3741 ( .A(n403), .B(n402), .Z(n407) );
  NANDN U3742 ( .A(n405), .B(n404), .Z(n406) );
  AND U3743 ( .A(n407), .B(n406), .Z(n3381) );
  XNOR U3744 ( .A(n3382), .B(n3381), .Z(n3384) );
  NANDN U3745 ( .A(n409), .B(n408), .Z(n413) );
  NANDN U3746 ( .A(n411), .B(n410), .Z(n412) );
  AND U3747 ( .A(n413), .B(n412), .Z(n3383) );
  XNOR U3748 ( .A(n3384), .B(n3383), .Z(n3559) );
  XNOR U3749 ( .A(n3561), .B(n3562), .Z(n3777) );
  NANDN U3750 ( .A(n415), .B(n414), .Z(n419) );
  NAND U3751 ( .A(n417), .B(n416), .Z(n418) );
  AND U3752 ( .A(n419), .B(n418), .Z(n4296) );
  NANDN U3753 ( .A(n421), .B(n420), .Z(n425) );
  NAND U3754 ( .A(n423), .B(n422), .Z(n424) );
  AND U3755 ( .A(n425), .B(n424), .Z(n4297) );
  NANDN U3756 ( .A(n427), .B(n426), .Z(n431) );
  NAND U3757 ( .A(n429), .B(n428), .Z(n430) );
  AND U3758 ( .A(n431), .B(n430), .Z(n4298) );
  XNOR U3759 ( .A(n4299), .B(n4298), .Z(n3801) );
  NANDN U3760 ( .A(n433), .B(n432), .Z(n437) );
  NANDN U3761 ( .A(n435), .B(n434), .Z(n436) );
  AND U3762 ( .A(n437), .B(n436), .Z(n3800) );
  NANDN U3763 ( .A(n439), .B(n438), .Z(n443) );
  NANDN U3764 ( .A(n441), .B(n440), .Z(n442) );
  AND U3765 ( .A(n443), .B(n442), .Z(n3803) );
  NANDN U3766 ( .A(n445), .B(n444), .Z(n449) );
  NAND U3767 ( .A(n447), .B(n446), .Z(n448) );
  NAND U3768 ( .A(n449), .B(n448), .Z(n4083) );
  NANDN U3769 ( .A(n451), .B(n450), .Z(n455) );
  NAND U3770 ( .A(n453), .B(n452), .Z(n454) );
  NAND U3771 ( .A(n455), .B(n454), .Z(n4082) );
  NANDN U3772 ( .A(n457), .B(n456), .Z(n461) );
  NAND U3773 ( .A(n459), .B(n458), .Z(n460) );
  AND U3774 ( .A(n461), .B(n460), .Z(n4081) );
  XOR U3775 ( .A(n4082), .B(n4081), .Z(n462) );
  XNOR U3776 ( .A(n4083), .B(n462), .Z(n3366) );
  NANDN U3777 ( .A(n464), .B(n463), .Z(n468) );
  NAND U3778 ( .A(n466), .B(n465), .Z(n467) );
  AND U3779 ( .A(n468), .B(n467), .Z(n3812) );
  NANDN U3780 ( .A(n470), .B(n469), .Z(n474) );
  NAND U3781 ( .A(n472), .B(n471), .Z(n473) );
  AND U3782 ( .A(n474), .B(n473), .Z(n3813) );
  NANDN U3783 ( .A(n476), .B(n475), .Z(n480) );
  NAND U3784 ( .A(n478), .B(n477), .Z(n479) );
  AND U3785 ( .A(n480), .B(n479), .Z(n3814) );
  XNOR U3786 ( .A(n3815), .B(n3814), .Z(n3364) );
  NANDN U3787 ( .A(n482), .B(n481), .Z(n486) );
  NANDN U3788 ( .A(n484), .B(n483), .Z(n485) );
  AND U3789 ( .A(n486), .B(n485), .Z(n3363) );
  XOR U3790 ( .A(n3366), .B(n3365), .Z(n3518) );
  NANDN U3791 ( .A(n488), .B(n487), .Z(n492) );
  NAND U3792 ( .A(n490), .B(n489), .Z(n491) );
  AND U3793 ( .A(n492), .B(n491), .Z(n3973) );
  NANDN U3794 ( .A(n494), .B(n493), .Z(n498) );
  NAND U3795 ( .A(n496), .B(n495), .Z(n497) );
  AND U3796 ( .A(n498), .B(n497), .Z(n3974) );
  NANDN U3797 ( .A(n500), .B(n499), .Z(n504) );
  NAND U3798 ( .A(n502), .B(n501), .Z(n503) );
  AND U3799 ( .A(n504), .B(n503), .Z(n3975) );
  XOR U3800 ( .A(n3976), .B(n3975), .Z(n3354) );
  NANDN U3801 ( .A(n506), .B(n505), .Z(n510) );
  NAND U3802 ( .A(n508), .B(n507), .Z(n509) );
  AND U3803 ( .A(n510), .B(n509), .Z(n4080) );
  NANDN U3804 ( .A(n512), .B(n511), .Z(n516) );
  NAND U3805 ( .A(n514), .B(n513), .Z(n515) );
  AND U3806 ( .A(n516), .B(n515), .Z(n4079) );
  NANDN U3807 ( .A(n518), .B(n517), .Z(n522) );
  NAND U3808 ( .A(n520), .B(n519), .Z(n521) );
  AND U3809 ( .A(n522), .B(n521), .Z(n4078) );
  NAND U3810 ( .A(n524), .B(n523), .Z(n528) );
  NAND U3811 ( .A(n526), .B(n525), .Z(n527) );
  NAND U3812 ( .A(n528), .B(n527), .Z(n3294) );
  NANDN U3813 ( .A(n530), .B(n529), .Z(n534) );
  NAND U3814 ( .A(n532), .B(n531), .Z(n533) );
  NAND U3815 ( .A(n534), .B(n533), .Z(n3293) );
  NANDN U3816 ( .A(n536), .B(n535), .Z(n540) );
  NAND U3817 ( .A(n538), .B(n537), .Z(n539) );
  AND U3818 ( .A(n540), .B(n539), .Z(n3292) );
  XOR U3819 ( .A(n3293), .B(n3292), .Z(n541) );
  XNOR U3820 ( .A(n3294), .B(n541), .Z(n3352) );
  XOR U3821 ( .A(n3351), .B(n3352), .Z(n3353) );
  XOR U3822 ( .A(n3354), .B(n3353), .Z(n3517) );
  XNOR U3823 ( .A(n3518), .B(n3517), .Z(n3519) );
  XOR U3824 ( .A(n3520), .B(n3519), .Z(n3776) );
  XNOR U3825 ( .A(n3777), .B(n3776), .Z(n542) );
  XNOR U3826 ( .A(n3775), .B(n542), .Z(n4034) );
  NANDN U3827 ( .A(n544), .B(n543), .Z(n548) );
  NANDN U3828 ( .A(n546), .B(n545), .Z(n547) );
  AND U3829 ( .A(n548), .B(n547), .Z(n3797) );
  NANDN U3830 ( .A(n550), .B(n549), .Z(n554) );
  NAND U3831 ( .A(n552), .B(n551), .Z(n553) );
  AND U3832 ( .A(n554), .B(n553), .Z(n3818) );
  NANDN U3833 ( .A(n556), .B(n555), .Z(n560) );
  NAND U3834 ( .A(n558), .B(n557), .Z(n559) );
  AND U3835 ( .A(n560), .B(n559), .Z(n3819) );
  NANDN U3836 ( .A(n562), .B(n561), .Z(n566) );
  NAND U3837 ( .A(n564), .B(n563), .Z(n565) );
  AND U3838 ( .A(n566), .B(n565), .Z(n3820) );
  XOR U3839 ( .A(n3821), .B(n3820), .Z(n3795) );
  NANDN U3840 ( .A(n568), .B(n567), .Z(n572) );
  NANDN U3841 ( .A(n570), .B(n569), .Z(n571) );
  AND U3842 ( .A(n572), .B(n571), .Z(n3794) );
  XNOR U3843 ( .A(n3795), .B(n3794), .Z(n3796) );
  XNOR U3844 ( .A(n3797), .B(n3796), .Z(n3629) );
  NANDN U3845 ( .A(n574), .B(n573), .Z(n578) );
  NANDN U3846 ( .A(n576), .B(n575), .Z(n577) );
  AND U3847 ( .A(n578), .B(n577), .Z(n3378) );
  NANDN U3848 ( .A(n580), .B(n579), .Z(n584) );
  NAND U3849 ( .A(n582), .B(n581), .Z(n583) );
  AND U3850 ( .A(n584), .B(n583), .Z(n4181) );
  NANDN U3851 ( .A(n586), .B(n585), .Z(n590) );
  NAND U3852 ( .A(n588), .B(n587), .Z(n589) );
  AND U3853 ( .A(n590), .B(n589), .Z(n4182) );
  NANDN U3854 ( .A(n592), .B(n591), .Z(n596) );
  NAND U3855 ( .A(n594), .B(n593), .Z(n595) );
  AND U3856 ( .A(n596), .B(n595), .Z(n4183) );
  XOR U3857 ( .A(n4184), .B(n4183), .Z(n3376) );
  NANDN U3858 ( .A(n598), .B(n597), .Z(n602) );
  NANDN U3859 ( .A(n600), .B(n599), .Z(n601) );
  AND U3860 ( .A(n602), .B(n601), .Z(n3375) );
  XNOR U3861 ( .A(n3376), .B(n3375), .Z(n3377) );
  XNOR U3862 ( .A(n3378), .B(n3377), .Z(n3627) );
  NANDN U3863 ( .A(n608), .B(n607), .Z(n612) );
  NAND U3864 ( .A(n610), .B(n609), .Z(n611) );
  AND U3865 ( .A(n612), .B(n611), .Z(n4344) );
  NANDN U3866 ( .A(n614), .B(n613), .Z(n618) );
  NAND U3867 ( .A(n616), .B(n615), .Z(n617) );
  NAND U3868 ( .A(n618), .B(n617), .Z(n4345) );
  XNOR U3869 ( .A(n4344), .B(n4345), .Z(n4347) );
  NANDN U3870 ( .A(n620), .B(n619), .Z(n624) );
  NAND U3871 ( .A(n622), .B(n621), .Z(n623) );
  AND U3872 ( .A(n624), .B(n623), .Z(n4346) );
  XOR U3873 ( .A(n4347), .B(n4346), .Z(n4585) );
  NANDN U3874 ( .A(n626), .B(n625), .Z(n630) );
  NANDN U3875 ( .A(n628), .B(n627), .Z(n629) );
  AND U3876 ( .A(n630), .B(n629), .Z(n4584) );
  XNOR U3877 ( .A(n4585), .B(n4584), .Z(n4586) );
  XOR U3878 ( .A(n4587), .B(n4586), .Z(n3626) );
  XNOR U3879 ( .A(n3629), .B(n3628), .Z(n3778) );
  NAND U3880 ( .A(n632), .B(n631), .Z(n636) );
  NAND U3881 ( .A(n634), .B(n633), .Z(n635) );
  AND U3882 ( .A(n636), .B(n635), .Z(n4425) );
  NANDN U3883 ( .A(n638), .B(n637), .Z(n642) );
  NAND U3884 ( .A(n640), .B(n639), .Z(n641) );
  AND U3885 ( .A(n642), .B(n641), .Z(n4320) );
  NANDN U3886 ( .A(n644), .B(n643), .Z(n648) );
  NAND U3887 ( .A(n646), .B(n645), .Z(n647) );
  NAND U3888 ( .A(n648), .B(n647), .Z(n4321) );
  XNOR U3889 ( .A(n4320), .B(n4321), .Z(n4323) );
  NANDN U3890 ( .A(n650), .B(n649), .Z(n654) );
  NAND U3891 ( .A(n652), .B(n651), .Z(n653) );
  AND U3892 ( .A(n654), .B(n653), .Z(n4322) );
  XOR U3893 ( .A(n4323), .B(n4322), .Z(n4423) );
  NANDN U3894 ( .A(n656), .B(n655), .Z(n660) );
  NANDN U3895 ( .A(n658), .B(n657), .Z(n659) );
  AND U3896 ( .A(n660), .B(n659), .Z(n4422) );
  XNOR U3897 ( .A(n4423), .B(n4422), .Z(n4424) );
  XOR U3898 ( .A(n4425), .B(n4424), .Z(n4195) );
  NANDN U3899 ( .A(n662), .B(n661), .Z(n666) );
  NANDN U3900 ( .A(n664), .B(n663), .Z(n665) );
  AND U3901 ( .A(n666), .B(n665), .Z(n4431) );
  NANDN U3902 ( .A(n668), .B(n667), .Z(n672) );
  NAND U3903 ( .A(n670), .B(n669), .Z(n671) );
  AND U3904 ( .A(n672), .B(n671), .Z(n4350) );
  NANDN U3905 ( .A(n674), .B(n673), .Z(n678) );
  NAND U3906 ( .A(n676), .B(n675), .Z(n677) );
  NAND U3907 ( .A(n678), .B(n677), .Z(n4351) );
  XNOR U3908 ( .A(n4350), .B(n4351), .Z(n4353) );
  NANDN U3909 ( .A(n680), .B(n679), .Z(n684) );
  NAND U3910 ( .A(n682), .B(n681), .Z(n683) );
  AND U3911 ( .A(n684), .B(n683), .Z(n4352) );
  XOR U3912 ( .A(n4353), .B(n4352), .Z(n4429) );
  NANDN U3913 ( .A(n686), .B(n685), .Z(n690) );
  NANDN U3914 ( .A(n688), .B(n687), .Z(n689) );
  AND U3915 ( .A(n690), .B(n689), .Z(n4428) );
  XNOR U3916 ( .A(n4429), .B(n4428), .Z(n4430) );
  XNOR U3917 ( .A(n4431), .B(n4430), .Z(n4194) );
  NANDN U3918 ( .A(n692), .B(n691), .Z(n696) );
  NANDN U3919 ( .A(n694), .B(n693), .Z(n695) );
  AND U3920 ( .A(n696), .B(n695), .Z(n4443) );
  NANDN U3921 ( .A(n698), .B(n697), .Z(n702) );
  NAND U3922 ( .A(n700), .B(n699), .Z(n701) );
  AND U3923 ( .A(n702), .B(n701), .Z(n4290) );
  NANDN U3924 ( .A(n704), .B(n703), .Z(n708) );
  NAND U3925 ( .A(n706), .B(n705), .Z(n707) );
  NAND U3926 ( .A(n708), .B(n707), .Z(n4291) );
  XNOR U3927 ( .A(n4290), .B(n4291), .Z(n4293) );
  NANDN U3928 ( .A(n710), .B(n709), .Z(n714) );
  NAND U3929 ( .A(n712), .B(n711), .Z(n713) );
  AND U3930 ( .A(n714), .B(n713), .Z(n4292) );
  XOR U3931 ( .A(n4293), .B(n4292), .Z(n4441) );
  NAND U3932 ( .A(n716), .B(n715), .Z(n720) );
  NAND U3933 ( .A(n718), .B(n717), .Z(n719) );
  AND U3934 ( .A(n720), .B(n719), .Z(n4440) );
  XNOR U3935 ( .A(n4441), .B(n4440), .Z(n4442) );
  XNOR U3936 ( .A(n4443), .B(n4442), .Z(n4193) );
  XOR U3937 ( .A(n4195), .B(n4196), .Z(n3780) );
  NANDN U3938 ( .A(n722), .B(n721), .Z(n726) );
  NANDN U3939 ( .A(n724), .B(n723), .Z(n725) );
  AND U3940 ( .A(n726), .B(n725), .Z(n4592) );
  NAND U3941 ( .A(n728), .B(n727), .Z(n732) );
  NAND U3942 ( .A(n730), .B(n729), .Z(n731) );
  AND U3943 ( .A(n732), .B(n731), .Z(n4338) );
  NAND U3944 ( .A(n734), .B(n733), .Z(n738) );
  NAND U3945 ( .A(n736), .B(n735), .Z(n737) );
  NAND U3946 ( .A(n738), .B(n737), .Z(n4339) );
  XNOR U3947 ( .A(n4338), .B(n4339), .Z(n4340) );
  NANDN U3948 ( .A(n740), .B(n739), .Z(n744) );
  NAND U3949 ( .A(n742), .B(n741), .Z(n743) );
  NAND U3950 ( .A(n744), .B(n743), .Z(n4341) );
  XNOR U3951 ( .A(n4340), .B(n4341), .Z(n4591) );
  NANDN U3952 ( .A(n746), .B(n745), .Z(n750) );
  NANDN U3953 ( .A(n748), .B(n747), .Z(n749) );
  AND U3954 ( .A(n750), .B(n749), .Z(n4590) );
  XNOR U3955 ( .A(n4591), .B(n4590), .Z(n751) );
  XNOR U3956 ( .A(n4592), .B(n751), .Z(n4090) );
  NANDN U3957 ( .A(n753), .B(n752), .Z(n757) );
  NANDN U3958 ( .A(n755), .B(n754), .Z(n756) );
  AND U3959 ( .A(n757), .B(n756), .Z(n4603) );
  NANDN U3960 ( .A(n759), .B(n758), .Z(n763) );
  NAND U3961 ( .A(n761), .B(n760), .Z(n762) );
  AND U3962 ( .A(n763), .B(n762), .Z(n4063) );
  NANDN U3963 ( .A(n765), .B(n764), .Z(n769) );
  NAND U3964 ( .A(n767), .B(n766), .Z(n768) );
  AND U3965 ( .A(n769), .B(n768), .Z(n4064) );
  NAND U3966 ( .A(n771), .B(n770), .Z(n775) );
  NAND U3967 ( .A(n773), .B(n772), .Z(n774) );
  AND U3968 ( .A(n775), .B(n774), .Z(n4065) );
  XOR U3969 ( .A(n4066), .B(n4065), .Z(n4601) );
  NANDN U3970 ( .A(n777), .B(n776), .Z(n781) );
  NANDN U3971 ( .A(n779), .B(n778), .Z(n780) );
  AND U3972 ( .A(n781), .B(n780), .Z(n4600) );
  XNOR U3973 ( .A(n4601), .B(n4600), .Z(n4602) );
  XNOR U3974 ( .A(n4603), .B(n4602), .Z(n4089) );
  NANDN U3975 ( .A(n783), .B(n782), .Z(n787) );
  NANDN U3976 ( .A(n785), .B(n784), .Z(n786) );
  AND U3977 ( .A(n787), .B(n786), .Z(n4608) );
  NANDN U3978 ( .A(n789), .B(n788), .Z(n793) );
  NAND U3979 ( .A(n791), .B(n790), .Z(n792) );
  AND U3980 ( .A(n793), .B(n792), .Z(n4051) );
  NANDN U3981 ( .A(n795), .B(n794), .Z(n799) );
  NAND U3982 ( .A(n797), .B(n796), .Z(n798) );
  AND U3983 ( .A(n799), .B(n798), .Z(n4052) );
  NANDN U3984 ( .A(n801), .B(n800), .Z(n805) );
  NAND U3985 ( .A(n803), .B(n802), .Z(n804) );
  AND U3986 ( .A(n805), .B(n804), .Z(n4054) );
  NANDN U3987 ( .A(n807), .B(n806), .Z(n811) );
  NANDN U3988 ( .A(n809), .B(n808), .Z(n810) );
  AND U3989 ( .A(n811), .B(n810), .Z(n4606) );
  XNOR U3990 ( .A(n4607), .B(n4606), .Z(n812) );
  XNOR U3991 ( .A(n4608), .B(n812), .Z(n4088) );
  XOR U3992 ( .A(n4090), .B(n4091), .Z(n3779) );
  XNOR U3993 ( .A(n3780), .B(n3779), .Z(n813) );
  XNOR U3994 ( .A(n3778), .B(n813), .Z(n4030) );
  IV U3995 ( .A(n4030), .Z(n4033) );
  NAND U3996 ( .A(n815), .B(n814), .Z(n819) );
  NAND U3997 ( .A(n817), .B(n816), .Z(n818) );
  AND U3998 ( .A(n819), .B(n818), .Z(n3413) );
  NAND U3999 ( .A(n821), .B(n820), .Z(n825) );
  NAND U4000 ( .A(n823), .B(n822), .Z(n824) );
  AND U4001 ( .A(n825), .B(n824), .Z(n3410) );
  NANDN U4002 ( .A(n827), .B(n826), .Z(n831) );
  NAND U4003 ( .A(n829), .B(n828), .Z(n830) );
  AND U4004 ( .A(n831), .B(n830), .Z(n4118) );
  NANDN U4005 ( .A(n833), .B(n832), .Z(n837) );
  NANDN U4006 ( .A(n835), .B(n834), .Z(n836) );
  AND U4007 ( .A(n837), .B(n836), .Z(n4119) );
  NANDN U4008 ( .A(n839), .B(n838), .Z(n843) );
  NAND U4009 ( .A(n841), .B(n840), .Z(n842) );
  AND U4010 ( .A(n843), .B(n842), .Z(n4120) );
  XNOR U4011 ( .A(n4121), .B(n4120), .Z(n4467) );
  NAND U4012 ( .A(n845), .B(n844), .Z(n849) );
  NAND U4013 ( .A(n847), .B(n846), .Z(n848) );
  AND U4014 ( .A(n849), .B(n848), .Z(n3836) );
  NAND U4015 ( .A(n851), .B(n850), .Z(n855) );
  NAND U4016 ( .A(n853), .B(n852), .Z(n854) );
  AND U4017 ( .A(n855), .B(n854), .Z(n3837) );
  NAND U4018 ( .A(n857), .B(n856), .Z(n861) );
  NAND U4019 ( .A(n859), .B(n858), .Z(n860) );
  AND U4020 ( .A(n861), .B(n860), .Z(n3838) );
  XNOR U4021 ( .A(n3839), .B(n3838), .Z(n4465) );
  NANDN U4022 ( .A(n863), .B(n862), .Z(n867) );
  NAND U4023 ( .A(n865), .B(n864), .Z(n866) );
  NAND U4024 ( .A(n867), .B(n866), .Z(n4145) );
  NANDN U4025 ( .A(n869), .B(n868), .Z(n873) );
  NAND U4026 ( .A(n871), .B(n870), .Z(n872) );
  NAND U4027 ( .A(n873), .B(n872), .Z(n4143) );
  NANDN U4028 ( .A(n874), .B(oglobal[0]), .Z(n878) );
  NANDN U4029 ( .A(n876), .B(n875), .Z(n877) );
  NAND U4030 ( .A(n878), .B(n877), .Z(n4142) );
  NANDN U4031 ( .A(n880), .B(n879), .Z(n884) );
  NAND U4032 ( .A(n882), .B(n881), .Z(n883) );
  AND U4033 ( .A(n884), .B(n883), .Z(n4130) );
  NANDN U4034 ( .A(n886), .B(n885), .Z(n890) );
  NAND U4035 ( .A(n888), .B(n887), .Z(n889) );
  AND U4036 ( .A(n890), .B(n889), .Z(n4131) );
  NANDN U4037 ( .A(n892), .B(n891), .Z(n896) );
  NAND U4038 ( .A(n894), .B(n893), .Z(n895) );
  AND U4039 ( .A(n896), .B(n895), .Z(n4132) );
  XNOR U4040 ( .A(n4133), .B(n4132), .Z(n3732) );
  NAND U4041 ( .A(n898), .B(n897), .Z(n902) );
  NAND U4042 ( .A(n900), .B(n899), .Z(n901) );
  AND U4043 ( .A(n902), .B(n901), .Z(n4217) );
  NAND U4044 ( .A(n904), .B(n903), .Z(n908) );
  NAND U4045 ( .A(n906), .B(n905), .Z(n907) );
  NAND U4046 ( .A(n908), .B(n907), .Z(n4218) );
  XNOR U4047 ( .A(n4217), .B(n4218), .Z(n4220) );
  NAND U4048 ( .A(n910), .B(n909), .Z(n914) );
  NAND U4049 ( .A(n912), .B(n911), .Z(n913) );
  AND U4050 ( .A(n914), .B(n913), .Z(n4219) );
  XNOR U4051 ( .A(n4220), .B(n4219), .Z(n3730) );
  NANDN U4052 ( .A(n916), .B(n915), .Z(n920) );
  NAND U4053 ( .A(n918), .B(n917), .Z(n919) );
  AND U4054 ( .A(n920), .B(n919), .Z(n4112) );
  NANDN U4055 ( .A(n922), .B(n921), .Z(n926) );
  NAND U4056 ( .A(n924), .B(n923), .Z(n925) );
  AND U4057 ( .A(n926), .B(n925), .Z(n4113) );
  NANDN U4058 ( .A(n928), .B(n927), .Z(n932) );
  NAND U4059 ( .A(n930), .B(n929), .Z(n931) );
  AND U4060 ( .A(n932), .B(n931), .Z(n4114) );
  XNOR U4061 ( .A(n4115), .B(n4114), .Z(n3729) );
  NANDN U4062 ( .A(n934), .B(n933), .Z(n938) );
  NAND U4063 ( .A(n936), .B(n935), .Z(n937) );
  AND U4064 ( .A(n938), .B(n937), .Z(n4100) );
  NANDN U4065 ( .A(n940), .B(n939), .Z(n944) );
  NAND U4066 ( .A(n942), .B(n941), .Z(n943) );
  AND U4067 ( .A(n944), .B(n943), .Z(n4101) );
  NANDN U4068 ( .A(n946), .B(n945), .Z(n950) );
  NAND U4069 ( .A(n948), .B(n947), .Z(n949) );
  AND U4070 ( .A(n950), .B(n949), .Z(n4102) );
  XOR U4071 ( .A(n4103), .B(n4102), .Z(n3756) );
  NAND U4072 ( .A(n952), .B(n951), .Z(n956) );
  NAND U4073 ( .A(n954), .B(n953), .Z(n955) );
  AND U4074 ( .A(n956), .B(n955), .Z(n4506) );
  NANDN U4075 ( .A(n958), .B(n957), .Z(n962) );
  NAND U4076 ( .A(n960), .B(n959), .Z(n961) );
  AND U4077 ( .A(n962), .B(n961), .Z(n4507) );
  NANDN U4078 ( .A(n964), .B(n963), .Z(n968) );
  NAND U4079 ( .A(n966), .B(n965), .Z(n967) );
  AND U4080 ( .A(n968), .B(n967), .Z(n4508) );
  XNOR U4081 ( .A(n4509), .B(n4508), .Z(n3754) );
  NANDN U4082 ( .A(n970), .B(n969), .Z(n974) );
  NANDN U4083 ( .A(n972), .B(n971), .Z(n973) );
  AND U4084 ( .A(n974), .B(n973), .Z(n3931) );
  NAND U4085 ( .A(n976), .B(n975), .Z(n980) );
  NAND U4086 ( .A(n978), .B(n977), .Z(n979) );
  AND U4087 ( .A(n980), .B(n979), .Z(n3932) );
  NANDN U4088 ( .A(n982), .B(n981), .Z(n986) );
  NAND U4089 ( .A(n984), .B(n983), .Z(n985) );
  AND U4090 ( .A(n986), .B(n985), .Z(n3933) );
  XNOR U4091 ( .A(n3934), .B(n3933), .Z(n3753) );
  XOR U4092 ( .A(n3756), .B(n3755), .Z(n3782) );
  XOR U4093 ( .A(n3783), .B(n3782), .Z(n3785) );
  XNOR U4094 ( .A(n3784), .B(n3785), .Z(n3411) );
  XNOR U4095 ( .A(n3413), .B(n3412), .Z(n4032) );
  IV U4096 ( .A(n4032), .Z(n4031) );
  XNOR U4097 ( .A(n4033), .B(n4031), .Z(n987) );
  XNOR U4098 ( .A(n4034), .B(n987), .Z(n3489) );
  NANDN U4099 ( .A(n989), .B(n988), .Z(n993) );
  NANDN U4100 ( .A(n991), .B(n990), .Z(n992) );
  AND U4101 ( .A(n993), .B(n992), .Z(n4311) );
  NANDN U4102 ( .A(n995), .B(n994), .Z(n999) );
  NAND U4103 ( .A(n997), .B(n996), .Z(n998) );
  NAND U4104 ( .A(n999), .B(n998), .Z(n3347) );
  NANDN U4105 ( .A(n1001), .B(n1000), .Z(n1005) );
  NAND U4106 ( .A(n1003), .B(n1002), .Z(n1004) );
  NAND U4107 ( .A(n1005), .B(n1004), .Z(n3346) );
  NANDN U4108 ( .A(n1007), .B(n1006), .Z(n1011) );
  NAND U4109 ( .A(n1009), .B(n1008), .Z(n1010) );
  AND U4110 ( .A(n1011), .B(n1010), .Z(n3345) );
  XOR U4111 ( .A(n3346), .B(n3345), .Z(n1012) );
  XOR U4112 ( .A(n3347), .B(n1012), .Z(n4309) );
  NANDN U4113 ( .A(n1014), .B(n1013), .Z(n1018) );
  NANDN U4114 ( .A(n1016), .B(n1015), .Z(n1017) );
  AND U4115 ( .A(n1018), .B(n1017), .Z(n4308) );
  XNOR U4116 ( .A(n4309), .B(n4308), .Z(n4310) );
  XNOR U4117 ( .A(n4311), .B(n4310), .Z(n3556) );
  NAND U4118 ( .A(n1020), .B(n1019), .Z(n1024) );
  NAND U4119 ( .A(n1022), .B(n1021), .Z(n1023) );
  AND U4120 ( .A(n1024), .B(n1023), .Z(n4536) );
  NANDN U4121 ( .A(n1026), .B(n1025), .Z(n1030) );
  NAND U4122 ( .A(n1028), .B(n1027), .Z(n1029) );
  AND U4123 ( .A(n1030), .B(n1029), .Z(n4537) );
  NANDN U4124 ( .A(n1032), .B(n1031), .Z(n1036) );
  NAND U4125 ( .A(n1034), .B(n1033), .Z(n1035) );
  AND U4126 ( .A(n1036), .B(n1035), .Z(n4538) );
  XOR U4127 ( .A(n4539), .B(n4538), .Z(n4377) );
  NANDN U4128 ( .A(n1038), .B(n1037), .Z(n1042) );
  NAND U4129 ( .A(n1040), .B(n1039), .Z(n1041) );
  AND U4130 ( .A(n1042), .B(n1041), .Z(n3907) );
  NANDN U4131 ( .A(n1044), .B(n1043), .Z(n1048) );
  NAND U4132 ( .A(n1046), .B(n1045), .Z(n1047) );
  AND U4133 ( .A(n1048), .B(n1047), .Z(n3908) );
  NANDN U4134 ( .A(n1050), .B(n1049), .Z(n1054) );
  NAND U4135 ( .A(n1052), .B(n1051), .Z(n1053) );
  AND U4136 ( .A(n1054), .B(n1053), .Z(n3909) );
  XOR U4137 ( .A(n3910), .B(n3909), .Z(n4375) );
  NANDN U4138 ( .A(n1056), .B(n1055), .Z(n1060) );
  NANDN U4139 ( .A(n1058), .B(n1057), .Z(n1059) );
  AND U4140 ( .A(n1060), .B(n1059), .Z(n4374) );
  XNOR U4141 ( .A(n4375), .B(n4374), .Z(n4376) );
  XOR U4142 ( .A(n4377), .B(n4376), .Z(n3554) );
  XOR U4143 ( .A(n3554), .B(n3553), .Z(n3555) );
  XOR U4144 ( .A(n3556), .B(n3555), .Z(n3393) );
  NANDN U4145 ( .A(n1066), .B(n1065), .Z(n1070) );
  NANDN U4146 ( .A(n1068), .B(n1067), .Z(n1069) );
  AND U4147 ( .A(n1070), .B(n1069), .Z(n4251) );
  NANDN U4148 ( .A(n1072), .B(n1071), .Z(n1076) );
  NAND U4149 ( .A(n1074), .B(n1073), .Z(n1075) );
  AND U4150 ( .A(n1076), .B(n1075), .Z(n3440) );
  NAND U4151 ( .A(n1078), .B(n1077), .Z(n1082) );
  NAND U4152 ( .A(n1080), .B(n1079), .Z(n1081) );
  NAND U4153 ( .A(n1082), .B(n1081), .Z(n3441) );
  XNOR U4154 ( .A(n3440), .B(n3441), .Z(n3443) );
  NANDN U4155 ( .A(n1084), .B(n1083), .Z(n1088) );
  NAND U4156 ( .A(n1086), .B(n1085), .Z(n1087) );
  AND U4157 ( .A(n1088), .B(n1087), .Z(n3442) );
  XNOR U4158 ( .A(n3443), .B(n3442), .Z(n4249) );
  NANDN U4159 ( .A(n1090), .B(n1089), .Z(n1094) );
  NANDN U4160 ( .A(n1092), .B(n1091), .Z(n1093) );
  AND U4161 ( .A(n1094), .B(n1093), .Z(n4248) );
  XNOR U4162 ( .A(n4251), .B(n4250), .Z(n3568) );
  NAND U4163 ( .A(n1096), .B(n1095), .Z(n1100) );
  NAND U4164 ( .A(n1098), .B(n1097), .Z(n1099) );
  NAND U4165 ( .A(n1100), .B(n1099), .Z(n3566) );
  NAND U4166 ( .A(n1102), .B(n1101), .Z(n1106) );
  NAND U4167 ( .A(n1104), .B(n1103), .Z(n1105) );
  AND U4168 ( .A(n1106), .B(n1105), .Z(n3691) );
  NAND U4169 ( .A(n1108), .B(n1107), .Z(n1112) );
  NAND U4170 ( .A(n1110), .B(n1109), .Z(n1111) );
  NAND U4171 ( .A(n1112), .B(n1111), .Z(n3689) );
  NANDN U4172 ( .A(n1114), .B(n1113), .Z(n1118) );
  NAND U4173 ( .A(n1116), .B(n1115), .Z(n1117) );
  AND U4174 ( .A(n1118), .B(n1117), .Z(n4404) );
  NANDN U4175 ( .A(n1120), .B(n1119), .Z(n1124) );
  NAND U4176 ( .A(n1122), .B(n1121), .Z(n1123) );
  AND U4177 ( .A(n1124), .B(n1123), .Z(n4405) );
  NANDN U4178 ( .A(n1126), .B(n1125), .Z(n1130) );
  NAND U4179 ( .A(n1128), .B(n1127), .Z(n1129) );
  AND U4180 ( .A(n1130), .B(n1129), .Z(n4406) );
  XNOR U4181 ( .A(n4407), .B(n4406), .Z(n3690) );
  XNOR U4182 ( .A(n3689), .B(n3690), .Z(n1131) );
  XNOR U4183 ( .A(n3691), .B(n1131), .Z(n3565) );
  NAND U4184 ( .A(n1133), .B(n1132), .Z(n1137) );
  NAND U4185 ( .A(n1135), .B(n1134), .Z(n1136) );
  NAND U4186 ( .A(n1137), .B(n1136), .Z(n3635) );
  NAND U4187 ( .A(n1139), .B(n1138), .Z(n1143) );
  NAND U4188 ( .A(n1141), .B(n1140), .Z(n1142) );
  NAND U4189 ( .A(n1143), .B(n1142), .Z(n3633) );
  NAND U4190 ( .A(n1145), .B(n1144), .Z(n1149) );
  NAND U4191 ( .A(n1147), .B(n1146), .Z(n1148) );
  NAND U4192 ( .A(n1149), .B(n1148), .Z(n3632) );
  XNOR U4193 ( .A(n3395), .B(n3394), .Z(n1150) );
  XOR U4194 ( .A(n3393), .B(n1150), .Z(n4029) );
  NANDN U4195 ( .A(n1152), .B(n1151), .Z(n1156) );
  NANDN U4196 ( .A(n1154), .B(n1153), .Z(n1155) );
  AND U4197 ( .A(n1156), .B(n1155), .Z(n3470) );
  NANDN U4198 ( .A(n1158), .B(n1157), .Z(n1162) );
  NAND U4199 ( .A(n1160), .B(n1159), .Z(n1161) );
  AND U4200 ( .A(n1162), .B(n1161), .Z(n4205) );
  NANDN U4201 ( .A(n1164), .B(n1163), .Z(n1168) );
  NAND U4202 ( .A(n1166), .B(n1165), .Z(n1167) );
  AND U4203 ( .A(n1168), .B(n1167), .Z(n4206) );
  NANDN U4204 ( .A(n1170), .B(n1169), .Z(n1174) );
  NAND U4205 ( .A(n1172), .B(n1171), .Z(n1173) );
  AND U4206 ( .A(n1174), .B(n1173), .Z(n4208) );
  NANDN U4207 ( .A(n1176), .B(n1175), .Z(n1180) );
  NANDN U4208 ( .A(n1178), .B(n1177), .Z(n1179) );
  AND U4209 ( .A(n1180), .B(n1179), .Z(n3468) );
  XNOR U4210 ( .A(n3469), .B(n3468), .Z(n1181) );
  XNOR U4211 ( .A(n3470), .B(n1181), .Z(n3670) );
  NANDN U4212 ( .A(n1183), .B(n1182), .Z(n1187) );
  NANDN U4213 ( .A(n1185), .B(n1184), .Z(n1186) );
  AND U4214 ( .A(n1187), .B(n1186), .Z(n4485) );
  NANDN U4215 ( .A(n1189), .B(n1188), .Z(n1193) );
  NAND U4216 ( .A(n1191), .B(n1190), .Z(n1192) );
  AND U4217 ( .A(n1193), .B(n1192), .Z(n4057) );
  NAND U4218 ( .A(n1195), .B(n1194), .Z(n1199) );
  NAND U4219 ( .A(n1197), .B(n1196), .Z(n1198) );
  AND U4220 ( .A(n1199), .B(n1198), .Z(n4058) );
  NAND U4221 ( .A(n1201), .B(n1200), .Z(n1205) );
  NAND U4222 ( .A(n1203), .B(n1202), .Z(n1204) );
  AND U4223 ( .A(n1205), .B(n1204), .Z(n4059) );
  XOR U4224 ( .A(n4060), .B(n4059), .Z(n4483) );
  NANDN U4225 ( .A(n1207), .B(n1206), .Z(n1211) );
  NANDN U4226 ( .A(n1209), .B(n1208), .Z(n1210) );
  AND U4227 ( .A(n1211), .B(n1210), .Z(n4482) );
  XNOR U4228 ( .A(n4483), .B(n4482), .Z(n4484) );
  XNOR U4229 ( .A(n4485), .B(n4484), .Z(n3669) );
  NANDN U4230 ( .A(n1213), .B(n1212), .Z(n1217) );
  NAND U4231 ( .A(n1215), .B(n1214), .Z(n1216) );
  NAND U4232 ( .A(n1217), .B(n1216), .Z(n3454) );
  NANDN U4233 ( .A(n1219), .B(n1218), .Z(n1223) );
  NAND U4234 ( .A(n1221), .B(n1220), .Z(n1222) );
  AND U4235 ( .A(n1223), .B(n1222), .Z(n3453) );
  NANDN U4236 ( .A(n1225), .B(n1224), .Z(n1229) );
  NAND U4237 ( .A(n1227), .B(n1226), .Z(n1228) );
  AND U4238 ( .A(n1229), .B(n1228), .Z(n3452) );
  XNOR U4239 ( .A(n3453), .B(n3452), .Z(n1230) );
  XNOR U4240 ( .A(n3454), .B(n1230), .Z(n3969) );
  NAND U4241 ( .A(n1232), .B(n1231), .Z(n1236) );
  NAND U4242 ( .A(n1234), .B(n1233), .Z(n1235) );
  AND U4243 ( .A(n1236), .B(n1235), .Z(n4155) );
  NANDN U4244 ( .A(n1238), .B(n1237), .Z(n1242) );
  NAND U4245 ( .A(n1240), .B(n1239), .Z(n1241) );
  AND U4246 ( .A(n1242), .B(n1241), .Z(n4156) );
  NAND U4247 ( .A(n1244), .B(n1243), .Z(n1248) );
  NAND U4248 ( .A(n1246), .B(n1245), .Z(n1247) );
  AND U4249 ( .A(n1248), .B(n1247), .Z(n4157) );
  XOR U4250 ( .A(n4158), .B(n4157), .Z(n3968) );
  NANDN U4251 ( .A(n1250), .B(n1249), .Z(n1254) );
  NANDN U4252 ( .A(n1252), .B(n1251), .Z(n1253) );
  AND U4253 ( .A(n1254), .B(n1253), .Z(n3967) );
  XNOR U4254 ( .A(n3968), .B(n3967), .Z(n3970) );
  XNOR U4255 ( .A(n3969), .B(n3970), .Z(n3668) );
  XOR U4256 ( .A(n3670), .B(n3671), .Z(n3657) );
  NANDN U4257 ( .A(n1256), .B(n1255), .Z(n1260) );
  NAND U4258 ( .A(n1258), .B(n1257), .Z(n1259) );
  AND U4259 ( .A(n1260), .B(n1259), .Z(n4015) );
  NANDN U4260 ( .A(n1262), .B(n1261), .Z(n1266) );
  NAND U4261 ( .A(n1264), .B(n1263), .Z(n1265) );
  AND U4262 ( .A(n1266), .B(n1265), .Z(n4016) );
  NAND U4263 ( .A(n1268), .B(n1267), .Z(n1272) );
  NAND U4264 ( .A(n1270), .B(n1269), .Z(n1271) );
  AND U4265 ( .A(n1272), .B(n1271), .Z(n4017) );
  XOR U4266 ( .A(n4018), .B(n4017), .Z(n3994) );
  NANDN U4267 ( .A(n1274), .B(n1273), .Z(n1278) );
  NAND U4268 ( .A(n1276), .B(n1275), .Z(n1277) );
  AND U4269 ( .A(n1278), .B(n1277), .Z(n3943) );
  NAND U4270 ( .A(n1280), .B(n1279), .Z(n1284) );
  NAND U4271 ( .A(n1282), .B(n1281), .Z(n1283) );
  NAND U4272 ( .A(n1284), .B(n1283), .Z(n3944) );
  XNOR U4273 ( .A(n3943), .B(n3944), .Z(n3946) );
  NANDN U4274 ( .A(n1286), .B(n1285), .Z(n1290) );
  NAND U4275 ( .A(n1288), .B(n1287), .Z(n1289) );
  AND U4276 ( .A(n1290), .B(n1289), .Z(n3945) );
  XOR U4277 ( .A(n3946), .B(n3945), .Z(n3992) );
  NANDN U4278 ( .A(n1292), .B(n1291), .Z(n1296) );
  NANDN U4279 ( .A(n1294), .B(n1293), .Z(n1295) );
  AND U4280 ( .A(n1296), .B(n1295), .Z(n3991) );
  XNOR U4281 ( .A(n3992), .B(n3991), .Z(n3993) );
  XOR U4282 ( .A(n3994), .B(n3993), .Z(n3676) );
  NAND U4283 ( .A(n1298), .B(n1297), .Z(n1302) );
  NAND U4284 ( .A(n1300), .B(n1299), .Z(n1301) );
  AND U4285 ( .A(n1302), .B(n1301), .Z(n3762) );
  NAND U4286 ( .A(n1304), .B(n1303), .Z(n1308) );
  NAND U4287 ( .A(n1306), .B(n1305), .Z(n1307) );
  NAND U4288 ( .A(n1308), .B(n1307), .Z(n4192) );
  NAND U4289 ( .A(n1310), .B(n1309), .Z(n1314) );
  NAND U4290 ( .A(n1312), .B(n1311), .Z(n1313) );
  NAND U4291 ( .A(n1314), .B(n1313), .Z(n4191) );
  NAND U4292 ( .A(n1316), .B(n1315), .Z(n1320) );
  NAND U4293 ( .A(n1318), .B(n1317), .Z(n1319) );
  AND U4294 ( .A(n1320), .B(n1319), .Z(n4190) );
  XOR U4295 ( .A(n4191), .B(n4190), .Z(n1321) );
  XOR U4296 ( .A(n4192), .B(n1321), .Z(n3760) );
  NANDN U4297 ( .A(n1323), .B(n1322), .Z(n1327) );
  NANDN U4298 ( .A(n1325), .B(n1324), .Z(n1326) );
  AND U4299 ( .A(n1327), .B(n1326), .Z(n3759) );
  XNOR U4300 ( .A(n3760), .B(n3759), .Z(n3761) );
  XNOR U4301 ( .A(n3762), .B(n3761), .Z(n3675) );
  NANDN U4302 ( .A(n1329), .B(n1328), .Z(n1333) );
  NANDN U4303 ( .A(n1331), .B(n1330), .Z(n1332) );
  NAND U4304 ( .A(n1333), .B(n1332), .Z(n3460) );
  NANDN U4305 ( .A(n1335), .B(n1334), .Z(n1339) );
  NAND U4306 ( .A(n1337), .B(n1336), .Z(n1338) );
  NAND U4307 ( .A(n1339), .B(n1338), .Z(n3291) );
  NANDN U4308 ( .A(n1341), .B(n1340), .Z(n1345) );
  NAND U4309 ( .A(n1343), .B(n1342), .Z(n1344) );
  NAND U4310 ( .A(n1345), .B(n1344), .Z(n3290) );
  NANDN U4311 ( .A(n1347), .B(n1346), .Z(n1351) );
  NAND U4312 ( .A(n1349), .B(n1348), .Z(n1350) );
  AND U4313 ( .A(n1351), .B(n1350), .Z(n3289) );
  XOR U4314 ( .A(n3290), .B(n3289), .Z(n1352) );
  XNOR U4315 ( .A(n3291), .B(n1352), .Z(n3459) );
  NAND U4316 ( .A(n1354), .B(n1353), .Z(n1358) );
  NAND U4317 ( .A(n1356), .B(n1355), .Z(n1357) );
  AND U4318 ( .A(n1358), .B(n1357), .Z(n3985) );
  NAND U4319 ( .A(n1360), .B(n1359), .Z(n1364) );
  NAND U4320 ( .A(n1362), .B(n1361), .Z(n1363) );
  AND U4321 ( .A(n1364), .B(n1363), .Z(n3986) );
  NAND U4322 ( .A(n1366), .B(n1365), .Z(n1370) );
  NAND U4323 ( .A(n1368), .B(n1367), .Z(n1369) );
  AND U4324 ( .A(n1370), .B(n1369), .Z(n3987) );
  XOR U4325 ( .A(n3988), .B(n3987), .Z(n3458) );
  XOR U4326 ( .A(n3459), .B(n3458), .Z(n1371) );
  XNOR U4327 ( .A(n3460), .B(n1371), .Z(n3674) );
  XOR U4328 ( .A(n3676), .B(n3677), .Z(n3656) );
  XOR U4329 ( .A(n3657), .B(n3656), .Z(n3659) );
  NANDN U4330 ( .A(n1373), .B(n1372), .Z(n1377) );
  NANDN U4331 ( .A(n1375), .B(n1374), .Z(n1376) );
  NAND U4332 ( .A(n1377), .B(n1376), .Z(n4177) );
  NANDN U4333 ( .A(n1379), .B(n1378), .Z(n1383) );
  NAND U4334 ( .A(n1381), .B(n1380), .Z(n1382) );
  AND U4335 ( .A(n1383), .B(n1382), .Z(n3949) );
  NANDN U4336 ( .A(n1385), .B(n1384), .Z(n1389) );
  NAND U4337 ( .A(n1387), .B(n1386), .Z(n1388) );
  AND U4338 ( .A(n1389), .B(n1388), .Z(n3950) );
  NANDN U4339 ( .A(n1391), .B(n1390), .Z(n1395) );
  NAND U4340 ( .A(n1393), .B(n1392), .Z(n1394) );
  AND U4341 ( .A(n1395), .B(n1394), .Z(n3952) );
  IV U4342 ( .A(n4173), .Z(n4176) );
  NANDN U4343 ( .A(n1397), .B(n1396), .Z(n1401) );
  NANDN U4344 ( .A(n1399), .B(n1398), .Z(n1400) );
  NAND U4345 ( .A(n1401), .B(n1400), .Z(n4175) );
  IV U4346 ( .A(n4175), .Z(n4174) );
  XNOR U4347 ( .A(n4176), .B(n4174), .Z(n1402) );
  XOR U4348 ( .A(n4177), .B(n1402), .Z(n3513) );
  NANDN U4349 ( .A(n1404), .B(n1403), .Z(n1408) );
  NANDN U4350 ( .A(n1406), .B(n1405), .Z(n1407) );
  AND U4351 ( .A(n1408), .B(n1407), .Z(n3726) );
  NANDN U4352 ( .A(n1410), .B(n1409), .Z(n1414) );
  NAND U4353 ( .A(n1412), .B(n1411), .Z(n1413) );
  AND U4354 ( .A(n1414), .B(n1413), .Z(n3298) );
  NANDN U4355 ( .A(n1416), .B(n1415), .Z(n1420) );
  NAND U4356 ( .A(n1418), .B(n1417), .Z(n1419) );
  AND U4357 ( .A(n1420), .B(n1419), .Z(n3299) );
  NAND U4358 ( .A(n1422), .B(n1421), .Z(n1426) );
  NAND U4359 ( .A(n1424), .B(n1423), .Z(n1425) );
  AND U4360 ( .A(n1426), .B(n1425), .Z(n3300) );
  XNOR U4361 ( .A(n3301), .B(n3300), .Z(n3724) );
  NANDN U4362 ( .A(n1428), .B(n1427), .Z(n1432) );
  NANDN U4363 ( .A(n1430), .B(n1429), .Z(n1431) );
  AND U4364 ( .A(n1432), .B(n1431), .Z(n3723) );
  XOR U4365 ( .A(n3726), .B(n3725), .Z(n3512) );
  NANDN U4366 ( .A(n1434), .B(n1433), .Z(n1438) );
  NANDN U4367 ( .A(n1436), .B(n1435), .Z(n1437) );
  NAND U4368 ( .A(n1438), .B(n1437), .Z(n3335) );
  NANDN U4369 ( .A(n1440), .B(n1439), .Z(n1444) );
  NAND U4370 ( .A(n1442), .B(n1441), .Z(n1443) );
  AND U4371 ( .A(n1444), .B(n1443), .Z(n4161) );
  NANDN U4372 ( .A(n1446), .B(n1445), .Z(n1450) );
  NAND U4373 ( .A(n1448), .B(n1447), .Z(n1449) );
  AND U4374 ( .A(n1450), .B(n1449), .Z(n4162) );
  NANDN U4375 ( .A(n1452), .B(n1451), .Z(n1456) );
  NAND U4376 ( .A(n1454), .B(n1453), .Z(n1455) );
  AND U4377 ( .A(n1456), .B(n1455), .Z(n4164) );
  IV U4378 ( .A(n3331), .Z(n3334) );
  NANDN U4379 ( .A(n1458), .B(n1457), .Z(n1462) );
  NANDN U4380 ( .A(n1460), .B(n1459), .Z(n1461) );
  NAND U4381 ( .A(n1462), .B(n1461), .Z(n3333) );
  IV U4382 ( .A(n3333), .Z(n3332) );
  XNOR U4383 ( .A(n3512), .B(n3511), .Z(n3514) );
  XOR U4384 ( .A(n3513), .B(n3514), .Z(n3658) );
  XNOR U4385 ( .A(n3659), .B(n3658), .Z(n4028) );
  NANDN U4386 ( .A(n1464), .B(n1463), .Z(n1468) );
  NANDN U4387 ( .A(n1466), .B(n1465), .Z(n1467) );
  AND U4388 ( .A(n1468), .B(n1467), .Z(n4527) );
  NAND U4389 ( .A(n1470), .B(n1469), .Z(n1474) );
  NAND U4390 ( .A(n1472), .B(n1471), .Z(n1473) );
  AND U4391 ( .A(n1474), .B(n1473), .Z(n4167) );
  NAND U4392 ( .A(n1476), .B(n1475), .Z(n1480) );
  NAND U4393 ( .A(n1478), .B(n1477), .Z(n1479) );
  NAND U4394 ( .A(n1480), .B(n1479), .Z(n4168) );
  XNOR U4395 ( .A(n4167), .B(n4168), .Z(n4170) );
  NAND U4396 ( .A(n1482), .B(n1481), .Z(n1486) );
  NAND U4397 ( .A(n1484), .B(n1483), .Z(n1485) );
  AND U4398 ( .A(n1486), .B(n1485), .Z(n4169) );
  XOR U4399 ( .A(n4170), .B(n4169), .Z(n4525) );
  NANDN U4400 ( .A(n1488), .B(n1487), .Z(n1492) );
  NANDN U4401 ( .A(n1490), .B(n1489), .Z(n1491) );
  AND U4402 ( .A(n1492), .B(n1491), .Z(n4524) );
  XNOR U4403 ( .A(n4525), .B(n4524), .Z(n4526) );
  XOR U4404 ( .A(n4527), .B(n4526), .Z(n4287) );
  NANDN U4405 ( .A(n1494), .B(n1493), .Z(n1498) );
  OR U4406 ( .A(n1496), .B(n1495), .Z(n1497) );
  AND U4407 ( .A(n1498), .B(n1497), .Z(n4285) );
  NAND U4408 ( .A(n1500), .B(n1499), .Z(n1504) );
  NAND U4409 ( .A(n1502), .B(n1501), .Z(n1503) );
  AND U4410 ( .A(n1504), .B(n1503), .Z(n4272) );
  NANDN U4411 ( .A(n1506), .B(n1505), .Z(n1510) );
  NAND U4412 ( .A(n1508), .B(n1507), .Z(n1509) );
  AND U4413 ( .A(n1510), .B(n1509), .Z(n4273) );
  NANDN U4414 ( .A(n1512), .B(n1511), .Z(n1516) );
  NAND U4415 ( .A(n1514), .B(n1513), .Z(n1515) );
  AND U4416 ( .A(n1516), .B(n1515), .Z(n4274) );
  XOR U4417 ( .A(n4275), .B(n4274), .Z(n4401) );
  NANDN U4418 ( .A(n1518), .B(n1517), .Z(n1522) );
  NAND U4419 ( .A(n1520), .B(n1519), .Z(n1521) );
  AND U4420 ( .A(n1522), .B(n1521), .Z(n4229) );
  NANDN U4421 ( .A(n1524), .B(n1523), .Z(n1528) );
  NAND U4422 ( .A(n1526), .B(n1525), .Z(n1527) );
  NAND U4423 ( .A(n1528), .B(n1527), .Z(n4230) );
  XNOR U4424 ( .A(n4229), .B(n4230), .Z(n4232) );
  NANDN U4425 ( .A(n1530), .B(n1529), .Z(n1534) );
  NAND U4426 ( .A(n1532), .B(n1531), .Z(n1533) );
  AND U4427 ( .A(n1534), .B(n1533), .Z(n4231) );
  XOR U4428 ( .A(n4232), .B(n4231), .Z(n4399) );
  NANDN U4429 ( .A(n1536), .B(n1535), .Z(n1540) );
  NANDN U4430 ( .A(n1538), .B(n1537), .Z(n1539) );
  AND U4431 ( .A(n1540), .B(n1539), .Z(n4398) );
  XNOR U4432 ( .A(n4399), .B(n4398), .Z(n4400) );
  XOR U4433 ( .A(n4401), .B(n4400), .Z(n4284) );
  XNOR U4434 ( .A(n4285), .B(n4284), .Z(n4286) );
  XNOR U4435 ( .A(n4287), .B(n4286), .Z(n3574) );
  NANDN U4436 ( .A(n1542), .B(n1541), .Z(n1546) );
  NAND U4437 ( .A(n1544), .B(n1543), .Z(n1545) );
  AND U4438 ( .A(n1546), .B(n1545), .Z(n3602) );
  NANDN U4439 ( .A(n1548), .B(n1547), .Z(n1552) );
  NAND U4440 ( .A(n1550), .B(n1549), .Z(n1551) );
  AND U4441 ( .A(n1552), .B(n1551), .Z(n3603) );
  NANDN U4442 ( .A(n1554), .B(n1553), .Z(n1558) );
  NAND U4443 ( .A(n1556), .B(n1555), .Z(n1557) );
  AND U4444 ( .A(n1558), .B(n1557), .Z(n3604) );
  XNOR U4445 ( .A(n3605), .B(n3604), .Z(n4000) );
  NANDN U4446 ( .A(n1560), .B(n1559), .Z(n1564) );
  NAND U4447 ( .A(n1562), .B(n1561), .Z(n1563) );
  AND U4448 ( .A(n1564), .B(n1563), .Z(n4106) );
  NAND U4449 ( .A(n1566), .B(n1565), .Z(n1570) );
  NAND U4450 ( .A(n1568), .B(n1567), .Z(n1569) );
  AND U4451 ( .A(n1570), .B(n1569), .Z(n4107) );
  NANDN U4452 ( .A(n1572), .B(n1571), .Z(n1576) );
  NAND U4453 ( .A(n1574), .B(n1573), .Z(n1575) );
  AND U4454 ( .A(n1576), .B(n1575), .Z(n4108) );
  XNOR U4455 ( .A(n4109), .B(n4108), .Z(n3998) );
  NANDN U4456 ( .A(n1578), .B(n1577), .Z(n1582) );
  NANDN U4457 ( .A(n1580), .B(n1579), .Z(n1581) );
  AND U4458 ( .A(n1582), .B(n1581), .Z(n3997) );
  NANDN U4459 ( .A(n1584), .B(n1583), .Z(n1588) );
  NANDN U4460 ( .A(n1586), .B(n1585), .Z(n1587) );
  AND U4461 ( .A(n1588), .B(n1587), .Z(n4245) );
  NAND U4462 ( .A(n1590), .B(n1589), .Z(n1594) );
  NAND U4463 ( .A(n1592), .B(n1591), .Z(n1593) );
  AND U4464 ( .A(n1594), .B(n1593), .Z(n3588) );
  NAND U4465 ( .A(n1596), .B(n1595), .Z(n1600) );
  NAND U4466 ( .A(n1598), .B(n1597), .Z(n1599) );
  AND U4467 ( .A(n1600), .B(n1599), .Z(n3587) );
  NANDN U4468 ( .A(n1602), .B(n1601), .Z(n1606) );
  NAND U4469 ( .A(n1604), .B(n1603), .Z(n1605) );
  AND U4470 ( .A(n1606), .B(n1605), .Z(n3586) );
  NANDN U4471 ( .A(n1608), .B(n1607), .Z(n1612) );
  NANDN U4472 ( .A(n1610), .B(n1609), .Z(n1611) );
  AND U4473 ( .A(n1612), .B(n1611), .Z(n4243) );
  XOR U4474 ( .A(n4242), .B(n4243), .Z(n4244) );
  XOR U4475 ( .A(n4245), .B(n4244), .Z(n3872) );
  NANDN U4476 ( .A(n1614), .B(n1613), .Z(n1618) );
  NAND U4477 ( .A(n1616), .B(n1615), .Z(n1617) );
  AND U4478 ( .A(n1618), .B(n1617), .Z(n3865) );
  NAND U4479 ( .A(n1620), .B(n1619), .Z(n1624) );
  NAND U4480 ( .A(n1622), .B(n1621), .Z(n1623) );
  NAND U4481 ( .A(n1624), .B(n1623), .Z(n3866) );
  XNOR U4482 ( .A(n3865), .B(n3866), .Z(n3868) );
  NAND U4483 ( .A(n1626), .B(n1625), .Z(n1630) );
  NAND U4484 ( .A(n1628), .B(n1627), .Z(n1629) );
  AND U4485 ( .A(n1630), .B(n1629), .Z(n3867) );
  XNOR U4486 ( .A(n3868), .B(n3867), .Z(n3896) );
  NANDN U4487 ( .A(n1632), .B(n1631), .Z(n1636) );
  NANDN U4488 ( .A(n1634), .B(n1633), .Z(n1635) );
  AND U4489 ( .A(n1636), .B(n1635), .Z(n3895) );
  NAND U4490 ( .A(n1638), .B(n1637), .Z(n1642) );
  NAND U4491 ( .A(n1640), .B(n1639), .Z(n1641) );
  AND U4492 ( .A(n1642), .B(n1641), .Z(n3854) );
  XNOR U4493 ( .A(oglobal[1]), .B(n3854), .Z(n3856) );
  NAND U4494 ( .A(n1644), .B(n1643), .Z(n1648) );
  NAND U4495 ( .A(n1646), .B(n1645), .Z(n1647) );
  AND U4496 ( .A(n1648), .B(n1647), .Z(n3855) );
  XOR U4497 ( .A(n3856), .B(n3855), .Z(n3845) );
  NANDN U4498 ( .A(n1650), .B(n1649), .Z(n1654) );
  NAND U4499 ( .A(n1652), .B(n1651), .Z(n1653) );
  AND U4500 ( .A(n1654), .B(n1653), .Z(n3843) );
  NANDN U4501 ( .A(n1656), .B(n1655), .Z(n1660) );
  NAND U4502 ( .A(n1658), .B(n1657), .Z(n1659) );
  NAND U4503 ( .A(n1660), .B(n1659), .Z(n3842) );
  XNOR U4504 ( .A(n3843), .B(n3842), .Z(n3844) );
  XNOR U4505 ( .A(n3845), .B(n3844), .Z(n3897) );
  XNOR U4506 ( .A(n3898), .B(n3897), .Z(n3871) );
  XNOR U4507 ( .A(n3872), .B(n3871), .Z(n3874) );
  XOR U4508 ( .A(n3873), .B(n3874), .Z(n3572) );
  NAND U4509 ( .A(n1662), .B(n1661), .Z(n1666) );
  NAND U4510 ( .A(n1664), .B(n1663), .Z(n1665) );
  AND U4511 ( .A(n1666), .B(n1665), .Z(n3848) );
  NANDN U4512 ( .A(n1668), .B(n1667), .Z(n1672) );
  NAND U4513 ( .A(n1670), .B(n1669), .Z(n1671) );
  NAND U4514 ( .A(n1672), .B(n1671), .Z(n3849) );
  XNOR U4515 ( .A(n3848), .B(n3849), .Z(n3851) );
  NANDN U4516 ( .A(n1674), .B(n1673), .Z(n1678) );
  NAND U4517 ( .A(n1676), .B(n1675), .Z(n1677) );
  AND U4518 ( .A(n1678), .B(n1677), .Z(n3850) );
  XOR U4519 ( .A(n3851), .B(n3850), .Z(n3928) );
  NANDN U4520 ( .A(n1680), .B(n1679), .Z(n1684) );
  NANDN U4521 ( .A(n1682), .B(n1681), .Z(n1683) );
  AND U4522 ( .A(n1684), .B(n1683), .Z(n3859) );
  NAND U4523 ( .A(n1686), .B(n1685), .Z(n1690) );
  NAND U4524 ( .A(n1688), .B(n1687), .Z(n1689) );
  NAND U4525 ( .A(n1690), .B(n1689), .Z(n3860) );
  XNOR U4526 ( .A(n3859), .B(n3860), .Z(n3862) );
  NANDN U4527 ( .A(n1692), .B(n1691), .Z(n1696) );
  NAND U4528 ( .A(n1694), .B(n1693), .Z(n1695) );
  AND U4529 ( .A(n1696), .B(n1695), .Z(n3861) );
  XOR U4530 ( .A(n3862), .B(n3861), .Z(n3926) );
  NANDN U4531 ( .A(n1698), .B(n1697), .Z(n1702) );
  NAND U4532 ( .A(n1700), .B(n1699), .Z(n1701) );
  NAND U4533 ( .A(n1702), .B(n1701), .Z(n3925) );
  XNOR U4534 ( .A(n3926), .B(n3925), .Z(n3927) );
  XOR U4535 ( .A(n3928), .B(n3927), .Z(n4201) );
  NANDN U4536 ( .A(n1704), .B(n1703), .Z(n1708) );
  NANDN U4537 ( .A(n1706), .B(n1705), .Z(n1707) );
  AND U4538 ( .A(n1708), .B(n1707), .Z(n4071) );
  NAND U4539 ( .A(n1710), .B(n1709), .Z(n1714) );
  NAND U4540 ( .A(n1712), .B(n1711), .Z(n1713) );
  AND U4541 ( .A(n1714), .B(n1713), .Z(n3434) );
  NAND U4542 ( .A(n1716), .B(n1715), .Z(n1720) );
  NAND U4543 ( .A(n1718), .B(n1717), .Z(n1719) );
  NAND U4544 ( .A(n1720), .B(n1719), .Z(n3435) );
  XNOR U4545 ( .A(n3434), .B(n3435), .Z(n3436) );
  NAND U4546 ( .A(n1722), .B(n1721), .Z(n1726) );
  NAND U4547 ( .A(n1724), .B(n1723), .Z(n1725) );
  NAND U4548 ( .A(n1726), .B(n1725), .Z(n3437) );
  XNOR U4549 ( .A(n3436), .B(n3437), .Z(n4070) );
  NANDN U4550 ( .A(n1728), .B(n1727), .Z(n1732) );
  NANDN U4551 ( .A(n1730), .B(n1729), .Z(n1731) );
  AND U4552 ( .A(n1732), .B(n1731), .Z(n4069) );
  XNOR U4553 ( .A(n4070), .B(n4069), .Z(n1733) );
  XNOR U4554 ( .A(n4071), .B(n1733), .Z(n4200) );
  NANDN U4555 ( .A(n1735), .B(n1734), .Z(n1739) );
  NANDN U4556 ( .A(n1737), .B(n1736), .Z(n1738) );
  AND U4557 ( .A(n1739), .B(n1738), .Z(n4643) );
  NANDN U4558 ( .A(n1741), .B(n1740), .Z(n1745) );
  NANDN U4559 ( .A(n1743), .B(n1742), .Z(n1744) );
  NAND U4560 ( .A(n1745), .B(n1744), .Z(n4641) );
  NAND U4561 ( .A(n1747), .B(n1746), .Z(n1751) );
  NAND U4562 ( .A(n1749), .B(n1748), .Z(n1750) );
  AND U4563 ( .A(n1751), .B(n1750), .Z(n4380) );
  NAND U4564 ( .A(n1753), .B(n1752), .Z(n1757) );
  NAND U4565 ( .A(n1755), .B(n1754), .Z(n1756) );
  AND U4566 ( .A(n1757), .B(n1756), .Z(n4381) );
  NAND U4567 ( .A(n1759), .B(n1758), .Z(n1763) );
  NAND U4568 ( .A(n1761), .B(n1760), .Z(n1762) );
  AND U4569 ( .A(n1763), .B(n1762), .Z(n4382) );
  XNOR U4570 ( .A(n4383), .B(n4382), .Z(n4642) );
  XNOR U4571 ( .A(n4641), .B(n4642), .Z(n1764) );
  XNOR U4572 ( .A(n4643), .B(n1764), .Z(n4199) );
  XOR U4573 ( .A(n4200), .B(n4199), .Z(n4202) );
  XOR U4574 ( .A(n4201), .B(n4202), .Z(n3571) );
  XOR U4575 ( .A(n3572), .B(n3571), .Z(n3573) );
  XOR U4576 ( .A(n3574), .B(n3573), .Z(n4027) );
  XOR U4577 ( .A(n4028), .B(n4027), .Z(n1765) );
  XNOR U4578 ( .A(n4029), .B(n1765), .Z(n3487) );
  NANDN U4579 ( .A(n1767), .B(n1766), .Z(n1771) );
  NAND U4580 ( .A(n1769), .B(n1768), .Z(n1770) );
  AND U4581 ( .A(n1771), .B(n1770), .Z(n3961) );
  NANDN U4582 ( .A(n1773), .B(n1772), .Z(n1777) );
  NAND U4583 ( .A(n1775), .B(n1774), .Z(n1776) );
  AND U4584 ( .A(n1777), .B(n1776), .Z(n3962) );
  NANDN U4585 ( .A(n1779), .B(n1778), .Z(n1783) );
  NAND U4586 ( .A(n1781), .B(n1780), .Z(n1782) );
  AND U4587 ( .A(n1783), .B(n1782), .Z(n3963) );
  XNOR U4588 ( .A(n3964), .B(n3963), .Z(n3297) );
  NANDN U4589 ( .A(n1785), .B(n1784), .Z(n1789) );
  NANDN U4590 ( .A(n1787), .B(n1786), .Z(n1788) );
  NAND U4591 ( .A(n1789), .B(n1788), .Z(n3295) );
  NANDN U4592 ( .A(n1791), .B(n1790), .Z(n1795) );
  NAND U4593 ( .A(n1793), .B(n1792), .Z(n1794) );
  AND U4594 ( .A(n1795), .B(n1794), .Z(n3955) );
  NANDN U4595 ( .A(n1797), .B(n1796), .Z(n1801) );
  NAND U4596 ( .A(n1799), .B(n1798), .Z(n1800) );
  AND U4597 ( .A(n1801), .B(n1800), .Z(n3956) );
  NANDN U4598 ( .A(n1803), .B(n1802), .Z(n1807) );
  NAND U4599 ( .A(n1805), .B(n1804), .Z(n1806) );
  AND U4600 ( .A(n1807), .B(n1806), .Z(n3957) );
  XNOR U4601 ( .A(n3958), .B(n3957), .Z(n3296) );
  XNOR U4602 ( .A(n3295), .B(n3296), .Z(n1808) );
  XNOR U4603 ( .A(n3297), .B(n1808), .Z(n3507) );
  NANDN U4604 ( .A(n1810), .B(n1809), .Z(n1814) );
  NAND U4605 ( .A(n1812), .B(n1811), .Z(n1813) );
  NAND U4606 ( .A(n1814), .B(n1813), .Z(n3506) );
  NANDN U4607 ( .A(n1816), .B(n1815), .Z(n1820) );
  NANDN U4608 ( .A(n1818), .B(n1817), .Z(n1819) );
  AND U4609 ( .A(n1820), .B(n1819), .Z(n4631) );
  NANDN U4610 ( .A(n1822), .B(n1821), .Z(n1826) );
  NANDN U4611 ( .A(n1824), .B(n1823), .Z(n1825) );
  AND U4612 ( .A(n1826), .B(n1825), .Z(n4630) );
  NAND U4613 ( .A(n1828), .B(n1827), .Z(n1832) );
  NAND U4614 ( .A(n1830), .B(n1829), .Z(n1831) );
  NAND U4615 ( .A(n1832), .B(n1831), .Z(n3309) );
  NAND U4616 ( .A(n1834), .B(n1833), .Z(n1838) );
  NAND U4617 ( .A(n1836), .B(n1835), .Z(n1837) );
  NAND U4618 ( .A(n1838), .B(n1837), .Z(n3308) );
  NAND U4619 ( .A(n1840), .B(n1839), .Z(n1844) );
  NAND U4620 ( .A(n1842), .B(n1841), .Z(n1843) );
  AND U4621 ( .A(n1844), .B(n1843), .Z(n3307) );
  XOR U4622 ( .A(n3308), .B(n3307), .Z(n1845) );
  XNOR U4623 ( .A(n3309), .B(n1845), .Z(n4629) );
  XNOR U4624 ( .A(n4630), .B(n4629), .Z(n1846) );
  XOR U4625 ( .A(n4631), .B(n1846), .Z(n3505) );
  XNOR U4626 ( .A(n3506), .B(n3505), .Z(n3508) );
  XNOR U4627 ( .A(n3507), .B(n3508), .Z(n3499) );
  NAND U4628 ( .A(n1848), .B(n1847), .Z(n1852) );
  NAND U4629 ( .A(n1850), .B(n1849), .Z(n1851) );
  NAND U4630 ( .A(n1852), .B(n1851), .Z(n3532) );
  NANDN U4631 ( .A(n1854), .B(n1853), .Z(n1858) );
  NAND U4632 ( .A(n1856), .B(n1855), .Z(n1857) );
  NAND U4633 ( .A(n1858), .B(n1857), .Z(n3530) );
  NANDN U4634 ( .A(n1860), .B(n1859), .Z(n1864) );
  NANDN U4635 ( .A(n1862), .B(n1861), .Z(n1863) );
  NAND U4636 ( .A(n1864), .B(n1863), .Z(n3742) );
  NANDN U4637 ( .A(n1866), .B(n1865), .Z(n1870) );
  NAND U4638 ( .A(n1868), .B(n1867), .Z(n1869) );
  AND U4639 ( .A(n1870), .B(n1869), .Z(n4416) );
  NANDN U4640 ( .A(n1872), .B(n1871), .Z(n1876) );
  NAND U4641 ( .A(n1874), .B(n1873), .Z(n1875) );
  AND U4642 ( .A(n1876), .B(n1875), .Z(n4417) );
  NANDN U4643 ( .A(n1878), .B(n1877), .Z(n1882) );
  NAND U4644 ( .A(n1880), .B(n1879), .Z(n1881) );
  AND U4645 ( .A(n1882), .B(n1881), .Z(n4419) );
  IV U4646 ( .A(n3738), .Z(n3741) );
  NANDN U4647 ( .A(n1884), .B(n1883), .Z(n1888) );
  NANDN U4648 ( .A(n1886), .B(n1885), .Z(n1887) );
  NAND U4649 ( .A(n1888), .B(n1887), .Z(n3740) );
  IV U4650 ( .A(n3740), .Z(n3739) );
  XNOR U4651 ( .A(n3499), .B(n3500), .Z(n3502) );
  NANDN U4652 ( .A(n1890), .B(n1889), .Z(n1894) );
  NAND U4653 ( .A(n1892), .B(n1891), .Z(n1893) );
  NAND U4654 ( .A(n1894), .B(n1893), .Z(n3538) );
  NANDN U4655 ( .A(n1896), .B(n1895), .Z(n1900) );
  NANDN U4656 ( .A(n1898), .B(n1897), .Z(n1899) );
  AND U4657 ( .A(n1900), .B(n1899), .Z(n4473) );
  NANDN U4658 ( .A(n1902), .B(n1901), .Z(n1906) );
  NAND U4659 ( .A(n1904), .B(n1903), .Z(n1905) );
  AND U4660 ( .A(n1906), .B(n1905), .Z(n4392) );
  NANDN U4661 ( .A(n1908), .B(n1907), .Z(n1912) );
  NAND U4662 ( .A(n1910), .B(n1909), .Z(n1911) );
  AND U4663 ( .A(n1912), .B(n1911), .Z(n4393) );
  NAND U4664 ( .A(n1914), .B(n1913), .Z(n1918) );
  NAND U4665 ( .A(n1916), .B(n1915), .Z(n1917) );
  AND U4666 ( .A(n1918), .B(n1917), .Z(n4394) );
  XNOR U4667 ( .A(n4395), .B(n4394), .Z(n4471) );
  NANDN U4668 ( .A(n1920), .B(n1919), .Z(n1924) );
  NANDN U4669 ( .A(n1922), .B(n1921), .Z(n1923) );
  AND U4670 ( .A(n1924), .B(n1923), .Z(n4470) );
  XNOR U4671 ( .A(n4473), .B(n4472), .Z(n3536) );
  XNOR U4672 ( .A(n3502), .B(n3501), .Z(n4024) );
  NAND U4673 ( .A(n1930), .B(n1929), .Z(n1934) );
  NAND U4674 ( .A(n1932), .B(n1931), .Z(n1933) );
  AND U4675 ( .A(n1934), .B(n1933), .Z(n3544) );
  NANDN U4676 ( .A(n1936), .B(n1935), .Z(n1940) );
  NANDN U4677 ( .A(n1938), .B(n1937), .Z(n1939) );
  AND U4678 ( .A(n1940), .B(n1939), .Z(n4455) );
  NAND U4679 ( .A(n1942), .B(n1941), .Z(n1946) );
  NAND U4680 ( .A(n1944), .B(n1943), .Z(n1945) );
  NAND U4681 ( .A(n1946), .B(n1945), .Z(n3306) );
  NANDN U4682 ( .A(n1948), .B(n1947), .Z(n1952) );
  NAND U4683 ( .A(n1950), .B(n1949), .Z(n1951) );
  NAND U4684 ( .A(n1952), .B(n1951), .Z(n3305) );
  NAND U4685 ( .A(n1954), .B(n1953), .Z(n1958) );
  NAND U4686 ( .A(n1956), .B(n1955), .Z(n1957) );
  AND U4687 ( .A(n1958), .B(n1957), .Z(n3304) );
  XOR U4688 ( .A(n3305), .B(n3304), .Z(n1959) );
  XNOR U4689 ( .A(n3306), .B(n1959), .Z(n4453) );
  NAND U4690 ( .A(n1961), .B(n1960), .Z(n1965) );
  NANDN U4691 ( .A(n1963), .B(n1962), .Z(n1964) );
  AND U4692 ( .A(n1965), .B(n1964), .Z(n4452) );
  XOR U4693 ( .A(n4455), .B(n4454), .Z(n3542) );
  XNOR U4694 ( .A(n3542), .B(n3541), .Z(n3543) );
  XNOR U4695 ( .A(n3544), .B(n3543), .Z(n3475) );
  NANDN U4696 ( .A(n1971), .B(n1970), .Z(n1975) );
  NANDN U4697 ( .A(n1973), .B(n1972), .Z(n1974) );
  AND U4698 ( .A(n1975), .B(n1974), .Z(n3550) );
  NANDN U4699 ( .A(n1977), .B(n1976), .Z(n1981) );
  NANDN U4700 ( .A(n1979), .B(n1978), .Z(n1980) );
  AND U4701 ( .A(n1981), .B(n1980), .Z(n4437) );
  NAND U4702 ( .A(n1983), .B(n1982), .Z(n1987) );
  NAND U4703 ( .A(n1985), .B(n1984), .Z(n1986) );
  NAND U4704 ( .A(n1987), .B(n1986), .Z(n4189) );
  NANDN U4705 ( .A(n1989), .B(n1988), .Z(n1993) );
  NAND U4706 ( .A(n1991), .B(n1990), .Z(n1992) );
  NAND U4707 ( .A(n1993), .B(n1992), .Z(n4188) );
  NAND U4708 ( .A(n1995), .B(n1994), .Z(n1999) );
  NAND U4709 ( .A(n1997), .B(n1996), .Z(n1998) );
  AND U4710 ( .A(n1999), .B(n1998), .Z(n4187) );
  XOR U4711 ( .A(n4188), .B(n4187), .Z(n2000) );
  XNOR U4712 ( .A(n4189), .B(n2000), .Z(n4435) );
  NAND U4713 ( .A(n2002), .B(n2001), .Z(n2006) );
  NAND U4714 ( .A(n2004), .B(n2003), .Z(n2005) );
  AND U4715 ( .A(n2006), .B(n2005), .Z(n4434) );
  XOR U4716 ( .A(n4437), .B(n4436), .Z(n3548) );
  NANDN U4717 ( .A(n2008), .B(n2007), .Z(n2012) );
  NAND U4718 ( .A(n2010), .B(n2009), .Z(n2011) );
  NAND U4719 ( .A(n2012), .B(n2011), .Z(n3547) );
  XNOR U4720 ( .A(n3548), .B(n3547), .Z(n3549) );
  XOR U4721 ( .A(n3550), .B(n3549), .Z(n3476) );
  XNOR U4722 ( .A(n3475), .B(n3476), .Z(n3478) );
  NANDN U4723 ( .A(n2022), .B(n2021), .Z(n2026) );
  NANDN U4724 ( .A(n2024), .B(n2023), .Z(n2025) );
  NAND U4725 ( .A(n2026), .B(n2025), .Z(n4613) );
  NAND U4726 ( .A(n2028), .B(n2027), .Z(n2032) );
  NAND U4727 ( .A(n2030), .B(n2029), .Z(n2031) );
  AND U4728 ( .A(n2032), .B(n2031), .Z(n4362) );
  NAND U4729 ( .A(n2034), .B(n2033), .Z(n2038) );
  NAND U4730 ( .A(n2036), .B(n2035), .Z(n2037) );
  AND U4731 ( .A(n2038), .B(n2037), .Z(n4363) );
  NAND U4732 ( .A(n2040), .B(n2039), .Z(n2044) );
  NAND U4733 ( .A(n2042), .B(n2041), .Z(n2043) );
  AND U4734 ( .A(n2044), .B(n2043), .Z(n4365) );
  IV U4735 ( .A(n4609), .Z(n4612) );
  NAND U4736 ( .A(n2046), .B(n2045), .Z(n2050) );
  NAND U4737 ( .A(n2048), .B(n2047), .Z(n2049) );
  NAND U4738 ( .A(n2050), .B(n2049), .Z(n4611) );
  IV U4739 ( .A(n4611), .Z(n4610) );
  XNOR U4740 ( .A(n3478), .B(n3477), .Z(n4022) );
  NANDN U4741 ( .A(n2052), .B(n2051), .Z(n2056) );
  NANDN U4742 ( .A(n2054), .B(n2053), .Z(n2055) );
  NAND U4743 ( .A(n2056), .B(n2055), .Z(n3641) );
  NANDN U4744 ( .A(n2058), .B(n2057), .Z(n2062) );
  NANDN U4745 ( .A(n2060), .B(n2059), .Z(n2061) );
  AND U4746 ( .A(n2062), .B(n2061), .Z(n3372) );
  NANDN U4747 ( .A(n2064), .B(n2063), .Z(n2068) );
  NAND U4748 ( .A(n2066), .B(n2065), .Z(n2067) );
  AND U4749 ( .A(n2068), .B(n2067), .Z(n4326) );
  NANDN U4750 ( .A(n2070), .B(n2069), .Z(n2074) );
  NAND U4751 ( .A(n2072), .B(n2071), .Z(n2073) );
  NAND U4752 ( .A(n2074), .B(n2073), .Z(n4327) );
  XNOR U4753 ( .A(n4326), .B(n4327), .Z(n4329) );
  NANDN U4754 ( .A(n2076), .B(n2075), .Z(n2080) );
  NAND U4755 ( .A(n2078), .B(n2077), .Z(n2079) );
  AND U4756 ( .A(n2080), .B(n2079), .Z(n4328) );
  XOR U4757 ( .A(n4329), .B(n4328), .Z(n3370) );
  NANDN U4758 ( .A(n2082), .B(n2081), .Z(n2086) );
  NANDN U4759 ( .A(n2084), .B(n2083), .Z(n2085) );
  AND U4760 ( .A(n2086), .B(n2085), .Z(n3369) );
  XNOR U4761 ( .A(n3370), .B(n3369), .Z(n3371) );
  XNOR U4762 ( .A(n3372), .B(n3371), .Z(n3639) );
  NANDN U4763 ( .A(n2088), .B(n2087), .Z(n2092) );
  NAND U4764 ( .A(n2090), .B(n2089), .Z(n2091) );
  NAND U4765 ( .A(n2092), .B(n2091), .Z(n3638) );
  XOR U4766 ( .A(n3641), .B(n3640), .Z(n3403) );
  NANDN U4767 ( .A(n2094), .B(n2093), .Z(n2098) );
  NANDN U4768 ( .A(n2096), .B(n2095), .Z(n2097) );
  AND U4769 ( .A(n2098), .B(n2097), .Z(n3526) );
  NANDN U4770 ( .A(n2100), .B(n2099), .Z(n2104) );
  NANDN U4771 ( .A(n2102), .B(n2101), .Z(n2103) );
  AND U4772 ( .A(n2104), .B(n2103), .Z(n4491) );
  NANDN U4773 ( .A(n2106), .B(n2105), .Z(n2110) );
  NAND U4774 ( .A(n2108), .B(n2107), .Z(n2109) );
  AND U4775 ( .A(n2110), .B(n2109), .Z(n4314) );
  NANDN U4776 ( .A(n2112), .B(n2111), .Z(n2116) );
  NAND U4777 ( .A(n2114), .B(n2113), .Z(n2115) );
  AND U4778 ( .A(n2116), .B(n2115), .Z(n4315) );
  NANDN U4779 ( .A(n2118), .B(n2117), .Z(n2122) );
  NAND U4780 ( .A(n2120), .B(n2119), .Z(n2121) );
  AND U4781 ( .A(n2122), .B(n2121), .Z(n4316) );
  XNOR U4782 ( .A(n4317), .B(n4316), .Z(n4489) );
  NANDN U4783 ( .A(n2124), .B(n2123), .Z(n2128) );
  NANDN U4784 ( .A(n2126), .B(n2125), .Z(n2127) );
  AND U4785 ( .A(n2128), .B(n2127), .Z(n4488) );
  XOR U4786 ( .A(n4491), .B(n4490), .Z(n3524) );
  NANDN U4787 ( .A(n2130), .B(n2129), .Z(n2134) );
  NANDN U4788 ( .A(n2132), .B(n2131), .Z(n2133) );
  NAND U4789 ( .A(n2134), .B(n2133), .Z(n3523) );
  XNOR U4790 ( .A(n3524), .B(n3523), .Z(n3525) );
  XOR U4791 ( .A(n3526), .B(n3525), .Z(n3405) );
  NANDN U4792 ( .A(n2140), .B(n2139), .Z(n2144) );
  NAND U4793 ( .A(n2142), .B(n2141), .Z(n2143) );
  NAND U4794 ( .A(n2144), .B(n2143), .Z(n3645) );
  NAND U4795 ( .A(n2146), .B(n2145), .Z(n2150) );
  NAND U4796 ( .A(n2148), .B(n2147), .Z(n2149) );
  AND U4797 ( .A(n2150), .B(n2149), .Z(n4595) );
  NANDN U4798 ( .A(n2152), .B(n2151), .Z(n2156) );
  NANDN U4799 ( .A(n2154), .B(n2153), .Z(n2155) );
  NAND U4800 ( .A(n2156), .B(n2155), .Z(n4593) );
  NAND U4801 ( .A(n2158), .B(n2157), .Z(n2162) );
  NAND U4802 ( .A(n2160), .B(n2159), .Z(n2161) );
  AND U4803 ( .A(n2162), .B(n2161), .Z(n4356) );
  NANDN U4804 ( .A(n2164), .B(n2163), .Z(n2168) );
  NAND U4805 ( .A(n2166), .B(n2165), .Z(n2167) );
  NAND U4806 ( .A(n2168), .B(n2167), .Z(n4357) );
  XNOR U4807 ( .A(n4356), .B(n4357), .Z(n4359) );
  NANDN U4808 ( .A(n2170), .B(n2169), .Z(n2174) );
  NAND U4809 ( .A(n2172), .B(n2171), .Z(n2173) );
  AND U4810 ( .A(n2174), .B(n2173), .Z(n4358) );
  XNOR U4811 ( .A(n4359), .B(n4358), .Z(n4594) );
  XNOR U4812 ( .A(n4593), .B(n4594), .Z(n2175) );
  XNOR U4813 ( .A(n4595), .B(n2175), .Z(n3644) );
  XNOR U4814 ( .A(n3405), .B(n3404), .Z(n2176) );
  XOR U4815 ( .A(n3403), .B(n2176), .Z(n4021) );
  XOR U4816 ( .A(n3487), .B(n3488), .Z(n3490) );
  XOR U4817 ( .A(n3489), .B(n3490), .Z(n3495) );
  NANDN U4818 ( .A(n2178), .B(n2177), .Z(n2182) );
  OR U4819 ( .A(n2180), .B(n2179), .Z(n2181) );
  NAND U4820 ( .A(n2182), .B(n2181), .Z(n4046) );
  IV U4821 ( .A(n4046), .Z(n4044) );
  NAND U4822 ( .A(n2184), .B(n2183), .Z(n2188) );
  NAND U4823 ( .A(n2186), .B(n2185), .Z(n2187) );
  AND U4824 ( .A(n2188), .B(n2187), .Z(n3608) );
  NAND U4825 ( .A(n2190), .B(n2189), .Z(n2194) );
  NAND U4826 ( .A(n2192), .B(n2191), .Z(n2193) );
  AND U4827 ( .A(n2194), .B(n2193), .Z(n3609) );
  NAND U4828 ( .A(n2196), .B(n2195), .Z(n2200) );
  NAND U4829 ( .A(n2198), .B(n2197), .Z(n2199) );
  AND U4830 ( .A(n2200), .B(n2199), .Z(n3610) );
  XOR U4831 ( .A(n3611), .B(n3610), .Z(n4623) );
  NAND U4832 ( .A(n2202), .B(n2201), .Z(n2206) );
  NAND U4833 ( .A(n2204), .B(n2203), .Z(n2205) );
  AND U4834 ( .A(n2206), .B(n2205), .Z(n4530) );
  NAND U4835 ( .A(n2208), .B(n2207), .Z(n2212) );
  NAND U4836 ( .A(n2210), .B(n2209), .Z(n2211) );
  AND U4837 ( .A(n2212), .B(n2211), .Z(n4531) );
  NAND U4838 ( .A(n2214), .B(n2213), .Z(n2218) );
  NAND U4839 ( .A(n2216), .B(n2215), .Z(n2217) );
  AND U4840 ( .A(n2218), .B(n2217), .Z(n4532) );
  XOR U4841 ( .A(n4533), .B(n4532), .Z(n4621) );
  NAND U4842 ( .A(n2220), .B(n2219), .Z(n2224) );
  NAND U4843 ( .A(n2222), .B(n2221), .Z(n2223) );
  AND U4844 ( .A(n2224), .B(n2223), .Z(n4566) );
  NAND U4845 ( .A(n2226), .B(n2225), .Z(n2230) );
  NAND U4846 ( .A(n2228), .B(n2227), .Z(n2229) );
  AND U4847 ( .A(n2230), .B(n2229), .Z(n4567) );
  NAND U4848 ( .A(n2232), .B(n2231), .Z(n2236) );
  NAND U4849 ( .A(n2234), .B(n2233), .Z(n2235) );
  AND U4850 ( .A(n2236), .B(n2235), .Z(n4568) );
  XNOR U4851 ( .A(n4569), .B(n4568), .Z(n4620) );
  XNOR U4852 ( .A(n4621), .B(n4620), .Z(n4622) );
  XOR U4853 ( .A(n4623), .B(n4622), .Z(n4619) );
  NANDN U4854 ( .A(n2238), .B(n2237), .Z(n2242) );
  NAND U4855 ( .A(n2240), .B(n2239), .Z(n2241) );
  AND U4856 ( .A(n2242), .B(n2241), .Z(n4009) );
  NAND U4857 ( .A(n2244), .B(n2243), .Z(n2248) );
  NAND U4858 ( .A(n2246), .B(n2245), .Z(n2247) );
  AND U4859 ( .A(n2248), .B(n2247), .Z(n4010) );
  NAND U4860 ( .A(n2250), .B(n2249), .Z(n2254) );
  NAND U4861 ( .A(n2252), .B(n2251), .Z(n2253) );
  AND U4862 ( .A(n2254), .B(n2253), .Z(n4011) );
  XNOR U4863 ( .A(n4012), .B(n4011), .Z(n4628) );
  NAND U4864 ( .A(n2256), .B(n2255), .Z(n2260) );
  NAND U4865 ( .A(n2258), .B(n2257), .Z(n2259) );
  NAND U4866 ( .A(n2260), .B(n2259), .Z(n4626) );
  NAND U4867 ( .A(n2262), .B(n2261), .Z(n2266) );
  NAND U4868 ( .A(n2264), .B(n2263), .Z(n2265) );
  AND U4869 ( .A(n2266), .B(n2265), .Z(n4560) );
  NAND U4870 ( .A(n2268), .B(n2267), .Z(n2272) );
  NAND U4871 ( .A(n2270), .B(n2269), .Z(n2271) );
  AND U4872 ( .A(n2272), .B(n2271), .Z(n4561) );
  NAND U4873 ( .A(n2274), .B(n2273), .Z(n2278) );
  NAND U4874 ( .A(n2276), .B(n2275), .Z(n2277) );
  AND U4875 ( .A(n2278), .B(n2277), .Z(n4562) );
  XNOR U4876 ( .A(n4563), .B(n4562), .Z(n4627) );
  XNOR U4877 ( .A(n4626), .B(n4627), .Z(n2279) );
  XOR U4878 ( .A(n4628), .B(n2279), .Z(n4617) );
  NAND U4879 ( .A(n2281), .B(n2280), .Z(n2285) );
  NAND U4880 ( .A(n2283), .B(n2282), .Z(n2284) );
  AND U4881 ( .A(n2285), .B(n2284), .Z(n3585) );
  NANDN U4882 ( .A(n2287), .B(n2286), .Z(n2291) );
  NAND U4883 ( .A(n2289), .B(n2288), .Z(n2290) );
  AND U4884 ( .A(n2291), .B(n2290), .Z(n3584) );
  NAND U4885 ( .A(n2293), .B(n2292), .Z(n2297) );
  NAND U4886 ( .A(n2295), .B(n2294), .Z(n2296) );
  AND U4887 ( .A(n2297), .B(n2296), .Z(n3583) );
  NANDN U4888 ( .A(n2299), .B(n2298), .Z(n2303) );
  NAND U4889 ( .A(n2301), .B(n2300), .Z(n2302) );
  AND U4890 ( .A(n2303), .B(n2302), .Z(n3937) );
  NAND U4891 ( .A(n2305), .B(n2304), .Z(n2309) );
  NAND U4892 ( .A(n2307), .B(n2306), .Z(n2308) );
  AND U4893 ( .A(n2309), .B(n2308), .Z(n3938) );
  NAND U4894 ( .A(n2311), .B(n2310), .Z(n2315) );
  NAND U4895 ( .A(n2313), .B(n2312), .Z(n2314) );
  AND U4896 ( .A(n2315), .B(n2314), .Z(n3939) );
  XOR U4897 ( .A(n3940), .B(n3939), .Z(n4633) );
  NAND U4898 ( .A(n2317), .B(n2316), .Z(n2321) );
  NAND U4899 ( .A(n2319), .B(n2318), .Z(n2320) );
  NAND U4900 ( .A(n2321), .B(n2320), .Z(n3350) );
  NAND U4901 ( .A(n2323), .B(n2322), .Z(n2327) );
  NAND U4902 ( .A(n2325), .B(n2324), .Z(n2326) );
  NAND U4903 ( .A(n2327), .B(n2326), .Z(n3349) );
  NAND U4904 ( .A(n2329), .B(n2328), .Z(n2333) );
  NAND U4905 ( .A(n2331), .B(n2330), .Z(n2332) );
  AND U4906 ( .A(n2333), .B(n2332), .Z(n3348) );
  XOR U4907 ( .A(n3349), .B(n3348), .Z(n2334) );
  XNOR U4908 ( .A(n3350), .B(n2334), .Z(n4632) );
  XNOR U4909 ( .A(n4633), .B(n4632), .Z(n4635) );
  XOR U4910 ( .A(n4634), .B(n4635), .Z(n4618) );
  NANDN U4911 ( .A(n2336), .B(n2335), .Z(n2340) );
  OR U4912 ( .A(n2338), .B(n2337), .Z(n2339) );
  AND U4913 ( .A(n2340), .B(n2339), .Z(n3417) );
  XOR U4914 ( .A(n3416), .B(n3417), .Z(n3419) );
  NANDN U4915 ( .A(n2346), .B(n2345), .Z(n2350) );
  NANDN U4916 ( .A(n2348), .B(n2347), .Z(n2349) );
  NAND U4917 ( .A(n2350), .B(n2349), .Z(n4279) );
  NANDN U4918 ( .A(n2352), .B(n2351), .Z(n2356) );
  NANDN U4919 ( .A(n2354), .B(n2353), .Z(n2355) );
  AND U4920 ( .A(n2356), .B(n2355), .Z(n3462) );
  NANDN U4921 ( .A(n2358), .B(n2357), .Z(n2362) );
  NANDN U4922 ( .A(n2360), .B(n2359), .Z(n2361) );
  NAND U4923 ( .A(n2362), .B(n2361), .Z(n3463) );
  XNOR U4924 ( .A(n3462), .B(n3463), .Z(n3465) );
  NANDN U4925 ( .A(n2364), .B(n2363), .Z(n2368) );
  NANDN U4926 ( .A(n2366), .B(n2365), .Z(n2367) );
  AND U4927 ( .A(n2368), .B(n2367), .Z(n3464) );
  XNOR U4928 ( .A(n3465), .B(n3464), .Z(n4278) );
  XOR U4929 ( .A(n3419), .B(n3418), .Z(n4047) );
  NANDN U4930 ( .A(n2370), .B(n2369), .Z(n2374) );
  NAND U4931 ( .A(n2372), .B(n2371), .Z(n2373) );
  AND U4932 ( .A(n2374), .B(n2373), .Z(n4266) );
  NANDN U4933 ( .A(n2376), .B(n2375), .Z(n2380) );
  NAND U4934 ( .A(n2378), .B(n2377), .Z(n2379) );
  AND U4935 ( .A(n2380), .B(n2379), .Z(n4267) );
  NANDN U4936 ( .A(n2382), .B(n2381), .Z(n2386) );
  NAND U4937 ( .A(n2384), .B(n2383), .Z(n2385) );
  AND U4938 ( .A(n2386), .B(n2385), .Z(n4269) );
  NAND U4939 ( .A(n2388), .B(n2387), .Z(n2392) );
  NAND U4940 ( .A(n2390), .B(n2389), .Z(n2391) );
  AND U4941 ( .A(n2392), .B(n2391), .Z(n3877) );
  NANDN U4942 ( .A(n2394), .B(n2393), .Z(n2398) );
  NAND U4943 ( .A(n2396), .B(n2395), .Z(n2397) );
  AND U4944 ( .A(n2398), .B(n2397), .Z(n3878) );
  NAND U4945 ( .A(n2400), .B(n2399), .Z(n2404) );
  NAND U4946 ( .A(n2402), .B(n2401), .Z(n2403) );
  AND U4947 ( .A(n2404), .B(n2403), .Z(n3880) );
  XNOR U4948 ( .A(n3879), .B(n3880), .Z(n4638) );
  NANDN U4949 ( .A(n2406), .B(n2405), .Z(n2410) );
  NAND U4950 ( .A(n2408), .B(n2407), .Z(n2409) );
  AND U4951 ( .A(n2410), .B(n2409), .Z(n4235) );
  NAND U4952 ( .A(n2412), .B(n2411), .Z(n2416) );
  NAND U4953 ( .A(n2414), .B(n2413), .Z(n2415) );
  AND U4954 ( .A(n2416), .B(n2415), .Z(n4236) );
  NANDN U4955 ( .A(n2418), .B(n2417), .Z(n2422) );
  NAND U4956 ( .A(n2420), .B(n2419), .Z(n2421) );
  AND U4957 ( .A(n2422), .B(n2421), .Z(n4238) );
  XOR U4958 ( .A(n4638), .B(n4639), .Z(n2423) );
  XNOR U4959 ( .A(n4640), .B(n2423), .Z(n3280) );
  NAND U4960 ( .A(n2425), .B(n2424), .Z(n2429) );
  NAND U4961 ( .A(n2427), .B(n2426), .Z(n2428) );
  AND U4962 ( .A(n2429), .B(n2428), .Z(n3339) );
  NANDN U4963 ( .A(n2431), .B(n2430), .Z(n2435) );
  NAND U4964 ( .A(n2433), .B(n2432), .Z(n2434) );
  AND U4965 ( .A(n2435), .B(n2434), .Z(n3340) );
  NAND U4966 ( .A(n2437), .B(n2436), .Z(n2441) );
  NAND U4967 ( .A(n2439), .B(n2438), .Z(n2440) );
  AND U4968 ( .A(n2441), .B(n2440), .Z(n3341) );
  XOR U4969 ( .A(n3342), .B(n3341), .Z(n4659) );
  NAND U4970 ( .A(n2443), .B(n2442), .Z(n2447) );
  NAND U4971 ( .A(n2445), .B(n2444), .Z(n2446) );
  AND U4972 ( .A(n2447), .B(n2446), .Z(n4542) );
  NANDN U4973 ( .A(n2449), .B(n2448), .Z(n2453) );
  NAND U4974 ( .A(n2451), .B(n2450), .Z(n2452) );
  AND U4975 ( .A(n2453), .B(n2452), .Z(n4543) );
  NAND U4976 ( .A(n2455), .B(n2454), .Z(n2459) );
  NAND U4977 ( .A(n2457), .B(n2456), .Z(n2458) );
  AND U4978 ( .A(n2459), .B(n2458), .Z(n4544) );
  XOR U4979 ( .A(n4545), .B(n4544), .Z(n4657) );
  NAND U4980 ( .A(n2461), .B(n2460), .Z(n2465) );
  NAND U4981 ( .A(n2463), .B(n2462), .Z(n2464) );
  AND U4982 ( .A(n2465), .B(n2464), .Z(n3325) );
  NAND U4983 ( .A(n2467), .B(n2466), .Z(n2471) );
  NAND U4984 ( .A(n2469), .B(n2468), .Z(n2470) );
  AND U4985 ( .A(n2471), .B(n2470), .Z(n3326) );
  NANDN U4986 ( .A(n2473), .B(n2472), .Z(n2477) );
  NAND U4987 ( .A(n2475), .B(n2474), .Z(n2476) );
  AND U4988 ( .A(n2477), .B(n2476), .Z(n3327) );
  XNOR U4989 ( .A(n3328), .B(n3327), .Z(n4656) );
  XNOR U4990 ( .A(n4657), .B(n4656), .Z(n4658) );
  XNOR U4991 ( .A(n4659), .B(n4658), .Z(n3278) );
  NANDN U4992 ( .A(n2479), .B(n2478), .Z(n2483) );
  NAND U4993 ( .A(n2481), .B(n2480), .Z(n2482) );
  AND U4994 ( .A(n2483), .B(n2482), .Z(n4223) );
  NAND U4995 ( .A(n2485), .B(n2484), .Z(n2489) );
  NAND U4996 ( .A(n2487), .B(n2486), .Z(n2488) );
  AND U4997 ( .A(n2489), .B(n2488), .Z(n4224) );
  NAND U4998 ( .A(n2491), .B(n2490), .Z(n2495) );
  NAND U4999 ( .A(n2493), .B(n2492), .Z(n2494) );
  AND U5000 ( .A(n2495), .B(n2494), .Z(n4225) );
  XOR U5001 ( .A(n4226), .B(n4225), .Z(n4647) );
  NAND U5002 ( .A(n2497), .B(n2496), .Z(n2501) );
  NAND U5003 ( .A(n2499), .B(n2498), .Z(n2500) );
  AND U5004 ( .A(n2501), .B(n2500), .Z(n3883) );
  NAND U5005 ( .A(n2503), .B(n2502), .Z(n2507) );
  NAND U5006 ( .A(n2505), .B(n2504), .Z(n2506) );
  AND U5007 ( .A(n2507), .B(n2506), .Z(n3884) );
  NANDN U5008 ( .A(n2509), .B(n2508), .Z(n2513) );
  NAND U5009 ( .A(n2511), .B(n2510), .Z(n2512) );
  AND U5010 ( .A(n2513), .B(n2512), .Z(n3885) );
  XOR U5011 ( .A(n3886), .B(n3885), .Z(n4645) );
  NAND U5012 ( .A(n2515), .B(n2514), .Z(n2519) );
  NAND U5013 ( .A(n2517), .B(n2516), .Z(n2518) );
  AND U5014 ( .A(n2519), .B(n2518), .Z(n4644) );
  XNOR U5015 ( .A(n4645), .B(n4644), .Z(n4646) );
  XOR U5016 ( .A(n4647), .B(n4646), .Z(n3277) );
  XNOR U5017 ( .A(n3278), .B(n3277), .Z(n3279) );
  XOR U5018 ( .A(n3280), .B(n3279), .Z(n3765) );
  NAND U5019 ( .A(n2521), .B(n2520), .Z(n2525) );
  NAND U5020 ( .A(n2523), .B(n2522), .Z(n2524) );
  AND U5021 ( .A(n2525), .B(n2524), .Z(n4003) );
  NAND U5022 ( .A(n2527), .B(n2526), .Z(n2531) );
  NAND U5023 ( .A(n2529), .B(n2528), .Z(n2530) );
  AND U5024 ( .A(n2531), .B(n2530), .Z(n4004) );
  NAND U5025 ( .A(n2533), .B(n2532), .Z(n2537) );
  NAND U5026 ( .A(n2535), .B(n2534), .Z(n2536) );
  AND U5027 ( .A(n2537), .B(n2536), .Z(n4005) );
  XOR U5028 ( .A(n4006), .B(n4005), .Z(n3683) );
  NANDN U5029 ( .A(n2539), .B(n2538), .Z(n2543) );
  NANDN U5030 ( .A(n2541), .B(n2540), .Z(n2542) );
  AND U5031 ( .A(n2543), .B(n2542), .Z(n3680) );
  NAND U5032 ( .A(n2545), .B(n2544), .Z(n2549) );
  NAND U5033 ( .A(n2547), .B(n2546), .Z(n2548) );
  NAND U5034 ( .A(n2549), .B(n2548), .Z(n3681) );
  XNOR U5035 ( .A(n3680), .B(n3681), .Z(n3682) );
  XNOR U5036 ( .A(n3683), .B(n3682), .Z(n3425) );
  NANDN U5037 ( .A(n2551), .B(n2550), .Z(n2555) );
  NANDN U5038 ( .A(n2553), .B(n2552), .Z(n2554) );
  AND U5039 ( .A(n2555), .B(n2554), .Z(n3696) );
  NANDN U5040 ( .A(n2557), .B(n2556), .Z(n2561) );
  NANDN U5041 ( .A(n2559), .B(n2558), .Z(n2560) );
  AND U5042 ( .A(n2561), .B(n2560), .Z(n3693) );
  NANDN U5043 ( .A(n2563), .B(n2562), .Z(n2567) );
  NANDN U5044 ( .A(n2565), .B(n2564), .Z(n2566) );
  NAND U5045 ( .A(n2567), .B(n2566), .Z(n3694) );
  XNOR U5046 ( .A(n3693), .B(n3694), .Z(n3695) );
  XOR U5047 ( .A(n3696), .B(n3695), .Z(n3423) );
  NAND U5048 ( .A(n2569), .B(n2568), .Z(n2573) );
  NAND U5049 ( .A(n2571), .B(n2570), .Z(n2572) );
  NAND U5050 ( .A(n2573), .B(n2572), .Z(n3688) );
  NAND U5051 ( .A(n2575), .B(n2574), .Z(n2579) );
  NAND U5052 ( .A(n2577), .B(n2576), .Z(n2578) );
  NAND U5053 ( .A(n2579), .B(n2578), .Z(n3687) );
  NANDN U5054 ( .A(n2581), .B(n2580), .Z(n2585) );
  NANDN U5055 ( .A(n2583), .B(n2582), .Z(n2584) );
  AND U5056 ( .A(n2585), .B(n2584), .Z(n3686) );
  XOR U5057 ( .A(n3687), .B(n3686), .Z(n2586) );
  XNOR U5058 ( .A(n3688), .B(n2586), .Z(n3422) );
  XNOR U5059 ( .A(n3423), .B(n3422), .Z(n3424) );
  XOR U5060 ( .A(n3425), .B(n3424), .Z(n3767) );
  NAND U5061 ( .A(n2592), .B(n2591), .Z(n2596) );
  NAND U5062 ( .A(n2594), .B(n2593), .Z(n2595) );
  NAND U5063 ( .A(n2596), .B(n2595), .Z(n3473) );
  NANDN U5064 ( .A(n2598), .B(n2597), .Z(n2602) );
  NANDN U5065 ( .A(n2600), .B(n2599), .Z(n2601) );
  NAND U5066 ( .A(n2602), .B(n2601), .Z(n3472) );
  NANDN U5067 ( .A(n2604), .B(n2603), .Z(n2608) );
  NANDN U5068 ( .A(n2606), .B(n2605), .Z(n2607) );
  AND U5069 ( .A(n2608), .B(n2607), .Z(n3471) );
  XOR U5070 ( .A(n3472), .B(n3471), .Z(n2609) );
  XOR U5071 ( .A(n3473), .B(n2609), .Z(n3706) );
  NANDN U5072 ( .A(n2611), .B(n2610), .Z(n2615) );
  NANDN U5073 ( .A(n2613), .B(n2612), .Z(n2614) );
  NAND U5074 ( .A(n2615), .B(n2614), .Z(n3701) );
  NANDN U5075 ( .A(n2617), .B(n2616), .Z(n2621) );
  NANDN U5076 ( .A(n2619), .B(n2618), .Z(n2620) );
  NAND U5077 ( .A(n2621), .B(n2620), .Z(n3700) );
  NANDN U5078 ( .A(n2623), .B(n2622), .Z(n2627) );
  NANDN U5079 ( .A(n2625), .B(n2624), .Z(n2626) );
  AND U5080 ( .A(n2627), .B(n2626), .Z(n3699) );
  XOR U5081 ( .A(n3700), .B(n3699), .Z(n2628) );
  XNOR U5082 ( .A(n3701), .B(n2628), .Z(n3705) );
  XNOR U5083 ( .A(n3706), .B(n3705), .Z(n3707) );
  XOR U5084 ( .A(n3708), .B(n3707), .Z(n3766) );
  XNOR U5085 ( .A(n3767), .B(n3766), .Z(n2629) );
  XNOR U5086 ( .A(n3765), .B(n2629), .Z(n4045) );
  XNOR U5087 ( .A(n4047), .B(n4045), .Z(n2630) );
  XNOR U5088 ( .A(n4044), .B(n2630), .Z(n3493) );
  XNOR U5089 ( .A(n3493), .B(n3494), .Z(n3496) );
  XOR U5090 ( .A(n3495), .B(n3496), .Z(n3481) );
  XNOR U5091 ( .A(n3482), .B(n3481), .Z(n3484) );
  NANDN U5092 ( .A(n2636), .B(n2635), .Z(n2640) );
  NANDN U5093 ( .A(n2638), .B(n2637), .Z(n2639) );
  AND U5094 ( .A(n2640), .B(n2639), .Z(n3772) );
  NAND U5095 ( .A(n2642), .B(n2641), .Z(n2646) );
  NANDN U5096 ( .A(n2644), .B(n2643), .Z(n2645) );
  AND U5097 ( .A(n2646), .B(n2645), .Z(n3770) );
  NANDN U5098 ( .A(n2648), .B(n2647), .Z(n2652) );
  NAND U5099 ( .A(n2650), .B(n2649), .Z(n2651) );
  NAND U5100 ( .A(n2652), .B(n2651), .Z(n4479) );
  NANDN U5101 ( .A(n2654), .B(n2653), .Z(n2658) );
  NAND U5102 ( .A(n2656), .B(n2655), .Z(n2657) );
  AND U5103 ( .A(n2658), .B(n2657), .Z(n4094) );
  NAND U5104 ( .A(n2660), .B(n2659), .Z(n2664) );
  NAND U5105 ( .A(n2662), .B(n2661), .Z(n2663) );
  AND U5106 ( .A(n2664), .B(n2663), .Z(n4095) );
  NAND U5107 ( .A(n2666), .B(n2665), .Z(n2670) );
  NAND U5108 ( .A(n2668), .B(n2667), .Z(n2669) );
  AND U5109 ( .A(n2670), .B(n2669), .Z(n4097) );
  NAND U5110 ( .A(n2672), .B(n2671), .Z(n2676) );
  NAND U5111 ( .A(n2674), .B(n2673), .Z(n2675) );
  AND U5112 ( .A(n2676), .B(n2675), .Z(n3596) );
  NAND U5113 ( .A(n2678), .B(n2677), .Z(n2682) );
  NAND U5114 ( .A(n2680), .B(n2679), .Z(n2681) );
  AND U5115 ( .A(n2682), .B(n2681), .Z(n3597) );
  NAND U5116 ( .A(n2684), .B(n2683), .Z(n2688) );
  NAND U5117 ( .A(n2686), .B(n2685), .Z(n2687) );
  AND U5118 ( .A(n2688), .B(n2687), .Z(n3599) );
  XNOR U5119 ( .A(n3598), .B(n3599), .Z(n3735) );
  NAND U5120 ( .A(n2690), .B(n2689), .Z(n2694) );
  NAND U5121 ( .A(n2692), .B(n2691), .Z(n2693) );
  AND U5122 ( .A(n2694), .B(n2693), .Z(n3901) );
  NAND U5123 ( .A(n2696), .B(n2695), .Z(n2700) );
  NAND U5124 ( .A(n2698), .B(n2697), .Z(n2699) );
  NAND U5125 ( .A(n2700), .B(n2699), .Z(n3902) );
  XNOR U5126 ( .A(n3901), .B(n3902), .Z(n3903) );
  NANDN U5127 ( .A(n2702), .B(n2701), .Z(n2706) );
  NAND U5128 ( .A(n2704), .B(n2703), .Z(n2705) );
  NAND U5129 ( .A(n2706), .B(n2705), .Z(n3904) );
  XNOR U5130 ( .A(n3903), .B(n3904), .Z(n3736) );
  XOR U5131 ( .A(n3735), .B(n3736), .Z(n2707) );
  XNOR U5132 ( .A(n3737), .B(n2707), .Z(n4476) );
  NANDN U5133 ( .A(n2709), .B(n2708), .Z(n2713) );
  NAND U5134 ( .A(n2711), .B(n2710), .Z(n2712) );
  NAND U5135 ( .A(n2713), .B(n2712), .Z(n4477) );
  XOR U5136 ( .A(n3770), .B(n3769), .Z(n3771) );
  XOR U5137 ( .A(n3772), .B(n3771), .Z(n3274) );
  NANDN U5138 ( .A(n2715), .B(n2714), .Z(n2719) );
  NANDN U5139 ( .A(n2717), .B(n2716), .Z(n2718) );
  AND U5140 ( .A(n2719), .B(n2718), .Z(n3400) );
  NAND U5141 ( .A(n2721), .B(n2720), .Z(n2725) );
  NAND U5142 ( .A(n2723), .B(n2722), .Z(n2724) );
  NAND U5143 ( .A(n2725), .B(n2724), .Z(n4503) );
  NAND U5144 ( .A(n2727), .B(n2726), .Z(n2731) );
  NAND U5145 ( .A(n2729), .B(n2728), .Z(n2730) );
  NAND U5146 ( .A(n2731), .B(n2730), .Z(n4501) );
  NAND U5147 ( .A(n2733), .B(n2732), .Z(n2737) );
  NAND U5148 ( .A(n2735), .B(n2734), .Z(n2736) );
  AND U5149 ( .A(n2737), .B(n2736), .Z(n3590) );
  NAND U5150 ( .A(n2739), .B(n2738), .Z(n2743) );
  NAND U5151 ( .A(n2741), .B(n2740), .Z(n2742) );
  AND U5152 ( .A(n2743), .B(n2742), .Z(n3591) );
  NAND U5153 ( .A(n2745), .B(n2744), .Z(n2749) );
  NAND U5154 ( .A(n2747), .B(n2746), .Z(n2748) );
  AND U5155 ( .A(n2749), .B(n2748), .Z(n3592) );
  XOR U5156 ( .A(n3593), .B(n3592), .Z(n3750) );
  NAND U5157 ( .A(n2751), .B(n2750), .Z(n2755) );
  NAND U5158 ( .A(n2753), .B(n2752), .Z(n2754) );
  AND U5159 ( .A(n2755), .B(n2754), .Z(n3913) );
  NAND U5160 ( .A(n2757), .B(n2756), .Z(n2761) );
  NAND U5161 ( .A(n2759), .B(n2758), .Z(n2760) );
  NAND U5162 ( .A(n2761), .B(n2760), .Z(n3914) );
  XNOR U5163 ( .A(n3913), .B(n3914), .Z(n3916) );
  NANDN U5164 ( .A(n2763), .B(n2762), .Z(n2767) );
  NAND U5165 ( .A(n2765), .B(n2764), .Z(n2766) );
  AND U5166 ( .A(n2767), .B(n2766), .Z(n3915) );
  XOR U5167 ( .A(n3916), .B(n3915), .Z(n3748) );
  NANDN U5168 ( .A(n2769), .B(n2768), .Z(n2773) );
  NANDN U5169 ( .A(n2771), .B(n2770), .Z(n2772) );
  AND U5170 ( .A(n2773), .B(n2772), .Z(n3747) );
  XNOR U5171 ( .A(n3748), .B(n3747), .Z(n3749) );
  XOR U5172 ( .A(n3750), .B(n3749), .Z(n4500) );
  NAND U5173 ( .A(n2775), .B(n2774), .Z(n2779) );
  NAND U5174 ( .A(n2777), .B(n2776), .Z(n2778) );
  NAND U5175 ( .A(n2779), .B(n2778), .Z(n3398) );
  XNOR U5176 ( .A(n3397), .B(n3398), .Z(n3399) );
  XOR U5177 ( .A(n3400), .B(n3399), .Z(n3272) );
  NAND U5178 ( .A(n2781), .B(n2780), .Z(n2785) );
  NAND U5179 ( .A(n2783), .B(n2782), .Z(n2784) );
  NAND U5180 ( .A(n2785), .B(n2784), .Z(n4663) );
  NAND U5181 ( .A(n2787), .B(n2786), .Z(n2791) );
  NAND U5182 ( .A(n2789), .B(n2788), .Z(n2790) );
  NAND U5183 ( .A(n2791), .B(n2790), .Z(n3809) );
  NANDN U5184 ( .A(n2793), .B(n2792), .Z(n2797) );
  NANDN U5185 ( .A(n2795), .B(n2794), .Z(n2796) );
  AND U5186 ( .A(n2797), .B(n2796), .Z(n4449) );
  NAND U5187 ( .A(n2799), .B(n2798), .Z(n2803) );
  NAND U5188 ( .A(n2801), .B(n2800), .Z(n2802) );
  AND U5189 ( .A(n2803), .B(n2802), .Z(n4368) );
  NAND U5190 ( .A(n2805), .B(n2804), .Z(n2809) );
  NAND U5191 ( .A(n2807), .B(n2806), .Z(n2808) );
  NAND U5192 ( .A(n2809), .B(n2808), .Z(n4369) );
  XNOR U5193 ( .A(n4368), .B(n4369), .Z(n4371) );
  NAND U5194 ( .A(n2811), .B(n2810), .Z(n2815) );
  NAND U5195 ( .A(n2813), .B(n2812), .Z(n2814) );
  AND U5196 ( .A(n2815), .B(n2814), .Z(n4370) );
  XNOR U5197 ( .A(n4371), .B(n4370), .Z(n4447) );
  NANDN U5198 ( .A(n2817), .B(n2816), .Z(n2821) );
  NANDN U5199 ( .A(n2819), .B(n2818), .Z(n2820) );
  AND U5200 ( .A(n2821), .B(n2820), .Z(n4446) );
  XNOR U5201 ( .A(n4449), .B(n4448), .Z(n3807) );
  NANDN U5202 ( .A(n2823), .B(n2822), .Z(n2827) );
  NAND U5203 ( .A(n2825), .B(n2824), .Z(n2826) );
  AND U5204 ( .A(n2827), .B(n2826), .Z(n4211) );
  NANDN U5205 ( .A(n2829), .B(n2828), .Z(n2833) );
  NAND U5206 ( .A(n2831), .B(n2830), .Z(n2832) );
  AND U5207 ( .A(n2833), .B(n2832), .Z(n4212) );
  NAND U5208 ( .A(n2835), .B(n2834), .Z(n2839) );
  NAND U5209 ( .A(n2837), .B(n2836), .Z(n2838) );
  AND U5210 ( .A(n2839), .B(n2838), .Z(n4213) );
  XOR U5211 ( .A(n4214), .B(n4213), .Z(n4461) );
  NAND U5212 ( .A(n2841), .B(n2840), .Z(n2845) );
  NAND U5213 ( .A(n2843), .B(n2842), .Z(n2844) );
  NAND U5214 ( .A(n2845), .B(n2844), .Z(n4459) );
  NAND U5215 ( .A(n2847), .B(n2846), .Z(n2851) );
  NAND U5216 ( .A(n2849), .B(n2848), .Z(n2850) );
  AND U5217 ( .A(n2851), .B(n2850), .Z(n3824) );
  NAND U5218 ( .A(n2853), .B(n2852), .Z(n2857) );
  NAND U5219 ( .A(n2855), .B(n2854), .Z(n2856) );
  AND U5220 ( .A(n2857), .B(n2856), .Z(n3825) );
  NAND U5221 ( .A(n2859), .B(n2858), .Z(n2863) );
  NAND U5222 ( .A(n2861), .B(n2860), .Z(n2862) );
  AND U5223 ( .A(n2863), .B(n2862), .Z(n3826) );
  XNOR U5224 ( .A(n3827), .B(n3826), .Z(n4458) );
  XOR U5225 ( .A(n4461), .B(n4460), .Z(n3806) );
  NANDN U5226 ( .A(n2865), .B(n2864), .Z(n2869) );
  NANDN U5227 ( .A(n2867), .B(n2866), .Z(n2868) );
  NAND U5228 ( .A(n2869), .B(n2868), .Z(n4662) );
  XOR U5229 ( .A(n4664), .B(n4662), .Z(n2870) );
  XOR U5230 ( .A(n4663), .B(n2870), .Z(n3271) );
  XNOR U5231 ( .A(n3272), .B(n3271), .Z(n3273) );
  XOR U5232 ( .A(n3274), .B(n3273), .Z(n3259) );
  NAND U5233 ( .A(n2872), .B(n2871), .Z(n2876) );
  NAND U5234 ( .A(n2874), .B(n2873), .Z(n2875) );
  AND U5235 ( .A(n2876), .B(n2875), .Z(n4041) );
  NAND U5236 ( .A(n2878), .B(n2877), .Z(n2882) );
  NAND U5237 ( .A(n2880), .B(n2879), .Z(n2881) );
  AND U5238 ( .A(n2882), .B(n2881), .Z(n3704) );
  NANDN U5239 ( .A(n2884), .B(n2883), .Z(n2888) );
  NANDN U5240 ( .A(n2886), .B(n2885), .Z(n2887) );
  NAND U5241 ( .A(n2888), .B(n2887), .Z(n3702) );
  NANDN U5242 ( .A(n2890), .B(n2889), .Z(n2894) );
  NAND U5243 ( .A(n2892), .B(n2891), .Z(n2893) );
  AND U5244 ( .A(n2894), .B(n2893), .Z(n4410) );
  NANDN U5245 ( .A(n2896), .B(n2895), .Z(n2900) );
  NAND U5246 ( .A(n2898), .B(n2897), .Z(n2899) );
  AND U5247 ( .A(n2900), .B(n2899), .Z(n4411) );
  NANDN U5248 ( .A(n2902), .B(n2901), .Z(n2906) );
  NAND U5249 ( .A(n2904), .B(n2903), .Z(n2905) );
  AND U5250 ( .A(n2906), .B(n2905), .Z(n4412) );
  XNOR U5251 ( .A(n4413), .B(n4412), .Z(n3703) );
  XNOR U5252 ( .A(n3702), .B(n3703), .Z(n2907) );
  XOR U5253 ( .A(n3704), .B(n2907), .Z(n4335) );
  NAND U5254 ( .A(n2909), .B(n2908), .Z(n2913) );
  NAND U5255 ( .A(n2911), .B(n2910), .Z(n2912) );
  AND U5256 ( .A(n2913), .B(n2912), .Z(n4551) );
  NAND U5257 ( .A(n2915), .B(n2914), .Z(n2919) );
  NAND U5258 ( .A(n2917), .B(n2916), .Z(n2918) );
  AND U5259 ( .A(n2919), .B(n2918), .Z(n4518) );
  NANDN U5260 ( .A(n2921), .B(n2920), .Z(n2925) );
  NAND U5261 ( .A(n2923), .B(n2922), .Z(n2924) );
  NAND U5262 ( .A(n2925), .B(n2924), .Z(n4519) );
  XNOR U5263 ( .A(n4518), .B(n4519), .Z(n4521) );
  NANDN U5264 ( .A(n2927), .B(n2926), .Z(n2931) );
  NAND U5265 ( .A(n2929), .B(n2928), .Z(n2930) );
  AND U5266 ( .A(n2931), .B(n2930), .Z(n4520) );
  XOR U5267 ( .A(n4521), .B(n4520), .Z(n4549) );
  NAND U5268 ( .A(n2933), .B(n2932), .Z(n2937) );
  NAND U5269 ( .A(n2935), .B(n2934), .Z(n2936) );
  AND U5270 ( .A(n2937), .B(n2936), .Z(n4548) );
  XNOR U5271 ( .A(n4549), .B(n4548), .Z(n4550) );
  XOR U5272 ( .A(n4551), .B(n4550), .Z(n4333) );
  NANDN U5273 ( .A(n2939), .B(n2938), .Z(n2943) );
  NANDN U5274 ( .A(n2941), .B(n2940), .Z(n2942) );
  AND U5275 ( .A(n2943), .B(n2942), .Z(n4653) );
  NAND U5276 ( .A(n2945), .B(n2944), .Z(n2949) );
  NAND U5277 ( .A(n2947), .B(n2946), .Z(n2948) );
  AND U5278 ( .A(n2949), .B(n2948), .Z(n4386) );
  NAND U5279 ( .A(n2951), .B(n2950), .Z(n2955) );
  NAND U5280 ( .A(n2953), .B(n2952), .Z(n2954) );
  AND U5281 ( .A(n2955), .B(n2954), .Z(n4387) );
  NANDN U5282 ( .A(n2957), .B(n2956), .Z(n2961) );
  NAND U5283 ( .A(n2959), .B(n2958), .Z(n2960) );
  AND U5284 ( .A(n2961), .B(n2960), .Z(n4388) );
  XOR U5285 ( .A(n4389), .B(n4388), .Z(n4651) );
  NANDN U5286 ( .A(n2963), .B(n2962), .Z(n2967) );
  NANDN U5287 ( .A(n2965), .B(n2964), .Z(n2966) );
  AND U5288 ( .A(n2967), .B(n2966), .Z(n4650) );
  XNOR U5289 ( .A(n4651), .B(n4650), .Z(n4652) );
  XNOR U5290 ( .A(n4653), .B(n4652), .Z(n4332) );
  XNOR U5291 ( .A(n4333), .B(n4332), .Z(n4334) );
  XOR U5292 ( .A(n4335), .B(n4334), .Z(n4149) );
  NAND U5293 ( .A(n2969), .B(n2968), .Z(n2973) );
  NAND U5294 ( .A(n2971), .B(n2970), .Z(n2972) );
  NAND U5295 ( .A(n2973), .B(n2972), .Z(n4580) );
  NAND U5296 ( .A(n2975), .B(n2974), .Z(n2979) );
  NAND U5297 ( .A(n2977), .B(n2976), .Z(n2978) );
  AND U5298 ( .A(n2979), .B(n2978), .Z(n3620) );
  NAND U5299 ( .A(n2981), .B(n2980), .Z(n2985) );
  NAND U5300 ( .A(n2983), .B(n2982), .Z(n2984) );
  AND U5301 ( .A(n2985), .B(n2984), .Z(n3621) );
  NAND U5302 ( .A(n2987), .B(n2986), .Z(n2991) );
  NAND U5303 ( .A(n2989), .B(n2988), .Z(n2990) );
  AND U5304 ( .A(n2991), .B(n2990), .Z(n3622) );
  XOR U5305 ( .A(n3623), .B(n3622), .Z(n4557) );
  NAND U5306 ( .A(n2993), .B(n2992), .Z(n2997) );
  NAND U5307 ( .A(n2995), .B(n2994), .Z(n2996) );
  AND U5308 ( .A(n2997), .B(n2996), .Z(n4572) );
  NAND U5309 ( .A(n2999), .B(n2998), .Z(n3003) );
  NAND U5310 ( .A(n3001), .B(n3000), .Z(n3002) );
  AND U5311 ( .A(n3003), .B(n3002), .Z(n4573) );
  NAND U5312 ( .A(n3005), .B(n3004), .Z(n3009) );
  NAND U5313 ( .A(n3007), .B(n3006), .Z(n3008) );
  AND U5314 ( .A(n3009), .B(n3008), .Z(n4574) );
  XOR U5315 ( .A(n4575), .B(n4574), .Z(n4555) );
  NAND U5316 ( .A(n3011), .B(n3010), .Z(n3015) );
  NAND U5317 ( .A(n3013), .B(n3012), .Z(n3014) );
  AND U5318 ( .A(n3015), .B(n3014), .Z(n4554) );
  XNOR U5319 ( .A(n4555), .B(n4554), .Z(n4556) );
  XNOR U5320 ( .A(n4557), .B(n4556), .Z(n4579) );
  NAND U5321 ( .A(n3017), .B(n3016), .Z(n3021) );
  NAND U5322 ( .A(n3019), .B(n3018), .Z(n3020) );
  AND U5323 ( .A(n3021), .B(n3020), .Z(n4136) );
  NANDN U5324 ( .A(n3023), .B(n3022), .Z(n3027) );
  NAND U5325 ( .A(n3025), .B(n3024), .Z(n3026) );
  AND U5326 ( .A(n3027), .B(n3026), .Z(n4137) );
  NAND U5327 ( .A(n3029), .B(n3028), .Z(n3033) );
  NAND U5328 ( .A(n3031), .B(n3030), .Z(n3032) );
  AND U5329 ( .A(n3033), .B(n3032), .Z(n4138) );
  XNOR U5330 ( .A(n4139), .B(n4138), .Z(n3922) );
  NAND U5331 ( .A(n3035), .B(n3034), .Z(n3039) );
  NAND U5332 ( .A(n3037), .B(n3036), .Z(n3038) );
  AND U5333 ( .A(n3039), .B(n3038), .Z(n4124) );
  NAND U5334 ( .A(n3041), .B(n3040), .Z(n3045) );
  NAND U5335 ( .A(n3043), .B(n3042), .Z(n3044) );
  AND U5336 ( .A(n3045), .B(n3044), .Z(n4125) );
  NAND U5337 ( .A(n3047), .B(n3046), .Z(n3051) );
  NAND U5338 ( .A(n3049), .B(n3048), .Z(n3050) );
  AND U5339 ( .A(n3051), .B(n3050), .Z(n4126) );
  XOR U5340 ( .A(n4127), .B(n4126), .Z(n3920) );
  NAND U5341 ( .A(n3053), .B(n3052), .Z(n3057) );
  NAND U5342 ( .A(n3055), .B(n3054), .Z(n3056) );
  AND U5343 ( .A(n3057), .B(n3056), .Z(n3919) );
  XNOR U5344 ( .A(n3920), .B(n3919), .Z(n3921) );
  XNOR U5345 ( .A(n3922), .B(n3921), .Z(n4578) );
  XOR U5346 ( .A(n4579), .B(n4578), .Z(n4581) );
  XOR U5347 ( .A(n4580), .B(n4581), .Z(n4151) );
  NANDN U5348 ( .A(n3059), .B(n3058), .Z(n3063) );
  NAND U5349 ( .A(n3061), .B(n3060), .Z(n3062) );
  AND U5350 ( .A(n3063), .B(n3062), .Z(n3889) );
  NAND U5351 ( .A(n3065), .B(n3064), .Z(n3069) );
  NAND U5352 ( .A(n3067), .B(n3066), .Z(n3068) );
  NAND U5353 ( .A(n3069), .B(n3068), .Z(n3890) );
  XNOR U5354 ( .A(n3889), .B(n3890), .Z(n3892) );
  NANDN U5355 ( .A(n3071), .B(n3070), .Z(n3075) );
  NAND U5356 ( .A(n3073), .B(n3072), .Z(n3074) );
  AND U5357 ( .A(n3075), .B(n3074), .Z(n3891) );
  XOR U5358 ( .A(n3892), .B(n3891), .Z(n4257) );
  NAND U5359 ( .A(n3077), .B(n3076), .Z(n3081) );
  NAND U5360 ( .A(n3079), .B(n3078), .Z(n3080) );
  AND U5361 ( .A(n3081), .B(n3080), .Z(n3319) );
  NAND U5362 ( .A(n3083), .B(n3082), .Z(n3087) );
  NAND U5363 ( .A(n3085), .B(n3084), .Z(n3086) );
  NAND U5364 ( .A(n3087), .B(n3086), .Z(n3320) );
  XNOR U5365 ( .A(n3319), .B(n3320), .Z(n3322) );
  NAND U5366 ( .A(n3089), .B(n3088), .Z(n3093) );
  NAND U5367 ( .A(n3091), .B(n3090), .Z(n3092) );
  AND U5368 ( .A(n3093), .B(n3092), .Z(n3321) );
  XOR U5369 ( .A(n3322), .B(n3321), .Z(n4255) );
  NAND U5370 ( .A(n3095), .B(n3094), .Z(n3099) );
  NAND U5371 ( .A(n3097), .B(n3096), .Z(n3098) );
  AND U5372 ( .A(n3099), .B(n3098), .Z(n4254) );
  XNOR U5373 ( .A(n4255), .B(n4254), .Z(n4256) );
  XNOR U5374 ( .A(n4257), .B(n4256), .Z(n4154) );
  NAND U5375 ( .A(n3101), .B(n3100), .Z(n3105) );
  NAND U5376 ( .A(n3103), .B(n3102), .Z(n3104) );
  AND U5377 ( .A(n3105), .B(n3104), .Z(n4153) );
  NAND U5378 ( .A(n3107), .B(n3106), .Z(n3111) );
  NAND U5379 ( .A(n3109), .B(n3108), .Z(n3110) );
  AND U5380 ( .A(n3111), .B(n3110), .Z(n4152) );
  XNOR U5381 ( .A(n4153), .B(n4152), .Z(n3112) );
  XNOR U5382 ( .A(n4154), .B(n3112), .Z(n4150) );
  IV U5383 ( .A(n4150), .Z(n4148) );
  XNOR U5384 ( .A(n4151), .B(n4148), .Z(n3113) );
  XNOR U5385 ( .A(n4149), .B(n3113), .Z(n4038) );
  NANDN U5386 ( .A(n3115), .B(n3114), .Z(n3119) );
  NANDN U5387 ( .A(n3117), .B(n3116), .Z(n3118) );
  AND U5388 ( .A(n3119), .B(n3118), .Z(n4039) );
  XNOR U5389 ( .A(n4038), .B(n4039), .Z(n4040) );
  XOR U5390 ( .A(n4041), .B(n4040), .Z(n3260) );
  XOR U5391 ( .A(n3259), .B(n3260), .Z(n3262) );
  NANDN U5392 ( .A(n3121), .B(n3120), .Z(n3125) );
  NAND U5393 ( .A(n3123), .B(n3122), .Z(n3124) );
  AND U5394 ( .A(n3125), .B(n3124), .Z(n3268) );
  NAND U5395 ( .A(n3127), .B(n3126), .Z(n3131) );
  NAND U5396 ( .A(n3129), .B(n3128), .Z(n3130) );
  AND U5397 ( .A(n3131), .B(n3130), .Z(n3390) );
  NAND U5398 ( .A(n3133), .B(n3132), .Z(n3137) );
  NAND U5399 ( .A(n3135), .B(n3134), .Z(n3136) );
  AND U5400 ( .A(n3137), .B(n3136), .Z(n3313) );
  NANDN U5401 ( .A(n3139), .B(n3138), .Z(n3143) );
  NAND U5402 ( .A(n3141), .B(n3140), .Z(n3142) );
  NAND U5403 ( .A(n3143), .B(n3142), .Z(n3314) );
  XNOR U5404 ( .A(n3313), .B(n3314), .Z(n3316) );
  NAND U5405 ( .A(n3145), .B(n3144), .Z(n3149) );
  NAND U5406 ( .A(n3147), .B(n3146), .Z(n3148) );
  AND U5407 ( .A(n3149), .B(n3148), .Z(n3315) );
  XNOR U5408 ( .A(n3316), .B(n3315), .Z(n3714) );
  NANDN U5409 ( .A(n3151), .B(n3150), .Z(n3155) );
  NAND U5410 ( .A(n3153), .B(n3152), .Z(n3154) );
  AND U5411 ( .A(n3155), .B(n3154), .Z(n4512) );
  NANDN U5412 ( .A(n3157), .B(n3156), .Z(n3161) );
  NAND U5413 ( .A(n3159), .B(n3158), .Z(n3160) );
  AND U5414 ( .A(n3161), .B(n3160), .Z(n4513) );
  NAND U5415 ( .A(n3163), .B(n3162), .Z(n3167) );
  NAND U5416 ( .A(n3165), .B(n3164), .Z(n3166) );
  AND U5417 ( .A(n3167), .B(n3166), .Z(n4514) );
  XNOR U5418 ( .A(n4515), .B(n4514), .Z(n3712) );
  NAND U5419 ( .A(n3169), .B(n3168), .Z(n3173) );
  NAND U5420 ( .A(n3171), .B(n3170), .Z(n3172) );
  AND U5421 ( .A(n3173), .B(n3172), .Z(n3446) );
  NAND U5422 ( .A(n3175), .B(n3174), .Z(n3179) );
  NAND U5423 ( .A(n3177), .B(n3176), .Z(n3178) );
  NAND U5424 ( .A(n3179), .B(n3178), .Z(n3447) );
  XNOR U5425 ( .A(n3446), .B(n3447), .Z(n3449) );
  NAND U5426 ( .A(n3181), .B(n3180), .Z(n3185) );
  NAND U5427 ( .A(n3183), .B(n3182), .Z(n3184) );
  AND U5428 ( .A(n3185), .B(n3184), .Z(n3448) );
  XNOR U5429 ( .A(n3449), .B(n3448), .Z(n3711) );
  NAND U5430 ( .A(n3187), .B(n3186), .Z(n3191) );
  NAND U5431 ( .A(n3189), .B(n3188), .Z(n3190) );
  AND U5432 ( .A(n3191), .B(n3190), .Z(n3614) );
  NAND U5433 ( .A(n3193), .B(n3192), .Z(n3197) );
  NAND U5434 ( .A(n3195), .B(n3194), .Z(n3196) );
  AND U5435 ( .A(n3197), .B(n3196), .Z(n3615) );
  NAND U5436 ( .A(n3199), .B(n3198), .Z(n3203) );
  NAND U5437 ( .A(n3201), .B(n3200), .Z(n3202) );
  AND U5438 ( .A(n3203), .B(n3202), .Z(n3616) );
  XOR U5439 ( .A(n3617), .B(n3616), .Z(n3720) );
  NAND U5440 ( .A(n3205), .B(n3204), .Z(n3209) );
  NAND U5441 ( .A(n3207), .B(n3206), .Z(n3208) );
  AND U5442 ( .A(n3209), .B(n3208), .Z(n4260) );
  NAND U5443 ( .A(n3211), .B(n3210), .Z(n3215) );
  NAND U5444 ( .A(n3213), .B(n3212), .Z(n3214) );
  AND U5445 ( .A(n3215), .B(n3214), .Z(n4261) );
  NAND U5446 ( .A(n3217), .B(n3216), .Z(n3221) );
  NAND U5447 ( .A(n3219), .B(n3218), .Z(n3220) );
  AND U5448 ( .A(n3221), .B(n3220), .Z(n4262) );
  XNOR U5449 ( .A(n4263), .B(n4262), .Z(n3718) );
  NAND U5450 ( .A(n3223), .B(n3222), .Z(n3227) );
  NAND U5451 ( .A(n3225), .B(n3224), .Z(n3226) );
  AND U5452 ( .A(n3227), .B(n3226), .Z(n3577) );
  NAND U5453 ( .A(n3229), .B(n3228), .Z(n3233) );
  NAND U5454 ( .A(n3231), .B(n3230), .Z(n3232) );
  NAND U5455 ( .A(n3233), .B(n3232), .Z(n3578) );
  XNOR U5456 ( .A(n3577), .B(n3578), .Z(n3580) );
  NAND U5457 ( .A(n3235), .B(n3234), .Z(n3239) );
  NAND U5458 ( .A(n3237), .B(n3236), .Z(n3238) );
  AND U5459 ( .A(n3239), .B(n3238), .Z(n3579) );
  XNOR U5460 ( .A(n3580), .B(n3579), .Z(n3717) );
  XOR U5461 ( .A(n3720), .B(n3719), .Z(n3387) );
  XOR U5462 ( .A(n3388), .B(n3387), .Z(n3389) );
  XOR U5463 ( .A(n3390), .B(n3389), .Z(n3407) );
  NANDN U5464 ( .A(n3241), .B(n3240), .Z(n3245) );
  NANDN U5465 ( .A(n3243), .B(n3242), .Z(n3244) );
  AND U5466 ( .A(n3245), .B(n3244), .Z(n3408) );
  NANDN U5467 ( .A(n3247), .B(n3246), .Z(n3251) );
  NAND U5468 ( .A(n3249), .B(n3248), .Z(n3250) );
  AND U5469 ( .A(n3251), .B(n3250), .Z(n3406) );
  XNOR U5470 ( .A(n3408), .B(n3406), .Z(n3252) );
  XOR U5471 ( .A(n3407), .B(n3252), .Z(n3265) );
  NANDN U5472 ( .A(n3254), .B(n3253), .Z(n3258) );
  NAND U5473 ( .A(n3256), .B(n3255), .Z(n3257) );
  NAND U5474 ( .A(n3258), .B(n3257), .Z(n3266) );
  XNOR U5475 ( .A(n3265), .B(n3266), .Z(n3267) );
  XNOR U5476 ( .A(n3268), .B(n3267), .Z(n3261) );
  XOR U5477 ( .A(n3262), .B(n3261), .Z(n3483) );
  XNOR U5478 ( .A(n3484), .B(n3483), .Z(o[1]) );
  NAND U5479 ( .A(n3260), .B(n3259), .Z(n3264) );
  NAND U5480 ( .A(n3262), .B(n3261), .Z(n3263) );
  AND U5481 ( .A(n3264), .B(n3263), .Z(n5359) );
  NANDN U5482 ( .A(n3266), .B(n3265), .Z(n3270) );
  NANDN U5483 ( .A(n3268), .B(n3267), .Z(n3269) );
  AND U5484 ( .A(n3270), .B(n3269), .Z(n4677) );
  NANDN U5485 ( .A(n3272), .B(n3271), .Z(n3276) );
  NANDN U5486 ( .A(n3274), .B(n3273), .Z(n3275) );
  AND U5487 ( .A(n3276), .B(n3275), .Z(n4675) );
  NANDN U5488 ( .A(n3278), .B(n3277), .Z(n3282) );
  NAND U5489 ( .A(n3280), .B(n3279), .Z(n3281) );
  AND U5490 ( .A(n3282), .B(n3281), .Z(n4732) );
  NAND U5491 ( .A(n3284), .B(n3283), .Z(n3288) );
  NAND U5492 ( .A(n3286), .B(n3285), .Z(n3287) );
  NAND U5493 ( .A(n3288), .B(n3287), .Z(n5279) );
  XNOR U5494 ( .A(n5277), .B(n5276), .Z(n5278) );
  NAND U5495 ( .A(n3299), .B(n3298), .Z(n3303) );
  NAND U5496 ( .A(n3301), .B(n3300), .Z(n3302) );
  NAND U5497 ( .A(n3303), .B(n3302), .Z(n4807) );
  IV U5498 ( .A(n4807), .Z(n3311) );
  XOR U5499 ( .A(n4806), .B(n4805), .Z(n3310) );
  XNOR U5500 ( .A(n3311), .B(n3310), .Z(n5008) );
  XNOR U5501 ( .A(n5006), .B(n5008), .Z(n3312) );
  XOR U5502 ( .A(n5007), .B(n3312), .Z(n4730) );
  NANDN U5503 ( .A(n3314), .B(n3313), .Z(n3318) );
  NAND U5504 ( .A(n3316), .B(n3315), .Z(n3317) );
  NAND U5505 ( .A(n3318), .B(n3317), .Z(n4909) );
  NANDN U5506 ( .A(n3320), .B(n3319), .Z(n3324) );
  NAND U5507 ( .A(n3322), .B(n3321), .Z(n3323) );
  NAND U5508 ( .A(n3324), .B(n3323), .Z(n4907) );
  NAND U5509 ( .A(n3326), .B(n3325), .Z(n3330) );
  NAND U5510 ( .A(n3328), .B(n3327), .Z(n3329) );
  NAND U5511 ( .A(n3330), .B(n3329), .Z(n4906) );
  NAND U5512 ( .A(n3332), .B(n3331), .Z(n3338) );
  AND U5513 ( .A(n3334), .B(n3333), .Z(n3336) );
  OR U5514 ( .A(n3336), .B(n3335), .Z(n3337) );
  AND U5515 ( .A(n3338), .B(n3337), .Z(n4998) );
  NAND U5516 ( .A(n3340), .B(n3339), .Z(n3344) );
  NAND U5517 ( .A(n3342), .B(n3341), .Z(n3343) );
  NAND U5518 ( .A(n3344), .B(n3343), .Z(n5302) );
  XNOR U5519 ( .A(n5301), .B(n5300), .Z(n5303) );
  XOR U5520 ( .A(n5302), .B(n5303), .Z(n4997) );
  XNOR U5521 ( .A(n4998), .B(n4997), .Z(n5000) );
  XOR U5522 ( .A(n4999), .B(n5000), .Z(n4729) );
  XNOR U5523 ( .A(n4730), .B(n4729), .Z(n4731) );
  XOR U5524 ( .A(n4732), .B(n4731), .Z(n4830) );
  NAND U5525 ( .A(n3352), .B(n3351), .Z(n3356) );
  NANDN U5526 ( .A(n3354), .B(n3353), .Z(n3355) );
  AND U5527 ( .A(n3356), .B(n3355), .Z(n4750) );
  NANDN U5528 ( .A(n3358), .B(n3357), .Z(n3362) );
  NANDN U5529 ( .A(n3360), .B(n3359), .Z(n3361) );
  AND U5530 ( .A(n3362), .B(n3361), .Z(n4748) );
  NAND U5531 ( .A(n3364), .B(n3363), .Z(n3368) );
  NAND U5532 ( .A(n3366), .B(n3365), .Z(n3367) );
  NAND U5533 ( .A(n3368), .B(n3367), .Z(n4747) );
  XNOR U5534 ( .A(n4748), .B(n4747), .Z(n4749) );
  XOR U5535 ( .A(n4750), .B(n4749), .Z(n5150) );
  NANDN U5536 ( .A(n3370), .B(n3369), .Z(n3374) );
  NAND U5537 ( .A(n3372), .B(n3371), .Z(n3373) );
  AND U5538 ( .A(n3374), .B(n3373), .Z(n4713) );
  NANDN U5539 ( .A(n3376), .B(n3375), .Z(n3380) );
  NAND U5540 ( .A(n3378), .B(n3377), .Z(n3379) );
  AND U5541 ( .A(n3380), .B(n3379), .Z(n4711) );
  NANDN U5542 ( .A(n3382), .B(n3381), .Z(n3386) );
  NAND U5543 ( .A(n3384), .B(n3383), .Z(n3385) );
  NAND U5544 ( .A(n3386), .B(n3385), .Z(n4710) );
  XNOR U5545 ( .A(n4711), .B(n4710), .Z(n4712) );
  XOR U5546 ( .A(n4713), .B(n4712), .Z(n5149) );
  NAND U5547 ( .A(n3388), .B(n3387), .Z(n3392) );
  NANDN U5548 ( .A(n3390), .B(n3389), .Z(n3391) );
  NAND U5549 ( .A(n3392), .B(n3391), .Z(n5148) );
  XOR U5550 ( .A(n5149), .B(n5148), .Z(n5151) );
  XOR U5551 ( .A(n5150), .B(n5151), .Z(n4831) );
  XNOR U5552 ( .A(n4831), .B(n4829), .Z(n3396) );
  XOR U5553 ( .A(n4830), .B(n3396), .Z(n4674) );
  XNOR U5554 ( .A(n4675), .B(n4674), .Z(n4676) );
  XOR U5555 ( .A(n4677), .B(n4676), .Z(n5357) );
  NANDN U5556 ( .A(n3398), .B(n3397), .Z(n3402) );
  NAND U5557 ( .A(n3400), .B(n3399), .Z(n3401) );
  NAND U5558 ( .A(n3402), .B(n3401), .Z(n4926) );
  XNOR U5559 ( .A(n4925), .B(n4924), .Z(n3409) );
  XOR U5560 ( .A(n4926), .B(n3409), .Z(n5338) );
  NAND U5561 ( .A(n3411), .B(n3410), .Z(n3415) );
  NAND U5562 ( .A(n3413), .B(n3412), .Z(n3414) );
  AND U5563 ( .A(n3415), .B(n3414), .Z(n5337) );
  XNOR U5564 ( .A(n5338), .B(n5337), .Z(n5340) );
  NAND U5565 ( .A(n3417), .B(n3416), .Z(n3421) );
  NAND U5566 ( .A(n3419), .B(n3418), .Z(n3420) );
  NAND U5567 ( .A(n3421), .B(n3420), .Z(n4725) );
  NANDN U5568 ( .A(n3423), .B(n3422), .Z(n3427) );
  NANDN U5569 ( .A(n3425), .B(n3424), .Z(n3426) );
  AND U5570 ( .A(n3427), .B(n3426), .Z(n4737) );
  NANDN U5571 ( .A(n3429), .B(n3428), .Z(n3433) );
  NAND U5572 ( .A(n3431), .B(n3430), .Z(n3432) );
  NAND U5573 ( .A(n3433), .B(n3432), .Z(n4850) );
  NANDN U5574 ( .A(n3435), .B(n3434), .Z(n3439) );
  NANDN U5575 ( .A(n3437), .B(n3436), .Z(n3438) );
  NAND U5576 ( .A(n3439), .B(n3438), .Z(n4848) );
  NANDN U5577 ( .A(n3441), .B(n3440), .Z(n3445) );
  NAND U5578 ( .A(n3443), .B(n3442), .Z(n3444) );
  NAND U5579 ( .A(n3445), .B(n3444), .Z(n4847) );
  NANDN U5580 ( .A(n3447), .B(n3446), .Z(n3451) );
  NAND U5581 ( .A(n3449), .B(n3448), .Z(n3450) );
  NAND U5582 ( .A(n3451), .B(n3450), .Z(n4856) );
  XOR U5583 ( .A(n4854), .B(n4853), .Z(n4855) );
  IV U5584 ( .A(n4789), .Z(n4791) );
  XNOR U5585 ( .A(n4791), .B(n4790), .Z(n3461) );
  XNOR U5586 ( .A(n4792), .B(n3461), .Z(n4736) );
  NANDN U5587 ( .A(n3463), .B(n3462), .Z(n3467) );
  NAND U5588 ( .A(n3465), .B(n3464), .Z(n3466) );
  NAND U5589 ( .A(n3467), .B(n3466), .Z(n4788) );
  XNOR U5590 ( .A(n4787), .B(n4786), .Z(n3474) );
  XNOR U5591 ( .A(n4788), .B(n3474), .Z(n4735) );
  XNOR U5592 ( .A(n4737), .B(n4738), .Z(n4724) );
  NANDN U5593 ( .A(n3476), .B(n3475), .Z(n3480) );
  NAND U5594 ( .A(n3478), .B(n3477), .Z(n3479) );
  NAND U5595 ( .A(n3480), .B(n3479), .Z(n4723) );
  XNOR U5596 ( .A(n4724), .B(n4723), .Z(n4726) );
  XOR U5597 ( .A(n4725), .B(n4726), .Z(n5339) );
  XOR U5598 ( .A(n5340), .B(n5339), .Z(n5356) );
  XNOR U5599 ( .A(n5357), .B(n5356), .Z(n5358) );
  XOR U5600 ( .A(n5359), .B(n5358), .Z(n5355) );
  NANDN U5601 ( .A(n3482), .B(n3481), .Z(n3486) );
  NAND U5602 ( .A(n3484), .B(n3483), .Z(n3485) );
  NAND U5603 ( .A(n3486), .B(n3485), .Z(n5353) );
  NANDN U5604 ( .A(n3488), .B(n3487), .Z(n3492) );
  NANDN U5605 ( .A(n3490), .B(n3489), .Z(n3491) );
  AND U5606 ( .A(n3492), .B(n3491), .Z(n5349) );
  NANDN U5607 ( .A(n3494), .B(n3493), .Z(n3498) );
  NAND U5608 ( .A(n3496), .B(n3495), .Z(n3497) );
  AND U5609 ( .A(n3498), .B(n3497), .Z(n5371) );
  NANDN U5610 ( .A(n3500), .B(n3499), .Z(n3504) );
  NAND U5611 ( .A(n3502), .B(n3501), .Z(n3503) );
  NAND U5612 ( .A(n3504), .B(n3503), .Z(n4686) );
  NAND U5613 ( .A(n3506), .B(n3505), .Z(n3510) );
  NANDN U5614 ( .A(n3508), .B(n3507), .Z(n3509) );
  NAND U5615 ( .A(n3510), .B(n3509), .Z(n4920) );
  NANDN U5616 ( .A(n3512), .B(n3511), .Z(n3516) );
  NAND U5617 ( .A(n3514), .B(n3513), .Z(n3515) );
  NAND U5618 ( .A(n3516), .B(n3515), .Z(n4919) );
  NANDN U5619 ( .A(n3518), .B(n3517), .Z(n3522) );
  NANDN U5620 ( .A(n3520), .B(n3519), .Z(n3521) );
  NAND U5621 ( .A(n3522), .B(n3521), .Z(n4918) );
  XOR U5622 ( .A(n4919), .B(n4918), .Z(n4921) );
  XOR U5623 ( .A(n4920), .B(n4921), .Z(n4687) );
  XOR U5624 ( .A(n4686), .B(n4687), .Z(n4688) );
  NANDN U5625 ( .A(n3524), .B(n3523), .Z(n3528) );
  NANDN U5626 ( .A(n3526), .B(n3525), .Z(n3527) );
  AND U5627 ( .A(n3528), .B(n3527), .Z(n5107) );
  NAND U5628 ( .A(n3530), .B(n3529), .Z(n3534) );
  NAND U5629 ( .A(n3532), .B(n3531), .Z(n3533) );
  AND U5630 ( .A(n3534), .B(n3533), .Z(n5106) );
  XOR U5631 ( .A(n5107), .B(n5106), .Z(n5109) );
  NAND U5632 ( .A(n3536), .B(n3535), .Z(n3540) );
  NAND U5633 ( .A(n3538), .B(n3537), .Z(n3539) );
  AND U5634 ( .A(n3540), .B(n3539), .Z(n5108) );
  XNOR U5635 ( .A(n5109), .B(n5108), .Z(n4955) );
  NANDN U5636 ( .A(n3542), .B(n3541), .Z(n3546) );
  NANDN U5637 ( .A(n3544), .B(n3543), .Z(n3545) );
  NAND U5638 ( .A(n3546), .B(n3545), .Z(n4953) );
  NANDN U5639 ( .A(n3548), .B(n3547), .Z(n3552) );
  NANDN U5640 ( .A(n3550), .B(n3549), .Z(n3551) );
  NAND U5641 ( .A(n3552), .B(n3551), .Z(n4952) );
  XNOR U5642 ( .A(n4688), .B(n4689), .Z(n4683) );
  NAND U5643 ( .A(n3554), .B(n3553), .Z(n3558) );
  NAND U5644 ( .A(n3556), .B(n3555), .Z(n3557) );
  AND U5645 ( .A(n3558), .B(n3557), .Z(n5192) );
  NAND U5646 ( .A(n3560), .B(n3559), .Z(n3564) );
  NAND U5647 ( .A(n3562), .B(n3561), .Z(n3563) );
  AND U5648 ( .A(n3564), .B(n3563), .Z(n5193) );
  NAND U5649 ( .A(n3566), .B(n3565), .Z(n3570) );
  NAND U5650 ( .A(n3568), .B(n3567), .Z(n3569) );
  AND U5651 ( .A(n3570), .B(n3569), .Z(n5194) );
  XNOR U5652 ( .A(n5195), .B(n5194), .Z(n5237) );
  NAND U5653 ( .A(n3572), .B(n3571), .Z(n3576) );
  NAND U5654 ( .A(n3574), .B(n3573), .Z(n3575) );
  NAND U5655 ( .A(n3576), .B(n3575), .Z(n5235) );
  NANDN U5656 ( .A(n3578), .B(n3577), .Z(n3582) );
  NAND U5657 ( .A(n3580), .B(n3579), .Z(n3581) );
  AND U5658 ( .A(n3582), .B(n3581), .Z(n4804) );
  XNOR U5659 ( .A(n4803), .B(n4802), .Z(n3589) );
  XNOR U5660 ( .A(n4804), .B(n3589), .Z(n5183) );
  NAND U5661 ( .A(n3591), .B(n3590), .Z(n3595) );
  NAND U5662 ( .A(n3593), .B(n3592), .Z(n3594) );
  NAND U5663 ( .A(n3595), .B(n3594), .Z(n5159) );
  NAND U5664 ( .A(n3597), .B(n3596), .Z(n3601) );
  NAND U5665 ( .A(n3599), .B(n3598), .Z(n3600) );
  NAND U5666 ( .A(n3601), .B(n3600), .Z(n5157) );
  NAND U5667 ( .A(n3603), .B(n3602), .Z(n3607) );
  NAND U5668 ( .A(n3605), .B(n3604), .Z(n3606) );
  NAND U5669 ( .A(n3607), .B(n3606), .Z(n5156) );
  NAND U5670 ( .A(n3609), .B(n3608), .Z(n3613) );
  NAND U5671 ( .A(n3611), .B(n3610), .Z(n3612) );
  AND U5672 ( .A(n3613), .B(n3612), .Z(n5036) );
  NAND U5673 ( .A(n3615), .B(n3614), .Z(n3619) );
  NAND U5674 ( .A(n3617), .B(n3616), .Z(n3618) );
  AND U5675 ( .A(n3619), .B(n3618), .Z(n5034) );
  NAND U5676 ( .A(n3621), .B(n3620), .Z(n3625) );
  NAND U5677 ( .A(n3623), .B(n3622), .Z(n3624) );
  NAND U5678 ( .A(n3625), .B(n3624), .Z(n5033) );
  XNOR U5679 ( .A(n5034), .B(n5033), .Z(n5035) );
  XOR U5680 ( .A(n5036), .B(n5035), .Z(n5180) );
  XOR U5681 ( .A(n5181), .B(n5180), .Z(n5182) );
  XOR U5682 ( .A(n5183), .B(n5182), .Z(n5228) );
  NAND U5683 ( .A(n3627), .B(n3626), .Z(n3631) );
  NAND U5684 ( .A(n3629), .B(n3628), .Z(n3630) );
  AND U5685 ( .A(n3631), .B(n3630), .Z(n5229) );
  NAND U5686 ( .A(n3633), .B(n3632), .Z(n3637) );
  NAND U5687 ( .A(n3635), .B(n3634), .Z(n3636) );
  AND U5688 ( .A(n3637), .B(n3636), .Z(n5230) );
  XNOR U5689 ( .A(n5231), .B(n5230), .Z(n5234) );
  NAND U5690 ( .A(n3639), .B(n3638), .Z(n3643) );
  NAND U5691 ( .A(n3641), .B(n3640), .Z(n3642) );
  AND U5692 ( .A(n3643), .B(n3642), .Z(n5319) );
  NAND U5693 ( .A(n3645), .B(n3644), .Z(n3649) );
  NAND U5694 ( .A(n3647), .B(n3646), .Z(n3648) );
  AND U5695 ( .A(n3649), .B(n3648), .Z(n5320) );
  NAND U5696 ( .A(n3651), .B(n3650), .Z(n3655) );
  NAND U5697 ( .A(n3653), .B(n3652), .Z(n3654) );
  AND U5698 ( .A(n3655), .B(n3654), .Z(n5321) );
  XOR U5699 ( .A(n5322), .B(n5321), .Z(n5243) );
  NAND U5700 ( .A(n3657), .B(n3656), .Z(n3661) );
  NAND U5701 ( .A(n3659), .B(n3658), .Z(n3660) );
  NAND U5702 ( .A(n3661), .B(n3660), .Z(n5241) );
  NAND U5703 ( .A(n3663), .B(n3662), .Z(n3667) );
  NAND U5704 ( .A(n3665), .B(n3664), .Z(n3666) );
  AND U5705 ( .A(n3667), .B(n3666), .Z(n5142) );
  NAND U5706 ( .A(n3669), .B(n3668), .Z(n3673) );
  NAND U5707 ( .A(n3671), .B(n3670), .Z(n3672) );
  AND U5708 ( .A(n3673), .B(n3672), .Z(n5143) );
  NAND U5709 ( .A(n3675), .B(n3674), .Z(n3679) );
  NAND U5710 ( .A(n3677), .B(n3676), .Z(n3678) );
  AND U5711 ( .A(n3679), .B(n3678), .Z(n5144) );
  XNOR U5712 ( .A(n5145), .B(n5144), .Z(n5240) );
  XOR U5713 ( .A(n5243), .B(n5242), .Z(n4680) );
  XNOR U5714 ( .A(n4681), .B(n4680), .Z(n4682) );
  XNOR U5715 ( .A(n4683), .B(n4682), .Z(n5369) );
  NANDN U5716 ( .A(n3681), .B(n3680), .Z(n3685) );
  NANDN U5717 ( .A(n3683), .B(n3682), .Z(n3684) );
  AND U5718 ( .A(n3685), .B(n3684), .Z(n5005) );
  XNOR U5719 ( .A(n5004), .B(n5003), .Z(n3692) );
  XOR U5720 ( .A(n5005), .B(n3692), .Z(n4693) );
  NANDN U5721 ( .A(n3694), .B(n3693), .Z(n3698) );
  NAND U5722 ( .A(n3696), .B(n3695), .Z(n3697) );
  NAND U5723 ( .A(n3698), .B(n3697), .Z(n4799) );
  XNOR U5724 ( .A(n4797), .B(n4796), .Z(n4798) );
  XNOR U5725 ( .A(n4693), .B(n4692), .Z(n4695) );
  NANDN U5726 ( .A(n3706), .B(n3705), .Z(n3710) );
  NANDN U5727 ( .A(n3708), .B(n3707), .Z(n3709) );
  AND U5728 ( .A(n3710), .B(n3709), .Z(n4694) );
  XOR U5729 ( .A(n4695), .B(n4694), .Z(n4833) );
  NAND U5730 ( .A(n3712), .B(n3711), .Z(n3716) );
  NAND U5731 ( .A(n3714), .B(n3713), .Z(n3715) );
  NAND U5732 ( .A(n3716), .B(n3715), .Z(n4885) );
  NAND U5733 ( .A(n3718), .B(n3717), .Z(n3722) );
  NANDN U5734 ( .A(n3720), .B(n3719), .Z(n3721) );
  NAND U5735 ( .A(n3722), .B(n3721), .Z(n4883) );
  NAND U5736 ( .A(n3724), .B(n3723), .Z(n3728) );
  NAND U5737 ( .A(n3726), .B(n3725), .Z(n3727) );
  NAND U5738 ( .A(n3728), .B(n3727), .Z(n4882) );
  NAND U5739 ( .A(n3730), .B(n3729), .Z(n3734) );
  NAND U5740 ( .A(n3732), .B(n3731), .Z(n3733) );
  AND U5741 ( .A(n3734), .B(n3733), .Z(n4932) );
  NAND U5742 ( .A(n3739), .B(n3738), .Z(n3745) );
  AND U5743 ( .A(n3741), .B(n3740), .Z(n3743) );
  OR U5744 ( .A(n3743), .B(n3742), .Z(n3744) );
  AND U5745 ( .A(n3745), .B(n3744), .Z(n4930) );
  XNOR U5746 ( .A(n4931), .B(n4930), .Z(n3746) );
  XNOR U5747 ( .A(n4932), .B(n3746), .Z(n4947) );
  NANDN U5748 ( .A(n3748), .B(n3747), .Z(n3752) );
  NANDN U5749 ( .A(n3750), .B(n3749), .Z(n3751) );
  NAND U5750 ( .A(n3752), .B(n3751), .Z(n5139) );
  NAND U5751 ( .A(n3754), .B(n3753), .Z(n3758) );
  NANDN U5752 ( .A(n3756), .B(n3755), .Z(n3757) );
  NAND U5753 ( .A(n3758), .B(n3757), .Z(n5137) );
  NANDN U5754 ( .A(n3760), .B(n3759), .Z(n3764) );
  NAND U5755 ( .A(n3762), .B(n3761), .Z(n3763) );
  NAND U5756 ( .A(n3764), .B(n3763), .Z(n5136) );
  XOR U5757 ( .A(n4947), .B(n4946), .Z(n4949) );
  XOR U5758 ( .A(n4948), .B(n4949), .Z(n4834) );
  XNOR U5759 ( .A(n4834), .B(n4832), .Z(n3768) );
  XOR U5760 ( .A(n4833), .B(n3768), .Z(n5345) );
  NAND U5761 ( .A(n3770), .B(n3769), .Z(n3774) );
  NAND U5762 ( .A(n3772), .B(n3771), .Z(n3773) );
  AND U5763 ( .A(n3774), .B(n3773), .Z(n4972) );
  XNOR U5764 ( .A(n4971), .B(n4970), .Z(n3781) );
  XOR U5765 ( .A(n4972), .B(n3781), .Z(n5343) );
  NAND U5766 ( .A(n3783), .B(n3782), .Z(n3787) );
  NAND U5767 ( .A(n3785), .B(n3784), .Z(n3786) );
  AND U5768 ( .A(n3787), .B(n3786), .Z(n4959) );
  NAND U5769 ( .A(n3789), .B(n3788), .Z(n3793) );
  NAND U5770 ( .A(n3791), .B(n3790), .Z(n3792) );
  AND U5771 ( .A(n3793), .B(n3792), .Z(n4756) );
  NANDN U5772 ( .A(n3795), .B(n3794), .Z(n3799) );
  NAND U5773 ( .A(n3797), .B(n3796), .Z(n3798) );
  AND U5774 ( .A(n3799), .B(n3798), .Z(n4754) );
  NAND U5775 ( .A(n3801), .B(n3800), .Z(n3805) );
  NAND U5776 ( .A(n3803), .B(n3802), .Z(n3804) );
  NAND U5777 ( .A(n3805), .B(n3804), .Z(n4753) );
  XNOR U5778 ( .A(n4754), .B(n4753), .Z(n4755) );
  XNOR U5779 ( .A(n4756), .B(n4755), .Z(n4958) );
  XOR U5780 ( .A(n4959), .B(n4958), .Z(n4960) );
  NAND U5781 ( .A(n3807), .B(n3806), .Z(n3811) );
  NAND U5782 ( .A(n3809), .B(n3808), .Z(n3810) );
  AND U5783 ( .A(n3811), .B(n3810), .Z(n4961) );
  NAND U5784 ( .A(n3813), .B(n3812), .Z(n3817) );
  NAND U5785 ( .A(n3815), .B(n3814), .Z(n3816) );
  NAND U5786 ( .A(n3817), .B(n3816), .Z(n5048) );
  NAND U5787 ( .A(n3819), .B(n3818), .Z(n3823) );
  NAND U5788 ( .A(n3821), .B(n3820), .Z(n3822) );
  NAND U5789 ( .A(n3823), .B(n3822), .Z(n5046) );
  NAND U5790 ( .A(n3825), .B(n3824), .Z(n3829) );
  NAND U5791 ( .A(n3827), .B(n3826), .Z(n3828) );
  NAND U5792 ( .A(n3829), .B(n3828), .Z(n5045) );
  NAND U5793 ( .A(n3831), .B(n3830), .Z(n3835) );
  NAND U5794 ( .A(n3833), .B(n3832), .Z(n3834) );
  NAND U5795 ( .A(n3835), .B(n3834), .Z(n4866) );
  NAND U5796 ( .A(n3837), .B(n3836), .Z(n3841) );
  NAND U5797 ( .A(n3839), .B(n3838), .Z(n3840) );
  NAND U5798 ( .A(n3841), .B(n3840), .Z(n4865) );
  XOR U5799 ( .A(n4868), .B(n4867), .Z(n4897) );
  NANDN U5800 ( .A(n3843), .B(n3842), .Z(n3847) );
  NANDN U5801 ( .A(n3845), .B(n3844), .Z(n3846) );
  NAND U5802 ( .A(n3847), .B(n3846), .Z(n5285) );
  NANDN U5803 ( .A(n3849), .B(n3848), .Z(n3853) );
  NAND U5804 ( .A(n3851), .B(n3850), .Z(n3852) );
  AND U5805 ( .A(n3853), .B(n3852), .Z(n5282) );
  NANDN U5806 ( .A(oglobal[1]), .B(n3854), .Z(n3858) );
  NAND U5807 ( .A(n3856), .B(n3855), .Z(n3857) );
  AND U5808 ( .A(n3858), .B(n3857), .Z(n5283) );
  NANDN U5809 ( .A(n3860), .B(n3859), .Z(n3864) );
  NAND U5810 ( .A(n3862), .B(n3861), .Z(n3863) );
  NAND U5811 ( .A(n3864), .B(n3863), .Z(n4879) );
  NANDN U5812 ( .A(n3866), .B(n3865), .Z(n3870) );
  NAND U5813 ( .A(n3868), .B(n3867), .Z(n3869) );
  NAND U5814 ( .A(n3870), .B(n3869), .Z(n4877) );
  XNOR U5815 ( .A(oglobal[2]), .B(n4877), .Z(n4878) );
  XOR U5816 ( .A(n4894), .B(n4895), .Z(n4896) );
  XNOR U5817 ( .A(n4897), .B(n4896), .Z(n5199) );
  NANDN U5818 ( .A(n3872), .B(n3871), .Z(n3876) );
  NAND U5819 ( .A(n3874), .B(n3873), .Z(n3875) );
  AND U5820 ( .A(n3876), .B(n3875), .Z(n5198) );
  NAND U5821 ( .A(n3878), .B(n3877), .Z(n3882) );
  NAND U5822 ( .A(n3880), .B(n3879), .Z(n3881) );
  NAND U5823 ( .A(n3882), .B(n3881), .Z(n4844) );
  NAND U5824 ( .A(n3884), .B(n3883), .Z(n3888) );
  NAND U5825 ( .A(n3886), .B(n3885), .Z(n3887) );
  NAND U5826 ( .A(n3888), .B(n3887), .Z(n4842) );
  NANDN U5827 ( .A(n3890), .B(n3889), .Z(n3894) );
  NAND U5828 ( .A(n3892), .B(n3891), .Z(n3893) );
  NAND U5829 ( .A(n3894), .B(n3893), .Z(n4841) );
  NAND U5830 ( .A(n3896), .B(n3895), .Z(n3900) );
  NAND U5831 ( .A(n3898), .B(n3897), .Z(n3899) );
  NAND U5832 ( .A(n3900), .B(n3899), .Z(n5307) );
  NANDN U5833 ( .A(n3902), .B(n3901), .Z(n3906) );
  NANDN U5834 ( .A(n3904), .B(n3903), .Z(n3905) );
  AND U5835 ( .A(n3906), .B(n3905), .Z(n4862) );
  NAND U5836 ( .A(n3908), .B(n3907), .Z(n3912) );
  NAND U5837 ( .A(n3910), .B(n3909), .Z(n3911) );
  NAND U5838 ( .A(n3912), .B(n3911), .Z(n4860) );
  NANDN U5839 ( .A(n3914), .B(n3913), .Z(n3918) );
  NAND U5840 ( .A(n3916), .B(n3915), .Z(n3917) );
  NAND U5841 ( .A(n3918), .B(n3917), .Z(n4859) );
  XOR U5842 ( .A(n4862), .B(n4861), .Z(n5306) );
  XOR U5843 ( .A(n5308), .B(n5309), .Z(n5200) );
  XNOR U5844 ( .A(n5201), .B(n5200), .Z(n4823) );
  XNOR U5845 ( .A(n4824), .B(n4823), .Z(n4826) );
  NANDN U5846 ( .A(n3920), .B(n3919), .Z(n3924) );
  NAND U5847 ( .A(n3922), .B(n3921), .Z(n3923) );
  NAND U5848 ( .A(n3924), .B(n3923), .Z(n5133) );
  NANDN U5849 ( .A(n3926), .B(n3925), .Z(n3930) );
  NANDN U5850 ( .A(n3928), .B(n3927), .Z(n3929) );
  NAND U5851 ( .A(n3930), .B(n3929), .Z(n5131) );
  NAND U5852 ( .A(n3932), .B(n3931), .Z(n3936) );
  NAND U5853 ( .A(n3934), .B(n3933), .Z(n3935) );
  AND U5854 ( .A(n3936), .B(n3935), .Z(n5102) );
  NAND U5855 ( .A(n3938), .B(n3937), .Z(n3942) );
  NAND U5856 ( .A(n3940), .B(n3939), .Z(n3941) );
  NAND U5857 ( .A(n3942), .B(n3941), .Z(n5100) );
  NANDN U5858 ( .A(n3944), .B(n3943), .Z(n3948) );
  NAND U5859 ( .A(n3946), .B(n3945), .Z(n3947) );
  NAND U5860 ( .A(n3948), .B(n3947), .Z(n5099) );
  XOR U5861 ( .A(n5102), .B(n5101), .Z(n5130) );
  NAND U5862 ( .A(n3950), .B(n3949), .Z(n3954) );
  NAND U5863 ( .A(n3952), .B(n3951), .Z(n3953) );
  AND U5864 ( .A(n3954), .B(n3953), .Z(n4765) );
  NAND U5865 ( .A(n3956), .B(n3955), .Z(n3960) );
  NAND U5866 ( .A(n3958), .B(n3957), .Z(n3959) );
  AND U5867 ( .A(n3960), .B(n3959), .Z(n4763) );
  NAND U5868 ( .A(n3962), .B(n3961), .Z(n3966) );
  NAND U5869 ( .A(n3964), .B(n3963), .Z(n3965) );
  NAND U5870 ( .A(n3966), .B(n3965), .Z(n4762) );
  XNOR U5871 ( .A(n4763), .B(n4762), .Z(n4764) );
  XOR U5872 ( .A(n4765), .B(n4764), .Z(n4981) );
  NANDN U5873 ( .A(n3968), .B(n3967), .Z(n3972) );
  NAND U5874 ( .A(n3970), .B(n3969), .Z(n3971) );
  NAND U5875 ( .A(n3972), .B(n3971), .Z(n4980) );
  NAND U5876 ( .A(n3974), .B(n3973), .Z(n3978) );
  NAND U5877 ( .A(n3976), .B(n3975), .Z(n3977) );
  AND U5878 ( .A(n3978), .B(n3977), .Z(n5297) );
  NAND U5879 ( .A(n3980), .B(n3979), .Z(n3984) );
  NAND U5880 ( .A(n3982), .B(n3981), .Z(n3983) );
  NAND U5881 ( .A(n3984), .B(n3983), .Z(n5295) );
  NAND U5882 ( .A(n3986), .B(n3985), .Z(n3990) );
  NAND U5883 ( .A(n3988), .B(n3987), .Z(n3989) );
  NAND U5884 ( .A(n3990), .B(n3989), .Z(n5294) );
  XOR U5885 ( .A(n5297), .B(n5296), .Z(n4979) );
  XNOR U5886 ( .A(n4981), .B(n4982), .Z(n5187) );
  NANDN U5887 ( .A(n3992), .B(n3991), .Z(n3996) );
  NANDN U5888 ( .A(n3994), .B(n3993), .Z(n3995) );
  AND U5889 ( .A(n3996), .B(n3995), .Z(n5127) );
  NAND U5890 ( .A(n3998), .B(n3997), .Z(n4002) );
  NAND U5891 ( .A(n4000), .B(n3999), .Z(n4001) );
  NAND U5892 ( .A(n4002), .B(n4001), .Z(n5125) );
  NAND U5893 ( .A(n4004), .B(n4003), .Z(n4008) );
  NAND U5894 ( .A(n4006), .B(n4005), .Z(n4007) );
  AND U5895 ( .A(n4008), .B(n4007), .Z(n5090) );
  NAND U5896 ( .A(n4010), .B(n4009), .Z(n4014) );
  NAND U5897 ( .A(n4012), .B(n4011), .Z(n4013) );
  NAND U5898 ( .A(n4014), .B(n4013), .Z(n5088) );
  NAND U5899 ( .A(n4016), .B(n4015), .Z(n4020) );
  NAND U5900 ( .A(n4018), .B(n4017), .Z(n4019) );
  NAND U5901 ( .A(n4020), .B(n4019), .Z(n5087) );
  XOR U5902 ( .A(n5090), .B(n5089), .Z(n5124) );
  XOR U5903 ( .A(n5127), .B(n5126), .Z(n5186) );
  XOR U5904 ( .A(n5187), .B(n5186), .Z(n5189) );
  XOR U5905 ( .A(n5188), .B(n5189), .Z(n4825) );
  XNOR U5906 ( .A(n4826), .B(n4825), .Z(n5344) );
  XOR U5907 ( .A(n5345), .B(n5346), .Z(n5368) );
  XOR U5908 ( .A(n5369), .B(n5368), .Z(n5370) );
  XOR U5909 ( .A(n5371), .B(n5370), .Z(n5351) );
  NAND U5910 ( .A(n4022), .B(n4021), .Z(n4026) );
  NAND U5911 ( .A(n4024), .B(n4023), .Z(n4025) );
  AND U5912 ( .A(n4026), .B(n4025), .Z(n5333) );
  NAND U5913 ( .A(n4031), .B(n4030), .Z(n4037) );
  AND U5914 ( .A(n4033), .B(n4032), .Z(n4035) );
  OR U5915 ( .A(n4035), .B(n4034), .Z(n4036) );
  AND U5916 ( .A(n4037), .B(n4036), .Z(n5331) );
  XNOR U5917 ( .A(n5332), .B(n5331), .Z(n5334) );
  NANDN U5918 ( .A(n4039), .B(n4038), .Z(n4043) );
  NAND U5919 ( .A(n4041), .B(n4040), .Z(n4042) );
  NAND U5920 ( .A(n4043), .B(n4042), .Z(n5327) );
  NAND U5921 ( .A(n4044), .B(n4045), .Z(n4050) );
  ANDN U5922 ( .B(n4046), .A(n4045), .Z(n4048) );
  NANDN U5923 ( .A(n4048), .B(n4047), .Z(n4049) );
  AND U5924 ( .A(n4050), .B(n4049), .Z(n5326) );
  NAND U5925 ( .A(n4052), .B(n4051), .Z(n4056) );
  NAND U5926 ( .A(n4054), .B(n4053), .Z(n4055) );
  AND U5927 ( .A(n4056), .B(n4055), .Z(n5261) );
  NAND U5928 ( .A(n4058), .B(n4057), .Z(n4062) );
  NAND U5929 ( .A(n4060), .B(n4059), .Z(n4061) );
  NAND U5930 ( .A(n4062), .B(n4061), .Z(n5259) );
  NAND U5931 ( .A(n4064), .B(n4063), .Z(n4068) );
  NAND U5932 ( .A(n4066), .B(n4065), .Z(n4067) );
  NAND U5933 ( .A(n4068), .B(n4067), .Z(n5258) );
  XOR U5934 ( .A(n5261), .B(n5260), .Z(n4929) );
  NAND U5935 ( .A(n4073), .B(n4072), .Z(n4077) );
  NAND U5936 ( .A(n4075), .B(n4074), .Z(n4076) );
  NAND U5937 ( .A(n4077), .B(n4076), .Z(n5255) );
  NANDN U5938 ( .A(n4081), .B(n4082), .Z(n4086) );
  NANDN U5939 ( .A(n4082), .B(n4081), .Z(n4084) );
  NAND U5940 ( .A(n4084), .B(n4083), .Z(n4085) );
  AND U5941 ( .A(n4086), .B(n4085), .Z(n5253) );
  XOR U5942 ( .A(n4927), .B(n4928), .Z(n4087) );
  XNOR U5943 ( .A(n4929), .B(n4087), .Z(n5223) );
  NAND U5944 ( .A(n4089), .B(n4088), .Z(n4093) );
  NAND U5945 ( .A(n4091), .B(n4090), .Z(n4092) );
  AND U5946 ( .A(n4093), .B(n4092), .Z(n5222) );
  NAND U5947 ( .A(n4095), .B(n4094), .Z(n4099) );
  NAND U5948 ( .A(n4097), .B(n4096), .Z(n4098) );
  NAND U5949 ( .A(n4099), .B(n4098), .Z(n5165) );
  NAND U5950 ( .A(n4101), .B(n4100), .Z(n4105) );
  NAND U5951 ( .A(n4103), .B(n4102), .Z(n4104) );
  NAND U5952 ( .A(n4105), .B(n4104), .Z(n5163) );
  NAND U5953 ( .A(n4107), .B(n4106), .Z(n4111) );
  NAND U5954 ( .A(n4109), .B(n4108), .Z(n4110) );
  NAND U5955 ( .A(n4111), .B(n4110), .Z(n5162) );
  NAND U5956 ( .A(n4113), .B(n4112), .Z(n4117) );
  NAND U5957 ( .A(n4115), .B(n4114), .Z(n4116) );
  NAND U5958 ( .A(n4117), .B(n4116), .Z(n5072) );
  NAND U5959 ( .A(n4119), .B(n4118), .Z(n4123) );
  NAND U5960 ( .A(n4121), .B(n4120), .Z(n4122) );
  NAND U5961 ( .A(n4123), .B(n4122), .Z(n5070) );
  NAND U5962 ( .A(n4125), .B(n4124), .Z(n4129) );
  NAND U5963 ( .A(n4127), .B(n4126), .Z(n4128) );
  NAND U5964 ( .A(n4129), .B(n4128), .Z(n5069) );
  NAND U5965 ( .A(n4131), .B(n4130), .Z(n4135) );
  NAND U5966 ( .A(n4133), .B(n4132), .Z(n4134) );
  NAND U5967 ( .A(n4135), .B(n4134), .Z(n5064) );
  NAND U5968 ( .A(n4137), .B(n4136), .Z(n4141) );
  NAND U5969 ( .A(n4139), .B(n4138), .Z(n4140) );
  NAND U5970 ( .A(n4141), .B(n4140), .Z(n5063) );
  NAND U5971 ( .A(n4143), .B(n4142), .Z(n4147) );
  NAND U5972 ( .A(n4145), .B(n4144), .Z(n4146) );
  AND U5973 ( .A(n4147), .B(n4146), .Z(n5065) );
  XNOR U5974 ( .A(n5066), .B(n5065), .Z(n4888) );
  XOR U5975 ( .A(n4889), .B(n4888), .Z(n4891) );
  XOR U5976 ( .A(n4890), .B(n4891), .Z(n5224) );
  XNOR U5977 ( .A(n5225), .B(n5224), .Z(n5121) );
  NAND U5978 ( .A(n4156), .B(n4155), .Z(n4160) );
  NAND U5979 ( .A(n4158), .B(n4157), .Z(n4159) );
  NAND U5980 ( .A(n4160), .B(n4159), .Z(n5291) );
  NAND U5981 ( .A(n4162), .B(n4161), .Z(n4166) );
  NAND U5982 ( .A(n4164), .B(n4163), .Z(n4165) );
  NAND U5983 ( .A(n4166), .B(n4165), .Z(n5289) );
  NANDN U5984 ( .A(n4168), .B(n4167), .Z(n4172) );
  NAND U5985 ( .A(n4170), .B(n4169), .Z(n4171) );
  NAND U5986 ( .A(n4172), .B(n4171), .Z(n5288) );
  NAND U5987 ( .A(n4174), .B(n4173), .Z(n4180) );
  AND U5988 ( .A(n4176), .B(n4175), .Z(n4178) );
  OR U5989 ( .A(n4178), .B(n4177), .Z(n4179) );
  AND U5990 ( .A(n4180), .B(n4179), .Z(n4974) );
  NAND U5991 ( .A(n4182), .B(n4181), .Z(n4186) );
  NAND U5992 ( .A(n4184), .B(n4183), .Z(n4185) );
  NAND U5993 ( .A(n4186), .B(n4185), .Z(n5170) );
  XNOR U5994 ( .A(n5169), .B(n5168), .Z(n5171) );
  XOR U5995 ( .A(n5170), .B(n5171), .Z(n4973) );
  XNOR U5996 ( .A(n4974), .B(n4973), .Z(n4976) );
  XOR U5997 ( .A(n4975), .B(n4976), .Z(n5216) );
  XOR U5998 ( .A(n5217), .B(n5216), .Z(n5219) );
  NAND U5999 ( .A(n4194), .B(n4193), .Z(n4198) );
  NAND U6000 ( .A(n4196), .B(n4195), .Z(n4197) );
  AND U6001 ( .A(n4198), .B(n4197), .Z(n5218) );
  XNOR U6002 ( .A(n5219), .B(n5218), .Z(n5118) );
  XNOR U6003 ( .A(n5119), .B(n5118), .Z(n5120) );
  XOR U6004 ( .A(n5326), .B(n5325), .Z(n5328) );
  XOR U6005 ( .A(n5327), .B(n5328), .Z(n5362) );
  NAND U6006 ( .A(n4200), .B(n4199), .Z(n4204) );
  NAND U6007 ( .A(n4202), .B(n4201), .Z(n4203) );
  AND U6008 ( .A(n4204), .B(n4203), .Z(n5028) );
  NAND U6009 ( .A(n4206), .B(n4205), .Z(n4210) );
  NAND U6010 ( .A(n4208), .B(n4207), .Z(n4209) );
  NAND U6011 ( .A(n4210), .B(n4209), .Z(n5273) );
  NAND U6012 ( .A(n4212), .B(n4211), .Z(n4216) );
  NAND U6013 ( .A(n4214), .B(n4213), .Z(n4215) );
  NAND U6014 ( .A(n4216), .B(n4215), .Z(n5271) );
  NANDN U6015 ( .A(n4218), .B(n4217), .Z(n4222) );
  NAND U6016 ( .A(n4220), .B(n4219), .Z(n4221) );
  NAND U6017 ( .A(n4222), .B(n4221), .Z(n5270) );
  NAND U6018 ( .A(n4224), .B(n4223), .Z(n4228) );
  NAND U6019 ( .A(n4226), .B(n4225), .Z(n4227) );
  AND U6020 ( .A(n4228), .B(n4227), .Z(n4773) );
  NANDN U6021 ( .A(n4230), .B(n4229), .Z(n4234) );
  NAND U6022 ( .A(n4232), .B(n4231), .Z(n4233) );
  NAND U6023 ( .A(n4234), .B(n4233), .Z(n4772) );
  NAND U6024 ( .A(n4236), .B(n4235), .Z(n4240) );
  NAND U6025 ( .A(n4238), .B(n4237), .Z(n4239) );
  AND U6026 ( .A(n4240), .B(n4239), .Z(n4771) );
  XOR U6027 ( .A(n4772), .B(n4771), .Z(n4241) );
  XNOR U6028 ( .A(n4773), .B(n4241), .Z(n4780) );
  NAND U6029 ( .A(n4243), .B(n4242), .Z(n4247) );
  NAND U6030 ( .A(n4245), .B(n4244), .Z(n4246) );
  AND U6031 ( .A(n4247), .B(n4246), .Z(n4781) );
  XNOR U6032 ( .A(n4780), .B(n4781), .Z(n4783) );
  XOR U6033 ( .A(n4782), .B(n4783), .Z(n5027) );
  XOR U6034 ( .A(n5028), .B(n5027), .Z(n5030) );
  NAND U6035 ( .A(n4249), .B(n4248), .Z(n4253) );
  NAND U6036 ( .A(n4251), .B(n4250), .Z(n4252) );
  NAND U6037 ( .A(n4253), .B(n4252), .Z(n5084) );
  NANDN U6038 ( .A(n4255), .B(n4254), .Z(n4259) );
  NANDN U6039 ( .A(n4257), .B(n4256), .Z(n4258) );
  NAND U6040 ( .A(n4259), .B(n4258), .Z(n5082) );
  NAND U6041 ( .A(n4261), .B(n4260), .Z(n4265) );
  NAND U6042 ( .A(n4263), .B(n4262), .Z(n4264) );
  AND U6043 ( .A(n4265), .B(n4264), .Z(n4915) );
  NAND U6044 ( .A(n4267), .B(n4266), .Z(n4271) );
  NAND U6045 ( .A(n4269), .B(n4268), .Z(n4270) );
  AND U6046 ( .A(n4271), .B(n4270), .Z(n4913) );
  NAND U6047 ( .A(n4273), .B(n4272), .Z(n4277) );
  NAND U6048 ( .A(n4275), .B(n4274), .Z(n4276) );
  NAND U6049 ( .A(n4277), .B(n4276), .Z(n4912) );
  XNOR U6050 ( .A(n4913), .B(n4912), .Z(n4914) );
  XOR U6051 ( .A(n4915), .B(n4914), .Z(n5081) );
  XNOR U6052 ( .A(n5030), .B(n5029), .Z(n5018) );
  NAND U6053 ( .A(n4279), .B(n4278), .Z(n4283) );
  NAND U6054 ( .A(n4281), .B(n4280), .Z(n4282) );
  AND U6055 ( .A(n4283), .B(n4282), .Z(n5213) );
  NANDN U6056 ( .A(n4285), .B(n4284), .Z(n4289) );
  NANDN U6057 ( .A(n4287), .B(n4286), .Z(n4288) );
  AND U6058 ( .A(n4289), .B(n4288), .Z(n5211) );
  NANDN U6059 ( .A(n4291), .B(n4290), .Z(n4295) );
  NAND U6060 ( .A(n4293), .B(n4292), .Z(n4294) );
  NAND U6061 ( .A(n4295), .B(n4294), .Z(n5042) );
  NAND U6062 ( .A(n4297), .B(n4296), .Z(n4301) );
  NAND U6063 ( .A(n4299), .B(n4298), .Z(n4300) );
  NAND U6064 ( .A(n4301), .B(n4300), .Z(n5040) );
  NANDN U6065 ( .A(n4303), .B(n4302), .Z(n4307) );
  NAND U6066 ( .A(n4305), .B(n4304), .Z(n4306) );
  NAND U6067 ( .A(n4307), .B(n4306), .Z(n5039) );
  NANDN U6068 ( .A(n4309), .B(n4308), .Z(n4313) );
  NAND U6069 ( .A(n4311), .B(n4310), .Z(n4312) );
  AND U6070 ( .A(n4313), .B(n4312), .Z(n4699) );
  NAND U6071 ( .A(n4315), .B(n4314), .Z(n4319) );
  NAND U6072 ( .A(n4317), .B(n4316), .Z(n4318) );
  AND U6073 ( .A(n4319), .B(n4318), .Z(n4811) );
  NANDN U6074 ( .A(n4321), .B(n4320), .Z(n4325) );
  NAND U6075 ( .A(n4323), .B(n4322), .Z(n4324) );
  NAND U6076 ( .A(n4325), .B(n4324), .Z(n4809) );
  NANDN U6077 ( .A(n4327), .B(n4326), .Z(n4331) );
  NAND U6078 ( .A(n4329), .B(n4328), .Z(n4330) );
  NAND U6079 ( .A(n4331), .B(n4330), .Z(n4808) );
  XOR U6080 ( .A(n4811), .B(n4810), .Z(n4698) );
  XNOR U6081 ( .A(n4699), .B(n4698), .Z(n4701) );
  XOR U6082 ( .A(n4700), .B(n4701), .Z(n5210) );
  XOR U6083 ( .A(n5211), .B(n5210), .Z(n5212) );
  XOR U6084 ( .A(n5213), .B(n5212), .Z(n5016) );
  NANDN U6085 ( .A(n4333), .B(n4332), .Z(n4337) );
  NANDN U6086 ( .A(n4335), .B(n4334), .Z(n4336) );
  AND U6087 ( .A(n4337), .B(n4336), .Z(n5022) );
  NANDN U6088 ( .A(n4339), .B(n4338), .Z(n4343) );
  NANDN U6089 ( .A(n4341), .B(n4340), .Z(n4342) );
  NAND U6090 ( .A(n4343), .B(n4342), .Z(n5096) );
  NANDN U6091 ( .A(n4345), .B(n4344), .Z(n4349) );
  NAND U6092 ( .A(n4347), .B(n4346), .Z(n4348) );
  NAND U6093 ( .A(n4349), .B(n4348), .Z(n5094) );
  NANDN U6094 ( .A(n4351), .B(n4350), .Z(n4355) );
  NAND U6095 ( .A(n4353), .B(n4352), .Z(n4354) );
  NAND U6096 ( .A(n4355), .B(n4354), .Z(n5093) );
  NANDN U6097 ( .A(n4357), .B(n4356), .Z(n4361) );
  NAND U6098 ( .A(n4359), .B(n4358), .Z(n4360) );
  NAND U6099 ( .A(n4361), .B(n4360), .Z(n4770) );
  NAND U6100 ( .A(n4363), .B(n4362), .Z(n4367) );
  NAND U6101 ( .A(n4365), .B(n4364), .Z(n4366) );
  NAND U6102 ( .A(n4367), .B(n4366), .Z(n4769) );
  NANDN U6103 ( .A(n4369), .B(n4368), .Z(n4373) );
  NAND U6104 ( .A(n4371), .B(n4370), .Z(n4372) );
  AND U6105 ( .A(n4373), .B(n4372), .Z(n4768) );
  NANDN U6106 ( .A(n4375), .B(n4374), .Z(n4379) );
  NANDN U6107 ( .A(n4377), .B(n4376), .Z(n4378) );
  AND U6108 ( .A(n4379), .B(n4378), .Z(n4742) );
  XNOR U6109 ( .A(n4741), .B(n4742), .Z(n4744) );
  XOR U6110 ( .A(n4743), .B(n4744), .Z(n5021) );
  XOR U6111 ( .A(n5022), .B(n5021), .Z(n5024) );
  NAND U6112 ( .A(n4381), .B(n4380), .Z(n4385) );
  NAND U6113 ( .A(n4383), .B(n4382), .Z(n4384) );
  NAND U6114 ( .A(n4385), .B(n4384), .Z(n5078) );
  NAND U6115 ( .A(n4387), .B(n4386), .Z(n4391) );
  NAND U6116 ( .A(n4389), .B(n4388), .Z(n4390) );
  NAND U6117 ( .A(n4391), .B(n4390), .Z(n5076) );
  NAND U6118 ( .A(n4393), .B(n4392), .Z(n4397) );
  NAND U6119 ( .A(n4395), .B(n4394), .Z(n4396) );
  NAND U6120 ( .A(n4397), .B(n4396), .Z(n5075) );
  NANDN U6121 ( .A(n4399), .B(n4398), .Z(n4403) );
  NANDN U6122 ( .A(n4401), .B(n4400), .Z(n4402) );
  AND U6123 ( .A(n4403), .B(n4402), .Z(n4818) );
  NAND U6124 ( .A(n4405), .B(n4404), .Z(n4409) );
  NAND U6125 ( .A(n4407), .B(n4406), .Z(n4408) );
  AND U6126 ( .A(n4409), .B(n4408), .Z(n4874) );
  NAND U6127 ( .A(n4411), .B(n4410), .Z(n4415) );
  NAND U6128 ( .A(n4413), .B(n4412), .Z(n4414) );
  NAND U6129 ( .A(n4415), .B(n4414), .Z(n4872) );
  NAND U6130 ( .A(n4417), .B(n4416), .Z(n4421) );
  NAND U6131 ( .A(n4419), .B(n4418), .Z(n4420) );
  NAND U6132 ( .A(n4421), .B(n4420), .Z(n4871) );
  XOR U6133 ( .A(n4874), .B(n4873), .Z(n4817) );
  XNOR U6134 ( .A(n4818), .B(n4817), .Z(n4820) );
  XOR U6135 ( .A(n4819), .B(n4820), .Z(n5023) );
  XNOR U6136 ( .A(n5024), .B(n5023), .Z(n5015) );
  XNOR U6137 ( .A(n5016), .B(n5015), .Z(n5017) );
  XNOR U6138 ( .A(n5018), .B(n5017), .Z(n4670) );
  NANDN U6139 ( .A(n4423), .B(n4422), .Z(n4427) );
  NANDN U6140 ( .A(n4425), .B(n4424), .Z(n4426) );
  NAND U6141 ( .A(n4427), .B(n4426), .Z(n5315) );
  NANDN U6142 ( .A(n4429), .B(n4428), .Z(n4433) );
  NAND U6143 ( .A(n4431), .B(n4430), .Z(n4432) );
  NAND U6144 ( .A(n4433), .B(n4432), .Z(n5313) );
  NAND U6145 ( .A(n4435), .B(n4434), .Z(n4439) );
  NAND U6146 ( .A(n4437), .B(n4436), .Z(n4438) );
  NAND U6147 ( .A(n4439), .B(n4438), .Z(n5312) );
  NANDN U6148 ( .A(n4441), .B(n4440), .Z(n4445) );
  NAND U6149 ( .A(n4443), .B(n4442), .Z(n4444) );
  NAND U6150 ( .A(n4445), .B(n4444), .Z(n5267) );
  NAND U6151 ( .A(n4447), .B(n4446), .Z(n4451) );
  NAND U6152 ( .A(n4449), .B(n4448), .Z(n4450) );
  NAND U6153 ( .A(n4451), .B(n4450), .Z(n5265) );
  NAND U6154 ( .A(n4453), .B(n4452), .Z(n4457) );
  NAND U6155 ( .A(n4455), .B(n4454), .Z(n4456) );
  NAND U6156 ( .A(n4457), .B(n4456), .Z(n5264) );
  XOR U6157 ( .A(n4965), .B(n4964), .Z(n4967) );
  NAND U6158 ( .A(n4459), .B(n4458), .Z(n4463) );
  NANDN U6159 ( .A(n4461), .B(n4460), .Z(n4462) );
  NAND U6160 ( .A(n4463), .B(n4462), .Z(n5054) );
  NAND U6161 ( .A(n4465), .B(n4464), .Z(n4469) );
  NAND U6162 ( .A(n4467), .B(n4466), .Z(n4468) );
  NAND U6163 ( .A(n4469), .B(n4468), .Z(n5052) );
  NAND U6164 ( .A(n4471), .B(n4470), .Z(n4475) );
  NAND U6165 ( .A(n4473), .B(n4472), .Z(n4474) );
  NAND U6166 ( .A(n4475), .B(n4474), .Z(n5051) );
  XOR U6167 ( .A(n4967), .B(n4966), .Z(n5012) );
  NAND U6168 ( .A(n4477), .B(n4476), .Z(n4481) );
  NAND U6169 ( .A(n4479), .B(n4478), .Z(n4480) );
  AND U6170 ( .A(n4481), .B(n4480), .Z(n5113) );
  NANDN U6171 ( .A(n4483), .B(n4482), .Z(n4487) );
  NAND U6172 ( .A(n4485), .B(n4484), .Z(n4486) );
  AND U6173 ( .A(n4487), .B(n4486), .Z(n4707) );
  NAND U6174 ( .A(n4489), .B(n4488), .Z(n4493) );
  NAND U6175 ( .A(n4491), .B(n4490), .Z(n4492) );
  AND U6176 ( .A(n4493), .B(n4492), .Z(n4705) );
  NANDN U6177 ( .A(n4495), .B(n4494), .Z(n4499) );
  NANDN U6178 ( .A(n4497), .B(n4496), .Z(n4498) );
  NAND U6179 ( .A(n4499), .B(n4498), .Z(n4704) );
  XNOR U6180 ( .A(n4705), .B(n4704), .Z(n4706) );
  XNOR U6181 ( .A(n4707), .B(n4706), .Z(n5112) );
  XOR U6182 ( .A(n5113), .B(n5112), .Z(n5114) );
  NAND U6183 ( .A(n4501), .B(n4500), .Z(n4505) );
  NAND U6184 ( .A(n4503), .B(n4502), .Z(n4504) );
  AND U6185 ( .A(n4505), .B(n4504), .Z(n5115) );
  NAND U6186 ( .A(n4507), .B(n4506), .Z(n4511) );
  NAND U6187 ( .A(n4509), .B(n4508), .Z(n4510) );
  AND U6188 ( .A(n4511), .B(n4510), .Z(n4838) );
  NAND U6189 ( .A(n4513), .B(n4512), .Z(n4517) );
  NAND U6190 ( .A(n4515), .B(n4514), .Z(n4516) );
  AND U6191 ( .A(n4517), .B(n4516), .Z(n4836) );
  NANDN U6192 ( .A(n4519), .B(n4518), .Z(n4523) );
  NAND U6193 ( .A(n4521), .B(n4520), .Z(n4522) );
  NAND U6194 ( .A(n4523), .B(n4522), .Z(n4835) );
  XNOR U6195 ( .A(n4836), .B(n4835), .Z(n4837) );
  XOR U6196 ( .A(n4838), .B(n4837), .Z(n5059) );
  NANDN U6197 ( .A(n4525), .B(n4524), .Z(n4529) );
  NAND U6198 ( .A(n4527), .B(n4526), .Z(n4528) );
  NAND U6199 ( .A(n4529), .B(n4528), .Z(n5058) );
  NAND U6200 ( .A(n4531), .B(n4530), .Z(n4535) );
  NAND U6201 ( .A(n4533), .B(n4532), .Z(n4534) );
  AND U6202 ( .A(n4535), .B(n4534), .Z(n4903) );
  NAND U6203 ( .A(n4537), .B(n4536), .Z(n4541) );
  NAND U6204 ( .A(n4539), .B(n4538), .Z(n4540) );
  AND U6205 ( .A(n4541), .B(n4540), .Z(n4901) );
  NAND U6206 ( .A(n4543), .B(n4542), .Z(n4547) );
  NAND U6207 ( .A(n4545), .B(n4544), .Z(n4546) );
  NAND U6208 ( .A(n4547), .B(n4546), .Z(n4900) );
  XNOR U6209 ( .A(n4901), .B(n4900), .Z(n4902) );
  XOR U6210 ( .A(n4903), .B(n4902), .Z(n5057) );
  XNOR U6211 ( .A(n5059), .B(n5060), .Z(n5206) );
  NANDN U6212 ( .A(n4549), .B(n4548), .Z(n4553) );
  NAND U6213 ( .A(n4551), .B(n4550), .Z(n4552) );
  NAND U6214 ( .A(n4553), .B(n4552), .Z(n5177) );
  NANDN U6215 ( .A(n4555), .B(n4554), .Z(n4559) );
  NANDN U6216 ( .A(n4557), .B(n4556), .Z(n4558) );
  NAND U6217 ( .A(n4559), .B(n4558), .Z(n5175) );
  NAND U6218 ( .A(n4561), .B(n4560), .Z(n4565) );
  NAND U6219 ( .A(n4563), .B(n4562), .Z(n4564) );
  AND U6220 ( .A(n4565), .B(n4564), .Z(n5249) );
  NAND U6221 ( .A(n4567), .B(n4566), .Z(n4571) );
  NAND U6222 ( .A(n4569), .B(n4568), .Z(n4570) );
  NAND U6223 ( .A(n4571), .B(n4570), .Z(n5247) );
  NAND U6224 ( .A(n4573), .B(n4572), .Z(n4577) );
  NAND U6225 ( .A(n4575), .B(n4574), .Z(n4576) );
  NAND U6226 ( .A(n4577), .B(n4576), .Z(n5246) );
  XOR U6227 ( .A(n5249), .B(n5248), .Z(n5174) );
  NANDN U6228 ( .A(n4579), .B(n4578), .Z(n4583) );
  NANDN U6229 ( .A(n4581), .B(n4580), .Z(n4582) );
  NAND U6230 ( .A(n4583), .B(n4582), .Z(n5204) );
  XOR U6231 ( .A(n5205), .B(n5204), .Z(n5207) );
  XOR U6232 ( .A(n5206), .B(n5207), .Z(n5009) );
  XNOR U6233 ( .A(n5010), .B(n5009), .Z(n5011) );
  XNOR U6234 ( .A(n5012), .B(n5011), .Z(n4669) );
  NANDN U6235 ( .A(n4585), .B(n4584), .Z(n4589) );
  NANDN U6236 ( .A(n4587), .B(n4586), .Z(n4588) );
  AND U6237 ( .A(n4589), .B(n4588), .Z(n4816) );
  NANDN U6238 ( .A(n4594), .B(n4593), .Z(n4598) );
  ANDN U6239 ( .B(n4594), .A(n4593), .Z(n4596) );
  OR U6240 ( .A(n4596), .B(n4595), .Z(n4597) );
  AND U6241 ( .A(n4598), .B(n4597), .Z(n4814) );
  XNOR U6242 ( .A(n4815), .B(n4814), .Z(n4599) );
  XNOR U6243 ( .A(n4816), .B(n4599), .Z(n4942) );
  NANDN U6244 ( .A(n4601), .B(n4600), .Z(n4605) );
  NAND U6245 ( .A(n4603), .B(n4602), .Z(n4604) );
  NAND U6246 ( .A(n4605), .B(n4604), .Z(n4777) );
  NAND U6247 ( .A(n4610), .B(n4609), .Z(n4616) );
  AND U6248 ( .A(n4612), .B(n4611), .Z(n4614) );
  OR U6249 ( .A(n4614), .B(n4613), .Z(n4615) );
  AND U6250 ( .A(n4616), .B(n4615), .Z(n4774) );
  XOR U6251 ( .A(n4775), .B(n4774), .Z(n4776) );
  IV U6252 ( .A(n4939), .Z(n4941) );
  NANDN U6253 ( .A(n4621), .B(n4620), .Z(n4625) );
  NANDN U6254 ( .A(n4623), .B(n4622), .Z(n4624) );
  NAND U6255 ( .A(n4625), .B(n4624), .Z(n4936) );
  XOR U6256 ( .A(n4934), .B(n4933), .Z(n4935) );
  NANDN U6257 ( .A(n4633), .B(n4632), .Z(n4637) );
  NAND U6258 ( .A(n4635), .B(n4634), .Z(n4636) );
  NAND U6259 ( .A(n4637), .B(n4636), .Z(n4988) );
  XNOR U6260 ( .A(n4986), .B(n4985), .Z(n4987) );
  XOR U6261 ( .A(n4717), .B(n4716), .Z(n4719) );
  NANDN U6262 ( .A(n4645), .B(n4644), .Z(n4649) );
  NANDN U6263 ( .A(n4647), .B(n4646), .Z(n4648) );
  NAND U6264 ( .A(n4649), .B(n4648), .Z(n4992) );
  NANDN U6265 ( .A(n4651), .B(n4650), .Z(n4655) );
  NAND U6266 ( .A(n4653), .B(n4652), .Z(n4654) );
  NAND U6267 ( .A(n4655), .B(n4654), .Z(n4991) );
  XOR U6268 ( .A(n4992), .B(n4991), .Z(n4994) );
  NANDN U6269 ( .A(n4657), .B(n4656), .Z(n4661) );
  NANDN U6270 ( .A(n4659), .B(n4658), .Z(n4660) );
  NAND U6271 ( .A(n4661), .B(n4660), .Z(n4993) );
  XOR U6272 ( .A(n4994), .B(n4993), .Z(n4718) );
  XOR U6273 ( .A(n4719), .B(n4718), .Z(n4760) );
  XNOR U6274 ( .A(n4760), .B(n4759), .Z(n4665) );
  XOR U6275 ( .A(n4761), .B(n4665), .Z(n4668) );
  XOR U6276 ( .A(n4669), .B(n4668), .Z(n4671) );
  XOR U6277 ( .A(n4670), .B(n4671), .Z(n5365) );
  XNOR U6278 ( .A(n5364), .B(n5365), .Z(n5350) );
  XNOR U6279 ( .A(n5351), .B(n5350), .Z(n4666) );
  XOR U6280 ( .A(n5349), .B(n4666), .Z(n5354) );
  XOR U6281 ( .A(n5353), .B(n5354), .Z(n4667) );
  XNOR U6282 ( .A(n5355), .B(n4667), .Z(o[2]) );
  NANDN U6283 ( .A(n4669), .B(n4668), .Z(n4673) );
  NANDN U6284 ( .A(n4671), .B(n4670), .Z(n4672) );
  NAND U6285 ( .A(n4673), .B(n4672), .Z(n5395) );
  NANDN U6286 ( .A(n4675), .B(n4674), .Z(n4679) );
  NAND U6287 ( .A(n4677), .B(n4676), .Z(n4678) );
  NAND U6288 ( .A(n4679), .B(n4678), .Z(n5394) );
  NANDN U6289 ( .A(n4681), .B(n4680), .Z(n4685) );
  NANDN U6290 ( .A(n4683), .B(n4682), .Z(n4684) );
  NAND U6291 ( .A(n4685), .B(n4684), .Z(n5393) );
  XOR U6292 ( .A(n5394), .B(n5393), .Z(n5396) );
  XNOR U6293 ( .A(n5395), .B(n5396), .Z(n5724) );
  NAND U6294 ( .A(n4687), .B(n4686), .Z(n4691) );
  NANDN U6295 ( .A(n4689), .B(n4688), .Z(n4690) );
  NAND U6296 ( .A(n4691), .B(n4690), .Z(n5428) );
  NANDN U6297 ( .A(n4693), .B(n4692), .Z(n4697) );
  NAND U6298 ( .A(n4695), .B(n4694), .Z(n4696) );
  AND U6299 ( .A(n4697), .B(n4696), .Z(n5537) );
  NANDN U6300 ( .A(n4699), .B(n4698), .Z(n4703) );
  NAND U6301 ( .A(n4701), .B(n4700), .Z(n4702) );
  AND U6302 ( .A(n4703), .B(n4702), .Z(n5629) );
  NANDN U6303 ( .A(n4705), .B(n4704), .Z(n4709) );
  NANDN U6304 ( .A(n4707), .B(n4706), .Z(n4708) );
  AND U6305 ( .A(n4709), .B(n4708), .Z(n5630) );
  NANDN U6306 ( .A(n4711), .B(n4710), .Z(n4715) );
  NANDN U6307 ( .A(n4713), .B(n4712), .Z(n4714) );
  AND U6308 ( .A(n4715), .B(n4714), .Z(n5632) );
  IV U6309 ( .A(n5534), .Z(n5536) );
  NAND U6310 ( .A(n4717), .B(n4716), .Z(n4721) );
  NAND U6311 ( .A(n4719), .B(n4718), .Z(n4720) );
  AND U6312 ( .A(n4721), .B(n4720), .Z(n5535) );
  XNOR U6313 ( .A(n5536), .B(n5535), .Z(n4722) );
  XNOR U6314 ( .A(n5537), .B(n4722), .Z(n5427) );
  NANDN U6315 ( .A(n4724), .B(n4723), .Z(n4728) );
  NAND U6316 ( .A(n4726), .B(n4725), .Z(n4727) );
  NAND U6317 ( .A(n4728), .B(n4727), .Z(n5426) );
  XOR U6318 ( .A(n5427), .B(n5426), .Z(n5429) );
  XNOR U6319 ( .A(n5428), .B(n5429), .Z(n5390) );
  NANDN U6320 ( .A(n4730), .B(n4729), .Z(n4734) );
  NAND U6321 ( .A(n4732), .B(n4731), .Z(n4733) );
  NAND U6322 ( .A(n4734), .B(n4733), .Z(n5506) );
  NAND U6323 ( .A(n4736), .B(n4735), .Z(n4740) );
  NANDN U6324 ( .A(n4738), .B(n4737), .Z(n4739) );
  NAND U6325 ( .A(n4740), .B(n4739), .Z(n5505) );
  NANDN U6326 ( .A(n4742), .B(n4741), .Z(n4746) );
  NAND U6327 ( .A(n4744), .B(n4743), .Z(n4745) );
  AND U6328 ( .A(n4746), .B(n4745), .Z(n5663) );
  NANDN U6329 ( .A(n4748), .B(n4747), .Z(n4752) );
  NANDN U6330 ( .A(n4750), .B(n4749), .Z(n4751) );
  AND U6331 ( .A(n4752), .B(n4751), .Z(n5664) );
  NANDN U6332 ( .A(n4754), .B(n4753), .Z(n4758) );
  NANDN U6333 ( .A(n4756), .B(n4755), .Z(n4757) );
  AND U6334 ( .A(n4758), .B(n4757), .Z(n5665) );
  XNOR U6335 ( .A(n5666), .B(n5665), .Z(n5504) );
  XOR U6336 ( .A(n5505), .B(n5504), .Z(n5507) );
  XNOR U6337 ( .A(n5506), .B(n5507), .Z(n5423) );
  NANDN U6338 ( .A(n4763), .B(n4762), .Z(n4767) );
  NANDN U6339 ( .A(n4765), .B(n4764), .Z(n4766) );
  AND U6340 ( .A(n4767), .B(n4766), .Z(n5656) );
  XOR U6341 ( .A(n5654), .B(n5653), .Z(n5655) );
  XNOR U6342 ( .A(n5656), .B(n5655), .Z(n5699) );
  OR U6343 ( .A(n4775), .B(n4774), .Z(n4779) );
  NAND U6344 ( .A(n4777), .B(n4776), .Z(n4778) );
  AND U6345 ( .A(n4779), .B(n4778), .Z(n5698) );
  NANDN U6346 ( .A(n4781), .B(n4780), .Z(n4785) );
  NAND U6347 ( .A(n4783), .B(n4782), .Z(n4784) );
  AND U6348 ( .A(n4785), .B(n4784), .Z(n5701) );
  NAND U6349 ( .A(n4789), .B(n4790), .Z(n4795) );
  ANDN U6350 ( .B(n4791), .A(n4790), .Z(n4793) );
  OR U6351 ( .A(n4793), .B(n4792), .Z(n4794) );
  AND U6352 ( .A(n4795), .B(n4794), .Z(n5593) );
  XNOR U6353 ( .A(n5594), .B(n5593), .Z(n5595) );
  NANDN U6354 ( .A(n4797), .B(n4796), .Z(n4801) );
  NAND U6355 ( .A(n4799), .B(n4798), .Z(n4800) );
  AND U6356 ( .A(n4801), .B(n4800), .Z(n5596) );
  NAND U6357 ( .A(n4809), .B(n4808), .Z(n4813) );
  NANDN U6358 ( .A(n4811), .B(n4810), .Z(n4812) );
  AND U6359 ( .A(n4813), .B(n4812), .Z(n5643) );
  XNOR U6360 ( .A(n5644), .B(n5643), .Z(n5705) );
  NANDN U6361 ( .A(n4818), .B(n4817), .Z(n4822) );
  NAND U6362 ( .A(n4820), .B(n4819), .Z(n4821) );
  AND U6363 ( .A(n4822), .B(n4821), .Z(n5707) );
  XOR U6364 ( .A(n5579), .B(n5578), .Z(n5580) );
  XOR U6365 ( .A(n5581), .B(n5580), .Z(n5420) );
  XNOR U6366 ( .A(n5421), .B(n5420), .Z(n5422) );
  NANDN U6367 ( .A(n4824), .B(n4823), .Z(n4828) );
  NAND U6368 ( .A(n4826), .B(n4825), .Z(n4827) );
  NAND U6369 ( .A(n4828), .B(n4827), .Z(n5434) );
  XOR U6370 ( .A(n5433), .B(n5432), .Z(n5435) );
  XNOR U6371 ( .A(n5434), .B(n5435), .Z(n5387) );
  NANDN U6372 ( .A(n4836), .B(n4835), .Z(n4840) );
  NANDN U6373 ( .A(n4838), .B(n4837), .Z(n4839) );
  AND U6374 ( .A(n4840), .B(n4839), .Z(n5568) );
  NAND U6375 ( .A(n4842), .B(n4841), .Z(n4846) );
  NAND U6376 ( .A(n4844), .B(n4843), .Z(n4845) );
  AND U6377 ( .A(n4846), .B(n4845), .Z(n5565) );
  NAND U6378 ( .A(n4848), .B(n4847), .Z(n4852) );
  NAND U6379 ( .A(n4850), .B(n4849), .Z(n4851) );
  AND U6380 ( .A(n4852), .B(n4851), .Z(n5566) );
  XNOR U6381 ( .A(n5568), .B(n5567), .Z(n5602) );
  NAND U6382 ( .A(n4854), .B(n4853), .Z(n4858) );
  NAND U6383 ( .A(n4856), .B(n4855), .Z(n4857) );
  NAND U6384 ( .A(n4858), .B(n4857), .Z(n5600) );
  NAND U6385 ( .A(n4860), .B(n4859), .Z(n4864) );
  NANDN U6386 ( .A(n4862), .B(n4861), .Z(n4863) );
  NAND U6387 ( .A(n4864), .B(n4863), .Z(n5599) );
  NAND U6388 ( .A(n4866), .B(n4865), .Z(n4870) );
  NAND U6389 ( .A(n4868), .B(n4867), .Z(n4869) );
  AND U6390 ( .A(n4870), .B(n4869), .Z(n5608) );
  NAND U6391 ( .A(n4872), .B(n4871), .Z(n4876) );
  NANDN U6392 ( .A(n4874), .B(n4873), .Z(n4875) );
  AND U6393 ( .A(n4876), .B(n4875), .Z(n5605) );
  NANDN U6394 ( .A(oglobal[2]), .B(n4877), .Z(n4881) );
  NAND U6395 ( .A(n4879), .B(n4878), .Z(n4880) );
  AND U6396 ( .A(n4881), .B(n4880), .Z(n5606) );
  XNOR U6397 ( .A(n5608), .B(n5607), .Z(n5670) );
  NAND U6398 ( .A(n4883), .B(n4882), .Z(n4887) );
  NAND U6399 ( .A(n4885), .B(n4884), .Z(n4886) );
  AND U6400 ( .A(n4887), .B(n4886), .Z(n5669) );
  XOR U6401 ( .A(n5672), .B(n5671), .Z(n5512) );
  NAND U6402 ( .A(n4889), .B(n4888), .Z(n4893) );
  NAND U6403 ( .A(n4891), .B(n4890), .Z(n4892) );
  NAND U6404 ( .A(n4893), .B(n4892), .Z(n5477) );
  NAND U6405 ( .A(n4895), .B(n4894), .Z(n4899) );
  NAND U6406 ( .A(n4897), .B(n4896), .Z(n4898) );
  AND U6407 ( .A(n4899), .B(n4898), .Z(n5475) );
  NANDN U6408 ( .A(n4901), .B(n4900), .Z(n4905) );
  NANDN U6409 ( .A(n4903), .B(n4902), .Z(n4904) );
  AND U6410 ( .A(n4905), .B(n4904), .Z(n5465) );
  NAND U6411 ( .A(n4907), .B(n4906), .Z(n4911) );
  NAND U6412 ( .A(n4909), .B(n4908), .Z(n4910) );
  AND U6413 ( .A(n4911), .B(n4910), .Z(n5462) );
  NANDN U6414 ( .A(n4913), .B(n4912), .Z(n4917) );
  NANDN U6415 ( .A(n4915), .B(n4914), .Z(n4916) );
  AND U6416 ( .A(n4917), .B(n4916), .Z(n5463) );
  XOR U6417 ( .A(n5465), .B(n5464), .Z(n5474) );
  XOR U6418 ( .A(n5475), .B(n5474), .Z(n5476) );
  NAND U6419 ( .A(n4919), .B(n4918), .Z(n4923) );
  NAND U6420 ( .A(n4921), .B(n4920), .Z(n4922) );
  NAND U6421 ( .A(n4923), .B(n4922), .Z(n5510) );
  XOR U6422 ( .A(n5512), .B(n5513), .Z(n5417) );
  XNOR U6423 ( .A(n5624), .B(n5623), .Z(n5626) );
  NAND U6424 ( .A(n4934), .B(n4933), .Z(n4938) );
  NAND U6425 ( .A(n4936), .B(n4935), .Z(n4937) );
  AND U6426 ( .A(n4938), .B(n4937), .Z(n5625) );
  XNOR U6427 ( .A(n5626), .B(n5625), .Z(n5445) );
  NAND U6428 ( .A(n4939), .B(n4940), .Z(n4945) );
  ANDN U6429 ( .B(n4941), .A(n4940), .Z(n4943) );
  OR U6430 ( .A(n4943), .B(n4942), .Z(n4944) );
  AND U6431 ( .A(n4945), .B(n4944), .Z(n5444) );
  NAND U6432 ( .A(n4947), .B(n4946), .Z(n4951) );
  NAND U6433 ( .A(n4949), .B(n4948), .Z(n4950) );
  AND U6434 ( .A(n4951), .B(n4950), .Z(n5447) );
  XNOR U6435 ( .A(n5415), .B(n5414), .Z(n5416) );
  NAND U6436 ( .A(n4953), .B(n4952), .Z(n4957) );
  NAND U6437 ( .A(n4955), .B(n4954), .Z(n4956) );
  NAND U6438 ( .A(n4957), .B(n4956), .Z(n5453) );
  NAND U6439 ( .A(n4959), .B(n4958), .Z(n4963) );
  NAND U6440 ( .A(n4961), .B(n4960), .Z(n4962) );
  AND U6441 ( .A(n4963), .B(n4962), .Z(n5450) );
  NAND U6442 ( .A(n4965), .B(n4964), .Z(n4969) );
  NAND U6443 ( .A(n4967), .B(n4966), .Z(n4968) );
  AND U6444 ( .A(n4969), .B(n4968), .Z(n5451) );
  NANDN U6445 ( .A(n4974), .B(n4973), .Z(n4978) );
  NAND U6446 ( .A(n4976), .B(n4975), .Z(n4977) );
  AND U6447 ( .A(n4978), .B(n4977), .Z(n5562) );
  NAND U6448 ( .A(n4980), .B(n4979), .Z(n4984) );
  NAND U6449 ( .A(n4982), .B(n4981), .Z(n4983) );
  AND U6450 ( .A(n4984), .B(n4983), .Z(n5559) );
  NANDN U6451 ( .A(n4986), .B(n4985), .Z(n4990) );
  NAND U6452 ( .A(n4988), .B(n4987), .Z(n4989) );
  AND U6453 ( .A(n4990), .B(n4989), .Z(n5560) );
  XNOR U6454 ( .A(n5562), .B(n5561), .Z(n5678) );
  NAND U6455 ( .A(n4992), .B(n4991), .Z(n4996) );
  NAND U6456 ( .A(n4994), .B(n4993), .Z(n4995) );
  NAND U6457 ( .A(n4996), .B(n4995), .Z(n5676) );
  NANDN U6458 ( .A(n4998), .B(n4997), .Z(n5002) );
  NAND U6459 ( .A(n5000), .B(n4999), .Z(n5001) );
  NAND U6460 ( .A(n5002), .B(n5001), .Z(n5550) );
  XOR U6461 ( .A(n5548), .B(n5547), .Z(n5549) );
  XOR U6462 ( .A(n5682), .B(n5681), .Z(n5683) );
  XOR U6463 ( .A(n5684), .B(n5683), .Z(n5408) );
  NANDN U6464 ( .A(n5010), .B(n5009), .Z(n5014) );
  NANDN U6465 ( .A(n5012), .B(n5011), .Z(n5013) );
  NAND U6466 ( .A(n5014), .B(n5013), .Z(n5530) );
  NANDN U6467 ( .A(n5016), .B(n5015), .Z(n5020) );
  NAND U6468 ( .A(n5018), .B(n5017), .Z(n5019) );
  NAND U6469 ( .A(n5020), .B(n5019), .Z(n5529) );
  NAND U6470 ( .A(n5022), .B(n5021), .Z(n5026) );
  NAND U6471 ( .A(n5024), .B(n5023), .Z(n5025) );
  AND U6472 ( .A(n5026), .B(n5025), .Z(n5590) );
  NAND U6473 ( .A(n5028), .B(n5027), .Z(n5032) );
  NAND U6474 ( .A(n5030), .B(n5029), .Z(n5031) );
  NAND U6475 ( .A(n5032), .B(n5031), .Z(n5588) );
  NANDN U6476 ( .A(n5034), .B(n5033), .Z(n5038) );
  NANDN U6477 ( .A(n5036), .B(n5035), .Z(n5037) );
  AND U6478 ( .A(n5038), .B(n5037), .Z(n5574) );
  NAND U6479 ( .A(n5040), .B(n5039), .Z(n5044) );
  NAND U6480 ( .A(n5042), .B(n5041), .Z(n5043) );
  AND U6481 ( .A(n5044), .B(n5043), .Z(n5571) );
  NAND U6482 ( .A(n5046), .B(n5045), .Z(n5050) );
  NAND U6483 ( .A(n5048), .B(n5047), .Z(n5049) );
  AND U6484 ( .A(n5050), .B(n5049), .Z(n5572) );
  XNOR U6485 ( .A(n5574), .B(n5573), .Z(n5618) );
  NAND U6486 ( .A(n5052), .B(n5051), .Z(n5056) );
  NAND U6487 ( .A(n5054), .B(n5053), .Z(n5055) );
  AND U6488 ( .A(n5056), .B(n5055), .Z(n5617) );
  NAND U6489 ( .A(n5058), .B(n5057), .Z(n5062) );
  NAND U6490 ( .A(n5060), .B(n5059), .Z(n5061) );
  AND U6491 ( .A(n5062), .B(n5061), .Z(n5619) );
  XNOR U6492 ( .A(n5620), .B(n5619), .Z(n5587) );
  XOR U6493 ( .A(n5590), .B(n5589), .Z(n5528) );
  XOR U6494 ( .A(n5529), .B(n5528), .Z(n5531) );
  XOR U6495 ( .A(n5530), .B(n5531), .Z(n5410) );
  XOR U6496 ( .A(n5411), .B(n5410), .Z(n5722) );
  XOR U6497 ( .A(n5723), .B(n5722), .Z(n5725) );
  XOR U6498 ( .A(n5724), .B(n5725), .Z(n5719) );
  NAND U6499 ( .A(n5064), .B(n5063), .Z(n5068) );
  NAND U6500 ( .A(n5066), .B(n5065), .Z(n5067) );
  NAND U6501 ( .A(n5068), .B(n5067), .Z(n5459) );
  NAND U6502 ( .A(n5070), .B(n5069), .Z(n5074) );
  NAND U6503 ( .A(n5072), .B(n5071), .Z(n5073) );
  NAND U6504 ( .A(n5074), .B(n5073), .Z(n5457) );
  NAND U6505 ( .A(n5076), .B(n5075), .Z(n5080) );
  NAND U6506 ( .A(n5078), .B(n5077), .Z(n5079) );
  NAND U6507 ( .A(n5080), .B(n5079), .Z(n5456) );
  NAND U6508 ( .A(n5082), .B(n5081), .Z(n5086) );
  NAND U6509 ( .A(n5084), .B(n5083), .Z(n5085) );
  NAND U6510 ( .A(n5086), .B(n5085), .Z(n5544) );
  NAND U6511 ( .A(n5088), .B(n5087), .Z(n5092) );
  NANDN U6512 ( .A(n5090), .B(n5089), .Z(n5091) );
  AND U6513 ( .A(n5092), .B(n5091), .Z(n5650) );
  NAND U6514 ( .A(n5094), .B(n5093), .Z(n5098) );
  NAND U6515 ( .A(n5096), .B(n5095), .Z(n5097) );
  AND U6516 ( .A(n5098), .B(n5097), .Z(n5647) );
  NAND U6517 ( .A(n5100), .B(n5099), .Z(n5104) );
  NANDN U6518 ( .A(n5102), .B(n5101), .Z(n5103) );
  AND U6519 ( .A(n5104), .B(n5103), .Z(n5648) );
  XNOR U6520 ( .A(n5650), .B(n5649), .Z(n5545) );
  XNOR U6521 ( .A(n5544), .B(n5545), .Z(n5105) );
  XNOR U6522 ( .A(n5546), .B(n5105), .Z(n5519) );
  NAND U6523 ( .A(n5107), .B(n5106), .Z(n5111) );
  NAND U6524 ( .A(n5109), .B(n5108), .Z(n5110) );
  NAND U6525 ( .A(n5111), .B(n5110), .Z(n5517) );
  NAND U6526 ( .A(n5113), .B(n5112), .Z(n5117) );
  NAND U6527 ( .A(n5115), .B(n5114), .Z(n5116) );
  NAND U6528 ( .A(n5117), .B(n5116), .Z(n5516) );
  XOR U6529 ( .A(n5517), .B(n5516), .Z(n5518) );
  IV U6530 ( .A(n5689), .Z(n5687) );
  NANDN U6531 ( .A(n5119), .B(n5118), .Z(n5123) );
  NAND U6532 ( .A(n5121), .B(n5120), .Z(n5122) );
  NAND U6533 ( .A(n5123), .B(n5122), .Z(n5691) );
  NAND U6534 ( .A(n5125), .B(n5124), .Z(n5129) );
  NANDN U6535 ( .A(n5127), .B(n5126), .Z(n5128) );
  AND U6536 ( .A(n5129), .B(n5128), .Z(n5483) );
  NAND U6537 ( .A(n5131), .B(n5130), .Z(n5135) );
  NAND U6538 ( .A(n5133), .B(n5132), .Z(n5134) );
  NAND U6539 ( .A(n5135), .B(n5134), .Z(n5481) );
  NAND U6540 ( .A(n5137), .B(n5136), .Z(n5141) );
  NAND U6541 ( .A(n5139), .B(n5138), .Z(n5140) );
  NAND U6542 ( .A(n5141), .B(n5140), .Z(n5480) );
  XOR U6543 ( .A(n5483), .B(n5482), .Z(n5697) );
  NAND U6544 ( .A(n5143), .B(n5142), .Z(n5147) );
  NAND U6545 ( .A(n5145), .B(n5144), .Z(n5146) );
  NAND U6546 ( .A(n5147), .B(n5146), .Z(n5695) );
  NAND U6547 ( .A(n5149), .B(n5148), .Z(n5153) );
  NAND U6548 ( .A(n5151), .B(n5150), .Z(n5152) );
  NAND U6549 ( .A(n5153), .B(n5152), .Z(n5696) );
  XNOR U6550 ( .A(n5695), .B(n5696), .Z(n5154) );
  XNOR U6551 ( .A(n5697), .B(n5154), .Z(n5688) );
  IV U6552 ( .A(n5688), .Z(n5690) );
  XNOR U6553 ( .A(n5691), .B(n5690), .Z(n5155) );
  XOR U6554 ( .A(n5687), .B(n5155), .Z(n5489) );
  NAND U6555 ( .A(n5157), .B(n5156), .Z(n5161) );
  NAND U6556 ( .A(n5159), .B(n5158), .Z(n5160) );
  AND U6557 ( .A(n5161), .B(n5160), .Z(n5661) );
  NAND U6558 ( .A(n5163), .B(n5162), .Z(n5167) );
  NAND U6559 ( .A(n5165), .B(n5164), .Z(n5166) );
  AND U6560 ( .A(n5167), .B(n5166), .Z(n5660) );
  OR U6561 ( .A(n5169), .B(n5168), .Z(n5173) );
  NANDN U6562 ( .A(n5171), .B(n5170), .Z(n5172) );
  AND U6563 ( .A(n5173), .B(n5172), .Z(n5659) );
  NAND U6564 ( .A(n5175), .B(n5174), .Z(n5179) );
  NAND U6565 ( .A(n5177), .B(n5176), .Z(n5178) );
  AND U6566 ( .A(n5179), .B(n5178), .Z(n5554) );
  XOR U6567 ( .A(n5553), .B(n5554), .Z(n5555) );
  NAND U6568 ( .A(n5181), .B(n5180), .Z(n5185) );
  NAND U6569 ( .A(n5183), .B(n5182), .Z(n5184) );
  AND U6570 ( .A(n5185), .B(n5184), .Z(n5556) );
  NAND U6571 ( .A(n5187), .B(n5186), .Z(n5191) );
  NAND U6572 ( .A(n5189), .B(n5188), .Z(n5190) );
  AND U6573 ( .A(n5191), .B(n5190), .Z(n5492) );
  NAND U6574 ( .A(n5193), .B(n5192), .Z(n5197) );
  NAND U6575 ( .A(n5195), .B(n5194), .Z(n5196) );
  NAND U6576 ( .A(n5197), .B(n5196), .Z(n5494) );
  XNOR U6577 ( .A(n5495), .B(n5494), .Z(n5525) );
  NAND U6578 ( .A(n5199), .B(n5198), .Z(n5203) );
  NAND U6579 ( .A(n5201), .B(n5200), .Z(n5202) );
  NAND U6580 ( .A(n5203), .B(n5202), .Z(n5498) );
  NAND U6581 ( .A(n5205), .B(n5204), .Z(n5209) );
  NAND U6582 ( .A(n5207), .B(n5206), .Z(n5208) );
  AND U6583 ( .A(n5209), .B(n5208), .Z(n5499) );
  XOR U6584 ( .A(n5498), .B(n5499), .Z(n5501) );
  NAND U6585 ( .A(n5211), .B(n5210), .Z(n5215) );
  NAND U6586 ( .A(n5213), .B(n5212), .Z(n5214) );
  NAND U6587 ( .A(n5215), .B(n5214), .Z(n5500) );
  XNOR U6588 ( .A(n5501), .B(n5500), .Z(n5523) );
  NAND U6589 ( .A(n5217), .B(n5216), .Z(n5221) );
  NAND U6590 ( .A(n5219), .B(n5218), .Z(n5220) );
  AND U6591 ( .A(n5221), .B(n5220), .Z(n5716) );
  NAND U6592 ( .A(n5223), .B(n5222), .Z(n5227) );
  NAND U6593 ( .A(n5225), .B(n5224), .Z(n5226) );
  NAND U6594 ( .A(n5227), .B(n5226), .Z(n5714) );
  NAND U6595 ( .A(n5229), .B(n5228), .Z(n5233) );
  NAND U6596 ( .A(n5231), .B(n5230), .Z(n5232) );
  NAND U6597 ( .A(n5233), .B(n5232), .Z(n5713) );
  XOR U6598 ( .A(n5716), .B(n5715), .Z(n5522) );
  NAND U6599 ( .A(n5235), .B(n5234), .Z(n5239) );
  NAND U6600 ( .A(n5237), .B(n5236), .Z(n5238) );
  NAND U6601 ( .A(n5239), .B(n5238), .Z(n5440) );
  NAND U6602 ( .A(n5241), .B(n5240), .Z(n5245) );
  NANDN U6603 ( .A(n5243), .B(n5242), .Z(n5244) );
  NAND U6604 ( .A(n5245), .B(n5244), .Z(n5438) );
  NAND U6605 ( .A(n5247), .B(n5246), .Z(n5251) );
  NANDN U6606 ( .A(n5249), .B(n5248), .Z(n5250) );
  AND U6607 ( .A(n5251), .B(n5250), .Z(n5638) );
  NAND U6608 ( .A(n5253), .B(n5252), .Z(n5257) );
  NAND U6609 ( .A(n5255), .B(n5254), .Z(n5256) );
  AND U6610 ( .A(n5257), .B(n5256), .Z(n5635) );
  NAND U6611 ( .A(n5259), .B(n5258), .Z(n5263) );
  NANDN U6612 ( .A(n5261), .B(n5260), .Z(n5262) );
  AND U6613 ( .A(n5263), .B(n5262), .Z(n5636) );
  XNOR U6614 ( .A(n5638), .B(n5637), .Z(n5539) );
  NAND U6615 ( .A(n5265), .B(n5264), .Z(n5269) );
  NAND U6616 ( .A(n5267), .B(n5266), .Z(n5268) );
  AND U6617 ( .A(n5269), .B(n5268), .Z(n5538) );
  NAND U6618 ( .A(n5271), .B(n5270), .Z(n5275) );
  NAND U6619 ( .A(n5273), .B(n5272), .Z(n5274) );
  AND U6620 ( .A(n5275), .B(n5274), .Z(n5577) );
  XNOR U6621 ( .A(n5577), .B(oglobal[3]), .Z(n5614) );
  NANDN U6622 ( .A(n5277), .B(n5276), .Z(n5281) );
  NAND U6623 ( .A(n5279), .B(n5278), .Z(n5280) );
  NAND U6624 ( .A(n5281), .B(n5280), .Z(n5612) );
  NAND U6625 ( .A(n5283), .B(n5282), .Z(n5287) );
  NAND U6626 ( .A(n5285), .B(n5284), .Z(n5286) );
  AND U6627 ( .A(n5287), .B(n5286), .Z(n5611) );
  XOR U6628 ( .A(n5541), .B(n5540), .Z(n5586) );
  NAND U6629 ( .A(n5289), .B(n5288), .Z(n5293) );
  NAND U6630 ( .A(n5291), .B(n5290), .Z(n5292) );
  AND U6631 ( .A(n5293), .B(n5292), .Z(n5471) );
  NAND U6632 ( .A(n5295), .B(n5294), .Z(n5299) );
  NANDN U6633 ( .A(n5297), .B(n5296), .Z(n5298) );
  AND U6634 ( .A(n5299), .B(n5298), .Z(n5468) );
  OR U6635 ( .A(n5301), .B(n5300), .Z(n5305) );
  NANDN U6636 ( .A(n5303), .B(n5302), .Z(n5304) );
  AND U6637 ( .A(n5305), .B(n5304), .Z(n5469) );
  XNOR U6638 ( .A(n5471), .B(n5470), .Z(n5712) );
  NAND U6639 ( .A(n5307), .B(n5306), .Z(n5311) );
  NAND U6640 ( .A(n5309), .B(n5308), .Z(n5310) );
  AND U6641 ( .A(n5311), .B(n5310), .Z(n5711) );
  NAND U6642 ( .A(n5313), .B(n5312), .Z(n5317) );
  NAND U6643 ( .A(n5315), .B(n5314), .Z(n5316) );
  AND U6644 ( .A(n5317), .B(n5316), .Z(n5710) );
  XNOR U6645 ( .A(n5711), .B(n5710), .Z(n5318) );
  XNOR U6646 ( .A(n5712), .B(n5318), .Z(n5585) );
  NAND U6647 ( .A(n5320), .B(n5319), .Z(n5324) );
  NAND U6648 ( .A(n5322), .B(n5321), .Z(n5323) );
  AND U6649 ( .A(n5324), .B(n5323), .Z(n5584) );
  XOR U6650 ( .A(n5438), .B(n5439), .Z(n5441) );
  XNOR U6651 ( .A(n5486), .B(n5487), .Z(n5488) );
  NANDN U6652 ( .A(n5326), .B(n5325), .Z(n5330) );
  NANDN U6653 ( .A(n5328), .B(n5327), .Z(n5329) );
  NAND U6654 ( .A(n5330), .B(n5329), .Z(n5383) );
  NANDN U6655 ( .A(n5332), .B(n5331), .Z(n5336) );
  NAND U6656 ( .A(n5334), .B(n5333), .Z(n5335) );
  NAND U6657 ( .A(n5336), .B(n5335), .Z(n5382) );
  NANDN U6658 ( .A(n5338), .B(n5337), .Z(n5342) );
  NAND U6659 ( .A(n5340), .B(n5339), .Z(n5341) );
  NAND U6660 ( .A(n5342), .B(n5341), .Z(n5381) );
  XOR U6661 ( .A(n5382), .B(n5381), .Z(n5384) );
  XNOR U6662 ( .A(n5383), .B(n5384), .Z(n5400) );
  NAND U6663 ( .A(n5344), .B(n5343), .Z(n5348) );
  NAND U6664 ( .A(n5346), .B(n5345), .Z(n5347) );
  NAND U6665 ( .A(n5348), .B(n5347), .Z(n5399) );
  XNOR U6666 ( .A(n5721), .B(n5720), .Z(n5352) );
  XOR U6667 ( .A(n5719), .B(n5352), .Z(n5407) );
  NANDN U6668 ( .A(n5357), .B(n5356), .Z(n5361) );
  NANDN U6669 ( .A(n5359), .B(n5358), .Z(n5360) );
  AND U6670 ( .A(n5361), .B(n5360), .Z(n5376) );
  NAND U6671 ( .A(n5363), .B(n5362), .Z(n5367) );
  NANDN U6672 ( .A(n5365), .B(n5364), .Z(n5366) );
  NAND U6673 ( .A(n5367), .B(n5366), .Z(n5375) );
  XOR U6674 ( .A(n5376), .B(n5375), .Z(n5378) );
  NAND U6675 ( .A(n5369), .B(n5368), .Z(n5373) );
  NAND U6676 ( .A(n5371), .B(n5370), .Z(n5372) );
  NAND U6677 ( .A(n5373), .B(n5372), .Z(n5377) );
  XNOR U6678 ( .A(n5378), .B(n5377), .Z(n5406) );
  XNOR U6679 ( .A(n5405), .B(n5406), .Z(n5374) );
  XNOR U6680 ( .A(n5407), .B(n5374), .Z(o[3]) );
  NAND U6681 ( .A(n5376), .B(n5375), .Z(n5380) );
  NAND U6682 ( .A(n5378), .B(n5377), .Z(n5379) );
  NAND U6683 ( .A(n5380), .B(n5379), .Z(n5882) );
  NAND U6684 ( .A(n5382), .B(n5381), .Z(n5386) );
  NAND U6685 ( .A(n5384), .B(n5383), .Z(n5385) );
  NAND U6686 ( .A(n5386), .B(n5385), .Z(n5894) );
  NAND U6687 ( .A(n5388), .B(n5387), .Z(n5392) );
  NAND U6688 ( .A(n5390), .B(n5389), .Z(n5391) );
  AND U6689 ( .A(n5392), .B(n5391), .Z(n5893) );
  NAND U6690 ( .A(n5394), .B(n5393), .Z(n5398) );
  NAND U6691 ( .A(n5396), .B(n5395), .Z(n5397) );
  AND U6692 ( .A(n5398), .B(n5397), .Z(n5892) );
  XOR U6693 ( .A(n5893), .B(n5892), .Z(n5895) );
  XNOR U6694 ( .A(n5894), .B(n5895), .Z(n5881) );
  NAND U6695 ( .A(n5400), .B(n5399), .Z(n5404) );
  NAND U6696 ( .A(n5402), .B(n5401), .Z(n5403) );
  NAND U6697 ( .A(n5404), .B(n5403), .Z(n5880) );
  XOR U6698 ( .A(n5882), .B(n5883), .Z(n5907) );
  NAND U6699 ( .A(n5409), .B(n5408), .Z(n5413) );
  NAND U6700 ( .A(n5411), .B(n5410), .Z(n5412) );
  NAND U6701 ( .A(n5413), .B(n5412), .Z(n5731) );
  NANDN U6702 ( .A(n5415), .B(n5414), .Z(n5419) );
  NAND U6703 ( .A(n5417), .B(n5416), .Z(n5418) );
  NAND U6704 ( .A(n5419), .B(n5418), .Z(n5735) );
  NANDN U6705 ( .A(n5421), .B(n5420), .Z(n5425) );
  NAND U6706 ( .A(n5423), .B(n5422), .Z(n5424) );
  AND U6707 ( .A(n5425), .B(n5424), .Z(n5736) );
  XOR U6708 ( .A(n5735), .B(n5736), .Z(n5738) );
  NAND U6709 ( .A(n5427), .B(n5426), .Z(n5431) );
  NAND U6710 ( .A(n5429), .B(n5428), .Z(n5430) );
  AND U6711 ( .A(n5431), .B(n5430), .Z(n5737) );
  XNOR U6712 ( .A(n5738), .B(n5737), .Z(n5730) );
  OR U6713 ( .A(n5433), .B(n5432), .Z(n5437) );
  NAND U6714 ( .A(n5435), .B(n5434), .Z(n5436) );
  NAND U6715 ( .A(n5437), .B(n5436), .Z(n5870) );
  NAND U6716 ( .A(n5439), .B(n5438), .Z(n5443) );
  NAND U6717 ( .A(n5441), .B(n5440), .Z(n5442) );
  NAND U6718 ( .A(n5443), .B(n5442), .Z(n5868) );
  NAND U6719 ( .A(n5445), .B(n5444), .Z(n5449) );
  NAND U6720 ( .A(n5447), .B(n5446), .Z(n5448) );
  AND U6721 ( .A(n5449), .B(n5448), .Z(n5786) );
  NAND U6722 ( .A(n5451), .B(n5450), .Z(n5455) );
  NAND U6723 ( .A(n5453), .B(n5452), .Z(n5454) );
  NAND U6724 ( .A(n5455), .B(n5454), .Z(n5784) );
  NAND U6725 ( .A(n5457), .B(n5456), .Z(n5461) );
  NAND U6726 ( .A(n5459), .B(n5458), .Z(n5460) );
  AND U6727 ( .A(n5461), .B(n5460), .Z(n5847) );
  NAND U6728 ( .A(n5463), .B(n5462), .Z(n5467) );
  NAND U6729 ( .A(n5465), .B(n5464), .Z(n5466) );
  NAND U6730 ( .A(n5467), .B(n5466), .Z(n5845) );
  NAND U6731 ( .A(n5469), .B(n5468), .Z(n5473) );
  NAND U6732 ( .A(n5471), .B(n5470), .Z(n5472) );
  NAND U6733 ( .A(n5473), .B(n5472), .Z(n5844) );
  XNOR U6734 ( .A(n5847), .B(n5846), .Z(n5857) );
  NAND U6735 ( .A(n5475), .B(n5474), .Z(n5479) );
  NAND U6736 ( .A(n5477), .B(n5476), .Z(n5478) );
  AND U6737 ( .A(n5479), .B(n5478), .Z(n5856) );
  NAND U6738 ( .A(n5481), .B(n5480), .Z(n5485) );
  NANDN U6739 ( .A(n5483), .B(n5482), .Z(n5484) );
  AND U6740 ( .A(n5485), .B(n5484), .Z(n5859) );
  XOR U6741 ( .A(n5786), .B(n5785), .Z(n5869) );
  XOR U6742 ( .A(n5868), .B(n5869), .Z(n5871) );
  XOR U6743 ( .A(n5870), .B(n5871), .Z(n5729) );
  XOR U6744 ( .A(n5731), .B(n5732), .Z(n5889) );
  NANDN U6745 ( .A(n5487), .B(n5486), .Z(n5491) );
  NAND U6746 ( .A(n5489), .B(n5488), .Z(n5490) );
  NAND U6747 ( .A(n5491), .B(n5490), .Z(n5886) );
  NAND U6748 ( .A(n5493), .B(n5492), .Z(n5497) );
  NAND U6749 ( .A(n5495), .B(n5494), .Z(n5496) );
  AND U6750 ( .A(n5497), .B(n5496), .Z(n5772) );
  NAND U6751 ( .A(n5499), .B(n5498), .Z(n5503) );
  NAND U6752 ( .A(n5501), .B(n5500), .Z(n5502) );
  AND U6753 ( .A(n5503), .B(n5502), .Z(n5771) );
  XOR U6754 ( .A(n5772), .B(n5771), .Z(n5774) );
  NAND U6755 ( .A(n5505), .B(n5504), .Z(n5509) );
  NAND U6756 ( .A(n5507), .B(n5506), .Z(n5508) );
  AND U6757 ( .A(n5509), .B(n5508), .Z(n5773) );
  XOR U6758 ( .A(n5774), .B(n5773), .Z(n5749) );
  NAND U6759 ( .A(n5511), .B(n5510), .Z(n5515) );
  NANDN U6760 ( .A(n5513), .B(n5512), .Z(n5514) );
  NAND U6761 ( .A(n5515), .B(n5514), .Z(n5747) );
  NAND U6762 ( .A(n5517), .B(n5516), .Z(n5521) );
  NAND U6763 ( .A(n5519), .B(n5518), .Z(n5520) );
  AND U6764 ( .A(n5521), .B(n5520), .Z(n5748) );
  XOR U6765 ( .A(n5747), .B(n5748), .Z(n5750) );
  NAND U6766 ( .A(n5523), .B(n5522), .Z(n5527) );
  NAND U6767 ( .A(n5525), .B(n5524), .Z(n5526) );
  AND U6768 ( .A(n5527), .B(n5526), .Z(n5863) );
  NAND U6769 ( .A(n5529), .B(n5528), .Z(n5533) );
  NAND U6770 ( .A(n5531), .B(n5530), .Z(n5532) );
  AND U6771 ( .A(n5533), .B(n5532), .Z(n5862) );
  XOR U6772 ( .A(n5863), .B(n5862), .Z(n5864) );
  NAND U6773 ( .A(n5539), .B(n5538), .Z(n5543) );
  NAND U6774 ( .A(n5541), .B(n5540), .Z(n5542) );
  AND U6775 ( .A(n5543), .B(n5542), .Z(n5852) );
  OR U6776 ( .A(n5548), .B(n5547), .Z(n5552) );
  NAND U6777 ( .A(n5550), .B(n5549), .Z(n5551) );
  NAND U6778 ( .A(n5552), .B(n5551), .Z(n5850) );
  XNOR U6779 ( .A(n5851), .B(n5850), .Z(n5853) );
  XNOR U6780 ( .A(n5778), .B(n5777), .Z(n5780) );
  NAND U6781 ( .A(n5554), .B(n5553), .Z(n5558) );
  NAND U6782 ( .A(n5556), .B(n5555), .Z(n5557) );
  AND U6783 ( .A(n5558), .B(n5557), .Z(n5768) );
  NAND U6784 ( .A(n5560), .B(n5559), .Z(n5564) );
  NAND U6785 ( .A(n5562), .B(n5561), .Z(n5563) );
  AND U6786 ( .A(n5564), .B(n5563), .Z(n5766) );
  NAND U6787 ( .A(n5566), .B(n5565), .Z(n5570) );
  NAND U6788 ( .A(n5568), .B(n5567), .Z(n5569) );
  NAND U6789 ( .A(n5570), .B(n5569), .Z(n5834) );
  NAND U6790 ( .A(n5572), .B(n5571), .Z(n5576) );
  NAND U6791 ( .A(n5574), .B(n5573), .Z(n5575) );
  NAND U6792 ( .A(n5576), .B(n5575), .Z(n5832) );
  AND U6793 ( .A(n5577), .B(oglobal[3]), .Z(n5837) );
  XOR U6794 ( .A(n5766), .B(n5765), .Z(n5767) );
  XOR U6795 ( .A(n5768), .B(n5767), .Z(n5779) );
  XNOR U6796 ( .A(n5780), .B(n5779), .Z(n5875) );
  NAND U6797 ( .A(n5579), .B(n5578), .Z(n5583) );
  NAND U6798 ( .A(n5581), .B(n5580), .Z(n5582) );
  NAND U6799 ( .A(n5583), .B(n5582), .Z(n5796) );
  NAND U6800 ( .A(n5588), .B(n5587), .Z(n5592) );
  NANDN U6801 ( .A(n5590), .B(n5589), .Z(n5591) );
  AND U6802 ( .A(n5592), .B(n5591), .Z(n5798) );
  NANDN U6803 ( .A(n5594), .B(n5593), .Z(n5598) );
  NAND U6804 ( .A(n5596), .B(n5595), .Z(n5597) );
  NAND U6805 ( .A(n5598), .B(n5597), .Z(n5814) );
  NAND U6806 ( .A(n5600), .B(n5599), .Z(n5604) );
  NAND U6807 ( .A(n5602), .B(n5601), .Z(n5603) );
  AND U6808 ( .A(n5604), .B(n5603), .Z(n5822) );
  NAND U6809 ( .A(n5606), .B(n5605), .Z(n5610) );
  NAND U6810 ( .A(n5608), .B(n5607), .Z(n5609) );
  NAND U6811 ( .A(n5610), .B(n5609), .Z(n5820) );
  NAND U6812 ( .A(n5612), .B(n5611), .Z(n5616) );
  NAND U6813 ( .A(n5614), .B(n5613), .Z(n5615) );
  AND U6814 ( .A(n5616), .B(n5615), .Z(n5819) );
  XNOR U6815 ( .A(n5822), .B(n5821), .Z(n5813) );
  XOR U6816 ( .A(n5814), .B(n5813), .Z(n5816) );
  NAND U6817 ( .A(n5618), .B(n5617), .Z(n5622) );
  NAND U6818 ( .A(n5620), .B(n5619), .Z(n5621) );
  NAND U6819 ( .A(n5622), .B(n5621), .Z(n5815) );
  XNOR U6820 ( .A(n5816), .B(n5815), .Z(n5756) );
  NANDN U6821 ( .A(n5624), .B(n5623), .Z(n5628) );
  NAND U6822 ( .A(n5626), .B(n5625), .Z(n5627) );
  AND U6823 ( .A(n5628), .B(n5627), .Z(n5753) );
  NAND U6824 ( .A(n5630), .B(n5629), .Z(n5634) );
  NAND U6825 ( .A(n5632), .B(n5631), .Z(n5633) );
  AND U6826 ( .A(n5634), .B(n5633), .Z(n5754) );
  NAND U6827 ( .A(n5636), .B(n5635), .Z(n5640) );
  NAND U6828 ( .A(n5638), .B(n5637), .Z(n5639) );
  NAND U6829 ( .A(n5640), .B(n5639), .Z(n5841) );
  NAND U6830 ( .A(n5642), .B(n5641), .Z(n5646) );
  NAND U6831 ( .A(n5644), .B(n5643), .Z(n5645) );
  NAND U6832 ( .A(n5646), .B(n5645), .Z(n5839) );
  NAND U6833 ( .A(n5648), .B(n5647), .Z(n5652) );
  NAND U6834 ( .A(n5650), .B(n5649), .Z(n5651) );
  NAND U6835 ( .A(n5652), .B(n5651), .Z(n5828) );
  IV U6836 ( .A(n5828), .Z(n5662) );
  OR U6837 ( .A(n5654), .B(n5653), .Z(n5658) );
  NAND U6838 ( .A(n5656), .B(n5655), .Z(n5657) );
  NAND U6839 ( .A(n5658), .B(n5657), .Z(n5826) );
  XNOR U6840 ( .A(n5662), .B(n5827), .Z(n5838) );
  NAND U6841 ( .A(n5664), .B(n5663), .Z(n5668) );
  NAND U6842 ( .A(n5666), .B(n5665), .Z(n5667) );
  AND U6843 ( .A(n5668), .B(n5667), .Z(n5759) );
  NAND U6844 ( .A(n5670), .B(n5669), .Z(n5674) );
  NAND U6845 ( .A(n5672), .B(n5671), .Z(n5673) );
  AND U6846 ( .A(n5674), .B(n5673), .Z(n5760) );
  XNOR U6847 ( .A(n5762), .B(n5761), .Z(n5790) );
  NAND U6848 ( .A(n5676), .B(n5675), .Z(n5680) );
  NAND U6849 ( .A(n5678), .B(n5677), .Z(n5679) );
  AND U6850 ( .A(n5680), .B(n5679), .Z(n5789) );
  XOR U6851 ( .A(n5791), .B(n5792), .Z(n5877) );
  NAND U6852 ( .A(n5682), .B(n5681), .Z(n5686) );
  NANDN U6853 ( .A(n5684), .B(n5683), .Z(n5685) );
  AND U6854 ( .A(n5686), .B(n5685), .Z(n5744) );
  NAND U6855 ( .A(n5688), .B(n5687), .Z(n5694) );
  AND U6856 ( .A(n5690), .B(n5689), .Z(n5692) );
  OR U6857 ( .A(n5692), .B(n5691), .Z(n5693) );
  AND U6858 ( .A(n5694), .B(n5693), .Z(n5742) );
  NAND U6859 ( .A(n5699), .B(n5698), .Z(n5703) );
  NAND U6860 ( .A(n5701), .B(n5700), .Z(n5702) );
  NAND U6861 ( .A(n5703), .B(n5702), .Z(n5810) );
  NAND U6862 ( .A(n5705), .B(n5704), .Z(n5709) );
  NAND U6863 ( .A(n5707), .B(n5706), .Z(n5708) );
  NAND U6864 ( .A(n5709), .B(n5708), .Z(n5808) );
  XOR U6865 ( .A(n5802), .B(n5801), .Z(n5804) );
  NAND U6866 ( .A(n5714), .B(n5713), .Z(n5718) );
  NANDN U6867 ( .A(n5716), .B(n5715), .Z(n5717) );
  AND U6868 ( .A(n5718), .B(n5717), .Z(n5803) );
  XOR U6869 ( .A(n5804), .B(n5803), .Z(n5741) );
  XOR U6870 ( .A(n5742), .B(n5741), .Z(n5743) );
  XOR U6871 ( .A(n5744), .B(n5743), .Z(n5898) );
  XOR U6872 ( .A(n5899), .B(n5898), .Z(n5900) );
  XOR U6873 ( .A(n5886), .B(n5887), .Z(n5888) );
  XOR U6874 ( .A(n5889), .B(n5888), .Z(n5914) );
  NANDN U6875 ( .A(n5723), .B(n5722), .Z(n5727) );
  NANDN U6876 ( .A(n5725), .B(n5724), .Z(n5726) );
  NAND U6877 ( .A(n5727), .B(n5726), .Z(n5912) );
  XNOR U6878 ( .A(n5911), .B(n5912), .Z(n5913) );
  XOR U6879 ( .A(n5914), .B(n5913), .Z(n5905) );
  IV U6880 ( .A(n5905), .Z(n5904) );
  XNOR U6881 ( .A(n5906), .B(n5904), .Z(n5728) );
  XNOR U6882 ( .A(n5907), .B(n5728), .Z(o[4]) );
  NAND U6883 ( .A(n5730), .B(n5729), .Z(n5734) );
  NAND U6884 ( .A(n5732), .B(n5731), .Z(n5733) );
  NAND U6885 ( .A(n5734), .B(n5733), .Z(n5942) );
  NAND U6886 ( .A(n5736), .B(n5735), .Z(n5740) );
  NAND U6887 ( .A(n5738), .B(n5737), .Z(n5739) );
  AND U6888 ( .A(n5740), .B(n5739), .Z(n5926) );
  NAND U6889 ( .A(n5742), .B(n5741), .Z(n5746) );
  NAND U6890 ( .A(n5744), .B(n5743), .Z(n5745) );
  NAND U6891 ( .A(n5746), .B(n5745), .Z(n5924) );
  NAND U6892 ( .A(n5748), .B(n5747), .Z(n5752) );
  NAND U6893 ( .A(n5750), .B(n5749), .Z(n5751) );
  AND U6894 ( .A(n5752), .B(n5751), .Z(n5933) );
  NAND U6895 ( .A(n5754), .B(n5753), .Z(n5758) );
  NAND U6896 ( .A(n5756), .B(n5755), .Z(n5757) );
  NAND U6897 ( .A(n5758), .B(n5757), .Z(n5986) );
  NAND U6898 ( .A(n5760), .B(n5759), .Z(n5764) );
  NAND U6899 ( .A(n5762), .B(n5761), .Z(n5763) );
  NAND U6900 ( .A(n5764), .B(n5763), .Z(n5984) );
  NAND U6901 ( .A(n5766), .B(n5765), .Z(n5770) );
  NAND U6902 ( .A(n5768), .B(n5767), .Z(n5769) );
  NAND U6903 ( .A(n5770), .B(n5769), .Z(n5983) );
  NAND U6904 ( .A(n5772), .B(n5771), .Z(n5776) );
  NAND U6905 ( .A(n5774), .B(n5773), .Z(n5775) );
  AND U6906 ( .A(n5776), .B(n5775), .Z(n5930) );
  XOR U6907 ( .A(n5931), .B(n5930), .Z(n5932) );
  XNOR U6908 ( .A(n5933), .B(n5932), .Z(n5925) );
  XNOR U6909 ( .A(n5926), .B(n5927), .Z(n5943) );
  XOR U6910 ( .A(n5942), .B(n5943), .Z(n5944) );
  NANDN U6911 ( .A(n5778), .B(n5777), .Z(n5782) );
  NAND U6912 ( .A(n5780), .B(n5779), .Z(n5781) );
  NAND U6913 ( .A(n5782), .B(n5781), .Z(n5990) );
  NAND U6914 ( .A(n5784), .B(n5783), .Z(n5788) );
  NAND U6915 ( .A(n5786), .B(n5785), .Z(n5787) );
  AND U6916 ( .A(n5788), .B(n5787), .Z(n5989) );
  NAND U6917 ( .A(n5790), .B(n5789), .Z(n5794) );
  NAND U6918 ( .A(n5792), .B(n5791), .Z(n5793) );
  AND U6919 ( .A(n5794), .B(n5793), .Z(n5992) );
  NAND U6920 ( .A(n5796), .B(n5795), .Z(n5800) );
  NAND U6921 ( .A(n5798), .B(n5797), .Z(n5799) );
  AND U6922 ( .A(n5800), .B(n5799), .Z(n5995) );
  NAND U6923 ( .A(n5802), .B(n5801), .Z(n5806) );
  NAND U6924 ( .A(n5804), .B(n5803), .Z(n5805) );
  AND U6925 ( .A(n5806), .B(n5805), .Z(n5996) );
  NAND U6926 ( .A(n5808), .B(n5807), .Z(n5812) );
  NAND U6927 ( .A(n5810), .B(n5809), .Z(n5811) );
  AND U6928 ( .A(n5812), .B(n5811), .Z(n5954) );
  NAND U6929 ( .A(n5814), .B(n5813), .Z(n5818) );
  NAND U6930 ( .A(n5816), .B(n5815), .Z(n5817) );
  AND U6931 ( .A(n5818), .B(n5817), .Z(n5955) );
  NAND U6932 ( .A(n5820), .B(n5819), .Z(n5824) );
  NAND U6933 ( .A(n5822), .B(n5821), .Z(n5823) );
  NAND U6934 ( .A(n5824), .B(n5823), .Z(n5966) );
  NAND U6935 ( .A(n5826), .B(n5825), .Z(n5830) );
  NAND U6936 ( .A(n5828), .B(n5827), .Z(n5829) );
  NAND U6937 ( .A(n5830), .B(n5829), .Z(n5965) );
  NAND U6938 ( .A(n5832), .B(n5831), .Z(n5836) );
  NAND U6939 ( .A(n5834), .B(n5833), .Z(n5835) );
  NAND U6940 ( .A(n5836), .B(n5835), .Z(n5962) );
  AND U6941 ( .A(oglobal[4]), .B(n5837), .Z(n5960) );
  XOR U6942 ( .A(oglobal[5]), .B(n5960), .Z(n5961) );
  XNOR U6943 ( .A(n5968), .B(n5967), .Z(n5974) );
  NAND U6944 ( .A(n5839), .B(n5838), .Z(n5843) );
  NAND U6945 ( .A(n5841), .B(n5840), .Z(n5842) );
  AND U6946 ( .A(n5843), .B(n5842), .Z(n5971) );
  NAND U6947 ( .A(n5845), .B(n5844), .Z(n5849) );
  NAND U6948 ( .A(n5847), .B(n5846), .Z(n5848) );
  AND U6949 ( .A(n5849), .B(n5848), .Z(n5972) );
  NANDN U6950 ( .A(n5851), .B(n5850), .Z(n5855) );
  NAND U6951 ( .A(n5853), .B(n5852), .Z(n5854) );
  NAND U6952 ( .A(n5855), .B(n5854), .Z(n5978) );
  NAND U6953 ( .A(n5857), .B(n5856), .Z(n5861) );
  NAND U6954 ( .A(n5859), .B(n5858), .Z(n5860) );
  AND U6955 ( .A(n5861), .B(n5860), .Z(n5977) );
  XOR U6956 ( .A(n5979), .B(n5980), .Z(n5956) );
  XOR U6957 ( .A(n5957), .B(n5956), .Z(n5997) );
  XOR U6958 ( .A(n5998), .B(n5997), .Z(n5936) );
  XOR U6959 ( .A(n5937), .B(n5936), .Z(n5939) );
  NAND U6960 ( .A(n5863), .B(n5862), .Z(n5867) );
  NAND U6961 ( .A(n5865), .B(n5864), .Z(n5866) );
  NAND U6962 ( .A(n5867), .B(n5866), .Z(n5938) );
  XNOR U6963 ( .A(n5939), .B(n5938), .Z(n5950) );
  NAND U6964 ( .A(n5869), .B(n5868), .Z(n5873) );
  NAND U6965 ( .A(n5871), .B(n5870), .Z(n5872) );
  NAND U6966 ( .A(n5873), .B(n5872), .Z(n5949) );
  NAND U6967 ( .A(n5875), .B(n5874), .Z(n5879) );
  NAND U6968 ( .A(n5877), .B(n5876), .Z(n5878) );
  NAND U6969 ( .A(n5879), .B(n5878), .Z(n5948) );
  XOR U6970 ( .A(n5949), .B(n5948), .Z(n5951) );
  XNOR U6971 ( .A(n5944), .B(n5945), .Z(n6009) );
  NAND U6972 ( .A(n5881), .B(n5880), .Z(n5885) );
  NANDN U6973 ( .A(n5883), .B(n5882), .Z(n5884) );
  AND U6974 ( .A(n5885), .B(n5884), .Z(n6008) );
  XOR U6975 ( .A(n6009), .B(n6008), .Z(n6011) );
  NAND U6976 ( .A(n5887), .B(n5886), .Z(n5891) );
  NAND U6977 ( .A(n5889), .B(n5888), .Z(n5890) );
  NAND U6978 ( .A(n5891), .B(n5890), .Z(n5920) );
  NAND U6979 ( .A(n5893), .B(n5892), .Z(n5897) );
  NAND U6980 ( .A(n5895), .B(n5894), .Z(n5896) );
  NAND U6981 ( .A(n5897), .B(n5896), .Z(n5919) );
  NAND U6982 ( .A(n5899), .B(n5898), .Z(n5903) );
  NAND U6983 ( .A(n5901), .B(n5900), .Z(n5902) );
  NAND U6984 ( .A(n5903), .B(n5902), .Z(n5918) );
  XOR U6985 ( .A(n5919), .B(n5918), .Z(n5921) );
  XOR U6986 ( .A(n5920), .B(n5921), .Z(n6010) );
  XNOR U6987 ( .A(n6011), .B(n6010), .Z(n6004) );
  NANDN U6988 ( .A(n5906), .B(n5904), .Z(n5910) );
  AND U6989 ( .A(n5906), .B(n5905), .Z(n5908) );
  OR U6990 ( .A(n5908), .B(n5907), .Z(n5909) );
  AND U6991 ( .A(n5910), .B(n5909), .Z(n6002) );
  NANDN U6992 ( .A(n5912), .B(n5911), .Z(n5916) );
  NANDN U6993 ( .A(n5914), .B(n5913), .Z(n5915) );
  NAND U6994 ( .A(n5916), .B(n5915), .Z(n6003) );
  IV U6995 ( .A(n6003), .Z(n6001) );
  XNOR U6996 ( .A(n6002), .B(n6001), .Z(n5917) );
  XNOR U6997 ( .A(n6004), .B(n5917), .Z(o[5]) );
  NAND U6998 ( .A(n5919), .B(n5918), .Z(n5923) );
  NAND U6999 ( .A(n5921), .B(n5920), .Z(n5922) );
  NAND U7000 ( .A(n5923), .B(n5922), .Z(n6053) );
  NAND U7001 ( .A(n5925), .B(n5924), .Z(n5929) );
  NANDN U7002 ( .A(n5927), .B(n5926), .Z(n5928) );
  NAND U7003 ( .A(n5929), .B(n5928), .Z(n6017) );
  NAND U7004 ( .A(n5931), .B(n5930), .Z(n5935) );
  NAND U7005 ( .A(n5933), .B(n5932), .Z(n5934) );
  AND U7006 ( .A(n5935), .B(n5934), .Z(n6016) );
  NAND U7007 ( .A(n5937), .B(n5936), .Z(n5941) );
  NAND U7008 ( .A(n5939), .B(n5938), .Z(n5940) );
  AND U7009 ( .A(n5941), .B(n5940), .Z(n6015) );
  XOR U7010 ( .A(n6016), .B(n6015), .Z(n6018) );
  XOR U7011 ( .A(n6017), .B(n6018), .Z(n6054) );
  XOR U7012 ( .A(n6053), .B(n6054), .Z(n6056) );
  NAND U7013 ( .A(n5943), .B(n5942), .Z(n5947) );
  NANDN U7014 ( .A(n5945), .B(n5944), .Z(n5946) );
  NAND U7015 ( .A(n5947), .B(n5946), .Z(n6046) );
  NAND U7016 ( .A(n5949), .B(n5948), .Z(n5953) );
  NAND U7017 ( .A(n5951), .B(n5950), .Z(n5952) );
  NAND U7018 ( .A(n5953), .B(n5952), .Z(n6044) );
  NAND U7019 ( .A(n5955), .B(n5954), .Z(n5959) );
  NAND U7020 ( .A(n5957), .B(n5956), .Z(n5958) );
  NAND U7021 ( .A(n5959), .B(n5958), .Z(n6041) );
  NAND U7022 ( .A(n5960), .B(oglobal[5]), .Z(n5964) );
  NAND U7023 ( .A(n5962), .B(n5961), .Z(n5963) );
  NAND U7024 ( .A(n5964), .B(n5963), .Z(n6033) );
  XOR U7025 ( .A(n6033), .B(oglobal[6]), .Z(n6035) );
  NAND U7026 ( .A(n5966), .B(n5965), .Z(n5970) );
  NAND U7027 ( .A(n5968), .B(n5967), .Z(n5969) );
  NAND U7028 ( .A(n5970), .B(n5969), .Z(n6034) );
  XNOR U7029 ( .A(n6035), .B(n6034), .Z(n6029) );
  NAND U7030 ( .A(n5972), .B(n5971), .Z(n5976) );
  NAND U7031 ( .A(n5974), .B(n5973), .Z(n5975) );
  NAND U7032 ( .A(n5976), .B(n5975), .Z(n6027) );
  NAND U7033 ( .A(n5978), .B(n5977), .Z(n5982) );
  NAND U7034 ( .A(n5980), .B(n5979), .Z(n5981) );
  AND U7035 ( .A(n5982), .B(n5981), .Z(n6028) );
  XOR U7036 ( .A(n6027), .B(n6028), .Z(n6030) );
  NAND U7037 ( .A(n5984), .B(n5983), .Z(n5988) );
  NAND U7038 ( .A(n5986), .B(n5985), .Z(n5987) );
  NAND U7039 ( .A(n5988), .B(n5987), .Z(n6038) );
  XOR U7040 ( .A(n6039), .B(n6038), .Z(n6040) );
  NAND U7041 ( .A(n5990), .B(n5989), .Z(n5994) );
  NAND U7042 ( .A(n5992), .B(n5991), .Z(n5993) );
  AND U7043 ( .A(n5994), .B(n5993), .Z(n6021) );
  NAND U7044 ( .A(n5996), .B(n5995), .Z(n6000) );
  NAND U7045 ( .A(n5998), .B(n5997), .Z(n5999) );
  AND U7046 ( .A(n6000), .B(n5999), .Z(n6022) );
  XOR U7047 ( .A(n6023), .B(n6024), .Z(n6045) );
  XOR U7048 ( .A(n6044), .B(n6045), .Z(n6047) );
  XOR U7049 ( .A(n6046), .B(n6047), .Z(n6055) );
  XNOR U7050 ( .A(n6056), .B(n6055), .Z(n6050) );
  NAND U7051 ( .A(n6001), .B(n6002), .Z(n6007) );
  ANDN U7052 ( .B(n6003), .A(n6002), .Z(n6005) );
  OR U7053 ( .A(n6005), .B(n6004), .Z(n6006) );
  AND U7054 ( .A(n6007), .B(n6006), .Z(n6051) );
  NAND U7055 ( .A(n6009), .B(n6008), .Z(n6013) );
  NAND U7056 ( .A(n6011), .B(n6010), .Z(n6012) );
  AND U7057 ( .A(n6013), .B(n6012), .Z(n6052) );
  XNOR U7058 ( .A(n6051), .B(n6052), .Z(n6014) );
  XNOR U7059 ( .A(n6050), .B(n6014), .Z(o[6]) );
  NAND U7060 ( .A(n6016), .B(n6015), .Z(n6020) );
  NAND U7061 ( .A(n6018), .B(n6017), .Z(n6019) );
  NAND U7062 ( .A(n6020), .B(n6019), .Z(n6060) );
  NAND U7063 ( .A(n6022), .B(n6021), .Z(n6026) );
  NAND U7064 ( .A(n6024), .B(n6023), .Z(n6025) );
  NAND U7065 ( .A(n6026), .B(n6025), .Z(n6069) );
  NAND U7066 ( .A(n6028), .B(n6027), .Z(n6032) );
  NAND U7067 ( .A(n6030), .B(n6029), .Z(n6031) );
  AND U7068 ( .A(n6032), .B(n6031), .Z(n6072) );
  XOR U7069 ( .A(oglobal[7]), .B(n6072), .Z(n6074) );
  NAND U7070 ( .A(oglobal[6]), .B(n6033), .Z(n6037) );
  NAND U7071 ( .A(n6035), .B(n6034), .Z(n6036) );
  NAND U7072 ( .A(n6037), .B(n6036), .Z(n6073) );
  XNOR U7073 ( .A(n6074), .B(n6073), .Z(n6067) );
  NAND U7074 ( .A(n6039), .B(n6038), .Z(n6043) );
  NAND U7075 ( .A(n6041), .B(n6040), .Z(n6042) );
  AND U7076 ( .A(n6043), .B(n6042), .Z(n6066) );
  XOR U7077 ( .A(n6060), .B(n6061), .Z(n6063) );
  NAND U7078 ( .A(n6045), .B(n6044), .Z(n6049) );
  NAND U7079 ( .A(n6047), .B(n6046), .Z(n6048) );
  NAND U7080 ( .A(n6049), .B(n6048), .Z(n6062) );
  XNOR U7081 ( .A(n6063), .B(n6062), .Z(n6077) );
  NAND U7082 ( .A(n6054), .B(n6053), .Z(n6058) );
  NAND U7083 ( .A(n6056), .B(n6055), .Z(n6057) );
  AND U7084 ( .A(n6058), .B(n6057), .Z(n6079) );
  XNOR U7085 ( .A(n6078), .B(n6079), .Z(n6059) );
  XNOR U7086 ( .A(n6077), .B(n6059), .Z(o[7]) );
  NAND U7087 ( .A(n6061), .B(n6060), .Z(n6065) );
  NAND U7088 ( .A(n6063), .B(n6062), .Z(n6064) );
  AND U7089 ( .A(n6065), .B(n6064), .Z(n6088) );
  NAND U7090 ( .A(n6067), .B(n6066), .Z(n6071) );
  NAND U7091 ( .A(n6069), .B(n6068), .Z(n6070) );
  AND U7092 ( .A(n6071), .B(n6070), .Z(n6083) );
  NAND U7093 ( .A(n6072), .B(oglobal[7]), .Z(n6076) );
  NAND U7094 ( .A(n6074), .B(n6073), .Z(n6075) );
  NAND U7095 ( .A(n6076), .B(n6075), .Z(n6081) );
  XOR U7096 ( .A(oglobal[8]), .B(n6081), .Z(n6082) );
  XOR U7097 ( .A(n6083), .B(n6082), .Z(n6087) );
  XNOR U7098 ( .A(n6087), .B(n6086), .Z(n6080) );
  XNOR U7099 ( .A(n6088), .B(n6080), .Z(o[8]) );
  NAND U7100 ( .A(oglobal[8]), .B(n6081), .Z(n6085) );
  NAND U7101 ( .A(n6083), .B(n6082), .Z(n6084) );
  NAND U7102 ( .A(n6085), .B(n6084), .Z(n6091) );
  XNOR U7103 ( .A(oglobal[9]), .B(n6090), .Z(n6089) );
  XNOR U7104 ( .A(n6091), .B(n6089), .Z(o[9]) );
  XOR U7105 ( .A(n6092), .B(oglobal[10]), .Z(o[10]) );
  AND U7106 ( .A(n6092), .B(oglobal[10]), .Z(n6093) );
  XOR U7107 ( .A(n6093), .B(oglobal[11]), .Z(o[11]) );
  NAND U7108 ( .A(n6093), .B(oglobal[11]), .Z(n6094) );
  XNOR U7109 ( .A(oglobal[12]), .B(n6094), .Z(o[12]) );
  NANDN U7110 ( .A(n6094), .B(oglobal[12]), .Z(n6095) );
  XNOR U7111 ( .A(oglobal[13]), .B(n6095), .Z(o[13]) );
endmodule

