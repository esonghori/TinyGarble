
module hamming_N1600_CC2 ( clk, rst, x, y, o );
  input [799:0] x;
  input [799:0] y;
  output [10:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845;
  wire   [10:0] oglobal;

  DFF \oglobal_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .Q(oglobal[10]) );
  DFF \oglobal_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .Q(oglobal[9]) );
  DFF \oglobal_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .Q(oglobal[8]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(oglobal[7]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(oglobal[6]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(oglobal[5]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(oglobal[4]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(oglobal[3]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(oglobal[2]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(oglobal[1]) );
  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(oglobal[0]) );
  NAND U803 ( .A(n3532), .B(n3533), .Z(n1) );
  XOR U804 ( .A(n3532), .B(n3533), .Z(n2) );
  NANDN U805 ( .A(n3531), .B(n2), .Z(n3) );
  NAND U806 ( .A(n1), .B(n3), .Z(n3786) );
  XOR U807 ( .A(n4218), .B(n4217), .Z(n3854) );
  XOR U808 ( .A(n1158), .B(n1157), .Z(n1159) );
  XOR U809 ( .A(n2871), .B(n2870), .Z(n2872) );
  XOR U810 ( .A(n2630), .B(n2629), .Z(n2632) );
  NAND U811 ( .A(n579), .B(n580), .Z(n4) );
  NANDN U812 ( .A(n577), .B(n578), .Z(n5) );
  NAND U813 ( .A(n4), .B(n5), .Z(n3487) );
  XOR U814 ( .A(n3569), .B(n3568), .Z(n3570) );
  XOR U815 ( .A(n3545), .B(n3544), .Z(n6) );
  NANDN U816 ( .A(n3543), .B(n6), .Z(n7) );
  NAND U817 ( .A(n3545), .B(n3544), .Z(n8) );
  AND U818 ( .A(n7), .B(n8), .Z(n4221) );
  NAND U819 ( .A(n3006), .B(n3005), .Z(n9) );
  XOR U820 ( .A(n3006), .B(n3005), .Z(n10) );
  NANDN U821 ( .A(n3007), .B(n10), .Z(n11) );
  NAND U822 ( .A(n9), .B(n11), .Z(n3853) );
  XOR U823 ( .A(n3789), .B(n3788), .Z(n4118) );
  NAND U824 ( .A(n3356), .B(n3357), .Z(n12) );
  XOR U825 ( .A(n3356), .B(n3357), .Z(n13) );
  NANDN U826 ( .A(n3355), .B(n13), .Z(n14) );
  NAND U827 ( .A(n12), .B(n14), .Z(n3859) );
  XOR U828 ( .A(n4497), .B(n4496), .Z(n15) );
  XNOR U829 ( .A(n4499), .B(n15), .Z(n4318) );
  NAND U830 ( .A(n3857), .B(n3858), .Z(n16) );
  XOR U831 ( .A(n3857), .B(n3858), .Z(n17) );
  NANDN U832 ( .A(n3856), .B(n17), .Z(n18) );
  NAND U833 ( .A(n16), .B(n18), .Z(n4458) );
  XOR U834 ( .A(n4382), .B(n4381), .Z(n4387) );
  XOR U835 ( .A(n369), .B(n368), .Z(n370) );
  XOR U836 ( .A(n634), .B(n633), .Z(n635) );
  XOR U837 ( .A(n893), .B(n892), .Z(n894) );
  XOR U838 ( .A(n3657), .B(n3656), .Z(n3658) );
  XOR U839 ( .A(n3310), .B(n3309), .Z(n3312) );
  XOR U840 ( .A(n3046), .B(n3045), .Z(n3048) );
  XOR U841 ( .A(n3022), .B(n3021), .Z(n3024) );
  XOR U842 ( .A(n2684), .B(n2683), .Z(n2685) );
  NAND U843 ( .A(n1089), .B(n1090), .Z(n19) );
  NANDN U844 ( .A(n1087), .B(n1088), .Z(n20) );
  NAND U845 ( .A(n19), .B(n20), .Z(n3384) );
  NAND U846 ( .A(n420), .B(n419), .Z(n21) );
  NANDN U847 ( .A(n417), .B(n418), .Z(n22) );
  AND U848 ( .A(n21), .B(n22), .Z(n3513) );
  XOR U849 ( .A(n3487), .B(n3486), .Z(n3488) );
  XOR U850 ( .A(n2873), .B(n2872), .Z(n3354) );
  NAND U851 ( .A(n2825), .B(n2827), .Z(n23) );
  XOR U852 ( .A(n2825), .B(n2827), .Z(n24) );
  NAND U853 ( .A(n24), .B(n2826), .Z(n25) );
  NAND U854 ( .A(n23), .B(n25), .Z(n3771) );
  NAND U855 ( .A(n3632), .B(n3633), .Z(n26) );
  XOR U856 ( .A(n3632), .B(n3633), .Z(n27) );
  NANDN U857 ( .A(n3631), .B(n27), .Z(n28) );
  NAND U858 ( .A(n26), .B(n28), .Z(n4160) );
  XOR U859 ( .A(n4210), .B(n4209), .Z(n4211) );
  NAND U860 ( .A(n3318), .B(n3320), .Z(n29) );
  XOR U861 ( .A(n3318), .B(n3320), .Z(n30) );
  NAND U862 ( .A(n30), .B(n3319), .Z(n31) );
  NAND U863 ( .A(n29), .B(n31), .Z(n4111) );
  XNOR U864 ( .A(n3970), .B(n3969), .Z(n4205) );
  XOR U865 ( .A(n4152), .B(n4153), .Z(n32) );
  XNOR U866 ( .A(n4151), .B(n32), .Z(n3795) );
  XOR U867 ( .A(n3528), .B(n3529), .Z(n33) );
  NANDN U868 ( .A(n3530), .B(n33), .Z(n34) );
  NAND U869 ( .A(n3528), .B(n3529), .Z(n35) );
  AND U870 ( .A(n34), .B(n35), .Z(n3787) );
  NAND U871 ( .A(n3547), .B(n3548), .Z(n36) );
  XOR U872 ( .A(n3547), .B(n3548), .Z(n37) );
  NANDN U873 ( .A(n3546), .B(n37), .Z(n38) );
  NAND U874 ( .A(n36), .B(n38), .Z(n4117) );
  XOR U875 ( .A(n4141), .B(n4140), .Z(n3875) );
  XOR U876 ( .A(n4467), .B(n4466), .Z(n4468) );
  XOR U877 ( .A(n4114), .B(n4115), .Z(n39) );
  NANDN U878 ( .A(n4116), .B(n39), .Z(n40) );
  NAND U879 ( .A(n4114), .B(n4115), .Z(n41) );
  AND U880 ( .A(n40), .B(n41), .Z(n4481) );
  XNOR U881 ( .A(n4463), .B(n4462), .Z(n4320) );
  NAND U882 ( .A(n4103), .B(n4104), .Z(n42) );
  XOR U883 ( .A(n4103), .B(n4104), .Z(n43) );
  NANDN U884 ( .A(n4102), .B(n43), .Z(n44) );
  NAND U885 ( .A(n42), .B(n44), .Z(n4455) );
  NAND U886 ( .A(n4473), .B(n4474), .Z(n45) );
  XOR U887 ( .A(n4473), .B(n4474), .Z(n46) );
  NANDN U888 ( .A(n4472), .B(n46), .Z(n47) );
  NAND U889 ( .A(n45), .B(n47), .Z(n4606) );
  NAND U890 ( .A(n4328), .B(n4329), .Z(n48) );
  XOR U891 ( .A(n4328), .B(n4329), .Z(n49) );
  NANDN U892 ( .A(n4327), .B(n49), .Z(n50) );
  NAND U893 ( .A(n48), .B(n50), .Z(n4644) );
  XNOR U894 ( .A(n4620), .B(n4619), .Z(n4648) );
  NAND U895 ( .A(n4457), .B(n4456), .Z(n51) );
  XOR U896 ( .A(n4457), .B(n4456), .Z(n52) );
  NANDN U897 ( .A(n4458), .B(n52), .Z(n53) );
  NAND U898 ( .A(n51), .B(n53), .Z(n4654) );
  XOR U899 ( .A(n4018), .B(n4017), .Z(n3706) );
  XOR U900 ( .A(n4362), .B(n4361), .Z(n4363) );
  XNOR U901 ( .A(n4804), .B(n4803), .Z(n4806) );
  NAND U902 ( .A(n4672), .B(n4673), .Z(n54) );
  XOR U903 ( .A(n4672), .B(n4673), .Z(n55) );
  NAND U904 ( .A(n55), .B(n4671), .Z(n56) );
  NAND U905 ( .A(n54), .B(n56), .Z(n4711) );
  XOR U906 ( .A(n562), .B(n561), .Z(n563) );
  XOR U907 ( .A(n2072), .B(n2071), .Z(n2073) );
  XOR U908 ( .A(n1805), .B(n1804), .Z(n1806) );
  XOR U909 ( .A(n640), .B(n639), .Z(n641) );
  XOR U910 ( .A(n2371), .B(n2370), .Z(n2372) );
  XOR U911 ( .A(n1505), .B(n1504), .Z(n1506) );
  XOR U912 ( .A(n716), .B(n715), .Z(n717) );
  XOR U913 ( .A(n1499), .B(n1498), .Z(n1500) );
  XOR U914 ( .A(n2365), .B(n2364), .Z(n2366) );
  XOR U915 ( .A(n1823), .B(n1822), .Z(n1824) );
  XOR U916 ( .A(n2261), .B(n2260), .Z(n2262) );
  XOR U917 ( .A(n2273), .B(n2272), .Z(n2274) );
  XOR U918 ( .A(n2865), .B(n2864), .Z(n2867) );
  XOR U919 ( .A(n2624), .B(n2623), .Z(n2626) );
  XOR U920 ( .A(n2636), .B(n2635), .Z(n2638) );
  XOR U921 ( .A(n3335), .B(n3334), .Z(n3337) );
  XOR U922 ( .A(n2799), .B(n2798), .Z(n2801) );
  XOR U923 ( .A(n2793), .B(n2792), .Z(n2795) );
  XOR U924 ( .A(n3557), .B(n3556), .Z(n3559) );
  XOR U925 ( .A(n3040), .B(n3039), .Z(n3042) );
  XOR U926 ( .A(n3010), .B(n3009), .Z(n3012) );
  XOR U927 ( .A(n2757), .B(n2756), .Z(n2759) );
  XOR U928 ( .A(n2763), .B(n2762), .Z(n2765) );
  XOR U929 ( .A(n2751), .B(n2750), .Z(n2753) );
  NAND U930 ( .A(n308), .B(n309), .Z(n57) );
  NANDN U931 ( .A(n306), .B(n307), .Z(n58) );
  NAND U932 ( .A(n57), .B(n58), .Z(n3475) );
  XNOR U933 ( .A(n3529), .B(n3528), .Z(n59) );
  XNOR U934 ( .A(n3530), .B(n59), .Z(n2643) );
  XOR U935 ( .A(n3366), .B(n3365), .Z(n3368) );
  XOR U936 ( .A(n3360), .B(n3359), .Z(n3361) );
  NAND U937 ( .A(n484), .B(n483), .Z(n60) );
  NANDN U938 ( .A(n481), .B(n482), .Z(n61) );
  AND U939 ( .A(n60), .B(n61), .Z(n3499) );
  XOR U940 ( .A(n899), .B(n898), .Z(n900) );
  XOR U941 ( .A(n2267), .B(n2266), .Z(n2268) );
  XOR U942 ( .A(n2907), .B(n2906), .Z(n2908) );
  XOR U943 ( .A(n3456), .B(n3455), .Z(n3457) );
  NAND U944 ( .A(n366), .B(n367), .Z(n62) );
  NANDN U945 ( .A(n364), .B(n365), .Z(n63) );
  NAND U946 ( .A(n62), .B(n63), .Z(n3450) );
  NAND U947 ( .A(n575), .B(n576), .Z(n64) );
  NANDN U948 ( .A(n573), .B(n574), .Z(n65) );
  NAND U949 ( .A(n64), .B(n65), .Z(n3489) );
  XOR U950 ( .A(n2722), .B(n2723), .Z(n66) );
  XNOR U951 ( .A(n2724), .B(n66), .Z(n3379) );
  XOR U952 ( .A(n3347), .B(n3346), .Z(n3348) );
  NANDN U953 ( .A(n695), .B(n696), .Z(n67) );
  NANDN U954 ( .A(n693), .B(n694), .Z(n68) );
  AND U955 ( .A(n67), .B(n68), .Z(n3298) );
  XOR U956 ( .A(n3386), .B(n3385), .Z(n3516) );
  XOR U957 ( .A(n3778), .B(n3777), .Z(n3779) );
  NAND U958 ( .A(n2823), .B(n2824), .Z(n69) );
  XOR U959 ( .A(n2823), .B(n2824), .Z(n70) );
  NANDN U960 ( .A(n2822), .B(n70), .Z(n71) );
  NAND U961 ( .A(n69), .B(n71), .Z(n3772) );
  XOR U962 ( .A(n3882), .B(n3881), .Z(n3883) );
  NAND U963 ( .A(n3541), .B(n3542), .Z(n72) );
  XOR U964 ( .A(n3541), .B(n3542), .Z(n73) );
  NANDN U965 ( .A(n3540), .B(n73), .Z(n74) );
  NAND U966 ( .A(n72), .B(n74), .Z(n4222) );
  XOR U967 ( .A(n4134), .B(n4133), .Z(n4135) );
  XOR U968 ( .A(n3760), .B(n3759), .Z(n3761) );
  XOR U969 ( .A(n3766), .B(n3765), .Z(n3767) );
  NAND U970 ( .A(n2714), .B(n2715), .Z(n75) );
  XOR U971 ( .A(n2714), .B(n2715), .Z(n76) );
  NANDN U972 ( .A(n2713), .B(n76), .Z(n77) );
  NAND U973 ( .A(n75), .B(n77), .Z(n4114) );
  NAND U974 ( .A(n3316), .B(n3317), .Z(n78) );
  XOR U975 ( .A(n3316), .B(n3317), .Z(n79) );
  NANDN U976 ( .A(n3315), .B(n79), .Z(n80) );
  NAND U977 ( .A(n78), .B(n80), .Z(n4112) );
  XOR U978 ( .A(n3974), .B(n3973), .Z(n3975) );
  XOR U979 ( .A(n3937), .B(n3936), .Z(n3939) );
  XOR U980 ( .A(n3811), .B(n3810), .Z(n3812) );
  XOR U981 ( .A(n3817), .B(n3816), .Z(n3818) );
  XOR U982 ( .A(n4254), .B(n4253), .Z(n3869) );
  NAND U983 ( .A(n3636), .B(n3637), .Z(n81) );
  XOR U984 ( .A(n3636), .B(n3637), .Z(n82) );
  NANDN U985 ( .A(n3635), .B(n82), .Z(n83) );
  NAND U986 ( .A(n81), .B(n83), .Z(n3876) );
  XOR U987 ( .A(n353), .B(n352), .Z(n354) );
  XOR U988 ( .A(n331), .B(n330), .Z(n2218) );
  XOR U989 ( .A(n3374), .B(n3373), .Z(n3159) );
  XOR U990 ( .A(n3462), .B(n3461), .Z(n3463) );
  NAND U991 ( .A(n3353), .B(n3354), .Z(n84) );
  XOR U992 ( .A(n3353), .B(n3354), .Z(n85) );
  NANDN U993 ( .A(n3352), .B(n85), .Z(n86) );
  NAND U994 ( .A(n84), .B(n86), .Z(n3860) );
  XOR U995 ( .A(n3931), .B(n3930), .Z(n3933) );
  NANDN U996 ( .A(n931), .B(n932), .Z(n87) );
  NANDN U997 ( .A(n929), .B(n930), .Z(n88) );
  AND U998 ( .A(n87), .B(n88), .Z(n3100) );
  XOR U999 ( .A(n4295), .B(n4294), .Z(n4296) );
  XOR U1000 ( .A(n4319), .B(n4318), .Z(n4321) );
  XOR U1001 ( .A(n4434), .B(n4433), .Z(n4435) );
  NAND U1002 ( .A(n3854), .B(n3855), .Z(n89) );
  XOR U1003 ( .A(n3854), .B(n3855), .Z(n90) );
  NAND U1004 ( .A(n90), .B(n3853), .Z(n91) );
  NAND U1005 ( .A(n89), .B(n91), .Z(n4456) );
  XNOR U1006 ( .A(n4303), .B(n4302), .Z(n4513) );
  NAND U1007 ( .A(n4494), .B(n4495), .Z(n92) );
  XOR U1008 ( .A(n4494), .B(n4495), .Z(n93) );
  NANDN U1009 ( .A(n4493), .B(n93), .Z(n94) );
  NAND U1010 ( .A(n92), .B(n94), .Z(n4613) );
  XOR U1011 ( .A(n4607), .B(n4606), .Z(n4608) );
  XOR U1012 ( .A(n4601), .B(n4600), .Z(n4603) );
  NAND U1013 ( .A(n4325), .B(n4326), .Z(n95) );
  XOR U1014 ( .A(n4325), .B(n4326), .Z(n96) );
  NANDN U1015 ( .A(n4324), .B(n96), .Z(n97) );
  NAND U1016 ( .A(n95), .B(n97), .Z(n4645) );
  XOR U1017 ( .A(n4455), .B(n4453), .Z(n98) );
  NANDN U1018 ( .A(n4454), .B(n98), .Z(n99) );
  NAND U1019 ( .A(n4455), .B(n4453), .Z(n100) );
  AND U1020 ( .A(n99), .B(n100), .Z(n4653) );
  XNOR U1021 ( .A(n1481), .B(n1480), .Z(n1483) );
  XOR U1022 ( .A(n4751), .B(n4750), .Z(n4752) );
  XOR U1023 ( .A(n4798), .B(n4797), .Z(n4799) );
  XNOR U1024 ( .A(n4022), .B(n4021), .Z(n4024) );
  XOR U1025 ( .A(n4270), .B(n4269), .Z(n4272) );
  XNOR U1026 ( .A(n4567), .B(n4566), .Z(n4559) );
  XOR U1027 ( .A(n3699), .B(n3698), .Z(n3701) );
  XNOR U1028 ( .A(n4666), .B(n4665), .Z(n4668) );
  XOR U1029 ( .A(n4555), .B(n4554), .Z(n101) );
  NANDN U1030 ( .A(n4556), .B(n101), .Z(n102) );
  NAND U1031 ( .A(n4555), .B(n4554), .Z(n103) );
  AND U1032 ( .A(n102), .B(n103), .Z(n4671) );
  NAND U1033 ( .A(n4783), .B(n4784), .Z(n104) );
  XOR U1034 ( .A(n4783), .B(n4784), .Z(n105) );
  NANDN U1035 ( .A(n4782), .B(n105), .Z(n106) );
  NAND U1036 ( .A(n104), .B(n106), .Z(n4819) );
  XOR U1037 ( .A(n2437), .B(n2436), .Z(n2438) );
  XOR U1038 ( .A(n2449), .B(n2448), .Z(n2450) );
  XOR U1039 ( .A(n2419), .B(n2418), .Z(n2420) );
  XOR U1040 ( .A(n2127), .B(n2126), .Z(n2128) );
  XOR U1041 ( .A(n1817), .B(n1816), .Z(n1818) );
  XOR U1042 ( .A(n1565), .B(n1564), .Z(n1566) );
  XOR U1043 ( .A(n510), .B(n509), .Z(n511) );
  XOR U1044 ( .A(n2249), .B(n2248), .Z(n2250) );
  XOR U1045 ( .A(n2389), .B(n2388), .Z(n2390) );
  XOR U1046 ( .A(n2383), .B(n2382), .Z(n2384) );
  XOR U1047 ( .A(n2395), .B(n2394), .Z(n2396) );
  XOR U1048 ( .A(n582), .B(n581), .Z(n583) );
  XOR U1049 ( .A(n2401), .B(n2400), .Z(n2402) );
  XOR U1050 ( .A(n2353), .B(n2352), .Z(n2354) );
  XOR U1051 ( .A(n1956), .B(n1955), .Z(n1957) );
  XOR U1052 ( .A(n1914), .B(n1913), .Z(n1915) );
  XOR U1053 ( .A(n1920), .B(n1919), .Z(n1921) );
  XOR U1054 ( .A(n1583), .B(n1582), .Z(n1584) );
  XOR U1055 ( .A(n2310), .B(n2309), .Z(n2311) );
  XOR U1056 ( .A(n2304), .B(n2303), .Z(n2305) );
  XOR U1057 ( .A(n604), .B(n603), .Z(n605) );
  XOR U1058 ( .A(n2485), .B(n2484), .Z(n2486) );
  XOR U1059 ( .A(n646), .B(n645), .Z(n647) );
  XOR U1060 ( .A(n2377), .B(n2376), .Z(n2378) );
  XOR U1061 ( .A(n1321), .B(n1320), .Z(n1322) );
  XOR U1062 ( .A(n2102), .B(n2101), .Z(n2103) );
  XOR U1063 ( .A(n2108), .B(n2107), .Z(n2109) );
  XOR U1064 ( .A(n1363), .B(n1362), .Z(n1364) );
  XOR U1065 ( .A(n1369), .B(n1368), .Z(n1370) );
  XOR U1066 ( .A(n2527), .B(n2526), .Z(n2528) );
  XOR U1067 ( .A(n1751), .B(n1750), .Z(n1752) );
  XOR U1068 ( .A(n856), .B(n855), .Z(n857) );
  XOR U1069 ( .A(n458), .B(n457), .Z(n459) );
  XOR U1070 ( .A(n1883), .B(n1882), .Z(n1884) );
  XOR U1071 ( .A(n1950), .B(n1949), .Z(n1951) );
  XOR U1072 ( .A(n1908), .B(n1907), .Z(n1909) );
  XOR U1073 ( .A(n2121), .B(n2120), .Z(n2122) );
  XOR U1074 ( .A(n1242), .B(n1241), .Z(n1243) );
  XOR U1075 ( .A(n1787), .B(n1786), .Z(n1788) );
  XOR U1076 ( .A(n2359), .B(n2358), .Z(n2360) );
  XOR U1077 ( .A(n2431), .B(n2430), .Z(n2432) );
  XOR U1078 ( .A(n2407), .B(n2406), .Z(n2408) );
  XOR U1079 ( .A(n2425), .B(n2424), .Z(n2426) );
  XOR U1080 ( .A(n1327), .B(n1326), .Z(n1328) );
  XOR U1081 ( .A(n1841), .B(n1840), .Z(n1842) );
  XOR U1082 ( .A(n1835), .B(n1834), .Z(n1836) );
  XOR U1083 ( .A(n1589), .B(n1588), .Z(n1590) );
  XOR U1084 ( .A(n2243), .B(n2242), .Z(n2244) );
  XOR U1085 ( .A(n1733), .B(n1732), .Z(n1734) );
  XOR U1086 ( .A(n2066), .B(n2065), .Z(n2067) );
  XOR U1087 ( .A(n1811), .B(n1810), .Z(n1812) );
  XOR U1088 ( .A(n2096), .B(n2095), .Z(n2097) );
  XOR U1089 ( .A(n2413), .B(n2412), .Z(n2414) );
  XOR U1090 ( .A(n2297), .B(n2296), .Z(n2298) );
  XOR U1091 ( .A(n2316), .B(n2315), .Z(n2317) );
  XOR U1092 ( .A(n2255), .B(n2254), .Z(n2256) );
  XOR U1093 ( .A(n1974), .B(n1973), .Z(n1975) );
  XOR U1094 ( .A(n550), .B(n549), .Z(n551) );
  XOR U1095 ( .A(n2285), .B(n2284), .Z(n2286) );
  XOR U1096 ( .A(n2291), .B(n2290), .Z(n2292) );
  XOR U1097 ( .A(n588), .B(n587), .Z(n589) );
  XOR U1098 ( .A(n2817), .B(n2816), .Z(n2819) );
  XOR U1099 ( .A(n3623), .B(n3622), .Z(n3625) );
  XOR U1100 ( .A(n2859), .B(n2858), .Z(n2861) );
  XOR U1101 ( .A(n2805), .B(n2804), .Z(n2807) );
  XOR U1102 ( .A(n3645), .B(n3644), .Z(n3646) );
  XOR U1103 ( .A(n2678), .B(n2677), .Z(n2680) );
  XOR U1104 ( .A(n2672), .B(n2671), .Z(n2674) );
  XOR U1105 ( .A(n2666), .B(n2665), .Z(n2668) );
  XOR U1106 ( .A(n2660), .B(n2659), .Z(n2662) );
  XOR U1107 ( .A(n2717), .B(n2716), .Z(n2719) );
  XOR U1108 ( .A(n2642), .B(n2641), .Z(n2644) );
  XOR U1109 ( .A(n3319), .B(n3320), .Z(n107) );
  XNOR U1110 ( .A(n3318), .B(n107), .Z(n3367) );
  XOR U1111 ( .A(n2925), .B(n2924), .Z(n2926) );
  XOR U1112 ( .A(n3384), .B(n3383), .Z(n3385) );
  XOR U1113 ( .A(n3659), .B(n3658), .Z(n3637) );
  XOR U1114 ( .A(n862), .B(n861), .Z(n863) );
  XOR U1115 ( .A(n1944), .B(n1943), .Z(n1945) );
  XOR U1116 ( .A(n2151), .B(n2150), .Z(n2152) );
  XOR U1117 ( .A(n1775), .B(n1774), .Z(n1776) );
  XOR U1118 ( .A(n2443), .B(n2442), .Z(n2444) );
  XOR U1119 ( .A(n1757), .B(n1756), .Z(n1758) );
  XOR U1120 ( .A(n1571), .B(n1570), .Z(n1572) );
  XOR U1121 ( .A(n1595), .B(n1594), .Z(n1596) );
  XOR U1122 ( .A(n329), .B(n328), .Z(n330) );
  XOR U1123 ( .A(n1493), .B(n1492), .Z(n1495) );
  XOR U1124 ( .A(n1619), .B(n1618), .Z(n1621) );
  XOR U1125 ( .A(n1932), .B(n1931), .Z(n1934) );
  XOR U1126 ( .A(n1938), .B(n1937), .Z(n1940) );
  XOR U1127 ( .A(n1727), .B(n1726), .Z(n1728) );
  XOR U1128 ( .A(n2060), .B(n2059), .Z(n2061) );
  XOR U1129 ( .A(n3372), .B(n3371), .Z(n3373) );
  XOR U1130 ( .A(n2901), .B(n2900), .Z(n2903) );
  XOR U1131 ( .A(n3481), .B(n3480), .Z(n3482) );
  XOR U1132 ( .A(n3475), .B(n3474), .Z(n3476) );
  NAND U1133 ( .A(n602), .B(n601), .Z(n108) );
  NANDN U1134 ( .A(n599), .B(n600), .Z(n109) );
  AND U1135 ( .A(n108), .B(n109), .Z(n3507) );
  XOR U1136 ( .A(n3378), .B(n3377), .Z(n3380) );
  XOR U1137 ( .A(n3432), .B(n3431), .Z(n3433) );
  XOR U1138 ( .A(n2686), .B(n2685), .Z(n3201) );
  XOR U1139 ( .A(n3349), .B(n3348), .Z(n3517) );
  XOR U1140 ( .A(n3362), .B(n3361), .Z(n2556) );
  NANDN U1141 ( .A(n935), .B(n936), .Z(n110) );
  NANDN U1142 ( .A(n933), .B(n934), .Z(n111) );
  AND U1143 ( .A(n110), .B(n111), .Z(n3682) );
  XOR U1144 ( .A(n4252), .B(n4251), .Z(n4253) );
  NAND U1145 ( .A(n3629), .B(n3630), .Z(n112) );
  XOR U1146 ( .A(n3629), .B(n3630), .Z(n113) );
  NANDN U1147 ( .A(n3628), .B(n113), .Z(n114) );
  NAND U1148 ( .A(n112), .B(n114), .Z(n4161) );
  XOR U1149 ( .A(n4155), .B(n4154), .Z(n4156) );
  NAND U1150 ( .A(n2979), .B(n2980), .Z(n115) );
  XOR U1151 ( .A(n2979), .B(n2980), .Z(n116) );
  NANDN U1152 ( .A(n2978), .B(n116), .Z(n117) );
  NAND U1153 ( .A(n115), .B(n117), .Z(n4216) );
  NAND U1154 ( .A(n2722), .B(n2724), .Z(n118) );
  XOR U1155 ( .A(n2722), .B(n2724), .Z(n119) );
  NAND U1156 ( .A(n119), .B(n2723), .Z(n120) );
  NAND U1157 ( .A(n118), .B(n120), .Z(n4115) );
  XOR U1158 ( .A(n4106), .B(n4105), .Z(n4107) );
  XOR U1159 ( .A(n3968), .B(n3967), .Z(n3969) );
  XOR U1160 ( .A(n3962), .B(n3961), .Z(n3963) );
  XNOR U1161 ( .A(n3976), .B(n3975), .Z(n3938) );
  XNOR U1162 ( .A(n3780), .B(n3779), .Z(n3736) );
  XOR U1163 ( .A(n4212), .B(n4211), .Z(n3855) );
  XOR U1164 ( .A(n3884), .B(n3883), .Z(n3870) );
  XOR U1165 ( .A(n4136), .B(n4135), .Z(n3877) );
  XOR U1166 ( .A(n2163), .B(n2162), .Z(n2164) );
  XOR U1167 ( .A(n1763), .B(n1762), .Z(n1764) );
  XOR U1168 ( .A(n1577), .B(n1576), .Z(n1578) );
  XOR U1169 ( .A(n1517), .B(n1516), .Z(n1519) );
  XOR U1170 ( .A(n1721), .B(n1720), .Z(n1723) );
  XOR U1171 ( .A(n2825), .B(n2826), .Z(n121) );
  XNOR U1172 ( .A(n2827), .B(n121), .Z(n3574) );
  XOR U1173 ( .A(n2909), .B(n2908), .Z(n3160) );
  XOR U1174 ( .A(n3458), .B(n3457), .Z(n3190) );
  XOR U1175 ( .A(n3450), .B(n3449), .Z(n3451) );
  XOR U1176 ( .A(n3489), .B(n3488), .Z(n3167) );
  XNOR U1177 ( .A(n3762), .B(n3761), .Z(n3932) );
  XNOR U1178 ( .A(n3813), .B(n3812), .Z(n3863) );
  XOR U1179 ( .A(n3819), .B(n3818), .Z(n4227) );
  NAND U1180 ( .A(n3784), .B(n3785), .Z(n122) );
  XOR U1181 ( .A(n3784), .B(n3785), .Z(n123) );
  NANDN U1182 ( .A(n3783), .B(n123), .Z(n124) );
  NAND U1183 ( .A(n122), .B(n124), .Z(n4497) );
  NAND U1184 ( .A(n4151), .B(n4153), .Z(n125) );
  XOR U1185 ( .A(n4151), .B(n4153), .Z(n126) );
  NAND U1186 ( .A(n126), .B(n4152), .Z(n127) );
  NAND U1187 ( .A(n125), .B(n127), .Z(n4493) );
  XOR U1188 ( .A(n4488), .B(n4487), .Z(n4489) );
  XOR U1189 ( .A(n4461), .B(n4460), .Z(n4462) );
  NAND U1190 ( .A(n4111), .B(n4113), .Z(n128) );
  XOR U1191 ( .A(n4111), .B(n4113), .Z(n129) );
  NAND U1192 ( .A(n129), .B(n4112), .Z(n130) );
  NAND U1193 ( .A(n128), .B(n130), .Z(n4482) );
  XOR U1194 ( .A(n4301), .B(n4300), .Z(n4302) );
  NAND U1195 ( .A(n3860), .B(n3861), .Z(n131) );
  XOR U1196 ( .A(n3860), .B(n3861), .Z(n132) );
  NANDN U1197 ( .A(n3859), .B(n132), .Z(n133) );
  NAND U1198 ( .A(n131), .B(n133), .Z(n4457) );
  NAND U1199 ( .A(n4118), .B(n4119), .Z(n134) );
  XOR U1200 ( .A(n4118), .B(n4119), .Z(n135) );
  NAND U1201 ( .A(n135), .B(n4117), .Z(n136) );
  NAND U1202 ( .A(n134), .B(n136), .Z(n4453) );
  XNOR U1203 ( .A(n1469), .B(n1468), .Z(n1471) );
  XOR U1204 ( .A(n355), .B(n354), .Z(n2220) );
  XOR U1205 ( .A(n3464), .B(n3463), .Z(n3143) );
  NAND U1206 ( .A(n161), .B(n160), .Z(n137) );
  NANDN U1207 ( .A(n158), .B(n159), .Z(n138) );
  AND U1208 ( .A(n137), .B(n138), .Z(n2547) );
  XOR U1209 ( .A(n4016), .B(n4015), .Z(n4017) );
  XNOR U1210 ( .A(n4091), .B(n4090), .Z(n4093) );
  XOR U1211 ( .A(n4436), .B(n4435), .Z(n4515) );
  XOR U1212 ( .A(n4297), .B(n4296), .Z(n4508) );
  XOR U1213 ( .A(n4332), .B(n4331), .Z(n4334) );
  XOR U1214 ( .A(n4618), .B(oglobal[4]), .Z(n4619) );
  NAND U1215 ( .A(n4504), .B(n4505), .Z(n139) );
  XOR U1216 ( .A(n4504), .B(n4505), .Z(n140) );
  NANDN U1217 ( .A(n4503), .B(n140), .Z(n141) );
  NAND U1218 ( .A(n139), .B(n141), .Z(n4638) );
  NAND U1219 ( .A(n536), .B(n535), .Z(n142) );
  NANDN U1220 ( .A(n533), .B(n534), .Z(n143) );
  AND U1221 ( .A(n142), .B(n143), .Z(n3084) );
  NAND U1222 ( .A(n1381), .B(n1380), .Z(n144) );
  NANDN U1223 ( .A(n1382), .B(n1383), .Z(n145) );
  AND U1224 ( .A(n144), .B(n145), .Z(n3060) );
  XOR U1225 ( .A(n4766), .B(n4765), .Z(n4757) );
  NAND U1226 ( .A(n4644), .B(n4646), .Z(n146) );
  XOR U1227 ( .A(n4644), .B(n4646), .Z(n147) );
  NAND U1228 ( .A(n147), .B(n4645), .Z(n148) );
  NAND U1229 ( .A(n146), .B(n148), .Z(n4769) );
  XOR U1230 ( .A(n3986), .B(n3985), .Z(n3988) );
  XOR U1231 ( .A(n4571), .B(n4570), .Z(n4572) );
  XOR U1232 ( .A(n4753), .B(n4752), .Z(n4746) );
  XOR U1233 ( .A(n4800), .B(n4799), .Z(n4793) );
  XOR U1234 ( .A(n4386), .B(n4385), .Z(n4388) );
  XOR U1235 ( .A(n4549), .B(n4548), .Z(n4550) );
  XOR U1236 ( .A(n4559), .B(n4558), .Z(n4561) );
  NAND U1237 ( .A(n4082), .B(n4083), .Z(n149) );
  XOR U1238 ( .A(n4082), .B(n4083), .Z(n150) );
  NANDN U1239 ( .A(n4081), .B(n150), .Z(n151) );
  NAND U1240 ( .A(n149), .B(n151), .Z(n4555) );
  NAND U1241 ( .A(n4712), .B(n4713), .Z(n152) );
  XOR U1242 ( .A(n4712), .B(n4713), .Z(n153) );
  NANDN U1243 ( .A(n4711), .B(n153), .Z(n154) );
  NAND U1244 ( .A(n152), .B(n154), .Z(n4783) );
  NAND U1245 ( .A(n4833), .B(n4834), .Z(n155) );
  XOR U1246 ( .A(n4833), .B(n4834), .Z(n156) );
  NANDN U1247 ( .A(n4832), .B(n156), .Z(n157) );
  NAND U1248 ( .A(n155), .B(n157), .Z(n4840) );
  XOR U1249 ( .A(x[196]), .B(y[196]), .Z(n1675) );
  XOR U1250 ( .A(x[198]), .B(y[198]), .Z(n1672) );
  XNOR U1251 ( .A(x[206]), .B(y[206]), .Z(n1673) );
  XNOR U1252 ( .A(n1672), .B(n1673), .Z(n1674) );
  XOR U1253 ( .A(n1675), .B(n1674), .Z(n2141) );
  XOR U1254 ( .A(x[186]), .B(y[186]), .Z(n1166) );
  XOR U1255 ( .A(x[188]), .B(y[188]), .Z(n1163) );
  XNOR U1256 ( .A(x[192]), .B(y[192]), .Z(n1164) );
  XNOR U1257 ( .A(n1163), .B(n1164), .Z(n1165) );
  XOR U1258 ( .A(n1166), .B(n1165), .Z(n2139) );
  XOR U1259 ( .A(x[178]), .B(y[178]), .Z(n1154) );
  XOR U1260 ( .A(x[115]), .B(y[115]), .Z(n1151) );
  XNOR U1261 ( .A(x[180]), .B(y[180]), .Z(n1152) );
  XNOR U1262 ( .A(n1151), .B(n1152), .Z(n1153) );
  XNOR U1263 ( .A(n1154), .B(n1153), .Z(n2138) );
  XNOR U1264 ( .A(n2139), .B(n2138), .Z(n2140) );
  XNOR U1265 ( .A(n2141), .B(n2140), .Z(n2341) );
  XOR U1266 ( .A(x[162]), .B(y[162]), .Z(n1048) );
  XOR U1267 ( .A(x[164]), .B(y[164]), .Z(n1045) );
  XNOR U1268 ( .A(x[166]), .B(y[166]), .Z(n1046) );
  XNOR U1269 ( .A(n1045), .B(n1046), .Z(n1047) );
  XOR U1270 ( .A(n1048), .B(n1047), .Z(n2117) );
  XOR U1271 ( .A(x[150]), .B(y[150]), .Z(n183) );
  XOR U1272 ( .A(x[133]), .B(y[133]), .Z(n180) );
  XNOR U1273 ( .A(x[152]), .B(y[152]), .Z(n181) );
  XNOR U1274 ( .A(n180), .B(n181), .Z(n182) );
  XOR U1275 ( .A(n183), .B(n182), .Z(n2115) );
  XOR U1276 ( .A(x[134]), .B(y[134]), .Z(n201) );
  XOR U1277 ( .A(x[138]), .B(y[138]), .Z(n198) );
  XNOR U1278 ( .A(x[142]), .B(y[142]), .Z(n199) );
  XNOR U1279 ( .A(n198), .B(n199), .Z(n200) );
  XNOR U1280 ( .A(n201), .B(n200), .Z(n2114) );
  XNOR U1281 ( .A(n2115), .B(n2114), .Z(n2116) );
  XNOR U1282 ( .A(n2117), .B(n2116), .Z(n2340) );
  XOR U1283 ( .A(n2341), .B(n2340), .Z(n2343) );
  XOR U1284 ( .A(x[126]), .B(y[126]), .Z(n870) );
  XOR U1285 ( .A(x[128]), .B(y[128]), .Z(n867) );
  XNOR U1286 ( .A(x[151]), .B(y[151]), .Z(n868) );
  XNOR U1287 ( .A(n867), .B(n868), .Z(n869) );
  XOR U1288 ( .A(n870), .B(n869), .Z(n2535) );
  XOR U1289 ( .A(x[110]), .B(y[110]), .Z(n889) );
  XOR U1290 ( .A(x[112]), .B(y[112]), .Z(n886) );
  XNOR U1291 ( .A(x[114]), .B(y[114]), .Z(n887) );
  XNOR U1292 ( .A(n886), .B(n887), .Z(n888) );
  XOR U1293 ( .A(n889), .B(n888), .Z(n2533) );
  XOR U1294 ( .A(x[98]), .B(y[98]), .Z(n852) );
  XOR U1295 ( .A(x[102]), .B(y[102]), .Z(n849) );
  XNOR U1296 ( .A(x[169]), .B(y[169]), .Z(n850) );
  XNOR U1297 ( .A(n849), .B(n850), .Z(n851) );
  XNOR U1298 ( .A(n852), .B(n851), .Z(n2532) );
  XNOR U1299 ( .A(n2533), .B(n2532), .Z(n2534) );
  XNOR U1300 ( .A(n2535), .B(n2534), .Z(n2342) );
  XOR U1301 ( .A(n2343), .B(n2342), .Z(n1477) );
  XOR U1302 ( .A(x[42]), .B(y[42]), .Z(n2080) );
  XOR U1303 ( .A(x[44]), .B(y[44]), .Z(n2077) );
  XNOR U1304 ( .A(x[795]), .B(y[795]), .Z(n2078) );
  XNOR U1305 ( .A(n2077), .B(n2078), .Z(n2079) );
  XOR U1306 ( .A(n2080), .B(n2079), .Z(n472) );
  XOR U1307 ( .A(x[38]), .B(y[38]), .Z(n2086) );
  XOR U1308 ( .A(x[40]), .B(y[40]), .Z(n2083) );
  XNOR U1309 ( .A(x[403]), .B(y[403]), .Z(n2084) );
  XNOR U1310 ( .A(n2083), .B(n2084), .Z(n2085) );
  XOR U1311 ( .A(n2086), .B(n2085), .Z(n470) );
  XOR U1312 ( .A(x[34]), .B(y[34]), .Z(n2104) );
  XOR U1313 ( .A(x[36]), .B(y[36]), .Z(n2101) );
  XOR U1314 ( .A(x[793]), .B(y[793]), .Z(n2102) );
  XNOR U1315 ( .A(n2104), .B(n2103), .Z(n469) );
  XNOR U1316 ( .A(n470), .B(n469), .Z(n471) );
  XNOR U1317 ( .A(n472), .B(n471), .Z(n1558) );
  XOR U1318 ( .A(x[26]), .B(y[26]), .Z(n2098) );
  XOR U1319 ( .A(x[30]), .B(y[30]), .Z(n2095) );
  XOR U1320 ( .A(x[407]), .B(y[407]), .Z(n2096) );
  XOR U1321 ( .A(n2098), .B(n2097), .Z(n834) );
  XOR U1322 ( .A(x[22]), .B(y[22]), .Z(n2110) );
  XOR U1323 ( .A(x[24]), .B(y[24]), .Z(n2107) );
  XOR U1324 ( .A(x[791]), .B(y[791]), .Z(n2108) );
  XOR U1325 ( .A(n2110), .B(n2109), .Z(n832) );
  XOR U1326 ( .A(x[18]), .B(y[18]), .Z(n2074) );
  XOR U1327 ( .A(x[20]), .B(y[20]), .Z(n2071) );
  XOR U1328 ( .A(x[411]), .B(y[411]), .Z(n2072) );
  XNOR U1329 ( .A(n2074), .B(n2073), .Z(n831) );
  XNOR U1330 ( .A(n832), .B(n831), .Z(n833) );
  XOR U1331 ( .A(n834), .B(n833), .Z(n1559) );
  XNOR U1332 ( .A(n1558), .B(n1559), .Z(n1561) );
  XOR U1333 ( .A(x[84]), .B(y[84]), .Z(n736) );
  XOR U1334 ( .A(x[88]), .B(y[88]), .Z(n733) );
  XNOR U1335 ( .A(x[90]), .B(y[90]), .Z(n734) );
  XNOR U1336 ( .A(n733), .B(n734), .Z(n735) );
  XOR U1337 ( .A(n736), .B(n735), .Z(n448) );
  XOR U1338 ( .A(x[74]), .B(y[74]), .Z(n242) );
  XOR U1339 ( .A(x[76]), .B(y[76]), .Z(n239) );
  XNOR U1340 ( .A(x[187]), .B(y[187]), .Z(n240) );
  XNOR U1341 ( .A(n239), .B(n240), .Z(n241) );
  XOR U1342 ( .A(n242), .B(n241), .Z(n446) );
  XOR U1343 ( .A(x[58]), .B(y[58]), .Z(n940) );
  XOR U1344 ( .A(x[60]), .B(y[60]), .Z(n937) );
  XNOR U1345 ( .A(x[62]), .B(y[62]), .Z(n938) );
  XNOR U1346 ( .A(n937), .B(n938), .Z(n939) );
  XNOR U1347 ( .A(n940), .B(n939), .Z(n445) );
  XNOR U1348 ( .A(n446), .B(n445), .Z(n447) );
  XNOR U1349 ( .A(n448), .B(n447), .Z(n1560) );
  XOR U1350 ( .A(n1561), .B(n1560), .Z(n1475) );
  XOR U1351 ( .A(x[1]), .B(y[1]), .Z(n1813) );
  XOR U1352 ( .A(x[0]), .B(y[0]), .Z(n1810) );
  XOR U1353 ( .A(x[419]), .B(y[419]), .Z(n1811) );
  XOR U1354 ( .A(n1813), .B(n1812), .Z(n754) );
  XOR U1355 ( .A(x[9]), .B(y[9]), .Z(n1819) );
  XOR U1356 ( .A(x[5]), .B(y[5]), .Z(n1816) );
  XOR U1357 ( .A(x[785]), .B(y[785]), .Z(n1817) );
  XOR U1358 ( .A(n1819), .B(n1818), .Z(n752) );
  XOR U1359 ( .A(x[13]), .B(y[13]), .Z(n1807) );
  XOR U1360 ( .A(x[11]), .B(y[11]), .Z(n1804) );
  XOR U1361 ( .A(x[423]), .B(y[423]), .Z(n1805) );
  XNOR U1362 ( .A(n1807), .B(n1806), .Z(n751) );
  XNOR U1363 ( .A(n752), .B(n751), .Z(n753) );
  XNOR U1364 ( .A(n754), .B(n753), .Z(n1522) );
  XOR U1365 ( .A(x[17]), .B(y[17]), .Z(n1795) );
  XOR U1366 ( .A(x[15]), .B(y[15]), .Z(n1792) );
  XNOR U1367 ( .A(x[783]), .B(y[783]), .Z(n1793) );
  XNOR U1368 ( .A(n1792), .B(n1793), .Z(n1794) );
  XOR U1369 ( .A(n1795), .B(n1794), .Z(n1377) );
  XOR U1370 ( .A(x[23]), .B(y[23]), .Z(n1801) );
  XOR U1371 ( .A(x[19]), .B(y[19]), .Z(n1798) );
  XNOR U1372 ( .A(x[427]), .B(y[427]), .Z(n1799) );
  XNOR U1373 ( .A(n1798), .B(n1799), .Z(n1800) );
  XOR U1374 ( .A(n1801), .B(n1800), .Z(n1375) );
  XOR U1375 ( .A(x[29]), .B(y[29]), .Z(n1783) );
  XOR U1376 ( .A(x[27]), .B(y[27]), .Z(n1780) );
  XNOR U1377 ( .A(x[781]), .B(y[781]), .Z(n1781) );
  XNOR U1378 ( .A(n1780), .B(n1781), .Z(n1782) );
  XNOR U1379 ( .A(n1783), .B(n1782), .Z(n1374) );
  XNOR U1380 ( .A(n1375), .B(n1374), .Z(n1376) );
  XOR U1381 ( .A(n1377), .B(n1376), .Z(n1523) );
  XNOR U1382 ( .A(n1522), .B(n1523), .Z(n1525) );
  XOR U1383 ( .A(x[12]), .B(y[12]), .Z(n2062) );
  XOR U1384 ( .A(x[16]), .B(y[16]), .Z(n2059) );
  XOR U1385 ( .A(x[789]), .B(y[789]), .Z(n2060) );
  XOR U1386 ( .A(n2062), .B(n2061), .Z(n778) );
  XOR U1387 ( .A(x[6]), .B(y[6]), .Z(n2068) );
  XOR U1388 ( .A(x[8]), .B(y[8]), .Z(n2065) );
  XOR U1389 ( .A(x[415]), .B(y[415]), .Z(n2066) );
  XOR U1390 ( .A(n2068), .B(n2067), .Z(n776) );
  XOR U1391 ( .A(x[2]), .B(y[2]), .Z(n1825) );
  XOR U1392 ( .A(x[4]), .B(y[4]), .Z(n1822) );
  XOR U1393 ( .A(x[787]), .B(y[787]), .Z(n1823) );
  XNOR U1394 ( .A(n1825), .B(n1824), .Z(n775) );
  XNOR U1395 ( .A(n776), .B(n775), .Z(n777) );
  XNOR U1396 ( .A(n778), .B(n777), .Z(n1524) );
  XNOR U1397 ( .A(n1525), .B(n1524), .Z(n1474) );
  XNOR U1398 ( .A(n1475), .B(n1474), .Z(n1476) );
  XOR U1399 ( .A(n1477), .B(n1476), .Z(n1648) );
  XOR U1400 ( .A(x[189]), .B(y[189]), .Z(n1729) );
  XOR U1401 ( .A(x[185]), .B(y[185]), .Z(n1726) );
  XOR U1402 ( .A(x[491]), .B(y[491]), .Z(n1727) );
  XOR U1403 ( .A(n1729), .B(n1728), .Z(n1897) );
  XOR U1404 ( .A(x[193]), .B(y[193]), .Z(n1735) );
  XOR U1405 ( .A(x[191]), .B(y[191]), .Z(n1732) );
  XOR U1406 ( .A(x[749]), .B(y[749]), .Z(n1733) );
  XOR U1407 ( .A(n1735), .B(n1734), .Z(n1895) );
  XOR U1408 ( .A(x[197]), .B(y[197]), .Z(n1705) );
  XOR U1409 ( .A(x[195]), .B(y[195]), .Z(n1702) );
  XNOR U1410 ( .A(x[495]), .B(y[495]), .Z(n1703) );
  XNOR U1411 ( .A(n1702), .B(n1703), .Z(n1704) );
  XNOR U1412 ( .A(n1705), .B(n1704), .Z(n1894) );
  XNOR U1413 ( .A(n1895), .B(n1894), .Z(n1896) );
  XNOR U1414 ( .A(n1897), .B(n1896), .Z(n1553) );
  XOR U1415 ( .A(x[173]), .B(y[173]), .Z(n1873) );
  XOR U1416 ( .A(x[171]), .B(y[171]), .Z(n1870) );
  XNOR U1417 ( .A(x[753]), .B(y[753]), .Z(n1871) );
  XNOR U1418 ( .A(n1870), .B(n1871), .Z(n1872) );
  XOR U1419 ( .A(n1873), .B(n1872), .Z(n1717) );
  XOR U1420 ( .A(x[177]), .B(y[177]), .Z(n1879) );
  XOR U1421 ( .A(x[175]), .B(y[175]), .Z(n1876) );
  XNOR U1422 ( .A(x[487]), .B(y[487]), .Z(n1877) );
  XNOR U1423 ( .A(n1876), .B(n1877), .Z(n1878) );
  XOR U1424 ( .A(n1879), .B(n1878), .Z(n1715) );
  XOR U1425 ( .A(x[181]), .B(y[181]), .Z(n1741) );
  XOR U1426 ( .A(x[179]), .B(y[179]), .Z(n1738) );
  XNOR U1427 ( .A(x[751]), .B(y[751]), .Z(n1739) );
  XNOR U1428 ( .A(n1738), .B(n1739), .Z(n1740) );
  XNOR U1429 ( .A(n1741), .B(n1740), .Z(n1714) );
  XNOR U1430 ( .A(n1715), .B(n1714), .Z(n1716) );
  XNOR U1431 ( .A(n1717), .B(n1716), .Z(n1552) );
  XOR U1432 ( .A(n1553), .B(n1552), .Z(n1555) );
  XOR U1433 ( .A(x[203]), .B(y[203]), .Z(n1693) );
  XOR U1434 ( .A(x[199]), .B(y[199]), .Z(n1690) );
  XNOR U1435 ( .A(x[747]), .B(y[747]), .Z(n1691) );
  XNOR U1436 ( .A(n1690), .B(n1691), .Z(n1692) );
  XOR U1437 ( .A(n1693), .B(n1692), .Z(n1891) );
  XOR U1438 ( .A(x[207]), .B(y[207]), .Z(n1699) );
  XOR U1439 ( .A(x[205]), .B(y[205]), .Z(n1696) );
  XNOR U1440 ( .A(x[499]), .B(y[499]), .Z(n1697) );
  XNOR U1441 ( .A(n1696), .B(n1697), .Z(n1698) );
  XOR U1442 ( .A(n1699), .B(n1698), .Z(n1889) );
  XOR U1443 ( .A(x[211]), .B(y[211]), .Z(n1184) );
  XOR U1444 ( .A(x[209]), .B(y[209]), .Z(n1181) );
  XNOR U1445 ( .A(x[745]), .B(y[745]), .Z(n1182) );
  XNOR U1446 ( .A(n1181), .B(n1182), .Z(n1183) );
  XNOR U1447 ( .A(n1184), .B(n1183), .Z(n1888) );
  XNOR U1448 ( .A(n1889), .B(n1888), .Z(n1890) );
  XNOR U1449 ( .A(n1891), .B(n1890), .Z(n1554) );
  XOR U1450 ( .A(n1555), .B(n1554), .Z(n1531) );
  XOR U1451 ( .A(x[247]), .B(y[247]), .Z(n1225) );
  XOR U1452 ( .A(x[245]), .B(y[245]), .Z(n1223) );
  XNOR U1453 ( .A(x[519]), .B(y[519]), .Z(n1224) );
  XOR U1454 ( .A(n1223), .B(n1224), .Z(n1226) );
  XNOR U1455 ( .A(n1225), .B(n1226), .Z(n1720) );
  XOR U1456 ( .A(x[243]), .B(y[243]), .Z(n1346) );
  XOR U1457 ( .A(x[241]), .B(y[241]), .Z(n1344) );
  XNOR U1458 ( .A(x[737]), .B(y[737]), .Z(n1345) );
  XOR U1459 ( .A(n1344), .B(n1345), .Z(n1347) );
  XNOR U1460 ( .A(n1346), .B(n1347), .Z(n1721) );
  XOR U1461 ( .A(x[239]), .B(y[239]), .Z(n1340) );
  XOR U1462 ( .A(x[237]), .B(y[237]), .Z(n1338) );
  XNOR U1463 ( .A(x[515]), .B(y[515]), .Z(n1339) );
  XOR U1464 ( .A(n1338), .B(n1339), .Z(n1341) );
  XNOR U1465 ( .A(n1340), .B(n1341), .Z(n1722) );
  XOR U1466 ( .A(n1723), .B(n1722), .Z(n1411) );
  XOR U1467 ( .A(x[235]), .B(y[235]), .Z(n1352) );
  XOR U1468 ( .A(x[233]), .B(y[233]), .Z(n1350) );
  XNOR U1469 ( .A(x[739]), .B(y[739]), .Z(n1351) );
  XOR U1470 ( .A(n1350), .B(n1351), .Z(n1353) );
  XNOR U1471 ( .A(n1352), .B(n1353), .Z(n1937) );
  XOR U1472 ( .A(x[231]), .B(y[231]), .Z(n1268) );
  XOR U1473 ( .A(x[229]), .B(y[229]), .Z(n1266) );
  XNOR U1474 ( .A(x[511]), .B(y[511]), .Z(n1267) );
  XOR U1475 ( .A(n1266), .B(n1267), .Z(n1269) );
  XNOR U1476 ( .A(n1268), .B(n1269), .Z(n1938) );
  XOR U1477 ( .A(x[227]), .B(y[227]), .Z(n1262) );
  XOR U1478 ( .A(x[225]), .B(y[225]), .Z(n1260) );
  XNOR U1479 ( .A(x[741]), .B(y[741]), .Z(n1261) );
  XOR U1480 ( .A(n1260), .B(n1261), .Z(n1263) );
  XNOR U1481 ( .A(n1262), .B(n1263), .Z(n1939) );
  XOR U1482 ( .A(n1940), .B(n1939), .Z(n1409) );
  XOR U1483 ( .A(x[223]), .B(y[223]), .Z(n1274) );
  XOR U1484 ( .A(x[221]), .B(y[221]), .Z(n1272) );
  XNOR U1485 ( .A(x[507]), .B(y[507]), .Z(n1273) );
  XOR U1486 ( .A(n1272), .B(n1273), .Z(n1275) );
  XNOR U1487 ( .A(n1274), .B(n1275), .Z(n1931) );
  XOR U1488 ( .A(x[219]), .B(y[219]), .Z(n1177) );
  XOR U1489 ( .A(x[217]), .B(y[217]), .Z(n1175) );
  XNOR U1490 ( .A(x[743]), .B(y[743]), .Z(n1176) );
  XOR U1491 ( .A(n1175), .B(n1176), .Z(n1178) );
  XNOR U1492 ( .A(n1177), .B(n1178), .Z(n1932) );
  XOR U1493 ( .A(x[215]), .B(y[215]), .Z(n1171) );
  XOR U1494 ( .A(x[213]), .B(y[213]), .Z(n1169) );
  XNOR U1495 ( .A(x[503]), .B(y[503]), .Z(n1170) );
  XOR U1496 ( .A(n1169), .B(n1170), .Z(n1172) );
  XNOR U1497 ( .A(n1171), .B(n1172), .Z(n1933) );
  XNOR U1498 ( .A(n1934), .B(n1933), .Z(n1408) );
  XNOR U1499 ( .A(n1409), .B(n1408), .Z(n1410) );
  XNOR U1500 ( .A(n1411), .B(n1410), .Z(n1528) );
  XOR U1501 ( .A(x[291]), .B(y[291]), .Z(n1292) );
  XOR U1502 ( .A(x[287]), .B(y[287]), .Z(n1290) );
  XNOR U1503 ( .A(x[289]), .B(y[289]), .Z(n1291) );
  XOR U1504 ( .A(n1290), .B(n1291), .Z(n1293) );
  XNOR U1505 ( .A(n1292), .B(n1293), .Z(n1516) );
  XOR U1506 ( .A(x[285]), .B(y[285]), .Z(n1304) );
  XOR U1507 ( .A(x[281]), .B(y[281]), .Z(n1302) );
  XNOR U1508 ( .A(x[283]), .B(y[283]), .Z(n1303) );
  XOR U1509 ( .A(n1302), .B(n1303), .Z(n1305) );
  XNOR U1510 ( .A(n1304), .B(n1305), .Z(n1517) );
  XOR U1511 ( .A(x[279]), .B(y[279]), .Z(n1316) );
  XOR U1512 ( .A(x[275]), .B(y[275]), .Z(n1314) );
  XNOR U1513 ( .A(x[277]), .B(y[277]), .Z(n1315) );
  XOR U1514 ( .A(n1314), .B(n1315), .Z(n1317) );
  XNOR U1515 ( .A(n1316), .B(n1317), .Z(n1518) );
  XOR U1516 ( .A(n1519), .B(n1518), .Z(n1405) );
  XOR U1517 ( .A(x[259]), .B(y[259]), .Z(n1207) );
  XOR U1518 ( .A(x[257]), .B(y[257]), .Z(n1205) );
  XNOR U1519 ( .A(x[733]), .B(y[733]), .Z(n1206) );
  XOR U1520 ( .A(n1205), .B(n1206), .Z(n1208) );
  XNOR U1521 ( .A(n1207), .B(n1208), .Z(n1618) );
  XOR U1522 ( .A(x[255]), .B(y[255]), .Z(n1219) );
  XOR U1523 ( .A(x[253]), .B(y[253]), .Z(n1217) );
  XNOR U1524 ( .A(x[523]), .B(y[523]), .Z(n1218) );
  XOR U1525 ( .A(n1217), .B(n1218), .Z(n1220) );
  XNOR U1526 ( .A(n1219), .B(n1220), .Z(n1619) );
  XOR U1527 ( .A(x[251]), .B(y[251]), .Z(n1213) );
  XOR U1528 ( .A(x[249]), .B(y[249]), .Z(n1211) );
  XNOR U1529 ( .A(x[735]), .B(y[735]), .Z(n1212) );
  XOR U1530 ( .A(n1211), .B(n1212), .Z(n1214) );
  XNOR U1531 ( .A(n1213), .B(n1214), .Z(n1620) );
  XOR U1532 ( .A(n1621), .B(n1620), .Z(n1403) );
  XOR U1533 ( .A(x[273]), .B(y[273]), .Z(n1358) );
  XOR U1534 ( .A(x[269]), .B(y[269]), .Z(n1356) );
  XNOR U1535 ( .A(x[271]), .B(y[271]), .Z(n1357) );
  XOR U1536 ( .A(n1356), .B(n1357), .Z(n1359) );
  XNOR U1537 ( .A(n1358), .B(n1359), .Z(n1492) );
  XOR U1538 ( .A(x[267]), .B(y[267]), .Z(n1195) );
  XOR U1539 ( .A(x[265]), .B(y[265]), .Z(n1193) );
  XNOR U1540 ( .A(x[731]), .B(y[731]), .Z(n1194) );
  XOR U1541 ( .A(n1193), .B(n1194), .Z(n1196) );
  XNOR U1542 ( .A(n1195), .B(n1196), .Z(n1493) );
  XOR U1543 ( .A(x[263]), .B(y[263]), .Z(n1201) );
  XOR U1544 ( .A(x[261]), .B(y[261]), .Z(n1199) );
  XNOR U1545 ( .A(x[527]), .B(y[527]), .Z(n1200) );
  XOR U1546 ( .A(n1199), .B(n1200), .Z(n1202) );
  XNOR U1547 ( .A(n1201), .B(n1202), .Z(n1494) );
  XNOR U1548 ( .A(n1495), .B(n1494), .Z(n1402) );
  XNOR U1549 ( .A(n1403), .B(n1402), .Z(n1404) );
  XOR U1550 ( .A(n1405), .B(n1404), .Z(n1529) );
  XNOR U1551 ( .A(n1528), .B(n1529), .Z(n1530) );
  XOR U1552 ( .A(n1531), .B(n1530), .Z(n1649) );
  XOR U1553 ( .A(n1648), .B(n1649), .Z(n1651) );
  XOR U1554 ( .A(x[484]), .B(y[484]), .Z(n1615) );
  XOR U1555 ( .A(x[486]), .B(y[486]), .Z(n1612) );
  XNOR U1556 ( .A(x[488]), .B(y[488]), .Z(n1613) );
  XNOR U1557 ( .A(n1612), .B(n1613), .Z(n1614) );
  XOR U1558 ( .A(n1615), .B(n1614), .Z(n1012) );
  XOR U1559 ( .A(x[714]), .B(y[714]), .Z(n2367) );
  XOR U1560 ( .A(x[326]), .B(y[326]), .Z(n2364) );
  XOR U1561 ( .A(x[716]), .B(y[716]), .Z(n2365) );
  XOR U1562 ( .A(n2367), .B(n2366), .Z(n1010) );
  XOR U1563 ( .A(x[478]), .B(y[478]), .Z(n1609) );
  XOR U1564 ( .A(x[480]), .B(y[480]), .Z(n1606) );
  XNOR U1565 ( .A(x[482]), .B(y[482]), .Z(n1607) );
  XNOR U1566 ( .A(n1606), .B(n1607), .Z(n1608) );
  XNOR U1567 ( .A(n1609), .B(n1608), .Z(n1009) );
  XNOR U1568 ( .A(n1010), .B(n1009), .Z(n1011) );
  XNOR U1569 ( .A(n1012), .B(n1011), .Z(n538) );
  XOR U1570 ( .A(x[474]), .B(y[474]), .Z(n1597) );
  XOR U1571 ( .A(x[104]), .B(y[104]), .Z(n1594) );
  XOR U1572 ( .A(x[476]), .B(y[476]), .Z(n1595) );
  XOR U1573 ( .A(n1597), .B(n1596), .Z(n1024) );
  XOR U1574 ( .A(x[718]), .B(y[718]), .Z(n2349) );
  XOR U1575 ( .A(x[720]), .B(y[720]), .Z(n2346) );
  XNOR U1576 ( .A(x[722]), .B(y[722]), .Z(n2347) );
  XNOR U1577 ( .A(n2346), .B(n2347), .Z(n2348) );
  XOR U1578 ( .A(n2349), .B(n2348), .Z(n1022) );
  XOR U1579 ( .A(x[470]), .B(y[470]), .Z(n1591) );
  XOR U1580 ( .A(x[100]), .B(y[100]), .Z(n1588) );
  XOR U1581 ( .A(x[472]), .B(y[472]), .Z(n1589) );
  XNOR U1582 ( .A(n1591), .B(n1590), .Z(n1021) );
  XNOR U1583 ( .A(n1022), .B(n1021), .Z(n1023) );
  XNOR U1584 ( .A(n1024), .B(n1023), .Z(n537) );
  XOR U1585 ( .A(n538), .B(n537), .Z(n540) );
  XOR U1586 ( .A(x[464]), .B(y[464]), .Z(n1579) );
  XOR U1587 ( .A(x[466]), .B(y[466]), .Z(n1576) );
  XOR U1588 ( .A(x[468]), .B(y[468]), .Z(n1577) );
  XOR U1589 ( .A(n1579), .B(n1578), .Z(n1018) );
  XOR U1590 ( .A(x[724]), .B(y[724]), .Z(n1603) );
  XOR U1591 ( .A(x[726]), .B(y[726]), .Z(n1600) );
  XNOR U1592 ( .A(x[728]), .B(y[728]), .Z(n1601) );
  XNOR U1593 ( .A(n1600), .B(n1601), .Z(n1602) );
  XOR U1594 ( .A(n1603), .B(n1602), .Z(n1016) );
  XOR U1595 ( .A(x[458]), .B(y[458]), .Z(n1573) );
  XOR U1596 ( .A(x[460]), .B(y[460]), .Z(n1570) );
  XOR U1597 ( .A(x[462]), .B(y[462]), .Z(n1571) );
  XNOR U1598 ( .A(n1573), .B(n1572), .Z(n1015) );
  XNOR U1599 ( .A(n1016), .B(n1015), .Z(n1017) );
  XNOR U1600 ( .A(n1018), .B(n1017), .Z(n539) );
  XOR U1601 ( .A(n540), .B(n539), .Z(n265) );
  XOR U1602 ( .A(x[424]), .B(y[424]), .Z(n2227) );
  XOR U1603 ( .A(x[426]), .B(y[426]), .Z(n2224) );
  XNOR U1604 ( .A(x[428]), .B(y[428]), .Z(n2225) );
  XNOR U1605 ( .A(n2224), .B(n2225), .Z(n2226) );
  XOR U1606 ( .A(n2227), .B(n2226), .Z(n171) );
  XOR U1607 ( .A(x[418]), .B(y[418]), .Z(n2233) );
  XOR U1608 ( .A(x[420]), .B(y[420]), .Z(n2230) );
  XNOR U1609 ( .A(x[422]), .B(y[422]), .Z(n2231) );
  XNOR U1610 ( .A(n2230), .B(n2231), .Z(n2232) );
  XOR U1611 ( .A(n2233), .B(n2232), .Z(n169) );
  XOR U1612 ( .A(x[414]), .B(y[414]), .Z(n2487) );
  XOR U1613 ( .A(x[50]), .B(y[50]), .Z(n2484) );
  XOR U1614 ( .A(x[416]), .B(y[416]), .Z(n2485) );
  XNOR U1615 ( .A(n2487), .B(n2486), .Z(n168) );
  XNOR U1616 ( .A(n169), .B(n168), .Z(n170) );
  XNOR U1617 ( .A(n171), .B(n170), .Z(n2219) );
  XOR U1618 ( .A(x[410]), .B(y[410]), .Z(n2475) );
  XOR U1619 ( .A(x[46]), .B(y[46]), .Z(n2472) );
  XNOR U1620 ( .A(x[412]), .B(y[412]), .Z(n2473) );
  XNOR U1621 ( .A(n2472), .B(n2473), .Z(n2474) );
  XNOR U1622 ( .A(n2475), .B(n2474), .Z(n331) );
  XOR U1623 ( .A(x[404]), .B(y[404]), .Z(n2481) );
  XOR U1624 ( .A(x[406]), .B(y[406]), .Z(n2478) );
  XNOR U1625 ( .A(x[408]), .B(y[408]), .Z(n2479) );
  XNOR U1626 ( .A(n2478), .B(n2479), .Z(n2480) );
  XNOR U1627 ( .A(n2481), .B(n2480), .Z(n329) );
  XOR U1628 ( .A(x[398]), .B(y[398]), .Z(n2505) );
  XOR U1629 ( .A(x[400]), .B(y[400]), .Z(n2502) );
  XNOR U1630 ( .A(x[402]), .B(y[402]), .Z(n2503) );
  XNOR U1631 ( .A(n2502), .B(n2503), .Z(n2504) );
  XNOR U1632 ( .A(n2505), .B(n2504), .Z(n328) );
  XOR U1633 ( .A(n2219), .B(n2218), .Z(n2221) );
  XOR U1634 ( .A(x[392]), .B(y[392]), .Z(n2493) );
  XOR U1635 ( .A(x[32]), .B(y[32]), .Z(n2490) );
  XNOR U1636 ( .A(x[396]), .B(y[396]), .Z(n2491) );
  XNOR U1637 ( .A(n2490), .B(n2491), .Z(n2492) );
  XNOR U1638 ( .A(n2493), .B(n2492), .Z(n355) );
  XOR U1639 ( .A(x[388]), .B(y[388]), .Z(n2499) );
  XOR U1640 ( .A(x[28]), .B(y[28]), .Z(n2496) );
  XNOR U1641 ( .A(x[390]), .B(y[390]), .Z(n2497) );
  XNOR U1642 ( .A(n2496), .B(n2497), .Z(n2498) );
  XNOR U1643 ( .A(n2499), .B(n2498), .Z(n353) );
  XOR U1644 ( .A(x[382]), .B(y[382]), .Z(n2469) );
  XOR U1645 ( .A(x[384]), .B(y[384]), .Z(n2466) );
  XNOR U1646 ( .A(x[386]), .B(y[386]), .Z(n2467) );
  XNOR U1647 ( .A(n2466), .B(n2467), .Z(n2468) );
  XNOR U1648 ( .A(n2469), .B(n2468), .Z(n352) );
  XOR U1649 ( .A(n2221), .B(n2220), .Z(n264) );
  XOR U1650 ( .A(x[444]), .B(y[444]), .Z(n2263) );
  XOR U1651 ( .A(x[446]), .B(y[446]), .Z(n2260) );
  XOR U1652 ( .A(x[448]), .B(y[448]), .Z(n2261) );
  XOR U1653 ( .A(n2263), .B(n2262), .Z(n1006) );
  XOR U1654 ( .A(x[734]), .B(y[734]), .Z(n1567) );
  XOR U1655 ( .A(x[344]), .B(y[344]), .Z(n1564) );
  XOR U1656 ( .A(x[736]), .B(y[736]), .Z(n1565) );
  XOR U1657 ( .A(n1567), .B(n1566), .Z(n1004) );
  XOR U1658 ( .A(x[438]), .B(y[438]), .Z(n2275) );
  XOR U1659 ( .A(x[440]), .B(y[440]), .Z(n2272) );
  XOR U1660 ( .A(x[442]), .B(y[442]), .Z(n2273) );
  XNOR U1661 ( .A(n2275), .B(n2274), .Z(n1003) );
  XNOR U1662 ( .A(n1004), .B(n1003), .Z(n1005) );
  XNOR U1663 ( .A(n1006), .B(n1005), .Z(n658) );
  XOR U1664 ( .A(x[454]), .B(y[454]), .Z(n2257) );
  XOR U1665 ( .A(x[86]), .B(y[86]), .Z(n2254) );
  XOR U1666 ( .A(x[456]), .B(y[456]), .Z(n2255) );
  XOR U1667 ( .A(n2257), .B(n2256), .Z(n666) );
  XOR U1668 ( .A(x[730]), .B(y[730]), .Z(n1585) );
  XOR U1669 ( .A(x[340]), .B(y[340]), .Z(n1582) );
  XOR U1670 ( .A(x[732]), .B(y[732]), .Z(n1583) );
  XOR U1671 ( .A(n1585), .B(n1584), .Z(n664) );
  XOR U1672 ( .A(x[450]), .B(y[450]), .Z(n2251) );
  XOR U1673 ( .A(x[82]), .B(y[82]), .Z(n2248) );
  XOR U1674 ( .A(x[452]), .B(y[452]), .Z(n2249) );
  XNOR U1675 ( .A(n2251), .B(n2250), .Z(n663) );
  XNOR U1676 ( .A(n664), .B(n663), .Z(n665) );
  XNOR U1677 ( .A(n666), .B(n665), .Z(n657) );
  XOR U1678 ( .A(n658), .B(n657), .Z(n660) );
  XOR U1679 ( .A(x[434]), .B(y[434]), .Z(n2269) );
  XOR U1680 ( .A(x[68]), .B(y[68]), .Z(n2266) );
  XOR U1681 ( .A(x[436]), .B(y[436]), .Z(n2267) );
  XOR U1682 ( .A(n2269), .B(n2268), .Z(n1000) );
  XOR U1683 ( .A(x[738]), .B(y[738]), .Z(n2245) );
  XOR U1684 ( .A(x[740]), .B(y[740]), .Z(n2242) );
  XOR U1685 ( .A(x[742]), .B(y[742]), .Z(n2243) );
  XOR U1686 ( .A(n2245), .B(n2244), .Z(n998) );
  XOR U1687 ( .A(x[430]), .B(y[430]), .Z(n2239) );
  XOR U1688 ( .A(x[64]), .B(y[64]), .Z(n2236) );
  XNOR U1689 ( .A(x[432]), .B(y[432]), .Z(n2237) );
  XNOR U1690 ( .A(n2236), .B(n2237), .Z(n2238) );
  XNOR U1691 ( .A(n2239), .B(n2238), .Z(n997) );
  XNOR U1692 ( .A(n998), .B(n997), .Z(n999) );
  XNOR U1693 ( .A(n1000), .B(n999), .Z(n659) );
  XNOR U1694 ( .A(n660), .B(n659), .Z(n263) );
  XOR U1695 ( .A(n264), .B(n263), .Z(n266) );
  XOR U1696 ( .A(n265), .B(n266), .Z(n1453) );
  XOR U1697 ( .A(x[574]), .B(y[574]), .Z(n2012) );
  XOR U1698 ( .A(x[194]), .B(y[194]), .Z(n2009) );
  XNOR U1699 ( .A(x[576]), .B(y[576]), .Z(n2010) );
  XNOR U1700 ( .A(n2009), .B(n2010), .Z(n2011) );
  XOR U1701 ( .A(n2012), .B(n2011), .Z(n1771) );
  XOR U1702 ( .A(x[670]), .B(y[670]), .Z(n1849) );
  XOR U1703 ( .A(x[286]), .B(y[286]), .Z(n1846) );
  XNOR U1704 ( .A(x[672]), .B(y[672]), .Z(n1847) );
  XNOR U1705 ( .A(n1846), .B(n1847), .Z(n1848) );
  XOR U1706 ( .A(n1849), .B(n1848), .Z(n1769) );
  XOR U1707 ( .A(x[570]), .B(y[570]), .Z(n2196) );
  XOR U1708 ( .A(x[190]), .B(y[190]), .Z(n2193) );
  XNOR U1709 ( .A(x[572]), .B(y[572]), .Z(n2194) );
  XNOR U1710 ( .A(n2193), .B(n2194), .Z(n2195) );
  XNOR U1711 ( .A(n2196), .B(n2195), .Z(n1768) );
  XNOR U1712 ( .A(n1769), .B(n1768), .Z(n1770) );
  XNOR U1713 ( .A(n1771), .B(n1770), .Z(n694) );
  XOR U1714 ( .A(x[564]), .B(y[564]), .Z(n1970) );
  XOR U1715 ( .A(x[566]), .B(y[566]), .Z(n1967) );
  XNOR U1716 ( .A(x[568]), .B(y[568]), .Z(n1968) );
  XNOR U1717 ( .A(n1967), .B(n1968), .Z(n1969) );
  XOR U1718 ( .A(n1970), .B(n1969), .Z(n712) );
  XOR U1719 ( .A(x[674]), .B(y[674]), .Z(n1837) );
  XOR U1720 ( .A(x[290]), .B(y[290]), .Z(n1834) );
  XOR U1721 ( .A(x[676]), .B(y[676]), .Z(n1835) );
  XOR U1722 ( .A(n1837), .B(n1836), .Z(n710) );
  XOR U1723 ( .A(x[558]), .B(y[558]), .Z(n1843) );
  XOR U1724 ( .A(x[560]), .B(y[560]), .Z(n1840) );
  XOR U1725 ( .A(x[562]), .B(y[562]), .Z(n1841) );
  XNOR U1726 ( .A(n1843), .B(n1842), .Z(n709) );
  XNOR U1727 ( .A(n710), .B(n709), .Z(n711) );
  XOR U1728 ( .A(n712), .B(n711), .Z(n693) );
  XNOR U1729 ( .A(n694), .B(n693), .Z(n696) );
  XOR U1730 ( .A(x[554]), .B(y[554]), .Z(n1765) );
  XOR U1731 ( .A(x[176]), .B(y[176]), .Z(n1762) );
  XOR U1732 ( .A(x[556]), .B(y[556]), .Z(n1763) );
  XOR U1733 ( .A(n1765), .B(n1764), .Z(n1831) );
  XOR U1734 ( .A(x[678]), .B(y[678]), .Z(n1759) );
  XOR U1735 ( .A(x[680]), .B(y[680]), .Z(n1756) );
  XOR U1736 ( .A(x[682]), .B(y[682]), .Z(n1757) );
  XOR U1737 ( .A(n1759), .B(n1758), .Z(n1829) );
  XOR U1738 ( .A(x[550]), .B(y[550]), .Z(n1867) );
  XOR U1739 ( .A(x[172]), .B(y[172]), .Z(n1864) );
  XNOR U1740 ( .A(x[552]), .B(y[552]), .Z(n1865) );
  XNOR U1741 ( .A(n1864), .B(n1865), .Z(n1866) );
  XNOR U1742 ( .A(n1867), .B(n1866), .Z(n1828) );
  XNOR U1743 ( .A(n1829), .B(n1828), .Z(n1830) );
  XOR U1744 ( .A(n1831), .B(n1830), .Z(n695) );
  XNOR U1745 ( .A(n696), .B(n695), .Z(n1451) );
  XOR U1746 ( .A(x[624]), .B(y[624]), .Z(n2043) );
  XOR U1747 ( .A(x[626]), .B(y[626]), .Z(n2040) );
  XNOR U1748 ( .A(x[628]), .B(y[628]), .Z(n2041) );
  XNOR U1749 ( .A(n2040), .B(n2041), .Z(n2042) );
  XOR U1750 ( .A(n2043), .B(n2042), .Z(n177) );
  XOR U1751 ( .A(x[638]), .B(y[638]), .Z(n2202) );
  XOR U1752 ( .A(x[640]), .B(y[640]), .Z(n2199) );
  XNOR U1753 ( .A(x[642]), .B(y[642]), .Z(n2200) );
  XNOR U1754 ( .A(n2199), .B(n2200), .Z(n2201) );
  XOR U1755 ( .A(n2202), .B(n2201), .Z(n175) );
  XOR U1756 ( .A(x[634]), .B(y[634]), .Z(n2208) );
  XOR U1757 ( .A(x[254]), .B(y[254]), .Z(n2205) );
  XNOR U1758 ( .A(x[636]), .B(y[636]), .Z(n2206) );
  XNOR U1759 ( .A(n2205), .B(n2206), .Z(n2207) );
  XNOR U1760 ( .A(n2208), .B(n2207), .Z(n174) );
  XNOR U1761 ( .A(n175), .B(n174), .Z(n176) );
  XNOR U1762 ( .A(n177), .B(n176), .Z(n934) );
  XOR U1763 ( .A(x[594]), .B(y[594]), .Z(n1982) );
  XOR U1764 ( .A(x[218]), .B(y[218]), .Z(n1979) );
  XNOR U1765 ( .A(x[596]), .B(y[596]), .Z(n1980) );
  XNOR U1766 ( .A(n1979), .B(n1980), .Z(n1981) );
  XOR U1767 ( .A(n1982), .B(n1981), .Z(n2000) );
  XOR U1768 ( .A(x[658]), .B(y[658]), .Z(n1994) );
  XOR U1769 ( .A(x[660]), .B(y[660]), .Z(n1991) );
  XNOR U1770 ( .A(x[662]), .B(y[662]), .Z(n1992) );
  XNOR U1771 ( .A(n1991), .B(n1992), .Z(n1993) );
  XOR U1772 ( .A(n1994), .B(n1993), .Z(n1998) );
  XOR U1773 ( .A(x[590]), .B(y[590]), .Z(n2037) );
  XOR U1774 ( .A(x[214]), .B(y[214]), .Z(n2034) );
  XNOR U1775 ( .A(x[592]), .B(y[592]), .Z(n2035) );
  XNOR U1776 ( .A(n2034), .B(n2035), .Z(n2036) );
  XNOR U1777 ( .A(n2037), .B(n2036), .Z(n1997) );
  XNOR U1778 ( .A(n1998), .B(n1997), .Z(n1999) );
  XOR U1779 ( .A(n2000), .B(n1999), .Z(n933) );
  XNOR U1780 ( .A(n934), .B(n933), .Z(n936) );
  XOR U1781 ( .A(x[584]), .B(y[584]), .Z(n1964) );
  XOR U1782 ( .A(x[586]), .B(y[586]), .Z(n1961) );
  XNOR U1783 ( .A(x[588]), .B(y[588]), .Z(n1962) );
  XNOR U1784 ( .A(n1961), .B(n1962), .Z(n1963) );
  XOR U1785 ( .A(n1964), .B(n1963), .Z(n1747) );
  XOR U1786 ( .A(x[664]), .B(y[664]), .Z(n1988) );
  XOR U1787 ( .A(x[666]), .B(y[666]), .Z(n1985) );
  XNOR U1788 ( .A(x[668]), .B(y[668]), .Z(n1986) );
  XNOR U1789 ( .A(n1985), .B(n1986), .Z(n1987) );
  XOR U1790 ( .A(n1988), .B(n1987), .Z(n1745) );
  XOR U1791 ( .A(x[578]), .B(y[578]), .Z(n2178) );
  XOR U1792 ( .A(x[580]), .B(y[580]), .Z(n2175) );
  XNOR U1793 ( .A(x[582]), .B(y[582]), .Z(n2176) );
  XNOR U1794 ( .A(n2175), .B(n2176), .Z(n2177) );
  XNOR U1795 ( .A(n2178), .B(n2177), .Z(n1744) );
  XNOR U1796 ( .A(n1745), .B(n1744), .Z(n1746) );
  XOR U1797 ( .A(n1747), .B(n1746), .Z(n935) );
  XNOR U1798 ( .A(n936), .B(n935), .Z(n1450) );
  XOR U1799 ( .A(n1451), .B(n1450), .Z(n1452) );
  XNOR U1800 ( .A(n1453), .B(n1452), .Z(n1650) );
  XOR U1801 ( .A(n1651), .B(n1650), .Z(n1447) );
  XOR U1802 ( .A(x[320]), .B(y[320]), .Z(n2330) );
  XOR U1803 ( .A(x[324]), .B(y[324]), .Z(n2327) );
  XNOR U1804 ( .A(x[328]), .B(y[328]), .Z(n2328) );
  XNOR U1805 ( .A(n2327), .B(n2328), .Z(n2329) );
  XOR U1806 ( .A(n2330), .B(n2329), .Z(n307) );
  XOR U1807 ( .A(x[330]), .B(y[330]), .Z(n2324) );
  XOR U1808 ( .A(x[332]), .B(y[332]), .Z(n2321) );
  XNOR U1809 ( .A(x[334]), .B(y[334]), .Z(n2322) );
  XNOR U1810 ( .A(n2321), .B(n2322), .Z(n2323) );
  XNOR U1811 ( .A(n2324), .B(n2323), .Z(n306) );
  XNOR U1812 ( .A(n307), .B(n306), .Z(n309) );
  XOR U1813 ( .A(x[336]), .B(y[336]), .Z(n2336) );
  XOR U1814 ( .A(x[7]), .B(y[7]), .Z(n2333) );
  XNOR U1815 ( .A(x[338]), .B(y[338]), .Z(n2334) );
  XNOR U1816 ( .A(n2333), .B(n2334), .Z(n2335) );
  XOR U1817 ( .A(n2336), .B(n2335), .Z(n308) );
  XOR U1818 ( .A(n309), .B(n308), .Z(n2056) );
  XOR U1819 ( .A(x[372]), .B(y[372]), .Z(n2457) );
  XOR U1820 ( .A(x[374]), .B(y[374]), .Z(n2454) );
  XNOR U1821 ( .A(x[378]), .B(y[378]), .Z(n2455) );
  XNOR U1822 ( .A(n2454), .B(n2455), .Z(n2456) );
  XOR U1823 ( .A(n2457), .B(n2456), .Z(n976) );
  XOR U1824 ( .A(x[368]), .B(y[368]), .Z(n2463) );
  XOR U1825 ( .A(x[14]), .B(y[14]), .Z(n2460) );
  XNOR U1826 ( .A(x[370]), .B(y[370]), .Z(n2461) );
  XNOR U1827 ( .A(n2460), .B(n2461), .Z(n2462) );
  XOR U1828 ( .A(n2463), .B(n2462), .Z(n974) );
  XOR U1829 ( .A(x[364]), .B(y[364]), .Z(n1365) );
  XOR U1830 ( .A(x[10]), .B(y[10]), .Z(n1362) );
  XOR U1831 ( .A(x[366]), .B(y[366]), .Z(n1363) );
  XNOR U1832 ( .A(n1365), .B(n1364), .Z(n973) );
  XNOR U1833 ( .A(n974), .B(n973), .Z(n975) );
  XNOR U1834 ( .A(n976), .B(n975), .Z(n2053) );
  XOR U1835 ( .A(x[354]), .B(y[354]), .Z(n1329) );
  XOR U1836 ( .A(x[356]), .B(y[356]), .Z(n1326) );
  XOR U1837 ( .A(x[360]), .B(y[360]), .Z(n1327) );
  XOR U1838 ( .A(n1329), .B(n1328), .Z(n219) );
  XOR U1839 ( .A(x[348]), .B(y[348]), .Z(n1323) );
  XOR U1840 ( .A(x[350]), .B(y[350]), .Z(n1320) );
  XOR U1841 ( .A(x[352]), .B(y[352]), .Z(n1321) );
  XOR U1842 ( .A(n1323), .B(n1322), .Z(n217) );
  XOR U1843 ( .A(x[342]), .B(y[342]), .Z(n1371) );
  XOR U1844 ( .A(x[3]), .B(y[3]), .Z(n1368) );
  XOR U1845 ( .A(x[346]), .B(y[346]), .Z(n1369) );
  XNOR U1846 ( .A(n1371), .B(n1370), .Z(n216) );
  XNOR U1847 ( .A(n217), .B(n216), .Z(n218) );
  XOR U1848 ( .A(n219), .B(n218), .Z(n2054) );
  XNOR U1849 ( .A(n2053), .B(n2054), .Z(n2055) );
  XNOR U1850 ( .A(n2056), .B(n2055), .Z(n536) );
  XOR U1851 ( .A(x[260]), .B(y[260]), .Z(n402) );
  XOR U1852 ( .A(x[61]), .B(y[61]), .Z(n399) );
  XNOR U1853 ( .A(x[262]), .B(y[262]), .Z(n400) );
  XNOR U1854 ( .A(n399), .B(n400), .Z(n401) );
  XOR U1855 ( .A(n402), .B(n401), .Z(n2511) );
  XOR U1856 ( .A(x[252]), .B(y[252]), .Z(n430) );
  XOR U1857 ( .A(x[256]), .B(y[256]), .Z(n427) );
  XNOR U1858 ( .A(x[258]), .B(y[258]), .Z(n428) );
  XNOR U1859 ( .A(n427), .B(n428), .Z(n429) );
  XOR U1860 ( .A(n430), .B(n429), .Z(n2509) );
  XOR U1861 ( .A(x[244]), .B(y[244]), .Z(n383) );
  XOR U1862 ( .A(x[246]), .B(y[246]), .Z(n380) );
  XNOR U1863 ( .A(x[248]), .B(y[248]), .Z(n381) );
  XNOR U1864 ( .A(n380), .B(n381), .Z(n382) );
  XNOR U1865 ( .A(n383), .B(n382), .Z(n2508) );
  XNOR U1866 ( .A(n2509), .B(n2508), .Z(n2510) );
  XNOR U1867 ( .A(n2511), .B(n2510), .Z(n2539) );
  XOR U1868 ( .A(x[240]), .B(y[240]), .Z(n612) );
  XOR U1869 ( .A(x[75]), .B(y[75]), .Z(n609) );
  XNOR U1870 ( .A(x[242]), .B(y[242]), .Z(n610) );
  XNOR U1871 ( .A(n609), .B(n610), .Z(n611) );
  XOR U1872 ( .A(n612), .B(n611), .Z(n2147) );
  XOR U1873 ( .A(x[234]), .B(y[234]), .Z(n648) );
  XOR U1874 ( .A(x[79]), .B(y[79]), .Z(n645) );
  XOR U1875 ( .A(x[238]), .B(y[238]), .Z(n646) );
  XOR U1876 ( .A(n648), .B(n647), .Z(n2145) );
  XOR U1877 ( .A(x[226]), .B(y[226]), .Z(n642) );
  XOR U1878 ( .A(x[228]), .B(y[228]), .Z(n639) );
  XOR U1879 ( .A(x[230]), .B(y[230]), .Z(n640) );
  XNOR U1880 ( .A(n642), .B(n641), .Z(n2144) );
  XNOR U1881 ( .A(n2145), .B(n2144), .Z(n2146) );
  XNOR U1882 ( .A(n2147), .B(n2146), .Z(n2538) );
  XOR U1883 ( .A(n2539), .B(n2538), .Z(n2541) );
  XOR U1884 ( .A(x[220]), .B(y[220]), .Z(n590) );
  XOR U1885 ( .A(x[222]), .B(y[222]), .Z(n587) );
  XOR U1886 ( .A(x[224]), .B(y[224]), .Z(n588) );
  XOR U1887 ( .A(n590), .B(n589), .Z(n2172) );
  XOR U1888 ( .A(x[212]), .B(y[212]), .Z(n1669) );
  XOR U1889 ( .A(x[93]), .B(y[93]), .Z(n1666) );
  XNOR U1890 ( .A(x[216]), .B(y[216]), .Z(n1667) );
  XNOR U1891 ( .A(n1666), .B(n1667), .Z(n1668) );
  XOR U1892 ( .A(n1669), .B(n1668), .Z(n2170) );
  XOR U1893 ( .A(x[208]), .B(y[208]), .Z(n1142) );
  XOR U1894 ( .A(x[97]), .B(y[97]), .Z(n1139) );
  XNOR U1895 ( .A(x[210]), .B(y[210]), .Z(n1140) );
  XNOR U1896 ( .A(n1139), .B(n1140), .Z(n1141) );
  XNOR U1897 ( .A(n1142), .B(n1141), .Z(n2169) );
  XNOR U1898 ( .A(n2170), .B(n2169), .Z(n2171) );
  XNOR U1899 ( .A(n2172), .B(n2171), .Z(n2540) );
  XOR U1900 ( .A(n2541), .B(n2540), .Z(n534) );
  XOR U1901 ( .A(x[316]), .B(y[316]), .Z(n2318) );
  XOR U1902 ( .A(x[21]), .B(y[21]), .Z(n2315) );
  XOR U1903 ( .A(x[318]), .B(y[318]), .Z(n2316) );
  XOR U1904 ( .A(n2318), .B(n2317), .Z(n260) );
  XOR U1905 ( .A(x[312]), .B(y[312]), .Z(n2306) );
  XOR U1906 ( .A(x[25]), .B(y[25]), .Z(n2303) );
  XOR U1907 ( .A(x[314]), .B(y[314]), .Z(n2304) );
  XOR U1908 ( .A(n2306), .B(n2305), .Z(n258) );
  XOR U1909 ( .A(x[302]), .B(y[302]), .Z(n2312) );
  XOR U1910 ( .A(x[306]), .B(y[306]), .Z(n2309) );
  XOR U1911 ( .A(x[310]), .B(y[310]), .Z(n2310) );
  XNOR U1912 ( .A(n2312), .B(n2311), .Z(n257) );
  XNOR U1913 ( .A(n258), .B(n257), .Z(n259) );
  XNOR U1914 ( .A(n260), .B(n259), .Z(n2278) );
  XOR U1915 ( .A(x[296]), .B(y[296]), .Z(n2293) );
  XOR U1916 ( .A(x[298]), .B(y[298]), .Z(n2290) );
  XOR U1917 ( .A(x[300]), .B(y[300]), .Z(n2291) );
  XOR U1918 ( .A(n2293), .B(n2292), .Z(n272) );
  XOR U1919 ( .A(x[292]), .B(y[292]), .Z(n2287) );
  XOR U1920 ( .A(x[39]), .B(y[39]), .Z(n2284) );
  XOR U1921 ( .A(x[294]), .B(y[294]), .Z(n2285) );
  XOR U1922 ( .A(n2287), .B(n2286), .Z(n270) );
  XOR U1923 ( .A(x[284]), .B(y[284]), .Z(n500) );
  XOR U1924 ( .A(x[43]), .B(y[43]), .Z(n497) );
  XNOR U1925 ( .A(x[288]), .B(y[288]), .Z(n498) );
  XNOR U1926 ( .A(n497), .B(n498), .Z(n499) );
  XNOR U1927 ( .A(n500), .B(n499), .Z(n269) );
  XNOR U1928 ( .A(n270), .B(n269), .Z(n271) );
  XOR U1929 ( .A(n272), .B(n271), .Z(n2279) );
  XNOR U1930 ( .A(n2278), .B(n2279), .Z(n2280) );
  XOR U1931 ( .A(x[278]), .B(y[278]), .Z(n518) );
  XOR U1932 ( .A(x[280]), .B(y[280]), .Z(n515) );
  XNOR U1933 ( .A(x[282]), .B(y[282]), .Z(n516) );
  XNOR U1934 ( .A(n515), .B(n516), .Z(n517) );
  XOR U1935 ( .A(n518), .B(n517), .Z(n297) );
  XOR U1936 ( .A(x[270]), .B(y[270]), .Z(n408) );
  XOR U1937 ( .A(x[274]), .B(y[274]), .Z(n405) );
  XNOR U1938 ( .A(x[276]), .B(y[276]), .Z(n406) );
  XNOR U1939 ( .A(n405), .B(n406), .Z(n407) );
  XOR U1940 ( .A(n408), .B(n407), .Z(n295) );
  XOR U1941 ( .A(x[264]), .B(y[264]), .Z(n524) );
  XOR U1942 ( .A(x[57]), .B(y[57]), .Z(n521) );
  XNOR U1943 ( .A(x[266]), .B(y[266]), .Z(n522) );
  XNOR U1944 ( .A(n521), .B(n522), .Z(n523) );
  XNOR U1945 ( .A(n524), .B(n523), .Z(n294) );
  XNOR U1946 ( .A(n295), .B(n294), .Z(n296) );
  XOR U1947 ( .A(n297), .B(n296), .Z(n2281) );
  XOR U1948 ( .A(n2280), .B(n2281), .Z(n533) );
  XNOR U1949 ( .A(n534), .B(n533), .Z(n535) );
  XOR U1950 ( .A(n536), .B(n535), .Z(n1439) );
  XOR U1951 ( .A(x[534]), .B(y[534]), .Z(n2427) );
  XOR U1952 ( .A(x[158]), .B(y[158]), .Z(n2424) );
  XOR U1953 ( .A(x[536]), .B(y[536]), .Z(n2425) );
  XOR U1954 ( .A(n2427), .B(n2426), .Z(n678) );
  XOR U1955 ( .A(x[690]), .B(y[690]), .Z(n2451) );
  XOR U1956 ( .A(x[304]), .B(y[304]), .Z(n2448) );
  XOR U1957 ( .A(x[692]), .B(y[692]), .Z(n2449) );
  XOR U1958 ( .A(n2451), .B(n2450), .Z(n676) );
  XOR U1959 ( .A(x[530]), .B(y[530]), .Z(n2415) );
  XOR U1960 ( .A(x[154]), .B(y[154]), .Z(n2412) );
  XOR U1961 ( .A(x[532]), .B(y[532]), .Z(n2413) );
  XNOR U1962 ( .A(n2415), .B(n2414), .Z(n675) );
  XNOR U1963 ( .A(n676), .B(n675), .Z(n677) );
  XNOR U1964 ( .A(n678), .B(n677), .Z(n980) );
  XOR U1965 ( .A(x[524]), .B(y[524]), .Z(n2409) );
  XOR U1966 ( .A(x[526]), .B(y[526]), .Z(n2406) );
  XOR U1967 ( .A(x[528]), .B(y[528]), .Z(n2407) );
  XOR U1968 ( .A(n2409), .B(n2408), .Z(n690) );
  XOR U1969 ( .A(x[694]), .B(y[694]), .Z(n2439) );
  XOR U1970 ( .A(x[308]), .B(y[308]), .Z(n2436) );
  XOR U1971 ( .A(x[696]), .B(y[696]), .Z(n2437) );
  XOR U1972 ( .A(n2439), .B(n2438), .Z(n688) );
  XOR U1973 ( .A(x[518]), .B(y[518]), .Z(n2397) );
  XOR U1974 ( .A(x[520]), .B(y[520]), .Z(n2394) );
  XOR U1975 ( .A(x[522]), .B(y[522]), .Z(n2395) );
  XNOR U1976 ( .A(n2397), .B(n2396), .Z(n687) );
  XNOR U1977 ( .A(n688), .B(n687), .Z(n689) );
  XNOR U1978 ( .A(n690), .B(n689), .Z(n979) );
  XOR U1979 ( .A(n980), .B(n979), .Z(n982) );
  XOR U1980 ( .A(x[544]), .B(y[544]), .Z(n2445) );
  XOR U1981 ( .A(x[546]), .B(y[546]), .Z(n2442) );
  XOR U1982 ( .A(x[548]), .B(y[548]), .Z(n2443) );
  XOR U1983 ( .A(n2445), .B(n2444), .Z(n700) );
  XOR U1984 ( .A(x[684]), .B(y[684]), .Z(n1861) );
  XOR U1985 ( .A(x[686]), .B(y[686]), .Z(n1858) );
  XNOR U1986 ( .A(x[688]), .B(y[688]), .Z(n1859) );
  XNOR U1987 ( .A(n1858), .B(n1859), .Z(n1860) );
  XOR U1988 ( .A(n1861), .B(n1860), .Z(n698) );
  XOR U1989 ( .A(x[538]), .B(y[538]), .Z(n2433) );
  XOR U1990 ( .A(x[540]), .B(y[540]), .Z(n2430) );
  XOR U1991 ( .A(x[542]), .B(y[542]), .Z(n2431) );
  XNOR U1992 ( .A(n2433), .B(n2432), .Z(n697) );
  XNOR U1993 ( .A(n698), .B(n697), .Z(n699) );
  XNOR U1994 ( .A(n700), .B(n699), .Z(n981) );
  XOR U1995 ( .A(n982), .B(n981), .Z(n161) );
  XOR U1996 ( .A(x[498]), .B(y[498]), .Z(n2373) );
  XOR U1997 ( .A(x[500]), .B(y[500]), .Z(n2370) );
  XOR U1998 ( .A(x[502]), .B(y[502]), .Z(n2371) );
  XOR U1999 ( .A(n2373), .B(n2372), .Z(n704) );
  XOR U2000 ( .A(x[704]), .B(y[704]), .Z(n2403) );
  XOR U2001 ( .A(x[706]), .B(y[706]), .Z(n2400) );
  XOR U2002 ( .A(x[708]), .B(y[708]), .Z(n2401) );
  XOR U2003 ( .A(n2403), .B(n2402), .Z(n703) );
  XOR U2004 ( .A(n704), .B(n703), .Z(n706) );
  XOR U2005 ( .A(x[504]), .B(y[504]), .Z(n2379) );
  XOR U2006 ( .A(x[506]), .B(y[506]), .Z(n2376) );
  XOR U2007 ( .A(x[508]), .B(y[508]), .Z(n2377) );
  XOR U2008 ( .A(n2379), .B(n2378), .Z(n705) );
  XOR U2009 ( .A(n706), .B(n705), .Z(n838) );
  XOR U2010 ( .A(x[514]), .B(y[514]), .Z(n2391) );
  XOR U2011 ( .A(x[140]), .B(y[140]), .Z(n2388) );
  XOR U2012 ( .A(x[516]), .B(y[516]), .Z(n2389) );
  XOR U2013 ( .A(n2391), .B(n2390), .Z(n672) );
  XOR U2014 ( .A(x[698]), .B(y[698]), .Z(n2421) );
  XOR U2015 ( .A(x[700]), .B(y[700]), .Z(n2418) );
  XOR U2016 ( .A(x[702]), .B(y[702]), .Z(n2419) );
  XOR U2017 ( .A(n2421), .B(n2420), .Z(n670) );
  XOR U2018 ( .A(x[510]), .B(y[510]), .Z(n371) );
  XOR U2019 ( .A(x[136]), .B(y[136]), .Z(n368) );
  XOR U2020 ( .A(x[512]), .B(y[512]), .Z(n369) );
  XNOR U2021 ( .A(n371), .B(n370), .Z(n669) );
  XNOR U2022 ( .A(n670), .B(n669), .Z(n671) );
  XNOR U2023 ( .A(n672), .B(n671), .Z(n837) );
  XNOR U2024 ( .A(n838), .B(n837), .Z(n840) );
  XOR U2025 ( .A(x[494]), .B(y[494]), .Z(n2361) );
  XOR U2026 ( .A(x[122]), .B(y[122]), .Z(n2358) );
  XOR U2027 ( .A(x[496]), .B(y[496]), .Z(n2359) );
  XOR U2028 ( .A(n2361), .B(n2360), .Z(n684) );
  XOR U2029 ( .A(x[710]), .B(y[710]), .Z(n2385) );
  XOR U2030 ( .A(x[322]), .B(y[322]), .Z(n2382) );
  XOR U2031 ( .A(x[712]), .B(y[712]), .Z(n2383) );
  XOR U2032 ( .A(n2385), .B(n2384), .Z(n682) );
  XOR U2033 ( .A(x[490]), .B(y[490]), .Z(n2355) );
  XOR U2034 ( .A(x[118]), .B(y[118]), .Z(n2352) );
  XOR U2035 ( .A(x[492]), .B(y[492]), .Z(n2353) );
  XNOR U2036 ( .A(n2355), .B(n2354), .Z(n681) );
  XNOR U2037 ( .A(n682), .B(n681), .Z(n683) );
  XNOR U2038 ( .A(n684), .B(n683), .Z(n839) );
  XOR U2039 ( .A(n840), .B(n839), .Z(n159) );
  XOR U2040 ( .A(x[614]), .B(y[614]), .Z(n1855) );
  XOR U2041 ( .A(x[236]), .B(y[236]), .Z(n1852) );
  XNOR U2042 ( .A(x[616]), .B(y[616]), .Z(n1853) );
  XNOR U2043 ( .A(n1852), .B(n1853), .Z(n1854) );
  XOR U2044 ( .A(n1855), .B(n1854), .Z(n994) );
  XOR U2045 ( .A(x[630]), .B(y[630]), .Z(n2184) );
  XOR U2046 ( .A(x[250]), .B(y[250]), .Z(n2181) );
  XNOR U2047 ( .A(x[632]), .B(y[632]), .Z(n2182) );
  XNOR U2048 ( .A(n2181), .B(n2182), .Z(n2183) );
  XOR U2049 ( .A(n2184), .B(n2183), .Z(n992) );
  XOR U2050 ( .A(x[610]), .B(y[610]), .Z(n1753) );
  XOR U2051 ( .A(x[232]), .B(y[232]), .Z(n1750) );
  XOR U2052 ( .A(x[612]), .B(y[612]), .Z(n1751) );
  XNOR U2053 ( .A(n1753), .B(n1752), .Z(n991) );
  XNOR U2054 ( .A(n992), .B(n991), .Z(n993) );
  XNOR U2055 ( .A(n994), .B(n993), .Z(n2004) );
  XOR U2056 ( .A(x[618]), .B(y[618]), .Z(n2214) );
  XOR U2057 ( .A(x[620]), .B(y[620]), .Z(n2211) );
  XNOR U2058 ( .A(x[622]), .B(y[622]), .Z(n2212) );
  XNOR U2059 ( .A(n2211), .B(n2212), .Z(n2213) );
  XOR U2060 ( .A(n2214), .B(n2213), .Z(n165) );
  XOR U2061 ( .A(x[650]), .B(y[650]), .Z(n2024) );
  XOR U2062 ( .A(x[268]), .B(y[268]), .Z(n2021) );
  XNOR U2063 ( .A(x[652]), .B(y[652]), .Z(n2022) );
  XNOR U2064 ( .A(n2021), .B(n2022), .Z(n2023) );
  XOR U2065 ( .A(n2024), .B(n2023), .Z(n163) );
  XOR U2066 ( .A(x[644]), .B(y[644]), .Z(n2018) );
  XOR U2067 ( .A(x[646]), .B(y[646]), .Z(n2015) );
  XNOR U2068 ( .A(x[648]), .B(y[648]), .Z(n2016) );
  XNOR U2069 ( .A(n2015), .B(n2016), .Z(n2017) );
  XNOR U2070 ( .A(n2018), .B(n2017), .Z(n162) );
  XNOR U2071 ( .A(n163), .B(n162), .Z(n164) );
  XNOR U2072 ( .A(n165), .B(n164), .Z(n2003) );
  XOR U2073 ( .A(n2004), .B(n2003), .Z(n2006) );
  XOR U2074 ( .A(x[604]), .B(y[604]), .Z(n2190) );
  XOR U2075 ( .A(x[606]), .B(y[606]), .Z(n2187) );
  XNOR U2076 ( .A(x[608]), .B(y[608]), .Z(n2188) );
  XNOR U2077 ( .A(n2187), .B(n2188), .Z(n2189) );
  XOR U2078 ( .A(n2190), .B(n2189), .Z(n2031) );
  XOR U2079 ( .A(x[654]), .B(y[654]), .Z(n1976) );
  XOR U2080 ( .A(x[272]), .B(y[272]), .Z(n1973) );
  XOR U2081 ( .A(x[656]), .B(y[656]), .Z(n1974) );
  XOR U2082 ( .A(n1976), .B(n1975), .Z(n2029) );
  XOR U2083 ( .A(x[598]), .B(y[598]), .Z(n2049) );
  XOR U2084 ( .A(x[600]), .B(y[600]), .Z(n2046) );
  XNOR U2085 ( .A(x[602]), .B(y[602]), .Z(n2047) );
  XNOR U2086 ( .A(n2046), .B(n2047), .Z(n2048) );
  XNOR U2087 ( .A(n2049), .B(n2048), .Z(n2028) );
  XNOR U2088 ( .A(n2029), .B(n2028), .Z(n2030) );
  XNOR U2089 ( .A(n2031), .B(n2030), .Z(n2005) );
  XNOR U2090 ( .A(n2006), .B(n2005), .Z(n158) );
  XNOR U2091 ( .A(n159), .B(n158), .Z(n160) );
  XNOR U2092 ( .A(n161), .B(n160), .Z(n1438) );
  XNOR U2093 ( .A(n1439), .B(n1438), .Z(n1441) );
  XOR U2094 ( .A(x[33]), .B(y[33]), .Z(n1777) );
  XOR U2095 ( .A(x[31]), .B(y[31]), .Z(n1774) );
  XOR U2096 ( .A(x[431]), .B(y[431]), .Z(n1775) );
  XOR U2097 ( .A(n1777), .B(n1776), .Z(n926) );
  XOR U2098 ( .A(x[37]), .B(y[37]), .Z(n1789) );
  XOR U2099 ( .A(x[35]), .B(y[35]), .Z(n1786) );
  XOR U2100 ( .A(x[779]), .B(y[779]), .Z(n1787) );
  XOR U2101 ( .A(n1789), .B(n1788), .Z(n924) );
  XOR U2102 ( .A(x[45]), .B(y[45]), .Z(n1244) );
  XOR U2103 ( .A(x[41]), .B(y[41]), .Z(n1241) );
  XOR U2104 ( .A(x[435]), .B(y[435]), .Z(n1242) );
  XNOR U2105 ( .A(n1244), .B(n1243), .Z(n923) );
  XNOR U2106 ( .A(n924), .B(n923), .Z(n925) );
  XNOR U2107 ( .A(n926), .B(n925), .Z(n1462) );
  XOR U2108 ( .A(x[49]), .B(y[49]), .Z(n1238) );
  XOR U2109 ( .A(x[47]), .B(y[47]), .Z(n1235) );
  XNOR U2110 ( .A(x[777]), .B(y[777]), .Z(n1236) );
  XNOR U2111 ( .A(n1235), .B(n1236), .Z(n1237) );
  XOR U2112 ( .A(n1238), .B(n1237), .Z(n1311) );
  XOR U2113 ( .A(x[53]), .B(y[53]), .Z(n1250) );
  XOR U2114 ( .A(x[51]), .B(y[51]), .Z(n1247) );
  XNOR U2115 ( .A(x[439]), .B(y[439]), .Z(n1248) );
  XNOR U2116 ( .A(n1247), .B(n1248), .Z(n1249) );
  XOR U2117 ( .A(n1250), .B(n1249), .Z(n1309) );
  XOR U2118 ( .A(x[59]), .B(y[59]), .Z(n2159) );
  XOR U2119 ( .A(x[55]), .B(y[55]), .Z(n2156) );
  XNOR U2120 ( .A(x[775]), .B(y[775]), .Z(n2157) );
  XNOR U2121 ( .A(n2156), .B(n2157), .Z(n2158) );
  XNOR U2122 ( .A(n2159), .B(n2158), .Z(n1308) );
  XNOR U2123 ( .A(n1309), .B(n1308), .Z(n1310) );
  XOR U2124 ( .A(n1311), .B(n1310), .Z(n1463) );
  XNOR U2125 ( .A(n1462), .B(n1463), .Z(n1465) );
  XOR U2126 ( .A(x[65]), .B(y[65]), .Z(n2165) );
  XOR U2127 ( .A(x[63]), .B(y[63]), .Z(n2162) );
  XOR U2128 ( .A(x[443]), .B(y[443]), .Z(n2163) );
  XOR U2129 ( .A(n2165), .B(n2164), .Z(n846) );
  XOR U2130 ( .A(x[69]), .B(y[69]), .Z(n2153) );
  XOR U2131 ( .A(x[67]), .B(y[67]), .Z(n2150) );
  XOR U2132 ( .A(x[773]), .B(y[773]), .Z(n2151) );
  XOR U2133 ( .A(n2153), .B(n2152), .Z(n844) );
  XOR U2134 ( .A(x[73]), .B(y[73]), .Z(n2135) );
  XOR U2135 ( .A(x[71]), .B(y[71]), .Z(n2132) );
  XNOR U2136 ( .A(x[447]), .B(y[447]), .Z(n2133) );
  XNOR U2137 ( .A(n2132), .B(n2133), .Z(n2134) );
  XNOR U2138 ( .A(n2135), .B(n2134), .Z(n843) );
  XNOR U2139 ( .A(n844), .B(n843), .Z(n845) );
  XNOR U2140 ( .A(n846), .B(n845), .Z(n1464) );
  XOR U2141 ( .A(n1465), .B(n1464), .Z(n1417) );
  XOR U2142 ( .A(x[81]), .B(y[81]), .Z(n2123) );
  XOR U2143 ( .A(x[77]), .B(y[77]), .Z(n2120) );
  XOR U2144 ( .A(x[771]), .B(y[771]), .Z(n2121) );
  XOR U2145 ( .A(n2123), .B(n2122), .Z(n1066) );
  XOR U2146 ( .A(x[85]), .B(y[85]), .Z(n2129) );
  XOR U2147 ( .A(x[83]), .B(y[83]), .Z(n2126) );
  XOR U2148 ( .A(x[451]), .B(y[451]), .Z(n2127) );
  XOR U2149 ( .A(n2129), .B(n2128), .Z(n1064) );
  XOR U2150 ( .A(x[89]), .B(y[89]), .Z(n2529) );
  XOR U2151 ( .A(x[87]), .B(y[87]), .Z(n2526) );
  XOR U2152 ( .A(x[769]), .B(y[769]), .Z(n2527) );
  XNOR U2153 ( .A(n2529), .B(n2528), .Z(n1063) );
  XNOR U2154 ( .A(n1064), .B(n1063), .Z(n1065) );
  XNOR U2155 ( .A(n1066), .B(n1065), .Z(n1432) );
  XOR U2156 ( .A(x[95]), .B(y[95]), .Z(n2517) );
  XOR U2157 ( .A(x[91]), .B(y[91]), .Z(n2514) );
  XNOR U2158 ( .A(x[455]), .B(y[455]), .Z(n2515) );
  XNOR U2159 ( .A(n2514), .B(n2515), .Z(n2516) );
  XOR U2160 ( .A(n2517), .B(n2516), .Z(n1335) );
  XOR U2161 ( .A(x[101]), .B(y[101]), .Z(n2523) );
  XOR U2162 ( .A(x[99]), .B(y[99]), .Z(n2520) );
  XNOR U2163 ( .A(x[767]), .B(y[767]), .Z(n2521) );
  XNOR U2164 ( .A(n2520), .B(n2521), .Z(n2522) );
  XOR U2165 ( .A(n2523), .B(n2522), .Z(n1333) );
  XOR U2166 ( .A(x[105]), .B(y[105]), .Z(n1639) );
  XOR U2167 ( .A(x[103]), .B(y[103]), .Z(n1636) );
  XNOR U2168 ( .A(x[459]), .B(y[459]), .Z(n1637) );
  XNOR U2169 ( .A(n1636), .B(n1637), .Z(n1638) );
  XNOR U2170 ( .A(n1639), .B(n1638), .Z(n1332) );
  XNOR U2171 ( .A(n1333), .B(n1332), .Z(n1334) );
  XOR U2172 ( .A(n1335), .B(n1334), .Z(n1433) );
  XNOR U2173 ( .A(n1432), .B(n1433), .Z(n1435) );
  XOR U2174 ( .A(x[109]), .B(y[109]), .Z(n1627) );
  XOR U2175 ( .A(x[107]), .B(y[107]), .Z(n1624) );
  XNOR U2176 ( .A(x[765]), .B(y[765]), .Z(n1625) );
  XNOR U2177 ( .A(n1624), .B(n1625), .Z(n1626) );
  XOR U2178 ( .A(n1627), .B(n1626), .Z(n1281) );
  XOR U2179 ( .A(x[117]), .B(y[117]), .Z(n1633) );
  XOR U2180 ( .A(x[113]), .B(y[113]), .Z(n1630) );
  XNOR U2181 ( .A(x[463]), .B(y[463]), .Z(n1631) );
  XNOR U2182 ( .A(n1630), .B(n1631), .Z(n1632) );
  XOR U2183 ( .A(n1633), .B(n1632), .Z(n1279) );
  XOR U2184 ( .A(x[121]), .B(y[121]), .Z(n1513) );
  XOR U2185 ( .A(x[119]), .B(y[119]), .Z(n1510) );
  XNOR U2186 ( .A(x[763]), .B(y[763]), .Z(n1511) );
  XNOR U2187 ( .A(n1510), .B(n1511), .Z(n1512) );
  XNOR U2188 ( .A(n1513), .B(n1512), .Z(n1278) );
  XNOR U2189 ( .A(n1279), .B(n1278), .Z(n1280) );
  XNOR U2190 ( .A(n1281), .B(n1280), .Z(n1434) );
  XOR U2191 ( .A(n1435), .B(n1434), .Z(n1415) );
  XOR U2192 ( .A(x[167]), .B(y[167]), .Z(n1885) );
  XOR U2193 ( .A(x[163]), .B(y[163]), .Z(n1882) );
  XOR U2194 ( .A(x[483]), .B(y[483]), .Z(n1883) );
  XOR U2195 ( .A(n1885), .B(n1884), .Z(n1088) );
  XOR U2196 ( .A(x[161]), .B(y[161]), .Z(n1952) );
  XOR U2197 ( .A(x[159]), .B(y[159]), .Z(n1949) );
  XOR U2198 ( .A(x[755]), .B(y[755]), .Z(n1950) );
  XNOR U2199 ( .A(n1952), .B(n1951), .Z(n1087) );
  XNOR U2200 ( .A(n1088), .B(n1087), .Z(n1090) );
  XOR U2201 ( .A(x[157]), .B(y[157]), .Z(n1946) );
  XOR U2202 ( .A(x[155]), .B(y[155]), .Z(n1943) );
  XOR U2203 ( .A(x[479]), .B(y[479]), .Z(n1944) );
  XOR U2204 ( .A(n1946), .B(n1945), .Z(n1089) );
  XOR U2205 ( .A(n1090), .B(n1089), .Z(n1398) );
  XOR U2206 ( .A(x[153]), .B(y[153]), .Z(n1958) );
  XOR U2207 ( .A(x[149]), .B(y[149]), .Z(n1955) );
  XOR U2208 ( .A(x[757]), .B(y[757]), .Z(n1956) );
  XOR U2209 ( .A(n1958), .B(n1957), .Z(n1685) );
  XOR U2210 ( .A(x[145]), .B(y[145]), .Z(n1916) );
  XOR U2211 ( .A(x[143]), .B(y[143]), .Z(n1913) );
  XOR U2212 ( .A(x[475]), .B(y[475]), .Z(n1914) );
  XOR U2213 ( .A(n1916), .B(n1915), .Z(n1684) );
  XOR U2214 ( .A(n1685), .B(n1684), .Z(n1687) );
  XOR U2215 ( .A(x[141]), .B(y[141]), .Z(n1910) );
  XOR U2216 ( .A(x[139]), .B(y[139]), .Z(n1907) );
  XOR U2217 ( .A(x[759]), .B(y[759]), .Z(n1908) );
  XOR U2218 ( .A(n1910), .B(n1909), .Z(n1686) );
  XOR U2219 ( .A(n1687), .B(n1686), .Z(n1397) );
  XOR U2220 ( .A(x[137]), .B(y[137]), .Z(n1922) );
  XOR U2221 ( .A(x[135]), .B(y[135]), .Z(n1919) );
  XOR U2222 ( .A(x[471]), .B(y[471]), .Z(n1920) );
  XOR U2223 ( .A(n1922), .B(n1921), .Z(n1284) );
  XOR U2224 ( .A(x[131]), .B(y[131]), .Z(n1507) );
  XOR U2225 ( .A(x[127]), .B(y[127]), .Z(n1504) );
  XOR U2226 ( .A(x[761]), .B(y[761]), .Z(n1505) );
  XOR U2227 ( .A(n1507), .B(n1506), .Z(n1285) );
  XOR U2228 ( .A(n1284), .B(n1285), .Z(n1287) );
  XOR U2229 ( .A(x[125]), .B(y[125]), .Z(n1501) );
  XOR U2230 ( .A(x[123]), .B(y[123]), .Z(n1498) );
  XOR U2231 ( .A(x[467]), .B(y[467]), .Z(n1499) );
  XOR U2232 ( .A(n1501), .B(n1500), .Z(n1286) );
  XNOR U2233 ( .A(n1287), .B(n1286), .Z(n1396) );
  XOR U2234 ( .A(n1397), .B(n1396), .Z(n1399) );
  XNOR U2235 ( .A(n1398), .B(n1399), .Z(n1414) );
  XNOR U2236 ( .A(n1415), .B(n1414), .Z(n1416) );
  XNOR U2237 ( .A(n1417), .B(n1416), .Z(n1440) );
  XOR U2238 ( .A(n1441), .B(n1440), .Z(n1445) );
  XOR U2239 ( .A(x[297]), .B(y[297]), .Z(n1299) );
  XOR U2240 ( .A(x[293]), .B(y[293]), .Z(n1296) );
  XNOR U2241 ( .A(x[295]), .B(y[295]), .Z(n1297) );
  XNOR U2242 ( .A(n1296), .B(n1297), .Z(n1298) );
  XOR U2243 ( .A(n1299), .B(n1298), .Z(n1645) );
  XOR U2244 ( .A(x[303]), .B(y[303]), .Z(n1106) );
  XOR U2245 ( .A(x[299]), .B(y[299]), .Z(n1103) );
  XNOR U2246 ( .A(x[301]), .B(y[301]), .Z(n1104) );
  XNOR U2247 ( .A(n1103), .B(n1104), .Z(n1105) );
  XOR U2248 ( .A(n1106), .B(n1105), .Z(n1643) );
  XOR U2249 ( .A(x[309]), .B(y[309]), .Z(n1094) );
  XOR U2250 ( .A(x[305]), .B(y[305]), .Z(n1091) );
  XNOR U2251 ( .A(x[307]), .B(y[307]), .Z(n1092) );
  XNOR U2252 ( .A(n1091), .B(n1092), .Z(n1093) );
  XNOR U2253 ( .A(n1094), .B(n1093), .Z(n1642) );
  XNOR U2254 ( .A(n1643), .B(n1642), .Z(n1644) );
  XNOR U2255 ( .A(n1645), .B(n1644), .Z(n1541) );
  XOR U2256 ( .A(x[315]), .B(y[315]), .Z(n1100) );
  XOR U2257 ( .A(x[311]), .B(y[311]), .Z(n1097) );
  XNOR U2258 ( .A(x[313]), .B(y[313]), .Z(n1098) );
  XNOR U2259 ( .A(n1097), .B(n1098), .Z(n1099) );
  XOR U2260 ( .A(n1100), .B(n1099), .Z(n1904) );
  XOR U2261 ( .A(x[321]), .B(y[321]), .Z(n349) );
  XOR U2262 ( .A(x[317]), .B(y[317]), .Z(n346) );
  XNOR U2263 ( .A(x[319]), .B(y[319]), .Z(n347) );
  XNOR U2264 ( .A(n346), .B(n347), .Z(n348) );
  XOR U2265 ( .A(n349), .B(n348), .Z(n1902) );
  XOR U2266 ( .A(x[327]), .B(y[327]), .Z(n337) );
  XOR U2267 ( .A(x[323]), .B(y[323]), .Z(n334) );
  XNOR U2268 ( .A(x[325]), .B(y[325]), .Z(n335) );
  XNOR U2269 ( .A(n334), .B(n335), .Z(n336) );
  XNOR U2270 ( .A(n337), .B(n336), .Z(n1901) );
  XNOR U2271 ( .A(n1902), .B(n1901), .Z(n1903) );
  XNOR U2272 ( .A(n1904), .B(n1903), .Z(n1540) );
  XOR U2273 ( .A(n1541), .B(n1540), .Z(n1543) );
  XOR U2274 ( .A(x[333]), .B(y[333]), .Z(n343) );
  XOR U2275 ( .A(x[329]), .B(y[329]), .Z(n340) );
  XNOR U2276 ( .A(x[331]), .B(y[331]), .Z(n341) );
  XNOR U2277 ( .A(n340), .B(n341), .Z(n342) );
  XOR U2278 ( .A(n343), .B(n342), .Z(n1928) );
  XOR U2279 ( .A(x[339]), .B(y[339]), .Z(n325) );
  XOR U2280 ( .A(x[335]), .B(y[335]), .Z(n322) );
  XNOR U2281 ( .A(x[337]), .B(y[337]), .Z(n323) );
  XNOR U2282 ( .A(n322), .B(n323), .Z(n324) );
  XOR U2283 ( .A(n325), .B(n324), .Z(n1926) );
  XOR U2284 ( .A(x[345]), .B(y[345]), .Z(n313) );
  XOR U2285 ( .A(x[341]), .B(y[341]), .Z(n310) );
  XNOR U2286 ( .A(x[343]), .B(y[343]), .Z(n311) );
  XNOR U2287 ( .A(n310), .B(n311), .Z(n312) );
  XNOR U2288 ( .A(n313), .B(n312), .Z(n1925) );
  XNOR U2289 ( .A(n1926), .B(n1925), .Z(n1927) );
  XNOR U2290 ( .A(n1928), .B(n1927), .Z(n1542) );
  XNOR U2291 ( .A(n1543), .B(n1542), .Z(n1482) );
  XOR U2292 ( .A(x[351]), .B(y[351]), .Z(n319) );
  XOR U2293 ( .A(x[347]), .B(y[347]), .Z(n316) );
  XNOR U2294 ( .A(x[349]), .B(y[349]), .Z(n317) );
  XNOR U2295 ( .A(n316), .B(n317), .Z(n318) );
  XOR U2296 ( .A(n319), .B(n318), .Z(n1711) );
  XOR U2297 ( .A(x[357]), .B(y[357]), .Z(n278) );
  XOR U2298 ( .A(x[353]), .B(y[353]), .Z(n275) );
  XNOR U2299 ( .A(x[355]), .B(y[355]), .Z(n276) );
  XNOR U2300 ( .A(n275), .B(n276), .Z(n277) );
  XOR U2301 ( .A(n278), .B(n277), .Z(n1709) );
  XOR U2302 ( .A(x[363]), .B(y[363]), .Z(n290) );
  XOR U2303 ( .A(x[359]), .B(y[359]), .Z(n287) );
  XNOR U2304 ( .A(x[361]), .B(y[361]), .Z(n288) );
  XNOR U2305 ( .A(n287), .B(n288), .Z(n289) );
  XNOR U2306 ( .A(n290), .B(n289), .Z(n1708) );
  XNOR U2307 ( .A(n1709), .B(n1708), .Z(n1710) );
  XNOR U2308 ( .A(n1711), .B(n1710), .Z(n1546) );
  XOR U2309 ( .A(x[369]), .B(y[369]), .Z(n284) );
  XOR U2310 ( .A(x[365]), .B(y[365]), .Z(n281) );
  XNOR U2311 ( .A(x[367]), .B(y[367]), .Z(n282) );
  XNOR U2312 ( .A(n281), .B(n282), .Z(n283) );
  XOR U2313 ( .A(n284), .B(n283), .Z(n1148) );
  XOR U2314 ( .A(x[375]), .B(y[375]), .Z(n466) );
  XOR U2315 ( .A(x[371]), .B(y[371]), .Z(n463) );
  XNOR U2316 ( .A(x[373]), .B(y[373]), .Z(n464) );
  XNOR U2317 ( .A(n463), .B(n464), .Z(n465) );
  XOR U2318 ( .A(n466), .B(n465), .Z(n1146) );
  XOR U2319 ( .A(x[381]), .B(y[381]), .Z(n454) );
  XOR U2320 ( .A(x[377]), .B(y[377]), .Z(n451) );
  XNOR U2321 ( .A(x[379]), .B(y[379]), .Z(n452) );
  XNOR U2322 ( .A(n451), .B(n452), .Z(n453) );
  XNOR U2323 ( .A(n454), .B(n453), .Z(n1145) );
  XNOR U2324 ( .A(n1146), .B(n1145), .Z(n1147) );
  XOR U2325 ( .A(n1148), .B(n1147), .Z(n1547) );
  XNOR U2326 ( .A(n1546), .B(n1547), .Z(n1548) );
  XOR U2327 ( .A(x[387]), .B(y[387]), .Z(n488) );
  XOR U2328 ( .A(x[383]), .B(y[383]), .Z(n485) );
  XNOR U2329 ( .A(x[385]), .B(y[385]), .Z(n486) );
  XNOR U2330 ( .A(n485), .B(n486), .Z(n487) );
  XOR U2331 ( .A(n488), .B(n487), .Z(n478) );
  XOR U2332 ( .A(x[393]), .B(y[393]), .Z(n512) );
  XOR U2333 ( .A(x[389]), .B(y[389]), .Z(n509) );
  XOR U2334 ( .A(x[391]), .B(y[391]), .Z(n510) );
  XOR U2335 ( .A(n512), .B(n511), .Z(n476) );
  XOR U2336 ( .A(x[401]), .B(y[401]), .Z(n396) );
  XOR U2337 ( .A(x[395]), .B(y[395]), .Z(n393) );
  XNOR U2338 ( .A(x[397]), .B(y[397]), .Z(n394) );
  XNOR U2339 ( .A(n393), .B(n394), .Z(n395) );
  XNOR U2340 ( .A(n396), .B(n395), .Z(n475) );
  XNOR U2341 ( .A(n476), .B(n475), .Z(n477) );
  XOR U2342 ( .A(n478), .B(n477), .Z(n1549) );
  XOR U2343 ( .A(n1548), .B(n1549), .Z(n1481) );
  XOR U2344 ( .A(x[750]), .B(y[750]), .Z(n1130) );
  XOR U2345 ( .A(x[358]), .B(y[358]), .Z(n1127) );
  XNOR U2346 ( .A(x[752]), .B(y[752]), .Z(n1128) );
  XNOR U2347 ( .A(n1127), .B(n1128), .Z(n1129) );
  XOR U2348 ( .A(n1130), .B(n1129), .Z(n387) );
  XOR U2349 ( .A(x[461]), .B(y[461]), .Z(n584) );
  XOR U2350 ( .A(x[453]), .B(y[453]), .Z(n581) );
  XOR U2351 ( .A(x[457]), .B(y[457]), .Z(n582) );
  XOR U2352 ( .A(n584), .B(n583), .Z(n388) );
  XOR U2353 ( .A(n387), .B(n388), .Z(n390) );
  XOR U2354 ( .A(x[473]), .B(y[473]), .Z(n460) );
  XOR U2355 ( .A(x[465]), .B(y[465]), .Z(n457) );
  XOR U2356 ( .A(x[469]), .B(y[469]), .Z(n458) );
  XOR U2357 ( .A(n460), .B(n459), .Z(n389) );
  XNOR U2358 ( .A(n390), .B(n389), .Z(n1387) );
  XOR U2359 ( .A(x[449]), .B(y[449]), .Z(n636) );
  XOR U2360 ( .A(x[441]), .B(y[441]), .Z(n633) );
  XOR U2361 ( .A(x[445]), .B(y[445]), .Z(n634) );
  XOR U2362 ( .A(n636), .B(n635), .Z(n482) );
  XOR U2363 ( .A(x[182]), .B(y[182]), .Z(n1160) );
  XOR U2364 ( .A(x[111]), .B(y[111]), .Z(n1157) );
  XOR U2365 ( .A(x[184]), .B(y[184]), .Z(n1158) );
  XNOR U2366 ( .A(n1160), .B(n1159), .Z(n481) );
  XNOR U2367 ( .A(n482), .B(n481), .Z(n484) );
  XOR U2368 ( .A(x[437]), .B(y[437]), .Z(n606) );
  XOR U2369 ( .A(x[429]), .B(y[429]), .Z(n603) );
  XOR U2370 ( .A(x[433]), .B(y[433]), .Z(n604) );
  XOR U2371 ( .A(n606), .B(n605), .Z(n483) );
  XOR U2372 ( .A(n484), .B(n483), .Z(n1385) );
  XOR U2373 ( .A(x[425]), .B(y[425]), .Z(n376) );
  XOR U2374 ( .A(x[417]), .B(y[417]), .Z(n374) );
  XNOR U2375 ( .A(x[421]), .B(y[421]), .Z(n375) );
  XOR U2376 ( .A(n374), .B(n375), .Z(n377) );
  XNOR U2377 ( .A(n376), .B(n377), .Z(n503) );
  XOR U2378 ( .A(x[744]), .B(y[744]), .Z(n552) );
  XOR U2379 ( .A(x[746]), .B(y[746]), .Z(n549) );
  XOR U2380 ( .A(x[748]), .B(y[748]), .Z(n550) );
  XOR U2381 ( .A(n552), .B(n551), .Z(n504) );
  XOR U2382 ( .A(n503), .B(n504), .Z(n506) );
  XOR U2383 ( .A(x[413]), .B(y[413]), .Z(n423) );
  XOR U2384 ( .A(x[405]), .B(y[405]), .Z(n421) );
  XNOR U2385 ( .A(x[409]), .B(y[409]), .Z(n422) );
  XOR U2386 ( .A(n421), .B(n422), .Z(n424) );
  XNOR U2387 ( .A(n423), .B(n424), .Z(n505) );
  XNOR U2388 ( .A(n506), .B(n505), .Z(n1384) );
  XNOR U2389 ( .A(n1385), .B(n1384), .Z(n1386) );
  XNOR U2390 ( .A(n1387), .B(n1386), .Z(n1480) );
  XOR U2391 ( .A(n1482), .B(n1483), .Z(n1381) );
  XOR U2392 ( .A(x[681]), .B(y[681]), .Z(n236) );
  XOR U2393 ( .A(x[675]), .B(y[675]), .Z(n233) );
  XNOR U2394 ( .A(x[689]), .B(y[689]), .Z(n234) );
  XNOR U2395 ( .A(n233), .B(n234), .Z(n235) );
  XOR U2396 ( .A(n236), .B(n235), .Z(n1232) );
  XOR U2397 ( .A(x[48]), .B(y[48]), .Z(n2092) );
  XOR U2398 ( .A(x[52]), .B(y[52]), .Z(n2089) );
  XNOR U2399 ( .A(x[399]), .B(y[399]), .Z(n2090) );
  XNOR U2400 ( .A(n2089), .B(n2090), .Z(n2091) );
  XOR U2401 ( .A(n2092), .B(n2091), .Z(n1230) );
  XOR U2402 ( .A(x[687]), .B(y[687]), .Z(n230) );
  XOR U2403 ( .A(x[683]), .B(y[683]), .Z(n227) );
  XNOR U2404 ( .A(x[685]), .B(y[685]), .Z(n228) );
  XNOR U2405 ( .A(n227), .B(n228), .Z(n229) );
  XNOR U2406 ( .A(n230), .B(n229), .Z(n1229) );
  XNOR U2407 ( .A(n1230), .B(n1229), .Z(n1231) );
  XNOR U2408 ( .A(n1232), .B(n1231), .Z(n1420) );
  XOR U2409 ( .A(x[531]), .B(y[531]), .Z(n1112) );
  XOR U2410 ( .A(x[525]), .B(y[525]), .Z(n1109) );
  XNOR U2411 ( .A(x[529]), .B(y[529]), .Z(n1110) );
  XNOR U2412 ( .A(n1109), .B(n1110), .Z(n1111) );
  XOR U2413 ( .A(n1112), .B(n1111), .Z(n442) );
  XOR U2414 ( .A(x[156]), .B(y[156]), .Z(n564) );
  XOR U2415 ( .A(x[129]), .B(y[129]), .Z(n561) );
  XOR U2416 ( .A(x[160]), .B(y[160]), .Z(n562) );
  XOR U2417 ( .A(n564), .B(n563), .Z(n440) );
  XOR U2418 ( .A(x[537]), .B(y[537]), .Z(n1118) );
  XOR U2419 ( .A(x[533]), .B(y[533]), .Z(n1115) );
  XNOR U2420 ( .A(x[535]), .B(y[535]), .Z(n1116) );
  XNOR U2421 ( .A(n1115), .B(n1116), .Z(n1117) );
  XNOR U2422 ( .A(n1118), .B(n1117), .Z(n439) );
  XNOR U2423 ( .A(n440), .B(n439), .Z(n441) );
  XOR U2424 ( .A(n442), .B(n441), .Z(n1421) );
  XNOR U2425 ( .A(n1420), .B(n1421), .Z(n1422) );
  XOR U2426 ( .A(x[543]), .B(y[543]), .Z(n195) );
  XOR U2427 ( .A(x[539]), .B(y[539]), .Z(n192) );
  XNOR U2428 ( .A(x[541]), .B(y[541]), .Z(n193) );
  XNOR U2429 ( .A(n192), .B(n193), .Z(n194) );
  XOR U2430 ( .A(n195), .B(n194), .Z(n361) );
  XOR U2431 ( .A(x[758]), .B(y[758]), .Z(n1124) );
  XOR U2432 ( .A(x[760]), .B(y[760]), .Z(n1121) );
  XNOR U2433 ( .A(x[762]), .B(y[762]), .Z(n1122) );
  XNOR U2434 ( .A(n1121), .B(n1122), .Z(n1123) );
  XOR U2435 ( .A(n1124), .B(n1123), .Z(n359) );
  XOR U2436 ( .A(x[549]), .B(y[549]), .Z(n189) );
  XOR U2437 ( .A(x[545]), .B(y[545]), .Z(n186) );
  XNOR U2438 ( .A(x[547]), .B(y[547]), .Z(n187) );
  XNOR U2439 ( .A(n186), .B(n187), .Z(n188) );
  XNOR U2440 ( .A(n189), .B(n188), .Z(n358) );
  XNOR U2441 ( .A(n359), .B(n358), .Z(n360) );
  XOR U2442 ( .A(n361), .B(n360), .Z(n1423) );
  XNOR U2443 ( .A(n1422), .B(n1423), .Z(n932) );
  XOR U2444 ( .A(x[643]), .B(y[643]), .Z(n821) );
  XOR U2445 ( .A(x[665]), .B(y[665]), .Z(n818) );
  XNOR U2446 ( .A(x[705]), .B(y[705]), .Z(n819) );
  XNOR U2447 ( .A(n818), .B(n819), .Z(n820) );
  XOR U2448 ( .A(n821), .B(n820), .Z(n570) );
  XOR U2449 ( .A(x[78]), .B(y[78]), .Z(n494) );
  XOR U2450 ( .A(x[80]), .B(y[80]), .Z(n491) );
  XNOR U2451 ( .A(x[183]), .B(y[183]), .Z(n492) );
  XNOR U2452 ( .A(n491), .B(n492), .Z(n493) );
  XOR U2453 ( .A(n494), .B(n493), .Z(n568) );
  XOR U2454 ( .A(x[703]), .B(y[703]), .Z(n827) );
  XOR U2455 ( .A(x[645]), .B(y[645]), .Z(n824) );
  XNOR U2456 ( .A(x[663]), .B(y[663]), .Z(n825) );
  XNOR U2457 ( .A(n824), .B(n825), .Z(n826) );
  XNOR U2458 ( .A(n827), .B(n826), .Z(n567) );
  XNOR U2459 ( .A(n568), .B(n567), .Z(n569) );
  XNOR U2460 ( .A(n570), .B(n569), .Z(n1486) );
  XOR U2461 ( .A(x[711]), .B(y[711]), .Z(n748) );
  XOR U2462 ( .A(x[653]), .B(y[653]), .Z(n745) );
  XNOR U2463 ( .A(x[713]), .B(y[713]), .Z(n746) );
  XNOR U2464 ( .A(n745), .B(n746), .Z(n747) );
  XOR U2465 ( .A(n748), .B(n747), .Z(n546) );
  XOR U2466 ( .A(x[784]), .B(y[784]), .Z(n907) );
  XOR U2467 ( .A(x[786]), .B(y[786]), .Z(n904) );
  XNOR U2468 ( .A(x[788]), .B(y[788]), .Z(n905) );
  XNOR U2469 ( .A(n904), .B(n905), .Z(n906) );
  XOR U2470 ( .A(n907), .B(n906), .Z(n544) );
  XOR U2471 ( .A(x[707]), .B(y[707]), .Z(n742) );
  XOR U2472 ( .A(x[671]), .B(y[671]), .Z(n739) );
  XNOR U2473 ( .A(x[709]), .B(y[709]), .Z(n740) );
  XNOR U2474 ( .A(n739), .B(n740), .Z(n741) );
  XNOR U2475 ( .A(n742), .B(n741), .Z(n543) );
  XNOR U2476 ( .A(n544), .B(n543), .Z(n545) );
  XOR U2477 ( .A(n546), .B(n545), .Z(n1487) );
  XNOR U2478 ( .A(n1486), .B(n1487), .Z(n1489) );
  XOR U2479 ( .A(x[621]), .B(y[621]), .Z(n730) );
  XOR U2480 ( .A(x[619]), .B(y[619]), .Z(n727) );
  XNOR U2481 ( .A(x[725]), .B(y[725]), .Z(n728) );
  XNOR U2482 ( .A(n727), .B(n728), .Z(n729) );
  XOR U2483 ( .A(n730), .B(n729), .Z(n1190) );
  XOR U2484 ( .A(x[106]), .B(y[106]), .Z(n618) );
  XOR U2485 ( .A(x[108]), .B(y[108]), .Z(n615) );
  XNOR U2486 ( .A(x[165]), .B(y[165]), .Z(n616) );
  XNOR U2487 ( .A(n615), .B(n616), .Z(n617) );
  XOR U2488 ( .A(n618), .B(n617), .Z(n1188) );
  XOR U2489 ( .A(x[625]), .B(y[625]), .Z(n724) );
  XOR U2490 ( .A(x[623]), .B(y[623]), .Z(n721) );
  XNOR U2491 ( .A(x[723]), .B(y[723]), .Z(n722) );
  XNOR U2492 ( .A(n721), .B(n722), .Z(n723) );
  XNOR U2493 ( .A(n724), .B(n723), .Z(n1187) );
  XNOR U2494 ( .A(n1188), .B(n1187), .Z(n1189) );
  XNOR U2495 ( .A(n1190), .B(n1189), .Z(n1488) );
  XOR U2496 ( .A(n1489), .B(n1488), .Z(n930) );
  XOR U2497 ( .A(x[597]), .B(y[597]), .Z(n876) );
  XOR U2498 ( .A(x[593]), .B(y[593]), .Z(n873) );
  XNOR U2499 ( .A(x[595]), .B(y[595]), .Z(n874) );
  XNOR U2500 ( .A(n873), .B(n874), .Z(n875) );
  XOR U2501 ( .A(n876), .B(n875), .Z(n574) );
  XOR U2502 ( .A(x[770]), .B(y[770]), .Z(n760) );
  XOR U2503 ( .A(x[376]), .B(y[376]), .Z(n757) );
  XNOR U2504 ( .A(x[772]), .B(y[772]), .Z(n758) );
  XNOR U2505 ( .A(n757), .B(n758), .Z(n759) );
  XNOR U2506 ( .A(n760), .B(n759), .Z(n573) );
  XNOR U2507 ( .A(n574), .B(n573), .Z(n576) );
  XOR U2508 ( .A(x[591]), .B(y[591]), .Z(n882) );
  XOR U2509 ( .A(x[587]), .B(y[587]), .Z(n879) );
  XNOR U2510 ( .A(x[589]), .B(y[589]), .Z(n880) );
  XNOR U2511 ( .A(n879), .B(n880), .Z(n881) );
  XOR U2512 ( .A(n882), .B(n881), .Z(n575) );
  XOR U2513 ( .A(n576), .B(n575), .Z(n1459) );
  XOR U2514 ( .A(x[693]), .B(y[693]), .Z(n807) );
  XOR U2515 ( .A(x[657]), .B(y[657]), .Z(n805) );
  XNOR U2516 ( .A(x[695]), .B(y[695]), .Z(n806) );
  XOR U2517 ( .A(n805), .B(n806), .Z(n808) );
  XNOR U2518 ( .A(n807), .B(n808), .Z(n1655) );
  XOR U2519 ( .A(x[66]), .B(y[66]), .Z(n2299) );
  XOR U2520 ( .A(x[70]), .B(y[70]), .Z(n2296) );
  XOR U2521 ( .A(x[72]), .B(y[72]), .Z(n2297) );
  XOR U2522 ( .A(n2299), .B(n2298), .Z(n1654) );
  XOR U2523 ( .A(n1655), .B(n1654), .Z(n1657) );
  XOR U2524 ( .A(x[651]), .B(y[651]), .Z(n795) );
  XOR U2525 ( .A(x[655]), .B(y[655]), .Z(n793) );
  XNOR U2526 ( .A(x[697]), .B(y[697]), .Z(n794) );
  XOR U2527 ( .A(n793), .B(n794), .Z(n796) );
  XNOR U2528 ( .A(n795), .B(n796), .Z(n1656) );
  XOR U2529 ( .A(n1657), .B(n1656), .Z(n1457) );
  XOR U2530 ( .A(x[579]), .B(y[579]), .Z(n772) );
  XOR U2531 ( .A(x[575]), .B(y[575]), .Z(n769) );
  XNOR U2532 ( .A(x[577]), .B(y[577]), .Z(n770) );
  XNOR U2533 ( .A(n769), .B(n770), .Z(n771) );
  XOR U2534 ( .A(n772), .B(n771), .Z(n654) );
  XOR U2535 ( .A(x[130]), .B(y[130]), .Z(n558) );
  XOR U2536 ( .A(x[132]), .B(y[132]), .Z(n555) );
  XNOR U2537 ( .A(x[147]), .B(y[147]), .Z(n556) );
  XNOR U2538 ( .A(n555), .B(n556), .Z(n557) );
  XOR U2539 ( .A(n558), .B(n557), .Z(n652) );
  XOR U2540 ( .A(x[585]), .B(y[585]), .Z(n766) );
  XOR U2541 ( .A(x[581]), .B(y[581]), .Z(n763) );
  XNOR U2542 ( .A(x[583]), .B(y[583]), .Z(n764) );
  XNOR U2543 ( .A(n763), .B(n764), .Z(n765) );
  XNOR U2544 ( .A(n766), .B(n765), .Z(n651) );
  XNOR U2545 ( .A(n652), .B(n651), .Z(n653) );
  XNOR U2546 ( .A(n654), .B(n653), .Z(n1456) );
  XNOR U2547 ( .A(n1457), .B(n1456), .Z(n1458) );
  XOR U2548 ( .A(n1459), .B(n1458), .Z(n929) );
  XOR U2549 ( .A(n930), .B(n929), .Z(n931) );
  XNOR U2550 ( .A(n932), .B(n931), .Z(n1380) );
  XOR U2551 ( .A(n1381), .B(n1380), .Z(n1383) );
  XOR U2552 ( .A(x[617]), .B(y[617]), .Z(n895) );
  XOR U2553 ( .A(x[615]), .B(y[615]), .Z(n892) );
  XOR U2554 ( .A(x[727]), .B(y[727]), .Z(n893) );
  XOR U2555 ( .A(n895), .B(n894), .Z(n600) );
  XOR U2556 ( .A(x[774]), .B(y[774]), .Z(n1030) );
  XOR U2557 ( .A(x[380]), .B(y[380]), .Z(n1027) );
  XNOR U2558 ( .A(x[776]), .B(y[776]), .Z(n1028) );
  XNOR U2559 ( .A(n1027), .B(n1028), .Z(n1029) );
  XNOR U2560 ( .A(n1030), .B(n1029), .Z(n599) );
  XNOR U2561 ( .A(n600), .B(n599), .Z(n601) );
  XOR U2562 ( .A(x[613]), .B(y[613]), .Z(n901) );
  XOR U2563 ( .A(x[611]), .B(y[611]), .Z(n898) );
  XOR U2564 ( .A(x[729]), .B(y[729]), .Z(n899) );
  XOR U2565 ( .A(n901), .B(n900), .Z(n602) );
  XNOR U2566 ( .A(n601), .B(n602), .Z(n1470) );
  XOR U2567 ( .A(x[699]), .B(y[699]), .Z(n247) );
  XOR U2568 ( .A(x[661]), .B(y[661]), .Z(n245) );
  XNOR U2569 ( .A(x[701]), .B(y[701]), .Z(n246) );
  XOR U2570 ( .A(n245), .B(n246), .Z(n248) );
  XNOR U2571 ( .A(n247), .B(n248), .Z(n1678) );
  XOR U2572 ( .A(x[790]), .B(y[790]), .Z(n814) );
  XOR U2573 ( .A(x[394]), .B(y[394]), .Z(n812) );
  XNOR U2574 ( .A(x[792]), .B(y[792]), .Z(n813) );
  XOR U2575 ( .A(n812), .B(n813), .Z(n815) );
  XOR U2576 ( .A(n814), .B(n815), .Z(n1679) );
  XNOR U2577 ( .A(n1678), .B(n1679), .Z(n1680) );
  XOR U2578 ( .A(x[649]), .B(y[649]), .Z(n253) );
  XOR U2579 ( .A(x[647]), .B(y[647]), .Z(n251) );
  XNOR U2580 ( .A(x[659]), .B(y[659]), .Z(n252) );
  XOR U2581 ( .A(n251), .B(n252), .Z(n254) );
  XOR U2582 ( .A(n253), .B(n254), .Z(n1681) );
  XOR U2583 ( .A(n1680), .B(n1681), .Z(n1469) );
  XOR U2584 ( .A(x[609]), .B(y[609]), .Z(n1036) );
  XOR U2585 ( .A(x[605]), .B(y[605]), .Z(n1033) );
  XNOR U2586 ( .A(x[607]), .B(y[607]), .Z(n1034) );
  XNOR U2587 ( .A(n1033), .B(n1034), .Z(n1035) );
  XOR U2588 ( .A(n1036), .B(n1035), .Z(n578) );
  XOR U2589 ( .A(x[116]), .B(y[116]), .Z(n596) );
  XOR U2590 ( .A(x[120]), .B(y[120]), .Z(n593) );
  XNOR U2591 ( .A(x[124]), .B(y[124]), .Z(n594) );
  XNOR U2592 ( .A(n593), .B(n594), .Z(n595) );
  XNOR U2593 ( .A(n596), .B(n595), .Z(n577) );
  XNOR U2594 ( .A(n578), .B(n577), .Z(n579) );
  XOR U2595 ( .A(x[603]), .B(y[603]), .Z(n1042) );
  XOR U2596 ( .A(x[599]), .B(y[599]), .Z(n1039) );
  XNOR U2597 ( .A(x[601]), .B(y[601]), .Z(n1040) );
  XNOR U2598 ( .A(n1039), .B(n1040), .Z(n1041) );
  XOR U2599 ( .A(n1042), .B(n1041), .Z(n580) );
  XNOR U2600 ( .A(n579), .B(n580), .Z(n1468) );
  XOR U2601 ( .A(n1470), .B(n1471), .Z(n987) );
  XOR U2602 ( .A(x[637]), .B(y[637]), .Z(n913) );
  XOR U2603 ( .A(x[635]), .B(y[635]), .Z(n910) );
  XNOR U2604 ( .A(x[717]), .B(y[717]), .Z(n911) );
  XNOR U2605 ( .A(n910), .B(n911), .Z(n912) );
  XOR U2606 ( .A(n913), .B(n912), .Z(n302) );
  XOR U2607 ( .A(x[92]), .B(y[92]), .Z(n436) );
  XOR U2608 ( .A(x[94]), .B(y[94]), .Z(n433) );
  XNOR U2609 ( .A(x[96]), .B(y[96]), .Z(n434) );
  XNOR U2610 ( .A(n433), .B(n434), .Z(n435) );
  XOR U2611 ( .A(n436), .B(n435), .Z(n301) );
  XOR U2612 ( .A(x[641]), .B(y[641]), .Z(n919) );
  XOR U2613 ( .A(x[639]), .B(y[639]), .Z(n916) );
  XNOR U2614 ( .A(x[715]), .B(y[715]), .Z(n917) );
  XNOR U2615 ( .A(n916), .B(n917), .Z(n918) );
  XNOR U2616 ( .A(n919), .B(n918), .Z(n300) );
  XOR U2617 ( .A(n301), .B(n300), .Z(n303) );
  XOR U2618 ( .A(n302), .B(n303), .Z(n986) );
  XOR U2619 ( .A(x[629]), .B(y[629]), .Z(n864) );
  XOR U2620 ( .A(x[627]), .B(y[627]), .Z(n861) );
  XOR U2621 ( .A(x[721]), .B(y[721]), .Z(n862) );
  XOR U2622 ( .A(n864), .B(n863), .Z(n623) );
  XOR U2623 ( .A(x[778]), .B(y[778]), .Z(n718) );
  XOR U2624 ( .A(x[780]), .B(y[780]), .Z(n715) );
  XOR U2625 ( .A(x[782]), .B(y[782]), .Z(n716) );
  XOR U2626 ( .A(n718), .B(n717), .Z(n622) );
  XOR U2627 ( .A(x[633]), .B(y[633]), .Z(n858) );
  XOR U2628 ( .A(x[631]), .B(y[631]), .Z(n855) );
  XOR U2629 ( .A(x[719]), .B(y[719]), .Z(n856) );
  XNOR U2630 ( .A(n858), .B(n857), .Z(n621) );
  XOR U2631 ( .A(n622), .B(n621), .Z(n624) );
  XNOR U2632 ( .A(n623), .B(n624), .Z(n985) );
  XOR U2633 ( .A(n986), .B(n985), .Z(n988) );
  XOR U2634 ( .A(n987), .B(n988), .Z(n1536) );
  XOR U2635 ( .A(x[521]), .B(y[521]), .Z(n1054) );
  XOR U2636 ( .A(x[513]), .B(y[513]), .Z(n1051) );
  XNOR U2637 ( .A(x[517]), .B(y[517]), .Z(n1052) );
  XNOR U2638 ( .A(n1051), .B(n1052), .Z(n1053) );
  XOR U2639 ( .A(n1054), .B(n1053), .Z(n418) );
  XOR U2640 ( .A(x[754]), .B(y[754]), .Z(n1072) );
  XOR U2641 ( .A(x[362]), .B(y[362]), .Z(n1069) );
  XNOR U2642 ( .A(x[756]), .B(y[756]), .Z(n1070) );
  XNOR U2643 ( .A(n1069), .B(n1070), .Z(n1071) );
  XNOR U2644 ( .A(n1072), .B(n1071), .Z(n417) );
  XNOR U2645 ( .A(n418), .B(n417), .Z(n420) );
  XOR U2646 ( .A(x[509]), .B(y[509]), .Z(n1060) );
  XOR U2647 ( .A(x[501]), .B(y[501]), .Z(n1057) );
  XNOR U2648 ( .A(x[505]), .B(y[505]), .Z(n1058) );
  XNOR U2649 ( .A(n1057), .B(n1058), .Z(n1059) );
  XOR U2650 ( .A(n1060), .B(n1059), .Z(n419) );
  XOR U2651 ( .A(n420), .B(n419), .Z(n1393) );
  XOR U2652 ( .A(x[54]), .B(y[54]), .Z(n783) );
  XOR U2653 ( .A(x[56]), .B(y[56]), .Z(n781) );
  XNOR U2654 ( .A(x[201]), .B(y[201]), .Z(n782) );
  XOR U2655 ( .A(n781), .B(n782), .Z(n784) );
  XNOR U2656 ( .A(n783), .B(n784), .Z(n1254) );
  XOR U2657 ( .A(x[200]), .B(y[200]), .Z(n789) );
  XOR U2658 ( .A(x[202]), .B(y[202]), .Z(n787) );
  XNOR U2659 ( .A(x[799]), .B(y[799]), .Z(n788) );
  XOR U2660 ( .A(n787), .B(n788), .Z(n790) );
  XOR U2661 ( .A(n789), .B(n790), .Z(n1255) );
  XNOR U2662 ( .A(n1254), .B(n1255), .Z(n1257) );
  XOR U2663 ( .A(x[798]), .B(y[798]), .Z(n223) );
  XNOR U2664 ( .A(x[204]), .B(y[204]), .Z(n222) );
  XOR U2665 ( .A(oglobal[0]), .B(n222), .Z(n224) );
  XNOR U2666 ( .A(n223), .B(n224), .Z(n1256) );
  XOR U2667 ( .A(n1257), .B(n1256), .Z(n1391) );
  XOR U2668 ( .A(x[497]), .B(y[497]), .Z(n1078) );
  XOR U2669 ( .A(x[489]), .B(y[489]), .Z(n1075) );
  XNOR U2670 ( .A(x[493]), .B(y[493]), .Z(n1076) );
  XNOR U2671 ( .A(n1075), .B(n1076), .Z(n1077) );
  XOR U2672 ( .A(n1078), .B(n1077), .Z(n411) );
  XOR U2673 ( .A(x[168]), .B(y[168]), .Z(n1136) );
  XOR U2674 ( .A(x[170]), .B(y[170]), .Z(n1133) );
  XNOR U2675 ( .A(x[174]), .B(y[174]), .Z(n1134) );
  XNOR U2676 ( .A(n1133), .B(n1134), .Z(n1135) );
  XOR U2677 ( .A(n1136), .B(n1135), .Z(n412) );
  XOR U2678 ( .A(n411), .B(n412), .Z(n414) );
  XOR U2679 ( .A(x[485]), .B(y[485]), .Z(n1084) );
  XOR U2680 ( .A(x[477]), .B(y[477]), .Z(n1081) );
  XNOR U2681 ( .A(x[481]), .B(y[481]), .Z(n1082) );
  XNOR U2682 ( .A(n1081), .B(n1082), .Z(n1083) );
  XOR U2683 ( .A(n1084), .B(n1083), .Z(n413) );
  XNOR U2684 ( .A(n414), .B(n413), .Z(n1390) );
  XNOR U2685 ( .A(n1391), .B(n1390), .Z(n1392) );
  XNOR U2686 ( .A(n1393), .B(n1392), .Z(n1535) );
  XOR U2687 ( .A(x[567]), .B(y[567]), .Z(n213) );
  XOR U2688 ( .A(x[563]), .B(y[563]), .Z(n210) );
  XNOR U2689 ( .A(x[565]), .B(y[565]), .Z(n211) );
  XNOR U2690 ( .A(n210), .B(n211), .Z(n212) );
  XOR U2691 ( .A(n213), .B(n212), .Z(n630) );
  XOR U2692 ( .A(x[764]), .B(y[764]), .Z(n958) );
  XOR U2693 ( .A(x[766]), .B(y[766]), .Z(n955) );
  XNOR U2694 ( .A(x[768]), .B(y[768]), .Z(n956) );
  XNOR U2695 ( .A(n955), .B(n956), .Z(n957) );
  XOR U2696 ( .A(n958), .B(n957), .Z(n628) );
  XOR U2697 ( .A(x[573]), .B(y[573]), .Z(n207) );
  XOR U2698 ( .A(x[569]), .B(y[569]), .Z(n204) );
  XNOR U2699 ( .A(x[571]), .B(y[571]), .Z(n205) );
  XNOR U2700 ( .A(n204), .B(n205), .Z(n206) );
  XNOR U2701 ( .A(n207), .B(n206), .Z(n627) );
  XNOR U2702 ( .A(n628), .B(n627), .Z(n629) );
  XNOR U2703 ( .A(n630), .B(n629), .Z(n1429) );
  XOR U2704 ( .A(x[561]), .B(y[561]), .Z(n964) );
  XOR U2705 ( .A(x[557]), .B(y[557]), .Z(n961) );
  XNOR U2706 ( .A(x[559]), .B(y[559]), .Z(n962) );
  XNOR U2707 ( .A(n961), .B(n962), .Z(n963) );
  XOR U2708 ( .A(n964), .B(n963), .Z(n365) );
  XOR U2709 ( .A(x[144]), .B(y[144]), .Z(n1663) );
  XOR U2710 ( .A(x[146]), .B(y[146]), .Z(n1660) );
  XNOR U2711 ( .A(x[148]), .B(y[148]), .Z(n1661) );
  XNOR U2712 ( .A(n1660), .B(n1661), .Z(n1662) );
  XNOR U2713 ( .A(n1663), .B(n1662), .Z(n364) );
  XNOR U2714 ( .A(n365), .B(n364), .Z(n367) );
  XOR U2715 ( .A(x[555]), .B(y[555]), .Z(n970) );
  XOR U2716 ( .A(x[551]), .B(y[551]), .Z(n967) );
  XNOR U2717 ( .A(x[553]), .B(y[553]), .Z(n968) );
  XNOR U2718 ( .A(n967), .B(n968), .Z(n969) );
  XOR U2719 ( .A(n970), .B(n969), .Z(n366) );
  XOR U2720 ( .A(n367), .B(n366), .Z(n1427) );
  XOR U2721 ( .A(x[669]), .B(y[669]), .Z(n952) );
  XOR U2722 ( .A(x[667]), .B(y[667]), .Z(n949) );
  XNOR U2723 ( .A(x[679]), .B(y[679]), .Z(n950) );
  XNOR U2724 ( .A(n949), .B(n950), .Z(n951) );
  XOR U2725 ( .A(n952), .B(n951), .Z(n530) );
  XOR U2726 ( .A(x[794]), .B(y[794]), .Z(n802) );
  XOR U2727 ( .A(x[796]), .B(y[796]), .Z(n799) );
  XNOR U2728 ( .A(x[797]), .B(y[797]), .Z(n800) );
  XNOR U2729 ( .A(n799), .B(n800), .Z(n801) );
  XOR U2730 ( .A(n802), .B(n801), .Z(n528) );
  XOR U2731 ( .A(x[691]), .B(y[691]), .Z(n946) );
  XOR U2732 ( .A(x[673]), .B(y[673]), .Z(n943) );
  XNOR U2733 ( .A(x[677]), .B(y[677]), .Z(n944) );
  XNOR U2734 ( .A(n943), .B(n944), .Z(n945) );
  XNOR U2735 ( .A(n946), .B(n945), .Z(n527) );
  XNOR U2736 ( .A(n528), .B(n527), .Z(n529) );
  XNOR U2737 ( .A(n530), .B(n529), .Z(n1426) );
  XNOR U2738 ( .A(n1427), .B(n1426), .Z(n1428) );
  XOR U2739 ( .A(n1429), .B(n1428), .Z(n1534) );
  XOR U2740 ( .A(n1535), .B(n1534), .Z(n1537) );
  XNOR U2741 ( .A(n1536), .B(n1537), .Z(n1382) );
  XNOR U2742 ( .A(n1383), .B(n1382), .Z(n1444) );
  XNOR U2743 ( .A(n1445), .B(n1444), .Z(n1446) );
  XNOR U2744 ( .A(n1447), .B(n1446), .Z(o[0]) );
  NANDN U2745 ( .A(n163), .B(n162), .Z(n167) );
  NANDN U2746 ( .A(n165), .B(n164), .Z(n166) );
  AND U2747 ( .A(n167), .B(n166), .Z(n3404) );
  NANDN U2748 ( .A(n169), .B(n168), .Z(n173) );
  NANDN U2749 ( .A(n171), .B(n170), .Z(n172) );
  AND U2750 ( .A(n173), .B(n172), .Z(n3401) );
  NANDN U2751 ( .A(n175), .B(n174), .Z(n179) );
  NANDN U2752 ( .A(n177), .B(n176), .Z(n178) );
  NAND U2753 ( .A(n179), .B(n178), .Z(n3402) );
  XNOR U2754 ( .A(n3401), .B(n3402), .Z(n3403) );
  XOR U2755 ( .A(n3404), .B(n3403), .Z(n2889) );
  NANDN U2756 ( .A(n181), .B(n180), .Z(n185) );
  NAND U2757 ( .A(n183), .B(n182), .Z(n184) );
  AND U2758 ( .A(n185), .B(n184), .Z(n2732) );
  NANDN U2759 ( .A(n187), .B(n186), .Z(n191) );
  NAND U2760 ( .A(n189), .B(n188), .Z(n190) );
  NAND U2761 ( .A(n191), .B(n190), .Z(n2733) );
  XNOR U2762 ( .A(n2732), .B(n2733), .Z(n2735) );
  NANDN U2763 ( .A(n193), .B(n192), .Z(n197) );
  NAND U2764 ( .A(n195), .B(n194), .Z(n196) );
  AND U2765 ( .A(n197), .B(n196), .Z(n2734) );
  XOR U2766 ( .A(n2735), .B(n2734), .Z(n3288) );
  NANDN U2767 ( .A(n199), .B(n198), .Z(n203) );
  NAND U2768 ( .A(n201), .B(n200), .Z(n202) );
  AND U2769 ( .A(n203), .B(n202), .Z(n2786) );
  NANDN U2770 ( .A(n205), .B(n204), .Z(n209) );
  NAND U2771 ( .A(n207), .B(n206), .Z(n208) );
  NAND U2772 ( .A(n209), .B(n208), .Z(n2787) );
  XNOR U2773 ( .A(n2786), .B(n2787), .Z(n2789) );
  NANDN U2774 ( .A(n211), .B(n210), .Z(n215) );
  NAND U2775 ( .A(n213), .B(n212), .Z(n214) );
  AND U2776 ( .A(n215), .B(n214), .Z(n2788) );
  XOR U2777 ( .A(n2789), .B(n2788), .Z(n3286) );
  NANDN U2778 ( .A(n217), .B(n216), .Z(n221) );
  NANDN U2779 ( .A(n219), .B(n218), .Z(n220) );
  AND U2780 ( .A(n221), .B(n220), .Z(n3285) );
  XNOR U2781 ( .A(n3286), .B(n3285), .Z(n3287) );
  XNOR U2782 ( .A(n3288), .B(n3287), .Z(n2888) );
  XOR U2783 ( .A(n2889), .B(n2888), .Z(n2891) );
  NANDN U2784 ( .A(n222), .B(oglobal[0]), .Z(n226) );
  NANDN U2785 ( .A(n224), .B(n223), .Z(n225) );
  AND U2786 ( .A(n226), .B(n225), .Z(n2972) );
  NANDN U2787 ( .A(n228), .B(n227), .Z(n232) );
  NAND U2788 ( .A(n230), .B(n229), .Z(n231) );
  NAND U2789 ( .A(n232), .B(n231), .Z(n2973) );
  XNOR U2790 ( .A(n2972), .B(n2973), .Z(n2975) );
  NANDN U2791 ( .A(n234), .B(n233), .Z(n238) );
  NAND U2792 ( .A(n236), .B(n235), .Z(n237) );
  AND U2793 ( .A(n238), .B(n237), .Z(n2974) );
  XOR U2794 ( .A(n2975), .B(n2974), .Z(n3282) );
  NANDN U2795 ( .A(n240), .B(n239), .Z(n244) );
  NAND U2796 ( .A(n242), .B(n241), .Z(n243) );
  AND U2797 ( .A(n244), .B(n243), .Z(n2993) );
  NANDN U2798 ( .A(n246), .B(n245), .Z(n250) );
  NANDN U2799 ( .A(n248), .B(n247), .Z(n249) );
  NAND U2800 ( .A(n250), .B(n249), .Z(n2994) );
  XNOR U2801 ( .A(n2993), .B(n2994), .Z(n2996) );
  NANDN U2802 ( .A(n252), .B(n251), .Z(n256) );
  NANDN U2803 ( .A(n254), .B(n253), .Z(n255) );
  AND U2804 ( .A(n256), .B(n255), .Z(n2995) );
  XOR U2805 ( .A(n2996), .B(n2995), .Z(n3280) );
  NANDN U2806 ( .A(n258), .B(n257), .Z(n262) );
  NANDN U2807 ( .A(n260), .B(n259), .Z(n261) );
  AND U2808 ( .A(n262), .B(n261), .Z(n3279) );
  XNOR U2809 ( .A(n3280), .B(n3279), .Z(n3281) );
  XNOR U2810 ( .A(n3282), .B(n3281), .Z(n2890) );
  XOR U2811 ( .A(n2891), .B(n2890), .Z(n2545) );
  NANDN U2812 ( .A(n264), .B(n263), .Z(n268) );
  OR U2813 ( .A(n266), .B(n265), .Z(n267) );
  AND U2814 ( .A(n268), .B(n267), .Z(n2544) );
  XNOR U2815 ( .A(n2545), .B(n2544), .Z(n2546) );
  XNOR U2816 ( .A(n2547), .B(n2546), .Z(n3088) );
  NANDN U2817 ( .A(n270), .B(n269), .Z(n274) );
  NANDN U2818 ( .A(n272), .B(n271), .Z(n273) );
  AND U2819 ( .A(n274), .B(n273), .Z(n2571) );
  NANDN U2820 ( .A(n276), .B(n275), .Z(n280) );
  NAND U2821 ( .A(n278), .B(n277), .Z(n279) );
  NAND U2822 ( .A(n280), .B(n279), .Z(n3545) );
  NANDN U2823 ( .A(n282), .B(n281), .Z(n286) );
  NAND U2824 ( .A(n284), .B(n283), .Z(n285) );
  NAND U2825 ( .A(n286), .B(n285), .Z(n3544) );
  NANDN U2826 ( .A(n288), .B(n287), .Z(n292) );
  NAND U2827 ( .A(n290), .B(n289), .Z(n291) );
  AND U2828 ( .A(n292), .B(n291), .Z(n3543) );
  XOR U2829 ( .A(n3544), .B(n3543), .Z(n293) );
  XNOR U2830 ( .A(n3545), .B(n293), .Z(n2568) );
  NANDN U2831 ( .A(n295), .B(n294), .Z(n299) );
  NANDN U2832 ( .A(n297), .B(n296), .Z(n298) );
  NAND U2833 ( .A(n299), .B(n298), .Z(n2569) );
  XNOR U2834 ( .A(n2568), .B(n2569), .Z(n2570) );
  XOR U2835 ( .A(n2571), .B(n2570), .Z(n3210) );
  NANDN U2836 ( .A(n301), .B(n300), .Z(n305) );
  OR U2837 ( .A(n303), .B(n302), .Z(n304) );
  AND U2838 ( .A(n305), .B(n304), .Z(n3477) );
  NANDN U2839 ( .A(n311), .B(n310), .Z(n315) );
  NAND U2840 ( .A(n313), .B(n312), .Z(n314) );
  AND U2841 ( .A(n315), .B(n314), .Z(n3534) );
  NANDN U2842 ( .A(n317), .B(n316), .Z(n321) );
  NAND U2843 ( .A(n319), .B(n318), .Z(n320) );
  NAND U2844 ( .A(n321), .B(n320), .Z(n3535) );
  XNOR U2845 ( .A(n3534), .B(n3535), .Z(n3537) );
  NANDN U2846 ( .A(n323), .B(n322), .Z(n327) );
  NAND U2847 ( .A(n325), .B(n324), .Z(n326) );
  AND U2848 ( .A(n327), .B(n326), .Z(n3536) );
  XNOR U2849 ( .A(n3537), .B(n3536), .Z(n3474) );
  XOR U2850 ( .A(n3477), .B(n3476), .Z(n3208) );
  NAND U2851 ( .A(n329), .B(n328), .Z(n333) );
  NAND U2852 ( .A(n331), .B(n330), .Z(n332) );
  AND U2853 ( .A(n333), .B(n332), .Z(n3483) );
  NANDN U2854 ( .A(n335), .B(n334), .Z(n339) );
  NAND U2855 ( .A(n337), .B(n336), .Z(n338) );
  AND U2856 ( .A(n339), .B(n338), .Z(n2635) );
  NANDN U2857 ( .A(n341), .B(n340), .Z(n345) );
  NAND U2858 ( .A(n343), .B(n342), .Z(n344) );
  AND U2859 ( .A(n345), .B(n344), .Z(n2636) );
  NANDN U2860 ( .A(n347), .B(n346), .Z(n351) );
  NAND U2861 ( .A(n349), .B(n348), .Z(n350) );
  AND U2862 ( .A(n351), .B(n350), .Z(n2637) );
  XNOR U2863 ( .A(n2638), .B(n2637), .Z(n3481) );
  NAND U2864 ( .A(n353), .B(n352), .Z(n357) );
  NAND U2865 ( .A(n355), .B(n354), .Z(n356) );
  AND U2866 ( .A(n357), .B(n356), .Z(n3480) );
  XNOR U2867 ( .A(n3483), .B(n3482), .Z(n3207) );
  XNOR U2868 ( .A(n3208), .B(n3207), .Z(n3209) );
  XNOR U2869 ( .A(n3210), .B(n3209), .Z(n3072) );
  NANDN U2870 ( .A(n359), .B(n358), .Z(n363) );
  NANDN U2871 ( .A(n361), .B(n360), .Z(n362) );
  AND U2872 ( .A(n363), .B(n362), .Z(n3452) );
  NAND U2873 ( .A(n369), .B(n368), .Z(n373) );
  NAND U2874 ( .A(n371), .B(n370), .Z(n372) );
  NAND U2875 ( .A(n373), .B(n372), .Z(n2824) );
  NANDN U2876 ( .A(n375), .B(n374), .Z(n379) );
  NANDN U2877 ( .A(n377), .B(n376), .Z(n378) );
  NAND U2878 ( .A(n379), .B(n378), .Z(n2823) );
  NANDN U2879 ( .A(n381), .B(n380), .Z(n385) );
  NAND U2880 ( .A(n383), .B(n382), .Z(n384) );
  AND U2881 ( .A(n385), .B(n384), .Z(n2822) );
  XOR U2882 ( .A(n2823), .B(n2822), .Z(n386) );
  XNOR U2883 ( .A(n2824), .B(n386), .Z(n3449) );
  XOR U2884 ( .A(n3452), .B(n3451), .Z(n3192) );
  NAND U2885 ( .A(n388), .B(n387), .Z(n392) );
  NAND U2886 ( .A(n390), .B(n389), .Z(n391) );
  NAND U2887 ( .A(n392), .B(n391), .Z(n3458) );
  NANDN U2888 ( .A(n394), .B(n393), .Z(n398) );
  NAND U2889 ( .A(n396), .B(n395), .Z(n397) );
  AND U2890 ( .A(n398), .B(n397), .Z(n2840) );
  NANDN U2891 ( .A(n400), .B(n399), .Z(n404) );
  NAND U2892 ( .A(n402), .B(n401), .Z(n403) );
  NAND U2893 ( .A(n404), .B(n403), .Z(n2841) );
  XNOR U2894 ( .A(n2840), .B(n2841), .Z(n2843) );
  NANDN U2895 ( .A(n406), .B(n405), .Z(n410) );
  NAND U2896 ( .A(n408), .B(n407), .Z(n409) );
  AND U2897 ( .A(n410), .B(n409), .Z(n2842) );
  XNOR U2898 ( .A(n2843), .B(n2842), .Z(n3456) );
  NAND U2899 ( .A(n412), .B(n411), .Z(n416) );
  NAND U2900 ( .A(n414), .B(n413), .Z(n415) );
  NAND U2901 ( .A(n416), .B(n415), .Z(n3455) );
  NANDN U2902 ( .A(n422), .B(n421), .Z(n426) );
  NANDN U2903 ( .A(n424), .B(n423), .Z(n425) );
  AND U2904 ( .A(n426), .B(n425), .Z(n2816) );
  NANDN U2905 ( .A(n428), .B(n427), .Z(n432) );
  NAND U2906 ( .A(n430), .B(n429), .Z(n431) );
  AND U2907 ( .A(n432), .B(n431), .Z(n2817) );
  NANDN U2908 ( .A(n434), .B(n433), .Z(n438) );
  NAND U2909 ( .A(n436), .B(n435), .Z(n437) );
  AND U2910 ( .A(n438), .B(n437), .Z(n2818) );
  XOR U2911 ( .A(n2819), .B(n2818), .Z(n3511) );
  NANDN U2912 ( .A(n440), .B(n439), .Z(n444) );
  NANDN U2913 ( .A(n442), .B(n441), .Z(n443) );
  AND U2914 ( .A(n444), .B(n443), .Z(n3510) );
  XNOR U2915 ( .A(n3511), .B(n3510), .Z(n3512) );
  XNOR U2916 ( .A(n3513), .B(n3512), .Z(n3189) );
  XOR U2917 ( .A(n3190), .B(n3189), .Z(n3191) );
  XOR U2918 ( .A(n3192), .B(n3191), .Z(n3070) );
  NANDN U2919 ( .A(n446), .B(n445), .Z(n450) );
  NANDN U2920 ( .A(n448), .B(n447), .Z(n449) );
  AND U2921 ( .A(n450), .B(n449), .Z(n2577) );
  NANDN U2922 ( .A(n452), .B(n451), .Z(n456) );
  NAND U2923 ( .A(n454), .B(n453), .Z(n455) );
  AND U2924 ( .A(n456), .B(n455), .Z(n3523) );
  NAND U2925 ( .A(n458), .B(n457), .Z(n462) );
  NAND U2926 ( .A(n460), .B(n459), .Z(n461) );
  AND U2927 ( .A(n462), .B(n461), .Z(n3522) );
  XOR U2928 ( .A(n3523), .B(n3522), .Z(n3525) );
  NANDN U2929 ( .A(n464), .B(n463), .Z(n468) );
  NAND U2930 ( .A(n466), .B(n465), .Z(n467) );
  AND U2931 ( .A(n468), .B(n467), .Z(n3524) );
  XOR U2932 ( .A(n3525), .B(n3524), .Z(n2575) );
  NANDN U2933 ( .A(n470), .B(n469), .Z(n474) );
  NANDN U2934 ( .A(n472), .B(n471), .Z(n473) );
  AND U2935 ( .A(n474), .B(n473), .Z(n2574) );
  XNOR U2936 ( .A(n2575), .B(n2574), .Z(n2576) );
  XOR U2937 ( .A(n2577), .B(n2576), .Z(n3142) );
  NANDN U2938 ( .A(n476), .B(n475), .Z(n480) );
  NANDN U2939 ( .A(n478), .B(n477), .Z(n479) );
  AND U2940 ( .A(n480), .B(n479), .Z(n3501) );
  NANDN U2941 ( .A(n486), .B(n485), .Z(n490) );
  NAND U2942 ( .A(n488), .B(n487), .Z(n489) );
  AND U2943 ( .A(n490), .B(n489), .Z(n2804) );
  NANDN U2944 ( .A(n492), .B(n491), .Z(n496) );
  NAND U2945 ( .A(n494), .B(n493), .Z(n495) );
  AND U2946 ( .A(n496), .B(n495), .Z(n2805) );
  NANDN U2947 ( .A(n498), .B(n497), .Z(n502) );
  NAND U2948 ( .A(n500), .B(n499), .Z(n501) );
  AND U2949 ( .A(n502), .B(n501), .Z(n2806) );
  XNOR U2950 ( .A(n2807), .B(n2806), .Z(n3498) );
  XNOR U2951 ( .A(n3499), .B(n3498), .Z(n3500) );
  XOR U2952 ( .A(n3501), .B(n3500), .Z(n3141) );
  XOR U2953 ( .A(n3142), .B(n3141), .Z(n3144) );
  NAND U2954 ( .A(n504), .B(n503), .Z(n508) );
  NAND U2955 ( .A(n506), .B(n505), .Z(n507) );
  NAND U2956 ( .A(n508), .B(n507), .Z(n3464) );
  NAND U2957 ( .A(n510), .B(n509), .Z(n514) );
  NAND U2958 ( .A(n512), .B(n511), .Z(n513) );
  AND U2959 ( .A(n514), .B(n513), .Z(n2834) );
  NANDN U2960 ( .A(n516), .B(n515), .Z(n520) );
  NAND U2961 ( .A(n518), .B(n517), .Z(n519) );
  NAND U2962 ( .A(n520), .B(n519), .Z(n2835) );
  XNOR U2963 ( .A(n2834), .B(n2835), .Z(n2837) );
  NANDN U2964 ( .A(n522), .B(n521), .Z(n526) );
  NAND U2965 ( .A(n524), .B(n523), .Z(n525) );
  AND U2966 ( .A(n526), .B(n525), .Z(n2836) );
  XNOR U2967 ( .A(n2837), .B(n2836), .Z(n3462) );
  NANDN U2968 ( .A(n528), .B(n527), .Z(n532) );
  NANDN U2969 ( .A(n530), .B(n529), .Z(n531) );
  AND U2970 ( .A(n532), .B(n531), .Z(n3461) );
  XNOR U2971 ( .A(n3144), .B(n3143), .Z(n3069) );
  XNOR U2972 ( .A(n3070), .B(n3069), .Z(n3071) );
  XOR U2973 ( .A(n3072), .B(n3071), .Z(n3087) );
  XOR U2974 ( .A(n3088), .B(n3087), .Z(n3090) );
  NAND U2975 ( .A(n538), .B(n537), .Z(n542) );
  NAND U2976 ( .A(n540), .B(n539), .Z(n541) );
  AND U2977 ( .A(n542), .B(n541), .Z(n3166) );
  NANDN U2978 ( .A(n544), .B(n543), .Z(n548) );
  NANDN U2979 ( .A(n546), .B(n545), .Z(n547) );
  AND U2980 ( .A(n548), .B(n547), .Z(n2927) );
  NAND U2981 ( .A(n550), .B(n549), .Z(n554) );
  NAND U2982 ( .A(n552), .B(n551), .Z(n553) );
  AND U2983 ( .A(n554), .B(n553), .Z(n2604) );
  NANDN U2984 ( .A(n556), .B(n555), .Z(n560) );
  NAND U2985 ( .A(n558), .B(n557), .Z(n559) );
  NAND U2986 ( .A(n560), .B(n559), .Z(n2605) );
  XNOR U2987 ( .A(n2604), .B(n2605), .Z(n2607) );
  NAND U2988 ( .A(n562), .B(n561), .Z(n566) );
  NAND U2989 ( .A(n564), .B(n563), .Z(n565) );
  AND U2990 ( .A(n566), .B(n565), .Z(n2606) );
  XNOR U2991 ( .A(n2607), .B(n2606), .Z(n2925) );
  NANDN U2992 ( .A(n568), .B(n567), .Z(n572) );
  NANDN U2993 ( .A(n570), .B(n569), .Z(n571) );
  AND U2994 ( .A(n572), .B(n571), .Z(n2924) );
  XOR U2995 ( .A(n2927), .B(n2926), .Z(n3165) );
  XOR U2996 ( .A(n3166), .B(n3165), .Z(n3168) );
  NAND U2997 ( .A(n582), .B(n581), .Z(n586) );
  NAND U2998 ( .A(n584), .B(n583), .Z(n585) );
  AND U2999 ( .A(n586), .B(n585), .Z(n2580) );
  NAND U3000 ( .A(n588), .B(n587), .Z(n592) );
  NAND U3001 ( .A(n590), .B(n589), .Z(n591) );
  NAND U3002 ( .A(n592), .B(n591), .Z(n2581) );
  XNOR U3003 ( .A(n2580), .B(n2581), .Z(n2583) );
  NANDN U3004 ( .A(n594), .B(n593), .Z(n598) );
  NAND U3005 ( .A(n596), .B(n595), .Z(n597) );
  AND U3006 ( .A(n598), .B(n597), .Z(n2582) );
  XNOR U3007 ( .A(n2583), .B(n2582), .Z(n3486) );
  XOR U3008 ( .A(n3168), .B(n3167), .Z(n3082) );
  NAND U3009 ( .A(n604), .B(n603), .Z(n608) );
  NAND U3010 ( .A(n606), .B(n605), .Z(n607) );
  AND U3011 ( .A(n608), .B(n607), .Z(n3556) );
  NANDN U3012 ( .A(n610), .B(n609), .Z(n614) );
  NAND U3013 ( .A(n612), .B(n611), .Z(n613) );
  AND U3014 ( .A(n614), .B(n613), .Z(n3557) );
  NANDN U3015 ( .A(n616), .B(n615), .Z(n620) );
  NAND U3016 ( .A(n618), .B(n617), .Z(n619) );
  AND U3017 ( .A(n620), .B(n619), .Z(n3558) );
  XOR U3018 ( .A(n3559), .B(n3558), .Z(n3505) );
  NANDN U3019 ( .A(n622), .B(n621), .Z(n626) );
  OR U3020 ( .A(n624), .B(n623), .Z(n625) );
  AND U3021 ( .A(n626), .B(n625), .Z(n3504) );
  XNOR U3022 ( .A(n3505), .B(n3504), .Z(n3506) );
  XOR U3023 ( .A(n3507), .B(n3506), .Z(n3185) );
  NANDN U3024 ( .A(n628), .B(n627), .Z(n632) );
  NANDN U3025 ( .A(n630), .B(n629), .Z(n631) );
  AND U3026 ( .A(n632), .B(n631), .Z(n2565) );
  NAND U3027 ( .A(n634), .B(n633), .Z(n638) );
  NAND U3028 ( .A(n636), .B(n635), .Z(n637) );
  AND U3029 ( .A(n638), .B(n637), .Z(n2671) );
  NAND U3030 ( .A(n640), .B(n639), .Z(n644) );
  NAND U3031 ( .A(n642), .B(n641), .Z(n643) );
  AND U3032 ( .A(n644), .B(n643), .Z(n2672) );
  NAND U3033 ( .A(n646), .B(n645), .Z(n650) );
  NAND U3034 ( .A(n648), .B(n647), .Z(n649) );
  AND U3035 ( .A(n650), .B(n649), .Z(n2673) );
  XOR U3036 ( .A(n2674), .B(n2673), .Z(n2563) );
  NANDN U3037 ( .A(n652), .B(n651), .Z(n656) );
  NANDN U3038 ( .A(n654), .B(n653), .Z(n655) );
  AND U3039 ( .A(n656), .B(n655), .Z(n2562) );
  XNOR U3040 ( .A(n2563), .B(n2562), .Z(n2564) );
  XOR U3041 ( .A(n2565), .B(n2564), .Z(n3184) );
  NAND U3042 ( .A(n658), .B(n657), .Z(n662) );
  NAND U3043 ( .A(n660), .B(n659), .Z(n661) );
  NAND U3044 ( .A(n662), .B(n661), .Z(n3183) );
  XNOR U3045 ( .A(n3184), .B(n3183), .Z(n3186) );
  XOR U3046 ( .A(n3185), .B(n3186), .Z(n3081) );
  XNOR U3047 ( .A(n3082), .B(n3081), .Z(n3083) );
  XNOR U3048 ( .A(n3084), .B(n3083), .Z(n3089) );
  XOR U3049 ( .A(n3090), .B(n3089), .Z(n3120) );
  NANDN U3050 ( .A(n664), .B(n663), .Z(n668) );
  NANDN U3051 ( .A(n666), .B(n665), .Z(n667) );
  AND U3052 ( .A(n668), .B(n667), .Z(n3434) );
  NANDN U3053 ( .A(n670), .B(n669), .Z(n674) );
  NANDN U3054 ( .A(n672), .B(n671), .Z(n673) );
  AND U3055 ( .A(n674), .B(n673), .Z(n3431) );
  NANDN U3056 ( .A(n676), .B(n675), .Z(n680) );
  NANDN U3057 ( .A(n678), .B(n677), .Z(n679) );
  AND U3058 ( .A(n680), .B(n679), .Z(n3432) );
  XOR U3059 ( .A(n3434), .B(n3433), .Z(n2933) );
  NANDN U3060 ( .A(n682), .B(n681), .Z(n686) );
  NANDN U3061 ( .A(n684), .B(n683), .Z(n685) );
  AND U3062 ( .A(n686), .B(n685), .Z(n2931) );
  NANDN U3063 ( .A(n688), .B(n687), .Z(n692) );
  NANDN U3064 ( .A(n690), .B(n689), .Z(n691) );
  NAND U3065 ( .A(n692), .B(n691), .Z(n2930) );
  XNOR U3066 ( .A(n2931), .B(n2930), .Z(n2932) );
  XOR U3067 ( .A(n2933), .B(n2932), .Z(n3299) );
  NANDN U3068 ( .A(n698), .B(n697), .Z(n702) );
  NANDN U3069 ( .A(n700), .B(n699), .Z(n701) );
  AND U3070 ( .A(n702), .B(n701), .Z(n3422) );
  NAND U3071 ( .A(n704), .B(n703), .Z(n708) );
  NAND U3072 ( .A(n706), .B(n705), .Z(n707) );
  AND U3073 ( .A(n708), .B(n707), .Z(n3420) );
  NANDN U3074 ( .A(n710), .B(n709), .Z(n714) );
  NANDN U3075 ( .A(n712), .B(n711), .Z(n713) );
  AND U3076 ( .A(n714), .B(n713), .Z(n3419) );
  XNOR U3077 ( .A(n3420), .B(n3419), .Z(n3421) );
  XOR U3078 ( .A(n3422), .B(n3421), .Z(n3297) );
  XOR U3079 ( .A(n3298), .B(n3297), .Z(n3300) );
  XOR U3080 ( .A(n3299), .B(n3300), .Z(n3096) );
  NAND U3081 ( .A(n716), .B(n715), .Z(n720) );
  NAND U3082 ( .A(n718), .B(n717), .Z(n719) );
  AND U3083 ( .A(n720), .B(n719), .Z(n2858) );
  NANDN U3084 ( .A(n722), .B(n721), .Z(n726) );
  NAND U3085 ( .A(n724), .B(n723), .Z(n725) );
  AND U3086 ( .A(n726), .B(n725), .Z(n2859) );
  NANDN U3087 ( .A(n728), .B(n727), .Z(n732) );
  NAND U3088 ( .A(n730), .B(n729), .Z(n731) );
  AND U3089 ( .A(n732), .B(n731), .Z(n2860) );
  XOR U3090 ( .A(n2861), .B(n2860), .Z(n3252) );
  NANDN U3091 ( .A(n734), .B(n733), .Z(n738) );
  NAND U3092 ( .A(n736), .B(n735), .Z(n737) );
  AND U3093 ( .A(n738), .B(n737), .Z(n2987) );
  NANDN U3094 ( .A(n740), .B(n739), .Z(n744) );
  NAND U3095 ( .A(n742), .B(n741), .Z(n743) );
  NAND U3096 ( .A(n744), .B(n743), .Z(n2988) );
  XNOR U3097 ( .A(n2987), .B(n2988), .Z(n2990) );
  NANDN U3098 ( .A(n746), .B(n745), .Z(n750) );
  NAND U3099 ( .A(n748), .B(n747), .Z(n749) );
  AND U3100 ( .A(n750), .B(n749), .Z(n2989) );
  XOR U3101 ( .A(n2990), .B(n2989), .Z(n3250) );
  NANDN U3102 ( .A(n752), .B(n751), .Z(n756) );
  NANDN U3103 ( .A(n754), .B(n753), .Z(n755) );
  AND U3104 ( .A(n756), .B(n755), .Z(n3249) );
  XNOR U3105 ( .A(n3250), .B(n3249), .Z(n3251) );
  XOR U3106 ( .A(n3252), .B(n3251), .Z(n3470) );
  NANDN U3107 ( .A(n758), .B(n757), .Z(n762) );
  NAND U3108 ( .A(n760), .B(n759), .Z(n761) );
  AND U3109 ( .A(n762), .B(n761), .Z(n3598) );
  NANDN U3110 ( .A(n764), .B(n763), .Z(n768) );
  NAND U3111 ( .A(n766), .B(n765), .Z(n767) );
  NAND U3112 ( .A(n768), .B(n767), .Z(n3599) );
  XNOR U3113 ( .A(n3598), .B(n3599), .Z(n3601) );
  NANDN U3114 ( .A(n770), .B(n769), .Z(n774) );
  NAND U3115 ( .A(n772), .B(n771), .Z(n773) );
  AND U3116 ( .A(n774), .B(n773), .Z(n3600) );
  XOR U3117 ( .A(n3601), .B(n3600), .Z(n3264) );
  NANDN U3118 ( .A(n776), .B(n775), .Z(n780) );
  NANDN U3119 ( .A(n778), .B(n777), .Z(n779) );
  AND U3120 ( .A(n780), .B(n779), .Z(n3262) );
  NANDN U3121 ( .A(n782), .B(n781), .Z(n786) );
  NANDN U3122 ( .A(n784), .B(n783), .Z(n785) );
  AND U3123 ( .A(n786), .B(n785), .Z(n3664) );
  NANDN U3124 ( .A(n788), .B(n787), .Z(n792) );
  NANDN U3125 ( .A(n790), .B(n789), .Z(n791) );
  AND U3126 ( .A(n792), .B(n791), .Z(n3662) );
  XNOR U3127 ( .A(n3662), .B(oglobal[1]), .Z(n3663) );
  XNOR U3128 ( .A(n3664), .B(n3663), .Z(n3261) );
  XOR U3129 ( .A(n3262), .B(n3261), .Z(n3263) );
  XOR U3130 ( .A(n3264), .B(n3263), .Z(n3469) );
  NANDN U3131 ( .A(n794), .B(n793), .Z(n798) );
  NANDN U3132 ( .A(n796), .B(n795), .Z(n797) );
  NAND U3133 ( .A(n798), .B(n797), .Z(n2980) );
  NANDN U3134 ( .A(n800), .B(n799), .Z(n804) );
  NAND U3135 ( .A(n802), .B(n801), .Z(n803) );
  NAND U3136 ( .A(n804), .B(n803), .Z(n2979) );
  NANDN U3137 ( .A(n806), .B(n805), .Z(n810) );
  NANDN U3138 ( .A(n808), .B(n807), .Z(n809) );
  AND U3139 ( .A(n810), .B(n809), .Z(n2978) );
  XOR U3140 ( .A(n2979), .B(n2978), .Z(n811) );
  XOR U3141 ( .A(n2980), .B(n811), .Z(n3270) );
  NANDN U3142 ( .A(n813), .B(n812), .Z(n817) );
  NANDN U3143 ( .A(n815), .B(n814), .Z(n816) );
  NAND U3144 ( .A(n817), .B(n816), .Z(n3628) );
  NANDN U3145 ( .A(n819), .B(n818), .Z(n823) );
  NAND U3146 ( .A(n821), .B(n820), .Z(n822) );
  AND U3147 ( .A(n823), .B(n822), .Z(n3630) );
  NANDN U3148 ( .A(n825), .B(n824), .Z(n829) );
  NAND U3149 ( .A(n827), .B(n826), .Z(n828) );
  AND U3150 ( .A(n829), .B(n828), .Z(n3629) );
  XNOR U3151 ( .A(n3630), .B(n3629), .Z(n830) );
  XNOR U3152 ( .A(n3628), .B(n830), .Z(n3267) );
  NANDN U3153 ( .A(n832), .B(n831), .Z(n836) );
  NANDN U3154 ( .A(n834), .B(n833), .Z(n835) );
  AND U3155 ( .A(n836), .B(n835), .Z(n3268) );
  XOR U3156 ( .A(n3267), .B(n3268), .Z(n3269) );
  XOR U3157 ( .A(n3270), .B(n3269), .Z(n3468) );
  XOR U3158 ( .A(n3469), .B(n3468), .Z(n3471) );
  XNOR U3159 ( .A(n3470), .B(n3471), .Z(n3094) );
  NANDN U3160 ( .A(n838), .B(n837), .Z(n842) );
  NAND U3161 ( .A(n840), .B(n839), .Z(n841) );
  AND U3162 ( .A(n842), .B(n841), .Z(n2553) );
  NANDN U3163 ( .A(n844), .B(n843), .Z(n848) );
  NANDN U3164 ( .A(n846), .B(n845), .Z(n847) );
  AND U3165 ( .A(n848), .B(n847), .Z(n3352) );
  NANDN U3166 ( .A(n850), .B(n849), .Z(n854) );
  NAND U3167 ( .A(n852), .B(n851), .Z(n853) );
  AND U3168 ( .A(n854), .B(n853), .Z(n2870) );
  NAND U3169 ( .A(n856), .B(n855), .Z(n860) );
  NAND U3170 ( .A(n858), .B(n857), .Z(n859) );
  AND U3171 ( .A(n860), .B(n859), .Z(n2871) );
  NAND U3172 ( .A(n862), .B(n861), .Z(n866) );
  NAND U3173 ( .A(n864), .B(n863), .Z(n865) );
  AND U3174 ( .A(n866), .B(n865), .Z(n2873) );
  NANDN U3175 ( .A(n868), .B(n867), .Z(n872) );
  NAND U3176 ( .A(n870), .B(n869), .Z(n871) );
  AND U3177 ( .A(n872), .B(n871), .Z(n3610) );
  NANDN U3178 ( .A(n874), .B(n873), .Z(n878) );
  NAND U3179 ( .A(n876), .B(n875), .Z(n877) );
  NAND U3180 ( .A(n878), .B(n877), .Z(n3611) );
  XNOR U3181 ( .A(n3610), .B(n3611), .Z(n3612) );
  NANDN U3182 ( .A(n880), .B(n879), .Z(n884) );
  NAND U3183 ( .A(n882), .B(n881), .Z(n883) );
  NAND U3184 ( .A(n884), .B(n883), .Z(n3613) );
  XNOR U3185 ( .A(n3612), .B(n3613), .Z(n3353) );
  XNOR U3186 ( .A(n3354), .B(n3353), .Z(n885) );
  XOR U3187 ( .A(n3352), .B(n885), .Z(n2551) );
  NANDN U3188 ( .A(n887), .B(n886), .Z(n891) );
  NAND U3189 ( .A(n889), .B(n888), .Z(n890) );
  AND U3190 ( .A(n891), .B(n890), .Z(n2756) );
  NAND U3191 ( .A(n893), .B(n892), .Z(n897) );
  NAND U3192 ( .A(n895), .B(n894), .Z(n896) );
  AND U3193 ( .A(n897), .B(n896), .Z(n2757) );
  NAND U3194 ( .A(n899), .B(n898), .Z(n903) );
  NAND U3195 ( .A(n901), .B(n900), .Z(n902) );
  AND U3196 ( .A(n903), .B(n902), .Z(n2758) );
  XOR U3197 ( .A(n2759), .B(n2758), .Z(n3246) );
  NANDN U3198 ( .A(n905), .B(n904), .Z(n909) );
  NAND U3199 ( .A(n907), .B(n906), .Z(n908) );
  NAND U3200 ( .A(n909), .B(n908), .Z(n3631) );
  NANDN U3201 ( .A(n911), .B(n910), .Z(n915) );
  NAND U3202 ( .A(n913), .B(n912), .Z(n914) );
  AND U3203 ( .A(n915), .B(n914), .Z(n3633) );
  NANDN U3204 ( .A(n917), .B(n916), .Z(n921) );
  NAND U3205 ( .A(n919), .B(n918), .Z(n920) );
  AND U3206 ( .A(n921), .B(n920), .Z(n3632) );
  XNOR U3207 ( .A(n3633), .B(n3632), .Z(n922) );
  XNOR U3208 ( .A(n3631), .B(n922), .Z(n3243) );
  NANDN U3209 ( .A(n924), .B(n923), .Z(n928) );
  NANDN U3210 ( .A(n926), .B(n925), .Z(n927) );
  AND U3211 ( .A(n928), .B(n927), .Z(n3244) );
  XOR U3212 ( .A(n3243), .B(n3244), .Z(n3245) );
  XOR U3213 ( .A(n3246), .B(n3245), .Z(n2550) );
  XOR U3214 ( .A(n2551), .B(n2550), .Z(n2552) );
  XOR U3215 ( .A(n2553), .B(n2552), .Z(n3093) );
  XOR U3216 ( .A(n3094), .B(n3093), .Z(n3095) );
  XOR U3217 ( .A(n3096), .B(n3095), .Z(n3064) );
  NANDN U3218 ( .A(n938), .B(n937), .Z(n942) );
  NAND U3219 ( .A(n940), .B(n939), .Z(n941) );
  AND U3220 ( .A(n942), .B(n941), .Z(n3650) );
  NANDN U3221 ( .A(n944), .B(n943), .Z(n948) );
  NAND U3222 ( .A(n946), .B(n945), .Z(n947) );
  NAND U3223 ( .A(n948), .B(n947), .Z(n3651) );
  XNOR U3224 ( .A(n3650), .B(n3651), .Z(n3653) );
  NANDN U3225 ( .A(n950), .B(n949), .Z(n954) );
  NAND U3226 ( .A(n952), .B(n951), .Z(n953) );
  AND U3227 ( .A(n954), .B(n953), .Z(n3652) );
  XOR U3228 ( .A(n3653), .B(n3652), .Z(n3398) );
  NANDN U3229 ( .A(n956), .B(n955), .Z(n960) );
  NAND U3230 ( .A(n958), .B(n957), .Z(n959) );
  AND U3231 ( .A(n960), .B(n959), .Z(n2738) );
  NANDN U3232 ( .A(n962), .B(n961), .Z(n966) );
  NAND U3233 ( .A(n964), .B(n963), .Z(n965) );
  NAND U3234 ( .A(n966), .B(n965), .Z(n2739) );
  XNOR U3235 ( .A(n2738), .B(n2739), .Z(n2741) );
  NANDN U3236 ( .A(n968), .B(n967), .Z(n972) );
  NAND U3237 ( .A(n970), .B(n969), .Z(n971) );
  AND U3238 ( .A(n972), .B(n971), .Z(n2740) );
  XOR U3239 ( .A(n2741), .B(n2740), .Z(n3396) );
  NANDN U3240 ( .A(n974), .B(n973), .Z(n978) );
  NANDN U3241 ( .A(n976), .B(n975), .Z(n977) );
  AND U3242 ( .A(n978), .B(n977), .Z(n3395) );
  XNOR U3243 ( .A(n3396), .B(n3395), .Z(n3397) );
  XOR U3244 ( .A(n3398), .B(n3397), .Z(n3680) );
  NAND U3245 ( .A(n980), .B(n979), .Z(n984) );
  NAND U3246 ( .A(n982), .B(n981), .Z(n983) );
  NAND U3247 ( .A(n984), .B(n983), .Z(n3679) );
  XOR U3248 ( .A(n3680), .B(n3679), .Z(n3681) );
  XNOR U3249 ( .A(n3682), .B(n3681), .Z(n3099) );
  XNOR U3250 ( .A(n3100), .B(n3099), .Z(n3102) );
  NANDN U3251 ( .A(n986), .B(n985), .Z(n990) );
  NANDN U3252 ( .A(n988), .B(n987), .Z(n989) );
  AND U3253 ( .A(n990), .B(n989), .Z(n3670) );
  NANDN U3254 ( .A(n992), .B(n991), .Z(n996) );
  NANDN U3255 ( .A(n994), .B(n993), .Z(n995) );
  AND U3256 ( .A(n996), .B(n995), .Z(n3416) );
  NANDN U3257 ( .A(n998), .B(n997), .Z(n1002) );
  NANDN U3258 ( .A(n1000), .B(n999), .Z(n1001) );
  AND U3259 ( .A(n1002), .B(n1001), .Z(n3413) );
  NANDN U3260 ( .A(n1004), .B(n1003), .Z(n1008) );
  NANDN U3261 ( .A(n1006), .B(n1005), .Z(n1007) );
  NAND U3262 ( .A(n1008), .B(n1007), .Z(n3414) );
  XNOR U3263 ( .A(n3413), .B(n3414), .Z(n3415) );
  XOR U3264 ( .A(n3416), .B(n3415), .Z(n3668) );
  NANDN U3265 ( .A(n1010), .B(n1009), .Z(n1014) );
  NANDN U3266 ( .A(n1012), .B(n1011), .Z(n1013) );
  AND U3267 ( .A(n1014), .B(n1013), .Z(n3440) );
  NANDN U3268 ( .A(n1016), .B(n1015), .Z(n1020) );
  NANDN U3269 ( .A(n1018), .B(n1017), .Z(n1019) );
  AND U3270 ( .A(n1020), .B(n1019), .Z(n3437) );
  NANDN U3271 ( .A(n1022), .B(n1021), .Z(n1026) );
  NANDN U3272 ( .A(n1024), .B(n1023), .Z(n1025) );
  NAND U3273 ( .A(n1026), .B(n1025), .Z(n3438) );
  XNOR U3274 ( .A(n3437), .B(n3438), .Z(n3439) );
  XNOR U3275 ( .A(n3440), .B(n3439), .Z(n3667) );
  XNOR U3276 ( .A(n3668), .B(n3667), .Z(n3669) );
  XOR U3277 ( .A(n3670), .B(n3669), .Z(n3101) );
  XOR U3278 ( .A(n3102), .B(n3101), .Z(n3063) );
  XNOR U3279 ( .A(n3064), .B(n3063), .Z(n3066) );
  NANDN U3280 ( .A(n1028), .B(n1027), .Z(n1032) );
  NAND U3281 ( .A(n1030), .B(n1029), .Z(n1031) );
  AND U3282 ( .A(n1032), .B(n1031), .Z(n2750) );
  NANDN U3283 ( .A(n1034), .B(n1033), .Z(n1038) );
  NAND U3284 ( .A(n1036), .B(n1035), .Z(n1037) );
  AND U3285 ( .A(n1038), .B(n1037), .Z(n2751) );
  NANDN U3286 ( .A(n1040), .B(n1039), .Z(n1044) );
  NAND U3287 ( .A(n1042), .B(n1041), .Z(n1043) );
  AND U3288 ( .A(n1044), .B(n1043), .Z(n2752) );
  XNOR U3289 ( .A(n2753), .B(n2752), .Z(n3349) );
  NANDN U3290 ( .A(n1046), .B(n1045), .Z(n1050) );
  NAND U3291 ( .A(n1048), .B(n1047), .Z(n1049) );
  AND U3292 ( .A(n1050), .B(n1049), .Z(n2716) );
  NANDN U3293 ( .A(n1052), .B(n1051), .Z(n1056) );
  NAND U3294 ( .A(n1054), .B(n1053), .Z(n1055) );
  AND U3295 ( .A(n1056), .B(n1055), .Z(n2717) );
  NANDN U3296 ( .A(n1058), .B(n1057), .Z(n1062) );
  NAND U3297 ( .A(n1060), .B(n1059), .Z(n1061) );
  AND U3298 ( .A(n1062), .B(n1061), .Z(n2718) );
  XNOR U3299 ( .A(n2719), .B(n2718), .Z(n3347) );
  NANDN U3300 ( .A(n1064), .B(n1063), .Z(n1068) );
  NANDN U3301 ( .A(n1066), .B(n1065), .Z(n1067) );
  AND U3302 ( .A(n1068), .B(n1067), .Z(n3346) );
  NANDN U3303 ( .A(n1070), .B(n1069), .Z(n1074) );
  NAND U3304 ( .A(n1072), .B(n1071), .Z(n1073) );
  AND U3305 ( .A(n1074), .B(n1073), .Z(n3309) );
  NANDN U3306 ( .A(n1076), .B(n1075), .Z(n1080) );
  NAND U3307 ( .A(n1078), .B(n1077), .Z(n1079) );
  AND U3308 ( .A(n1080), .B(n1079), .Z(n3310) );
  NANDN U3309 ( .A(n1082), .B(n1081), .Z(n1086) );
  NAND U3310 ( .A(n1084), .B(n1083), .Z(n1085) );
  AND U3311 ( .A(n1086), .B(n1085), .Z(n3311) );
  XNOR U3312 ( .A(n3312), .B(n3311), .Z(n3386) );
  NANDN U3313 ( .A(n1092), .B(n1091), .Z(n1096) );
  NAND U3314 ( .A(n1094), .B(n1093), .Z(n1095) );
  AND U3315 ( .A(n1096), .B(n1095), .Z(n2629) );
  NANDN U3316 ( .A(n1098), .B(n1097), .Z(n1102) );
  NAND U3317 ( .A(n1100), .B(n1099), .Z(n1101) );
  AND U3318 ( .A(n1102), .B(n1101), .Z(n2630) );
  NANDN U3319 ( .A(n1104), .B(n1103), .Z(n1108) );
  NAND U3320 ( .A(n1106), .B(n1105), .Z(n1107) );
  AND U3321 ( .A(n1108), .B(n1107), .Z(n2631) );
  XNOR U3322 ( .A(n2632), .B(n2631), .Z(n3383) );
  XOR U3323 ( .A(n3517), .B(n3516), .Z(n3519) );
  NANDN U3324 ( .A(n1110), .B(n1109), .Z(n1114) );
  NAND U3325 ( .A(n1112), .B(n1111), .Z(n1113) );
  AND U3326 ( .A(n1114), .B(n1113), .Z(n2724) );
  NANDN U3327 ( .A(n1116), .B(n1115), .Z(n1120) );
  NAND U3328 ( .A(n1118), .B(n1117), .Z(n1119) );
  AND U3329 ( .A(n1120), .B(n1119), .Z(n2723) );
  NANDN U3330 ( .A(n1122), .B(n1121), .Z(n1126) );
  NAND U3331 ( .A(n1124), .B(n1123), .Z(n1125) );
  AND U3332 ( .A(n1126), .B(n1125), .Z(n2722) );
  NANDN U3333 ( .A(n1128), .B(n1127), .Z(n1132) );
  NAND U3334 ( .A(n1130), .B(n1129), .Z(n1131) );
  AND U3335 ( .A(n1132), .B(n1131), .Z(n3334) );
  NANDN U3336 ( .A(n1134), .B(n1133), .Z(n1138) );
  NAND U3337 ( .A(n1136), .B(n1135), .Z(n1137) );
  AND U3338 ( .A(n1138), .B(n1137), .Z(n3335) );
  NANDN U3339 ( .A(n1140), .B(n1139), .Z(n1144) );
  NAND U3340 ( .A(n1142), .B(n1141), .Z(n1143) );
  AND U3341 ( .A(n1144), .B(n1143), .Z(n3336) );
  XNOR U3342 ( .A(n3337), .B(n3336), .Z(n3378) );
  NANDN U3343 ( .A(n1146), .B(n1145), .Z(n1150) );
  NANDN U3344 ( .A(n1148), .B(n1147), .Z(n1149) );
  AND U3345 ( .A(n1150), .B(n1149), .Z(n3377) );
  XOR U3346 ( .A(n3379), .B(n3380), .Z(n3518) );
  XOR U3347 ( .A(n3519), .B(n3518), .Z(n3078) );
  NANDN U3348 ( .A(n1152), .B(n1151), .Z(n1156) );
  NAND U3349 ( .A(n1154), .B(n1153), .Z(n1155) );
  AND U3350 ( .A(n1156), .B(n1155), .Z(n3318) );
  NAND U3351 ( .A(n1158), .B(n1157), .Z(n1162) );
  NAND U3352 ( .A(n1160), .B(n1159), .Z(n1161) );
  AND U3353 ( .A(n1162), .B(n1161), .Z(n3320) );
  NANDN U3354 ( .A(n1164), .B(n1163), .Z(n1168) );
  NAND U3355 ( .A(n1166), .B(n1165), .Z(n1167) );
  AND U3356 ( .A(n1168), .B(n1167), .Z(n3319) );
  NANDN U3357 ( .A(n1170), .B(n1169), .Z(n1174) );
  NANDN U3358 ( .A(n1172), .B(n1171), .Z(n1173) );
  AND U3359 ( .A(n1174), .B(n1173), .Z(n3592) );
  NANDN U3360 ( .A(n1176), .B(n1175), .Z(n1180) );
  NANDN U3361 ( .A(n1178), .B(n1177), .Z(n1179) );
  NAND U3362 ( .A(n1180), .B(n1179), .Z(n3593) );
  XNOR U3363 ( .A(n3592), .B(n3593), .Z(n3595) );
  NANDN U3364 ( .A(n1182), .B(n1181), .Z(n1186) );
  NAND U3365 ( .A(n1184), .B(n1183), .Z(n1185) );
  AND U3366 ( .A(n1186), .B(n1185), .Z(n3594) );
  XNOR U3367 ( .A(n3595), .B(n3594), .Z(n3366) );
  NANDN U3368 ( .A(n1188), .B(n1187), .Z(n1192) );
  NANDN U3369 ( .A(n1190), .B(n1189), .Z(n1191) );
  AND U3370 ( .A(n1192), .B(n1191), .Z(n3365) );
  XOR U3371 ( .A(n3367), .B(n3368), .Z(n2557) );
  NANDN U3372 ( .A(n1194), .B(n1193), .Z(n1198) );
  NANDN U3373 ( .A(n1196), .B(n1195), .Z(n1197) );
  AND U3374 ( .A(n1198), .B(n1197), .Z(n3009) );
  NANDN U3375 ( .A(n1200), .B(n1199), .Z(n1204) );
  NANDN U3376 ( .A(n1202), .B(n1201), .Z(n1203) );
  AND U3377 ( .A(n1204), .B(n1203), .Z(n3010) );
  NANDN U3378 ( .A(n1206), .B(n1205), .Z(n1210) );
  NANDN U3379 ( .A(n1208), .B(n1207), .Z(n1209) );
  AND U3380 ( .A(n1210), .B(n1209), .Z(n3011) );
  XNOR U3381 ( .A(n3012), .B(n3011), .Z(n3362) );
  NANDN U3382 ( .A(n1212), .B(n1211), .Z(n1216) );
  NANDN U3383 ( .A(n1214), .B(n1213), .Z(n1215) );
  AND U3384 ( .A(n1216), .B(n1215), .Z(n3045) );
  NANDN U3385 ( .A(n1218), .B(n1217), .Z(n1222) );
  NANDN U3386 ( .A(n1220), .B(n1219), .Z(n1221) );
  AND U3387 ( .A(n1222), .B(n1221), .Z(n3046) );
  NANDN U3388 ( .A(n1224), .B(n1223), .Z(n1228) );
  NANDN U3389 ( .A(n1226), .B(n1225), .Z(n1227) );
  AND U3390 ( .A(n1228), .B(n1227), .Z(n3047) );
  XNOR U3391 ( .A(n3048), .B(n3047), .Z(n3360) );
  NANDN U3392 ( .A(n1230), .B(n1229), .Z(n1234) );
  NANDN U3393 ( .A(n1232), .B(n1231), .Z(n1233) );
  AND U3394 ( .A(n1234), .B(n1233), .Z(n3359) );
  XOR U3395 ( .A(n2557), .B(n2556), .Z(n2559) );
  NANDN U3396 ( .A(n1236), .B(n1235), .Z(n1240) );
  NAND U3397 ( .A(n1238), .B(n1237), .Z(n1239) );
  AND U3398 ( .A(n1240), .B(n1239), .Z(n3532) );
  NAND U3399 ( .A(n1242), .B(n1241), .Z(n1246) );
  NAND U3400 ( .A(n1244), .B(n1243), .Z(n1245) );
  AND U3401 ( .A(n1246), .B(n1245), .Z(n3533) );
  NANDN U3402 ( .A(n1248), .B(n1247), .Z(n1252) );
  NAND U3403 ( .A(n1250), .B(n1249), .Z(n1251) );
  NAND U3404 ( .A(n1252), .B(n1251), .Z(n3531) );
  XOR U3405 ( .A(n3533), .B(n3531), .Z(n1253) );
  XOR U3406 ( .A(n3532), .B(n1253), .Z(n2902) );
  NANDN U3407 ( .A(n1255), .B(n1254), .Z(n1259) );
  NAND U3408 ( .A(n1257), .B(n1256), .Z(n1258) );
  NAND U3409 ( .A(n1259), .B(n1258), .Z(n2901) );
  NANDN U3410 ( .A(n1261), .B(n1260), .Z(n1265) );
  NANDN U3411 ( .A(n1263), .B(n1262), .Z(n1264) );
  AND U3412 ( .A(n1265), .B(n1264), .Z(n2966) );
  NANDN U3413 ( .A(n1267), .B(n1266), .Z(n1271) );
  NANDN U3414 ( .A(n1269), .B(n1268), .Z(n1270) );
  NAND U3415 ( .A(n1271), .B(n1270), .Z(n2967) );
  XNOR U3416 ( .A(n2966), .B(n2967), .Z(n2969) );
  NANDN U3417 ( .A(n1273), .B(n1272), .Z(n1277) );
  NANDN U3418 ( .A(n1275), .B(n1274), .Z(n1276) );
  AND U3419 ( .A(n1277), .B(n1276), .Z(n2968) );
  XNOR U3420 ( .A(n2969), .B(n2968), .Z(n2900) );
  XOR U3421 ( .A(n2902), .B(n2903), .Z(n2558) );
  XOR U3422 ( .A(n2559), .B(n2558), .Z(n3076) );
  NANDN U3423 ( .A(n1279), .B(n1278), .Z(n1283) );
  NANDN U3424 ( .A(n1281), .B(n1280), .Z(n1282) );
  AND U3425 ( .A(n1283), .B(n1282), .Z(n2915) );
  NAND U3426 ( .A(n1285), .B(n1284), .Z(n1289) );
  NAND U3427 ( .A(n1287), .B(n1286), .Z(n1288) );
  AND U3428 ( .A(n1289), .B(n1288), .Z(n2913) );
  NANDN U3429 ( .A(n1291), .B(n1290), .Z(n1295) );
  NANDN U3430 ( .A(n1293), .B(n1292), .Z(n1294) );
  AND U3431 ( .A(n1295), .B(n1294), .Z(n2653) );
  NANDN U3432 ( .A(n1297), .B(n1296), .Z(n1301) );
  NAND U3433 ( .A(n1299), .B(n1298), .Z(n1300) );
  NAND U3434 ( .A(n1301), .B(n1300), .Z(n2654) );
  XNOR U3435 ( .A(n2653), .B(n2654), .Z(n2656) );
  NANDN U3436 ( .A(n1303), .B(n1302), .Z(n1307) );
  NANDN U3437 ( .A(n1305), .B(n1304), .Z(n1306) );
  AND U3438 ( .A(n1307), .B(n1306), .Z(n2655) );
  XNOR U3439 ( .A(n2656), .B(n2655), .Z(n2912) );
  XNOR U3440 ( .A(n2913), .B(n2912), .Z(n2914) );
  XOR U3441 ( .A(n2915), .B(n2914), .Z(n3228) );
  NANDN U3442 ( .A(n1309), .B(n1308), .Z(n1313) );
  NANDN U3443 ( .A(n1311), .B(n1310), .Z(n1312) );
  AND U3444 ( .A(n1313), .B(n1312), .Z(n2921) );
  NANDN U3445 ( .A(n1315), .B(n1314), .Z(n1319) );
  NANDN U3446 ( .A(n1317), .B(n1316), .Z(n1318) );
  AND U3447 ( .A(n1319), .B(n1318), .Z(n2647) );
  NAND U3448 ( .A(n1321), .B(n1320), .Z(n1325) );
  NAND U3449 ( .A(n1323), .B(n1322), .Z(n1324) );
  NAND U3450 ( .A(n1325), .B(n1324), .Z(n2648) );
  XNOR U3451 ( .A(n2647), .B(n2648), .Z(n2650) );
  NAND U3452 ( .A(n1327), .B(n1326), .Z(n1331) );
  NAND U3453 ( .A(n1329), .B(n1328), .Z(n1330) );
  AND U3454 ( .A(n1331), .B(n1330), .Z(n2649) );
  XOR U3455 ( .A(n2650), .B(n2649), .Z(n2919) );
  NANDN U3456 ( .A(n1333), .B(n1332), .Z(n1337) );
  NANDN U3457 ( .A(n1335), .B(n1334), .Z(n1336) );
  AND U3458 ( .A(n1337), .B(n1336), .Z(n2918) );
  XNOR U3459 ( .A(n2919), .B(n2918), .Z(n2920) );
  XOR U3460 ( .A(n2921), .B(n2920), .Z(n3226) );
  NANDN U3461 ( .A(n1339), .B(n1338), .Z(n1343) );
  NANDN U3462 ( .A(n1341), .B(n1340), .Z(n1342) );
  AND U3463 ( .A(n1343), .B(n1342), .Z(n3033) );
  NANDN U3464 ( .A(n1345), .B(n1344), .Z(n1349) );
  NANDN U3465 ( .A(n1347), .B(n1346), .Z(n1348) );
  NAND U3466 ( .A(n1349), .B(n1348), .Z(n3034) );
  XNOR U3467 ( .A(n3033), .B(n3034), .Z(n3036) );
  NANDN U3468 ( .A(n1351), .B(n1350), .Z(n1355) );
  NANDN U3469 ( .A(n1353), .B(n1352), .Z(n1354) );
  AND U3470 ( .A(n1355), .B(n1354), .Z(n3035) );
  XOR U3471 ( .A(n3036), .B(n3035), .Z(n2897) );
  NANDN U3472 ( .A(n1357), .B(n1356), .Z(n1361) );
  NANDN U3473 ( .A(n1359), .B(n1358), .Z(n1360) );
  AND U3474 ( .A(n1361), .B(n1360), .Z(n3015) );
  NAND U3475 ( .A(n1363), .B(n1362), .Z(n1367) );
  NAND U3476 ( .A(n1365), .B(n1364), .Z(n1366) );
  NAND U3477 ( .A(n1367), .B(n1366), .Z(n3016) );
  XNOR U3478 ( .A(n3015), .B(n3016), .Z(n3018) );
  NAND U3479 ( .A(n1369), .B(n1368), .Z(n1373) );
  NAND U3480 ( .A(n1371), .B(n1370), .Z(n1372) );
  AND U3481 ( .A(n1373), .B(n1372), .Z(n3017) );
  XOR U3482 ( .A(n3018), .B(n3017), .Z(n2895) );
  NANDN U3483 ( .A(n1375), .B(n1374), .Z(n1379) );
  NANDN U3484 ( .A(n1377), .B(n1376), .Z(n1378) );
  AND U3485 ( .A(n1379), .B(n1378), .Z(n2894) );
  XNOR U3486 ( .A(n2895), .B(n2894), .Z(n2896) );
  XOR U3487 ( .A(n2897), .B(n2896), .Z(n3225) );
  XNOR U3488 ( .A(n3226), .B(n3225), .Z(n3227) );
  XNOR U3489 ( .A(n3228), .B(n3227), .Z(n3075) );
  XNOR U3490 ( .A(n3076), .B(n3075), .Z(n3077) );
  XNOR U3491 ( .A(n3078), .B(n3077), .Z(n3065) );
  XOR U3492 ( .A(n3066), .B(n3065), .Z(n3118) );
  NANDN U3493 ( .A(n1385), .B(n1384), .Z(n1389) );
  NAND U3494 ( .A(n1387), .B(n1386), .Z(n1388) );
  AND U3495 ( .A(n1389), .B(n1388), .Z(n3676) );
  NANDN U3496 ( .A(n1391), .B(n1390), .Z(n1395) );
  NANDN U3497 ( .A(n1393), .B(n1392), .Z(n1394) );
  AND U3498 ( .A(n1395), .B(n1394), .Z(n3674) );
  NANDN U3499 ( .A(n1397), .B(n1396), .Z(n1401) );
  OR U3500 ( .A(n1399), .B(n1398), .Z(n1400) );
  AND U3501 ( .A(n1401), .B(n1400), .Z(n3673) );
  XOR U3502 ( .A(n3674), .B(n3673), .Z(n3675) );
  XOR U3503 ( .A(n3676), .B(n3675), .Z(n3495) );
  NANDN U3504 ( .A(n1403), .B(n1402), .Z(n1407) );
  NANDN U3505 ( .A(n1405), .B(n1404), .Z(n1406) );
  AND U3506 ( .A(n1407), .B(n1406), .Z(n3493) );
  NANDN U3507 ( .A(n1409), .B(n1408), .Z(n1413) );
  NANDN U3508 ( .A(n1411), .B(n1410), .Z(n1412) );
  NAND U3509 ( .A(n1413), .B(n1412), .Z(n3492) );
  XNOR U3510 ( .A(n3493), .B(n3492), .Z(n3494) );
  XNOR U3511 ( .A(n3495), .B(n3494), .Z(n2879) );
  NANDN U3512 ( .A(n1415), .B(n1414), .Z(n1419) );
  NANDN U3513 ( .A(n1417), .B(n1416), .Z(n1418) );
  AND U3514 ( .A(n1419), .B(n1418), .Z(n2877) );
  NANDN U3515 ( .A(n1421), .B(n1420), .Z(n1425) );
  NANDN U3516 ( .A(n1423), .B(n1422), .Z(n1424) );
  AND U3517 ( .A(n1425), .B(n1424), .Z(n3234) );
  NANDN U3518 ( .A(n1427), .B(n1426), .Z(n1431) );
  NAND U3519 ( .A(n1429), .B(n1428), .Z(n1430) );
  AND U3520 ( .A(n1431), .B(n1430), .Z(n3232) );
  NANDN U3521 ( .A(n1433), .B(n1432), .Z(n1437) );
  NAND U3522 ( .A(n1435), .B(n1434), .Z(n1436) );
  NAND U3523 ( .A(n1437), .B(n1436), .Z(n3231) );
  XNOR U3524 ( .A(n3232), .B(n3231), .Z(n3233) );
  XNOR U3525 ( .A(n3234), .B(n3233), .Z(n2876) );
  XOR U3526 ( .A(n2877), .B(n2876), .Z(n2878) );
  XOR U3527 ( .A(n2879), .B(n2878), .Z(n3057) );
  NANDN U3528 ( .A(n1439), .B(n1438), .Z(n1443) );
  NAND U3529 ( .A(n1441), .B(n1440), .Z(n1442) );
  NAND U3530 ( .A(n1443), .B(n1442), .Z(n3058) );
  XNOR U3531 ( .A(n3057), .B(n3058), .Z(n3059) );
  XOR U3532 ( .A(n3060), .B(n3059), .Z(n3117) );
  XNOR U3533 ( .A(n3118), .B(n3117), .Z(n3119) );
  XOR U3534 ( .A(n3120), .B(n3119), .Z(n3692) );
  NANDN U3535 ( .A(n1445), .B(n1444), .Z(n1449) );
  NAND U3536 ( .A(n1447), .B(n1446), .Z(n1448) );
  NAND U3537 ( .A(n1449), .B(n1448), .Z(n3691) );
  XOR U3538 ( .A(n3692), .B(n3691), .Z(n3694) );
  NAND U3539 ( .A(n1451), .B(n1450), .Z(n1455) );
  NANDN U3540 ( .A(n1453), .B(n1452), .Z(n1454) );
  NAND U3541 ( .A(n1455), .B(n1454), .Z(n3239) );
  NANDN U3542 ( .A(n1457), .B(n1456), .Z(n1461) );
  NANDN U3543 ( .A(n1459), .B(n1458), .Z(n1460) );
  AND U3544 ( .A(n1461), .B(n1460), .Z(n3222) );
  NANDN U3545 ( .A(n1463), .B(n1462), .Z(n1467) );
  NAND U3546 ( .A(n1465), .B(n1464), .Z(n1466) );
  AND U3547 ( .A(n1467), .B(n1466), .Z(n3220) );
  NAND U3548 ( .A(n1469), .B(n1468), .Z(n1473) );
  NANDN U3549 ( .A(n1471), .B(n1470), .Z(n1472) );
  NAND U3550 ( .A(n1473), .B(n1472), .Z(n3219) );
  XNOR U3551 ( .A(n3220), .B(n3219), .Z(n3221) );
  XNOR U3552 ( .A(n3222), .B(n3221), .Z(n3238) );
  NANDN U3553 ( .A(n1475), .B(n1474), .Z(n1479) );
  NANDN U3554 ( .A(n1477), .B(n1476), .Z(n1478) );
  AND U3555 ( .A(n1479), .B(n1478), .Z(n3237) );
  XOR U3556 ( .A(n3238), .B(n3237), .Z(n3240) );
  XNOR U3557 ( .A(n3239), .B(n3240), .Z(n3053) );
  NAND U3558 ( .A(n1481), .B(n1480), .Z(n1485) );
  NANDN U3559 ( .A(n1483), .B(n1482), .Z(n1484) );
  NAND U3560 ( .A(n1485), .B(n1484), .Z(n3130) );
  NANDN U3561 ( .A(n1487), .B(n1486), .Z(n1491) );
  NAND U3562 ( .A(n1489), .B(n1488), .Z(n1490) );
  AND U3563 ( .A(n1491), .B(n1490), .Z(n2831) );
  NAND U3564 ( .A(n1493), .B(n1492), .Z(n1497) );
  NAND U3565 ( .A(n1495), .B(n1494), .Z(n1496) );
  AND U3566 ( .A(n1497), .B(n1496), .Z(n3294) );
  NAND U3567 ( .A(n1499), .B(n1498), .Z(n1503) );
  NAND U3568 ( .A(n1501), .B(n1500), .Z(n1502) );
  AND U3569 ( .A(n1503), .B(n1502), .Z(n2659) );
  NAND U3570 ( .A(n1505), .B(n1504), .Z(n1509) );
  NAND U3571 ( .A(n1507), .B(n1506), .Z(n1508) );
  AND U3572 ( .A(n1509), .B(n1508), .Z(n2660) );
  NANDN U3573 ( .A(n1511), .B(n1510), .Z(n1515) );
  NAND U3574 ( .A(n1513), .B(n1512), .Z(n1514) );
  AND U3575 ( .A(n1515), .B(n1514), .Z(n2661) );
  XOR U3576 ( .A(n2662), .B(n2661), .Z(n3292) );
  NAND U3577 ( .A(n1517), .B(n1516), .Z(n1521) );
  NAND U3578 ( .A(n1519), .B(n1518), .Z(n1520) );
  NAND U3579 ( .A(n1521), .B(n1520), .Z(n3291) );
  XNOR U3580 ( .A(n3292), .B(n3291), .Z(n3293) );
  XOR U3581 ( .A(n3294), .B(n3293), .Z(n2829) );
  NANDN U3582 ( .A(n1523), .B(n1522), .Z(n1527) );
  NAND U3583 ( .A(n1525), .B(n1524), .Z(n1526) );
  NAND U3584 ( .A(n1527), .B(n1526), .Z(n2828) );
  XOR U3585 ( .A(n2829), .B(n2828), .Z(n2830) );
  XOR U3586 ( .A(n2831), .B(n2830), .Z(n3129) );
  XOR U3587 ( .A(n3130), .B(n3129), .Z(n3132) );
  NANDN U3588 ( .A(n1529), .B(n1528), .Z(n1533) );
  NAND U3589 ( .A(n1531), .B(n1530), .Z(n1532) );
  AND U3590 ( .A(n1533), .B(n1532), .Z(n3131) );
  XOR U3591 ( .A(n3132), .B(n3131), .Z(n3052) );
  NAND U3592 ( .A(n1535), .B(n1534), .Z(n1539) );
  NAND U3593 ( .A(n1537), .B(n1536), .Z(n1538) );
  AND U3594 ( .A(n1539), .B(n1538), .Z(n3174) );
  NAND U3595 ( .A(n1541), .B(n1540), .Z(n1545) );
  NAND U3596 ( .A(n1543), .B(n1542), .Z(n1544) );
  AND U3597 ( .A(n1545), .B(n1544), .Z(n3688) );
  NANDN U3598 ( .A(n1547), .B(n1546), .Z(n1551) );
  NANDN U3599 ( .A(n1549), .B(n1548), .Z(n1550) );
  AND U3600 ( .A(n1551), .B(n1550), .Z(n3686) );
  NAND U3601 ( .A(n1553), .B(n1552), .Z(n1557) );
  NAND U3602 ( .A(n1555), .B(n1554), .Z(n1556) );
  NAND U3603 ( .A(n1557), .B(n1556), .Z(n3685) );
  XNOR U3604 ( .A(n3686), .B(n3685), .Z(n3687) );
  XOR U3605 ( .A(n3688), .B(n3687), .Z(n3171) );
  NANDN U3606 ( .A(n1559), .B(n1558), .Z(n1563) );
  NAND U3607 ( .A(n1561), .B(n1560), .Z(n1562) );
  AND U3608 ( .A(n1563), .B(n1562), .Z(n2708) );
  NAND U3609 ( .A(n1565), .B(n1564), .Z(n1569) );
  NAND U3610 ( .A(n1567), .B(n1566), .Z(n1568) );
  AND U3611 ( .A(n1569), .B(n1568), .Z(n2846) );
  NAND U3612 ( .A(n1571), .B(n1570), .Z(n1575) );
  NAND U3613 ( .A(n1573), .B(n1572), .Z(n1574) );
  NAND U3614 ( .A(n1575), .B(n1574), .Z(n2847) );
  XNOR U3615 ( .A(n2846), .B(n2847), .Z(n2849) );
  NAND U3616 ( .A(n1577), .B(n1576), .Z(n1581) );
  NAND U3617 ( .A(n1579), .B(n1578), .Z(n1580) );
  AND U3618 ( .A(n1581), .B(n1580), .Z(n2848) );
  XOR U3619 ( .A(n2849), .B(n2848), .Z(n2813) );
  NAND U3620 ( .A(n1583), .B(n1582), .Z(n1587) );
  NAND U3621 ( .A(n1585), .B(n1584), .Z(n1586) );
  AND U3622 ( .A(n1587), .B(n1586), .Z(n3562) );
  NAND U3623 ( .A(n1589), .B(n1588), .Z(n1593) );
  NAND U3624 ( .A(n1591), .B(n1590), .Z(n1592) );
  NAND U3625 ( .A(n1593), .B(n1592), .Z(n3563) );
  XNOR U3626 ( .A(n3562), .B(n3563), .Z(n3565) );
  NAND U3627 ( .A(n1595), .B(n1594), .Z(n1599) );
  NAND U3628 ( .A(n1597), .B(n1596), .Z(n1598) );
  AND U3629 ( .A(n1599), .B(n1598), .Z(n3564) );
  XOR U3630 ( .A(n3565), .B(n3564), .Z(n2811) );
  NANDN U3631 ( .A(n1601), .B(n1600), .Z(n1605) );
  NAND U3632 ( .A(n1603), .B(n1602), .Z(n1604) );
  AND U3633 ( .A(n1605), .B(n1604), .Z(n2689) );
  NANDN U3634 ( .A(n1607), .B(n1606), .Z(n1611) );
  NAND U3635 ( .A(n1609), .B(n1608), .Z(n1610) );
  NAND U3636 ( .A(n1611), .B(n1610), .Z(n2690) );
  XNOR U3637 ( .A(n2689), .B(n2690), .Z(n2692) );
  NANDN U3638 ( .A(n1613), .B(n1612), .Z(n1617) );
  NAND U3639 ( .A(n1615), .B(n1614), .Z(n1616) );
  AND U3640 ( .A(n1617), .B(n1616), .Z(n2691) );
  XNOR U3641 ( .A(n2692), .B(n2691), .Z(n2810) );
  XNOR U3642 ( .A(n2811), .B(n2810), .Z(n2812) );
  XNOR U3643 ( .A(n2813), .B(n2812), .Z(n2707) );
  XOR U3644 ( .A(n2708), .B(n2707), .Z(n2710) );
  NAND U3645 ( .A(n1619), .B(n1618), .Z(n1623) );
  NAND U3646 ( .A(n1621), .B(n1620), .Z(n1622) );
  AND U3647 ( .A(n1623), .B(n1622), .Z(n3410) );
  NANDN U3648 ( .A(n1625), .B(n1624), .Z(n1629) );
  NAND U3649 ( .A(n1627), .B(n1626), .Z(n1628) );
  AND U3650 ( .A(n1629), .B(n1628), .Z(n2960) );
  NANDN U3651 ( .A(n1631), .B(n1630), .Z(n1635) );
  NAND U3652 ( .A(n1633), .B(n1632), .Z(n1634) );
  NAND U3653 ( .A(n1635), .B(n1634), .Z(n2961) );
  XNOR U3654 ( .A(n2960), .B(n2961), .Z(n2963) );
  NANDN U3655 ( .A(n1637), .B(n1636), .Z(n1641) );
  NAND U3656 ( .A(n1639), .B(n1638), .Z(n1640) );
  AND U3657 ( .A(n1641), .B(n1640), .Z(n2962) );
  XOR U3658 ( .A(n2963), .B(n2962), .Z(n3408) );
  NANDN U3659 ( .A(n1643), .B(n1642), .Z(n1647) );
  NANDN U3660 ( .A(n1645), .B(n1644), .Z(n1646) );
  AND U3661 ( .A(n1647), .B(n1646), .Z(n3407) );
  XNOR U3662 ( .A(n3408), .B(n3407), .Z(n3409) );
  XNOR U3663 ( .A(n3410), .B(n3409), .Z(n2709) );
  XOR U3664 ( .A(n2710), .B(n2709), .Z(n3172) );
  XOR U3665 ( .A(n3171), .B(n3172), .Z(n3173) );
  XOR U3666 ( .A(n3174), .B(n3173), .Z(n3051) );
  XOR U3667 ( .A(n3052), .B(n3051), .Z(n3054) );
  XNOR U3668 ( .A(n3053), .B(n3054), .Z(n3112) );
  NAND U3669 ( .A(n1649), .B(n1648), .Z(n1653) );
  NAND U3670 ( .A(n1651), .B(n1650), .Z(n1652) );
  NAND U3671 ( .A(n1653), .B(n1652), .Z(n3111) );
  XOR U3672 ( .A(n3112), .B(n3111), .Z(n3114) );
  NAND U3673 ( .A(n1655), .B(n1654), .Z(n1659) );
  NAND U3674 ( .A(n1657), .B(n1656), .Z(n1658) );
  NAND U3675 ( .A(n1659), .B(n1658), .Z(n2909) );
  NANDN U3676 ( .A(n1661), .B(n1660), .Z(n1665) );
  NAND U3677 ( .A(n1663), .B(n1662), .Z(n1664) );
  AND U3678 ( .A(n1665), .B(n1664), .Z(n3328) );
  NANDN U3679 ( .A(n1667), .B(n1666), .Z(n1671) );
  NAND U3680 ( .A(n1669), .B(n1668), .Z(n1670) );
  NAND U3681 ( .A(n1671), .B(n1670), .Z(n3329) );
  XNOR U3682 ( .A(n3328), .B(n3329), .Z(n3331) );
  NANDN U3683 ( .A(n1673), .B(n1672), .Z(n1677) );
  NAND U3684 ( .A(n1675), .B(n1674), .Z(n1676) );
  AND U3685 ( .A(n1677), .B(n1676), .Z(n3330) );
  XNOR U3686 ( .A(n3331), .B(n3330), .Z(n2907) );
  NANDN U3687 ( .A(n1679), .B(n1678), .Z(n1683) );
  NANDN U3688 ( .A(n1681), .B(n1680), .Z(n1682) );
  NAND U3689 ( .A(n1683), .B(n1682), .Z(n2906) );
  NAND U3690 ( .A(n1685), .B(n1684), .Z(n1689) );
  NAND U3691 ( .A(n1687), .B(n1686), .Z(n1688) );
  NAND U3692 ( .A(n1689), .B(n1688), .Z(n3374) );
  NANDN U3693 ( .A(n1691), .B(n1690), .Z(n1695) );
  NAND U3694 ( .A(n1693), .B(n1692), .Z(n1694) );
  AND U3695 ( .A(n1695), .B(n1694), .Z(n2942) );
  NANDN U3696 ( .A(n1697), .B(n1696), .Z(n1701) );
  NAND U3697 ( .A(n1699), .B(n1698), .Z(n1700) );
  NAND U3698 ( .A(n1701), .B(n1700), .Z(n2943) );
  XNOR U3699 ( .A(n2942), .B(n2943), .Z(n2945) );
  NANDN U3700 ( .A(n1703), .B(n1702), .Z(n1707) );
  NAND U3701 ( .A(n1705), .B(n1704), .Z(n1706) );
  AND U3702 ( .A(n1707), .B(n1706), .Z(n2944) );
  XNOR U3703 ( .A(n2945), .B(n2944), .Z(n3372) );
  NANDN U3704 ( .A(n1709), .B(n1708), .Z(n1713) );
  NANDN U3705 ( .A(n1711), .B(n1710), .Z(n1712) );
  AND U3706 ( .A(n1713), .B(n1712), .Z(n3371) );
  XOR U3707 ( .A(n3160), .B(n3159), .Z(n3162) );
  NANDN U3708 ( .A(n1715), .B(n1714), .Z(n1719) );
  NANDN U3709 ( .A(n1717), .B(n1716), .Z(n1718) );
  AND U3710 ( .A(n1719), .B(n1718), .Z(n3392) );
  NAND U3711 ( .A(n1721), .B(n1720), .Z(n1725) );
  NAND U3712 ( .A(n1723), .B(n1722), .Z(n1724) );
  AND U3713 ( .A(n1725), .B(n1724), .Z(n3390) );
  NAND U3714 ( .A(n1727), .B(n1726), .Z(n1731) );
  NAND U3715 ( .A(n1729), .B(n1728), .Z(n1730) );
  AND U3716 ( .A(n1731), .B(n1730), .Z(n3039) );
  NAND U3717 ( .A(n1733), .B(n1732), .Z(n1737) );
  NAND U3718 ( .A(n1735), .B(n1734), .Z(n1736) );
  AND U3719 ( .A(n1737), .B(n1736), .Z(n3040) );
  NANDN U3720 ( .A(n1739), .B(n1738), .Z(n1743) );
  NAND U3721 ( .A(n1741), .B(n1740), .Z(n1742) );
  AND U3722 ( .A(n1743), .B(n1742), .Z(n3041) );
  XNOR U3723 ( .A(n3042), .B(n3041), .Z(n3389) );
  XNOR U3724 ( .A(n3390), .B(n3389), .Z(n3391) );
  XOR U3725 ( .A(n3392), .B(n3391), .Z(n3161) );
  XOR U3726 ( .A(n3162), .B(n3161), .Z(n3108) );
  NANDN U3727 ( .A(n1745), .B(n1744), .Z(n1749) );
  NANDN U3728 ( .A(n1747), .B(n1746), .Z(n1748) );
  AND U3729 ( .A(n1749), .B(n1748), .Z(n2771) );
  NAND U3730 ( .A(n1751), .B(n1750), .Z(n1755) );
  NAND U3731 ( .A(n1753), .B(n1752), .Z(n1754) );
  AND U3732 ( .A(n1755), .B(n1754), .Z(n2762) );
  NAND U3733 ( .A(n1757), .B(n1756), .Z(n1761) );
  NAND U3734 ( .A(n1759), .B(n1758), .Z(n1760) );
  AND U3735 ( .A(n1761), .B(n1760), .Z(n2763) );
  NAND U3736 ( .A(n1763), .B(n1762), .Z(n1767) );
  NAND U3737 ( .A(n1765), .B(n1764), .Z(n1766) );
  AND U3738 ( .A(n1767), .B(n1766), .Z(n2764) );
  XOR U3739 ( .A(n2765), .B(n2764), .Z(n2769) );
  NANDN U3740 ( .A(n1769), .B(n1768), .Z(n1773) );
  NANDN U3741 ( .A(n1771), .B(n1770), .Z(n1772) );
  AND U3742 ( .A(n1773), .B(n1772), .Z(n2768) );
  XNOR U3743 ( .A(n2769), .B(n2768), .Z(n2770) );
  XOR U3744 ( .A(n2771), .B(n2770), .Z(n3196) );
  NAND U3745 ( .A(n1775), .B(n1774), .Z(n1779) );
  NAND U3746 ( .A(n1777), .B(n1776), .Z(n1778) );
  AND U3747 ( .A(n1779), .B(n1778), .Z(n3528) );
  NANDN U3748 ( .A(n1781), .B(n1780), .Z(n1785) );
  NAND U3749 ( .A(n1783), .B(n1782), .Z(n1784) );
  NAND U3750 ( .A(n1785), .B(n1784), .Z(n3530) );
  NAND U3751 ( .A(n1787), .B(n1786), .Z(n1791) );
  NAND U3752 ( .A(n1789), .B(n1788), .Z(n1790) );
  AND U3753 ( .A(n1791), .B(n1790), .Z(n3529) );
  NANDN U3754 ( .A(n1793), .B(n1792), .Z(n1797) );
  NAND U3755 ( .A(n1795), .B(n1794), .Z(n1796) );
  AND U3756 ( .A(n1797), .B(n1796), .Z(n2792) );
  NANDN U3757 ( .A(n1799), .B(n1798), .Z(n1803) );
  NAND U3758 ( .A(n1801), .B(n1800), .Z(n1802) );
  AND U3759 ( .A(n1803), .B(n1802), .Z(n2793) );
  NAND U3760 ( .A(n1805), .B(n1804), .Z(n1809) );
  NAND U3761 ( .A(n1807), .B(n1806), .Z(n1808) );
  AND U3762 ( .A(n1809), .B(n1808), .Z(n2794) );
  XNOR U3763 ( .A(n2795), .B(n2794), .Z(n2642) );
  NAND U3764 ( .A(n1811), .B(n1810), .Z(n1815) );
  NAND U3765 ( .A(n1813), .B(n1812), .Z(n1814) );
  AND U3766 ( .A(n1815), .B(n1814), .Z(n2744) );
  NAND U3767 ( .A(n1817), .B(n1816), .Z(n1821) );
  NAND U3768 ( .A(n1819), .B(n1818), .Z(n1820) );
  NAND U3769 ( .A(n1821), .B(n1820), .Z(n2745) );
  XNOR U3770 ( .A(n2744), .B(n2745), .Z(n2747) );
  NAND U3771 ( .A(n1823), .B(n1822), .Z(n1827) );
  NAND U3772 ( .A(n1825), .B(n1824), .Z(n1826) );
  AND U3773 ( .A(n1827), .B(n1826), .Z(n2746) );
  XNOR U3774 ( .A(n2747), .B(n2746), .Z(n2641) );
  XOR U3775 ( .A(n2643), .B(n2644), .Z(n3195) );
  XOR U3776 ( .A(n3196), .B(n3195), .Z(n3198) );
  NANDN U3777 ( .A(n1829), .B(n1828), .Z(n1833) );
  NANDN U3778 ( .A(n1831), .B(n1830), .Z(n1832) );
  AND U3779 ( .A(n1833), .B(n1832), .Z(n2729) );
  NAND U3780 ( .A(n1835), .B(n1834), .Z(n1839) );
  NAND U3781 ( .A(n1837), .B(n1836), .Z(n1838) );
  AND U3782 ( .A(n1839), .B(n1838), .Z(n2864) );
  NAND U3783 ( .A(n1841), .B(n1840), .Z(n1845) );
  NAND U3784 ( .A(n1843), .B(n1842), .Z(n1844) );
  AND U3785 ( .A(n1845), .B(n1844), .Z(n2865) );
  NANDN U3786 ( .A(n1847), .B(n1846), .Z(n1851) );
  NAND U3787 ( .A(n1849), .B(n1848), .Z(n1850) );
  AND U3788 ( .A(n1851), .B(n1850), .Z(n2866) );
  XOR U3789 ( .A(n2867), .B(n2866), .Z(n2727) );
  NANDN U3790 ( .A(n1853), .B(n1852), .Z(n1857) );
  NAND U3791 ( .A(n1855), .B(n1854), .Z(n1856) );
  AND U3792 ( .A(n1857), .B(n1856), .Z(n3604) );
  NANDN U3793 ( .A(n1859), .B(n1858), .Z(n1863) );
  NAND U3794 ( .A(n1861), .B(n1860), .Z(n1862) );
  NAND U3795 ( .A(n1863), .B(n1862), .Z(n3605) );
  XNOR U3796 ( .A(n3604), .B(n3605), .Z(n3607) );
  NANDN U3797 ( .A(n1865), .B(n1864), .Z(n1869) );
  NAND U3798 ( .A(n1867), .B(n1866), .Z(n1868) );
  AND U3799 ( .A(n1869), .B(n1868), .Z(n3606) );
  XNOR U3800 ( .A(n3607), .B(n3606), .Z(n2726) );
  XNOR U3801 ( .A(n2727), .B(n2726), .Z(n2728) );
  XOR U3802 ( .A(n2729), .B(n2728), .Z(n3197) );
  XOR U3803 ( .A(n3198), .B(n3197), .Z(n3106) );
  NANDN U3804 ( .A(n1871), .B(n1870), .Z(n1875) );
  NAND U3805 ( .A(n1873), .B(n1872), .Z(n1874) );
  AND U3806 ( .A(n1875), .B(n1874), .Z(n2623) );
  NANDN U3807 ( .A(n1877), .B(n1876), .Z(n1881) );
  NAND U3808 ( .A(n1879), .B(n1878), .Z(n1880) );
  AND U3809 ( .A(n1881), .B(n1880), .Z(n2624) );
  NAND U3810 ( .A(n1883), .B(n1882), .Z(n1887) );
  NAND U3811 ( .A(n1885), .B(n1884), .Z(n1886) );
  AND U3812 ( .A(n1887), .B(n1886), .Z(n2625) );
  XNOR U3813 ( .A(n2626), .B(n2625), .Z(n3356) );
  NANDN U3814 ( .A(n1889), .B(n1888), .Z(n1893) );
  NANDN U3815 ( .A(n1891), .B(n1890), .Z(n1892) );
  AND U3816 ( .A(n1893), .B(n1892), .Z(n3357) );
  NANDN U3817 ( .A(n1895), .B(n1894), .Z(n1899) );
  NANDN U3818 ( .A(n1897), .B(n1896), .Z(n1898) );
  NAND U3819 ( .A(n1899), .B(n1898), .Z(n3355) );
  XOR U3820 ( .A(n3357), .B(n3355), .Z(n1900) );
  XNOR U3821 ( .A(n3356), .B(n1900), .Z(n3156) );
  NANDN U3822 ( .A(n1902), .B(n1901), .Z(n1906) );
  NANDN U3823 ( .A(n1904), .B(n1903), .Z(n1905) );
  AND U3824 ( .A(n1906), .B(n1905), .Z(n3276) );
  NAND U3825 ( .A(n1908), .B(n1907), .Z(n1912) );
  NAND U3826 ( .A(n1910), .B(n1909), .Z(n1911) );
  AND U3827 ( .A(n1912), .B(n1911), .Z(n2936) );
  NAND U3828 ( .A(n1914), .B(n1913), .Z(n1918) );
  NAND U3829 ( .A(n1916), .B(n1915), .Z(n1917) );
  NAND U3830 ( .A(n1918), .B(n1917), .Z(n2937) );
  XNOR U3831 ( .A(n2936), .B(n2937), .Z(n2939) );
  NAND U3832 ( .A(n1920), .B(n1919), .Z(n1924) );
  NAND U3833 ( .A(n1922), .B(n1921), .Z(n1923) );
  AND U3834 ( .A(n1924), .B(n1923), .Z(n2938) );
  XOR U3835 ( .A(n2939), .B(n2938), .Z(n3274) );
  NANDN U3836 ( .A(n1926), .B(n1925), .Z(n1930) );
  NANDN U3837 ( .A(n1928), .B(n1927), .Z(n1929) );
  AND U3838 ( .A(n1930), .B(n1929), .Z(n3273) );
  XNOR U3839 ( .A(n3274), .B(n3273), .Z(n3275) );
  XOR U3840 ( .A(n3276), .B(n3275), .Z(n3154) );
  NAND U3841 ( .A(n1932), .B(n1931), .Z(n1936) );
  NAND U3842 ( .A(n1934), .B(n1933), .Z(n1935) );
  AND U3843 ( .A(n1936), .B(n1935), .Z(n3258) );
  NAND U3844 ( .A(n1938), .B(n1937), .Z(n1942) );
  NAND U3845 ( .A(n1940), .B(n1939), .Z(n1941) );
  AND U3846 ( .A(n1942), .B(n1941), .Z(n3256) );
  NAND U3847 ( .A(n1944), .B(n1943), .Z(n1948) );
  NAND U3848 ( .A(n1946), .B(n1945), .Z(n1947) );
  AND U3849 ( .A(n1948), .B(n1947), .Z(n2948) );
  NAND U3850 ( .A(n1950), .B(n1949), .Z(n1954) );
  NAND U3851 ( .A(n1952), .B(n1951), .Z(n1953) );
  NAND U3852 ( .A(n1954), .B(n1953), .Z(n2949) );
  XNOR U3853 ( .A(n2948), .B(n2949), .Z(n2951) );
  NAND U3854 ( .A(n1956), .B(n1955), .Z(n1960) );
  NAND U3855 ( .A(n1958), .B(n1957), .Z(n1959) );
  AND U3856 ( .A(n1960), .B(n1959), .Z(n2950) );
  XNOR U3857 ( .A(n2951), .B(n2950), .Z(n3255) );
  XNOR U3858 ( .A(n3256), .B(n3255), .Z(n3257) );
  XNOR U3859 ( .A(n3258), .B(n3257), .Z(n3153) );
  XOR U3860 ( .A(n3154), .B(n3153), .Z(n3155) );
  XNOR U3861 ( .A(n3156), .B(n3155), .Z(n3105) );
  XNOR U3862 ( .A(n3106), .B(n3105), .Z(n3107) );
  XNOR U3863 ( .A(n3108), .B(n3107), .Z(n3124) );
  NANDN U3864 ( .A(n1962), .B(n1961), .Z(n1966) );
  NAND U3865 ( .A(n1964), .B(n1963), .Z(n1965) );
  AND U3866 ( .A(n1966), .B(n1965), .Z(n2999) );
  NANDN U3867 ( .A(n1968), .B(n1967), .Z(n1972) );
  NAND U3868 ( .A(n1970), .B(n1969), .Z(n1971) );
  NAND U3869 ( .A(n1972), .B(n1971), .Z(n3000) );
  XNOR U3870 ( .A(n2999), .B(n3000), .Z(n3002) );
  NAND U3871 ( .A(n1974), .B(n1973), .Z(n1978) );
  NAND U3872 ( .A(n1976), .B(n1975), .Z(n1977) );
  AND U3873 ( .A(n1978), .B(n1977), .Z(n3001) );
  XOR U3874 ( .A(n3002), .B(n3001), .Z(n3619) );
  NANDN U3875 ( .A(n1980), .B(n1979), .Z(n1984) );
  NAND U3876 ( .A(n1982), .B(n1981), .Z(n1983) );
  AND U3877 ( .A(n1984), .B(n1983), .Z(n3622) );
  NANDN U3878 ( .A(n1986), .B(n1985), .Z(n1990) );
  NAND U3879 ( .A(n1988), .B(n1987), .Z(n1989) );
  AND U3880 ( .A(n1990), .B(n1989), .Z(n3623) );
  NANDN U3881 ( .A(n1992), .B(n1991), .Z(n1996) );
  NAND U3882 ( .A(n1994), .B(n1993), .Z(n1995) );
  AND U3883 ( .A(n1996), .B(n1995), .Z(n3624) );
  XOR U3884 ( .A(n3625), .B(n3624), .Z(n3617) );
  NANDN U3885 ( .A(n1998), .B(n1997), .Z(n2002) );
  NANDN U3886 ( .A(n2000), .B(n1999), .Z(n2001) );
  AND U3887 ( .A(n2002), .B(n2001), .Z(n3616) );
  XNOR U3888 ( .A(n3617), .B(n3616), .Z(n3618) );
  XOR U3889 ( .A(n3619), .B(n3618), .Z(n3137) );
  NAND U3890 ( .A(n2004), .B(n2003), .Z(n2008) );
  NAND U3891 ( .A(n2006), .B(n2005), .Z(n2007) );
  AND U3892 ( .A(n2008), .B(n2007), .Z(n3136) );
  NANDN U3893 ( .A(n2010), .B(n2009), .Z(n2014) );
  NAND U3894 ( .A(n2012), .B(n2011), .Z(n2013) );
  NAND U3895 ( .A(n2014), .B(n2013), .Z(n2981) );
  NANDN U3896 ( .A(n2016), .B(n2015), .Z(n2020) );
  NAND U3897 ( .A(n2018), .B(n2017), .Z(n2019) );
  AND U3898 ( .A(n2020), .B(n2019), .Z(n2984) );
  NANDN U3899 ( .A(n2022), .B(n2021), .Z(n2026) );
  NAND U3900 ( .A(n2024), .B(n2023), .Z(n2025) );
  AND U3901 ( .A(n2026), .B(n2025), .Z(n2982) );
  XNOR U3902 ( .A(n2984), .B(n2982), .Z(n2027) );
  XOR U3903 ( .A(n2981), .B(n2027), .Z(n3005) );
  NANDN U3904 ( .A(n2029), .B(n2028), .Z(n2033) );
  NANDN U3905 ( .A(n2031), .B(n2030), .Z(n2032) );
  AND U3906 ( .A(n2033), .B(n2032), .Z(n3007) );
  NANDN U3907 ( .A(n2035), .B(n2034), .Z(n2039) );
  NAND U3908 ( .A(n2037), .B(n2036), .Z(n2038) );
  AND U3909 ( .A(n2039), .B(n2038), .Z(n3638) );
  NANDN U3910 ( .A(n2041), .B(n2040), .Z(n2045) );
  NAND U3911 ( .A(n2043), .B(n2042), .Z(n2044) );
  NAND U3912 ( .A(n2045), .B(n2044), .Z(n3639) );
  XNOR U3913 ( .A(n3638), .B(n3639), .Z(n3640) );
  NANDN U3914 ( .A(n2047), .B(n2046), .Z(n2051) );
  NAND U3915 ( .A(n2049), .B(n2048), .Z(n2050) );
  NAND U3916 ( .A(n2051), .B(n2050), .Z(n3641) );
  XNOR U3917 ( .A(n3640), .B(n3641), .Z(n3006) );
  XNOR U3918 ( .A(n3007), .B(n3006), .Z(n2052) );
  XOR U3919 ( .A(n3005), .B(n2052), .Z(n3135) );
  XNOR U3920 ( .A(n3136), .B(n3135), .Z(n3138) );
  XOR U3921 ( .A(n3137), .B(n3138), .Z(n2885) );
  NANDN U3922 ( .A(n2054), .B(n2053), .Z(n2058) );
  NANDN U3923 ( .A(n2056), .B(n2055), .Z(n2057) );
  AND U3924 ( .A(n2058), .B(n2057), .Z(n3202) );
  NAND U3925 ( .A(n2060), .B(n2059), .Z(n2064) );
  NAND U3926 ( .A(n2062), .B(n2061), .Z(n2063) );
  AND U3927 ( .A(n2064), .B(n2063), .Z(n2798) );
  NAND U3928 ( .A(n2066), .B(n2065), .Z(n2070) );
  NAND U3929 ( .A(n2068), .B(n2067), .Z(n2069) );
  AND U3930 ( .A(n2070), .B(n2069), .Z(n2799) );
  NAND U3931 ( .A(n2072), .B(n2071), .Z(n2076) );
  NAND U3932 ( .A(n2074), .B(n2073), .Z(n2075) );
  AND U3933 ( .A(n2076), .B(n2075), .Z(n2800) );
  XNOR U3934 ( .A(n2801), .B(n2800), .Z(n2686) );
  NANDN U3935 ( .A(n2078), .B(n2077), .Z(n2082) );
  NAND U3936 ( .A(n2080), .B(n2079), .Z(n2081) );
  AND U3937 ( .A(n2082), .B(n2081), .Z(n3580) );
  NANDN U3938 ( .A(n2084), .B(n2083), .Z(n2088) );
  NAND U3939 ( .A(n2086), .B(n2085), .Z(n2087) );
  NAND U3940 ( .A(n2088), .B(n2087), .Z(n3581) );
  XNOR U3941 ( .A(n3580), .B(n3581), .Z(n3583) );
  NANDN U3942 ( .A(n2090), .B(n2089), .Z(n2094) );
  NAND U3943 ( .A(n2092), .B(n2091), .Z(n2093) );
  AND U3944 ( .A(n2094), .B(n2093), .Z(n3582) );
  XNOR U3945 ( .A(n3583), .B(n3582), .Z(n2684) );
  NAND U3946 ( .A(n2096), .B(n2095), .Z(n2100) );
  NAND U3947 ( .A(n2098), .B(n2097), .Z(n2099) );
  NAND U3948 ( .A(n2100), .B(n2099), .Z(n2713) );
  NAND U3949 ( .A(n2102), .B(n2101), .Z(n2106) );
  NAND U3950 ( .A(n2104), .B(n2103), .Z(n2105) );
  AND U3951 ( .A(n2106), .B(n2105), .Z(n2715) );
  NAND U3952 ( .A(n2108), .B(n2107), .Z(n2112) );
  NAND U3953 ( .A(n2110), .B(n2109), .Z(n2111) );
  AND U3954 ( .A(n2112), .B(n2111), .Z(n2714) );
  XNOR U3955 ( .A(n2715), .B(n2714), .Z(n2113) );
  XNOR U3956 ( .A(n2713), .B(n2113), .Z(n2683) );
  XOR U3957 ( .A(n3202), .B(n3201), .Z(n3204) );
  NANDN U3958 ( .A(n2115), .B(n2114), .Z(n2119) );
  NANDN U3959 ( .A(n2117), .B(n2116), .Z(n2118) );
  AND U3960 ( .A(n2119), .B(n2118), .Z(n3446) );
  NAND U3961 ( .A(n2121), .B(n2120), .Z(n2125) );
  NAND U3962 ( .A(n2123), .B(n2122), .Z(n2124) );
  AND U3963 ( .A(n2125), .B(n2124), .Z(n2954) );
  NAND U3964 ( .A(n2127), .B(n2126), .Z(n2131) );
  NAND U3965 ( .A(n2129), .B(n2128), .Z(n2130) );
  NAND U3966 ( .A(n2131), .B(n2130), .Z(n2955) );
  XNOR U3967 ( .A(n2954), .B(n2955), .Z(n2957) );
  NANDN U3968 ( .A(n2133), .B(n2132), .Z(n2137) );
  NAND U3969 ( .A(n2135), .B(n2134), .Z(n2136) );
  AND U3970 ( .A(n2137), .B(n2136), .Z(n2956) );
  XOR U3971 ( .A(n2957), .B(n2956), .Z(n3444) );
  NANDN U3972 ( .A(n2139), .B(n2138), .Z(n2143) );
  NANDN U3973 ( .A(n2141), .B(n2140), .Z(n2142) );
  AND U3974 ( .A(n2143), .B(n2142), .Z(n3443) );
  XNOR U3975 ( .A(n3444), .B(n3443), .Z(n3445) );
  XOR U3976 ( .A(n3446), .B(n3445), .Z(n3203) );
  XOR U3977 ( .A(n3204), .B(n3203), .Z(n2883) );
  NANDN U3978 ( .A(n2145), .B(n2144), .Z(n2149) );
  NANDN U3979 ( .A(n2147), .B(n2146), .Z(n2148) );
  AND U3980 ( .A(n2149), .B(n2148), .Z(n2620) );
  NAND U3981 ( .A(n2151), .B(n2150), .Z(n2155) );
  NAND U3982 ( .A(n2153), .B(n2152), .Z(n2154) );
  AND U3983 ( .A(n2155), .B(n2154), .Z(n3540) );
  NANDN U3984 ( .A(n2157), .B(n2156), .Z(n2161) );
  NAND U3985 ( .A(n2159), .B(n2158), .Z(n2160) );
  NAND U3986 ( .A(n2161), .B(n2160), .Z(n3542) );
  NAND U3987 ( .A(n2163), .B(n2162), .Z(n2167) );
  NAND U3988 ( .A(n2165), .B(n2164), .Z(n2166) );
  NAND U3989 ( .A(n2167), .B(n2166), .Z(n3541) );
  XNOR U3990 ( .A(n3542), .B(n3541), .Z(n2168) );
  XOR U3991 ( .A(n3540), .B(n2168), .Z(n2617) );
  NANDN U3992 ( .A(n2170), .B(n2169), .Z(n2174) );
  NANDN U3993 ( .A(n2172), .B(n2171), .Z(n2173) );
  AND U3994 ( .A(n2174), .B(n2173), .Z(n2618) );
  XOR U3995 ( .A(n2617), .B(n2618), .Z(n2619) );
  XOR U3996 ( .A(n2620), .B(n2619), .Z(n3150) );
  NANDN U3997 ( .A(n2176), .B(n2175), .Z(n2180) );
  NAND U3998 ( .A(n2178), .B(n2177), .Z(n2179) );
  AND U3999 ( .A(n2180), .B(n2179), .Z(n3644) );
  NANDN U4000 ( .A(n2182), .B(n2181), .Z(n2186) );
  NAND U4001 ( .A(n2184), .B(n2183), .Z(n2185) );
  AND U4002 ( .A(n2186), .B(n2185), .Z(n3645) );
  NANDN U4003 ( .A(n2188), .B(n2187), .Z(n2192) );
  NAND U4004 ( .A(n2190), .B(n2189), .Z(n2191) );
  AND U4005 ( .A(n2192), .B(n2191), .Z(n3647) );
  XNOR U4006 ( .A(n3646), .B(n3647), .Z(n3635) );
  NANDN U4007 ( .A(n2194), .B(n2193), .Z(n2198) );
  NAND U4008 ( .A(n2196), .B(n2195), .Z(n2197) );
  AND U4009 ( .A(n2198), .B(n2197), .Z(n3656) );
  NANDN U4010 ( .A(n2200), .B(n2199), .Z(n2204) );
  NAND U4011 ( .A(n2202), .B(n2201), .Z(n2203) );
  AND U4012 ( .A(n2204), .B(n2203), .Z(n3657) );
  NANDN U4013 ( .A(n2206), .B(n2205), .Z(n2210) );
  NAND U4014 ( .A(n2208), .B(n2207), .Z(n2209) );
  AND U4015 ( .A(n2210), .B(n2209), .Z(n3659) );
  NANDN U4016 ( .A(n2212), .B(n2211), .Z(n2216) );
  NAND U4017 ( .A(n2214), .B(n2213), .Z(n2215) );
  AND U4018 ( .A(n2216), .B(n2215), .Z(n3636) );
  XNOR U4019 ( .A(n3637), .B(n3636), .Z(n2217) );
  XOR U4020 ( .A(n3635), .B(n2217), .Z(n3147) );
  NAND U4021 ( .A(n2219), .B(n2218), .Z(n2223) );
  NAND U4022 ( .A(n2221), .B(n2220), .Z(n2222) );
  AND U4023 ( .A(n2223), .B(n2222), .Z(n3148) );
  XNOR U4024 ( .A(n3147), .B(n3148), .Z(n3149) );
  XNOR U4025 ( .A(n3150), .B(n3149), .Z(n2882) );
  XNOR U4026 ( .A(n2883), .B(n2882), .Z(n2884) );
  XOR U4027 ( .A(n2885), .B(n2884), .Z(n3123) );
  XOR U4028 ( .A(n3124), .B(n3123), .Z(n3126) );
  NANDN U4029 ( .A(n2225), .B(n2224), .Z(n2229) );
  NAND U4030 ( .A(n2227), .B(n2226), .Z(n2228) );
  AND U4031 ( .A(n2229), .B(n2228), .Z(n2695) );
  NANDN U4032 ( .A(n2231), .B(n2230), .Z(n2235) );
  NAND U4033 ( .A(n2233), .B(n2232), .Z(n2234) );
  NAND U4034 ( .A(n2235), .B(n2234), .Z(n2696) );
  XNOR U4035 ( .A(n2695), .B(n2696), .Z(n2698) );
  NANDN U4036 ( .A(n2237), .B(n2236), .Z(n2241) );
  NAND U4037 ( .A(n2239), .B(n2238), .Z(n2240) );
  AND U4038 ( .A(n2241), .B(n2240), .Z(n2697) );
  XOR U4039 ( .A(n2698), .B(n2697), .Z(n3577) );
  NAND U4040 ( .A(n2243), .B(n2242), .Z(n2247) );
  NAND U4041 ( .A(n2245), .B(n2244), .Z(n2246) );
  AND U4042 ( .A(n2247), .B(n2246), .Z(n3586) );
  NAND U4043 ( .A(n2249), .B(n2248), .Z(n2253) );
  NAND U4044 ( .A(n2251), .B(n2250), .Z(n2252) );
  NAND U4045 ( .A(n2253), .B(n2252), .Z(n3587) );
  XNOR U4046 ( .A(n3586), .B(n3587), .Z(n3589) );
  NAND U4047 ( .A(n2255), .B(n2254), .Z(n2259) );
  NAND U4048 ( .A(n2257), .B(n2256), .Z(n2258) );
  AND U4049 ( .A(n2259), .B(n2258), .Z(n3588) );
  XOR U4050 ( .A(n3589), .B(n3588), .Z(n3575) );
  NAND U4051 ( .A(n2261), .B(n2260), .Z(n2265) );
  NAND U4052 ( .A(n2263), .B(n2262), .Z(n2264) );
  AND U4053 ( .A(n2265), .B(n2264), .Z(n2827) );
  NAND U4054 ( .A(n2267), .B(n2266), .Z(n2271) );
  NAND U4055 ( .A(n2269), .B(n2268), .Z(n2270) );
  AND U4056 ( .A(n2271), .B(n2270), .Z(n2826) );
  NAND U4057 ( .A(n2273), .B(n2272), .Z(n2277) );
  NAND U4058 ( .A(n2275), .B(n2274), .Z(n2276) );
  AND U4059 ( .A(n2277), .B(n2276), .Z(n2825) );
  XNOR U4060 ( .A(n3575), .B(n3574), .Z(n3576) );
  XOR U4061 ( .A(n3577), .B(n3576), .Z(n3215) );
  NANDN U4062 ( .A(n2279), .B(n2278), .Z(n2283) );
  NANDN U4063 ( .A(n2281), .B(n2280), .Z(n2282) );
  AND U4064 ( .A(n2283), .B(n2282), .Z(n3214) );
  NAND U4065 ( .A(n2285), .B(n2284), .Z(n2289) );
  NAND U4066 ( .A(n2287), .B(n2286), .Z(n2288) );
  NAND U4067 ( .A(n2289), .B(n2288), .Z(n3315) );
  NAND U4068 ( .A(n2291), .B(n2290), .Z(n2295) );
  NAND U4069 ( .A(n2293), .B(n2292), .Z(n2294) );
  AND U4070 ( .A(n2295), .B(n2294), .Z(n3317) );
  NAND U4071 ( .A(n2297), .B(n2296), .Z(n2301) );
  NAND U4072 ( .A(n2299), .B(n2298), .Z(n2300) );
  AND U4073 ( .A(n2301), .B(n2300), .Z(n3316) );
  XNOR U4074 ( .A(n3317), .B(n3316), .Z(n2302) );
  XOR U4075 ( .A(n3315), .B(n2302), .Z(n3548) );
  NAND U4076 ( .A(n2304), .B(n2303), .Z(n2308) );
  NAND U4077 ( .A(n2306), .B(n2305), .Z(n2307) );
  AND U4078 ( .A(n2308), .B(n2307), .Z(n3568) );
  NAND U4079 ( .A(n2310), .B(n2309), .Z(n2314) );
  NAND U4080 ( .A(n2312), .B(n2311), .Z(n2313) );
  AND U4081 ( .A(n2314), .B(n2313), .Z(n3569) );
  NAND U4082 ( .A(n2316), .B(n2315), .Z(n2320) );
  NAND U4083 ( .A(n2318), .B(n2317), .Z(n2319) );
  AND U4084 ( .A(n2320), .B(n2319), .Z(n3571) );
  XNOR U4085 ( .A(n3570), .B(n3571), .Z(n3546) );
  NANDN U4086 ( .A(n2322), .B(n2321), .Z(n2326) );
  NAND U4087 ( .A(n2324), .B(n2323), .Z(n2325) );
  AND U4088 ( .A(n2326), .B(n2325), .Z(n3340) );
  NANDN U4089 ( .A(n2328), .B(n2327), .Z(n2332) );
  NAND U4090 ( .A(n2330), .B(n2329), .Z(n2331) );
  NAND U4091 ( .A(n2332), .B(n2331), .Z(n3341) );
  XNOR U4092 ( .A(n3340), .B(n3341), .Z(n3342) );
  NANDN U4093 ( .A(n2334), .B(n2333), .Z(n2338) );
  NAND U4094 ( .A(n2336), .B(n2335), .Z(n2337) );
  NAND U4095 ( .A(n2338), .B(n2337), .Z(n3343) );
  XNOR U4096 ( .A(n3342), .B(n3343), .Z(n3547) );
  XOR U4097 ( .A(n3546), .B(n3547), .Z(n2339) );
  XNOR U4098 ( .A(n3548), .B(n2339), .Z(n3213) );
  XNOR U4099 ( .A(n3214), .B(n3213), .Z(n3216) );
  XOR U4100 ( .A(n3215), .B(n3216), .Z(n3180) );
  NAND U4101 ( .A(n2341), .B(n2340), .Z(n2345) );
  NAND U4102 ( .A(n2343), .B(n2342), .Z(n2344) );
  AND U4103 ( .A(n2345), .B(n2344), .Z(n3304) );
  NANDN U4104 ( .A(n2347), .B(n2346), .Z(n2351) );
  NAND U4105 ( .A(n2349), .B(n2348), .Z(n2350) );
  AND U4106 ( .A(n2351), .B(n2350), .Z(n2701) );
  NAND U4107 ( .A(n2353), .B(n2352), .Z(n2357) );
  NAND U4108 ( .A(n2355), .B(n2354), .Z(n2356) );
  NAND U4109 ( .A(n2357), .B(n2356), .Z(n2702) );
  XNOR U4110 ( .A(n2701), .B(n2702), .Z(n2704) );
  NAND U4111 ( .A(n2359), .B(n2358), .Z(n2363) );
  NAND U4112 ( .A(n2361), .B(n2360), .Z(n2362) );
  AND U4113 ( .A(n2363), .B(n2362), .Z(n2703) );
  XOR U4114 ( .A(n2704), .B(n2703), .Z(n2855) );
  NAND U4115 ( .A(n2365), .B(n2364), .Z(n2369) );
  NAND U4116 ( .A(n2367), .B(n2366), .Z(n2368) );
  AND U4117 ( .A(n2369), .B(n2368), .Z(n2665) );
  NAND U4118 ( .A(n2371), .B(n2370), .Z(n2375) );
  NAND U4119 ( .A(n2373), .B(n2372), .Z(n2374) );
  AND U4120 ( .A(n2375), .B(n2374), .Z(n2666) );
  NAND U4121 ( .A(n2377), .B(n2376), .Z(n2381) );
  NAND U4122 ( .A(n2379), .B(n2378), .Z(n2380) );
  AND U4123 ( .A(n2381), .B(n2380), .Z(n2667) );
  XOR U4124 ( .A(n2668), .B(n2667), .Z(n2853) );
  NAND U4125 ( .A(n2383), .B(n2382), .Z(n2387) );
  NAND U4126 ( .A(n2385), .B(n2384), .Z(n2386) );
  AND U4127 ( .A(n2387), .B(n2386), .Z(n2586) );
  NAND U4128 ( .A(n2389), .B(n2388), .Z(n2393) );
  NAND U4129 ( .A(n2391), .B(n2390), .Z(n2392) );
  NAND U4130 ( .A(n2393), .B(n2392), .Z(n2587) );
  XNOR U4131 ( .A(n2586), .B(n2587), .Z(n2589) );
  NAND U4132 ( .A(n2395), .B(n2394), .Z(n2399) );
  NAND U4133 ( .A(n2397), .B(n2396), .Z(n2398) );
  AND U4134 ( .A(n2399), .B(n2398), .Z(n2588) );
  XNOR U4135 ( .A(n2589), .B(n2588), .Z(n2852) );
  XNOR U4136 ( .A(n2853), .B(n2852), .Z(n2854) );
  XNOR U4137 ( .A(n2855), .B(n2854), .Z(n3303) );
  XOR U4138 ( .A(n3304), .B(n3303), .Z(n3306) );
  NAND U4139 ( .A(n2401), .B(n2400), .Z(n2405) );
  NAND U4140 ( .A(n2403), .B(n2402), .Z(n2404) );
  AND U4141 ( .A(n2405), .B(n2404), .Z(n2610) );
  NAND U4142 ( .A(n2407), .B(n2406), .Z(n2411) );
  NAND U4143 ( .A(n2409), .B(n2408), .Z(n2410) );
  NAND U4144 ( .A(n2411), .B(n2410), .Z(n2611) );
  XNOR U4145 ( .A(n2610), .B(n2611), .Z(n2613) );
  NAND U4146 ( .A(n2413), .B(n2412), .Z(n2417) );
  NAND U4147 ( .A(n2415), .B(n2414), .Z(n2416) );
  AND U4148 ( .A(n2417), .B(n2416), .Z(n2612) );
  XOR U4149 ( .A(n2613), .B(n2612), .Z(n3325) );
  NAND U4150 ( .A(n2419), .B(n2418), .Z(n2423) );
  NAND U4151 ( .A(n2421), .B(n2420), .Z(n2422) );
  AND U4152 ( .A(n2423), .B(n2422), .Z(n2774) );
  NAND U4153 ( .A(n2425), .B(n2424), .Z(n2429) );
  NAND U4154 ( .A(n2427), .B(n2426), .Z(n2428) );
  NAND U4155 ( .A(n2429), .B(n2428), .Z(n2775) );
  XNOR U4156 ( .A(n2774), .B(n2775), .Z(n2777) );
  NAND U4157 ( .A(n2431), .B(n2430), .Z(n2435) );
  NAND U4158 ( .A(n2433), .B(n2432), .Z(n2434) );
  AND U4159 ( .A(n2435), .B(n2434), .Z(n2776) );
  XOR U4160 ( .A(n2777), .B(n2776), .Z(n3323) );
  NAND U4161 ( .A(n2437), .B(n2436), .Z(n2441) );
  NAND U4162 ( .A(n2439), .B(n2438), .Z(n2440) );
  AND U4163 ( .A(n2441), .B(n2440), .Z(n2780) );
  NAND U4164 ( .A(n2443), .B(n2442), .Z(n2447) );
  NAND U4165 ( .A(n2445), .B(n2444), .Z(n2446) );
  NAND U4166 ( .A(n2447), .B(n2446), .Z(n2781) );
  XNOR U4167 ( .A(n2780), .B(n2781), .Z(n2783) );
  NAND U4168 ( .A(n2449), .B(n2448), .Z(n2453) );
  NAND U4169 ( .A(n2451), .B(n2450), .Z(n2452) );
  AND U4170 ( .A(n2453), .B(n2452), .Z(n2782) );
  XNOR U4171 ( .A(n2783), .B(n2782), .Z(n3322) );
  XNOR U4172 ( .A(n3323), .B(n3322), .Z(n3324) );
  XNOR U4173 ( .A(n3325), .B(n3324), .Z(n3305) );
  XOR U4174 ( .A(n3306), .B(n3305), .Z(n3178) );
  NANDN U4175 ( .A(n2455), .B(n2454), .Z(n2459) );
  NAND U4176 ( .A(n2457), .B(n2456), .Z(n2458) );
  AND U4177 ( .A(n2459), .B(n2458), .Z(n2592) );
  NANDN U4178 ( .A(n2461), .B(n2460), .Z(n2465) );
  NAND U4179 ( .A(n2463), .B(n2462), .Z(n2464) );
  NAND U4180 ( .A(n2465), .B(n2464), .Z(n2593) );
  XNOR U4181 ( .A(n2592), .B(n2593), .Z(n2595) );
  NANDN U4182 ( .A(n2467), .B(n2466), .Z(n2471) );
  NAND U4183 ( .A(n2469), .B(n2468), .Z(n2470) );
  AND U4184 ( .A(n2471), .B(n2470), .Z(n2594) );
  XOR U4185 ( .A(n2595), .B(n2594), .Z(n3030) );
  NANDN U4186 ( .A(n2473), .B(n2472), .Z(n2477) );
  NAND U4187 ( .A(n2475), .B(n2474), .Z(n2476) );
  AND U4188 ( .A(n2477), .B(n2476), .Z(n2677) );
  NANDN U4189 ( .A(n2479), .B(n2478), .Z(n2483) );
  NAND U4190 ( .A(n2481), .B(n2480), .Z(n2482) );
  AND U4191 ( .A(n2483), .B(n2482), .Z(n2678) );
  NAND U4192 ( .A(n2485), .B(n2484), .Z(n2489) );
  NAND U4193 ( .A(n2487), .B(n2486), .Z(n2488) );
  AND U4194 ( .A(n2489), .B(n2488), .Z(n2679) );
  XOR U4195 ( .A(n2680), .B(n2679), .Z(n3028) );
  NANDN U4196 ( .A(n2491), .B(n2490), .Z(n2495) );
  NAND U4197 ( .A(n2493), .B(n2492), .Z(n2494) );
  AND U4198 ( .A(n2495), .B(n2494), .Z(n2598) );
  NANDN U4199 ( .A(n2497), .B(n2496), .Z(n2501) );
  NAND U4200 ( .A(n2499), .B(n2498), .Z(n2500) );
  NAND U4201 ( .A(n2501), .B(n2500), .Z(n2599) );
  XNOR U4202 ( .A(n2598), .B(n2599), .Z(n2601) );
  NANDN U4203 ( .A(n2503), .B(n2502), .Z(n2507) );
  NAND U4204 ( .A(n2505), .B(n2504), .Z(n2506) );
  AND U4205 ( .A(n2507), .B(n2506), .Z(n2600) );
  XNOR U4206 ( .A(n2601), .B(n2600), .Z(n3027) );
  XNOR U4207 ( .A(n3028), .B(n3027), .Z(n3029) );
  XOR U4208 ( .A(n3030), .B(n3029), .Z(n3552) );
  NANDN U4209 ( .A(n2509), .B(n2508), .Z(n2513) );
  NANDN U4210 ( .A(n2511), .B(n2510), .Z(n2512) );
  AND U4211 ( .A(n2513), .B(n2512), .Z(n3428) );
  NANDN U4212 ( .A(n2515), .B(n2514), .Z(n2519) );
  NAND U4213 ( .A(n2517), .B(n2516), .Z(n2518) );
  AND U4214 ( .A(n2519), .B(n2518), .Z(n3021) );
  NANDN U4215 ( .A(n2521), .B(n2520), .Z(n2525) );
  NAND U4216 ( .A(n2523), .B(n2522), .Z(n2524) );
  AND U4217 ( .A(n2525), .B(n2524), .Z(n3022) );
  NAND U4218 ( .A(n2527), .B(n2526), .Z(n2531) );
  NAND U4219 ( .A(n2529), .B(n2528), .Z(n2530) );
  AND U4220 ( .A(n2531), .B(n2530), .Z(n3023) );
  XOR U4221 ( .A(n3024), .B(n3023), .Z(n3426) );
  NANDN U4222 ( .A(n2533), .B(n2532), .Z(n2537) );
  NANDN U4223 ( .A(n2535), .B(n2534), .Z(n2536) );
  AND U4224 ( .A(n2537), .B(n2536), .Z(n3425) );
  XNOR U4225 ( .A(n3426), .B(n3425), .Z(n3427) );
  XOR U4226 ( .A(n3428), .B(n3427), .Z(n3551) );
  NAND U4227 ( .A(n2539), .B(n2538), .Z(n2543) );
  NAND U4228 ( .A(n2541), .B(n2540), .Z(n2542) );
  NAND U4229 ( .A(n2543), .B(n2542), .Z(n3550) );
  XNOR U4230 ( .A(n3551), .B(n3550), .Z(n3553) );
  XOR U4231 ( .A(n3552), .B(n3553), .Z(n3177) );
  XNOR U4232 ( .A(n3178), .B(n3177), .Z(n3179) );
  XOR U4233 ( .A(n3180), .B(n3179), .Z(n3125) );
  XOR U4234 ( .A(n3126), .B(n3125), .Z(n3113) );
  XOR U4235 ( .A(n3114), .B(n3113), .Z(n3693) );
  XNOR U4236 ( .A(n3694), .B(n3693), .Z(o[1]) );
  NANDN U4237 ( .A(n2545), .B(n2544), .Z(n2549) );
  NANDN U4238 ( .A(n2547), .B(n2546), .Z(n2548) );
  AND U4239 ( .A(n2549), .B(n2548), .Z(n3901) );
  NAND U4240 ( .A(n2551), .B(n2550), .Z(n2555) );
  NANDN U4241 ( .A(n2553), .B(n2552), .Z(n2554) );
  AND U4242 ( .A(n2555), .B(n2554), .Z(n4230) );
  NAND U4243 ( .A(n2557), .B(n2556), .Z(n2561) );
  NAND U4244 ( .A(n2559), .B(n2558), .Z(n2560) );
  AND U4245 ( .A(n2561), .B(n2560), .Z(n4228) );
  NANDN U4246 ( .A(n2563), .B(n2562), .Z(n2567) );
  NAND U4247 ( .A(n2565), .B(n2564), .Z(n2566) );
  NAND U4248 ( .A(n2567), .B(n2566), .Z(n3819) );
  NANDN U4249 ( .A(n2569), .B(n2568), .Z(n2573) );
  NAND U4250 ( .A(n2571), .B(n2570), .Z(n2572) );
  NAND U4251 ( .A(n2573), .B(n2572), .Z(n3817) );
  NANDN U4252 ( .A(n2575), .B(n2574), .Z(n2579) );
  NAND U4253 ( .A(n2577), .B(n2576), .Z(n2578) );
  NAND U4254 ( .A(n2579), .B(n2578), .Z(n3816) );
  XNOR U4255 ( .A(n4228), .B(n4227), .Z(n4229) );
  XOR U4256 ( .A(n4230), .B(n4229), .Z(n3900) );
  XOR U4257 ( .A(n3901), .B(n3900), .Z(n3903) );
  NANDN U4258 ( .A(n2581), .B(n2580), .Z(n2585) );
  NAND U4259 ( .A(n2583), .B(n2582), .Z(n2584) );
  NAND U4260 ( .A(n2585), .B(n2584), .Z(n3780) );
  NANDN U4261 ( .A(n2587), .B(n2586), .Z(n2591) );
  NAND U4262 ( .A(n2589), .B(n2588), .Z(n2590) );
  NAND U4263 ( .A(n2591), .B(n2590), .Z(n3778) );
  NANDN U4264 ( .A(n2593), .B(n2592), .Z(n2597) );
  NAND U4265 ( .A(n2595), .B(n2594), .Z(n2596) );
  NAND U4266 ( .A(n2597), .B(n2596), .Z(n3777) );
  NANDN U4267 ( .A(n2599), .B(n2598), .Z(n2603) );
  NAND U4268 ( .A(n2601), .B(n2600), .Z(n2602) );
  NAND U4269 ( .A(n2603), .B(n2602), .Z(n3783) );
  NANDN U4270 ( .A(n2605), .B(n2604), .Z(n2609) );
  NAND U4271 ( .A(n2607), .B(n2606), .Z(n2608) );
  AND U4272 ( .A(n2609), .B(n2608), .Z(n3785) );
  NANDN U4273 ( .A(n2611), .B(n2610), .Z(n2615) );
  NAND U4274 ( .A(n2613), .B(n2612), .Z(n2614) );
  AND U4275 ( .A(n2615), .B(n2614), .Z(n3784) );
  XNOR U4276 ( .A(n3785), .B(n3784), .Z(n2616) );
  XOR U4277 ( .A(n3783), .B(n2616), .Z(n3734) );
  NAND U4278 ( .A(n2618), .B(n2617), .Z(n2622) );
  NAND U4279 ( .A(n2620), .B(n2619), .Z(n2621) );
  AND U4280 ( .A(n2622), .B(n2621), .Z(n3735) );
  XNOR U4281 ( .A(n3734), .B(n3735), .Z(n3737) );
  XOR U4282 ( .A(n3736), .B(n3737), .Z(n4028) );
  NAND U4283 ( .A(n2624), .B(n2623), .Z(n2628) );
  NAND U4284 ( .A(n2626), .B(n2625), .Z(n2627) );
  NAND U4285 ( .A(n2628), .B(n2627), .Z(n4151) );
  NAND U4286 ( .A(n2630), .B(n2629), .Z(n2634) );
  NAND U4287 ( .A(n2632), .B(n2631), .Z(n2633) );
  NAND U4288 ( .A(n2634), .B(n2633), .Z(n4153) );
  NAND U4289 ( .A(n2636), .B(n2635), .Z(n2640) );
  NAND U4290 ( .A(n2638), .B(n2637), .Z(n2639) );
  NAND U4291 ( .A(n2640), .B(n2639), .Z(n4152) );
  NAND U4292 ( .A(n2642), .B(n2641), .Z(n2646) );
  NAND U4293 ( .A(n2644), .B(n2643), .Z(n2645) );
  AND U4294 ( .A(n2646), .B(n2645), .Z(n3793) );
  NANDN U4295 ( .A(n2648), .B(n2647), .Z(n2652) );
  NAND U4296 ( .A(n2650), .B(n2649), .Z(n2651) );
  AND U4297 ( .A(n2652), .B(n2651), .Z(n3768) );
  NANDN U4298 ( .A(n2654), .B(n2653), .Z(n2658) );
  NAND U4299 ( .A(n2656), .B(n2655), .Z(n2657) );
  NAND U4300 ( .A(n2658), .B(n2657), .Z(n3766) );
  NAND U4301 ( .A(n2660), .B(n2659), .Z(n2664) );
  NAND U4302 ( .A(n2662), .B(n2661), .Z(n2663) );
  NAND U4303 ( .A(n2664), .B(n2663), .Z(n3765) );
  XOR U4304 ( .A(n3768), .B(n3767), .Z(n3792) );
  XNOR U4305 ( .A(n3793), .B(n3792), .Z(n3794) );
  XOR U4306 ( .A(n3795), .B(n3794), .Z(n4027) );
  XOR U4307 ( .A(n4028), .B(n4027), .Z(n4030) );
  NAND U4308 ( .A(n2666), .B(n2665), .Z(n2670) );
  NAND U4309 ( .A(n2668), .B(n2667), .Z(n2669) );
  AND U4310 ( .A(n2670), .B(n2669), .Z(n3756) );
  NAND U4311 ( .A(n2672), .B(n2671), .Z(n2676) );
  NAND U4312 ( .A(n2674), .B(n2673), .Z(n2675) );
  AND U4313 ( .A(n2676), .B(n2675), .Z(n3754) );
  NAND U4314 ( .A(n2678), .B(n2677), .Z(n2682) );
  NAND U4315 ( .A(n2680), .B(n2679), .Z(n2681) );
  NAND U4316 ( .A(n2682), .B(n2681), .Z(n3753) );
  XNOR U4317 ( .A(n3754), .B(n3753), .Z(n3755) );
  XOR U4318 ( .A(n3756), .B(n3755), .Z(n3824) );
  NAND U4319 ( .A(n2684), .B(n2683), .Z(n2688) );
  NAND U4320 ( .A(n2686), .B(n2685), .Z(n2687) );
  AND U4321 ( .A(n2688), .B(n2687), .Z(n3823) );
  NANDN U4322 ( .A(n2690), .B(n2689), .Z(n2694) );
  NAND U4323 ( .A(n2692), .B(n2691), .Z(n2693) );
  AND U4324 ( .A(n2694), .B(n2693), .Z(n3890) );
  NANDN U4325 ( .A(n2696), .B(n2695), .Z(n2700) );
  NAND U4326 ( .A(n2698), .B(n2697), .Z(n2699) );
  AND U4327 ( .A(n2700), .B(n2699), .Z(n3888) );
  NANDN U4328 ( .A(n2702), .B(n2701), .Z(n2706) );
  NAND U4329 ( .A(n2704), .B(n2703), .Z(n2705) );
  NAND U4330 ( .A(n2706), .B(n2705), .Z(n3887) );
  XNOR U4331 ( .A(n3888), .B(n3887), .Z(n3889) );
  XOR U4332 ( .A(n3890), .B(n3889), .Z(n3822) );
  XNOR U4333 ( .A(n3823), .B(n3822), .Z(n3825) );
  XOR U4334 ( .A(n3824), .B(n3825), .Z(n4029) );
  XOR U4335 ( .A(n4030), .B(n4029), .Z(n3902) );
  XOR U4336 ( .A(n3903), .B(n3902), .Z(n3719) );
  NAND U4337 ( .A(n2708), .B(n2707), .Z(n2712) );
  NAND U4338 ( .A(n2710), .B(n2709), .Z(n2711) );
  AND U4339 ( .A(n2712), .B(n2711), .Z(n4046) );
  NAND U4340 ( .A(n2717), .B(n2716), .Z(n2721) );
  NAND U4341 ( .A(n2719), .B(n2718), .Z(n2720) );
  AND U4342 ( .A(n2721), .B(n2720), .Z(n4116) );
  XNOR U4343 ( .A(n4116), .B(n4115), .Z(n2725) );
  XNOR U4344 ( .A(n4114), .B(n2725), .Z(n4200) );
  NANDN U4345 ( .A(n2727), .B(n2726), .Z(n2731) );
  NAND U4346 ( .A(n2729), .B(n2728), .Z(n2730) );
  AND U4347 ( .A(n2731), .B(n2730), .Z(n4198) );
  NANDN U4348 ( .A(n2733), .B(n2732), .Z(n2737) );
  NAND U4349 ( .A(n2735), .B(n2734), .Z(n2736) );
  AND U4350 ( .A(n2737), .B(n2736), .Z(n4248) );
  NANDN U4351 ( .A(n2739), .B(n2738), .Z(n2743) );
  NAND U4352 ( .A(n2741), .B(n2740), .Z(n2742) );
  AND U4353 ( .A(n2743), .B(n2742), .Z(n4246) );
  NANDN U4354 ( .A(n2745), .B(n2744), .Z(n2749) );
  NAND U4355 ( .A(n2747), .B(n2746), .Z(n2748) );
  NAND U4356 ( .A(n2749), .B(n2748), .Z(n4245) );
  XNOR U4357 ( .A(n4246), .B(n4245), .Z(n4247) );
  XOR U4358 ( .A(n4248), .B(n4247), .Z(n4197) );
  XNOR U4359 ( .A(n4198), .B(n4197), .Z(n4199) );
  XOR U4360 ( .A(n4200), .B(n4199), .Z(n4045) );
  XNOR U4361 ( .A(n4046), .B(n4045), .Z(n4048) );
  NAND U4362 ( .A(n2751), .B(n2750), .Z(n2755) );
  NAND U4363 ( .A(n2753), .B(n2752), .Z(n2754) );
  NAND U4364 ( .A(n2755), .B(n2754), .Z(n3970) );
  NAND U4365 ( .A(n2757), .B(n2756), .Z(n2761) );
  NAND U4366 ( .A(n2759), .B(n2758), .Z(n2760) );
  NAND U4367 ( .A(n2761), .B(n2760), .Z(n3968) );
  NAND U4368 ( .A(n2763), .B(n2762), .Z(n2767) );
  NAND U4369 ( .A(n2765), .B(n2764), .Z(n2766) );
  NAND U4370 ( .A(n2767), .B(n2766), .Z(n3967) );
  NANDN U4371 ( .A(n2769), .B(n2768), .Z(n2773) );
  NAND U4372 ( .A(n2771), .B(n2770), .Z(n2772) );
  AND U4373 ( .A(n2773), .B(n2772), .Z(n4204) );
  NANDN U4374 ( .A(n2775), .B(n2774), .Z(n2779) );
  NAND U4375 ( .A(n2777), .B(n2776), .Z(n2778) );
  AND U4376 ( .A(n2779), .B(n2778), .Z(n4260) );
  NANDN U4377 ( .A(n2781), .B(n2780), .Z(n2785) );
  NAND U4378 ( .A(n2783), .B(n2782), .Z(n2784) );
  AND U4379 ( .A(n2785), .B(n2784), .Z(n4258) );
  NANDN U4380 ( .A(n2787), .B(n2786), .Z(n2791) );
  NAND U4381 ( .A(n2789), .B(n2788), .Z(n2790) );
  NAND U4382 ( .A(n2791), .B(n2790), .Z(n4257) );
  XNOR U4383 ( .A(n4258), .B(n4257), .Z(n4259) );
  XOR U4384 ( .A(n4260), .B(n4259), .Z(n4203) );
  XNOR U4385 ( .A(n4204), .B(n4203), .Z(n4206) );
  XOR U4386 ( .A(n4205), .B(n4206), .Z(n4047) );
  XNOR U4387 ( .A(n4048), .B(n4047), .Z(n4092) );
  NAND U4388 ( .A(n2793), .B(n2792), .Z(n2797) );
  NAND U4389 ( .A(n2795), .B(n2794), .Z(n2796) );
  AND U4390 ( .A(n2797), .B(n2796), .Z(n4130) );
  NAND U4391 ( .A(n2799), .B(n2798), .Z(n2803) );
  NAND U4392 ( .A(n2801), .B(n2800), .Z(n2802) );
  AND U4393 ( .A(n2803), .B(n2802), .Z(n4128) );
  NAND U4394 ( .A(n2805), .B(n2804), .Z(n2809) );
  NAND U4395 ( .A(n2807), .B(n2806), .Z(n2808) );
  NAND U4396 ( .A(n2809), .B(n2808), .Z(n4127) );
  XNOR U4397 ( .A(n4128), .B(n4127), .Z(n4129) );
  XNOR U4398 ( .A(n4130), .B(n4129), .Z(n3955) );
  NANDN U4399 ( .A(n2811), .B(n2810), .Z(n2815) );
  NANDN U4400 ( .A(n2813), .B(n2812), .Z(n2814) );
  NAND U4401 ( .A(n2815), .B(n2814), .Z(n3956) );
  XNOR U4402 ( .A(n3955), .B(n3956), .Z(n3958) );
  NAND U4403 ( .A(n2817), .B(n2816), .Z(n2821) );
  NAND U4404 ( .A(n2819), .B(n2818), .Z(n2820) );
  AND U4405 ( .A(n2821), .B(n2820), .Z(n3774) );
  XNOR U4406 ( .A(n3772), .B(n3771), .Z(n3773) );
  XNOR U4407 ( .A(n3774), .B(n3773), .Z(n3957) );
  XOR U4408 ( .A(n3958), .B(n3957), .Z(n4058) );
  NAND U4409 ( .A(n2829), .B(n2828), .Z(n2833) );
  NANDN U4410 ( .A(n2831), .B(n2830), .Z(n2832) );
  AND U4411 ( .A(n2833), .B(n2832), .Z(n4057) );
  XNOR U4412 ( .A(n4058), .B(n4057), .Z(n4060) );
  NANDN U4413 ( .A(n2835), .B(n2834), .Z(n2839) );
  NAND U4414 ( .A(n2837), .B(n2836), .Z(n2838) );
  AND U4415 ( .A(n2839), .B(n2838), .Z(n4242) );
  NANDN U4416 ( .A(n2841), .B(n2840), .Z(n2845) );
  NAND U4417 ( .A(n2843), .B(n2842), .Z(n2844) );
  AND U4418 ( .A(n2845), .B(n2844), .Z(n4240) );
  NANDN U4419 ( .A(n2847), .B(n2846), .Z(n2851) );
  NAND U4420 ( .A(n2849), .B(n2848), .Z(n2850) );
  NAND U4421 ( .A(n2851), .B(n2850), .Z(n4239) );
  XNOR U4422 ( .A(n4240), .B(n4239), .Z(n4241) );
  XOR U4423 ( .A(n4242), .B(n4241), .Z(n4265) );
  NANDN U4424 ( .A(n2853), .B(n2852), .Z(n2857) );
  NANDN U4425 ( .A(n2855), .B(n2854), .Z(n2856) );
  AND U4426 ( .A(n2857), .B(n2856), .Z(n4264) );
  NAND U4427 ( .A(n2859), .B(n2858), .Z(n2863) );
  NAND U4428 ( .A(n2861), .B(n2860), .Z(n2862) );
  AND U4429 ( .A(n2863), .B(n2862), .Z(n4157) );
  NAND U4430 ( .A(n2865), .B(n2864), .Z(n2869) );
  NAND U4431 ( .A(n2867), .B(n2866), .Z(n2868) );
  NAND U4432 ( .A(n2869), .B(n2868), .Z(n4155) );
  NAND U4433 ( .A(n2871), .B(n2870), .Z(n2875) );
  NAND U4434 ( .A(n2873), .B(n2872), .Z(n2874) );
  NAND U4435 ( .A(n2875), .B(n2874), .Z(n4154) );
  XOR U4436 ( .A(n4157), .B(n4156), .Z(n4263) );
  XNOR U4437 ( .A(n4264), .B(n4263), .Z(n4266) );
  XOR U4438 ( .A(n4265), .B(n4266), .Z(n4059) );
  XNOR U4439 ( .A(n4060), .B(n4059), .Z(n4091) );
  NAND U4440 ( .A(n2877), .B(n2876), .Z(n2881) );
  NAND U4441 ( .A(n2879), .B(n2878), .Z(n2880) );
  NAND U4442 ( .A(n2881), .B(n2880), .Z(n4090) );
  XOR U4443 ( .A(n4092), .B(n4093), .Z(n3716) );
  NANDN U4444 ( .A(n2883), .B(n2882), .Z(n2887) );
  NAND U4445 ( .A(n2885), .B(n2884), .Z(n2886) );
  AND U4446 ( .A(n2887), .B(n2886), .Z(n3907) );
  NAND U4447 ( .A(n2889), .B(n2888), .Z(n2893) );
  NAND U4448 ( .A(n2891), .B(n2890), .Z(n2892) );
  AND U4449 ( .A(n2893), .B(n2892), .Z(n3830) );
  NANDN U4450 ( .A(n2895), .B(n2894), .Z(n2899) );
  NANDN U4451 ( .A(n2897), .B(n2896), .Z(n2898) );
  AND U4452 ( .A(n2899), .B(n2898), .Z(n3982) );
  NAND U4453 ( .A(n2901), .B(n2900), .Z(n2905) );
  NAND U4454 ( .A(n2903), .B(n2902), .Z(n2904) );
  AND U4455 ( .A(n2905), .B(n2904), .Z(n3980) );
  NAND U4456 ( .A(n2907), .B(n2906), .Z(n2911) );
  NAND U4457 ( .A(n2909), .B(n2908), .Z(n2910) );
  NAND U4458 ( .A(n2911), .B(n2910), .Z(n3979) );
  XNOR U4459 ( .A(n3980), .B(n3979), .Z(n3981) );
  XNOR U4460 ( .A(n3982), .B(n3981), .Z(n3829) );
  XNOR U4461 ( .A(n3830), .B(n3829), .Z(n3832) );
  NANDN U4462 ( .A(n2913), .B(n2912), .Z(n2917) );
  NAND U4463 ( .A(n2915), .B(n2914), .Z(n2916) );
  AND U4464 ( .A(n2917), .B(n2916), .Z(n3945) );
  NANDN U4465 ( .A(n2919), .B(n2918), .Z(n2923) );
  NAND U4466 ( .A(n2921), .B(n2920), .Z(n2922) );
  AND U4467 ( .A(n2923), .B(n2922), .Z(n3943) );
  NAND U4468 ( .A(n2925), .B(n2924), .Z(n2929) );
  NAND U4469 ( .A(n2927), .B(n2926), .Z(n2928) );
  NAND U4470 ( .A(n2929), .B(n2928), .Z(n3942) );
  XNOR U4471 ( .A(n3943), .B(n3942), .Z(n3944) );
  XNOR U4472 ( .A(n3945), .B(n3944), .Z(n3831) );
  XOR U4473 ( .A(n3832), .B(n3831), .Z(n3906) );
  XOR U4474 ( .A(n3907), .B(n3906), .Z(n3909) );
  NANDN U4475 ( .A(n2931), .B(n2930), .Z(n2935) );
  NANDN U4476 ( .A(n2933), .B(n2932), .Z(n2934) );
  AND U4477 ( .A(n2935), .B(n2934), .Z(n3872) );
  NANDN U4478 ( .A(n2937), .B(n2936), .Z(n2941) );
  NAND U4479 ( .A(n2939), .B(n2938), .Z(n2940) );
  NAND U4480 ( .A(n2941), .B(n2940), .Z(n3884) );
  NANDN U4481 ( .A(n2943), .B(n2942), .Z(n2947) );
  NAND U4482 ( .A(n2945), .B(n2944), .Z(n2946) );
  NAND U4483 ( .A(n2947), .B(n2946), .Z(n3882) );
  NANDN U4484 ( .A(n2949), .B(n2948), .Z(n2953) );
  NAND U4485 ( .A(n2951), .B(n2950), .Z(n2952) );
  NAND U4486 ( .A(n2953), .B(n2952), .Z(n3881) );
  NANDN U4487 ( .A(n2955), .B(n2954), .Z(n2959) );
  NAND U4488 ( .A(n2957), .B(n2956), .Z(n2958) );
  NAND U4489 ( .A(n2959), .B(n2958), .Z(n4254) );
  NANDN U4490 ( .A(n2961), .B(n2960), .Z(n2965) );
  NAND U4491 ( .A(n2963), .B(n2962), .Z(n2964) );
  NAND U4492 ( .A(n2965), .B(n2964), .Z(n4252) );
  NANDN U4493 ( .A(n2967), .B(n2966), .Z(n2971) );
  NAND U4494 ( .A(n2969), .B(n2968), .Z(n2970) );
  NAND U4495 ( .A(n2971), .B(n2970), .Z(n4251) );
  XOR U4496 ( .A(n3870), .B(n3869), .Z(n3871) );
  XOR U4497 ( .A(n3872), .B(n3871), .Z(n4011) );
  NANDN U4498 ( .A(n2973), .B(n2972), .Z(n2977) );
  NAND U4499 ( .A(n2975), .B(n2974), .Z(n2976) );
  NAND U4500 ( .A(n2977), .B(n2976), .Z(n4218) );
  NANDN U4501 ( .A(n2982), .B(n2981), .Z(n2986) );
  ANDN U4502 ( .B(n2982), .A(n2981), .Z(n2983) );
  OR U4503 ( .A(n2984), .B(n2983), .Z(n2985) );
  AND U4504 ( .A(n2986), .B(n2985), .Z(n4215) );
  XNOR U4505 ( .A(n4216), .B(n4215), .Z(n4217) );
  NANDN U4506 ( .A(n2988), .B(n2987), .Z(n2992) );
  NAND U4507 ( .A(n2990), .B(n2989), .Z(n2991) );
  NAND U4508 ( .A(n2992), .B(n2991), .Z(n4212) );
  NANDN U4509 ( .A(n2994), .B(n2993), .Z(n2998) );
  NAND U4510 ( .A(n2996), .B(n2995), .Z(n2997) );
  NAND U4511 ( .A(n2998), .B(n2997), .Z(n4210) );
  NANDN U4512 ( .A(n3000), .B(n2999), .Z(n3004) );
  NAND U4513 ( .A(n3002), .B(n3001), .Z(n3003) );
  NAND U4514 ( .A(n3004), .B(n3003), .Z(n4209) );
  XNOR U4515 ( .A(n3855), .B(n3853), .Z(n3008) );
  XOR U4516 ( .A(n3854), .B(n3008), .Z(n4009) );
  NAND U4517 ( .A(n3010), .B(n3009), .Z(n3014) );
  NAND U4518 ( .A(n3012), .B(n3011), .Z(n3013) );
  NAND U4519 ( .A(n3014), .B(n3013), .Z(n3976) );
  NANDN U4520 ( .A(n3016), .B(n3015), .Z(n3020) );
  NAND U4521 ( .A(n3018), .B(n3017), .Z(n3019) );
  NAND U4522 ( .A(n3020), .B(n3019), .Z(n3974) );
  NAND U4523 ( .A(n3022), .B(n3021), .Z(n3026) );
  NAND U4524 ( .A(n3024), .B(n3023), .Z(n3025) );
  NAND U4525 ( .A(n3026), .B(n3025), .Z(n3973) );
  NANDN U4526 ( .A(n3028), .B(n3027), .Z(n3032) );
  NANDN U4527 ( .A(n3030), .B(n3029), .Z(n3031) );
  NAND U4528 ( .A(n3032), .B(n3031), .Z(n3937) );
  NANDN U4529 ( .A(n3034), .B(n3033), .Z(n3038) );
  NAND U4530 ( .A(n3036), .B(n3035), .Z(n3037) );
  AND U4531 ( .A(n3038), .B(n3037), .Z(n4108) );
  NAND U4532 ( .A(n3040), .B(n3039), .Z(n3044) );
  NAND U4533 ( .A(n3042), .B(n3041), .Z(n3043) );
  NAND U4534 ( .A(n3044), .B(n3043), .Z(n4106) );
  NAND U4535 ( .A(n3046), .B(n3045), .Z(n3050) );
  NAND U4536 ( .A(n3048), .B(n3047), .Z(n3049) );
  NAND U4537 ( .A(n3050), .B(n3049), .Z(n4105) );
  XOR U4538 ( .A(n4108), .B(n4107), .Z(n3936) );
  XOR U4539 ( .A(n3938), .B(n3939), .Z(n4010) );
  XOR U4540 ( .A(n4009), .B(n4010), .Z(n4012) );
  XOR U4541 ( .A(n4011), .B(n4012), .Z(n3908) );
  XOR U4542 ( .A(n3909), .B(n3908), .Z(n3717) );
  XOR U4543 ( .A(n3716), .B(n3717), .Z(n3718) );
  XNOR U4544 ( .A(n3719), .B(n3718), .Z(n3699) );
  NAND U4545 ( .A(n3052), .B(n3051), .Z(n3056) );
  NAND U4546 ( .A(n3054), .B(n3053), .Z(n3055) );
  AND U4547 ( .A(n3056), .B(n3055), .Z(n3713) );
  NANDN U4548 ( .A(n3058), .B(n3057), .Z(n3062) );
  NANDN U4549 ( .A(n3060), .B(n3059), .Z(n3061) );
  AND U4550 ( .A(n3062), .B(n3061), .Z(n3711) );
  NANDN U4551 ( .A(n3064), .B(n3063), .Z(n3068) );
  NAND U4552 ( .A(n3066), .B(n3065), .Z(n3067) );
  NAND U4553 ( .A(n3068), .B(n3067), .Z(n3710) );
  XNOR U4554 ( .A(n3711), .B(n3710), .Z(n3712) );
  XOR U4555 ( .A(n3713), .B(n3712), .Z(n3698) );
  NANDN U4556 ( .A(n3070), .B(n3069), .Z(n3074) );
  NAND U4557 ( .A(n3072), .B(n3071), .Z(n3073) );
  AND U4558 ( .A(n3074), .B(n3073), .Z(n4099) );
  NANDN U4559 ( .A(n3076), .B(n3075), .Z(n3080) );
  NANDN U4560 ( .A(n3078), .B(n3077), .Z(n3079) );
  AND U4561 ( .A(n3080), .B(n3079), .Z(n4097) );
  NANDN U4562 ( .A(n3082), .B(n3081), .Z(n3086) );
  NANDN U4563 ( .A(n3084), .B(n3083), .Z(n3085) );
  NAND U4564 ( .A(n3086), .B(n3085), .Z(n4096) );
  XNOR U4565 ( .A(n4097), .B(n4096), .Z(n4098) );
  XNOR U4566 ( .A(n4099), .B(n4098), .Z(n4023) );
  NAND U4567 ( .A(n3088), .B(n3087), .Z(n3092) );
  NAND U4568 ( .A(n3090), .B(n3089), .Z(n3091) );
  NAND U4569 ( .A(n3092), .B(n3091), .Z(n4021) );
  NAND U4570 ( .A(n3094), .B(n3093), .Z(n3098) );
  NAND U4571 ( .A(n3096), .B(n3095), .Z(n3097) );
  AND U4572 ( .A(n3098), .B(n3097), .Z(n4194) );
  NANDN U4573 ( .A(n3100), .B(n3099), .Z(n3104) );
  NAND U4574 ( .A(n3102), .B(n3101), .Z(n3103) );
  AND U4575 ( .A(n3104), .B(n3103), .Z(n4191) );
  NANDN U4576 ( .A(n3106), .B(n3105), .Z(n3110) );
  NANDN U4577 ( .A(n3108), .B(n3107), .Z(n3109) );
  NAND U4578 ( .A(n3110), .B(n3109), .Z(n4192) );
  XNOR U4579 ( .A(n4191), .B(n4192), .Z(n4193) );
  XOR U4580 ( .A(n4194), .B(n4193), .Z(n4022) );
  XNOR U4581 ( .A(n4023), .B(n4024), .Z(n3700) );
  XOR U4582 ( .A(n3701), .B(n3700), .Z(n4083) );
  NAND U4583 ( .A(n3112), .B(n3111), .Z(n3116) );
  NAND U4584 ( .A(n3114), .B(n3113), .Z(n3115) );
  AND U4585 ( .A(n3116), .B(n3115), .Z(n4085) );
  NANDN U4586 ( .A(n3118), .B(n3117), .Z(n3122) );
  NANDN U4587 ( .A(n3120), .B(n3119), .Z(n3121) );
  AND U4588 ( .A(n3122), .B(n3121), .Z(n4084) );
  XNOR U4589 ( .A(n4085), .B(n4084), .Z(n4087) );
  NAND U4590 ( .A(n3124), .B(n3123), .Z(n3128) );
  NAND U4591 ( .A(n3126), .B(n3125), .Z(n3127) );
  NAND U4592 ( .A(n3128), .B(n3127), .Z(n4270) );
  NAND U4593 ( .A(n3130), .B(n3129), .Z(n3134) );
  NAND U4594 ( .A(n3132), .B(n3131), .Z(n3133) );
  NAND U4595 ( .A(n3134), .B(n3133), .Z(n3991) );
  NANDN U4596 ( .A(n3136), .B(n3135), .Z(n3140) );
  NAND U4597 ( .A(n3138), .B(n3137), .Z(n3139) );
  AND U4598 ( .A(n3140), .B(n3139), .Z(n4072) );
  NAND U4599 ( .A(n3142), .B(n3141), .Z(n3146) );
  NAND U4600 ( .A(n3144), .B(n3143), .Z(n3145) );
  AND U4601 ( .A(n3146), .B(n3145), .Z(n4070) );
  NANDN U4602 ( .A(n3148), .B(n3147), .Z(n3152) );
  NANDN U4603 ( .A(n3150), .B(n3149), .Z(n3151) );
  AND U4604 ( .A(n3152), .B(n3151), .Z(n4069) );
  XNOR U4605 ( .A(n4070), .B(n4069), .Z(n4071) );
  XOR U4606 ( .A(n4072), .B(n4071), .Z(n3992) );
  XOR U4607 ( .A(n3991), .B(n3992), .Z(n3994) );
  NAND U4608 ( .A(n3154), .B(n3153), .Z(n3158) );
  NAND U4609 ( .A(n3156), .B(n3155), .Z(n3157) );
  AND U4610 ( .A(n3158), .B(n3157), .Z(n4182) );
  NAND U4611 ( .A(n3160), .B(n3159), .Z(n3164) );
  NAND U4612 ( .A(n3162), .B(n3161), .Z(n3163) );
  AND U4613 ( .A(n3164), .B(n3163), .Z(n4180) );
  NAND U4614 ( .A(n3166), .B(n3165), .Z(n3170) );
  NAND U4615 ( .A(n3168), .B(n3167), .Z(n3169) );
  NAND U4616 ( .A(n3170), .B(n3169), .Z(n4179) );
  XNOR U4617 ( .A(n4180), .B(n4179), .Z(n4181) );
  XNOR U4618 ( .A(n4182), .B(n4181), .Z(n3993) );
  XOR U4619 ( .A(n3994), .B(n3993), .Z(n3705) );
  NAND U4620 ( .A(n3172), .B(n3171), .Z(n3176) );
  NAND U4621 ( .A(n3174), .B(n3173), .Z(n3175) );
  AND U4622 ( .A(n3176), .B(n3175), .Z(n4170) );
  NANDN U4623 ( .A(n3178), .B(n3177), .Z(n3182) );
  NAND U4624 ( .A(n3180), .B(n3179), .Z(n3181) );
  AND U4625 ( .A(n3182), .B(n3181), .Z(n4168) );
  NANDN U4626 ( .A(n3184), .B(n3183), .Z(n3188) );
  NAND U4627 ( .A(n3186), .B(n3185), .Z(n3187) );
  AND U4628 ( .A(n3188), .B(n3187), .Z(n4176) );
  NAND U4629 ( .A(n3190), .B(n3189), .Z(n3194) );
  NAND U4630 ( .A(n3192), .B(n3191), .Z(n3193) );
  AND U4631 ( .A(n3194), .B(n3193), .Z(n4174) );
  NAND U4632 ( .A(n3196), .B(n3195), .Z(n3200) );
  NAND U4633 ( .A(n3198), .B(n3197), .Z(n3199) );
  NAND U4634 ( .A(n3200), .B(n3199), .Z(n4173) );
  XNOR U4635 ( .A(n4174), .B(n4173), .Z(n4175) );
  XOR U4636 ( .A(n4176), .B(n4175), .Z(n4167) );
  XOR U4637 ( .A(n4168), .B(n4167), .Z(n4169) );
  XOR U4638 ( .A(n4170), .B(n4169), .Z(n3704) );
  XNOR U4639 ( .A(n3705), .B(n3704), .Z(n3707) );
  NAND U4640 ( .A(n3202), .B(n3201), .Z(n3206) );
  NAND U4641 ( .A(n3204), .B(n3203), .Z(n3205) );
  AND U4642 ( .A(n3206), .B(n3205), .Z(n4066) );
  NANDN U4643 ( .A(n3208), .B(n3207), .Z(n3212) );
  NANDN U4644 ( .A(n3210), .B(n3209), .Z(n3211) );
  AND U4645 ( .A(n3212), .B(n3211), .Z(n4063) );
  NANDN U4646 ( .A(n3214), .B(n3213), .Z(n3218) );
  NAND U4647 ( .A(n3216), .B(n3215), .Z(n3217) );
  NAND U4648 ( .A(n3218), .B(n3217), .Z(n4064) );
  XNOR U4649 ( .A(n4063), .B(n4064), .Z(n4065) );
  XOR U4650 ( .A(n4066), .B(n4065), .Z(n4018) );
  NANDN U4651 ( .A(n3220), .B(n3219), .Z(n3224) );
  NANDN U4652 ( .A(n3222), .B(n3221), .Z(n3223) );
  AND U4653 ( .A(n3224), .B(n3223), .Z(n4036) );
  NANDN U4654 ( .A(n3226), .B(n3225), .Z(n3230) );
  NANDN U4655 ( .A(n3228), .B(n3227), .Z(n3229) );
  AND U4656 ( .A(n3230), .B(n3229), .Z(n4033) );
  NANDN U4657 ( .A(n3232), .B(n3231), .Z(n3236) );
  NANDN U4658 ( .A(n3234), .B(n3233), .Z(n3235) );
  NAND U4659 ( .A(n3236), .B(n3235), .Z(n4034) );
  XNOR U4660 ( .A(n4033), .B(n4034), .Z(n4035) );
  XNOR U4661 ( .A(n4036), .B(n4035), .Z(n4016) );
  NAND U4662 ( .A(n3238), .B(n3237), .Z(n3242) );
  NAND U4663 ( .A(n3240), .B(n3239), .Z(n3241) );
  NAND U4664 ( .A(n3242), .B(n3241), .Z(n4015) );
  XOR U4665 ( .A(n3707), .B(n3706), .Z(n4269) );
  NAND U4666 ( .A(n3244), .B(n3243), .Z(n3248) );
  NANDN U4667 ( .A(n3246), .B(n3245), .Z(n3247) );
  AND U4668 ( .A(n3248), .B(n3247), .Z(n3750) );
  NANDN U4669 ( .A(n3250), .B(n3249), .Z(n3254) );
  NANDN U4670 ( .A(n3252), .B(n3251), .Z(n3253) );
  AND U4671 ( .A(n3254), .B(n3253), .Z(n3748) );
  NANDN U4672 ( .A(n3256), .B(n3255), .Z(n3260) );
  NANDN U4673 ( .A(n3258), .B(n3257), .Z(n3259) );
  NAND U4674 ( .A(n3260), .B(n3259), .Z(n3747) );
  XNOR U4675 ( .A(n3748), .B(n3747), .Z(n3749) );
  XNOR U4676 ( .A(n3750), .B(n3749), .Z(n4186) );
  NAND U4677 ( .A(n3262), .B(n3261), .Z(n3266) );
  NANDN U4678 ( .A(n3264), .B(n3263), .Z(n3265) );
  AND U4679 ( .A(n3266), .B(n3265), .Z(n3744) );
  NAND U4680 ( .A(n3268), .B(n3267), .Z(n3272) );
  NANDN U4681 ( .A(n3270), .B(n3269), .Z(n3271) );
  AND U4682 ( .A(n3272), .B(n3271), .Z(n3742) );
  NANDN U4683 ( .A(n3274), .B(n3273), .Z(n3278) );
  NAND U4684 ( .A(n3276), .B(n3275), .Z(n3277) );
  NAND U4685 ( .A(n3278), .B(n3277), .Z(n3741) );
  XNOR U4686 ( .A(n3742), .B(n3741), .Z(n3743) );
  XNOR U4687 ( .A(n3744), .B(n3743), .Z(n4185) );
  XOR U4688 ( .A(n4186), .B(n4185), .Z(n4188) );
  NANDN U4689 ( .A(n3280), .B(n3279), .Z(n3284) );
  NANDN U4690 ( .A(n3282), .B(n3281), .Z(n3283) );
  AND U4691 ( .A(n3284), .B(n3283), .Z(n3850) );
  NANDN U4692 ( .A(n3286), .B(n3285), .Z(n3290) );
  NANDN U4693 ( .A(n3288), .B(n3287), .Z(n3289) );
  AND U4694 ( .A(n3290), .B(n3289), .Z(n3848) );
  NANDN U4695 ( .A(n3292), .B(n3291), .Z(n3296) );
  NANDN U4696 ( .A(n3294), .B(n3293), .Z(n3295) );
  NAND U4697 ( .A(n3296), .B(n3295), .Z(n3847) );
  XNOR U4698 ( .A(n3848), .B(n3847), .Z(n3849) );
  XNOR U4699 ( .A(n3850), .B(n3849), .Z(n4187) );
  XOR U4700 ( .A(n4188), .B(n4187), .Z(n3919) );
  NAND U4701 ( .A(n3298), .B(n3297), .Z(n3302) );
  NAND U4702 ( .A(n3300), .B(n3299), .Z(n3301) );
  AND U4703 ( .A(n3302), .B(n3301), .Z(n4054) );
  NAND U4704 ( .A(n3304), .B(n3303), .Z(n3308) );
  NAND U4705 ( .A(n3306), .B(n3305), .Z(n3307) );
  AND U4706 ( .A(n3308), .B(n3307), .Z(n4052) );
  NAND U4707 ( .A(n3310), .B(n3309), .Z(n3314) );
  NAND U4708 ( .A(n3312), .B(n3311), .Z(n3313) );
  NAND U4709 ( .A(n3314), .B(n3313), .Z(n4113) );
  XNOR U4710 ( .A(n4112), .B(n4111), .Z(n3321) );
  XOR U4711 ( .A(n4113), .B(n3321), .Z(n4148) );
  NANDN U4712 ( .A(n3323), .B(n3322), .Z(n3327) );
  NANDN U4713 ( .A(n3325), .B(n3324), .Z(n3326) );
  AND U4714 ( .A(n3327), .B(n3326), .Z(n4146) );
  NANDN U4715 ( .A(n3329), .B(n3328), .Z(n3333) );
  NAND U4716 ( .A(n3331), .B(n3330), .Z(n3332) );
  AND U4717 ( .A(n3333), .B(n3332), .Z(n3896) );
  NAND U4718 ( .A(n3335), .B(n3334), .Z(n3339) );
  NAND U4719 ( .A(n3337), .B(n3336), .Z(n3338) );
  AND U4720 ( .A(n3339), .B(n3338), .Z(n3894) );
  NANDN U4721 ( .A(n3341), .B(n3340), .Z(n3345) );
  NANDN U4722 ( .A(n3343), .B(n3342), .Z(n3344) );
  NAND U4723 ( .A(n3345), .B(n3344), .Z(n3893) );
  XNOR U4724 ( .A(n3894), .B(n3893), .Z(n3895) );
  XNOR U4725 ( .A(n3896), .B(n3895), .Z(n4145) );
  XOR U4726 ( .A(n4146), .B(n4145), .Z(n4147) );
  XOR U4727 ( .A(n4148), .B(n4147), .Z(n4051) );
  XNOR U4728 ( .A(n4052), .B(n4051), .Z(n4053) );
  XNOR U4729 ( .A(n4054), .B(n4053), .Z(n3918) );
  XOR U4730 ( .A(n3919), .B(n3918), .Z(n3921) );
  NAND U4731 ( .A(n3347), .B(n3346), .Z(n3351) );
  NAND U4732 ( .A(n3349), .B(n3348), .Z(n3350) );
  AND U4733 ( .A(n3351), .B(n3350), .Z(n3861) );
  XNOR U4734 ( .A(n3860), .B(n3859), .Z(n3358) );
  XOR U4735 ( .A(n3861), .B(n3358), .Z(n3952) );
  NAND U4736 ( .A(n3360), .B(n3359), .Z(n3364) );
  NAND U4737 ( .A(n3362), .B(n3361), .Z(n3363) );
  AND U4738 ( .A(n3364), .B(n3363), .Z(n3807) );
  NAND U4739 ( .A(n3366), .B(n3365), .Z(n3370) );
  NAND U4740 ( .A(n3368), .B(n3367), .Z(n3369) );
  AND U4741 ( .A(n3370), .B(n3369), .Z(n3805) );
  NAND U4742 ( .A(n3372), .B(n3371), .Z(n3376) );
  NAND U4743 ( .A(n3374), .B(n3373), .Z(n3375) );
  NAND U4744 ( .A(n3376), .B(n3375), .Z(n3804) );
  XNOR U4745 ( .A(n3805), .B(n3804), .Z(n3806) );
  XNOR U4746 ( .A(n3807), .B(n3806), .Z(n3950) );
  NAND U4747 ( .A(n3378), .B(n3377), .Z(n3382) );
  NAND U4748 ( .A(n3380), .B(n3379), .Z(n3381) );
  AND U4749 ( .A(n3382), .B(n3381), .Z(n3838) );
  NAND U4750 ( .A(n3384), .B(n3383), .Z(n3388) );
  NAND U4751 ( .A(n3386), .B(n3385), .Z(n3387) );
  AND U4752 ( .A(n3388), .B(n3387), .Z(n3836) );
  NANDN U4753 ( .A(n3390), .B(n3389), .Z(n3394) );
  NAND U4754 ( .A(n3392), .B(n3391), .Z(n3393) );
  NAND U4755 ( .A(n3394), .B(n3393), .Z(n3835) );
  XNOR U4756 ( .A(n3836), .B(n3835), .Z(n3837) );
  XNOR U4757 ( .A(n3838), .B(n3837), .Z(n3949) );
  XOR U4758 ( .A(n3950), .B(n3949), .Z(n3951) );
  XNOR U4759 ( .A(n3952), .B(n3951), .Z(n3920) );
  XNOR U4760 ( .A(n3921), .B(n3920), .Z(n3986) );
  NANDN U4761 ( .A(n3396), .B(n3395), .Z(n3400) );
  NANDN U4762 ( .A(n3398), .B(n3397), .Z(n3399) );
  AND U4763 ( .A(n3400), .B(n3399), .Z(n3844) );
  NANDN U4764 ( .A(n3402), .B(n3401), .Z(n3406) );
  NAND U4765 ( .A(n3404), .B(n3403), .Z(n3405) );
  AND U4766 ( .A(n3406), .B(n3405), .Z(n3842) );
  NANDN U4767 ( .A(n3408), .B(n3407), .Z(n3412) );
  NANDN U4768 ( .A(n3410), .B(n3409), .Z(n3411) );
  NAND U4769 ( .A(n3412), .B(n3411), .Z(n3841) );
  XNOR U4770 ( .A(n3842), .B(n3841), .Z(n3843) );
  XNOR U4771 ( .A(n3844), .B(n3843), .Z(n4076) );
  NANDN U4772 ( .A(n3414), .B(n3413), .Z(n3418) );
  NAND U4773 ( .A(n3416), .B(n3415), .Z(n3417) );
  AND U4774 ( .A(n3418), .B(n3417), .Z(n3731) );
  NANDN U4775 ( .A(n3420), .B(n3419), .Z(n3424) );
  NAND U4776 ( .A(n3422), .B(n3421), .Z(n3423) );
  AND U4777 ( .A(n3424), .B(n3423), .Z(n3729) );
  NANDN U4778 ( .A(n3426), .B(n3425), .Z(n3430) );
  NAND U4779 ( .A(n3428), .B(n3427), .Z(n3429) );
  NAND U4780 ( .A(n3430), .B(n3429), .Z(n3728) );
  XNOR U4781 ( .A(n3729), .B(n3728), .Z(n3730) );
  XNOR U4782 ( .A(n3731), .B(n3730), .Z(n4075) );
  XOR U4783 ( .A(n4076), .B(n4075), .Z(n4078) );
  NAND U4784 ( .A(n3432), .B(n3431), .Z(n3436) );
  NAND U4785 ( .A(n3434), .B(n3433), .Z(n3435) );
  AND U4786 ( .A(n3436), .B(n3435), .Z(n3725) );
  NANDN U4787 ( .A(n3438), .B(n3437), .Z(n3442) );
  NAND U4788 ( .A(n3440), .B(n3439), .Z(n3441) );
  AND U4789 ( .A(n3442), .B(n3441), .Z(n3723) );
  NANDN U4790 ( .A(n3444), .B(n3443), .Z(n3448) );
  NAND U4791 ( .A(n3446), .B(n3445), .Z(n3447) );
  NAND U4792 ( .A(n3448), .B(n3447), .Z(n3722) );
  XNOR U4793 ( .A(n3723), .B(n3722), .Z(n3724) );
  XNOR U4794 ( .A(n3725), .B(n3724), .Z(n4077) );
  XOR U4795 ( .A(n4078), .B(n4077), .Z(n3915) );
  NAND U4796 ( .A(n3450), .B(n3449), .Z(n3454) );
  NAND U4797 ( .A(n3452), .B(n3451), .Z(n3453) );
  NAND U4798 ( .A(n3454), .B(n3453), .Z(n4102) );
  NAND U4799 ( .A(n3456), .B(n3455), .Z(n3460) );
  NAND U4800 ( .A(n3458), .B(n3457), .Z(n3459) );
  AND U4801 ( .A(n3460), .B(n3459), .Z(n4104) );
  NAND U4802 ( .A(n3462), .B(n3461), .Z(n3466) );
  NAND U4803 ( .A(n3464), .B(n3463), .Z(n3465) );
  AND U4804 ( .A(n3466), .B(n3465), .Z(n4103) );
  XNOR U4805 ( .A(n4104), .B(n4103), .Z(n3467) );
  XNOR U4806 ( .A(n4102), .B(n3467), .Z(n4123) );
  NAND U4807 ( .A(n3469), .B(n3468), .Z(n3473) );
  NAND U4808 ( .A(n3471), .B(n3470), .Z(n3472) );
  AND U4809 ( .A(n3473), .B(n3472), .Z(n4122) );
  NAND U4810 ( .A(n3475), .B(n3474), .Z(n3479) );
  NAND U4811 ( .A(n3477), .B(n3476), .Z(n3478) );
  AND U4812 ( .A(n3479), .B(n3478), .Z(n3801) );
  NAND U4813 ( .A(n3481), .B(n3480), .Z(n3485) );
  NAND U4814 ( .A(n3483), .B(n3482), .Z(n3484) );
  AND U4815 ( .A(n3485), .B(n3484), .Z(n3799) );
  NAND U4816 ( .A(n3487), .B(n3486), .Z(n3491) );
  NAND U4817 ( .A(n3489), .B(n3488), .Z(n3490) );
  NAND U4818 ( .A(n3491), .B(n3490), .Z(n3798) );
  XNOR U4819 ( .A(n3799), .B(n3798), .Z(n3800) );
  XNOR U4820 ( .A(n3801), .B(n3800), .Z(n4121) );
  XOR U4821 ( .A(n4122), .B(n4121), .Z(n4124) );
  XNOR U4822 ( .A(n4123), .B(n4124), .Z(n3912) );
  NANDN U4823 ( .A(n3493), .B(n3492), .Z(n3497) );
  NANDN U4824 ( .A(n3495), .B(n3494), .Z(n3496) );
  AND U4825 ( .A(n3497), .B(n3496), .Z(n3866) );
  NANDN U4826 ( .A(n3499), .B(n3498), .Z(n3503) );
  NAND U4827 ( .A(n3501), .B(n3500), .Z(n3502) );
  NAND U4828 ( .A(n3503), .B(n3502), .Z(n3813) );
  NANDN U4829 ( .A(n3505), .B(n3504), .Z(n3509) );
  NANDN U4830 ( .A(n3507), .B(n3506), .Z(n3508) );
  NAND U4831 ( .A(n3509), .B(n3508), .Z(n3811) );
  NANDN U4832 ( .A(n3511), .B(n3510), .Z(n3515) );
  NANDN U4833 ( .A(n3513), .B(n3512), .Z(n3514) );
  NAND U4834 ( .A(n3515), .B(n3514), .Z(n3810) );
  NAND U4835 ( .A(n3517), .B(n3516), .Z(n3521) );
  NAND U4836 ( .A(n3519), .B(n3518), .Z(n3520) );
  AND U4837 ( .A(n3521), .B(n3520), .Z(n3864) );
  XOR U4838 ( .A(n3863), .B(n3864), .Z(n3865) );
  XNOR U4839 ( .A(n3866), .B(n3865), .Z(n3913) );
  XOR U4840 ( .A(n3912), .B(n3913), .Z(n3914) );
  XNOR U4841 ( .A(n3915), .B(n3914), .Z(n3985) );
  NAND U4842 ( .A(n3523), .B(n3522), .Z(n3527) );
  NAND U4843 ( .A(n3525), .B(n3524), .Z(n3526) );
  NAND U4844 ( .A(n3527), .B(n3526), .Z(n3789) );
  XNOR U4845 ( .A(n3787), .B(n3786), .Z(n3788) );
  NANDN U4846 ( .A(n3535), .B(n3534), .Z(n3539) );
  NAND U4847 ( .A(n3537), .B(n3536), .Z(n3538) );
  AND U4848 ( .A(n3539), .B(n3538), .Z(n4224) );
  XNOR U4849 ( .A(n4222), .B(n4221), .Z(n4223) );
  XNOR U4850 ( .A(n4224), .B(n4223), .Z(n4119) );
  XNOR U4851 ( .A(n4119), .B(n4117), .Z(n3549) );
  XOR U4852 ( .A(n4118), .B(n3549), .Z(n3997) );
  NANDN U4853 ( .A(n3551), .B(n3550), .Z(n3555) );
  NAND U4854 ( .A(n3553), .B(n3552), .Z(n3554) );
  AND U4855 ( .A(n3555), .B(n3554), .Z(n3998) );
  XOR U4856 ( .A(n3997), .B(n3998), .Z(n4000) );
  NAND U4857 ( .A(n3557), .B(n3556), .Z(n3561) );
  NAND U4858 ( .A(n3559), .B(n3558), .Z(n3560) );
  NAND U4859 ( .A(n3561), .B(n3560), .Z(n3762) );
  NANDN U4860 ( .A(n3563), .B(n3562), .Z(n3567) );
  NAND U4861 ( .A(n3565), .B(n3564), .Z(n3566) );
  NAND U4862 ( .A(n3567), .B(n3566), .Z(n3760) );
  NAND U4863 ( .A(n3569), .B(n3568), .Z(n3573) );
  NAND U4864 ( .A(n3571), .B(n3570), .Z(n3572) );
  NAND U4865 ( .A(n3573), .B(n3572), .Z(n3759) );
  NANDN U4866 ( .A(n3575), .B(n3574), .Z(n3579) );
  NANDN U4867 ( .A(n3577), .B(n3576), .Z(n3578) );
  NAND U4868 ( .A(n3579), .B(n3578), .Z(n3931) );
  NANDN U4869 ( .A(n3581), .B(n3580), .Z(n3585) );
  NAND U4870 ( .A(n3583), .B(n3582), .Z(n3584) );
  AND U4871 ( .A(n3585), .B(n3584), .Z(n4236) );
  NANDN U4872 ( .A(n3587), .B(n3586), .Z(n3591) );
  NAND U4873 ( .A(n3589), .B(n3588), .Z(n3590) );
  AND U4874 ( .A(n3591), .B(n3590), .Z(n4234) );
  NANDN U4875 ( .A(n3593), .B(n3592), .Z(n3597) );
  NAND U4876 ( .A(n3595), .B(n3594), .Z(n3596) );
  NAND U4877 ( .A(n3597), .B(n3596), .Z(n4233) );
  XNOR U4878 ( .A(n4234), .B(n4233), .Z(n4235) );
  XOR U4879 ( .A(n4236), .B(n4235), .Z(n3930) );
  XOR U4880 ( .A(n3932), .B(n3933), .Z(n3999) );
  XOR U4881 ( .A(n4000), .B(n3999), .Z(n3927) );
  NANDN U4882 ( .A(n3599), .B(n3598), .Z(n3603) );
  NAND U4883 ( .A(n3601), .B(n3600), .Z(n3602) );
  AND U4884 ( .A(n3603), .B(n3602), .Z(n3964) );
  NANDN U4885 ( .A(n3605), .B(n3604), .Z(n3609) );
  NAND U4886 ( .A(n3607), .B(n3606), .Z(n3608) );
  NAND U4887 ( .A(n3609), .B(n3608), .Z(n3962) );
  NANDN U4888 ( .A(n3611), .B(n3610), .Z(n3615) );
  NANDN U4889 ( .A(n3613), .B(n3612), .Z(n3614) );
  NAND U4890 ( .A(n3615), .B(n3614), .Z(n3961) );
  XOR U4891 ( .A(n3964), .B(n3963), .Z(n3858) );
  NANDN U4892 ( .A(n3617), .B(n3616), .Z(n3621) );
  NANDN U4893 ( .A(n3619), .B(n3618), .Z(n3620) );
  NAND U4894 ( .A(n3621), .B(n3620), .Z(n3857) );
  NAND U4895 ( .A(n3623), .B(n3622), .Z(n3627) );
  NAND U4896 ( .A(n3625), .B(n3624), .Z(n3626) );
  NAND U4897 ( .A(n3627), .B(n3626), .Z(n4162) );
  XOR U4898 ( .A(n4161), .B(n4160), .Z(n4163) );
  XOR U4899 ( .A(n4162), .B(n4163), .Z(n3856) );
  XOR U4900 ( .A(n3857), .B(n3856), .Z(n3634) );
  XOR U4901 ( .A(n3858), .B(n3634), .Z(n4006) );
  NANDN U4902 ( .A(n3639), .B(n3638), .Z(n3643) );
  NANDN U4903 ( .A(n3641), .B(n3640), .Z(n3642) );
  NAND U4904 ( .A(n3643), .B(n3642), .Z(n4141) );
  NAND U4905 ( .A(n3645), .B(n3644), .Z(n3649) );
  NAND U4906 ( .A(n3647), .B(n3646), .Z(n3648) );
  NAND U4907 ( .A(n3649), .B(n3648), .Z(n4139) );
  XNOR U4908 ( .A(oglobal[2]), .B(n4139), .Z(n4140) );
  XOR U4909 ( .A(n3876), .B(n3875), .Z(n3878) );
  NANDN U4910 ( .A(n3651), .B(n3650), .Z(n3655) );
  NAND U4911 ( .A(n3653), .B(n3652), .Z(n3654) );
  NAND U4912 ( .A(n3655), .B(n3654), .Z(n4136) );
  NAND U4913 ( .A(n3657), .B(n3656), .Z(n3661) );
  NAND U4914 ( .A(n3659), .B(n3658), .Z(n3660) );
  NAND U4915 ( .A(n3661), .B(n3660), .Z(n4134) );
  NANDN U4916 ( .A(n3662), .B(oglobal[1]), .Z(n3666) );
  NANDN U4917 ( .A(n3664), .B(n3663), .Z(n3665) );
  AND U4918 ( .A(n3666), .B(n3665), .Z(n4133) );
  XOR U4919 ( .A(n3878), .B(n3877), .Z(n4004) );
  NANDN U4920 ( .A(n3668), .B(n3667), .Z(n3672) );
  NAND U4921 ( .A(n3670), .B(n3669), .Z(n3671) );
  AND U4922 ( .A(n3672), .B(n3671), .Z(n4003) );
  XNOR U4923 ( .A(n4004), .B(n4003), .Z(n4005) );
  XOR U4924 ( .A(n4006), .B(n4005), .Z(n3925) );
  NAND U4925 ( .A(n3674), .B(n3673), .Z(n3678) );
  NAND U4926 ( .A(n3676), .B(n3675), .Z(n3677) );
  AND U4927 ( .A(n3678), .B(n3677), .Z(n4042) );
  NAND U4928 ( .A(n3680), .B(n3679), .Z(n3684) );
  NANDN U4929 ( .A(n3682), .B(n3681), .Z(n3683) );
  AND U4930 ( .A(n3684), .B(n3683), .Z(n4039) );
  NANDN U4931 ( .A(n3686), .B(n3685), .Z(n3690) );
  NANDN U4932 ( .A(n3688), .B(n3687), .Z(n3689) );
  NAND U4933 ( .A(n3690), .B(n3689), .Z(n4040) );
  XNOR U4934 ( .A(n4039), .B(n4040), .Z(n4041) );
  XOR U4935 ( .A(n4042), .B(n4041), .Z(n3924) );
  XOR U4936 ( .A(n3925), .B(n3924), .Z(n3926) );
  XNOR U4937 ( .A(n3927), .B(n3926), .Z(n3987) );
  XOR U4938 ( .A(n3988), .B(n3987), .Z(n4271) );
  XOR U4939 ( .A(n4272), .B(n4271), .Z(n4086) );
  XOR U4940 ( .A(n4087), .B(n4086), .Z(n4082) );
  NAND U4941 ( .A(n3692), .B(n3691), .Z(n3696) );
  NAND U4942 ( .A(n3694), .B(n3693), .Z(n3695) );
  AND U4943 ( .A(n3696), .B(n3695), .Z(n4081) );
  XNOR U4944 ( .A(n4082), .B(n4081), .Z(n3697) );
  XNOR U4945 ( .A(n4083), .B(n3697), .Z(o[2]) );
  NAND U4946 ( .A(n3699), .B(n3698), .Z(n3703) );
  NAND U4947 ( .A(n3701), .B(n3700), .Z(n3702) );
  NAND U4948 ( .A(n3703), .B(n3702), .Z(n4386) );
  NANDN U4949 ( .A(n3705), .B(n3704), .Z(n3709) );
  NAND U4950 ( .A(n3707), .B(n3706), .Z(n3708) );
  AND U4951 ( .A(n3709), .B(n3708), .Z(n4358) );
  NANDN U4952 ( .A(n3711), .B(n3710), .Z(n3715) );
  NAND U4953 ( .A(n3713), .B(n3712), .Z(n3714) );
  AND U4954 ( .A(n3715), .B(n3714), .Z(n4356) );
  NAND U4955 ( .A(n3717), .B(n3716), .Z(n3721) );
  NAND U4956 ( .A(n3719), .B(n3718), .Z(n3720) );
  AND U4957 ( .A(n3721), .B(n3720), .Z(n4355) );
  XNOR U4958 ( .A(n4356), .B(n4355), .Z(n4357) );
  XNOR U4959 ( .A(n4358), .B(n4357), .Z(n4385) );
  NANDN U4960 ( .A(n3723), .B(n3722), .Z(n3727) );
  NANDN U4961 ( .A(n3725), .B(n3724), .Z(n3726) );
  AND U4962 ( .A(n3727), .B(n3726), .Z(n4324) );
  NANDN U4963 ( .A(n3729), .B(n3728), .Z(n3733) );
  NANDN U4964 ( .A(n3731), .B(n3730), .Z(n3732) );
  NAND U4965 ( .A(n3733), .B(n3732), .Z(n4326) );
  NANDN U4966 ( .A(n3735), .B(n3734), .Z(n3739) );
  NAND U4967 ( .A(n3737), .B(n3736), .Z(n3738) );
  NAND U4968 ( .A(n3739), .B(n3738), .Z(n4325) );
  XNOR U4969 ( .A(n4326), .B(n4325), .Z(n3740) );
  XOR U4970 ( .A(n4324), .B(n3740), .Z(n4527) );
  NANDN U4971 ( .A(n3742), .B(n3741), .Z(n3746) );
  NANDN U4972 ( .A(n3744), .B(n3743), .Z(n3745) );
  AND U4973 ( .A(n3746), .B(n3745), .Z(n4526) );
  NANDN U4974 ( .A(n3748), .B(n3747), .Z(n3752) );
  NANDN U4975 ( .A(n3750), .B(n3749), .Z(n3751) );
  NAND U4976 ( .A(n3752), .B(n3751), .Z(n4525) );
  XNOR U4977 ( .A(n4526), .B(n4525), .Z(n4528) );
  XNOR U4978 ( .A(n4527), .B(n4528), .Z(n4509) );
  NANDN U4979 ( .A(n3754), .B(n3753), .Z(n3758) );
  NANDN U4980 ( .A(n3756), .B(n3755), .Z(n3757) );
  NAND U4981 ( .A(n3758), .B(n3757), .Z(n4463) );
  NAND U4982 ( .A(n3760), .B(n3759), .Z(n3764) );
  NAND U4983 ( .A(n3762), .B(n3761), .Z(n3763) );
  NAND U4984 ( .A(n3764), .B(n3763), .Z(n4461) );
  NAND U4985 ( .A(n3766), .B(n3765), .Z(n3770) );
  NANDN U4986 ( .A(n3768), .B(n3767), .Z(n3769) );
  NAND U4987 ( .A(n3770), .B(n3769), .Z(n4460) );
  NANDN U4988 ( .A(n3772), .B(n3771), .Z(n3776) );
  NANDN U4989 ( .A(n3774), .B(n3773), .Z(n3775) );
  NAND U4990 ( .A(n3776), .B(n3775), .Z(n4498) );
  IV U4991 ( .A(n4498), .Z(n4496) );
  NAND U4992 ( .A(n3778), .B(n3777), .Z(n3782) );
  NAND U4993 ( .A(n3780), .B(n3779), .Z(n3781) );
  NAND U4994 ( .A(n3782), .B(n3781), .Z(n4499) );
  NANDN U4995 ( .A(n3787), .B(n3786), .Z(n3791) );
  NAND U4996 ( .A(n3789), .B(n3788), .Z(n3790) );
  AND U4997 ( .A(n3791), .B(n3790), .Z(n4319) );
  XNOR U4998 ( .A(n4320), .B(n4321), .Z(n4507) );
  NANDN U4999 ( .A(n3793), .B(n3792), .Z(n3797) );
  NAND U5000 ( .A(n3795), .B(n3794), .Z(n3796) );
  AND U5001 ( .A(n3797), .B(n3796), .Z(n4294) );
  NANDN U5002 ( .A(n3799), .B(n3798), .Z(n3803) );
  NANDN U5003 ( .A(n3801), .B(n3800), .Z(n3802) );
  AND U5004 ( .A(n3803), .B(n3802), .Z(n4295) );
  NANDN U5005 ( .A(n3805), .B(n3804), .Z(n3809) );
  NANDN U5006 ( .A(n3807), .B(n3806), .Z(n3808) );
  AND U5007 ( .A(n3809), .B(n3808), .Z(n4297) );
  XOR U5008 ( .A(n4507), .B(n4508), .Z(n4510) );
  XOR U5009 ( .A(n4509), .B(n4510), .Z(n4394) );
  NAND U5010 ( .A(n3811), .B(n3810), .Z(n3815) );
  NAND U5011 ( .A(n3813), .B(n3812), .Z(n3814) );
  AND U5012 ( .A(n3815), .B(n3814), .Z(n4503) );
  NAND U5013 ( .A(n3817), .B(n3816), .Z(n3821) );
  NAND U5014 ( .A(n3819), .B(n3818), .Z(n3820) );
  NAND U5015 ( .A(n3821), .B(n3820), .Z(n4505) );
  NANDN U5016 ( .A(n3823), .B(n3822), .Z(n3827) );
  NAND U5017 ( .A(n3825), .B(n3824), .Z(n3826) );
  NAND U5018 ( .A(n3827), .B(n3826), .Z(n4504) );
  XNOR U5019 ( .A(n4505), .B(n4504), .Z(n3828) );
  XOR U5020 ( .A(n4503), .B(n3828), .Z(n4278) );
  NANDN U5021 ( .A(n3830), .B(n3829), .Z(n3834) );
  NAND U5022 ( .A(n3832), .B(n3831), .Z(n3833) );
  AND U5023 ( .A(n3834), .B(n3833), .Z(n4277) );
  NANDN U5024 ( .A(n3836), .B(n3835), .Z(n3840) );
  NANDN U5025 ( .A(n3838), .B(n3837), .Z(n3839) );
  AND U5026 ( .A(n3840), .B(n3839), .Z(n4542) );
  NANDN U5027 ( .A(n3842), .B(n3841), .Z(n3846) );
  NANDN U5028 ( .A(n3844), .B(n3843), .Z(n3845) );
  NAND U5029 ( .A(n3846), .B(n3845), .Z(n4543) );
  XNOR U5030 ( .A(n4542), .B(n4543), .Z(n4545) );
  NANDN U5031 ( .A(n3848), .B(n3847), .Z(n3852) );
  NANDN U5032 ( .A(n3850), .B(n3849), .Z(n3851) );
  AND U5033 ( .A(n3852), .B(n3851), .Z(n4544) );
  XNOR U5034 ( .A(n4545), .B(n4544), .Z(n4276) );
  XNOR U5035 ( .A(n4277), .B(n4276), .Z(n4279) );
  XNOR U5036 ( .A(n4278), .B(n4279), .Z(n4391) );
  XOR U5037 ( .A(n4458), .B(n4457), .Z(n3862) );
  XOR U5038 ( .A(n4456), .B(n3862), .Z(n4522) );
  NAND U5039 ( .A(n3864), .B(n3863), .Z(n3868) );
  NANDN U5040 ( .A(n3866), .B(n3865), .Z(n3867) );
  AND U5041 ( .A(n3868), .B(n3867), .Z(n4520) );
  NAND U5042 ( .A(n3870), .B(n3869), .Z(n3874) );
  NANDN U5043 ( .A(n3872), .B(n3871), .Z(n3873) );
  AND U5044 ( .A(n3874), .B(n3873), .Z(n4447) );
  IV U5045 ( .A(n4447), .Z(n4445) );
  NAND U5046 ( .A(n3876), .B(n3875), .Z(n3880) );
  NAND U5047 ( .A(n3878), .B(n3877), .Z(n3879) );
  AND U5048 ( .A(n3880), .B(n3879), .Z(n4450) );
  NAND U5049 ( .A(n3882), .B(n3881), .Z(n3886) );
  NAND U5050 ( .A(n3884), .B(n3883), .Z(n3885) );
  AND U5051 ( .A(n3886), .B(n3885), .Z(n4490) );
  NANDN U5052 ( .A(n3888), .B(n3887), .Z(n3892) );
  NANDN U5053 ( .A(n3890), .B(n3889), .Z(n3891) );
  AND U5054 ( .A(n3892), .B(n3891), .Z(n4487) );
  NANDN U5055 ( .A(n3894), .B(n3893), .Z(n3898) );
  NANDN U5056 ( .A(n3896), .B(n3895), .Z(n3897) );
  AND U5057 ( .A(n3898), .B(n3897), .Z(n4488) );
  XNOR U5058 ( .A(n4490), .B(n4489), .Z(n4446) );
  IV U5059 ( .A(n4446), .Z(n4448) );
  XNOR U5060 ( .A(n4450), .B(n4448), .Z(n3899) );
  XNOR U5061 ( .A(n4445), .B(n3899), .Z(n4519) );
  XNOR U5062 ( .A(n4520), .B(n4519), .Z(n4521) );
  XNOR U5063 ( .A(n4522), .B(n4521), .Z(n4392) );
  XOR U5064 ( .A(n4391), .B(n4392), .Z(n4393) );
  XNOR U5065 ( .A(n4394), .B(n4393), .Z(n4362) );
  NAND U5066 ( .A(n3901), .B(n3900), .Z(n3905) );
  NAND U5067 ( .A(n3903), .B(n3902), .Z(n3904) );
  AND U5068 ( .A(n3905), .B(n3904), .Z(n4400) );
  NAND U5069 ( .A(n3907), .B(n3906), .Z(n3911) );
  NAND U5070 ( .A(n3909), .B(n3908), .Z(n3910) );
  AND U5071 ( .A(n3911), .B(n3910), .Z(n4398) );
  NAND U5072 ( .A(n3913), .B(n3912), .Z(n3917) );
  NANDN U5073 ( .A(n3915), .B(n3914), .Z(n3916) );
  AND U5074 ( .A(n3917), .B(n3916), .Z(n4397) );
  XNOR U5075 ( .A(n4398), .B(n4397), .Z(n4399) );
  XNOR U5076 ( .A(n4400), .B(n4399), .Z(n4361) );
  NAND U5077 ( .A(n3919), .B(n3918), .Z(n3923) );
  NAND U5078 ( .A(n3921), .B(n3920), .Z(n3922) );
  AND U5079 ( .A(n3923), .B(n3922), .Z(n4352) );
  NAND U5080 ( .A(n3925), .B(n3924), .Z(n3929) );
  NANDN U5081 ( .A(n3927), .B(n3926), .Z(n3928) );
  AND U5082 ( .A(n3929), .B(n3928), .Z(n4350) );
  NAND U5083 ( .A(n3931), .B(n3930), .Z(n3935) );
  NAND U5084 ( .A(n3933), .B(n3932), .Z(n3934) );
  AND U5085 ( .A(n3935), .B(n3934), .Z(n4327) );
  NAND U5086 ( .A(n3937), .B(n3936), .Z(n3941) );
  NAND U5087 ( .A(n3939), .B(n3938), .Z(n3940) );
  NAND U5088 ( .A(n3941), .B(n3940), .Z(n4329) );
  NANDN U5089 ( .A(n3943), .B(n3942), .Z(n3947) );
  NANDN U5090 ( .A(n3945), .B(n3944), .Z(n3946) );
  NAND U5091 ( .A(n3947), .B(n3946), .Z(n4328) );
  XNOR U5092 ( .A(n4329), .B(n4328), .Z(n3948) );
  XOR U5093 ( .A(n4327), .B(n3948), .Z(n4314) );
  NAND U5094 ( .A(n3950), .B(n3949), .Z(n3954) );
  NANDN U5095 ( .A(n3952), .B(n3951), .Z(n3953) );
  AND U5096 ( .A(n3954), .B(n3953), .Z(n4313) );
  NANDN U5097 ( .A(n3956), .B(n3955), .Z(n3960) );
  NAND U5098 ( .A(n3958), .B(n3957), .Z(n3959) );
  AND U5099 ( .A(n3960), .B(n3959), .Z(n4291) );
  NAND U5100 ( .A(n3962), .B(n3961), .Z(n3966) );
  NANDN U5101 ( .A(n3964), .B(n3963), .Z(n3965) );
  AND U5102 ( .A(n3966), .B(n3965), .Z(n4478) );
  NAND U5103 ( .A(n3968), .B(n3967), .Z(n3972) );
  NAND U5104 ( .A(n3970), .B(n3969), .Z(n3971) );
  AND U5105 ( .A(n3972), .B(n3971), .Z(n4475) );
  NAND U5106 ( .A(n3974), .B(n3973), .Z(n3978) );
  NAND U5107 ( .A(n3976), .B(n3975), .Z(n3977) );
  NAND U5108 ( .A(n3978), .B(n3977), .Z(n4476) );
  XNOR U5109 ( .A(n4475), .B(n4476), .Z(n4477) );
  XOR U5110 ( .A(n4478), .B(n4477), .Z(n4289) );
  NANDN U5111 ( .A(n3980), .B(n3979), .Z(n3984) );
  NANDN U5112 ( .A(n3982), .B(n3981), .Z(n3983) );
  AND U5113 ( .A(n3984), .B(n3983), .Z(n4288) );
  XNOR U5114 ( .A(n4289), .B(n4288), .Z(n4290) );
  XOR U5115 ( .A(n4291), .B(n4290), .Z(n4312) );
  XNOR U5116 ( .A(n4313), .B(n4312), .Z(n4315) );
  XOR U5117 ( .A(n4314), .B(n4315), .Z(n4349) );
  XOR U5118 ( .A(n4350), .B(n4349), .Z(n4351) );
  XOR U5119 ( .A(n4352), .B(n4351), .Z(n4364) );
  XOR U5120 ( .A(n4363), .B(n4364), .Z(n4382) );
  NAND U5121 ( .A(n3986), .B(n3985), .Z(n3990) );
  NAND U5122 ( .A(n3988), .B(n3987), .Z(n3989) );
  NAND U5123 ( .A(n3990), .B(n3989), .Z(n4380) );
  NAND U5124 ( .A(n3992), .B(n3991), .Z(n3996) );
  NAND U5125 ( .A(n3994), .B(n3993), .Z(n3995) );
  AND U5126 ( .A(n3996), .B(n3995), .Z(n4428) );
  NAND U5127 ( .A(n3998), .B(n3997), .Z(n4002) );
  NAND U5128 ( .A(n4000), .B(n3999), .Z(n4001) );
  AND U5129 ( .A(n4002), .B(n4001), .Z(n4412) );
  NANDN U5130 ( .A(n4004), .B(n4003), .Z(n4008) );
  NANDN U5131 ( .A(n4006), .B(n4005), .Z(n4007) );
  AND U5132 ( .A(n4008), .B(n4007), .Z(n4410) );
  NAND U5133 ( .A(n4010), .B(n4009), .Z(n4014) );
  NAND U5134 ( .A(n4012), .B(n4011), .Z(n4013) );
  NAND U5135 ( .A(n4014), .B(n4013), .Z(n4409) );
  XNOR U5136 ( .A(n4410), .B(n4409), .Z(n4411) );
  XNOR U5137 ( .A(n4412), .B(n4411), .Z(n4427) );
  XNOR U5138 ( .A(n4428), .B(n4427), .Z(n4429) );
  NAND U5139 ( .A(n4016), .B(n4015), .Z(n4020) );
  NAND U5140 ( .A(n4018), .B(n4017), .Z(n4019) );
  NAND U5141 ( .A(n4020), .B(n4019), .Z(n4430) );
  XNOR U5142 ( .A(n4429), .B(n4430), .Z(n4374) );
  NAND U5143 ( .A(n4022), .B(n4021), .Z(n4026) );
  NANDN U5144 ( .A(n4024), .B(n4023), .Z(n4025) );
  AND U5145 ( .A(n4026), .B(n4025), .Z(n4373) );
  XOR U5146 ( .A(n4374), .B(n4373), .Z(n4376) );
  NAND U5147 ( .A(n4028), .B(n4027), .Z(n4032) );
  NAND U5148 ( .A(n4030), .B(n4029), .Z(n4031) );
  AND U5149 ( .A(n4032), .B(n4031), .Z(n4331) );
  NANDN U5150 ( .A(n4034), .B(n4033), .Z(n4038) );
  NAND U5151 ( .A(n4036), .B(n4035), .Z(n4037) );
  AND U5152 ( .A(n4038), .B(n4037), .Z(n4332) );
  NANDN U5153 ( .A(n4040), .B(n4039), .Z(n4044) );
  NANDN U5154 ( .A(n4042), .B(n4041), .Z(n4043) );
  AND U5155 ( .A(n4044), .B(n4043), .Z(n4333) );
  XOR U5156 ( .A(n4334), .B(n4333), .Z(n4404) );
  NANDN U5157 ( .A(n4046), .B(n4045), .Z(n4050) );
  NAND U5158 ( .A(n4048), .B(n4047), .Z(n4049) );
  AND U5159 ( .A(n4050), .B(n4049), .Z(n4309) );
  NANDN U5160 ( .A(n4052), .B(n4051), .Z(n4056) );
  NANDN U5161 ( .A(n4054), .B(n4053), .Z(n4055) );
  AND U5162 ( .A(n4056), .B(n4055), .Z(n4307) );
  NANDN U5163 ( .A(n4058), .B(n4057), .Z(n4062) );
  NAND U5164 ( .A(n4060), .B(n4059), .Z(n4061) );
  NAND U5165 ( .A(n4062), .B(n4061), .Z(n4306) );
  XNOR U5166 ( .A(n4307), .B(n4306), .Z(n4308) );
  XNOR U5167 ( .A(n4309), .B(n4308), .Z(n4403) );
  XNOR U5168 ( .A(n4404), .B(n4403), .Z(n4406) );
  NANDN U5169 ( .A(n4064), .B(n4063), .Z(n4068) );
  NANDN U5170 ( .A(n4066), .B(n4065), .Z(n4067) );
  AND U5171 ( .A(n4068), .B(n4067), .Z(n4424) );
  NANDN U5172 ( .A(n4070), .B(n4069), .Z(n4074) );
  NAND U5173 ( .A(n4072), .B(n4071), .Z(n4073) );
  AND U5174 ( .A(n4074), .B(n4073), .Z(n4422) );
  NAND U5175 ( .A(n4076), .B(n4075), .Z(n4080) );
  NAND U5176 ( .A(n4078), .B(n4077), .Z(n4079) );
  NAND U5177 ( .A(n4080), .B(n4079), .Z(n4421) );
  XNOR U5178 ( .A(n4422), .B(n4421), .Z(n4423) );
  XNOR U5179 ( .A(n4424), .B(n4423), .Z(n4405) );
  XOR U5180 ( .A(n4406), .B(n4405), .Z(n4375) );
  XNOR U5181 ( .A(n4376), .B(n4375), .Z(n4379) );
  XOR U5182 ( .A(n4380), .B(n4379), .Z(n4381) );
  XNOR U5183 ( .A(n4388), .B(n4387), .Z(n4556) );
  NANDN U5184 ( .A(n4085), .B(n4084), .Z(n4089) );
  NAND U5185 ( .A(n4087), .B(n4086), .Z(n4088) );
  AND U5186 ( .A(n4089), .B(n4088), .Z(n4551) );
  NAND U5187 ( .A(n4091), .B(n4090), .Z(n4095) );
  NANDN U5188 ( .A(n4093), .B(n4092), .Z(n4094) );
  NAND U5189 ( .A(n4095), .B(n4094), .Z(n4367) );
  NANDN U5190 ( .A(n4097), .B(n4096), .Z(n4101) );
  NANDN U5191 ( .A(n4099), .B(n4098), .Z(n4100) );
  AND U5192 ( .A(n4101), .B(n4100), .Z(n4346) );
  NAND U5193 ( .A(n4106), .B(n4105), .Z(n4110) );
  NANDN U5194 ( .A(n4108), .B(n4107), .Z(n4109) );
  AND U5195 ( .A(n4110), .B(n4109), .Z(n4483) );
  XOR U5196 ( .A(n4482), .B(n4481), .Z(n4484) );
  XNOR U5197 ( .A(n4483), .B(n4484), .Z(n4454) );
  XNOR U5198 ( .A(n4454), .B(n4453), .Z(n4120) );
  XOR U5199 ( .A(n4455), .B(n4120), .Z(n4285) );
  NAND U5200 ( .A(n4122), .B(n4121), .Z(n4126) );
  NAND U5201 ( .A(n4124), .B(n4123), .Z(n4125) );
  AND U5202 ( .A(n4126), .B(n4125), .Z(n4283) );
  NANDN U5203 ( .A(n4128), .B(n4127), .Z(n4132) );
  NANDN U5204 ( .A(n4130), .B(n4129), .Z(n4131) );
  NAND U5205 ( .A(n4132), .B(n4131), .Z(n4472) );
  NAND U5206 ( .A(n4134), .B(n4133), .Z(n4138) );
  NAND U5207 ( .A(n4136), .B(n4135), .Z(n4137) );
  AND U5208 ( .A(n4138), .B(n4137), .Z(n4474) );
  NANDN U5209 ( .A(oglobal[2]), .B(n4139), .Z(n4143) );
  NAND U5210 ( .A(n4141), .B(n4140), .Z(n4142) );
  AND U5211 ( .A(n4143), .B(n4142), .Z(n4473) );
  XNOR U5212 ( .A(n4474), .B(n4473), .Z(n4144) );
  XNOR U5213 ( .A(n4472), .B(n4144), .Z(n4441) );
  NAND U5214 ( .A(n4146), .B(n4145), .Z(n4150) );
  NANDN U5215 ( .A(n4148), .B(n4147), .Z(n4149) );
  AND U5216 ( .A(n4150), .B(n4149), .Z(n4440) );
  NAND U5217 ( .A(n4155), .B(n4154), .Z(n4159) );
  NANDN U5218 ( .A(n4157), .B(n4156), .Z(n4158) );
  AND U5219 ( .A(n4159), .B(n4158), .Z(n4495) );
  NAND U5220 ( .A(n4161), .B(n4160), .Z(n4165) );
  NAND U5221 ( .A(n4163), .B(n4162), .Z(n4164) );
  AND U5222 ( .A(n4165), .B(n4164), .Z(n4494) );
  XNOR U5223 ( .A(n4495), .B(n4494), .Z(n4166) );
  XNOR U5224 ( .A(n4493), .B(n4166), .Z(n4439) );
  XNOR U5225 ( .A(n4440), .B(n4439), .Z(n4442) );
  XNOR U5226 ( .A(n4441), .B(n4442), .Z(n4282) );
  XNOR U5227 ( .A(n4283), .B(n4282), .Z(n4284) );
  XOR U5228 ( .A(n4285), .B(n4284), .Z(n4343) );
  NAND U5229 ( .A(n4168), .B(n4167), .Z(n4172) );
  NANDN U5230 ( .A(n4170), .B(n4169), .Z(n4171) );
  AND U5231 ( .A(n4172), .B(n4171), .Z(n4344) );
  XOR U5232 ( .A(n4343), .B(n4344), .Z(n4345) );
  XNOR U5233 ( .A(n4346), .B(n4345), .Z(n4368) );
  XOR U5234 ( .A(n4367), .B(n4368), .Z(n4370) );
  NANDN U5235 ( .A(n4174), .B(n4173), .Z(n4178) );
  NAND U5236 ( .A(n4176), .B(n4175), .Z(n4177) );
  AND U5237 ( .A(n4178), .B(n4177), .Z(n4418) );
  NANDN U5238 ( .A(n4180), .B(n4179), .Z(n4184) );
  NANDN U5239 ( .A(n4182), .B(n4181), .Z(n4183) );
  AND U5240 ( .A(n4184), .B(n4183), .Z(n4416) );
  NAND U5241 ( .A(n4186), .B(n4185), .Z(n4190) );
  NAND U5242 ( .A(n4188), .B(n4187), .Z(n4189) );
  NAND U5243 ( .A(n4190), .B(n4189), .Z(n4415) );
  XNOR U5244 ( .A(n4416), .B(n4415), .Z(n4417) );
  XOR U5245 ( .A(n4418), .B(n4417), .Z(n4337) );
  NANDN U5246 ( .A(n4192), .B(n4191), .Z(n4196) );
  NANDN U5247 ( .A(n4194), .B(n4193), .Z(n4195) );
  AND U5248 ( .A(n4196), .B(n4195), .Z(n4338) );
  XOR U5249 ( .A(n4337), .B(n4338), .Z(n4340) );
  NANDN U5250 ( .A(n4198), .B(n4197), .Z(n4202) );
  NAND U5251 ( .A(n4200), .B(n4199), .Z(n4201) );
  NAND U5252 ( .A(n4202), .B(n4201), .Z(n4303) );
  NANDN U5253 ( .A(n4204), .B(n4203), .Z(n4208) );
  NAND U5254 ( .A(n4206), .B(n4205), .Z(n4207) );
  NAND U5255 ( .A(n4208), .B(n4207), .Z(n4301) );
  NAND U5256 ( .A(n4210), .B(n4209), .Z(n4214) );
  NAND U5257 ( .A(n4212), .B(n4211), .Z(n4213) );
  AND U5258 ( .A(n4214), .B(n4213), .Z(n4469) );
  NANDN U5259 ( .A(n4216), .B(n4215), .Z(n4220) );
  NAND U5260 ( .A(n4218), .B(n4217), .Z(n4219) );
  AND U5261 ( .A(n4220), .B(n4219), .Z(n4466) );
  NANDN U5262 ( .A(n4222), .B(n4221), .Z(n4226) );
  NANDN U5263 ( .A(n4224), .B(n4223), .Z(n4225) );
  AND U5264 ( .A(n4226), .B(n4225), .Z(n4467) );
  XOR U5265 ( .A(n4469), .B(n4468), .Z(n4300) );
  NANDN U5266 ( .A(n4228), .B(n4227), .Z(n4232) );
  NAND U5267 ( .A(n4230), .B(n4229), .Z(n4231) );
  AND U5268 ( .A(n4232), .B(n4231), .Z(n4514) );
  XOR U5269 ( .A(n4513), .B(n4514), .Z(n4516) );
  NANDN U5270 ( .A(n4234), .B(n4233), .Z(n4238) );
  NANDN U5271 ( .A(n4236), .B(n4235), .Z(n4237) );
  AND U5272 ( .A(n4238), .B(n4237), .Z(n4533) );
  NANDN U5273 ( .A(n4240), .B(n4239), .Z(n4244) );
  NANDN U5274 ( .A(n4242), .B(n4241), .Z(n4243) );
  NAND U5275 ( .A(n4244), .B(n4243), .Z(n4531) );
  XNOR U5276 ( .A(oglobal[3]), .B(n4531), .Z(n4532) );
  XNOR U5277 ( .A(n4533), .B(n4532), .Z(n4436) );
  NANDN U5278 ( .A(n4246), .B(n4245), .Z(n4250) );
  NANDN U5279 ( .A(n4248), .B(n4247), .Z(n4249) );
  AND U5280 ( .A(n4250), .B(n4249), .Z(n4539) );
  NAND U5281 ( .A(n4252), .B(n4251), .Z(n4256) );
  NAND U5282 ( .A(n4254), .B(n4253), .Z(n4255) );
  AND U5283 ( .A(n4256), .B(n4255), .Z(n4536) );
  NANDN U5284 ( .A(n4258), .B(n4257), .Z(n4262) );
  NANDN U5285 ( .A(n4260), .B(n4259), .Z(n4261) );
  NAND U5286 ( .A(n4262), .B(n4261), .Z(n4537) );
  XNOR U5287 ( .A(n4536), .B(n4537), .Z(n4538) );
  XNOR U5288 ( .A(n4539), .B(n4538), .Z(n4434) );
  NANDN U5289 ( .A(n4264), .B(n4263), .Z(n4268) );
  NAND U5290 ( .A(n4266), .B(n4265), .Z(n4267) );
  AND U5291 ( .A(n4268), .B(n4267), .Z(n4433) );
  XOR U5292 ( .A(n4516), .B(n4515), .Z(n4339) );
  XOR U5293 ( .A(n4340), .B(n4339), .Z(n4369) );
  XNOR U5294 ( .A(n4370), .B(n4369), .Z(n4549) );
  NAND U5295 ( .A(n4270), .B(n4269), .Z(n4274) );
  NAND U5296 ( .A(n4272), .B(n4271), .Z(n4273) );
  AND U5297 ( .A(n4274), .B(n4273), .Z(n4548) );
  XNOR U5298 ( .A(n4551), .B(n4550), .Z(n4554) );
  XNOR U5299 ( .A(n4555), .B(n4554), .Z(n4275) );
  XNOR U5300 ( .A(n4556), .B(n4275), .Z(o[3]) );
  NANDN U5301 ( .A(n4277), .B(n4276), .Z(n4281) );
  NAND U5302 ( .A(n4279), .B(n4278), .Z(n4280) );
  AND U5303 ( .A(n4281), .B(n4280), .Z(n4662) );
  NANDN U5304 ( .A(n4283), .B(n4282), .Z(n4287) );
  NANDN U5305 ( .A(n4285), .B(n4284), .Z(n4286) );
  AND U5306 ( .A(n4287), .B(n4286), .Z(n4660) );
  NANDN U5307 ( .A(n4289), .B(n4288), .Z(n4293) );
  NANDN U5308 ( .A(n4291), .B(n4290), .Z(n4292) );
  AND U5309 ( .A(n4293), .B(n4292), .Z(n4597) );
  NAND U5310 ( .A(n4295), .B(n4294), .Z(n4299) );
  NAND U5311 ( .A(n4297), .B(n4296), .Z(n4298) );
  AND U5312 ( .A(n4299), .B(n4298), .Z(n4595) );
  NAND U5313 ( .A(n4301), .B(n4300), .Z(n4305) );
  NAND U5314 ( .A(n4303), .B(n4302), .Z(n4304) );
  AND U5315 ( .A(n4305), .B(n4304), .Z(n4594) );
  XNOR U5316 ( .A(n4595), .B(n4594), .Z(n4596) );
  XOR U5317 ( .A(n4597), .B(n4596), .Z(n4659) );
  XNOR U5318 ( .A(n4660), .B(n4659), .Z(n4661) );
  XOR U5319 ( .A(n4662), .B(n4661), .Z(n4694) );
  NANDN U5320 ( .A(n4307), .B(n4306), .Z(n4311) );
  NANDN U5321 ( .A(n4309), .B(n4308), .Z(n4310) );
  AND U5322 ( .A(n4311), .B(n4310), .Z(n4626) );
  NANDN U5323 ( .A(n4313), .B(n4312), .Z(n4317) );
  NAND U5324 ( .A(n4315), .B(n4314), .Z(n4316) );
  AND U5325 ( .A(n4317), .B(n4316), .Z(n4624) );
  NAND U5326 ( .A(n4319), .B(n4318), .Z(n4323) );
  NAND U5327 ( .A(n4321), .B(n4320), .Z(n4322) );
  NAND U5328 ( .A(n4323), .B(n4322), .Z(n4646) );
  XNOR U5329 ( .A(n4645), .B(n4644), .Z(n4330) );
  XNOR U5330 ( .A(n4646), .B(n4330), .Z(n4623) );
  XNOR U5331 ( .A(n4624), .B(n4623), .Z(n4625) );
  XOR U5332 ( .A(n4626), .B(n4625), .Z(n4693) );
  NAND U5333 ( .A(n4332), .B(n4331), .Z(n4336) );
  NAND U5334 ( .A(n4334), .B(n4333), .Z(n4335) );
  NAND U5335 ( .A(n4336), .B(n4335), .Z(n4692) );
  XOR U5336 ( .A(n4693), .B(n4692), .Z(n4695) );
  XNOR U5337 ( .A(n4694), .B(n4695), .Z(n4675) );
  NAND U5338 ( .A(n4338), .B(n4337), .Z(n4342) );
  NAND U5339 ( .A(n4340), .B(n4339), .Z(n4341) );
  AND U5340 ( .A(n4342), .B(n4341), .Z(n4701) );
  NAND U5341 ( .A(n4344), .B(n4343), .Z(n4348) );
  NANDN U5342 ( .A(n4346), .B(n4345), .Z(n4347) );
  AND U5343 ( .A(n4348), .B(n4347), .Z(n4699) );
  NAND U5344 ( .A(n4350), .B(n4349), .Z(n4354) );
  NANDN U5345 ( .A(n4352), .B(n4351), .Z(n4353) );
  AND U5346 ( .A(n4354), .B(n4353), .Z(n4698) );
  XNOR U5347 ( .A(n4699), .B(n4698), .Z(n4700) );
  XOR U5348 ( .A(n4701), .B(n4700), .Z(n4674) );
  XOR U5349 ( .A(n4675), .B(n4674), .Z(n4676) );
  NANDN U5350 ( .A(n4356), .B(n4355), .Z(n4360) );
  NANDN U5351 ( .A(n4358), .B(n4357), .Z(n4359) );
  NAND U5352 ( .A(n4360), .B(n4359), .Z(n4677) );
  XNOR U5353 ( .A(n4676), .B(n4677), .Z(n4558) );
  NAND U5354 ( .A(n4362), .B(n4361), .Z(n4366) );
  NANDN U5355 ( .A(n4364), .B(n4363), .Z(n4365) );
  AND U5356 ( .A(n4366), .B(n4365), .Z(n4566) );
  NAND U5357 ( .A(n4368), .B(n4367), .Z(n4372) );
  NAND U5358 ( .A(n4370), .B(n4369), .Z(n4371) );
  NAND U5359 ( .A(n4372), .B(n4371), .Z(n4564) );
  NAND U5360 ( .A(n4374), .B(n4373), .Z(n4378) );
  NAND U5361 ( .A(n4376), .B(n4375), .Z(n4377) );
  AND U5362 ( .A(n4378), .B(n4377), .Z(n4565) );
  XOR U5363 ( .A(n4564), .B(n4565), .Z(n4567) );
  NAND U5364 ( .A(n4380), .B(n4379), .Z(n4384) );
  NAND U5365 ( .A(n4382), .B(n4381), .Z(n4383) );
  AND U5366 ( .A(n4384), .B(n4383), .Z(n4560) );
  XOR U5367 ( .A(n4561), .B(n4560), .Z(n4673) );
  NAND U5368 ( .A(n4386), .B(n4385), .Z(n4390) );
  NAND U5369 ( .A(n4388), .B(n4387), .Z(n4389) );
  AND U5370 ( .A(n4390), .B(n4389), .Z(n4667) );
  NAND U5371 ( .A(n4392), .B(n4391), .Z(n4396) );
  NAND U5372 ( .A(n4394), .B(n4393), .Z(n4395) );
  AND U5373 ( .A(n4396), .B(n4395), .Z(n4681) );
  NANDN U5374 ( .A(n4398), .B(n4397), .Z(n4402) );
  NANDN U5375 ( .A(n4400), .B(n4399), .Z(n4401) );
  AND U5376 ( .A(n4402), .B(n4401), .Z(n4689) );
  NANDN U5377 ( .A(n4404), .B(n4403), .Z(n4408) );
  NAND U5378 ( .A(n4406), .B(n4405), .Z(n4407) );
  AND U5379 ( .A(n4408), .B(n4407), .Z(n4687) );
  NANDN U5380 ( .A(n4410), .B(n4409), .Z(n4414) );
  NANDN U5381 ( .A(n4412), .B(n4411), .Z(n4413) );
  AND U5382 ( .A(n4414), .B(n4413), .Z(n4588) );
  NANDN U5383 ( .A(n4416), .B(n4415), .Z(n4420) );
  NANDN U5384 ( .A(n4418), .B(n4417), .Z(n4419) );
  NAND U5385 ( .A(n4420), .B(n4419), .Z(n4589) );
  XNOR U5386 ( .A(n4588), .B(n4589), .Z(n4591) );
  NANDN U5387 ( .A(n4422), .B(n4421), .Z(n4426) );
  NANDN U5388 ( .A(n4424), .B(n4423), .Z(n4425) );
  AND U5389 ( .A(n4426), .B(n4425), .Z(n4590) );
  XNOR U5390 ( .A(n4591), .B(n4590), .Z(n4686) );
  XNOR U5391 ( .A(n4687), .B(n4686), .Z(n4688) );
  XOR U5392 ( .A(n4689), .B(n4688), .Z(n4680) );
  XNOR U5393 ( .A(n4681), .B(n4680), .Z(n4683) );
  NANDN U5394 ( .A(n4428), .B(n4427), .Z(n4432) );
  NANDN U5395 ( .A(n4430), .B(n4429), .Z(n4431) );
  AND U5396 ( .A(n4432), .B(n4431), .Z(n4570) );
  NAND U5397 ( .A(n4434), .B(n4433), .Z(n4438) );
  NAND U5398 ( .A(n4436), .B(n4435), .Z(n4437) );
  AND U5399 ( .A(n4438), .B(n4437), .Z(n4631) );
  IV U5400 ( .A(n4631), .Z(n4629) );
  NANDN U5401 ( .A(n4440), .B(n4439), .Z(n4444) );
  NAND U5402 ( .A(n4442), .B(n4441), .Z(n4443) );
  AND U5403 ( .A(n4444), .B(n4443), .Z(n4634) );
  NAND U5404 ( .A(n4446), .B(n4445), .Z(n4452) );
  AND U5405 ( .A(n4448), .B(n4447), .Z(n4449) );
  OR U5406 ( .A(n4450), .B(n4449), .Z(n4451) );
  AND U5407 ( .A(n4452), .B(n4451), .Z(n4656) );
  XNOR U5408 ( .A(n4653), .B(n4654), .Z(n4655) );
  XNOR U5409 ( .A(n4656), .B(n4655), .Z(n4630) );
  IV U5410 ( .A(n4630), .Z(n4632) );
  XNOR U5411 ( .A(n4634), .B(n4632), .Z(n4459) );
  XNOR U5412 ( .A(n4629), .B(n4459), .Z(n4578) );
  NAND U5413 ( .A(n4461), .B(n4460), .Z(n4465) );
  NAND U5414 ( .A(n4463), .B(n4462), .Z(n4464) );
  AND U5415 ( .A(n4465), .B(n4464), .Z(n4609) );
  NAND U5416 ( .A(n4467), .B(n4466), .Z(n4471) );
  NAND U5417 ( .A(n4469), .B(n4468), .Z(n4470) );
  NAND U5418 ( .A(n4471), .B(n4470), .Z(n4607) );
  XNOR U5419 ( .A(n4609), .B(n4608), .Z(n4639) );
  IV U5420 ( .A(n4639), .Z(n4637) );
  NANDN U5421 ( .A(n4476), .B(n4475), .Z(n4480) );
  NAND U5422 ( .A(n4478), .B(n4477), .Z(n4479) );
  AND U5423 ( .A(n4480), .B(n4479), .Z(n4600) );
  NANDN U5424 ( .A(n4482), .B(n4481), .Z(n4486) );
  NANDN U5425 ( .A(n4484), .B(n4483), .Z(n4485) );
  AND U5426 ( .A(n4486), .B(n4485), .Z(n4601) );
  NAND U5427 ( .A(n4488), .B(n4487), .Z(n4492) );
  NAND U5428 ( .A(n4490), .B(n4489), .Z(n4491) );
  AND U5429 ( .A(n4492), .B(n4491), .Z(n4615) );
  NAND U5430 ( .A(n4496), .B(n4497), .Z(n4502) );
  ANDN U5431 ( .B(n4498), .A(n4497), .Z(n4500) );
  OR U5432 ( .A(n4500), .B(n4499), .Z(n4501) );
  AND U5433 ( .A(n4502), .B(n4501), .Z(n4612) );
  XNOR U5434 ( .A(n4613), .B(n4612), .Z(n4614) );
  XOR U5435 ( .A(n4615), .B(n4614), .Z(n4602) );
  XOR U5436 ( .A(n4603), .B(n4602), .Z(n4641) );
  XNOR U5437 ( .A(n4641), .B(n4638), .Z(n4506) );
  XNOR U5438 ( .A(n4637), .B(n4506), .Z(n4576) );
  NAND U5439 ( .A(n4508), .B(n4507), .Z(n4512) );
  NAND U5440 ( .A(n4510), .B(n4509), .Z(n4511) );
  AND U5441 ( .A(n4512), .B(n4511), .Z(n4577) );
  XNOR U5442 ( .A(n4576), .B(n4577), .Z(n4579) );
  XOR U5443 ( .A(n4578), .B(n4579), .Z(n4571) );
  NAND U5444 ( .A(n4514), .B(n4513), .Z(n4518) );
  NAND U5445 ( .A(n4516), .B(n4515), .Z(n4517) );
  AND U5446 ( .A(n4518), .B(n4517), .Z(n4585) );
  NANDN U5447 ( .A(n4520), .B(n4519), .Z(n4524) );
  NANDN U5448 ( .A(n4522), .B(n4521), .Z(n4523) );
  AND U5449 ( .A(n4524), .B(n4523), .Z(n4583) );
  NANDN U5450 ( .A(n4526), .B(n4525), .Z(n4530) );
  NAND U5451 ( .A(n4528), .B(n4527), .Z(n4529) );
  AND U5452 ( .A(n4530), .B(n4529), .Z(n4650) );
  NANDN U5453 ( .A(n4531), .B(oglobal[3]), .Z(n4535) );
  NAND U5454 ( .A(n4533), .B(n4532), .Z(n4534) );
  NAND U5455 ( .A(n4535), .B(n4534), .Z(n4620) );
  NANDN U5456 ( .A(n4537), .B(n4536), .Z(n4541) );
  NAND U5457 ( .A(n4539), .B(n4538), .Z(n4540) );
  NAND U5458 ( .A(n4541), .B(n4540), .Z(n4618) );
  NANDN U5459 ( .A(n4543), .B(n4542), .Z(n4547) );
  NAND U5460 ( .A(n4545), .B(n4544), .Z(n4546) );
  NAND U5461 ( .A(n4547), .B(n4546), .Z(n4647) );
  XOR U5462 ( .A(n4648), .B(n4647), .Z(n4649) );
  XOR U5463 ( .A(n4650), .B(n4649), .Z(n4582) );
  XNOR U5464 ( .A(n4583), .B(n4582), .Z(n4584) );
  XOR U5465 ( .A(n4585), .B(n4584), .Z(n4573) );
  XNOR U5466 ( .A(n4572), .B(n4573), .Z(n4682) );
  XNOR U5467 ( .A(n4683), .B(n4682), .Z(n4666) );
  NAND U5468 ( .A(n4549), .B(n4548), .Z(n4553) );
  NAND U5469 ( .A(n4551), .B(n4550), .Z(n4552) );
  NAND U5470 ( .A(n4553), .B(n4552), .Z(n4665) );
  XNOR U5471 ( .A(n4667), .B(n4668), .Z(n4672) );
  XNOR U5472 ( .A(n4672), .B(n4671), .Z(n4557) );
  XNOR U5473 ( .A(n4673), .B(n4557), .Z(o[4]) );
  NAND U5474 ( .A(n4559), .B(n4558), .Z(n4563) );
  NAND U5475 ( .A(n4561), .B(n4560), .Z(n4562) );
  NAND U5476 ( .A(n4563), .B(n4562), .Z(n4706) );
  NAND U5477 ( .A(n4565), .B(n4564), .Z(n4569) );
  NAND U5478 ( .A(n4567), .B(n4566), .Z(n4568) );
  NAND U5479 ( .A(n4569), .B(n4568), .Z(n4722) );
  NAND U5480 ( .A(n4571), .B(n4570), .Z(n4575) );
  NANDN U5481 ( .A(n4573), .B(n4572), .Z(n4574) );
  NAND U5482 ( .A(n4575), .B(n4574), .Z(n4720) );
  NANDN U5483 ( .A(n4577), .B(n4576), .Z(n4581) );
  NAND U5484 ( .A(n4579), .B(n4578), .Z(n4580) );
  AND U5485 ( .A(n4581), .B(n4580), .Z(n4741) );
  NANDN U5486 ( .A(n4583), .B(n4582), .Z(n4587) );
  NANDN U5487 ( .A(n4585), .B(n4584), .Z(n4586) );
  AND U5488 ( .A(n4587), .B(n4586), .Z(n4739) );
  NANDN U5489 ( .A(n4589), .B(n4588), .Z(n4593) );
  NAND U5490 ( .A(n4591), .B(n4590), .Z(n4592) );
  NAND U5491 ( .A(n4593), .B(n4592), .Z(n4738) );
  XNOR U5492 ( .A(n4739), .B(n4738), .Z(n4740) );
  XNOR U5493 ( .A(n4741), .B(n4740), .Z(n4735) );
  NANDN U5494 ( .A(n4595), .B(n4594), .Z(n4599) );
  NANDN U5495 ( .A(n4597), .B(n4596), .Z(n4598) );
  AND U5496 ( .A(n4599), .B(n4598), .Z(n4759) );
  NAND U5497 ( .A(n4601), .B(n4600), .Z(n4605) );
  NAND U5498 ( .A(n4603), .B(n4602), .Z(n4604) );
  AND U5499 ( .A(n4605), .B(n4604), .Z(n4765) );
  NAND U5500 ( .A(n4607), .B(n4606), .Z(n4611) );
  NAND U5501 ( .A(n4609), .B(n4608), .Z(n4610) );
  NAND U5502 ( .A(n4611), .B(n4610), .Z(n4763) );
  NANDN U5503 ( .A(n4613), .B(n4612), .Z(n4617) );
  NAND U5504 ( .A(n4615), .B(n4614), .Z(n4616) );
  AND U5505 ( .A(n4617), .B(n4616), .Z(n4764) );
  XOR U5506 ( .A(n4763), .B(n4764), .Z(n4766) );
  NAND U5507 ( .A(n4618), .B(oglobal[4]), .Z(n4622) );
  NAND U5508 ( .A(n4620), .B(n4619), .Z(n4621) );
  NAND U5509 ( .A(n4622), .B(n4621), .Z(n4762) );
  XOR U5510 ( .A(n4762), .B(oglobal[5]), .Z(n4756) );
  XOR U5511 ( .A(n4757), .B(n4756), .Z(n4758) );
  XOR U5512 ( .A(n4759), .B(n4758), .Z(n4745) );
  NANDN U5513 ( .A(n4624), .B(n4623), .Z(n4628) );
  NANDN U5514 ( .A(n4626), .B(n4625), .Z(n4627) );
  AND U5515 ( .A(n4628), .B(n4627), .Z(n4744) );
  XNOR U5516 ( .A(n4745), .B(n4744), .Z(n4747) );
  NAND U5517 ( .A(n4630), .B(n4629), .Z(n4636) );
  AND U5518 ( .A(n4632), .B(n4631), .Z(n4633) );
  OR U5519 ( .A(n4634), .B(n4633), .Z(n4635) );
  AND U5520 ( .A(n4636), .B(n4635), .Z(n4772) );
  NAND U5521 ( .A(n4637), .B(n4638), .Z(n4643) );
  ANDN U5522 ( .B(n4639), .A(n4638), .Z(n4640) );
  OR U5523 ( .A(n4641), .B(n4640), .Z(n4642) );
  AND U5524 ( .A(n4643), .B(n4642), .Z(n4770) );
  XNOR U5525 ( .A(n4770), .B(n4769), .Z(n4771) );
  XNOR U5526 ( .A(n4772), .B(n4771), .Z(n4751) );
  NAND U5527 ( .A(n4648), .B(n4647), .Z(n4652) );
  NAND U5528 ( .A(n4650), .B(n4649), .Z(n4651) );
  NAND U5529 ( .A(n4652), .B(n4651), .Z(n4750) );
  NANDN U5530 ( .A(n4654), .B(n4653), .Z(n4658) );
  NAND U5531 ( .A(n4656), .B(n4655), .Z(n4657) );
  AND U5532 ( .A(n4658), .B(n4657), .Z(n4753) );
  XOR U5533 ( .A(n4747), .B(n4746), .Z(n4732) );
  NANDN U5534 ( .A(n4660), .B(n4659), .Z(n4664) );
  NANDN U5535 ( .A(n4662), .B(n4661), .Z(n4663) );
  NAND U5536 ( .A(n4664), .B(n4663), .Z(n4733) );
  XNOR U5537 ( .A(n4732), .B(n4733), .Z(n4734) );
  XOR U5538 ( .A(n4735), .B(n4734), .Z(n4721) );
  XNOR U5539 ( .A(n4720), .B(n4721), .Z(n4723) );
  XOR U5540 ( .A(n4722), .B(n4723), .Z(n4705) );
  XOR U5541 ( .A(n4706), .B(n4705), .Z(n4708) );
  NAND U5542 ( .A(n4666), .B(n4665), .Z(n4670) );
  NANDN U5543 ( .A(n4668), .B(n4667), .Z(n4669) );
  NAND U5544 ( .A(n4670), .B(n4669), .Z(n4707) );
  XNOR U5545 ( .A(n4708), .B(n4707), .Z(n4713) );
  NAND U5546 ( .A(n4675), .B(n4674), .Z(n4679) );
  NANDN U5547 ( .A(n4677), .B(n4676), .Z(n4678) );
  NAND U5548 ( .A(n4679), .B(n4678), .Z(n4716) );
  NANDN U5549 ( .A(n4681), .B(n4680), .Z(n4685) );
  NAND U5550 ( .A(n4683), .B(n4682), .Z(n4684) );
  AND U5551 ( .A(n4685), .B(n4684), .Z(n4715) );
  NANDN U5552 ( .A(n4687), .B(n4686), .Z(n4691) );
  NANDN U5553 ( .A(n4689), .B(n4688), .Z(n4690) );
  AND U5554 ( .A(n4691), .B(n4690), .Z(n4727) );
  NAND U5555 ( .A(n4693), .B(n4692), .Z(n4697) );
  NAND U5556 ( .A(n4695), .B(n4694), .Z(n4696) );
  AND U5557 ( .A(n4697), .B(n4696), .Z(n4726) );
  XNOR U5558 ( .A(n4727), .B(n4726), .Z(n4728) );
  NANDN U5559 ( .A(n4699), .B(n4698), .Z(n4703) );
  NANDN U5560 ( .A(n4701), .B(n4700), .Z(n4702) );
  NAND U5561 ( .A(n4703), .B(n4702), .Z(n4729) );
  XNOR U5562 ( .A(n4728), .B(n4729), .Z(n4714) );
  XOR U5563 ( .A(n4715), .B(n4714), .Z(n4717) );
  XNOR U5564 ( .A(n4716), .B(n4717), .Z(n4712) );
  XNOR U5565 ( .A(n4711), .B(n4712), .Z(n4704) );
  XNOR U5566 ( .A(n4713), .B(n4704), .Z(o[5]) );
  NAND U5567 ( .A(n4706), .B(n4705), .Z(n4710) );
  NAND U5568 ( .A(n4708), .B(n4707), .Z(n4709) );
  AND U5569 ( .A(n4710), .B(n4709), .Z(n4784) );
  NAND U5570 ( .A(n4715), .B(n4714), .Z(n4719) );
  NAND U5571 ( .A(n4717), .B(n4716), .Z(n4718) );
  NAND U5572 ( .A(n4719), .B(n4718), .Z(n4778) );
  NAND U5573 ( .A(n4721), .B(n4720), .Z(n4725) );
  NANDN U5574 ( .A(n4723), .B(n4722), .Z(n4724) );
  AND U5575 ( .A(n4725), .B(n4724), .Z(n4777) );
  NANDN U5576 ( .A(n4727), .B(n4726), .Z(n4731) );
  NANDN U5577 ( .A(n4729), .B(n4728), .Z(n4730) );
  AND U5578 ( .A(n4731), .B(n4730), .Z(n4788) );
  NANDN U5579 ( .A(n4733), .B(n4732), .Z(n4737) );
  NAND U5580 ( .A(n4735), .B(n4734), .Z(n4736) );
  AND U5581 ( .A(n4737), .B(n4736), .Z(n4786) );
  NANDN U5582 ( .A(n4739), .B(n4738), .Z(n4743) );
  NANDN U5583 ( .A(n4741), .B(n4740), .Z(n4742) );
  AND U5584 ( .A(n4743), .B(n4742), .Z(n4792) );
  NANDN U5585 ( .A(n4745), .B(n4744), .Z(n4749) );
  NAND U5586 ( .A(n4747), .B(n4746), .Z(n4748) );
  NAND U5587 ( .A(n4749), .B(n4748), .Z(n4791) );
  XNOR U5588 ( .A(n4792), .B(n4791), .Z(n4794) );
  NAND U5589 ( .A(n4751), .B(n4750), .Z(n4755) );
  NAND U5590 ( .A(n4753), .B(n4752), .Z(n4754) );
  NAND U5591 ( .A(n4755), .B(n4754), .Z(n4800) );
  NAND U5592 ( .A(n4757), .B(n4756), .Z(n4761) );
  NAND U5593 ( .A(n4759), .B(n4758), .Z(n4760) );
  AND U5594 ( .A(n4761), .B(n4760), .Z(n4805) );
  AND U5595 ( .A(oglobal[5]), .B(n4762), .Z(n4809) );
  XNOR U5596 ( .A(oglobal[6]), .B(n4809), .Z(n4804) );
  NAND U5597 ( .A(n4764), .B(n4763), .Z(n4768) );
  NAND U5598 ( .A(n4766), .B(n4765), .Z(n4767) );
  AND U5599 ( .A(n4768), .B(n4767), .Z(n4803) );
  XNOR U5600 ( .A(n4805), .B(n4806), .Z(n4797) );
  NANDN U5601 ( .A(n4770), .B(n4769), .Z(n4774) );
  NAND U5602 ( .A(n4772), .B(n4771), .Z(n4773) );
  AND U5603 ( .A(n4774), .B(n4773), .Z(n4798) );
  XOR U5604 ( .A(n4794), .B(n4793), .Z(n4785) );
  XNOR U5605 ( .A(n4786), .B(n4785), .Z(n4787) );
  XNOR U5606 ( .A(n4788), .B(n4787), .Z(n4776) );
  XOR U5607 ( .A(n4777), .B(n4776), .Z(n4779) );
  XOR U5608 ( .A(n4778), .B(n4779), .Z(n4782) );
  XNOR U5609 ( .A(n4783), .B(n4782), .Z(n4775) );
  XNOR U5610 ( .A(n4784), .B(n4775), .Z(o[6]) );
  NAND U5611 ( .A(n4777), .B(n4776), .Z(n4781) );
  NAND U5612 ( .A(n4779), .B(n4778), .Z(n4780) );
  NAND U5613 ( .A(n4781), .B(n4780), .Z(n4821) );
  NANDN U5614 ( .A(n4786), .B(n4785), .Z(n4790) );
  NAND U5615 ( .A(n4788), .B(n4787), .Z(n4789) );
  AND U5616 ( .A(n4790), .B(n4789), .Z(n4828) );
  NANDN U5617 ( .A(n4792), .B(n4791), .Z(n4796) );
  NAND U5618 ( .A(n4794), .B(n4793), .Z(n4795) );
  AND U5619 ( .A(n4796), .B(n4795), .Z(n4826) );
  NAND U5620 ( .A(n4798), .B(n4797), .Z(n4802) );
  NAND U5621 ( .A(n4800), .B(n4799), .Z(n4801) );
  NAND U5622 ( .A(n4802), .B(n4801), .Z(n4814) );
  NAND U5623 ( .A(n4804), .B(n4803), .Z(n4808) );
  NANDN U5624 ( .A(n4806), .B(n4805), .Z(n4807) );
  NAND U5625 ( .A(n4808), .B(n4807), .Z(n4813) );
  AND U5626 ( .A(n4809), .B(oglobal[6]), .Z(n4811) );
  XNOR U5627 ( .A(n4811), .B(oglobal[7]), .Z(n4812) );
  XOR U5628 ( .A(n4813), .B(n4812), .Z(n4815) );
  XOR U5629 ( .A(n4814), .B(n4815), .Z(n4825) );
  XNOR U5630 ( .A(n4826), .B(n4825), .Z(n4827) );
  XOR U5631 ( .A(n4828), .B(n4827), .Z(n4820) );
  IV U5632 ( .A(n4820), .Z(n4818) );
  XNOR U5633 ( .A(n4819), .B(n4818), .Z(n4810) );
  XNOR U5634 ( .A(n4821), .B(n4810), .Z(o[7]) );
  AND U5635 ( .A(n4811), .B(oglobal[7]), .Z(n4835) );
  XOR U5636 ( .A(oglobal[8]), .B(n4835), .Z(n4837) );
  NAND U5637 ( .A(n4813), .B(n4812), .Z(n4817) );
  NAND U5638 ( .A(n4815), .B(n4814), .Z(n4816) );
  AND U5639 ( .A(n4817), .B(n4816), .Z(n4836) );
  XNOR U5640 ( .A(n4837), .B(n4836), .Z(n4834) );
  NAND U5641 ( .A(n4818), .B(n4819), .Z(n4824) );
  ANDN U5642 ( .B(n4820), .A(n4819), .Z(n4822) );
  OR U5643 ( .A(n4822), .B(n4821), .Z(n4823) );
  AND U5644 ( .A(n4824), .B(n4823), .Z(n4832) );
  NANDN U5645 ( .A(n4826), .B(n4825), .Z(n4830) );
  NANDN U5646 ( .A(n4828), .B(n4827), .Z(n4829) );
  NAND U5647 ( .A(n4830), .B(n4829), .Z(n4833) );
  XNOR U5648 ( .A(n4832), .B(n4833), .Z(n4831) );
  XNOR U5649 ( .A(n4834), .B(n4831), .Z(o[8]) );
  XNOR U5650 ( .A(n4840), .B(oglobal[9]), .Z(n4842) );
  NAND U5651 ( .A(n4835), .B(oglobal[8]), .Z(n4839) );
  NAND U5652 ( .A(n4837), .B(n4836), .Z(n4838) );
  NAND U5653 ( .A(n4839), .B(n4838), .Z(n4841) );
  XOR U5654 ( .A(n4842), .B(n4841), .Z(o[9]) );
  ANDN U5655 ( .B(oglobal[9]), .A(n4840), .Z(n4844) );
  AND U5656 ( .A(n4842), .B(n4841), .Z(n4843) );
  NOR U5657 ( .A(n4844), .B(n4843), .Z(n4845) );
  XNOR U5658 ( .A(oglobal[10]), .B(n4845), .Z(o[10]) );
endmodule

