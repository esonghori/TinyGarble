
module first_nns_comb_W15_N128 ( q, DB, min_val_out );
  input [14:0] q;
  input [1919:0] DB;
  output [14:0] min_val_out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622;

  XOR U1921 ( .A(DB[1914]), .B(n1), .Z(min_val_out[9]) );
  AND U1922 ( .A(n2), .B(n3), .Z(n1) );
  XOR U1923 ( .A(n4), .B(n5), .Z(n3) );
  XOR U1924 ( .A(DB[1914]), .B(DB[1899]), .Z(n5) );
  AND U1925 ( .A(n6), .B(n7), .Z(n4) );
  XOR U1926 ( .A(n8), .B(n9), .Z(n7) );
  XOR U1927 ( .A(DB[1899]), .B(DB[1884]), .Z(n9) );
  AND U1928 ( .A(n10), .B(n11), .Z(n8) );
  XOR U1929 ( .A(n12), .B(n13), .Z(n11) );
  XOR U1930 ( .A(DB[1884]), .B(DB[1869]), .Z(n13) );
  AND U1931 ( .A(n14), .B(n15), .Z(n12) );
  XOR U1932 ( .A(n16), .B(n17), .Z(n15) );
  XOR U1933 ( .A(DB[1869]), .B(DB[1854]), .Z(n17) );
  AND U1934 ( .A(n18), .B(n19), .Z(n16) );
  XOR U1935 ( .A(n20), .B(n21), .Z(n19) );
  XOR U1936 ( .A(DB[1854]), .B(DB[1839]), .Z(n21) );
  AND U1937 ( .A(n22), .B(n23), .Z(n20) );
  XOR U1938 ( .A(n24), .B(n25), .Z(n23) );
  XOR U1939 ( .A(DB[1839]), .B(DB[1824]), .Z(n25) );
  AND U1940 ( .A(n26), .B(n27), .Z(n24) );
  XOR U1941 ( .A(n28), .B(n29), .Z(n27) );
  XOR U1942 ( .A(DB[1824]), .B(DB[1809]), .Z(n29) );
  AND U1943 ( .A(n30), .B(n31), .Z(n28) );
  XOR U1944 ( .A(n32), .B(n33), .Z(n31) );
  XOR U1945 ( .A(DB[1809]), .B(DB[1794]), .Z(n33) );
  AND U1946 ( .A(n34), .B(n35), .Z(n32) );
  XOR U1947 ( .A(n36), .B(n37), .Z(n35) );
  XOR U1948 ( .A(DB[1794]), .B(DB[1779]), .Z(n37) );
  AND U1949 ( .A(n38), .B(n39), .Z(n36) );
  XOR U1950 ( .A(n40), .B(n41), .Z(n39) );
  XOR U1951 ( .A(DB[1779]), .B(DB[1764]), .Z(n41) );
  AND U1952 ( .A(n42), .B(n43), .Z(n40) );
  XOR U1953 ( .A(n44), .B(n45), .Z(n43) );
  XOR U1954 ( .A(DB[1764]), .B(DB[1749]), .Z(n45) );
  AND U1955 ( .A(n46), .B(n47), .Z(n44) );
  XOR U1956 ( .A(n48), .B(n49), .Z(n47) );
  XOR U1957 ( .A(DB[1749]), .B(DB[1734]), .Z(n49) );
  AND U1958 ( .A(n50), .B(n51), .Z(n48) );
  XOR U1959 ( .A(n52), .B(n53), .Z(n51) );
  XOR U1960 ( .A(DB[1734]), .B(DB[1719]), .Z(n53) );
  AND U1961 ( .A(n54), .B(n55), .Z(n52) );
  XOR U1962 ( .A(n56), .B(n57), .Z(n55) );
  XOR U1963 ( .A(DB[1719]), .B(DB[1704]), .Z(n57) );
  AND U1964 ( .A(n58), .B(n59), .Z(n56) );
  XOR U1965 ( .A(n60), .B(n61), .Z(n59) );
  XOR U1966 ( .A(DB[1704]), .B(DB[1689]), .Z(n61) );
  AND U1967 ( .A(n62), .B(n63), .Z(n60) );
  XOR U1968 ( .A(n64), .B(n65), .Z(n63) );
  XOR U1969 ( .A(DB[1689]), .B(DB[1674]), .Z(n65) );
  AND U1970 ( .A(n66), .B(n67), .Z(n64) );
  XOR U1971 ( .A(n68), .B(n69), .Z(n67) );
  XOR U1972 ( .A(DB[1674]), .B(DB[1659]), .Z(n69) );
  AND U1973 ( .A(n70), .B(n71), .Z(n68) );
  XOR U1974 ( .A(n72), .B(n73), .Z(n71) );
  XOR U1975 ( .A(DB[1659]), .B(DB[1644]), .Z(n73) );
  AND U1976 ( .A(n74), .B(n75), .Z(n72) );
  XOR U1977 ( .A(n76), .B(n77), .Z(n75) );
  XOR U1978 ( .A(DB[1644]), .B(DB[1629]), .Z(n77) );
  AND U1979 ( .A(n78), .B(n79), .Z(n76) );
  XOR U1980 ( .A(n80), .B(n81), .Z(n79) );
  XOR U1981 ( .A(DB[1629]), .B(DB[1614]), .Z(n81) );
  AND U1982 ( .A(n82), .B(n83), .Z(n80) );
  XOR U1983 ( .A(n84), .B(n85), .Z(n83) );
  XOR U1984 ( .A(DB[1614]), .B(DB[1599]), .Z(n85) );
  AND U1985 ( .A(n86), .B(n87), .Z(n84) );
  XOR U1986 ( .A(n88), .B(n89), .Z(n87) );
  XOR U1987 ( .A(DB[1599]), .B(DB[1584]), .Z(n89) );
  AND U1988 ( .A(n90), .B(n91), .Z(n88) );
  XOR U1989 ( .A(n92), .B(n93), .Z(n91) );
  XOR U1990 ( .A(DB[1584]), .B(DB[1569]), .Z(n93) );
  AND U1991 ( .A(n94), .B(n95), .Z(n92) );
  XOR U1992 ( .A(n96), .B(n97), .Z(n95) );
  XOR U1993 ( .A(DB[1569]), .B(DB[1554]), .Z(n97) );
  AND U1994 ( .A(n98), .B(n99), .Z(n96) );
  XOR U1995 ( .A(n100), .B(n101), .Z(n99) );
  XOR U1996 ( .A(DB[1554]), .B(DB[1539]), .Z(n101) );
  AND U1997 ( .A(n102), .B(n103), .Z(n100) );
  XOR U1998 ( .A(n104), .B(n105), .Z(n103) );
  XOR U1999 ( .A(DB[1539]), .B(DB[1524]), .Z(n105) );
  AND U2000 ( .A(n106), .B(n107), .Z(n104) );
  XOR U2001 ( .A(n108), .B(n109), .Z(n107) );
  XOR U2002 ( .A(DB[1524]), .B(DB[1509]), .Z(n109) );
  AND U2003 ( .A(n110), .B(n111), .Z(n108) );
  XOR U2004 ( .A(n112), .B(n113), .Z(n111) );
  XOR U2005 ( .A(DB[1509]), .B(DB[1494]), .Z(n113) );
  AND U2006 ( .A(n114), .B(n115), .Z(n112) );
  XOR U2007 ( .A(n116), .B(n117), .Z(n115) );
  XOR U2008 ( .A(DB[1494]), .B(DB[1479]), .Z(n117) );
  AND U2009 ( .A(n118), .B(n119), .Z(n116) );
  XOR U2010 ( .A(n120), .B(n121), .Z(n119) );
  XOR U2011 ( .A(DB[1479]), .B(DB[1464]), .Z(n121) );
  AND U2012 ( .A(n122), .B(n123), .Z(n120) );
  XOR U2013 ( .A(n124), .B(n125), .Z(n123) );
  XOR U2014 ( .A(DB[1464]), .B(DB[1449]), .Z(n125) );
  AND U2015 ( .A(n126), .B(n127), .Z(n124) );
  XOR U2016 ( .A(n128), .B(n129), .Z(n127) );
  XOR U2017 ( .A(DB[1449]), .B(DB[1434]), .Z(n129) );
  AND U2018 ( .A(n130), .B(n131), .Z(n128) );
  XOR U2019 ( .A(n132), .B(n133), .Z(n131) );
  XOR U2020 ( .A(DB[1434]), .B(DB[1419]), .Z(n133) );
  AND U2021 ( .A(n134), .B(n135), .Z(n132) );
  XOR U2022 ( .A(n136), .B(n137), .Z(n135) );
  XOR U2023 ( .A(DB[1419]), .B(DB[1404]), .Z(n137) );
  AND U2024 ( .A(n138), .B(n139), .Z(n136) );
  XOR U2025 ( .A(n140), .B(n141), .Z(n139) );
  XOR U2026 ( .A(DB[1404]), .B(DB[1389]), .Z(n141) );
  AND U2027 ( .A(n142), .B(n143), .Z(n140) );
  XOR U2028 ( .A(n144), .B(n145), .Z(n143) );
  XOR U2029 ( .A(DB[1389]), .B(DB[1374]), .Z(n145) );
  AND U2030 ( .A(n146), .B(n147), .Z(n144) );
  XOR U2031 ( .A(n148), .B(n149), .Z(n147) );
  XOR U2032 ( .A(DB[1374]), .B(DB[1359]), .Z(n149) );
  AND U2033 ( .A(n150), .B(n151), .Z(n148) );
  XOR U2034 ( .A(n152), .B(n153), .Z(n151) );
  XOR U2035 ( .A(DB[1359]), .B(DB[1344]), .Z(n153) );
  AND U2036 ( .A(n154), .B(n155), .Z(n152) );
  XOR U2037 ( .A(n156), .B(n157), .Z(n155) );
  XOR U2038 ( .A(DB[1344]), .B(DB[1329]), .Z(n157) );
  AND U2039 ( .A(n158), .B(n159), .Z(n156) );
  XOR U2040 ( .A(n160), .B(n161), .Z(n159) );
  XOR U2041 ( .A(DB[1329]), .B(DB[1314]), .Z(n161) );
  AND U2042 ( .A(n162), .B(n163), .Z(n160) );
  XOR U2043 ( .A(n164), .B(n165), .Z(n163) );
  XOR U2044 ( .A(DB[1314]), .B(DB[1299]), .Z(n165) );
  AND U2045 ( .A(n166), .B(n167), .Z(n164) );
  XOR U2046 ( .A(n168), .B(n169), .Z(n167) );
  XOR U2047 ( .A(DB[1299]), .B(DB[1284]), .Z(n169) );
  AND U2048 ( .A(n170), .B(n171), .Z(n168) );
  XOR U2049 ( .A(n172), .B(n173), .Z(n171) );
  XOR U2050 ( .A(DB[1284]), .B(DB[1269]), .Z(n173) );
  AND U2051 ( .A(n174), .B(n175), .Z(n172) );
  XOR U2052 ( .A(n176), .B(n177), .Z(n175) );
  XOR U2053 ( .A(DB[1269]), .B(DB[1254]), .Z(n177) );
  AND U2054 ( .A(n178), .B(n179), .Z(n176) );
  XOR U2055 ( .A(n180), .B(n181), .Z(n179) );
  XOR U2056 ( .A(DB[1254]), .B(DB[1239]), .Z(n181) );
  AND U2057 ( .A(n182), .B(n183), .Z(n180) );
  XOR U2058 ( .A(n184), .B(n185), .Z(n183) );
  XOR U2059 ( .A(DB[1239]), .B(DB[1224]), .Z(n185) );
  AND U2060 ( .A(n186), .B(n187), .Z(n184) );
  XOR U2061 ( .A(n188), .B(n189), .Z(n187) );
  XOR U2062 ( .A(DB[1224]), .B(DB[1209]), .Z(n189) );
  AND U2063 ( .A(n190), .B(n191), .Z(n188) );
  XOR U2064 ( .A(n192), .B(n193), .Z(n191) );
  XOR U2065 ( .A(DB[1209]), .B(DB[1194]), .Z(n193) );
  AND U2066 ( .A(n194), .B(n195), .Z(n192) );
  XOR U2067 ( .A(n196), .B(n197), .Z(n195) );
  XOR U2068 ( .A(DB[1194]), .B(DB[1179]), .Z(n197) );
  AND U2069 ( .A(n198), .B(n199), .Z(n196) );
  XOR U2070 ( .A(n200), .B(n201), .Z(n199) );
  XOR U2071 ( .A(DB[1179]), .B(DB[1164]), .Z(n201) );
  AND U2072 ( .A(n202), .B(n203), .Z(n200) );
  XOR U2073 ( .A(n204), .B(n205), .Z(n203) );
  XOR U2074 ( .A(DB[1164]), .B(DB[1149]), .Z(n205) );
  AND U2075 ( .A(n206), .B(n207), .Z(n204) );
  XOR U2076 ( .A(n208), .B(n209), .Z(n207) );
  XOR U2077 ( .A(DB[1149]), .B(DB[1134]), .Z(n209) );
  AND U2078 ( .A(n210), .B(n211), .Z(n208) );
  XOR U2079 ( .A(n212), .B(n213), .Z(n211) );
  XOR U2080 ( .A(DB[1134]), .B(DB[1119]), .Z(n213) );
  AND U2081 ( .A(n214), .B(n215), .Z(n212) );
  XOR U2082 ( .A(n216), .B(n217), .Z(n215) );
  XOR U2083 ( .A(DB[1119]), .B(DB[1104]), .Z(n217) );
  AND U2084 ( .A(n218), .B(n219), .Z(n216) );
  XOR U2085 ( .A(n220), .B(n221), .Z(n219) );
  XOR U2086 ( .A(DB[1104]), .B(DB[1089]), .Z(n221) );
  AND U2087 ( .A(n222), .B(n223), .Z(n220) );
  XOR U2088 ( .A(n224), .B(n225), .Z(n223) );
  XOR U2089 ( .A(DB[1089]), .B(DB[1074]), .Z(n225) );
  AND U2090 ( .A(n226), .B(n227), .Z(n224) );
  XOR U2091 ( .A(n228), .B(n229), .Z(n227) );
  XOR U2092 ( .A(DB[1074]), .B(DB[1059]), .Z(n229) );
  AND U2093 ( .A(n230), .B(n231), .Z(n228) );
  XOR U2094 ( .A(n232), .B(n233), .Z(n231) );
  XOR U2095 ( .A(DB[1059]), .B(DB[1044]), .Z(n233) );
  AND U2096 ( .A(n234), .B(n235), .Z(n232) );
  XOR U2097 ( .A(n236), .B(n237), .Z(n235) );
  XOR U2098 ( .A(DB[1044]), .B(DB[1029]), .Z(n237) );
  AND U2099 ( .A(n238), .B(n239), .Z(n236) );
  XOR U2100 ( .A(n240), .B(n241), .Z(n239) );
  XOR U2101 ( .A(DB[1029]), .B(DB[1014]), .Z(n241) );
  AND U2102 ( .A(n242), .B(n243), .Z(n240) );
  XOR U2103 ( .A(n244), .B(n245), .Z(n243) );
  XOR U2104 ( .A(DB[999]), .B(DB[1014]), .Z(n245) );
  AND U2105 ( .A(n246), .B(n247), .Z(n244) );
  XOR U2106 ( .A(n248), .B(n249), .Z(n247) );
  XOR U2107 ( .A(DB[999]), .B(DB[984]), .Z(n249) );
  AND U2108 ( .A(n250), .B(n251), .Z(n248) );
  XOR U2109 ( .A(n252), .B(n253), .Z(n251) );
  XOR U2110 ( .A(DB[984]), .B(DB[969]), .Z(n253) );
  AND U2111 ( .A(n254), .B(n255), .Z(n252) );
  XOR U2112 ( .A(n256), .B(n257), .Z(n255) );
  XOR U2113 ( .A(DB[969]), .B(DB[954]), .Z(n257) );
  AND U2114 ( .A(n258), .B(n259), .Z(n256) );
  XOR U2115 ( .A(n260), .B(n261), .Z(n259) );
  XOR U2116 ( .A(DB[954]), .B(DB[939]), .Z(n261) );
  AND U2117 ( .A(n262), .B(n263), .Z(n260) );
  XOR U2118 ( .A(n264), .B(n265), .Z(n263) );
  XOR U2119 ( .A(DB[939]), .B(DB[924]), .Z(n265) );
  AND U2120 ( .A(n266), .B(n267), .Z(n264) );
  XOR U2121 ( .A(n268), .B(n269), .Z(n267) );
  XOR U2122 ( .A(DB[924]), .B(DB[909]), .Z(n269) );
  AND U2123 ( .A(n270), .B(n271), .Z(n268) );
  XOR U2124 ( .A(n272), .B(n273), .Z(n271) );
  XOR U2125 ( .A(DB[909]), .B(DB[894]), .Z(n273) );
  AND U2126 ( .A(n274), .B(n275), .Z(n272) );
  XOR U2127 ( .A(n276), .B(n277), .Z(n275) );
  XOR U2128 ( .A(DB[894]), .B(DB[879]), .Z(n277) );
  AND U2129 ( .A(n278), .B(n279), .Z(n276) );
  XOR U2130 ( .A(n280), .B(n281), .Z(n279) );
  XOR U2131 ( .A(DB[879]), .B(DB[864]), .Z(n281) );
  AND U2132 ( .A(n282), .B(n283), .Z(n280) );
  XOR U2133 ( .A(n284), .B(n285), .Z(n283) );
  XOR U2134 ( .A(DB[864]), .B(DB[849]), .Z(n285) );
  AND U2135 ( .A(n286), .B(n287), .Z(n284) );
  XOR U2136 ( .A(n288), .B(n289), .Z(n287) );
  XOR U2137 ( .A(DB[849]), .B(DB[834]), .Z(n289) );
  AND U2138 ( .A(n290), .B(n291), .Z(n288) );
  XOR U2139 ( .A(n292), .B(n293), .Z(n291) );
  XOR U2140 ( .A(DB[834]), .B(DB[819]), .Z(n293) );
  AND U2141 ( .A(n294), .B(n295), .Z(n292) );
  XOR U2142 ( .A(n296), .B(n297), .Z(n295) );
  XOR U2143 ( .A(DB[819]), .B(DB[804]), .Z(n297) );
  AND U2144 ( .A(n298), .B(n299), .Z(n296) );
  XOR U2145 ( .A(n300), .B(n301), .Z(n299) );
  XOR U2146 ( .A(DB[804]), .B(DB[789]), .Z(n301) );
  AND U2147 ( .A(n302), .B(n303), .Z(n300) );
  XOR U2148 ( .A(n304), .B(n305), .Z(n303) );
  XOR U2149 ( .A(DB[789]), .B(DB[774]), .Z(n305) );
  AND U2150 ( .A(n306), .B(n307), .Z(n304) );
  XOR U2151 ( .A(n308), .B(n309), .Z(n307) );
  XOR U2152 ( .A(DB[774]), .B(DB[759]), .Z(n309) );
  AND U2153 ( .A(n310), .B(n311), .Z(n308) );
  XOR U2154 ( .A(n312), .B(n313), .Z(n311) );
  XOR U2155 ( .A(DB[759]), .B(DB[744]), .Z(n313) );
  AND U2156 ( .A(n314), .B(n315), .Z(n312) );
  XOR U2157 ( .A(n316), .B(n317), .Z(n315) );
  XOR U2158 ( .A(DB[744]), .B(DB[729]), .Z(n317) );
  AND U2159 ( .A(n318), .B(n319), .Z(n316) );
  XOR U2160 ( .A(n320), .B(n321), .Z(n319) );
  XOR U2161 ( .A(DB[729]), .B(DB[714]), .Z(n321) );
  AND U2162 ( .A(n322), .B(n323), .Z(n320) );
  XOR U2163 ( .A(n324), .B(n325), .Z(n323) );
  XOR U2164 ( .A(DB[714]), .B(DB[699]), .Z(n325) );
  AND U2165 ( .A(n326), .B(n327), .Z(n324) );
  XOR U2166 ( .A(n328), .B(n329), .Z(n327) );
  XOR U2167 ( .A(DB[699]), .B(DB[684]), .Z(n329) );
  AND U2168 ( .A(n330), .B(n331), .Z(n328) );
  XOR U2169 ( .A(n332), .B(n333), .Z(n331) );
  XOR U2170 ( .A(DB[684]), .B(DB[669]), .Z(n333) );
  AND U2171 ( .A(n334), .B(n335), .Z(n332) );
  XOR U2172 ( .A(n336), .B(n337), .Z(n335) );
  XOR U2173 ( .A(DB[669]), .B(DB[654]), .Z(n337) );
  AND U2174 ( .A(n338), .B(n339), .Z(n336) );
  XOR U2175 ( .A(n340), .B(n341), .Z(n339) );
  XOR U2176 ( .A(DB[654]), .B(DB[639]), .Z(n341) );
  AND U2177 ( .A(n342), .B(n343), .Z(n340) );
  XOR U2178 ( .A(n344), .B(n345), .Z(n343) );
  XOR U2179 ( .A(DB[639]), .B(DB[624]), .Z(n345) );
  AND U2180 ( .A(n346), .B(n347), .Z(n344) );
  XOR U2181 ( .A(n348), .B(n349), .Z(n347) );
  XOR U2182 ( .A(DB[624]), .B(DB[609]), .Z(n349) );
  AND U2183 ( .A(n350), .B(n351), .Z(n348) );
  XOR U2184 ( .A(n352), .B(n353), .Z(n351) );
  XOR U2185 ( .A(DB[609]), .B(DB[594]), .Z(n353) );
  AND U2186 ( .A(n354), .B(n355), .Z(n352) );
  XOR U2187 ( .A(n356), .B(n357), .Z(n355) );
  XOR U2188 ( .A(DB[594]), .B(DB[579]), .Z(n357) );
  AND U2189 ( .A(n358), .B(n359), .Z(n356) );
  XOR U2190 ( .A(n360), .B(n361), .Z(n359) );
  XOR U2191 ( .A(DB[579]), .B(DB[564]), .Z(n361) );
  AND U2192 ( .A(n362), .B(n363), .Z(n360) );
  XOR U2193 ( .A(n364), .B(n365), .Z(n363) );
  XOR U2194 ( .A(DB[564]), .B(DB[549]), .Z(n365) );
  AND U2195 ( .A(n366), .B(n367), .Z(n364) );
  XOR U2196 ( .A(n368), .B(n369), .Z(n367) );
  XOR U2197 ( .A(DB[549]), .B(DB[534]), .Z(n369) );
  AND U2198 ( .A(n370), .B(n371), .Z(n368) );
  XOR U2199 ( .A(n372), .B(n373), .Z(n371) );
  XOR U2200 ( .A(DB[534]), .B(DB[519]), .Z(n373) );
  AND U2201 ( .A(n374), .B(n375), .Z(n372) );
  XOR U2202 ( .A(n376), .B(n377), .Z(n375) );
  XOR U2203 ( .A(DB[519]), .B(DB[504]), .Z(n377) );
  AND U2204 ( .A(n378), .B(n379), .Z(n376) );
  XOR U2205 ( .A(n380), .B(n381), .Z(n379) );
  XOR U2206 ( .A(DB[504]), .B(DB[489]), .Z(n381) );
  AND U2207 ( .A(n382), .B(n383), .Z(n380) );
  XOR U2208 ( .A(n384), .B(n385), .Z(n383) );
  XOR U2209 ( .A(DB[489]), .B(DB[474]), .Z(n385) );
  AND U2210 ( .A(n386), .B(n387), .Z(n384) );
  XOR U2211 ( .A(n388), .B(n389), .Z(n387) );
  XOR U2212 ( .A(DB[474]), .B(DB[459]), .Z(n389) );
  AND U2213 ( .A(n390), .B(n391), .Z(n388) );
  XOR U2214 ( .A(n392), .B(n393), .Z(n391) );
  XOR U2215 ( .A(DB[459]), .B(DB[444]), .Z(n393) );
  AND U2216 ( .A(n394), .B(n395), .Z(n392) );
  XOR U2217 ( .A(n396), .B(n397), .Z(n395) );
  XOR U2218 ( .A(DB[444]), .B(DB[429]), .Z(n397) );
  AND U2219 ( .A(n398), .B(n399), .Z(n396) );
  XOR U2220 ( .A(n400), .B(n401), .Z(n399) );
  XOR U2221 ( .A(DB[429]), .B(DB[414]), .Z(n401) );
  AND U2222 ( .A(n402), .B(n403), .Z(n400) );
  XOR U2223 ( .A(n404), .B(n405), .Z(n403) );
  XOR U2224 ( .A(DB[414]), .B(DB[399]), .Z(n405) );
  AND U2225 ( .A(n406), .B(n407), .Z(n404) );
  XOR U2226 ( .A(n408), .B(n409), .Z(n407) );
  XOR U2227 ( .A(DB[399]), .B(DB[384]), .Z(n409) );
  AND U2228 ( .A(n410), .B(n411), .Z(n408) );
  XOR U2229 ( .A(n412), .B(n413), .Z(n411) );
  XOR U2230 ( .A(DB[384]), .B(DB[369]), .Z(n413) );
  AND U2231 ( .A(n414), .B(n415), .Z(n412) );
  XOR U2232 ( .A(n416), .B(n417), .Z(n415) );
  XOR U2233 ( .A(DB[369]), .B(DB[354]), .Z(n417) );
  AND U2234 ( .A(n418), .B(n419), .Z(n416) );
  XOR U2235 ( .A(n420), .B(n421), .Z(n419) );
  XOR U2236 ( .A(DB[354]), .B(DB[339]), .Z(n421) );
  AND U2237 ( .A(n422), .B(n423), .Z(n420) );
  XOR U2238 ( .A(n424), .B(n425), .Z(n423) );
  XOR U2239 ( .A(DB[339]), .B(DB[324]), .Z(n425) );
  AND U2240 ( .A(n426), .B(n427), .Z(n424) );
  XOR U2241 ( .A(n428), .B(n429), .Z(n427) );
  XOR U2242 ( .A(DB[324]), .B(DB[309]), .Z(n429) );
  AND U2243 ( .A(n430), .B(n431), .Z(n428) );
  XOR U2244 ( .A(n432), .B(n433), .Z(n431) );
  XOR U2245 ( .A(DB[309]), .B(DB[294]), .Z(n433) );
  AND U2246 ( .A(n434), .B(n435), .Z(n432) );
  XOR U2247 ( .A(n436), .B(n437), .Z(n435) );
  XOR U2248 ( .A(DB[294]), .B(DB[279]), .Z(n437) );
  AND U2249 ( .A(n438), .B(n439), .Z(n436) );
  XOR U2250 ( .A(n440), .B(n441), .Z(n439) );
  XOR U2251 ( .A(DB[279]), .B(DB[264]), .Z(n441) );
  AND U2252 ( .A(n442), .B(n443), .Z(n440) );
  XOR U2253 ( .A(n444), .B(n445), .Z(n443) );
  XOR U2254 ( .A(DB[264]), .B(DB[249]), .Z(n445) );
  AND U2255 ( .A(n446), .B(n447), .Z(n444) );
  XOR U2256 ( .A(n448), .B(n449), .Z(n447) );
  XOR U2257 ( .A(DB[249]), .B(DB[234]), .Z(n449) );
  AND U2258 ( .A(n450), .B(n451), .Z(n448) );
  XOR U2259 ( .A(n452), .B(n453), .Z(n451) );
  XOR U2260 ( .A(DB[234]), .B(DB[219]), .Z(n453) );
  AND U2261 ( .A(n454), .B(n455), .Z(n452) );
  XOR U2262 ( .A(n456), .B(n457), .Z(n455) );
  XOR U2263 ( .A(DB[219]), .B(DB[204]), .Z(n457) );
  AND U2264 ( .A(n458), .B(n459), .Z(n456) );
  XOR U2265 ( .A(n460), .B(n461), .Z(n459) );
  XOR U2266 ( .A(DB[204]), .B(DB[189]), .Z(n461) );
  AND U2267 ( .A(n462), .B(n463), .Z(n460) );
  XOR U2268 ( .A(n464), .B(n465), .Z(n463) );
  XOR U2269 ( .A(DB[189]), .B(DB[174]), .Z(n465) );
  AND U2270 ( .A(n466), .B(n467), .Z(n464) );
  XOR U2271 ( .A(n468), .B(n469), .Z(n467) );
  XOR U2272 ( .A(DB[174]), .B(DB[159]), .Z(n469) );
  AND U2273 ( .A(n470), .B(n471), .Z(n468) );
  XOR U2274 ( .A(n472), .B(n473), .Z(n471) );
  XOR U2275 ( .A(DB[159]), .B(DB[144]), .Z(n473) );
  AND U2276 ( .A(n474), .B(n475), .Z(n472) );
  XOR U2277 ( .A(n476), .B(n477), .Z(n475) );
  XOR U2278 ( .A(DB[144]), .B(DB[129]), .Z(n477) );
  AND U2279 ( .A(n478), .B(n479), .Z(n476) );
  XOR U2280 ( .A(n480), .B(n481), .Z(n479) );
  XOR U2281 ( .A(DB[129]), .B(DB[114]), .Z(n481) );
  AND U2282 ( .A(n482), .B(n483), .Z(n480) );
  XOR U2283 ( .A(n484), .B(n485), .Z(n483) );
  XOR U2284 ( .A(DB[99]), .B(DB[114]), .Z(n485) );
  AND U2285 ( .A(n486), .B(n487), .Z(n484) );
  XOR U2286 ( .A(n488), .B(n489), .Z(n487) );
  XOR U2287 ( .A(DB[99]), .B(DB[84]), .Z(n489) );
  AND U2288 ( .A(n490), .B(n491), .Z(n488) );
  XOR U2289 ( .A(n492), .B(n493), .Z(n491) );
  XOR U2290 ( .A(DB[84]), .B(DB[69]), .Z(n493) );
  AND U2291 ( .A(n494), .B(n495), .Z(n492) );
  XOR U2292 ( .A(n496), .B(n497), .Z(n495) );
  XOR U2293 ( .A(DB[69]), .B(DB[54]), .Z(n497) );
  AND U2294 ( .A(n498), .B(n499), .Z(n496) );
  XOR U2295 ( .A(n500), .B(n501), .Z(n499) );
  XOR U2296 ( .A(DB[54]), .B(DB[39]), .Z(n501) );
  AND U2297 ( .A(n502), .B(n503), .Z(n500) );
  XOR U2298 ( .A(n504), .B(n505), .Z(n503) );
  XOR U2299 ( .A(DB[39]), .B(DB[24]), .Z(n505) );
  AND U2300 ( .A(n506), .B(n507), .Z(n504) );
  XOR U2301 ( .A(DB[9]), .B(DB[24]), .Z(n507) );
  XOR U2302 ( .A(DB[1913]), .B(n508), .Z(min_val_out[8]) );
  AND U2303 ( .A(n2), .B(n509), .Z(n508) );
  XOR U2304 ( .A(n510), .B(n511), .Z(n509) );
  XOR U2305 ( .A(DB[1913]), .B(DB[1898]), .Z(n511) );
  AND U2306 ( .A(n6), .B(n512), .Z(n510) );
  XOR U2307 ( .A(n513), .B(n514), .Z(n512) );
  XOR U2308 ( .A(DB[1898]), .B(DB[1883]), .Z(n514) );
  AND U2309 ( .A(n10), .B(n515), .Z(n513) );
  XOR U2310 ( .A(n516), .B(n517), .Z(n515) );
  XOR U2311 ( .A(DB[1883]), .B(DB[1868]), .Z(n517) );
  AND U2312 ( .A(n14), .B(n518), .Z(n516) );
  XOR U2313 ( .A(n519), .B(n520), .Z(n518) );
  XOR U2314 ( .A(DB[1868]), .B(DB[1853]), .Z(n520) );
  AND U2315 ( .A(n18), .B(n521), .Z(n519) );
  XOR U2316 ( .A(n522), .B(n523), .Z(n521) );
  XOR U2317 ( .A(DB[1853]), .B(DB[1838]), .Z(n523) );
  AND U2318 ( .A(n22), .B(n524), .Z(n522) );
  XOR U2319 ( .A(n525), .B(n526), .Z(n524) );
  XOR U2320 ( .A(DB[1838]), .B(DB[1823]), .Z(n526) );
  AND U2321 ( .A(n26), .B(n527), .Z(n525) );
  XOR U2322 ( .A(n528), .B(n529), .Z(n527) );
  XOR U2323 ( .A(DB[1823]), .B(DB[1808]), .Z(n529) );
  AND U2324 ( .A(n30), .B(n530), .Z(n528) );
  XOR U2325 ( .A(n531), .B(n532), .Z(n530) );
  XOR U2326 ( .A(DB[1808]), .B(DB[1793]), .Z(n532) );
  AND U2327 ( .A(n34), .B(n533), .Z(n531) );
  XOR U2328 ( .A(n534), .B(n535), .Z(n533) );
  XOR U2329 ( .A(DB[1793]), .B(DB[1778]), .Z(n535) );
  AND U2330 ( .A(n38), .B(n536), .Z(n534) );
  XOR U2331 ( .A(n537), .B(n538), .Z(n536) );
  XOR U2332 ( .A(DB[1778]), .B(DB[1763]), .Z(n538) );
  AND U2333 ( .A(n42), .B(n539), .Z(n537) );
  XOR U2334 ( .A(n540), .B(n541), .Z(n539) );
  XOR U2335 ( .A(DB[1763]), .B(DB[1748]), .Z(n541) );
  AND U2336 ( .A(n46), .B(n542), .Z(n540) );
  XOR U2337 ( .A(n543), .B(n544), .Z(n542) );
  XOR U2338 ( .A(DB[1748]), .B(DB[1733]), .Z(n544) );
  AND U2339 ( .A(n50), .B(n545), .Z(n543) );
  XOR U2340 ( .A(n546), .B(n547), .Z(n545) );
  XOR U2341 ( .A(DB[1733]), .B(DB[1718]), .Z(n547) );
  AND U2342 ( .A(n54), .B(n548), .Z(n546) );
  XOR U2343 ( .A(n549), .B(n550), .Z(n548) );
  XOR U2344 ( .A(DB[1718]), .B(DB[1703]), .Z(n550) );
  AND U2345 ( .A(n58), .B(n551), .Z(n549) );
  XOR U2346 ( .A(n552), .B(n553), .Z(n551) );
  XOR U2347 ( .A(DB[1703]), .B(DB[1688]), .Z(n553) );
  AND U2348 ( .A(n62), .B(n554), .Z(n552) );
  XOR U2349 ( .A(n555), .B(n556), .Z(n554) );
  XOR U2350 ( .A(DB[1688]), .B(DB[1673]), .Z(n556) );
  AND U2351 ( .A(n66), .B(n557), .Z(n555) );
  XOR U2352 ( .A(n558), .B(n559), .Z(n557) );
  XOR U2353 ( .A(DB[1673]), .B(DB[1658]), .Z(n559) );
  AND U2354 ( .A(n70), .B(n560), .Z(n558) );
  XOR U2355 ( .A(n561), .B(n562), .Z(n560) );
  XOR U2356 ( .A(DB[1658]), .B(DB[1643]), .Z(n562) );
  AND U2357 ( .A(n74), .B(n563), .Z(n561) );
  XOR U2358 ( .A(n564), .B(n565), .Z(n563) );
  XOR U2359 ( .A(DB[1643]), .B(DB[1628]), .Z(n565) );
  AND U2360 ( .A(n78), .B(n566), .Z(n564) );
  XOR U2361 ( .A(n567), .B(n568), .Z(n566) );
  XOR U2362 ( .A(DB[1628]), .B(DB[1613]), .Z(n568) );
  AND U2363 ( .A(n82), .B(n569), .Z(n567) );
  XOR U2364 ( .A(n570), .B(n571), .Z(n569) );
  XOR U2365 ( .A(DB[1613]), .B(DB[1598]), .Z(n571) );
  AND U2366 ( .A(n86), .B(n572), .Z(n570) );
  XOR U2367 ( .A(n573), .B(n574), .Z(n572) );
  XOR U2368 ( .A(DB[1598]), .B(DB[1583]), .Z(n574) );
  AND U2369 ( .A(n90), .B(n575), .Z(n573) );
  XOR U2370 ( .A(n576), .B(n577), .Z(n575) );
  XOR U2371 ( .A(DB[1583]), .B(DB[1568]), .Z(n577) );
  AND U2372 ( .A(n94), .B(n578), .Z(n576) );
  XOR U2373 ( .A(n579), .B(n580), .Z(n578) );
  XOR U2374 ( .A(DB[1568]), .B(DB[1553]), .Z(n580) );
  AND U2375 ( .A(n98), .B(n581), .Z(n579) );
  XOR U2376 ( .A(n582), .B(n583), .Z(n581) );
  XOR U2377 ( .A(DB[1553]), .B(DB[1538]), .Z(n583) );
  AND U2378 ( .A(n102), .B(n584), .Z(n582) );
  XOR U2379 ( .A(n585), .B(n586), .Z(n584) );
  XOR U2380 ( .A(DB[1538]), .B(DB[1523]), .Z(n586) );
  AND U2381 ( .A(n106), .B(n587), .Z(n585) );
  XOR U2382 ( .A(n588), .B(n589), .Z(n587) );
  XOR U2383 ( .A(DB[1523]), .B(DB[1508]), .Z(n589) );
  AND U2384 ( .A(n110), .B(n590), .Z(n588) );
  XOR U2385 ( .A(n591), .B(n592), .Z(n590) );
  XOR U2386 ( .A(DB[1508]), .B(DB[1493]), .Z(n592) );
  AND U2387 ( .A(n114), .B(n593), .Z(n591) );
  XOR U2388 ( .A(n594), .B(n595), .Z(n593) );
  XOR U2389 ( .A(DB[1493]), .B(DB[1478]), .Z(n595) );
  AND U2390 ( .A(n118), .B(n596), .Z(n594) );
  XOR U2391 ( .A(n597), .B(n598), .Z(n596) );
  XOR U2392 ( .A(DB[1478]), .B(DB[1463]), .Z(n598) );
  AND U2393 ( .A(n122), .B(n599), .Z(n597) );
  XOR U2394 ( .A(n600), .B(n601), .Z(n599) );
  XOR U2395 ( .A(DB[1463]), .B(DB[1448]), .Z(n601) );
  AND U2396 ( .A(n126), .B(n602), .Z(n600) );
  XOR U2397 ( .A(n603), .B(n604), .Z(n602) );
  XOR U2398 ( .A(DB[1448]), .B(DB[1433]), .Z(n604) );
  AND U2399 ( .A(n130), .B(n605), .Z(n603) );
  XOR U2400 ( .A(n606), .B(n607), .Z(n605) );
  XOR U2401 ( .A(DB[1433]), .B(DB[1418]), .Z(n607) );
  AND U2402 ( .A(n134), .B(n608), .Z(n606) );
  XOR U2403 ( .A(n609), .B(n610), .Z(n608) );
  XOR U2404 ( .A(DB[1418]), .B(DB[1403]), .Z(n610) );
  AND U2405 ( .A(n138), .B(n611), .Z(n609) );
  XOR U2406 ( .A(n612), .B(n613), .Z(n611) );
  XOR U2407 ( .A(DB[1403]), .B(DB[1388]), .Z(n613) );
  AND U2408 ( .A(n142), .B(n614), .Z(n612) );
  XOR U2409 ( .A(n615), .B(n616), .Z(n614) );
  XOR U2410 ( .A(DB[1388]), .B(DB[1373]), .Z(n616) );
  AND U2411 ( .A(n146), .B(n617), .Z(n615) );
  XOR U2412 ( .A(n618), .B(n619), .Z(n617) );
  XOR U2413 ( .A(DB[1373]), .B(DB[1358]), .Z(n619) );
  AND U2414 ( .A(n150), .B(n620), .Z(n618) );
  XOR U2415 ( .A(n621), .B(n622), .Z(n620) );
  XOR U2416 ( .A(DB[1358]), .B(DB[1343]), .Z(n622) );
  AND U2417 ( .A(n154), .B(n623), .Z(n621) );
  XOR U2418 ( .A(n624), .B(n625), .Z(n623) );
  XOR U2419 ( .A(DB[1343]), .B(DB[1328]), .Z(n625) );
  AND U2420 ( .A(n158), .B(n626), .Z(n624) );
  XOR U2421 ( .A(n627), .B(n628), .Z(n626) );
  XOR U2422 ( .A(DB[1328]), .B(DB[1313]), .Z(n628) );
  AND U2423 ( .A(n162), .B(n629), .Z(n627) );
  XOR U2424 ( .A(n630), .B(n631), .Z(n629) );
  XOR U2425 ( .A(DB[1313]), .B(DB[1298]), .Z(n631) );
  AND U2426 ( .A(n166), .B(n632), .Z(n630) );
  XOR U2427 ( .A(n633), .B(n634), .Z(n632) );
  XOR U2428 ( .A(DB[1298]), .B(DB[1283]), .Z(n634) );
  AND U2429 ( .A(n170), .B(n635), .Z(n633) );
  XOR U2430 ( .A(n636), .B(n637), .Z(n635) );
  XOR U2431 ( .A(DB[1283]), .B(DB[1268]), .Z(n637) );
  AND U2432 ( .A(n174), .B(n638), .Z(n636) );
  XOR U2433 ( .A(n639), .B(n640), .Z(n638) );
  XOR U2434 ( .A(DB[1268]), .B(DB[1253]), .Z(n640) );
  AND U2435 ( .A(n178), .B(n641), .Z(n639) );
  XOR U2436 ( .A(n642), .B(n643), .Z(n641) );
  XOR U2437 ( .A(DB[1253]), .B(DB[1238]), .Z(n643) );
  AND U2438 ( .A(n182), .B(n644), .Z(n642) );
  XOR U2439 ( .A(n645), .B(n646), .Z(n644) );
  XOR U2440 ( .A(DB[1238]), .B(DB[1223]), .Z(n646) );
  AND U2441 ( .A(n186), .B(n647), .Z(n645) );
  XOR U2442 ( .A(n648), .B(n649), .Z(n647) );
  XOR U2443 ( .A(DB[1223]), .B(DB[1208]), .Z(n649) );
  AND U2444 ( .A(n190), .B(n650), .Z(n648) );
  XOR U2445 ( .A(n651), .B(n652), .Z(n650) );
  XOR U2446 ( .A(DB[1208]), .B(DB[1193]), .Z(n652) );
  AND U2447 ( .A(n194), .B(n653), .Z(n651) );
  XOR U2448 ( .A(n654), .B(n655), .Z(n653) );
  XOR U2449 ( .A(DB[1193]), .B(DB[1178]), .Z(n655) );
  AND U2450 ( .A(n198), .B(n656), .Z(n654) );
  XOR U2451 ( .A(n657), .B(n658), .Z(n656) );
  XOR U2452 ( .A(DB[1178]), .B(DB[1163]), .Z(n658) );
  AND U2453 ( .A(n202), .B(n659), .Z(n657) );
  XOR U2454 ( .A(n660), .B(n661), .Z(n659) );
  XOR U2455 ( .A(DB[1163]), .B(DB[1148]), .Z(n661) );
  AND U2456 ( .A(n206), .B(n662), .Z(n660) );
  XOR U2457 ( .A(n663), .B(n664), .Z(n662) );
  XOR U2458 ( .A(DB[1148]), .B(DB[1133]), .Z(n664) );
  AND U2459 ( .A(n210), .B(n665), .Z(n663) );
  XOR U2460 ( .A(n666), .B(n667), .Z(n665) );
  XOR U2461 ( .A(DB[1133]), .B(DB[1118]), .Z(n667) );
  AND U2462 ( .A(n214), .B(n668), .Z(n666) );
  XOR U2463 ( .A(n669), .B(n670), .Z(n668) );
  XOR U2464 ( .A(DB[1118]), .B(DB[1103]), .Z(n670) );
  AND U2465 ( .A(n218), .B(n671), .Z(n669) );
  XOR U2466 ( .A(n672), .B(n673), .Z(n671) );
  XOR U2467 ( .A(DB[1103]), .B(DB[1088]), .Z(n673) );
  AND U2468 ( .A(n222), .B(n674), .Z(n672) );
  XOR U2469 ( .A(n675), .B(n676), .Z(n674) );
  XOR U2470 ( .A(DB[1088]), .B(DB[1073]), .Z(n676) );
  AND U2471 ( .A(n226), .B(n677), .Z(n675) );
  XOR U2472 ( .A(n678), .B(n679), .Z(n677) );
  XOR U2473 ( .A(DB[1073]), .B(DB[1058]), .Z(n679) );
  AND U2474 ( .A(n230), .B(n680), .Z(n678) );
  XOR U2475 ( .A(n681), .B(n682), .Z(n680) );
  XOR U2476 ( .A(DB[1058]), .B(DB[1043]), .Z(n682) );
  AND U2477 ( .A(n234), .B(n683), .Z(n681) );
  XOR U2478 ( .A(n684), .B(n685), .Z(n683) );
  XOR U2479 ( .A(DB[1043]), .B(DB[1028]), .Z(n685) );
  AND U2480 ( .A(n238), .B(n686), .Z(n684) );
  XOR U2481 ( .A(n687), .B(n688), .Z(n686) );
  XOR U2482 ( .A(DB[1028]), .B(DB[1013]), .Z(n688) );
  AND U2483 ( .A(n242), .B(n689), .Z(n687) );
  XOR U2484 ( .A(n690), .B(n691), .Z(n689) );
  XOR U2485 ( .A(DB[998]), .B(DB[1013]), .Z(n691) );
  AND U2486 ( .A(n246), .B(n692), .Z(n690) );
  XOR U2487 ( .A(n693), .B(n694), .Z(n692) );
  XOR U2488 ( .A(DB[998]), .B(DB[983]), .Z(n694) );
  AND U2489 ( .A(n250), .B(n695), .Z(n693) );
  XOR U2490 ( .A(n696), .B(n697), .Z(n695) );
  XOR U2491 ( .A(DB[983]), .B(DB[968]), .Z(n697) );
  AND U2492 ( .A(n254), .B(n698), .Z(n696) );
  XOR U2493 ( .A(n699), .B(n700), .Z(n698) );
  XOR U2494 ( .A(DB[968]), .B(DB[953]), .Z(n700) );
  AND U2495 ( .A(n258), .B(n701), .Z(n699) );
  XOR U2496 ( .A(n702), .B(n703), .Z(n701) );
  XOR U2497 ( .A(DB[953]), .B(DB[938]), .Z(n703) );
  AND U2498 ( .A(n262), .B(n704), .Z(n702) );
  XOR U2499 ( .A(n705), .B(n706), .Z(n704) );
  XOR U2500 ( .A(DB[938]), .B(DB[923]), .Z(n706) );
  AND U2501 ( .A(n266), .B(n707), .Z(n705) );
  XOR U2502 ( .A(n708), .B(n709), .Z(n707) );
  XOR U2503 ( .A(DB[923]), .B(DB[908]), .Z(n709) );
  AND U2504 ( .A(n270), .B(n710), .Z(n708) );
  XOR U2505 ( .A(n711), .B(n712), .Z(n710) );
  XOR U2506 ( .A(DB[908]), .B(DB[893]), .Z(n712) );
  AND U2507 ( .A(n274), .B(n713), .Z(n711) );
  XOR U2508 ( .A(n714), .B(n715), .Z(n713) );
  XOR U2509 ( .A(DB[893]), .B(DB[878]), .Z(n715) );
  AND U2510 ( .A(n278), .B(n716), .Z(n714) );
  XOR U2511 ( .A(n717), .B(n718), .Z(n716) );
  XOR U2512 ( .A(DB[878]), .B(DB[863]), .Z(n718) );
  AND U2513 ( .A(n282), .B(n719), .Z(n717) );
  XOR U2514 ( .A(n720), .B(n721), .Z(n719) );
  XOR U2515 ( .A(DB[863]), .B(DB[848]), .Z(n721) );
  AND U2516 ( .A(n286), .B(n722), .Z(n720) );
  XOR U2517 ( .A(n723), .B(n724), .Z(n722) );
  XOR U2518 ( .A(DB[848]), .B(DB[833]), .Z(n724) );
  AND U2519 ( .A(n290), .B(n725), .Z(n723) );
  XOR U2520 ( .A(n726), .B(n727), .Z(n725) );
  XOR U2521 ( .A(DB[833]), .B(DB[818]), .Z(n727) );
  AND U2522 ( .A(n294), .B(n728), .Z(n726) );
  XOR U2523 ( .A(n729), .B(n730), .Z(n728) );
  XOR U2524 ( .A(DB[818]), .B(DB[803]), .Z(n730) );
  AND U2525 ( .A(n298), .B(n731), .Z(n729) );
  XOR U2526 ( .A(n732), .B(n733), .Z(n731) );
  XOR U2527 ( .A(DB[803]), .B(DB[788]), .Z(n733) );
  AND U2528 ( .A(n302), .B(n734), .Z(n732) );
  XOR U2529 ( .A(n735), .B(n736), .Z(n734) );
  XOR U2530 ( .A(DB[788]), .B(DB[773]), .Z(n736) );
  AND U2531 ( .A(n306), .B(n737), .Z(n735) );
  XOR U2532 ( .A(n738), .B(n739), .Z(n737) );
  XOR U2533 ( .A(DB[773]), .B(DB[758]), .Z(n739) );
  AND U2534 ( .A(n310), .B(n740), .Z(n738) );
  XOR U2535 ( .A(n741), .B(n742), .Z(n740) );
  XOR U2536 ( .A(DB[758]), .B(DB[743]), .Z(n742) );
  AND U2537 ( .A(n314), .B(n743), .Z(n741) );
  XOR U2538 ( .A(n744), .B(n745), .Z(n743) );
  XOR U2539 ( .A(DB[743]), .B(DB[728]), .Z(n745) );
  AND U2540 ( .A(n318), .B(n746), .Z(n744) );
  XOR U2541 ( .A(n747), .B(n748), .Z(n746) );
  XOR U2542 ( .A(DB[728]), .B(DB[713]), .Z(n748) );
  AND U2543 ( .A(n322), .B(n749), .Z(n747) );
  XOR U2544 ( .A(n750), .B(n751), .Z(n749) );
  XOR U2545 ( .A(DB[713]), .B(DB[698]), .Z(n751) );
  AND U2546 ( .A(n326), .B(n752), .Z(n750) );
  XOR U2547 ( .A(n753), .B(n754), .Z(n752) );
  XOR U2548 ( .A(DB[698]), .B(DB[683]), .Z(n754) );
  AND U2549 ( .A(n330), .B(n755), .Z(n753) );
  XOR U2550 ( .A(n756), .B(n757), .Z(n755) );
  XOR U2551 ( .A(DB[683]), .B(DB[668]), .Z(n757) );
  AND U2552 ( .A(n334), .B(n758), .Z(n756) );
  XOR U2553 ( .A(n759), .B(n760), .Z(n758) );
  XOR U2554 ( .A(DB[668]), .B(DB[653]), .Z(n760) );
  AND U2555 ( .A(n338), .B(n761), .Z(n759) );
  XOR U2556 ( .A(n762), .B(n763), .Z(n761) );
  XOR U2557 ( .A(DB[653]), .B(DB[638]), .Z(n763) );
  AND U2558 ( .A(n342), .B(n764), .Z(n762) );
  XOR U2559 ( .A(n765), .B(n766), .Z(n764) );
  XOR U2560 ( .A(DB[638]), .B(DB[623]), .Z(n766) );
  AND U2561 ( .A(n346), .B(n767), .Z(n765) );
  XOR U2562 ( .A(n768), .B(n769), .Z(n767) );
  XOR U2563 ( .A(DB[623]), .B(DB[608]), .Z(n769) );
  AND U2564 ( .A(n350), .B(n770), .Z(n768) );
  XOR U2565 ( .A(n771), .B(n772), .Z(n770) );
  XOR U2566 ( .A(DB[608]), .B(DB[593]), .Z(n772) );
  AND U2567 ( .A(n354), .B(n773), .Z(n771) );
  XOR U2568 ( .A(n774), .B(n775), .Z(n773) );
  XOR U2569 ( .A(DB[593]), .B(DB[578]), .Z(n775) );
  AND U2570 ( .A(n358), .B(n776), .Z(n774) );
  XOR U2571 ( .A(n777), .B(n778), .Z(n776) );
  XOR U2572 ( .A(DB[578]), .B(DB[563]), .Z(n778) );
  AND U2573 ( .A(n362), .B(n779), .Z(n777) );
  XOR U2574 ( .A(n780), .B(n781), .Z(n779) );
  XOR U2575 ( .A(DB[563]), .B(DB[548]), .Z(n781) );
  AND U2576 ( .A(n366), .B(n782), .Z(n780) );
  XOR U2577 ( .A(n783), .B(n784), .Z(n782) );
  XOR U2578 ( .A(DB[548]), .B(DB[533]), .Z(n784) );
  AND U2579 ( .A(n370), .B(n785), .Z(n783) );
  XOR U2580 ( .A(n786), .B(n787), .Z(n785) );
  XOR U2581 ( .A(DB[533]), .B(DB[518]), .Z(n787) );
  AND U2582 ( .A(n374), .B(n788), .Z(n786) );
  XOR U2583 ( .A(n789), .B(n790), .Z(n788) );
  XOR U2584 ( .A(DB[518]), .B(DB[503]), .Z(n790) );
  AND U2585 ( .A(n378), .B(n791), .Z(n789) );
  XOR U2586 ( .A(n792), .B(n793), .Z(n791) );
  XOR U2587 ( .A(DB[503]), .B(DB[488]), .Z(n793) );
  AND U2588 ( .A(n382), .B(n794), .Z(n792) );
  XOR U2589 ( .A(n795), .B(n796), .Z(n794) );
  XOR U2590 ( .A(DB[488]), .B(DB[473]), .Z(n796) );
  AND U2591 ( .A(n386), .B(n797), .Z(n795) );
  XOR U2592 ( .A(n798), .B(n799), .Z(n797) );
  XOR U2593 ( .A(DB[473]), .B(DB[458]), .Z(n799) );
  AND U2594 ( .A(n390), .B(n800), .Z(n798) );
  XOR U2595 ( .A(n801), .B(n802), .Z(n800) );
  XOR U2596 ( .A(DB[458]), .B(DB[443]), .Z(n802) );
  AND U2597 ( .A(n394), .B(n803), .Z(n801) );
  XOR U2598 ( .A(n804), .B(n805), .Z(n803) );
  XOR U2599 ( .A(DB[443]), .B(DB[428]), .Z(n805) );
  AND U2600 ( .A(n398), .B(n806), .Z(n804) );
  XOR U2601 ( .A(n807), .B(n808), .Z(n806) );
  XOR U2602 ( .A(DB[428]), .B(DB[413]), .Z(n808) );
  AND U2603 ( .A(n402), .B(n809), .Z(n807) );
  XOR U2604 ( .A(n810), .B(n811), .Z(n809) );
  XOR U2605 ( .A(DB[413]), .B(DB[398]), .Z(n811) );
  AND U2606 ( .A(n406), .B(n812), .Z(n810) );
  XOR U2607 ( .A(n813), .B(n814), .Z(n812) );
  XOR U2608 ( .A(DB[398]), .B(DB[383]), .Z(n814) );
  AND U2609 ( .A(n410), .B(n815), .Z(n813) );
  XOR U2610 ( .A(n816), .B(n817), .Z(n815) );
  XOR U2611 ( .A(DB[383]), .B(DB[368]), .Z(n817) );
  AND U2612 ( .A(n414), .B(n818), .Z(n816) );
  XOR U2613 ( .A(n819), .B(n820), .Z(n818) );
  XOR U2614 ( .A(DB[368]), .B(DB[353]), .Z(n820) );
  AND U2615 ( .A(n418), .B(n821), .Z(n819) );
  XOR U2616 ( .A(n822), .B(n823), .Z(n821) );
  XOR U2617 ( .A(DB[353]), .B(DB[338]), .Z(n823) );
  AND U2618 ( .A(n422), .B(n824), .Z(n822) );
  XOR U2619 ( .A(n825), .B(n826), .Z(n824) );
  XOR U2620 ( .A(DB[338]), .B(DB[323]), .Z(n826) );
  AND U2621 ( .A(n426), .B(n827), .Z(n825) );
  XOR U2622 ( .A(n828), .B(n829), .Z(n827) );
  XOR U2623 ( .A(DB[323]), .B(DB[308]), .Z(n829) );
  AND U2624 ( .A(n430), .B(n830), .Z(n828) );
  XOR U2625 ( .A(n831), .B(n832), .Z(n830) );
  XOR U2626 ( .A(DB[308]), .B(DB[293]), .Z(n832) );
  AND U2627 ( .A(n434), .B(n833), .Z(n831) );
  XOR U2628 ( .A(n834), .B(n835), .Z(n833) );
  XOR U2629 ( .A(DB[293]), .B(DB[278]), .Z(n835) );
  AND U2630 ( .A(n438), .B(n836), .Z(n834) );
  XOR U2631 ( .A(n837), .B(n838), .Z(n836) );
  XOR U2632 ( .A(DB[278]), .B(DB[263]), .Z(n838) );
  AND U2633 ( .A(n442), .B(n839), .Z(n837) );
  XOR U2634 ( .A(n840), .B(n841), .Z(n839) );
  XOR U2635 ( .A(DB[263]), .B(DB[248]), .Z(n841) );
  AND U2636 ( .A(n446), .B(n842), .Z(n840) );
  XOR U2637 ( .A(n843), .B(n844), .Z(n842) );
  XOR U2638 ( .A(DB[248]), .B(DB[233]), .Z(n844) );
  AND U2639 ( .A(n450), .B(n845), .Z(n843) );
  XOR U2640 ( .A(n846), .B(n847), .Z(n845) );
  XOR U2641 ( .A(DB[233]), .B(DB[218]), .Z(n847) );
  AND U2642 ( .A(n454), .B(n848), .Z(n846) );
  XOR U2643 ( .A(n849), .B(n850), .Z(n848) );
  XOR U2644 ( .A(DB[218]), .B(DB[203]), .Z(n850) );
  AND U2645 ( .A(n458), .B(n851), .Z(n849) );
  XOR U2646 ( .A(n852), .B(n853), .Z(n851) );
  XOR U2647 ( .A(DB[203]), .B(DB[188]), .Z(n853) );
  AND U2648 ( .A(n462), .B(n854), .Z(n852) );
  XOR U2649 ( .A(n855), .B(n856), .Z(n854) );
  XOR U2650 ( .A(DB[188]), .B(DB[173]), .Z(n856) );
  AND U2651 ( .A(n466), .B(n857), .Z(n855) );
  XOR U2652 ( .A(n858), .B(n859), .Z(n857) );
  XOR U2653 ( .A(DB[173]), .B(DB[158]), .Z(n859) );
  AND U2654 ( .A(n470), .B(n860), .Z(n858) );
  XOR U2655 ( .A(n861), .B(n862), .Z(n860) );
  XOR U2656 ( .A(DB[158]), .B(DB[143]), .Z(n862) );
  AND U2657 ( .A(n474), .B(n863), .Z(n861) );
  XOR U2658 ( .A(n864), .B(n865), .Z(n863) );
  XOR U2659 ( .A(DB[143]), .B(DB[128]), .Z(n865) );
  AND U2660 ( .A(n478), .B(n866), .Z(n864) );
  XOR U2661 ( .A(n867), .B(n868), .Z(n866) );
  XOR U2662 ( .A(DB[128]), .B(DB[113]), .Z(n868) );
  AND U2663 ( .A(n482), .B(n869), .Z(n867) );
  XOR U2664 ( .A(n870), .B(n871), .Z(n869) );
  XOR U2665 ( .A(DB[98]), .B(DB[113]), .Z(n871) );
  AND U2666 ( .A(n486), .B(n872), .Z(n870) );
  XOR U2667 ( .A(n873), .B(n874), .Z(n872) );
  XOR U2668 ( .A(DB[98]), .B(DB[83]), .Z(n874) );
  AND U2669 ( .A(n490), .B(n875), .Z(n873) );
  XOR U2670 ( .A(n876), .B(n877), .Z(n875) );
  XOR U2671 ( .A(DB[83]), .B(DB[68]), .Z(n877) );
  AND U2672 ( .A(n494), .B(n878), .Z(n876) );
  XOR U2673 ( .A(n879), .B(n880), .Z(n878) );
  XOR U2674 ( .A(DB[68]), .B(DB[53]), .Z(n880) );
  AND U2675 ( .A(n498), .B(n881), .Z(n879) );
  XOR U2676 ( .A(n882), .B(n883), .Z(n881) );
  XOR U2677 ( .A(DB[53]), .B(DB[38]), .Z(n883) );
  AND U2678 ( .A(n502), .B(n884), .Z(n882) );
  XOR U2679 ( .A(n885), .B(n886), .Z(n884) );
  XOR U2680 ( .A(DB[38]), .B(DB[23]), .Z(n886) );
  AND U2681 ( .A(n506), .B(n887), .Z(n885) );
  XOR U2682 ( .A(DB[8]), .B(DB[23]), .Z(n887) );
  XOR U2683 ( .A(DB[1912]), .B(n888), .Z(min_val_out[7]) );
  AND U2684 ( .A(n2), .B(n889), .Z(n888) );
  XOR U2685 ( .A(n890), .B(n891), .Z(n889) );
  XOR U2686 ( .A(DB[1912]), .B(DB[1897]), .Z(n891) );
  AND U2687 ( .A(n6), .B(n892), .Z(n890) );
  XOR U2688 ( .A(n893), .B(n894), .Z(n892) );
  XOR U2689 ( .A(DB[1897]), .B(DB[1882]), .Z(n894) );
  AND U2690 ( .A(n10), .B(n895), .Z(n893) );
  XOR U2691 ( .A(n896), .B(n897), .Z(n895) );
  XOR U2692 ( .A(DB[1882]), .B(DB[1867]), .Z(n897) );
  AND U2693 ( .A(n14), .B(n898), .Z(n896) );
  XOR U2694 ( .A(n899), .B(n900), .Z(n898) );
  XOR U2695 ( .A(DB[1867]), .B(DB[1852]), .Z(n900) );
  AND U2696 ( .A(n18), .B(n901), .Z(n899) );
  XOR U2697 ( .A(n902), .B(n903), .Z(n901) );
  XOR U2698 ( .A(DB[1852]), .B(DB[1837]), .Z(n903) );
  AND U2699 ( .A(n22), .B(n904), .Z(n902) );
  XOR U2700 ( .A(n905), .B(n906), .Z(n904) );
  XOR U2701 ( .A(DB[1837]), .B(DB[1822]), .Z(n906) );
  AND U2702 ( .A(n26), .B(n907), .Z(n905) );
  XOR U2703 ( .A(n908), .B(n909), .Z(n907) );
  XOR U2704 ( .A(DB[1822]), .B(DB[1807]), .Z(n909) );
  AND U2705 ( .A(n30), .B(n910), .Z(n908) );
  XOR U2706 ( .A(n911), .B(n912), .Z(n910) );
  XOR U2707 ( .A(DB[1807]), .B(DB[1792]), .Z(n912) );
  AND U2708 ( .A(n34), .B(n913), .Z(n911) );
  XOR U2709 ( .A(n914), .B(n915), .Z(n913) );
  XOR U2710 ( .A(DB[1792]), .B(DB[1777]), .Z(n915) );
  AND U2711 ( .A(n38), .B(n916), .Z(n914) );
  XOR U2712 ( .A(n917), .B(n918), .Z(n916) );
  XOR U2713 ( .A(DB[1777]), .B(DB[1762]), .Z(n918) );
  AND U2714 ( .A(n42), .B(n919), .Z(n917) );
  XOR U2715 ( .A(n920), .B(n921), .Z(n919) );
  XOR U2716 ( .A(DB[1762]), .B(DB[1747]), .Z(n921) );
  AND U2717 ( .A(n46), .B(n922), .Z(n920) );
  XOR U2718 ( .A(n923), .B(n924), .Z(n922) );
  XOR U2719 ( .A(DB[1747]), .B(DB[1732]), .Z(n924) );
  AND U2720 ( .A(n50), .B(n925), .Z(n923) );
  XOR U2721 ( .A(n926), .B(n927), .Z(n925) );
  XOR U2722 ( .A(DB[1732]), .B(DB[1717]), .Z(n927) );
  AND U2723 ( .A(n54), .B(n928), .Z(n926) );
  XOR U2724 ( .A(n929), .B(n930), .Z(n928) );
  XOR U2725 ( .A(DB[1717]), .B(DB[1702]), .Z(n930) );
  AND U2726 ( .A(n58), .B(n931), .Z(n929) );
  XOR U2727 ( .A(n932), .B(n933), .Z(n931) );
  XOR U2728 ( .A(DB[1702]), .B(DB[1687]), .Z(n933) );
  AND U2729 ( .A(n62), .B(n934), .Z(n932) );
  XOR U2730 ( .A(n935), .B(n936), .Z(n934) );
  XOR U2731 ( .A(DB[1687]), .B(DB[1672]), .Z(n936) );
  AND U2732 ( .A(n66), .B(n937), .Z(n935) );
  XOR U2733 ( .A(n938), .B(n939), .Z(n937) );
  XOR U2734 ( .A(DB[1672]), .B(DB[1657]), .Z(n939) );
  AND U2735 ( .A(n70), .B(n940), .Z(n938) );
  XOR U2736 ( .A(n941), .B(n942), .Z(n940) );
  XOR U2737 ( .A(DB[1657]), .B(DB[1642]), .Z(n942) );
  AND U2738 ( .A(n74), .B(n943), .Z(n941) );
  XOR U2739 ( .A(n944), .B(n945), .Z(n943) );
  XOR U2740 ( .A(DB[1642]), .B(DB[1627]), .Z(n945) );
  AND U2741 ( .A(n78), .B(n946), .Z(n944) );
  XOR U2742 ( .A(n947), .B(n948), .Z(n946) );
  XOR U2743 ( .A(DB[1627]), .B(DB[1612]), .Z(n948) );
  AND U2744 ( .A(n82), .B(n949), .Z(n947) );
  XOR U2745 ( .A(n950), .B(n951), .Z(n949) );
  XOR U2746 ( .A(DB[1612]), .B(DB[1597]), .Z(n951) );
  AND U2747 ( .A(n86), .B(n952), .Z(n950) );
  XOR U2748 ( .A(n953), .B(n954), .Z(n952) );
  XOR U2749 ( .A(DB[1597]), .B(DB[1582]), .Z(n954) );
  AND U2750 ( .A(n90), .B(n955), .Z(n953) );
  XOR U2751 ( .A(n956), .B(n957), .Z(n955) );
  XOR U2752 ( .A(DB[1582]), .B(DB[1567]), .Z(n957) );
  AND U2753 ( .A(n94), .B(n958), .Z(n956) );
  XOR U2754 ( .A(n959), .B(n960), .Z(n958) );
  XOR U2755 ( .A(DB[1567]), .B(DB[1552]), .Z(n960) );
  AND U2756 ( .A(n98), .B(n961), .Z(n959) );
  XOR U2757 ( .A(n962), .B(n963), .Z(n961) );
  XOR U2758 ( .A(DB[1552]), .B(DB[1537]), .Z(n963) );
  AND U2759 ( .A(n102), .B(n964), .Z(n962) );
  XOR U2760 ( .A(n965), .B(n966), .Z(n964) );
  XOR U2761 ( .A(DB[1537]), .B(DB[1522]), .Z(n966) );
  AND U2762 ( .A(n106), .B(n967), .Z(n965) );
  XOR U2763 ( .A(n968), .B(n969), .Z(n967) );
  XOR U2764 ( .A(DB[1522]), .B(DB[1507]), .Z(n969) );
  AND U2765 ( .A(n110), .B(n970), .Z(n968) );
  XOR U2766 ( .A(n971), .B(n972), .Z(n970) );
  XOR U2767 ( .A(DB[1507]), .B(DB[1492]), .Z(n972) );
  AND U2768 ( .A(n114), .B(n973), .Z(n971) );
  XOR U2769 ( .A(n974), .B(n975), .Z(n973) );
  XOR U2770 ( .A(DB[1492]), .B(DB[1477]), .Z(n975) );
  AND U2771 ( .A(n118), .B(n976), .Z(n974) );
  XOR U2772 ( .A(n977), .B(n978), .Z(n976) );
  XOR U2773 ( .A(DB[1477]), .B(DB[1462]), .Z(n978) );
  AND U2774 ( .A(n122), .B(n979), .Z(n977) );
  XOR U2775 ( .A(n980), .B(n981), .Z(n979) );
  XOR U2776 ( .A(DB[1462]), .B(DB[1447]), .Z(n981) );
  AND U2777 ( .A(n126), .B(n982), .Z(n980) );
  XOR U2778 ( .A(n983), .B(n984), .Z(n982) );
  XOR U2779 ( .A(DB[1447]), .B(DB[1432]), .Z(n984) );
  AND U2780 ( .A(n130), .B(n985), .Z(n983) );
  XOR U2781 ( .A(n986), .B(n987), .Z(n985) );
  XOR U2782 ( .A(DB[1432]), .B(DB[1417]), .Z(n987) );
  AND U2783 ( .A(n134), .B(n988), .Z(n986) );
  XOR U2784 ( .A(n989), .B(n990), .Z(n988) );
  XOR U2785 ( .A(DB[1417]), .B(DB[1402]), .Z(n990) );
  AND U2786 ( .A(n138), .B(n991), .Z(n989) );
  XOR U2787 ( .A(n992), .B(n993), .Z(n991) );
  XOR U2788 ( .A(DB[1402]), .B(DB[1387]), .Z(n993) );
  AND U2789 ( .A(n142), .B(n994), .Z(n992) );
  XOR U2790 ( .A(n995), .B(n996), .Z(n994) );
  XOR U2791 ( .A(DB[1387]), .B(DB[1372]), .Z(n996) );
  AND U2792 ( .A(n146), .B(n997), .Z(n995) );
  XOR U2793 ( .A(n998), .B(n999), .Z(n997) );
  XOR U2794 ( .A(DB[1372]), .B(DB[1357]), .Z(n999) );
  AND U2795 ( .A(n150), .B(n1000), .Z(n998) );
  XOR U2796 ( .A(n1001), .B(n1002), .Z(n1000) );
  XOR U2797 ( .A(DB[1357]), .B(DB[1342]), .Z(n1002) );
  AND U2798 ( .A(n154), .B(n1003), .Z(n1001) );
  XOR U2799 ( .A(n1004), .B(n1005), .Z(n1003) );
  XOR U2800 ( .A(DB[1342]), .B(DB[1327]), .Z(n1005) );
  AND U2801 ( .A(n158), .B(n1006), .Z(n1004) );
  XOR U2802 ( .A(n1007), .B(n1008), .Z(n1006) );
  XOR U2803 ( .A(DB[1327]), .B(DB[1312]), .Z(n1008) );
  AND U2804 ( .A(n162), .B(n1009), .Z(n1007) );
  XOR U2805 ( .A(n1010), .B(n1011), .Z(n1009) );
  XOR U2806 ( .A(DB[1312]), .B(DB[1297]), .Z(n1011) );
  AND U2807 ( .A(n166), .B(n1012), .Z(n1010) );
  XOR U2808 ( .A(n1013), .B(n1014), .Z(n1012) );
  XOR U2809 ( .A(DB[1297]), .B(DB[1282]), .Z(n1014) );
  AND U2810 ( .A(n170), .B(n1015), .Z(n1013) );
  XOR U2811 ( .A(n1016), .B(n1017), .Z(n1015) );
  XOR U2812 ( .A(DB[1282]), .B(DB[1267]), .Z(n1017) );
  AND U2813 ( .A(n174), .B(n1018), .Z(n1016) );
  XOR U2814 ( .A(n1019), .B(n1020), .Z(n1018) );
  XOR U2815 ( .A(DB[1267]), .B(DB[1252]), .Z(n1020) );
  AND U2816 ( .A(n178), .B(n1021), .Z(n1019) );
  XOR U2817 ( .A(n1022), .B(n1023), .Z(n1021) );
  XOR U2818 ( .A(DB[1252]), .B(DB[1237]), .Z(n1023) );
  AND U2819 ( .A(n182), .B(n1024), .Z(n1022) );
  XOR U2820 ( .A(n1025), .B(n1026), .Z(n1024) );
  XOR U2821 ( .A(DB[1237]), .B(DB[1222]), .Z(n1026) );
  AND U2822 ( .A(n186), .B(n1027), .Z(n1025) );
  XOR U2823 ( .A(n1028), .B(n1029), .Z(n1027) );
  XOR U2824 ( .A(DB[1222]), .B(DB[1207]), .Z(n1029) );
  AND U2825 ( .A(n190), .B(n1030), .Z(n1028) );
  XOR U2826 ( .A(n1031), .B(n1032), .Z(n1030) );
  XOR U2827 ( .A(DB[1207]), .B(DB[1192]), .Z(n1032) );
  AND U2828 ( .A(n194), .B(n1033), .Z(n1031) );
  XOR U2829 ( .A(n1034), .B(n1035), .Z(n1033) );
  XOR U2830 ( .A(DB[1192]), .B(DB[1177]), .Z(n1035) );
  AND U2831 ( .A(n198), .B(n1036), .Z(n1034) );
  XOR U2832 ( .A(n1037), .B(n1038), .Z(n1036) );
  XOR U2833 ( .A(DB[1177]), .B(DB[1162]), .Z(n1038) );
  AND U2834 ( .A(n202), .B(n1039), .Z(n1037) );
  XOR U2835 ( .A(n1040), .B(n1041), .Z(n1039) );
  XOR U2836 ( .A(DB[1162]), .B(DB[1147]), .Z(n1041) );
  AND U2837 ( .A(n206), .B(n1042), .Z(n1040) );
  XOR U2838 ( .A(n1043), .B(n1044), .Z(n1042) );
  XOR U2839 ( .A(DB[1147]), .B(DB[1132]), .Z(n1044) );
  AND U2840 ( .A(n210), .B(n1045), .Z(n1043) );
  XOR U2841 ( .A(n1046), .B(n1047), .Z(n1045) );
  XOR U2842 ( .A(DB[1132]), .B(DB[1117]), .Z(n1047) );
  AND U2843 ( .A(n214), .B(n1048), .Z(n1046) );
  XOR U2844 ( .A(n1049), .B(n1050), .Z(n1048) );
  XOR U2845 ( .A(DB[1117]), .B(DB[1102]), .Z(n1050) );
  AND U2846 ( .A(n218), .B(n1051), .Z(n1049) );
  XOR U2847 ( .A(n1052), .B(n1053), .Z(n1051) );
  XOR U2848 ( .A(DB[1102]), .B(DB[1087]), .Z(n1053) );
  AND U2849 ( .A(n222), .B(n1054), .Z(n1052) );
  XOR U2850 ( .A(n1055), .B(n1056), .Z(n1054) );
  XOR U2851 ( .A(DB[1087]), .B(DB[1072]), .Z(n1056) );
  AND U2852 ( .A(n226), .B(n1057), .Z(n1055) );
  XOR U2853 ( .A(n1058), .B(n1059), .Z(n1057) );
  XOR U2854 ( .A(DB[1072]), .B(DB[1057]), .Z(n1059) );
  AND U2855 ( .A(n230), .B(n1060), .Z(n1058) );
  XOR U2856 ( .A(n1061), .B(n1062), .Z(n1060) );
  XOR U2857 ( .A(DB[1057]), .B(DB[1042]), .Z(n1062) );
  AND U2858 ( .A(n234), .B(n1063), .Z(n1061) );
  XOR U2859 ( .A(n1064), .B(n1065), .Z(n1063) );
  XOR U2860 ( .A(DB[1042]), .B(DB[1027]), .Z(n1065) );
  AND U2861 ( .A(n238), .B(n1066), .Z(n1064) );
  XOR U2862 ( .A(n1067), .B(n1068), .Z(n1066) );
  XOR U2863 ( .A(DB[1027]), .B(DB[1012]), .Z(n1068) );
  AND U2864 ( .A(n242), .B(n1069), .Z(n1067) );
  XOR U2865 ( .A(n1070), .B(n1071), .Z(n1069) );
  XOR U2866 ( .A(DB[997]), .B(DB[1012]), .Z(n1071) );
  AND U2867 ( .A(n246), .B(n1072), .Z(n1070) );
  XOR U2868 ( .A(n1073), .B(n1074), .Z(n1072) );
  XOR U2869 ( .A(DB[997]), .B(DB[982]), .Z(n1074) );
  AND U2870 ( .A(n250), .B(n1075), .Z(n1073) );
  XOR U2871 ( .A(n1076), .B(n1077), .Z(n1075) );
  XOR U2872 ( .A(DB[982]), .B(DB[967]), .Z(n1077) );
  AND U2873 ( .A(n254), .B(n1078), .Z(n1076) );
  XOR U2874 ( .A(n1079), .B(n1080), .Z(n1078) );
  XOR U2875 ( .A(DB[967]), .B(DB[952]), .Z(n1080) );
  AND U2876 ( .A(n258), .B(n1081), .Z(n1079) );
  XOR U2877 ( .A(n1082), .B(n1083), .Z(n1081) );
  XOR U2878 ( .A(DB[952]), .B(DB[937]), .Z(n1083) );
  AND U2879 ( .A(n262), .B(n1084), .Z(n1082) );
  XOR U2880 ( .A(n1085), .B(n1086), .Z(n1084) );
  XOR U2881 ( .A(DB[937]), .B(DB[922]), .Z(n1086) );
  AND U2882 ( .A(n266), .B(n1087), .Z(n1085) );
  XOR U2883 ( .A(n1088), .B(n1089), .Z(n1087) );
  XOR U2884 ( .A(DB[922]), .B(DB[907]), .Z(n1089) );
  AND U2885 ( .A(n270), .B(n1090), .Z(n1088) );
  XOR U2886 ( .A(n1091), .B(n1092), .Z(n1090) );
  XOR U2887 ( .A(DB[907]), .B(DB[892]), .Z(n1092) );
  AND U2888 ( .A(n274), .B(n1093), .Z(n1091) );
  XOR U2889 ( .A(n1094), .B(n1095), .Z(n1093) );
  XOR U2890 ( .A(DB[892]), .B(DB[877]), .Z(n1095) );
  AND U2891 ( .A(n278), .B(n1096), .Z(n1094) );
  XOR U2892 ( .A(n1097), .B(n1098), .Z(n1096) );
  XOR U2893 ( .A(DB[877]), .B(DB[862]), .Z(n1098) );
  AND U2894 ( .A(n282), .B(n1099), .Z(n1097) );
  XOR U2895 ( .A(n1100), .B(n1101), .Z(n1099) );
  XOR U2896 ( .A(DB[862]), .B(DB[847]), .Z(n1101) );
  AND U2897 ( .A(n286), .B(n1102), .Z(n1100) );
  XOR U2898 ( .A(n1103), .B(n1104), .Z(n1102) );
  XOR U2899 ( .A(DB[847]), .B(DB[832]), .Z(n1104) );
  AND U2900 ( .A(n290), .B(n1105), .Z(n1103) );
  XOR U2901 ( .A(n1106), .B(n1107), .Z(n1105) );
  XOR U2902 ( .A(DB[832]), .B(DB[817]), .Z(n1107) );
  AND U2903 ( .A(n294), .B(n1108), .Z(n1106) );
  XOR U2904 ( .A(n1109), .B(n1110), .Z(n1108) );
  XOR U2905 ( .A(DB[817]), .B(DB[802]), .Z(n1110) );
  AND U2906 ( .A(n298), .B(n1111), .Z(n1109) );
  XOR U2907 ( .A(n1112), .B(n1113), .Z(n1111) );
  XOR U2908 ( .A(DB[802]), .B(DB[787]), .Z(n1113) );
  AND U2909 ( .A(n302), .B(n1114), .Z(n1112) );
  XOR U2910 ( .A(n1115), .B(n1116), .Z(n1114) );
  XOR U2911 ( .A(DB[787]), .B(DB[772]), .Z(n1116) );
  AND U2912 ( .A(n306), .B(n1117), .Z(n1115) );
  XOR U2913 ( .A(n1118), .B(n1119), .Z(n1117) );
  XOR U2914 ( .A(DB[772]), .B(DB[757]), .Z(n1119) );
  AND U2915 ( .A(n310), .B(n1120), .Z(n1118) );
  XOR U2916 ( .A(n1121), .B(n1122), .Z(n1120) );
  XOR U2917 ( .A(DB[757]), .B(DB[742]), .Z(n1122) );
  AND U2918 ( .A(n314), .B(n1123), .Z(n1121) );
  XOR U2919 ( .A(n1124), .B(n1125), .Z(n1123) );
  XOR U2920 ( .A(DB[742]), .B(DB[727]), .Z(n1125) );
  AND U2921 ( .A(n318), .B(n1126), .Z(n1124) );
  XOR U2922 ( .A(n1127), .B(n1128), .Z(n1126) );
  XOR U2923 ( .A(DB[727]), .B(DB[712]), .Z(n1128) );
  AND U2924 ( .A(n322), .B(n1129), .Z(n1127) );
  XOR U2925 ( .A(n1130), .B(n1131), .Z(n1129) );
  XOR U2926 ( .A(DB[712]), .B(DB[697]), .Z(n1131) );
  AND U2927 ( .A(n326), .B(n1132), .Z(n1130) );
  XOR U2928 ( .A(n1133), .B(n1134), .Z(n1132) );
  XOR U2929 ( .A(DB[697]), .B(DB[682]), .Z(n1134) );
  AND U2930 ( .A(n330), .B(n1135), .Z(n1133) );
  XOR U2931 ( .A(n1136), .B(n1137), .Z(n1135) );
  XOR U2932 ( .A(DB[682]), .B(DB[667]), .Z(n1137) );
  AND U2933 ( .A(n334), .B(n1138), .Z(n1136) );
  XOR U2934 ( .A(n1139), .B(n1140), .Z(n1138) );
  XOR U2935 ( .A(DB[667]), .B(DB[652]), .Z(n1140) );
  AND U2936 ( .A(n338), .B(n1141), .Z(n1139) );
  XOR U2937 ( .A(n1142), .B(n1143), .Z(n1141) );
  XOR U2938 ( .A(DB[652]), .B(DB[637]), .Z(n1143) );
  AND U2939 ( .A(n342), .B(n1144), .Z(n1142) );
  XOR U2940 ( .A(n1145), .B(n1146), .Z(n1144) );
  XOR U2941 ( .A(DB[637]), .B(DB[622]), .Z(n1146) );
  AND U2942 ( .A(n346), .B(n1147), .Z(n1145) );
  XOR U2943 ( .A(n1148), .B(n1149), .Z(n1147) );
  XOR U2944 ( .A(DB[622]), .B(DB[607]), .Z(n1149) );
  AND U2945 ( .A(n350), .B(n1150), .Z(n1148) );
  XOR U2946 ( .A(n1151), .B(n1152), .Z(n1150) );
  XOR U2947 ( .A(DB[607]), .B(DB[592]), .Z(n1152) );
  AND U2948 ( .A(n354), .B(n1153), .Z(n1151) );
  XOR U2949 ( .A(n1154), .B(n1155), .Z(n1153) );
  XOR U2950 ( .A(DB[592]), .B(DB[577]), .Z(n1155) );
  AND U2951 ( .A(n358), .B(n1156), .Z(n1154) );
  XOR U2952 ( .A(n1157), .B(n1158), .Z(n1156) );
  XOR U2953 ( .A(DB[577]), .B(DB[562]), .Z(n1158) );
  AND U2954 ( .A(n362), .B(n1159), .Z(n1157) );
  XOR U2955 ( .A(n1160), .B(n1161), .Z(n1159) );
  XOR U2956 ( .A(DB[562]), .B(DB[547]), .Z(n1161) );
  AND U2957 ( .A(n366), .B(n1162), .Z(n1160) );
  XOR U2958 ( .A(n1163), .B(n1164), .Z(n1162) );
  XOR U2959 ( .A(DB[547]), .B(DB[532]), .Z(n1164) );
  AND U2960 ( .A(n370), .B(n1165), .Z(n1163) );
  XOR U2961 ( .A(n1166), .B(n1167), .Z(n1165) );
  XOR U2962 ( .A(DB[532]), .B(DB[517]), .Z(n1167) );
  AND U2963 ( .A(n374), .B(n1168), .Z(n1166) );
  XOR U2964 ( .A(n1169), .B(n1170), .Z(n1168) );
  XOR U2965 ( .A(DB[517]), .B(DB[502]), .Z(n1170) );
  AND U2966 ( .A(n378), .B(n1171), .Z(n1169) );
  XOR U2967 ( .A(n1172), .B(n1173), .Z(n1171) );
  XOR U2968 ( .A(DB[502]), .B(DB[487]), .Z(n1173) );
  AND U2969 ( .A(n382), .B(n1174), .Z(n1172) );
  XOR U2970 ( .A(n1175), .B(n1176), .Z(n1174) );
  XOR U2971 ( .A(DB[487]), .B(DB[472]), .Z(n1176) );
  AND U2972 ( .A(n386), .B(n1177), .Z(n1175) );
  XOR U2973 ( .A(n1178), .B(n1179), .Z(n1177) );
  XOR U2974 ( .A(DB[472]), .B(DB[457]), .Z(n1179) );
  AND U2975 ( .A(n390), .B(n1180), .Z(n1178) );
  XOR U2976 ( .A(n1181), .B(n1182), .Z(n1180) );
  XOR U2977 ( .A(DB[457]), .B(DB[442]), .Z(n1182) );
  AND U2978 ( .A(n394), .B(n1183), .Z(n1181) );
  XOR U2979 ( .A(n1184), .B(n1185), .Z(n1183) );
  XOR U2980 ( .A(DB[442]), .B(DB[427]), .Z(n1185) );
  AND U2981 ( .A(n398), .B(n1186), .Z(n1184) );
  XOR U2982 ( .A(n1187), .B(n1188), .Z(n1186) );
  XOR U2983 ( .A(DB[427]), .B(DB[412]), .Z(n1188) );
  AND U2984 ( .A(n402), .B(n1189), .Z(n1187) );
  XOR U2985 ( .A(n1190), .B(n1191), .Z(n1189) );
  XOR U2986 ( .A(DB[412]), .B(DB[397]), .Z(n1191) );
  AND U2987 ( .A(n406), .B(n1192), .Z(n1190) );
  XOR U2988 ( .A(n1193), .B(n1194), .Z(n1192) );
  XOR U2989 ( .A(DB[397]), .B(DB[382]), .Z(n1194) );
  AND U2990 ( .A(n410), .B(n1195), .Z(n1193) );
  XOR U2991 ( .A(n1196), .B(n1197), .Z(n1195) );
  XOR U2992 ( .A(DB[382]), .B(DB[367]), .Z(n1197) );
  AND U2993 ( .A(n414), .B(n1198), .Z(n1196) );
  XOR U2994 ( .A(n1199), .B(n1200), .Z(n1198) );
  XOR U2995 ( .A(DB[367]), .B(DB[352]), .Z(n1200) );
  AND U2996 ( .A(n418), .B(n1201), .Z(n1199) );
  XOR U2997 ( .A(n1202), .B(n1203), .Z(n1201) );
  XOR U2998 ( .A(DB[352]), .B(DB[337]), .Z(n1203) );
  AND U2999 ( .A(n422), .B(n1204), .Z(n1202) );
  XOR U3000 ( .A(n1205), .B(n1206), .Z(n1204) );
  XOR U3001 ( .A(DB[337]), .B(DB[322]), .Z(n1206) );
  AND U3002 ( .A(n426), .B(n1207), .Z(n1205) );
  XOR U3003 ( .A(n1208), .B(n1209), .Z(n1207) );
  XOR U3004 ( .A(DB[322]), .B(DB[307]), .Z(n1209) );
  AND U3005 ( .A(n430), .B(n1210), .Z(n1208) );
  XOR U3006 ( .A(n1211), .B(n1212), .Z(n1210) );
  XOR U3007 ( .A(DB[307]), .B(DB[292]), .Z(n1212) );
  AND U3008 ( .A(n434), .B(n1213), .Z(n1211) );
  XOR U3009 ( .A(n1214), .B(n1215), .Z(n1213) );
  XOR U3010 ( .A(DB[292]), .B(DB[277]), .Z(n1215) );
  AND U3011 ( .A(n438), .B(n1216), .Z(n1214) );
  XOR U3012 ( .A(n1217), .B(n1218), .Z(n1216) );
  XOR U3013 ( .A(DB[277]), .B(DB[262]), .Z(n1218) );
  AND U3014 ( .A(n442), .B(n1219), .Z(n1217) );
  XOR U3015 ( .A(n1220), .B(n1221), .Z(n1219) );
  XOR U3016 ( .A(DB[262]), .B(DB[247]), .Z(n1221) );
  AND U3017 ( .A(n446), .B(n1222), .Z(n1220) );
  XOR U3018 ( .A(n1223), .B(n1224), .Z(n1222) );
  XOR U3019 ( .A(DB[247]), .B(DB[232]), .Z(n1224) );
  AND U3020 ( .A(n450), .B(n1225), .Z(n1223) );
  XOR U3021 ( .A(n1226), .B(n1227), .Z(n1225) );
  XOR U3022 ( .A(DB[232]), .B(DB[217]), .Z(n1227) );
  AND U3023 ( .A(n454), .B(n1228), .Z(n1226) );
  XOR U3024 ( .A(n1229), .B(n1230), .Z(n1228) );
  XOR U3025 ( .A(DB[217]), .B(DB[202]), .Z(n1230) );
  AND U3026 ( .A(n458), .B(n1231), .Z(n1229) );
  XOR U3027 ( .A(n1232), .B(n1233), .Z(n1231) );
  XOR U3028 ( .A(DB[202]), .B(DB[187]), .Z(n1233) );
  AND U3029 ( .A(n462), .B(n1234), .Z(n1232) );
  XOR U3030 ( .A(n1235), .B(n1236), .Z(n1234) );
  XOR U3031 ( .A(DB[187]), .B(DB[172]), .Z(n1236) );
  AND U3032 ( .A(n466), .B(n1237), .Z(n1235) );
  XOR U3033 ( .A(n1238), .B(n1239), .Z(n1237) );
  XOR U3034 ( .A(DB[172]), .B(DB[157]), .Z(n1239) );
  AND U3035 ( .A(n470), .B(n1240), .Z(n1238) );
  XOR U3036 ( .A(n1241), .B(n1242), .Z(n1240) );
  XOR U3037 ( .A(DB[157]), .B(DB[142]), .Z(n1242) );
  AND U3038 ( .A(n474), .B(n1243), .Z(n1241) );
  XOR U3039 ( .A(n1244), .B(n1245), .Z(n1243) );
  XOR U3040 ( .A(DB[142]), .B(DB[127]), .Z(n1245) );
  AND U3041 ( .A(n478), .B(n1246), .Z(n1244) );
  XOR U3042 ( .A(n1247), .B(n1248), .Z(n1246) );
  XOR U3043 ( .A(DB[127]), .B(DB[112]), .Z(n1248) );
  AND U3044 ( .A(n482), .B(n1249), .Z(n1247) );
  XOR U3045 ( .A(n1250), .B(n1251), .Z(n1249) );
  XOR U3046 ( .A(DB[97]), .B(DB[112]), .Z(n1251) );
  AND U3047 ( .A(n486), .B(n1252), .Z(n1250) );
  XOR U3048 ( .A(n1253), .B(n1254), .Z(n1252) );
  XOR U3049 ( .A(DB[97]), .B(DB[82]), .Z(n1254) );
  AND U3050 ( .A(n490), .B(n1255), .Z(n1253) );
  XOR U3051 ( .A(n1256), .B(n1257), .Z(n1255) );
  XOR U3052 ( .A(DB[82]), .B(DB[67]), .Z(n1257) );
  AND U3053 ( .A(n494), .B(n1258), .Z(n1256) );
  XOR U3054 ( .A(n1259), .B(n1260), .Z(n1258) );
  XOR U3055 ( .A(DB[67]), .B(DB[52]), .Z(n1260) );
  AND U3056 ( .A(n498), .B(n1261), .Z(n1259) );
  XOR U3057 ( .A(n1262), .B(n1263), .Z(n1261) );
  XOR U3058 ( .A(DB[52]), .B(DB[37]), .Z(n1263) );
  AND U3059 ( .A(n502), .B(n1264), .Z(n1262) );
  XOR U3060 ( .A(n1265), .B(n1266), .Z(n1264) );
  XOR U3061 ( .A(DB[37]), .B(DB[22]), .Z(n1266) );
  AND U3062 ( .A(n506), .B(n1267), .Z(n1265) );
  XOR U3063 ( .A(DB[7]), .B(DB[22]), .Z(n1267) );
  XOR U3064 ( .A(DB[1911]), .B(n1268), .Z(min_val_out[6]) );
  AND U3065 ( .A(n2), .B(n1269), .Z(n1268) );
  XOR U3066 ( .A(n1270), .B(n1271), .Z(n1269) );
  XOR U3067 ( .A(DB[1911]), .B(DB[1896]), .Z(n1271) );
  AND U3068 ( .A(n6), .B(n1272), .Z(n1270) );
  XOR U3069 ( .A(n1273), .B(n1274), .Z(n1272) );
  XOR U3070 ( .A(DB[1896]), .B(DB[1881]), .Z(n1274) );
  AND U3071 ( .A(n10), .B(n1275), .Z(n1273) );
  XOR U3072 ( .A(n1276), .B(n1277), .Z(n1275) );
  XOR U3073 ( .A(DB[1881]), .B(DB[1866]), .Z(n1277) );
  AND U3074 ( .A(n14), .B(n1278), .Z(n1276) );
  XOR U3075 ( .A(n1279), .B(n1280), .Z(n1278) );
  XOR U3076 ( .A(DB[1866]), .B(DB[1851]), .Z(n1280) );
  AND U3077 ( .A(n18), .B(n1281), .Z(n1279) );
  XOR U3078 ( .A(n1282), .B(n1283), .Z(n1281) );
  XOR U3079 ( .A(DB[1851]), .B(DB[1836]), .Z(n1283) );
  AND U3080 ( .A(n22), .B(n1284), .Z(n1282) );
  XOR U3081 ( .A(n1285), .B(n1286), .Z(n1284) );
  XOR U3082 ( .A(DB[1836]), .B(DB[1821]), .Z(n1286) );
  AND U3083 ( .A(n26), .B(n1287), .Z(n1285) );
  XOR U3084 ( .A(n1288), .B(n1289), .Z(n1287) );
  XOR U3085 ( .A(DB[1821]), .B(DB[1806]), .Z(n1289) );
  AND U3086 ( .A(n30), .B(n1290), .Z(n1288) );
  XOR U3087 ( .A(n1291), .B(n1292), .Z(n1290) );
  XOR U3088 ( .A(DB[1806]), .B(DB[1791]), .Z(n1292) );
  AND U3089 ( .A(n34), .B(n1293), .Z(n1291) );
  XOR U3090 ( .A(n1294), .B(n1295), .Z(n1293) );
  XOR U3091 ( .A(DB[1791]), .B(DB[1776]), .Z(n1295) );
  AND U3092 ( .A(n38), .B(n1296), .Z(n1294) );
  XOR U3093 ( .A(n1297), .B(n1298), .Z(n1296) );
  XOR U3094 ( .A(DB[1776]), .B(DB[1761]), .Z(n1298) );
  AND U3095 ( .A(n42), .B(n1299), .Z(n1297) );
  XOR U3096 ( .A(n1300), .B(n1301), .Z(n1299) );
  XOR U3097 ( .A(DB[1761]), .B(DB[1746]), .Z(n1301) );
  AND U3098 ( .A(n46), .B(n1302), .Z(n1300) );
  XOR U3099 ( .A(n1303), .B(n1304), .Z(n1302) );
  XOR U3100 ( .A(DB[1746]), .B(DB[1731]), .Z(n1304) );
  AND U3101 ( .A(n50), .B(n1305), .Z(n1303) );
  XOR U3102 ( .A(n1306), .B(n1307), .Z(n1305) );
  XOR U3103 ( .A(DB[1731]), .B(DB[1716]), .Z(n1307) );
  AND U3104 ( .A(n54), .B(n1308), .Z(n1306) );
  XOR U3105 ( .A(n1309), .B(n1310), .Z(n1308) );
  XOR U3106 ( .A(DB[1716]), .B(DB[1701]), .Z(n1310) );
  AND U3107 ( .A(n58), .B(n1311), .Z(n1309) );
  XOR U3108 ( .A(n1312), .B(n1313), .Z(n1311) );
  XOR U3109 ( .A(DB[1701]), .B(DB[1686]), .Z(n1313) );
  AND U3110 ( .A(n62), .B(n1314), .Z(n1312) );
  XOR U3111 ( .A(n1315), .B(n1316), .Z(n1314) );
  XOR U3112 ( .A(DB[1686]), .B(DB[1671]), .Z(n1316) );
  AND U3113 ( .A(n66), .B(n1317), .Z(n1315) );
  XOR U3114 ( .A(n1318), .B(n1319), .Z(n1317) );
  XOR U3115 ( .A(DB[1671]), .B(DB[1656]), .Z(n1319) );
  AND U3116 ( .A(n70), .B(n1320), .Z(n1318) );
  XOR U3117 ( .A(n1321), .B(n1322), .Z(n1320) );
  XOR U3118 ( .A(DB[1656]), .B(DB[1641]), .Z(n1322) );
  AND U3119 ( .A(n74), .B(n1323), .Z(n1321) );
  XOR U3120 ( .A(n1324), .B(n1325), .Z(n1323) );
  XOR U3121 ( .A(DB[1641]), .B(DB[1626]), .Z(n1325) );
  AND U3122 ( .A(n78), .B(n1326), .Z(n1324) );
  XOR U3123 ( .A(n1327), .B(n1328), .Z(n1326) );
  XOR U3124 ( .A(DB[1626]), .B(DB[1611]), .Z(n1328) );
  AND U3125 ( .A(n82), .B(n1329), .Z(n1327) );
  XOR U3126 ( .A(n1330), .B(n1331), .Z(n1329) );
  XOR U3127 ( .A(DB[1611]), .B(DB[1596]), .Z(n1331) );
  AND U3128 ( .A(n86), .B(n1332), .Z(n1330) );
  XOR U3129 ( .A(n1333), .B(n1334), .Z(n1332) );
  XOR U3130 ( .A(DB[1596]), .B(DB[1581]), .Z(n1334) );
  AND U3131 ( .A(n90), .B(n1335), .Z(n1333) );
  XOR U3132 ( .A(n1336), .B(n1337), .Z(n1335) );
  XOR U3133 ( .A(DB[1581]), .B(DB[1566]), .Z(n1337) );
  AND U3134 ( .A(n94), .B(n1338), .Z(n1336) );
  XOR U3135 ( .A(n1339), .B(n1340), .Z(n1338) );
  XOR U3136 ( .A(DB[1566]), .B(DB[1551]), .Z(n1340) );
  AND U3137 ( .A(n98), .B(n1341), .Z(n1339) );
  XOR U3138 ( .A(n1342), .B(n1343), .Z(n1341) );
  XOR U3139 ( .A(DB[1551]), .B(DB[1536]), .Z(n1343) );
  AND U3140 ( .A(n102), .B(n1344), .Z(n1342) );
  XOR U3141 ( .A(n1345), .B(n1346), .Z(n1344) );
  XOR U3142 ( .A(DB[1536]), .B(DB[1521]), .Z(n1346) );
  AND U3143 ( .A(n106), .B(n1347), .Z(n1345) );
  XOR U3144 ( .A(n1348), .B(n1349), .Z(n1347) );
  XOR U3145 ( .A(DB[1521]), .B(DB[1506]), .Z(n1349) );
  AND U3146 ( .A(n110), .B(n1350), .Z(n1348) );
  XOR U3147 ( .A(n1351), .B(n1352), .Z(n1350) );
  XOR U3148 ( .A(DB[1506]), .B(DB[1491]), .Z(n1352) );
  AND U3149 ( .A(n114), .B(n1353), .Z(n1351) );
  XOR U3150 ( .A(n1354), .B(n1355), .Z(n1353) );
  XOR U3151 ( .A(DB[1491]), .B(DB[1476]), .Z(n1355) );
  AND U3152 ( .A(n118), .B(n1356), .Z(n1354) );
  XOR U3153 ( .A(n1357), .B(n1358), .Z(n1356) );
  XOR U3154 ( .A(DB[1476]), .B(DB[1461]), .Z(n1358) );
  AND U3155 ( .A(n122), .B(n1359), .Z(n1357) );
  XOR U3156 ( .A(n1360), .B(n1361), .Z(n1359) );
  XOR U3157 ( .A(DB[1461]), .B(DB[1446]), .Z(n1361) );
  AND U3158 ( .A(n126), .B(n1362), .Z(n1360) );
  XOR U3159 ( .A(n1363), .B(n1364), .Z(n1362) );
  XOR U3160 ( .A(DB[1446]), .B(DB[1431]), .Z(n1364) );
  AND U3161 ( .A(n130), .B(n1365), .Z(n1363) );
  XOR U3162 ( .A(n1366), .B(n1367), .Z(n1365) );
  XOR U3163 ( .A(DB[1431]), .B(DB[1416]), .Z(n1367) );
  AND U3164 ( .A(n134), .B(n1368), .Z(n1366) );
  XOR U3165 ( .A(n1369), .B(n1370), .Z(n1368) );
  XOR U3166 ( .A(DB[1416]), .B(DB[1401]), .Z(n1370) );
  AND U3167 ( .A(n138), .B(n1371), .Z(n1369) );
  XOR U3168 ( .A(n1372), .B(n1373), .Z(n1371) );
  XOR U3169 ( .A(DB[1401]), .B(DB[1386]), .Z(n1373) );
  AND U3170 ( .A(n142), .B(n1374), .Z(n1372) );
  XOR U3171 ( .A(n1375), .B(n1376), .Z(n1374) );
  XOR U3172 ( .A(DB[1386]), .B(DB[1371]), .Z(n1376) );
  AND U3173 ( .A(n146), .B(n1377), .Z(n1375) );
  XOR U3174 ( .A(n1378), .B(n1379), .Z(n1377) );
  XOR U3175 ( .A(DB[1371]), .B(DB[1356]), .Z(n1379) );
  AND U3176 ( .A(n150), .B(n1380), .Z(n1378) );
  XOR U3177 ( .A(n1381), .B(n1382), .Z(n1380) );
  XOR U3178 ( .A(DB[1356]), .B(DB[1341]), .Z(n1382) );
  AND U3179 ( .A(n154), .B(n1383), .Z(n1381) );
  XOR U3180 ( .A(n1384), .B(n1385), .Z(n1383) );
  XOR U3181 ( .A(DB[1341]), .B(DB[1326]), .Z(n1385) );
  AND U3182 ( .A(n158), .B(n1386), .Z(n1384) );
  XOR U3183 ( .A(n1387), .B(n1388), .Z(n1386) );
  XOR U3184 ( .A(DB[1326]), .B(DB[1311]), .Z(n1388) );
  AND U3185 ( .A(n162), .B(n1389), .Z(n1387) );
  XOR U3186 ( .A(n1390), .B(n1391), .Z(n1389) );
  XOR U3187 ( .A(DB[1311]), .B(DB[1296]), .Z(n1391) );
  AND U3188 ( .A(n166), .B(n1392), .Z(n1390) );
  XOR U3189 ( .A(n1393), .B(n1394), .Z(n1392) );
  XOR U3190 ( .A(DB[1296]), .B(DB[1281]), .Z(n1394) );
  AND U3191 ( .A(n170), .B(n1395), .Z(n1393) );
  XOR U3192 ( .A(n1396), .B(n1397), .Z(n1395) );
  XOR U3193 ( .A(DB[1281]), .B(DB[1266]), .Z(n1397) );
  AND U3194 ( .A(n174), .B(n1398), .Z(n1396) );
  XOR U3195 ( .A(n1399), .B(n1400), .Z(n1398) );
  XOR U3196 ( .A(DB[1266]), .B(DB[1251]), .Z(n1400) );
  AND U3197 ( .A(n178), .B(n1401), .Z(n1399) );
  XOR U3198 ( .A(n1402), .B(n1403), .Z(n1401) );
  XOR U3199 ( .A(DB[1251]), .B(DB[1236]), .Z(n1403) );
  AND U3200 ( .A(n182), .B(n1404), .Z(n1402) );
  XOR U3201 ( .A(n1405), .B(n1406), .Z(n1404) );
  XOR U3202 ( .A(DB[1236]), .B(DB[1221]), .Z(n1406) );
  AND U3203 ( .A(n186), .B(n1407), .Z(n1405) );
  XOR U3204 ( .A(n1408), .B(n1409), .Z(n1407) );
  XOR U3205 ( .A(DB[1221]), .B(DB[1206]), .Z(n1409) );
  AND U3206 ( .A(n190), .B(n1410), .Z(n1408) );
  XOR U3207 ( .A(n1411), .B(n1412), .Z(n1410) );
  XOR U3208 ( .A(DB[1206]), .B(DB[1191]), .Z(n1412) );
  AND U3209 ( .A(n194), .B(n1413), .Z(n1411) );
  XOR U3210 ( .A(n1414), .B(n1415), .Z(n1413) );
  XOR U3211 ( .A(DB[1191]), .B(DB[1176]), .Z(n1415) );
  AND U3212 ( .A(n198), .B(n1416), .Z(n1414) );
  XOR U3213 ( .A(n1417), .B(n1418), .Z(n1416) );
  XOR U3214 ( .A(DB[1176]), .B(DB[1161]), .Z(n1418) );
  AND U3215 ( .A(n202), .B(n1419), .Z(n1417) );
  XOR U3216 ( .A(n1420), .B(n1421), .Z(n1419) );
  XOR U3217 ( .A(DB[1161]), .B(DB[1146]), .Z(n1421) );
  AND U3218 ( .A(n206), .B(n1422), .Z(n1420) );
  XOR U3219 ( .A(n1423), .B(n1424), .Z(n1422) );
  XOR U3220 ( .A(DB[1146]), .B(DB[1131]), .Z(n1424) );
  AND U3221 ( .A(n210), .B(n1425), .Z(n1423) );
  XOR U3222 ( .A(n1426), .B(n1427), .Z(n1425) );
  XOR U3223 ( .A(DB[1131]), .B(DB[1116]), .Z(n1427) );
  AND U3224 ( .A(n214), .B(n1428), .Z(n1426) );
  XOR U3225 ( .A(n1429), .B(n1430), .Z(n1428) );
  XOR U3226 ( .A(DB[1116]), .B(DB[1101]), .Z(n1430) );
  AND U3227 ( .A(n218), .B(n1431), .Z(n1429) );
  XOR U3228 ( .A(n1432), .B(n1433), .Z(n1431) );
  XOR U3229 ( .A(DB[1101]), .B(DB[1086]), .Z(n1433) );
  AND U3230 ( .A(n222), .B(n1434), .Z(n1432) );
  XOR U3231 ( .A(n1435), .B(n1436), .Z(n1434) );
  XOR U3232 ( .A(DB[1086]), .B(DB[1071]), .Z(n1436) );
  AND U3233 ( .A(n226), .B(n1437), .Z(n1435) );
  XOR U3234 ( .A(n1438), .B(n1439), .Z(n1437) );
  XOR U3235 ( .A(DB[1071]), .B(DB[1056]), .Z(n1439) );
  AND U3236 ( .A(n230), .B(n1440), .Z(n1438) );
  XOR U3237 ( .A(n1441), .B(n1442), .Z(n1440) );
  XOR U3238 ( .A(DB[1056]), .B(DB[1041]), .Z(n1442) );
  AND U3239 ( .A(n234), .B(n1443), .Z(n1441) );
  XOR U3240 ( .A(n1444), .B(n1445), .Z(n1443) );
  XOR U3241 ( .A(DB[1041]), .B(DB[1026]), .Z(n1445) );
  AND U3242 ( .A(n238), .B(n1446), .Z(n1444) );
  XOR U3243 ( .A(n1447), .B(n1448), .Z(n1446) );
  XOR U3244 ( .A(DB[1026]), .B(DB[1011]), .Z(n1448) );
  AND U3245 ( .A(n242), .B(n1449), .Z(n1447) );
  XOR U3246 ( .A(n1450), .B(n1451), .Z(n1449) );
  XOR U3247 ( .A(DB[996]), .B(DB[1011]), .Z(n1451) );
  AND U3248 ( .A(n246), .B(n1452), .Z(n1450) );
  XOR U3249 ( .A(n1453), .B(n1454), .Z(n1452) );
  XOR U3250 ( .A(DB[996]), .B(DB[981]), .Z(n1454) );
  AND U3251 ( .A(n250), .B(n1455), .Z(n1453) );
  XOR U3252 ( .A(n1456), .B(n1457), .Z(n1455) );
  XOR U3253 ( .A(DB[981]), .B(DB[966]), .Z(n1457) );
  AND U3254 ( .A(n254), .B(n1458), .Z(n1456) );
  XOR U3255 ( .A(n1459), .B(n1460), .Z(n1458) );
  XOR U3256 ( .A(DB[966]), .B(DB[951]), .Z(n1460) );
  AND U3257 ( .A(n258), .B(n1461), .Z(n1459) );
  XOR U3258 ( .A(n1462), .B(n1463), .Z(n1461) );
  XOR U3259 ( .A(DB[951]), .B(DB[936]), .Z(n1463) );
  AND U3260 ( .A(n262), .B(n1464), .Z(n1462) );
  XOR U3261 ( .A(n1465), .B(n1466), .Z(n1464) );
  XOR U3262 ( .A(DB[936]), .B(DB[921]), .Z(n1466) );
  AND U3263 ( .A(n266), .B(n1467), .Z(n1465) );
  XOR U3264 ( .A(n1468), .B(n1469), .Z(n1467) );
  XOR U3265 ( .A(DB[921]), .B(DB[906]), .Z(n1469) );
  AND U3266 ( .A(n270), .B(n1470), .Z(n1468) );
  XOR U3267 ( .A(n1471), .B(n1472), .Z(n1470) );
  XOR U3268 ( .A(DB[906]), .B(DB[891]), .Z(n1472) );
  AND U3269 ( .A(n274), .B(n1473), .Z(n1471) );
  XOR U3270 ( .A(n1474), .B(n1475), .Z(n1473) );
  XOR U3271 ( .A(DB[891]), .B(DB[876]), .Z(n1475) );
  AND U3272 ( .A(n278), .B(n1476), .Z(n1474) );
  XOR U3273 ( .A(n1477), .B(n1478), .Z(n1476) );
  XOR U3274 ( .A(DB[876]), .B(DB[861]), .Z(n1478) );
  AND U3275 ( .A(n282), .B(n1479), .Z(n1477) );
  XOR U3276 ( .A(n1480), .B(n1481), .Z(n1479) );
  XOR U3277 ( .A(DB[861]), .B(DB[846]), .Z(n1481) );
  AND U3278 ( .A(n286), .B(n1482), .Z(n1480) );
  XOR U3279 ( .A(n1483), .B(n1484), .Z(n1482) );
  XOR U3280 ( .A(DB[846]), .B(DB[831]), .Z(n1484) );
  AND U3281 ( .A(n290), .B(n1485), .Z(n1483) );
  XOR U3282 ( .A(n1486), .B(n1487), .Z(n1485) );
  XOR U3283 ( .A(DB[831]), .B(DB[816]), .Z(n1487) );
  AND U3284 ( .A(n294), .B(n1488), .Z(n1486) );
  XOR U3285 ( .A(n1489), .B(n1490), .Z(n1488) );
  XOR U3286 ( .A(DB[816]), .B(DB[801]), .Z(n1490) );
  AND U3287 ( .A(n298), .B(n1491), .Z(n1489) );
  XOR U3288 ( .A(n1492), .B(n1493), .Z(n1491) );
  XOR U3289 ( .A(DB[801]), .B(DB[786]), .Z(n1493) );
  AND U3290 ( .A(n302), .B(n1494), .Z(n1492) );
  XOR U3291 ( .A(n1495), .B(n1496), .Z(n1494) );
  XOR U3292 ( .A(DB[786]), .B(DB[771]), .Z(n1496) );
  AND U3293 ( .A(n306), .B(n1497), .Z(n1495) );
  XOR U3294 ( .A(n1498), .B(n1499), .Z(n1497) );
  XOR U3295 ( .A(DB[771]), .B(DB[756]), .Z(n1499) );
  AND U3296 ( .A(n310), .B(n1500), .Z(n1498) );
  XOR U3297 ( .A(n1501), .B(n1502), .Z(n1500) );
  XOR U3298 ( .A(DB[756]), .B(DB[741]), .Z(n1502) );
  AND U3299 ( .A(n314), .B(n1503), .Z(n1501) );
  XOR U3300 ( .A(n1504), .B(n1505), .Z(n1503) );
  XOR U3301 ( .A(DB[741]), .B(DB[726]), .Z(n1505) );
  AND U3302 ( .A(n318), .B(n1506), .Z(n1504) );
  XOR U3303 ( .A(n1507), .B(n1508), .Z(n1506) );
  XOR U3304 ( .A(DB[726]), .B(DB[711]), .Z(n1508) );
  AND U3305 ( .A(n322), .B(n1509), .Z(n1507) );
  XOR U3306 ( .A(n1510), .B(n1511), .Z(n1509) );
  XOR U3307 ( .A(DB[711]), .B(DB[696]), .Z(n1511) );
  AND U3308 ( .A(n326), .B(n1512), .Z(n1510) );
  XOR U3309 ( .A(n1513), .B(n1514), .Z(n1512) );
  XOR U3310 ( .A(DB[696]), .B(DB[681]), .Z(n1514) );
  AND U3311 ( .A(n330), .B(n1515), .Z(n1513) );
  XOR U3312 ( .A(n1516), .B(n1517), .Z(n1515) );
  XOR U3313 ( .A(DB[681]), .B(DB[666]), .Z(n1517) );
  AND U3314 ( .A(n334), .B(n1518), .Z(n1516) );
  XOR U3315 ( .A(n1519), .B(n1520), .Z(n1518) );
  XOR U3316 ( .A(DB[666]), .B(DB[651]), .Z(n1520) );
  AND U3317 ( .A(n338), .B(n1521), .Z(n1519) );
  XOR U3318 ( .A(n1522), .B(n1523), .Z(n1521) );
  XOR U3319 ( .A(DB[651]), .B(DB[636]), .Z(n1523) );
  AND U3320 ( .A(n342), .B(n1524), .Z(n1522) );
  XOR U3321 ( .A(n1525), .B(n1526), .Z(n1524) );
  XOR U3322 ( .A(DB[636]), .B(DB[621]), .Z(n1526) );
  AND U3323 ( .A(n346), .B(n1527), .Z(n1525) );
  XOR U3324 ( .A(n1528), .B(n1529), .Z(n1527) );
  XOR U3325 ( .A(DB[621]), .B(DB[606]), .Z(n1529) );
  AND U3326 ( .A(n350), .B(n1530), .Z(n1528) );
  XOR U3327 ( .A(n1531), .B(n1532), .Z(n1530) );
  XOR U3328 ( .A(DB[606]), .B(DB[591]), .Z(n1532) );
  AND U3329 ( .A(n354), .B(n1533), .Z(n1531) );
  XOR U3330 ( .A(n1534), .B(n1535), .Z(n1533) );
  XOR U3331 ( .A(DB[591]), .B(DB[576]), .Z(n1535) );
  AND U3332 ( .A(n358), .B(n1536), .Z(n1534) );
  XOR U3333 ( .A(n1537), .B(n1538), .Z(n1536) );
  XOR U3334 ( .A(DB[576]), .B(DB[561]), .Z(n1538) );
  AND U3335 ( .A(n362), .B(n1539), .Z(n1537) );
  XOR U3336 ( .A(n1540), .B(n1541), .Z(n1539) );
  XOR U3337 ( .A(DB[561]), .B(DB[546]), .Z(n1541) );
  AND U3338 ( .A(n366), .B(n1542), .Z(n1540) );
  XOR U3339 ( .A(n1543), .B(n1544), .Z(n1542) );
  XOR U3340 ( .A(DB[546]), .B(DB[531]), .Z(n1544) );
  AND U3341 ( .A(n370), .B(n1545), .Z(n1543) );
  XOR U3342 ( .A(n1546), .B(n1547), .Z(n1545) );
  XOR U3343 ( .A(DB[531]), .B(DB[516]), .Z(n1547) );
  AND U3344 ( .A(n374), .B(n1548), .Z(n1546) );
  XOR U3345 ( .A(n1549), .B(n1550), .Z(n1548) );
  XOR U3346 ( .A(DB[516]), .B(DB[501]), .Z(n1550) );
  AND U3347 ( .A(n378), .B(n1551), .Z(n1549) );
  XOR U3348 ( .A(n1552), .B(n1553), .Z(n1551) );
  XOR U3349 ( .A(DB[501]), .B(DB[486]), .Z(n1553) );
  AND U3350 ( .A(n382), .B(n1554), .Z(n1552) );
  XOR U3351 ( .A(n1555), .B(n1556), .Z(n1554) );
  XOR U3352 ( .A(DB[486]), .B(DB[471]), .Z(n1556) );
  AND U3353 ( .A(n386), .B(n1557), .Z(n1555) );
  XOR U3354 ( .A(n1558), .B(n1559), .Z(n1557) );
  XOR U3355 ( .A(DB[471]), .B(DB[456]), .Z(n1559) );
  AND U3356 ( .A(n390), .B(n1560), .Z(n1558) );
  XOR U3357 ( .A(n1561), .B(n1562), .Z(n1560) );
  XOR U3358 ( .A(DB[456]), .B(DB[441]), .Z(n1562) );
  AND U3359 ( .A(n394), .B(n1563), .Z(n1561) );
  XOR U3360 ( .A(n1564), .B(n1565), .Z(n1563) );
  XOR U3361 ( .A(DB[441]), .B(DB[426]), .Z(n1565) );
  AND U3362 ( .A(n398), .B(n1566), .Z(n1564) );
  XOR U3363 ( .A(n1567), .B(n1568), .Z(n1566) );
  XOR U3364 ( .A(DB[426]), .B(DB[411]), .Z(n1568) );
  AND U3365 ( .A(n402), .B(n1569), .Z(n1567) );
  XOR U3366 ( .A(n1570), .B(n1571), .Z(n1569) );
  XOR U3367 ( .A(DB[411]), .B(DB[396]), .Z(n1571) );
  AND U3368 ( .A(n406), .B(n1572), .Z(n1570) );
  XOR U3369 ( .A(n1573), .B(n1574), .Z(n1572) );
  XOR U3370 ( .A(DB[396]), .B(DB[381]), .Z(n1574) );
  AND U3371 ( .A(n410), .B(n1575), .Z(n1573) );
  XOR U3372 ( .A(n1576), .B(n1577), .Z(n1575) );
  XOR U3373 ( .A(DB[381]), .B(DB[366]), .Z(n1577) );
  AND U3374 ( .A(n414), .B(n1578), .Z(n1576) );
  XOR U3375 ( .A(n1579), .B(n1580), .Z(n1578) );
  XOR U3376 ( .A(DB[366]), .B(DB[351]), .Z(n1580) );
  AND U3377 ( .A(n418), .B(n1581), .Z(n1579) );
  XOR U3378 ( .A(n1582), .B(n1583), .Z(n1581) );
  XOR U3379 ( .A(DB[351]), .B(DB[336]), .Z(n1583) );
  AND U3380 ( .A(n422), .B(n1584), .Z(n1582) );
  XOR U3381 ( .A(n1585), .B(n1586), .Z(n1584) );
  XOR U3382 ( .A(DB[336]), .B(DB[321]), .Z(n1586) );
  AND U3383 ( .A(n426), .B(n1587), .Z(n1585) );
  XOR U3384 ( .A(n1588), .B(n1589), .Z(n1587) );
  XOR U3385 ( .A(DB[321]), .B(DB[306]), .Z(n1589) );
  AND U3386 ( .A(n430), .B(n1590), .Z(n1588) );
  XOR U3387 ( .A(n1591), .B(n1592), .Z(n1590) );
  XOR U3388 ( .A(DB[306]), .B(DB[291]), .Z(n1592) );
  AND U3389 ( .A(n434), .B(n1593), .Z(n1591) );
  XOR U3390 ( .A(n1594), .B(n1595), .Z(n1593) );
  XOR U3391 ( .A(DB[291]), .B(DB[276]), .Z(n1595) );
  AND U3392 ( .A(n438), .B(n1596), .Z(n1594) );
  XOR U3393 ( .A(n1597), .B(n1598), .Z(n1596) );
  XOR U3394 ( .A(DB[276]), .B(DB[261]), .Z(n1598) );
  AND U3395 ( .A(n442), .B(n1599), .Z(n1597) );
  XOR U3396 ( .A(n1600), .B(n1601), .Z(n1599) );
  XOR U3397 ( .A(DB[261]), .B(DB[246]), .Z(n1601) );
  AND U3398 ( .A(n446), .B(n1602), .Z(n1600) );
  XOR U3399 ( .A(n1603), .B(n1604), .Z(n1602) );
  XOR U3400 ( .A(DB[246]), .B(DB[231]), .Z(n1604) );
  AND U3401 ( .A(n450), .B(n1605), .Z(n1603) );
  XOR U3402 ( .A(n1606), .B(n1607), .Z(n1605) );
  XOR U3403 ( .A(DB[231]), .B(DB[216]), .Z(n1607) );
  AND U3404 ( .A(n454), .B(n1608), .Z(n1606) );
  XOR U3405 ( .A(n1609), .B(n1610), .Z(n1608) );
  XOR U3406 ( .A(DB[216]), .B(DB[201]), .Z(n1610) );
  AND U3407 ( .A(n458), .B(n1611), .Z(n1609) );
  XOR U3408 ( .A(n1612), .B(n1613), .Z(n1611) );
  XOR U3409 ( .A(DB[201]), .B(DB[186]), .Z(n1613) );
  AND U3410 ( .A(n462), .B(n1614), .Z(n1612) );
  XOR U3411 ( .A(n1615), .B(n1616), .Z(n1614) );
  XOR U3412 ( .A(DB[186]), .B(DB[171]), .Z(n1616) );
  AND U3413 ( .A(n466), .B(n1617), .Z(n1615) );
  XOR U3414 ( .A(n1618), .B(n1619), .Z(n1617) );
  XOR U3415 ( .A(DB[171]), .B(DB[156]), .Z(n1619) );
  AND U3416 ( .A(n470), .B(n1620), .Z(n1618) );
  XOR U3417 ( .A(n1621), .B(n1622), .Z(n1620) );
  XOR U3418 ( .A(DB[156]), .B(DB[141]), .Z(n1622) );
  AND U3419 ( .A(n474), .B(n1623), .Z(n1621) );
  XOR U3420 ( .A(n1624), .B(n1625), .Z(n1623) );
  XOR U3421 ( .A(DB[141]), .B(DB[126]), .Z(n1625) );
  AND U3422 ( .A(n478), .B(n1626), .Z(n1624) );
  XOR U3423 ( .A(n1627), .B(n1628), .Z(n1626) );
  XOR U3424 ( .A(DB[126]), .B(DB[111]), .Z(n1628) );
  AND U3425 ( .A(n482), .B(n1629), .Z(n1627) );
  XOR U3426 ( .A(n1630), .B(n1631), .Z(n1629) );
  XOR U3427 ( .A(DB[96]), .B(DB[111]), .Z(n1631) );
  AND U3428 ( .A(n486), .B(n1632), .Z(n1630) );
  XOR U3429 ( .A(n1633), .B(n1634), .Z(n1632) );
  XOR U3430 ( .A(DB[96]), .B(DB[81]), .Z(n1634) );
  AND U3431 ( .A(n490), .B(n1635), .Z(n1633) );
  XOR U3432 ( .A(n1636), .B(n1637), .Z(n1635) );
  XOR U3433 ( .A(DB[81]), .B(DB[66]), .Z(n1637) );
  AND U3434 ( .A(n494), .B(n1638), .Z(n1636) );
  XOR U3435 ( .A(n1639), .B(n1640), .Z(n1638) );
  XOR U3436 ( .A(DB[66]), .B(DB[51]), .Z(n1640) );
  AND U3437 ( .A(n498), .B(n1641), .Z(n1639) );
  XOR U3438 ( .A(n1642), .B(n1643), .Z(n1641) );
  XOR U3439 ( .A(DB[51]), .B(DB[36]), .Z(n1643) );
  AND U3440 ( .A(n502), .B(n1644), .Z(n1642) );
  XOR U3441 ( .A(n1645), .B(n1646), .Z(n1644) );
  XOR U3442 ( .A(DB[36]), .B(DB[21]), .Z(n1646) );
  AND U3443 ( .A(n506), .B(n1647), .Z(n1645) );
  XOR U3444 ( .A(DB[6]), .B(DB[21]), .Z(n1647) );
  XOR U3445 ( .A(DB[1910]), .B(n1648), .Z(min_val_out[5]) );
  AND U3446 ( .A(n2), .B(n1649), .Z(n1648) );
  XOR U3447 ( .A(n1650), .B(n1651), .Z(n1649) );
  XOR U3448 ( .A(DB[1910]), .B(DB[1895]), .Z(n1651) );
  AND U3449 ( .A(n6), .B(n1652), .Z(n1650) );
  XOR U3450 ( .A(n1653), .B(n1654), .Z(n1652) );
  XOR U3451 ( .A(DB[1895]), .B(DB[1880]), .Z(n1654) );
  AND U3452 ( .A(n10), .B(n1655), .Z(n1653) );
  XOR U3453 ( .A(n1656), .B(n1657), .Z(n1655) );
  XOR U3454 ( .A(DB[1880]), .B(DB[1865]), .Z(n1657) );
  AND U3455 ( .A(n14), .B(n1658), .Z(n1656) );
  XOR U3456 ( .A(n1659), .B(n1660), .Z(n1658) );
  XOR U3457 ( .A(DB[1865]), .B(DB[1850]), .Z(n1660) );
  AND U3458 ( .A(n18), .B(n1661), .Z(n1659) );
  XOR U3459 ( .A(n1662), .B(n1663), .Z(n1661) );
  XOR U3460 ( .A(DB[1850]), .B(DB[1835]), .Z(n1663) );
  AND U3461 ( .A(n22), .B(n1664), .Z(n1662) );
  XOR U3462 ( .A(n1665), .B(n1666), .Z(n1664) );
  XOR U3463 ( .A(DB[1835]), .B(DB[1820]), .Z(n1666) );
  AND U3464 ( .A(n26), .B(n1667), .Z(n1665) );
  XOR U3465 ( .A(n1668), .B(n1669), .Z(n1667) );
  XOR U3466 ( .A(DB[1820]), .B(DB[1805]), .Z(n1669) );
  AND U3467 ( .A(n30), .B(n1670), .Z(n1668) );
  XOR U3468 ( .A(n1671), .B(n1672), .Z(n1670) );
  XOR U3469 ( .A(DB[1805]), .B(DB[1790]), .Z(n1672) );
  AND U3470 ( .A(n34), .B(n1673), .Z(n1671) );
  XOR U3471 ( .A(n1674), .B(n1675), .Z(n1673) );
  XOR U3472 ( .A(DB[1790]), .B(DB[1775]), .Z(n1675) );
  AND U3473 ( .A(n38), .B(n1676), .Z(n1674) );
  XOR U3474 ( .A(n1677), .B(n1678), .Z(n1676) );
  XOR U3475 ( .A(DB[1775]), .B(DB[1760]), .Z(n1678) );
  AND U3476 ( .A(n42), .B(n1679), .Z(n1677) );
  XOR U3477 ( .A(n1680), .B(n1681), .Z(n1679) );
  XOR U3478 ( .A(DB[1760]), .B(DB[1745]), .Z(n1681) );
  AND U3479 ( .A(n46), .B(n1682), .Z(n1680) );
  XOR U3480 ( .A(n1683), .B(n1684), .Z(n1682) );
  XOR U3481 ( .A(DB[1745]), .B(DB[1730]), .Z(n1684) );
  AND U3482 ( .A(n50), .B(n1685), .Z(n1683) );
  XOR U3483 ( .A(n1686), .B(n1687), .Z(n1685) );
  XOR U3484 ( .A(DB[1730]), .B(DB[1715]), .Z(n1687) );
  AND U3485 ( .A(n54), .B(n1688), .Z(n1686) );
  XOR U3486 ( .A(n1689), .B(n1690), .Z(n1688) );
  XOR U3487 ( .A(DB[1715]), .B(DB[1700]), .Z(n1690) );
  AND U3488 ( .A(n58), .B(n1691), .Z(n1689) );
  XOR U3489 ( .A(n1692), .B(n1693), .Z(n1691) );
  XOR U3490 ( .A(DB[1700]), .B(DB[1685]), .Z(n1693) );
  AND U3491 ( .A(n62), .B(n1694), .Z(n1692) );
  XOR U3492 ( .A(n1695), .B(n1696), .Z(n1694) );
  XOR U3493 ( .A(DB[1685]), .B(DB[1670]), .Z(n1696) );
  AND U3494 ( .A(n66), .B(n1697), .Z(n1695) );
  XOR U3495 ( .A(n1698), .B(n1699), .Z(n1697) );
  XOR U3496 ( .A(DB[1670]), .B(DB[1655]), .Z(n1699) );
  AND U3497 ( .A(n70), .B(n1700), .Z(n1698) );
  XOR U3498 ( .A(n1701), .B(n1702), .Z(n1700) );
  XOR U3499 ( .A(DB[1655]), .B(DB[1640]), .Z(n1702) );
  AND U3500 ( .A(n74), .B(n1703), .Z(n1701) );
  XOR U3501 ( .A(n1704), .B(n1705), .Z(n1703) );
  XOR U3502 ( .A(DB[1640]), .B(DB[1625]), .Z(n1705) );
  AND U3503 ( .A(n78), .B(n1706), .Z(n1704) );
  XOR U3504 ( .A(n1707), .B(n1708), .Z(n1706) );
  XOR U3505 ( .A(DB[1625]), .B(DB[1610]), .Z(n1708) );
  AND U3506 ( .A(n82), .B(n1709), .Z(n1707) );
  XOR U3507 ( .A(n1710), .B(n1711), .Z(n1709) );
  XOR U3508 ( .A(DB[1610]), .B(DB[1595]), .Z(n1711) );
  AND U3509 ( .A(n86), .B(n1712), .Z(n1710) );
  XOR U3510 ( .A(n1713), .B(n1714), .Z(n1712) );
  XOR U3511 ( .A(DB[1595]), .B(DB[1580]), .Z(n1714) );
  AND U3512 ( .A(n90), .B(n1715), .Z(n1713) );
  XOR U3513 ( .A(n1716), .B(n1717), .Z(n1715) );
  XOR U3514 ( .A(DB[1580]), .B(DB[1565]), .Z(n1717) );
  AND U3515 ( .A(n94), .B(n1718), .Z(n1716) );
  XOR U3516 ( .A(n1719), .B(n1720), .Z(n1718) );
  XOR U3517 ( .A(DB[1565]), .B(DB[1550]), .Z(n1720) );
  AND U3518 ( .A(n98), .B(n1721), .Z(n1719) );
  XOR U3519 ( .A(n1722), .B(n1723), .Z(n1721) );
  XOR U3520 ( .A(DB[1550]), .B(DB[1535]), .Z(n1723) );
  AND U3521 ( .A(n102), .B(n1724), .Z(n1722) );
  XOR U3522 ( .A(n1725), .B(n1726), .Z(n1724) );
  XOR U3523 ( .A(DB[1535]), .B(DB[1520]), .Z(n1726) );
  AND U3524 ( .A(n106), .B(n1727), .Z(n1725) );
  XOR U3525 ( .A(n1728), .B(n1729), .Z(n1727) );
  XOR U3526 ( .A(DB[1520]), .B(DB[1505]), .Z(n1729) );
  AND U3527 ( .A(n110), .B(n1730), .Z(n1728) );
  XOR U3528 ( .A(n1731), .B(n1732), .Z(n1730) );
  XOR U3529 ( .A(DB[1505]), .B(DB[1490]), .Z(n1732) );
  AND U3530 ( .A(n114), .B(n1733), .Z(n1731) );
  XOR U3531 ( .A(n1734), .B(n1735), .Z(n1733) );
  XOR U3532 ( .A(DB[1490]), .B(DB[1475]), .Z(n1735) );
  AND U3533 ( .A(n118), .B(n1736), .Z(n1734) );
  XOR U3534 ( .A(n1737), .B(n1738), .Z(n1736) );
  XOR U3535 ( .A(DB[1475]), .B(DB[1460]), .Z(n1738) );
  AND U3536 ( .A(n122), .B(n1739), .Z(n1737) );
  XOR U3537 ( .A(n1740), .B(n1741), .Z(n1739) );
  XOR U3538 ( .A(DB[1460]), .B(DB[1445]), .Z(n1741) );
  AND U3539 ( .A(n126), .B(n1742), .Z(n1740) );
  XOR U3540 ( .A(n1743), .B(n1744), .Z(n1742) );
  XOR U3541 ( .A(DB[1445]), .B(DB[1430]), .Z(n1744) );
  AND U3542 ( .A(n130), .B(n1745), .Z(n1743) );
  XOR U3543 ( .A(n1746), .B(n1747), .Z(n1745) );
  XOR U3544 ( .A(DB[1430]), .B(DB[1415]), .Z(n1747) );
  AND U3545 ( .A(n134), .B(n1748), .Z(n1746) );
  XOR U3546 ( .A(n1749), .B(n1750), .Z(n1748) );
  XOR U3547 ( .A(DB[1415]), .B(DB[1400]), .Z(n1750) );
  AND U3548 ( .A(n138), .B(n1751), .Z(n1749) );
  XOR U3549 ( .A(n1752), .B(n1753), .Z(n1751) );
  XOR U3550 ( .A(DB[1400]), .B(DB[1385]), .Z(n1753) );
  AND U3551 ( .A(n142), .B(n1754), .Z(n1752) );
  XOR U3552 ( .A(n1755), .B(n1756), .Z(n1754) );
  XOR U3553 ( .A(DB[1385]), .B(DB[1370]), .Z(n1756) );
  AND U3554 ( .A(n146), .B(n1757), .Z(n1755) );
  XOR U3555 ( .A(n1758), .B(n1759), .Z(n1757) );
  XOR U3556 ( .A(DB[1370]), .B(DB[1355]), .Z(n1759) );
  AND U3557 ( .A(n150), .B(n1760), .Z(n1758) );
  XOR U3558 ( .A(n1761), .B(n1762), .Z(n1760) );
  XOR U3559 ( .A(DB[1355]), .B(DB[1340]), .Z(n1762) );
  AND U3560 ( .A(n154), .B(n1763), .Z(n1761) );
  XOR U3561 ( .A(n1764), .B(n1765), .Z(n1763) );
  XOR U3562 ( .A(DB[1340]), .B(DB[1325]), .Z(n1765) );
  AND U3563 ( .A(n158), .B(n1766), .Z(n1764) );
  XOR U3564 ( .A(n1767), .B(n1768), .Z(n1766) );
  XOR U3565 ( .A(DB[1325]), .B(DB[1310]), .Z(n1768) );
  AND U3566 ( .A(n162), .B(n1769), .Z(n1767) );
  XOR U3567 ( .A(n1770), .B(n1771), .Z(n1769) );
  XOR U3568 ( .A(DB[1310]), .B(DB[1295]), .Z(n1771) );
  AND U3569 ( .A(n166), .B(n1772), .Z(n1770) );
  XOR U3570 ( .A(n1773), .B(n1774), .Z(n1772) );
  XOR U3571 ( .A(DB[1295]), .B(DB[1280]), .Z(n1774) );
  AND U3572 ( .A(n170), .B(n1775), .Z(n1773) );
  XOR U3573 ( .A(n1776), .B(n1777), .Z(n1775) );
  XOR U3574 ( .A(DB[1280]), .B(DB[1265]), .Z(n1777) );
  AND U3575 ( .A(n174), .B(n1778), .Z(n1776) );
  XOR U3576 ( .A(n1779), .B(n1780), .Z(n1778) );
  XOR U3577 ( .A(DB[1265]), .B(DB[1250]), .Z(n1780) );
  AND U3578 ( .A(n178), .B(n1781), .Z(n1779) );
  XOR U3579 ( .A(n1782), .B(n1783), .Z(n1781) );
  XOR U3580 ( .A(DB[1250]), .B(DB[1235]), .Z(n1783) );
  AND U3581 ( .A(n182), .B(n1784), .Z(n1782) );
  XOR U3582 ( .A(n1785), .B(n1786), .Z(n1784) );
  XOR U3583 ( .A(DB[1235]), .B(DB[1220]), .Z(n1786) );
  AND U3584 ( .A(n186), .B(n1787), .Z(n1785) );
  XOR U3585 ( .A(n1788), .B(n1789), .Z(n1787) );
  XOR U3586 ( .A(DB[1220]), .B(DB[1205]), .Z(n1789) );
  AND U3587 ( .A(n190), .B(n1790), .Z(n1788) );
  XOR U3588 ( .A(n1791), .B(n1792), .Z(n1790) );
  XOR U3589 ( .A(DB[1205]), .B(DB[1190]), .Z(n1792) );
  AND U3590 ( .A(n194), .B(n1793), .Z(n1791) );
  XOR U3591 ( .A(n1794), .B(n1795), .Z(n1793) );
  XOR U3592 ( .A(DB[1190]), .B(DB[1175]), .Z(n1795) );
  AND U3593 ( .A(n198), .B(n1796), .Z(n1794) );
  XOR U3594 ( .A(n1797), .B(n1798), .Z(n1796) );
  XOR U3595 ( .A(DB[1175]), .B(DB[1160]), .Z(n1798) );
  AND U3596 ( .A(n202), .B(n1799), .Z(n1797) );
  XOR U3597 ( .A(n1800), .B(n1801), .Z(n1799) );
  XOR U3598 ( .A(DB[1160]), .B(DB[1145]), .Z(n1801) );
  AND U3599 ( .A(n206), .B(n1802), .Z(n1800) );
  XOR U3600 ( .A(n1803), .B(n1804), .Z(n1802) );
  XOR U3601 ( .A(DB[1145]), .B(DB[1130]), .Z(n1804) );
  AND U3602 ( .A(n210), .B(n1805), .Z(n1803) );
  XOR U3603 ( .A(n1806), .B(n1807), .Z(n1805) );
  XOR U3604 ( .A(DB[1130]), .B(DB[1115]), .Z(n1807) );
  AND U3605 ( .A(n214), .B(n1808), .Z(n1806) );
  XOR U3606 ( .A(n1809), .B(n1810), .Z(n1808) );
  XOR U3607 ( .A(DB[1115]), .B(DB[1100]), .Z(n1810) );
  AND U3608 ( .A(n218), .B(n1811), .Z(n1809) );
  XOR U3609 ( .A(n1812), .B(n1813), .Z(n1811) );
  XOR U3610 ( .A(DB[1100]), .B(DB[1085]), .Z(n1813) );
  AND U3611 ( .A(n222), .B(n1814), .Z(n1812) );
  XOR U3612 ( .A(n1815), .B(n1816), .Z(n1814) );
  XOR U3613 ( .A(DB[1085]), .B(DB[1070]), .Z(n1816) );
  AND U3614 ( .A(n226), .B(n1817), .Z(n1815) );
  XOR U3615 ( .A(n1818), .B(n1819), .Z(n1817) );
  XOR U3616 ( .A(DB[1070]), .B(DB[1055]), .Z(n1819) );
  AND U3617 ( .A(n230), .B(n1820), .Z(n1818) );
  XOR U3618 ( .A(n1821), .B(n1822), .Z(n1820) );
  XOR U3619 ( .A(DB[1055]), .B(DB[1040]), .Z(n1822) );
  AND U3620 ( .A(n234), .B(n1823), .Z(n1821) );
  XOR U3621 ( .A(n1824), .B(n1825), .Z(n1823) );
  XOR U3622 ( .A(DB[1040]), .B(DB[1025]), .Z(n1825) );
  AND U3623 ( .A(n238), .B(n1826), .Z(n1824) );
  XOR U3624 ( .A(n1827), .B(n1828), .Z(n1826) );
  XOR U3625 ( .A(DB[1025]), .B(DB[1010]), .Z(n1828) );
  AND U3626 ( .A(n242), .B(n1829), .Z(n1827) );
  XOR U3627 ( .A(n1830), .B(n1831), .Z(n1829) );
  XOR U3628 ( .A(DB[995]), .B(DB[1010]), .Z(n1831) );
  AND U3629 ( .A(n246), .B(n1832), .Z(n1830) );
  XOR U3630 ( .A(n1833), .B(n1834), .Z(n1832) );
  XOR U3631 ( .A(DB[995]), .B(DB[980]), .Z(n1834) );
  AND U3632 ( .A(n250), .B(n1835), .Z(n1833) );
  XOR U3633 ( .A(n1836), .B(n1837), .Z(n1835) );
  XOR U3634 ( .A(DB[980]), .B(DB[965]), .Z(n1837) );
  AND U3635 ( .A(n254), .B(n1838), .Z(n1836) );
  XOR U3636 ( .A(n1839), .B(n1840), .Z(n1838) );
  XOR U3637 ( .A(DB[965]), .B(DB[950]), .Z(n1840) );
  AND U3638 ( .A(n258), .B(n1841), .Z(n1839) );
  XOR U3639 ( .A(n1842), .B(n1843), .Z(n1841) );
  XOR U3640 ( .A(DB[950]), .B(DB[935]), .Z(n1843) );
  AND U3641 ( .A(n262), .B(n1844), .Z(n1842) );
  XOR U3642 ( .A(n1845), .B(n1846), .Z(n1844) );
  XOR U3643 ( .A(DB[935]), .B(DB[920]), .Z(n1846) );
  AND U3644 ( .A(n266), .B(n1847), .Z(n1845) );
  XOR U3645 ( .A(n1848), .B(n1849), .Z(n1847) );
  XOR U3646 ( .A(DB[920]), .B(DB[905]), .Z(n1849) );
  AND U3647 ( .A(n270), .B(n1850), .Z(n1848) );
  XOR U3648 ( .A(n1851), .B(n1852), .Z(n1850) );
  XOR U3649 ( .A(DB[905]), .B(DB[890]), .Z(n1852) );
  AND U3650 ( .A(n274), .B(n1853), .Z(n1851) );
  XOR U3651 ( .A(n1854), .B(n1855), .Z(n1853) );
  XOR U3652 ( .A(DB[890]), .B(DB[875]), .Z(n1855) );
  AND U3653 ( .A(n278), .B(n1856), .Z(n1854) );
  XOR U3654 ( .A(n1857), .B(n1858), .Z(n1856) );
  XOR U3655 ( .A(DB[875]), .B(DB[860]), .Z(n1858) );
  AND U3656 ( .A(n282), .B(n1859), .Z(n1857) );
  XOR U3657 ( .A(n1860), .B(n1861), .Z(n1859) );
  XOR U3658 ( .A(DB[860]), .B(DB[845]), .Z(n1861) );
  AND U3659 ( .A(n286), .B(n1862), .Z(n1860) );
  XOR U3660 ( .A(n1863), .B(n1864), .Z(n1862) );
  XOR U3661 ( .A(DB[845]), .B(DB[830]), .Z(n1864) );
  AND U3662 ( .A(n290), .B(n1865), .Z(n1863) );
  XOR U3663 ( .A(n1866), .B(n1867), .Z(n1865) );
  XOR U3664 ( .A(DB[830]), .B(DB[815]), .Z(n1867) );
  AND U3665 ( .A(n294), .B(n1868), .Z(n1866) );
  XOR U3666 ( .A(n1869), .B(n1870), .Z(n1868) );
  XOR U3667 ( .A(DB[815]), .B(DB[800]), .Z(n1870) );
  AND U3668 ( .A(n298), .B(n1871), .Z(n1869) );
  XOR U3669 ( .A(n1872), .B(n1873), .Z(n1871) );
  XOR U3670 ( .A(DB[800]), .B(DB[785]), .Z(n1873) );
  AND U3671 ( .A(n302), .B(n1874), .Z(n1872) );
  XOR U3672 ( .A(n1875), .B(n1876), .Z(n1874) );
  XOR U3673 ( .A(DB[785]), .B(DB[770]), .Z(n1876) );
  AND U3674 ( .A(n306), .B(n1877), .Z(n1875) );
  XOR U3675 ( .A(n1878), .B(n1879), .Z(n1877) );
  XOR U3676 ( .A(DB[770]), .B(DB[755]), .Z(n1879) );
  AND U3677 ( .A(n310), .B(n1880), .Z(n1878) );
  XOR U3678 ( .A(n1881), .B(n1882), .Z(n1880) );
  XOR U3679 ( .A(DB[755]), .B(DB[740]), .Z(n1882) );
  AND U3680 ( .A(n314), .B(n1883), .Z(n1881) );
  XOR U3681 ( .A(n1884), .B(n1885), .Z(n1883) );
  XOR U3682 ( .A(DB[740]), .B(DB[725]), .Z(n1885) );
  AND U3683 ( .A(n318), .B(n1886), .Z(n1884) );
  XOR U3684 ( .A(n1887), .B(n1888), .Z(n1886) );
  XOR U3685 ( .A(DB[725]), .B(DB[710]), .Z(n1888) );
  AND U3686 ( .A(n322), .B(n1889), .Z(n1887) );
  XOR U3687 ( .A(n1890), .B(n1891), .Z(n1889) );
  XOR U3688 ( .A(DB[710]), .B(DB[695]), .Z(n1891) );
  AND U3689 ( .A(n326), .B(n1892), .Z(n1890) );
  XOR U3690 ( .A(n1893), .B(n1894), .Z(n1892) );
  XOR U3691 ( .A(DB[695]), .B(DB[680]), .Z(n1894) );
  AND U3692 ( .A(n330), .B(n1895), .Z(n1893) );
  XOR U3693 ( .A(n1896), .B(n1897), .Z(n1895) );
  XOR U3694 ( .A(DB[680]), .B(DB[665]), .Z(n1897) );
  AND U3695 ( .A(n334), .B(n1898), .Z(n1896) );
  XOR U3696 ( .A(n1899), .B(n1900), .Z(n1898) );
  XOR U3697 ( .A(DB[665]), .B(DB[650]), .Z(n1900) );
  AND U3698 ( .A(n338), .B(n1901), .Z(n1899) );
  XOR U3699 ( .A(n1902), .B(n1903), .Z(n1901) );
  XOR U3700 ( .A(DB[650]), .B(DB[635]), .Z(n1903) );
  AND U3701 ( .A(n342), .B(n1904), .Z(n1902) );
  XOR U3702 ( .A(n1905), .B(n1906), .Z(n1904) );
  XOR U3703 ( .A(DB[635]), .B(DB[620]), .Z(n1906) );
  AND U3704 ( .A(n346), .B(n1907), .Z(n1905) );
  XOR U3705 ( .A(n1908), .B(n1909), .Z(n1907) );
  XOR U3706 ( .A(DB[620]), .B(DB[605]), .Z(n1909) );
  AND U3707 ( .A(n350), .B(n1910), .Z(n1908) );
  XOR U3708 ( .A(n1911), .B(n1912), .Z(n1910) );
  XOR U3709 ( .A(DB[605]), .B(DB[590]), .Z(n1912) );
  AND U3710 ( .A(n354), .B(n1913), .Z(n1911) );
  XOR U3711 ( .A(n1914), .B(n1915), .Z(n1913) );
  XOR U3712 ( .A(DB[590]), .B(DB[575]), .Z(n1915) );
  AND U3713 ( .A(n358), .B(n1916), .Z(n1914) );
  XOR U3714 ( .A(n1917), .B(n1918), .Z(n1916) );
  XOR U3715 ( .A(DB[575]), .B(DB[560]), .Z(n1918) );
  AND U3716 ( .A(n362), .B(n1919), .Z(n1917) );
  XOR U3717 ( .A(n1920), .B(n1921), .Z(n1919) );
  XOR U3718 ( .A(DB[560]), .B(DB[545]), .Z(n1921) );
  AND U3719 ( .A(n366), .B(n1922), .Z(n1920) );
  XOR U3720 ( .A(n1923), .B(n1924), .Z(n1922) );
  XOR U3721 ( .A(DB[545]), .B(DB[530]), .Z(n1924) );
  AND U3722 ( .A(n370), .B(n1925), .Z(n1923) );
  XOR U3723 ( .A(n1926), .B(n1927), .Z(n1925) );
  XOR U3724 ( .A(DB[530]), .B(DB[515]), .Z(n1927) );
  AND U3725 ( .A(n374), .B(n1928), .Z(n1926) );
  XOR U3726 ( .A(n1929), .B(n1930), .Z(n1928) );
  XOR U3727 ( .A(DB[515]), .B(DB[500]), .Z(n1930) );
  AND U3728 ( .A(n378), .B(n1931), .Z(n1929) );
  XOR U3729 ( .A(n1932), .B(n1933), .Z(n1931) );
  XOR U3730 ( .A(DB[500]), .B(DB[485]), .Z(n1933) );
  AND U3731 ( .A(n382), .B(n1934), .Z(n1932) );
  XOR U3732 ( .A(n1935), .B(n1936), .Z(n1934) );
  XOR U3733 ( .A(DB[485]), .B(DB[470]), .Z(n1936) );
  AND U3734 ( .A(n386), .B(n1937), .Z(n1935) );
  XOR U3735 ( .A(n1938), .B(n1939), .Z(n1937) );
  XOR U3736 ( .A(DB[470]), .B(DB[455]), .Z(n1939) );
  AND U3737 ( .A(n390), .B(n1940), .Z(n1938) );
  XOR U3738 ( .A(n1941), .B(n1942), .Z(n1940) );
  XOR U3739 ( .A(DB[455]), .B(DB[440]), .Z(n1942) );
  AND U3740 ( .A(n394), .B(n1943), .Z(n1941) );
  XOR U3741 ( .A(n1944), .B(n1945), .Z(n1943) );
  XOR U3742 ( .A(DB[440]), .B(DB[425]), .Z(n1945) );
  AND U3743 ( .A(n398), .B(n1946), .Z(n1944) );
  XOR U3744 ( .A(n1947), .B(n1948), .Z(n1946) );
  XOR U3745 ( .A(DB[425]), .B(DB[410]), .Z(n1948) );
  AND U3746 ( .A(n402), .B(n1949), .Z(n1947) );
  XOR U3747 ( .A(n1950), .B(n1951), .Z(n1949) );
  XOR U3748 ( .A(DB[410]), .B(DB[395]), .Z(n1951) );
  AND U3749 ( .A(n406), .B(n1952), .Z(n1950) );
  XOR U3750 ( .A(n1953), .B(n1954), .Z(n1952) );
  XOR U3751 ( .A(DB[395]), .B(DB[380]), .Z(n1954) );
  AND U3752 ( .A(n410), .B(n1955), .Z(n1953) );
  XOR U3753 ( .A(n1956), .B(n1957), .Z(n1955) );
  XOR U3754 ( .A(DB[380]), .B(DB[365]), .Z(n1957) );
  AND U3755 ( .A(n414), .B(n1958), .Z(n1956) );
  XOR U3756 ( .A(n1959), .B(n1960), .Z(n1958) );
  XOR U3757 ( .A(DB[365]), .B(DB[350]), .Z(n1960) );
  AND U3758 ( .A(n418), .B(n1961), .Z(n1959) );
  XOR U3759 ( .A(n1962), .B(n1963), .Z(n1961) );
  XOR U3760 ( .A(DB[350]), .B(DB[335]), .Z(n1963) );
  AND U3761 ( .A(n422), .B(n1964), .Z(n1962) );
  XOR U3762 ( .A(n1965), .B(n1966), .Z(n1964) );
  XOR U3763 ( .A(DB[335]), .B(DB[320]), .Z(n1966) );
  AND U3764 ( .A(n426), .B(n1967), .Z(n1965) );
  XOR U3765 ( .A(n1968), .B(n1969), .Z(n1967) );
  XOR U3766 ( .A(DB[320]), .B(DB[305]), .Z(n1969) );
  AND U3767 ( .A(n430), .B(n1970), .Z(n1968) );
  XOR U3768 ( .A(n1971), .B(n1972), .Z(n1970) );
  XOR U3769 ( .A(DB[305]), .B(DB[290]), .Z(n1972) );
  AND U3770 ( .A(n434), .B(n1973), .Z(n1971) );
  XOR U3771 ( .A(n1974), .B(n1975), .Z(n1973) );
  XOR U3772 ( .A(DB[290]), .B(DB[275]), .Z(n1975) );
  AND U3773 ( .A(n438), .B(n1976), .Z(n1974) );
  XOR U3774 ( .A(n1977), .B(n1978), .Z(n1976) );
  XOR U3775 ( .A(DB[275]), .B(DB[260]), .Z(n1978) );
  AND U3776 ( .A(n442), .B(n1979), .Z(n1977) );
  XOR U3777 ( .A(n1980), .B(n1981), .Z(n1979) );
  XOR U3778 ( .A(DB[260]), .B(DB[245]), .Z(n1981) );
  AND U3779 ( .A(n446), .B(n1982), .Z(n1980) );
  XOR U3780 ( .A(n1983), .B(n1984), .Z(n1982) );
  XOR U3781 ( .A(DB[245]), .B(DB[230]), .Z(n1984) );
  AND U3782 ( .A(n450), .B(n1985), .Z(n1983) );
  XOR U3783 ( .A(n1986), .B(n1987), .Z(n1985) );
  XOR U3784 ( .A(DB[230]), .B(DB[215]), .Z(n1987) );
  AND U3785 ( .A(n454), .B(n1988), .Z(n1986) );
  XOR U3786 ( .A(n1989), .B(n1990), .Z(n1988) );
  XOR U3787 ( .A(DB[215]), .B(DB[200]), .Z(n1990) );
  AND U3788 ( .A(n458), .B(n1991), .Z(n1989) );
  XOR U3789 ( .A(n1992), .B(n1993), .Z(n1991) );
  XOR U3790 ( .A(DB[200]), .B(DB[185]), .Z(n1993) );
  AND U3791 ( .A(n462), .B(n1994), .Z(n1992) );
  XOR U3792 ( .A(n1995), .B(n1996), .Z(n1994) );
  XOR U3793 ( .A(DB[185]), .B(DB[170]), .Z(n1996) );
  AND U3794 ( .A(n466), .B(n1997), .Z(n1995) );
  XOR U3795 ( .A(n1998), .B(n1999), .Z(n1997) );
  XOR U3796 ( .A(DB[170]), .B(DB[155]), .Z(n1999) );
  AND U3797 ( .A(n470), .B(n2000), .Z(n1998) );
  XOR U3798 ( .A(n2001), .B(n2002), .Z(n2000) );
  XOR U3799 ( .A(DB[155]), .B(DB[140]), .Z(n2002) );
  AND U3800 ( .A(n474), .B(n2003), .Z(n2001) );
  XOR U3801 ( .A(n2004), .B(n2005), .Z(n2003) );
  XOR U3802 ( .A(DB[140]), .B(DB[125]), .Z(n2005) );
  AND U3803 ( .A(n478), .B(n2006), .Z(n2004) );
  XOR U3804 ( .A(n2007), .B(n2008), .Z(n2006) );
  XOR U3805 ( .A(DB[125]), .B(DB[110]), .Z(n2008) );
  AND U3806 ( .A(n482), .B(n2009), .Z(n2007) );
  XOR U3807 ( .A(n2010), .B(n2011), .Z(n2009) );
  XOR U3808 ( .A(DB[95]), .B(DB[110]), .Z(n2011) );
  AND U3809 ( .A(n486), .B(n2012), .Z(n2010) );
  XOR U3810 ( .A(n2013), .B(n2014), .Z(n2012) );
  XOR U3811 ( .A(DB[95]), .B(DB[80]), .Z(n2014) );
  AND U3812 ( .A(n490), .B(n2015), .Z(n2013) );
  XOR U3813 ( .A(n2016), .B(n2017), .Z(n2015) );
  XOR U3814 ( .A(DB[80]), .B(DB[65]), .Z(n2017) );
  AND U3815 ( .A(n494), .B(n2018), .Z(n2016) );
  XOR U3816 ( .A(n2019), .B(n2020), .Z(n2018) );
  XOR U3817 ( .A(DB[65]), .B(DB[50]), .Z(n2020) );
  AND U3818 ( .A(n498), .B(n2021), .Z(n2019) );
  XOR U3819 ( .A(n2022), .B(n2023), .Z(n2021) );
  XOR U3820 ( .A(DB[50]), .B(DB[35]), .Z(n2023) );
  AND U3821 ( .A(n502), .B(n2024), .Z(n2022) );
  XOR U3822 ( .A(n2025), .B(n2026), .Z(n2024) );
  XOR U3823 ( .A(DB[35]), .B(DB[20]), .Z(n2026) );
  AND U3824 ( .A(n506), .B(n2027), .Z(n2025) );
  XOR U3825 ( .A(DB[5]), .B(DB[20]), .Z(n2027) );
  XOR U3826 ( .A(DB[1909]), .B(n2028), .Z(min_val_out[4]) );
  AND U3827 ( .A(n2), .B(n2029), .Z(n2028) );
  XOR U3828 ( .A(n2030), .B(n2031), .Z(n2029) );
  XOR U3829 ( .A(DB[1909]), .B(DB[1894]), .Z(n2031) );
  AND U3830 ( .A(n6), .B(n2032), .Z(n2030) );
  XOR U3831 ( .A(n2033), .B(n2034), .Z(n2032) );
  XOR U3832 ( .A(DB[1894]), .B(DB[1879]), .Z(n2034) );
  AND U3833 ( .A(n10), .B(n2035), .Z(n2033) );
  XOR U3834 ( .A(n2036), .B(n2037), .Z(n2035) );
  XOR U3835 ( .A(DB[1879]), .B(DB[1864]), .Z(n2037) );
  AND U3836 ( .A(n14), .B(n2038), .Z(n2036) );
  XOR U3837 ( .A(n2039), .B(n2040), .Z(n2038) );
  XOR U3838 ( .A(DB[1864]), .B(DB[1849]), .Z(n2040) );
  AND U3839 ( .A(n18), .B(n2041), .Z(n2039) );
  XOR U3840 ( .A(n2042), .B(n2043), .Z(n2041) );
  XOR U3841 ( .A(DB[1849]), .B(DB[1834]), .Z(n2043) );
  AND U3842 ( .A(n22), .B(n2044), .Z(n2042) );
  XOR U3843 ( .A(n2045), .B(n2046), .Z(n2044) );
  XOR U3844 ( .A(DB[1834]), .B(DB[1819]), .Z(n2046) );
  AND U3845 ( .A(n26), .B(n2047), .Z(n2045) );
  XOR U3846 ( .A(n2048), .B(n2049), .Z(n2047) );
  XOR U3847 ( .A(DB[1819]), .B(DB[1804]), .Z(n2049) );
  AND U3848 ( .A(n30), .B(n2050), .Z(n2048) );
  XOR U3849 ( .A(n2051), .B(n2052), .Z(n2050) );
  XOR U3850 ( .A(DB[1804]), .B(DB[1789]), .Z(n2052) );
  AND U3851 ( .A(n34), .B(n2053), .Z(n2051) );
  XOR U3852 ( .A(n2054), .B(n2055), .Z(n2053) );
  XOR U3853 ( .A(DB[1789]), .B(DB[1774]), .Z(n2055) );
  AND U3854 ( .A(n38), .B(n2056), .Z(n2054) );
  XOR U3855 ( .A(n2057), .B(n2058), .Z(n2056) );
  XOR U3856 ( .A(DB[1774]), .B(DB[1759]), .Z(n2058) );
  AND U3857 ( .A(n42), .B(n2059), .Z(n2057) );
  XOR U3858 ( .A(n2060), .B(n2061), .Z(n2059) );
  XOR U3859 ( .A(DB[1759]), .B(DB[1744]), .Z(n2061) );
  AND U3860 ( .A(n46), .B(n2062), .Z(n2060) );
  XOR U3861 ( .A(n2063), .B(n2064), .Z(n2062) );
  XOR U3862 ( .A(DB[1744]), .B(DB[1729]), .Z(n2064) );
  AND U3863 ( .A(n50), .B(n2065), .Z(n2063) );
  XOR U3864 ( .A(n2066), .B(n2067), .Z(n2065) );
  XOR U3865 ( .A(DB[1729]), .B(DB[1714]), .Z(n2067) );
  AND U3866 ( .A(n54), .B(n2068), .Z(n2066) );
  XOR U3867 ( .A(n2069), .B(n2070), .Z(n2068) );
  XOR U3868 ( .A(DB[1714]), .B(DB[1699]), .Z(n2070) );
  AND U3869 ( .A(n58), .B(n2071), .Z(n2069) );
  XOR U3870 ( .A(n2072), .B(n2073), .Z(n2071) );
  XOR U3871 ( .A(DB[1699]), .B(DB[1684]), .Z(n2073) );
  AND U3872 ( .A(n62), .B(n2074), .Z(n2072) );
  XOR U3873 ( .A(n2075), .B(n2076), .Z(n2074) );
  XOR U3874 ( .A(DB[1684]), .B(DB[1669]), .Z(n2076) );
  AND U3875 ( .A(n66), .B(n2077), .Z(n2075) );
  XOR U3876 ( .A(n2078), .B(n2079), .Z(n2077) );
  XOR U3877 ( .A(DB[1669]), .B(DB[1654]), .Z(n2079) );
  AND U3878 ( .A(n70), .B(n2080), .Z(n2078) );
  XOR U3879 ( .A(n2081), .B(n2082), .Z(n2080) );
  XOR U3880 ( .A(DB[1654]), .B(DB[1639]), .Z(n2082) );
  AND U3881 ( .A(n74), .B(n2083), .Z(n2081) );
  XOR U3882 ( .A(n2084), .B(n2085), .Z(n2083) );
  XOR U3883 ( .A(DB[1639]), .B(DB[1624]), .Z(n2085) );
  AND U3884 ( .A(n78), .B(n2086), .Z(n2084) );
  XOR U3885 ( .A(n2087), .B(n2088), .Z(n2086) );
  XOR U3886 ( .A(DB[1624]), .B(DB[1609]), .Z(n2088) );
  AND U3887 ( .A(n82), .B(n2089), .Z(n2087) );
  XOR U3888 ( .A(n2090), .B(n2091), .Z(n2089) );
  XOR U3889 ( .A(DB[1609]), .B(DB[1594]), .Z(n2091) );
  AND U3890 ( .A(n86), .B(n2092), .Z(n2090) );
  XOR U3891 ( .A(n2093), .B(n2094), .Z(n2092) );
  XOR U3892 ( .A(DB[1594]), .B(DB[1579]), .Z(n2094) );
  AND U3893 ( .A(n90), .B(n2095), .Z(n2093) );
  XOR U3894 ( .A(n2096), .B(n2097), .Z(n2095) );
  XOR U3895 ( .A(DB[1579]), .B(DB[1564]), .Z(n2097) );
  AND U3896 ( .A(n94), .B(n2098), .Z(n2096) );
  XOR U3897 ( .A(n2099), .B(n2100), .Z(n2098) );
  XOR U3898 ( .A(DB[1564]), .B(DB[1549]), .Z(n2100) );
  AND U3899 ( .A(n98), .B(n2101), .Z(n2099) );
  XOR U3900 ( .A(n2102), .B(n2103), .Z(n2101) );
  XOR U3901 ( .A(DB[1549]), .B(DB[1534]), .Z(n2103) );
  AND U3902 ( .A(n102), .B(n2104), .Z(n2102) );
  XOR U3903 ( .A(n2105), .B(n2106), .Z(n2104) );
  XOR U3904 ( .A(DB[1534]), .B(DB[1519]), .Z(n2106) );
  AND U3905 ( .A(n106), .B(n2107), .Z(n2105) );
  XOR U3906 ( .A(n2108), .B(n2109), .Z(n2107) );
  XOR U3907 ( .A(DB[1519]), .B(DB[1504]), .Z(n2109) );
  AND U3908 ( .A(n110), .B(n2110), .Z(n2108) );
  XOR U3909 ( .A(n2111), .B(n2112), .Z(n2110) );
  XOR U3910 ( .A(DB[1504]), .B(DB[1489]), .Z(n2112) );
  AND U3911 ( .A(n114), .B(n2113), .Z(n2111) );
  XOR U3912 ( .A(n2114), .B(n2115), .Z(n2113) );
  XOR U3913 ( .A(DB[1489]), .B(DB[1474]), .Z(n2115) );
  AND U3914 ( .A(n118), .B(n2116), .Z(n2114) );
  XOR U3915 ( .A(n2117), .B(n2118), .Z(n2116) );
  XOR U3916 ( .A(DB[1474]), .B(DB[1459]), .Z(n2118) );
  AND U3917 ( .A(n122), .B(n2119), .Z(n2117) );
  XOR U3918 ( .A(n2120), .B(n2121), .Z(n2119) );
  XOR U3919 ( .A(DB[1459]), .B(DB[1444]), .Z(n2121) );
  AND U3920 ( .A(n126), .B(n2122), .Z(n2120) );
  XOR U3921 ( .A(n2123), .B(n2124), .Z(n2122) );
  XOR U3922 ( .A(DB[1444]), .B(DB[1429]), .Z(n2124) );
  AND U3923 ( .A(n130), .B(n2125), .Z(n2123) );
  XOR U3924 ( .A(n2126), .B(n2127), .Z(n2125) );
  XOR U3925 ( .A(DB[1429]), .B(DB[1414]), .Z(n2127) );
  AND U3926 ( .A(n134), .B(n2128), .Z(n2126) );
  XOR U3927 ( .A(n2129), .B(n2130), .Z(n2128) );
  XOR U3928 ( .A(DB[1414]), .B(DB[1399]), .Z(n2130) );
  AND U3929 ( .A(n138), .B(n2131), .Z(n2129) );
  XOR U3930 ( .A(n2132), .B(n2133), .Z(n2131) );
  XOR U3931 ( .A(DB[1399]), .B(DB[1384]), .Z(n2133) );
  AND U3932 ( .A(n142), .B(n2134), .Z(n2132) );
  XOR U3933 ( .A(n2135), .B(n2136), .Z(n2134) );
  XOR U3934 ( .A(DB[1384]), .B(DB[1369]), .Z(n2136) );
  AND U3935 ( .A(n146), .B(n2137), .Z(n2135) );
  XOR U3936 ( .A(n2138), .B(n2139), .Z(n2137) );
  XOR U3937 ( .A(DB[1369]), .B(DB[1354]), .Z(n2139) );
  AND U3938 ( .A(n150), .B(n2140), .Z(n2138) );
  XOR U3939 ( .A(n2141), .B(n2142), .Z(n2140) );
  XOR U3940 ( .A(DB[1354]), .B(DB[1339]), .Z(n2142) );
  AND U3941 ( .A(n154), .B(n2143), .Z(n2141) );
  XOR U3942 ( .A(n2144), .B(n2145), .Z(n2143) );
  XOR U3943 ( .A(DB[1339]), .B(DB[1324]), .Z(n2145) );
  AND U3944 ( .A(n158), .B(n2146), .Z(n2144) );
  XOR U3945 ( .A(n2147), .B(n2148), .Z(n2146) );
  XOR U3946 ( .A(DB[1324]), .B(DB[1309]), .Z(n2148) );
  AND U3947 ( .A(n162), .B(n2149), .Z(n2147) );
  XOR U3948 ( .A(n2150), .B(n2151), .Z(n2149) );
  XOR U3949 ( .A(DB[1309]), .B(DB[1294]), .Z(n2151) );
  AND U3950 ( .A(n166), .B(n2152), .Z(n2150) );
  XOR U3951 ( .A(n2153), .B(n2154), .Z(n2152) );
  XOR U3952 ( .A(DB[1294]), .B(DB[1279]), .Z(n2154) );
  AND U3953 ( .A(n170), .B(n2155), .Z(n2153) );
  XOR U3954 ( .A(n2156), .B(n2157), .Z(n2155) );
  XOR U3955 ( .A(DB[1279]), .B(DB[1264]), .Z(n2157) );
  AND U3956 ( .A(n174), .B(n2158), .Z(n2156) );
  XOR U3957 ( .A(n2159), .B(n2160), .Z(n2158) );
  XOR U3958 ( .A(DB[1264]), .B(DB[1249]), .Z(n2160) );
  AND U3959 ( .A(n178), .B(n2161), .Z(n2159) );
  XOR U3960 ( .A(n2162), .B(n2163), .Z(n2161) );
  XOR U3961 ( .A(DB[1249]), .B(DB[1234]), .Z(n2163) );
  AND U3962 ( .A(n182), .B(n2164), .Z(n2162) );
  XOR U3963 ( .A(n2165), .B(n2166), .Z(n2164) );
  XOR U3964 ( .A(DB[1234]), .B(DB[1219]), .Z(n2166) );
  AND U3965 ( .A(n186), .B(n2167), .Z(n2165) );
  XOR U3966 ( .A(n2168), .B(n2169), .Z(n2167) );
  XOR U3967 ( .A(DB[1219]), .B(DB[1204]), .Z(n2169) );
  AND U3968 ( .A(n190), .B(n2170), .Z(n2168) );
  XOR U3969 ( .A(n2171), .B(n2172), .Z(n2170) );
  XOR U3970 ( .A(DB[1204]), .B(DB[1189]), .Z(n2172) );
  AND U3971 ( .A(n194), .B(n2173), .Z(n2171) );
  XOR U3972 ( .A(n2174), .B(n2175), .Z(n2173) );
  XOR U3973 ( .A(DB[1189]), .B(DB[1174]), .Z(n2175) );
  AND U3974 ( .A(n198), .B(n2176), .Z(n2174) );
  XOR U3975 ( .A(n2177), .B(n2178), .Z(n2176) );
  XOR U3976 ( .A(DB[1174]), .B(DB[1159]), .Z(n2178) );
  AND U3977 ( .A(n202), .B(n2179), .Z(n2177) );
  XOR U3978 ( .A(n2180), .B(n2181), .Z(n2179) );
  XOR U3979 ( .A(DB[1159]), .B(DB[1144]), .Z(n2181) );
  AND U3980 ( .A(n206), .B(n2182), .Z(n2180) );
  XOR U3981 ( .A(n2183), .B(n2184), .Z(n2182) );
  XOR U3982 ( .A(DB[1144]), .B(DB[1129]), .Z(n2184) );
  AND U3983 ( .A(n210), .B(n2185), .Z(n2183) );
  XOR U3984 ( .A(n2186), .B(n2187), .Z(n2185) );
  XOR U3985 ( .A(DB[1129]), .B(DB[1114]), .Z(n2187) );
  AND U3986 ( .A(n214), .B(n2188), .Z(n2186) );
  XOR U3987 ( .A(n2189), .B(n2190), .Z(n2188) );
  XOR U3988 ( .A(DB[1114]), .B(DB[1099]), .Z(n2190) );
  AND U3989 ( .A(n218), .B(n2191), .Z(n2189) );
  XOR U3990 ( .A(n2192), .B(n2193), .Z(n2191) );
  XOR U3991 ( .A(DB[1099]), .B(DB[1084]), .Z(n2193) );
  AND U3992 ( .A(n222), .B(n2194), .Z(n2192) );
  XOR U3993 ( .A(n2195), .B(n2196), .Z(n2194) );
  XOR U3994 ( .A(DB[1084]), .B(DB[1069]), .Z(n2196) );
  AND U3995 ( .A(n226), .B(n2197), .Z(n2195) );
  XOR U3996 ( .A(n2198), .B(n2199), .Z(n2197) );
  XOR U3997 ( .A(DB[1069]), .B(DB[1054]), .Z(n2199) );
  AND U3998 ( .A(n230), .B(n2200), .Z(n2198) );
  XOR U3999 ( .A(n2201), .B(n2202), .Z(n2200) );
  XOR U4000 ( .A(DB[1054]), .B(DB[1039]), .Z(n2202) );
  AND U4001 ( .A(n234), .B(n2203), .Z(n2201) );
  XOR U4002 ( .A(n2204), .B(n2205), .Z(n2203) );
  XOR U4003 ( .A(DB[1039]), .B(DB[1024]), .Z(n2205) );
  AND U4004 ( .A(n238), .B(n2206), .Z(n2204) );
  XOR U4005 ( .A(n2207), .B(n2208), .Z(n2206) );
  XOR U4006 ( .A(DB[1024]), .B(DB[1009]), .Z(n2208) );
  AND U4007 ( .A(n242), .B(n2209), .Z(n2207) );
  XOR U4008 ( .A(n2210), .B(n2211), .Z(n2209) );
  XOR U4009 ( .A(DB[994]), .B(DB[1009]), .Z(n2211) );
  AND U4010 ( .A(n246), .B(n2212), .Z(n2210) );
  XOR U4011 ( .A(n2213), .B(n2214), .Z(n2212) );
  XOR U4012 ( .A(DB[994]), .B(DB[979]), .Z(n2214) );
  AND U4013 ( .A(n250), .B(n2215), .Z(n2213) );
  XOR U4014 ( .A(n2216), .B(n2217), .Z(n2215) );
  XOR U4015 ( .A(DB[979]), .B(DB[964]), .Z(n2217) );
  AND U4016 ( .A(n254), .B(n2218), .Z(n2216) );
  XOR U4017 ( .A(n2219), .B(n2220), .Z(n2218) );
  XOR U4018 ( .A(DB[964]), .B(DB[949]), .Z(n2220) );
  AND U4019 ( .A(n258), .B(n2221), .Z(n2219) );
  XOR U4020 ( .A(n2222), .B(n2223), .Z(n2221) );
  XOR U4021 ( .A(DB[949]), .B(DB[934]), .Z(n2223) );
  AND U4022 ( .A(n262), .B(n2224), .Z(n2222) );
  XOR U4023 ( .A(n2225), .B(n2226), .Z(n2224) );
  XOR U4024 ( .A(DB[934]), .B(DB[919]), .Z(n2226) );
  AND U4025 ( .A(n266), .B(n2227), .Z(n2225) );
  XOR U4026 ( .A(n2228), .B(n2229), .Z(n2227) );
  XOR U4027 ( .A(DB[919]), .B(DB[904]), .Z(n2229) );
  AND U4028 ( .A(n270), .B(n2230), .Z(n2228) );
  XOR U4029 ( .A(n2231), .B(n2232), .Z(n2230) );
  XOR U4030 ( .A(DB[904]), .B(DB[889]), .Z(n2232) );
  AND U4031 ( .A(n274), .B(n2233), .Z(n2231) );
  XOR U4032 ( .A(n2234), .B(n2235), .Z(n2233) );
  XOR U4033 ( .A(DB[889]), .B(DB[874]), .Z(n2235) );
  AND U4034 ( .A(n278), .B(n2236), .Z(n2234) );
  XOR U4035 ( .A(n2237), .B(n2238), .Z(n2236) );
  XOR U4036 ( .A(DB[874]), .B(DB[859]), .Z(n2238) );
  AND U4037 ( .A(n282), .B(n2239), .Z(n2237) );
  XOR U4038 ( .A(n2240), .B(n2241), .Z(n2239) );
  XOR U4039 ( .A(DB[859]), .B(DB[844]), .Z(n2241) );
  AND U4040 ( .A(n286), .B(n2242), .Z(n2240) );
  XOR U4041 ( .A(n2243), .B(n2244), .Z(n2242) );
  XOR U4042 ( .A(DB[844]), .B(DB[829]), .Z(n2244) );
  AND U4043 ( .A(n290), .B(n2245), .Z(n2243) );
  XOR U4044 ( .A(n2246), .B(n2247), .Z(n2245) );
  XOR U4045 ( .A(DB[829]), .B(DB[814]), .Z(n2247) );
  AND U4046 ( .A(n294), .B(n2248), .Z(n2246) );
  XOR U4047 ( .A(n2249), .B(n2250), .Z(n2248) );
  XOR U4048 ( .A(DB[814]), .B(DB[799]), .Z(n2250) );
  AND U4049 ( .A(n298), .B(n2251), .Z(n2249) );
  XOR U4050 ( .A(n2252), .B(n2253), .Z(n2251) );
  XOR U4051 ( .A(DB[799]), .B(DB[784]), .Z(n2253) );
  AND U4052 ( .A(n302), .B(n2254), .Z(n2252) );
  XOR U4053 ( .A(n2255), .B(n2256), .Z(n2254) );
  XOR U4054 ( .A(DB[784]), .B(DB[769]), .Z(n2256) );
  AND U4055 ( .A(n306), .B(n2257), .Z(n2255) );
  XOR U4056 ( .A(n2258), .B(n2259), .Z(n2257) );
  XOR U4057 ( .A(DB[769]), .B(DB[754]), .Z(n2259) );
  AND U4058 ( .A(n310), .B(n2260), .Z(n2258) );
  XOR U4059 ( .A(n2261), .B(n2262), .Z(n2260) );
  XOR U4060 ( .A(DB[754]), .B(DB[739]), .Z(n2262) );
  AND U4061 ( .A(n314), .B(n2263), .Z(n2261) );
  XOR U4062 ( .A(n2264), .B(n2265), .Z(n2263) );
  XOR U4063 ( .A(DB[739]), .B(DB[724]), .Z(n2265) );
  AND U4064 ( .A(n318), .B(n2266), .Z(n2264) );
  XOR U4065 ( .A(n2267), .B(n2268), .Z(n2266) );
  XOR U4066 ( .A(DB[724]), .B(DB[709]), .Z(n2268) );
  AND U4067 ( .A(n322), .B(n2269), .Z(n2267) );
  XOR U4068 ( .A(n2270), .B(n2271), .Z(n2269) );
  XOR U4069 ( .A(DB[709]), .B(DB[694]), .Z(n2271) );
  AND U4070 ( .A(n326), .B(n2272), .Z(n2270) );
  XOR U4071 ( .A(n2273), .B(n2274), .Z(n2272) );
  XOR U4072 ( .A(DB[694]), .B(DB[679]), .Z(n2274) );
  AND U4073 ( .A(n330), .B(n2275), .Z(n2273) );
  XOR U4074 ( .A(n2276), .B(n2277), .Z(n2275) );
  XOR U4075 ( .A(DB[679]), .B(DB[664]), .Z(n2277) );
  AND U4076 ( .A(n334), .B(n2278), .Z(n2276) );
  XOR U4077 ( .A(n2279), .B(n2280), .Z(n2278) );
  XOR U4078 ( .A(DB[664]), .B(DB[649]), .Z(n2280) );
  AND U4079 ( .A(n338), .B(n2281), .Z(n2279) );
  XOR U4080 ( .A(n2282), .B(n2283), .Z(n2281) );
  XOR U4081 ( .A(DB[649]), .B(DB[634]), .Z(n2283) );
  AND U4082 ( .A(n342), .B(n2284), .Z(n2282) );
  XOR U4083 ( .A(n2285), .B(n2286), .Z(n2284) );
  XOR U4084 ( .A(DB[634]), .B(DB[619]), .Z(n2286) );
  AND U4085 ( .A(n346), .B(n2287), .Z(n2285) );
  XOR U4086 ( .A(n2288), .B(n2289), .Z(n2287) );
  XOR U4087 ( .A(DB[619]), .B(DB[604]), .Z(n2289) );
  AND U4088 ( .A(n350), .B(n2290), .Z(n2288) );
  XOR U4089 ( .A(n2291), .B(n2292), .Z(n2290) );
  XOR U4090 ( .A(DB[604]), .B(DB[589]), .Z(n2292) );
  AND U4091 ( .A(n354), .B(n2293), .Z(n2291) );
  XOR U4092 ( .A(n2294), .B(n2295), .Z(n2293) );
  XOR U4093 ( .A(DB[589]), .B(DB[574]), .Z(n2295) );
  AND U4094 ( .A(n358), .B(n2296), .Z(n2294) );
  XOR U4095 ( .A(n2297), .B(n2298), .Z(n2296) );
  XOR U4096 ( .A(DB[574]), .B(DB[559]), .Z(n2298) );
  AND U4097 ( .A(n362), .B(n2299), .Z(n2297) );
  XOR U4098 ( .A(n2300), .B(n2301), .Z(n2299) );
  XOR U4099 ( .A(DB[559]), .B(DB[544]), .Z(n2301) );
  AND U4100 ( .A(n366), .B(n2302), .Z(n2300) );
  XOR U4101 ( .A(n2303), .B(n2304), .Z(n2302) );
  XOR U4102 ( .A(DB[544]), .B(DB[529]), .Z(n2304) );
  AND U4103 ( .A(n370), .B(n2305), .Z(n2303) );
  XOR U4104 ( .A(n2306), .B(n2307), .Z(n2305) );
  XOR U4105 ( .A(DB[529]), .B(DB[514]), .Z(n2307) );
  AND U4106 ( .A(n374), .B(n2308), .Z(n2306) );
  XOR U4107 ( .A(n2309), .B(n2310), .Z(n2308) );
  XOR U4108 ( .A(DB[514]), .B(DB[499]), .Z(n2310) );
  AND U4109 ( .A(n378), .B(n2311), .Z(n2309) );
  XOR U4110 ( .A(n2312), .B(n2313), .Z(n2311) );
  XOR U4111 ( .A(DB[499]), .B(DB[484]), .Z(n2313) );
  AND U4112 ( .A(n382), .B(n2314), .Z(n2312) );
  XOR U4113 ( .A(n2315), .B(n2316), .Z(n2314) );
  XOR U4114 ( .A(DB[484]), .B(DB[469]), .Z(n2316) );
  AND U4115 ( .A(n386), .B(n2317), .Z(n2315) );
  XOR U4116 ( .A(n2318), .B(n2319), .Z(n2317) );
  XOR U4117 ( .A(DB[469]), .B(DB[454]), .Z(n2319) );
  AND U4118 ( .A(n390), .B(n2320), .Z(n2318) );
  XOR U4119 ( .A(n2321), .B(n2322), .Z(n2320) );
  XOR U4120 ( .A(DB[454]), .B(DB[439]), .Z(n2322) );
  AND U4121 ( .A(n394), .B(n2323), .Z(n2321) );
  XOR U4122 ( .A(n2324), .B(n2325), .Z(n2323) );
  XOR U4123 ( .A(DB[439]), .B(DB[424]), .Z(n2325) );
  AND U4124 ( .A(n398), .B(n2326), .Z(n2324) );
  XOR U4125 ( .A(n2327), .B(n2328), .Z(n2326) );
  XOR U4126 ( .A(DB[424]), .B(DB[409]), .Z(n2328) );
  AND U4127 ( .A(n402), .B(n2329), .Z(n2327) );
  XOR U4128 ( .A(n2330), .B(n2331), .Z(n2329) );
  XOR U4129 ( .A(DB[409]), .B(DB[394]), .Z(n2331) );
  AND U4130 ( .A(n406), .B(n2332), .Z(n2330) );
  XOR U4131 ( .A(n2333), .B(n2334), .Z(n2332) );
  XOR U4132 ( .A(DB[394]), .B(DB[379]), .Z(n2334) );
  AND U4133 ( .A(n410), .B(n2335), .Z(n2333) );
  XOR U4134 ( .A(n2336), .B(n2337), .Z(n2335) );
  XOR U4135 ( .A(DB[379]), .B(DB[364]), .Z(n2337) );
  AND U4136 ( .A(n414), .B(n2338), .Z(n2336) );
  XOR U4137 ( .A(n2339), .B(n2340), .Z(n2338) );
  XOR U4138 ( .A(DB[364]), .B(DB[349]), .Z(n2340) );
  AND U4139 ( .A(n418), .B(n2341), .Z(n2339) );
  XOR U4140 ( .A(n2342), .B(n2343), .Z(n2341) );
  XOR U4141 ( .A(DB[349]), .B(DB[334]), .Z(n2343) );
  AND U4142 ( .A(n422), .B(n2344), .Z(n2342) );
  XOR U4143 ( .A(n2345), .B(n2346), .Z(n2344) );
  XOR U4144 ( .A(DB[334]), .B(DB[319]), .Z(n2346) );
  AND U4145 ( .A(n426), .B(n2347), .Z(n2345) );
  XOR U4146 ( .A(n2348), .B(n2349), .Z(n2347) );
  XOR U4147 ( .A(DB[319]), .B(DB[304]), .Z(n2349) );
  AND U4148 ( .A(n430), .B(n2350), .Z(n2348) );
  XOR U4149 ( .A(n2351), .B(n2352), .Z(n2350) );
  XOR U4150 ( .A(DB[304]), .B(DB[289]), .Z(n2352) );
  AND U4151 ( .A(n434), .B(n2353), .Z(n2351) );
  XOR U4152 ( .A(n2354), .B(n2355), .Z(n2353) );
  XOR U4153 ( .A(DB[289]), .B(DB[274]), .Z(n2355) );
  AND U4154 ( .A(n438), .B(n2356), .Z(n2354) );
  XOR U4155 ( .A(n2357), .B(n2358), .Z(n2356) );
  XOR U4156 ( .A(DB[274]), .B(DB[259]), .Z(n2358) );
  AND U4157 ( .A(n442), .B(n2359), .Z(n2357) );
  XOR U4158 ( .A(n2360), .B(n2361), .Z(n2359) );
  XOR U4159 ( .A(DB[259]), .B(DB[244]), .Z(n2361) );
  AND U4160 ( .A(n446), .B(n2362), .Z(n2360) );
  XOR U4161 ( .A(n2363), .B(n2364), .Z(n2362) );
  XOR U4162 ( .A(DB[244]), .B(DB[229]), .Z(n2364) );
  AND U4163 ( .A(n450), .B(n2365), .Z(n2363) );
  XOR U4164 ( .A(n2366), .B(n2367), .Z(n2365) );
  XOR U4165 ( .A(DB[229]), .B(DB[214]), .Z(n2367) );
  AND U4166 ( .A(n454), .B(n2368), .Z(n2366) );
  XOR U4167 ( .A(n2369), .B(n2370), .Z(n2368) );
  XOR U4168 ( .A(DB[214]), .B(DB[199]), .Z(n2370) );
  AND U4169 ( .A(n458), .B(n2371), .Z(n2369) );
  XOR U4170 ( .A(n2372), .B(n2373), .Z(n2371) );
  XOR U4171 ( .A(DB[199]), .B(DB[184]), .Z(n2373) );
  AND U4172 ( .A(n462), .B(n2374), .Z(n2372) );
  XOR U4173 ( .A(n2375), .B(n2376), .Z(n2374) );
  XOR U4174 ( .A(DB[184]), .B(DB[169]), .Z(n2376) );
  AND U4175 ( .A(n466), .B(n2377), .Z(n2375) );
  XOR U4176 ( .A(n2378), .B(n2379), .Z(n2377) );
  XOR U4177 ( .A(DB[169]), .B(DB[154]), .Z(n2379) );
  AND U4178 ( .A(n470), .B(n2380), .Z(n2378) );
  XOR U4179 ( .A(n2381), .B(n2382), .Z(n2380) );
  XOR U4180 ( .A(DB[154]), .B(DB[139]), .Z(n2382) );
  AND U4181 ( .A(n474), .B(n2383), .Z(n2381) );
  XOR U4182 ( .A(n2384), .B(n2385), .Z(n2383) );
  XOR U4183 ( .A(DB[139]), .B(DB[124]), .Z(n2385) );
  AND U4184 ( .A(n478), .B(n2386), .Z(n2384) );
  XOR U4185 ( .A(n2387), .B(n2388), .Z(n2386) );
  XOR U4186 ( .A(DB[124]), .B(DB[109]), .Z(n2388) );
  AND U4187 ( .A(n482), .B(n2389), .Z(n2387) );
  XOR U4188 ( .A(n2390), .B(n2391), .Z(n2389) );
  XOR U4189 ( .A(DB[94]), .B(DB[109]), .Z(n2391) );
  AND U4190 ( .A(n486), .B(n2392), .Z(n2390) );
  XOR U4191 ( .A(n2393), .B(n2394), .Z(n2392) );
  XOR U4192 ( .A(DB[94]), .B(DB[79]), .Z(n2394) );
  AND U4193 ( .A(n490), .B(n2395), .Z(n2393) );
  XOR U4194 ( .A(n2396), .B(n2397), .Z(n2395) );
  XOR U4195 ( .A(DB[79]), .B(DB[64]), .Z(n2397) );
  AND U4196 ( .A(n494), .B(n2398), .Z(n2396) );
  XOR U4197 ( .A(n2399), .B(n2400), .Z(n2398) );
  XOR U4198 ( .A(DB[64]), .B(DB[49]), .Z(n2400) );
  AND U4199 ( .A(n498), .B(n2401), .Z(n2399) );
  XOR U4200 ( .A(n2402), .B(n2403), .Z(n2401) );
  XOR U4201 ( .A(DB[49]), .B(DB[34]), .Z(n2403) );
  AND U4202 ( .A(n502), .B(n2404), .Z(n2402) );
  XOR U4203 ( .A(n2405), .B(n2406), .Z(n2404) );
  XOR U4204 ( .A(DB[34]), .B(DB[19]), .Z(n2406) );
  AND U4205 ( .A(n506), .B(n2407), .Z(n2405) );
  XOR U4206 ( .A(DB[4]), .B(DB[19]), .Z(n2407) );
  XOR U4207 ( .A(DB[1908]), .B(n2408), .Z(min_val_out[3]) );
  AND U4208 ( .A(n2), .B(n2409), .Z(n2408) );
  XOR U4209 ( .A(n2410), .B(n2411), .Z(n2409) );
  XOR U4210 ( .A(DB[1908]), .B(DB[1893]), .Z(n2411) );
  AND U4211 ( .A(n6), .B(n2412), .Z(n2410) );
  XOR U4212 ( .A(n2413), .B(n2414), .Z(n2412) );
  XOR U4213 ( .A(DB[1893]), .B(DB[1878]), .Z(n2414) );
  AND U4214 ( .A(n10), .B(n2415), .Z(n2413) );
  XOR U4215 ( .A(n2416), .B(n2417), .Z(n2415) );
  XOR U4216 ( .A(DB[1878]), .B(DB[1863]), .Z(n2417) );
  AND U4217 ( .A(n14), .B(n2418), .Z(n2416) );
  XOR U4218 ( .A(n2419), .B(n2420), .Z(n2418) );
  XOR U4219 ( .A(DB[1863]), .B(DB[1848]), .Z(n2420) );
  AND U4220 ( .A(n18), .B(n2421), .Z(n2419) );
  XOR U4221 ( .A(n2422), .B(n2423), .Z(n2421) );
  XOR U4222 ( .A(DB[1848]), .B(DB[1833]), .Z(n2423) );
  AND U4223 ( .A(n22), .B(n2424), .Z(n2422) );
  XOR U4224 ( .A(n2425), .B(n2426), .Z(n2424) );
  XOR U4225 ( .A(DB[1833]), .B(DB[1818]), .Z(n2426) );
  AND U4226 ( .A(n26), .B(n2427), .Z(n2425) );
  XOR U4227 ( .A(n2428), .B(n2429), .Z(n2427) );
  XOR U4228 ( .A(DB[1818]), .B(DB[1803]), .Z(n2429) );
  AND U4229 ( .A(n30), .B(n2430), .Z(n2428) );
  XOR U4230 ( .A(n2431), .B(n2432), .Z(n2430) );
  XOR U4231 ( .A(DB[1803]), .B(DB[1788]), .Z(n2432) );
  AND U4232 ( .A(n34), .B(n2433), .Z(n2431) );
  XOR U4233 ( .A(n2434), .B(n2435), .Z(n2433) );
  XOR U4234 ( .A(DB[1788]), .B(DB[1773]), .Z(n2435) );
  AND U4235 ( .A(n38), .B(n2436), .Z(n2434) );
  XOR U4236 ( .A(n2437), .B(n2438), .Z(n2436) );
  XOR U4237 ( .A(DB[1773]), .B(DB[1758]), .Z(n2438) );
  AND U4238 ( .A(n42), .B(n2439), .Z(n2437) );
  XOR U4239 ( .A(n2440), .B(n2441), .Z(n2439) );
  XOR U4240 ( .A(DB[1758]), .B(DB[1743]), .Z(n2441) );
  AND U4241 ( .A(n46), .B(n2442), .Z(n2440) );
  XOR U4242 ( .A(n2443), .B(n2444), .Z(n2442) );
  XOR U4243 ( .A(DB[1743]), .B(DB[1728]), .Z(n2444) );
  AND U4244 ( .A(n50), .B(n2445), .Z(n2443) );
  XOR U4245 ( .A(n2446), .B(n2447), .Z(n2445) );
  XOR U4246 ( .A(DB[1728]), .B(DB[1713]), .Z(n2447) );
  AND U4247 ( .A(n54), .B(n2448), .Z(n2446) );
  XOR U4248 ( .A(n2449), .B(n2450), .Z(n2448) );
  XOR U4249 ( .A(DB[1713]), .B(DB[1698]), .Z(n2450) );
  AND U4250 ( .A(n58), .B(n2451), .Z(n2449) );
  XOR U4251 ( .A(n2452), .B(n2453), .Z(n2451) );
  XOR U4252 ( .A(DB[1698]), .B(DB[1683]), .Z(n2453) );
  AND U4253 ( .A(n62), .B(n2454), .Z(n2452) );
  XOR U4254 ( .A(n2455), .B(n2456), .Z(n2454) );
  XOR U4255 ( .A(DB[1683]), .B(DB[1668]), .Z(n2456) );
  AND U4256 ( .A(n66), .B(n2457), .Z(n2455) );
  XOR U4257 ( .A(n2458), .B(n2459), .Z(n2457) );
  XOR U4258 ( .A(DB[1668]), .B(DB[1653]), .Z(n2459) );
  AND U4259 ( .A(n70), .B(n2460), .Z(n2458) );
  XOR U4260 ( .A(n2461), .B(n2462), .Z(n2460) );
  XOR U4261 ( .A(DB[1653]), .B(DB[1638]), .Z(n2462) );
  AND U4262 ( .A(n74), .B(n2463), .Z(n2461) );
  XOR U4263 ( .A(n2464), .B(n2465), .Z(n2463) );
  XOR U4264 ( .A(DB[1638]), .B(DB[1623]), .Z(n2465) );
  AND U4265 ( .A(n78), .B(n2466), .Z(n2464) );
  XOR U4266 ( .A(n2467), .B(n2468), .Z(n2466) );
  XOR U4267 ( .A(DB[1623]), .B(DB[1608]), .Z(n2468) );
  AND U4268 ( .A(n82), .B(n2469), .Z(n2467) );
  XOR U4269 ( .A(n2470), .B(n2471), .Z(n2469) );
  XOR U4270 ( .A(DB[1608]), .B(DB[1593]), .Z(n2471) );
  AND U4271 ( .A(n86), .B(n2472), .Z(n2470) );
  XOR U4272 ( .A(n2473), .B(n2474), .Z(n2472) );
  XOR U4273 ( .A(DB[1593]), .B(DB[1578]), .Z(n2474) );
  AND U4274 ( .A(n90), .B(n2475), .Z(n2473) );
  XOR U4275 ( .A(n2476), .B(n2477), .Z(n2475) );
  XOR U4276 ( .A(DB[1578]), .B(DB[1563]), .Z(n2477) );
  AND U4277 ( .A(n94), .B(n2478), .Z(n2476) );
  XOR U4278 ( .A(n2479), .B(n2480), .Z(n2478) );
  XOR U4279 ( .A(DB[1563]), .B(DB[1548]), .Z(n2480) );
  AND U4280 ( .A(n98), .B(n2481), .Z(n2479) );
  XOR U4281 ( .A(n2482), .B(n2483), .Z(n2481) );
  XOR U4282 ( .A(DB[1548]), .B(DB[1533]), .Z(n2483) );
  AND U4283 ( .A(n102), .B(n2484), .Z(n2482) );
  XOR U4284 ( .A(n2485), .B(n2486), .Z(n2484) );
  XOR U4285 ( .A(DB[1533]), .B(DB[1518]), .Z(n2486) );
  AND U4286 ( .A(n106), .B(n2487), .Z(n2485) );
  XOR U4287 ( .A(n2488), .B(n2489), .Z(n2487) );
  XOR U4288 ( .A(DB[1518]), .B(DB[1503]), .Z(n2489) );
  AND U4289 ( .A(n110), .B(n2490), .Z(n2488) );
  XOR U4290 ( .A(n2491), .B(n2492), .Z(n2490) );
  XOR U4291 ( .A(DB[1503]), .B(DB[1488]), .Z(n2492) );
  AND U4292 ( .A(n114), .B(n2493), .Z(n2491) );
  XOR U4293 ( .A(n2494), .B(n2495), .Z(n2493) );
  XOR U4294 ( .A(DB[1488]), .B(DB[1473]), .Z(n2495) );
  AND U4295 ( .A(n118), .B(n2496), .Z(n2494) );
  XOR U4296 ( .A(n2497), .B(n2498), .Z(n2496) );
  XOR U4297 ( .A(DB[1473]), .B(DB[1458]), .Z(n2498) );
  AND U4298 ( .A(n122), .B(n2499), .Z(n2497) );
  XOR U4299 ( .A(n2500), .B(n2501), .Z(n2499) );
  XOR U4300 ( .A(DB[1458]), .B(DB[1443]), .Z(n2501) );
  AND U4301 ( .A(n126), .B(n2502), .Z(n2500) );
  XOR U4302 ( .A(n2503), .B(n2504), .Z(n2502) );
  XOR U4303 ( .A(DB[1443]), .B(DB[1428]), .Z(n2504) );
  AND U4304 ( .A(n130), .B(n2505), .Z(n2503) );
  XOR U4305 ( .A(n2506), .B(n2507), .Z(n2505) );
  XOR U4306 ( .A(DB[1428]), .B(DB[1413]), .Z(n2507) );
  AND U4307 ( .A(n134), .B(n2508), .Z(n2506) );
  XOR U4308 ( .A(n2509), .B(n2510), .Z(n2508) );
  XOR U4309 ( .A(DB[1413]), .B(DB[1398]), .Z(n2510) );
  AND U4310 ( .A(n138), .B(n2511), .Z(n2509) );
  XOR U4311 ( .A(n2512), .B(n2513), .Z(n2511) );
  XOR U4312 ( .A(DB[1398]), .B(DB[1383]), .Z(n2513) );
  AND U4313 ( .A(n142), .B(n2514), .Z(n2512) );
  XOR U4314 ( .A(n2515), .B(n2516), .Z(n2514) );
  XOR U4315 ( .A(DB[1383]), .B(DB[1368]), .Z(n2516) );
  AND U4316 ( .A(n146), .B(n2517), .Z(n2515) );
  XOR U4317 ( .A(n2518), .B(n2519), .Z(n2517) );
  XOR U4318 ( .A(DB[1368]), .B(DB[1353]), .Z(n2519) );
  AND U4319 ( .A(n150), .B(n2520), .Z(n2518) );
  XOR U4320 ( .A(n2521), .B(n2522), .Z(n2520) );
  XOR U4321 ( .A(DB[1353]), .B(DB[1338]), .Z(n2522) );
  AND U4322 ( .A(n154), .B(n2523), .Z(n2521) );
  XOR U4323 ( .A(n2524), .B(n2525), .Z(n2523) );
  XOR U4324 ( .A(DB[1338]), .B(DB[1323]), .Z(n2525) );
  AND U4325 ( .A(n158), .B(n2526), .Z(n2524) );
  XOR U4326 ( .A(n2527), .B(n2528), .Z(n2526) );
  XOR U4327 ( .A(DB[1323]), .B(DB[1308]), .Z(n2528) );
  AND U4328 ( .A(n162), .B(n2529), .Z(n2527) );
  XOR U4329 ( .A(n2530), .B(n2531), .Z(n2529) );
  XOR U4330 ( .A(DB[1308]), .B(DB[1293]), .Z(n2531) );
  AND U4331 ( .A(n166), .B(n2532), .Z(n2530) );
  XOR U4332 ( .A(n2533), .B(n2534), .Z(n2532) );
  XOR U4333 ( .A(DB[1293]), .B(DB[1278]), .Z(n2534) );
  AND U4334 ( .A(n170), .B(n2535), .Z(n2533) );
  XOR U4335 ( .A(n2536), .B(n2537), .Z(n2535) );
  XOR U4336 ( .A(DB[1278]), .B(DB[1263]), .Z(n2537) );
  AND U4337 ( .A(n174), .B(n2538), .Z(n2536) );
  XOR U4338 ( .A(n2539), .B(n2540), .Z(n2538) );
  XOR U4339 ( .A(DB[1263]), .B(DB[1248]), .Z(n2540) );
  AND U4340 ( .A(n178), .B(n2541), .Z(n2539) );
  XOR U4341 ( .A(n2542), .B(n2543), .Z(n2541) );
  XOR U4342 ( .A(DB[1248]), .B(DB[1233]), .Z(n2543) );
  AND U4343 ( .A(n182), .B(n2544), .Z(n2542) );
  XOR U4344 ( .A(n2545), .B(n2546), .Z(n2544) );
  XOR U4345 ( .A(DB[1233]), .B(DB[1218]), .Z(n2546) );
  AND U4346 ( .A(n186), .B(n2547), .Z(n2545) );
  XOR U4347 ( .A(n2548), .B(n2549), .Z(n2547) );
  XOR U4348 ( .A(DB[1218]), .B(DB[1203]), .Z(n2549) );
  AND U4349 ( .A(n190), .B(n2550), .Z(n2548) );
  XOR U4350 ( .A(n2551), .B(n2552), .Z(n2550) );
  XOR U4351 ( .A(DB[1203]), .B(DB[1188]), .Z(n2552) );
  AND U4352 ( .A(n194), .B(n2553), .Z(n2551) );
  XOR U4353 ( .A(n2554), .B(n2555), .Z(n2553) );
  XOR U4354 ( .A(DB[1188]), .B(DB[1173]), .Z(n2555) );
  AND U4355 ( .A(n198), .B(n2556), .Z(n2554) );
  XOR U4356 ( .A(n2557), .B(n2558), .Z(n2556) );
  XOR U4357 ( .A(DB[1173]), .B(DB[1158]), .Z(n2558) );
  AND U4358 ( .A(n202), .B(n2559), .Z(n2557) );
  XOR U4359 ( .A(n2560), .B(n2561), .Z(n2559) );
  XOR U4360 ( .A(DB[1158]), .B(DB[1143]), .Z(n2561) );
  AND U4361 ( .A(n206), .B(n2562), .Z(n2560) );
  XOR U4362 ( .A(n2563), .B(n2564), .Z(n2562) );
  XOR U4363 ( .A(DB[1143]), .B(DB[1128]), .Z(n2564) );
  AND U4364 ( .A(n210), .B(n2565), .Z(n2563) );
  XOR U4365 ( .A(n2566), .B(n2567), .Z(n2565) );
  XOR U4366 ( .A(DB[1128]), .B(DB[1113]), .Z(n2567) );
  AND U4367 ( .A(n214), .B(n2568), .Z(n2566) );
  XOR U4368 ( .A(n2569), .B(n2570), .Z(n2568) );
  XOR U4369 ( .A(DB[1113]), .B(DB[1098]), .Z(n2570) );
  AND U4370 ( .A(n218), .B(n2571), .Z(n2569) );
  XOR U4371 ( .A(n2572), .B(n2573), .Z(n2571) );
  XOR U4372 ( .A(DB[1098]), .B(DB[1083]), .Z(n2573) );
  AND U4373 ( .A(n222), .B(n2574), .Z(n2572) );
  XOR U4374 ( .A(n2575), .B(n2576), .Z(n2574) );
  XOR U4375 ( .A(DB[1083]), .B(DB[1068]), .Z(n2576) );
  AND U4376 ( .A(n226), .B(n2577), .Z(n2575) );
  XOR U4377 ( .A(n2578), .B(n2579), .Z(n2577) );
  XOR U4378 ( .A(DB[1068]), .B(DB[1053]), .Z(n2579) );
  AND U4379 ( .A(n230), .B(n2580), .Z(n2578) );
  XOR U4380 ( .A(n2581), .B(n2582), .Z(n2580) );
  XOR U4381 ( .A(DB[1053]), .B(DB[1038]), .Z(n2582) );
  AND U4382 ( .A(n234), .B(n2583), .Z(n2581) );
  XOR U4383 ( .A(n2584), .B(n2585), .Z(n2583) );
  XOR U4384 ( .A(DB[1038]), .B(DB[1023]), .Z(n2585) );
  AND U4385 ( .A(n238), .B(n2586), .Z(n2584) );
  XOR U4386 ( .A(n2587), .B(n2588), .Z(n2586) );
  XOR U4387 ( .A(DB[1023]), .B(DB[1008]), .Z(n2588) );
  AND U4388 ( .A(n242), .B(n2589), .Z(n2587) );
  XOR U4389 ( .A(n2590), .B(n2591), .Z(n2589) );
  XOR U4390 ( .A(DB[993]), .B(DB[1008]), .Z(n2591) );
  AND U4391 ( .A(n246), .B(n2592), .Z(n2590) );
  XOR U4392 ( .A(n2593), .B(n2594), .Z(n2592) );
  XOR U4393 ( .A(DB[993]), .B(DB[978]), .Z(n2594) );
  AND U4394 ( .A(n250), .B(n2595), .Z(n2593) );
  XOR U4395 ( .A(n2596), .B(n2597), .Z(n2595) );
  XOR U4396 ( .A(DB[978]), .B(DB[963]), .Z(n2597) );
  AND U4397 ( .A(n254), .B(n2598), .Z(n2596) );
  XOR U4398 ( .A(n2599), .B(n2600), .Z(n2598) );
  XOR U4399 ( .A(DB[963]), .B(DB[948]), .Z(n2600) );
  AND U4400 ( .A(n258), .B(n2601), .Z(n2599) );
  XOR U4401 ( .A(n2602), .B(n2603), .Z(n2601) );
  XOR U4402 ( .A(DB[948]), .B(DB[933]), .Z(n2603) );
  AND U4403 ( .A(n262), .B(n2604), .Z(n2602) );
  XOR U4404 ( .A(n2605), .B(n2606), .Z(n2604) );
  XOR U4405 ( .A(DB[933]), .B(DB[918]), .Z(n2606) );
  AND U4406 ( .A(n266), .B(n2607), .Z(n2605) );
  XOR U4407 ( .A(n2608), .B(n2609), .Z(n2607) );
  XOR U4408 ( .A(DB[918]), .B(DB[903]), .Z(n2609) );
  AND U4409 ( .A(n270), .B(n2610), .Z(n2608) );
  XOR U4410 ( .A(n2611), .B(n2612), .Z(n2610) );
  XOR U4411 ( .A(DB[903]), .B(DB[888]), .Z(n2612) );
  AND U4412 ( .A(n274), .B(n2613), .Z(n2611) );
  XOR U4413 ( .A(n2614), .B(n2615), .Z(n2613) );
  XOR U4414 ( .A(DB[888]), .B(DB[873]), .Z(n2615) );
  AND U4415 ( .A(n278), .B(n2616), .Z(n2614) );
  XOR U4416 ( .A(n2617), .B(n2618), .Z(n2616) );
  XOR U4417 ( .A(DB[873]), .B(DB[858]), .Z(n2618) );
  AND U4418 ( .A(n282), .B(n2619), .Z(n2617) );
  XOR U4419 ( .A(n2620), .B(n2621), .Z(n2619) );
  XOR U4420 ( .A(DB[858]), .B(DB[843]), .Z(n2621) );
  AND U4421 ( .A(n286), .B(n2622), .Z(n2620) );
  XOR U4422 ( .A(n2623), .B(n2624), .Z(n2622) );
  XOR U4423 ( .A(DB[843]), .B(DB[828]), .Z(n2624) );
  AND U4424 ( .A(n290), .B(n2625), .Z(n2623) );
  XOR U4425 ( .A(n2626), .B(n2627), .Z(n2625) );
  XOR U4426 ( .A(DB[828]), .B(DB[813]), .Z(n2627) );
  AND U4427 ( .A(n294), .B(n2628), .Z(n2626) );
  XOR U4428 ( .A(n2629), .B(n2630), .Z(n2628) );
  XOR U4429 ( .A(DB[813]), .B(DB[798]), .Z(n2630) );
  AND U4430 ( .A(n298), .B(n2631), .Z(n2629) );
  XOR U4431 ( .A(n2632), .B(n2633), .Z(n2631) );
  XOR U4432 ( .A(DB[798]), .B(DB[783]), .Z(n2633) );
  AND U4433 ( .A(n302), .B(n2634), .Z(n2632) );
  XOR U4434 ( .A(n2635), .B(n2636), .Z(n2634) );
  XOR U4435 ( .A(DB[783]), .B(DB[768]), .Z(n2636) );
  AND U4436 ( .A(n306), .B(n2637), .Z(n2635) );
  XOR U4437 ( .A(n2638), .B(n2639), .Z(n2637) );
  XOR U4438 ( .A(DB[768]), .B(DB[753]), .Z(n2639) );
  AND U4439 ( .A(n310), .B(n2640), .Z(n2638) );
  XOR U4440 ( .A(n2641), .B(n2642), .Z(n2640) );
  XOR U4441 ( .A(DB[753]), .B(DB[738]), .Z(n2642) );
  AND U4442 ( .A(n314), .B(n2643), .Z(n2641) );
  XOR U4443 ( .A(n2644), .B(n2645), .Z(n2643) );
  XOR U4444 ( .A(DB[738]), .B(DB[723]), .Z(n2645) );
  AND U4445 ( .A(n318), .B(n2646), .Z(n2644) );
  XOR U4446 ( .A(n2647), .B(n2648), .Z(n2646) );
  XOR U4447 ( .A(DB[723]), .B(DB[708]), .Z(n2648) );
  AND U4448 ( .A(n322), .B(n2649), .Z(n2647) );
  XOR U4449 ( .A(n2650), .B(n2651), .Z(n2649) );
  XOR U4450 ( .A(DB[708]), .B(DB[693]), .Z(n2651) );
  AND U4451 ( .A(n326), .B(n2652), .Z(n2650) );
  XOR U4452 ( .A(n2653), .B(n2654), .Z(n2652) );
  XOR U4453 ( .A(DB[693]), .B(DB[678]), .Z(n2654) );
  AND U4454 ( .A(n330), .B(n2655), .Z(n2653) );
  XOR U4455 ( .A(n2656), .B(n2657), .Z(n2655) );
  XOR U4456 ( .A(DB[678]), .B(DB[663]), .Z(n2657) );
  AND U4457 ( .A(n334), .B(n2658), .Z(n2656) );
  XOR U4458 ( .A(n2659), .B(n2660), .Z(n2658) );
  XOR U4459 ( .A(DB[663]), .B(DB[648]), .Z(n2660) );
  AND U4460 ( .A(n338), .B(n2661), .Z(n2659) );
  XOR U4461 ( .A(n2662), .B(n2663), .Z(n2661) );
  XOR U4462 ( .A(DB[648]), .B(DB[633]), .Z(n2663) );
  AND U4463 ( .A(n342), .B(n2664), .Z(n2662) );
  XOR U4464 ( .A(n2665), .B(n2666), .Z(n2664) );
  XOR U4465 ( .A(DB[633]), .B(DB[618]), .Z(n2666) );
  AND U4466 ( .A(n346), .B(n2667), .Z(n2665) );
  XOR U4467 ( .A(n2668), .B(n2669), .Z(n2667) );
  XOR U4468 ( .A(DB[618]), .B(DB[603]), .Z(n2669) );
  AND U4469 ( .A(n350), .B(n2670), .Z(n2668) );
  XOR U4470 ( .A(n2671), .B(n2672), .Z(n2670) );
  XOR U4471 ( .A(DB[603]), .B(DB[588]), .Z(n2672) );
  AND U4472 ( .A(n354), .B(n2673), .Z(n2671) );
  XOR U4473 ( .A(n2674), .B(n2675), .Z(n2673) );
  XOR U4474 ( .A(DB[588]), .B(DB[573]), .Z(n2675) );
  AND U4475 ( .A(n358), .B(n2676), .Z(n2674) );
  XOR U4476 ( .A(n2677), .B(n2678), .Z(n2676) );
  XOR U4477 ( .A(DB[573]), .B(DB[558]), .Z(n2678) );
  AND U4478 ( .A(n362), .B(n2679), .Z(n2677) );
  XOR U4479 ( .A(n2680), .B(n2681), .Z(n2679) );
  XOR U4480 ( .A(DB[558]), .B(DB[543]), .Z(n2681) );
  AND U4481 ( .A(n366), .B(n2682), .Z(n2680) );
  XOR U4482 ( .A(n2683), .B(n2684), .Z(n2682) );
  XOR U4483 ( .A(DB[543]), .B(DB[528]), .Z(n2684) );
  AND U4484 ( .A(n370), .B(n2685), .Z(n2683) );
  XOR U4485 ( .A(n2686), .B(n2687), .Z(n2685) );
  XOR U4486 ( .A(DB[528]), .B(DB[513]), .Z(n2687) );
  AND U4487 ( .A(n374), .B(n2688), .Z(n2686) );
  XOR U4488 ( .A(n2689), .B(n2690), .Z(n2688) );
  XOR U4489 ( .A(DB[513]), .B(DB[498]), .Z(n2690) );
  AND U4490 ( .A(n378), .B(n2691), .Z(n2689) );
  XOR U4491 ( .A(n2692), .B(n2693), .Z(n2691) );
  XOR U4492 ( .A(DB[498]), .B(DB[483]), .Z(n2693) );
  AND U4493 ( .A(n382), .B(n2694), .Z(n2692) );
  XOR U4494 ( .A(n2695), .B(n2696), .Z(n2694) );
  XOR U4495 ( .A(DB[483]), .B(DB[468]), .Z(n2696) );
  AND U4496 ( .A(n386), .B(n2697), .Z(n2695) );
  XOR U4497 ( .A(n2698), .B(n2699), .Z(n2697) );
  XOR U4498 ( .A(DB[468]), .B(DB[453]), .Z(n2699) );
  AND U4499 ( .A(n390), .B(n2700), .Z(n2698) );
  XOR U4500 ( .A(n2701), .B(n2702), .Z(n2700) );
  XOR U4501 ( .A(DB[453]), .B(DB[438]), .Z(n2702) );
  AND U4502 ( .A(n394), .B(n2703), .Z(n2701) );
  XOR U4503 ( .A(n2704), .B(n2705), .Z(n2703) );
  XOR U4504 ( .A(DB[438]), .B(DB[423]), .Z(n2705) );
  AND U4505 ( .A(n398), .B(n2706), .Z(n2704) );
  XOR U4506 ( .A(n2707), .B(n2708), .Z(n2706) );
  XOR U4507 ( .A(DB[423]), .B(DB[408]), .Z(n2708) );
  AND U4508 ( .A(n402), .B(n2709), .Z(n2707) );
  XOR U4509 ( .A(n2710), .B(n2711), .Z(n2709) );
  XOR U4510 ( .A(DB[408]), .B(DB[393]), .Z(n2711) );
  AND U4511 ( .A(n406), .B(n2712), .Z(n2710) );
  XOR U4512 ( .A(n2713), .B(n2714), .Z(n2712) );
  XOR U4513 ( .A(DB[393]), .B(DB[378]), .Z(n2714) );
  AND U4514 ( .A(n410), .B(n2715), .Z(n2713) );
  XOR U4515 ( .A(n2716), .B(n2717), .Z(n2715) );
  XOR U4516 ( .A(DB[378]), .B(DB[363]), .Z(n2717) );
  AND U4517 ( .A(n414), .B(n2718), .Z(n2716) );
  XOR U4518 ( .A(n2719), .B(n2720), .Z(n2718) );
  XOR U4519 ( .A(DB[363]), .B(DB[348]), .Z(n2720) );
  AND U4520 ( .A(n418), .B(n2721), .Z(n2719) );
  XOR U4521 ( .A(n2722), .B(n2723), .Z(n2721) );
  XOR U4522 ( .A(DB[348]), .B(DB[333]), .Z(n2723) );
  AND U4523 ( .A(n422), .B(n2724), .Z(n2722) );
  XOR U4524 ( .A(n2725), .B(n2726), .Z(n2724) );
  XOR U4525 ( .A(DB[333]), .B(DB[318]), .Z(n2726) );
  AND U4526 ( .A(n426), .B(n2727), .Z(n2725) );
  XOR U4527 ( .A(n2728), .B(n2729), .Z(n2727) );
  XOR U4528 ( .A(DB[318]), .B(DB[303]), .Z(n2729) );
  AND U4529 ( .A(n430), .B(n2730), .Z(n2728) );
  XOR U4530 ( .A(n2731), .B(n2732), .Z(n2730) );
  XOR U4531 ( .A(DB[303]), .B(DB[288]), .Z(n2732) );
  AND U4532 ( .A(n434), .B(n2733), .Z(n2731) );
  XOR U4533 ( .A(n2734), .B(n2735), .Z(n2733) );
  XOR U4534 ( .A(DB[288]), .B(DB[273]), .Z(n2735) );
  AND U4535 ( .A(n438), .B(n2736), .Z(n2734) );
  XOR U4536 ( .A(n2737), .B(n2738), .Z(n2736) );
  XOR U4537 ( .A(DB[273]), .B(DB[258]), .Z(n2738) );
  AND U4538 ( .A(n442), .B(n2739), .Z(n2737) );
  XOR U4539 ( .A(n2740), .B(n2741), .Z(n2739) );
  XOR U4540 ( .A(DB[258]), .B(DB[243]), .Z(n2741) );
  AND U4541 ( .A(n446), .B(n2742), .Z(n2740) );
  XOR U4542 ( .A(n2743), .B(n2744), .Z(n2742) );
  XOR U4543 ( .A(DB[243]), .B(DB[228]), .Z(n2744) );
  AND U4544 ( .A(n450), .B(n2745), .Z(n2743) );
  XOR U4545 ( .A(n2746), .B(n2747), .Z(n2745) );
  XOR U4546 ( .A(DB[228]), .B(DB[213]), .Z(n2747) );
  AND U4547 ( .A(n454), .B(n2748), .Z(n2746) );
  XOR U4548 ( .A(n2749), .B(n2750), .Z(n2748) );
  XOR U4549 ( .A(DB[213]), .B(DB[198]), .Z(n2750) );
  AND U4550 ( .A(n458), .B(n2751), .Z(n2749) );
  XOR U4551 ( .A(n2752), .B(n2753), .Z(n2751) );
  XOR U4552 ( .A(DB[198]), .B(DB[183]), .Z(n2753) );
  AND U4553 ( .A(n462), .B(n2754), .Z(n2752) );
  XOR U4554 ( .A(n2755), .B(n2756), .Z(n2754) );
  XOR U4555 ( .A(DB[183]), .B(DB[168]), .Z(n2756) );
  AND U4556 ( .A(n466), .B(n2757), .Z(n2755) );
  XOR U4557 ( .A(n2758), .B(n2759), .Z(n2757) );
  XOR U4558 ( .A(DB[168]), .B(DB[153]), .Z(n2759) );
  AND U4559 ( .A(n470), .B(n2760), .Z(n2758) );
  XOR U4560 ( .A(n2761), .B(n2762), .Z(n2760) );
  XOR U4561 ( .A(DB[153]), .B(DB[138]), .Z(n2762) );
  AND U4562 ( .A(n474), .B(n2763), .Z(n2761) );
  XOR U4563 ( .A(n2764), .B(n2765), .Z(n2763) );
  XOR U4564 ( .A(DB[138]), .B(DB[123]), .Z(n2765) );
  AND U4565 ( .A(n478), .B(n2766), .Z(n2764) );
  XOR U4566 ( .A(n2767), .B(n2768), .Z(n2766) );
  XOR U4567 ( .A(DB[123]), .B(DB[108]), .Z(n2768) );
  AND U4568 ( .A(n482), .B(n2769), .Z(n2767) );
  XOR U4569 ( .A(n2770), .B(n2771), .Z(n2769) );
  XOR U4570 ( .A(DB[93]), .B(DB[108]), .Z(n2771) );
  AND U4571 ( .A(n486), .B(n2772), .Z(n2770) );
  XOR U4572 ( .A(n2773), .B(n2774), .Z(n2772) );
  XOR U4573 ( .A(DB[93]), .B(DB[78]), .Z(n2774) );
  AND U4574 ( .A(n490), .B(n2775), .Z(n2773) );
  XOR U4575 ( .A(n2776), .B(n2777), .Z(n2775) );
  XOR U4576 ( .A(DB[78]), .B(DB[63]), .Z(n2777) );
  AND U4577 ( .A(n494), .B(n2778), .Z(n2776) );
  XOR U4578 ( .A(n2779), .B(n2780), .Z(n2778) );
  XOR U4579 ( .A(DB[63]), .B(DB[48]), .Z(n2780) );
  AND U4580 ( .A(n498), .B(n2781), .Z(n2779) );
  XOR U4581 ( .A(n2782), .B(n2783), .Z(n2781) );
  XOR U4582 ( .A(DB[48]), .B(DB[33]), .Z(n2783) );
  AND U4583 ( .A(n502), .B(n2784), .Z(n2782) );
  XOR U4584 ( .A(n2785), .B(n2786), .Z(n2784) );
  XOR U4585 ( .A(DB[33]), .B(DB[18]), .Z(n2786) );
  AND U4586 ( .A(n506), .B(n2787), .Z(n2785) );
  XOR U4587 ( .A(DB[3]), .B(DB[18]), .Z(n2787) );
  XOR U4588 ( .A(DB[1907]), .B(n2788), .Z(min_val_out[2]) );
  AND U4589 ( .A(n2), .B(n2789), .Z(n2788) );
  XOR U4590 ( .A(n2790), .B(n2791), .Z(n2789) );
  XOR U4591 ( .A(DB[1907]), .B(DB[1892]), .Z(n2791) );
  AND U4592 ( .A(n6), .B(n2792), .Z(n2790) );
  XOR U4593 ( .A(n2793), .B(n2794), .Z(n2792) );
  XOR U4594 ( .A(DB[1892]), .B(DB[1877]), .Z(n2794) );
  AND U4595 ( .A(n10), .B(n2795), .Z(n2793) );
  XOR U4596 ( .A(n2796), .B(n2797), .Z(n2795) );
  XOR U4597 ( .A(DB[1877]), .B(DB[1862]), .Z(n2797) );
  AND U4598 ( .A(n14), .B(n2798), .Z(n2796) );
  XOR U4599 ( .A(n2799), .B(n2800), .Z(n2798) );
  XOR U4600 ( .A(DB[1862]), .B(DB[1847]), .Z(n2800) );
  AND U4601 ( .A(n18), .B(n2801), .Z(n2799) );
  XOR U4602 ( .A(n2802), .B(n2803), .Z(n2801) );
  XOR U4603 ( .A(DB[1847]), .B(DB[1832]), .Z(n2803) );
  AND U4604 ( .A(n22), .B(n2804), .Z(n2802) );
  XOR U4605 ( .A(n2805), .B(n2806), .Z(n2804) );
  XOR U4606 ( .A(DB[1832]), .B(DB[1817]), .Z(n2806) );
  AND U4607 ( .A(n26), .B(n2807), .Z(n2805) );
  XOR U4608 ( .A(n2808), .B(n2809), .Z(n2807) );
  XOR U4609 ( .A(DB[1817]), .B(DB[1802]), .Z(n2809) );
  AND U4610 ( .A(n30), .B(n2810), .Z(n2808) );
  XOR U4611 ( .A(n2811), .B(n2812), .Z(n2810) );
  XOR U4612 ( .A(DB[1802]), .B(DB[1787]), .Z(n2812) );
  AND U4613 ( .A(n34), .B(n2813), .Z(n2811) );
  XOR U4614 ( .A(n2814), .B(n2815), .Z(n2813) );
  XOR U4615 ( .A(DB[1787]), .B(DB[1772]), .Z(n2815) );
  AND U4616 ( .A(n38), .B(n2816), .Z(n2814) );
  XOR U4617 ( .A(n2817), .B(n2818), .Z(n2816) );
  XOR U4618 ( .A(DB[1772]), .B(DB[1757]), .Z(n2818) );
  AND U4619 ( .A(n42), .B(n2819), .Z(n2817) );
  XOR U4620 ( .A(n2820), .B(n2821), .Z(n2819) );
  XOR U4621 ( .A(DB[1757]), .B(DB[1742]), .Z(n2821) );
  AND U4622 ( .A(n46), .B(n2822), .Z(n2820) );
  XOR U4623 ( .A(n2823), .B(n2824), .Z(n2822) );
  XOR U4624 ( .A(DB[1742]), .B(DB[1727]), .Z(n2824) );
  AND U4625 ( .A(n50), .B(n2825), .Z(n2823) );
  XOR U4626 ( .A(n2826), .B(n2827), .Z(n2825) );
  XOR U4627 ( .A(DB[1727]), .B(DB[1712]), .Z(n2827) );
  AND U4628 ( .A(n54), .B(n2828), .Z(n2826) );
  XOR U4629 ( .A(n2829), .B(n2830), .Z(n2828) );
  XOR U4630 ( .A(DB[1712]), .B(DB[1697]), .Z(n2830) );
  AND U4631 ( .A(n58), .B(n2831), .Z(n2829) );
  XOR U4632 ( .A(n2832), .B(n2833), .Z(n2831) );
  XOR U4633 ( .A(DB[1697]), .B(DB[1682]), .Z(n2833) );
  AND U4634 ( .A(n62), .B(n2834), .Z(n2832) );
  XOR U4635 ( .A(n2835), .B(n2836), .Z(n2834) );
  XOR U4636 ( .A(DB[1682]), .B(DB[1667]), .Z(n2836) );
  AND U4637 ( .A(n66), .B(n2837), .Z(n2835) );
  XOR U4638 ( .A(n2838), .B(n2839), .Z(n2837) );
  XOR U4639 ( .A(DB[1667]), .B(DB[1652]), .Z(n2839) );
  AND U4640 ( .A(n70), .B(n2840), .Z(n2838) );
  XOR U4641 ( .A(n2841), .B(n2842), .Z(n2840) );
  XOR U4642 ( .A(DB[1652]), .B(DB[1637]), .Z(n2842) );
  AND U4643 ( .A(n74), .B(n2843), .Z(n2841) );
  XOR U4644 ( .A(n2844), .B(n2845), .Z(n2843) );
  XOR U4645 ( .A(DB[1637]), .B(DB[1622]), .Z(n2845) );
  AND U4646 ( .A(n78), .B(n2846), .Z(n2844) );
  XOR U4647 ( .A(n2847), .B(n2848), .Z(n2846) );
  XOR U4648 ( .A(DB[1622]), .B(DB[1607]), .Z(n2848) );
  AND U4649 ( .A(n82), .B(n2849), .Z(n2847) );
  XOR U4650 ( .A(n2850), .B(n2851), .Z(n2849) );
  XOR U4651 ( .A(DB[1607]), .B(DB[1592]), .Z(n2851) );
  AND U4652 ( .A(n86), .B(n2852), .Z(n2850) );
  XOR U4653 ( .A(n2853), .B(n2854), .Z(n2852) );
  XOR U4654 ( .A(DB[1592]), .B(DB[1577]), .Z(n2854) );
  AND U4655 ( .A(n90), .B(n2855), .Z(n2853) );
  XOR U4656 ( .A(n2856), .B(n2857), .Z(n2855) );
  XOR U4657 ( .A(DB[1577]), .B(DB[1562]), .Z(n2857) );
  AND U4658 ( .A(n94), .B(n2858), .Z(n2856) );
  XOR U4659 ( .A(n2859), .B(n2860), .Z(n2858) );
  XOR U4660 ( .A(DB[1562]), .B(DB[1547]), .Z(n2860) );
  AND U4661 ( .A(n98), .B(n2861), .Z(n2859) );
  XOR U4662 ( .A(n2862), .B(n2863), .Z(n2861) );
  XOR U4663 ( .A(DB[1547]), .B(DB[1532]), .Z(n2863) );
  AND U4664 ( .A(n102), .B(n2864), .Z(n2862) );
  XOR U4665 ( .A(n2865), .B(n2866), .Z(n2864) );
  XOR U4666 ( .A(DB[1532]), .B(DB[1517]), .Z(n2866) );
  AND U4667 ( .A(n106), .B(n2867), .Z(n2865) );
  XOR U4668 ( .A(n2868), .B(n2869), .Z(n2867) );
  XOR U4669 ( .A(DB[1517]), .B(DB[1502]), .Z(n2869) );
  AND U4670 ( .A(n110), .B(n2870), .Z(n2868) );
  XOR U4671 ( .A(n2871), .B(n2872), .Z(n2870) );
  XOR U4672 ( .A(DB[1502]), .B(DB[1487]), .Z(n2872) );
  AND U4673 ( .A(n114), .B(n2873), .Z(n2871) );
  XOR U4674 ( .A(n2874), .B(n2875), .Z(n2873) );
  XOR U4675 ( .A(DB[1487]), .B(DB[1472]), .Z(n2875) );
  AND U4676 ( .A(n118), .B(n2876), .Z(n2874) );
  XOR U4677 ( .A(n2877), .B(n2878), .Z(n2876) );
  XOR U4678 ( .A(DB[1472]), .B(DB[1457]), .Z(n2878) );
  AND U4679 ( .A(n122), .B(n2879), .Z(n2877) );
  XOR U4680 ( .A(n2880), .B(n2881), .Z(n2879) );
  XOR U4681 ( .A(DB[1457]), .B(DB[1442]), .Z(n2881) );
  AND U4682 ( .A(n126), .B(n2882), .Z(n2880) );
  XOR U4683 ( .A(n2883), .B(n2884), .Z(n2882) );
  XOR U4684 ( .A(DB[1442]), .B(DB[1427]), .Z(n2884) );
  AND U4685 ( .A(n130), .B(n2885), .Z(n2883) );
  XOR U4686 ( .A(n2886), .B(n2887), .Z(n2885) );
  XOR U4687 ( .A(DB[1427]), .B(DB[1412]), .Z(n2887) );
  AND U4688 ( .A(n134), .B(n2888), .Z(n2886) );
  XOR U4689 ( .A(n2889), .B(n2890), .Z(n2888) );
  XOR U4690 ( .A(DB[1412]), .B(DB[1397]), .Z(n2890) );
  AND U4691 ( .A(n138), .B(n2891), .Z(n2889) );
  XOR U4692 ( .A(n2892), .B(n2893), .Z(n2891) );
  XOR U4693 ( .A(DB[1397]), .B(DB[1382]), .Z(n2893) );
  AND U4694 ( .A(n142), .B(n2894), .Z(n2892) );
  XOR U4695 ( .A(n2895), .B(n2896), .Z(n2894) );
  XOR U4696 ( .A(DB[1382]), .B(DB[1367]), .Z(n2896) );
  AND U4697 ( .A(n146), .B(n2897), .Z(n2895) );
  XOR U4698 ( .A(n2898), .B(n2899), .Z(n2897) );
  XOR U4699 ( .A(DB[1367]), .B(DB[1352]), .Z(n2899) );
  AND U4700 ( .A(n150), .B(n2900), .Z(n2898) );
  XOR U4701 ( .A(n2901), .B(n2902), .Z(n2900) );
  XOR U4702 ( .A(DB[1352]), .B(DB[1337]), .Z(n2902) );
  AND U4703 ( .A(n154), .B(n2903), .Z(n2901) );
  XOR U4704 ( .A(n2904), .B(n2905), .Z(n2903) );
  XOR U4705 ( .A(DB[1337]), .B(DB[1322]), .Z(n2905) );
  AND U4706 ( .A(n158), .B(n2906), .Z(n2904) );
  XOR U4707 ( .A(n2907), .B(n2908), .Z(n2906) );
  XOR U4708 ( .A(DB[1322]), .B(DB[1307]), .Z(n2908) );
  AND U4709 ( .A(n162), .B(n2909), .Z(n2907) );
  XOR U4710 ( .A(n2910), .B(n2911), .Z(n2909) );
  XOR U4711 ( .A(DB[1307]), .B(DB[1292]), .Z(n2911) );
  AND U4712 ( .A(n166), .B(n2912), .Z(n2910) );
  XOR U4713 ( .A(n2913), .B(n2914), .Z(n2912) );
  XOR U4714 ( .A(DB[1292]), .B(DB[1277]), .Z(n2914) );
  AND U4715 ( .A(n170), .B(n2915), .Z(n2913) );
  XOR U4716 ( .A(n2916), .B(n2917), .Z(n2915) );
  XOR U4717 ( .A(DB[1277]), .B(DB[1262]), .Z(n2917) );
  AND U4718 ( .A(n174), .B(n2918), .Z(n2916) );
  XOR U4719 ( .A(n2919), .B(n2920), .Z(n2918) );
  XOR U4720 ( .A(DB[1262]), .B(DB[1247]), .Z(n2920) );
  AND U4721 ( .A(n178), .B(n2921), .Z(n2919) );
  XOR U4722 ( .A(n2922), .B(n2923), .Z(n2921) );
  XOR U4723 ( .A(DB[1247]), .B(DB[1232]), .Z(n2923) );
  AND U4724 ( .A(n182), .B(n2924), .Z(n2922) );
  XOR U4725 ( .A(n2925), .B(n2926), .Z(n2924) );
  XOR U4726 ( .A(DB[1232]), .B(DB[1217]), .Z(n2926) );
  AND U4727 ( .A(n186), .B(n2927), .Z(n2925) );
  XOR U4728 ( .A(n2928), .B(n2929), .Z(n2927) );
  XOR U4729 ( .A(DB[1217]), .B(DB[1202]), .Z(n2929) );
  AND U4730 ( .A(n190), .B(n2930), .Z(n2928) );
  XOR U4731 ( .A(n2931), .B(n2932), .Z(n2930) );
  XOR U4732 ( .A(DB[1202]), .B(DB[1187]), .Z(n2932) );
  AND U4733 ( .A(n194), .B(n2933), .Z(n2931) );
  XOR U4734 ( .A(n2934), .B(n2935), .Z(n2933) );
  XOR U4735 ( .A(DB[1187]), .B(DB[1172]), .Z(n2935) );
  AND U4736 ( .A(n198), .B(n2936), .Z(n2934) );
  XOR U4737 ( .A(n2937), .B(n2938), .Z(n2936) );
  XOR U4738 ( .A(DB[1172]), .B(DB[1157]), .Z(n2938) );
  AND U4739 ( .A(n202), .B(n2939), .Z(n2937) );
  XOR U4740 ( .A(n2940), .B(n2941), .Z(n2939) );
  XOR U4741 ( .A(DB[1157]), .B(DB[1142]), .Z(n2941) );
  AND U4742 ( .A(n206), .B(n2942), .Z(n2940) );
  XOR U4743 ( .A(n2943), .B(n2944), .Z(n2942) );
  XOR U4744 ( .A(DB[1142]), .B(DB[1127]), .Z(n2944) );
  AND U4745 ( .A(n210), .B(n2945), .Z(n2943) );
  XOR U4746 ( .A(n2946), .B(n2947), .Z(n2945) );
  XOR U4747 ( .A(DB[1127]), .B(DB[1112]), .Z(n2947) );
  AND U4748 ( .A(n214), .B(n2948), .Z(n2946) );
  XOR U4749 ( .A(n2949), .B(n2950), .Z(n2948) );
  XOR U4750 ( .A(DB[1112]), .B(DB[1097]), .Z(n2950) );
  AND U4751 ( .A(n218), .B(n2951), .Z(n2949) );
  XOR U4752 ( .A(n2952), .B(n2953), .Z(n2951) );
  XOR U4753 ( .A(DB[1097]), .B(DB[1082]), .Z(n2953) );
  AND U4754 ( .A(n222), .B(n2954), .Z(n2952) );
  XOR U4755 ( .A(n2955), .B(n2956), .Z(n2954) );
  XOR U4756 ( .A(DB[1082]), .B(DB[1067]), .Z(n2956) );
  AND U4757 ( .A(n226), .B(n2957), .Z(n2955) );
  XOR U4758 ( .A(n2958), .B(n2959), .Z(n2957) );
  XOR U4759 ( .A(DB[1067]), .B(DB[1052]), .Z(n2959) );
  AND U4760 ( .A(n230), .B(n2960), .Z(n2958) );
  XOR U4761 ( .A(n2961), .B(n2962), .Z(n2960) );
  XOR U4762 ( .A(DB[1052]), .B(DB[1037]), .Z(n2962) );
  AND U4763 ( .A(n234), .B(n2963), .Z(n2961) );
  XOR U4764 ( .A(n2964), .B(n2965), .Z(n2963) );
  XOR U4765 ( .A(DB[1037]), .B(DB[1022]), .Z(n2965) );
  AND U4766 ( .A(n238), .B(n2966), .Z(n2964) );
  XOR U4767 ( .A(n2967), .B(n2968), .Z(n2966) );
  XOR U4768 ( .A(DB[1022]), .B(DB[1007]), .Z(n2968) );
  AND U4769 ( .A(n242), .B(n2969), .Z(n2967) );
  XOR U4770 ( .A(n2970), .B(n2971), .Z(n2969) );
  XOR U4771 ( .A(DB[992]), .B(DB[1007]), .Z(n2971) );
  AND U4772 ( .A(n246), .B(n2972), .Z(n2970) );
  XOR U4773 ( .A(n2973), .B(n2974), .Z(n2972) );
  XOR U4774 ( .A(DB[992]), .B(DB[977]), .Z(n2974) );
  AND U4775 ( .A(n250), .B(n2975), .Z(n2973) );
  XOR U4776 ( .A(n2976), .B(n2977), .Z(n2975) );
  XOR U4777 ( .A(DB[977]), .B(DB[962]), .Z(n2977) );
  AND U4778 ( .A(n254), .B(n2978), .Z(n2976) );
  XOR U4779 ( .A(n2979), .B(n2980), .Z(n2978) );
  XOR U4780 ( .A(DB[962]), .B(DB[947]), .Z(n2980) );
  AND U4781 ( .A(n258), .B(n2981), .Z(n2979) );
  XOR U4782 ( .A(n2982), .B(n2983), .Z(n2981) );
  XOR U4783 ( .A(DB[947]), .B(DB[932]), .Z(n2983) );
  AND U4784 ( .A(n262), .B(n2984), .Z(n2982) );
  XOR U4785 ( .A(n2985), .B(n2986), .Z(n2984) );
  XOR U4786 ( .A(DB[932]), .B(DB[917]), .Z(n2986) );
  AND U4787 ( .A(n266), .B(n2987), .Z(n2985) );
  XOR U4788 ( .A(n2988), .B(n2989), .Z(n2987) );
  XOR U4789 ( .A(DB[917]), .B(DB[902]), .Z(n2989) );
  AND U4790 ( .A(n270), .B(n2990), .Z(n2988) );
  XOR U4791 ( .A(n2991), .B(n2992), .Z(n2990) );
  XOR U4792 ( .A(DB[902]), .B(DB[887]), .Z(n2992) );
  AND U4793 ( .A(n274), .B(n2993), .Z(n2991) );
  XOR U4794 ( .A(n2994), .B(n2995), .Z(n2993) );
  XOR U4795 ( .A(DB[887]), .B(DB[872]), .Z(n2995) );
  AND U4796 ( .A(n278), .B(n2996), .Z(n2994) );
  XOR U4797 ( .A(n2997), .B(n2998), .Z(n2996) );
  XOR U4798 ( .A(DB[872]), .B(DB[857]), .Z(n2998) );
  AND U4799 ( .A(n282), .B(n2999), .Z(n2997) );
  XOR U4800 ( .A(n3000), .B(n3001), .Z(n2999) );
  XOR U4801 ( .A(DB[857]), .B(DB[842]), .Z(n3001) );
  AND U4802 ( .A(n286), .B(n3002), .Z(n3000) );
  XOR U4803 ( .A(n3003), .B(n3004), .Z(n3002) );
  XOR U4804 ( .A(DB[842]), .B(DB[827]), .Z(n3004) );
  AND U4805 ( .A(n290), .B(n3005), .Z(n3003) );
  XOR U4806 ( .A(n3006), .B(n3007), .Z(n3005) );
  XOR U4807 ( .A(DB[827]), .B(DB[812]), .Z(n3007) );
  AND U4808 ( .A(n294), .B(n3008), .Z(n3006) );
  XOR U4809 ( .A(n3009), .B(n3010), .Z(n3008) );
  XOR U4810 ( .A(DB[812]), .B(DB[797]), .Z(n3010) );
  AND U4811 ( .A(n298), .B(n3011), .Z(n3009) );
  XOR U4812 ( .A(n3012), .B(n3013), .Z(n3011) );
  XOR U4813 ( .A(DB[797]), .B(DB[782]), .Z(n3013) );
  AND U4814 ( .A(n302), .B(n3014), .Z(n3012) );
  XOR U4815 ( .A(n3015), .B(n3016), .Z(n3014) );
  XOR U4816 ( .A(DB[782]), .B(DB[767]), .Z(n3016) );
  AND U4817 ( .A(n306), .B(n3017), .Z(n3015) );
  XOR U4818 ( .A(n3018), .B(n3019), .Z(n3017) );
  XOR U4819 ( .A(DB[767]), .B(DB[752]), .Z(n3019) );
  AND U4820 ( .A(n310), .B(n3020), .Z(n3018) );
  XOR U4821 ( .A(n3021), .B(n3022), .Z(n3020) );
  XOR U4822 ( .A(DB[752]), .B(DB[737]), .Z(n3022) );
  AND U4823 ( .A(n314), .B(n3023), .Z(n3021) );
  XOR U4824 ( .A(n3024), .B(n3025), .Z(n3023) );
  XOR U4825 ( .A(DB[737]), .B(DB[722]), .Z(n3025) );
  AND U4826 ( .A(n318), .B(n3026), .Z(n3024) );
  XOR U4827 ( .A(n3027), .B(n3028), .Z(n3026) );
  XOR U4828 ( .A(DB[722]), .B(DB[707]), .Z(n3028) );
  AND U4829 ( .A(n322), .B(n3029), .Z(n3027) );
  XOR U4830 ( .A(n3030), .B(n3031), .Z(n3029) );
  XOR U4831 ( .A(DB[707]), .B(DB[692]), .Z(n3031) );
  AND U4832 ( .A(n326), .B(n3032), .Z(n3030) );
  XOR U4833 ( .A(n3033), .B(n3034), .Z(n3032) );
  XOR U4834 ( .A(DB[692]), .B(DB[677]), .Z(n3034) );
  AND U4835 ( .A(n330), .B(n3035), .Z(n3033) );
  XOR U4836 ( .A(n3036), .B(n3037), .Z(n3035) );
  XOR U4837 ( .A(DB[677]), .B(DB[662]), .Z(n3037) );
  AND U4838 ( .A(n334), .B(n3038), .Z(n3036) );
  XOR U4839 ( .A(n3039), .B(n3040), .Z(n3038) );
  XOR U4840 ( .A(DB[662]), .B(DB[647]), .Z(n3040) );
  AND U4841 ( .A(n338), .B(n3041), .Z(n3039) );
  XOR U4842 ( .A(n3042), .B(n3043), .Z(n3041) );
  XOR U4843 ( .A(DB[647]), .B(DB[632]), .Z(n3043) );
  AND U4844 ( .A(n342), .B(n3044), .Z(n3042) );
  XOR U4845 ( .A(n3045), .B(n3046), .Z(n3044) );
  XOR U4846 ( .A(DB[632]), .B(DB[617]), .Z(n3046) );
  AND U4847 ( .A(n346), .B(n3047), .Z(n3045) );
  XOR U4848 ( .A(n3048), .B(n3049), .Z(n3047) );
  XOR U4849 ( .A(DB[617]), .B(DB[602]), .Z(n3049) );
  AND U4850 ( .A(n350), .B(n3050), .Z(n3048) );
  XOR U4851 ( .A(n3051), .B(n3052), .Z(n3050) );
  XOR U4852 ( .A(DB[602]), .B(DB[587]), .Z(n3052) );
  AND U4853 ( .A(n354), .B(n3053), .Z(n3051) );
  XOR U4854 ( .A(n3054), .B(n3055), .Z(n3053) );
  XOR U4855 ( .A(DB[587]), .B(DB[572]), .Z(n3055) );
  AND U4856 ( .A(n358), .B(n3056), .Z(n3054) );
  XOR U4857 ( .A(n3057), .B(n3058), .Z(n3056) );
  XOR U4858 ( .A(DB[572]), .B(DB[557]), .Z(n3058) );
  AND U4859 ( .A(n362), .B(n3059), .Z(n3057) );
  XOR U4860 ( .A(n3060), .B(n3061), .Z(n3059) );
  XOR U4861 ( .A(DB[557]), .B(DB[542]), .Z(n3061) );
  AND U4862 ( .A(n366), .B(n3062), .Z(n3060) );
  XOR U4863 ( .A(n3063), .B(n3064), .Z(n3062) );
  XOR U4864 ( .A(DB[542]), .B(DB[527]), .Z(n3064) );
  AND U4865 ( .A(n370), .B(n3065), .Z(n3063) );
  XOR U4866 ( .A(n3066), .B(n3067), .Z(n3065) );
  XOR U4867 ( .A(DB[527]), .B(DB[512]), .Z(n3067) );
  AND U4868 ( .A(n374), .B(n3068), .Z(n3066) );
  XOR U4869 ( .A(n3069), .B(n3070), .Z(n3068) );
  XOR U4870 ( .A(DB[512]), .B(DB[497]), .Z(n3070) );
  AND U4871 ( .A(n378), .B(n3071), .Z(n3069) );
  XOR U4872 ( .A(n3072), .B(n3073), .Z(n3071) );
  XOR U4873 ( .A(DB[497]), .B(DB[482]), .Z(n3073) );
  AND U4874 ( .A(n382), .B(n3074), .Z(n3072) );
  XOR U4875 ( .A(n3075), .B(n3076), .Z(n3074) );
  XOR U4876 ( .A(DB[482]), .B(DB[467]), .Z(n3076) );
  AND U4877 ( .A(n386), .B(n3077), .Z(n3075) );
  XOR U4878 ( .A(n3078), .B(n3079), .Z(n3077) );
  XOR U4879 ( .A(DB[467]), .B(DB[452]), .Z(n3079) );
  AND U4880 ( .A(n390), .B(n3080), .Z(n3078) );
  XOR U4881 ( .A(n3081), .B(n3082), .Z(n3080) );
  XOR U4882 ( .A(DB[452]), .B(DB[437]), .Z(n3082) );
  AND U4883 ( .A(n394), .B(n3083), .Z(n3081) );
  XOR U4884 ( .A(n3084), .B(n3085), .Z(n3083) );
  XOR U4885 ( .A(DB[437]), .B(DB[422]), .Z(n3085) );
  AND U4886 ( .A(n398), .B(n3086), .Z(n3084) );
  XOR U4887 ( .A(n3087), .B(n3088), .Z(n3086) );
  XOR U4888 ( .A(DB[422]), .B(DB[407]), .Z(n3088) );
  AND U4889 ( .A(n402), .B(n3089), .Z(n3087) );
  XOR U4890 ( .A(n3090), .B(n3091), .Z(n3089) );
  XOR U4891 ( .A(DB[407]), .B(DB[392]), .Z(n3091) );
  AND U4892 ( .A(n406), .B(n3092), .Z(n3090) );
  XOR U4893 ( .A(n3093), .B(n3094), .Z(n3092) );
  XOR U4894 ( .A(DB[392]), .B(DB[377]), .Z(n3094) );
  AND U4895 ( .A(n410), .B(n3095), .Z(n3093) );
  XOR U4896 ( .A(n3096), .B(n3097), .Z(n3095) );
  XOR U4897 ( .A(DB[377]), .B(DB[362]), .Z(n3097) );
  AND U4898 ( .A(n414), .B(n3098), .Z(n3096) );
  XOR U4899 ( .A(n3099), .B(n3100), .Z(n3098) );
  XOR U4900 ( .A(DB[362]), .B(DB[347]), .Z(n3100) );
  AND U4901 ( .A(n418), .B(n3101), .Z(n3099) );
  XOR U4902 ( .A(n3102), .B(n3103), .Z(n3101) );
  XOR U4903 ( .A(DB[347]), .B(DB[332]), .Z(n3103) );
  AND U4904 ( .A(n422), .B(n3104), .Z(n3102) );
  XOR U4905 ( .A(n3105), .B(n3106), .Z(n3104) );
  XOR U4906 ( .A(DB[332]), .B(DB[317]), .Z(n3106) );
  AND U4907 ( .A(n426), .B(n3107), .Z(n3105) );
  XOR U4908 ( .A(n3108), .B(n3109), .Z(n3107) );
  XOR U4909 ( .A(DB[317]), .B(DB[302]), .Z(n3109) );
  AND U4910 ( .A(n430), .B(n3110), .Z(n3108) );
  XOR U4911 ( .A(n3111), .B(n3112), .Z(n3110) );
  XOR U4912 ( .A(DB[302]), .B(DB[287]), .Z(n3112) );
  AND U4913 ( .A(n434), .B(n3113), .Z(n3111) );
  XOR U4914 ( .A(n3114), .B(n3115), .Z(n3113) );
  XOR U4915 ( .A(DB[287]), .B(DB[272]), .Z(n3115) );
  AND U4916 ( .A(n438), .B(n3116), .Z(n3114) );
  XOR U4917 ( .A(n3117), .B(n3118), .Z(n3116) );
  XOR U4918 ( .A(DB[272]), .B(DB[257]), .Z(n3118) );
  AND U4919 ( .A(n442), .B(n3119), .Z(n3117) );
  XOR U4920 ( .A(n3120), .B(n3121), .Z(n3119) );
  XOR U4921 ( .A(DB[257]), .B(DB[242]), .Z(n3121) );
  AND U4922 ( .A(n446), .B(n3122), .Z(n3120) );
  XOR U4923 ( .A(n3123), .B(n3124), .Z(n3122) );
  XOR U4924 ( .A(DB[242]), .B(DB[227]), .Z(n3124) );
  AND U4925 ( .A(n450), .B(n3125), .Z(n3123) );
  XOR U4926 ( .A(n3126), .B(n3127), .Z(n3125) );
  XOR U4927 ( .A(DB[227]), .B(DB[212]), .Z(n3127) );
  AND U4928 ( .A(n454), .B(n3128), .Z(n3126) );
  XOR U4929 ( .A(n3129), .B(n3130), .Z(n3128) );
  XOR U4930 ( .A(DB[212]), .B(DB[197]), .Z(n3130) );
  AND U4931 ( .A(n458), .B(n3131), .Z(n3129) );
  XOR U4932 ( .A(n3132), .B(n3133), .Z(n3131) );
  XOR U4933 ( .A(DB[197]), .B(DB[182]), .Z(n3133) );
  AND U4934 ( .A(n462), .B(n3134), .Z(n3132) );
  XOR U4935 ( .A(n3135), .B(n3136), .Z(n3134) );
  XOR U4936 ( .A(DB[182]), .B(DB[167]), .Z(n3136) );
  AND U4937 ( .A(n466), .B(n3137), .Z(n3135) );
  XOR U4938 ( .A(n3138), .B(n3139), .Z(n3137) );
  XOR U4939 ( .A(DB[167]), .B(DB[152]), .Z(n3139) );
  AND U4940 ( .A(n470), .B(n3140), .Z(n3138) );
  XOR U4941 ( .A(n3141), .B(n3142), .Z(n3140) );
  XOR U4942 ( .A(DB[152]), .B(DB[137]), .Z(n3142) );
  AND U4943 ( .A(n474), .B(n3143), .Z(n3141) );
  XOR U4944 ( .A(n3144), .B(n3145), .Z(n3143) );
  XOR U4945 ( .A(DB[137]), .B(DB[122]), .Z(n3145) );
  AND U4946 ( .A(n478), .B(n3146), .Z(n3144) );
  XOR U4947 ( .A(n3147), .B(n3148), .Z(n3146) );
  XOR U4948 ( .A(DB[122]), .B(DB[107]), .Z(n3148) );
  AND U4949 ( .A(n482), .B(n3149), .Z(n3147) );
  XOR U4950 ( .A(n3150), .B(n3151), .Z(n3149) );
  XOR U4951 ( .A(DB[92]), .B(DB[107]), .Z(n3151) );
  AND U4952 ( .A(n486), .B(n3152), .Z(n3150) );
  XOR U4953 ( .A(n3153), .B(n3154), .Z(n3152) );
  XOR U4954 ( .A(DB[92]), .B(DB[77]), .Z(n3154) );
  AND U4955 ( .A(n490), .B(n3155), .Z(n3153) );
  XOR U4956 ( .A(n3156), .B(n3157), .Z(n3155) );
  XOR U4957 ( .A(DB[77]), .B(DB[62]), .Z(n3157) );
  AND U4958 ( .A(n494), .B(n3158), .Z(n3156) );
  XOR U4959 ( .A(n3159), .B(n3160), .Z(n3158) );
  XOR U4960 ( .A(DB[62]), .B(DB[47]), .Z(n3160) );
  AND U4961 ( .A(n498), .B(n3161), .Z(n3159) );
  XOR U4962 ( .A(n3162), .B(n3163), .Z(n3161) );
  XOR U4963 ( .A(DB[47]), .B(DB[32]), .Z(n3163) );
  AND U4964 ( .A(n502), .B(n3164), .Z(n3162) );
  XOR U4965 ( .A(n3165), .B(n3166), .Z(n3164) );
  XOR U4966 ( .A(DB[32]), .B(DB[17]), .Z(n3166) );
  AND U4967 ( .A(n506), .B(n3167), .Z(n3165) );
  XOR U4968 ( .A(DB[2]), .B(DB[17]), .Z(n3167) );
  XOR U4969 ( .A(DB[1906]), .B(n3168), .Z(min_val_out[1]) );
  AND U4970 ( .A(n2), .B(n3169), .Z(n3168) );
  XOR U4971 ( .A(n3170), .B(n3171), .Z(n3169) );
  XOR U4972 ( .A(DB[1906]), .B(DB[1891]), .Z(n3171) );
  AND U4973 ( .A(n6), .B(n3172), .Z(n3170) );
  XOR U4974 ( .A(n3173), .B(n3174), .Z(n3172) );
  XOR U4975 ( .A(DB[1891]), .B(DB[1876]), .Z(n3174) );
  AND U4976 ( .A(n10), .B(n3175), .Z(n3173) );
  XOR U4977 ( .A(n3176), .B(n3177), .Z(n3175) );
  XOR U4978 ( .A(DB[1876]), .B(DB[1861]), .Z(n3177) );
  AND U4979 ( .A(n14), .B(n3178), .Z(n3176) );
  XOR U4980 ( .A(n3179), .B(n3180), .Z(n3178) );
  XOR U4981 ( .A(DB[1861]), .B(DB[1846]), .Z(n3180) );
  AND U4982 ( .A(n18), .B(n3181), .Z(n3179) );
  XOR U4983 ( .A(n3182), .B(n3183), .Z(n3181) );
  XOR U4984 ( .A(DB[1846]), .B(DB[1831]), .Z(n3183) );
  AND U4985 ( .A(n22), .B(n3184), .Z(n3182) );
  XOR U4986 ( .A(n3185), .B(n3186), .Z(n3184) );
  XOR U4987 ( .A(DB[1831]), .B(DB[1816]), .Z(n3186) );
  AND U4988 ( .A(n26), .B(n3187), .Z(n3185) );
  XOR U4989 ( .A(n3188), .B(n3189), .Z(n3187) );
  XOR U4990 ( .A(DB[1816]), .B(DB[1801]), .Z(n3189) );
  AND U4991 ( .A(n30), .B(n3190), .Z(n3188) );
  XOR U4992 ( .A(n3191), .B(n3192), .Z(n3190) );
  XOR U4993 ( .A(DB[1801]), .B(DB[1786]), .Z(n3192) );
  AND U4994 ( .A(n34), .B(n3193), .Z(n3191) );
  XOR U4995 ( .A(n3194), .B(n3195), .Z(n3193) );
  XOR U4996 ( .A(DB[1786]), .B(DB[1771]), .Z(n3195) );
  AND U4997 ( .A(n38), .B(n3196), .Z(n3194) );
  XOR U4998 ( .A(n3197), .B(n3198), .Z(n3196) );
  XOR U4999 ( .A(DB[1771]), .B(DB[1756]), .Z(n3198) );
  AND U5000 ( .A(n42), .B(n3199), .Z(n3197) );
  XOR U5001 ( .A(n3200), .B(n3201), .Z(n3199) );
  XOR U5002 ( .A(DB[1756]), .B(DB[1741]), .Z(n3201) );
  AND U5003 ( .A(n46), .B(n3202), .Z(n3200) );
  XOR U5004 ( .A(n3203), .B(n3204), .Z(n3202) );
  XOR U5005 ( .A(DB[1741]), .B(DB[1726]), .Z(n3204) );
  AND U5006 ( .A(n50), .B(n3205), .Z(n3203) );
  XOR U5007 ( .A(n3206), .B(n3207), .Z(n3205) );
  XOR U5008 ( .A(DB[1726]), .B(DB[1711]), .Z(n3207) );
  AND U5009 ( .A(n54), .B(n3208), .Z(n3206) );
  XOR U5010 ( .A(n3209), .B(n3210), .Z(n3208) );
  XOR U5011 ( .A(DB[1711]), .B(DB[1696]), .Z(n3210) );
  AND U5012 ( .A(n58), .B(n3211), .Z(n3209) );
  XOR U5013 ( .A(n3212), .B(n3213), .Z(n3211) );
  XOR U5014 ( .A(DB[1696]), .B(DB[1681]), .Z(n3213) );
  AND U5015 ( .A(n62), .B(n3214), .Z(n3212) );
  XOR U5016 ( .A(n3215), .B(n3216), .Z(n3214) );
  XOR U5017 ( .A(DB[1681]), .B(DB[1666]), .Z(n3216) );
  AND U5018 ( .A(n66), .B(n3217), .Z(n3215) );
  XOR U5019 ( .A(n3218), .B(n3219), .Z(n3217) );
  XOR U5020 ( .A(DB[1666]), .B(DB[1651]), .Z(n3219) );
  AND U5021 ( .A(n70), .B(n3220), .Z(n3218) );
  XOR U5022 ( .A(n3221), .B(n3222), .Z(n3220) );
  XOR U5023 ( .A(DB[1651]), .B(DB[1636]), .Z(n3222) );
  AND U5024 ( .A(n74), .B(n3223), .Z(n3221) );
  XOR U5025 ( .A(n3224), .B(n3225), .Z(n3223) );
  XOR U5026 ( .A(DB[1636]), .B(DB[1621]), .Z(n3225) );
  AND U5027 ( .A(n78), .B(n3226), .Z(n3224) );
  XOR U5028 ( .A(n3227), .B(n3228), .Z(n3226) );
  XOR U5029 ( .A(DB[1621]), .B(DB[1606]), .Z(n3228) );
  AND U5030 ( .A(n82), .B(n3229), .Z(n3227) );
  XOR U5031 ( .A(n3230), .B(n3231), .Z(n3229) );
  XOR U5032 ( .A(DB[1606]), .B(DB[1591]), .Z(n3231) );
  AND U5033 ( .A(n86), .B(n3232), .Z(n3230) );
  XOR U5034 ( .A(n3233), .B(n3234), .Z(n3232) );
  XOR U5035 ( .A(DB[1591]), .B(DB[1576]), .Z(n3234) );
  AND U5036 ( .A(n90), .B(n3235), .Z(n3233) );
  XOR U5037 ( .A(n3236), .B(n3237), .Z(n3235) );
  XOR U5038 ( .A(DB[1576]), .B(DB[1561]), .Z(n3237) );
  AND U5039 ( .A(n94), .B(n3238), .Z(n3236) );
  XOR U5040 ( .A(n3239), .B(n3240), .Z(n3238) );
  XOR U5041 ( .A(DB[1561]), .B(DB[1546]), .Z(n3240) );
  AND U5042 ( .A(n98), .B(n3241), .Z(n3239) );
  XOR U5043 ( .A(n3242), .B(n3243), .Z(n3241) );
  XOR U5044 ( .A(DB[1546]), .B(DB[1531]), .Z(n3243) );
  AND U5045 ( .A(n102), .B(n3244), .Z(n3242) );
  XOR U5046 ( .A(n3245), .B(n3246), .Z(n3244) );
  XOR U5047 ( .A(DB[1531]), .B(DB[1516]), .Z(n3246) );
  AND U5048 ( .A(n106), .B(n3247), .Z(n3245) );
  XOR U5049 ( .A(n3248), .B(n3249), .Z(n3247) );
  XOR U5050 ( .A(DB[1516]), .B(DB[1501]), .Z(n3249) );
  AND U5051 ( .A(n110), .B(n3250), .Z(n3248) );
  XOR U5052 ( .A(n3251), .B(n3252), .Z(n3250) );
  XOR U5053 ( .A(DB[1501]), .B(DB[1486]), .Z(n3252) );
  AND U5054 ( .A(n114), .B(n3253), .Z(n3251) );
  XOR U5055 ( .A(n3254), .B(n3255), .Z(n3253) );
  XOR U5056 ( .A(DB[1486]), .B(DB[1471]), .Z(n3255) );
  AND U5057 ( .A(n118), .B(n3256), .Z(n3254) );
  XOR U5058 ( .A(n3257), .B(n3258), .Z(n3256) );
  XOR U5059 ( .A(DB[1471]), .B(DB[1456]), .Z(n3258) );
  AND U5060 ( .A(n122), .B(n3259), .Z(n3257) );
  XOR U5061 ( .A(n3260), .B(n3261), .Z(n3259) );
  XOR U5062 ( .A(DB[1456]), .B(DB[1441]), .Z(n3261) );
  AND U5063 ( .A(n126), .B(n3262), .Z(n3260) );
  XOR U5064 ( .A(n3263), .B(n3264), .Z(n3262) );
  XOR U5065 ( .A(DB[1441]), .B(DB[1426]), .Z(n3264) );
  AND U5066 ( .A(n130), .B(n3265), .Z(n3263) );
  XOR U5067 ( .A(n3266), .B(n3267), .Z(n3265) );
  XOR U5068 ( .A(DB[1426]), .B(DB[1411]), .Z(n3267) );
  AND U5069 ( .A(n134), .B(n3268), .Z(n3266) );
  XOR U5070 ( .A(n3269), .B(n3270), .Z(n3268) );
  XOR U5071 ( .A(DB[1411]), .B(DB[1396]), .Z(n3270) );
  AND U5072 ( .A(n138), .B(n3271), .Z(n3269) );
  XOR U5073 ( .A(n3272), .B(n3273), .Z(n3271) );
  XOR U5074 ( .A(DB[1396]), .B(DB[1381]), .Z(n3273) );
  AND U5075 ( .A(n142), .B(n3274), .Z(n3272) );
  XOR U5076 ( .A(n3275), .B(n3276), .Z(n3274) );
  XOR U5077 ( .A(DB[1381]), .B(DB[1366]), .Z(n3276) );
  AND U5078 ( .A(n146), .B(n3277), .Z(n3275) );
  XOR U5079 ( .A(n3278), .B(n3279), .Z(n3277) );
  XOR U5080 ( .A(DB[1366]), .B(DB[1351]), .Z(n3279) );
  AND U5081 ( .A(n150), .B(n3280), .Z(n3278) );
  XOR U5082 ( .A(n3281), .B(n3282), .Z(n3280) );
  XOR U5083 ( .A(DB[1351]), .B(DB[1336]), .Z(n3282) );
  AND U5084 ( .A(n154), .B(n3283), .Z(n3281) );
  XOR U5085 ( .A(n3284), .B(n3285), .Z(n3283) );
  XOR U5086 ( .A(DB[1336]), .B(DB[1321]), .Z(n3285) );
  AND U5087 ( .A(n158), .B(n3286), .Z(n3284) );
  XOR U5088 ( .A(n3287), .B(n3288), .Z(n3286) );
  XOR U5089 ( .A(DB[1321]), .B(DB[1306]), .Z(n3288) );
  AND U5090 ( .A(n162), .B(n3289), .Z(n3287) );
  XOR U5091 ( .A(n3290), .B(n3291), .Z(n3289) );
  XOR U5092 ( .A(DB[1306]), .B(DB[1291]), .Z(n3291) );
  AND U5093 ( .A(n166), .B(n3292), .Z(n3290) );
  XOR U5094 ( .A(n3293), .B(n3294), .Z(n3292) );
  XOR U5095 ( .A(DB[1291]), .B(DB[1276]), .Z(n3294) );
  AND U5096 ( .A(n170), .B(n3295), .Z(n3293) );
  XOR U5097 ( .A(n3296), .B(n3297), .Z(n3295) );
  XOR U5098 ( .A(DB[1276]), .B(DB[1261]), .Z(n3297) );
  AND U5099 ( .A(n174), .B(n3298), .Z(n3296) );
  XOR U5100 ( .A(n3299), .B(n3300), .Z(n3298) );
  XOR U5101 ( .A(DB[1261]), .B(DB[1246]), .Z(n3300) );
  AND U5102 ( .A(n178), .B(n3301), .Z(n3299) );
  XOR U5103 ( .A(n3302), .B(n3303), .Z(n3301) );
  XOR U5104 ( .A(DB[1246]), .B(DB[1231]), .Z(n3303) );
  AND U5105 ( .A(n182), .B(n3304), .Z(n3302) );
  XOR U5106 ( .A(n3305), .B(n3306), .Z(n3304) );
  XOR U5107 ( .A(DB[1231]), .B(DB[1216]), .Z(n3306) );
  AND U5108 ( .A(n186), .B(n3307), .Z(n3305) );
  XOR U5109 ( .A(n3308), .B(n3309), .Z(n3307) );
  XOR U5110 ( .A(DB[1216]), .B(DB[1201]), .Z(n3309) );
  AND U5111 ( .A(n190), .B(n3310), .Z(n3308) );
  XOR U5112 ( .A(n3311), .B(n3312), .Z(n3310) );
  XOR U5113 ( .A(DB[1201]), .B(DB[1186]), .Z(n3312) );
  AND U5114 ( .A(n194), .B(n3313), .Z(n3311) );
  XOR U5115 ( .A(n3314), .B(n3315), .Z(n3313) );
  XOR U5116 ( .A(DB[1186]), .B(DB[1171]), .Z(n3315) );
  AND U5117 ( .A(n198), .B(n3316), .Z(n3314) );
  XOR U5118 ( .A(n3317), .B(n3318), .Z(n3316) );
  XOR U5119 ( .A(DB[1171]), .B(DB[1156]), .Z(n3318) );
  AND U5120 ( .A(n202), .B(n3319), .Z(n3317) );
  XOR U5121 ( .A(n3320), .B(n3321), .Z(n3319) );
  XOR U5122 ( .A(DB[1156]), .B(DB[1141]), .Z(n3321) );
  AND U5123 ( .A(n206), .B(n3322), .Z(n3320) );
  XOR U5124 ( .A(n3323), .B(n3324), .Z(n3322) );
  XOR U5125 ( .A(DB[1141]), .B(DB[1126]), .Z(n3324) );
  AND U5126 ( .A(n210), .B(n3325), .Z(n3323) );
  XOR U5127 ( .A(n3326), .B(n3327), .Z(n3325) );
  XOR U5128 ( .A(DB[1126]), .B(DB[1111]), .Z(n3327) );
  AND U5129 ( .A(n214), .B(n3328), .Z(n3326) );
  XOR U5130 ( .A(n3329), .B(n3330), .Z(n3328) );
  XOR U5131 ( .A(DB[1111]), .B(DB[1096]), .Z(n3330) );
  AND U5132 ( .A(n218), .B(n3331), .Z(n3329) );
  XOR U5133 ( .A(n3332), .B(n3333), .Z(n3331) );
  XOR U5134 ( .A(DB[1096]), .B(DB[1081]), .Z(n3333) );
  AND U5135 ( .A(n222), .B(n3334), .Z(n3332) );
  XOR U5136 ( .A(n3335), .B(n3336), .Z(n3334) );
  XOR U5137 ( .A(DB[1081]), .B(DB[1066]), .Z(n3336) );
  AND U5138 ( .A(n226), .B(n3337), .Z(n3335) );
  XOR U5139 ( .A(n3338), .B(n3339), .Z(n3337) );
  XOR U5140 ( .A(DB[1066]), .B(DB[1051]), .Z(n3339) );
  AND U5141 ( .A(n230), .B(n3340), .Z(n3338) );
  XOR U5142 ( .A(n3341), .B(n3342), .Z(n3340) );
  XOR U5143 ( .A(DB[1051]), .B(DB[1036]), .Z(n3342) );
  AND U5144 ( .A(n234), .B(n3343), .Z(n3341) );
  XOR U5145 ( .A(n3344), .B(n3345), .Z(n3343) );
  XOR U5146 ( .A(DB[1036]), .B(DB[1021]), .Z(n3345) );
  AND U5147 ( .A(n238), .B(n3346), .Z(n3344) );
  XOR U5148 ( .A(n3347), .B(n3348), .Z(n3346) );
  XOR U5149 ( .A(DB[1021]), .B(DB[1006]), .Z(n3348) );
  AND U5150 ( .A(n242), .B(n3349), .Z(n3347) );
  XOR U5151 ( .A(n3350), .B(n3351), .Z(n3349) );
  XOR U5152 ( .A(DB[991]), .B(DB[1006]), .Z(n3351) );
  AND U5153 ( .A(n246), .B(n3352), .Z(n3350) );
  XOR U5154 ( .A(n3353), .B(n3354), .Z(n3352) );
  XOR U5155 ( .A(DB[991]), .B(DB[976]), .Z(n3354) );
  AND U5156 ( .A(n250), .B(n3355), .Z(n3353) );
  XOR U5157 ( .A(n3356), .B(n3357), .Z(n3355) );
  XOR U5158 ( .A(DB[976]), .B(DB[961]), .Z(n3357) );
  AND U5159 ( .A(n254), .B(n3358), .Z(n3356) );
  XOR U5160 ( .A(n3359), .B(n3360), .Z(n3358) );
  XOR U5161 ( .A(DB[961]), .B(DB[946]), .Z(n3360) );
  AND U5162 ( .A(n258), .B(n3361), .Z(n3359) );
  XOR U5163 ( .A(n3362), .B(n3363), .Z(n3361) );
  XOR U5164 ( .A(DB[946]), .B(DB[931]), .Z(n3363) );
  AND U5165 ( .A(n262), .B(n3364), .Z(n3362) );
  XOR U5166 ( .A(n3365), .B(n3366), .Z(n3364) );
  XOR U5167 ( .A(DB[931]), .B(DB[916]), .Z(n3366) );
  AND U5168 ( .A(n266), .B(n3367), .Z(n3365) );
  XOR U5169 ( .A(n3368), .B(n3369), .Z(n3367) );
  XOR U5170 ( .A(DB[916]), .B(DB[901]), .Z(n3369) );
  AND U5171 ( .A(n270), .B(n3370), .Z(n3368) );
  XOR U5172 ( .A(n3371), .B(n3372), .Z(n3370) );
  XOR U5173 ( .A(DB[901]), .B(DB[886]), .Z(n3372) );
  AND U5174 ( .A(n274), .B(n3373), .Z(n3371) );
  XOR U5175 ( .A(n3374), .B(n3375), .Z(n3373) );
  XOR U5176 ( .A(DB[886]), .B(DB[871]), .Z(n3375) );
  AND U5177 ( .A(n278), .B(n3376), .Z(n3374) );
  XOR U5178 ( .A(n3377), .B(n3378), .Z(n3376) );
  XOR U5179 ( .A(DB[871]), .B(DB[856]), .Z(n3378) );
  AND U5180 ( .A(n282), .B(n3379), .Z(n3377) );
  XOR U5181 ( .A(n3380), .B(n3381), .Z(n3379) );
  XOR U5182 ( .A(DB[856]), .B(DB[841]), .Z(n3381) );
  AND U5183 ( .A(n286), .B(n3382), .Z(n3380) );
  XOR U5184 ( .A(n3383), .B(n3384), .Z(n3382) );
  XOR U5185 ( .A(DB[841]), .B(DB[826]), .Z(n3384) );
  AND U5186 ( .A(n290), .B(n3385), .Z(n3383) );
  XOR U5187 ( .A(n3386), .B(n3387), .Z(n3385) );
  XOR U5188 ( .A(DB[826]), .B(DB[811]), .Z(n3387) );
  AND U5189 ( .A(n294), .B(n3388), .Z(n3386) );
  XOR U5190 ( .A(n3389), .B(n3390), .Z(n3388) );
  XOR U5191 ( .A(DB[811]), .B(DB[796]), .Z(n3390) );
  AND U5192 ( .A(n298), .B(n3391), .Z(n3389) );
  XOR U5193 ( .A(n3392), .B(n3393), .Z(n3391) );
  XOR U5194 ( .A(DB[796]), .B(DB[781]), .Z(n3393) );
  AND U5195 ( .A(n302), .B(n3394), .Z(n3392) );
  XOR U5196 ( .A(n3395), .B(n3396), .Z(n3394) );
  XOR U5197 ( .A(DB[781]), .B(DB[766]), .Z(n3396) );
  AND U5198 ( .A(n306), .B(n3397), .Z(n3395) );
  XOR U5199 ( .A(n3398), .B(n3399), .Z(n3397) );
  XOR U5200 ( .A(DB[766]), .B(DB[751]), .Z(n3399) );
  AND U5201 ( .A(n310), .B(n3400), .Z(n3398) );
  XOR U5202 ( .A(n3401), .B(n3402), .Z(n3400) );
  XOR U5203 ( .A(DB[751]), .B(DB[736]), .Z(n3402) );
  AND U5204 ( .A(n314), .B(n3403), .Z(n3401) );
  XOR U5205 ( .A(n3404), .B(n3405), .Z(n3403) );
  XOR U5206 ( .A(DB[736]), .B(DB[721]), .Z(n3405) );
  AND U5207 ( .A(n318), .B(n3406), .Z(n3404) );
  XOR U5208 ( .A(n3407), .B(n3408), .Z(n3406) );
  XOR U5209 ( .A(DB[721]), .B(DB[706]), .Z(n3408) );
  AND U5210 ( .A(n322), .B(n3409), .Z(n3407) );
  XOR U5211 ( .A(n3410), .B(n3411), .Z(n3409) );
  XOR U5212 ( .A(DB[706]), .B(DB[691]), .Z(n3411) );
  AND U5213 ( .A(n326), .B(n3412), .Z(n3410) );
  XOR U5214 ( .A(n3413), .B(n3414), .Z(n3412) );
  XOR U5215 ( .A(DB[691]), .B(DB[676]), .Z(n3414) );
  AND U5216 ( .A(n330), .B(n3415), .Z(n3413) );
  XOR U5217 ( .A(n3416), .B(n3417), .Z(n3415) );
  XOR U5218 ( .A(DB[676]), .B(DB[661]), .Z(n3417) );
  AND U5219 ( .A(n334), .B(n3418), .Z(n3416) );
  XOR U5220 ( .A(n3419), .B(n3420), .Z(n3418) );
  XOR U5221 ( .A(DB[661]), .B(DB[646]), .Z(n3420) );
  AND U5222 ( .A(n338), .B(n3421), .Z(n3419) );
  XOR U5223 ( .A(n3422), .B(n3423), .Z(n3421) );
  XOR U5224 ( .A(DB[646]), .B(DB[631]), .Z(n3423) );
  AND U5225 ( .A(n342), .B(n3424), .Z(n3422) );
  XOR U5226 ( .A(n3425), .B(n3426), .Z(n3424) );
  XOR U5227 ( .A(DB[631]), .B(DB[616]), .Z(n3426) );
  AND U5228 ( .A(n346), .B(n3427), .Z(n3425) );
  XOR U5229 ( .A(n3428), .B(n3429), .Z(n3427) );
  XOR U5230 ( .A(DB[616]), .B(DB[601]), .Z(n3429) );
  AND U5231 ( .A(n350), .B(n3430), .Z(n3428) );
  XOR U5232 ( .A(n3431), .B(n3432), .Z(n3430) );
  XOR U5233 ( .A(DB[601]), .B(DB[586]), .Z(n3432) );
  AND U5234 ( .A(n354), .B(n3433), .Z(n3431) );
  XOR U5235 ( .A(n3434), .B(n3435), .Z(n3433) );
  XOR U5236 ( .A(DB[586]), .B(DB[571]), .Z(n3435) );
  AND U5237 ( .A(n358), .B(n3436), .Z(n3434) );
  XOR U5238 ( .A(n3437), .B(n3438), .Z(n3436) );
  XOR U5239 ( .A(DB[571]), .B(DB[556]), .Z(n3438) );
  AND U5240 ( .A(n362), .B(n3439), .Z(n3437) );
  XOR U5241 ( .A(n3440), .B(n3441), .Z(n3439) );
  XOR U5242 ( .A(DB[556]), .B(DB[541]), .Z(n3441) );
  AND U5243 ( .A(n366), .B(n3442), .Z(n3440) );
  XOR U5244 ( .A(n3443), .B(n3444), .Z(n3442) );
  XOR U5245 ( .A(DB[541]), .B(DB[526]), .Z(n3444) );
  AND U5246 ( .A(n370), .B(n3445), .Z(n3443) );
  XOR U5247 ( .A(n3446), .B(n3447), .Z(n3445) );
  XOR U5248 ( .A(DB[526]), .B(DB[511]), .Z(n3447) );
  AND U5249 ( .A(n374), .B(n3448), .Z(n3446) );
  XOR U5250 ( .A(n3449), .B(n3450), .Z(n3448) );
  XOR U5251 ( .A(DB[511]), .B(DB[496]), .Z(n3450) );
  AND U5252 ( .A(n378), .B(n3451), .Z(n3449) );
  XOR U5253 ( .A(n3452), .B(n3453), .Z(n3451) );
  XOR U5254 ( .A(DB[496]), .B(DB[481]), .Z(n3453) );
  AND U5255 ( .A(n382), .B(n3454), .Z(n3452) );
  XOR U5256 ( .A(n3455), .B(n3456), .Z(n3454) );
  XOR U5257 ( .A(DB[481]), .B(DB[466]), .Z(n3456) );
  AND U5258 ( .A(n386), .B(n3457), .Z(n3455) );
  XOR U5259 ( .A(n3458), .B(n3459), .Z(n3457) );
  XOR U5260 ( .A(DB[466]), .B(DB[451]), .Z(n3459) );
  AND U5261 ( .A(n390), .B(n3460), .Z(n3458) );
  XOR U5262 ( .A(n3461), .B(n3462), .Z(n3460) );
  XOR U5263 ( .A(DB[451]), .B(DB[436]), .Z(n3462) );
  AND U5264 ( .A(n394), .B(n3463), .Z(n3461) );
  XOR U5265 ( .A(n3464), .B(n3465), .Z(n3463) );
  XOR U5266 ( .A(DB[436]), .B(DB[421]), .Z(n3465) );
  AND U5267 ( .A(n398), .B(n3466), .Z(n3464) );
  XOR U5268 ( .A(n3467), .B(n3468), .Z(n3466) );
  XOR U5269 ( .A(DB[421]), .B(DB[406]), .Z(n3468) );
  AND U5270 ( .A(n402), .B(n3469), .Z(n3467) );
  XOR U5271 ( .A(n3470), .B(n3471), .Z(n3469) );
  XOR U5272 ( .A(DB[406]), .B(DB[391]), .Z(n3471) );
  AND U5273 ( .A(n406), .B(n3472), .Z(n3470) );
  XOR U5274 ( .A(n3473), .B(n3474), .Z(n3472) );
  XOR U5275 ( .A(DB[391]), .B(DB[376]), .Z(n3474) );
  AND U5276 ( .A(n410), .B(n3475), .Z(n3473) );
  XOR U5277 ( .A(n3476), .B(n3477), .Z(n3475) );
  XOR U5278 ( .A(DB[376]), .B(DB[361]), .Z(n3477) );
  AND U5279 ( .A(n414), .B(n3478), .Z(n3476) );
  XOR U5280 ( .A(n3479), .B(n3480), .Z(n3478) );
  XOR U5281 ( .A(DB[361]), .B(DB[346]), .Z(n3480) );
  AND U5282 ( .A(n418), .B(n3481), .Z(n3479) );
  XOR U5283 ( .A(n3482), .B(n3483), .Z(n3481) );
  XOR U5284 ( .A(DB[346]), .B(DB[331]), .Z(n3483) );
  AND U5285 ( .A(n422), .B(n3484), .Z(n3482) );
  XOR U5286 ( .A(n3485), .B(n3486), .Z(n3484) );
  XOR U5287 ( .A(DB[331]), .B(DB[316]), .Z(n3486) );
  AND U5288 ( .A(n426), .B(n3487), .Z(n3485) );
  XOR U5289 ( .A(n3488), .B(n3489), .Z(n3487) );
  XOR U5290 ( .A(DB[316]), .B(DB[301]), .Z(n3489) );
  AND U5291 ( .A(n430), .B(n3490), .Z(n3488) );
  XOR U5292 ( .A(n3491), .B(n3492), .Z(n3490) );
  XOR U5293 ( .A(DB[301]), .B(DB[286]), .Z(n3492) );
  AND U5294 ( .A(n434), .B(n3493), .Z(n3491) );
  XOR U5295 ( .A(n3494), .B(n3495), .Z(n3493) );
  XOR U5296 ( .A(DB[286]), .B(DB[271]), .Z(n3495) );
  AND U5297 ( .A(n438), .B(n3496), .Z(n3494) );
  XOR U5298 ( .A(n3497), .B(n3498), .Z(n3496) );
  XOR U5299 ( .A(DB[271]), .B(DB[256]), .Z(n3498) );
  AND U5300 ( .A(n442), .B(n3499), .Z(n3497) );
  XOR U5301 ( .A(n3500), .B(n3501), .Z(n3499) );
  XOR U5302 ( .A(DB[256]), .B(DB[241]), .Z(n3501) );
  AND U5303 ( .A(n446), .B(n3502), .Z(n3500) );
  XOR U5304 ( .A(n3503), .B(n3504), .Z(n3502) );
  XOR U5305 ( .A(DB[241]), .B(DB[226]), .Z(n3504) );
  AND U5306 ( .A(n450), .B(n3505), .Z(n3503) );
  XOR U5307 ( .A(n3506), .B(n3507), .Z(n3505) );
  XOR U5308 ( .A(DB[226]), .B(DB[211]), .Z(n3507) );
  AND U5309 ( .A(n454), .B(n3508), .Z(n3506) );
  XOR U5310 ( .A(n3509), .B(n3510), .Z(n3508) );
  XOR U5311 ( .A(DB[211]), .B(DB[196]), .Z(n3510) );
  AND U5312 ( .A(n458), .B(n3511), .Z(n3509) );
  XOR U5313 ( .A(n3512), .B(n3513), .Z(n3511) );
  XOR U5314 ( .A(DB[196]), .B(DB[181]), .Z(n3513) );
  AND U5315 ( .A(n462), .B(n3514), .Z(n3512) );
  XOR U5316 ( .A(n3515), .B(n3516), .Z(n3514) );
  XOR U5317 ( .A(DB[181]), .B(DB[166]), .Z(n3516) );
  AND U5318 ( .A(n466), .B(n3517), .Z(n3515) );
  XOR U5319 ( .A(n3518), .B(n3519), .Z(n3517) );
  XOR U5320 ( .A(DB[166]), .B(DB[151]), .Z(n3519) );
  AND U5321 ( .A(n470), .B(n3520), .Z(n3518) );
  XOR U5322 ( .A(n3521), .B(n3522), .Z(n3520) );
  XOR U5323 ( .A(DB[151]), .B(DB[136]), .Z(n3522) );
  AND U5324 ( .A(n474), .B(n3523), .Z(n3521) );
  XOR U5325 ( .A(n3524), .B(n3525), .Z(n3523) );
  XOR U5326 ( .A(DB[136]), .B(DB[121]), .Z(n3525) );
  AND U5327 ( .A(n478), .B(n3526), .Z(n3524) );
  XOR U5328 ( .A(n3527), .B(n3528), .Z(n3526) );
  XOR U5329 ( .A(DB[121]), .B(DB[106]), .Z(n3528) );
  AND U5330 ( .A(n482), .B(n3529), .Z(n3527) );
  XOR U5331 ( .A(n3530), .B(n3531), .Z(n3529) );
  XOR U5332 ( .A(DB[91]), .B(DB[106]), .Z(n3531) );
  AND U5333 ( .A(n486), .B(n3532), .Z(n3530) );
  XOR U5334 ( .A(n3533), .B(n3534), .Z(n3532) );
  XOR U5335 ( .A(DB[91]), .B(DB[76]), .Z(n3534) );
  AND U5336 ( .A(n490), .B(n3535), .Z(n3533) );
  XOR U5337 ( .A(n3536), .B(n3537), .Z(n3535) );
  XOR U5338 ( .A(DB[76]), .B(DB[61]), .Z(n3537) );
  AND U5339 ( .A(n494), .B(n3538), .Z(n3536) );
  XOR U5340 ( .A(n3539), .B(n3540), .Z(n3538) );
  XOR U5341 ( .A(DB[61]), .B(DB[46]), .Z(n3540) );
  AND U5342 ( .A(n498), .B(n3541), .Z(n3539) );
  XOR U5343 ( .A(n3542), .B(n3543), .Z(n3541) );
  XOR U5344 ( .A(DB[46]), .B(DB[31]), .Z(n3543) );
  AND U5345 ( .A(n502), .B(n3544), .Z(n3542) );
  XOR U5346 ( .A(n3545), .B(n3546), .Z(n3544) );
  XOR U5347 ( .A(DB[31]), .B(DB[16]), .Z(n3546) );
  AND U5348 ( .A(n506), .B(n3547), .Z(n3545) );
  XOR U5349 ( .A(DB[1]), .B(DB[16]), .Z(n3547) );
  XOR U5350 ( .A(DB[1919]), .B(n3548), .Z(min_val_out[14]) );
  AND U5351 ( .A(n2), .B(n3549), .Z(n3548) );
  XOR U5352 ( .A(n3550), .B(n3551), .Z(n3549) );
  XOR U5353 ( .A(DB[1919]), .B(DB[1904]), .Z(n3551) );
  AND U5354 ( .A(n6), .B(n3552), .Z(n3550) );
  XOR U5355 ( .A(n3553), .B(n3554), .Z(n3552) );
  XOR U5356 ( .A(DB[1904]), .B(DB[1889]), .Z(n3554) );
  AND U5357 ( .A(n10), .B(n3555), .Z(n3553) );
  XOR U5358 ( .A(n3556), .B(n3557), .Z(n3555) );
  XOR U5359 ( .A(DB[1889]), .B(DB[1874]), .Z(n3557) );
  AND U5360 ( .A(n14), .B(n3558), .Z(n3556) );
  XOR U5361 ( .A(n3559), .B(n3560), .Z(n3558) );
  XOR U5362 ( .A(DB[1874]), .B(DB[1859]), .Z(n3560) );
  AND U5363 ( .A(n18), .B(n3561), .Z(n3559) );
  XOR U5364 ( .A(n3562), .B(n3563), .Z(n3561) );
  XOR U5365 ( .A(DB[1859]), .B(DB[1844]), .Z(n3563) );
  AND U5366 ( .A(n22), .B(n3564), .Z(n3562) );
  XOR U5367 ( .A(n3565), .B(n3566), .Z(n3564) );
  XOR U5368 ( .A(DB[1844]), .B(DB[1829]), .Z(n3566) );
  AND U5369 ( .A(n26), .B(n3567), .Z(n3565) );
  XOR U5370 ( .A(n3568), .B(n3569), .Z(n3567) );
  XOR U5371 ( .A(DB[1829]), .B(DB[1814]), .Z(n3569) );
  AND U5372 ( .A(n30), .B(n3570), .Z(n3568) );
  XOR U5373 ( .A(n3571), .B(n3572), .Z(n3570) );
  XOR U5374 ( .A(DB[1814]), .B(DB[1799]), .Z(n3572) );
  AND U5375 ( .A(n34), .B(n3573), .Z(n3571) );
  XOR U5376 ( .A(n3574), .B(n3575), .Z(n3573) );
  XOR U5377 ( .A(DB[1799]), .B(DB[1784]), .Z(n3575) );
  AND U5378 ( .A(n38), .B(n3576), .Z(n3574) );
  XOR U5379 ( .A(n3577), .B(n3578), .Z(n3576) );
  XOR U5380 ( .A(DB[1784]), .B(DB[1769]), .Z(n3578) );
  AND U5381 ( .A(n42), .B(n3579), .Z(n3577) );
  XOR U5382 ( .A(n3580), .B(n3581), .Z(n3579) );
  XOR U5383 ( .A(DB[1769]), .B(DB[1754]), .Z(n3581) );
  AND U5384 ( .A(n46), .B(n3582), .Z(n3580) );
  XOR U5385 ( .A(n3583), .B(n3584), .Z(n3582) );
  XOR U5386 ( .A(DB[1754]), .B(DB[1739]), .Z(n3584) );
  AND U5387 ( .A(n50), .B(n3585), .Z(n3583) );
  XOR U5388 ( .A(n3586), .B(n3587), .Z(n3585) );
  XOR U5389 ( .A(DB[1739]), .B(DB[1724]), .Z(n3587) );
  AND U5390 ( .A(n54), .B(n3588), .Z(n3586) );
  XOR U5391 ( .A(n3589), .B(n3590), .Z(n3588) );
  XOR U5392 ( .A(DB[1724]), .B(DB[1709]), .Z(n3590) );
  AND U5393 ( .A(n58), .B(n3591), .Z(n3589) );
  XOR U5394 ( .A(n3592), .B(n3593), .Z(n3591) );
  XOR U5395 ( .A(DB[1709]), .B(DB[1694]), .Z(n3593) );
  AND U5396 ( .A(n62), .B(n3594), .Z(n3592) );
  XOR U5397 ( .A(n3595), .B(n3596), .Z(n3594) );
  XOR U5398 ( .A(DB[1694]), .B(DB[1679]), .Z(n3596) );
  AND U5399 ( .A(n66), .B(n3597), .Z(n3595) );
  XOR U5400 ( .A(n3598), .B(n3599), .Z(n3597) );
  XOR U5401 ( .A(DB[1679]), .B(DB[1664]), .Z(n3599) );
  AND U5402 ( .A(n70), .B(n3600), .Z(n3598) );
  XOR U5403 ( .A(n3601), .B(n3602), .Z(n3600) );
  XOR U5404 ( .A(DB[1664]), .B(DB[1649]), .Z(n3602) );
  AND U5405 ( .A(n74), .B(n3603), .Z(n3601) );
  XOR U5406 ( .A(n3604), .B(n3605), .Z(n3603) );
  XOR U5407 ( .A(DB[1649]), .B(DB[1634]), .Z(n3605) );
  AND U5408 ( .A(n78), .B(n3606), .Z(n3604) );
  XOR U5409 ( .A(n3607), .B(n3608), .Z(n3606) );
  XOR U5410 ( .A(DB[1634]), .B(DB[1619]), .Z(n3608) );
  AND U5411 ( .A(n82), .B(n3609), .Z(n3607) );
  XOR U5412 ( .A(n3610), .B(n3611), .Z(n3609) );
  XOR U5413 ( .A(DB[1619]), .B(DB[1604]), .Z(n3611) );
  AND U5414 ( .A(n86), .B(n3612), .Z(n3610) );
  XOR U5415 ( .A(n3613), .B(n3614), .Z(n3612) );
  XOR U5416 ( .A(DB[1604]), .B(DB[1589]), .Z(n3614) );
  AND U5417 ( .A(n90), .B(n3615), .Z(n3613) );
  XOR U5418 ( .A(n3616), .B(n3617), .Z(n3615) );
  XOR U5419 ( .A(DB[1589]), .B(DB[1574]), .Z(n3617) );
  AND U5420 ( .A(n94), .B(n3618), .Z(n3616) );
  XOR U5421 ( .A(n3619), .B(n3620), .Z(n3618) );
  XOR U5422 ( .A(DB[1574]), .B(DB[1559]), .Z(n3620) );
  AND U5423 ( .A(n98), .B(n3621), .Z(n3619) );
  XOR U5424 ( .A(n3622), .B(n3623), .Z(n3621) );
  XOR U5425 ( .A(DB[1559]), .B(DB[1544]), .Z(n3623) );
  AND U5426 ( .A(n102), .B(n3624), .Z(n3622) );
  XOR U5427 ( .A(n3625), .B(n3626), .Z(n3624) );
  XOR U5428 ( .A(DB[1544]), .B(DB[1529]), .Z(n3626) );
  AND U5429 ( .A(n106), .B(n3627), .Z(n3625) );
  XOR U5430 ( .A(n3628), .B(n3629), .Z(n3627) );
  XOR U5431 ( .A(DB[1529]), .B(DB[1514]), .Z(n3629) );
  AND U5432 ( .A(n110), .B(n3630), .Z(n3628) );
  XOR U5433 ( .A(n3631), .B(n3632), .Z(n3630) );
  XOR U5434 ( .A(DB[1514]), .B(DB[1499]), .Z(n3632) );
  AND U5435 ( .A(n114), .B(n3633), .Z(n3631) );
  XOR U5436 ( .A(n3634), .B(n3635), .Z(n3633) );
  XOR U5437 ( .A(DB[1499]), .B(DB[1484]), .Z(n3635) );
  AND U5438 ( .A(n118), .B(n3636), .Z(n3634) );
  XOR U5439 ( .A(n3637), .B(n3638), .Z(n3636) );
  XOR U5440 ( .A(DB[1484]), .B(DB[1469]), .Z(n3638) );
  AND U5441 ( .A(n122), .B(n3639), .Z(n3637) );
  XOR U5442 ( .A(n3640), .B(n3641), .Z(n3639) );
  XOR U5443 ( .A(DB[1469]), .B(DB[1454]), .Z(n3641) );
  AND U5444 ( .A(n126), .B(n3642), .Z(n3640) );
  XOR U5445 ( .A(n3643), .B(n3644), .Z(n3642) );
  XOR U5446 ( .A(DB[1454]), .B(DB[1439]), .Z(n3644) );
  AND U5447 ( .A(n130), .B(n3645), .Z(n3643) );
  XOR U5448 ( .A(n3646), .B(n3647), .Z(n3645) );
  XOR U5449 ( .A(DB[1439]), .B(DB[1424]), .Z(n3647) );
  AND U5450 ( .A(n134), .B(n3648), .Z(n3646) );
  XOR U5451 ( .A(n3649), .B(n3650), .Z(n3648) );
  XOR U5452 ( .A(DB[1424]), .B(DB[1409]), .Z(n3650) );
  AND U5453 ( .A(n138), .B(n3651), .Z(n3649) );
  XOR U5454 ( .A(n3652), .B(n3653), .Z(n3651) );
  XOR U5455 ( .A(DB[1409]), .B(DB[1394]), .Z(n3653) );
  AND U5456 ( .A(n142), .B(n3654), .Z(n3652) );
  XOR U5457 ( .A(n3655), .B(n3656), .Z(n3654) );
  XOR U5458 ( .A(DB[1394]), .B(DB[1379]), .Z(n3656) );
  AND U5459 ( .A(n146), .B(n3657), .Z(n3655) );
  XOR U5460 ( .A(n3658), .B(n3659), .Z(n3657) );
  XOR U5461 ( .A(DB[1379]), .B(DB[1364]), .Z(n3659) );
  AND U5462 ( .A(n150), .B(n3660), .Z(n3658) );
  XOR U5463 ( .A(n3661), .B(n3662), .Z(n3660) );
  XOR U5464 ( .A(DB[1364]), .B(DB[1349]), .Z(n3662) );
  AND U5465 ( .A(n154), .B(n3663), .Z(n3661) );
  XOR U5466 ( .A(n3664), .B(n3665), .Z(n3663) );
  XOR U5467 ( .A(DB[1349]), .B(DB[1334]), .Z(n3665) );
  AND U5468 ( .A(n158), .B(n3666), .Z(n3664) );
  XOR U5469 ( .A(n3667), .B(n3668), .Z(n3666) );
  XOR U5470 ( .A(DB[1334]), .B(DB[1319]), .Z(n3668) );
  AND U5471 ( .A(n162), .B(n3669), .Z(n3667) );
  XOR U5472 ( .A(n3670), .B(n3671), .Z(n3669) );
  XOR U5473 ( .A(DB[1319]), .B(DB[1304]), .Z(n3671) );
  AND U5474 ( .A(n166), .B(n3672), .Z(n3670) );
  XOR U5475 ( .A(n3673), .B(n3674), .Z(n3672) );
  XOR U5476 ( .A(DB[1304]), .B(DB[1289]), .Z(n3674) );
  AND U5477 ( .A(n170), .B(n3675), .Z(n3673) );
  XOR U5478 ( .A(n3676), .B(n3677), .Z(n3675) );
  XOR U5479 ( .A(DB[1289]), .B(DB[1274]), .Z(n3677) );
  AND U5480 ( .A(n174), .B(n3678), .Z(n3676) );
  XOR U5481 ( .A(n3679), .B(n3680), .Z(n3678) );
  XOR U5482 ( .A(DB[1274]), .B(DB[1259]), .Z(n3680) );
  AND U5483 ( .A(n178), .B(n3681), .Z(n3679) );
  XOR U5484 ( .A(n3682), .B(n3683), .Z(n3681) );
  XOR U5485 ( .A(DB[1259]), .B(DB[1244]), .Z(n3683) );
  AND U5486 ( .A(n182), .B(n3684), .Z(n3682) );
  XOR U5487 ( .A(n3685), .B(n3686), .Z(n3684) );
  XOR U5488 ( .A(DB[1244]), .B(DB[1229]), .Z(n3686) );
  AND U5489 ( .A(n186), .B(n3687), .Z(n3685) );
  XOR U5490 ( .A(n3688), .B(n3689), .Z(n3687) );
  XOR U5491 ( .A(DB[1229]), .B(DB[1214]), .Z(n3689) );
  AND U5492 ( .A(n190), .B(n3690), .Z(n3688) );
  XOR U5493 ( .A(n3691), .B(n3692), .Z(n3690) );
  XOR U5494 ( .A(DB[1214]), .B(DB[1199]), .Z(n3692) );
  AND U5495 ( .A(n194), .B(n3693), .Z(n3691) );
  XOR U5496 ( .A(n3694), .B(n3695), .Z(n3693) );
  XOR U5497 ( .A(DB[1199]), .B(DB[1184]), .Z(n3695) );
  AND U5498 ( .A(n198), .B(n3696), .Z(n3694) );
  XOR U5499 ( .A(n3697), .B(n3698), .Z(n3696) );
  XOR U5500 ( .A(DB[1184]), .B(DB[1169]), .Z(n3698) );
  AND U5501 ( .A(n202), .B(n3699), .Z(n3697) );
  XOR U5502 ( .A(n3700), .B(n3701), .Z(n3699) );
  XOR U5503 ( .A(DB[1169]), .B(DB[1154]), .Z(n3701) );
  AND U5504 ( .A(n206), .B(n3702), .Z(n3700) );
  XOR U5505 ( .A(n3703), .B(n3704), .Z(n3702) );
  XOR U5506 ( .A(DB[1154]), .B(DB[1139]), .Z(n3704) );
  AND U5507 ( .A(n210), .B(n3705), .Z(n3703) );
  XOR U5508 ( .A(n3706), .B(n3707), .Z(n3705) );
  XOR U5509 ( .A(DB[1139]), .B(DB[1124]), .Z(n3707) );
  AND U5510 ( .A(n214), .B(n3708), .Z(n3706) );
  XOR U5511 ( .A(n3709), .B(n3710), .Z(n3708) );
  XOR U5512 ( .A(DB[1124]), .B(DB[1109]), .Z(n3710) );
  AND U5513 ( .A(n218), .B(n3711), .Z(n3709) );
  XOR U5514 ( .A(n3712), .B(n3713), .Z(n3711) );
  XOR U5515 ( .A(DB[1109]), .B(DB[1094]), .Z(n3713) );
  AND U5516 ( .A(n222), .B(n3714), .Z(n3712) );
  XOR U5517 ( .A(n3715), .B(n3716), .Z(n3714) );
  XOR U5518 ( .A(DB[1094]), .B(DB[1079]), .Z(n3716) );
  AND U5519 ( .A(n226), .B(n3717), .Z(n3715) );
  XOR U5520 ( .A(n3718), .B(n3719), .Z(n3717) );
  XOR U5521 ( .A(DB[1079]), .B(DB[1064]), .Z(n3719) );
  AND U5522 ( .A(n230), .B(n3720), .Z(n3718) );
  XOR U5523 ( .A(n3721), .B(n3722), .Z(n3720) );
  XOR U5524 ( .A(DB[1064]), .B(DB[1049]), .Z(n3722) );
  AND U5525 ( .A(n234), .B(n3723), .Z(n3721) );
  XOR U5526 ( .A(n3724), .B(n3725), .Z(n3723) );
  XOR U5527 ( .A(DB[1049]), .B(DB[1034]), .Z(n3725) );
  AND U5528 ( .A(n238), .B(n3726), .Z(n3724) );
  XOR U5529 ( .A(n3727), .B(n3728), .Z(n3726) );
  XOR U5530 ( .A(DB[1034]), .B(DB[1019]), .Z(n3728) );
  AND U5531 ( .A(n242), .B(n3729), .Z(n3727) );
  XOR U5532 ( .A(n3730), .B(n3731), .Z(n3729) );
  XOR U5533 ( .A(DB[1019]), .B(DB[1004]), .Z(n3731) );
  AND U5534 ( .A(n246), .B(n3732), .Z(n3730) );
  XOR U5535 ( .A(n3733), .B(n3734), .Z(n3732) );
  XOR U5536 ( .A(DB[989]), .B(DB[1004]), .Z(n3734) );
  AND U5537 ( .A(n250), .B(n3735), .Z(n3733) );
  XOR U5538 ( .A(n3736), .B(n3737), .Z(n3735) );
  XOR U5539 ( .A(DB[989]), .B(DB[974]), .Z(n3737) );
  AND U5540 ( .A(n254), .B(n3738), .Z(n3736) );
  XOR U5541 ( .A(n3739), .B(n3740), .Z(n3738) );
  XOR U5542 ( .A(DB[974]), .B(DB[959]), .Z(n3740) );
  AND U5543 ( .A(n258), .B(n3741), .Z(n3739) );
  XOR U5544 ( .A(n3742), .B(n3743), .Z(n3741) );
  XOR U5545 ( .A(DB[959]), .B(DB[944]), .Z(n3743) );
  AND U5546 ( .A(n262), .B(n3744), .Z(n3742) );
  XOR U5547 ( .A(n3745), .B(n3746), .Z(n3744) );
  XOR U5548 ( .A(DB[944]), .B(DB[929]), .Z(n3746) );
  AND U5549 ( .A(n266), .B(n3747), .Z(n3745) );
  XOR U5550 ( .A(n3748), .B(n3749), .Z(n3747) );
  XOR U5551 ( .A(DB[929]), .B(DB[914]), .Z(n3749) );
  AND U5552 ( .A(n270), .B(n3750), .Z(n3748) );
  XOR U5553 ( .A(n3751), .B(n3752), .Z(n3750) );
  XOR U5554 ( .A(DB[914]), .B(DB[899]), .Z(n3752) );
  AND U5555 ( .A(n274), .B(n3753), .Z(n3751) );
  XOR U5556 ( .A(n3754), .B(n3755), .Z(n3753) );
  XOR U5557 ( .A(DB[899]), .B(DB[884]), .Z(n3755) );
  AND U5558 ( .A(n278), .B(n3756), .Z(n3754) );
  XOR U5559 ( .A(n3757), .B(n3758), .Z(n3756) );
  XOR U5560 ( .A(DB[884]), .B(DB[869]), .Z(n3758) );
  AND U5561 ( .A(n282), .B(n3759), .Z(n3757) );
  XOR U5562 ( .A(n3760), .B(n3761), .Z(n3759) );
  XOR U5563 ( .A(DB[869]), .B(DB[854]), .Z(n3761) );
  AND U5564 ( .A(n286), .B(n3762), .Z(n3760) );
  XOR U5565 ( .A(n3763), .B(n3764), .Z(n3762) );
  XOR U5566 ( .A(DB[854]), .B(DB[839]), .Z(n3764) );
  AND U5567 ( .A(n290), .B(n3765), .Z(n3763) );
  XOR U5568 ( .A(n3766), .B(n3767), .Z(n3765) );
  XOR U5569 ( .A(DB[839]), .B(DB[824]), .Z(n3767) );
  AND U5570 ( .A(n294), .B(n3768), .Z(n3766) );
  XOR U5571 ( .A(n3769), .B(n3770), .Z(n3768) );
  XOR U5572 ( .A(DB[824]), .B(DB[809]), .Z(n3770) );
  AND U5573 ( .A(n298), .B(n3771), .Z(n3769) );
  XOR U5574 ( .A(n3772), .B(n3773), .Z(n3771) );
  XOR U5575 ( .A(DB[809]), .B(DB[794]), .Z(n3773) );
  AND U5576 ( .A(n302), .B(n3774), .Z(n3772) );
  XOR U5577 ( .A(n3775), .B(n3776), .Z(n3774) );
  XOR U5578 ( .A(DB[794]), .B(DB[779]), .Z(n3776) );
  AND U5579 ( .A(n306), .B(n3777), .Z(n3775) );
  XOR U5580 ( .A(n3778), .B(n3779), .Z(n3777) );
  XOR U5581 ( .A(DB[779]), .B(DB[764]), .Z(n3779) );
  AND U5582 ( .A(n310), .B(n3780), .Z(n3778) );
  XOR U5583 ( .A(n3781), .B(n3782), .Z(n3780) );
  XOR U5584 ( .A(DB[764]), .B(DB[749]), .Z(n3782) );
  AND U5585 ( .A(n314), .B(n3783), .Z(n3781) );
  XOR U5586 ( .A(n3784), .B(n3785), .Z(n3783) );
  XOR U5587 ( .A(DB[749]), .B(DB[734]), .Z(n3785) );
  AND U5588 ( .A(n318), .B(n3786), .Z(n3784) );
  XOR U5589 ( .A(n3787), .B(n3788), .Z(n3786) );
  XOR U5590 ( .A(DB[734]), .B(DB[719]), .Z(n3788) );
  AND U5591 ( .A(n322), .B(n3789), .Z(n3787) );
  XOR U5592 ( .A(n3790), .B(n3791), .Z(n3789) );
  XOR U5593 ( .A(DB[719]), .B(DB[704]), .Z(n3791) );
  AND U5594 ( .A(n326), .B(n3792), .Z(n3790) );
  XOR U5595 ( .A(n3793), .B(n3794), .Z(n3792) );
  XOR U5596 ( .A(DB[704]), .B(DB[689]), .Z(n3794) );
  AND U5597 ( .A(n330), .B(n3795), .Z(n3793) );
  XOR U5598 ( .A(n3796), .B(n3797), .Z(n3795) );
  XOR U5599 ( .A(DB[689]), .B(DB[674]), .Z(n3797) );
  AND U5600 ( .A(n334), .B(n3798), .Z(n3796) );
  XOR U5601 ( .A(n3799), .B(n3800), .Z(n3798) );
  XOR U5602 ( .A(DB[674]), .B(DB[659]), .Z(n3800) );
  AND U5603 ( .A(n338), .B(n3801), .Z(n3799) );
  XOR U5604 ( .A(n3802), .B(n3803), .Z(n3801) );
  XOR U5605 ( .A(DB[659]), .B(DB[644]), .Z(n3803) );
  AND U5606 ( .A(n342), .B(n3804), .Z(n3802) );
  XOR U5607 ( .A(n3805), .B(n3806), .Z(n3804) );
  XOR U5608 ( .A(DB[644]), .B(DB[629]), .Z(n3806) );
  AND U5609 ( .A(n346), .B(n3807), .Z(n3805) );
  XOR U5610 ( .A(n3808), .B(n3809), .Z(n3807) );
  XOR U5611 ( .A(DB[629]), .B(DB[614]), .Z(n3809) );
  AND U5612 ( .A(n350), .B(n3810), .Z(n3808) );
  XOR U5613 ( .A(n3811), .B(n3812), .Z(n3810) );
  XOR U5614 ( .A(DB[614]), .B(DB[599]), .Z(n3812) );
  AND U5615 ( .A(n354), .B(n3813), .Z(n3811) );
  XOR U5616 ( .A(n3814), .B(n3815), .Z(n3813) );
  XOR U5617 ( .A(DB[599]), .B(DB[584]), .Z(n3815) );
  AND U5618 ( .A(n358), .B(n3816), .Z(n3814) );
  XOR U5619 ( .A(n3817), .B(n3818), .Z(n3816) );
  XOR U5620 ( .A(DB[584]), .B(DB[569]), .Z(n3818) );
  AND U5621 ( .A(n362), .B(n3819), .Z(n3817) );
  XOR U5622 ( .A(n3820), .B(n3821), .Z(n3819) );
  XOR U5623 ( .A(DB[569]), .B(DB[554]), .Z(n3821) );
  AND U5624 ( .A(n366), .B(n3822), .Z(n3820) );
  XOR U5625 ( .A(n3823), .B(n3824), .Z(n3822) );
  XOR U5626 ( .A(DB[554]), .B(DB[539]), .Z(n3824) );
  AND U5627 ( .A(n370), .B(n3825), .Z(n3823) );
  XOR U5628 ( .A(n3826), .B(n3827), .Z(n3825) );
  XOR U5629 ( .A(DB[539]), .B(DB[524]), .Z(n3827) );
  AND U5630 ( .A(n374), .B(n3828), .Z(n3826) );
  XOR U5631 ( .A(n3829), .B(n3830), .Z(n3828) );
  XOR U5632 ( .A(DB[524]), .B(DB[509]), .Z(n3830) );
  AND U5633 ( .A(n378), .B(n3831), .Z(n3829) );
  XOR U5634 ( .A(n3832), .B(n3833), .Z(n3831) );
  XOR U5635 ( .A(DB[509]), .B(DB[494]), .Z(n3833) );
  AND U5636 ( .A(n382), .B(n3834), .Z(n3832) );
  XOR U5637 ( .A(n3835), .B(n3836), .Z(n3834) );
  XOR U5638 ( .A(DB[494]), .B(DB[479]), .Z(n3836) );
  AND U5639 ( .A(n386), .B(n3837), .Z(n3835) );
  XOR U5640 ( .A(n3838), .B(n3839), .Z(n3837) );
  XOR U5641 ( .A(DB[479]), .B(DB[464]), .Z(n3839) );
  AND U5642 ( .A(n390), .B(n3840), .Z(n3838) );
  XOR U5643 ( .A(n3841), .B(n3842), .Z(n3840) );
  XOR U5644 ( .A(DB[464]), .B(DB[449]), .Z(n3842) );
  AND U5645 ( .A(n394), .B(n3843), .Z(n3841) );
  XOR U5646 ( .A(n3844), .B(n3845), .Z(n3843) );
  XOR U5647 ( .A(DB[449]), .B(DB[434]), .Z(n3845) );
  AND U5648 ( .A(n398), .B(n3846), .Z(n3844) );
  XOR U5649 ( .A(n3847), .B(n3848), .Z(n3846) );
  XOR U5650 ( .A(DB[434]), .B(DB[419]), .Z(n3848) );
  AND U5651 ( .A(n402), .B(n3849), .Z(n3847) );
  XOR U5652 ( .A(n3850), .B(n3851), .Z(n3849) );
  XOR U5653 ( .A(DB[419]), .B(DB[404]), .Z(n3851) );
  AND U5654 ( .A(n406), .B(n3852), .Z(n3850) );
  XOR U5655 ( .A(n3853), .B(n3854), .Z(n3852) );
  XOR U5656 ( .A(DB[404]), .B(DB[389]), .Z(n3854) );
  AND U5657 ( .A(n410), .B(n3855), .Z(n3853) );
  XOR U5658 ( .A(n3856), .B(n3857), .Z(n3855) );
  XOR U5659 ( .A(DB[389]), .B(DB[374]), .Z(n3857) );
  AND U5660 ( .A(n414), .B(n3858), .Z(n3856) );
  XOR U5661 ( .A(n3859), .B(n3860), .Z(n3858) );
  XOR U5662 ( .A(DB[374]), .B(DB[359]), .Z(n3860) );
  AND U5663 ( .A(n418), .B(n3861), .Z(n3859) );
  XOR U5664 ( .A(n3862), .B(n3863), .Z(n3861) );
  XOR U5665 ( .A(DB[359]), .B(DB[344]), .Z(n3863) );
  AND U5666 ( .A(n422), .B(n3864), .Z(n3862) );
  XOR U5667 ( .A(n3865), .B(n3866), .Z(n3864) );
  XOR U5668 ( .A(DB[344]), .B(DB[329]), .Z(n3866) );
  AND U5669 ( .A(n426), .B(n3867), .Z(n3865) );
  XOR U5670 ( .A(n3868), .B(n3869), .Z(n3867) );
  XOR U5671 ( .A(DB[329]), .B(DB[314]), .Z(n3869) );
  AND U5672 ( .A(n430), .B(n3870), .Z(n3868) );
  XOR U5673 ( .A(n3871), .B(n3872), .Z(n3870) );
  XOR U5674 ( .A(DB[314]), .B(DB[299]), .Z(n3872) );
  AND U5675 ( .A(n434), .B(n3873), .Z(n3871) );
  XOR U5676 ( .A(n3874), .B(n3875), .Z(n3873) );
  XOR U5677 ( .A(DB[299]), .B(DB[284]), .Z(n3875) );
  AND U5678 ( .A(n438), .B(n3876), .Z(n3874) );
  XOR U5679 ( .A(n3877), .B(n3878), .Z(n3876) );
  XOR U5680 ( .A(DB[284]), .B(DB[269]), .Z(n3878) );
  AND U5681 ( .A(n442), .B(n3879), .Z(n3877) );
  XOR U5682 ( .A(n3880), .B(n3881), .Z(n3879) );
  XOR U5683 ( .A(DB[269]), .B(DB[254]), .Z(n3881) );
  AND U5684 ( .A(n446), .B(n3882), .Z(n3880) );
  XOR U5685 ( .A(n3883), .B(n3884), .Z(n3882) );
  XOR U5686 ( .A(DB[254]), .B(DB[239]), .Z(n3884) );
  AND U5687 ( .A(n450), .B(n3885), .Z(n3883) );
  XOR U5688 ( .A(n3886), .B(n3887), .Z(n3885) );
  XOR U5689 ( .A(DB[239]), .B(DB[224]), .Z(n3887) );
  AND U5690 ( .A(n454), .B(n3888), .Z(n3886) );
  XOR U5691 ( .A(n3889), .B(n3890), .Z(n3888) );
  XOR U5692 ( .A(DB[224]), .B(DB[209]), .Z(n3890) );
  AND U5693 ( .A(n458), .B(n3891), .Z(n3889) );
  XOR U5694 ( .A(n3892), .B(n3893), .Z(n3891) );
  XOR U5695 ( .A(DB[209]), .B(DB[194]), .Z(n3893) );
  AND U5696 ( .A(n462), .B(n3894), .Z(n3892) );
  XOR U5697 ( .A(n3895), .B(n3896), .Z(n3894) );
  XOR U5698 ( .A(DB[194]), .B(DB[179]), .Z(n3896) );
  AND U5699 ( .A(n466), .B(n3897), .Z(n3895) );
  XOR U5700 ( .A(n3898), .B(n3899), .Z(n3897) );
  XOR U5701 ( .A(DB[179]), .B(DB[164]), .Z(n3899) );
  AND U5702 ( .A(n470), .B(n3900), .Z(n3898) );
  XOR U5703 ( .A(n3901), .B(n3902), .Z(n3900) );
  XOR U5704 ( .A(DB[164]), .B(DB[149]), .Z(n3902) );
  AND U5705 ( .A(n474), .B(n3903), .Z(n3901) );
  XOR U5706 ( .A(n3904), .B(n3905), .Z(n3903) );
  XOR U5707 ( .A(DB[149]), .B(DB[134]), .Z(n3905) );
  AND U5708 ( .A(n478), .B(n3906), .Z(n3904) );
  XOR U5709 ( .A(n3907), .B(n3908), .Z(n3906) );
  XOR U5710 ( .A(DB[134]), .B(DB[119]), .Z(n3908) );
  AND U5711 ( .A(n482), .B(n3909), .Z(n3907) );
  XOR U5712 ( .A(n3910), .B(n3911), .Z(n3909) );
  XOR U5713 ( .A(DB[119]), .B(DB[104]), .Z(n3911) );
  AND U5714 ( .A(n486), .B(n3912), .Z(n3910) );
  XOR U5715 ( .A(n3913), .B(n3914), .Z(n3912) );
  XOR U5716 ( .A(DB[89]), .B(DB[104]), .Z(n3914) );
  AND U5717 ( .A(n490), .B(n3915), .Z(n3913) );
  XOR U5718 ( .A(n3916), .B(n3917), .Z(n3915) );
  XOR U5719 ( .A(DB[89]), .B(DB[74]), .Z(n3917) );
  AND U5720 ( .A(n494), .B(n3918), .Z(n3916) );
  XOR U5721 ( .A(n3919), .B(n3920), .Z(n3918) );
  XOR U5722 ( .A(DB[74]), .B(DB[59]), .Z(n3920) );
  AND U5723 ( .A(n498), .B(n3921), .Z(n3919) );
  XOR U5724 ( .A(n3922), .B(n3923), .Z(n3921) );
  XOR U5725 ( .A(DB[59]), .B(DB[44]), .Z(n3923) );
  AND U5726 ( .A(n502), .B(n3924), .Z(n3922) );
  XOR U5727 ( .A(n3925), .B(n3926), .Z(n3924) );
  XOR U5728 ( .A(DB[44]), .B(DB[29]), .Z(n3926) );
  AND U5729 ( .A(n506), .B(n3927), .Z(n3925) );
  XOR U5730 ( .A(DB[29]), .B(DB[14]), .Z(n3927) );
  XOR U5731 ( .A(DB[1918]), .B(n3928), .Z(min_val_out[13]) );
  AND U5732 ( .A(n2), .B(n3929), .Z(n3928) );
  XOR U5733 ( .A(n3930), .B(n3931), .Z(n3929) );
  XOR U5734 ( .A(DB[1918]), .B(DB[1903]), .Z(n3931) );
  AND U5735 ( .A(n6), .B(n3932), .Z(n3930) );
  XOR U5736 ( .A(n3933), .B(n3934), .Z(n3932) );
  XOR U5737 ( .A(DB[1903]), .B(DB[1888]), .Z(n3934) );
  AND U5738 ( .A(n10), .B(n3935), .Z(n3933) );
  XOR U5739 ( .A(n3936), .B(n3937), .Z(n3935) );
  XOR U5740 ( .A(DB[1888]), .B(DB[1873]), .Z(n3937) );
  AND U5741 ( .A(n14), .B(n3938), .Z(n3936) );
  XOR U5742 ( .A(n3939), .B(n3940), .Z(n3938) );
  XOR U5743 ( .A(DB[1873]), .B(DB[1858]), .Z(n3940) );
  AND U5744 ( .A(n18), .B(n3941), .Z(n3939) );
  XOR U5745 ( .A(n3942), .B(n3943), .Z(n3941) );
  XOR U5746 ( .A(DB[1858]), .B(DB[1843]), .Z(n3943) );
  AND U5747 ( .A(n22), .B(n3944), .Z(n3942) );
  XOR U5748 ( .A(n3945), .B(n3946), .Z(n3944) );
  XOR U5749 ( .A(DB[1843]), .B(DB[1828]), .Z(n3946) );
  AND U5750 ( .A(n26), .B(n3947), .Z(n3945) );
  XOR U5751 ( .A(n3948), .B(n3949), .Z(n3947) );
  XOR U5752 ( .A(DB[1828]), .B(DB[1813]), .Z(n3949) );
  AND U5753 ( .A(n30), .B(n3950), .Z(n3948) );
  XOR U5754 ( .A(n3951), .B(n3952), .Z(n3950) );
  XOR U5755 ( .A(DB[1813]), .B(DB[1798]), .Z(n3952) );
  AND U5756 ( .A(n34), .B(n3953), .Z(n3951) );
  XOR U5757 ( .A(n3954), .B(n3955), .Z(n3953) );
  XOR U5758 ( .A(DB[1798]), .B(DB[1783]), .Z(n3955) );
  AND U5759 ( .A(n38), .B(n3956), .Z(n3954) );
  XOR U5760 ( .A(n3957), .B(n3958), .Z(n3956) );
  XOR U5761 ( .A(DB[1783]), .B(DB[1768]), .Z(n3958) );
  AND U5762 ( .A(n42), .B(n3959), .Z(n3957) );
  XOR U5763 ( .A(n3960), .B(n3961), .Z(n3959) );
  XOR U5764 ( .A(DB[1768]), .B(DB[1753]), .Z(n3961) );
  AND U5765 ( .A(n46), .B(n3962), .Z(n3960) );
  XOR U5766 ( .A(n3963), .B(n3964), .Z(n3962) );
  XOR U5767 ( .A(DB[1753]), .B(DB[1738]), .Z(n3964) );
  AND U5768 ( .A(n50), .B(n3965), .Z(n3963) );
  XOR U5769 ( .A(n3966), .B(n3967), .Z(n3965) );
  XOR U5770 ( .A(DB[1738]), .B(DB[1723]), .Z(n3967) );
  AND U5771 ( .A(n54), .B(n3968), .Z(n3966) );
  XOR U5772 ( .A(n3969), .B(n3970), .Z(n3968) );
  XOR U5773 ( .A(DB[1723]), .B(DB[1708]), .Z(n3970) );
  AND U5774 ( .A(n58), .B(n3971), .Z(n3969) );
  XOR U5775 ( .A(n3972), .B(n3973), .Z(n3971) );
  XOR U5776 ( .A(DB[1708]), .B(DB[1693]), .Z(n3973) );
  AND U5777 ( .A(n62), .B(n3974), .Z(n3972) );
  XOR U5778 ( .A(n3975), .B(n3976), .Z(n3974) );
  XOR U5779 ( .A(DB[1693]), .B(DB[1678]), .Z(n3976) );
  AND U5780 ( .A(n66), .B(n3977), .Z(n3975) );
  XOR U5781 ( .A(n3978), .B(n3979), .Z(n3977) );
  XOR U5782 ( .A(DB[1678]), .B(DB[1663]), .Z(n3979) );
  AND U5783 ( .A(n70), .B(n3980), .Z(n3978) );
  XOR U5784 ( .A(n3981), .B(n3982), .Z(n3980) );
  XOR U5785 ( .A(DB[1663]), .B(DB[1648]), .Z(n3982) );
  AND U5786 ( .A(n74), .B(n3983), .Z(n3981) );
  XOR U5787 ( .A(n3984), .B(n3985), .Z(n3983) );
  XOR U5788 ( .A(DB[1648]), .B(DB[1633]), .Z(n3985) );
  AND U5789 ( .A(n78), .B(n3986), .Z(n3984) );
  XOR U5790 ( .A(n3987), .B(n3988), .Z(n3986) );
  XOR U5791 ( .A(DB[1633]), .B(DB[1618]), .Z(n3988) );
  AND U5792 ( .A(n82), .B(n3989), .Z(n3987) );
  XOR U5793 ( .A(n3990), .B(n3991), .Z(n3989) );
  XOR U5794 ( .A(DB[1618]), .B(DB[1603]), .Z(n3991) );
  AND U5795 ( .A(n86), .B(n3992), .Z(n3990) );
  XOR U5796 ( .A(n3993), .B(n3994), .Z(n3992) );
  XOR U5797 ( .A(DB[1603]), .B(DB[1588]), .Z(n3994) );
  AND U5798 ( .A(n90), .B(n3995), .Z(n3993) );
  XOR U5799 ( .A(n3996), .B(n3997), .Z(n3995) );
  XOR U5800 ( .A(DB[1588]), .B(DB[1573]), .Z(n3997) );
  AND U5801 ( .A(n94), .B(n3998), .Z(n3996) );
  XOR U5802 ( .A(n3999), .B(n4000), .Z(n3998) );
  XOR U5803 ( .A(DB[1573]), .B(DB[1558]), .Z(n4000) );
  AND U5804 ( .A(n98), .B(n4001), .Z(n3999) );
  XOR U5805 ( .A(n4002), .B(n4003), .Z(n4001) );
  XOR U5806 ( .A(DB[1558]), .B(DB[1543]), .Z(n4003) );
  AND U5807 ( .A(n102), .B(n4004), .Z(n4002) );
  XOR U5808 ( .A(n4005), .B(n4006), .Z(n4004) );
  XOR U5809 ( .A(DB[1543]), .B(DB[1528]), .Z(n4006) );
  AND U5810 ( .A(n106), .B(n4007), .Z(n4005) );
  XOR U5811 ( .A(n4008), .B(n4009), .Z(n4007) );
  XOR U5812 ( .A(DB[1528]), .B(DB[1513]), .Z(n4009) );
  AND U5813 ( .A(n110), .B(n4010), .Z(n4008) );
  XOR U5814 ( .A(n4011), .B(n4012), .Z(n4010) );
  XOR U5815 ( .A(DB[1513]), .B(DB[1498]), .Z(n4012) );
  AND U5816 ( .A(n114), .B(n4013), .Z(n4011) );
  XOR U5817 ( .A(n4014), .B(n4015), .Z(n4013) );
  XOR U5818 ( .A(DB[1498]), .B(DB[1483]), .Z(n4015) );
  AND U5819 ( .A(n118), .B(n4016), .Z(n4014) );
  XOR U5820 ( .A(n4017), .B(n4018), .Z(n4016) );
  XOR U5821 ( .A(DB[1483]), .B(DB[1468]), .Z(n4018) );
  AND U5822 ( .A(n122), .B(n4019), .Z(n4017) );
  XOR U5823 ( .A(n4020), .B(n4021), .Z(n4019) );
  XOR U5824 ( .A(DB[1468]), .B(DB[1453]), .Z(n4021) );
  AND U5825 ( .A(n126), .B(n4022), .Z(n4020) );
  XOR U5826 ( .A(n4023), .B(n4024), .Z(n4022) );
  XOR U5827 ( .A(DB[1453]), .B(DB[1438]), .Z(n4024) );
  AND U5828 ( .A(n130), .B(n4025), .Z(n4023) );
  XOR U5829 ( .A(n4026), .B(n4027), .Z(n4025) );
  XOR U5830 ( .A(DB[1438]), .B(DB[1423]), .Z(n4027) );
  AND U5831 ( .A(n134), .B(n4028), .Z(n4026) );
  XOR U5832 ( .A(n4029), .B(n4030), .Z(n4028) );
  XOR U5833 ( .A(DB[1423]), .B(DB[1408]), .Z(n4030) );
  AND U5834 ( .A(n138), .B(n4031), .Z(n4029) );
  XOR U5835 ( .A(n4032), .B(n4033), .Z(n4031) );
  XOR U5836 ( .A(DB[1408]), .B(DB[1393]), .Z(n4033) );
  AND U5837 ( .A(n142), .B(n4034), .Z(n4032) );
  XOR U5838 ( .A(n4035), .B(n4036), .Z(n4034) );
  XOR U5839 ( .A(DB[1393]), .B(DB[1378]), .Z(n4036) );
  AND U5840 ( .A(n146), .B(n4037), .Z(n4035) );
  XOR U5841 ( .A(n4038), .B(n4039), .Z(n4037) );
  XOR U5842 ( .A(DB[1378]), .B(DB[1363]), .Z(n4039) );
  AND U5843 ( .A(n150), .B(n4040), .Z(n4038) );
  XOR U5844 ( .A(n4041), .B(n4042), .Z(n4040) );
  XOR U5845 ( .A(DB[1363]), .B(DB[1348]), .Z(n4042) );
  AND U5846 ( .A(n154), .B(n4043), .Z(n4041) );
  XOR U5847 ( .A(n4044), .B(n4045), .Z(n4043) );
  XOR U5848 ( .A(DB[1348]), .B(DB[1333]), .Z(n4045) );
  AND U5849 ( .A(n158), .B(n4046), .Z(n4044) );
  XOR U5850 ( .A(n4047), .B(n4048), .Z(n4046) );
  XOR U5851 ( .A(DB[1333]), .B(DB[1318]), .Z(n4048) );
  AND U5852 ( .A(n162), .B(n4049), .Z(n4047) );
  XOR U5853 ( .A(n4050), .B(n4051), .Z(n4049) );
  XOR U5854 ( .A(DB[1318]), .B(DB[1303]), .Z(n4051) );
  AND U5855 ( .A(n166), .B(n4052), .Z(n4050) );
  XOR U5856 ( .A(n4053), .B(n4054), .Z(n4052) );
  XOR U5857 ( .A(DB[1303]), .B(DB[1288]), .Z(n4054) );
  AND U5858 ( .A(n170), .B(n4055), .Z(n4053) );
  XOR U5859 ( .A(n4056), .B(n4057), .Z(n4055) );
  XOR U5860 ( .A(DB[1288]), .B(DB[1273]), .Z(n4057) );
  AND U5861 ( .A(n174), .B(n4058), .Z(n4056) );
  XOR U5862 ( .A(n4059), .B(n4060), .Z(n4058) );
  XOR U5863 ( .A(DB[1273]), .B(DB[1258]), .Z(n4060) );
  AND U5864 ( .A(n178), .B(n4061), .Z(n4059) );
  XOR U5865 ( .A(n4062), .B(n4063), .Z(n4061) );
  XOR U5866 ( .A(DB[1258]), .B(DB[1243]), .Z(n4063) );
  AND U5867 ( .A(n182), .B(n4064), .Z(n4062) );
  XOR U5868 ( .A(n4065), .B(n4066), .Z(n4064) );
  XOR U5869 ( .A(DB[1243]), .B(DB[1228]), .Z(n4066) );
  AND U5870 ( .A(n186), .B(n4067), .Z(n4065) );
  XOR U5871 ( .A(n4068), .B(n4069), .Z(n4067) );
  XOR U5872 ( .A(DB[1228]), .B(DB[1213]), .Z(n4069) );
  AND U5873 ( .A(n190), .B(n4070), .Z(n4068) );
  XOR U5874 ( .A(n4071), .B(n4072), .Z(n4070) );
  XOR U5875 ( .A(DB[1213]), .B(DB[1198]), .Z(n4072) );
  AND U5876 ( .A(n194), .B(n4073), .Z(n4071) );
  XOR U5877 ( .A(n4074), .B(n4075), .Z(n4073) );
  XOR U5878 ( .A(DB[1198]), .B(DB[1183]), .Z(n4075) );
  AND U5879 ( .A(n198), .B(n4076), .Z(n4074) );
  XOR U5880 ( .A(n4077), .B(n4078), .Z(n4076) );
  XOR U5881 ( .A(DB[1183]), .B(DB[1168]), .Z(n4078) );
  AND U5882 ( .A(n202), .B(n4079), .Z(n4077) );
  XOR U5883 ( .A(n4080), .B(n4081), .Z(n4079) );
  XOR U5884 ( .A(DB[1168]), .B(DB[1153]), .Z(n4081) );
  AND U5885 ( .A(n206), .B(n4082), .Z(n4080) );
  XOR U5886 ( .A(n4083), .B(n4084), .Z(n4082) );
  XOR U5887 ( .A(DB[1153]), .B(DB[1138]), .Z(n4084) );
  AND U5888 ( .A(n210), .B(n4085), .Z(n4083) );
  XOR U5889 ( .A(n4086), .B(n4087), .Z(n4085) );
  XOR U5890 ( .A(DB[1138]), .B(DB[1123]), .Z(n4087) );
  AND U5891 ( .A(n214), .B(n4088), .Z(n4086) );
  XOR U5892 ( .A(n4089), .B(n4090), .Z(n4088) );
  XOR U5893 ( .A(DB[1123]), .B(DB[1108]), .Z(n4090) );
  AND U5894 ( .A(n218), .B(n4091), .Z(n4089) );
  XOR U5895 ( .A(n4092), .B(n4093), .Z(n4091) );
  XOR U5896 ( .A(DB[1108]), .B(DB[1093]), .Z(n4093) );
  AND U5897 ( .A(n222), .B(n4094), .Z(n4092) );
  XOR U5898 ( .A(n4095), .B(n4096), .Z(n4094) );
  XOR U5899 ( .A(DB[1093]), .B(DB[1078]), .Z(n4096) );
  AND U5900 ( .A(n226), .B(n4097), .Z(n4095) );
  XOR U5901 ( .A(n4098), .B(n4099), .Z(n4097) );
  XOR U5902 ( .A(DB[1078]), .B(DB[1063]), .Z(n4099) );
  AND U5903 ( .A(n230), .B(n4100), .Z(n4098) );
  XOR U5904 ( .A(n4101), .B(n4102), .Z(n4100) );
  XOR U5905 ( .A(DB[1063]), .B(DB[1048]), .Z(n4102) );
  AND U5906 ( .A(n234), .B(n4103), .Z(n4101) );
  XOR U5907 ( .A(n4104), .B(n4105), .Z(n4103) );
  XOR U5908 ( .A(DB[1048]), .B(DB[1033]), .Z(n4105) );
  AND U5909 ( .A(n238), .B(n4106), .Z(n4104) );
  XOR U5910 ( .A(n4107), .B(n4108), .Z(n4106) );
  XOR U5911 ( .A(DB[1033]), .B(DB[1018]), .Z(n4108) );
  AND U5912 ( .A(n242), .B(n4109), .Z(n4107) );
  XOR U5913 ( .A(n4110), .B(n4111), .Z(n4109) );
  XOR U5914 ( .A(DB[1018]), .B(DB[1003]), .Z(n4111) );
  AND U5915 ( .A(n246), .B(n4112), .Z(n4110) );
  XOR U5916 ( .A(n4113), .B(n4114), .Z(n4112) );
  XOR U5917 ( .A(DB[988]), .B(DB[1003]), .Z(n4114) );
  AND U5918 ( .A(n250), .B(n4115), .Z(n4113) );
  XOR U5919 ( .A(n4116), .B(n4117), .Z(n4115) );
  XOR U5920 ( .A(DB[988]), .B(DB[973]), .Z(n4117) );
  AND U5921 ( .A(n254), .B(n4118), .Z(n4116) );
  XOR U5922 ( .A(n4119), .B(n4120), .Z(n4118) );
  XOR U5923 ( .A(DB[973]), .B(DB[958]), .Z(n4120) );
  AND U5924 ( .A(n258), .B(n4121), .Z(n4119) );
  XOR U5925 ( .A(n4122), .B(n4123), .Z(n4121) );
  XOR U5926 ( .A(DB[958]), .B(DB[943]), .Z(n4123) );
  AND U5927 ( .A(n262), .B(n4124), .Z(n4122) );
  XOR U5928 ( .A(n4125), .B(n4126), .Z(n4124) );
  XOR U5929 ( .A(DB[943]), .B(DB[928]), .Z(n4126) );
  AND U5930 ( .A(n266), .B(n4127), .Z(n4125) );
  XOR U5931 ( .A(n4128), .B(n4129), .Z(n4127) );
  XOR U5932 ( .A(DB[928]), .B(DB[913]), .Z(n4129) );
  AND U5933 ( .A(n270), .B(n4130), .Z(n4128) );
  XOR U5934 ( .A(n4131), .B(n4132), .Z(n4130) );
  XOR U5935 ( .A(DB[913]), .B(DB[898]), .Z(n4132) );
  AND U5936 ( .A(n274), .B(n4133), .Z(n4131) );
  XOR U5937 ( .A(n4134), .B(n4135), .Z(n4133) );
  XOR U5938 ( .A(DB[898]), .B(DB[883]), .Z(n4135) );
  AND U5939 ( .A(n278), .B(n4136), .Z(n4134) );
  XOR U5940 ( .A(n4137), .B(n4138), .Z(n4136) );
  XOR U5941 ( .A(DB[883]), .B(DB[868]), .Z(n4138) );
  AND U5942 ( .A(n282), .B(n4139), .Z(n4137) );
  XOR U5943 ( .A(n4140), .B(n4141), .Z(n4139) );
  XOR U5944 ( .A(DB[868]), .B(DB[853]), .Z(n4141) );
  AND U5945 ( .A(n286), .B(n4142), .Z(n4140) );
  XOR U5946 ( .A(n4143), .B(n4144), .Z(n4142) );
  XOR U5947 ( .A(DB[853]), .B(DB[838]), .Z(n4144) );
  AND U5948 ( .A(n290), .B(n4145), .Z(n4143) );
  XOR U5949 ( .A(n4146), .B(n4147), .Z(n4145) );
  XOR U5950 ( .A(DB[838]), .B(DB[823]), .Z(n4147) );
  AND U5951 ( .A(n294), .B(n4148), .Z(n4146) );
  XOR U5952 ( .A(n4149), .B(n4150), .Z(n4148) );
  XOR U5953 ( .A(DB[823]), .B(DB[808]), .Z(n4150) );
  AND U5954 ( .A(n298), .B(n4151), .Z(n4149) );
  XOR U5955 ( .A(n4152), .B(n4153), .Z(n4151) );
  XOR U5956 ( .A(DB[808]), .B(DB[793]), .Z(n4153) );
  AND U5957 ( .A(n302), .B(n4154), .Z(n4152) );
  XOR U5958 ( .A(n4155), .B(n4156), .Z(n4154) );
  XOR U5959 ( .A(DB[793]), .B(DB[778]), .Z(n4156) );
  AND U5960 ( .A(n306), .B(n4157), .Z(n4155) );
  XOR U5961 ( .A(n4158), .B(n4159), .Z(n4157) );
  XOR U5962 ( .A(DB[778]), .B(DB[763]), .Z(n4159) );
  AND U5963 ( .A(n310), .B(n4160), .Z(n4158) );
  XOR U5964 ( .A(n4161), .B(n4162), .Z(n4160) );
  XOR U5965 ( .A(DB[763]), .B(DB[748]), .Z(n4162) );
  AND U5966 ( .A(n314), .B(n4163), .Z(n4161) );
  XOR U5967 ( .A(n4164), .B(n4165), .Z(n4163) );
  XOR U5968 ( .A(DB[748]), .B(DB[733]), .Z(n4165) );
  AND U5969 ( .A(n318), .B(n4166), .Z(n4164) );
  XOR U5970 ( .A(n4167), .B(n4168), .Z(n4166) );
  XOR U5971 ( .A(DB[733]), .B(DB[718]), .Z(n4168) );
  AND U5972 ( .A(n322), .B(n4169), .Z(n4167) );
  XOR U5973 ( .A(n4170), .B(n4171), .Z(n4169) );
  XOR U5974 ( .A(DB[718]), .B(DB[703]), .Z(n4171) );
  AND U5975 ( .A(n326), .B(n4172), .Z(n4170) );
  XOR U5976 ( .A(n4173), .B(n4174), .Z(n4172) );
  XOR U5977 ( .A(DB[703]), .B(DB[688]), .Z(n4174) );
  AND U5978 ( .A(n330), .B(n4175), .Z(n4173) );
  XOR U5979 ( .A(n4176), .B(n4177), .Z(n4175) );
  XOR U5980 ( .A(DB[688]), .B(DB[673]), .Z(n4177) );
  AND U5981 ( .A(n334), .B(n4178), .Z(n4176) );
  XOR U5982 ( .A(n4179), .B(n4180), .Z(n4178) );
  XOR U5983 ( .A(DB[673]), .B(DB[658]), .Z(n4180) );
  AND U5984 ( .A(n338), .B(n4181), .Z(n4179) );
  XOR U5985 ( .A(n4182), .B(n4183), .Z(n4181) );
  XOR U5986 ( .A(DB[658]), .B(DB[643]), .Z(n4183) );
  AND U5987 ( .A(n342), .B(n4184), .Z(n4182) );
  XOR U5988 ( .A(n4185), .B(n4186), .Z(n4184) );
  XOR U5989 ( .A(DB[643]), .B(DB[628]), .Z(n4186) );
  AND U5990 ( .A(n346), .B(n4187), .Z(n4185) );
  XOR U5991 ( .A(n4188), .B(n4189), .Z(n4187) );
  XOR U5992 ( .A(DB[628]), .B(DB[613]), .Z(n4189) );
  AND U5993 ( .A(n350), .B(n4190), .Z(n4188) );
  XOR U5994 ( .A(n4191), .B(n4192), .Z(n4190) );
  XOR U5995 ( .A(DB[613]), .B(DB[598]), .Z(n4192) );
  AND U5996 ( .A(n354), .B(n4193), .Z(n4191) );
  XOR U5997 ( .A(n4194), .B(n4195), .Z(n4193) );
  XOR U5998 ( .A(DB[598]), .B(DB[583]), .Z(n4195) );
  AND U5999 ( .A(n358), .B(n4196), .Z(n4194) );
  XOR U6000 ( .A(n4197), .B(n4198), .Z(n4196) );
  XOR U6001 ( .A(DB[583]), .B(DB[568]), .Z(n4198) );
  AND U6002 ( .A(n362), .B(n4199), .Z(n4197) );
  XOR U6003 ( .A(n4200), .B(n4201), .Z(n4199) );
  XOR U6004 ( .A(DB[568]), .B(DB[553]), .Z(n4201) );
  AND U6005 ( .A(n366), .B(n4202), .Z(n4200) );
  XOR U6006 ( .A(n4203), .B(n4204), .Z(n4202) );
  XOR U6007 ( .A(DB[553]), .B(DB[538]), .Z(n4204) );
  AND U6008 ( .A(n370), .B(n4205), .Z(n4203) );
  XOR U6009 ( .A(n4206), .B(n4207), .Z(n4205) );
  XOR U6010 ( .A(DB[538]), .B(DB[523]), .Z(n4207) );
  AND U6011 ( .A(n374), .B(n4208), .Z(n4206) );
  XOR U6012 ( .A(n4209), .B(n4210), .Z(n4208) );
  XOR U6013 ( .A(DB[523]), .B(DB[508]), .Z(n4210) );
  AND U6014 ( .A(n378), .B(n4211), .Z(n4209) );
  XOR U6015 ( .A(n4212), .B(n4213), .Z(n4211) );
  XOR U6016 ( .A(DB[508]), .B(DB[493]), .Z(n4213) );
  AND U6017 ( .A(n382), .B(n4214), .Z(n4212) );
  XOR U6018 ( .A(n4215), .B(n4216), .Z(n4214) );
  XOR U6019 ( .A(DB[493]), .B(DB[478]), .Z(n4216) );
  AND U6020 ( .A(n386), .B(n4217), .Z(n4215) );
  XOR U6021 ( .A(n4218), .B(n4219), .Z(n4217) );
  XOR U6022 ( .A(DB[478]), .B(DB[463]), .Z(n4219) );
  AND U6023 ( .A(n390), .B(n4220), .Z(n4218) );
  XOR U6024 ( .A(n4221), .B(n4222), .Z(n4220) );
  XOR U6025 ( .A(DB[463]), .B(DB[448]), .Z(n4222) );
  AND U6026 ( .A(n394), .B(n4223), .Z(n4221) );
  XOR U6027 ( .A(n4224), .B(n4225), .Z(n4223) );
  XOR U6028 ( .A(DB[448]), .B(DB[433]), .Z(n4225) );
  AND U6029 ( .A(n398), .B(n4226), .Z(n4224) );
  XOR U6030 ( .A(n4227), .B(n4228), .Z(n4226) );
  XOR U6031 ( .A(DB[433]), .B(DB[418]), .Z(n4228) );
  AND U6032 ( .A(n402), .B(n4229), .Z(n4227) );
  XOR U6033 ( .A(n4230), .B(n4231), .Z(n4229) );
  XOR U6034 ( .A(DB[418]), .B(DB[403]), .Z(n4231) );
  AND U6035 ( .A(n406), .B(n4232), .Z(n4230) );
  XOR U6036 ( .A(n4233), .B(n4234), .Z(n4232) );
  XOR U6037 ( .A(DB[403]), .B(DB[388]), .Z(n4234) );
  AND U6038 ( .A(n410), .B(n4235), .Z(n4233) );
  XOR U6039 ( .A(n4236), .B(n4237), .Z(n4235) );
  XOR U6040 ( .A(DB[388]), .B(DB[373]), .Z(n4237) );
  AND U6041 ( .A(n414), .B(n4238), .Z(n4236) );
  XOR U6042 ( .A(n4239), .B(n4240), .Z(n4238) );
  XOR U6043 ( .A(DB[373]), .B(DB[358]), .Z(n4240) );
  AND U6044 ( .A(n418), .B(n4241), .Z(n4239) );
  XOR U6045 ( .A(n4242), .B(n4243), .Z(n4241) );
  XOR U6046 ( .A(DB[358]), .B(DB[343]), .Z(n4243) );
  AND U6047 ( .A(n422), .B(n4244), .Z(n4242) );
  XOR U6048 ( .A(n4245), .B(n4246), .Z(n4244) );
  XOR U6049 ( .A(DB[343]), .B(DB[328]), .Z(n4246) );
  AND U6050 ( .A(n426), .B(n4247), .Z(n4245) );
  XOR U6051 ( .A(n4248), .B(n4249), .Z(n4247) );
  XOR U6052 ( .A(DB[328]), .B(DB[313]), .Z(n4249) );
  AND U6053 ( .A(n430), .B(n4250), .Z(n4248) );
  XOR U6054 ( .A(n4251), .B(n4252), .Z(n4250) );
  XOR U6055 ( .A(DB[313]), .B(DB[298]), .Z(n4252) );
  AND U6056 ( .A(n434), .B(n4253), .Z(n4251) );
  XOR U6057 ( .A(n4254), .B(n4255), .Z(n4253) );
  XOR U6058 ( .A(DB[298]), .B(DB[283]), .Z(n4255) );
  AND U6059 ( .A(n438), .B(n4256), .Z(n4254) );
  XOR U6060 ( .A(n4257), .B(n4258), .Z(n4256) );
  XOR U6061 ( .A(DB[283]), .B(DB[268]), .Z(n4258) );
  AND U6062 ( .A(n442), .B(n4259), .Z(n4257) );
  XOR U6063 ( .A(n4260), .B(n4261), .Z(n4259) );
  XOR U6064 ( .A(DB[268]), .B(DB[253]), .Z(n4261) );
  AND U6065 ( .A(n446), .B(n4262), .Z(n4260) );
  XOR U6066 ( .A(n4263), .B(n4264), .Z(n4262) );
  XOR U6067 ( .A(DB[253]), .B(DB[238]), .Z(n4264) );
  AND U6068 ( .A(n450), .B(n4265), .Z(n4263) );
  XOR U6069 ( .A(n4266), .B(n4267), .Z(n4265) );
  XOR U6070 ( .A(DB[238]), .B(DB[223]), .Z(n4267) );
  AND U6071 ( .A(n454), .B(n4268), .Z(n4266) );
  XOR U6072 ( .A(n4269), .B(n4270), .Z(n4268) );
  XOR U6073 ( .A(DB[223]), .B(DB[208]), .Z(n4270) );
  AND U6074 ( .A(n458), .B(n4271), .Z(n4269) );
  XOR U6075 ( .A(n4272), .B(n4273), .Z(n4271) );
  XOR U6076 ( .A(DB[208]), .B(DB[193]), .Z(n4273) );
  AND U6077 ( .A(n462), .B(n4274), .Z(n4272) );
  XOR U6078 ( .A(n4275), .B(n4276), .Z(n4274) );
  XOR U6079 ( .A(DB[193]), .B(DB[178]), .Z(n4276) );
  AND U6080 ( .A(n466), .B(n4277), .Z(n4275) );
  XOR U6081 ( .A(n4278), .B(n4279), .Z(n4277) );
  XOR U6082 ( .A(DB[178]), .B(DB[163]), .Z(n4279) );
  AND U6083 ( .A(n470), .B(n4280), .Z(n4278) );
  XOR U6084 ( .A(n4281), .B(n4282), .Z(n4280) );
  XOR U6085 ( .A(DB[163]), .B(DB[148]), .Z(n4282) );
  AND U6086 ( .A(n474), .B(n4283), .Z(n4281) );
  XOR U6087 ( .A(n4284), .B(n4285), .Z(n4283) );
  XOR U6088 ( .A(DB[148]), .B(DB[133]), .Z(n4285) );
  AND U6089 ( .A(n478), .B(n4286), .Z(n4284) );
  XOR U6090 ( .A(n4287), .B(n4288), .Z(n4286) );
  XOR U6091 ( .A(DB[133]), .B(DB[118]), .Z(n4288) );
  AND U6092 ( .A(n482), .B(n4289), .Z(n4287) );
  XOR U6093 ( .A(n4290), .B(n4291), .Z(n4289) );
  XOR U6094 ( .A(DB[118]), .B(DB[103]), .Z(n4291) );
  AND U6095 ( .A(n486), .B(n4292), .Z(n4290) );
  XOR U6096 ( .A(n4293), .B(n4294), .Z(n4292) );
  XOR U6097 ( .A(DB[88]), .B(DB[103]), .Z(n4294) );
  AND U6098 ( .A(n490), .B(n4295), .Z(n4293) );
  XOR U6099 ( .A(n4296), .B(n4297), .Z(n4295) );
  XOR U6100 ( .A(DB[88]), .B(DB[73]), .Z(n4297) );
  AND U6101 ( .A(n494), .B(n4298), .Z(n4296) );
  XOR U6102 ( .A(n4299), .B(n4300), .Z(n4298) );
  XOR U6103 ( .A(DB[73]), .B(DB[58]), .Z(n4300) );
  AND U6104 ( .A(n498), .B(n4301), .Z(n4299) );
  XOR U6105 ( .A(n4302), .B(n4303), .Z(n4301) );
  XOR U6106 ( .A(DB[58]), .B(DB[43]), .Z(n4303) );
  AND U6107 ( .A(n502), .B(n4304), .Z(n4302) );
  XOR U6108 ( .A(n4305), .B(n4306), .Z(n4304) );
  XOR U6109 ( .A(DB[43]), .B(DB[28]), .Z(n4306) );
  AND U6110 ( .A(n506), .B(n4307), .Z(n4305) );
  XOR U6111 ( .A(DB[28]), .B(DB[13]), .Z(n4307) );
  XOR U6112 ( .A(DB[1917]), .B(n4308), .Z(min_val_out[12]) );
  AND U6113 ( .A(n2), .B(n4309), .Z(n4308) );
  XOR U6114 ( .A(n4310), .B(n4311), .Z(n4309) );
  XOR U6115 ( .A(n4312), .B(n4313), .Z(n4311) );
  IV U6116 ( .A(DB[1917]), .Z(n4312) );
  AND U6117 ( .A(n6), .B(n4314), .Z(n4310) );
  XOR U6118 ( .A(n4315), .B(n4316), .Z(n4314) );
  XOR U6119 ( .A(DB[1902]), .B(DB[1887]), .Z(n4316) );
  AND U6120 ( .A(n10), .B(n4317), .Z(n4315) );
  XOR U6121 ( .A(n4318), .B(n4319), .Z(n4317) );
  XOR U6122 ( .A(DB[1887]), .B(DB[1872]), .Z(n4319) );
  AND U6123 ( .A(n14), .B(n4320), .Z(n4318) );
  XOR U6124 ( .A(n4321), .B(n4322), .Z(n4320) );
  XOR U6125 ( .A(DB[1872]), .B(DB[1857]), .Z(n4322) );
  AND U6126 ( .A(n18), .B(n4323), .Z(n4321) );
  XOR U6127 ( .A(n4324), .B(n4325), .Z(n4323) );
  XOR U6128 ( .A(DB[1857]), .B(DB[1842]), .Z(n4325) );
  AND U6129 ( .A(n22), .B(n4326), .Z(n4324) );
  XOR U6130 ( .A(n4327), .B(n4328), .Z(n4326) );
  XOR U6131 ( .A(DB[1842]), .B(DB[1827]), .Z(n4328) );
  AND U6132 ( .A(n26), .B(n4329), .Z(n4327) );
  XOR U6133 ( .A(n4330), .B(n4331), .Z(n4329) );
  XOR U6134 ( .A(DB[1827]), .B(DB[1812]), .Z(n4331) );
  AND U6135 ( .A(n30), .B(n4332), .Z(n4330) );
  XOR U6136 ( .A(n4333), .B(n4334), .Z(n4332) );
  XOR U6137 ( .A(DB[1812]), .B(DB[1797]), .Z(n4334) );
  AND U6138 ( .A(n34), .B(n4335), .Z(n4333) );
  XOR U6139 ( .A(n4336), .B(n4337), .Z(n4335) );
  XOR U6140 ( .A(DB[1797]), .B(DB[1782]), .Z(n4337) );
  AND U6141 ( .A(n38), .B(n4338), .Z(n4336) );
  XOR U6142 ( .A(n4339), .B(n4340), .Z(n4338) );
  XOR U6143 ( .A(DB[1782]), .B(DB[1767]), .Z(n4340) );
  AND U6144 ( .A(n42), .B(n4341), .Z(n4339) );
  XOR U6145 ( .A(n4342), .B(n4343), .Z(n4341) );
  XOR U6146 ( .A(DB[1767]), .B(DB[1752]), .Z(n4343) );
  AND U6147 ( .A(n46), .B(n4344), .Z(n4342) );
  XOR U6148 ( .A(n4345), .B(n4346), .Z(n4344) );
  XOR U6149 ( .A(DB[1752]), .B(DB[1737]), .Z(n4346) );
  AND U6150 ( .A(n50), .B(n4347), .Z(n4345) );
  XOR U6151 ( .A(n4348), .B(n4349), .Z(n4347) );
  XOR U6152 ( .A(DB[1737]), .B(DB[1722]), .Z(n4349) );
  AND U6153 ( .A(n54), .B(n4350), .Z(n4348) );
  XOR U6154 ( .A(n4351), .B(n4352), .Z(n4350) );
  XOR U6155 ( .A(DB[1722]), .B(DB[1707]), .Z(n4352) );
  AND U6156 ( .A(n58), .B(n4353), .Z(n4351) );
  XOR U6157 ( .A(n4354), .B(n4355), .Z(n4353) );
  XOR U6158 ( .A(DB[1707]), .B(DB[1692]), .Z(n4355) );
  AND U6159 ( .A(n62), .B(n4356), .Z(n4354) );
  XOR U6160 ( .A(n4357), .B(n4358), .Z(n4356) );
  XOR U6161 ( .A(DB[1692]), .B(DB[1677]), .Z(n4358) );
  AND U6162 ( .A(n66), .B(n4359), .Z(n4357) );
  XOR U6163 ( .A(n4360), .B(n4361), .Z(n4359) );
  XOR U6164 ( .A(DB[1677]), .B(DB[1662]), .Z(n4361) );
  AND U6165 ( .A(n70), .B(n4362), .Z(n4360) );
  XOR U6166 ( .A(n4363), .B(n4364), .Z(n4362) );
  XOR U6167 ( .A(DB[1662]), .B(DB[1647]), .Z(n4364) );
  AND U6168 ( .A(n74), .B(n4365), .Z(n4363) );
  XOR U6169 ( .A(n4366), .B(n4367), .Z(n4365) );
  XOR U6170 ( .A(DB[1647]), .B(DB[1632]), .Z(n4367) );
  AND U6171 ( .A(n78), .B(n4368), .Z(n4366) );
  XOR U6172 ( .A(n4369), .B(n4370), .Z(n4368) );
  XOR U6173 ( .A(DB[1632]), .B(DB[1617]), .Z(n4370) );
  AND U6174 ( .A(n82), .B(n4371), .Z(n4369) );
  XOR U6175 ( .A(n4372), .B(n4373), .Z(n4371) );
  XOR U6176 ( .A(DB[1617]), .B(DB[1602]), .Z(n4373) );
  AND U6177 ( .A(n86), .B(n4374), .Z(n4372) );
  XOR U6178 ( .A(n4375), .B(n4376), .Z(n4374) );
  XOR U6179 ( .A(DB[1602]), .B(DB[1587]), .Z(n4376) );
  AND U6180 ( .A(n90), .B(n4377), .Z(n4375) );
  XOR U6181 ( .A(n4378), .B(n4379), .Z(n4377) );
  XOR U6182 ( .A(DB[1587]), .B(DB[1572]), .Z(n4379) );
  AND U6183 ( .A(n94), .B(n4380), .Z(n4378) );
  XOR U6184 ( .A(n4381), .B(n4382), .Z(n4380) );
  XOR U6185 ( .A(DB[1572]), .B(DB[1557]), .Z(n4382) );
  AND U6186 ( .A(n98), .B(n4383), .Z(n4381) );
  XOR U6187 ( .A(n4384), .B(n4385), .Z(n4383) );
  XOR U6188 ( .A(DB[1557]), .B(DB[1542]), .Z(n4385) );
  AND U6189 ( .A(n102), .B(n4386), .Z(n4384) );
  XOR U6190 ( .A(n4387), .B(n4388), .Z(n4386) );
  XOR U6191 ( .A(DB[1542]), .B(DB[1527]), .Z(n4388) );
  AND U6192 ( .A(n106), .B(n4389), .Z(n4387) );
  XOR U6193 ( .A(n4390), .B(n4391), .Z(n4389) );
  XOR U6194 ( .A(DB[1527]), .B(DB[1512]), .Z(n4391) );
  AND U6195 ( .A(n110), .B(n4392), .Z(n4390) );
  XOR U6196 ( .A(n4393), .B(n4394), .Z(n4392) );
  XOR U6197 ( .A(DB[1512]), .B(DB[1497]), .Z(n4394) );
  AND U6198 ( .A(n114), .B(n4395), .Z(n4393) );
  XOR U6199 ( .A(n4396), .B(n4397), .Z(n4395) );
  XOR U6200 ( .A(DB[1497]), .B(DB[1482]), .Z(n4397) );
  AND U6201 ( .A(n118), .B(n4398), .Z(n4396) );
  XOR U6202 ( .A(n4399), .B(n4400), .Z(n4398) );
  XOR U6203 ( .A(DB[1482]), .B(DB[1467]), .Z(n4400) );
  AND U6204 ( .A(n122), .B(n4401), .Z(n4399) );
  XOR U6205 ( .A(n4402), .B(n4403), .Z(n4401) );
  XOR U6206 ( .A(DB[1467]), .B(DB[1452]), .Z(n4403) );
  AND U6207 ( .A(n126), .B(n4404), .Z(n4402) );
  XOR U6208 ( .A(n4405), .B(n4406), .Z(n4404) );
  XOR U6209 ( .A(DB[1452]), .B(DB[1437]), .Z(n4406) );
  AND U6210 ( .A(n130), .B(n4407), .Z(n4405) );
  XOR U6211 ( .A(n4408), .B(n4409), .Z(n4407) );
  XOR U6212 ( .A(DB[1437]), .B(DB[1422]), .Z(n4409) );
  AND U6213 ( .A(n134), .B(n4410), .Z(n4408) );
  XOR U6214 ( .A(n4411), .B(n4412), .Z(n4410) );
  XOR U6215 ( .A(DB[1422]), .B(DB[1407]), .Z(n4412) );
  AND U6216 ( .A(n138), .B(n4413), .Z(n4411) );
  XOR U6217 ( .A(n4414), .B(n4415), .Z(n4413) );
  XOR U6218 ( .A(DB[1407]), .B(DB[1392]), .Z(n4415) );
  AND U6219 ( .A(n142), .B(n4416), .Z(n4414) );
  XOR U6220 ( .A(n4417), .B(n4418), .Z(n4416) );
  XOR U6221 ( .A(DB[1392]), .B(DB[1377]), .Z(n4418) );
  AND U6222 ( .A(n146), .B(n4419), .Z(n4417) );
  XOR U6223 ( .A(n4420), .B(n4421), .Z(n4419) );
  XOR U6224 ( .A(DB[1377]), .B(DB[1362]), .Z(n4421) );
  AND U6225 ( .A(n150), .B(n4422), .Z(n4420) );
  XOR U6226 ( .A(n4423), .B(n4424), .Z(n4422) );
  XOR U6227 ( .A(DB[1362]), .B(DB[1347]), .Z(n4424) );
  AND U6228 ( .A(n154), .B(n4425), .Z(n4423) );
  XOR U6229 ( .A(n4426), .B(n4427), .Z(n4425) );
  XOR U6230 ( .A(DB[1347]), .B(DB[1332]), .Z(n4427) );
  AND U6231 ( .A(n158), .B(n4428), .Z(n4426) );
  XOR U6232 ( .A(n4429), .B(n4430), .Z(n4428) );
  XOR U6233 ( .A(DB[1332]), .B(DB[1317]), .Z(n4430) );
  AND U6234 ( .A(n162), .B(n4431), .Z(n4429) );
  XOR U6235 ( .A(n4432), .B(n4433), .Z(n4431) );
  XOR U6236 ( .A(DB[1317]), .B(DB[1302]), .Z(n4433) );
  AND U6237 ( .A(n166), .B(n4434), .Z(n4432) );
  XOR U6238 ( .A(n4435), .B(n4436), .Z(n4434) );
  XOR U6239 ( .A(DB[1302]), .B(DB[1287]), .Z(n4436) );
  AND U6240 ( .A(n170), .B(n4437), .Z(n4435) );
  XOR U6241 ( .A(n4438), .B(n4439), .Z(n4437) );
  XOR U6242 ( .A(DB[1287]), .B(DB[1272]), .Z(n4439) );
  AND U6243 ( .A(n174), .B(n4440), .Z(n4438) );
  XOR U6244 ( .A(n4441), .B(n4442), .Z(n4440) );
  XOR U6245 ( .A(DB[1272]), .B(DB[1257]), .Z(n4442) );
  AND U6246 ( .A(n178), .B(n4443), .Z(n4441) );
  XOR U6247 ( .A(n4444), .B(n4445), .Z(n4443) );
  XOR U6248 ( .A(DB[1257]), .B(DB[1242]), .Z(n4445) );
  AND U6249 ( .A(n182), .B(n4446), .Z(n4444) );
  XOR U6250 ( .A(n4447), .B(n4448), .Z(n4446) );
  XOR U6251 ( .A(DB[1242]), .B(DB[1227]), .Z(n4448) );
  AND U6252 ( .A(n186), .B(n4449), .Z(n4447) );
  XOR U6253 ( .A(n4450), .B(n4451), .Z(n4449) );
  XOR U6254 ( .A(DB[1227]), .B(DB[1212]), .Z(n4451) );
  AND U6255 ( .A(n190), .B(n4452), .Z(n4450) );
  XOR U6256 ( .A(n4453), .B(n4454), .Z(n4452) );
  XOR U6257 ( .A(DB[1212]), .B(DB[1197]), .Z(n4454) );
  AND U6258 ( .A(n194), .B(n4455), .Z(n4453) );
  XOR U6259 ( .A(n4456), .B(n4457), .Z(n4455) );
  XOR U6260 ( .A(DB[1197]), .B(DB[1182]), .Z(n4457) );
  AND U6261 ( .A(n198), .B(n4458), .Z(n4456) );
  XOR U6262 ( .A(n4459), .B(n4460), .Z(n4458) );
  XOR U6263 ( .A(DB[1182]), .B(DB[1167]), .Z(n4460) );
  AND U6264 ( .A(n202), .B(n4461), .Z(n4459) );
  XOR U6265 ( .A(n4462), .B(n4463), .Z(n4461) );
  XOR U6266 ( .A(DB[1167]), .B(DB[1152]), .Z(n4463) );
  AND U6267 ( .A(n206), .B(n4464), .Z(n4462) );
  XOR U6268 ( .A(n4465), .B(n4466), .Z(n4464) );
  XOR U6269 ( .A(DB[1152]), .B(DB[1137]), .Z(n4466) );
  AND U6270 ( .A(n210), .B(n4467), .Z(n4465) );
  XOR U6271 ( .A(n4468), .B(n4469), .Z(n4467) );
  XOR U6272 ( .A(DB[1137]), .B(DB[1122]), .Z(n4469) );
  AND U6273 ( .A(n214), .B(n4470), .Z(n4468) );
  XOR U6274 ( .A(n4471), .B(n4472), .Z(n4470) );
  XOR U6275 ( .A(DB[1122]), .B(DB[1107]), .Z(n4472) );
  AND U6276 ( .A(n218), .B(n4473), .Z(n4471) );
  XOR U6277 ( .A(n4474), .B(n4475), .Z(n4473) );
  XOR U6278 ( .A(DB[1107]), .B(DB[1092]), .Z(n4475) );
  AND U6279 ( .A(n222), .B(n4476), .Z(n4474) );
  XOR U6280 ( .A(n4477), .B(n4478), .Z(n4476) );
  XOR U6281 ( .A(DB[1092]), .B(DB[1077]), .Z(n4478) );
  AND U6282 ( .A(n226), .B(n4479), .Z(n4477) );
  XOR U6283 ( .A(n4480), .B(n4481), .Z(n4479) );
  XOR U6284 ( .A(DB[1077]), .B(DB[1062]), .Z(n4481) );
  AND U6285 ( .A(n230), .B(n4482), .Z(n4480) );
  XOR U6286 ( .A(n4483), .B(n4484), .Z(n4482) );
  XOR U6287 ( .A(DB[1062]), .B(DB[1047]), .Z(n4484) );
  AND U6288 ( .A(n234), .B(n4485), .Z(n4483) );
  XOR U6289 ( .A(n4486), .B(n4487), .Z(n4485) );
  XOR U6290 ( .A(DB[1047]), .B(DB[1032]), .Z(n4487) );
  AND U6291 ( .A(n238), .B(n4488), .Z(n4486) );
  XOR U6292 ( .A(n4489), .B(n4490), .Z(n4488) );
  XOR U6293 ( .A(DB[1032]), .B(DB[1017]), .Z(n4490) );
  AND U6294 ( .A(n242), .B(n4491), .Z(n4489) );
  XOR U6295 ( .A(n4492), .B(n4493), .Z(n4491) );
  XOR U6296 ( .A(DB[1017]), .B(DB[1002]), .Z(n4493) );
  AND U6297 ( .A(n246), .B(n4494), .Z(n4492) );
  XOR U6298 ( .A(n4495), .B(n4496), .Z(n4494) );
  XOR U6299 ( .A(DB[987]), .B(DB[1002]), .Z(n4496) );
  AND U6300 ( .A(n250), .B(n4497), .Z(n4495) );
  XOR U6301 ( .A(n4498), .B(n4499), .Z(n4497) );
  XOR U6302 ( .A(DB[987]), .B(DB[972]), .Z(n4499) );
  AND U6303 ( .A(n254), .B(n4500), .Z(n4498) );
  XOR U6304 ( .A(n4501), .B(n4502), .Z(n4500) );
  XOR U6305 ( .A(DB[972]), .B(DB[957]), .Z(n4502) );
  AND U6306 ( .A(n258), .B(n4503), .Z(n4501) );
  XOR U6307 ( .A(n4504), .B(n4505), .Z(n4503) );
  XOR U6308 ( .A(DB[957]), .B(DB[942]), .Z(n4505) );
  AND U6309 ( .A(n262), .B(n4506), .Z(n4504) );
  XOR U6310 ( .A(n4507), .B(n4508), .Z(n4506) );
  XOR U6311 ( .A(DB[942]), .B(DB[927]), .Z(n4508) );
  AND U6312 ( .A(n266), .B(n4509), .Z(n4507) );
  XOR U6313 ( .A(n4510), .B(n4511), .Z(n4509) );
  XOR U6314 ( .A(DB[927]), .B(DB[912]), .Z(n4511) );
  AND U6315 ( .A(n270), .B(n4512), .Z(n4510) );
  XOR U6316 ( .A(n4513), .B(n4514), .Z(n4512) );
  XOR U6317 ( .A(DB[912]), .B(DB[897]), .Z(n4514) );
  AND U6318 ( .A(n274), .B(n4515), .Z(n4513) );
  XOR U6319 ( .A(n4516), .B(n4517), .Z(n4515) );
  XOR U6320 ( .A(DB[897]), .B(DB[882]), .Z(n4517) );
  AND U6321 ( .A(n278), .B(n4518), .Z(n4516) );
  XOR U6322 ( .A(n4519), .B(n4520), .Z(n4518) );
  XOR U6323 ( .A(DB[882]), .B(DB[867]), .Z(n4520) );
  AND U6324 ( .A(n282), .B(n4521), .Z(n4519) );
  XOR U6325 ( .A(n4522), .B(n4523), .Z(n4521) );
  XOR U6326 ( .A(DB[867]), .B(DB[852]), .Z(n4523) );
  AND U6327 ( .A(n286), .B(n4524), .Z(n4522) );
  XOR U6328 ( .A(n4525), .B(n4526), .Z(n4524) );
  XOR U6329 ( .A(DB[852]), .B(DB[837]), .Z(n4526) );
  AND U6330 ( .A(n290), .B(n4527), .Z(n4525) );
  XOR U6331 ( .A(n4528), .B(n4529), .Z(n4527) );
  XOR U6332 ( .A(DB[837]), .B(DB[822]), .Z(n4529) );
  AND U6333 ( .A(n294), .B(n4530), .Z(n4528) );
  XOR U6334 ( .A(n4531), .B(n4532), .Z(n4530) );
  XOR U6335 ( .A(DB[822]), .B(DB[807]), .Z(n4532) );
  AND U6336 ( .A(n298), .B(n4533), .Z(n4531) );
  XOR U6337 ( .A(n4534), .B(n4535), .Z(n4533) );
  XOR U6338 ( .A(DB[807]), .B(DB[792]), .Z(n4535) );
  AND U6339 ( .A(n302), .B(n4536), .Z(n4534) );
  XOR U6340 ( .A(n4537), .B(n4538), .Z(n4536) );
  XOR U6341 ( .A(DB[792]), .B(DB[777]), .Z(n4538) );
  AND U6342 ( .A(n306), .B(n4539), .Z(n4537) );
  XOR U6343 ( .A(n4540), .B(n4541), .Z(n4539) );
  XOR U6344 ( .A(DB[777]), .B(DB[762]), .Z(n4541) );
  AND U6345 ( .A(n310), .B(n4542), .Z(n4540) );
  XOR U6346 ( .A(n4543), .B(n4544), .Z(n4542) );
  XOR U6347 ( .A(DB[762]), .B(DB[747]), .Z(n4544) );
  AND U6348 ( .A(n314), .B(n4545), .Z(n4543) );
  XOR U6349 ( .A(n4546), .B(n4547), .Z(n4545) );
  XOR U6350 ( .A(DB[747]), .B(DB[732]), .Z(n4547) );
  AND U6351 ( .A(n318), .B(n4548), .Z(n4546) );
  XOR U6352 ( .A(n4549), .B(n4550), .Z(n4548) );
  XOR U6353 ( .A(DB[732]), .B(DB[717]), .Z(n4550) );
  AND U6354 ( .A(n322), .B(n4551), .Z(n4549) );
  XOR U6355 ( .A(n4552), .B(n4553), .Z(n4551) );
  XOR U6356 ( .A(DB[717]), .B(DB[702]), .Z(n4553) );
  AND U6357 ( .A(n326), .B(n4554), .Z(n4552) );
  XOR U6358 ( .A(n4555), .B(n4556), .Z(n4554) );
  XOR U6359 ( .A(DB[702]), .B(DB[687]), .Z(n4556) );
  AND U6360 ( .A(n330), .B(n4557), .Z(n4555) );
  XOR U6361 ( .A(n4558), .B(n4559), .Z(n4557) );
  XOR U6362 ( .A(DB[687]), .B(DB[672]), .Z(n4559) );
  AND U6363 ( .A(n334), .B(n4560), .Z(n4558) );
  XOR U6364 ( .A(n4561), .B(n4562), .Z(n4560) );
  XOR U6365 ( .A(DB[672]), .B(DB[657]), .Z(n4562) );
  AND U6366 ( .A(n338), .B(n4563), .Z(n4561) );
  XOR U6367 ( .A(n4564), .B(n4565), .Z(n4563) );
  XOR U6368 ( .A(DB[657]), .B(DB[642]), .Z(n4565) );
  AND U6369 ( .A(n342), .B(n4566), .Z(n4564) );
  XOR U6370 ( .A(n4567), .B(n4568), .Z(n4566) );
  XOR U6371 ( .A(DB[642]), .B(DB[627]), .Z(n4568) );
  AND U6372 ( .A(n346), .B(n4569), .Z(n4567) );
  XOR U6373 ( .A(n4570), .B(n4571), .Z(n4569) );
  XOR U6374 ( .A(DB[627]), .B(DB[612]), .Z(n4571) );
  AND U6375 ( .A(n350), .B(n4572), .Z(n4570) );
  XOR U6376 ( .A(n4573), .B(n4574), .Z(n4572) );
  XOR U6377 ( .A(DB[612]), .B(DB[597]), .Z(n4574) );
  AND U6378 ( .A(n354), .B(n4575), .Z(n4573) );
  XOR U6379 ( .A(n4576), .B(n4577), .Z(n4575) );
  XOR U6380 ( .A(DB[597]), .B(DB[582]), .Z(n4577) );
  AND U6381 ( .A(n358), .B(n4578), .Z(n4576) );
  XOR U6382 ( .A(n4579), .B(n4580), .Z(n4578) );
  XOR U6383 ( .A(DB[582]), .B(DB[567]), .Z(n4580) );
  AND U6384 ( .A(n362), .B(n4581), .Z(n4579) );
  XOR U6385 ( .A(n4582), .B(n4583), .Z(n4581) );
  XOR U6386 ( .A(DB[567]), .B(DB[552]), .Z(n4583) );
  AND U6387 ( .A(n366), .B(n4584), .Z(n4582) );
  XOR U6388 ( .A(n4585), .B(n4586), .Z(n4584) );
  XOR U6389 ( .A(DB[552]), .B(DB[537]), .Z(n4586) );
  AND U6390 ( .A(n370), .B(n4587), .Z(n4585) );
  XOR U6391 ( .A(n4588), .B(n4589), .Z(n4587) );
  XOR U6392 ( .A(DB[537]), .B(DB[522]), .Z(n4589) );
  AND U6393 ( .A(n374), .B(n4590), .Z(n4588) );
  XOR U6394 ( .A(n4591), .B(n4592), .Z(n4590) );
  XOR U6395 ( .A(DB[522]), .B(DB[507]), .Z(n4592) );
  AND U6396 ( .A(n378), .B(n4593), .Z(n4591) );
  XOR U6397 ( .A(n4594), .B(n4595), .Z(n4593) );
  XOR U6398 ( .A(DB[507]), .B(DB[492]), .Z(n4595) );
  AND U6399 ( .A(n382), .B(n4596), .Z(n4594) );
  XOR U6400 ( .A(n4597), .B(n4598), .Z(n4596) );
  XOR U6401 ( .A(DB[492]), .B(DB[477]), .Z(n4598) );
  AND U6402 ( .A(n386), .B(n4599), .Z(n4597) );
  XOR U6403 ( .A(n4600), .B(n4601), .Z(n4599) );
  XOR U6404 ( .A(DB[477]), .B(DB[462]), .Z(n4601) );
  AND U6405 ( .A(n390), .B(n4602), .Z(n4600) );
  XOR U6406 ( .A(n4603), .B(n4604), .Z(n4602) );
  XOR U6407 ( .A(DB[462]), .B(DB[447]), .Z(n4604) );
  AND U6408 ( .A(n394), .B(n4605), .Z(n4603) );
  XOR U6409 ( .A(n4606), .B(n4607), .Z(n4605) );
  XOR U6410 ( .A(DB[447]), .B(DB[432]), .Z(n4607) );
  AND U6411 ( .A(n398), .B(n4608), .Z(n4606) );
  XOR U6412 ( .A(n4609), .B(n4610), .Z(n4608) );
  XOR U6413 ( .A(DB[432]), .B(DB[417]), .Z(n4610) );
  AND U6414 ( .A(n402), .B(n4611), .Z(n4609) );
  XOR U6415 ( .A(n4612), .B(n4613), .Z(n4611) );
  XOR U6416 ( .A(DB[417]), .B(DB[402]), .Z(n4613) );
  AND U6417 ( .A(n406), .B(n4614), .Z(n4612) );
  XOR U6418 ( .A(n4615), .B(n4616), .Z(n4614) );
  XOR U6419 ( .A(DB[402]), .B(DB[387]), .Z(n4616) );
  AND U6420 ( .A(n410), .B(n4617), .Z(n4615) );
  XOR U6421 ( .A(n4618), .B(n4619), .Z(n4617) );
  XOR U6422 ( .A(DB[387]), .B(DB[372]), .Z(n4619) );
  AND U6423 ( .A(n414), .B(n4620), .Z(n4618) );
  XOR U6424 ( .A(n4621), .B(n4622), .Z(n4620) );
  XOR U6425 ( .A(DB[372]), .B(DB[357]), .Z(n4622) );
  AND U6426 ( .A(n418), .B(n4623), .Z(n4621) );
  XOR U6427 ( .A(n4624), .B(n4625), .Z(n4623) );
  XOR U6428 ( .A(DB[357]), .B(DB[342]), .Z(n4625) );
  AND U6429 ( .A(n422), .B(n4626), .Z(n4624) );
  XOR U6430 ( .A(n4627), .B(n4628), .Z(n4626) );
  XOR U6431 ( .A(DB[342]), .B(DB[327]), .Z(n4628) );
  AND U6432 ( .A(n426), .B(n4629), .Z(n4627) );
  XOR U6433 ( .A(n4630), .B(n4631), .Z(n4629) );
  XOR U6434 ( .A(DB[327]), .B(DB[312]), .Z(n4631) );
  AND U6435 ( .A(n430), .B(n4632), .Z(n4630) );
  XOR U6436 ( .A(n4633), .B(n4634), .Z(n4632) );
  XOR U6437 ( .A(DB[312]), .B(DB[297]), .Z(n4634) );
  AND U6438 ( .A(n434), .B(n4635), .Z(n4633) );
  XOR U6439 ( .A(n4636), .B(n4637), .Z(n4635) );
  XOR U6440 ( .A(DB[297]), .B(DB[282]), .Z(n4637) );
  AND U6441 ( .A(n438), .B(n4638), .Z(n4636) );
  XOR U6442 ( .A(n4639), .B(n4640), .Z(n4638) );
  XOR U6443 ( .A(DB[282]), .B(DB[267]), .Z(n4640) );
  AND U6444 ( .A(n442), .B(n4641), .Z(n4639) );
  XOR U6445 ( .A(n4642), .B(n4643), .Z(n4641) );
  XOR U6446 ( .A(DB[267]), .B(DB[252]), .Z(n4643) );
  AND U6447 ( .A(n446), .B(n4644), .Z(n4642) );
  XOR U6448 ( .A(n4645), .B(n4646), .Z(n4644) );
  XOR U6449 ( .A(DB[252]), .B(DB[237]), .Z(n4646) );
  AND U6450 ( .A(n450), .B(n4647), .Z(n4645) );
  XOR U6451 ( .A(n4648), .B(n4649), .Z(n4647) );
  XOR U6452 ( .A(DB[237]), .B(DB[222]), .Z(n4649) );
  AND U6453 ( .A(n454), .B(n4650), .Z(n4648) );
  XOR U6454 ( .A(n4651), .B(n4652), .Z(n4650) );
  XOR U6455 ( .A(DB[222]), .B(DB[207]), .Z(n4652) );
  AND U6456 ( .A(n458), .B(n4653), .Z(n4651) );
  XOR U6457 ( .A(n4654), .B(n4655), .Z(n4653) );
  XOR U6458 ( .A(DB[207]), .B(DB[192]), .Z(n4655) );
  AND U6459 ( .A(n462), .B(n4656), .Z(n4654) );
  XOR U6460 ( .A(n4657), .B(n4658), .Z(n4656) );
  XOR U6461 ( .A(DB[192]), .B(DB[177]), .Z(n4658) );
  AND U6462 ( .A(n466), .B(n4659), .Z(n4657) );
  XOR U6463 ( .A(n4660), .B(n4661), .Z(n4659) );
  XOR U6464 ( .A(DB[177]), .B(DB[162]), .Z(n4661) );
  AND U6465 ( .A(n470), .B(n4662), .Z(n4660) );
  XOR U6466 ( .A(n4663), .B(n4664), .Z(n4662) );
  XOR U6467 ( .A(DB[162]), .B(DB[147]), .Z(n4664) );
  AND U6468 ( .A(n474), .B(n4665), .Z(n4663) );
  XOR U6469 ( .A(n4666), .B(n4667), .Z(n4665) );
  XOR U6470 ( .A(DB[147]), .B(DB[132]), .Z(n4667) );
  AND U6471 ( .A(n478), .B(n4668), .Z(n4666) );
  XOR U6472 ( .A(n4669), .B(n4670), .Z(n4668) );
  XOR U6473 ( .A(DB[132]), .B(DB[117]), .Z(n4670) );
  AND U6474 ( .A(n482), .B(n4671), .Z(n4669) );
  XOR U6475 ( .A(n4672), .B(n4673), .Z(n4671) );
  XOR U6476 ( .A(DB[117]), .B(DB[102]), .Z(n4673) );
  AND U6477 ( .A(n486), .B(n4674), .Z(n4672) );
  XOR U6478 ( .A(n4675), .B(n4676), .Z(n4674) );
  XOR U6479 ( .A(DB[87]), .B(DB[102]), .Z(n4676) );
  AND U6480 ( .A(n490), .B(n4677), .Z(n4675) );
  XOR U6481 ( .A(n4678), .B(n4679), .Z(n4677) );
  XOR U6482 ( .A(DB[87]), .B(DB[72]), .Z(n4679) );
  AND U6483 ( .A(n494), .B(n4680), .Z(n4678) );
  XOR U6484 ( .A(n4681), .B(n4682), .Z(n4680) );
  XOR U6485 ( .A(DB[72]), .B(DB[57]), .Z(n4682) );
  AND U6486 ( .A(n498), .B(n4683), .Z(n4681) );
  XOR U6487 ( .A(n4684), .B(n4685), .Z(n4683) );
  XOR U6488 ( .A(DB[57]), .B(DB[42]), .Z(n4685) );
  AND U6489 ( .A(n502), .B(n4686), .Z(n4684) );
  XOR U6490 ( .A(n4687), .B(n4688), .Z(n4686) );
  XOR U6491 ( .A(DB[42]), .B(DB[27]), .Z(n4688) );
  AND U6492 ( .A(n506), .B(n4689), .Z(n4687) );
  XOR U6493 ( .A(DB[27]), .B(DB[12]), .Z(n4689) );
  XOR U6494 ( .A(DB[1916]), .B(n4690), .Z(min_val_out[11]) );
  AND U6495 ( .A(n2), .B(n4691), .Z(n4690) );
  XOR U6496 ( .A(n4692), .B(n4693), .Z(n4691) );
  XOR U6497 ( .A(n4694), .B(n4695), .Z(n4693) );
  IV U6498 ( .A(DB[1916]), .Z(n4694) );
  AND U6499 ( .A(n6), .B(n4696), .Z(n4692) );
  XOR U6500 ( .A(n4697), .B(n4698), .Z(n4696) );
  XOR U6501 ( .A(DB[1901]), .B(DB[1886]), .Z(n4698) );
  AND U6502 ( .A(n10), .B(n4699), .Z(n4697) );
  XOR U6503 ( .A(n4700), .B(n4701), .Z(n4699) );
  XOR U6504 ( .A(DB[1886]), .B(DB[1871]), .Z(n4701) );
  AND U6505 ( .A(n14), .B(n4702), .Z(n4700) );
  XOR U6506 ( .A(n4703), .B(n4704), .Z(n4702) );
  XOR U6507 ( .A(DB[1871]), .B(DB[1856]), .Z(n4704) );
  AND U6508 ( .A(n18), .B(n4705), .Z(n4703) );
  XOR U6509 ( .A(n4706), .B(n4707), .Z(n4705) );
  XOR U6510 ( .A(DB[1856]), .B(DB[1841]), .Z(n4707) );
  AND U6511 ( .A(n22), .B(n4708), .Z(n4706) );
  XOR U6512 ( .A(n4709), .B(n4710), .Z(n4708) );
  XOR U6513 ( .A(DB[1841]), .B(DB[1826]), .Z(n4710) );
  AND U6514 ( .A(n26), .B(n4711), .Z(n4709) );
  XOR U6515 ( .A(n4712), .B(n4713), .Z(n4711) );
  XOR U6516 ( .A(DB[1826]), .B(DB[1811]), .Z(n4713) );
  AND U6517 ( .A(n30), .B(n4714), .Z(n4712) );
  XOR U6518 ( .A(n4715), .B(n4716), .Z(n4714) );
  XOR U6519 ( .A(DB[1811]), .B(DB[1796]), .Z(n4716) );
  AND U6520 ( .A(n34), .B(n4717), .Z(n4715) );
  XOR U6521 ( .A(n4718), .B(n4719), .Z(n4717) );
  XOR U6522 ( .A(DB[1796]), .B(DB[1781]), .Z(n4719) );
  AND U6523 ( .A(n38), .B(n4720), .Z(n4718) );
  XOR U6524 ( .A(n4721), .B(n4722), .Z(n4720) );
  XOR U6525 ( .A(DB[1781]), .B(DB[1766]), .Z(n4722) );
  AND U6526 ( .A(n42), .B(n4723), .Z(n4721) );
  XOR U6527 ( .A(n4724), .B(n4725), .Z(n4723) );
  XOR U6528 ( .A(DB[1766]), .B(DB[1751]), .Z(n4725) );
  AND U6529 ( .A(n46), .B(n4726), .Z(n4724) );
  XOR U6530 ( .A(n4727), .B(n4728), .Z(n4726) );
  XOR U6531 ( .A(DB[1751]), .B(DB[1736]), .Z(n4728) );
  AND U6532 ( .A(n50), .B(n4729), .Z(n4727) );
  XOR U6533 ( .A(n4730), .B(n4731), .Z(n4729) );
  XOR U6534 ( .A(DB[1736]), .B(DB[1721]), .Z(n4731) );
  AND U6535 ( .A(n54), .B(n4732), .Z(n4730) );
  XOR U6536 ( .A(n4733), .B(n4734), .Z(n4732) );
  XOR U6537 ( .A(DB[1721]), .B(DB[1706]), .Z(n4734) );
  AND U6538 ( .A(n58), .B(n4735), .Z(n4733) );
  XOR U6539 ( .A(n4736), .B(n4737), .Z(n4735) );
  XOR U6540 ( .A(DB[1706]), .B(DB[1691]), .Z(n4737) );
  AND U6541 ( .A(n62), .B(n4738), .Z(n4736) );
  XOR U6542 ( .A(n4739), .B(n4740), .Z(n4738) );
  XOR U6543 ( .A(DB[1691]), .B(DB[1676]), .Z(n4740) );
  AND U6544 ( .A(n66), .B(n4741), .Z(n4739) );
  XOR U6545 ( .A(n4742), .B(n4743), .Z(n4741) );
  XOR U6546 ( .A(DB[1676]), .B(DB[1661]), .Z(n4743) );
  AND U6547 ( .A(n70), .B(n4744), .Z(n4742) );
  XOR U6548 ( .A(n4745), .B(n4746), .Z(n4744) );
  XOR U6549 ( .A(DB[1661]), .B(DB[1646]), .Z(n4746) );
  AND U6550 ( .A(n74), .B(n4747), .Z(n4745) );
  XOR U6551 ( .A(n4748), .B(n4749), .Z(n4747) );
  XOR U6552 ( .A(DB[1646]), .B(DB[1631]), .Z(n4749) );
  AND U6553 ( .A(n78), .B(n4750), .Z(n4748) );
  XOR U6554 ( .A(n4751), .B(n4752), .Z(n4750) );
  XOR U6555 ( .A(DB[1631]), .B(DB[1616]), .Z(n4752) );
  AND U6556 ( .A(n82), .B(n4753), .Z(n4751) );
  XOR U6557 ( .A(n4754), .B(n4755), .Z(n4753) );
  XOR U6558 ( .A(DB[1616]), .B(DB[1601]), .Z(n4755) );
  AND U6559 ( .A(n86), .B(n4756), .Z(n4754) );
  XOR U6560 ( .A(n4757), .B(n4758), .Z(n4756) );
  XOR U6561 ( .A(DB[1601]), .B(DB[1586]), .Z(n4758) );
  AND U6562 ( .A(n90), .B(n4759), .Z(n4757) );
  XOR U6563 ( .A(n4760), .B(n4761), .Z(n4759) );
  XOR U6564 ( .A(DB[1586]), .B(DB[1571]), .Z(n4761) );
  AND U6565 ( .A(n94), .B(n4762), .Z(n4760) );
  XOR U6566 ( .A(n4763), .B(n4764), .Z(n4762) );
  XOR U6567 ( .A(DB[1571]), .B(DB[1556]), .Z(n4764) );
  AND U6568 ( .A(n98), .B(n4765), .Z(n4763) );
  XOR U6569 ( .A(n4766), .B(n4767), .Z(n4765) );
  XOR U6570 ( .A(DB[1556]), .B(DB[1541]), .Z(n4767) );
  AND U6571 ( .A(n102), .B(n4768), .Z(n4766) );
  XOR U6572 ( .A(n4769), .B(n4770), .Z(n4768) );
  XOR U6573 ( .A(DB[1541]), .B(DB[1526]), .Z(n4770) );
  AND U6574 ( .A(n106), .B(n4771), .Z(n4769) );
  XOR U6575 ( .A(n4772), .B(n4773), .Z(n4771) );
  XOR U6576 ( .A(DB[1526]), .B(DB[1511]), .Z(n4773) );
  AND U6577 ( .A(n110), .B(n4774), .Z(n4772) );
  XOR U6578 ( .A(n4775), .B(n4776), .Z(n4774) );
  XOR U6579 ( .A(DB[1511]), .B(DB[1496]), .Z(n4776) );
  AND U6580 ( .A(n114), .B(n4777), .Z(n4775) );
  XOR U6581 ( .A(n4778), .B(n4779), .Z(n4777) );
  XOR U6582 ( .A(DB[1496]), .B(DB[1481]), .Z(n4779) );
  AND U6583 ( .A(n118), .B(n4780), .Z(n4778) );
  XOR U6584 ( .A(n4781), .B(n4782), .Z(n4780) );
  XOR U6585 ( .A(DB[1481]), .B(DB[1466]), .Z(n4782) );
  AND U6586 ( .A(n122), .B(n4783), .Z(n4781) );
  XOR U6587 ( .A(n4784), .B(n4785), .Z(n4783) );
  XOR U6588 ( .A(DB[1466]), .B(DB[1451]), .Z(n4785) );
  AND U6589 ( .A(n126), .B(n4786), .Z(n4784) );
  XOR U6590 ( .A(n4787), .B(n4788), .Z(n4786) );
  XOR U6591 ( .A(DB[1451]), .B(DB[1436]), .Z(n4788) );
  AND U6592 ( .A(n130), .B(n4789), .Z(n4787) );
  XOR U6593 ( .A(n4790), .B(n4791), .Z(n4789) );
  XOR U6594 ( .A(DB[1436]), .B(DB[1421]), .Z(n4791) );
  AND U6595 ( .A(n134), .B(n4792), .Z(n4790) );
  XOR U6596 ( .A(n4793), .B(n4794), .Z(n4792) );
  XOR U6597 ( .A(DB[1421]), .B(DB[1406]), .Z(n4794) );
  AND U6598 ( .A(n138), .B(n4795), .Z(n4793) );
  XOR U6599 ( .A(n4796), .B(n4797), .Z(n4795) );
  XOR U6600 ( .A(DB[1406]), .B(DB[1391]), .Z(n4797) );
  AND U6601 ( .A(n142), .B(n4798), .Z(n4796) );
  XOR U6602 ( .A(n4799), .B(n4800), .Z(n4798) );
  XOR U6603 ( .A(DB[1391]), .B(DB[1376]), .Z(n4800) );
  AND U6604 ( .A(n146), .B(n4801), .Z(n4799) );
  XOR U6605 ( .A(n4802), .B(n4803), .Z(n4801) );
  XOR U6606 ( .A(DB[1376]), .B(DB[1361]), .Z(n4803) );
  AND U6607 ( .A(n150), .B(n4804), .Z(n4802) );
  XOR U6608 ( .A(n4805), .B(n4806), .Z(n4804) );
  XOR U6609 ( .A(DB[1361]), .B(DB[1346]), .Z(n4806) );
  AND U6610 ( .A(n154), .B(n4807), .Z(n4805) );
  XOR U6611 ( .A(n4808), .B(n4809), .Z(n4807) );
  XOR U6612 ( .A(DB[1346]), .B(DB[1331]), .Z(n4809) );
  AND U6613 ( .A(n158), .B(n4810), .Z(n4808) );
  XOR U6614 ( .A(n4811), .B(n4812), .Z(n4810) );
  XOR U6615 ( .A(DB[1331]), .B(DB[1316]), .Z(n4812) );
  AND U6616 ( .A(n162), .B(n4813), .Z(n4811) );
  XOR U6617 ( .A(n4814), .B(n4815), .Z(n4813) );
  XOR U6618 ( .A(DB[1316]), .B(DB[1301]), .Z(n4815) );
  AND U6619 ( .A(n166), .B(n4816), .Z(n4814) );
  XOR U6620 ( .A(n4817), .B(n4818), .Z(n4816) );
  XOR U6621 ( .A(DB[1301]), .B(DB[1286]), .Z(n4818) );
  AND U6622 ( .A(n170), .B(n4819), .Z(n4817) );
  XOR U6623 ( .A(n4820), .B(n4821), .Z(n4819) );
  XOR U6624 ( .A(DB[1286]), .B(DB[1271]), .Z(n4821) );
  AND U6625 ( .A(n174), .B(n4822), .Z(n4820) );
  XOR U6626 ( .A(n4823), .B(n4824), .Z(n4822) );
  XOR U6627 ( .A(DB[1271]), .B(DB[1256]), .Z(n4824) );
  AND U6628 ( .A(n178), .B(n4825), .Z(n4823) );
  XOR U6629 ( .A(n4826), .B(n4827), .Z(n4825) );
  XOR U6630 ( .A(DB[1256]), .B(DB[1241]), .Z(n4827) );
  AND U6631 ( .A(n182), .B(n4828), .Z(n4826) );
  XOR U6632 ( .A(n4829), .B(n4830), .Z(n4828) );
  XOR U6633 ( .A(DB[1241]), .B(DB[1226]), .Z(n4830) );
  AND U6634 ( .A(n186), .B(n4831), .Z(n4829) );
  XOR U6635 ( .A(n4832), .B(n4833), .Z(n4831) );
  XOR U6636 ( .A(DB[1226]), .B(DB[1211]), .Z(n4833) );
  AND U6637 ( .A(n190), .B(n4834), .Z(n4832) );
  XOR U6638 ( .A(n4835), .B(n4836), .Z(n4834) );
  XOR U6639 ( .A(DB[1211]), .B(DB[1196]), .Z(n4836) );
  AND U6640 ( .A(n194), .B(n4837), .Z(n4835) );
  XOR U6641 ( .A(n4838), .B(n4839), .Z(n4837) );
  XOR U6642 ( .A(DB[1196]), .B(DB[1181]), .Z(n4839) );
  AND U6643 ( .A(n198), .B(n4840), .Z(n4838) );
  XOR U6644 ( .A(n4841), .B(n4842), .Z(n4840) );
  XOR U6645 ( .A(DB[1181]), .B(DB[1166]), .Z(n4842) );
  AND U6646 ( .A(n202), .B(n4843), .Z(n4841) );
  XOR U6647 ( .A(n4844), .B(n4845), .Z(n4843) );
  XOR U6648 ( .A(DB[1166]), .B(DB[1151]), .Z(n4845) );
  AND U6649 ( .A(n206), .B(n4846), .Z(n4844) );
  XOR U6650 ( .A(n4847), .B(n4848), .Z(n4846) );
  XOR U6651 ( .A(DB[1151]), .B(DB[1136]), .Z(n4848) );
  AND U6652 ( .A(n210), .B(n4849), .Z(n4847) );
  XOR U6653 ( .A(n4850), .B(n4851), .Z(n4849) );
  XOR U6654 ( .A(DB[1136]), .B(DB[1121]), .Z(n4851) );
  AND U6655 ( .A(n214), .B(n4852), .Z(n4850) );
  XOR U6656 ( .A(n4853), .B(n4854), .Z(n4852) );
  XOR U6657 ( .A(DB[1121]), .B(DB[1106]), .Z(n4854) );
  AND U6658 ( .A(n218), .B(n4855), .Z(n4853) );
  XOR U6659 ( .A(n4856), .B(n4857), .Z(n4855) );
  XOR U6660 ( .A(DB[1106]), .B(DB[1091]), .Z(n4857) );
  AND U6661 ( .A(n222), .B(n4858), .Z(n4856) );
  XOR U6662 ( .A(n4859), .B(n4860), .Z(n4858) );
  XOR U6663 ( .A(DB[1091]), .B(DB[1076]), .Z(n4860) );
  AND U6664 ( .A(n226), .B(n4861), .Z(n4859) );
  XOR U6665 ( .A(n4862), .B(n4863), .Z(n4861) );
  XOR U6666 ( .A(DB[1076]), .B(DB[1061]), .Z(n4863) );
  AND U6667 ( .A(n230), .B(n4864), .Z(n4862) );
  XOR U6668 ( .A(n4865), .B(n4866), .Z(n4864) );
  XOR U6669 ( .A(DB[1061]), .B(DB[1046]), .Z(n4866) );
  AND U6670 ( .A(n234), .B(n4867), .Z(n4865) );
  XOR U6671 ( .A(n4868), .B(n4869), .Z(n4867) );
  XOR U6672 ( .A(DB[1046]), .B(DB[1031]), .Z(n4869) );
  AND U6673 ( .A(n238), .B(n4870), .Z(n4868) );
  XOR U6674 ( .A(n4871), .B(n4872), .Z(n4870) );
  XOR U6675 ( .A(DB[1031]), .B(DB[1016]), .Z(n4872) );
  AND U6676 ( .A(n242), .B(n4873), .Z(n4871) );
  XOR U6677 ( .A(n4874), .B(n4875), .Z(n4873) );
  XOR U6678 ( .A(DB[1016]), .B(DB[1001]), .Z(n4875) );
  AND U6679 ( .A(n246), .B(n4876), .Z(n4874) );
  XOR U6680 ( .A(n4877), .B(n4878), .Z(n4876) );
  XOR U6681 ( .A(DB[986]), .B(DB[1001]), .Z(n4878) );
  AND U6682 ( .A(n250), .B(n4879), .Z(n4877) );
  XOR U6683 ( .A(n4880), .B(n4881), .Z(n4879) );
  XOR U6684 ( .A(DB[986]), .B(DB[971]), .Z(n4881) );
  AND U6685 ( .A(n254), .B(n4882), .Z(n4880) );
  XOR U6686 ( .A(n4883), .B(n4884), .Z(n4882) );
  XOR U6687 ( .A(DB[971]), .B(DB[956]), .Z(n4884) );
  AND U6688 ( .A(n258), .B(n4885), .Z(n4883) );
  XOR U6689 ( .A(n4886), .B(n4887), .Z(n4885) );
  XOR U6690 ( .A(DB[956]), .B(DB[941]), .Z(n4887) );
  AND U6691 ( .A(n262), .B(n4888), .Z(n4886) );
  XOR U6692 ( .A(n4889), .B(n4890), .Z(n4888) );
  XOR U6693 ( .A(DB[941]), .B(DB[926]), .Z(n4890) );
  AND U6694 ( .A(n266), .B(n4891), .Z(n4889) );
  XOR U6695 ( .A(n4892), .B(n4893), .Z(n4891) );
  XOR U6696 ( .A(DB[926]), .B(DB[911]), .Z(n4893) );
  AND U6697 ( .A(n270), .B(n4894), .Z(n4892) );
  XOR U6698 ( .A(n4895), .B(n4896), .Z(n4894) );
  XOR U6699 ( .A(DB[911]), .B(DB[896]), .Z(n4896) );
  AND U6700 ( .A(n274), .B(n4897), .Z(n4895) );
  XOR U6701 ( .A(n4898), .B(n4899), .Z(n4897) );
  XOR U6702 ( .A(DB[896]), .B(DB[881]), .Z(n4899) );
  AND U6703 ( .A(n278), .B(n4900), .Z(n4898) );
  XOR U6704 ( .A(n4901), .B(n4902), .Z(n4900) );
  XOR U6705 ( .A(DB[881]), .B(DB[866]), .Z(n4902) );
  AND U6706 ( .A(n282), .B(n4903), .Z(n4901) );
  XOR U6707 ( .A(n4904), .B(n4905), .Z(n4903) );
  XOR U6708 ( .A(DB[866]), .B(DB[851]), .Z(n4905) );
  AND U6709 ( .A(n286), .B(n4906), .Z(n4904) );
  XOR U6710 ( .A(n4907), .B(n4908), .Z(n4906) );
  XOR U6711 ( .A(DB[851]), .B(DB[836]), .Z(n4908) );
  AND U6712 ( .A(n290), .B(n4909), .Z(n4907) );
  XOR U6713 ( .A(n4910), .B(n4911), .Z(n4909) );
  XOR U6714 ( .A(DB[836]), .B(DB[821]), .Z(n4911) );
  AND U6715 ( .A(n294), .B(n4912), .Z(n4910) );
  XOR U6716 ( .A(n4913), .B(n4914), .Z(n4912) );
  XOR U6717 ( .A(DB[821]), .B(DB[806]), .Z(n4914) );
  AND U6718 ( .A(n298), .B(n4915), .Z(n4913) );
  XOR U6719 ( .A(n4916), .B(n4917), .Z(n4915) );
  XOR U6720 ( .A(DB[806]), .B(DB[791]), .Z(n4917) );
  AND U6721 ( .A(n302), .B(n4918), .Z(n4916) );
  XOR U6722 ( .A(n4919), .B(n4920), .Z(n4918) );
  XOR U6723 ( .A(DB[791]), .B(DB[776]), .Z(n4920) );
  AND U6724 ( .A(n306), .B(n4921), .Z(n4919) );
  XOR U6725 ( .A(n4922), .B(n4923), .Z(n4921) );
  XOR U6726 ( .A(DB[776]), .B(DB[761]), .Z(n4923) );
  AND U6727 ( .A(n310), .B(n4924), .Z(n4922) );
  XOR U6728 ( .A(n4925), .B(n4926), .Z(n4924) );
  XOR U6729 ( .A(DB[761]), .B(DB[746]), .Z(n4926) );
  AND U6730 ( .A(n314), .B(n4927), .Z(n4925) );
  XOR U6731 ( .A(n4928), .B(n4929), .Z(n4927) );
  XOR U6732 ( .A(DB[746]), .B(DB[731]), .Z(n4929) );
  AND U6733 ( .A(n318), .B(n4930), .Z(n4928) );
  XOR U6734 ( .A(n4931), .B(n4932), .Z(n4930) );
  XOR U6735 ( .A(DB[731]), .B(DB[716]), .Z(n4932) );
  AND U6736 ( .A(n322), .B(n4933), .Z(n4931) );
  XOR U6737 ( .A(n4934), .B(n4935), .Z(n4933) );
  XOR U6738 ( .A(DB[716]), .B(DB[701]), .Z(n4935) );
  AND U6739 ( .A(n326), .B(n4936), .Z(n4934) );
  XOR U6740 ( .A(n4937), .B(n4938), .Z(n4936) );
  XOR U6741 ( .A(DB[701]), .B(DB[686]), .Z(n4938) );
  AND U6742 ( .A(n330), .B(n4939), .Z(n4937) );
  XOR U6743 ( .A(n4940), .B(n4941), .Z(n4939) );
  XOR U6744 ( .A(DB[686]), .B(DB[671]), .Z(n4941) );
  AND U6745 ( .A(n334), .B(n4942), .Z(n4940) );
  XOR U6746 ( .A(n4943), .B(n4944), .Z(n4942) );
  XOR U6747 ( .A(DB[671]), .B(DB[656]), .Z(n4944) );
  AND U6748 ( .A(n338), .B(n4945), .Z(n4943) );
  XOR U6749 ( .A(n4946), .B(n4947), .Z(n4945) );
  XOR U6750 ( .A(DB[656]), .B(DB[641]), .Z(n4947) );
  AND U6751 ( .A(n342), .B(n4948), .Z(n4946) );
  XOR U6752 ( .A(n4949), .B(n4950), .Z(n4948) );
  XOR U6753 ( .A(DB[641]), .B(DB[626]), .Z(n4950) );
  AND U6754 ( .A(n346), .B(n4951), .Z(n4949) );
  XOR U6755 ( .A(n4952), .B(n4953), .Z(n4951) );
  XOR U6756 ( .A(DB[626]), .B(DB[611]), .Z(n4953) );
  AND U6757 ( .A(n350), .B(n4954), .Z(n4952) );
  XOR U6758 ( .A(n4955), .B(n4956), .Z(n4954) );
  XOR U6759 ( .A(DB[611]), .B(DB[596]), .Z(n4956) );
  AND U6760 ( .A(n354), .B(n4957), .Z(n4955) );
  XOR U6761 ( .A(n4958), .B(n4959), .Z(n4957) );
  XOR U6762 ( .A(DB[596]), .B(DB[581]), .Z(n4959) );
  AND U6763 ( .A(n358), .B(n4960), .Z(n4958) );
  XOR U6764 ( .A(n4961), .B(n4962), .Z(n4960) );
  XOR U6765 ( .A(DB[581]), .B(DB[566]), .Z(n4962) );
  AND U6766 ( .A(n362), .B(n4963), .Z(n4961) );
  XOR U6767 ( .A(n4964), .B(n4965), .Z(n4963) );
  XOR U6768 ( .A(DB[566]), .B(DB[551]), .Z(n4965) );
  AND U6769 ( .A(n366), .B(n4966), .Z(n4964) );
  XOR U6770 ( .A(n4967), .B(n4968), .Z(n4966) );
  XOR U6771 ( .A(DB[551]), .B(DB[536]), .Z(n4968) );
  AND U6772 ( .A(n370), .B(n4969), .Z(n4967) );
  XOR U6773 ( .A(n4970), .B(n4971), .Z(n4969) );
  XOR U6774 ( .A(DB[536]), .B(DB[521]), .Z(n4971) );
  AND U6775 ( .A(n374), .B(n4972), .Z(n4970) );
  XOR U6776 ( .A(n4973), .B(n4974), .Z(n4972) );
  XOR U6777 ( .A(DB[521]), .B(DB[506]), .Z(n4974) );
  AND U6778 ( .A(n378), .B(n4975), .Z(n4973) );
  XOR U6779 ( .A(n4976), .B(n4977), .Z(n4975) );
  XOR U6780 ( .A(DB[506]), .B(DB[491]), .Z(n4977) );
  AND U6781 ( .A(n382), .B(n4978), .Z(n4976) );
  XOR U6782 ( .A(n4979), .B(n4980), .Z(n4978) );
  XOR U6783 ( .A(DB[491]), .B(DB[476]), .Z(n4980) );
  AND U6784 ( .A(n386), .B(n4981), .Z(n4979) );
  XOR U6785 ( .A(n4982), .B(n4983), .Z(n4981) );
  XOR U6786 ( .A(DB[476]), .B(DB[461]), .Z(n4983) );
  AND U6787 ( .A(n390), .B(n4984), .Z(n4982) );
  XOR U6788 ( .A(n4985), .B(n4986), .Z(n4984) );
  XOR U6789 ( .A(DB[461]), .B(DB[446]), .Z(n4986) );
  AND U6790 ( .A(n394), .B(n4987), .Z(n4985) );
  XOR U6791 ( .A(n4988), .B(n4989), .Z(n4987) );
  XOR U6792 ( .A(DB[446]), .B(DB[431]), .Z(n4989) );
  AND U6793 ( .A(n398), .B(n4990), .Z(n4988) );
  XOR U6794 ( .A(n4991), .B(n4992), .Z(n4990) );
  XOR U6795 ( .A(DB[431]), .B(DB[416]), .Z(n4992) );
  AND U6796 ( .A(n402), .B(n4993), .Z(n4991) );
  XOR U6797 ( .A(n4994), .B(n4995), .Z(n4993) );
  XOR U6798 ( .A(DB[416]), .B(DB[401]), .Z(n4995) );
  AND U6799 ( .A(n406), .B(n4996), .Z(n4994) );
  XOR U6800 ( .A(n4997), .B(n4998), .Z(n4996) );
  XOR U6801 ( .A(DB[401]), .B(DB[386]), .Z(n4998) );
  AND U6802 ( .A(n410), .B(n4999), .Z(n4997) );
  XOR U6803 ( .A(n5000), .B(n5001), .Z(n4999) );
  XOR U6804 ( .A(DB[386]), .B(DB[371]), .Z(n5001) );
  AND U6805 ( .A(n414), .B(n5002), .Z(n5000) );
  XOR U6806 ( .A(n5003), .B(n5004), .Z(n5002) );
  XOR U6807 ( .A(DB[371]), .B(DB[356]), .Z(n5004) );
  AND U6808 ( .A(n418), .B(n5005), .Z(n5003) );
  XOR U6809 ( .A(n5006), .B(n5007), .Z(n5005) );
  XOR U6810 ( .A(DB[356]), .B(DB[341]), .Z(n5007) );
  AND U6811 ( .A(n422), .B(n5008), .Z(n5006) );
  XOR U6812 ( .A(n5009), .B(n5010), .Z(n5008) );
  XOR U6813 ( .A(DB[341]), .B(DB[326]), .Z(n5010) );
  AND U6814 ( .A(n426), .B(n5011), .Z(n5009) );
  XOR U6815 ( .A(n5012), .B(n5013), .Z(n5011) );
  XOR U6816 ( .A(DB[326]), .B(DB[311]), .Z(n5013) );
  AND U6817 ( .A(n430), .B(n5014), .Z(n5012) );
  XOR U6818 ( .A(n5015), .B(n5016), .Z(n5014) );
  XOR U6819 ( .A(DB[311]), .B(DB[296]), .Z(n5016) );
  AND U6820 ( .A(n434), .B(n5017), .Z(n5015) );
  XOR U6821 ( .A(n5018), .B(n5019), .Z(n5017) );
  XOR U6822 ( .A(DB[296]), .B(DB[281]), .Z(n5019) );
  AND U6823 ( .A(n438), .B(n5020), .Z(n5018) );
  XOR U6824 ( .A(n5021), .B(n5022), .Z(n5020) );
  XOR U6825 ( .A(DB[281]), .B(DB[266]), .Z(n5022) );
  AND U6826 ( .A(n442), .B(n5023), .Z(n5021) );
  XOR U6827 ( .A(n5024), .B(n5025), .Z(n5023) );
  XOR U6828 ( .A(DB[266]), .B(DB[251]), .Z(n5025) );
  AND U6829 ( .A(n446), .B(n5026), .Z(n5024) );
  XOR U6830 ( .A(n5027), .B(n5028), .Z(n5026) );
  XOR U6831 ( .A(DB[251]), .B(DB[236]), .Z(n5028) );
  AND U6832 ( .A(n450), .B(n5029), .Z(n5027) );
  XOR U6833 ( .A(n5030), .B(n5031), .Z(n5029) );
  XOR U6834 ( .A(DB[236]), .B(DB[221]), .Z(n5031) );
  AND U6835 ( .A(n454), .B(n5032), .Z(n5030) );
  XOR U6836 ( .A(n5033), .B(n5034), .Z(n5032) );
  XOR U6837 ( .A(DB[221]), .B(DB[206]), .Z(n5034) );
  AND U6838 ( .A(n458), .B(n5035), .Z(n5033) );
  XOR U6839 ( .A(n5036), .B(n5037), .Z(n5035) );
  XOR U6840 ( .A(DB[206]), .B(DB[191]), .Z(n5037) );
  AND U6841 ( .A(n462), .B(n5038), .Z(n5036) );
  XOR U6842 ( .A(n5039), .B(n5040), .Z(n5038) );
  XOR U6843 ( .A(DB[191]), .B(DB[176]), .Z(n5040) );
  AND U6844 ( .A(n466), .B(n5041), .Z(n5039) );
  XOR U6845 ( .A(n5042), .B(n5043), .Z(n5041) );
  XOR U6846 ( .A(DB[176]), .B(DB[161]), .Z(n5043) );
  AND U6847 ( .A(n470), .B(n5044), .Z(n5042) );
  XOR U6848 ( .A(n5045), .B(n5046), .Z(n5044) );
  XOR U6849 ( .A(DB[161]), .B(DB[146]), .Z(n5046) );
  AND U6850 ( .A(n474), .B(n5047), .Z(n5045) );
  XOR U6851 ( .A(n5048), .B(n5049), .Z(n5047) );
  XOR U6852 ( .A(DB[146]), .B(DB[131]), .Z(n5049) );
  AND U6853 ( .A(n478), .B(n5050), .Z(n5048) );
  XOR U6854 ( .A(n5051), .B(n5052), .Z(n5050) );
  XOR U6855 ( .A(DB[131]), .B(DB[116]), .Z(n5052) );
  AND U6856 ( .A(n482), .B(n5053), .Z(n5051) );
  XOR U6857 ( .A(n5054), .B(n5055), .Z(n5053) );
  XOR U6858 ( .A(DB[116]), .B(DB[101]), .Z(n5055) );
  AND U6859 ( .A(n486), .B(n5056), .Z(n5054) );
  XOR U6860 ( .A(n5057), .B(n5058), .Z(n5056) );
  XOR U6861 ( .A(DB[86]), .B(DB[101]), .Z(n5058) );
  AND U6862 ( .A(n490), .B(n5059), .Z(n5057) );
  XOR U6863 ( .A(n5060), .B(n5061), .Z(n5059) );
  XOR U6864 ( .A(DB[86]), .B(DB[71]), .Z(n5061) );
  AND U6865 ( .A(n494), .B(n5062), .Z(n5060) );
  XOR U6866 ( .A(n5063), .B(n5064), .Z(n5062) );
  XOR U6867 ( .A(DB[71]), .B(DB[56]), .Z(n5064) );
  AND U6868 ( .A(n498), .B(n5065), .Z(n5063) );
  XOR U6869 ( .A(n5066), .B(n5067), .Z(n5065) );
  XOR U6870 ( .A(DB[56]), .B(DB[41]), .Z(n5067) );
  AND U6871 ( .A(n502), .B(n5068), .Z(n5066) );
  XOR U6872 ( .A(n5069), .B(n5070), .Z(n5068) );
  XOR U6873 ( .A(DB[41]), .B(DB[26]), .Z(n5070) );
  AND U6874 ( .A(n506), .B(n5071), .Z(n5069) );
  XOR U6875 ( .A(DB[26]), .B(DB[11]), .Z(n5071) );
  XOR U6876 ( .A(DB[1915]), .B(n5072), .Z(min_val_out[10]) );
  AND U6877 ( .A(n2), .B(n5073), .Z(n5072) );
  XOR U6878 ( .A(n5074), .B(n5075), .Z(n5073) );
  XOR U6879 ( .A(DB[1915]), .B(DB[1900]), .Z(n5075) );
  AND U6880 ( .A(n6), .B(n5076), .Z(n5074) );
  XOR U6881 ( .A(n5077), .B(n5078), .Z(n5076) );
  XOR U6882 ( .A(DB[1900]), .B(DB[1885]), .Z(n5078) );
  AND U6883 ( .A(n10), .B(n5079), .Z(n5077) );
  XOR U6884 ( .A(n5080), .B(n5081), .Z(n5079) );
  XOR U6885 ( .A(DB[1885]), .B(DB[1870]), .Z(n5081) );
  AND U6886 ( .A(n14), .B(n5082), .Z(n5080) );
  XOR U6887 ( .A(n5083), .B(n5084), .Z(n5082) );
  XOR U6888 ( .A(DB[1870]), .B(DB[1855]), .Z(n5084) );
  AND U6889 ( .A(n18), .B(n5085), .Z(n5083) );
  XOR U6890 ( .A(n5086), .B(n5087), .Z(n5085) );
  XOR U6891 ( .A(DB[1855]), .B(DB[1840]), .Z(n5087) );
  AND U6892 ( .A(n22), .B(n5088), .Z(n5086) );
  XOR U6893 ( .A(n5089), .B(n5090), .Z(n5088) );
  XOR U6894 ( .A(DB[1840]), .B(DB[1825]), .Z(n5090) );
  AND U6895 ( .A(n26), .B(n5091), .Z(n5089) );
  XOR U6896 ( .A(n5092), .B(n5093), .Z(n5091) );
  XOR U6897 ( .A(DB[1825]), .B(DB[1810]), .Z(n5093) );
  AND U6898 ( .A(n30), .B(n5094), .Z(n5092) );
  XOR U6899 ( .A(n5095), .B(n5096), .Z(n5094) );
  XOR U6900 ( .A(DB[1810]), .B(DB[1795]), .Z(n5096) );
  AND U6901 ( .A(n34), .B(n5097), .Z(n5095) );
  XOR U6902 ( .A(n5098), .B(n5099), .Z(n5097) );
  XOR U6903 ( .A(DB[1795]), .B(DB[1780]), .Z(n5099) );
  AND U6904 ( .A(n38), .B(n5100), .Z(n5098) );
  XOR U6905 ( .A(n5101), .B(n5102), .Z(n5100) );
  XOR U6906 ( .A(DB[1780]), .B(DB[1765]), .Z(n5102) );
  AND U6907 ( .A(n42), .B(n5103), .Z(n5101) );
  XOR U6908 ( .A(n5104), .B(n5105), .Z(n5103) );
  XOR U6909 ( .A(DB[1765]), .B(DB[1750]), .Z(n5105) );
  AND U6910 ( .A(n46), .B(n5106), .Z(n5104) );
  XOR U6911 ( .A(n5107), .B(n5108), .Z(n5106) );
  XOR U6912 ( .A(DB[1750]), .B(DB[1735]), .Z(n5108) );
  AND U6913 ( .A(n50), .B(n5109), .Z(n5107) );
  XOR U6914 ( .A(n5110), .B(n5111), .Z(n5109) );
  XOR U6915 ( .A(DB[1735]), .B(DB[1720]), .Z(n5111) );
  AND U6916 ( .A(n54), .B(n5112), .Z(n5110) );
  XOR U6917 ( .A(n5113), .B(n5114), .Z(n5112) );
  XOR U6918 ( .A(DB[1720]), .B(DB[1705]), .Z(n5114) );
  AND U6919 ( .A(n58), .B(n5115), .Z(n5113) );
  XOR U6920 ( .A(n5116), .B(n5117), .Z(n5115) );
  XOR U6921 ( .A(DB[1705]), .B(DB[1690]), .Z(n5117) );
  AND U6922 ( .A(n62), .B(n5118), .Z(n5116) );
  XOR U6923 ( .A(n5119), .B(n5120), .Z(n5118) );
  XOR U6924 ( .A(DB[1690]), .B(DB[1675]), .Z(n5120) );
  AND U6925 ( .A(n66), .B(n5121), .Z(n5119) );
  XOR U6926 ( .A(n5122), .B(n5123), .Z(n5121) );
  XOR U6927 ( .A(DB[1675]), .B(DB[1660]), .Z(n5123) );
  AND U6928 ( .A(n70), .B(n5124), .Z(n5122) );
  XOR U6929 ( .A(n5125), .B(n5126), .Z(n5124) );
  XOR U6930 ( .A(DB[1660]), .B(DB[1645]), .Z(n5126) );
  AND U6931 ( .A(n74), .B(n5127), .Z(n5125) );
  XOR U6932 ( .A(n5128), .B(n5129), .Z(n5127) );
  XOR U6933 ( .A(DB[1645]), .B(DB[1630]), .Z(n5129) );
  AND U6934 ( .A(n78), .B(n5130), .Z(n5128) );
  XOR U6935 ( .A(n5131), .B(n5132), .Z(n5130) );
  XOR U6936 ( .A(DB[1630]), .B(DB[1615]), .Z(n5132) );
  AND U6937 ( .A(n82), .B(n5133), .Z(n5131) );
  XOR U6938 ( .A(n5134), .B(n5135), .Z(n5133) );
  XOR U6939 ( .A(DB[1615]), .B(DB[1600]), .Z(n5135) );
  AND U6940 ( .A(n86), .B(n5136), .Z(n5134) );
  XOR U6941 ( .A(n5137), .B(n5138), .Z(n5136) );
  XOR U6942 ( .A(DB[1600]), .B(DB[1585]), .Z(n5138) );
  AND U6943 ( .A(n90), .B(n5139), .Z(n5137) );
  XOR U6944 ( .A(n5140), .B(n5141), .Z(n5139) );
  XOR U6945 ( .A(DB[1585]), .B(DB[1570]), .Z(n5141) );
  AND U6946 ( .A(n94), .B(n5142), .Z(n5140) );
  XOR U6947 ( .A(n5143), .B(n5144), .Z(n5142) );
  XOR U6948 ( .A(DB[1570]), .B(DB[1555]), .Z(n5144) );
  AND U6949 ( .A(n98), .B(n5145), .Z(n5143) );
  XOR U6950 ( .A(n5146), .B(n5147), .Z(n5145) );
  XOR U6951 ( .A(DB[1555]), .B(DB[1540]), .Z(n5147) );
  AND U6952 ( .A(n102), .B(n5148), .Z(n5146) );
  XOR U6953 ( .A(n5149), .B(n5150), .Z(n5148) );
  XOR U6954 ( .A(DB[1540]), .B(DB[1525]), .Z(n5150) );
  AND U6955 ( .A(n106), .B(n5151), .Z(n5149) );
  XOR U6956 ( .A(n5152), .B(n5153), .Z(n5151) );
  XOR U6957 ( .A(DB[1525]), .B(DB[1510]), .Z(n5153) );
  AND U6958 ( .A(n110), .B(n5154), .Z(n5152) );
  XOR U6959 ( .A(n5155), .B(n5156), .Z(n5154) );
  XOR U6960 ( .A(DB[1510]), .B(DB[1495]), .Z(n5156) );
  AND U6961 ( .A(n114), .B(n5157), .Z(n5155) );
  XOR U6962 ( .A(n5158), .B(n5159), .Z(n5157) );
  XOR U6963 ( .A(DB[1495]), .B(DB[1480]), .Z(n5159) );
  AND U6964 ( .A(n118), .B(n5160), .Z(n5158) );
  XOR U6965 ( .A(n5161), .B(n5162), .Z(n5160) );
  XOR U6966 ( .A(DB[1480]), .B(DB[1465]), .Z(n5162) );
  AND U6967 ( .A(n122), .B(n5163), .Z(n5161) );
  XOR U6968 ( .A(n5164), .B(n5165), .Z(n5163) );
  XOR U6969 ( .A(DB[1465]), .B(DB[1450]), .Z(n5165) );
  AND U6970 ( .A(n126), .B(n5166), .Z(n5164) );
  XOR U6971 ( .A(n5167), .B(n5168), .Z(n5166) );
  XOR U6972 ( .A(DB[1450]), .B(DB[1435]), .Z(n5168) );
  AND U6973 ( .A(n130), .B(n5169), .Z(n5167) );
  XOR U6974 ( .A(n5170), .B(n5171), .Z(n5169) );
  XOR U6975 ( .A(DB[1435]), .B(DB[1420]), .Z(n5171) );
  AND U6976 ( .A(n134), .B(n5172), .Z(n5170) );
  XOR U6977 ( .A(n5173), .B(n5174), .Z(n5172) );
  XOR U6978 ( .A(DB[1420]), .B(DB[1405]), .Z(n5174) );
  AND U6979 ( .A(n138), .B(n5175), .Z(n5173) );
  XOR U6980 ( .A(n5176), .B(n5177), .Z(n5175) );
  XOR U6981 ( .A(DB[1405]), .B(DB[1390]), .Z(n5177) );
  AND U6982 ( .A(n142), .B(n5178), .Z(n5176) );
  XOR U6983 ( .A(n5179), .B(n5180), .Z(n5178) );
  XOR U6984 ( .A(DB[1390]), .B(DB[1375]), .Z(n5180) );
  AND U6985 ( .A(n146), .B(n5181), .Z(n5179) );
  XOR U6986 ( .A(n5182), .B(n5183), .Z(n5181) );
  XOR U6987 ( .A(DB[1375]), .B(DB[1360]), .Z(n5183) );
  AND U6988 ( .A(n150), .B(n5184), .Z(n5182) );
  XOR U6989 ( .A(n5185), .B(n5186), .Z(n5184) );
  XOR U6990 ( .A(DB[1360]), .B(DB[1345]), .Z(n5186) );
  AND U6991 ( .A(n154), .B(n5187), .Z(n5185) );
  XOR U6992 ( .A(n5188), .B(n5189), .Z(n5187) );
  XOR U6993 ( .A(DB[1345]), .B(DB[1330]), .Z(n5189) );
  AND U6994 ( .A(n158), .B(n5190), .Z(n5188) );
  XOR U6995 ( .A(n5191), .B(n5192), .Z(n5190) );
  XOR U6996 ( .A(DB[1330]), .B(DB[1315]), .Z(n5192) );
  AND U6997 ( .A(n162), .B(n5193), .Z(n5191) );
  XOR U6998 ( .A(n5194), .B(n5195), .Z(n5193) );
  XOR U6999 ( .A(DB[1315]), .B(DB[1300]), .Z(n5195) );
  AND U7000 ( .A(n166), .B(n5196), .Z(n5194) );
  XOR U7001 ( .A(n5197), .B(n5198), .Z(n5196) );
  XOR U7002 ( .A(DB[1300]), .B(DB[1285]), .Z(n5198) );
  AND U7003 ( .A(n170), .B(n5199), .Z(n5197) );
  XOR U7004 ( .A(n5200), .B(n5201), .Z(n5199) );
  XOR U7005 ( .A(DB[1285]), .B(DB[1270]), .Z(n5201) );
  AND U7006 ( .A(n174), .B(n5202), .Z(n5200) );
  XOR U7007 ( .A(n5203), .B(n5204), .Z(n5202) );
  XOR U7008 ( .A(DB[1270]), .B(DB[1255]), .Z(n5204) );
  AND U7009 ( .A(n178), .B(n5205), .Z(n5203) );
  XOR U7010 ( .A(n5206), .B(n5207), .Z(n5205) );
  XOR U7011 ( .A(DB[1255]), .B(DB[1240]), .Z(n5207) );
  AND U7012 ( .A(n182), .B(n5208), .Z(n5206) );
  XOR U7013 ( .A(n5209), .B(n5210), .Z(n5208) );
  XOR U7014 ( .A(DB[1240]), .B(DB[1225]), .Z(n5210) );
  AND U7015 ( .A(n186), .B(n5211), .Z(n5209) );
  XOR U7016 ( .A(n5212), .B(n5213), .Z(n5211) );
  XOR U7017 ( .A(DB[1225]), .B(DB[1210]), .Z(n5213) );
  AND U7018 ( .A(n190), .B(n5214), .Z(n5212) );
  XOR U7019 ( .A(n5215), .B(n5216), .Z(n5214) );
  XOR U7020 ( .A(DB[1210]), .B(DB[1195]), .Z(n5216) );
  AND U7021 ( .A(n194), .B(n5217), .Z(n5215) );
  XOR U7022 ( .A(n5218), .B(n5219), .Z(n5217) );
  XOR U7023 ( .A(DB[1195]), .B(DB[1180]), .Z(n5219) );
  AND U7024 ( .A(n198), .B(n5220), .Z(n5218) );
  XOR U7025 ( .A(n5221), .B(n5222), .Z(n5220) );
  XOR U7026 ( .A(DB[1180]), .B(DB[1165]), .Z(n5222) );
  AND U7027 ( .A(n202), .B(n5223), .Z(n5221) );
  XOR U7028 ( .A(n5224), .B(n5225), .Z(n5223) );
  XOR U7029 ( .A(DB[1165]), .B(DB[1150]), .Z(n5225) );
  AND U7030 ( .A(n206), .B(n5226), .Z(n5224) );
  XOR U7031 ( .A(n5227), .B(n5228), .Z(n5226) );
  XOR U7032 ( .A(DB[1150]), .B(DB[1135]), .Z(n5228) );
  AND U7033 ( .A(n210), .B(n5229), .Z(n5227) );
  XOR U7034 ( .A(n5230), .B(n5231), .Z(n5229) );
  XOR U7035 ( .A(DB[1135]), .B(DB[1120]), .Z(n5231) );
  AND U7036 ( .A(n214), .B(n5232), .Z(n5230) );
  XOR U7037 ( .A(n5233), .B(n5234), .Z(n5232) );
  XOR U7038 ( .A(DB[1120]), .B(DB[1105]), .Z(n5234) );
  AND U7039 ( .A(n218), .B(n5235), .Z(n5233) );
  XOR U7040 ( .A(n5236), .B(n5237), .Z(n5235) );
  XOR U7041 ( .A(DB[1105]), .B(DB[1090]), .Z(n5237) );
  AND U7042 ( .A(n222), .B(n5238), .Z(n5236) );
  XOR U7043 ( .A(n5239), .B(n5240), .Z(n5238) );
  XOR U7044 ( .A(DB[1090]), .B(DB[1075]), .Z(n5240) );
  AND U7045 ( .A(n226), .B(n5241), .Z(n5239) );
  XOR U7046 ( .A(n5242), .B(n5243), .Z(n5241) );
  XOR U7047 ( .A(DB[1075]), .B(DB[1060]), .Z(n5243) );
  AND U7048 ( .A(n230), .B(n5244), .Z(n5242) );
  XOR U7049 ( .A(n5245), .B(n5246), .Z(n5244) );
  XOR U7050 ( .A(DB[1060]), .B(DB[1045]), .Z(n5246) );
  AND U7051 ( .A(n234), .B(n5247), .Z(n5245) );
  XOR U7052 ( .A(n5248), .B(n5249), .Z(n5247) );
  XOR U7053 ( .A(DB[1045]), .B(DB[1030]), .Z(n5249) );
  AND U7054 ( .A(n238), .B(n5250), .Z(n5248) );
  XOR U7055 ( .A(n5251), .B(n5252), .Z(n5250) );
  XOR U7056 ( .A(DB[1030]), .B(DB[1015]), .Z(n5252) );
  AND U7057 ( .A(n242), .B(n5253), .Z(n5251) );
  XOR U7058 ( .A(n5254), .B(n5255), .Z(n5253) );
  XOR U7059 ( .A(DB[1015]), .B(DB[1000]), .Z(n5255) );
  AND U7060 ( .A(n246), .B(n5256), .Z(n5254) );
  XOR U7061 ( .A(n5257), .B(n5258), .Z(n5256) );
  XOR U7062 ( .A(DB[985]), .B(DB[1000]), .Z(n5258) );
  AND U7063 ( .A(n250), .B(n5259), .Z(n5257) );
  XOR U7064 ( .A(n5260), .B(n5261), .Z(n5259) );
  XOR U7065 ( .A(DB[985]), .B(DB[970]), .Z(n5261) );
  AND U7066 ( .A(n254), .B(n5262), .Z(n5260) );
  XOR U7067 ( .A(n5263), .B(n5264), .Z(n5262) );
  XOR U7068 ( .A(DB[970]), .B(DB[955]), .Z(n5264) );
  AND U7069 ( .A(n258), .B(n5265), .Z(n5263) );
  XOR U7070 ( .A(n5266), .B(n5267), .Z(n5265) );
  XOR U7071 ( .A(DB[955]), .B(DB[940]), .Z(n5267) );
  AND U7072 ( .A(n262), .B(n5268), .Z(n5266) );
  XOR U7073 ( .A(n5269), .B(n5270), .Z(n5268) );
  XOR U7074 ( .A(DB[940]), .B(DB[925]), .Z(n5270) );
  AND U7075 ( .A(n266), .B(n5271), .Z(n5269) );
  XOR U7076 ( .A(n5272), .B(n5273), .Z(n5271) );
  XOR U7077 ( .A(DB[925]), .B(DB[910]), .Z(n5273) );
  AND U7078 ( .A(n270), .B(n5274), .Z(n5272) );
  XOR U7079 ( .A(n5275), .B(n5276), .Z(n5274) );
  XOR U7080 ( .A(DB[910]), .B(DB[895]), .Z(n5276) );
  AND U7081 ( .A(n274), .B(n5277), .Z(n5275) );
  XOR U7082 ( .A(n5278), .B(n5279), .Z(n5277) );
  XOR U7083 ( .A(DB[895]), .B(DB[880]), .Z(n5279) );
  AND U7084 ( .A(n278), .B(n5280), .Z(n5278) );
  XOR U7085 ( .A(n5281), .B(n5282), .Z(n5280) );
  XOR U7086 ( .A(DB[880]), .B(DB[865]), .Z(n5282) );
  AND U7087 ( .A(n282), .B(n5283), .Z(n5281) );
  XOR U7088 ( .A(n5284), .B(n5285), .Z(n5283) );
  XOR U7089 ( .A(DB[865]), .B(DB[850]), .Z(n5285) );
  AND U7090 ( .A(n286), .B(n5286), .Z(n5284) );
  XOR U7091 ( .A(n5287), .B(n5288), .Z(n5286) );
  XOR U7092 ( .A(DB[850]), .B(DB[835]), .Z(n5288) );
  AND U7093 ( .A(n290), .B(n5289), .Z(n5287) );
  XOR U7094 ( .A(n5290), .B(n5291), .Z(n5289) );
  XOR U7095 ( .A(DB[835]), .B(DB[820]), .Z(n5291) );
  AND U7096 ( .A(n294), .B(n5292), .Z(n5290) );
  XOR U7097 ( .A(n5293), .B(n5294), .Z(n5292) );
  XOR U7098 ( .A(DB[820]), .B(DB[805]), .Z(n5294) );
  AND U7099 ( .A(n298), .B(n5295), .Z(n5293) );
  XOR U7100 ( .A(n5296), .B(n5297), .Z(n5295) );
  XOR U7101 ( .A(DB[805]), .B(DB[790]), .Z(n5297) );
  AND U7102 ( .A(n302), .B(n5298), .Z(n5296) );
  XOR U7103 ( .A(n5299), .B(n5300), .Z(n5298) );
  XOR U7104 ( .A(DB[790]), .B(DB[775]), .Z(n5300) );
  AND U7105 ( .A(n306), .B(n5301), .Z(n5299) );
  XOR U7106 ( .A(n5302), .B(n5303), .Z(n5301) );
  XOR U7107 ( .A(DB[775]), .B(DB[760]), .Z(n5303) );
  AND U7108 ( .A(n310), .B(n5304), .Z(n5302) );
  XOR U7109 ( .A(n5305), .B(n5306), .Z(n5304) );
  XOR U7110 ( .A(DB[760]), .B(DB[745]), .Z(n5306) );
  AND U7111 ( .A(n314), .B(n5307), .Z(n5305) );
  XOR U7112 ( .A(n5308), .B(n5309), .Z(n5307) );
  XOR U7113 ( .A(DB[745]), .B(DB[730]), .Z(n5309) );
  AND U7114 ( .A(n318), .B(n5310), .Z(n5308) );
  XOR U7115 ( .A(n5311), .B(n5312), .Z(n5310) );
  XOR U7116 ( .A(DB[730]), .B(DB[715]), .Z(n5312) );
  AND U7117 ( .A(n322), .B(n5313), .Z(n5311) );
  XOR U7118 ( .A(n5314), .B(n5315), .Z(n5313) );
  XOR U7119 ( .A(DB[715]), .B(DB[700]), .Z(n5315) );
  AND U7120 ( .A(n326), .B(n5316), .Z(n5314) );
  XOR U7121 ( .A(n5317), .B(n5318), .Z(n5316) );
  XOR U7122 ( .A(DB[700]), .B(DB[685]), .Z(n5318) );
  AND U7123 ( .A(n330), .B(n5319), .Z(n5317) );
  XOR U7124 ( .A(n5320), .B(n5321), .Z(n5319) );
  XOR U7125 ( .A(DB[685]), .B(DB[670]), .Z(n5321) );
  AND U7126 ( .A(n334), .B(n5322), .Z(n5320) );
  XOR U7127 ( .A(n5323), .B(n5324), .Z(n5322) );
  XOR U7128 ( .A(DB[670]), .B(DB[655]), .Z(n5324) );
  AND U7129 ( .A(n338), .B(n5325), .Z(n5323) );
  XOR U7130 ( .A(n5326), .B(n5327), .Z(n5325) );
  XOR U7131 ( .A(DB[655]), .B(DB[640]), .Z(n5327) );
  AND U7132 ( .A(n342), .B(n5328), .Z(n5326) );
  XOR U7133 ( .A(n5329), .B(n5330), .Z(n5328) );
  XOR U7134 ( .A(DB[640]), .B(DB[625]), .Z(n5330) );
  AND U7135 ( .A(n346), .B(n5331), .Z(n5329) );
  XOR U7136 ( .A(n5332), .B(n5333), .Z(n5331) );
  XOR U7137 ( .A(DB[625]), .B(DB[610]), .Z(n5333) );
  AND U7138 ( .A(n350), .B(n5334), .Z(n5332) );
  XOR U7139 ( .A(n5335), .B(n5336), .Z(n5334) );
  XOR U7140 ( .A(DB[610]), .B(DB[595]), .Z(n5336) );
  AND U7141 ( .A(n354), .B(n5337), .Z(n5335) );
  XOR U7142 ( .A(n5338), .B(n5339), .Z(n5337) );
  XOR U7143 ( .A(DB[595]), .B(DB[580]), .Z(n5339) );
  AND U7144 ( .A(n358), .B(n5340), .Z(n5338) );
  XOR U7145 ( .A(n5341), .B(n5342), .Z(n5340) );
  XOR U7146 ( .A(DB[580]), .B(DB[565]), .Z(n5342) );
  AND U7147 ( .A(n362), .B(n5343), .Z(n5341) );
  XOR U7148 ( .A(n5344), .B(n5345), .Z(n5343) );
  XOR U7149 ( .A(DB[565]), .B(DB[550]), .Z(n5345) );
  AND U7150 ( .A(n366), .B(n5346), .Z(n5344) );
  XOR U7151 ( .A(n5347), .B(n5348), .Z(n5346) );
  XOR U7152 ( .A(DB[550]), .B(DB[535]), .Z(n5348) );
  AND U7153 ( .A(n370), .B(n5349), .Z(n5347) );
  XOR U7154 ( .A(n5350), .B(n5351), .Z(n5349) );
  XOR U7155 ( .A(DB[535]), .B(DB[520]), .Z(n5351) );
  AND U7156 ( .A(n374), .B(n5352), .Z(n5350) );
  XOR U7157 ( .A(n5353), .B(n5354), .Z(n5352) );
  XOR U7158 ( .A(DB[520]), .B(DB[505]), .Z(n5354) );
  AND U7159 ( .A(n378), .B(n5355), .Z(n5353) );
  XOR U7160 ( .A(n5356), .B(n5357), .Z(n5355) );
  XOR U7161 ( .A(DB[505]), .B(DB[490]), .Z(n5357) );
  AND U7162 ( .A(n382), .B(n5358), .Z(n5356) );
  XOR U7163 ( .A(n5359), .B(n5360), .Z(n5358) );
  XOR U7164 ( .A(DB[490]), .B(DB[475]), .Z(n5360) );
  AND U7165 ( .A(n386), .B(n5361), .Z(n5359) );
  XOR U7166 ( .A(n5362), .B(n5363), .Z(n5361) );
  XOR U7167 ( .A(DB[475]), .B(DB[460]), .Z(n5363) );
  AND U7168 ( .A(n390), .B(n5364), .Z(n5362) );
  XOR U7169 ( .A(n5365), .B(n5366), .Z(n5364) );
  XOR U7170 ( .A(DB[460]), .B(DB[445]), .Z(n5366) );
  AND U7171 ( .A(n394), .B(n5367), .Z(n5365) );
  XOR U7172 ( .A(n5368), .B(n5369), .Z(n5367) );
  XOR U7173 ( .A(DB[445]), .B(DB[430]), .Z(n5369) );
  AND U7174 ( .A(n398), .B(n5370), .Z(n5368) );
  XOR U7175 ( .A(n5371), .B(n5372), .Z(n5370) );
  XOR U7176 ( .A(DB[430]), .B(DB[415]), .Z(n5372) );
  AND U7177 ( .A(n402), .B(n5373), .Z(n5371) );
  XOR U7178 ( .A(n5374), .B(n5375), .Z(n5373) );
  XOR U7179 ( .A(DB[415]), .B(DB[400]), .Z(n5375) );
  AND U7180 ( .A(n406), .B(n5376), .Z(n5374) );
  XOR U7181 ( .A(n5377), .B(n5378), .Z(n5376) );
  XOR U7182 ( .A(DB[400]), .B(DB[385]), .Z(n5378) );
  AND U7183 ( .A(n410), .B(n5379), .Z(n5377) );
  XOR U7184 ( .A(n5380), .B(n5381), .Z(n5379) );
  XOR U7185 ( .A(DB[385]), .B(DB[370]), .Z(n5381) );
  AND U7186 ( .A(n414), .B(n5382), .Z(n5380) );
  XOR U7187 ( .A(n5383), .B(n5384), .Z(n5382) );
  XOR U7188 ( .A(DB[370]), .B(DB[355]), .Z(n5384) );
  AND U7189 ( .A(n418), .B(n5385), .Z(n5383) );
  XOR U7190 ( .A(n5386), .B(n5387), .Z(n5385) );
  XOR U7191 ( .A(DB[355]), .B(DB[340]), .Z(n5387) );
  AND U7192 ( .A(n422), .B(n5388), .Z(n5386) );
  XOR U7193 ( .A(n5389), .B(n5390), .Z(n5388) );
  XOR U7194 ( .A(DB[340]), .B(DB[325]), .Z(n5390) );
  AND U7195 ( .A(n426), .B(n5391), .Z(n5389) );
  XOR U7196 ( .A(n5392), .B(n5393), .Z(n5391) );
  XOR U7197 ( .A(DB[325]), .B(DB[310]), .Z(n5393) );
  AND U7198 ( .A(n430), .B(n5394), .Z(n5392) );
  XOR U7199 ( .A(n5395), .B(n5396), .Z(n5394) );
  XOR U7200 ( .A(DB[310]), .B(DB[295]), .Z(n5396) );
  AND U7201 ( .A(n434), .B(n5397), .Z(n5395) );
  XOR U7202 ( .A(n5398), .B(n5399), .Z(n5397) );
  XOR U7203 ( .A(DB[295]), .B(DB[280]), .Z(n5399) );
  AND U7204 ( .A(n438), .B(n5400), .Z(n5398) );
  XOR U7205 ( .A(n5401), .B(n5402), .Z(n5400) );
  XOR U7206 ( .A(DB[280]), .B(DB[265]), .Z(n5402) );
  AND U7207 ( .A(n442), .B(n5403), .Z(n5401) );
  XOR U7208 ( .A(n5404), .B(n5405), .Z(n5403) );
  XOR U7209 ( .A(DB[265]), .B(DB[250]), .Z(n5405) );
  AND U7210 ( .A(n446), .B(n5406), .Z(n5404) );
  XOR U7211 ( .A(n5407), .B(n5408), .Z(n5406) );
  XOR U7212 ( .A(DB[250]), .B(DB[235]), .Z(n5408) );
  AND U7213 ( .A(n450), .B(n5409), .Z(n5407) );
  XOR U7214 ( .A(n5410), .B(n5411), .Z(n5409) );
  XOR U7215 ( .A(DB[235]), .B(DB[220]), .Z(n5411) );
  AND U7216 ( .A(n454), .B(n5412), .Z(n5410) );
  XOR U7217 ( .A(n5413), .B(n5414), .Z(n5412) );
  XOR U7218 ( .A(DB[220]), .B(DB[205]), .Z(n5414) );
  AND U7219 ( .A(n458), .B(n5415), .Z(n5413) );
  XOR U7220 ( .A(n5416), .B(n5417), .Z(n5415) );
  XOR U7221 ( .A(DB[205]), .B(DB[190]), .Z(n5417) );
  AND U7222 ( .A(n462), .B(n5418), .Z(n5416) );
  XOR U7223 ( .A(n5419), .B(n5420), .Z(n5418) );
  XOR U7224 ( .A(DB[190]), .B(DB[175]), .Z(n5420) );
  AND U7225 ( .A(n466), .B(n5421), .Z(n5419) );
  XOR U7226 ( .A(n5422), .B(n5423), .Z(n5421) );
  XOR U7227 ( .A(DB[175]), .B(DB[160]), .Z(n5423) );
  AND U7228 ( .A(n470), .B(n5424), .Z(n5422) );
  XOR U7229 ( .A(n5425), .B(n5426), .Z(n5424) );
  XOR U7230 ( .A(DB[160]), .B(DB[145]), .Z(n5426) );
  AND U7231 ( .A(n474), .B(n5427), .Z(n5425) );
  XOR U7232 ( .A(n5428), .B(n5429), .Z(n5427) );
  XOR U7233 ( .A(DB[145]), .B(DB[130]), .Z(n5429) );
  AND U7234 ( .A(n478), .B(n5430), .Z(n5428) );
  XOR U7235 ( .A(n5431), .B(n5432), .Z(n5430) );
  XOR U7236 ( .A(DB[130]), .B(DB[115]), .Z(n5432) );
  AND U7237 ( .A(n482), .B(n5433), .Z(n5431) );
  XOR U7238 ( .A(n5434), .B(n5435), .Z(n5433) );
  XOR U7239 ( .A(DB[115]), .B(DB[100]), .Z(n5435) );
  AND U7240 ( .A(n486), .B(n5436), .Z(n5434) );
  XOR U7241 ( .A(n5437), .B(n5438), .Z(n5436) );
  XOR U7242 ( .A(DB[85]), .B(DB[100]), .Z(n5438) );
  AND U7243 ( .A(n490), .B(n5439), .Z(n5437) );
  XOR U7244 ( .A(n5440), .B(n5441), .Z(n5439) );
  XOR U7245 ( .A(DB[85]), .B(DB[70]), .Z(n5441) );
  AND U7246 ( .A(n494), .B(n5442), .Z(n5440) );
  XOR U7247 ( .A(n5443), .B(n5444), .Z(n5442) );
  XOR U7248 ( .A(DB[70]), .B(DB[55]), .Z(n5444) );
  AND U7249 ( .A(n498), .B(n5445), .Z(n5443) );
  XOR U7250 ( .A(n5446), .B(n5447), .Z(n5445) );
  XOR U7251 ( .A(DB[55]), .B(DB[40]), .Z(n5447) );
  AND U7252 ( .A(n502), .B(n5448), .Z(n5446) );
  XOR U7253 ( .A(n5449), .B(n5450), .Z(n5448) );
  XOR U7254 ( .A(DB[40]), .B(DB[25]), .Z(n5450) );
  AND U7255 ( .A(n506), .B(n5451), .Z(n5449) );
  XOR U7256 ( .A(DB[25]), .B(DB[10]), .Z(n5451) );
  XOR U7257 ( .A(DB[1905]), .B(n5452), .Z(min_val_out[0]) );
  AND U7258 ( .A(n2), .B(n5453), .Z(n5452) );
  XOR U7259 ( .A(n5454), .B(n5455), .Z(n5453) );
  XOR U7260 ( .A(DB[1905]), .B(DB[1890]), .Z(n5455) );
  AND U7261 ( .A(n6), .B(n5456), .Z(n5454) );
  XOR U7262 ( .A(n5457), .B(n5458), .Z(n5456) );
  XOR U7263 ( .A(DB[1890]), .B(DB[1875]), .Z(n5458) );
  AND U7264 ( .A(n10), .B(n5459), .Z(n5457) );
  XOR U7265 ( .A(n5460), .B(n5461), .Z(n5459) );
  XOR U7266 ( .A(DB[1875]), .B(DB[1860]), .Z(n5461) );
  AND U7267 ( .A(n14), .B(n5462), .Z(n5460) );
  XOR U7268 ( .A(n5463), .B(n5464), .Z(n5462) );
  XOR U7269 ( .A(DB[1860]), .B(DB[1845]), .Z(n5464) );
  AND U7270 ( .A(n18), .B(n5465), .Z(n5463) );
  XOR U7271 ( .A(n5466), .B(n5467), .Z(n5465) );
  XOR U7272 ( .A(DB[1845]), .B(DB[1830]), .Z(n5467) );
  AND U7273 ( .A(n22), .B(n5468), .Z(n5466) );
  XOR U7274 ( .A(n5469), .B(n5470), .Z(n5468) );
  XOR U7275 ( .A(DB[1830]), .B(DB[1815]), .Z(n5470) );
  AND U7276 ( .A(n26), .B(n5471), .Z(n5469) );
  XOR U7277 ( .A(n5472), .B(n5473), .Z(n5471) );
  XOR U7278 ( .A(DB[1815]), .B(DB[1800]), .Z(n5473) );
  AND U7279 ( .A(n30), .B(n5474), .Z(n5472) );
  XOR U7280 ( .A(n5475), .B(n5476), .Z(n5474) );
  XOR U7281 ( .A(DB[1800]), .B(DB[1785]), .Z(n5476) );
  AND U7282 ( .A(n34), .B(n5477), .Z(n5475) );
  XOR U7283 ( .A(n5478), .B(n5479), .Z(n5477) );
  XOR U7284 ( .A(DB[1785]), .B(DB[1770]), .Z(n5479) );
  AND U7285 ( .A(n38), .B(n5480), .Z(n5478) );
  XOR U7286 ( .A(n5481), .B(n5482), .Z(n5480) );
  XOR U7287 ( .A(DB[1770]), .B(DB[1755]), .Z(n5482) );
  AND U7288 ( .A(n42), .B(n5483), .Z(n5481) );
  XOR U7289 ( .A(n5484), .B(n5485), .Z(n5483) );
  XOR U7290 ( .A(DB[1755]), .B(DB[1740]), .Z(n5485) );
  AND U7291 ( .A(n46), .B(n5486), .Z(n5484) );
  XOR U7292 ( .A(n5487), .B(n5488), .Z(n5486) );
  XOR U7293 ( .A(DB[1740]), .B(DB[1725]), .Z(n5488) );
  AND U7294 ( .A(n50), .B(n5489), .Z(n5487) );
  XOR U7295 ( .A(n5490), .B(n5491), .Z(n5489) );
  XOR U7296 ( .A(DB[1725]), .B(DB[1710]), .Z(n5491) );
  AND U7297 ( .A(n54), .B(n5492), .Z(n5490) );
  XOR U7298 ( .A(n5493), .B(n5494), .Z(n5492) );
  XOR U7299 ( .A(DB[1710]), .B(DB[1695]), .Z(n5494) );
  AND U7300 ( .A(n58), .B(n5495), .Z(n5493) );
  XOR U7301 ( .A(n5496), .B(n5497), .Z(n5495) );
  XOR U7302 ( .A(DB[1695]), .B(DB[1680]), .Z(n5497) );
  AND U7303 ( .A(n62), .B(n5498), .Z(n5496) );
  XOR U7304 ( .A(n5499), .B(n5500), .Z(n5498) );
  XOR U7305 ( .A(DB[1680]), .B(DB[1665]), .Z(n5500) );
  AND U7306 ( .A(n66), .B(n5501), .Z(n5499) );
  XOR U7307 ( .A(n5502), .B(n5503), .Z(n5501) );
  XOR U7308 ( .A(DB[1665]), .B(DB[1650]), .Z(n5503) );
  AND U7309 ( .A(n70), .B(n5504), .Z(n5502) );
  XOR U7310 ( .A(n5505), .B(n5506), .Z(n5504) );
  XOR U7311 ( .A(DB[1650]), .B(DB[1635]), .Z(n5506) );
  AND U7312 ( .A(n74), .B(n5507), .Z(n5505) );
  XOR U7313 ( .A(n5508), .B(n5509), .Z(n5507) );
  XOR U7314 ( .A(DB[1635]), .B(DB[1620]), .Z(n5509) );
  AND U7315 ( .A(n78), .B(n5510), .Z(n5508) );
  XOR U7316 ( .A(n5511), .B(n5512), .Z(n5510) );
  XOR U7317 ( .A(DB[1620]), .B(DB[1605]), .Z(n5512) );
  AND U7318 ( .A(n82), .B(n5513), .Z(n5511) );
  XOR U7319 ( .A(n5514), .B(n5515), .Z(n5513) );
  XOR U7320 ( .A(DB[1605]), .B(DB[1590]), .Z(n5515) );
  AND U7321 ( .A(n86), .B(n5516), .Z(n5514) );
  XOR U7322 ( .A(n5517), .B(n5518), .Z(n5516) );
  XOR U7323 ( .A(DB[1590]), .B(DB[1575]), .Z(n5518) );
  AND U7324 ( .A(n90), .B(n5519), .Z(n5517) );
  XOR U7325 ( .A(n5520), .B(n5521), .Z(n5519) );
  XOR U7326 ( .A(DB[1575]), .B(DB[1560]), .Z(n5521) );
  AND U7327 ( .A(n94), .B(n5522), .Z(n5520) );
  XOR U7328 ( .A(n5523), .B(n5524), .Z(n5522) );
  XOR U7329 ( .A(DB[1560]), .B(DB[1545]), .Z(n5524) );
  AND U7330 ( .A(n98), .B(n5525), .Z(n5523) );
  XOR U7331 ( .A(n5526), .B(n5527), .Z(n5525) );
  XOR U7332 ( .A(DB[1545]), .B(DB[1530]), .Z(n5527) );
  AND U7333 ( .A(n102), .B(n5528), .Z(n5526) );
  XOR U7334 ( .A(n5529), .B(n5530), .Z(n5528) );
  XOR U7335 ( .A(DB[1530]), .B(DB[1515]), .Z(n5530) );
  AND U7336 ( .A(n106), .B(n5531), .Z(n5529) );
  XOR U7337 ( .A(n5532), .B(n5533), .Z(n5531) );
  XOR U7338 ( .A(DB[1515]), .B(DB[1500]), .Z(n5533) );
  AND U7339 ( .A(n110), .B(n5534), .Z(n5532) );
  XOR U7340 ( .A(n5535), .B(n5536), .Z(n5534) );
  XOR U7341 ( .A(DB[1500]), .B(DB[1485]), .Z(n5536) );
  AND U7342 ( .A(n114), .B(n5537), .Z(n5535) );
  XOR U7343 ( .A(n5538), .B(n5539), .Z(n5537) );
  XOR U7344 ( .A(DB[1485]), .B(DB[1470]), .Z(n5539) );
  AND U7345 ( .A(n118), .B(n5540), .Z(n5538) );
  XOR U7346 ( .A(n5541), .B(n5542), .Z(n5540) );
  XOR U7347 ( .A(DB[1470]), .B(DB[1455]), .Z(n5542) );
  AND U7348 ( .A(n122), .B(n5543), .Z(n5541) );
  XOR U7349 ( .A(n5544), .B(n5545), .Z(n5543) );
  XOR U7350 ( .A(DB[1455]), .B(DB[1440]), .Z(n5545) );
  AND U7351 ( .A(n126), .B(n5546), .Z(n5544) );
  XOR U7352 ( .A(n5547), .B(n5548), .Z(n5546) );
  XOR U7353 ( .A(DB[1440]), .B(DB[1425]), .Z(n5548) );
  AND U7354 ( .A(n130), .B(n5549), .Z(n5547) );
  XOR U7355 ( .A(n5550), .B(n5551), .Z(n5549) );
  XOR U7356 ( .A(DB[1425]), .B(DB[1410]), .Z(n5551) );
  AND U7357 ( .A(n134), .B(n5552), .Z(n5550) );
  XOR U7358 ( .A(n5553), .B(n5554), .Z(n5552) );
  XOR U7359 ( .A(DB[1410]), .B(DB[1395]), .Z(n5554) );
  AND U7360 ( .A(n138), .B(n5555), .Z(n5553) );
  XOR U7361 ( .A(n5556), .B(n5557), .Z(n5555) );
  XOR U7362 ( .A(DB[1395]), .B(DB[1380]), .Z(n5557) );
  AND U7363 ( .A(n142), .B(n5558), .Z(n5556) );
  XOR U7364 ( .A(n5559), .B(n5560), .Z(n5558) );
  XOR U7365 ( .A(DB[1380]), .B(DB[1365]), .Z(n5560) );
  AND U7366 ( .A(n146), .B(n5561), .Z(n5559) );
  XOR U7367 ( .A(n5562), .B(n5563), .Z(n5561) );
  XOR U7368 ( .A(DB[1365]), .B(DB[1350]), .Z(n5563) );
  AND U7369 ( .A(n150), .B(n5564), .Z(n5562) );
  XOR U7370 ( .A(n5565), .B(n5566), .Z(n5564) );
  XOR U7371 ( .A(DB[1350]), .B(DB[1335]), .Z(n5566) );
  AND U7372 ( .A(n154), .B(n5567), .Z(n5565) );
  XOR U7373 ( .A(n5568), .B(n5569), .Z(n5567) );
  XOR U7374 ( .A(DB[1335]), .B(DB[1320]), .Z(n5569) );
  AND U7375 ( .A(n158), .B(n5570), .Z(n5568) );
  XOR U7376 ( .A(n5571), .B(n5572), .Z(n5570) );
  XOR U7377 ( .A(DB[1320]), .B(DB[1305]), .Z(n5572) );
  AND U7378 ( .A(n162), .B(n5573), .Z(n5571) );
  XOR U7379 ( .A(n5574), .B(n5575), .Z(n5573) );
  XOR U7380 ( .A(DB[1305]), .B(DB[1290]), .Z(n5575) );
  AND U7381 ( .A(n166), .B(n5576), .Z(n5574) );
  XOR U7382 ( .A(n5577), .B(n5578), .Z(n5576) );
  XOR U7383 ( .A(DB[1290]), .B(DB[1275]), .Z(n5578) );
  AND U7384 ( .A(n170), .B(n5579), .Z(n5577) );
  XOR U7385 ( .A(n5580), .B(n5581), .Z(n5579) );
  XOR U7386 ( .A(DB[1275]), .B(DB[1260]), .Z(n5581) );
  AND U7387 ( .A(n174), .B(n5582), .Z(n5580) );
  XOR U7388 ( .A(n5583), .B(n5584), .Z(n5582) );
  XOR U7389 ( .A(DB[1260]), .B(DB[1245]), .Z(n5584) );
  AND U7390 ( .A(n178), .B(n5585), .Z(n5583) );
  XOR U7391 ( .A(n5586), .B(n5587), .Z(n5585) );
  XOR U7392 ( .A(DB[1245]), .B(DB[1230]), .Z(n5587) );
  AND U7393 ( .A(n182), .B(n5588), .Z(n5586) );
  XOR U7394 ( .A(n5589), .B(n5590), .Z(n5588) );
  XOR U7395 ( .A(DB[1230]), .B(DB[1215]), .Z(n5590) );
  AND U7396 ( .A(n186), .B(n5591), .Z(n5589) );
  XOR U7397 ( .A(n5592), .B(n5593), .Z(n5591) );
  XOR U7398 ( .A(DB[1215]), .B(DB[1200]), .Z(n5593) );
  AND U7399 ( .A(n190), .B(n5594), .Z(n5592) );
  XOR U7400 ( .A(n5595), .B(n5596), .Z(n5594) );
  XOR U7401 ( .A(DB[1200]), .B(DB[1185]), .Z(n5596) );
  AND U7402 ( .A(n194), .B(n5597), .Z(n5595) );
  XOR U7403 ( .A(n5598), .B(n5599), .Z(n5597) );
  XOR U7404 ( .A(DB[1185]), .B(DB[1170]), .Z(n5599) );
  AND U7405 ( .A(n198), .B(n5600), .Z(n5598) );
  XOR U7406 ( .A(n5601), .B(n5602), .Z(n5600) );
  XOR U7407 ( .A(DB[1170]), .B(DB[1155]), .Z(n5602) );
  AND U7408 ( .A(n202), .B(n5603), .Z(n5601) );
  XOR U7409 ( .A(n5604), .B(n5605), .Z(n5603) );
  XOR U7410 ( .A(DB[1155]), .B(DB[1140]), .Z(n5605) );
  AND U7411 ( .A(n206), .B(n5606), .Z(n5604) );
  XOR U7412 ( .A(n5607), .B(n5608), .Z(n5606) );
  XOR U7413 ( .A(DB[1140]), .B(DB[1125]), .Z(n5608) );
  AND U7414 ( .A(n210), .B(n5609), .Z(n5607) );
  XOR U7415 ( .A(n5610), .B(n5611), .Z(n5609) );
  XOR U7416 ( .A(DB[1125]), .B(DB[1110]), .Z(n5611) );
  AND U7417 ( .A(n214), .B(n5612), .Z(n5610) );
  XOR U7418 ( .A(n5613), .B(n5614), .Z(n5612) );
  XOR U7419 ( .A(DB[1110]), .B(DB[1095]), .Z(n5614) );
  AND U7420 ( .A(n218), .B(n5615), .Z(n5613) );
  XOR U7421 ( .A(n5616), .B(n5617), .Z(n5615) );
  XOR U7422 ( .A(DB[1095]), .B(DB[1080]), .Z(n5617) );
  AND U7423 ( .A(n222), .B(n5618), .Z(n5616) );
  XOR U7424 ( .A(n5619), .B(n5620), .Z(n5618) );
  XOR U7425 ( .A(DB[1080]), .B(DB[1065]), .Z(n5620) );
  AND U7426 ( .A(n226), .B(n5621), .Z(n5619) );
  XOR U7427 ( .A(n5622), .B(n5623), .Z(n5621) );
  XOR U7428 ( .A(DB[1065]), .B(DB[1050]), .Z(n5623) );
  AND U7429 ( .A(n230), .B(n5624), .Z(n5622) );
  XOR U7430 ( .A(n5625), .B(n5626), .Z(n5624) );
  XOR U7431 ( .A(DB[1050]), .B(DB[1035]), .Z(n5626) );
  AND U7432 ( .A(n234), .B(n5627), .Z(n5625) );
  XOR U7433 ( .A(n5628), .B(n5629), .Z(n5627) );
  XOR U7434 ( .A(DB[1035]), .B(DB[1020]), .Z(n5629) );
  AND U7435 ( .A(n238), .B(n5630), .Z(n5628) );
  XOR U7436 ( .A(n5631), .B(n5632), .Z(n5630) );
  XOR U7437 ( .A(DB[1020]), .B(DB[1005]), .Z(n5632) );
  AND U7438 ( .A(n242), .B(n5633), .Z(n5631) );
  XOR U7439 ( .A(n5634), .B(n5635), .Z(n5633) );
  XOR U7440 ( .A(DB[990]), .B(DB[1005]), .Z(n5635) );
  AND U7441 ( .A(n246), .B(n5636), .Z(n5634) );
  XOR U7442 ( .A(n5637), .B(n5638), .Z(n5636) );
  XOR U7443 ( .A(DB[990]), .B(DB[975]), .Z(n5638) );
  AND U7444 ( .A(n250), .B(n5639), .Z(n5637) );
  XOR U7445 ( .A(n5640), .B(n5641), .Z(n5639) );
  XOR U7446 ( .A(DB[975]), .B(DB[960]), .Z(n5641) );
  AND U7447 ( .A(n254), .B(n5642), .Z(n5640) );
  XOR U7448 ( .A(n5643), .B(n5644), .Z(n5642) );
  XOR U7449 ( .A(DB[960]), .B(DB[945]), .Z(n5644) );
  AND U7450 ( .A(n258), .B(n5645), .Z(n5643) );
  XOR U7451 ( .A(n5646), .B(n5647), .Z(n5645) );
  XOR U7452 ( .A(DB[945]), .B(DB[930]), .Z(n5647) );
  AND U7453 ( .A(n262), .B(n5648), .Z(n5646) );
  XOR U7454 ( .A(n5649), .B(n5650), .Z(n5648) );
  XOR U7455 ( .A(DB[930]), .B(DB[915]), .Z(n5650) );
  AND U7456 ( .A(n266), .B(n5651), .Z(n5649) );
  XOR U7457 ( .A(n5652), .B(n5653), .Z(n5651) );
  XOR U7458 ( .A(DB[915]), .B(DB[900]), .Z(n5653) );
  AND U7459 ( .A(n270), .B(n5654), .Z(n5652) );
  XOR U7460 ( .A(n5655), .B(n5656), .Z(n5654) );
  XOR U7461 ( .A(DB[900]), .B(DB[885]), .Z(n5656) );
  AND U7462 ( .A(n274), .B(n5657), .Z(n5655) );
  XOR U7463 ( .A(n5658), .B(n5659), .Z(n5657) );
  XOR U7464 ( .A(DB[885]), .B(DB[870]), .Z(n5659) );
  AND U7465 ( .A(n278), .B(n5660), .Z(n5658) );
  XOR U7466 ( .A(n5661), .B(n5662), .Z(n5660) );
  XOR U7467 ( .A(DB[870]), .B(DB[855]), .Z(n5662) );
  AND U7468 ( .A(n282), .B(n5663), .Z(n5661) );
  XOR U7469 ( .A(n5664), .B(n5665), .Z(n5663) );
  XOR U7470 ( .A(DB[855]), .B(DB[840]), .Z(n5665) );
  AND U7471 ( .A(n286), .B(n5666), .Z(n5664) );
  XOR U7472 ( .A(n5667), .B(n5668), .Z(n5666) );
  XOR U7473 ( .A(DB[840]), .B(DB[825]), .Z(n5668) );
  AND U7474 ( .A(n290), .B(n5669), .Z(n5667) );
  XOR U7475 ( .A(n5670), .B(n5671), .Z(n5669) );
  XOR U7476 ( .A(DB[825]), .B(DB[810]), .Z(n5671) );
  AND U7477 ( .A(n294), .B(n5672), .Z(n5670) );
  XOR U7478 ( .A(n5673), .B(n5674), .Z(n5672) );
  XOR U7479 ( .A(DB[810]), .B(DB[795]), .Z(n5674) );
  AND U7480 ( .A(n298), .B(n5675), .Z(n5673) );
  XOR U7481 ( .A(n5676), .B(n5677), .Z(n5675) );
  XOR U7482 ( .A(DB[795]), .B(DB[780]), .Z(n5677) );
  AND U7483 ( .A(n302), .B(n5678), .Z(n5676) );
  XOR U7484 ( .A(n5679), .B(n5680), .Z(n5678) );
  XOR U7485 ( .A(DB[780]), .B(DB[765]), .Z(n5680) );
  AND U7486 ( .A(n306), .B(n5681), .Z(n5679) );
  XOR U7487 ( .A(n5682), .B(n5683), .Z(n5681) );
  XOR U7488 ( .A(DB[765]), .B(DB[750]), .Z(n5683) );
  AND U7489 ( .A(n310), .B(n5684), .Z(n5682) );
  XOR U7490 ( .A(n5685), .B(n5686), .Z(n5684) );
  XOR U7491 ( .A(DB[750]), .B(DB[735]), .Z(n5686) );
  AND U7492 ( .A(n314), .B(n5687), .Z(n5685) );
  XOR U7493 ( .A(n5688), .B(n5689), .Z(n5687) );
  XOR U7494 ( .A(DB[735]), .B(DB[720]), .Z(n5689) );
  AND U7495 ( .A(n318), .B(n5690), .Z(n5688) );
  XOR U7496 ( .A(n5691), .B(n5692), .Z(n5690) );
  XOR U7497 ( .A(DB[720]), .B(DB[705]), .Z(n5692) );
  AND U7498 ( .A(n322), .B(n5693), .Z(n5691) );
  XOR U7499 ( .A(n5694), .B(n5695), .Z(n5693) );
  XOR U7500 ( .A(DB[705]), .B(DB[690]), .Z(n5695) );
  AND U7501 ( .A(n326), .B(n5696), .Z(n5694) );
  XOR U7502 ( .A(n5697), .B(n5698), .Z(n5696) );
  XOR U7503 ( .A(DB[690]), .B(DB[675]), .Z(n5698) );
  AND U7504 ( .A(n330), .B(n5699), .Z(n5697) );
  XOR U7505 ( .A(n5700), .B(n5701), .Z(n5699) );
  XOR U7506 ( .A(DB[675]), .B(DB[660]), .Z(n5701) );
  AND U7507 ( .A(n334), .B(n5702), .Z(n5700) );
  XOR U7508 ( .A(n5703), .B(n5704), .Z(n5702) );
  XOR U7509 ( .A(DB[660]), .B(DB[645]), .Z(n5704) );
  AND U7510 ( .A(n338), .B(n5705), .Z(n5703) );
  XOR U7511 ( .A(n5706), .B(n5707), .Z(n5705) );
  XOR U7512 ( .A(DB[645]), .B(DB[630]), .Z(n5707) );
  AND U7513 ( .A(n342), .B(n5708), .Z(n5706) );
  XOR U7514 ( .A(n5709), .B(n5710), .Z(n5708) );
  XOR U7515 ( .A(DB[630]), .B(DB[615]), .Z(n5710) );
  AND U7516 ( .A(n346), .B(n5711), .Z(n5709) );
  XOR U7517 ( .A(n5712), .B(n5713), .Z(n5711) );
  XOR U7518 ( .A(DB[615]), .B(DB[600]), .Z(n5713) );
  AND U7519 ( .A(n350), .B(n5714), .Z(n5712) );
  XOR U7520 ( .A(n5715), .B(n5716), .Z(n5714) );
  XOR U7521 ( .A(DB[600]), .B(DB[585]), .Z(n5716) );
  AND U7522 ( .A(n354), .B(n5717), .Z(n5715) );
  XOR U7523 ( .A(n5718), .B(n5719), .Z(n5717) );
  XOR U7524 ( .A(DB[585]), .B(DB[570]), .Z(n5719) );
  AND U7525 ( .A(n358), .B(n5720), .Z(n5718) );
  XOR U7526 ( .A(n5721), .B(n5722), .Z(n5720) );
  XOR U7527 ( .A(DB[570]), .B(DB[555]), .Z(n5722) );
  AND U7528 ( .A(n362), .B(n5723), .Z(n5721) );
  XOR U7529 ( .A(n5724), .B(n5725), .Z(n5723) );
  XOR U7530 ( .A(DB[555]), .B(DB[540]), .Z(n5725) );
  AND U7531 ( .A(n366), .B(n5726), .Z(n5724) );
  XOR U7532 ( .A(n5727), .B(n5728), .Z(n5726) );
  XOR U7533 ( .A(DB[540]), .B(DB[525]), .Z(n5728) );
  AND U7534 ( .A(n370), .B(n5729), .Z(n5727) );
  XOR U7535 ( .A(n5730), .B(n5731), .Z(n5729) );
  XOR U7536 ( .A(DB[525]), .B(DB[510]), .Z(n5731) );
  AND U7537 ( .A(n374), .B(n5732), .Z(n5730) );
  XOR U7538 ( .A(n5733), .B(n5734), .Z(n5732) );
  XOR U7539 ( .A(DB[510]), .B(DB[495]), .Z(n5734) );
  AND U7540 ( .A(n378), .B(n5735), .Z(n5733) );
  XOR U7541 ( .A(n5736), .B(n5737), .Z(n5735) );
  XOR U7542 ( .A(DB[495]), .B(DB[480]), .Z(n5737) );
  AND U7543 ( .A(n382), .B(n5738), .Z(n5736) );
  XOR U7544 ( .A(n5739), .B(n5740), .Z(n5738) );
  XOR U7545 ( .A(DB[480]), .B(DB[465]), .Z(n5740) );
  AND U7546 ( .A(n386), .B(n5741), .Z(n5739) );
  XOR U7547 ( .A(n5742), .B(n5743), .Z(n5741) );
  XOR U7548 ( .A(DB[465]), .B(DB[450]), .Z(n5743) );
  AND U7549 ( .A(n390), .B(n5744), .Z(n5742) );
  XOR U7550 ( .A(n5745), .B(n5746), .Z(n5744) );
  XOR U7551 ( .A(DB[450]), .B(DB[435]), .Z(n5746) );
  AND U7552 ( .A(n394), .B(n5747), .Z(n5745) );
  XOR U7553 ( .A(n5748), .B(n5749), .Z(n5747) );
  XOR U7554 ( .A(DB[435]), .B(DB[420]), .Z(n5749) );
  AND U7555 ( .A(n398), .B(n5750), .Z(n5748) );
  XOR U7556 ( .A(n5751), .B(n5752), .Z(n5750) );
  XOR U7557 ( .A(DB[420]), .B(DB[405]), .Z(n5752) );
  AND U7558 ( .A(n402), .B(n5753), .Z(n5751) );
  XOR U7559 ( .A(n5754), .B(n5755), .Z(n5753) );
  XOR U7560 ( .A(DB[405]), .B(DB[390]), .Z(n5755) );
  AND U7561 ( .A(n406), .B(n5756), .Z(n5754) );
  XOR U7562 ( .A(n5757), .B(n5758), .Z(n5756) );
  XOR U7563 ( .A(DB[390]), .B(DB[375]), .Z(n5758) );
  AND U7564 ( .A(n410), .B(n5759), .Z(n5757) );
  XOR U7565 ( .A(n5760), .B(n5761), .Z(n5759) );
  XOR U7566 ( .A(DB[375]), .B(DB[360]), .Z(n5761) );
  AND U7567 ( .A(n414), .B(n5762), .Z(n5760) );
  XOR U7568 ( .A(n5763), .B(n5764), .Z(n5762) );
  XOR U7569 ( .A(DB[360]), .B(DB[345]), .Z(n5764) );
  AND U7570 ( .A(n418), .B(n5765), .Z(n5763) );
  XOR U7571 ( .A(n5766), .B(n5767), .Z(n5765) );
  XOR U7572 ( .A(DB[345]), .B(DB[330]), .Z(n5767) );
  AND U7573 ( .A(n422), .B(n5768), .Z(n5766) );
  XOR U7574 ( .A(n5769), .B(n5770), .Z(n5768) );
  XOR U7575 ( .A(DB[330]), .B(DB[315]), .Z(n5770) );
  AND U7576 ( .A(n426), .B(n5771), .Z(n5769) );
  XOR U7577 ( .A(n5772), .B(n5773), .Z(n5771) );
  XOR U7578 ( .A(DB[315]), .B(DB[300]), .Z(n5773) );
  AND U7579 ( .A(n430), .B(n5774), .Z(n5772) );
  XOR U7580 ( .A(n5775), .B(n5776), .Z(n5774) );
  XOR U7581 ( .A(DB[300]), .B(DB[285]), .Z(n5776) );
  AND U7582 ( .A(n434), .B(n5777), .Z(n5775) );
  XOR U7583 ( .A(n5778), .B(n5779), .Z(n5777) );
  XOR U7584 ( .A(DB[285]), .B(DB[270]), .Z(n5779) );
  AND U7585 ( .A(n438), .B(n5780), .Z(n5778) );
  XOR U7586 ( .A(n5781), .B(n5782), .Z(n5780) );
  XOR U7587 ( .A(DB[270]), .B(DB[255]), .Z(n5782) );
  AND U7588 ( .A(n442), .B(n5783), .Z(n5781) );
  XOR U7589 ( .A(n5784), .B(n5785), .Z(n5783) );
  XOR U7590 ( .A(DB[255]), .B(DB[240]), .Z(n5785) );
  AND U7591 ( .A(n446), .B(n5786), .Z(n5784) );
  XOR U7592 ( .A(n5787), .B(n5788), .Z(n5786) );
  XOR U7593 ( .A(DB[240]), .B(DB[225]), .Z(n5788) );
  AND U7594 ( .A(n450), .B(n5789), .Z(n5787) );
  XOR U7595 ( .A(n5790), .B(n5791), .Z(n5789) );
  XOR U7596 ( .A(DB[225]), .B(DB[210]), .Z(n5791) );
  AND U7597 ( .A(n454), .B(n5792), .Z(n5790) );
  XOR U7598 ( .A(n5793), .B(n5794), .Z(n5792) );
  XOR U7599 ( .A(DB[210]), .B(DB[195]), .Z(n5794) );
  AND U7600 ( .A(n458), .B(n5795), .Z(n5793) );
  XOR U7601 ( .A(n5796), .B(n5797), .Z(n5795) );
  XOR U7602 ( .A(DB[195]), .B(DB[180]), .Z(n5797) );
  AND U7603 ( .A(n462), .B(n5798), .Z(n5796) );
  XOR U7604 ( .A(n5799), .B(n5800), .Z(n5798) );
  XOR U7605 ( .A(DB[180]), .B(DB[165]), .Z(n5800) );
  AND U7606 ( .A(n466), .B(n5801), .Z(n5799) );
  XOR U7607 ( .A(n5802), .B(n5803), .Z(n5801) );
  XOR U7608 ( .A(DB[165]), .B(DB[150]), .Z(n5803) );
  AND U7609 ( .A(n470), .B(n5804), .Z(n5802) );
  XOR U7610 ( .A(n5805), .B(n5806), .Z(n5804) );
  XOR U7611 ( .A(DB[150]), .B(DB[135]), .Z(n5806) );
  AND U7612 ( .A(n474), .B(n5807), .Z(n5805) );
  XOR U7613 ( .A(n5808), .B(n5809), .Z(n5807) );
  XOR U7614 ( .A(DB[135]), .B(DB[120]), .Z(n5809) );
  AND U7615 ( .A(n478), .B(n5810), .Z(n5808) );
  XOR U7616 ( .A(n5811), .B(n5812), .Z(n5810) );
  XOR U7617 ( .A(DB[120]), .B(DB[105]), .Z(n5812) );
  AND U7618 ( .A(n482), .B(n5813), .Z(n5811) );
  XOR U7619 ( .A(n5814), .B(n5815), .Z(n5813) );
  XOR U7620 ( .A(DB[90]), .B(DB[105]), .Z(n5815) );
  AND U7621 ( .A(n486), .B(n5816), .Z(n5814) );
  XOR U7622 ( .A(n5817), .B(n5818), .Z(n5816) );
  XOR U7623 ( .A(DB[90]), .B(DB[75]), .Z(n5818) );
  AND U7624 ( .A(n490), .B(n5819), .Z(n5817) );
  XOR U7625 ( .A(n5820), .B(n5821), .Z(n5819) );
  XOR U7626 ( .A(DB[75]), .B(DB[60]), .Z(n5821) );
  AND U7627 ( .A(n494), .B(n5822), .Z(n5820) );
  XOR U7628 ( .A(n5823), .B(n5824), .Z(n5822) );
  XOR U7629 ( .A(DB[60]), .B(DB[45]), .Z(n5824) );
  AND U7630 ( .A(n498), .B(n5825), .Z(n5823) );
  XOR U7631 ( .A(n5826), .B(n5827), .Z(n5825) );
  XOR U7632 ( .A(DB[45]), .B(DB[30]), .Z(n5827) );
  AND U7633 ( .A(n502), .B(n5828), .Z(n5826) );
  XOR U7634 ( .A(n5829), .B(n5830), .Z(n5828) );
  XOR U7635 ( .A(DB[30]), .B(DB[15]), .Z(n5830) );
  AND U7636 ( .A(n506), .B(n5831), .Z(n5829) );
  XOR U7637 ( .A(DB[15]), .B(DB[0]), .Z(n5831) );
  XNOR U7638 ( .A(n5832), .B(n5833), .Z(n2) );
  AND U7639 ( .A(n5834), .B(n5835), .Z(n5832) );
  XOR U7640 ( .A(n5833), .B(n5836), .Z(n5835) );
  XOR U7641 ( .A(n5837), .B(n5838), .Z(n5836) );
  AND U7642 ( .A(n5839), .B(n5840), .Z(n5837) );
  XNOR U7643 ( .A(n5841), .B(n5842), .Z(n5840) );
  XOR U7644 ( .A(n5833), .B(n5843), .Z(n5834) );
  XNOR U7645 ( .A(n5844), .B(n5845), .Z(n5843) );
  AND U7646 ( .A(n6), .B(n5846), .Z(n5844) );
  XOR U7647 ( .A(n5847), .B(n5845), .Z(n5846) );
  XNOR U7648 ( .A(n5848), .B(n5849), .Z(n5833) );
  AND U7649 ( .A(n5850), .B(n5851), .Z(n5848) );
  XOR U7650 ( .A(n5839), .B(n5852), .Z(n5851) );
  XNOR U7651 ( .A(n5849), .B(n5841), .Z(n5852) );
  XNOR U7652 ( .A(n5853), .B(n5854), .Z(n5841) );
  ANDN U7653 ( .B(n5855), .A(n5856), .Z(n5853) );
  XOR U7654 ( .A(n5854), .B(n5857), .Z(n5855) );
  XNOR U7655 ( .A(n5838), .B(n5858), .Z(n5839) );
  XNOR U7656 ( .A(n5859), .B(n5860), .Z(n5858) );
  ANDN U7657 ( .B(n5861), .A(n5862), .Z(n5859) );
  XNOR U7658 ( .A(n5863), .B(n5864), .Z(n5861) );
  IV U7659 ( .A(n5842), .Z(n5838) );
  XOR U7660 ( .A(n5865), .B(n5866), .Z(n5842) );
  AND U7661 ( .A(n5867), .B(n5868), .Z(n5865) );
  XOR U7662 ( .A(n5869), .B(n5866), .Z(n5868) );
  XNOR U7663 ( .A(n5849), .B(n5870), .Z(n5850) );
  XOR U7664 ( .A(n5871), .B(n5872), .Z(n5870) );
  AND U7665 ( .A(n6), .B(n5873), .Z(n5871) );
  XNOR U7666 ( .A(n5874), .B(n5872), .Z(n5873) );
  XNOR U7667 ( .A(n5875), .B(n5876), .Z(n5849) );
  NAND U7668 ( .A(n5877), .B(n5878), .Z(n5876) );
  XOR U7669 ( .A(n5867), .B(n5879), .Z(n5878) );
  XOR U7670 ( .A(n5875), .B(n5869), .Z(n5879) );
  XOR U7671 ( .A(n5880), .B(n5857), .Z(n5869) );
  XNOR U7672 ( .A(n5881), .B(n5882), .Z(n5857) );
  ANDN U7673 ( .B(n5883), .A(n5884), .Z(n5881) );
  XNOR U7674 ( .A(n5882), .B(n5885), .Z(n5883) );
  IV U7675 ( .A(n5856), .Z(n5880) );
  XOR U7676 ( .A(n5886), .B(n5887), .Z(n5856) );
  XNOR U7677 ( .A(n5888), .B(n5889), .Z(n5887) );
  ANDN U7678 ( .B(n5890), .A(n5891), .Z(n5888) );
  XNOR U7679 ( .A(n5892), .B(n5893), .Z(n5890) );
  IV U7680 ( .A(n5889), .Z(n5893) );
  IV U7681 ( .A(n5854), .Z(n5886) );
  XNOR U7682 ( .A(n5894), .B(n5895), .Z(n5854) );
  ANDN U7683 ( .B(n5896), .A(n5897), .Z(n5894) );
  XNOR U7684 ( .A(n5895), .B(n5898), .Z(n5896) );
  XNOR U7685 ( .A(n5899), .B(n5900), .Z(n5867) );
  XNOR U7686 ( .A(n5863), .B(n5901), .Z(n5900) );
  IV U7687 ( .A(n5866), .Z(n5901) );
  XNOR U7688 ( .A(n5902), .B(n5903), .Z(n5866) );
  AND U7689 ( .A(n5904), .B(n5905), .Z(n5902) );
  XNOR U7690 ( .A(n5903), .B(n5906), .Z(n5905) );
  XOR U7691 ( .A(n5907), .B(n5908), .Z(n5863) );
  ANDN U7692 ( .B(n5909), .A(n5910), .Z(n5907) );
  XNOR U7693 ( .A(n5908), .B(n5911), .Z(n5909) );
  IV U7694 ( .A(n5862), .Z(n5899) );
  XOR U7695 ( .A(n5860), .B(n5912), .Z(n5862) );
  XNOR U7696 ( .A(n5913), .B(n5914), .Z(n5912) );
  ANDN U7697 ( .B(n5915), .A(n5916), .Z(n5913) );
  XNOR U7698 ( .A(n5917), .B(n5918), .Z(n5915) );
  IV U7699 ( .A(n5914), .Z(n5918) );
  IV U7700 ( .A(n5864), .Z(n5860) );
  XNOR U7701 ( .A(n5919), .B(n5920), .Z(n5864) );
  ANDN U7702 ( .B(n5921), .A(n5922), .Z(n5919) );
  XNOR U7703 ( .A(n5923), .B(n5920), .Z(n5921) );
  XOR U7704 ( .A(n5924), .B(n5925), .Z(n5877) );
  XNOR U7705 ( .A(n5875), .B(n5926), .Z(n5925) );
  NAND U7706 ( .A(n5927), .B(n6), .Z(n5926) );
  XOR U7707 ( .A(n5928), .B(n5924), .Z(n5927) );
  NAND U7708 ( .A(n5929), .B(n5930), .Z(n5875) );
  XNOR U7709 ( .A(n5904), .B(n5906), .Z(n5930) );
  XOR U7710 ( .A(n5931), .B(n5898), .Z(n5906) );
  XOR U7711 ( .A(n5932), .B(n5885), .Z(n5898) );
  XNOR U7712 ( .A(q[14]), .B(DB[1919]), .Z(n5885) );
  IV U7713 ( .A(n5884), .Z(n5932) );
  XOR U7714 ( .A(n5882), .B(n5933), .Z(n5884) );
  XNOR U7715 ( .A(q[13]), .B(DB[1918]), .Z(n5933) );
  XOR U7716 ( .A(q[12]), .B(DB[1917]), .Z(n5882) );
  IV U7717 ( .A(n5897), .Z(n5931) );
  XOR U7718 ( .A(n5934), .B(n5935), .Z(n5897) );
  XNOR U7719 ( .A(n5892), .B(n5895), .Z(n5935) );
  XOR U7720 ( .A(q[8]), .B(DB[1913]), .Z(n5895) );
  XOR U7721 ( .A(q[11]), .B(DB[1916]), .Z(n5892) );
  IV U7722 ( .A(n5891), .Z(n5934) );
  XOR U7723 ( .A(n5889), .B(n5936), .Z(n5891) );
  XNOR U7724 ( .A(q[10]), .B(DB[1915]), .Z(n5936) );
  XOR U7725 ( .A(q[9]), .B(DB[1914]), .Z(n5889) );
  XNOR U7726 ( .A(n5937), .B(n5938), .Z(n5904) );
  XOR U7727 ( .A(n5923), .B(n5903), .Z(n5938) );
  XOR U7728 ( .A(q[0]), .B(DB[1905]), .Z(n5903) );
  XOR U7729 ( .A(n5939), .B(n5911), .Z(n5923) );
  XNOR U7730 ( .A(q[7]), .B(DB[1912]), .Z(n5911) );
  IV U7731 ( .A(n5910), .Z(n5939) );
  XOR U7732 ( .A(n5908), .B(n5940), .Z(n5910) );
  XNOR U7733 ( .A(q[6]), .B(DB[1911]), .Z(n5940) );
  XOR U7734 ( .A(q[5]), .B(DB[1910]), .Z(n5908) );
  IV U7735 ( .A(n5922), .Z(n5937) );
  XOR U7736 ( .A(n5941), .B(n5942), .Z(n5922) );
  XNOR U7737 ( .A(n5917), .B(n5920), .Z(n5942) );
  XOR U7738 ( .A(q[1]), .B(DB[1906]), .Z(n5920) );
  XOR U7739 ( .A(q[4]), .B(DB[1909]), .Z(n5917) );
  IV U7740 ( .A(n5916), .Z(n5941) );
  XOR U7741 ( .A(n5914), .B(n5943), .Z(n5916) );
  XNOR U7742 ( .A(q[3]), .B(DB[1908]), .Z(n5943) );
  XOR U7743 ( .A(q[2]), .B(DB[1907]), .Z(n5914) );
  XOR U7744 ( .A(n5944), .B(n5945), .Z(n5929) );
  AND U7745 ( .A(n6), .B(n5946), .Z(n5944) );
  XOR U7746 ( .A(n5945), .B(n5947), .Z(n5946) );
  XNOR U7747 ( .A(n5948), .B(n5949), .Z(n6) );
  AND U7748 ( .A(n5950), .B(n5951), .Z(n5948) );
  XOR U7749 ( .A(n5949), .B(n5845), .Z(n5951) );
  XNOR U7750 ( .A(n5952), .B(n5953), .Z(n5845) );
  ANDN U7751 ( .B(n5954), .A(n5955), .Z(n5952) );
  XOR U7752 ( .A(n5953), .B(n5956), .Z(n5954) );
  XNOR U7753 ( .A(n5949), .B(n5847), .Z(n5950) );
  XOR U7754 ( .A(n5957), .B(n5958), .Z(n5847) );
  AND U7755 ( .A(n10), .B(n5959), .Z(n5957) );
  XOR U7756 ( .A(n5960), .B(n5958), .Z(n5959) );
  XNOR U7757 ( .A(n5961), .B(n5962), .Z(n5949) );
  AND U7758 ( .A(n5963), .B(n5964), .Z(n5961) );
  XOR U7759 ( .A(n5962), .B(n5872), .Z(n5964) );
  XOR U7760 ( .A(n5965), .B(n5956), .Z(n5872) );
  XNOR U7761 ( .A(n5966), .B(n5967), .Z(n5956) );
  ANDN U7762 ( .B(n5968), .A(n5969), .Z(n5966) );
  XOR U7763 ( .A(n5970), .B(n5971), .Z(n5968) );
  IV U7764 ( .A(n5955), .Z(n5965) );
  XOR U7765 ( .A(n5972), .B(n5973), .Z(n5955) );
  XNOR U7766 ( .A(n5974), .B(n5975), .Z(n5973) );
  ANDN U7767 ( .B(n5976), .A(n5977), .Z(n5974) );
  XNOR U7768 ( .A(n5978), .B(n5979), .Z(n5976) );
  IV U7769 ( .A(n5953), .Z(n5972) );
  XOR U7770 ( .A(n5980), .B(n5981), .Z(n5953) );
  ANDN U7771 ( .B(n5982), .A(n5983), .Z(n5980) );
  XOR U7772 ( .A(n5981), .B(n5984), .Z(n5982) );
  XOR U7773 ( .A(n5962), .B(n5874), .Z(n5963) );
  XOR U7774 ( .A(n5985), .B(n5986), .Z(n5874) );
  AND U7775 ( .A(n10), .B(n5987), .Z(n5985) );
  XOR U7776 ( .A(n5988), .B(n5986), .Z(n5987) );
  XNOR U7777 ( .A(n5989), .B(n5990), .Z(n5962) );
  NAND U7778 ( .A(n5991), .B(n5992), .Z(n5990) );
  XOR U7779 ( .A(n5993), .B(n5924), .Z(n5992) );
  XNOR U7780 ( .A(n5994), .B(n5984), .Z(n5924) );
  XOR U7781 ( .A(n5995), .B(n5971), .Z(n5984) );
  XOR U7782 ( .A(n5996), .B(n5997), .Z(n5971) );
  ANDN U7783 ( .B(n5998), .A(n5999), .Z(n5996) );
  XOR U7784 ( .A(n5997), .B(n6000), .Z(n5998) );
  IV U7785 ( .A(n5969), .Z(n5995) );
  XOR U7786 ( .A(n5967), .B(n6001), .Z(n5969) );
  XOR U7787 ( .A(n6002), .B(n6003), .Z(n6001) );
  ANDN U7788 ( .B(n6004), .A(n6005), .Z(n6002) );
  XOR U7789 ( .A(n6006), .B(n6003), .Z(n6004) );
  IV U7790 ( .A(n5970), .Z(n5967) );
  XOR U7791 ( .A(n6007), .B(n6008), .Z(n5970) );
  ANDN U7792 ( .B(n6009), .A(n6010), .Z(n6007) );
  XOR U7793 ( .A(n6008), .B(n6011), .Z(n6009) );
  IV U7794 ( .A(n5983), .Z(n5994) );
  XOR U7795 ( .A(n6012), .B(n6013), .Z(n5983) );
  XNOR U7796 ( .A(n5978), .B(n6014), .Z(n6013) );
  IV U7797 ( .A(n5981), .Z(n6014) );
  XOR U7798 ( .A(n6015), .B(n6016), .Z(n5981) );
  ANDN U7799 ( .B(n6017), .A(n6018), .Z(n6015) );
  XOR U7800 ( .A(n6016), .B(n6019), .Z(n6017) );
  XNOR U7801 ( .A(n6020), .B(n6021), .Z(n5978) );
  ANDN U7802 ( .B(n6022), .A(n6023), .Z(n6020) );
  XOR U7803 ( .A(n6021), .B(n6024), .Z(n6022) );
  IV U7804 ( .A(n5977), .Z(n6012) );
  XOR U7805 ( .A(n5975), .B(n6025), .Z(n5977) );
  XOR U7806 ( .A(n6026), .B(n6027), .Z(n6025) );
  ANDN U7807 ( .B(n6028), .A(n6029), .Z(n6026) );
  XOR U7808 ( .A(n6030), .B(n6027), .Z(n6028) );
  IV U7809 ( .A(n5979), .Z(n5975) );
  XOR U7810 ( .A(n6031), .B(n6032), .Z(n5979) );
  ANDN U7811 ( .B(n6033), .A(n6034), .Z(n6031) );
  XOR U7812 ( .A(n6035), .B(n6032), .Z(n6033) );
  IV U7813 ( .A(n5989), .Z(n5993) );
  XOR U7814 ( .A(n5989), .B(n5928), .Z(n5991) );
  XOR U7815 ( .A(n6036), .B(n6037), .Z(n5928) );
  AND U7816 ( .A(n10), .B(n6038), .Z(n6036) );
  XOR U7817 ( .A(n6039), .B(n6037), .Z(n6038) );
  NANDN U7818 ( .A(n5945), .B(n5947), .Z(n5989) );
  XOR U7819 ( .A(n6040), .B(n6041), .Z(n5947) );
  AND U7820 ( .A(n10), .B(n6042), .Z(n6040) );
  XOR U7821 ( .A(n6041), .B(n6043), .Z(n6042) );
  XNOR U7822 ( .A(n6044), .B(n6045), .Z(n10) );
  AND U7823 ( .A(n6046), .B(n6047), .Z(n6044) );
  XOR U7824 ( .A(n6045), .B(n5958), .Z(n6047) );
  XNOR U7825 ( .A(n6048), .B(n6049), .Z(n5958) );
  ANDN U7826 ( .B(n6050), .A(n6051), .Z(n6048) );
  XOR U7827 ( .A(n6049), .B(n6052), .Z(n6050) );
  XNOR U7828 ( .A(n6045), .B(n5960), .Z(n6046) );
  XOR U7829 ( .A(n6053), .B(n6054), .Z(n5960) );
  AND U7830 ( .A(n14), .B(n6055), .Z(n6053) );
  XOR U7831 ( .A(n6056), .B(n6054), .Z(n6055) );
  XNOR U7832 ( .A(n6057), .B(n6058), .Z(n6045) );
  AND U7833 ( .A(n6059), .B(n6060), .Z(n6057) );
  XNOR U7834 ( .A(n6058), .B(n5986), .Z(n6060) );
  XOR U7835 ( .A(n6051), .B(n6052), .Z(n5986) );
  XNOR U7836 ( .A(n6061), .B(n6062), .Z(n6052) );
  ANDN U7837 ( .B(n6063), .A(n6064), .Z(n6061) );
  XOR U7838 ( .A(n6065), .B(n6066), .Z(n6063) );
  XOR U7839 ( .A(n6067), .B(n6068), .Z(n6051) );
  XNOR U7840 ( .A(n6069), .B(n6070), .Z(n6068) );
  ANDN U7841 ( .B(n6071), .A(n6072), .Z(n6069) );
  XNOR U7842 ( .A(n6073), .B(n6074), .Z(n6071) );
  IV U7843 ( .A(n6049), .Z(n6067) );
  XOR U7844 ( .A(n6075), .B(n6076), .Z(n6049) );
  ANDN U7845 ( .B(n6077), .A(n6078), .Z(n6075) );
  XOR U7846 ( .A(n6076), .B(n6079), .Z(n6077) );
  XOR U7847 ( .A(n6058), .B(n5988), .Z(n6059) );
  XOR U7848 ( .A(n6080), .B(n6081), .Z(n5988) );
  AND U7849 ( .A(n14), .B(n6082), .Z(n6080) );
  XOR U7850 ( .A(n6083), .B(n6081), .Z(n6082) );
  XNOR U7851 ( .A(n6084), .B(n6085), .Z(n6058) );
  NAND U7852 ( .A(n6086), .B(n6087), .Z(n6085) );
  XOR U7853 ( .A(n6088), .B(n6037), .Z(n6087) );
  XOR U7854 ( .A(n6078), .B(n6079), .Z(n6037) );
  XOR U7855 ( .A(n6089), .B(n6066), .Z(n6079) );
  XOR U7856 ( .A(n6090), .B(n6091), .Z(n6066) );
  ANDN U7857 ( .B(n6092), .A(n6093), .Z(n6090) );
  XOR U7858 ( .A(n6091), .B(n6094), .Z(n6092) );
  IV U7859 ( .A(n6064), .Z(n6089) );
  XOR U7860 ( .A(n6062), .B(n6095), .Z(n6064) );
  XOR U7861 ( .A(n6096), .B(n6097), .Z(n6095) );
  ANDN U7862 ( .B(n6098), .A(n6099), .Z(n6096) );
  XOR U7863 ( .A(n6100), .B(n6097), .Z(n6098) );
  IV U7864 ( .A(n6065), .Z(n6062) );
  XOR U7865 ( .A(n6101), .B(n6102), .Z(n6065) );
  ANDN U7866 ( .B(n6103), .A(n6104), .Z(n6101) );
  XOR U7867 ( .A(n6102), .B(n6105), .Z(n6103) );
  XOR U7868 ( .A(n6106), .B(n6107), .Z(n6078) );
  XNOR U7869 ( .A(n6073), .B(n6108), .Z(n6107) );
  IV U7870 ( .A(n6076), .Z(n6108) );
  XOR U7871 ( .A(n6109), .B(n6110), .Z(n6076) );
  ANDN U7872 ( .B(n6111), .A(n6112), .Z(n6109) );
  XOR U7873 ( .A(n6110), .B(n6113), .Z(n6111) );
  XNOR U7874 ( .A(n6114), .B(n6115), .Z(n6073) );
  ANDN U7875 ( .B(n6116), .A(n6117), .Z(n6114) );
  XOR U7876 ( .A(n6115), .B(n6118), .Z(n6116) );
  IV U7877 ( .A(n6072), .Z(n6106) );
  XOR U7878 ( .A(n6070), .B(n6119), .Z(n6072) );
  XOR U7879 ( .A(n6120), .B(n6121), .Z(n6119) );
  ANDN U7880 ( .B(n6122), .A(n6123), .Z(n6120) );
  XOR U7881 ( .A(n6124), .B(n6121), .Z(n6122) );
  IV U7882 ( .A(n6074), .Z(n6070) );
  XOR U7883 ( .A(n6125), .B(n6126), .Z(n6074) );
  ANDN U7884 ( .B(n6127), .A(n6128), .Z(n6125) );
  XOR U7885 ( .A(n6129), .B(n6126), .Z(n6127) );
  IV U7886 ( .A(n6084), .Z(n6088) );
  XOR U7887 ( .A(n6084), .B(n6039), .Z(n6086) );
  XOR U7888 ( .A(n6130), .B(n6131), .Z(n6039) );
  AND U7889 ( .A(n14), .B(n6132), .Z(n6130) );
  XOR U7890 ( .A(n6133), .B(n6131), .Z(n6132) );
  NANDN U7891 ( .A(n6041), .B(n6043), .Z(n6084) );
  XOR U7892 ( .A(n6134), .B(n6135), .Z(n6043) );
  AND U7893 ( .A(n14), .B(n6136), .Z(n6134) );
  XOR U7894 ( .A(n6135), .B(n6137), .Z(n6136) );
  XNOR U7895 ( .A(n6138), .B(n6139), .Z(n14) );
  AND U7896 ( .A(n6140), .B(n6141), .Z(n6138) );
  XOR U7897 ( .A(n6139), .B(n6054), .Z(n6141) );
  XNOR U7898 ( .A(n6142), .B(n6143), .Z(n6054) );
  ANDN U7899 ( .B(n6144), .A(n6145), .Z(n6142) );
  XOR U7900 ( .A(n6143), .B(n6146), .Z(n6144) );
  XNOR U7901 ( .A(n6139), .B(n6056), .Z(n6140) );
  XOR U7902 ( .A(n6147), .B(n6148), .Z(n6056) );
  AND U7903 ( .A(n18), .B(n6149), .Z(n6147) );
  XOR U7904 ( .A(n6150), .B(n6148), .Z(n6149) );
  XNOR U7905 ( .A(n6151), .B(n6152), .Z(n6139) );
  AND U7906 ( .A(n6153), .B(n6154), .Z(n6151) );
  XNOR U7907 ( .A(n6152), .B(n6081), .Z(n6154) );
  XOR U7908 ( .A(n6145), .B(n6146), .Z(n6081) );
  XNOR U7909 ( .A(n6155), .B(n6156), .Z(n6146) );
  ANDN U7910 ( .B(n6157), .A(n6158), .Z(n6155) );
  XOR U7911 ( .A(n6159), .B(n6160), .Z(n6157) );
  XOR U7912 ( .A(n6161), .B(n6162), .Z(n6145) );
  XNOR U7913 ( .A(n6163), .B(n6164), .Z(n6162) );
  ANDN U7914 ( .B(n6165), .A(n6166), .Z(n6163) );
  XNOR U7915 ( .A(n6167), .B(n6168), .Z(n6165) );
  IV U7916 ( .A(n6143), .Z(n6161) );
  XOR U7917 ( .A(n6169), .B(n6170), .Z(n6143) );
  ANDN U7918 ( .B(n6171), .A(n6172), .Z(n6169) );
  XOR U7919 ( .A(n6170), .B(n6173), .Z(n6171) );
  XOR U7920 ( .A(n6152), .B(n6083), .Z(n6153) );
  XOR U7921 ( .A(n6174), .B(n6175), .Z(n6083) );
  AND U7922 ( .A(n18), .B(n6176), .Z(n6174) );
  XOR U7923 ( .A(n6177), .B(n6175), .Z(n6176) );
  XNOR U7924 ( .A(n6178), .B(n6179), .Z(n6152) );
  NAND U7925 ( .A(n6180), .B(n6181), .Z(n6179) );
  XOR U7926 ( .A(n6182), .B(n6131), .Z(n6181) );
  XOR U7927 ( .A(n6172), .B(n6173), .Z(n6131) );
  XOR U7928 ( .A(n6183), .B(n6160), .Z(n6173) );
  XOR U7929 ( .A(n6184), .B(n6185), .Z(n6160) );
  ANDN U7930 ( .B(n6186), .A(n6187), .Z(n6184) );
  XOR U7931 ( .A(n6185), .B(n6188), .Z(n6186) );
  IV U7932 ( .A(n6158), .Z(n6183) );
  XOR U7933 ( .A(n6156), .B(n6189), .Z(n6158) );
  XOR U7934 ( .A(n6190), .B(n6191), .Z(n6189) );
  ANDN U7935 ( .B(n6192), .A(n6193), .Z(n6190) );
  XOR U7936 ( .A(n6194), .B(n6191), .Z(n6192) );
  IV U7937 ( .A(n6159), .Z(n6156) );
  XOR U7938 ( .A(n6195), .B(n6196), .Z(n6159) );
  ANDN U7939 ( .B(n6197), .A(n6198), .Z(n6195) );
  XOR U7940 ( .A(n6196), .B(n6199), .Z(n6197) );
  XOR U7941 ( .A(n6200), .B(n6201), .Z(n6172) );
  XNOR U7942 ( .A(n6167), .B(n6202), .Z(n6201) );
  IV U7943 ( .A(n6170), .Z(n6202) );
  XOR U7944 ( .A(n6203), .B(n6204), .Z(n6170) );
  ANDN U7945 ( .B(n6205), .A(n6206), .Z(n6203) );
  XOR U7946 ( .A(n6204), .B(n6207), .Z(n6205) );
  XNOR U7947 ( .A(n6208), .B(n6209), .Z(n6167) );
  ANDN U7948 ( .B(n6210), .A(n6211), .Z(n6208) );
  XOR U7949 ( .A(n6209), .B(n6212), .Z(n6210) );
  IV U7950 ( .A(n6166), .Z(n6200) );
  XOR U7951 ( .A(n6164), .B(n6213), .Z(n6166) );
  XOR U7952 ( .A(n6214), .B(n6215), .Z(n6213) );
  ANDN U7953 ( .B(n6216), .A(n6217), .Z(n6214) );
  XOR U7954 ( .A(n6218), .B(n6215), .Z(n6216) );
  IV U7955 ( .A(n6168), .Z(n6164) );
  XOR U7956 ( .A(n6219), .B(n6220), .Z(n6168) );
  ANDN U7957 ( .B(n6221), .A(n6222), .Z(n6219) );
  XOR U7958 ( .A(n6223), .B(n6220), .Z(n6221) );
  IV U7959 ( .A(n6178), .Z(n6182) );
  XOR U7960 ( .A(n6178), .B(n6133), .Z(n6180) );
  XOR U7961 ( .A(n6224), .B(n6225), .Z(n6133) );
  AND U7962 ( .A(n18), .B(n6226), .Z(n6224) );
  XOR U7963 ( .A(n6227), .B(n6225), .Z(n6226) );
  NANDN U7964 ( .A(n6135), .B(n6137), .Z(n6178) );
  XOR U7965 ( .A(n6228), .B(n6229), .Z(n6137) );
  AND U7966 ( .A(n18), .B(n6230), .Z(n6228) );
  XOR U7967 ( .A(n6229), .B(n6231), .Z(n6230) );
  XNOR U7968 ( .A(n6232), .B(n6233), .Z(n18) );
  AND U7969 ( .A(n6234), .B(n6235), .Z(n6232) );
  XOR U7970 ( .A(n6233), .B(n6148), .Z(n6235) );
  XNOR U7971 ( .A(n6236), .B(n6237), .Z(n6148) );
  ANDN U7972 ( .B(n6238), .A(n6239), .Z(n6236) );
  XOR U7973 ( .A(n6237), .B(n6240), .Z(n6238) );
  XNOR U7974 ( .A(n6233), .B(n6150), .Z(n6234) );
  XOR U7975 ( .A(n6241), .B(n6242), .Z(n6150) );
  AND U7976 ( .A(n22), .B(n6243), .Z(n6241) );
  XOR U7977 ( .A(n6244), .B(n6242), .Z(n6243) );
  XNOR U7978 ( .A(n6245), .B(n6246), .Z(n6233) );
  AND U7979 ( .A(n6247), .B(n6248), .Z(n6245) );
  XNOR U7980 ( .A(n6246), .B(n6175), .Z(n6248) );
  XOR U7981 ( .A(n6239), .B(n6240), .Z(n6175) );
  XNOR U7982 ( .A(n6249), .B(n6250), .Z(n6240) );
  ANDN U7983 ( .B(n6251), .A(n6252), .Z(n6249) );
  XOR U7984 ( .A(n6253), .B(n6254), .Z(n6251) );
  XOR U7985 ( .A(n6255), .B(n6256), .Z(n6239) );
  XNOR U7986 ( .A(n6257), .B(n6258), .Z(n6256) );
  ANDN U7987 ( .B(n6259), .A(n6260), .Z(n6257) );
  XNOR U7988 ( .A(n6261), .B(n6262), .Z(n6259) );
  IV U7989 ( .A(n6237), .Z(n6255) );
  XOR U7990 ( .A(n6263), .B(n6264), .Z(n6237) );
  ANDN U7991 ( .B(n6265), .A(n6266), .Z(n6263) );
  XOR U7992 ( .A(n6264), .B(n6267), .Z(n6265) );
  XOR U7993 ( .A(n6246), .B(n6177), .Z(n6247) );
  XOR U7994 ( .A(n6268), .B(n6269), .Z(n6177) );
  AND U7995 ( .A(n22), .B(n6270), .Z(n6268) );
  XOR U7996 ( .A(n6271), .B(n6269), .Z(n6270) );
  XNOR U7997 ( .A(n6272), .B(n6273), .Z(n6246) );
  NAND U7998 ( .A(n6274), .B(n6275), .Z(n6273) );
  XOR U7999 ( .A(n6276), .B(n6225), .Z(n6275) );
  XOR U8000 ( .A(n6266), .B(n6267), .Z(n6225) );
  XOR U8001 ( .A(n6277), .B(n6254), .Z(n6267) );
  XOR U8002 ( .A(n6278), .B(n6279), .Z(n6254) );
  ANDN U8003 ( .B(n6280), .A(n6281), .Z(n6278) );
  XOR U8004 ( .A(n6279), .B(n6282), .Z(n6280) );
  IV U8005 ( .A(n6252), .Z(n6277) );
  XOR U8006 ( .A(n6250), .B(n6283), .Z(n6252) );
  XOR U8007 ( .A(n6284), .B(n6285), .Z(n6283) );
  ANDN U8008 ( .B(n6286), .A(n6287), .Z(n6284) );
  XOR U8009 ( .A(n6288), .B(n6285), .Z(n6286) );
  IV U8010 ( .A(n6253), .Z(n6250) );
  XOR U8011 ( .A(n6289), .B(n6290), .Z(n6253) );
  ANDN U8012 ( .B(n6291), .A(n6292), .Z(n6289) );
  XOR U8013 ( .A(n6290), .B(n6293), .Z(n6291) );
  XOR U8014 ( .A(n6294), .B(n6295), .Z(n6266) );
  XNOR U8015 ( .A(n6261), .B(n6296), .Z(n6295) );
  IV U8016 ( .A(n6264), .Z(n6296) );
  XOR U8017 ( .A(n6297), .B(n6298), .Z(n6264) );
  ANDN U8018 ( .B(n6299), .A(n6300), .Z(n6297) );
  XOR U8019 ( .A(n6298), .B(n6301), .Z(n6299) );
  XNOR U8020 ( .A(n6302), .B(n6303), .Z(n6261) );
  ANDN U8021 ( .B(n6304), .A(n6305), .Z(n6302) );
  XOR U8022 ( .A(n6303), .B(n6306), .Z(n6304) );
  IV U8023 ( .A(n6260), .Z(n6294) );
  XOR U8024 ( .A(n6258), .B(n6307), .Z(n6260) );
  XOR U8025 ( .A(n6308), .B(n6309), .Z(n6307) );
  ANDN U8026 ( .B(n6310), .A(n6311), .Z(n6308) );
  XOR U8027 ( .A(n6312), .B(n6309), .Z(n6310) );
  IV U8028 ( .A(n6262), .Z(n6258) );
  XOR U8029 ( .A(n6313), .B(n6314), .Z(n6262) );
  ANDN U8030 ( .B(n6315), .A(n6316), .Z(n6313) );
  XOR U8031 ( .A(n6317), .B(n6314), .Z(n6315) );
  IV U8032 ( .A(n6272), .Z(n6276) );
  XOR U8033 ( .A(n6272), .B(n6227), .Z(n6274) );
  XOR U8034 ( .A(n6318), .B(n6319), .Z(n6227) );
  AND U8035 ( .A(n22), .B(n6320), .Z(n6318) );
  XOR U8036 ( .A(n6321), .B(n6319), .Z(n6320) );
  NANDN U8037 ( .A(n6229), .B(n6231), .Z(n6272) );
  XOR U8038 ( .A(n6322), .B(n6323), .Z(n6231) );
  AND U8039 ( .A(n22), .B(n6324), .Z(n6322) );
  XOR U8040 ( .A(n6323), .B(n6325), .Z(n6324) );
  XNOR U8041 ( .A(n6326), .B(n6327), .Z(n22) );
  AND U8042 ( .A(n6328), .B(n6329), .Z(n6326) );
  XOR U8043 ( .A(n6327), .B(n6242), .Z(n6329) );
  XNOR U8044 ( .A(n6330), .B(n6331), .Z(n6242) );
  ANDN U8045 ( .B(n6332), .A(n6333), .Z(n6330) );
  XOR U8046 ( .A(n6331), .B(n6334), .Z(n6332) );
  XNOR U8047 ( .A(n6327), .B(n6244), .Z(n6328) );
  XOR U8048 ( .A(n6335), .B(n6336), .Z(n6244) );
  AND U8049 ( .A(n26), .B(n6337), .Z(n6335) );
  XOR U8050 ( .A(n6338), .B(n6336), .Z(n6337) );
  XNOR U8051 ( .A(n6339), .B(n6340), .Z(n6327) );
  AND U8052 ( .A(n6341), .B(n6342), .Z(n6339) );
  XNOR U8053 ( .A(n6340), .B(n6269), .Z(n6342) );
  XOR U8054 ( .A(n6333), .B(n6334), .Z(n6269) );
  XNOR U8055 ( .A(n6343), .B(n6344), .Z(n6334) );
  ANDN U8056 ( .B(n6345), .A(n6346), .Z(n6343) );
  XOR U8057 ( .A(n6347), .B(n6348), .Z(n6345) );
  XOR U8058 ( .A(n6349), .B(n6350), .Z(n6333) );
  XNOR U8059 ( .A(n6351), .B(n6352), .Z(n6350) );
  ANDN U8060 ( .B(n6353), .A(n6354), .Z(n6351) );
  XNOR U8061 ( .A(n6355), .B(n6356), .Z(n6353) );
  IV U8062 ( .A(n6331), .Z(n6349) );
  XOR U8063 ( .A(n6357), .B(n6358), .Z(n6331) );
  ANDN U8064 ( .B(n6359), .A(n6360), .Z(n6357) );
  XOR U8065 ( .A(n6358), .B(n6361), .Z(n6359) );
  XOR U8066 ( .A(n6340), .B(n6271), .Z(n6341) );
  XOR U8067 ( .A(n6362), .B(n6363), .Z(n6271) );
  AND U8068 ( .A(n26), .B(n6364), .Z(n6362) );
  XOR U8069 ( .A(n6365), .B(n6363), .Z(n6364) );
  XNOR U8070 ( .A(n6366), .B(n6367), .Z(n6340) );
  NAND U8071 ( .A(n6368), .B(n6369), .Z(n6367) );
  XOR U8072 ( .A(n6370), .B(n6319), .Z(n6369) );
  XOR U8073 ( .A(n6360), .B(n6361), .Z(n6319) );
  XOR U8074 ( .A(n6371), .B(n6348), .Z(n6361) );
  XOR U8075 ( .A(n6372), .B(n6373), .Z(n6348) );
  ANDN U8076 ( .B(n6374), .A(n6375), .Z(n6372) );
  XOR U8077 ( .A(n6373), .B(n6376), .Z(n6374) );
  IV U8078 ( .A(n6346), .Z(n6371) );
  XOR U8079 ( .A(n6344), .B(n6377), .Z(n6346) );
  XOR U8080 ( .A(n6378), .B(n6379), .Z(n6377) );
  ANDN U8081 ( .B(n6380), .A(n6381), .Z(n6378) );
  XOR U8082 ( .A(n6382), .B(n6379), .Z(n6380) );
  IV U8083 ( .A(n6347), .Z(n6344) );
  XOR U8084 ( .A(n6383), .B(n6384), .Z(n6347) );
  ANDN U8085 ( .B(n6385), .A(n6386), .Z(n6383) );
  XOR U8086 ( .A(n6384), .B(n6387), .Z(n6385) );
  XOR U8087 ( .A(n6388), .B(n6389), .Z(n6360) );
  XNOR U8088 ( .A(n6355), .B(n6390), .Z(n6389) );
  IV U8089 ( .A(n6358), .Z(n6390) );
  XOR U8090 ( .A(n6391), .B(n6392), .Z(n6358) );
  ANDN U8091 ( .B(n6393), .A(n6394), .Z(n6391) );
  XOR U8092 ( .A(n6392), .B(n6395), .Z(n6393) );
  XNOR U8093 ( .A(n6396), .B(n6397), .Z(n6355) );
  ANDN U8094 ( .B(n6398), .A(n6399), .Z(n6396) );
  XOR U8095 ( .A(n6397), .B(n6400), .Z(n6398) );
  IV U8096 ( .A(n6354), .Z(n6388) );
  XOR U8097 ( .A(n6352), .B(n6401), .Z(n6354) );
  XOR U8098 ( .A(n6402), .B(n6403), .Z(n6401) );
  ANDN U8099 ( .B(n6404), .A(n6405), .Z(n6402) );
  XOR U8100 ( .A(n6406), .B(n6403), .Z(n6404) );
  IV U8101 ( .A(n6356), .Z(n6352) );
  XOR U8102 ( .A(n6407), .B(n6408), .Z(n6356) );
  ANDN U8103 ( .B(n6409), .A(n6410), .Z(n6407) );
  XOR U8104 ( .A(n6411), .B(n6408), .Z(n6409) );
  IV U8105 ( .A(n6366), .Z(n6370) );
  XOR U8106 ( .A(n6366), .B(n6321), .Z(n6368) );
  XOR U8107 ( .A(n6412), .B(n6413), .Z(n6321) );
  AND U8108 ( .A(n26), .B(n6414), .Z(n6412) );
  XOR U8109 ( .A(n6415), .B(n6413), .Z(n6414) );
  NANDN U8110 ( .A(n6323), .B(n6325), .Z(n6366) );
  XOR U8111 ( .A(n6416), .B(n6417), .Z(n6325) );
  AND U8112 ( .A(n26), .B(n6418), .Z(n6416) );
  XOR U8113 ( .A(n6417), .B(n6419), .Z(n6418) );
  XNOR U8114 ( .A(n6420), .B(n6421), .Z(n26) );
  AND U8115 ( .A(n6422), .B(n6423), .Z(n6420) );
  XOR U8116 ( .A(n6421), .B(n6336), .Z(n6423) );
  XNOR U8117 ( .A(n6424), .B(n6425), .Z(n6336) );
  ANDN U8118 ( .B(n6426), .A(n6427), .Z(n6424) );
  XOR U8119 ( .A(n6425), .B(n6428), .Z(n6426) );
  XNOR U8120 ( .A(n6421), .B(n6338), .Z(n6422) );
  XOR U8121 ( .A(n6429), .B(n6430), .Z(n6338) );
  AND U8122 ( .A(n30), .B(n6431), .Z(n6429) );
  XOR U8123 ( .A(n6432), .B(n6430), .Z(n6431) );
  XNOR U8124 ( .A(n6433), .B(n6434), .Z(n6421) );
  AND U8125 ( .A(n6435), .B(n6436), .Z(n6433) );
  XNOR U8126 ( .A(n6434), .B(n6363), .Z(n6436) );
  XOR U8127 ( .A(n6427), .B(n6428), .Z(n6363) );
  XNOR U8128 ( .A(n6437), .B(n6438), .Z(n6428) );
  ANDN U8129 ( .B(n6439), .A(n6440), .Z(n6437) );
  XOR U8130 ( .A(n6441), .B(n6442), .Z(n6439) );
  XOR U8131 ( .A(n6443), .B(n6444), .Z(n6427) );
  XNOR U8132 ( .A(n6445), .B(n6446), .Z(n6444) );
  ANDN U8133 ( .B(n6447), .A(n6448), .Z(n6445) );
  XNOR U8134 ( .A(n6449), .B(n6450), .Z(n6447) );
  IV U8135 ( .A(n6425), .Z(n6443) );
  XOR U8136 ( .A(n6451), .B(n6452), .Z(n6425) );
  ANDN U8137 ( .B(n6453), .A(n6454), .Z(n6451) );
  XOR U8138 ( .A(n6452), .B(n6455), .Z(n6453) );
  XOR U8139 ( .A(n6434), .B(n6365), .Z(n6435) );
  XOR U8140 ( .A(n6456), .B(n6457), .Z(n6365) );
  AND U8141 ( .A(n30), .B(n6458), .Z(n6456) );
  XOR U8142 ( .A(n6459), .B(n6457), .Z(n6458) );
  XNOR U8143 ( .A(n6460), .B(n6461), .Z(n6434) );
  NAND U8144 ( .A(n6462), .B(n6463), .Z(n6461) );
  XOR U8145 ( .A(n6464), .B(n6413), .Z(n6463) );
  XOR U8146 ( .A(n6454), .B(n6455), .Z(n6413) );
  XOR U8147 ( .A(n6465), .B(n6442), .Z(n6455) );
  XOR U8148 ( .A(n6466), .B(n6467), .Z(n6442) );
  ANDN U8149 ( .B(n6468), .A(n6469), .Z(n6466) );
  XOR U8150 ( .A(n6467), .B(n6470), .Z(n6468) );
  IV U8151 ( .A(n6440), .Z(n6465) );
  XOR U8152 ( .A(n6438), .B(n6471), .Z(n6440) );
  XOR U8153 ( .A(n6472), .B(n6473), .Z(n6471) );
  ANDN U8154 ( .B(n6474), .A(n6475), .Z(n6472) );
  XOR U8155 ( .A(n6476), .B(n6473), .Z(n6474) );
  IV U8156 ( .A(n6441), .Z(n6438) );
  XOR U8157 ( .A(n6477), .B(n6478), .Z(n6441) );
  ANDN U8158 ( .B(n6479), .A(n6480), .Z(n6477) );
  XOR U8159 ( .A(n6478), .B(n6481), .Z(n6479) );
  XOR U8160 ( .A(n6482), .B(n6483), .Z(n6454) );
  XNOR U8161 ( .A(n6449), .B(n6484), .Z(n6483) );
  IV U8162 ( .A(n6452), .Z(n6484) );
  XOR U8163 ( .A(n6485), .B(n6486), .Z(n6452) );
  ANDN U8164 ( .B(n6487), .A(n6488), .Z(n6485) );
  XOR U8165 ( .A(n6486), .B(n6489), .Z(n6487) );
  XNOR U8166 ( .A(n6490), .B(n6491), .Z(n6449) );
  ANDN U8167 ( .B(n6492), .A(n6493), .Z(n6490) );
  XOR U8168 ( .A(n6491), .B(n6494), .Z(n6492) );
  IV U8169 ( .A(n6448), .Z(n6482) );
  XOR U8170 ( .A(n6446), .B(n6495), .Z(n6448) );
  XOR U8171 ( .A(n6496), .B(n6497), .Z(n6495) );
  ANDN U8172 ( .B(n6498), .A(n6499), .Z(n6496) );
  XOR U8173 ( .A(n6500), .B(n6497), .Z(n6498) );
  IV U8174 ( .A(n6450), .Z(n6446) );
  XOR U8175 ( .A(n6501), .B(n6502), .Z(n6450) );
  ANDN U8176 ( .B(n6503), .A(n6504), .Z(n6501) );
  XOR U8177 ( .A(n6505), .B(n6502), .Z(n6503) );
  IV U8178 ( .A(n6460), .Z(n6464) );
  XOR U8179 ( .A(n6460), .B(n6415), .Z(n6462) );
  XOR U8180 ( .A(n6506), .B(n6507), .Z(n6415) );
  AND U8181 ( .A(n30), .B(n6508), .Z(n6506) );
  XOR U8182 ( .A(n6509), .B(n6507), .Z(n6508) );
  NANDN U8183 ( .A(n6417), .B(n6419), .Z(n6460) );
  XOR U8184 ( .A(n6510), .B(n6511), .Z(n6419) );
  AND U8185 ( .A(n30), .B(n6512), .Z(n6510) );
  XOR U8186 ( .A(n6511), .B(n6513), .Z(n6512) );
  XNOR U8187 ( .A(n6514), .B(n6515), .Z(n30) );
  AND U8188 ( .A(n6516), .B(n6517), .Z(n6514) );
  XOR U8189 ( .A(n6515), .B(n6430), .Z(n6517) );
  XNOR U8190 ( .A(n6518), .B(n6519), .Z(n6430) );
  ANDN U8191 ( .B(n6520), .A(n6521), .Z(n6518) );
  XOR U8192 ( .A(n6519), .B(n6522), .Z(n6520) );
  XNOR U8193 ( .A(n6515), .B(n6432), .Z(n6516) );
  XOR U8194 ( .A(n6523), .B(n6524), .Z(n6432) );
  AND U8195 ( .A(n34), .B(n6525), .Z(n6523) );
  XOR U8196 ( .A(n6526), .B(n6524), .Z(n6525) );
  XNOR U8197 ( .A(n6527), .B(n6528), .Z(n6515) );
  AND U8198 ( .A(n6529), .B(n6530), .Z(n6527) );
  XNOR U8199 ( .A(n6528), .B(n6457), .Z(n6530) );
  XOR U8200 ( .A(n6521), .B(n6522), .Z(n6457) );
  XNOR U8201 ( .A(n6531), .B(n6532), .Z(n6522) );
  ANDN U8202 ( .B(n6533), .A(n6534), .Z(n6531) );
  XOR U8203 ( .A(n6535), .B(n6536), .Z(n6533) );
  XOR U8204 ( .A(n6537), .B(n6538), .Z(n6521) );
  XNOR U8205 ( .A(n6539), .B(n6540), .Z(n6538) );
  ANDN U8206 ( .B(n6541), .A(n6542), .Z(n6539) );
  XNOR U8207 ( .A(n6543), .B(n6544), .Z(n6541) );
  IV U8208 ( .A(n6519), .Z(n6537) );
  XOR U8209 ( .A(n6545), .B(n6546), .Z(n6519) );
  ANDN U8210 ( .B(n6547), .A(n6548), .Z(n6545) );
  XOR U8211 ( .A(n6546), .B(n6549), .Z(n6547) );
  XOR U8212 ( .A(n6528), .B(n6459), .Z(n6529) );
  XOR U8213 ( .A(n6550), .B(n6551), .Z(n6459) );
  AND U8214 ( .A(n34), .B(n6552), .Z(n6550) );
  XOR U8215 ( .A(n6553), .B(n6551), .Z(n6552) );
  XNOR U8216 ( .A(n6554), .B(n6555), .Z(n6528) );
  NAND U8217 ( .A(n6556), .B(n6557), .Z(n6555) );
  XOR U8218 ( .A(n6558), .B(n6507), .Z(n6557) );
  XOR U8219 ( .A(n6548), .B(n6549), .Z(n6507) );
  XOR U8220 ( .A(n6559), .B(n6536), .Z(n6549) );
  XOR U8221 ( .A(n6560), .B(n6561), .Z(n6536) );
  ANDN U8222 ( .B(n6562), .A(n6563), .Z(n6560) );
  XOR U8223 ( .A(n6561), .B(n6564), .Z(n6562) );
  IV U8224 ( .A(n6534), .Z(n6559) );
  XOR U8225 ( .A(n6532), .B(n6565), .Z(n6534) );
  XOR U8226 ( .A(n6566), .B(n6567), .Z(n6565) );
  ANDN U8227 ( .B(n6568), .A(n6569), .Z(n6566) );
  XOR U8228 ( .A(n6570), .B(n6567), .Z(n6568) );
  IV U8229 ( .A(n6535), .Z(n6532) );
  XOR U8230 ( .A(n6571), .B(n6572), .Z(n6535) );
  ANDN U8231 ( .B(n6573), .A(n6574), .Z(n6571) );
  XOR U8232 ( .A(n6572), .B(n6575), .Z(n6573) );
  XOR U8233 ( .A(n6576), .B(n6577), .Z(n6548) );
  XNOR U8234 ( .A(n6543), .B(n6578), .Z(n6577) );
  IV U8235 ( .A(n6546), .Z(n6578) );
  XOR U8236 ( .A(n6579), .B(n6580), .Z(n6546) );
  ANDN U8237 ( .B(n6581), .A(n6582), .Z(n6579) );
  XOR U8238 ( .A(n6580), .B(n6583), .Z(n6581) );
  XNOR U8239 ( .A(n6584), .B(n6585), .Z(n6543) );
  ANDN U8240 ( .B(n6586), .A(n6587), .Z(n6584) );
  XOR U8241 ( .A(n6585), .B(n6588), .Z(n6586) );
  IV U8242 ( .A(n6542), .Z(n6576) );
  XOR U8243 ( .A(n6540), .B(n6589), .Z(n6542) );
  XOR U8244 ( .A(n6590), .B(n6591), .Z(n6589) );
  ANDN U8245 ( .B(n6592), .A(n6593), .Z(n6590) );
  XOR U8246 ( .A(n6594), .B(n6591), .Z(n6592) );
  IV U8247 ( .A(n6544), .Z(n6540) );
  XOR U8248 ( .A(n6595), .B(n6596), .Z(n6544) );
  ANDN U8249 ( .B(n6597), .A(n6598), .Z(n6595) );
  XOR U8250 ( .A(n6599), .B(n6596), .Z(n6597) );
  IV U8251 ( .A(n6554), .Z(n6558) );
  XOR U8252 ( .A(n6554), .B(n6509), .Z(n6556) );
  XOR U8253 ( .A(n6600), .B(n6601), .Z(n6509) );
  AND U8254 ( .A(n34), .B(n6602), .Z(n6600) );
  XOR U8255 ( .A(n6603), .B(n6601), .Z(n6602) );
  NANDN U8256 ( .A(n6511), .B(n6513), .Z(n6554) );
  XOR U8257 ( .A(n6604), .B(n6605), .Z(n6513) );
  AND U8258 ( .A(n34), .B(n6606), .Z(n6604) );
  XOR U8259 ( .A(n6605), .B(n6607), .Z(n6606) );
  XNOR U8260 ( .A(n6608), .B(n6609), .Z(n34) );
  AND U8261 ( .A(n6610), .B(n6611), .Z(n6608) );
  XOR U8262 ( .A(n6609), .B(n6524), .Z(n6611) );
  XNOR U8263 ( .A(n6612), .B(n6613), .Z(n6524) );
  ANDN U8264 ( .B(n6614), .A(n6615), .Z(n6612) );
  XOR U8265 ( .A(n6613), .B(n6616), .Z(n6614) );
  XNOR U8266 ( .A(n6609), .B(n6526), .Z(n6610) );
  XOR U8267 ( .A(n6617), .B(n6618), .Z(n6526) );
  AND U8268 ( .A(n38), .B(n6619), .Z(n6617) );
  XOR U8269 ( .A(n6620), .B(n6618), .Z(n6619) );
  XNOR U8270 ( .A(n6621), .B(n6622), .Z(n6609) );
  AND U8271 ( .A(n6623), .B(n6624), .Z(n6621) );
  XNOR U8272 ( .A(n6622), .B(n6551), .Z(n6624) );
  XOR U8273 ( .A(n6615), .B(n6616), .Z(n6551) );
  XNOR U8274 ( .A(n6625), .B(n6626), .Z(n6616) );
  ANDN U8275 ( .B(n6627), .A(n6628), .Z(n6625) );
  XOR U8276 ( .A(n6629), .B(n6630), .Z(n6627) );
  XOR U8277 ( .A(n6631), .B(n6632), .Z(n6615) );
  XNOR U8278 ( .A(n6633), .B(n6634), .Z(n6632) );
  ANDN U8279 ( .B(n6635), .A(n6636), .Z(n6633) );
  XNOR U8280 ( .A(n6637), .B(n6638), .Z(n6635) );
  IV U8281 ( .A(n6613), .Z(n6631) );
  XOR U8282 ( .A(n6639), .B(n6640), .Z(n6613) );
  ANDN U8283 ( .B(n6641), .A(n6642), .Z(n6639) );
  XOR U8284 ( .A(n6640), .B(n6643), .Z(n6641) );
  XOR U8285 ( .A(n6622), .B(n6553), .Z(n6623) );
  XOR U8286 ( .A(n6644), .B(n6645), .Z(n6553) );
  AND U8287 ( .A(n38), .B(n6646), .Z(n6644) );
  XOR U8288 ( .A(n6647), .B(n6645), .Z(n6646) );
  XNOR U8289 ( .A(n6648), .B(n6649), .Z(n6622) );
  NAND U8290 ( .A(n6650), .B(n6651), .Z(n6649) );
  XOR U8291 ( .A(n6652), .B(n6601), .Z(n6651) );
  XOR U8292 ( .A(n6642), .B(n6643), .Z(n6601) );
  XOR U8293 ( .A(n6653), .B(n6630), .Z(n6643) );
  XOR U8294 ( .A(n6654), .B(n6655), .Z(n6630) );
  ANDN U8295 ( .B(n6656), .A(n6657), .Z(n6654) );
  XOR U8296 ( .A(n6655), .B(n6658), .Z(n6656) );
  IV U8297 ( .A(n6628), .Z(n6653) );
  XOR U8298 ( .A(n6626), .B(n6659), .Z(n6628) );
  XOR U8299 ( .A(n6660), .B(n6661), .Z(n6659) );
  ANDN U8300 ( .B(n6662), .A(n6663), .Z(n6660) );
  XOR U8301 ( .A(n6664), .B(n6661), .Z(n6662) );
  IV U8302 ( .A(n6629), .Z(n6626) );
  XOR U8303 ( .A(n6665), .B(n6666), .Z(n6629) );
  ANDN U8304 ( .B(n6667), .A(n6668), .Z(n6665) );
  XOR U8305 ( .A(n6666), .B(n6669), .Z(n6667) );
  XOR U8306 ( .A(n6670), .B(n6671), .Z(n6642) );
  XNOR U8307 ( .A(n6637), .B(n6672), .Z(n6671) );
  IV U8308 ( .A(n6640), .Z(n6672) );
  XOR U8309 ( .A(n6673), .B(n6674), .Z(n6640) );
  ANDN U8310 ( .B(n6675), .A(n6676), .Z(n6673) );
  XOR U8311 ( .A(n6674), .B(n6677), .Z(n6675) );
  XNOR U8312 ( .A(n6678), .B(n6679), .Z(n6637) );
  ANDN U8313 ( .B(n6680), .A(n6681), .Z(n6678) );
  XOR U8314 ( .A(n6679), .B(n6682), .Z(n6680) );
  IV U8315 ( .A(n6636), .Z(n6670) );
  XOR U8316 ( .A(n6634), .B(n6683), .Z(n6636) );
  XOR U8317 ( .A(n6684), .B(n6685), .Z(n6683) );
  ANDN U8318 ( .B(n6686), .A(n6687), .Z(n6684) );
  XOR U8319 ( .A(n6688), .B(n6685), .Z(n6686) );
  IV U8320 ( .A(n6638), .Z(n6634) );
  XOR U8321 ( .A(n6689), .B(n6690), .Z(n6638) );
  ANDN U8322 ( .B(n6691), .A(n6692), .Z(n6689) );
  XOR U8323 ( .A(n6693), .B(n6690), .Z(n6691) );
  IV U8324 ( .A(n6648), .Z(n6652) );
  XOR U8325 ( .A(n6648), .B(n6603), .Z(n6650) );
  XOR U8326 ( .A(n6694), .B(n6695), .Z(n6603) );
  AND U8327 ( .A(n38), .B(n6696), .Z(n6694) );
  XOR U8328 ( .A(n6697), .B(n6695), .Z(n6696) );
  NANDN U8329 ( .A(n6605), .B(n6607), .Z(n6648) );
  XOR U8330 ( .A(n6698), .B(n6699), .Z(n6607) );
  AND U8331 ( .A(n38), .B(n6700), .Z(n6698) );
  XOR U8332 ( .A(n6699), .B(n6701), .Z(n6700) );
  XNOR U8333 ( .A(n6702), .B(n6703), .Z(n38) );
  AND U8334 ( .A(n6704), .B(n6705), .Z(n6702) );
  XOR U8335 ( .A(n6703), .B(n6618), .Z(n6705) );
  XNOR U8336 ( .A(n6706), .B(n6707), .Z(n6618) );
  ANDN U8337 ( .B(n6708), .A(n6709), .Z(n6706) );
  XOR U8338 ( .A(n6707), .B(n6710), .Z(n6708) );
  XNOR U8339 ( .A(n6703), .B(n6620), .Z(n6704) );
  XOR U8340 ( .A(n6711), .B(n6712), .Z(n6620) );
  AND U8341 ( .A(n42), .B(n6713), .Z(n6711) );
  XOR U8342 ( .A(n6714), .B(n6712), .Z(n6713) );
  XNOR U8343 ( .A(n6715), .B(n6716), .Z(n6703) );
  AND U8344 ( .A(n6717), .B(n6718), .Z(n6715) );
  XNOR U8345 ( .A(n6716), .B(n6645), .Z(n6718) );
  XOR U8346 ( .A(n6709), .B(n6710), .Z(n6645) );
  XNOR U8347 ( .A(n6719), .B(n6720), .Z(n6710) );
  ANDN U8348 ( .B(n6721), .A(n6722), .Z(n6719) );
  XOR U8349 ( .A(n6723), .B(n6724), .Z(n6721) );
  XOR U8350 ( .A(n6725), .B(n6726), .Z(n6709) );
  XNOR U8351 ( .A(n6727), .B(n6728), .Z(n6726) );
  ANDN U8352 ( .B(n6729), .A(n6730), .Z(n6727) );
  XNOR U8353 ( .A(n6731), .B(n6732), .Z(n6729) );
  IV U8354 ( .A(n6707), .Z(n6725) );
  XOR U8355 ( .A(n6733), .B(n6734), .Z(n6707) );
  ANDN U8356 ( .B(n6735), .A(n6736), .Z(n6733) );
  XOR U8357 ( .A(n6734), .B(n6737), .Z(n6735) );
  XOR U8358 ( .A(n6716), .B(n6647), .Z(n6717) );
  XOR U8359 ( .A(n6738), .B(n6739), .Z(n6647) );
  AND U8360 ( .A(n42), .B(n6740), .Z(n6738) );
  XOR U8361 ( .A(n6741), .B(n6739), .Z(n6740) );
  XNOR U8362 ( .A(n6742), .B(n6743), .Z(n6716) );
  NAND U8363 ( .A(n6744), .B(n6745), .Z(n6743) );
  XOR U8364 ( .A(n6746), .B(n6695), .Z(n6745) );
  XOR U8365 ( .A(n6736), .B(n6737), .Z(n6695) );
  XOR U8366 ( .A(n6747), .B(n6724), .Z(n6737) );
  XOR U8367 ( .A(n6748), .B(n6749), .Z(n6724) );
  ANDN U8368 ( .B(n6750), .A(n6751), .Z(n6748) );
  XOR U8369 ( .A(n6749), .B(n6752), .Z(n6750) );
  IV U8370 ( .A(n6722), .Z(n6747) );
  XOR U8371 ( .A(n6720), .B(n6753), .Z(n6722) );
  XOR U8372 ( .A(n6754), .B(n6755), .Z(n6753) );
  ANDN U8373 ( .B(n6756), .A(n6757), .Z(n6754) );
  XOR U8374 ( .A(n6758), .B(n6755), .Z(n6756) );
  IV U8375 ( .A(n6723), .Z(n6720) );
  XOR U8376 ( .A(n6759), .B(n6760), .Z(n6723) );
  ANDN U8377 ( .B(n6761), .A(n6762), .Z(n6759) );
  XOR U8378 ( .A(n6760), .B(n6763), .Z(n6761) );
  XOR U8379 ( .A(n6764), .B(n6765), .Z(n6736) );
  XNOR U8380 ( .A(n6731), .B(n6766), .Z(n6765) );
  IV U8381 ( .A(n6734), .Z(n6766) );
  XOR U8382 ( .A(n6767), .B(n6768), .Z(n6734) );
  ANDN U8383 ( .B(n6769), .A(n6770), .Z(n6767) );
  XOR U8384 ( .A(n6768), .B(n6771), .Z(n6769) );
  XNOR U8385 ( .A(n6772), .B(n6773), .Z(n6731) );
  ANDN U8386 ( .B(n6774), .A(n6775), .Z(n6772) );
  XOR U8387 ( .A(n6773), .B(n6776), .Z(n6774) );
  IV U8388 ( .A(n6730), .Z(n6764) );
  XOR U8389 ( .A(n6728), .B(n6777), .Z(n6730) );
  XOR U8390 ( .A(n6778), .B(n6779), .Z(n6777) );
  ANDN U8391 ( .B(n6780), .A(n6781), .Z(n6778) );
  XOR U8392 ( .A(n6782), .B(n6779), .Z(n6780) );
  IV U8393 ( .A(n6732), .Z(n6728) );
  XOR U8394 ( .A(n6783), .B(n6784), .Z(n6732) );
  ANDN U8395 ( .B(n6785), .A(n6786), .Z(n6783) );
  XOR U8396 ( .A(n6787), .B(n6784), .Z(n6785) );
  IV U8397 ( .A(n6742), .Z(n6746) );
  XOR U8398 ( .A(n6742), .B(n6697), .Z(n6744) );
  XOR U8399 ( .A(n6788), .B(n6789), .Z(n6697) );
  AND U8400 ( .A(n42), .B(n6790), .Z(n6788) );
  XOR U8401 ( .A(n6791), .B(n6789), .Z(n6790) );
  NANDN U8402 ( .A(n6699), .B(n6701), .Z(n6742) );
  XOR U8403 ( .A(n6792), .B(n6793), .Z(n6701) );
  AND U8404 ( .A(n42), .B(n6794), .Z(n6792) );
  XOR U8405 ( .A(n6793), .B(n6795), .Z(n6794) );
  XNOR U8406 ( .A(n6796), .B(n6797), .Z(n42) );
  AND U8407 ( .A(n6798), .B(n6799), .Z(n6796) );
  XOR U8408 ( .A(n6797), .B(n6712), .Z(n6799) );
  XNOR U8409 ( .A(n6800), .B(n6801), .Z(n6712) );
  ANDN U8410 ( .B(n6802), .A(n6803), .Z(n6800) );
  XOR U8411 ( .A(n6801), .B(n6804), .Z(n6802) );
  XNOR U8412 ( .A(n6797), .B(n6714), .Z(n6798) );
  XOR U8413 ( .A(n6805), .B(n6806), .Z(n6714) );
  AND U8414 ( .A(n46), .B(n6807), .Z(n6805) );
  XOR U8415 ( .A(n6808), .B(n6806), .Z(n6807) );
  XNOR U8416 ( .A(n6809), .B(n6810), .Z(n6797) );
  AND U8417 ( .A(n6811), .B(n6812), .Z(n6809) );
  XNOR U8418 ( .A(n6810), .B(n6739), .Z(n6812) );
  XOR U8419 ( .A(n6803), .B(n6804), .Z(n6739) );
  XNOR U8420 ( .A(n6813), .B(n6814), .Z(n6804) );
  ANDN U8421 ( .B(n6815), .A(n6816), .Z(n6813) );
  XOR U8422 ( .A(n6817), .B(n6818), .Z(n6815) );
  XOR U8423 ( .A(n6819), .B(n6820), .Z(n6803) );
  XNOR U8424 ( .A(n6821), .B(n6822), .Z(n6820) );
  ANDN U8425 ( .B(n6823), .A(n6824), .Z(n6821) );
  XNOR U8426 ( .A(n6825), .B(n6826), .Z(n6823) );
  IV U8427 ( .A(n6801), .Z(n6819) );
  XOR U8428 ( .A(n6827), .B(n6828), .Z(n6801) );
  ANDN U8429 ( .B(n6829), .A(n6830), .Z(n6827) );
  XOR U8430 ( .A(n6828), .B(n6831), .Z(n6829) );
  XOR U8431 ( .A(n6810), .B(n6741), .Z(n6811) );
  XOR U8432 ( .A(n6832), .B(n6833), .Z(n6741) );
  AND U8433 ( .A(n46), .B(n6834), .Z(n6832) );
  XOR U8434 ( .A(n6835), .B(n6833), .Z(n6834) );
  XNOR U8435 ( .A(n6836), .B(n6837), .Z(n6810) );
  NAND U8436 ( .A(n6838), .B(n6839), .Z(n6837) );
  XOR U8437 ( .A(n6840), .B(n6789), .Z(n6839) );
  XOR U8438 ( .A(n6830), .B(n6831), .Z(n6789) );
  XOR U8439 ( .A(n6841), .B(n6818), .Z(n6831) );
  XOR U8440 ( .A(n6842), .B(n6843), .Z(n6818) );
  ANDN U8441 ( .B(n6844), .A(n6845), .Z(n6842) );
  XOR U8442 ( .A(n6843), .B(n6846), .Z(n6844) );
  IV U8443 ( .A(n6816), .Z(n6841) );
  XOR U8444 ( .A(n6814), .B(n6847), .Z(n6816) );
  XOR U8445 ( .A(n6848), .B(n6849), .Z(n6847) );
  ANDN U8446 ( .B(n6850), .A(n6851), .Z(n6848) );
  XOR U8447 ( .A(n6852), .B(n6849), .Z(n6850) );
  IV U8448 ( .A(n6817), .Z(n6814) );
  XOR U8449 ( .A(n6853), .B(n6854), .Z(n6817) );
  ANDN U8450 ( .B(n6855), .A(n6856), .Z(n6853) );
  XOR U8451 ( .A(n6854), .B(n6857), .Z(n6855) );
  XOR U8452 ( .A(n6858), .B(n6859), .Z(n6830) );
  XNOR U8453 ( .A(n6825), .B(n6860), .Z(n6859) );
  IV U8454 ( .A(n6828), .Z(n6860) );
  XOR U8455 ( .A(n6861), .B(n6862), .Z(n6828) );
  ANDN U8456 ( .B(n6863), .A(n6864), .Z(n6861) );
  XOR U8457 ( .A(n6862), .B(n6865), .Z(n6863) );
  XNOR U8458 ( .A(n6866), .B(n6867), .Z(n6825) );
  ANDN U8459 ( .B(n6868), .A(n6869), .Z(n6866) );
  XOR U8460 ( .A(n6867), .B(n6870), .Z(n6868) );
  IV U8461 ( .A(n6824), .Z(n6858) );
  XOR U8462 ( .A(n6822), .B(n6871), .Z(n6824) );
  XOR U8463 ( .A(n6872), .B(n6873), .Z(n6871) );
  ANDN U8464 ( .B(n6874), .A(n6875), .Z(n6872) );
  XOR U8465 ( .A(n6876), .B(n6873), .Z(n6874) );
  IV U8466 ( .A(n6826), .Z(n6822) );
  XOR U8467 ( .A(n6877), .B(n6878), .Z(n6826) );
  ANDN U8468 ( .B(n6879), .A(n6880), .Z(n6877) );
  XOR U8469 ( .A(n6881), .B(n6878), .Z(n6879) );
  IV U8470 ( .A(n6836), .Z(n6840) );
  XOR U8471 ( .A(n6836), .B(n6791), .Z(n6838) );
  XOR U8472 ( .A(n6882), .B(n6883), .Z(n6791) );
  AND U8473 ( .A(n46), .B(n6884), .Z(n6882) );
  XOR U8474 ( .A(n6885), .B(n6883), .Z(n6884) );
  NANDN U8475 ( .A(n6793), .B(n6795), .Z(n6836) );
  XOR U8476 ( .A(n6886), .B(n6887), .Z(n6795) );
  AND U8477 ( .A(n46), .B(n6888), .Z(n6886) );
  XOR U8478 ( .A(n6887), .B(n6889), .Z(n6888) );
  XNOR U8479 ( .A(n6890), .B(n6891), .Z(n46) );
  AND U8480 ( .A(n6892), .B(n6893), .Z(n6890) );
  XOR U8481 ( .A(n6891), .B(n6806), .Z(n6893) );
  XNOR U8482 ( .A(n6894), .B(n6895), .Z(n6806) );
  ANDN U8483 ( .B(n6896), .A(n6897), .Z(n6894) );
  XOR U8484 ( .A(n6895), .B(n6898), .Z(n6896) );
  XNOR U8485 ( .A(n6891), .B(n6808), .Z(n6892) );
  XOR U8486 ( .A(n6899), .B(n6900), .Z(n6808) );
  AND U8487 ( .A(n50), .B(n6901), .Z(n6899) );
  XOR U8488 ( .A(n6902), .B(n6900), .Z(n6901) );
  XNOR U8489 ( .A(n6903), .B(n6904), .Z(n6891) );
  AND U8490 ( .A(n6905), .B(n6906), .Z(n6903) );
  XNOR U8491 ( .A(n6904), .B(n6833), .Z(n6906) );
  XOR U8492 ( .A(n6897), .B(n6898), .Z(n6833) );
  XNOR U8493 ( .A(n6907), .B(n6908), .Z(n6898) );
  ANDN U8494 ( .B(n6909), .A(n6910), .Z(n6907) );
  XOR U8495 ( .A(n6911), .B(n6912), .Z(n6909) );
  XOR U8496 ( .A(n6913), .B(n6914), .Z(n6897) );
  XNOR U8497 ( .A(n6915), .B(n6916), .Z(n6914) );
  ANDN U8498 ( .B(n6917), .A(n6918), .Z(n6915) );
  XNOR U8499 ( .A(n6919), .B(n6920), .Z(n6917) );
  IV U8500 ( .A(n6895), .Z(n6913) );
  XOR U8501 ( .A(n6921), .B(n6922), .Z(n6895) );
  ANDN U8502 ( .B(n6923), .A(n6924), .Z(n6921) );
  XOR U8503 ( .A(n6922), .B(n6925), .Z(n6923) );
  XOR U8504 ( .A(n6904), .B(n6835), .Z(n6905) );
  XOR U8505 ( .A(n6926), .B(n6927), .Z(n6835) );
  AND U8506 ( .A(n50), .B(n6928), .Z(n6926) );
  XOR U8507 ( .A(n6929), .B(n6927), .Z(n6928) );
  XNOR U8508 ( .A(n6930), .B(n6931), .Z(n6904) );
  NAND U8509 ( .A(n6932), .B(n6933), .Z(n6931) );
  XOR U8510 ( .A(n6934), .B(n6883), .Z(n6933) );
  XOR U8511 ( .A(n6924), .B(n6925), .Z(n6883) );
  XOR U8512 ( .A(n6935), .B(n6912), .Z(n6925) );
  XOR U8513 ( .A(n6936), .B(n6937), .Z(n6912) );
  ANDN U8514 ( .B(n6938), .A(n6939), .Z(n6936) );
  XOR U8515 ( .A(n6937), .B(n6940), .Z(n6938) );
  IV U8516 ( .A(n6910), .Z(n6935) );
  XOR U8517 ( .A(n6908), .B(n6941), .Z(n6910) );
  XOR U8518 ( .A(n6942), .B(n6943), .Z(n6941) );
  ANDN U8519 ( .B(n6944), .A(n6945), .Z(n6942) );
  XOR U8520 ( .A(n6946), .B(n6943), .Z(n6944) );
  IV U8521 ( .A(n6911), .Z(n6908) );
  XOR U8522 ( .A(n6947), .B(n6948), .Z(n6911) );
  ANDN U8523 ( .B(n6949), .A(n6950), .Z(n6947) );
  XOR U8524 ( .A(n6948), .B(n6951), .Z(n6949) );
  XOR U8525 ( .A(n6952), .B(n6953), .Z(n6924) );
  XNOR U8526 ( .A(n6919), .B(n6954), .Z(n6953) );
  IV U8527 ( .A(n6922), .Z(n6954) );
  XOR U8528 ( .A(n6955), .B(n6956), .Z(n6922) );
  ANDN U8529 ( .B(n6957), .A(n6958), .Z(n6955) );
  XOR U8530 ( .A(n6956), .B(n6959), .Z(n6957) );
  XNOR U8531 ( .A(n6960), .B(n6961), .Z(n6919) );
  ANDN U8532 ( .B(n6962), .A(n6963), .Z(n6960) );
  XOR U8533 ( .A(n6961), .B(n6964), .Z(n6962) );
  IV U8534 ( .A(n6918), .Z(n6952) );
  XOR U8535 ( .A(n6916), .B(n6965), .Z(n6918) );
  XOR U8536 ( .A(n6966), .B(n6967), .Z(n6965) );
  ANDN U8537 ( .B(n6968), .A(n6969), .Z(n6966) );
  XOR U8538 ( .A(n6970), .B(n6967), .Z(n6968) );
  IV U8539 ( .A(n6920), .Z(n6916) );
  XOR U8540 ( .A(n6971), .B(n6972), .Z(n6920) );
  ANDN U8541 ( .B(n6973), .A(n6974), .Z(n6971) );
  XOR U8542 ( .A(n6975), .B(n6972), .Z(n6973) );
  IV U8543 ( .A(n6930), .Z(n6934) );
  XOR U8544 ( .A(n6930), .B(n6885), .Z(n6932) );
  XOR U8545 ( .A(n6976), .B(n6977), .Z(n6885) );
  AND U8546 ( .A(n50), .B(n6978), .Z(n6976) );
  XOR U8547 ( .A(n6979), .B(n6977), .Z(n6978) );
  NANDN U8548 ( .A(n6887), .B(n6889), .Z(n6930) );
  XOR U8549 ( .A(n6980), .B(n6981), .Z(n6889) );
  AND U8550 ( .A(n50), .B(n6982), .Z(n6980) );
  XOR U8551 ( .A(n6981), .B(n6983), .Z(n6982) );
  XNOR U8552 ( .A(n6984), .B(n6985), .Z(n50) );
  AND U8553 ( .A(n6986), .B(n6987), .Z(n6984) );
  XOR U8554 ( .A(n6985), .B(n6900), .Z(n6987) );
  XNOR U8555 ( .A(n6988), .B(n6989), .Z(n6900) );
  ANDN U8556 ( .B(n6990), .A(n6991), .Z(n6988) );
  XOR U8557 ( .A(n6989), .B(n6992), .Z(n6990) );
  XNOR U8558 ( .A(n6985), .B(n6902), .Z(n6986) );
  XOR U8559 ( .A(n6993), .B(n6994), .Z(n6902) );
  AND U8560 ( .A(n54), .B(n6995), .Z(n6993) );
  XOR U8561 ( .A(n6996), .B(n6994), .Z(n6995) );
  XNOR U8562 ( .A(n6997), .B(n6998), .Z(n6985) );
  AND U8563 ( .A(n6999), .B(n7000), .Z(n6997) );
  XNOR U8564 ( .A(n6998), .B(n6927), .Z(n7000) );
  XOR U8565 ( .A(n6991), .B(n6992), .Z(n6927) );
  XNOR U8566 ( .A(n7001), .B(n7002), .Z(n6992) );
  ANDN U8567 ( .B(n7003), .A(n7004), .Z(n7001) );
  XOR U8568 ( .A(n7005), .B(n7006), .Z(n7003) );
  XOR U8569 ( .A(n7007), .B(n7008), .Z(n6991) );
  XNOR U8570 ( .A(n7009), .B(n7010), .Z(n7008) );
  ANDN U8571 ( .B(n7011), .A(n7012), .Z(n7009) );
  XNOR U8572 ( .A(n7013), .B(n7014), .Z(n7011) );
  IV U8573 ( .A(n6989), .Z(n7007) );
  XOR U8574 ( .A(n7015), .B(n7016), .Z(n6989) );
  ANDN U8575 ( .B(n7017), .A(n7018), .Z(n7015) );
  XOR U8576 ( .A(n7016), .B(n7019), .Z(n7017) );
  XOR U8577 ( .A(n6998), .B(n6929), .Z(n6999) );
  XOR U8578 ( .A(n7020), .B(n7021), .Z(n6929) );
  AND U8579 ( .A(n54), .B(n7022), .Z(n7020) );
  XOR U8580 ( .A(n7023), .B(n7021), .Z(n7022) );
  XNOR U8581 ( .A(n7024), .B(n7025), .Z(n6998) );
  NAND U8582 ( .A(n7026), .B(n7027), .Z(n7025) );
  XOR U8583 ( .A(n7028), .B(n6977), .Z(n7027) );
  XOR U8584 ( .A(n7018), .B(n7019), .Z(n6977) );
  XOR U8585 ( .A(n7029), .B(n7006), .Z(n7019) );
  XOR U8586 ( .A(n7030), .B(n7031), .Z(n7006) );
  ANDN U8587 ( .B(n7032), .A(n7033), .Z(n7030) );
  XOR U8588 ( .A(n7031), .B(n7034), .Z(n7032) );
  IV U8589 ( .A(n7004), .Z(n7029) );
  XOR U8590 ( .A(n7002), .B(n7035), .Z(n7004) );
  XOR U8591 ( .A(n7036), .B(n7037), .Z(n7035) );
  ANDN U8592 ( .B(n7038), .A(n7039), .Z(n7036) );
  XOR U8593 ( .A(n7040), .B(n7037), .Z(n7038) );
  IV U8594 ( .A(n7005), .Z(n7002) );
  XOR U8595 ( .A(n7041), .B(n7042), .Z(n7005) );
  ANDN U8596 ( .B(n7043), .A(n7044), .Z(n7041) );
  XOR U8597 ( .A(n7042), .B(n7045), .Z(n7043) );
  XOR U8598 ( .A(n7046), .B(n7047), .Z(n7018) );
  XNOR U8599 ( .A(n7013), .B(n7048), .Z(n7047) );
  IV U8600 ( .A(n7016), .Z(n7048) );
  XOR U8601 ( .A(n7049), .B(n7050), .Z(n7016) );
  ANDN U8602 ( .B(n7051), .A(n7052), .Z(n7049) );
  XOR U8603 ( .A(n7050), .B(n7053), .Z(n7051) );
  XNOR U8604 ( .A(n7054), .B(n7055), .Z(n7013) );
  ANDN U8605 ( .B(n7056), .A(n7057), .Z(n7054) );
  XOR U8606 ( .A(n7055), .B(n7058), .Z(n7056) );
  IV U8607 ( .A(n7012), .Z(n7046) );
  XOR U8608 ( .A(n7010), .B(n7059), .Z(n7012) );
  XOR U8609 ( .A(n7060), .B(n7061), .Z(n7059) );
  ANDN U8610 ( .B(n7062), .A(n7063), .Z(n7060) );
  XOR U8611 ( .A(n7064), .B(n7061), .Z(n7062) );
  IV U8612 ( .A(n7014), .Z(n7010) );
  XOR U8613 ( .A(n7065), .B(n7066), .Z(n7014) );
  ANDN U8614 ( .B(n7067), .A(n7068), .Z(n7065) );
  XOR U8615 ( .A(n7069), .B(n7066), .Z(n7067) );
  IV U8616 ( .A(n7024), .Z(n7028) );
  XOR U8617 ( .A(n7024), .B(n6979), .Z(n7026) );
  XOR U8618 ( .A(n7070), .B(n7071), .Z(n6979) );
  AND U8619 ( .A(n54), .B(n7072), .Z(n7070) );
  XOR U8620 ( .A(n7073), .B(n7071), .Z(n7072) );
  NANDN U8621 ( .A(n6981), .B(n6983), .Z(n7024) );
  XOR U8622 ( .A(n7074), .B(n7075), .Z(n6983) );
  AND U8623 ( .A(n54), .B(n7076), .Z(n7074) );
  XOR U8624 ( .A(n7075), .B(n7077), .Z(n7076) );
  XNOR U8625 ( .A(n7078), .B(n7079), .Z(n54) );
  AND U8626 ( .A(n7080), .B(n7081), .Z(n7078) );
  XOR U8627 ( .A(n7079), .B(n6994), .Z(n7081) );
  XNOR U8628 ( .A(n7082), .B(n7083), .Z(n6994) );
  ANDN U8629 ( .B(n7084), .A(n7085), .Z(n7082) );
  XOR U8630 ( .A(n7083), .B(n7086), .Z(n7084) );
  XNOR U8631 ( .A(n7079), .B(n6996), .Z(n7080) );
  XOR U8632 ( .A(n7087), .B(n7088), .Z(n6996) );
  AND U8633 ( .A(n58), .B(n7089), .Z(n7087) );
  XOR U8634 ( .A(n7090), .B(n7088), .Z(n7089) );
  XNOR U8635 ( .A(n7091), .B(n7092), .Z(n7079) );
  AND U8636 ( .A(n7093), .B(n7094), .Z(n7091) );
  XNOR U8637 ( .A(n7092), .B(n7021), .Z(n7094) );
  XOR U8638 ( .A(n7085), .B(n7086), .Z(n7021) );
  XNOR U8639 ( .A(n7095), .B(n7096), .Z(n7086) );
  ANDN U8640 ( .B(n7097), .A(n7098), .Z(n7095) );
  XOR U8641 ( .A(n7099), .B(n7100), .Z(n7097) );
  XOR U8642 ( .A(n7101), .B(n7102), .Z(n7085) );
  XNOR U8643 ( .A(n7103), .B(n7104), .Z(n7102) );
  ANDN U8644 ( .B(n7105), .A(n7106), .Z(n7103) );
  XNOR U8645 ( .A(n7107), .B(n7108), .Z(n7105) );
  IV U8646 ( .A(n7083), .Z(n7101) );
  XOR U8647 ( .A(n7109), .B(n7110), .Z(n7083) );
  ANDN U8648 ( .B(n7111), .A(n7112), .Z(n7109) );
  XOR U8649 ( .A(n7110), .B(n7113), .Z(n7111) );
  XOR U8650 ( .A(n7092), .B(n7023), .Z(n7093) );
  XOR U8651 ( .A(n7114), .B(n7115), .Z(n7023) );
  AND U8652 ( .A(n58), .B(n7116), .Z(n7114) );
  XOR U8653 ( .A(n7117), .B(n7115), .Z(n7116) );
  XNOR U8654 ( .A(n7118), .B(n7119), .Z(n7092) );
  NAND U8655 ( .A(n7120), .B(n7121), .Z(n7119) );
  XOR U8656 ( .A(n7122), .B(n7071), .Z(n7121) );
  XOR U8657 ( .A(n7112), .B(n7113), .Z(n7071) );
  XOR U8658 ( .A(n7123), .B(n7100), .Z(n7113) );
  XOR U8659 ( .A(n7124), .B(n7125), .Z(n7100) );
  ANDN U8660 ( .B(n7126), .A(n7127), .Z(n7124) );
  XOR U8661 ( .A(n7125), .B(n7128), .Z(n7126) );
  IV U8662 ( .A(n7098), .Z(n7123) );
  XOR U8663 ( .A(n7096), .B(n7129), .Z(n7098) );
  XOR U8664 ( .A(n7130), .B(n7131), .Z(n7129) );
  ANDN U8665 ( .B(n7132), .A(n7133), .Z(n7130) );
  XOR U8666 ( .A(n7134), .B(n7131), .Z(n7132) );
  IV U8667 ( .A(n7099), .Z(n7096) );
  XOR U8668 ( .A(n7135), .B(n7136), .Z(n7099) );
  ANDN U8669 ( .B(n7137), .A(n7138), .Z(n7135) );
  XOR U8670 ( .A(n7136), .B(n7139), .Z(n7137) );
  XOR U8671 ( .A(n7140), .B(n7141), .Z(n7112) );
  XNOR U8672 ( .A(n7107), .B(n7142), .Z(n7141) );
  IV U8673 ( .A(n7110), .Z(n7142) );
  XOR U8674 ( .A(n7143), .B(n7144), .Z(n7110) );
  ANDN U8675 ( .B(n7145), .A(n7146), .Z(n7143) );
  XOR U8676 ( .A(n7144), .B(n7147), .Z(n7145) );
  XNOR U8677 ( .A(n7148), .B(n7149), .Z(n7107) );
  ANDN U8678 ( .B(n7150), .A(n7151), .Z(n7148) );
  XOR U8679 ( .A(n7149), .B(n7152), .Z(n7150) );
  IV U8680 ( .A(n7106), .Z(n7140) );
  XOR U8681 ( .A(n7104), .B(n7153), .Z(n7106) );
  XOR U8682 ( .A(n7154), .B(n7155), .Z(n7153) );
  ANDN U8683 ( .B(n7156), .A(n7157), .Z(n7154) );
  XOR U8684 ( .A(n7158), .B(n7155), .Z(n7156) );
  IV U8685 ( .A(n7108), .Z(n7104) );
  XOR U8686 ( .A(n7159), .B(n7160), .Z(n7108) );
  ANDN U8687 ( .B(n7161), .A(n7162), .Z(n7159) );
  XOR U8688 ( .A(n7163), .B(n7160), .Z(n7161) );
  IV U8689 ( .A(n7118), .Z(n7122) );
  XOR U8690 ( .A(n7118), .B(n7073), .Z(n7120) );
  XOR U8691 ( .A(n7164), .B(n7165), .Z(n7073) );
  AND U8692 ( .A(n58), .B(n7166), .Z(n7164) );
  XOR U8693 ( .A(n7167), .B(n7165), .Z(n7166) );
  NANDN U8694 ( .A(n7075), .B(n7077), .Z(n7118) );
  XOR U8695 ( .A(n7168), .B(n7169), .Z(n7077) );
  AND U8696 ( .A(n58), .B(n7170), .Z(n7168) );
  XOR U8697 ( .A(n7169), .B(n7171), .Z(n7170) );
  XNOR U8698 ( .A(n7172), .B(n7173), .Z(n58) );
  AND U8699 ( .A(n7174), .B(n7175), .Z(n7172) );
  XOR U8700 ( .A(n7173), .B(n7088), .Z(n7175) );
  XNOR U8701 ( .A(n7176), .B(n7177), .Z(n7088) );
  ANDN U8702 ( .B(n7178), .A(n7179), .Z(n7176) );
  XOR U8703 ( .A(n7177), .B(n7180), .Z(n7178) );
  XNOR U8704 ( .A(n7173), .B(n7090), .Z(n7174) );
  XOR U8705 ( .A(n7181), .B(n7182), .Z(n7090) );
  AND U8706 ( .A(n62), .B(n7183), .Z(n7181) );
  XOR U8707 ( .A(n7184), .B(n7182), .Z(n7183) );
  XNOR U8708 ( .A(n7185), .B(n7186), .Z(n7173) );
  AND U8709 ( .A(n7187), .B(n7188), .Z(n7185) );
  XNOR U8710 ( .A(n7186), .B(n7115), .Z(n7188) );
  XOR U8711 ( .A(n7179), .B(n7180), .Z(n7115) );
  XNOR U8712 ( .A(n7189), .B(n7190), .Z(n7180) );
  ANDN U8713 ( .B(n7191), .A(n7192), .Z(n7189) );
  XOR U8714 ( .A(n7193), .B(n7194), .Z(n7191) );
  XOR U8715 ( .A(n7195), .B(n7196), .Z(n7179) );
  XNOR U8716 ( .A(n7197), .B(n7198), .Z(n7196) );
  ANDN U8717 ( .B(n7199), .A(n7200), .Z(n7197) );
  XNOR U8718 ( .A(n7201), .B(n7202), .Z(n7199) );
  IV U8719 ( .A(n7177), .Z(n7195) );
  XOR U8720 ( .A(n7203), .B(n7204), .Z(n7177) );
  ANDN U8721 ( .B(n7205), .A(n7206), .Z(n7203) );
  XOR U8722 ( .A(n7204), .B(n7207), .Z(n7205) );
  XOR U8723 ( .A(n7186), .B(n7117), .Z(n7187) );
  XOR U8724 ( .A(n7208), .B(n7209), .Z(n7117) );
  AND U8725 ( .A(n62), .B(n7210), .Z(n7208) );
  XOR U8726 ( .A(n7211), .B(n7209), .Z(n7210) );
  XNOR U8727 ( .A(n7212), .B(n7213), .Z(n7186) );
  NAND U8728 ( .A(n7214), .B(n7215), .Z(n7213) );
  XOR U8729 ( .A(n7216), .B(n7165), .Z(n7215) );
  XOR U8730 ( .A(n7206), .B(n7207), .Z(n7165) );
  XOR U8731 ( .A(n7217), .B(n7194), .Z(n7207) );
  XOR U8732 ( .A(n7218), .B(n7219), .Z(n7194) );
  ANDN U8733 ( .B(n7220), .A(n7221), .Z(n7218) );
  XOR U8734 ( .A(n7219), .B(n7222), .Z(n7220) );
  IV U8735 ( .A(n7192), .Z(n7217) );
  XOR U8736 ( .A(n7190), .B(n7223), .Z(n7192) );
  XOR U8737 ( .A(n7224), .B(n7225), .Z(n7223) );
  ANDN U8738 ( .B(n7226), .A(n7227), .Z(n7224) );
  XOR U8739 ( .A(n7228), .B(n7225), .Z(n7226) );
  IV U8740 ( .A(n7193), .Z(n7190) );
  XOR U8741 ( .A(n7229), .B(n7230), .Z(n7193) );
  ANDN U8742 ( .B(n7231), .A(n7232), .Z(n7229) );
  XOR U8743 ( .A(n7230), .B(n7233), .Z(n7231) );
  XOR U8744 ( .A(n7234), .B(n7235), .Z(n7206) );
  XNOR U8745 ( .A(n7201), .B(n7236), .Z(n7235) );
  IV U8746 ( .A(n7204), .Z(n7236) );
  XOR U8747 ( .A(n7237), .B(n7238), .Z(n7204) );
  ANDN U8748 ( .B(n7239), .A(n7240), .Z(n7237) );
  XOR U8749 ( .A(n7238), .B(n7241), .Z(n7239) );
  XNOR U8750 ( .A(n7242), .B(n7243), .Z(n7201) );
  ANDN U8751 ( .B(n7244), .A(n7245), .Z(n7242) );
  XOR U8752 ( .A(n7243), .B(n7246), .Z(n7244) );
  IV U8753 ( .A(n7200), .Z(n7234) );
  XOR U8754 ( .A(n7198), .B(n7247), .Z(n7200) );
  XOR U8755 ( .A(n7248), .B(n7249), .Z(n7247) );
  ANDN U8756 ( .B(n7250), .A(n7251), .Z(n7248) );
  XOR U8757 ( .A(n7252), .B(n7249), .Z(n7250) );
  IV U8758 ( .A(n7202), .Z(n7198) );
  XOR U8759 ( .A(n7253), .B(n7254), .Z(n7202) );
  ANDN U8760 ( .B(n7255), .A(n7256), .Z(n7253) );
  XOR U8761 ( .A(n7257), .B(n7254), .Z(n7255) );
  IV U8762 ( .A(n7212), .Z(n7216) );
  XOR U8763 ( .A(n7212), .B(n7167), .Z(n7214) );
  XOR U8764 ( .A(n7258), .B(n7259), .Z(n7167) );
  AND U8765 ( .A(n62), .B(n7260), .Z(n7258) );
  XOR U8766 ( .A(n7261), .B(n7259), .Z(n7260) );
  NANDN U8767 ( .A(n7169), .B(n7171), .Z(n7212) );
  XOR U8768 ( .A(n7262), .B(n7263), .Z(n7171) );
  AND U8769 ( .A(n62), .B(n7264), .Z(n7262) );
  XOR U8770 ( .A(n7263), .B(n7265), .Z(n7264) );
  XNOR U8771 ( .A(n7266), .B(n7267), .Z(n62) );
  AND U8772 ( .A(n7268), .B(n7269), .Z(n7266) );
  XOR U8773 ( .A(n7267), .B(n7182), .Z(n7269) );
  XNOR U8774 ( .A(n7270), .B(n7271), .Z(n7182) );
  ANDN U8775 ( .B(n7272), .A(n7273), .Z(n7270) );
  XOR U8776 ( .A(n7271), .B(n7274), .Z(n7272) );
  XNOR U8777 ( .A(n7267), .B(n7184), .Z(n7268) );
  XOR U8778 ( .A(n7275), .B(n7276), .Z(n7184) );
  AND U8779 ( .A(n66), .B(n7277), .Z(n7275) );
  XOR U8780 ( .A(n7278), .B(n7276), .Z(n7277) );
  XNOR U8781 ( .A(n7279), .B(n7280), .Z(n7267) );
  AND U8782 ( .A(n7281), .B(n7282), .Z(n7279) );
  XNOR U8783 ( .A(n7280), .B(n7209), .Z(n7282) );
  XOR U8784 ( .A(n7273), .B(n7274), .Z(n7209) );
  XNOR U8785 ( .A(n7283), .B(n7284), .Z(n7274) );
  ANDN U8786 ( .B(n7285), .A(n7286), .Z(n7283) );
  XOR U8787 ( .A(n7287), .B(n7288), .Z(n7285) );
  XOR U8788 ( .A(n7289), .B(n7290), .Z(n7273) );
  XNOR U8789 ( .A(n7291), .B(n7292), .Z(n7290) );
  ANDN U8790 ( .B(n7293), .A(n7294), .Z(n7291) );
  XNOR U8791 ( .A(n7295), .B(n7296), .Z(n7293) );
  IV U8792 ( .A(n7271), .Z(n7289) );
  XOR U8793 ( .A(n7297), .B(n7298), .Z(n7271) );
  ANDN U8794 ( .B(n7299), .A(n7300), .Z(n7297) );
  XOR U8795 ( .A(n7298), .B(n7301), .Z(n7299) );
  XOR U8796 ( .A(n7280), .B(n7211), .Z(n7281) );
  XOR U8797 ( .A(n7302), .B(n7303), .Z(n7211) );
  AND U8798 ( .A(n66), .B(n7304), .Z(n7302) );
  XOR U8799 ( .A(n7305), .B(n7303), .Z(n7304) );
  XNOR U8800 ( .A(n7306), .B(n7307), .Z(n7280) );
  NAND U8801 ( .A(n7308), .B(n7309), .Z(n7307) );
  XOR U8802 ( .A(n7310), .B(n7259), .Z(n7309) );
  XOR U8803 ( .A(n7300), .B(n7301), .Z(n7259) );
  XOR U8804 ( .A(n7311), .B(n7288), .Z(n7301) );
  XOR U8805 ( .A(n7312), .B(n7313), .Z(n7288) );
  ANDN U8806 ( .B(n7314), .A(n7315), .Z(n7312) );
  XOR U8807 ( .A(n7313), .B(n7316), .Z(n7314) );
  IV U8808 ( .A(n7286), .Z(n7311) );
  XOR U8809 ( .A(n7284), .B(n7317), .Z(n7286) );
  XOR U8810 ( .A(n7318), .B(n7319), .Z(n7317) );
  ANDN U8811 ( .B(n7320), .A(n7321), .Z(n7318) );
  XOR U8812 ( .A(n7322), .B(n7319), .Z(n7320) );
  IV U8813 ( .A(n7287), .Z(n7284) );
  XOR U8814 ( .A(n7323), .B(n7324), .Z(n7287) );
  ANDN U8815 ( .B(n7325), .A(n7326), .Z(n7323) );
  XOR U8816 ( .A(n7324), .B(n7327), .Z(n7325) );
  XOR U8817 ( .A(n7328), .B(n7329), .Z(n7300) );
  XNOR U8818 ( .A(n7295), .B(n7330), .Z(n7329) );
  IV U8819 ( .A(n7298), .Z(n7330) );
  XOR U8820 ( .A(n7331), .B(n7332), .Z(n7298) );
  ANDN U8821 ( .B(n7333), .A(n7334), .Z(n7331) );
  XOR U8822 ( .A(n7332), .B(n7335), .Z(n7333) );
  XNOR U8823 ( .A(n7336), .B(n7337), .Z(n7295) );
  ANDN U8824 ( .B(n7338), .A(n7339), .Z(n7336) );
  XOR U8825 ( .A(n7337), .B(n7340), .Z(n7338) );
  IV U8826 ( .A(n7294), .Z(n7328) );
  XOR U8827 ( .A(n7292), .B(n7341), .Z(n7294) );
  XOR U8828 ( .A(n7342), .B(n7343), .Z(n7341) );
  ANDN U8829 ( .B(n7344), .A(n7345), .Z(n7342) );
  XOR U8830 ( .A(n7346), .B(n7343), .Z(n7344) );
  IV U8831 ( .A(n7296), .Z(n7292) );
  XOR U8832 ( .A(n7347), .B(n7348), .Z(n7296) );
  ANDN U8833 ( .B(n7349), .A(n7350), .Z(n7347) );
  XOR U8834 ( .A(n7351), .B(n7348), .Z(n7349) );
  IV U8835 ( .A(n7306), .Z(n7310) );
  XOR U8836 ( .A(n7306), .B(n7261), .Z(n7308) );
  XOR U8837 ( .A(n7352), .B(n7353), .Z(n7261) );
  AND U8838 ( .A(n66), .B(n7354), .Z(n7352) );
  XOR U8839 ( .A(n7355), .B(n7353), .Z(n7354) );
  NANDN U8840 ( .A(n7263), .B(n7265), .Z(n7306) );
  XOR U8841 ( .A(n7356), .B(n7357), .Z(n7265) );
  AND U8842 ( .A(n66), .B(n7358), .Z(n7356) );
  XOR U8843 ( .A(n7357), .B(n7359), .Z(n7358) );
  XNOR U8844 ( .A(n7360), .B(n7361), .Z(n66) );
  AND U8845 ( .A(n7362), .B(n7363), .Z(n7360) );
  XOR U8846 ( .A(n7361), .B(n7276), .Z(n7363) );
  XNOR U8847 ( .A(n7364), .B(n7365), .Z(n7276) );
  ANDN U8848 ( .B(n7366), .A(n7367), .Z(n7364) );
  XOR U8849 ( .A(n7365), .B(n7368), .Z(n7366) );
  XNOR U8850 ( .A(n7361), .B(n7278), .Z(n7362) );
  XOR U8851 ( .A(n7369), .B(n7370), .Z(n7278) );
  AND U8852 ( .A(n70), .B(n7371), .Z(n7369) );
  XOR U8853 ( .A(n7372), .B(n7370), .Z(n7371) );
  XNOR U8854 ( .A(n7373), .B(n7374), .Z(n7361) );
  AND U8855 ( .A(n7375), .B(n7376), .Z(n7373) );
  XNOR U8856 ( .A(n7374), .B(n7303), .Z(n7376) );
  XOR U8857 ( .A(n7367), .B(n7368), .Z(n7303) );
  XNOR U8858 ( .A(n7377), .B(n7378), .Z(n7368) );
  ANDN U8859 ( .B(n7379), .A(n7380), .Z(n7377) );
  XOR U8860 ( .A(n7381), .B(n7382), .Z(n7379) );
  XOR U8861 ( .A(n7383), .B(n7384), .Z(n7367) );
  XNOR U8862 ( .A(n7385), .B(n7386), .Z(n7384) );
  ANDN U8863 ( .B(n7387), .A(n7388), .Z(n7385) );
  XNOR U8864 ( .A(n7389), .B(n7390), .Z(n7387) );
  IV U8865 ( .A(n7365), .Z(n7383) );
  XOR U8866 ( .A(n7391), .B(n7392), .Z(n7365) );
  ANDN U8867 ( .B(n7393), .A(n7394), .Z(n7391) );
  XOR U8868 ( .A(n7392), .B(n7395), .Z(n7393) );
  XOR U8869 ( .A(n7374), .B(n7305), .Z(n7375) );
  XOR U8870 ( .A(n7396), .B(n7397), .Z(n7305) );
  AND U8871 ( .A(n70), .B(n7398), .Z(n7396) );
  XOR U8872 ( .A(n7399), .B(n7397), .Z(n7398) );
  XNOR U8873 ( .A(n7400), .B(n7401), .Z(n7374) );
  NAND U8874 ( .A(n7402), .B(n7403), .Z(n7401) );
  XOR U8875 ( .A(n7404), .B(n7353), .Z(n7403) );
  XOR U8876 ( .A(n7394), .B(n7395), .Z(n7353) );
  XOR U8877 ( .A(n7405), .B(n7382), .Z(n7395) );
  XOR U8878 ( .A(n7406), .B(n7407), .Z(n7382) );
  ANDN U8879 ( .B(n7408), .A(n7409), .Z(n7406) );
  XOR U8880 ( .A(n7407), .B(n7410), .Z(n7408) );
  IV U8881 ( .A(n7380), .Z(n7405) );
  XOR U8882 ( .A(n7378), .B(n7411), .Z(n7380) );
  XOR U8883 ( .A(n7412), .B(n7413), .Z(n7411) );
  ANDN U8884 ( .B(n7414), .A(n7415), .Z(n7412) );
  XOR U8885 ( .A(n7416), .B(n7413), .Z(n7414) );
  IV U8886 ( .A(n7381), .Z(n7378) );
  XOR U8887 ( .A(n7417), .B(n7418), .Z(n7381) );
  ANDN U8888 ( .B(n7419), .A(n7420), .Z(n7417) );
  XOR U8889 ( .A(n7418), .B(n7421), .Z(n7419) );
  XOR U8890 ( .A(n7422), .B(n7423), .Z(n7394) );
  XNOR U8891 ( .A(n7389), .B(n7424), .Z(n7423) );
  IV U8892 ( .A(n7392), .Z(n7424) );
  XOR U8893 ( .A(n7425), .B(n7426), .Z(n7392) );
  ANDN U8894 ( .B(n7427), .A(n7428), .Z(n7425) );
  XOR U8895 ( .A(n7426), .B(n7429), .Z(n7427) );
  XNOR U8896 ( .A(n7430), .B(n7431), .Z(n7389) );
  ANDN U8897 ( .B(n7432), .A(n7433), .Z(n7430) );
  XOR U8898 ( .A(n7431), .B(n7434), .Z(n7432) );
  IV U8899 ( .A(n7388), .Z(n7422) );
  XOR U8900 ( .A(n7386), .B(n7435), .Z(n7388) );
  XOR U8901 ( .A(n7436), .B(n7437), .Z(n7435) );
  ANDN U8902 ( .B(n7438), .A(n7439), .Z(n7436) );
  XOR U8903 ( .A(n7440), .B(n7437), .Z(n7438) );
  IV U8904 ( .A(n7390), .Z(n7386) );
  XOR U8905 ( .A(n7441), .B(n7442), .Z(n7390) );
  ANDN U8906 ( .B(n7443), .A(n7444), .Z(n7441) );
  XOR U8907 ( .A(n7445), .B(n7442), .Z(n7443) );
  IV U8908 ( .A(n7400), .Z(n7404) );
  XOR U8909 ( .A(n7400), .B(n7355), .Z(n7402) );
  XOR U8910 ( .A(n7446), .B(n7447), .Z(n7355) );
  AND U8911 ( .A(n70), .B(n7448), .Z(n7446) );
  XOR U8912 ( .A(n7449), .B(n7447), .Z(n7448) );
  NANDN U8913 ( .A(n7357), .B(n7359), .Z(n7400) );
  XOR U8914 ( .A(n7450), .B(n7451), .Z(n7359) );
  AND U8915 ( .A(n70), .B(n7452), .Z(n7450) );
  XOR U8916 ( .A(n7451), .B(n7453), .Z(n7452) );
  XNOR U8917 ( .A(n7454), .B(n7455), .Z(n70) );
  AND U8918 ( .A(n7456), .B(n7457), .Z(n7454) );
  XOR U8919 ( .A(n7455), .B(n7370), .Z(n7457) );
  XNOR U8920 ( .A(n7458), .B(n7459), .Z(n7370) );
  ANDN U8921 ( .B(n7460), .A(n7461), .Z(n7458) );
  XOR U8922 ( .A(n7459), .B(n7462), .Z(n7460) );
  XNOR U8923 ( .A(n7455), .B(n7372), .Z(n7456) );
  XOR U8924 ( .A(n7463), .B(n7464), .Z(n7372) );
  AND U8925 ( .A(n74), .B(n7465), .Z(n7463) );
  XOR U8926 ( .A(n7466), .B(n7464), .Z(n7465) );
  XNOR U8927 ( .A(n7467), .B(n7468), .Z(n7455) );
  AND U8928 ( .A(n7469), .B(n7470), .Z(n7467) );
  XNOR U8929 ( .A(n7468), .B(n7397), .Z(n7470) );
  XOR U8930 ( .A(n7461), .B(n7462), .Z(n7397) );
  XNOR U8931 ( .A(n7471), .B(n7472), .Z(n7462) );
  ANDN U8932 ( .B(n7473), .A(n7474), .Z(n7471) );
  XOR U8933 ( .A(n7475), .B(n7476), .Z(n7473) );
  XOR U8934 ( .A(n7477), .B(n7478), .Z(n7461) );
  XNOR U8935 ( .A(n7479), .B(n7480), .Z(n7478) );
  ANDN U8936 ( .B(n7481), .A(n7482), .Z(n7479) );
  XNOR U8937 ( .A(n7483), .B(n7484), .Z(n7481) );
  IV U8938 ( .A(n7459), .Z(n7477) );
  XOR U8939 ( .A(n7485), .B(n7486), .Z(n7459) );
  ANDN U8940 ( .B(n7487), .A(n7488), .Z(n7485) );
  XOR U8941 ( .A(n7486), .B(n7489), .Z(n7487) );
  XOR U8942 ( .A(n7468), .B(n7399), .Z(n7469) );
  XOR U8943 ( .A(n7490), .B(n7491), .Z(n7399) );
  AND U8944 ( .A(n74), .B(n7492), .Z(n7490) );
  XOR U8945 ( .A(n7493), .B(n7491), .Z(n7492) );
  XNOR U8946 ( .A(n7494), .B(n7495), .Z(n7468) );
  NAND U8947 ( .A(n7496), .B(n7497), .Z(n7495) );
  XOR U8948 ( .A(n7498), .B(n7447), .Z(n7497) );
  XOR U8949 ( .A(n7488), .B(n7489), .Z(n7447) );
  XOR U8950 ( .A(n7499), .B(n7476), .Z(n7489) );
  XOR U8951 ( .A(n7500), .B(n7501), .Z(n7476) );
  ANDN U8952 ( .B(n7502), .A(n7503), .Z(n7500) );
  XOR U8953 ( .A(n7501), .B(n7504), .Z(n7502) );
  IV U8954 ( .A(n7474), .Z(n7499) );
  XOR U8955 ( .A(n7472), .B(n7505), .Z(n7474) );
  XOR U8956 ( .A(n7506), .B(n7507), .Z(n7505) );
  ANDN U8957 ( .B(n7508), .A(n7509), .Z(n7506) );
  XOR U8958 ( .A(n7510), .B(n7507), .Z(n7508) );
  IV U8959 ( .A(n7475), .Z(n7472) );
  XOR U8960 ( .A(n7511), .B(n7512), .Z(n7475) );
  ANDN U8961 ( .B(n7513), .A(n7514), .Z(n7511) );
  XOR U8962 ( .A(n7512), .B(n7515), .Z(n7513) );
  XOR U8963 ( .A(n7516), .B(n7517), .Z(n7488) );
  XNOR U8964 ( .A(n7483), .B(n7518), .Z(n7517) );
  IV U8965 ( .A(n7486), .Z(n7518) );
  XOR U8966 ( .A(n7519), .B(n7520), .Z(n7486) );
  ANDN U8967 ( .B(n7521), .A(n7522), .Z(n7519) );
  XOR U8968 ( .A(n7520), .B(n7523), .Z(n7521) );
  XNOR U8969 ( .A(n7524), .B(n7525), .Z(n7483) );
  ANDN U8970 ( .B(n7526), .A(n7527), .Z(n7524) );
  XOR U8971 ( .A(n7525), .B(n7528), .Z(n7526) );
  IV U8972 ( .A(n7482), .Z(n7516) );
  XOR U8973 ( .A(n7480), .B(n7529), .Z(n7482) );
  XOR U8974 ( .A(n7530), .B(n7531), .Z(n7529) );
  ANDN U8975 ( .B(n7532), .A(n7533), .Z(n7530) );
  XOR U8976 ( .A(n7534), .B(n7531), .Z(n7532) );
  IV U8977 ( .A(n7484), .Z(n7480) );
  XOR U8978 ( .A(n7535), .B(n7536), .Z(n7484) );
  ANDN U8979 ( .B(n7537), .A(n7538), .Z(n7535) );
  XOR U8980 ( .A(n7539), .B(n7536), .Z(n7537) );
  IV U8981 ( .A(n7494), .Z(n7498) );
  XOR U8982 ( .A(n7494), .B(n7449), .Z(n7496) );
  XOR U8983 ( .A(n7540), .B(n7541), .Z(n7449) );
  AND U8984 ( .A(n74), .B(n7542), .Z(n7540) );
  XOR U8985 ( .A(n7543), .B(n7541), .Z(n7542) );
  NANDN U8986 ( .A(n7451), .B(n7453), .Z(n7494) );
  XOR U8987 ( .A(n7544), .B(n7545), .Z(n7453) );
  AND U8988 ( .A(n74), .B(n7546), .Z(n7544) );
  XOR U8989 ( .A(n7545), .B(n7547), .Z(n7546) );
  XNOR U8990 ( .A(n7548), .B(n7549), .Z(n74) );
  AND U8991 ( .A(n7550), .B(n7551), .Z(n7548) );
  XOR U8992 ( .A(n7549), .B(n7464), .Z(n7551) );
  XNOR U8993 ( .A(n7552), .B(n7553), .Z(n7464) );
  ANDN U8994 ( .B(n7554), .A(n7555), .Z(n7552) );
  XOR U8995 ( .A(n7553), .B(n7556), .Z(n7554) );
  XNOR U8996 ( .A(n7549), .B(n7466), .Z(n7550) );
  XOR U8997 ( .A(n7557), .B(n7558), .Z(n7466) );
  AND U8998 ( .A(n78), .B(n7559), .Z(n7557) );
  XOR U8999 ( .A(n7560), .B(n7558), .Z(n7559) );
  XNOR U9000 ( .A(n7561), .B(n7562), .Z(n7549) );
  AND U9001 ( .A(n7563), .B(n7564), .Z(n7561) );
  XNOR U9002 ( .A(n7562), .B(n7491), .Z(n7564) );
  XOR U9003 ( .A(n7555), .B(n7556), .Z(n7491) );
  XNOR U9004 ( .A(n7565), .B(n7566), .Z(n7556) );
  ANDN U9005 ( .B(n7567), .A(n7568), .Z(n7565) );
  XOR U9006 ( .A(n7569), .B(n7570), .Z(n7567) );
  XOR U9007 ( .A(n7571), .B(n7572), .Z(n7555) );
  XNOR U9008 ( .A(n7573), .B(n7574), .Z(n7572) );
  ANDN U9009 ( .B(n7575), .A(n7576), .Z(n7573) );
  XNOR U9010 ( .A(n7577), .B(n7578), .Z(n7575) );
  IV U9011 ( .A(n7553), .Z(n7571) );
  XOR U9012 ( .A(n7579), .B(n7580), .Z(n7553) );
  ANDN U9013 ( .B(n7581), .A(n7582), .Z(n7579) );
  XOR U9014 ( .A(n7580), .B(n7583), .Z(n7581) );
  XOR U9015 ( .A(n7562), .B(n7493), .Z(n7563) );
  XOR U9016 ( .A(n7584), .B(n7585), .Z(n7493) );
  AND U9017 ( .A(n78), .B(n7586), .Z(n7584) );
  XOR U9018 ( .A(n7587), .B(n7585), .Z(n7586) );
  XNOR U9019 ( .A(n7588), .B(n7589), .Z(n7562) );
  NAND U9020 ( .A(n7590), .B(n7591), .Z(n7589) );
  XOR U9021 ( .A(n7592), .B(n7541), .Z(n7591) );
  XOR U9022 ( .A(n7582), .B(n7583), .Z(n7541) );
  XOR U9023 ( .A(n7593), .B(n7570), .Z(n7583) );
  XOR U9024 ( .A(n7594), .B(n7595), .Z(n7570) );
  ANDN U9025 ( .B(n7596), .A(n7597), .Z(n7594) );
  XOR U9026 ( .A(n7595), .B(n7598), .Z(n7596) );
  IV U9027 ( .A(n7568), .Z(n7593) );
  XOR U9028 ( .A(n7566), .B(n7599), .Z(n7568) );
  XOR U9029 ( .A(n7600), .B(n7601), .Z(n7599) );
  ANDN U9030 ( .B(n7602), .A(n7603), .Z(n7600) );
  XOR U9031 ( .A(n7604), .B(n7601), .Z(n7602) );
  IV U9032 ( .A(n7569), .Z(n7566) );
  XOR U9033 ( .A(n7605), .B(n7606), .Z(n7569) );
  ANDN U9034 ( .B(n7607), .A(n7608), .Z(n7605) );
  XOR U9035 ( .A(n7606), .B(n7609), .Z(n7607) );
  XOR U9036 ( .A(n7610), .B(n7611), .Z(n7582) );
  XNOR U9037 ( .A(n7577), .B(n7612), .Z(n7611) );
  IV U9038 ( .A(n7580), .Z(n7612) );
  XOR U9039 ( .A(n7613), .B(n7614), .Z(n7580) );
  ANDN U9040 ( .B(n7615), .A(n7616), .Z(n7613) );
  XOR U9041 ( .A(n7614), .B(n7617), .Z(n7615) );
  XNOR U9042 ( .A(n7618), .B(n7619), .Z(n7577) );
  ANDN U9043 ( .B(n7620), .A(n7621), .Z(n7618) );
  XOR U9044 ( .A(n7619), .B(n7622), .Z(n7620) );
  IV U9045 ( .A(n7576), .Z(n7610) );
  XOR U9046 ( .A(n7574), .B(n7623), .Z(n7576) );
  XOR U9047 ( .A(n7624), .B(n7625), .Z(n7623) );
  ANDN U9048 ( .B(n7626), .A(n7627), .Z(n7624) );
  XOR U9049 ( .A(n7628), .B(n7625), .Z(n7626) );
  IV U9050 ( .A(n7578), .Z(n7574) );
  XOR U9051 ( .A(n7629), .B(n7630), .Z(n7578) );
  ANDN U9052 ( .B(n7631), .A(n7632), .Z(n7629) );
  XOR U9053 ( .A(n7633), .B(n7630), .Z(n7631) );
  IV U9054 ( .A(n7588), .Z(n7592) );
  XOR U9055 ( .A(n7588), .B(n7543), .Z(n7590) );
  XOR U9056 ( .A(n7634), .B(n7635), .Z(n7543) );
  AND U9057 ( .A(n78), .B(n7636), .Z(n7634) );
  XOR U9058 ( .A(n7637), .B(n7635), .Z(n7636) );
  NANDN U9059 ( .A(n7545), .B(n7547), .Z(n7588) );
  XOR U9060 ( .A(n7638), .B(n7639), .Z(n7547) );
  AND U9061 ( .A(n78), .B(n7640), .Z(n7638) );
  XOR U9062 ( .A(n7639), .B(n7641), .Z(n7640) );
  XNOR U9063 ( .A(n7642), .B(n7643), .Z(n78) );
  AND U9064 ( .A(n7644), .B(n7645), .Z(n7642) );
  XOR U9065 ( .A(n7643), .B(n7558), .Z(n7645) );
  XNOR U9066 ( .A(n7646), .B(n7647), .Z(n7558) );
  ANDN U9067 ( .B(n7648), .A(n7649), .Z(n7646) );
  XOR U9068 ( .A(n7647), .B(n7650), .Z(n7648) );
  XNOR U9069 ( .A(n7643), .B(n7560), .Z(n7644) );
  XOR U9070 ( .A(n7651), .B(n7652), .Z(n7560) );
  AND U9071 ( .A(n82), .B(n7653), .Z(n7651) );
  XOR U9072 ( .A(n7654), .B(n7652), .Z(n7653) );
  XNOR U9073 ( .A(n7655), .B(n7656), .Z(n7643) );
  AND U9074 ( .A(n7657), .B(n7658), .Z(n7655) );
  XNOR U9075 ( .A(n7656), .B(n7585), .Z(n7658) );
  XOR U9076 ( .A(n7649), .B(n7650), .Z(n7585) );
  XNOR U9077 ( .A(n7659), .B(n7660), .Z(n7650) );
  ANDN U9078 ( .B(n7661), .A(n7662), .Z(n7659) );
  XOR U9079 ( .A(n7663), .B(n7664), .Z(n7661) );
  XOR U9080 ( .A(n7665), .B(n7666), .Z(n7649) );
  XNOR U9081 ( .A(n7667), .B(n7668), .Z(n7666) );
  ANDN U9082 ( .B(n7669), .A(n7670), .Z(n7667) );
  XNOR U9083 ( .A(n7671), .B(n7672), .Z(n7669) );
  IV U9084 ( .A(n7647), .Z(n7665) );
  XOR U9085 ( .A(n7673), .B(n7674), .Z(n7647) );
  ANDN U9086 ( .B(n7675), .A(n7676), .Z(n7673) );
  XOR U9087 ( .A(n7674), .B(n7677), .Z(n7675) );
  XOR U9088 ( .A(n7656), .B(n7587), .Z(n7657) );
  XOR U9089 ( .A(n7678), .B(n7679), .Z(n7587) );
  AND U9090 ( .A(n82), .B(n7680), .Z(n7678) );
  XOR U9091 ( .A(n7681), .B(n7679), .Z(n7680) );
  XNOR U9092 ( .A(n7682), .B(n7683), .Z(n7656) );
  NAND U9093 ( .A(n7684), .B(n7685), .Z(n7683) );
  XOR U9094 ( .A(n7686), .B(n7635), .Z(n7685) );
  XOR U9095 ( .A(n7676), .B(n7677), .Z(n7635) );
  XOR U9096 ( .A(n7687), .B(n7664), .Z(n7677) );
  XOR U9097 ( .A(n7688), .B(n7689), .Z(n7664) );
  ANDN U9098 ( .B(n7690), .A(n7691), .Z(n7688) );
  XOR U9099 ( .A(n7689), .B(n7692), .Z(n7690) );
  IV U9100 ( .A(n7662), .Z(n7687) );
  XOR U9101 ( .A(n7660), .B(n7693), .Z(n7662) );
  XOR U9102 ( .A(n7694), .B(n7695), .Z(n7693) );
  ANDN U9103 ( .B(n7696), .A(n7697), .Z(n7694) );
  XOR U9104 ( .A(n7698), .B(n7695), .Z(n7696) );
  IV U9105 ( .A(n7663), .Z(n7660) );
  XOR U9106 ( .A(n7699), .B(n7700), .Z(n7663) );
  ANDN U9107 ( .B(n7701), .A(n7702), .Z(n7699) );
  XOR U9108 ( .A(n7700), .B(n7703), .Z(n7701) );
  XOR U9109 ( .A(n7704), .B(n7705), .Z(n7676) );
  XNOR U9110 ( .A(n7671), .B(n7706), .Z(n7705) );
  IV U9111 ( .A(n7674), .Z(n7706) );
  XOR U9112 ( .A(n7707), .B(n7708), .Z(n7674) );
  ANDN U9113 ( .B(n7709), .A(n7710), .Z(n7707) );
  XOR U9114 ( .A(n7708), .B(n7711), .Z(n7709) );
  XNOR U9115 ( .A(n7712), .B(n7713), .Z(n7671) );
  ANDN U9116 ( .B(n7714), .A(n7715), .Z(n7712) );
  XOR U9117 ( .A(n7713), .B(n7716), .Z(n7714) );
  IV U9118 ( .A(n7670), .Z(n7704) );
  XOR U9119 ( .A(n7668), .B(n7717), .Z(n7670) );
  XOR U9120 ( .A(n7718), .B(n7719), .Z(n7717) );
  ANDN U9121 ( .B(n7720), .A(n7721), .Z(n7718) );
  XOR U9122 ( .A(n7722), .B(n7719), .Z(n7720) );
  IV U9123 ( .A(n7672), .Z(n7668) );
  XOR U9124 ( .A(n7723), .B(n7724), .Z(n7672) );
  ANDN U9125 ( .B(n7725), .A(n7726), .Z(n7723) );
  XOR U9126 ( .A(n7727), .B(n7724), .Z(n7725) );
  IV U9127 ( .A(n7682), .Z(n7686) );
  XOR U9128 ( .A(n7682), .B(n7637), .Z(n7684) );
  XOR U9129 ( .A(n7728), .B(n7729), .Z(n7637) );
  AND U9130 ( .A(n82), .B(n7730), .Z(n7728) );
  XOR U9131 ( .A(n7731), .B(n7729), .Z(n7730) );
  NANDN U9132 ( .A(n7639), .B(n7641), .Z(n7682) );
  XOR U9133 ( .A(n7732), .B(n7733), .Z(n7641) );
  AND U9134 ( .A(n82), .B(n7734), .Z(n7732) );
  XOR U9135 ( .A(n7733), .B(n7735), .Z(n7734) );
  XNOR U9136 ( .A(n7736), .B(n7737), .Z(n82) );
  AND U9137 ( .A(n7738), .B(n7739), .Z(n7736) );
  XOR U9138 ( .A(n7737), .B(n7652), .Z(n7739) );
  XNOR U9139 ( .A(n7740), .B(n7741), .Z(n7652) );
  ANDN U9140 ( .B(n7742), .A(n7743), .Z(n7740) );
  XOR U9141 ( .A(n7741), .B(n7744), .Z(n7742) );
  XNOR U9142 ( .A(n7737), .B(n7654), .Z(n7738) );
  XOR U9143 ( .A(n7745), .B(n7746), .Z(n7654) );
  AND U9144 ( .A(n86), .B(n7747), .Z(n7745) );
  XOR U9145 ( .A(n7748), .B(n7746), .Z(n7747) );
  XNOR U9146 ( .A(n7749), .B(n7750), .Z(n7737) );
  AND U9147 ( .A(n7751), .B(n7752), .Z(n7749) );
  XNOR U9148 ( .A(n7750), .B(n7679), .Z(n7752) );
  XOR U9149 ( .A(n7743), .B(n7744), .Z(n7679) );
  XNOR U9150 ( .A(n7753), .B(n7754), .Z(n7744) );
  ANDN U9151 ( .B(n7755), .A(n7756), .Z(n7753) );
  XOR U9152 ( .A(n7757), .B(n7758), .Z(n7755) );
  XOR U9153 ( .A(n7759), .B(n7760), .Z(n7743) );
  XNOR U9154 ( .A(n7761), .B(n7762), .Z(n7760) );
  ANDN U9155 ( .B(n7763), .A(n7764), .Z(n7761) );
  XNOR U9156 ( .A(n7765), .B(n7766), .Z(n7763) );
  IV U9157 ( .A(n7741), .Z(n7759) );
  XOR U9158 ( .A(n7767), .B(n7768), .Z(n7741) );
  ANDN U9159 ( .B(n7769), .A(n7770), .Z(n7767) );
  XOR U9160 ( .A(n7768), .B(n7771), .Z(n7769) );
  XOR U9161 ( .A(n7750), .B(n7681), .Z(n7751) );
  XOR U9162 ( .A(n7772), .B(n7773), .Z(n7681) );
  AND U9163 ( .A(n86), .B(n7774), .Z(n7772) );
  XOR U9164 ( .A(n7775), .B(n7773), .Z(n7774) );
  XNOR U9165 ( .A(n7776), .B(n7777), .Z(n7750) );
  NAND U9166 ( .A(n7778), .B(n7779), .Z(n7777) );
  XOR U9167 ( .A(n7780), .B(n7729), .Z(n7779) );
  XOR U9168 ( .A(n7770), .B(n7771), .Z(n7729) );
  XOR U9169 ( .A(n7781), .B(n7758), .Z(n7771) );
  XOR U9170 ( .A(n7782), .B(n7783), .Z(n7758) );
  ANDN U9171 ( .B(n7784), .A(n7785), .Z(n7782) );
  XOR U9172 ( .A(n7783), .B(n7786), .Z(n7784) );
  IV U9173 ( .A(n7756), .Z(n7781) );
  XOR U9174 ( .A(n7754), .B(n7787), .Z(n7756) );
  XOR U9175 ( .A(n7788), .B(n7789), .Z(n7787) );
  ANDN U9176 ( .B(n7790), .A(n7791), .Z(n7788) );
  XOR U9177 ( .A(n7792), .B(n7789), .Z(n7790) );
  IV U9178 ( .A(n7757), .Z(n7754) );
  XOR U9179 ( .A(n7793), .B(n7794), .Z(n7757) );
  ANDN U9180 ( .B(n7795), .A(n7796), .Z(n7793) );
  XOR U9181 ( .A(n7794), .B(n7797), .Z(n7795) );
  XOR U9182 ( .A(n7798), .B(n7799), .Z(n7770) );
  XNOR U9183 ( .A(n7765), .B(n7800), .Z(n7799) );
  IV U9184 ( .A(n7768), .Z(n7800) );
  XOR U9185 ( .A(n7801), .B(n7802), .Z(n7768) );
  ANDN U9186 ( .B(n7803), .A(n7804), .Z(n7801) );
  XOR U9187 ( .A(n7802), .B(n7805), .Z(n7803) );
  XNOR U9188 ( .A(n7806), .B(n7807), .Z(n7765) );
  ANDN U9189 ( .B(n7808), .A(n7809), .Z(n7806) );
  XOR U9190 ( .A(n7807), .B(n7810), .Z(n7808) );
  IV U9191 ( .A(n7764), .Z(n7798) );
  XOR U9192 ( .A(n7762), .B(n7811), .Z(n7764) );
  XOR U9193 ( .A(n7812), .B(n7813), .Z(n7811) );
  ANDN U9194 ( .B(n7814), .A(n7815), .Z(n7812) );
  XOR U9195 ( .A(n7816), .B(n7813), .Z(n7814) );
  IV U9196 ( .A(n7766), .Z(n7762) );
  XOR U9197 ( .A(n7817), .B(n7818), .Z(n7766) );
  ANDN U9198 ( .B(n7819), .A(n7820), .Z(n7817) );
  XOR U9199 ( .A(n7821), .B(n7818), .Z(n7819) );
  IV U9200 ( .A(n7776), .Z(n7780) );
  XOR U9201 ( .A(n7776), .B(n7731), .Z(n7778) );
  XOR U9202 ( .A(n7822), .B(n7823), .Z(n7731) );
  AND U9203 ( .A(n86), .B(n7824), .Z(n7822) );
  XOR U9204 ( .A(n7825), .B(n7823), .Z(n7824) );
  NANDN U9205 ( .A(n7733), .B(n7735), .Z(n7776) );
  XOR U9206 ( .A(n7826), .B(n7827), .Z(n7735) );
  AND U9207 ( .A(n86), .B(n7828), .Z(n7826) );
  XOR U9208 ( .A(n7827), .B(n7829), .Z(n7828) );
  XNOR U9209 ( .A(n7830), .B(n7831), .Z(n86) );
  AND U9210 ( .A(n7832), .B(n7833), .Z(n7830) );
  XOR U9211 ( .A(n7831), .B(n7746), .Z(n7833) );
  XNOR U9212 ( .A(n7834), .B(n7835), .Z(n7746) );
  ANDN U9213 ( .B(n7836), .A(n7837), .Z(n7834) );
  XOR U9214 ( .A(n7835), .B(n7838), .Z(n7836) );
  XNOR U9215 ( .A(n7831), .B(n7748), .Z(n7832) );
  XOR U9216 ( .A(n7839), .B(n7840), .Z(n7748) );
  AND U9217 ( .A(n90), .B(n7841), .Z(n7839) );
  XOR U9218 ( .A(n7842), .B(n7840), .Z(n7841) );
  XNOR U9219 ( .A(n7843), .B(n7844), .Z(n7831) );
  AND U9220 ( .A(n7845), .B(n7846), .Z(n7843) );
  XNOR U9221 ( .A(n7844), .B(n7773), .Z(n7846) );
  XOR U9222 ( .A(n7837), .B(n7838), .Z(n7773) );
  XNOR U9223 ( .A(n7847), .B(n7848), .Z(n7838) );
  ANDN U9224 ( .B(n7849), .A(n7850), .Z(n7847) );
  XOR U9225 ( .A(n7851), .B(n7852), .Z(n7849) );
  XOR U9226 ( .A(n7853), .B(n7854), .Z(n7837) );
  XNOR U9227 ( .A(n7855), .B(n7856), .Z(n7854) );
  ANDN U9228 ( .B(n7857), .A(n7858), .Z(n7855) );
  XNOR U9229 ( .A(n7859), .B(n7860), .Z(n7857) );
  IV U9230 ( .A(n7835), .Z(n7853) );
  XOR U9231 ( .A(n7861), .B(n7862), .Z(n7835) );
  ANDN U9232 ( .B(n7863), .A(n7864), .Z(n7861) );
  XOR U9233 ( .A(n7862), .B(n7865), .Z(n7863) );
  XOR U9234 ( .A(n7844), .B(n7775), .Z(n7845) );
  XOR U9235 ( .A(n7866), .B(n7867), .Z(n7775) );
  AND U9236 ( .A(n90), .B(n7868), .Z(n7866) );
  XOR U9237 ( .A(n7869), .B(n7867), .Z(n7868) );
  XNOR U9238 ( .A(n7870), .B(n7871), .Z(n7844) );
  NAND U9239 ( .A(n7872), .B(n7873), .Z(n7871) );
  XOR U9240 ( .A(n7874), .B(n7823), .Z(n7873) );
  XOR U9241 ( .A(n7864), .B(n7865), .Z(n7823) );
  XOR U9242 ( .A(n7875), .B(n7852), .Z(n7865) );
  XOR U9243 ( .A(n7876), .B(n7877), .Z(n7852) );
  ANDN U9244 ( .B(n7878), .A(n7879), .Z(n7876) );
  XOR U9245 ( .A(n7877), .B(n7880), .Z(n7878) );
  IV U9246 ( .A(n7850), .Z(n7875) );
  XOR U9247 ( .A(n7848), .B(n7881), .Z(n7850) );
  XOR U9248 ( .A(n7882), .B(n7883), .Z(n7881) );
  ANDN U9249 ( .B(n7884), .A(n7885), .Z(n7882) );
  XOR U9250 ( .A(n7886), .B(n7883), .Z(n7884) );
  IV U9251 ( .A(n7851), .Z(n7848) );
  XOR U9252 ( .A(n7887), .B(n7888), .Z(n7851) );
  ANDN U9253 ( .B(n7889), .A(n7890), .Z(n7887) );
  XOR U9254 ( .A(n7888), .B(n7891), .Z(n7889) );
  XOR U9255 ( .A(n7892), .B(n7893), .Z(n7864) );
  XNOR U9256 ( .A(n7859), .B(n7894), .Z(n7893) );
  IV U9257 ( .A(n7862), .Z(n7894) );
  XOR U9258 ( .A(n7895), .B(n7896), .Z(n7862) );
  ANDN U9259 ( .B(n7897), .A(n7898), .Z(n7895) );
  XOR U9260 ( .A(n7896), .B(n7899), .Z(n7897) );
  XNOR U9261 ( .A(n7900), .B(n7901), .Z(n7859) );
  ANDN U9262 ( .B(n7902), .A(n7903), .Z(n7900) );
  XOR U9263 ( .A(n7901), .B(n7904), .Z(n7902) );
  IV U9264 ( .A(n7858), .Z(n7892) );
  XOR U9265 ( .A(n7856), .B(n7905), .Z(n7858) );
  XOR U9266 ( .A(n7906), .B(n7907), .Z(n7905) );
  ANDN U9267 ( .B(n7908), .A(n7909), .Z(n7906) );
  XOR U9268 ( .A(n7910), .B(n7907), .Z(n7908) );
  IV U9269 ( .A(n7860), .Z(n7856) );
  XOR U9270 ( .A(n7911), .B(n7912), .Z(n7860) );
  ANDN U9271 ( .B(n7913), .A(n7914), .Z(n7911) );
  XOR U9272 ( .A(n7915), .B(n7912), .Z(n7913) );
  IV U9273 ( .A(n7870), .Z(n7874) );
  XOR U9274 ( .A(n7870), .B(n7825), .Z(n7872) );
  XOR U9275 ( .A(n7916), .B(n7917), .Z(n7825) );
  AND U9276 ( .A(n90), .B(n7918), .Z(n7916) );
  XOR U9277 ( .A(n7919), .B(n7917), .Z(n7918) );
  NANDN U9278 ( .A(n7827), .B(n7829), .Z(n7870) );
  XOR U9279 ( .A(n7920), .B(n7921), .Z(n7829) );
  AND U9280 ( .A(n90), .B(n7922), .Z(n7920) );
  XOR U9281 ( .A(n7921), .B(n7923), .Z(n7922) );
  XNOR U9282 ( .A(n7924), .B(n7925), .Z(n90) );
  AND U9283 ( .A(n7926), .B(n7927), .Z(n7924) );
  XOR U9284 ( .A(n7925), .B(n7840), .Z(n7927) );
  XNOR U9285 ( .A(n7928), .B(n7929), .Z(n7840) );
  ANDN U9286 ( .B(n7930), .A(n7931), .Z(n7928) );
  XOR U9287 ( .A(n7929), .B(n7932), .Z(n7930) );
  XNOR U9288 ( .A(n7925), .B(n7842), .Z(n7926) );
  XOR U9289 ( .A(n7933), .B(n7934), .Z(n7842) );
  AND U9290 ( .A(n94), .B(n7935), .Z(n7933) );
  XOR U9291 ( .A(n7936), .B(n7934), .Z(n7935) );
  XNOR U9292 ( .A(n7937), .B(n7938), .Z(n7925) );
  AND U9293 ( .A(n7939), .B(n7940), .Z(n7937) );
  XNOR U9294 ( .A(n7938), .B(n7867), .Z(n7940) );
  XOR U9295 ( .A(n7931), .B(n7932), .Z(n7867) );
  XNOR U9296 ( .A(n7941), .B(n7942), .Z(n7932) );
  ANDN U9297 ( .B(n7943), .A(n7944), .Z(n7941) );
  XOR U9298 ( .A(n7945), .B(n7946), .Z(n7943) );
  XOR U9299 ( .A(n7947), .B(n7948), .Z(n7931) );
  XNOR U9300 ( .A(n7949), .B(n7950), .Z(n7948) );
  ANDN U9301 ( .B(n7951), .A(n7952), .Z(n7949) );
  XNOR U9302 ( .A(n7953), .B(n7954), .Z(n7951) );
  IV U9303 ( .A(n7929), .Z(n7947) );
  XOR U9304 ( .A(n7955), .B(n7956), .Z(n7929) );
  ANDN U9305 ( .B(n7957), .A(n7958), .Z(n7955) );
  XOR U9306 ( .A(n7956), .B(n7959), .Z(n7957) );
  XOR U9307 ( .A(n7938), .B(n7869), .Z(n7939) );
  XOR U9308 ( .A(n7960), .B(n7961), .Z(n7869) );
  AND U9309 ( .A(n94), .B(n7962), .Z(n7960) );
  XOR U9310 ( .A(n7963), .B(n7961), .Z(n7962) );
  XNOR U9311 ( .A(n7964), .B(n7965), .Z(n7938) );
  NAND U9312 ( .A(n7966), .B(n7967), .Z(n7965) );
  XOR U9313 ( .A(n7968), .B(n7917), .Z(n7967) );
  XOR U9314 ( .A(n7958), .B(n7959), .Z(n7917) );
  XOR U9315 ( .A(n7969), .B(n7946), .Z(n7959) );
  XOR U9316 ( .A(n7970), .B(n7971), .Z(n7946) );
  ANDN U9317 ( .B(n7972), .A(n7973), .Z(n7970) );
  XOR U9318 ( .A(n7971), .B(n7974), .Z(n7972) );
  IV U9319 ( .A(n7944), .Z(n7969) );
  XOR U9320 ( .A(n7942), .B(n7975), .Z(n7944) );
  XOR U9321 ( .A(n7976), .B(n7977), .Z(n7975) );
  ANDN U9322 ( .B(n7978), .A(n7979), .Z(n7976) );
  XOR U9323 ( .A(n7980), .B(n7977), .Z(n7978) );
  IV U9324 ( .A(n7945), .Z(n7942) );
  XOR U9325 ( .A(n7981), .B(n7982), .Z(n7945) );
  ANDN U9326 ( .B(n7983), .A(n7984), .Z(n7981) );
  XOR U9327 ( .A(n7982), .B(n7985), .Z(n7983) );
  XOR U9328 ( .A(n7986), .B(n7987), .Z(n7958) );
  XNOR U9329 ( .A(n7953), .B(n7988), .Z(n7987) );
  IV U9330 ( .A(n7956), .Z(n7988) );
  XOR U9331 ( .A(n7989), .B(n7990), .Z(n7956) );
  ANDN U9332 ( .B(n7991), .A(n7992), .Z(n7989) );
  XOR U9333 ( .A(n7990), .B(n7993), .Z(n7991) );
  XNOR U9334 ( .A(n7994), .B(n7995), .Z(n7953) );
  ANDN U9335 ( .B(n7996), .A(n7997), .Z(n7994) );
  XOR U9336 ( .A(n7995), .B(n7998), .Z(n7996) );
  IV U9337 ( .A(n7952), .Z(n7986) );
  XOR U9338 ( .A(n7950), .B(n7999), .Z(n7952) );
  XOR U9339 ( .A(n8000), .B(n8001), .Z(n7999) );
  ANDN U9340 ( .B(n8002), .A(n8003), .Z(n8000) );
  XOR U9341 ( .A(n8004), .B(n8001), .Z(n8002) );
  IV U9342 ( .A(n7954), .Z(n7950) );
  XOR U9343 ( .A(n8005), .B(n8006), .Z(n7954) );
  ANDN U9344 ( .B(n8007), .A(n8008), .Z(n8005) );
  XOR U9345 ( .A(n8009), .B(n8006), .Z(n8007) );
  IV U9346 ( .A(n7964), .Z(n7968) );
  XOR U9347 ( .A(n7964), .B(n7919), .Z(n7966) );
  XOR U9348 ( .A(n8010), .B(n8011), .Z(n7919) );
  AND U9349 ( .A(n94), .B(n8012), .Z(n8010) );
  XOR U9350 ( .A(n8013), .B(n8011), .Z(n8012) );
  NANDN U9351 ( .A(n7921), .B(n7923), .Z(n7964) );
  XOR U9352 ( .A(n8014), .B(n8015), .Z(n7923) );
  AND U9353 ( .A(n94), .B(n8016), .Z(n8014) );
  XOR U9354 ( .A(n8015), .B(n8017), .Z(n8016) );
  XNOR U9355 ( .A(n8018), .B(n8019), .Z(n94) );
  AND U9356 ( .A(n8020), .B(n8021), .Z(n8018) );
  XOR U9357 ( .A(n8019), .B(n7934), .Z(n8021) );
  XNOR U9358 ( .A(n8022), .B(n8023), .Z(n7934) );
  ANDN U9359 ( .B(n8024), .A(n8025), .Z(n8022) );
  XOR U9360 ( .A(n8023), .B(n8026), .Z(n8024) );
  XNOR U9361 ( .A(n8019), .B(n7936), .Z(n8020) );
  XOR U9362 ( .A(n8027), .B(n8028), .Z(n7936) );
  AND U9363 ( .A(n98), .B(n8029), .Z(n8027) );
  XOR U9364 ( .A(n8030), .B(n8028), .Z(n8029) );
  XNOR U9365 ( .A(n8031), .B(n8032), .Z(n8019) );
  AND U9366 ( .A(n8033), .B(n8034), .Z(n8031) );
  XNOR U9367 ( .A(n8032), .B(n7961), .Z(n8034) );
  XOR U9368 ( .A(n8025), .B(n8026), .Z(n7961) );
  XNOR U9369 ( .A(n8035), .B(n8036), .Z(n8026) );
  ANDN U9370 ( .B(n8037), .A(n8038), .Z(n8035) );
  XOR U9371 ( .A(n8039), .B(n8040), .Z(n8037) );
  XOR U9372 ( .A(n8041), .B(n8042), .Z(n8025) );
  XNOR U9373 ( .A(n8043), .B(n8044), .Z(n8042) );
  ANDN U9374 ( .B(n8045), .A(n8046), .Z(n8043) );
  XNOR U9375 ( .A(n8047), .B(n8048), .Z(n8045) );
  IV U9376 ( .A(n8023), .Z(n8041) );
  XOR U9377 ( .A(n8049), .B(n8050), .Z(n8023) );
  ANDN U9378 ( .B(n8051), .A(n8052), .Z(n8049) );
  XOR U9379 ( .A(n8050), .B(n8053), .Z(n8051) );
  XOR U9380 ( .A(n8032), .B(n7963), .Z(n8033) );
  XOR U9381 ( .A(n8054), .B(n8055), .Z(n7963) );
  AND U9382 ( .A(n98), .B(n8056), .Z(n8054) );
  XOR U9383 ( .A(n8057), .B(n8055), .Z(n8056) );
  XNOR U9384 ( .A(n8058), .B(n8059), .Z(n8032) );
  NAND U9385 ( .A(n8060), .B(n8061), .Z(n8059) );
  XOR U9386 ( .A(n8062), .B(n8011), .Z(n8061) );
  XOR U9387 ( .A(n8052), .B(n8053), .Z(n8011) );
  XOR U9388 ( .A(n8063), .B(n8040), .Z(n8053) );
  XOR U9389 ( .A(n8064), .B(n8065), .Z(n8040) );
  ANDN U9390 ( .B(n8066), .A(n8067), .Z(n8064) );
  XOR U9391 ( .A(n8065), .B(n8068), .Z(n8066) );
  IV U9392 ( .A(n8038), .Z(n8063) );
  XOR U9393 ( .A(n8036), .B(n8069), .Z(n8038) );
  XOR U9394 ( .A(n8070), .B(n8071), .Z(n8069) );
  ANDN U9395 ( .B(n8072), .A(n8073), .Z(n8070) );
  XOR U9396 ( .A(n8074), .B(n8071), .Z(n8072) );
  IV U9397 ( .A(n8039), .Z(n8036) );
  XOR U9398 ( .A(n8075), .B(n8076), .Z(n8039) );
  ANDN U9399 ( .B(n8077), .A(n8078), .Z(n8075) );
  XOR U9400 ( .A(n8076), .B(n8079), .Z(n8077) );
  XOR U9401 ( .A(n8080), .B(n8081), .Z(n8052) );
  XNOR U9402 ( .A(n8047), .B(n8082), .Z(n8081) );
  IV U9403 ( .A(n8050), .Z(n8082) );
  XOR U9404 ( .A(n8083), .B(n8084), .Z(n8050) );
  ANDN U9405 ( .B(n8085), .A(n8086), .Z(n8083) );
  XOR U9406 ( .A(n8084), .B(n8087), .Z(n8085) );
  XNOR U9407 ( .A(n8088), .B(n8089), .Z(n8047) );
  ANDN U9408 ( .B(n8090), .A(n8091), .Z(n8088) );
  XOR U9409 ( .A(n8089), .B(n8092), .Z(n8090) );
  IV U9410 ( .A(n8046), .Z(n8080) );
  XOR U9411 ( .A(n8044), .B(n8093), .Z(n8046) );
  XOR U9412 ( .A(n8094), .B(n8095), .Z(n8093) );
  ANDN U9413 ( .B(n8096), .A(n8097), .Z(n8094) );
  XOR U9414 ( .A(n8098), .B(n8095), .Z(n8096) );
  IV U9415 ( .A(n8048), .Z(n8044) );
  XOR U9416 ( .A(n8099), .B(n8100), .Z(n8048) );
  ANDN U9417 ( .B(n8101), .A(n8102), .Z(n8099) );
  XOR U9418 ( .A(n8103), .B(n8100), .Z(n8101) );
  IV U9419 ( .A(n8058), .Z(n8062) );
  XOR U9420 ( .A(n8058), .B(n8013), .Z(n8060) );
  XOR U9421 ( .A(n8104), .B(n8105), .Z(n8013) );
  AND U9422 ( .A(n98), .B(n8106), .Z(n8104) );
  XOR U9423 ( .A(n8107), .B(n8105), .Z(n8106) );
  NANDN U9424 ( .A(n8015), .B(n8017), .Z(n8058) );
  XOR U9425 ( .A(n8108), .B(n8109), .Z(n8017) );
  AND U9426 ( .A(n98), .B(n8110), .Z(n8108) );
  XOR U9427 ( .A(n8109), .B(n8111), .Z(n8110) );
  XNOR U9428 ( .A(n8112), .B(n8113), .Z(n98) );
  AND U9429 ( .A(n8114), .B(n8115), .Z(n8112) );
  XOR U9430 ( .A(n8113), .B(n8028), .Z(n8115) );
  XNOR U9431 ( .A(n8116), .B(n8117), .Z(n8028) );
  ANDN U9432 ( .B(n8118), .A(n8119), .Z(n8116) );
  XOR U9433 ( .A(n8117), .B(n8120), .Z(n8118) );
  XNOR U9434 ( .A(n8113), .B(n8030), .Z(n8114) );
  XOR U9435 ( .A(n8121), .B(n8122), .Z(n8030) );
  AND U9436 ( .A(n102), .B(n8123), .Z(n8121) );
  XOR U9437 ( .A(n8124), .B(n8122), .Z(n8123) );
  XNOR U9438 ( .A(n8125), .B(n8126), .Z(n8113) );
  AND U9439 ( .A(n8127), .B(n8128), .Z(n8125) );
  XNOR U9440 ( .A(n8126), .B(n8055), .Z(n8128) );
  XOR U9441 ( .A(n8119), .B(n8120), .Z(n8055) );
  XNOR U9442 ( .A(n8129), .B(n8130), .Z(n8120) );
  ANDN U9443 ( .B(n8131), .A(n8132), .Z(n8129) );
  XOR U9444 ( .A(n8133), .B(n8134), .Z(n8131) );
  XOR U9445 ( .A(n8135), .B(n8136), .Z(n8119) );
  XNOR U9446 ( .A(n8137), .B(n8138), .Z(n8136) );
  ANDN U9447 ( .B(n8139), .A(n8140), .Z(n8137) );
  XNOR U9448 ( .A(n8141), .B(n8142), .Z(n8139) );
  IV U9449 ( .A(n8117), .Z(n8135) );
  XOR U9450 ( .A(n8143), .B(n8144), .Z(n8117) );
  ANDN U9451 ( .B(n8145), .A(n8146), .Z(n8143) );
  XOR U9452 ( .A(n8144), .B(n8147), .Z(n8145) );
  XOR U9453 ( .A(n8126), .B(n8057), .Z(n8127) );
  XOR U9454 ( .A(n8148), .B(n8149), .Z(n8057) );
  AND U9455 ( .A(n102), .B(n8150), .Z(n8148) );
  XOR U9456 ( .A(n8151), .B(n8149), .Z(n8150) );
  XNOR U9457 ( .A(n8152), .B(n8153), .Z(n8126) );
  NAND U9458 ( .A(n8154), .B(n8155), .Z(n8153) );
  XOR U9459 ( .A(n8156), .B(n8105), .Z(n8155) );
  XOR U9460 ( .A(n8146), .B(n8147), .Z(n8105) );
  XOR U9461 ( .A(n8157), .B(n8134), .Z(n8147) );
  XOR U9462 ( .A(n8158), .B(n8159), .Z(n8134) );
  ANDN U9463 ( .B(n8160), .A(n8161), .Z(n8158) );
  XOR U9464 ( .A(n8159), .B(n8162), .Z(n8160) );
  IV U9465 ( .A(n8132), .Z(n8157) );
  XOR U9466 ( .A(n8130), .B(n8163), .Z(n8132) );
  XOR U9467 ( .A(n8164), .B(n8165), .Z(n8163) );
  ANDN U9468 ( .B(n8166), .A(n8167), .Z(n8164) );
  XOR U9469 ( .A(n8168), .B(n8165), .Z(n8166) );
  IV U9470 ( .A(n8133), .Z(n8130) );
  XOR U9471 ( .A(n8169), .B(n8170), .Z(n8133) );
  ANDN U9472 ( .B(n8171), .A(n8172), .Z(n8169) );
  XOR U9473 ( .A(n8170), .B(n8173), .Z(n8171) );
  XOR U9474 ( .A(n8174), .B(n8175), .Z(n8146) );
  XNOR U9475 ( .A(n8141), .B(n8176), .Z(n8175) );
  IV U9476 ( .A(n8144), .Z(n8176) );
  XOR U9477 ( .A(n8177), .B(n8178), .Z(n8144) );
  ANDN U9478 ( .B(n8179), .A(n8180), .Z(n8177) );
  XOR U9479 ( .A(n8178), .B(n8181), .Z(n8179) );
  XNOR U9480 ( .A(n8182), .B(n8183), .Z(n8141) );
  ANDN U9481 ( .B(n8184), .A(n8185), .Z(n8182) );
  XOR U9482 ( .A(n8183), .B(n8186), .Z(n8184) );
  IV U9483 ( .A(n8140), .Z(n8174) );
  XOR U9484 ( .A(n8138), .B(n8187), .Z(n8140) );
  XOR U9485 ( .A(n8188), .B(n8189), .Z(n8187) );
  ANDN U9486 ( .B(n8190), .A(n8191), .Z(n8188) );
  XOR U9487 ( .A(n8192), .B(n8189), .Z(n8190) );
  IV U9488 ( .A(n8142), .Z(n8138) );
  XOR U9489 ( .A(n8193), .B(n8194), .Z(n8142) );
  ANDN U9490 ( .B(n8195), .A(n8196), .Z(n8193) );
  XOR U9491 ( .A(n8197), .B(n8194), .Z(n8195) );
  IV U9492 ( .A(n8152), .Z(n8156) );
  XOR U9493 ( .A(n8152), .B(n8107), .Z(n8154) );
  XOR U9494 ( .A(n8198), .B(n8199), .Z(n8107) );
  AND U9495 ( .A(n102), .B(n8200), .Z(n8198) );
  XOR U9496 ( .A(n8201), .B(n8199), .Z(n8200) );
  NANDN U9497 ( .A(n8109), .B(n8111), .Z(n8152) );
  XOR U9498 ( .A(n8202), .B(n8203), .Z(n8111) );
  AND U9499 ( .A(n102), .B(n8204), .Z(n8202) );
  XOR U9500 ( .A(n8203), .B(n8205), .Z(n8204) );
  XNOR U9501 ( .A(n8206), .B(n8207), .Z(n102) );
  AND U9502 ( .A(n8208), .B(n8209), .Z(n8206) );
  XOR U9503 ( .A(n8207), .B(n8122), .Z(n8209) );
  XNOR U9504 ( .A(n8210), .B(n8211), .Z(n8122) );
  ANDN U9505 ( .B(n8212), .A(n8213), .Z(n8210) );
  XOR U9506 ( .A(n8211), .B(n8214), .Z(n8212) );
  XNOR U9507 ( .A(n8207), .B(n8124), .Z(n8208) );
  XOR U9508 ( .A(n8215), .B(n8216), .Z(n8124) );
  AND U9509 ( .A(n106), .B(n8217), .Z(n8215) );
  XOR U9510 ( .A(n8218), .B(n8216), .Z(n8217) );
  XNOR U9511 ( .A(n8219), .B(n8220), .Z(n8207) );
  AND U9512 ( .A(n8221), .B(n8222), .Z(n8219) );
  XNOR U9513 ( .A(n8220), .B(n8149), .Z(n8222) );
  XOR U9514 ( .A(n8213), .B(n8214), .Z(n8149) );
  XNOR U9515 ( .A(n8223), .B(n8224), .Z(n8214) );
  ANDN U9516 ( .B(n8225), .A(n8226), .Z(n8223) );
  XOR U9517 ( .A(n8227), .B(n8228), .Z(n8225) );
  XOR U9518 ( .A(n8229), .B(n8230), .Z(n8213) );
  XNOR U9519 ( .A(n8231), .B(n8232), .Z(n8230) );
  ANDN U9520 ( .B(n8233), .A(n8234), .Z(n8231) );
  XNOR U9521 ( .A(n8235), .B(n8236), .Z(n8233) );
  IV U9522 ( .A(n8211), .Z(n8229) );
  XOR U9523 ( .A(n8237), .B(n8238), .Z(n8211) );
  ANDN U9524 ( .B(n8239), .A(n8240), .Z(n8237) );
  XOR U9525 ( .A(n8238), .B(n8241), .Z(n8239) );
  XOR U9526 ( .A(n8220), .B(n8151), .Z(n8221) );
  XOR U9527 ( .A(n8242), .B(n8243), .Z(n8151) );
  AND U9528 ( .A(n106), .B(n8244), .Z(n8242) );
  XOR U9529 ( .A(n8245), .B(n8243), .Z(n8244) );
  XNOR U9530 ( .A(n8246), .B(n8247), .Z(n8220) );
  NAND U9531 ( .A(n8248), .B(n8249), .Z(n8247) );
  XOR U9532 ( .A(n8250), .B(n8199), .Z(n8249) );
  XOR U9533 ( .A(n8240), .B(n8241), .Z(n8199) );
  XOR U9534 ( .A(n8251), .B(n8228), .Z(n8241) );
  XOR U9535 ( .A(n8252), .B(n8253), .Z(n8228) );
  ANDN U9536 ( .B(n8254), .A(n8255), .Z(n8252) );
  XOR U9537 ( .A(n8253), .B(n8256), .Z(n8254) );
  IV U9538 ( .A(n8226), .Z(n8251) );
  XOR U9539 ( .A(n8224), .B(n8257), .Z(n8226) );
  XOR U9540 ( .A(n8258), .B(n8259), .Z(n8257) );
  ANDN U9541 ( .B(n8260), .A(n8261), .Z(n8258) );
  XOR U9542 ( .A(n8262), .B(n8259), .Z(n8260) );
  IV U9543 ( .A(n8227), .Z(n8224) );
  XOR U9544 ( .A(n8263), .B(n8264), .Z(n8227) );
  ANDN U9545 ( .B(n8265), .A(n8266), .Z(n8263) );
  XOR U9546 ( .A(n8264), .B(n8267), .Z(n8265) );
  XOR U9547 ( .A(n8268), .B(n8269), .Z(n8240) );
  XNOR U9548 ( .A(n8235), .B(n8270), .Z(n8269) );
  IV U9549 ( .A(n8238), .Z(n8270) );
  XOR U9550 ( .A(n8271), .B(n8272), .Z(n8238) );
  ANDN U9551 ( .B(n8273), .A(n8274), .Z(n8271) );
  XOR U9552 ( .A(n8272), .B(n8275), .Z(n8273) );
  XNOR U9553 ( .A(n8276), .B(n8277), .Z(n8235) );
  ANDN U9554 ( .B(n8278), .A(n8279), .Z(n8276) );
  XOR U9555 ( .A(n8277), .B(n8280), .Z(n8278) );
  IV U9556 ( .A(n8234), .Z(n8268) );
  XOR U9557 ( .A(n8232), .B(n8281), .Z(n8234) );
  XOR U9558 ( .A(n8282), .B(n8283), .Z(n8281) );
  ANDN U9559 ( .B(n8284), .A(n8285), .Z(n8282) );
  XOR U9560 ( .A(n8286), .B(n8283), .Z(n8284) );
  IV U9561 ( .A(n8236), .Z(n8232) );
  XOR U9562 ( .A(n8287), .B(n8288), .Z(n8236) );
  ANDN U9563 ( .B(n8289), .A(n8290), .Z(n8287) );
  XOR U9564 ( .A(n8291), .B(n8288), .Z(n8289) );
  IV U9565 ( .A(n8246), .Z(n8250) );
  XOR U9566 ( .A(n8246), .B(n8201), .Z(n8248) );
  XOR U9567 ( .A(n8292), .B(n8293), .Z(n8201) );
  AND U9568 ( .A(n106), .B(n8294), .Z(n8292) );
  XOR U9569 ( .A(n8295), .B(n8293), .Z(n8294) );
  NANDN U9570 ( .A(n8203), .B(n8205), .Z(n8246) );
  XOR U9571 ( .A(n8296), .B(n8297), .Z(n8205) );
  AND U9572 ( .A(n106), .B(n8298), .Z(n8296) );
  XOR U9573 ( .A(n8297), .B(n8299), .Z(n8298) );
  XNOR U9574 ( .A(n8300), .B(n8301), .Z(n106) );
  AND U9575 ( .A(n8302), .B(n8303), .Z(n8300) );
  XOR U9576 ( .A(n8301), .B(n8216), .Z(n8303) );
  XNOR U9577 ( .A(n8304), .B(n8305), .Z(n8216) );
  ANDN U9578 ( .B(n8306), .A(n8307), .Z(n8304) );
  XOR U9579 ( .A(n8305), .B(n8308), .Z(n8306) );
  XNOR U9580 ( .A(n8301), .B(n8218), .Z(n8302) );
  XOR U9581 ( .A(n8309), .B(n8310), .Z(n8218) );
  AND U9582 ( .A(n110), .B(n8311), .Z(n8309) );
  XOR U9583 ( .A(n8312), .B(n8310), .Z(n8311) );
  XNOR U9584 ( .A(n8313), .B(n8314), .Z(n8301) );
  AND U9585 ( .A(n8315), .B(n8316), .Z(n8313) );
  XNOR U9586 ( .A(n8314), .B(n8243), .Z(n8316) );
  XOR U9587 ( .A(n8307), .B(n8308), .Z(n8243) );
  XNOR U9588 ( .A(n8317), .B(n8318), .Z(n8308) );
  ANDN U9589 ( .B(n8319), .A(n8320), .Z(n8317) );
  XOR U9590 ( .A(n8321), .B(n8322), .Z(n8319) );
  XOR U9591 ( .A(n8323), .B(n8324), .Z(n8307) );
  XNOR U9592 ( .A(n8325), .B(n8326), .Z(n8324) );
  ANDN U9593 ( .B(n8327), .A(n8328), .Z(n8325) );
  XNOR U9594 ( .A(n8329), .B(n8330), .Z(n8327) );
  IV U9595 ( .A(n8305), .Z(n8323) );
  XOR U9596 ( .A(n8331), .B(n8332), .Z(n8305) );
  ANDN U9597 ( .B(n8333), .A(n8334), .Z(n8331) );
  XOR U9598 ( .A(n8332), .B(n8335), .Z(n8333) );
  XOR U9599 ( .A(n8314), .B(n8245), .Z(n8315) );
  XOR U9600 ( .A(n8336), .B(n8337), .Z(n8245) );
  AND U9601 ( .A(n110), .B(n8338), .Z(n8336) );
  XOR U9602 ( .A(n8339), .B(n8337), .Z(n8338) );
  XNOR U9603 ( .A(n8340), .B(n8341), .Z(n8314) );
  NAND U9604 ( .A(n8342), .B(n8343), .Z(n8341) );
  XOR U9605 ( .A(n8344), .B(n8293), .Z(n8343) );
  XOR U9606 ( .A(n8334), .B(n8335), .Z(n8293) );
  XOR U9607 ( .A(n8345), .B(n8322), .Z(n8335) );
  XOR U9608 ( .A(n8346), .B(n8347), .Z(n8322) );
  ANDN U9609 ( .B(n8348), .A(n8349), .Z(n8346) );
  XOR U9610 ( .A(n8347), .B(n8350), .Z(n8348) );
  IV U9611 ( .A(n8320), .Z(n8345) );
  XOR U9612 ( .A(n8318), .B(n8351), .Z(n8320) );
  XOR U9613 ( .A(n8352), .B(n8353), .Z(n8351) );
  ANDN U9614 ( .B(n8354), .A(n8355), .Z(n8352) );
  XOR U9615 ( .A(n8356), .B(n8353), .Z(n8354) );
  IV U9616 ( .A(n8321), .Z(n8318) );
  XOR U9617 ( .A(n8357), .B(n8358), .Z(n8321) );
  ANDN U9618 ( .B(n8359), .A(n8360), .Z(n8357) );
  XOR U9619 ( .A(n8358), .B(n8361), .Z(n8359) );
  XOR U9620 ( .A(n8362), .B(n8363), .Z(n8334) );
  XNOR U9621 ( .A(n8329), .B(n8364), .Z(n8363) );
  IV U9622 ( .A(n8332), .Z(n8364) );
  XOR U9623 ( .A(n8365), .B(n8366), .Z(n8332) );
  ANDN U9624 ( .B(n8367), .A(n8368), .Z(n8365) );
  XOR U9625 ( .A(n8366), .B(n8369), .Z(n8367) );
  XNOR U9626 ( .A(n8370), .B(n8371), .Z(n8329) );
  ANDN U9627 ( .B(n8372), .A(n8373), .Z(n8370) );
  XOR U9628 ( .A(n8371), .B(n8374), .Z(n8372) );
  IV U9629 ( .A(n8328), .Z(n8362) );
  XOR U9630 ( .A(n8326), .B(n8375), .Z(n8328) );
  XOR U9631 ( .A(n8376), .B(n8377), .Z(n8375) );
  ANDN U9632 ( .B(n8378), .A(n8379), .Z(n8376) );
  XOR U9633 ( .A(n8380), .B(n8377), .Z(n8378) );
  IV U9634 ( .A(n8330), .Z(n8326) );
  XOR U9635 ( .A(n8381), .B(n8382), .Z(n8330) );
  ANDN U9636 ( .B(n8383), .A(n8384), .Z(n8381) );
  XOR U9637 ( .A(n8385), .B(n8382), .Z(n8383) );
  IV U9638 ( .A(n8340), .Z(n8344) );
  XOR U9639 ( .A(n8340), .B(n8295), .Z(n8342) );
  XOR U9640 ( .A(n8386), .B(n8387), .Z(n8295) );
  AND U9641 ( .A(n110), .B(n8388), .Z(n8386) );
  XOR U9642 ( .A(n8389), .B(n8387), .Z(n8388) );
  NANDN U9643 ( .A(n8297), .B(n8299), .Z(n8340) );
  XOR U9644 ( .A(n8390), .B(n8391), .Z(n8299) );
  AND U9645 ( .A(n110), .B(n8392), .Z(n8390) );
  XOR U9646 ( .A(n8391), .B(n8393), .Z(n8392) );
  XNOR U9647 ( .A(n8394), .B(n8395), .Z(n110) );
  AND U9648 ( .A(n8396), .B(n8397), .Z(n8394) );
  XOR U9649 ( .A(n8395), .B(n8310), .Z(n8397) );
  XNOR U9650 ( .A(n8398), .B(n8399), .Z(n8310) );
  ANDN U9651 ( .B(n8400), .A(n8401), .Z(n8398) );
  XOR U9652 ( .A(n8399), .B(n8402), .Z(n8400) );
  XNOR U9653 ( .A(n8395), .B(n8312), .Z(n8396) );
  XOR U9654 ( .A(n8403), .B(n8404), .Z(n8312) );
  AND U9655 ( .A(n114), .B(n8405), .Z(n8403) );
  XOR U9656 ( .A(n8406), .B(n8404), .Z(n8405) );
  XNOR U9657 ( .A(n8407), .B(n8408), .Z(n8395) );
  AND U9658 ( .A(n8409), .B(n8410), .Z(n8407) );
  XNOR U9659 ( .A(n8408), .B(n8337), .Z(n8410) );
  XOR U9660 ( .A(n8401), .B(n8402), .Z(n8337) );
  XNOR U9661 ( .A(n8411), .B(n8412), .Z(n8402) );
  ANDN U9662 ( .B(n8413), .A(n8414), .Z(n8411) );
  XOR U9663 ( .A(n8415), .B(n8416), .Z(n8413) );
  XOR U9664 ( .A(n8417), .B(n8418), .Z(n8401) );
  XNOR U9665 ( .A(n8419), .B(n8420), .Z(n8418) );
  ANDN U9666 ( .B(n8421), .A(n8422), .Z(n8419) );
  XNOR U9667 ( .A(n8423), .B(n8424), .Z(n8421) );
  IV U9668 ( .A(n8399), .Z(n8417) );
  XOR U9669 ( .A(n8425), .B(n8426), .Z(n8399) );
  ANDN U9670 ( .B(n8427), .A(n8428), .Z(n8425) );
  XOR U9671 ( .A(n8426), .B(n8429), .Z(n8427) );
  XOR U9672 ( .A(n8408), .B(n8339), .Z(n8409) );
  XOR U9673 ( .A(n8430), .B(n8431), .Z(n8339) );
  AND U9674 ( .A(n114), .B(n8432), .Z(n8430) );
  XOR U9675 ( .A(n8433), .B(n8431), .Z(n8432) );
  XNOR U9676 ( .A(n8434), .B(n8435), .Z(n8408) );
  NAND U9677 ( .A(n8436), .B(n8437), .Z(n8435) );
  XOR U9678 ( .A(n8438), .B(n8387), .Z(n8437) );
  XOR U9679 ( .A(n8428), .B(n8429), .Z(n8387) );
  XOR U9680 ( .A(n8439), .B(n8416), .Z(n8429) );
  XOR U9681 ( .A(n8440), .B(n8441), .Z(n8416) );
  ANDN U9682 ( .B(n8442), .A(n8443), .Z(n8440) );
  XOR U9683 ( .A(n8441), .B(n8444), .Z(n8442) );
  IV U9684 ( .A(n8414), .Z(n8439) );
  XOR U9685 ( .A(n8412), .B(n8445), .Z(n8414) );
  XOR U9686 ( .A(n8446), .B(n8447), .Z(n8445) );
  ANDN U9687 ( .B(n8448), .A(n8449), .Z(n8446) );
  XOR U9688 ( .A(n8450), .B(n8447), .Z(n8448) );
  IV U9689 ( .A(n8415), .Z(n8412) );
  XOR U9690 ( .A(n8451), .B(n8452), .Z(n8415) );
  ANDN U9691 ( .B(n8453), .A(n8454), .Z(n8451) );
  XOR U9692 ( .A(n8452), .B(n8455), .Z(n8453) );
  XOR U9693 ( .A(n8456), .B(n8457), .Z(n8428) );
  XNOR U9694 ( .A(n8423), .B(n8458), .Z(n8457) );
  IV U9695 ( .A(n8426), .Z(n8458) );
  XOR U9696 ( .A(n8459), .B(n8460), .Z(n8426) );
  ANDN U9697 ( .B(n8461), .A(n8462), .Z(n8459) );
  XOR U9698 ( .A(n8460), .B(n8463), .Z(n8461) );
  XNOR U9699 ( .A(n8464), .B(n8465), .Z(n8423) );
  ANDN U9700 ( .B(n8466), .A(n8467), .Z(n8464) );
  XOR U9701 ( .A(n8465), .B(n8468), .Z(n8466) );
  IV U9702 ( .A(n8422), .Z(n8456) );
  XOR U9703 ( .A(n8420), .B(n8469), .Z(n8422) );
  XOR U9704 ( .A(n8470), .B(n8471), .Z(n8469) );
  ANDN U9705 ( .B(n8472), .A(n8473), .Z(n8470) );
  XOR U9706 ( .A(n8474), .B(n8471), .Z(n8472) );
  IV U9707 ( .A(n8424), .Z(n8420) );
  XOR U9708 ( .A(n8475), .B(n8476), .Z(n8424) );
  ANDN U9709 ( .B(n8477), .A(n8478), .Z(n8475) );
  XOR U9710 ( .A(n8479), .B(n8476), .Z(n8477) );
  IV U9711 ( .A(n8434), .Z(n8438) );
  XOR U9712 ( .A(n8434), .B(n8389), .Z(n8436) );
  XOR U9713 ( .A(n8480), .B(n8481), .Z(n8389) );
  AND U9714 ( .A(n114), .B(n8482), .Z(n8480) );
  XOR U9715 ( .A(n8483), .B(n8481), .Z(n8482) );
  NANDN U9716 ( .A(n8391), .B(n8393), .Z(n8434) );
  XOR U9717 ( .A(n8484), .B(n8485), .Z(n8393) );
  AND U9718 ( .A(n114), .B(n8486), .Z(n8484) );
  XOR U9719 ( .A(n8485), .B(n8487), .Z(n8486) );
  XNOR U9720 ( .A(n8488), .B(n8489), .Z(n114) );
  AND U9721 ( .A(n8490), .B(n8491), .Z(n8488) );
  XOR U9722 ( .A(n8489), .B(n8404), .Z(n8491) );
  XNOR U9723 ( .A(n8492), .B(n8493), .Z(n8404) );
  ANDN U9724 ( .B(n8494), .A(n8495), .Z(n8492) );
  XOR U9725 ( .A(n8493), .B(n8496), .Z(n8494) );
  XNOR U9726 ( .A(n8489), .B(n8406), .Z(n8490) );
  XOR U9727 ( .A(n8497), .B(n8498), .Z(n8406) );
  AND U9728 ( .A(n118), .B(n8499), .Z(n8497) );
  XOR U9729 ( .A(n8500), .B(n8498), .Z(n8499) );
  XNOR U9730 ( .A(n8501), .B(n8502), .Z(n8489) );
  AND U9731 ( .A(n8503), .B(n8504), .Z(n8501) );
  XNOR U9732 ( .A(n8502), .B(n8431), .Z(n8504) );
  XOR U9733 ( .A(n8495), .B(n8496), .Z(n8431) );
  XNOR U9734 ( .A(n8505), .B(n8506), .Z(n8496) );
  ANDN U9735 ( .B(n8507), .A(n8508), .Z(n8505) );
  XOR U9736 ( .A(n8509), .B(n8510), .Z(n8507) );
  XOR U9737 ( .A(n8511), .B(n8512), .Z(n8495) );
  XNOR U9738 ( .A(n8513), .B(n8514), .Z(n8512) );
  ANDN U9739 ( .B(n8515), .A(n8516), .Z(n8513) );
  XNOR U9740 ( .A(n8517), .B(n8518), .Z(n8515) );
  IV U9741 ( .A(n8493), .Z(n8511) );
  XOR U9742 ( .A(n8519), .B(n8520), .Z(n8493) );
  ANDN U9743 ( .B(n8521), .A(n8522), .Z(n8519) );
  XOR U9744 ( .A(n8520), .B(n8523), .Z(n8521) );
  XOR U9745 ( .A(n8502), .B(n8433), .Z(n8503) );
  XOR U9746 ( .A(n8524), .B(n8525), .Z(n8433) );
  AND U9747 ( .A(n118), .B(n8526), .Z(n8524) );
  XOR U9748 ( .A(n8527), .B(n8525), .Z(n8526) );
  XNOR U9749 ( .A(n8528), .B(n8529), .Z(n8502) );
  NAND U9750 ( .A(n8530), .B(n8531), .Z(n8529) );
  XOR U9751 ( .A(n8532), .B(n8481), .Z(n8531) );
  XOR U9752 ( .A(n8522), .B(n8523), .Z(n8481) );
  XOR U9753 ( .A(n8533), .B(n8510), .Z(n8523) );
  XOR U9754 ( .A(n8534), .B(n8535), .Z(n8510) );
  ANDN U9755 ( .B(n8536), .A(n8537), .Z(n8534) );
  XOR U9756 ( .A(n8535), .B(n8538), .Z(n8536) );
  IV U9757 ( .A(n8508), .Z(n8533) );
  XOR U9758 ( .A(n8506), .B(n8539), .Z(n8508) );
  XOR U9759 ( .A(n8540), .B(n8541), .Z(n8539) );
  ANDN U9760 ( .B(n8542), .A(n8543), .Z(n8540) );
  XOR U9761 ( .A(n8544), .B(n8541), .Z(n8542) );
  IV U9762 ( .A(n8509), .Z(n8506) );
  XOR U9763 ( .A(n8545), .B(n8546), .Z(n8509) );
  ANDN U9764 ( .B(n8547), .A(n8548), .Z(n8545) );
  XOR U9765 ( .A(n8546), .B(n8549), .Z(n8547) );
  XOR U9766 ( .A(n8550), .B(n8551), .Z(n8522) );
  XNOR U9767 ( .A(n8517), .B(n8552), .Z(n8551) );
  IV U9768 ( .A(n8520), .Z(n8552) );
  XOR U9769 ( .A(n8553), .B(n8554), .Z(n8520) );
  ANDN U9770 ( .B(n8555), .A(n8556), .Z(n8553) );
  XOR U9771 ( .A(n8554), .B(n8557), .Z(n8555) );
  XNOR U9772 ( .A(n8558), .B(n8559), .Z(n8517) );
  ANDN U9773 ( .B(n8560), .A(n8561), .Z(n8558) );
  XOR U9774 ( .A(n8559), .B(n8562), .Z(n8560) );
  IV U9775 ( .A(n8516), .Z(n8550) );
  XOR U9776 ( .A(n8514), .B(n8563), .Z(n8516) );
  XOR U9777 ( .A(n8564), .B(n8565), .Z(n8563) );
  ANDN U9778 ( .B(n8566), .A(n8567), .Z(n8564) );
  XOR U9779 ( .A(n8568), .B(n8565), .Z(n8566) );
  IV U9780 ( .A(n8518), .Z(n8514) );
  XOR U9781 ( .A(n8569), .B(n8570), .Z(n8518) );
  ANDN U9782 ( .B(n8571), .A(n8572), .Z(n8569) );
  XOR U9783 ( .A(n8573), .B(n8570), .Z(n8571) );
  IV U9784 ( .A(n8528), .Z(n8532) );
  XOR U9785 ( .A(n8528), .B(n8483), .Z(n8530) );
  XOR U9786 ( .A(n8574), .B(n8575), .Z(n8483) );
  AND U9787 ( .A(n118), .B(n8576), .Z(n8574) );
  XOR U9788 ( .A(n8577), .B(n8575), .Z(n8576) );
  NANDN U9789 ( .A(n8485), .B(n8487), .Z(n8528) );
  XOR U9790 ( .A(n8578), .B(n8579), .Z(n8487) );
  AND U9791 ( .A(n118), .B(n8580), .Z(n8578) );
  XOR U9792 ( .A(n8579), .B(n8581), .Z(n8580) );
  XNOR U9793 ( .A(n8582), .B(n8583), .Z(n118) );
  AND U9794 ( .A(n8584), .B(n8585), .Z(n8582) );
  XOR U9795 ( .A(n8583), .B(n8498), .Z(n8585) );
  XNOR U9796 ( .A(n8586), .B(n8587), .Z(n8498) );
  ANDN U9797 ( .B(n8588), .A(n8589), .Z(n8586) );
  XOR U9798 ( .A(n8587), .B(n8590), .Z(n8588) );
  XNOR U9799 ( .A(n8583), .B(n8500), .Z(n8584) );
  XOR U9800 ( .A(n8591), .B(n8592), .Z(n8500) );
  AND U9801 ( .A(n122), .B(n8593), .Z(n8591) );
  XOR U9802 ( .A(n8594), .B(n8592), .Z(n8593) );
  XNOR U9803 ( .A(n8595), .B(n8596), .Z(n8583) );
  AND U9804 ( .A(n8597), .B(n8598), .Z(n8595) );
  XNOR U9805 ( .A(n8596), .B(n8525), .Z(n8598) );
  XOR U9806 ( .A(n8589), .B(n8590), .Z(n8525) );
  XNOR U9807 ( .A(n8599), .B(n8600), .Z(n8590) );
  ANDN U9808 ( .B(n8601), .A(n8602), .Z(n8599) );
  XOR U9809 ( .A(n8603), .B(n8604), .Z(n8601) );
  XOR U9810 ( .A(n8605), .B(n8606), .Z(n8589) );
  XNOR U9811 ( .A(n8607), .B(n8608), .Z(n8606) );
  ANDN U9812 ( .B(n8609), .A(n8610), .Z(n8607) );
  XNOR U9813 ( .A(n8611), .B(n8612), .Z(n8609) );
  IV U9814 ( .A(n8587), .Z(n8605) );
  XOR U9815 ( .A(n8613), .B(n8614), .Z(n8587) );
  ANDN U9816 ( .B(n8615), .A(n8616), .Z(n8613) );
  XOR U9817 ( .A(n8614), .B(n8617), .Z(n8615) );
  XOR U9818 ( .A(n8596), .B(n8527), .Z(n8597) );
  XOR U9819 ( .A(n8618), .B(n8619), .Z(n8527) );
  AND U9820 ( .A(n122), .B(n8620), .Z(n8618) );
  XOR U9821 ( .A(n8621), .B(n8619), .Z(n8620) );
  XNOR U9822 ( .A(n8622), .B(n8623), .Z(n8596) );
  NAND U9823 ( .A(n8624), .B(n8625), .Z(n8623) );
  XOR U9824 ( .A(n8626), .B(n8575), .Z(n8625) );
  XOR U9825 ( .A(n8616), .B(n8617), .Z(n8575) );
  XOR U9826 ( .A(n8627), .B(n8604), .Z(n8617) );
  XOR U9827 ( .A(n8628), .B(n8629), .Z(n8604) );
  ANDN U9828 ( .B(n8630), .A(n8631), .Z(n8628) );
  XOR U9829 ( .A(n8629), .B(n8632), .Z(n8630) );
  IV U9830 ( .A(n8602), .Z(n8627) );
  XOR U9831 ( .A(n8600), .B(n8633), .Z(n8602) );
  XOR U9832 ( .A(n8634), .B(n8635), .Z(n8633) );
  ANDN U9833 ( .B(n8636), .A(n8637), .Z(n8634) );
  XOR U9834 ( .A(n8638), .B(n8635), .Z(n8636) );
  IV U9835 ( .A(n8603), .Z(n8600) );
  XOR U9836 ( .A(n8639), .B(n8640), .Z(n8603) );
  ANDN U9837 ( .B(n8641), .A(n8642), .Z(n8639) );
  XOR U9838 ( .A(n8640), .B(n8643), .Z(n8641) );
  XOR U9839 ( .A(n8644), .B(n8645), .Z(n8616) );
  XNOR U9840 ( .A(n8611), .B(n8646), .Z(n8645) );
  IV U9841 ( .A(n8614), .Z(n8646) );
  XOR U9842 ( .A(n8647), .B(n8648), .Z(n8614) );
  ANDN U9843 ( .B(n8649), .A(n8650), .Z(n8647) );
  XOR U9844 ( .A(n8648), .B(n8651), .Z(n8649) );
  XNOR U9845 ( .A(n8652), .B(n8653), .Z(n8611) );
  ANDN U9846 ( .B(n8654), .A(n8655), .Z(n8652) );
  XOR U9847 ( .A(n8653), .B(n8656), .Z(n8654) );
  IV U9848 ( .A(n8610), .Z(n8644) );
  XOR U9849 ( .A(n8608), .B(n8657), .Z(n8610) );
  XOR U9850 ( .A(n8658), .B(n8659), .Z(n8657) );
  ANDN U9851 ( .B(n8660), .A(n8661), .Z(n8658) );
  XOR U9852 ( .A(n8662), .B(n8659), .Z(n8660) );
  IV U9853 ( .A(n8612), .Z(n8608) );
  XOR U9854 ( .A(n8663), .B(n8664), .Z(n8612) );
  ANDN U9855 ( .B(n8665), .A(n8666), .Z(n8663) );
  XOR U9856 ( .A(n8667), .B(n8664), .Z(n8665) );
  IV U9857 ( .A(n8622), .Z(n8626) );
  XOR U9858 ( .A(n8622), .B(n8577), .Z(n8624) );
  XOR U9859 ( .A(n8668), .B(n8669), .Z(n8577) );
  AND U9860 ( .A(n122), .B(n8670), .Z(n8668) );
  XOR U9861 ( .A(n8671), .B(n8669), .Z(n8670) );
  NANDN U9862 ( .A(n8579), .B(n8581), .Z(n8622) );
  XOR U9863 ( .A(n8672), .B(n8673), .Z(n8581) );
  AND U9864 ( .A(n122), .B(n8674), .Z(n8672) );
  XOR U9865 ( .A(n8673), .B(n8675), .Z(n8674) );
  XNOR U9866 ( .A(n8676), .B(n8677), .Z(n122) );
  AND U9867 ( .A(n8678), .B(n8679), .Z(n8676) );
  XOR U9868 ( .A(n8677), .B(n8592), .Z(n8679) );
  XNOR U9869 ( .A(n8680), .B(n8681), .Z(n8592) );
  ANDN U9870 ( .B(n8682), .A(n8683), .Z(n8680) );
  XOR U9871 ( .A(n8681), .B(n8684), .Z(n8682) );
  XNOR U9872 ( .A(n8677), .B(n8594), .Z(n8678) );
  XOR U9873 ( .A(n8685), .B(n8686), .Z(n8594) );
  AND U9874 ( .A(n126), .B(n8687), .Z(n8685) );
  XOR U9875 ( .A(n8688), .B(n8686), .Z(n8687) );
  XNOR U9876 ( .A(n8689), .B(n8690), .Z(n8677) );
  AND U9877 ( .A(n8691), .B(n8692), .Z(n8689) );
  XNOR U9878 ( .A(n8690), .B(n8619), .Z(n8692) );
  XOR U9879 ( .A(n8683), .B(n8684), .Z(n8619) );
  XNOR U9880 ( .A(n8693), .B(n8694), .Z(n8684) );
  ANDN U9881 ( .B(n8695), .A(n8696), .Z(n8693) );
  XOR U9882 ( .A(n8697), .B(n8698), .Z(n8695) );
  XOR U9883 ( .A(n8699), .B(n8700), .Z(n8683) );
  XNOR U9884 ( .A(n8701), .B(n8702), .Z(n8700) );
  ANDN U9885 ( .B(n8703), .A(n8704), .Z(n8701) );
  XNOR U9886 ( .A(n8705), .B(n8706), .Z(n8703) );
  IV U9887 ( .A(n8681), .Z(n8699) );
  XOR U9888 ( .A(n8707), .B(n8708), .Z(n8681) );
  ANDN U9889 ( .B(n8709), .A(n8710), .Z(n8707) );
  XOR U9890 ( .A(n8708), .B(n8711), .Z(n8709) );
  XOR U9891 ( .A(n8690), .B(n8621), .Z(n8691) );
  XOR U9892 ( .A(n8712), .B(n8713), .Z(n8621) );
  AND U9893 ( .A(n126), .B(n8714), .Z(n8712) );
  XOR U9894 ( .A(n8715), .B(n8713), .Z(n8714) );
  XNOR U9895 ( .A(n8716), .B(n8717), .Z(n8690) );
  NAND U9896 ( .A(n8718), .B(n8719), .Z(n8717) );
  XOR U9897 ( .A(n8720), .B(n8669), .Z(n8719) );
  XOR U9898 ( .A(n8710), .B(n8711), .Z(n8669) );
  XOR U9899 ( .A(n8721), .B(n8698), .Z(n8711) );
  XOR U9900 ( .A(n8722), .B(n8723), .Z(n8698) );
  ANDN U9901 ( .B(n8724), .A(n8725), .Z(n8722) );
  XOR U9902 ( .A(n8723), .B(n8726), .Z(n8724) );
  IV U9903 ( .A(n8696), .Z(n8721) );
  XOR U9904 ( .A(n8694), .B(n8727), .Z(n8696) );
  XOR U9905 ( .A(n8728), .B(n8729), .Z(n8727) );
  ANDN U9906 ( .B(n8730), .A(n8731), .Z(n8728) );
  XOR U9907 ( .A(n8732), .B(n8729), .Z(n8730) );
  IV U9908 ( .A(n8697), .Z(n8694) );
  XOR U9909 ( .A(n8733), .B(n8734), .Z(n8697) );
  ANDN U9910 ( .B(n8735), .A(n8736), .Z(n8733) );
  XOR U9911 ( .A(n8734), .B(n8737), .Z(n8735) );
  XOR U9912 ( .A(n8738), .B(n8739), .Z(n8710) );
  XNOR U9913 ( .A(n8705), .B(n8740), .Z(n8739) );
  IV U9914 ( .A(n8708), .Z(n8740) );
  XOR U9915 ( .A(n8741), .B(n8742), .Z(n8708) );
  ANDN U9916 ( .B(n8743), .A(n8744), .Z(n8741) );
  XOR U9917 ( .A(n8742), .B(n8745), .Z(n8743) );
  XNOR U9918 ( .A(n8746), .B(n8747), .Z(n8705) );
  ANDN U9919 ( .B(n8748), .A(n8749), .Z(n8746) );
  XOR U9920 ( .A(n8747), .B(n8750), .Z(n8748) );
  IV U9921 ( .A(n8704), .Z(n8738) );
  XOR U9922 ( .A(n8702), .B(n8751), .Z(n8704) );
  XOR U9923 ( .A(n8752), .B(n8753), .Z(n8751) );
  ANDN U9924 ( .B(n8754), .A(n8755), .Z(n8752) );
  XOR U9925 ( .A(n8756), .B(n8753), .Z(n8754) );
  IV U9926 ( .A(n8706), .Z(n8702) );
  XOR U9927 ( .A(n8757), .B(n8758), .Z(n8706) );
  ANDN U9928 ( .B(n8759), .A(n8760), .Z(n8757) );
  XOR U9929 ( .A(n8761), .B(n8758), .Z(n8759) );
  IV U9930 ( .A(n8716), .Z(n8720) );
  XOR U9931 ( .A(n8716), .B(n8671), .Z(n8718) );
  XOR U9932 ( .A(n8762), .B(n8763), .Z(n8671) );
  AND U9933 ( .A(n126), .B(n8764), .Z(n8762) );
  XOR U9934 ( .A(n8765), .B(n8763), .Z(n8764) );
  NANDN U9935 ( .A(n8673), .B(n8675), .Z(n8716) );
  XOR U9936 ( .A(n8766), .B(n8767), .Z(n8675) );
  AND U9937 ( .A(n126), .B(n8768), .Z(n8766) );
  XOR U9938 ( .A(n8767), .B(n8769), .Z(n8768) );
  XNOR U9939 ( .A(n8770), .B(n8771), .Z(n126) );
  AND U9940 ( .A(n8772), .B(n8773), .Z(n8770) );
  XOR U9941 ( .A(n8771), .B(n8686), .Z(n8773) );
  XNOR U9942 ( .A(n8774), .B(n8775), .Z(n8686) );
  ANDN U9943 ( .B(n8776), .A(n8777), .Z(n8774) );
  XOR U9944 ( .A(n8775), .B(n8778), .Z(n8776) );
  XNOR U9945 ( .A(n8771), .B(n8688), .Z(n8772) );
  XOR U9946 ( .A(n8779), .B(n8780), .Z(n8688) );
  AND U9947 ( .A(n130), .B(n8781), .Z(n8779) );
  XOR U9948 ( .A(n8782), .B(n8780), .Z(n8781) );
  XNOR U9949 ( .A(n8783), .B(n8784), .Z(n8771) );
  AND U9950 ( .A(n8785), .B(n8786), .Z(n8783) );
  XNOR U9951 ( .A(n8784), .B(n8713), .Z(n8786) );
  XOR U9952 ( .A(n8777), .B(n8778), .Z(n8713) );
  XNOR U9953 ( .A(n8787), .B(n8788), .Z(n8778) );
  ANDN U9954 ( .B(n8789), .A(n8790), .Z(n8787) );
  XOR U9955 ( .A(n8791), .B(n8792), .Z(n8789) );
  XOR U9956 ( .A(n8793), .B(n8794), .Z(n8777) );
  XNOR U9957 ( .A(n8795), .B(n8796), .Z(n8794) );
  ANDN U9958 ( .B(n8797), .A(n8798), .Z(n8795) );
  XNOR U9959 ( .A(n8799), .B(n8800), .Z(n8797) );
  IV U9960 ( .A(n8775), .Z(n8793) );
  XOR U9961 ( .A(n8801), .B(n8802), .Z(n8775) );
  ANDN U9962 ( .B(n8803), .A(n8804), .Z(n8801) );
  XOR U9963 ( .A(n8802), .B(n8805), .Z(n8803) );
  XOR U9964 ( .A(n8784), .B(n8715), .Z(n8785) );
  XOR U9965 ( .A(n8806), .B(n8807), .Z(n8715) );
  AND U9966 ( .A(n130), .B(n8808), .Z(n8806) );
  XOR U9967 ( .A(n8809), .B(n8807), .Z(n8808) );
  XNOR U9968 ( .A(n8810), .B(n8811), .Z(n8784) );
  NAND U9969 ( .A(n8812), .B(n8813), .Z(n8811) );
  XOR U9970 ( .A(n8814), .B(n8763), .Z(n8813) );
  XOR U9971 ( .A(n8804), .B(n8805), .Z(n8763) );
  XOR U9972 ( .A(n8815), .B(n8792), .Z(n8805) );
  XOR U9973 ( .A(n8816), .B(n8817), .Z(n8792) );
  ANDN U9974 ( .B(n8818), .A(n8819), .Z(n8816) );
  XOR U9975 ( .A(n8817), .B(n8820), .Z(n8818) );
  IV U9976 ( .A(n8790), .Z(n8815) );
  XOR U9977 ( .A(n8788), .B(n8821), .Z(n8790) );
  XOR U9978 ( .A(n8822), .B(n8823), .Z(n8821) );
  ANDN U9979 ( .B(n8824), .A(n8825), .Z(n8822) );
  XOR U9980 ( .A(n8826), .B(n8823), .Z(n8824) );
  IV U9981 ( .A(n8791), .Z(n8788) );
  XOR U9982 ( .A(n8827), .B(n8828), .Z(n8791) );
  ANDN U9983 ( .B(n8829), .A(n8830), .Z(n8827) );
  XOR U9984 ( .A(n8828), .B(n8831), .Z(n8829) );
  XOR U9985 ( .A(n8832), .B(n8833), .Z(n8804) );
  XNOR U9986 ( .A(n8799), .B(n8834), .Z(n8833) );
  IV U9987 ( .A(n8802), .Z(n8834) );
  XOR U9988 ( .A(n8835), .B(n8836), .Z(n8802) );
  ANDN U9989 ( .B(n8837), .A(n8838), .Z(n8835) );
  XOR U9990 ( .A(n8836), .B(n8839), .Z(n8837) );
  XNOR U9991 ( .A(n8840), .B(n8841), .Z(n8799) );
  ANDN U9992 ( .B(n8842), .A(n8843), .Z(n8840) );
  XOR U9993 ( .A(n8841), .B(n8844), .Z(n8842) );
  IV U9994 ( .A(n8798), .Z(n8832) );
  XOR U9995 ( .A(n8796), .B(n8845), .Z(n8798) );
  XOR U9996 ( .A(n8846), .B(n8847), .Z(n8845) );
  ANDN U9997 ( .B(n8848), .A(n8849), .Z(n8846) );
  XOR U9998 ( .A(n8850), .B(n8847), .Z(n8848) );
  IV U9999 ( .A(n8800), .Z(n8796) );
  XOR U10000 ( .A(n8851), .B(n8852), .Z(n8800) );
  ANDN U10001 ( .B(n8853), .A(n8854), .Z(n8851) );
  XOR U10002 ( .A(n8855), .B(n8852), .Z(n8853) );
  IV U10003 ( .A(n8810), .Z(n8814) );
  XOR U10004 ( .A(n8810), .B(n8765), .Z(n8812) );
  XOR U10005 ( .A(n8856), .B(n8857), .Z(n8765) );
  AND U10006 ( .A(n130), .B(n8858), .Z(n8856) );
  XOR U10007 ( .A(n8859), .B(n8857), .Z(n8858) );
  NANDN U10008 ( .A(n8767), .B(n8769), .Z(n8810) );
  XOR U10009 ( .A(n8860), .B(n8861), .Z(n8769) );
  AND U10010 ( .A(n130), .B(n8862), .Z(n8860) );
  XOR U10011 ( .A(n8861), .B(n8863), .Z(n8862) );
  XNOR U10012 ( .A(n8864), .B(n8865), .Z(n130) );
  AND U10013 ( .A(n8866), .B(n8867), .Z(n8864) );
  XOR U10014 ( .A(n8865), .B(n8780), .Z(n8867) );
  XNOR U10015 ( .A(n8868), .B(n8869), .Z(n8780) );
  ANDN U10016 ( .B(n8870), .A(n8871), .Z(n8868) );
  XOR U10017 ( .A(n8869), .B(n8872), .Z(n8870) );
  XNOR U10018 ( .A(n8865), .B(n8782), .Z(n8866) );
  XOR U10019 ( .A(n8873), .B(n8874), .Z(n8782) );
  AND U10020 ( .A(n134), .B(n8875), .Z(n8873) );
  XOR U10021 ( .A(n8876), .B(n8874), .Z(n8875) );
  XNOR U10022 ( .A(n8877), .B(n8878), .Z(n8865) );
  AND U10023 ( .A(n8879), .B(n8880), .Z(n8877) );
  XNOR U10024 ( .A(n8878), .B(n8807), .Z(n8880) );
  XOR U10025 ( .A(n8871), .B(n8872), .Z(n8807) );
  XNOR U10026 ( .A(n8881), .B(n8882), .Z(n8872) );
  ANDN U10027 ( .B(n8883), .A(n8884), .Z(n8881) );
  XOR U10028 ( .A(n8885), .B(n8886), .Z(n8883) );
  XOR U10029 ( .A(n8887), .B(n8888), .Z(n8871) );
  XNOR U10030 ( .A(n8889), .B(n8890), .Z(n8888) );
  ANDN U10031 ( .B(n8891), .A(n8892), .Z(n8889) );
  XNOR U10032 ( .A(n8893), .B(n8894), .Z(n8891) );
  IV U10033 ( .A(n8869), .Z(n8887) );
  XOR U10034 ( .A(n8895), .B(n8896), .Z(n8869) );
  ANDN U10035 ( .B(n8897), .A(n8898), .Z(n8895) );
  XOR U10036 ( .A(n8896), .B(n8899), .Z(n8897) );
  XOR U10037 ( .A(n8878), .B(n8809), .Z(n8879) );
  XOR U10038 ( .A(n8900), .B(n8901), .Z(n8809) );
  AND U10039 ( .A(n134), .B(n8902), .Z(n8900) );
  XOR U10040 ( .A(n8903), .B(n8901), .Z(n8902) );
  XNOR U10041 ( .A(n8904), .B(n8905), .Z(n8878) );
  NAND U10042 ( .A(n8906), .B(n8907), .Z(n8905) );
  XOR U10043 ( .A(n8908), .B(n8857), .Z(n8907) );
  XOR U10044 ( .A(n8898), .B(n8899), .Z(n8857) );
  XOR U10045 ( .A(n8909), .B(n8886), .Z(n8899) );
  XOR U10046 ( .A(n8910), .B(n8911), .Z(n8886) );
  ANDN U10047 ( .B(n8912), .A(n8913), .Z(n8910) );
  XOR U10048 ( .A(n8911), .B(n8914), .Z(n8912) );
  IV U10049 ( .A(n8884), .Z(n8909) );
  XOR U10050 ( .A(n8882), .B(n8915), .Z(n8884) );
  XOR U10051 ( .A(n8916), .B(n8917), .Z(n8915) );
  ANDN U10052 ( .B(n8918), .A(n8919), .Z(n8916) );
  XOR U10053 ( .A(n8920), .B(n8917), .Z(n8918) );
  IV U10054 ( .A(n8885), .Z(n8882) );
  XOR U10055 ( .A(n8921), .B(n8922), .Z(n8885) );
  ANDN U10056 ( .B(n8923), .A(n8924), .Z(n8921) );
  XOR U10057 ( .A(n8922), .B(n8925), .Z(n8923) );
  XOR U10058 ( .A(n8926), .B(n8927), .Z(n8898) );
  XNOR U10059 ( .A(n8893), .B(n8928), .Z(n8927) );
  IV U10060 ( .A(n8896), .Z(n8928) );
  XOR U10061 ( .A(n8929), .B(n8930), .Z(n8896) );
  ANDN U10062 ( .B(n8931), .A(n8932), .Z(n8929) );
  XOR U10063 ( .A(n8930), .B(n8933), .Z(n8931) );
  XNOR U10064 ( .A(n8934), .B(n8935), .Z(n8893) );
  ANDN U10065 ( .B(n8936), .A(n8937), .Z(n8934) );
  XOR U10066 ( .A(n8935), .B(n8938), .Z(n8936) );
  IV U10067 ( .A(n8892), .Z(n8926) );
  XOR U10068 ( .A(n8890), .B(n8939), .Z(n8892) );
  XOR U10069 ( .A(n8940), .B(n8941), .Z(n8939) );
  ANDN U10070 ( .B(n8942), .A(n8943), .Z(n8940) );
  XOR U10071 ( .A(n8944), .B(n8941), .Z(n8942) );
  IV U10072 ( .A(n8894), .Z(n8890) );
  XOR U10073 ( .A(n8945), .B(n8946), .Z(n8894) );
  ANDN U10074 ( .B(n8947), .A(n8948), .Z(n8945) );
  XOR U10075 ( .A(n8949), .B(n8946), .Z(n8947) );
  IV U10076 ( .A(n8904), .Z(n8908) );
  XOR U10077 ( .A(n8904), .B(n8859), .Z(n8906) );
  XOR U10078 ( .A(n8950), .B(n8951), .Z(n8859) );
  AND U10079 ( .A(n134), .B(n8952), .Z(n8950) );
  XOR U10080 ( .A(n8953), .B(n8951), .Z(n8952) );
  NANDN U10081 ( .A(n8861), .B(n8863), .Z(n8904) );
  XOR U10082 ( .A(n8954), .B(n8955), .Z(n8863) );
  AND U10083 ( .A(n134), .B(n8956), .Z(n8954) );
  XOR U10084 ( .A(n8955), .B(n8957), .Z(n8956) );
  XNOR U10085 ( .A(n8958), .B(n8959), .Z(n134) );
  AND U10086 ( .A(n8960), .B(n8961), .Z(n8958) );
  XOR U10087 ( .A(n8959), .B(n8874), .Z(n8961) );
  XNOR U10088 ( .A(n8962), .B(n8963), .Z(n8874) );
  ANDN U10089 ( .B(n8964), .A(n8965), .Z(n8962) );
  XOR U10090 ( .A(n8963), .B(n8966), .Z(n8964) );
  XNOR U10091 ( .A(n8959), .B(n8876), .Z(n8960) );
  XOR U10092 ( .A(n8967), .B(n8968), .Z(n8876) );
  AND U10093 ( .A(n138), .B(n8969), .Z(n8967) );
  XOR U10094 ( .A(n8970), .B(n8968), .Z(n8969) );
  XNOR U10095 ( .A(n8971), .B(n8972), .Z(n8959) );
  AND U10096 ( .A(n8973), .B(n8974), .Z(n8971) );
  XNOR U10097 ( .A(n8972), .B(n8901), .Z(n8974) );
  XOR U10098 ( .A(n8965), .B(n8966), .Z(n8901) );
  XNOR U10099 ( .A(n8975), .B(n8976), .Z(n8966) );
  ANDN U10100 ( .B(n8977), .A(n8978), .Z(n8975) );
  XOR U10101 ( .A(n8979), .B(n8980), .Z(n8977) );
  XOR U10102 ( .A(n8981), .B(n8982), .Z(n8965) );
  XNOR U10103 ( .A(n8983), .B(n8984), .Z(n8982) );
  ANDN U10104 ( .B(n8985), .A(n8986), .Z(n8983) );
  XNOR U10105 ( .A(n8987), .B(n8988), .Z(n8985) );
  IV U10106 ( .A(n8963), .Z(n8981) );
  XOR U10107 ( .A(n8989), .B(n8990), .Z(n8963) );
  ANDN U10108 ( .B(n8991), .A(n8992), .Z(n8989) );
  XOR U10109 ( .A(n8990), .B(n8993), .Z(n8991) );
  XOR U10110 ( .A(n8972), .B(n8903), .Z(n8973) );
  XOR U10111 ( .A(n8994), .B(n8995), .Z(n8903) );
  AND U10112 ( .A(n138), .B(n8996), .Z(n8994) );
  XOR U10113 ( .A(n8997), .B(n8995), .Z(n8996) );
  XNOR U10114 ( .A(n8998), .B(n8999), .Z(n8972) );
  NAND U10115 ( .A(n9000), .B(n9001), .Z(n8999) );
  XOR U10116 ( .A(n9002), .B(n8951), .Z(n9001) );
  XOR U10117 ( .A(n8992), .B(n8993), .Z(n8951) );
  XOR U10118 ( .A(n9003), .B(n8980), .Z(n8993) );
  XOR U10119 ( .A(n9004), .B(n9005), .Z(n8980) );
  ANDN U10120 ( .B(n9006), .A(n9007), .Z(n9004) );
  XOR U10121 ( .A(n9005), .B(n9008), .Z(n9006) );
  IV U10122 ( .A(n8978), .Z(n9003) );
  XOR U10123 ( .A(n8976), .B(n9009), .Z(n8978) );
  XOR U10124 ( .A(n9010), .B(n9011), .Z(n9009) );
  ANDN U10125 ( .B(n9012), .A(n9013), .Z(n9010) );
  XOR U10126 ( .A(n9014), .B(n9011), .Z(n9012) );
  IV U10127 ( .A(n8979), .Z(n8976) );
  XOR U10128 ( .A(n9015), .B(n9016), .Z(n8979) );
  ANDN U10129 ( .B(n9017), .A(n9018), .Z(n9015) );
  XOR U10130 ( .A(n9016), .B(n9019), .Z(n9017) );
  XOR U10131 ( .A(n9020), .B(n9021), .Z(n8992) );
  XNOR U10132 ( .A(n8987), .B(n9022), .Z(n9021) );
  IV U10133 ( .A(n8990), .Z(n9022) );
  XOR U10134 ( .A(n9023), .B(n9024), .Z(n8990) );
  ANDN U10135 ( .B(n9025), .A(n9026), .Z(n9023) );
  XOR U10136 ( .A(n9024), .B(n9027), .Z(n9025) );
  XNOR U10137 ( .A(n9028), .B(n9029), .Z(n8987) );
  ANDN U10138 ( .B(n9030), .A(n9031), .Z(n9028) );
  XOR U10139 ( .A(n9029), .B(n9032), .Z(n9030) );
  IV U10140 ( .A(n8986), .Z(n9020) );
  XOR U10141 ( .A(n8984), .B(n9033), .Z(n8986) );
  XOR U10142 ( .A(n9034), .B(n9035), .Z(n9033) );
  ANDN U10143 ( .B(n9036), .A(n9037), .Z(n9034) );
  XOR U10144 ( .A(n9038), .B(n9035), .Z(n9036) );
  IV U10145 ( .A(n8988), .Z(n8984) );
  XOR U10146 ( .A(n9039), .B(n9040), .Z(n8988) );
  ANDN U10147 ( .B(n9041), .A(n9042), .Z(n9039) );
  XOR U10148 ( .A(n9043), .B(n9040), .Z(n9041) );
  IV U10149 ( .A(n8998), .Z(n9002) );
  XOR U10150 ( .A(n8998), .B(n8953), .Z(n9000) );
  XOR U10151 ( .A(n9044), .B(n9045), .Z(n8953) );
  AND U10152 ( .A(n138), .B(n9046), .Z(n9044) );
  XOR U10153 ( .A(n9047), .B(n9045), .Z(n9046) );
  NANDN U10154 ( .A(n8955), .B(n8957), .Z(n8998) );
  XOR U10155 ( .A(n9048), .B(n9049), .Z(n8957) );
  AND U10156 ( .A(n138), .B(n9050), .Z(n9048) );
  XOR U10157 ( .A(n9049), .B(n9051), .Z(n9050) );
  XNOR U10158 ( .A(n9052), .B(n9053), .Z(n138) );
  AND U10159 ( .A(n9054), .B(n9055), .Z(n9052) );
  XOR U10160 ( .A(n9053), .B(n8968), .Z(n9055) );
  XNOR U10161 ( .A(n9056), .B(n9057), .Z(n8968) );
  ANDN U10162 ( .B(n9058), .A(n9059), .Z(n9056) );
  XOR U10163 ( .A(n9057), .B(n9060), .Z(n9058) );
  XNOR U10164 ( .A(n9053), .B(n8970), .Z(n9054) );
  XOR U10165 ( .A(n9061), .B(n9062), .Z(n8970) );
  AND U10166 ( .A(n142), .B(n9063), .Z(n9061) );
  XOR U10167 ( .A(n9064), .B(n9062), .Z(n9063) );
  XNOR U10168 ( .A(n9065), .B(n9066), .Z(n9053) );
  AND U10169 ( .A(n9067), .B(n9068), .Z(n9065) );
  XNOR U10170 ( .A(n9066), .B(n8995), .Z(n9068) );
  XOR U10171 ( .A(n9059), .B(n9060), .Z(n8995) );
  XNOR U10172 ( .A(n9069), .B(n9070), .Z(n9060) );
  ANDN U10173 ( .B(n9071), .A(n9072), .Z(n9069) );
  XOR U10174 ( .A(n9073), .B(n9074), .Z(n9071) );
  XOR U10175 ( .A(n9075), .B(n9076), .Z(n9059) );
  XNOR U10176 ( .A(n9077), .B(n9078), .Z(n9076) );
  ANDN U10177 ( .B(n9079), .A(n9080), .Z(n9077) );
  XNOR U10178 ( .A(n9081), .B(n9082), .Z(n9079) );
  IV U10179 ( .A(n9057), .Z(n9075) );
  XOR U10180 ( .A(n9083), .B(n9084), .Z(n9057) );
  ANDN U10181 ( .B(n9085), .A(n9086), .Z(n9083) );
  XOR U10182 ( .A(n9084), .B(n9087), .Z(n9085) );
  XOR U10183 ( .A(n9066), .B(n8997), .Z(n9067) );
  XOR U10184 ( .A(n9088), .B(n9089), .Z(n8997) );
  AND U10185 ( .A(n142), .B(n9090), .Z(n9088) );
  XOR U10186 ( .A(n9091), .B(n9089), .Z(n9090) );
  XNOR U10187 ( .A(n9092), .B(n9093), .Z(n9066) );
  NAND U10188 ( .A(n9094), .B(n9095), .Z(n9093) );
  XOR U10189 ( .A(n9096), .B(n9045), .Z(n9095) );
  XOR U10190 ( .A(n9086), .B(n9087), .Z(n9045) );
  XOR U10191 ( .A(n9097), .B(n9074), .Z(n9087) );
  XOR U10192 ( .A(n9098), .B(n9099), .Z(n9074) );
  ANDN U10193 ( .B(n9100), .A(n9101), .Z(n9098) );
  XOR U10194 ( .A(n9099), .B(n9102), .Z(n9100) );
  IV U10195 ( .A(n9072), .Z(n9097) );
  XOR U10196 ( .A(n9070), .B(n9103), .Z(n9072) );
  XOR U10197 ( .A(n9104), .B(n9105), .Z(n9103) );
  ANDN U10198 ( .B(n9106), .A(n9107), .Z(n9104) );
  XOR U10199 ( .A(n9108), .B(n9105), .Z(n9106) );
  IV U10200 ( .A(n9073), .Z(n9070) );
  XOR U10201 ( .A(n9109), .B(n9110), .Z(n9073) );
  ANDN U10202 ( .B(n9111), .A(n9112), .Z(n9109) );
  XOR U10203 ( .A(n9110), .B(n9113), .Z(n9111) );
  XOR U10204 ( .A(n9114), .B(n9115), .Z(n9086) );
  XNOR U10205 ( .A(n9081), .B(n9116), .Z(n9115) );
  IV U10206 ( .A(n9084), .Z(n9116) );
  XOR U10207 ( .A(n9117), .B(n9118), .Z(n9084) );
  ANDN U10208 ( .B(n9119), .A(n9120), .Z(n9117) );
  XOR U10209 ( .A(n9118), .B(n9121), .Z(n9119) );
  XNOR U10210 ( .A(n9122), .B(n9123), .Z(n9081) );
  ANDN U10211 ( .B(n9124), .A(n9125), .Z(n9122) );
  XOR U10212 ( .A(n9123), .B(n9126), .Z(n9124) );
  IV U10213 ( .A(n9080), .Z(n9114) );
  XOR U10214 ( .A(n9078), .B(n9127), .Z(n9080) );
  XOR U10215 ( .A(n9128), .B(n9129), .Z(n9127) );
  ANDN U10216 ( .B(n9130), .A(n9131), .Z(n9128) );
  XOR U10217 ( .A(n9132), .B(n9129), .Z(n9130) );
  IV U10218 ( .A(n9082), .Z(n9078) );
  XOR U10219 ( .A(n9133), .B(n9134), .Z(n9082) );
  ANDN U10220 ( .B(n9135), .A(n9136), .Z(n9133) );
  XOR U10221 ( .A(n9137), .B(n9134), .Z(n9135) );
  IV U10222 ( .A(n9092), .Z(n9096) );
  XOR U10223 ( .A(n9092), .B(n9047), .Z(n9094) );
  XOR U10224 ( .A(n9138), .B(n9139), .Z(n9047) );
  AND U10225 ( .A(n142), .B(n9140), .Z(n9138) );
  XOR U10226 ( .A(n9141), .B(n9139), .Z(n9140) );
  NANDN U10227 ( .A(n9049), .B(n9051), .Z(n9092) );
  XOR U10228 ( .A(n9142), .B(n9143), .Z(n9051) );
  AND U10229 ( .A(n142), .B(n9144), .Z(n9142) );
  XOR U10230 ( .A(n9143), .B(n9145), .Z(n9144) );
  XNOR U10231 ( .A(n9146), .B(n9147), .Z(n142) );
  AND U10232 ( .A(n9148), .B(n9149), .Z(n9146) );
  XOR U10233 ( .A(n9147), .B(n9062), .Z(n9149) );
  XNOR U10234 ( .A(n9150), .B(n9151), .Z(n9062) );
  ANDN U10235 ( .B(n9152), .A(n9153), .Z(n9150) );
  XOR U10236 ( .A(n9151), .B(n9154), .Z(n9152) );
  XNOR U10237 ( .A(n9147), .B(n9064), .Z(n9148) );
  XOR U10238 ( .A(n9155), .B(n9156), .Z(n9064) );
  AND U10239 ( .A(n146), .B(n9157), .Z(n9155) );
  XOR U10240 ( .A(n9158), .B(n9156), .Z(n9157) );
  XNOR U10241 ( .A(n9159), .B(n9160), .Z(n9147) );
  AND U10242 ( .A(n9161), .B(n9162), .Z(n9159) );
  XNOR U10243 ( .A(n9160), .B(n9089), .Z(n9162) );
  XOR U10244 ( .A(n9153), .B(n9154), .Z(n9089) );
  XNOR U10245 ( .A(n9163), .B(n9164), .Z(n9154) );
  ANDN U10246 ( .B(n9165), .A(n9166), .Z(n9163) );
  XOR U10247 ( .A(n9167), .B(n9168), .Z(n9165) );
  XOR U10248 ( .A(n9169), .B(n9170), .Z(n9153) );
  XNOR U10249 ( .A(n9171), .B(n9172), .Z(n9170) );
  ANDN U10250 ( .B(n9173), .A(n9174), .Z(n9171) );
  XNOR U10251 ( .A(n9175), .B(n9176), .Z(n9173) );
  IV U10252 ( .A(n9151), .Z(n9169) );
  XOR U10253 ( .A(n9177), .B(n9178), .Z(n9151) );
  ANDN U10254 ( .B(n9179), .A(n9180), .Z(n9177) );
  XOR U10255 ( .A(n9178), .B(n9181), .Z(n9179) );
  XOR U10256 ( .A(n9160), .B(n9091), .Z(n9161) );
  XOR U10257 ( .A(n9182), .B(n9183), .Z(n9091) );
  AND U10258 ( .A(n146), .B(n9184), .Z(n9182) );
  XOR U10259 ( .A(n9185), .B(n9183), .Z(n9184) );
  XNOR U10260 ( .A(n9186), .B(n9187), .Z(n9160) );
  NAND U10261 ( .A(n9188), .B(n9189), .Z(n9187) );
  XOR U10262 ( .A(n9190), .B(n9139), .Z(n9189) );
  XOR U10263 ( .A(n9180), .B(n9181), .Z(n9139) );
  XOR U10264 ( .A(n9191), .B(n9168), .Z(n9181) );
  XOR U10265 ( .A(n9192), .B(n9193), .Z(n9168) );
  ANDN U10266 ( .B(n9194), .A(n9195), .Z(n9192) );
  XOR U10267 ( .A(n9193), .B(n9196), .Z(n9194) );
  IV U10268 ( .A(n9166), .Z(n9191) );
  XOR U10269 ( .A(n9164), .B(n9197), .Z(n9166) );
  XOR U10270 ( .A(n9198), .B(n9199), .Z(n9197) );
  ANDN U10271 ( .B(n9200), .A(n9201), .Z(n9198) );
  XOR U10272 ( .A(n9202), .B(n9199), .Z(n9200) );
  IV U10273 ( .A(n9167), .Z(n9164) );
  XOR U10274 ( .A(n9203), .B(n9204), .Z(n9167) );
  ANDN U10275 ( .B(n9205), .A(n9206), .Z(n9203) );
  XOR U10276 ( .A(n9204), .B(n9207), .Z(n9205) );
  XOR U10277 ( .A(n9208), .B(n9209), .Z(n9180) );
  XNOR U10278 ( .A(n9175), .B(n9210), .Z(n9209) );
  IV U10279 ( .A(n9178), .Z(n9210) );
  XOR U10280 ( .A(n9211), .B(n9212), .Z(n9178) );
  ANDN U10281 ( .B(n9213), .A(n9214), .Z(n9211) );
  XOR U10282 ( .A(n9212), .B(n9215), .Z(n9213) );
  XNOR U10283 ( .A(n9216), .B(n9217), .Z(n9175) );
  ANDN U10284 ( .B(n9218), .A(n9219), .Z(n9216) );
  XOR U10285 ( .A(n9217), .B(n9220), .Z(n9218) );
  IV U10286 ( .A(n9174), .Z(n9208) );
  XOR U10287 ( .A(n9172), .B(n9221), .Z(n9174) );
  XOR U10288 ( .A(n9222), .B(n9223), .Z(n9221) );
  ANDN U10289 ( .B(n9224), .A(n9225), .Z(n9222) );
  XOR U10290 ( .A(n9226), .B(n9223), .Z(n9224) );
  IV U10291 ( .A(n9176), .Z(n9172) );
  XOR U10292 ( .A(n9227), .B(n9228), .Z(n9176) );
  ANDN U10293 ( .B(n9229), .A(n9230), .Z(n9227) );
  XOR U10294 ( .A(n9231), .B(n9228), .Z(n9229) );
  IV U10295 ( .A(n9186), .Z(n9190) );
  XOR U10296 ( .A(n9186), .B(n9141), .Z(n9188) );
  XOR U10297 ( .A(n9232), .B(n9233), .Z(n9141) );
  AND U10298 ( .A(n146), .B(n9234), .Z(n9232) );
  XOR U10299 ( .A(n9235), .B(n9233), .Z(n9234) );
  NANDN U10300 ( .A(n9143), .B(n9145), .Z(n9186) );
  XOR U10301 ( .A(n9236), .B(n9237), .Z(n9145) );
  AND U10302 ( .A(n146), .B(n9238), .Z(n9236) );
  XOR U10303 ( .A(n9237), .B(n9239), .Z(n9238) );
  XNOR U10304 ( .A(n9240), .B(n9241), .Z(n146) );
  AND U10305 ( .A(n9242), .B(n9243), .Z(n9240) );
  XOR U10306 ( .A(n9241), .B(n9156), .Z(n9243) );
  XNOR U10307 ( .A(n9244), .B(n9245), .Z(n9156) );
  ANDN U10308 ( .B(n9246), .A(n9247), .Z(n9244) );
  XOR U10309 ( .A(n9245), .B(n9248), .Z(n9246) );
  XNOR U10310 ( .A(n9241), .B(n9158), .Z(n9242) );
  XOR U10311 ( .A(n9249), .B(n9250), .Z(n9158) );
  AND U10312 ( .A(n150), .B(n9251), .Z(n9249) );
  XOR U10313 ( .A(n9252), .B(n9250), .Z(n9251) );
  XNOR U10314 ( .A(n9253), .B(n9254), .Z(n9241) );
  AND U10315 ( .A(n9255), .B(n9256), .Z(n9253) );
  XNOR U10316 ( .A(n9254), .B(n9183), .Z(n9256) );
  XOR U10317 ( .A(n9247), .B(n9248), .Z(n9183) );
  XNOR U10318 ( .A(n9257), .B(n9258), .Z(n9248) );
  ANDN U10319 ( .B(n9259), .A(n9260), .Z(n9257) );
  XOR U10320 ( .A(n9261), .B(n9262), .Z(n9259) );
  XOR U10321 ( .A(n9263), .B(n9264), .Z(n9247) );
  XNOR U10322 ( .A(n9265), .B(n9266), .Z(n9264) );
  ANDN U10323 ( .B(n9267), .A(n9268), .Z(n9265) );
  XNOR U10324 ( .A(n9269), .B(n9270), .Z(n9267) );
  IV U10325 ( .A(n9245), .Z(n9263) );
  XOR U10326 ( .A(n9271), .B(n9272), .Z(n9245) );
  ANDN U10327 ( .B(n9273), .A(n9274), .Z(n9271) );
  XOR U10328 ( .A(n9272), .B(n9275), .Z(n9273) );
  XOR U10329 ( .A(n9254), .B(n9185), .Z(n9255) );
  XOR U10330 ( .A(n9276), .B(n9277), .Z(n9185) );
  AND U10331 ( .A(n150), .B(n9278), .Z(n9276) );
  XOR U10332 ( .A(n9279), .B(n9277), .Z(n9278) );
  XNOR U10333 ( .A(n9280), .B(n9281), .Z(n9254) );
  NAND U10334 ( .A(n9282), .B(n9283), .Z(n9281) );
  XOR U10335 ( .A(n9284), .B(n9233), .Z(n9283) );
  XOR U10336 ( .A(n9274), .B(n9275), .Z(n9233) );
  XOR U10337 ( .A(n9285), .B(n9262), .Z(n9275) );
  XOR U10338 ( .A(n9286), .B(n9287), .Z(n9262) );
  ANDN U10339 ( .B(n9288), .A(n9289), .Z(n9286) );
  XOR U10340 ( .A(n9287), .B(n9290), .Z(n9288) );
  IV U10341 ( .A(n9260), .Z(n9285) );
  XOR U10342 ( .A(n9258), .B(n9291), .Z(n9260) );
  XOR U10343 ( .A(n9292), .B(n9293), .Z(n9291) );
  ANDN U10344 ( .B(n9294), .A(n9295), .Z(n9292) );
  XOR U10345 ( .A(n9296), .B(n9293), .Z(n9294) );
  IV U10346 ( .A(n9261), .Z(n9258) );
  XOR U10347 ( .A(n9297), .B(n9298), .Z(n9261) );
  ANDN U10348 ( .B(n9299), .A(n9300), .Z(n9297) );
  XOR U10349 ( .A(n9298), .B(n9301), .Z(n9299) );
  XOR U10350 ( .A(n9302), .B(n9303), .Z(n9274) );
  XNOR U10351 ( .A(n9269), .B(n9304), .Z(n9303) );
  IV U10352 ( .A(n9272), .Z(n9304) );
  XOR U10353 ( .A(n9305), .B(n9306), .Z(n9272) );
  ANDN U10354 ( .B(n9307), .A(n9308), .Z(n9305) );
  XOR U10355 ( .A(n9306), .B(n9309), .Z(n9307) );
  XNOR U10356 ( .A(n9310), .B(n9311), .Z(n9269) );
  ANDN U10357 ( .B(n9312), .A(n9313), .Z(n9310) );
  XOR U10358 ( .A(n9311), .B(n9314), .Z(n9312) );
  IV U10359 ( .A(n9268), .Z(n9302) );
  XOR U10360 ( .A(n9266), .B(n9315), .Z(n9268) );
  XOR U10361 ( .A(n9316), .B(n9317), .Z(n9315) );
  ANDN U10362 ( .B(n9318), .A(n9319), .Z(n9316) );
  XOR U10363 ( .A(n9320), .B(n9317), .Z(n9318) );
  IV U10364 ( .A(n9270), .Z(n9266) );
  XOR U10365 ( .A(n9321), .B(n9322), .Z(n9270) );
  ANDN U10366 ( .B(n9323), .A(n9324), .Z(n9321) );
  XOR U10367 ( .A(n9325), .B(n9322), .Z(n9323) );
  IV U10368 ( .A(n9280), .Z(n9284) );
  XOR U10369 ( .A(n9280), .B(n9235), .Z(n9282) );
  XOR U10370 ( .A(n9326), .B(n9327), .Z(n9235) );
  AND U10371 ( .A(n150), .B(n9328), .Z(n9326) );
  XOR U10372 ( .A(n9329), .B(n9327), .Z(n9328) );
  NANDN U10373 ( .A(n9237), .B(n9239), .Z(n9280) );
  XOR U10374 ( .A(n9330), .B(n9331), .Z(n9239) );
  AND U10375 ( .A(n150), .B(n9332), .Z(n9330) );
  XOR U10376 ( .A(n9331), .B(n9333), .Z(n9332) );
  XNOR U10377 ( .A(n9334), .B(n9335), .Z(n150) );
  AND U10378 ( .A(n9336), .B(n9337), .Z(n9334) );
  XOR U10379 ( .A(n9335), .B(n9250), .Z(n9337) );
  XNOR U10380 ( .A(n9338), .B(n9339), .Z(n9250) );
  ANDN U10381 ( .B(n9340), .A(n9341), .Z(n9338) );
  XOR U10382 ( .A(n9339), .B(n9342), .Z(n9340) );
  XNOR U10383 ( .A(n9335), .B(n9252), .Z(n9336) );
  XOR U10384 ( .A(n9343), .B(n9344), .Z(n9252) );
  AND U10385 ( .A(n154), .B(n9345), .Z(n9343) );
  XOR U10386 ( .A(n9346), .B(n9344), .Z(n9345) );
  XNOR U10387 ( .A(n9347), .B(n9348), .Z(n9335) );
  AND U10388 ( .A(n9349), .B(n9350), .Z(n9347) );
  XNOR U10389 ( .A(n9348), .B(n9277), .Z(n9350) );
  XOR U10390 ( .A(n9341), .B(n9342), .Z(n9277) );
  XNOR U10391 ( .A(n9351), .B(n9352), .Z(n9342) );
  ANDN U10392 ( .B(n9353), .A(n9354), .Z(n9351) );
  XOR U10393 ( .A(n9355), .B(n9356), .Z(n9353) );
  XOR U10394 ( .A(n9357), .B(n9358), .Z(n9341) );
  XNOR U10395 ( .A(n9359), .B(n9360), .Z(n9358) );
  ANDN U10396 ( .B(n9361), .A(n9362), .Z(n9359) );
  XNOR U10397 ( .A(n9363), .B(n9364), .Z(n9361) );
  IV U10398 ( .A(n9339), .Z(n9357) );
  XOR U10399 ( .A(n9365), .B(n9366), .Z(n9339) );
  ANDN U10400 ( .B(n9367), .A(n9368), .Z(n9365) );
  XOR U10401 ( .A(n9366), .B(n9369), .Z(n9367) );
  XOR U10402 ( .A(n9348), .B(n9279), .Z(n9349) );
  XOR U10403 ( .A(n9370), .B(n9371), .Z(n9279) );
  AND U10404 ( .A(n154), .B(n9372), .Z(n9370) );
  XOR U10405 ( .A(n9373), .B(n9371), .Z(n9372) );
  XNOR U10406 ( .A(n9374), .B(n9375), .Z(n9348) );
  NAND U10407 ( .A(n9376), .B(n9377), .Z(n9375) );
  XOR U10408 ( .A(n9378), .B(n9327), .Z(n9377) );
  XOR U10409 ( .A(n9368), .B(n9369), .Z(n9327) );
  XOR U10410 ( .A(n9379), .B(n9356), .Z(n9369) );
  XOR U10411 ( .A(n9380), .B(n9381), .Z(n9356) );
  ANDN U10412 ( .B(n9382), .A(n9383), .Z(n9380) );
  XOR U10413 ( .A(n9381), .B(n9384), .Z(n9382) );
  IV U10414 ( .A(n9354), .Z(n9379) );
  XOR U10415 ( .A(n9352), .B(n9385), .Z(n9354) );
  XOR U10416 ( .A(n9386), .B(n9387), .Z(n9385) );
  ANDN U10417 ( .B(n9388), .A(n9389), .Z(n9386) );
  XOR U10418 ( .A(n9390), .B(n9387), .Z(n9388) );
  IV U10419 ( .A(n9355), .Z(n9352) );
  XOR U10420 ( .A(n9391), .B(n9392), .Z(n9355) );
  ANDN U10421 ( .B(n9393), .A(n9394), .Z(n9391) );
  XOR U10422 ( .A(n9392), .B(n9395), .Z(n9393) );
  XOR U10423 ( .A(n9396), .B(n9397), .Z(n9368) );
  XNOR U10424 ( .A(n9363), .B(n9398), .Z(n9397) );
  IV U10425 ( .A(n9366), .Z(n9398) );
  XOR U10426 ( .A(n9399), .B(n9400), .Z(n9366) );
  ANDN U10427 ( .B(n9401), .A(n9402), .Z(n9399) );
  XOR U10428 ( .A(n9400), .B(n9403), .Z(n9401) );
  XNOR U10429 ( .A(n9404), .B(n9405), .Z(n9363) );
  ANDN U10430 ( .B(n9406), .A(n9407), .Z(n9404) );
  XOR U10431 ( .A(n9405), .B(n9408), .Z(n9406) );
  IV U10432 ( .A(n9362), .Z(n9396) );
  XOR U10433 ( .A(n9360), .B(n9409), .Z(n9362) );
  XOR U10434 ( .A(n9410), .B(n9411), .Z(n9409) );
  ANDN U10435 ( .B(n9412), .A(n9413), .Z(n9410) );
  XOR U10436 ( .A(n9414), .B(n9411), .Z(n9412) );
  IV U10437 ( .A(n9364), .Z(n9360) );
  XOR U10438 ( .A(n9415), .B(n9416), .Z(n9364) );
  ANDN U10439 ( .B(n9417), .A(n9418), .Z(n9415) );
  XOR U10440 ( .A(n9419), .B(n9416), .Z(n9417) );
  IV U10441 ( .A(n9374), .Z(n9378) );
  XOR U10442 ( .A(n9374), .B(n9329), .Z(n9376) );
  XOR U10443 ( .A(n9420), .B(n9421), .Z(n9329) );
  AND U10444 ( .A(n154), .B(n9422), .Z(n9420) );
  XOR U10445 ( .A(n9423), .B(n9421), .Z(n9422) );
  NANDN U10446 ( .A(n9331), .B(n9333), .Z(n9374) );
  XOR U10447 ( .A(n9424), .B(n9425), .Z(n9333) );
  AND U10448 ( .A(n154), .B(n9426), .Z(n9424) );
  XOR U10449 ( .A(n9425), .B(n9427), .Z(n9426) );
  XNOR U10450 ( .A(n9428), .B(n9429), .Z(n154) );
  AND U10451 ( .A(n9430), .B(n9431), .Z(n9428) );
  XOR U10452 ( .A(n9429), .B(n9344), .Z(n9431) );
  XNOR U10453 ( .A(n9432), .B(n9433), .Z(n9344) );
  ANDN U10454 ( .B(n9434), .A(n9435), .Z(n9432) );
  XOR U10455 ( .A(n9433), .B(n9436), .Z(n9434) );
  XNOR U10456 ( .A(n9429), .B(n9346), .Z(n9430) );
  XOR U10457 ( .A(n9437), .B(n9438), .Z(n9346) );
  AND U10458 ( .A(n158), .B(n9439), .Z(n9437) );
  XOR U10459 ( .A(n9440), .B(n9438), .Z(n9439) );
  XNOR U10460 ( .A(n9441), .B(n9442), .Z(n9429) );
  AND U10461 ( .A(n9443), .B(n9444), .Z(n9441) );
  XNOR U10462 ( .A(n9442), .B(n9371), .Z(n9444) );
  XOR U10463 ( .A(n9435), .B(n9436), .Z(n9371) );
  XNOR U10464 ( .A(n9445), .B(n9446), .Z(n9436) );
  ANDN U10465 ( .B(n9447), .A(n9448), .Z(n9445) );
  XOR U10466 ( .A(n9449), .B(n9450), .Z(n9447) );
  XOR U10467 ( .A(n9451), .B(n9452), .Z(n9435) );
  XNOR U10468 ( .A(n9453), .B(n9454), .Z(n9452) );
  ANDN U10469 ( .B(n9455), .A(n9456), .Z(n9453) );
  XNOR U10470 ( .A(n9457), .B(n9458), .Z(n9455) );
  IV U10471 ( .A(n9433), .Z(n9451) );
  XOR U10472 ( .A(n9459), .B(n9460), .Z(n9433) );
  ANDN U10473 ( .B(n9461), .A(n9462), .Z(n9459) );
  XOR U10474 ( .A(n9460), .B(n9463), .Z(n9461) );
  XOR U10475 ( .A(n9442), .B(n9373), .Z(n9443) );
  XOR U10476 ( .A(n9464), .B(n9465), .Z(n9373) );
  AND U10477 ( .A(n158), .B(n9466), .Z(n9464) );
  XOR U10478 ( .A(n9467), .B(n9465), .Z(n9466) );
  XNOR U10479 ( .A(n9468), .B(n9469), .Z(n9442) );
  NAND U10480 ( .A(n9470), .B(n9471), .Z(n9469) );
  XOR U10481 ( .A(n9472), .B(n9421), .Z(n9471) );
  XOR U10482 ( .A(n9462), .B(n9463), .Z(n9421) );
  XOR U10483 ( .A(n9473), .B(n9450), .Z(n9463) );
  XOR U10484 ( .A(n9474), .B(n9475), .Z(n9450) );
  ANDN U10485 ( .B(n9476), .A(n9477), .Z(n9474) );
  XOR U10486 ( .A(n9475), .B(n9478), .Z(n9476) );
  IV U10487 ( .A(n9448), .Z(n9473) );
  XOR U10488 ( .A(n9446), .B(n9479), .Z(n9448) );
  XOR U10489 ( .A(n9480), .B(n9481), .Z(n9479) );
  ANDN U10490 ( .B(n9482), .A(n9483), .Z(n9480) );
  XOR U10491 ( .A(n9484), .B(n9481), .Z(n9482) );
  IV U10492 ( .A(n9449), .Z(n9446) );
  XOR U10493 ( .A(n9485), .B(n9486), .Z(n9449) );
  ANDN U10494 ( .B(n9487), .A(n9488), .Z(n9485) );
  XOR U10495 ( .A(n9486), .B(n9489), .Z(n9487) );
  XOR U10496 ( .A(n9490), .B(n9491), .Z(n9462) );
  XNOR U10497 ( .A(n9457), .B(n9492), .Z(n9491) );
  IV U10498 ( .A(n9460), .Z(n9492) );
  XOR U10499 ( .A(n9493), .B(n9494), .Z(n9460) );
  ANDN U10500 ( .B(n9495), .A(n9496), .Z(n9493) );
  XOR U10501 ( .A(n9494), .B(n9497), .Z(n9495) );
  XNOR U10502 ( .A(n9498), .B(n9499), .Z(n9457) );
  ANDN U10503 ( .B(n9500), .A(n9501), .Z(n9498) );
  XOR U10504 ( .A(n9499), .B(n9502), .Z(n9500) );
  IV U10505 ( .A(n9456), .Z(n9490) );
  XOR U10506 ( .A(n9454), .B(n9503), .Z(n9456) );
  XOR U10507 ( .A(n9504), .B(n9505), .Z(n9503) );
  ANDN U10508 ( .B(n9506), .A(n9507), .Z(n9504) );
  XOR U10509 ( .A(n9508), .B(n9505), .Z(n9506) );
  IV U10510 ( .A(n9458), .Z(n9454) );
  XOR U10511 ( .A(n9509), .B(n9510), .Z(n9458) );
  ANDN U10512 ( .B(n9511), .A(n9512), .Z(n9509) );
  XOR U10513 ( .A(n9513), .B(n9510), .Z(n9511) );
  IV U10514 ( .A(n9468), .Z(n9472) );
  XOR U10515 ( .A(n9468), .B(n9423), .Z(n9470) );
  XOR U10516 ( .A(n9514), .B(n9515), .Z(n9423) );
  AND U10517 ( .A(n158), .B(n9516), .Z(n9514) );
  XOR U10518 ( .A(n9517), .B(n9515), .Z(n9516) );
  NANDN U10519 ( .A(n9425), .B(n9427), .Z(n9468) );
  XOR U10520 ( .A(n9518), .B(n9519), .Z(n9427) );
  AND U10521 ( .A(n158), .B(n9520), .Z(n9518) );
  XOR U10522 ( .A(n9519), .B(n9521), .Z(n9520) );
  XNOR U10523 ( .A(n9522), .B(n9523), .Z(n158) );
  AND U10524 ( .A(n9524), .B(n9525), .Z(n9522) );
  XOR U10525 ( .A(n9523), .B(n9438), .Z(n9525) );
  XNOR U10526 ( .A(n9526), .B(n9527), .Z(n9438) );
  ANDN U10527 ( .B(n9528), .A(n9529), .Z(n9526) );
  XOR U10528 ( .A(n9527), .B(n9530), .Z(n9528) );
  XNOR U10529 ( .A(n9523), .B(n9440), .Z(n9524) );
  XOR U10530 ( .A(n9531), .B(n9532), .Z(n9440) );
  AND U10531 ( .A(n162), .B(n9533), .Z(n9531) );
  XOR U10532 ( .A(n9534), .B(n9532), .Z(n9533) );
  XNOR U10533 ( .A(n9535), .B(n9536), .Z(n9523) );
  AND U10534 ( .A(n9537), .B(n9538), .Z(n9535) );
  XNOR U10535 ( .A(n9536), .B(n9465), .Z(n9538) );
  XOR U10536 ( .A(n9529), .B(n9530), .Z(n9465) );
  XNOR U10537 ( .A(n9539), .B(n9540), .Z(n9530) );
  ANDN U10538 ( .B(n9541), .A(n9542), .Z(n9539) );
  XOR U10539 ( .A(n9543), .B(n9544), .Z(n9541) );
  XOR U10540 ( .A(n9545), .B(n9546), .Z(n9529) );
  XNOR U10541 ( .A(n9547), .B(n9548), .Z(n9546) );
  ANDN U10542 ( .B(n9549), .A(n9550), .Z(n9547) );
  XNOR U10543 ( .A(n9551), .B(n9552), .Z(n9549) );
  IV U10544 ( .A(n9527), .Z(n9545) );
  XOR U10545 ( .A(n9553), .B(n9554), .Z(n9527) );
  ANDN U10546 ( .B(n9555), .A(n9556), .Z(n9553) );
  XOR U10547 ( .A(n9554), .B(n9557), .Z(n9555) );
  XOR U10548 ( .A(n9536), .B(n9467), .Z(n9537) );
  XOR U10549 ( .A(n9558), .B(n9559), .Z(n9467) );
  AND U10550 ( .A(n162), .B(n9560), .Z(n9558) );
  XOR U10551 ( .A(n9561), .B(n9559), .Z(n9560) );
  XNOR U10552 ( .A(n9562), .B(n9563), .Z(n9536) );
  NAND U10553 ( .A(n9564), .B(n9565), .Z(n9563) );
  XOR U10554 ( .A(n9566), .B(n9515), .Z(n9565) );
  XOR U10555 ( .A(n9556), .B(n9557), .Z(n9515) );
  XOR U10556 ( .A(n9567), .B(n9544), .Z(n9557) );
  XOR U10557 ( .A(n9568), .B(n9569), .Z(n9544) );
  ANDN U10558 ( .B(n9570), .A(n9571), .Z(n9568) );
  XOR U10559 ( .A(n9569), .B(n9572), .Z(n9570) );
  IV U10560 ( .A(n9542), .Z(n9567) );
  XOR U10561 ( .A(n9540), .B(n9573), .Z(n9542) );
  XOR U10562 ( .A(n9574), .B(n9575), .Z(n9573) );
  ANDN U10563 ( .B(n9576), .A(n9577), .Z(n9574) );
  XOR U10564 ( .A(n9578), .B(n9575), .Z(n9576) );
  IV U10565 ( .A(n9543), .Z(n9540) );
  XOR U10566 ( .A(n9579), .B(n9580), .Z(n9543) );
  ANDN U10567 ( .B(n9581), .A(n9582), .Z(n9579) );
  XOR U10568 ( .A(n9580), .B(n9583), .Z(n9581) );
  XOR U10569 ( .A(n9584), .B(n9585), .Z(n9556) );
  XNOR U10570 ( .A(n9551), .B(n9586), .Z(n9585) );
  IV U10571 ( .A(n9554), .Z(n9586) );
  XOR U10572 ( .A(n9587), .B(n9588), .Z(n9554) );
  ANDN U10573 ( .B(n9589), .A(n9590), .Z(n9587) );
  XOR U10574 ( .A(n9588), .B(n9591), .Z(n9589) );
  XNOR U10575 ( .A(n9592), .B(n9593), .Z(n9551) );
  ANDN U10576 ( .B(n9594), .A(n9595), .Z(n9592) );
  XOR U10577 ( .A(n9593), .B(n9596), .Z(n9594) );
  IV U10578 ( .A(n9550), .Z(n9584) );
  XOR U10579 ( .A(n9548), .B(n9597), .Z(n9550) );
  XOR U10580 ( .A(n9598), .B(n9599), .Z(n9597) );
  ANDN U10581 ( .B(n9600), .A(n9601), .Z(n9598) );
  XOR U10582 ( .A(n9602), .B(n9599), .Z(n9600) );
  IV U10583 ( .A(n9552), .Z(n9548) );
  XOR U10584 ( .A(n9603), .B(n9604), .Z(n9552) );
  ANDN U10585 ( .B(n9605), .A(n9606), .Z(n9603) );
  XOR U10586 ( .A(n9607), .B(n9604), .Z(n9605) );
  IV U10587 ( .A(n9562), .Z(n9566) );
  XOR U10588 ( .A(n9562), .B(n9517), .Z(n9564) );
  XOR U10589 ( .A(n9608), .B(n9609), .Z(n9517) );
  AND U10590 ( .A(n162), .B(n9610), .Z(n9608) );
  XOR U10591 ( .A(n9611), .B(n9609), .Z(n9610) );
  NANDN U10592 ( .A(n9519), .B(n9521), .Z(n9562) );
  XOR U10593 ( .A(n9612), .B(n9613), .Z(n9521) );
  AND U10594 ( .A(n162), .B(n9614), .Z(n9612) );
  XOR U10595 ( .A(n9613), .B(n9615), .Z(n9614) );
  XNOR U10596 ( .A(n9616), .B(n9617), .Z(n162) );
  AND U10597 ( .A(n9618), .B(n9619), .Z(n9616) );
  XOR U10598 ( .A(n9617), .B(n9532), .Z(n9619) );
  XNOR U10599 ( .A(n9620), .B(n9621), .Z(n9532) );
  ANDN U10600 ( .B(n9622), .A(n9623), .Z(n9620) );
  XOR U10601 ( .A(n9621), .B(n9624), .Z(n9622) );
  XNOR U10602 ( .A(n9617), .B(n9534), .Z(n9618) );
  XOR U10603 ( .A(n9625), .B(n9626), .Z(n9534) );
  AND U10604 ( .A(n166), .B(n9627), .Z(n9625) );
  XOR U10605 ( .A(n9628), .B(n9626), .Z(n9627) );
  XNOR U10606 ( .A(n9629), .B(n9630), .Z(n9617) );
  AND U10607 ( .A(n9631), .B(n9632), .Z(n9629) );
  XNOR U10608 ( .A(n9630), .B(n9559), .Z(n9632) );
  XOR U10609 ( .A(n9623), .B(n9624), .Z(n9559) );
  XNOR U10610 ( .A(n9633), .B(n9634), .Z(n9624) );
  ANDN U10611 ( .B(n9635), .A(n9636), .Z(n9633) );
  XOR U10612 ( .A(n9637), .B(n9638), .Z(n9635) );
  XOR U10613 ( .A(n9639), .B(n9640), .Z(n9623) );
  XNOR U10614 ( .A(n9641), .B(n9642), .Z(n9640) );
  ANDN U10615 ( .B(n9643), .A(n9644), .Z(n9641) );
  XNOR U10616 ( .A(n9645), .B(n9646), .Z(n9643) );
  IV U10617 ( .A(n9621), .Z(n9639) );
  XOR U10618 ( .A(n9647), .B(n9648), .Z(n9621) );
  ANDN U10619 ( .B(n9649), .A(n9650), .Z(n9647) );
  XOR U10620 ( .A(n9648), .B(n9651), .Z(n9649) );
  XOR U10621 ( .A(n9630), .B(n9561), .Z(n9631) );
  XOR U10622 ( .A(n9652), .B(n9653), .Z(n9561) );
  AND U10623 ( .A(n166), .B(n9654), .Z(n9652) );
  XOR U10624 ( .A(n9655), .B(n9653), .Z(n9654) );
  XNOR U10625 ( .A(n9656), .B(n9657), .Z(n9630) );
  NAND U10626 ( .A(n9658), .B(n9659), .Z(n9657) );
  XOR U10627 ( .A(n9660), .B(n9609), .Z(n9659) );
  XOR U10628 ( .A(n9650), .B(n9651), .Z(n9609) );
  XOR U10629 ( .A(n9661), .B(n9638), .Z(n9651) );
  XOR U10630 ( .A(n9662), .B(n9663), .Z(n9638) );
  ANDN U10631 ( .B(n9664), .A(n9665), .Z(n9662) );
  XOR U10632 ( .A(n9663), .B(n9666), .Z(n9664) );
  IV U10633 ( .A(n9636), .Z(n9661) );
  XOR U10634 ( .A(n9634), .B(n9667), .Z(n9636) );
  XOR U10635 ( .A(n9668), .B(n9669), .Z(n9667) );
  ANDN U10636 ( .B(n9670), .A(n9671), .Z(n9668) );
  XOR U10637 ( .A(n9672), .B(n9669), .Z(n9670) );
  IV U10638 ( .A(n9637), .Z(n9634) );
  XOR U10639 ( .A(n9673), .B(n9674), .Z(n9637) );
  ANDN U10640 ( .B(n9675), .A(n9676), .Z(n9673) );
  XOR U10641 ( .A(n9674), .B(n9677), .Z(n9675) );
  XOR U10642 ( .A(n9678), .B(n9679), .Z(n9650) );
  XNOR U10643 ( .A(n9645), .B(n9680), .Z(n9679) );
  IV U10644 ( .A(n9648), .Z(n9680) );
  XOR U10645 ( .A(n9681), .B(n9682), .Z(n9648) );
  ANDN U10646 ( .B(n9683), .A(n9684), .Z(n9681) );
  XOR U10647 ( .A(n9682), .B(n9685), .Z(n9683) );
  XNOR U10648 ( .A(n9686), .B(n9687), .Z(n9645) );
  ANDN U10649 ( .B(n9688), .A(n9689), .Z(n9686) );
  XOR U10650 ( .A(n9687), .B(n9690), .Z(n9688) );
  IV U10651 ( .A(n9644), .Z(n9678) );
  XOR U10652 ( .A(n9642), .B(n9691), .Z(n9644) );
  XOR U10653 ( .A(n9692), .B(n9693), .Z(n9691) );
  ANDN U10654 ( .B(n9694), .A(n9695), .Z(n9692) );
  XOR U10655 ( .A(n9696), .B(n9693), .Z(n9694) );
  IV U10656 ( .A(n9646), .Z(n9642) );
  XOR U10657 ( .A(n9697), .B(n9698), .Z(n9646) );
  ANDN U10658 ( .B(n9699), .A(n9700), .Z(n9697) );
  XOR U10659 ( .A(n9701), .B(n9698), .Z(n9699) );
  IV U10660 ( .A(n9656), .Z(n9660) );
  XOR U10661 ( .A(n9656), .B(n9611), .Z(n9658) );
  XOR U10662 ( .A(n9702), .B(n9703), .Z(n9611) );
  AND U10663 ( .A(n166), .B(n9704), .Z(n9702) );
  XOR U10664 ( .A(n9705), .B(n9703), .Z(n9704) );
  NANDN U10665 ( .A(n9613), .B(n9615), .Z(n9656) );
  XOR U10666 ( .A(n9706), .B(n9707), .Z(n9615) );
  AND U10667 ( .A(n166), .B(n9708), .Z(n9706) );
  XOR U10668 ( .A(n9707), .B(n9709), .Z(n9708) );
  XNOR U10669 ( .A(n9710), .B(n9711), .Z(n166) );
  AND U10670 ( .A(n9712), .B(n9713), .Z(n9710) );
  XOR U10671 ( .A(n9711), .B(n9626), .Z(n9713) );
  XNOR U10672 ( .A(n9714), .B(n9715), .Z(n9626) );
  ANDN U10673 ( .B(n9716), .A(n9717), .Z(n9714) );
  XOR U10674 ( .A(n9715), .B(n9718), .Z(n9716) );
  XNOR U10675 ( .A(n9711), .B(n9628), .Z(n9712) );
  XOR U10676 ( .A(n9719), .B(n9720), .Z(n9628) );
  AND U10677 ( .A(n170), .B(n9721), .Z(n9719) );
  XOR U10678 ( .A(n9722), .B(n9720), .Z(n9721) );
  XNOR U10679 ( .A(n9723), .B(n9724), .Z(n9711) );
  AND U10680 ( .A(n9725), .B(n9726), .Z(n9723) );
  XNOR U10681 ( .A(n9724), .B(n9653), .Z(n9726) );
  XOR U10682 ( .A(n9717), .B(n9718), .Z(n9653) );
  XNOR U10683 ( .A(n9727), .B(n9728), .Z(n9718) );
  ANDN U10684 ( .B(n9729), .A(n9730), .Z(n9727) );
  XOR U10685 ( .A(n9731), .B(n9732), .Z(n9729) );
  XOR U10686 ( .A(n9733), .B(n9734), .Z(n9717) );
  XNOR U10687 ( .A(n9735), .B(n9736), .Z(n9734) );
  ANDN U10688 ( .B(n9737), .A(n9738), .Z(n9735) );
  XNOR U10689 ( .A(n9739), .B(n9740), .Z(n9737) );
  IV U10690 ( .A(n9715), .Z(n9733) );
  XOR U10691 ( .A(n9741), .B(n9742), .Z(n9715) );
  ANDN U10692 ( .B(n9743), .A(n9744), .Z(n9741) );
  XOR U10693 ( .A(n9742), .B(n9745), .Z(n9743) );
  XOR U10694 ( .A(n9724), .B(n9655), .Z(n9725) );
  XOR U10695 ( .A(n9746), .B(n9747), .Z(n9655) );
  AND U10696 ( .A(n170), .B(n9748), .Z(n9746) );
  XOR U10697 ( .A(n9749), .B(n9747), .Z(n9748) );
  XNOR U10698 ( .A(n9750), .B(n9751), .Z(n9724) );
  NAND U10699 ( .A(n9752), .B(n9753), .Z(n9751) );
  XOR U10700 ( .A(n9754), .B(n9703), .Z(n9753) );
  XOR U10701 ( .A(n9744), .B(n9745), .Z(n9703) );
  XOR U10702 ( .A(n9755), .B(n9732), .Z(n9745) );
  XOR U10703 ( .A(n9756), .B(n9757), .Z(n9732) );
  ANDN U10704 ( .B(n9758), .A(n9759), .Z(n9756) );
  XOR U10705 ( .A(n9757), .B(n9760), .Z(n9758) );
  IV U10706 ( .A(n9730), .Z(n9755) );
  XOR U10707 ( .A(n9728), .B(n9761), .Z(n9730) );
  XOR U10708 ( .A(n9762), .B(n9763), .Z(n9761) );
  ANDN U10709 ( .B(n9764), .A(n9765), .Z(n9762) );
  XOR U10710 ( .A(n9766), .B(n9763), .Z(n9764) );
  IV U10711 ( .A(n9731), .Z(n9728) );
  XOR U10712 ( .A(n9767), .B(n9768), .Z(n9731) );
  ANDN U10713 ( .B(n9769), .A(n9770), .Z(n9767) );
  XOR U10714 ( .A(n9768), .B(n9771), .Z(n9769) );
  XOR U10715 ( .A(n9772), .B(n9773), .Z(n9744) );
  XNOR U10716 ( .A(n9739), .B(n9774), .Z(n9773) );
  IV U10717 ( .A(n9742), .Z(n9774) );
  XOR U10718 ( .A(n9775), .B(n9776), .Z(n9742) );
  ANDN U10719 ( .B(n9777), .A(n9778), .Z(n9775) );
  XOR U10720 ( .A(n9776), .B(n9779), .Z(n9777) );
  XNOR U10721 ( .A(n9780), .B(n9781), .Z(n9739) );
  ANDN U10722 ( .B(n9782), .A(n9783), .Z(n9780) );
  XOR U10723 ( .A(n9781), .B(n9784), .Z(n9782) );
  IV U10724 ( .A(n9738), .Z(n9772) );
  XOR U10725 ( .A(n9736), .B(n9785), .Z(n9738) );
  XOR U10726 ( .A(n9786), .B(n9787), .Z(n9785) );
  ANDN U10727 ( .B(n9788), .A(n9789), .Z(n9786) );
  XOR U10728 ( .A(n9790), .B(n9787), .Z(n9788) );
  IV U10729 ( .A(n9740), .Z(n9736) );
  XOR U10730 ( .A(n9791), .B(n9792), .Z(n9740) );
  ANDN U10731 ( .B(n9793), .A(n9794), .Z(n9791) );
  XOR U10732 ( .A(n9795), .B(n9792), .Z(n9793) );
  IV U10733 ( .A(n9750), .Z(n9754) );
  XOR U10734 ( .A(n9750), .B(n9705), .Z(n9752) );
  XOR U10735 ( .A(n9796), .B(n9797), .Z(n9705) );
  AND U10736 ( .A(n170), .B(n9798), .Z(n9796) );
  XOR U10737 ( .A(n9799), .B(n9797), .Z(n9798) );
  NANDN U10738 ( .A(n9707), .B(n9709), .Z(n9750) );
  XOR U10739 ( .A(n9800), .B(n9801), .Z(n9709) );
  AND U10740 ( .A(n170), .B(n9802), .Z(n9800) );
  XOR U10741 ( .A(n9801), .B(n9803), .Z(n9802) );
  XNOR U10742 ( .A(n9804), .B(n9805), .Z(n170) );
  AND U10743 ( .A(n9806), .B(n9807), .Z(n9804) );
  XOR U10744 ( .A(n9805), .B(n9720), .Z(n9807) );
  XNOR U10745 ( .A(n9808), .B(n9809), .Z(n9720) );
  ANDN U10746 ( .B(n9810), .A(n9811), .Z(n9808) );
  XOR U10747 ( .A(n9809), .B(n9812), .Z(n9810) );
  XNOR U10748 ( .A(n9805), .B(n9722), .Z(n9806) );
  XOR U10749 ( .A(n9813), .B(n9814), .Z(n9722) );
  AND U10750 ( .A(n174), .B(n9815), .Z(n9813) );
  XOR U10751 ( .A(n9816), .B(n9814), .Z(n9815) );
  XNOR U10752 ( .A(n9817), .B(n9818), .Z(n9805) );
  AND U10753 ( .A(n9819), .B(n9820), .Z(n9817) );
  XNOR U10754 ( .A(n9818), .B(n9747), .Z(n9820) );
  XOR U10755 ( .A(n9811), .B(n9812), .Z(n9747) );
  XNOR U10756 ( .A(n9821), .B(n9822), .Z(n9812) );
  ANDN U10757 ( .B(n9823), .A(n9824), .Z(n9821) );
  XOR U10758 ( .A(n9825), .B(n9826), .Z(n9823) );
  XOR U10759 ( .A(n9827), .B(n9828), .Z(n9811) );
  XNOR U10760 ( .A(n9829), .B(n9830), .Z(n9828) );
  ANDN U10761 ( .B(n9831), .A(n9832), .Z(n9829) );
  XNOR U10762 ( .A(n9833), .B(n9834), .Z(n9831) );
  IV U10763 ( .A(n9809), .Z(n9827) );
  XOR U10764 ( .A(n9835), .B(n9836), .Z(n9809) );
  ANDN U10765 ( .B(n9837), .A(n9838), .Z(n9835) );
  XOR U10766 ( .A(n9836), .B(n9839), .Z(n9837) );
  XOR U10767 ( .A(n9818), .B(n9749), .Z(n9819) );
  XOR U10768 ( .A(n9840), .B(n9841), .Z(n9749) );
  AND U10769 ( .A(n174), .B(n9842), .Z(n9840) );
  XOR U10770 ( .A(n9843), .B(n9841), .Z(n9842) );
  XNOR U10771 ( .A(n9844), .B(n9845), .Z(n9818) );
  NAND U10772 ( .A(n9846), .B(n9847), .Z(n9845) );
  XOR U10773 ( .A(n9848), .B(n9797), .Z(n9847) );
  XOR U10774 ( .A(n9838), .B(n9839), .Z(n9797) );
  XOR U10775 ( .A(n9849), .B(n9826), .Z(n9839) );
  XOR U10776 ( .A(n9850), .B(n9851), .Z(n9826) );
  ANDN U10777 ( .B(n9852), .A(n9853), .Z(n9850) );
  XOR U10778 ( .A(n9851), .B(n9854), .Z(n9852) );
  IV U10779 ( .A(n9824), .Z(n9849) );
  XOR U10780 ( .A(n9822), .B(n9855), .Z(n9824) );
  XOR U10781 ( .A(n9856), .B(n9857), .Z(n9855) );
  ANDN U10782 ( .B(n9858), .A(n9859), .Z(n9856) );
  XOR U10783 ( .A(n9860), .B(n9857), .Z(n9858) );
  IV U10784 ( .A(n9825), .Z(n9822) );
  XOR U10785 ( .A(n9861), .B(n9862), .Z(n9825) );
  ANDN U10786 ( .B(n9863), .A(n9864), .Z(n9861) );
  XOR U10787 ( .A(n9862), .B(n9865), .Z(n9863) );
  XOR U10788 ( .A(n9866), .B(n9867), .Z(n9838) );
  XNOR U10789 ( .A(n9833), .B(n9868), .Z(n9867) );
  IV U10790 ( .A(n9836), .Z(n9868) );
  XOR U10791 ( .A(n9869), .B(n9870), .Z(n9836) );
  ANDN U10792 ( .B(n9871), .A(n9872), .Z(n9869) );
  XOR U10793 ( .A(n9870), .B(n9873), .Z(n9871) );
  XNOR U10794 ( .A(n9874), .B(n9875), .Z(n9833) );
  ANDN U10795 ( .B(n9876), .A(n9877), .Z(n9874) );
  XOR U10796 ( .A(n9875), .B(n9878), .Z(n9876) );
  IV U10797 ( .A(n9832), .Z(n9866) );
  XOR U10798 ( .A(n9830), .B(n9879), .Z(n9832) );
  XOR U10799 ( .A(n9880), .B(n9881), .Z(n9879) );
  ANDN U10800 ( .B(n9882), .A(n9883), .Z(n9880) );
  XOR U10801 ( .A(n9884), .B(n9881), .Z(n9882) );
  IV U10802 ( .A(n9834), .Z(n9830) );
  XOR U10803 ( .A(n9885), .B(n9886), .Z(n9834) );
  ANDN U10804 ( .B(n9887), .A(n9888), .Z(n9885) );
  XOR U10805 ( .A(n9889), .B(n9886), .Z(n9887) );
  IV U10806 ( .A(n9844), .Z(n9848) );
  XOR U10807 ( .A(n9844), .B(n9799), .Z(n9846) );
  XOR U10808 ( .A(n9890), .B(n9891), .Z(n9799) );
  AND U10809 ( .A(n174), .B(n9892), .Z(n9890) );
  XOR U10810 ( .A(n9893), .B(n9891), .Z(n9892) );
  NANDN U10811 ( .A(n9801), .B(n9803), .Z(n9844) );
  XOR U10812 ( .A(n9894), .B(n9895), .Z(n9803) );
  AND U10813 ( .A(n174), .B(n9896), .Z(n9894) );
  XOR U10814 ( .A(n9895), .B(n9897), .Z(n9896) );
  XNOR U10815 ( .A(n9898), .B(n9899), .Z(n174) );
  AND U10816 ( .A(n9900), .B(n9901), .Z(n9898) );
  XOR U10817 ( .A(n9899), .B(n9814), .Z(n9901) );
  XNOR U10818 ( .A(n9902), .B(n9903), .Z(n9814) );
  ANDN U10819 ( .B(n9904), .A(n9905), .Z(n9902) );
  XOR U10820 ( .A(n9903), .B(n9906), .Z(n9904) );
  XNOR U10821 ( .A(n9899), .B(n9816), .Z(n9900) );
  XOR U10822 ( .A(n9907), .B(n9908), .Z(n9816) );
  AND U10823 ( .A(n178), .B(n9909), .Z(n9907) );
  XOR U10824 ( .A(n9910), .B(n9908), .Z(n9909) );
  XNOR U10825 ( .A(n9911), .B(n9912), .Z(n9899) );
  AND U10826 ( .A(n9913), .B(n9914), .Z(n9911) );
  XNOR U10827 ( .A(n9912), .B(n9841), .Z(n9914) );
  XOR U10828 ( .A(n9905), .B(n9906), .Z(n9841) );
  XNOR U10829 ( .A(n9915), .B(n9916), .Z(n9906) );
  ANDN U10830 ( .B(n9917), .A(n9918), .Z(n9915) );
  XOR U10831 ( .A(n9919), .B(n9920), .Z(n9917) );
  XOR U10832 ( .A(n9921), .B(n9922), .Z(n9905) );
  XNOR U10833 ( .A(n9923), .B(n9924), .Z(n9922) );
  ANDN U10834 ( .B(n9925), .A(n9926), .Z(n9923) );
  XNOR U10835 ( .A(n9927), .B(n9928), .Z(n9925) );
  IV U10836 ( .A(n9903), .Z(n9921) );
  XOR U10837 ( .A(n9929), .B(n9930), .Z(n9903) );
  ANDN U10838 ( .B(n9931), .A(n9932), .Z(n9929) );
  XOR U10839 ( .A(n9930), .B(n9933), .Z(n9931) );
  XOR U10840 ( .A(n9912), .B(n9843), .Z(n9913) );
  XOR U10841 ( .A(n9934), .B(n9935), .Z(n9843) );
  AND U10842 ( .A(n178), .B(n9936), .Z(n9934) );
  XOR U10843 ( .A(n9937), .B(n9935), .Z(n9936) );
  XNOR U10844 ( .A(n9938), .B(n9939), .Z(n9912) );
  NAND U10845 ( .A(n9940), .B(n9941), .Z(n9939) );
  XOR U10846 ( .A(n9942), .B(n9891), .Z(n9941) );
  XOR U10847 ( .A(n9932), .B(n9933), .Z(n9891) );
  XOR U10848 ( .A(n9943), .B(n9920), .Z(n9933) );
  XOR U10849 ( .A(n9944), .B(n9945), .Z(n9920) );
  ANDN U10850 ( .B(n9946), .A(n9947), .Z(n9944) );
  XOR U10851 ( .A(n9945), .B(n9948), .Z(n9946) );
  IV U10852 ( .A(n9918), .Z(n9943) );
  XOR U10853 ( .A(n9916), .B(n9949), .Z(n9918) );
  XOR U10854 ( .A(n9950), .B(n9951), .Z(n9949) );
  ANDN U10855 ( .B(n9952), .A(n9953), .Z(n9950) );
  XOR U10856 ( .A(n9954), .B(n9951), .Z(n9952) );
  IV U10857 ( .A(n9919), .Z(n9916) );
  XOR U10858 ( .A(n9955), .B(n9956), .Z(n9919) );
  ANDN U10859 ( .B(n9957), .A(n9958), .Z(n9955) );
  XOR U10860 ( .A(n9956), .B(n9959), .Z(n9957) );
  XOR U10861 ( .A(n9960), .B(n9961), .Z(n9932) );
  XNOR U10862 ( .A(n9927), .B(n9962), .Z(n9961) );
  IV U10863 ( .A(n9930), .Z(n9962) );
  XOR U10864 ( .A(n9963), .B(n9964), .Z(n9930) );
  ANDN U10865 ( .B(n9965), .A(n9966), .Z(n9963) );
  XOR U10866 ( .A(n9964), .B(n9967), .Z(n9965) );
  XNOR U10867 ( .A(n9968), .B(n9969), .Z(n9927) );
  ANDN U10868 ( .B(n9970), .A(n9971), .Z(n9968) );
  XOR U10869 ( .A(n9969), .B(n9972), .Z(n9970) );
  IV U10870 ( .A(n9926), .Z(n9960) );
  XOR U10871 ( .A(n9924), .B(n9973), .Z(n9926) );
  XOR U10872 ( .A(n9974), .B(n9975), .Z(n9973) );
  ANDN U10873 ( .B(n9976), .A(n9977), .Z(n9974) );
  XOR U10874 ( .A(n9978), .B(n9975), .Z(n9976) );
  IV U10875 ( .A(n9928), .Z(n9924) );
  XOR U10876 ( .A(n9979), .B(n9980), .Z(n9928) );
  ANDN U10877 ( .B(n9981), .A(n9982), .Z(n9979) );
  XOR U10878 ( .A(n9983), .B(n9980), .Z(n9981) );
  IV U10879 ( .A(n9938), .Z(n9942) );
  XOR U10880 ( .A(n9938), .B(n9893), .Z(n9940) );
  XOR U10881 ( .A(n9984), .B(n9985), .Z(n9893) );
  AND U10882 ( .A(n178), .B(n9986), .Z(n9984) );
  XOR U10883 ( .A(n9987), .B(n9985), .Z(n9986) );
  NANDN U10884 ( .A(n9895), .B(n9897), .Z(n9938) );
  XOR U10885 ( .A(n9988), .B(n9989), .Z(n9897) );
  AND U10886 ( .A(n178), .B(n9990), .Z(n9988) );
  XOR U10887 ( .A(n9989), .B(n9991), .Z(n9990) );
  XNOR U10888 ( .A(n9992), .B(n9993), .Z(n178) );
  AND U10889 ( .A(n9994), .B(n9995), .Z(n9992) );
  XOR U10890 ( .A(n9993), .B(n9908), .Z(n9995) );
  XNOR U10891 ( .A(n9996), .B(n9997), .Z(n9908) );
  ANDN U10892 ( .B(n9998), .A(n9999), .Z(n9996) );
  XOR U10893 ( .A(n9997), .B(n10000), .Z(n9998) );
  XNOR U10894 ( .A(n9993), .B(n9910), .Z(n9994) );
  XOR U10895 ( .A(n10001), .B(n10002), .Z(n9910) );
  AND U10896 ( .A(n182), .B(n10003), .Z(n10001) );
  XOR U10897 ( .A(n10004), .B(n10002), .Z(n10003) );
  XNOR U10898 ( .A(n10005), .B(n10006), .Z(n9993) );
  AND U10899 ( .A(n10007), .B(n10008), .Z(n10005) );
  XNOR U10900 ( .A(n10006), .B(n9935), .Z(n10008) );
  XOR U10901 ( .A(n9999), .B(n10000), .Z(n9935) );
  XNOR U10902 ( .A(n10009), .B(n10010), .Z(n10000) );
  ANDN U10903 ( .B(n10011), .A(n10012), .Z(n10009) );
  XOR U10904 ( .A(n10013), .B(n10014), .Z(n10011) );
  XOR U10905 ( .A(n10015), .B(n10016), .Z(n9999) );
  XNOR U10906 ( .A(n10017), .B(n10018), .Z(n10016) );
  ANDN U10907 ( .B(n10019), .A(n10020), .Z(n10017) );
  XNOR U10908 ( .A(n10021), .B(n10022), .Z(n10019) );
  IV U10909 ( .A(n9997), .Z(n10015) );
  XOR U10910 ( .A(n10023), .B(n10024), .Z(n9997) );
  ANDN U10911 ( .B(n10025), .A(n10026), .Z(n10023) );
  XOR U10912 ( .A(n10024), .B(n10027), .Z(n10025) );
  XOR U10913 ( .A(n10006), .B(n9937), .Z(n10007) );
  XOR U10914 ( .A(n10028), .B(n10029), .Z(n9937) );
  AND U10915 ( .A(n182), .B(n10030), .Z(n10028) );
  XOR U10916 ( .A(n10031), .B(n10029), .Z(n10030) );
  XNOR U10917 ( .A(n10032), .B(n10033), .Z(n10006) );
  NAND U10918 ( .A(n10034), .B(n10035), .Z(n10033) );
  XOR U10919 ( .A(n10036), .B(n9985), .Z(n10035) );
  XOR U10920 ( .A(n10026), .B(n10027), .Z(n9985) );
  XOR U10921 ( .A(n10037), .B(n10014), .Z(n10027) );
  XOR U10922 ( .A(n10038), .B(n10039), .Z(n10014) );
  ANDN U10923 ( .B(n10040), .A(n10041), .Z(n10038) );
  XOR U10924 ( .A(n10039), .B(n10042), .Z(n10040) );
  IV U10925 ( .A(n10012), .Z(n10037) );
  XOR U10926 ( .A(n10010), .B(n10043), .Z(n10012) );
  XOR U10927 ( .A(n10044), .B(n10045), .Z(n10043) );
  ANDN U10928 ( .B(n10046), .A(n10047), .Z(n10044) );
  XOR U10929 ( .A(n10048), .B(n10045), .Z(n10046) );
  IV U10930 ( .A(n10013), .Z(n10010) );
  XOR U10931 ( .A(n10049), .B(n10050), .Z(n10013) );
  ANDN U10932 ( .B(n10051), .A(n10052), .Z(n10049) );
  XOR U10933 ( .A(n10050), .B(n10053), .Z(n10051) );
  XOR U10934 ( .A(n10054), .B(n10055), .Z(n10026) );
  XNOR U10935 ( .A(n10021), .B(n10056), .Z(n10055) );
  IV U10936 ( .A(n10024), .Z(n10056) );
  XOR U10937 ( .A(n10057), .B(n10058), .Z(n10024) );
  ANDN U10938 ( .B(n10059), .A(n10060), .Z(n10057) );
  XOR U10939 ( .A(n10058), .B(n10061), .Z(n10059) );
  XNOR U10940 ( .A(n10062), .B(n10063), .Z(n10021) );
  ANDN U10941 ( .B(n10064), .A(n10065), .Z(n10062) );
  XOR U10942 ( .A(n10063), .B(n10066), .Z(n10064) );
  IV U10943 ( .A(n10020), .Z(n10054) );
  XOR U10944 ( .A(n10018), .B(n10067), .Z(n10020) );
  XOR U10945 ( .A(n10068), .B(n10069), .Z(n10067) );
  ANDN U10946 ( .B(n10070), .A(n10071), .Z(n10068) );
  XOR U10947 ( .A(n10072), .B(n10069), .Z(n10070) );
  IV U10948 ( .A(n10022), .Z(n10018) );
  XOR U10949 ( .A(n10073), .B(n10074), .Z(n10022) );
  ANDN U10950 ( .B(n10075), .A(n10076), .Z(n10073) );
  XOR U10951 ( .A(n10077), .B(n10074), .Z(n10075) );
  IV U10952 ( .A(n10032), .Z(n10036) );
  XOR U10953 ( .A(n10032), .B(n9987), .Z(n10034) );
  XOR U10954 ( .A(n10078), .B(n10079), .Z(n9987) );
  AND U10955 ( .A(n182), .B(n10080), .Z(n10078) );
  XOR U10956 ( .A(n10081), .B(n10079), .Z(n10080) );
  NANDN U10957 ( .A(n9989), .B(n9991), .Z(n10032) );
  XOR U10958 ( .A(n10082), .B(n10083), .Z(n9991) );
  AND U10959 ( .A(n182), .B(n10084), .Z(n10082) );
  XOR U10960 ( .A(n10083), .B(n10085), .Z(n10084) );
  XNOR U10961 ( .A(n10086), .B(n10087), .Z(n182) );
  AND U10962 ( .A(n10088), .B(n10089), .Z(n10086) );
  XOR U10963 ( .A(n10087), .B(n10002), .Z(n10089) );
  XNOR U10964 ( .A(n10090), .B(n10091), .Z(n10002) );
  ANDN U10965 ( .B(n10092), .A(n10093), .Z(n10090) );
  XOR U10966 ( .A(n10091), .B(n10094), .Z(n10092) );
  XNOR U10967 ( .A(n10087), .B(n10004), .Z(n10088) );
  XOR U10968 ( .A(n10095), .B(n10096), .Z(n10004) );
  AND U10969 ( .A(n186), .B(n10097), .Z(n10095) );
  XOR U10970 ( .A(n10098), .B(n10096), .Z(n10097) );
  XNOR U10971 ( .A(n10099), .B(n10100), .Z(n10087) );
  AND U10972 ( .A(n10101), .B(n10102), .Z(n10099) );
  XNOR U10973 ( .A(n10100), .B(n10029), .Z(n10102) );
  XOR U10974 ( .A(n10093), .B(n10094), .Z(n10029) );
  XNOR U10975 ( .A(n10103), .B(n10104), .Z(n10094) );
  ANDN U10976 ( .B(n10105), .A(n10106), .Z(n10103) );
  XOR U10977 ( .A(n10107), .B(n10108), .Z(n10105) );
  XOR U10978 ( .A(n10109), .B(n10110), .Z(n10093) );
  XNOR U10979 ( .A(n10111), .B(n10112), .Z(n10110) );
  ANDN U10980 ( .B(n10113), .A(n10114), .Z(n10111) );
  XNOR U10981 ( .A(n10115), .B(n10116), .Z(n10113) );
  IV U10982 ( .A(n10091), .Z(n10109) );
  XOR U10983 ( .A(n10117), .B(n10118), .Z(n10091) );
  ANDN U10984 ( .B(n10119), .A(n10120), .Z(n10117) );
  XOR U10985 ( .A(n10118), .B(n10121), .Z(n10119) );
  XOR U10986 ( .A(n10100), .B(n10031), .Z(n10101) );
  XOR U10987 ( .A(n10122), .B(n10123), .Z(n10031) );
  AND U10988 ( .A(n186), .B(n10124), .Z(n10122) );
  XOR U10989 ( .A(n10125), .B(n10123), .Z(n10124) );
  XNOR U10990 ( .A(n10126), .B(n10127), .Z(n10100) );
  NAND U10991 ( .A(n10128), .B(n10129), .Z(n10127) );
  XOR U10992 ( .A(n10130), .B(n10079), .Z(n10129) );
  XOR U10993 ( .A(n10120), .B(n10121), .Z(n10079) );
  XOR U10994 ( .A(n10131), .B(n10108), .Z(n10121) );
  XOR U10995 ( .A(n10132), .B(n10133), .Z(n10108) );
  ANDN U10996 ( .B(n10134), .A(n10135), .Z(n10132) );
  XOR U10997 ( .A(n10133), .B(n10136), .Z(n10134) );
  IV U10998 ( .A(n10106), .Z(n10131) );
  XOR U10999 ( .A(n10104), .B(n10137), .Z(n10106) );
  XOR U11000 ( .A(n10138), .B(n10139), .Z(n10137) );
  ANDN U11001 ( .B(n10140), .A(n10141), .Z(n10138) );
  XOR U11002 ( .A(n10142), .B(n10139), .Z(n10140) );
  IV U11003 ( .A(n10107), .Z(n10104) );
  XOR U11004 ( .A(n10143), .B(n10144), .Z(n10107) );
  ANDN U11005 ( .B(n10145), .A(n10146), .Z(n10143) );
  XOR U11006 ( .A(n10144), .B(n10147), .Z(n10145) );
  XOR U11007 ( .A(n10148), .B(n10149), .Z(n10120) );
  XNOR U11008 ( .A(n10115), .B(n10150), .Z(n10149) );
  IV U11009 ( .A(n10118), .Z(n10150) );
  XOR U11010 ( .A(n10151), .B(n10152), .Z(n10118) );
  ANDN U11011 ( .B(n10153), .A(n10154), .Z(n10151) );
  XOR U11012 ( .A(n10152), .B(n10155), .Z(n10153) );
  XNOR U11013 ( .A(n10156), .B(n10157), .Z(n10115) );
  ANDN U11014 ( .B(n10158), .A(n10159), .Z(n10156) );
  XOR U11015 ( .A(n10157), .B(n10160), .Z(n10158) );
  IV U11016 ( .A(n10114), .Z(n10148) );
  XOR U11017 ( .A(n10112), .B(n10161), .Z(n10114) );
  XOR U11018 ( .A(n10162), .B(n10163), .Z(n10161) );
  ANDN U11019 ( .B(n10164), .A(n10165), .Z(n10162) );
  XOR U11020 ( .A(n10166), .B(n10163), .Z(n10164) );
  IV U11021 ( .A(n10116), .Z(n10112) );
  XOR U11022 ( .A(n10167), .B(n10168), .Z(n10116) );
  ANDN U11023 ( .B(n10169), .A(n10170), .Z(n10167) );
  XOR U11024 ( .A(n10171), .B(n10168), .Z(n10169) );
  IV U11025 ( .A(n10126), .Z(n10130) );
  XOR U11026 ( .A(n10126), .B(n10081), .Z(n10128) );
  XOR U11027 ( .A(n10172), .B(n10173), .Z(n10081) );
  AND U11028 ( .A(n186), .B(n10174), .Z(n10172) );
  XOR U11029 ( .A(n10175), .B(n10173), .Z(n10174) );
  NANDN U11030 ( .A(n10083), .B(n10085), .Z(n10126) );
  XOR U11031 ( .A(n10176), .B(n10177), .Z(n10085) );
  AND U11032 ( .A(n186), .B(n10178), .Z(n10176) );
  XOR U11033 ( .A(n10177), .B(n10179), .Z(n10178) );
  XNOR U11034 ( .A(n10180), .B(n10181), .Z(n186) );
  AND U11035 ( .A(n10182), .B(n10183), .Z(n10180) );
  XOR U11036 ( .A(n10181), .B(n10096), .Z(n10183) );
  XNOR U11037 ( .A(n10184), .B(n10185), .Z(n10096) );
  ANDN U11038 ( .B(n10186), .A(n10187), .Z(n10184) );
  XOR U11039 ( .A(n10185), .B(n10188), .Z(n10186) );
  XNOR U11040 ( .A(n10181), .B(n10098), .Z(n10182) );
  XOR U11041 ( .A(n10189), .B(n10190), .Z(n10098) );
  AND U11042 ( .A(n190), .B(n10191), .Z(n10189) );
  XOR U11043 ( .A(n10192), .B(n10190), .Z(n10191) );
  XNOR U11044 ( .A(n10193), .B(n10194), .Z(n10181) );
  AND U11045 ( .A(n10195), .B(n10196), .Z(n10193) );
  XNOR U11046 ( .A(n10194), .B(n10123), .Z(n10196) );
  XOR U11047 ( .A(n10187), .B(n10188), .Z(n10123) );
  XNOR U11048 ( .A(n10197), .B(n10198), .Z(n10188) );
  ANDN U11049 ( .B(n10199), .A(n10200), .Z(n10197) );
  XOR U11050 ( .A(n10201), .B(n10202), .Z(n10199) );
  XOR U11051 ( .A(n10203), .B(n10204), .Z(n10187) );
  XNOR U11052 ( .A(n10205), .B(n10206), .Z(n10204) );
  ANDN U11053 ( .B(n10207), .A(n10208), .Z(n10205) );
  XNOR U11054 ( .A(n10209), .B(n10210), .Z(n10207) );
  IV U11055 ( .A(n10185), .Z(n10203) );
  XOR U11056 ( .A(n10211), .B(n10212), .Z(n10185) );
  ANDN U11057 ( .B(n10213), .A(n10214), .Z(n10211) );
  XOR U11058 ( .A(n10212), .B(n10215), .Z(n10213) );
  XOR U11059 ( .A(n10194), .B(n10125), .Z(n10195) );
  XOR U11060 ( .A(n10216), .B(n10217), .Z(n10125) );
  AND U11061 ( .A(n190), .B(n10218), .Z(n10216) );
  XOR U11062 ( .A(n10219), .B(n10217), .Z(n10218) );
  XNOR U11063 ( .A(n10220), .B(n10221), .Z(n10194) );
  NAND U11064 ( .A(n10222), .B(n10223), .Z(n10221) );
  XOR U11065 ( .A(n10224), .B(n10173), .Z(n10223) );
  XOR U11066 ( .A(n10214), .B(n10215), .Z(n10173) );
  XOR U11067 ( .A(n10225), .B(n10202), .Z(n10215) );
  XOR U11068 ( .A(n10226), .B(n10227), .Z(n10202) );
  ANDN U11069 ( .B(n10228), .A(n10229), .Z(n10226) );
  XOR U11070 ( .A(n10227), .B(n10230), .Z(n10228) );
  IV U11071 ( .A(n10200), .Z(n10225) );
  XOR U11072 ( .A(n10198), .B(n10231), .Z(n10200) );
  XOR U11073 ( .A(n10232), .B(n10233), .Z(n10231) );
  ANDN U11074 ( .B(n10234), .A(n10235), .Z(n10232) );
  XOR U11075 ( .A(n10236), .B(n10233), .Z(n10234) );
  IV U11076 ( .A(n10201), .Z(n10198) );
  XOR U11077 ( .A(n10237), .B(n10238), .Z(n10201) );
  ANDN U11078 ( .B(n10239), .A(n10240), .Z(n10237) );
  XOR U11079 ( .A(n10238), .B(n10241), .Z(n10239) );
  XOR U11080 ( .A(n10242), .B(n10243), .Z(n10214) );
  XNOR U11081 ( .A(n10209), .B(n10244), .Z(n10243) );
  IV U11082 ( .A(n10212), .Z(n10244) );
  XOR U11083 ( .A(n10245), .B(n10246), .Z(n10212) );
  ANDN U11084 ( .B(n10247), .A(n10248), .Z(n10245) );
  XOR U11085 ( .A(n10246), .B(n10249), .Z(n10247) );
  XNOR U11086 ( .A(n10250), .B(n10251), .Z(n10209) );
  ANDN U11087 ( .B(n10252), .A(n10253), .Z(n10250) );
  XOR U11088 ( .A(n10251), .B(n10254), .Z(n10252) );
  IV U11089 ( .A(n10208), .Z(n10242) );
  XOR U11090 ( .A(n10206), .B(n10255), .Z(n10208) );
  XOR U11091 ( .A(n10256), .B(n10257), .Z(n10255) );
  ANDN U11092 ( .B(n10258), .A(n10259), .Z(n10256) );
  XOR U11093 ( .A(n10260), .B(n10257), .Z(n10258) );
  IV U11094 ( .A(n10210), .Z(n10206) );
  XOR U11095 ( .A(n10261), .B(n10262), .Z(n10210) );
  ANDN U11096 ( .B(n10263), .A(n10264), .Z(n10261) );
  XOR U11097 ( .A(n10265), .B(n10262), .Z(n10263) );
  IV U11098 ( .A(n10220), .Z(n10224) );
  XOR U11099 ( .A(n10220), .B(n10175), .Z(n10222) );
  XOR U11100 ( .A(n10266), .B(n10267), .Z(n10175) );
  AND U11101 ( .A(n190), .B(n10268), .Z(n10266) );
  XOR U11102 ( .A(n10269), .B(n10267), .Z(n10268) );
  NANDN U11103 ( .A(n10177), .B(n10179), .Z(n10220) );
  XOR U11104 ( .A(n10270), .B(n10271), .Z(n10179) );
  AND U11105 ( .A(n190), .B(n10272), .Z(n10270) );
  XOR U11106 ( .A(n10271), .B(n10273), .Z(n10272) );
  XNOR U11107 ( .A(n10274), .B(n10275), .Z(n190) );
  AND U11108 ( .A(n10276), .B(n10277), .Z(n10274) );
  XOR U11109 ( .A(n10275), .B(n10190), .Z(n10277) );
  XNOR U11110 ( .A(n10278), .B(n10279), .Z(n10190) );
  ANDN U11111 ( .B(n10280), .A(n10281), .Z(n10278) );
  XOR U11112 ( .A(n10279), .B(n10282), .Z(n10280) );
  XNOR U11113 ( .A(n10275), .B(n10192), .Z(n10276) );
  XOR U11114 ( .A(n10283), .B(n10284), .Z(n10192) );
  AND U11115 ( .A(n194), .B(n10285), .Z(n10283) );
  XOR U11116 ( .A(n10286), .B(n10284), .Z(n10285) );
  XNOR U11117 ( .A(n10287), .B(n10288), .Z(n10275) );
  AND U11118 ( .A(n10289), .B(n10290), .Z(n10287) );
  XNOR U11119 ( .A(n10288), .B(n10217), .Z(n10290) );
  XOR U11120 ( .A(n10281), .B(n10282), .Z(n10217) );
  XNOR U11121 ( .A(n10291), .B(n10292), .Z(n10282) );
  ANDN U11122 ( .B(n10293), .A(n10294), .Z(n10291) );
  XOR U11123 ( .A(n10295), .B(n10296), .Z(n10293) );
  XOR U11124 ( .A(n10297), .B(n10298), .Z(n10281) );
  XNOR U11125 ( .A(n10299), .B(n10300), .Z(n10298) );
  ANDN U11126 ( .B(n10301), .A(n10302), .Z(n10299) );
  XNOR U11127 ( .A(n10303), .B(n10304), .Z(n10301) );
  IV U11128 ( .A(n10279), .Z(n10297) );
  XOR U11129 ( .A(n10305), .B(n10306), .Z(n10279) );
  ANDN U11130 ( .B(n10307), .A(n10308), .Z(n10305) );
  XOR U11131 ( .A(n10306), .B(n10309), .Z(n10307) );
  XOR U11132 ( .A(n10288), .B(n10219), .Z(n10289) );
  XOR U11133 ( .A(n10310), .B(n10311), .Z(n10219) );
  AND U11134 ( .A(n194), .B(n10312), .Z(n10310) );
  XOR U11135 ( .A(n10313), .B(n10311), .Z(n10312) );
  XNOR U11136 ( .A(n10314), .B(n10315), .Z(n10288) );
  NAND U11137 ( .A(n10316), .B(n10317), .Z(n10315) );
  XOR U11138 ( .A(n10318), .B(n10267), .Z(n10317) );
  XOR U11139 ( .A(n10308), .B(n10309), .Z(n10267) );
  XOR U11140 ( .A(n10319), .B(n10296), .Z(n10309) );
  XOR U11141 ( .A(n10320), .B(n10321), .Z(n10296) );
  ANDN U11142 ( .B(n10322), .A(n10323), .Z(n10320) );
  XOR U11143 ( .A(n10321), .B(n10324), .Z(n10322) );
  IV U11144 ( .A(n10294), .Z(n10319) );
  XOR U11145 ( .A(n10292), .B(n10325), .Z(n10294) );
  XOR U11146 ( .A(n10326), .B(n10327), .Z(n10325) );
  ANDN U11147 ( .B(n10328), .A(n10329), .Z(n10326) );
  XOR U11148 ( .A(n10330), .B(n10327), .Z(n10328) );
  IV U11149 ( .A(n10295), .Z(n10292) );
  XOR U11150 ( .A(n10331), .B(n10332), .Z(n10295) );
  ANDN U11151 ( .B(n10333), .A(n10334), .Z(n10331) );
  XOR U11152 ( .A(n10332), .B(n10335), .Z(n10333) );
  XOR U11153 ( .A(n10336), .B(n10337), .Z(n10308) );
  XNOR U11154 ( .A(n10303), .B(n10338), .Z(n10337) );
  IV U11155 ( .A(n10306), .Z(n10338) );
  XOR U11156 ( .A(n10339), .B(n10340), .Z(n10306) );
  ANDN U11157 ( .B(n10341), .A(n10342), .Z(n10339) );
  XOR U11158 ( .A(n10340), .B(n10343), .Z(n10341) );
  XNOR U11159 ( .A(n10344), .B(n10345), .Z(n10303) );
  ANDN U11160 ( .B(n10346), .A(n10347), .Z(n10344) );
  XOR U11161 ( .A(n10345), .B(n10348), .Z(n10346) );
  IV U11162 ( .A(n10302), .Z(n10336) );
  XOR U11163 ( .A(n10300), .B(n10349), .Z(n10302) );
  XOR U11164 ( .A(n10350), .B(n10351), .Z(n10349) );
  ANDN U11165 ( .B(n10352), .A(n10353), .Z(n10350) );
  XOR U11166 ( .A(n10354), .B(n10351), .Z(n10352) );
  IV U11167 ( .A(n10304), .Z(n10300) );
  XOR U11168 ( .A(n10355), .B(n10356), .Z(n10304) );
  ANDN U11169 ( .B(n10357), .A(n10358), .Z(n10355) );
  XOR U11170 ( .A(n10359), .B(n10356), .Z(n10357) );
  IV U11171 ( .A(n10314), .Z(n10318) );
  XOR U11172 ( .A(n10314), .B(n10269), .Z(n10316) );
  XOR U11173 ( .A(n10360), .B(n10361), .Z(n10269) );
  AND U11174 ( .A(n194), .B(n10362), .Z(n10360) );
  XOR U11175 ( .A(n10363), .B(n10361), .Z(n10362) );
  NANDN U11176 ( .A(n10271), .B(n10273), .Z(n10314) );
  XOR U11177 ( .A(n10364), .B(n10365), .Z(n10273) );
  AND U11178 ( .A(n194), .B(n10366), .Z(n10364) );
  XOR U11179 ( .A(n10365), .B(n10367), .Z(n10366) );
  XNOR U11180 ( .A(n10368), .B(n10369), .Z(n194) );
  AND U11181 ( .A(n10370), .B(n10371), .Z(n10368) );
  XOR U11182 ( .A(n10369), .B(n10284), .Z(n10371) );
  XNOR U11183 ( .A(n10372), .B(n10373), .Z(n10284) );
  ANDN U11184 ( .B(n10374), .A(n10375), .Z(n10372) );
  XOR U11185 ( .A(n10373), .B(n10376), .Z(n10374) );
  XNOR U11186 ( .A(n10369), .B(n10286), .Z(n10370) );
  XOR U11187 ( .A(n10377), .B(n10378), .Z(n10286) );
  AND U11188 ( .A(n198), .B(n10379), .Z(n10377) );
  XOR U11189 ( .A(n10380), .B(n10378), .Z(n10379) );
  XNOR U11190 ( .A(n10381), .B(n10382), .Z(n10369) );
  AND U11191 ( .A(n10383), .B(n10384), .Z(n10381) );
  XNOR U11192 ( .A(n10382), .B(n10311), .Z(n10384) );
  XOR U11193 ( .A(n10375), .B(n10376), .Z(n10311) );
  XNOR U11194 ( .A(n10385), .B(n10386), .Z(n10376) );
  ANDN U11195 ( .B(n10387), .A(n10388), .Z(n10385) );
  XOR U11196 ( .A(n10389), .B(n10390), .Z(n10387) );
  XOR U11197 ( .A(n10391), .B(n10392), .Z(n10375) );
  XNOR U11198 ( .A(n10393), .B(n10394), .Z(n10392) );
  ANDN U11199 ( .B(n10395), .A(n10396), .Z(n10393) );
  XNOR U11200 ( .A(n10397), .B(n10398), .Z(n10395) );
  IV U11201 ( .A(n10373), .Z(n10391) );
  XOR U11202 ( .A(n10399), .B(n10400), .Z(n10373) );
  ANDN U11203 ( .B(n10401), .A(n10402), .Z(n10399) );
  XOR U11204 ( .A(n10400), .B(n10403), .Z(n10401) );
  XOR U11205 ( .A(n10382), .B(n10313), .Z(n10383) );
  XOR U11206 ( .A(n10404), .B(n10405), .Z(n10313) );
  AND U11207 ( .A(n198), .B(n10406), .Z(n10404) );
  XOR U11208 ( .A(n10407), .B(n10405), .Z(n10406) );
  XNOR U11209 ( .A(n10408), .B(n10409), .Z(n10382) );
  NAND U11210 ( .A(n10410), .B(n10411), .Z(n10409) );
  XOR U11211 ( .A(n10412), .B(n10361), .Z(n10411) );
  XOR U11212 ( .A(n10402), .B(n10403), .Z(n10361) );
  XOR U11213 ( .A(n10413), .B(n10390), .Z(n10403) );
  XOR U11214 ( .A(n10414), .B(n10415), .Z(n10390) );
  ANDN U11215 ( .B(n10416), .A(n10417), .Z(n10414) );
  XOR U11216 ( .A(n10415), .B(n10418), .Z(n10416) );
  IV U11217 ( .A(n10388), .Z(n10413) );
  XOR U11218 ( .A(n10386), .B(n10419), .Z(n10388) );
  XOR U11219 ( .A(n10420), .B(n10421), .Z(n10419) );
  ANDN U11220 ( .B(n10422), .A(n10423), .Z(n10420) );
  XOR U11221 ( .A(n10424), .B(n10421), .Z(n10422) );
  IV U11222 ( .A(n10389), .Z(n10386) );
  XOR U11223 ( .A(n10425), .B(n10426), .Z(n10389) );
  ANDN U11224 ( .B(n10427), .A(n10428), .Z(n10425) );
  XOR U11225 ( .A(n10426), .B(n10429), .Z(n10427) );
  XOR U11226 ( .A(n10430), .B(n10431), .Z(n10402) );
  XNOR U11227 ( .A(n10397), .B(n10432), .Z(n10431) );
  IV U11228 ( .A(n10400), .Z(n10432) );
  XOR U11229 ( .A(n10433), .B(n10434), .Z(n10400) );
  ANDN U11230 ( .B(n10435), .A(n10436), .Z(n10433) );
  XOR U11231 ( .A(n10434), .B(n10437), .Z(n10435) );
  XNOR U11232 ( .A(n10438), .B(n10439), .Z(n10397) );
  ANDN U11233 ( .B(n10440), .A(n10441), .Z(n10438) );
  XOR U11234 ( .A(n10439), .B(n10442), .Z(n10440) );
  IV U11235 ( .A(n10396), .Z(n10430) );
  XOR U11236 ( .A(n10394), .B(n10443), .Z(n10396) );
  XOR U11237 ( .A(n10444), .B(n10445), .Z(n10443) );
  ANDN U11238 ( .B(n10446), .A(n10447), .Z(n10444) );
  XOR U11239 ( .A(n10448), .B(n10445), .Z(n10446) );
  IV U11240 ( .A(n10398), .Z(n10394) );
  XOR U11241 ( .A(n10449), .B(n10450), .Z(n10398) );
  ANDN U11242 ( .B(n10451), .A(n10452), .Z(n10449) );
  XOR U11243 ( .A(n10453), .B(n10450), .Z(n10451) );
  IV U11244 ( .A(n10408), .Z(n10412) );
  XOR U11245 ( .A(n10408), .B(n10363), .Z(n10410) );
  XOR U11246 ( .A(n10454), .B(n10455), .Z(n10363) );
  AND U11247 ( .A(n198), .B(n10456), .Z(n10454) );
  XOR U11248 ( .A(n10457), .B(n10455), .Z(n10456) );
  NANDN U11249 ( .A(n10365), .B(n10367), .Z(n10408) );
  XOR U11250 ( .A(n10458), .B(n10459), .Z(n10367) );
  AND U11251 ( .A(n198), .B(n10460), .Z(n10458) );
  XOR U11252 ( .A(n10459), .B(n10461), .Z(n10460) );
  XNOR U11253 ( .A(n10462), .B(n10463), .Z(n198) );
  AND U11254 ( .A(n10464), .B(n10465), .Z(n10462) );
  XOR U11255 ( .A(n10463), .B(n10378), .Z(n10465) );
  XNOR U11256 ( .A(n10466), .B(n10467), .Z(n10378) );
  ANDN U11257 ( .B(n10468), .A(n10469), .Z(n10466) );
  XOR U11258 ( .A(n10467), .B(n10470), .Z(n10468) );
  XNOR U11259 ( .A(n10463), .B(n10380), .Z(n10464) );
  XOR U11260 ( .A(n10471), .B(n10472), .Z(n10380) );
  AND U11261 ( .A(n202), .B(n10473), .Z(n10471) );
  XOR U11262 ( .A(n10474), .B(n10472), .Z(n10473) );
  XNOR U11263 ( .A(n10475), .B(n10476), .Z(n10463) );
  AND U11264 ( .A(n10477), .B(n10478), .Z(n10475) );
  XNOR U11265 ( .A(n10476), .B(n10405), .Z(n10478) );
  XOR U11266 ( .A(n10469), .B(n10470), .Z(n10405) );
  XNOR U11267 ( .A(n10479), .B(n10480), .Z(n10470) );
  ANDN U11268 ( .B(n10481), .A(n10482), .Z(n10479) );
  XOR U11269 ( .A(n10483), .B(n10484), .Z(n10481) );
  XOR U11270 ( .A(n10485), .B(n10486), .Z(n10469) );
  XNOR U11271 ( .A(n10487), .B(n10488), .Z(n10486) );
  ANDN U11272 ( .B(n10489), .A(n10490), .Z(n10487) );
  XNOR U11273 ( .A(n10491), .B(n10492), .Z(n10489) );
  IV U11274 ( .A(n10467), .Z(n10485) );
  XOR U11275 ( .A(n10493), .B(n10494), .Z(n10467) );
  ANDN U11276 ( .B(n10495), .A(n10496), .Z(n10493) );
  XOR U11277 ( .A(n10494), .B(n10497), .Z(n10495) );
  XOR U11278 ( .A(n10476), .B(n10407), .Z(n10477) );
  XOR U11279 ( .A(n10498), .B(n10499), .Z(n10407) );
  AND U11280 ( .A(n202), .B(n10500), .Z(n10498) );
  XOR U11281 ( .A(n10501), .B(n10499), .Z(n10500) );
  XNOR U11282 ( .A(n10502), .B(n10503), .Z(n10476) );
  NAND U11283 ( .A(n10504), .B(n10505), .Z(n10503) );
  XOR U11284 ( .A(n10506), .B(n10455), .Z(n10505) );
  XOR U11285 ( .A(n10496), .B(n10497), .Z(n10455) );
  XOR U11286 ( .A(n10507), .B(n10484), .Z(n10497) );
  XOR U11287 ( .A(n10508), .B(n10509), .Z(n10484) );
  ANDN U11288 ( .B(n10510), .A(n10511), .Z(n10508) );
  XOR U11289 ( .A(n10509), .B(n10512), .Z(n10510) );
  IV U11290 ( .A(n10482), .Z(n10507) );
  XOR U11291 ( .A(n10480), .B(n10513), .Z(n10482) );
  XOR U11292 ( .A(n10514), .B(n10515), .Z(n10513) );
  ANDN U11293 ( .B(n10516), .A(n10517), .Z(n10514) );
  XOR U11294 ( .A(n10518), .B(n10515), .Z(n10516) );
  IV U11295 ( .A(n10483), .Z(n10480) );
  XOR U11296 ( .A(n10519), .B(n10520), .Z(n10483) );
  ANDN U11297 ( .B(n10521), .A(n10522), .Z(n10519) );
  XOR U11298 ( .A(n10520), .B(n10523), .Z(n10521) );
  XOR U11299 ( .A(n10524), .B(n10525), .Z(n10496) );
  XNOR U11300 ( .A(n10491), .B(n10526), .Z(n10525) );
  IV U11301 ( .A(n10494), .Z(n10526) );
  XOR U11302 ( .A(n10527), .B(n10528), .Z(n10494) );
  ANDN U11303 ( .B(n10529), .A(n10530), .Z(n10527) );
  XOR U11304 ( .A(n10528), .B(n10531), .Z(n10529) );
  XNOR U11305 ( .A(n10532), .B(n10533), .Z(n10491) );
  ANDN U11306 ( .B(n10534), .A(n10535), .Z(n10532) );
  XOR U11307 ( .A(n10533), .B(n10536), .Z(n10534) );
  IV U11308 ( .A(n10490), .Z(n10524) );
  XOR U11309 ( .A(n10488), .B(n10537), .Z(n10490) );
  XOR U11310 ( .A(n10538), .B(n10539), .Z(n10537) );
  ANDN U11311 ( .B(n10540), .A(n10541), .Z(n10538) );
  XOR U11312 ( .A(n10542), .B(n10539), .Z(n10540) );
  IV U11313 ( .A(n10492), .Z(n10488) );
  XOR U11314 ( .A(n10543), .B(n10544), .Z(n10492) );
  ANDN U11315 ( .B(n10545), .A(n10546), .Z(n10543) );
  XOR U11316 ( .A(n10547), .B(n10544), .Z(n10545) );
  IV U11317 ( .A(n10502), .Z(n10506) );
  XOR U11318 ( .A(n10502), .B(n10457), .Z(n10504) );
  XOR U11319 ( .A(n10548), .B(n10549), .Z(n10457) );
  AND U11320 ( .A(n202), .B(n10550), .Z(n10548) );
  XOR U11321 ( .A(n10551), .B(n10549), .Z(n10550) );
  NANDN U11322 ( .A(n10459), .B(n10461), .Z(n10502) );
  XOR U11323 ( .A(n10552), .B(n10553), .Z(n10461) );
  AND U11324 ( .A(n202), .B(n10554), .Z(n10552) );
  XOR U11325 ( .A(n10553), .B(n10555), .Z(n10554) );
  XNOR U11326 ( .A(n10556), .B(n10557), .Z(n202) );
  AND U11327 ( .A(n10558), .B(n10559), .Z(n10556) );
  XOR U11328 ( .A(n10557), .B(n10472), .Z(n10559) );
  XNOR U11329 ( .A(n10560), .B(n10561), .Z(n10472) );
  ANDN U11330 ( .B(n10562), .A(n10563), .Z(n10560) );
  XOR U11331 ( .A(n10561), .B(n10564), .Z(n10562) );
  XNOR U11332 ( .A(n10557), .B(n10474), .Z(n10558) );
  XOR U11333 ( .A(n10565), .B(n10566), .Z(n10474) );
  AND U11334 ( .A(n206), .B(n10567), .Z(n10565) );
  XOR U11335 ( .A(n10568), .B(n10566), .Z(n10567) );
  XNOR U11336 ( .A(n10569), .B(n10570), .Z(n10557) );
  AND U11337 ( .A(n10571), .B(n10572), .Z(n10569) );
  XNOR U11338 ( .A(n10570), .B(n10499), .Z(n10572) );
  XOR U11339 ( .A(n10563), .B(n10564), .Z(n10499) );
  XNOR U11340 ( .A(n10573), .B(n10574), .Z(n10564) );
  ANDN U11341 ( .B(n10575), .A(n10576), .Z(n10573) );
  XOR U11342 ( .A(n10577), .B(n10578), .Z(n10575) );
  XOR U11343 ( .A(n10579), .B(n10580), .Z(n10563) );
  XNOR U11344 ( .A(n10581), .B(n10582), .Z(n10580) );
  ANDN U11345 ( .B(n10583), .A(n10584), .Z(n10581) );
  XNOR U11346 ( .A(n10585), .B(n10586), .Z(n10583) );
  IV U11347 ( .A(n10561), .Z(n10579) );
  XOR U11348 ( .A(n10587), .B(n10588), .Z(n10561) );
  ANDN U11349 ( .B(n10589), .A(n10590), .Z(n10587) );
  XOR U11350 ( .A(n10588), .B(n10591), .Z(n10589) );
  XOR U11351 ( .A(n10570), .B(n10501), .Z(n10571) );
  XOR U11352 ( .A(n10592), .B(n10593), .Z(n10501) );
  AND U11353 ( .A(n206), .B(n10594), .Z(n10592) );
  XOR U11354 ( .A(n10595), .B(n10593), .Z(n10594) );
  XNOR U11355 ( .A(n10596), .B(n10597), .Z(n10570) );
  NAND U11356 ( .A(n10598), .B(n10599), .Z(n10597) );
  XOR U11357 ( .A(n10600), .B(n10549), .Z(n10599) );
  XOR U11358 ( .A(n10590), .B(n10591), .Z(n10549) );
  XOR U11359 ( .A(n10601), .B(n10578), .Z(n10591) );
  XOR U11360 ( .A(n10602), .B(n10603), .Z(n10578) );
  ANDN U11361 ( .B(n10604), .A(n10605), .Z(n10602) );
  XOR U11362 ( .A(n10603), .B(n10606), .Z(n10604) );
  IV U11363 ( .A(n10576), .Z(n10601) );
  XOR U11364 ( .A(n10574), .B(n10607), .Z(n10576) );
  XOR U11365 ( .A(n10608), .B(n10609), .Z(n10607) );
  ANDN U11366 ( .B(n10610), .A(n10611), .Z(n10608) );
  XOR U11367 ( .A(n10612), .B(n10609), .Z(n10610) );
  IV U11368 ( .A(n10577), .Z(n10574) );
  XOR U11369 ( .A(n10613), .B(n10614), .Z(n10577) );
  ANDN U11370 ( .B(n10615), .A(n10616), .Z(n10613) );
  XOR U11371 ( .A(n10614), .B(n10617), .Z(n10615) );
  XOR U11372 ( .A(n10618), .B(n10619), .Z(n10590) );
  XNOR U11373 ( .A(n10585), .B(n10620), .Z(n10619) );
  IV U11374 ( .A(n10588), .Z(n10620) );
  XOR U11375 ( .A(n10621), .B(n10622), .Z(n10588) );
  ANDN U11376 ( .B(n10623), .A(n10624), .Z(n10621) );
  XOR U11377 ( .A(n10622), .B(n10625), .Z(n10623) );
  XNOR U11378 ( .A(n10626), .B(n10627), .Z(n10585) );
  ANDN U11379 ( .B(n10628), .A(n10629), .Z(n10626) );
  XOR U11380 ( .A(n10627), .B(n10630), .Z(n10628) );
  IV U11381 ( .A(n10584), .Z(n10618) );
  XOR U11382 ( .A(n10582), .B(n10631), .Z(n10584) );
  XOR U11383 ( .A(n10632), .B(n10633), .Z(n10631) );
  ANDN U11384 ( .B(n10634), .A(n10635), .Z(n10632) );
  XOR U11385 ( .A(n10636), .B(n10633), .Z(n10634) );
  IV U11386 ( .A(n10586), .Z(n10582) );
  XOR U11387 ( .A(n10637), .B(n10638), .Z(n10586) );
  ANDN U11388 ( .B(n10639), .A(n10640), .Z(n10637) );
  XOR U11389 ( .A(n10641), .B(n10638), .Z(n10639) );
  IV U11390 ( .A(n10596), .Z(n10600) );
  XOR U11391 ( .A(n10596), .B(n10551), .Z(n10598) );
  XOR U11392 ( .A(n10642), .B(n10643), .Z(n10551) );
  AND U11393 ( .A(n206), .B(n10644), .Z(n10642) );
  XOR U11394 ( .A(n10645), .B(n10643), .Z(n10644) );
  NANDN U11395 ( .A(n10553), .B(n10555), .Z(n10596) );
  XOR U11396 ( .A(n10646), .B(n10647), .Z(n10555) );
  AND U11397 ( .A(n206), .B(n10648), .Z(n10646) );
  XOR U11398 ( .A(n10647), .B(n10649), .Z(n10648) );
  XNOR U11399 ( .A(n10650), .B(n10651), .Z(n206) );
  AND U11400 ( .A(n10652), .B(n10653), .Z(n10650) );
  XOR U11401 ( .A(n10651), .B(n10566), .Z(n10653) );
  XNOR U11402 ( .A(n10654), .B(n10655), .Z(n10566) );
  ANDN U11403 ( .B(n10656), .A(n10657), .Z(n10654) );
  XOR U11404 ( .A(n10655), .B(n10658), .Z(n10656) );
  XNOR U11405 ( .A(n10651), .B(n10568), .Z(n10652) );
  XOR U11406 ( .A(n10659), .B(n10660), .Z(n10568) );
  AND U11407 ( .A(n210), .B(n10661), .Z(n10659) );
  XOR U11408 ( .A(n10662), .B(n10660), .Z(n10661) );
  XNOR U11409 ( .A(n10663), .B(n10664), .Z(n10651) );
  AND U11410 ( .A(n10665), .B(n10666), .Z(n10663) );
  XNOR U11411 ( .A(n10664), .B(n10593), .Z(n10666) );
  XOR U11412 ( .A(n10657), .B(n10658), .Z(n10593) );
  XNOR U11413 ( .A(n10667), .B(n10668), .Z(n10658) );
  ANDN U11414 ( .B(n10669), .A(n10670), .Z(n10667) );
  XOR U11415 ( .A(n10671), .B(n10672), .Z(n10669) );
  XOR U11416 ( .A(n10673), .B(n10674), .Z(n10657) );
  XNOR U11417 ( .A(n10675), .B(n10676), .Z(n10674) );
  ANDN U11418 ( .B(n10677), .A(n10678), .Z(n10675) );
  XNOR U11419 ( .A(n10679), .B(n10680), .Z(n10677) );
  IV U11420 ( .A(n10655), .Z(n10673) );
  XOR U11421 ( .A(n10681), .B(n10682), .Z(n10655) );
  ANDN U11422 ( .B(n10683), .A(n10684), .Z(n10681) );
  XOR U11423 ( .A(n10682), .B(n10685), .Z(n10683) );
  XOR U11424 ( .A(n10664), .B(n10595), .Z(n10665) );
  XOR U11425 ( .A(n10686), .B(n10687), .Z(n10595) );
  AND U11426 ( .A(n210), .B(n10688), .Z(n10686) );
  XOR U11427 ( .A(n10689), .B(n10687), .Z(n10688) );
  XNOR U11428 ( .A(n10690), .B(n10691), .Z(n10664) );
  NAND U11429 ( .A(n10692), .B(n10693), .Z(n10691) );
  XOR U11430 ( .A(n10694), .B(n10643), .Z(n10693) );
  XOR U11431 ( .A(n10684), .B(n10685), .Z(n10643) );
  XOR U11432 ( .A(n10695), .B(n10672), .Z(n10685) );
  XOR U11433 ( .A(n10696), .B(n10697), .Z(n10672) );
  ANDN U11434 ( .B(n10698), .A(n10699), .Z(n10696) );
  XOR U11435 ( .A(n10697), .B(n10700), .Z(n10698) );
  IV U11436 ( .A(n10670), .Z(n10695) );
  XOR U11437 ( .A(n10668), .B(n10701), .Z(n10670) );
  XOR U11438 ( .A(n10702), .B(n10703), .Z(n10701) );
  ANDN U11439 ( .B(n10704), .A(n10705), .Z(n10702) );
  XOR U11440 ( .A(n10706), .B(n10703), .Z(n10704) );
  IV U11441 ( .A(n10671), .Z(n10668) );
  XOR U11442 ( .A(n10707), .B(n10708), .Z(n10671) );
  ANDN U11443 ( .B(n10709), .A(n10710), .Z(n10707) );
  XOR U11444 ( .A(n10708), .B(n10711), .Z(n10709) );
  XOR U11445 ( .A(n10712), .B(n10713), .Z(n10684) );
  XNOR U11446 ( .A(n10679), .B(n10714), .Z(n10713) );
  IV U11447 ( .A(n10682), .Z(n10714) );
  XOR U11448 ( .A(n10715), .B(n10716), .Z(n10682) );
  ANDN U11449 ( .B(n10717), .A(n10718), .Z(n10715) );
  XOR U11450 ( .A(n10716), .B(n10719), .Z(n10717) );
  XNOR U11451 ( .A(n10720), .B(n10721), .Z(n10679) );
  ANDN U11452 ( .B(n10722), .A(n10723), .Z(n10720) );
  XOR U11453 ( .A(n10721), .B(n10724), .Z(n10722) );
  IV U11454 ( .A(n10678), .Z(n10712) );
  XOR U11455 ( .A(n10676), .B(n10725), .Z(n10678) );
  XOR U11456 ( .A(n10726), .B(n10727), .Z(n10725) );
  ANDN U11457 ( .B(n10728), .A(n10729), .Z(n10726) );
  XOR U11458 ( .A(n10730), .B(n10727), .Z(n10728) );
  IV U11459 ( .A(n10680), .Z(n10676) );
  XOR U11460 ( .A(n10731), .B(n10732), .Z(n10680) );
  ANDN U11461 ( .B(n10733), .A(n10734), .Z(n10731) );
  XOR U11462 ( .A(n10735), .B(n10732), .Z(n10733) );
  IV U11463 ( .A(n10690), .Z(n10694) );
  XOR U11464 ( .A(n10690), .B(n10645), .Z(n10692) );
  XOR U11465 ( .A(n10736), .B(n10737), .Z(n10645) );
  AND U11466 ( .A(n210), .B(n10738), .Z(n10736) );
  XOR U11467 ( .A(n10739), .B(n10737), .Z(n10738) );
  NANDN U11468 ( .A(n10647), .B(n10649), .Z(n10690) );
  XOR U11469 ( .A(n10740), .B(n10741), .Z(n10649) );
  AND U11470 ( .A(n210), .B(n10742), .Z(n10740) );
  XOR U11471 ( .A(n10741), .B(n10743), .Z(n10742) );
  XNOR U11472 ( .A(n10744), .B(n10745), .Z(n210) );
  AND U11473 ( .A(n10746), .B(n10747), .Z(n10744) );
  XOR U11474 ( .A(n10745), .B(n10660), .Z(n10747) );
  XNOR U11475 ( .A(n10748), .B(n10749), .Z(n10660) );
  ANDN U11476 ( .B(n10750), .A(n10751), .Z(n10748) );
  XOR U11477 ( .A(n10749), .B(n10752), .Z(n10750) );
  XNOR U11478 ( .A(n10745), .B(n10662), .Z(n10746) );
  XOR U11479 ( .A(n10753), .B(n10754), .Z(n10662) );
  AND U11480 ( .A(n214), .B(n10755), .Z(n10753) );
  XOR U11481 ( .A(n10756), .B(n10754), .Z(n10755) );
  XNOR U11482 ( .A(n10757), .B(n10758), .Z(n10745) );
  AND U11483 ( .A(n10759), .B(n10760), .Z(n10757) );
  XNOR U11484 ( .A(n10758), .B(n10687), .Z(n10760) );
  XOR U11485 ( .A(n10751), .B(n10752), .Z(n10687) );
  XNOR U11486 ( .A(n10761), .B(n10762), .Z(n10752) );
  ANDN U11487 ( .B(n10763), .A(n10764), .Z(n10761) );
  XOR U11488 ( .A(n10765), .B(n10766), .Z(n10763) );
  XOR U11489 ( .A(n10767), .B(n10768), .Z(n10751) );
  XNOR U11490 ( .A(n10769), .B(n10770), .Z(n10768) );
  ANDN U11491 ( .B(n10771), .A(n10772), .Z(n10769) );
  XNOR U11492 ( .A(n10773), .B(n10774), .Z(n10771) );
  IV U11493 ( .A(n10749), .Z(n10767) );
  XOR U11494 ( .A(n10775), .B(n10776), .Z(n10749) );
  ANDN U11495 ( .B(n10777), .A(n10778), .Z(n10775) );
  XOR U11496 ( .A(n10776), .B(n10779), .Z(n10777) );
  XOR U11497 ( .A(n10758), .B(n10689), .Z(n10759) );
  XOR U11498 ( .A(n10780), .B(n10781), .Z(n10689) );
  AND U11499 ( .A(n214), .B(n10782), .Z(n10780) );
  XOR U11500 ( .A(n10783), .B(n10781), .Z(n10782) );
  XNOR U11501 ( .A(n10784), .B(n10785), .Z(n10758) );
  NAND U11502 ( .A(n10786), .B(n10787), .Z(n10785) );
  XOR U11503 ( .A(n10788), .B(n10737), .Z(n10787) );
  XOR U11504 ( .A(n10778), .B(n10779), .Z(n10737) );
  XOR U11505 ( .A(n10789), .B(n10766), .Z(n10779) );
  XOR U11506 ( .A(n10790), .B(n10791), .Z(n10766) );
  ANDN U11507 ( .B(n10792), .A(n10793), .Z(n10790) );
  XOR U11508 ( .A(n10791), .B(n10794), .Z(n10792) );
  IV U11509 ( .A(n10764), .Z(n10789) );
  XOR U11510 ( .A(n10762), .B(n10795), .Z(n10764) );
  XOR U11511 ( .A(n10796), .B(n10797), .Z(n10795) );
  ANDN U11512 ( .B(n10798), .A(n10799), .Z(n10796) );
  XOR U11513 ( .A(n10800), .B(n10797), .Z(n10798) );
  IV U11514 ( .A(n10765), .Z(n10762) );
  XOR U11515 ( .A(n10801), .B(n10802), .Z(n10765) );
  ANDN U11516 ( .B(n10803), .A(n10804), .Z(n10801) );
  XOR U11517 ( .A(n10802), .B(n10805), .Z(n10803) );
  XOR U11518 ( .A(n10806), .B(n10807), .Z(n10778) );
  XNOR U11519 ( .A(n10773), .B(n10808), .Z(n10807) );
  IV U11520 ( .A(n10776), .Z(n10808) );
  XOR U11521 ( .A(n10809), .B(n10810), .Z(n10776) );
  ANDN U11522 ( .B(n10811), .A(n10812), .Z(n10809) );
  XOR U11523 ( .A(n10810), .B(n10813), .Z(n10811) );
  XNOR U11524 ( .A(n10814), .B(n10815), .Z(n10773) );
  ANDN U11525 ( .B(n10816), .A(n10817), .Z(n10814) );
  XOR U11526 ( .A(n10815), .B(n10818), .Z(n10816) );
  IV U11527 ( .A(n10772), .Z(n10806) );
  XOR U11528 ( .A(n10770), .B(n10819), .Z(n10772) );
  XOR U11529 ( .A(n10820), .B(n10821), .Z(n10819) );
  ANDN U11530 ( .B(n10822), .A(n10823), .Z(n10820) );
  XOR U11531 ( .A(n10824), .B(n10821), .Z(n10822) );
  IV U11532 ( .A(n10774), .Z(n10770) );
  XOR U11533 ( .A(n10825), .B(n10826), .Z(n10774) );
  ANDN U11534 ( .B(n10827), .A(n10828), .Z(n10825) );
  XOR U11535 ( .A(n10829), .B(n10826), .Z(n10827) );
  IV U11536 ( .A(n10784), .Z(n10788) );
  XOR U11537 ( .A(n10784), .B(n10739), .Z(n10786) );
  XOR U11538 ( .A(n10830), .B(n10831), .Z(n10739) );
  AND U11539 ( .A(n214), .B(n10832), .Z(n10830) );
  XOR U11540 ( .A(n10833), .B(n10831), .Z(n10832) );
  NANDN U11541 ( .A(n10741), .B(n10743), .Z(n10784) );
  XOR U11542 ( .A(n10834), .B(n10835), .Z(n10743) );
  AND U11543 ( .A(n214), .B(n10836), .Z(n10834) );
  XOR U11544 ( .A(n10835), .B(n10837), .Z(n10836) );
  XNOR U11545 ( .A(n10838), .B(n10839), .Z(n214) );
  AND U11546 ( .A(n10840), .B(n10841), .Z(n10838) );
  XOR U11547 ( .A(n10839), .B(n10754), .Z(n10841) );
  XNOR U11548 ( .A(n10842), .B(n10843), .Z(n10754) );
  ANDN U11549 ( .B(n10844), .A(n10845), .Z(n10842) );
  XOR U11550 ( .A(n10843), .B(n10846), .Z(n10844) );
  XNOR U11551 ( .A(n10839), .B(n10756), .Z(n10840) );
  XOR U11552 ( .A(n10847), .B(n10848), .Z(n10756) );
  AND U11553 ( .A(n218), .B(n10849), .Z(n10847) );
  XOR U11554 ( .A(n10850), .B(n10848), .Z(n10849) );
  XNOR U11555 ( .A(n10851), .B(n10852), .Z(n10839) );
  AND U11556 ( .A(n10853), .B(n10854), .Z(n10851) );
  XNOR U11557 ( .A(n10852), .B(n10781), .Z(n10854) );
  XOR U11558 ( .A(n10845), .B(n10846), .Z(n10781) );
  XNOR U11559 ( .A(n10855), .B(n10856), .Z(n10846) );
  ANDN U11560 ( .B(n10857), .A(n10858), .Z(n10855) );
  XOR U11561 ( .A(n10859), .B(n10860), .Z(n10857) );
  XOR U11562 ( .A(n10861), .B(n10862), .Z(n10845) );
  XNOR U11563 ( .A(n10863), .B(n10864), .Z(n10862) );
  ANDN U11564 ( .B(n10865), .A(n10866), .Z(n10863) );
  XNOR U11565 ( .A(n10867), .B(n10868), .Z(n10865) );
  IV U11566 ( .A(n10843), .Z(n10861) );
  XOR U11567 ( .A(n10869), .B(n10870), .Z(n10843) );
  ANDN U11568 ( .B(n10871), .A(n10872), .Z(n10869) );
  XOR U11569 ( .A(n10870), .B(n10873), .Z(n10871) );
  XOR U11570 ( .A(n10852), .B(n10783), .Z(n10853) );
  XOR U11571 ( .A(n10874), .B(n10875), .Z(n10783) );
  AND U11572 ( .A(n218), .B(n10876), .Z(n10874) );
  XOR U11573 ( .A(n10877), .B(n10875), .Z(n10876) );
  XNOR U11574 ( .A(n10878), .B(n10879), .Z(n10852) );
  NAND U11575 ( .A(n10880), .B(n10881), .Z(n10879) );
  XOR U11576 ( .A(n10882), .B(n10831), .Z(n10881) );
  XOR U11577 ( .A(n10872), .B(n10873), .Z(n10831) );
  XOR U11578 ( .A(n10883), .B(n10860), .Z(n10873) );
  XOR U11579 ( .A(n10884), .B(n10885), .Z(n10860) );
  ANDN U11580 ( .B(n10886), .A(n10887), .Z(n10884) );
  XOR U11581 ( .A(n10885), .B(n10888), .Z(n10886) );
  IV U11582 ( .A(n10858), .Z(n10883) );
  XOR U11583 ( .A(n10856), .B(n10889), .Z(n10858) );
  XOR U11584 ( .A(n10890), .B(n10891), .Z(n10889) );
  ANDN U11585 ( .B(n10892), .A(n10893), .Z(n10890) );
  XOR U11586 ( .A(n10894), .B(n10891), .Z(n10892) );
  IV U11587 ( .A(n10859), .Z(n10856) );
  XOR U11588 ( .A(n10895), .B(n10896), .Z(n10859) );
  ANDN U11589 ( .B(n10897), .A(n10898), .Z(n10895) );
  XOR U11590 ( .A(n10896), .B(n10899), .Z(n10897) );
  XOR U11591 ( .A(n10900), .B(n10901), .Z(n10872) );
  XNOR U11592 ( .A(n10867), .B(n10902), .Z(n10901) );
  IV U11593 ( .A(n10870), .Z(n10902) );
  XOR U11594 ( .A(n10903), .B(n10904), .Z(n10870) );
  ANDN U11595 ( .B(n10905), .A(n10906), .Z(n10903) );
  XOR U11596 ( .A(n10904), .B(n10907), .Z(n10905) );
  XNOR U11597 ( .A(n10908), .B(n10909), .Z(n10867) );
  ANDN U11598 ( .B(n10910), .A(n10911), .Z(n10908) );
  XOR U11599 ( .A(n10909), .B(n10912), .Z(n10910) );
  IV U11600 ( .A(n10866), .Z(n10900) );
  XOR U11601 ( .A(n10864), .B(n10913), .Z(n10866) );
  XOR U11602 ( .A(n10914), .B(n10915), .Z(n10913) );
  ANDN U11603 ( .B(n10916), .A(n10917), .Z(n10914) );
  XOR U11604 ( .A(n10918), .B(n10915), .Z(n10916) );
  IV U11605 ( .A(n10868), .Z(n10864) );
  XOR U11606 ( .A(n10919), .B(n10920), .Z(n10868) );
  ANDN U11607 ( .B(n10921), .A(n10922), .Z(n10919) );
  XOR U11608 ( .A(n10923), .B(n10920), .Z(n10921) );
  IV U11609 ( .A(n10878), .Z(n10882) );
  XOR U11610 ( .A(n10878), .B(n10833), .Z(n10880) );
  XOR U11611 ( .A(n10924), .B(n10925), .Z(n10833) );
  AND U11612 ( .A(n218), .B(n10926), .Z(n10924) );
  XOR U11613 ( .A(n10927), .B(n10925), .Z(n10926) );
  NANDN U11614 ( .A(n10835), .B(n10837), .Z(n10878) );
  XOR U11615 ( .A(n10928), .B(n10929), .Z(n10837) );
  AND U11616 ( .A(n218), .B(n10930), .Z(n10928) );
  XOR U11617 ( .A(n10929), .B(n10931), .Z(n10930) );
  XNOR U11618 ( .A(n10932), .B(n10933), .Z(n218) );
  AND U11619 ( .A(n10934), .B(n10935), .Z(n10932) );
  XOR U11620 ( .A(n10933), .B(n10848), .Z(n10935) );
  XNOR U11621 ( .A(n10936), .B(n10937), .Z(n10848) );
  ANDN U11622 ( .B(n10938), .A(n10939), .Z(n10936) );
  XOR U11623 ( .A(n10937), .B(n10940), .Z(n10938) );
  XNOR U11624 ( .A(n10933), .B(n10850), .Z(n10934) );
  XOR U11625 ( .A(n10941), .B(n10942), .Z(n10850) );
  AND U11626 ( .A(n222), .B(n10943), .Z(n10941) );
  XOR U11627 ( .A(n10944), .B(n10942), .Z(n10943) );
  XNOR U11628 ( .A(n10945), .B(n10946), .Z(n10933) );
  AND U11629 ( .A(n10947), .B(n10948), .Z(n10945) );
  XNOR U11630 ( .A(n10946), .B(n10875), .Z(n10948) );
  XOR U11631 ( .A(n10939), .B(n10940), .Z(n10875) );
  XNOR U11632 ( .A(n10949), .B(n10950), .Z(n10940) );
  ANDN U11633 ( .B(n10951), .A(n10952), .Z(n10949) );
  XOR U11634 ( .A(n10953), .B(n10954), .Z(n10951) );
  XOR U11635 ( .A(n10955), .B(n10956), .Z(n10939) );
  XNOR U11636 ( .A(n10957), .B(n10958), .Z(n10956) );
  ANDN U11637 ( .B(n10959), .A(n10960), .Z(n10957) );
  XNOR U11638 ( .A(n10961), .B(n10962), .Z(n10959) );
  IV U11639 ( .A(n10937), .Z(n10955) );
  XOR U11640 ( .A(n10963), .B(n10964), .Z(n10937) );
  ANDN U11641 ( .B(n10965), .A(n10966), .Z(n10963) );
  XOR U11642 ( .A(n10964), .B(n10967), .Z(n10965) );
  XOR U11643 ( .A(n10946), .B(n10877), .Z(n10947) );
  XOR U11644 ( .A(n10968), .B(n10969), .Z(n10877) );
  AND U11645 ( .A(n222), .B(n10970), .Z(n10968) );
  XOR U11646 ( .A(n10971), .B(n10969), .Z(n10970) );
  XNOR U11647 ( .A(n10972), .B(n10973), .Z(n10946) );
  NAND U11648 ( .A(n10974), .B(n10975), .Z(n10973) );
  XOR U11649 ( .A(n10976), .B(n10925), .Z(n10975) );
  XOR U11650 ( .A(n10966), .B(n10967), .Z(n10925) );
  XOR U11651 ( .A(n10977), .B(n10954), .Z(n10967) );
  XOR U11652 ( .A(n10978), .B(n10979), .Z(n10954) );
  ANDN U11653 ( .B(n10980), .A(n10981), .Z(n10978) );
  XOR U11654 ( .A(n10979), .B(n10982), .Z(n10980) );
  IV U11655 ( .A(n10952), .Z(n10977) );
  XOR U11656 ( .A(n10950), .B(n10983), .Z(n10952) );
  XOR U11657 ( .A(n10984), .B(n10985), .Z(n10983) );
  ANDN U11658 ( .B(n10986), .A(n10987), .Z(n10984) );
  XOR U11659 ( .A(n10988), .B(n10985), .Z(n10986) );
  IV U11660 ( .A(n10953), .Z(n10950) );
  XOR U11661 ( .A(n10989), .B(n10990), .Z(n10953) );
  ANDN U11662 ( .B(n10991), .A(n10992), .Z(n10989) );
  XOR U11663 ( .A(n10990), .B(n10993), .Z(n10991) );
  XOR U11664 ( .A(n10994), .B(n10995), .Z(n10966) );
  XNOR U11665 ( .A(n10961), .B(n10996), .Z(n10995) );
  IV U11666 ( .A(n10964), .Z(n10996) );
  XOR U11667 ( .A(n10997), .B(n10998), .Z(n10964) );
  ANDN U11668 ( .B(n10999), .A(n11000), .Z(n10997) );
  XOR U11669 ( .A(n10998), .B(n11001), .Z(n10999) );
  XNOR U11670 ( .A(n11002), .B(n11003), .Z(n10961) );
  ANDN U11671 ( .B(n11004), .A(n11005), .Z(n11002) );
  XOR U11672 ( .A(n11003), .B(n11006), .Z(n11004) );
  IV U11673 ( .A(n10960), .Z(n10994) );
  XOR U11674 ( .A(n10958), .B(n11007), .Z(n10960) );
  XOR U11675 ( .A(n11008), .B(n11009), .Z(n11007) );
  ANDN U11676 ( .B(n11010), .A(n11011), .Z(n11008) );
  XOR U11677 ( .A(n11012), .B(n11009), .Z(n11010) );
  IV U11678 ( .A(n10962), .Z(n10958) );
  XOR U11679 ( .A(n11013), .B(n11014), .Z(n10962) );
  ANDN U11680 ( .B(n11015), .A(n11016), .Z(n11013) );
  XOR U11681 ( .A(n11017), .B(n11014), .Z(n11015) );
  IV U11682 ( .A(n10972), .Z(n10976) );
  XOR U11683 ( .A(n10972), .B(n10927), .Z(n10974) );
  XOR U11684 ( .A(n11018), .B(n11019), .Z(n10927) );
  AND U11685 ( .A(n222), .B(n11020), .Z(n11018) );
  XOR U11686 ( .A(n11021), .B(n11019), .Z(n11020) );
  NANDN U11687 ( .A(n10929), .B(n10931), .Z(n10972) );
  XOR U11688 ( .A(n11022), .B(n11023), .Z(n10931) );
  AND U11689 ( .A(n222), .B(n11024), .Z(n11022) );
  XOR U11690 ( .A(n11023), .B(n11025), .Z(n11024) );
  XNOR U11691 ( .A(n11026), .B(n11027), .Z(n222) );
  AND U11692 ( .A(n11028), .B(n11029), .Z(n11026) );
  XOR U11693 ( .A(n11027), .B(n10942), .Z(n11029) );
  XNOR U11694 ( .A(n11030), .B(n11031), .Z(n10942) );
  ANDN U11695 ( .B(n11032), .A(n11033), .Z(n11030) );
  XOR U11696 ( .A(n11031), .B(n11034), .Z(n11032) );
  XNOR U11697 ( .A(n11027), .B(n10944), .Z(n11028) );
  XOR U11698 ( .A(n11035), .B(n11036), .Z(n10944) );
  AND U11699 ( .A(n226), .B(n11037), .Z(n11035) );
  XOR U11700 ( .A(n11038), .B(n11036), .Z(n11037) );
  XNOR U11701 ( .A(n11039), .B(n11040), .Z(n11027) );
  AND U11702 ( .A(n11041), .B(n11042), .Z(n11039) );
  XNOR U11703 ( .A(n11040), .B(n10969), .Z(n11042) );
  XOR U11704 ( .A(n11033), .B(n11034), .Z(n10969) );
  XNOR U11705 ( .A(n11043), .B(n11044), .Z(n11034) );
  ANDN U11706 ( .B(n11045), .A(n11046), .Z(n11043) );
  XOR U11707 ( .A(n11047), .B(n11048), .Z(n11045) );
  XOR U11708 ( .A(n11049), .B(n11050), .Z(n11033) );
  XNOR U11709 ( .A(n11051), .B(n11052), .Z(n11050) );
  ANDN U11710 ( .B(n11053), .A(n11054), .Z(n11051) );
  XNOR U11711 ( .A(n11055), .B(n11056), .Z(n11053) );
  IV U11712 ( .A(n11031), .Z(n11049) );
  XOR U11713 ( .A(n11057), .B(n11058), .Z(n11031) );
  ANDN U11714 ( .B(n11059), .A(n11060), .Z(n11057) );
  XOR U11715 ( .A(n11058), .B(n11061), .Z(n11059) );
  XOR U11716 ( .A(n11040), .B(n10971), .Z(n11041) );
  XOR U11717 ( .A(n11062), .B(n11063), .Z(n10971) );
  AND U11718 ( .A(n226), .B(n11064), .Z(n11062) );
  XOR U11719 ( .A(n11065), .B(n11063), .Z(n11064) );
  XNOR U11720 ( .A(n11066), .B(n11067), .Z(n11040) );
  NAND U11721 ( .A(n11068), .B(n11069), .Z(n11067) );
  XOR U11722 ( .A(n11070), .B(n11019), .Z(n11069) );
  XOR U11723 ( .A(n11060), .B(n11061), .Z(n11019) );
  XOR U11724 ( .A(n11071), .B(n11048), .Z(n11061) );
  XOR U11725 ( .A(n11072), .B(n11073), .Z(n11048) );
  ANDN U11726 ( .B(n11074), .A(n11075), .Z(n11072) );
  XOR U11727 ( .A(n11073), .B(n11076), .Z(n11074) );
  IV U11728 ( .A(n11046), .Z(n11071) );
  XOR U11729 ( .A(n11044), .B(n11077), .Z(n11046) );
  XOR U11730 ( .A(n11078), .B(n11079), .Z(n11077) );
  ANDN U11731 ( .B(n11080), .A(n11081), .Z(n11078) );
  XOR U11732 ( .A(n11082), .B(n11079), .Z(n11080) );
  IV U11733 ( .A(n11047), .Z(n11044) );
  XOR U11734 ( .A(n11083), .B(n11084), .Z(n11047) );
  ANDN U11735 ( .B(n11085), .A(n11086), .Z(n11083) );
  XOR U11736 ( .A(n11084), .B(n11087), .Z(n11085) );
  XOR U11737 ( .A(n11088), .B(n11089), .Z(n11060) );
  XNOR U11738 ( .A(n11055), .B(n11090), .Z(n11089) );
  IV U11739 ( .A(n11058), .Z(n11090) );
  XOR U11740 ( .A(n11091), .B(n11092), .Z(n11058) );
  ANDN U11741 ( .B(n11093), .A(n11094), .Z(n11091) );
  XOR U11742 ( .A(n11092), .B(n11095), .Z(n11093) );
  XNOR U11743 ( .A(n11096), .B(n11097), .Z(n11055) );
  ANDN U11744 ( .B(n11098), .A(n11099), .Z(n11096) );
  XOR U11745 ( .A(n11097), .B(n11100), .Z(n11098) );
  IV U11746 ( .A(n11054), .Z(n11088) );
  XOR U11747 ( .A(n11052), .B(n11101), .Z(n11054) );
  XOR U11748 ( .A(n11102), .B(n11103), .Z(n11101) );
  ANDN U11749 ( .B(n11104), .A(n11105), .Z(n11102) );
  XOR U11750 ( .A(n11106), .B(n11103), .Z(n11104) );
  IV U11751 ( .A(n11056), .Z(n11052) );
  XOR U11752 ( .A(n11107), .B(n11108), .Z(n11056) );
  ANDN U11753 ( .B(n11109), .A(n11110), .Z(n11107) );
  XOR U11754 ( .A(n11111), .B(n11108), .Z(n11109) );
  IV U11755 ( .A(n11066), .Z(n11070) );
  XOR U11756 ( .A(n11066), .B(n11021), .Z(n11068) );
  XOR U11757 ( .A(n11112), .B(n11113), .Z(n11021) );
  AND U11758 ( .A(n226), .B(n11114), .Z(n11112) );
  XOR U11759 ( .A(n11115), .B(n11113), .Z(n11114) );
  NANDN U11760 ( .A(n11023), .B(n11025), .Z(n11066) );
  XOR U11761 ( .A(n11116), .B(n11117), .Z(n11025) );
  AND U11762 ( .A(n226), .B(n11118), .Z(n11116) );
  XOR U11763 ( .A(n11117), .B(n11119), .Z(n11118) );
  XNOR U11764 ( .A(n11120), .B(n11121), .Z(n226) );
  AND U11765 ( .A(n11122), .B(n11123), .Z(n11120) );
  XOR U11766 ( .A(n11121), .B(n11036), .Z(n11123) );
  XNOR U11767 ( .A(n11124), .B(n11125), .Z(n11036) );
  ANDN U11768 ( .B(n11126), .A(n11127), .Z(n11124) );
  XOR U11769 ( .A(n11125), .B(n11128), .Z(n11126) );
  XNOR U11770 ( .A(n11121), .B(n11038), .Z(n11122) );
  XOR U11771 ( .A(n11129), .B(n11130), .Z(n11038) );
  AND U11772 ( .A(n230), .B(n11131), .Z(n11129) );
  XOR U11773 ( .A(n11132), .B(n11130), .Z(n11131) );
  XNOR U11774 ( .A(n11133), .B(n11134), .Z(n11121) );
  AND U11775 ( .A(n11135), .B(n11136), .Z(n11133) );
  XNOR U11776 ( .A(n11134), .B(n11063), .Z(n11136) );
  XOR U11777 ( .A(n11127), .B(n11128), .Z(n11063) );
  XNOR U11778 ( .A(n11137), .B(n11138), .Z(n11128) );
  ANDN U11779 ( .B(n11139), .A(n11140), .Z(n11137) );
  XOR U11780 ( .A(n11141), .B(n11142), .Z(n11139) );
  XOR U11781 ( .A(n11143), .B(n11144), .Z(n11127) );
  XNOR U11782 ( .A(n11145), .B(n11146), .Z(n11144) );
  ANDN U11783 ( .B(n11147), .A(n11148), .Z(n11145) );
  XNOR U11784 ( .A(n11149), .B(n11150), .Z(n11147) );
  IV U11785 ( .A(n11125), .Z(n11143) );
  XOR U11786 ( .A(n11151), .B(n11152), .Z(n11125) );
  ANDN U11787 ( .B(n11153), .A(n11154), .Z(n11151) );
  XOR U11788 ( .A(n11152), .B(n11155), .Z(n11153) );
  XOR U11789 ( .A(n11134), .B(n11065), .Z(n11135) );
  XOR U11790 ( .A(n11156), .B(n11157), .Z(n11065) );
  AND U11791 ( .A(n230), .B(n11158), .Z(n11156) );
  XOR U11792 ( .A(n11159), .B(n11157), .Z(n11158) );
  XNOR U11793 ( .A(n11160), .B(n11161), .Z(n11134) );
  NAND U11794 ( .A(n11162), .B(n11163), .Z(n11161) );
  XOR U11795 ( .A(n11164), .B(n11113), .Z(n11163) );
  XOR U11796 ( .A(n11154), .B(n11155), .Z(n11113) );
  XOR U11797 ( .A(n11165), .B(n11142), .Z(n11155) );
  XOR U11798 ( .A(n11166), .B(n11167), .Z(n11142) );
  ANDN U11799 ( .B(n11168), .A(n11169), .Z(n11166) );
  XOR U11800 ( .A(n11167), .B(n11170), .Z(n11168) );
  IV U11801 ( .A(n11140), .Z(n11165) );
  XOR U11802 ( .A(n11138), .B(n11171), .Z(n11140) );
  XOR U11803 ( .A(n11172), .B(n11173), .Z(n11171) );
  ANDN U11804 ( .B(n11174), .A(n11175), .Z(n11172) );
  XOR U11805 ( .A(n11176), .B(n11173), .Z(n11174) );
  IV U11806 ( .A(n11141), .Z(n11138) );
  XOR U11807 ( .A(n11177), .B(n11178), .Z(n11141) );
  ANDN U11808 ( .B(n11179), .A(n11180), .Z(n11177) );
  XOR U11809 ( .A(n11178), .B(n11181), .Z(n11179) );
  XOR U11810 ( .A(n11182), .B(n11183), .Z(n11154) );
  XNOR U11811 ( .A(n11149), .B(n11184), .Z(n11183) );
  IV U11812 ( .A(n11152), .Z(n11184) );
  XOR U11813 ( .A(n11185), .B(n11186), .Z(n11152) );
  ANDN U11814 ( .B(n11187), .A(n11188), .Z(n11185) );
  XOR U11815 ( .A(n11186), .B(n11189), .Z(n11187) );
  XNOR U11816 ( .A(n11190), .B(n11191), .Z(n11149) );
  ANDN U11817 ( .B(n11192), .A(n11193), .Z(n11190) );
  XOR U11818 ( .A(n11191), .B(n11194), .Z(n11192) );
  IV U11819 ( .A(n11148), .Z(n11182) );
  XOR U11820 ( .A(n11146), .B(n11195), .Z(n11148) );
  XOR U11821 ( .A(n11196), .B(n11197), .Z(n11195) );
  ANDN U11822 ( .B(n11198), .A(n11199), .Z(n11196) );
  XOR U11823 ( .A(n11200), .B(n11197), .Z(n11198) );
  IV U11824 ( .A(n11150), .Z(n11146) );
  XOR U11825 ( .A(n11201), .B(n11202), .Z(n11150) );
  ANDN U11826 ( .B(n11203), .A(n11204), .Z(n11201) );
  XOR U11827 ( .A(n11205), .B(n11202), .Z(n11203) );
  IV U11828 ( .A(n11160), .Z(n11164) );
  XOR U11829 ( .A(n11160), .B(n11115), .Z(n11162) );
  XOR U11830 ( .A(n11206), .B(n11207), .Z(n11115) );
  AND U11831 ( .A(n230), .B(n11208), .Z(n11206) );
  XOR U11832 ( .A(n11209), .B(n11207), .Z(n11208) );
  NANDN U11833 ( .A(n11117), .B(n11119), .Z(n11160) );
  XOR U11834 ( .A(n11210), .B(n11211), .Z(n11119) );
  AND U11835 ( .A(n230), .B(n11212), .Z(n11210) );
  XOR U11836 ( .A(n11211), .B(n11213), .Z(n11212) );
  XNOR U11837 ( .A(n11214), .B(n11215), .Z(n230) );
  AND U11838 ( .A(n11216), .B(n11217), .Z(n11214) );
  XOR U11839 ( .A(n11215), .B(n11130), .Z(n11217) );
  XNOR U11840 ( .A(n11218), .B(n11219), .Z(n11130) );
  ANDN U11841 ( .B(n11220), .A(n11221), .Z(n11218) );
  XOR U11842 ( .A(n11219), .B(n11222), .Z(n11220) );
  XNOR U11843 ( .A(n11215), .B(n11132), .Z(n11216) );
  XOR U11844 ( .A(n11223), .B(n11224), .Z(n11132) );
  AND U11845 ( .A(n234), .B(n11225), .Z(n11223) );
  XOR U11846 ( .A(n11226), .B(n11224), .Z(n11225) );
  XNOR U11847 ( .A(n11227), .B(n11228), .Z(n11215) );
  AND U11848 ( .A(n11229), .B(n11230), .Z(n11227) );
  XNOR U11849 ( .A(n11228), .B(n11157), .Z(n11230) );
  XOR U11850 ( .A(n11221), .B(n11222), .Z(n11157) );
  XNOR U11851 ( .A(n11231), .B(n11232), .Z(n11222) );
  ANDN U11852 ( .B(n11233), .A(n11234), .Z(n11231) );
  XOR U11853 ( .A(n11235), .B(n11236), .Z(n11233) );
  XOR U11854 ( .A(n11237), .B(n11238), .Z(n11221) );
  XNOR U11855 ( .A(n11239), .B(n11240), .Z(n11238) );
  ANDN U11856 ( .B(n11241), .A(n11242), .Z(n11239) );
  XNOR U11857 ( .A(n11243), .B(n11244), .Z(n11241) );
  IV U11858 ( .A(n11219), .Z(n11237) );
  XOR U11859 ( .A(n11245), .B(n11246), .Z(n11219) );
  ANDN U11860 ( .B(n11247), .A(n11248), .Z(n11245) );
  XOR U11861 ( .A(n11246), .B(n11249), .Z(n11247) );
  XOR U11862 ( .A(n11228), .B(n11159), .Z(n11229) );
  XOR U11863 ( .A(n11250), .B(n11251), .Z(n11159) );
  AND U11864 ( .A(n234), .B(n11252), .Z(n11250) );
  XOR U11865 ( .A(n11253), .B(n11251), .Z(n11252) );
  XNOR U11866 ( .A(n11254), .B(n11255), .Z(n11228) );
  NAND U11867 ( .A(n11256), .B(n11257), .Z(n11255) );
  XOR U11868 ( .A(n11258), .B(n11207), .Z(n11257) );
  XOR U11869 ( .A(n11248), .B(n11249), .Z(n11207) );
  XOR U11870 ( .A(n11259), .B(n11236), .Z(n11249) );
  XOR U11871 ( .A(n11260), .B(n11261), .Z(n11236) );
  ANDN U11872 ( .B(n11262), .A(n11263), .Z(n11260) );
  XOR U11873 ( .A(n11261), .B(n11264), .Z(n11262) );
  IV U11874 ( .A(n11234), .Z(n11259) );
  XOR U11875 ( .A(n11232), .B(n11265), .Z(n11234) );
  XOR U11876 ( .A(n11266), .B(n11267), .Z(n11265) );
  ANDN U11877 ( .B(n11268), .A(n11269), .Z(n11266) );
  XOR U11878 ( .A(n11270), .B(n11267), .Z(n11268) );
  IV U11879 ( .A(n11235), .Z(n11232) );
  XOR U11880 ( .A(n11271), .B(n11272), .Z(n11235) );
  ANDN U11881 ( .B(n11273), .A(n11274), .Z(n11271) );
  XOR U11882 ( .A(n11272), .B(n11275), .Z(n11273) );
  XOR U11883 ( .A(n11276), .B(n11277), .Z(n11248) );
  XNOR U11884 ( .A(n11243), .B(n11278), .Z(n11277) );
  IV U11885 ( .A(n11246), .Z(n11278) );
  XOR U11886 ( .A(n11279), .B(n11280), .Z(n11246) );
  ANDN U11887 ( .B(n11281), .A(n11282), .Z(n11279) );
  XOR U11888 ( .A(n11280), .B(n11283), .Z(n11281) );
  XNOR U11889 ( .A(n11284), .B(n11285), .Z(n11243) );
  ANDN U11890 ( .B(n11286), .A(n11287), .Z(n11284) );
  XOR U11891 ( .A(n11285), .B(n11288), .Z(n11286) );
  IV U11892 ( .A(n11242), .Z(n11276) );
  XOR U11893 ( .A(n11240), .B(n11289), .Z(n11242) );
  XOR U11894 ( .A(n11290), .B(n11291), .Z(n11289) );
  ANDN U11895 ( .B(n11292), .A(n11293), .Z(n11290) );
  XOR U11896 ( .A(n11294), .B(n11291), .Z(n11292) );
  IV U11897 ( .A(n11244), .Z(n11240) );
  XOR U11898 ( .A(n11295), .B(n11296), .Z(n11244) );
  ANDN U11899 ( .B(n11297), .A(n11298), .Z(n11295) );
  XOR U11900 ( .A(n11299), .B(n11296), .Z(n11297) );
  IV U11901 ( .A(n11254), .Z(n11258) );
  XOR U11902 ( .A(n11254), .B(n11209), .Z(n11256) );
  XOR U11903 ( .A(n11300), .B(n11301), .Z(n11209) );
  AND U11904 ( .A(n234), .B(n11302), .Z(n11300) );
  XOR U11905 ( .A(n11303), .B(n11301), .Z(n11302) );
  NANDN U11906 ( .A(n11211), .B(n11213), .Z(n11254) );
  XOR U11907 ( .A(n11304), .B(n11305), .Z(n11213) );
  AND U11908 ( .A(n234), .B(n11306), .Z(n11304) );
  XOR U11909 ( .A(n11305), .B(n11307), .Z(n11306) );
  XNOR U11910 ( .A(n11308), .B(n11309), .Z(n234) );
  AND U11911 ( .A(n11310), .B(n11311), .Z(n11308) );
  XOR U11912 ( .A(n11309), .B(n11224), .Z(n11311) );
  XNOR U11913 ( .A(n11312), .B(n11313), .Z(n11224) );
  ANDN U11914 ( .B(n11314), .A(n11315), .Z(n11312) );
  XOR U11915 ( .A(n11313), .B(n11316), .Z(n11314) );
  XNOR U11916 ( .A(n11309), .B(n11226), .Z(n11310) );
  XOR U11917 ( .A(n11317), .B(n11318), .Z(n11226) );
  AND U11918 ( .A(n238), .B(n11319), .Z(n11317) );
  XOR U11919 ( .A(n11320), .B(n11318), .Z(n11319) );
  XNOR U11920 ( .A(n11321), .B(n11322), .Z(n11309) );
  AND U11921 ( .A(n11323), .B(n11324), .Z(n11321) );
  XNOR U11922 ( .A(n11322), .B(n11251), .Z(n11324) );
  XOR U11923 ( .A(n11315), .B(n11316), .Z(n11251) );
  XNOR U11924 ( .A(n11325), .B(n11326), .Z(n11316) );
  ANDN U11925 ( .B(n11327), .A(n11328), .Z(n11325) );
  XOR U11926 ( .A(n11329), .B(n11330), .Z(n11327) );
  XOR U11927 ( .A(n11331), .B(n11332), .Z(n11315) );
  XNOR U11928 ( .A(n11333), .B(n11334), .Z(n11332) );
  ANDN U11929 ( .B(n11335), .A(n11336), .Z(n11333) );
  XNOR U11930 ( .A(n11337), .B(n11338), .Z(n11335) );
  IV U11931 ( .A(n11313), .Z(n11331) );
  XOR U11932 ( .A(n11339), .B(n11340), .Z(n11313) );
  ANDN U11933 ( .B(n11341), .A(n11342), .Z(n11339) );
  XOR U11934 ( .A(n11340), .B(n11343), .Z(n11341) );
  XOR U11935 ( .A(n11322), .B(n11253), .Z(n11323) );
  XOR U11936 ( .A(n11344), .B(n11345), .Z(n11253) );
  AND U11937 ( .A(n238), .B(n11346), .Z(n11344) );
  XOR U11938 ( .A(n11347), .B(n11345), .Z(n11346) );
  XNOR U11939 ( .A(n11348), .B(n11349), .Z(n11322) );
  NAND U11940 ( .A(n11350), .B(n11351), .Z(n11349) );
  XOR U11941 ( .A(n11352), .B(n11301), .Z(n11351) );
  XOR U11942 ( .A(n11342), .B(n11343), .Z(n11301) );
  XOR U11943 ( .A(n11353), .B(n11330), .Z(n11343) );
  XOR U11944 ( .A(n11354), .B(n11355), .Z(n11330) );
  ANDN U11945 ( .B(n11356), .A(n11357), .Z(n11354) );
  XOR U11946 ( .A(n11355), .B(n11358), .Z(n11356) );
  IV U11947 ( .A(n11328), .Z(n11353) );
  XOR U11948 ( .A(n11326), .B(n11359), .Z(n11328) );
  XOR U11949 ( .A(n11360), .B(n11361), .Z(n11359) );
  ANDN U11950 ( .B(n11362), .A(n11363), .Z(n11360) );
  XOR U11951 ( .A(n11364), .B(n11361), .Z(n11362) );
  IV U11952 ( .A(n11329), .Z(n11326) );
  XOR U11953 ( .A(n11365), .B(n11366), .Z(n11329) );
  ANDN U11954 ( .B(n11367), .A(n11368), .Z(n11365) );
  XOR U11955 ( .A(n11366), .B(n11369), .Z(n11367) );
  XOR U11956 ( .A(n11370), .B(n11371), .Z(n11342) );
  XNOR U11957 ( .A(n11337), .B(n11372), .Z(n11371) );
  IV U11958 ( .A(n11340), .Z(n11372) );
  XOR U11959 ( .A(n11373), .B(n11374), .Z(n11340) );
  ANDN U11960 ( .B(n11375), .A(n11376), .Z(n11373) );
  XOR U11961 ( .A(n11374), .B(n11377), .Z(n11375) );
  XNOR U11962 ( .A(n11378), .B(n11379), .Z(n11337) );
  ANDN U11963 ( .B(n11380), .A(n11381), .Z(n11378) );
  XOR U11964 ( .A(n11379), .B(n11382), .Z(n11380) );
  IV U11965 ( .A(n11336), .Z(n11370) );
  XOR U11966 ( .A(n11334), .B(n11383), .Z(n11336) );
  XOR U11967 ( .A(n11384), .B(n11385), .Z(n11383) );
  ANDN U11968 ( .B(n11386), .A(n11387), .Z(n11384) );
  XOR U11969 ( .A(n11388), .B(n11385), .Z(n11386) );
  IV U11970 ( .A(n11338), .Z(n11334) );
  XOR U11971 ( .A(n11389), .B(n11390), .Z(n11338) );
  ANDN U11972 ( .B(n11391), .A(n11392), .Z(n11389) );
  XOR U11973 ( .A(n11393), .B(n11390), .Z(n11391) );
  IV U11974 ( .A(n11348), .Z(n11352) );
  XOR U11975 ( .A(n11348), .B(n11303), .Z(n11350) );
  XOR U11976 ( .A(n11394), .B(n11395), .Z(n11303) );
  AND U11977 ( .A(n238), .B(n11396), .Z(n11394) );
  XOR U11978 ( .A(n11397), .B(n11395), .Z(n11396) );
  NANDN U11979 ( .A(n11305), .B(n11307), .Z(n11348) );
  XOR U11980 ( .A(n11398), .B(n11399), .Z(n11307) );
  AND U11981 ( .A(n238), .B(n11400), .Z(n11398) );
  XOR U11982 ( .A(n11399), .B(n11401), .Z(n11400) );
  XNOR U11983 ( .A(n11402), .B(n11403), .Z(n238) );
  AND U11984 ( .A(n11404), .B(n11405), .Z(n11402) );
  XOR U11985 ( .A(n11403), .B(n11318), .Z(n11405) );
  XNOR U11986 ( .A(n11406), .B(n11407), .Z(n11318) );
  ANDN U11987 ( .B(n11408), .A(n11409), .Z(n11406) );
  XOR U11988 ( .A(n11407), .B(n11410), .Z(n11408) );
  XNOR U11989 ( .A(n11403), .B(n11320), .Z(n11404) );
  XOR U11990 ( .A(n11411), .B(n11412), .Z(n11320) );
  AND U11991 ( .A(n242), .B(n11413), .Z(n11411) );
  XOR U11992 ( .A(n11414), .B(n11412), .Z(n11413) );
  XNOR U11993 ( .A(n11415), .B(n11416), .Z(n11403) );
  AND U11994 ( .A(n11417), .B(n11418), .Z(n11415) );
  XNOR U11995 ( .A(n11416), .B(n11345), .Z(n11418) );
  XOR U11996 ( .A(n11409), .B(n11410), .Z(n11345) );
  XNOR U11997 ( .A(n11419), .B(n11420), .Z(n11410) );
  ANDN U11998 ( .B(n11421), .A(n11422), .Z(n11419) );
  XOR U11999 ( .A(n11423), .B(n11424), .Z(n11421) );
  XOR U12000 ( .A(n11425), .B(n11426), .Z(n11409) );
  XNOR U12001 ( .A(n11427), .B(n11428), .Z(n11426) );
  ANDN U12002 ( .B(n11429), .A(n11430), .Z(n11427) );
  XNOR U12003 ( .A(n11431), .B(n11432), .Z(n11429) );
  IV U12004 ( .A(n11407), .Z(n11425) );
  XOR U12005 ( .A(n11433), .B(n11434), .Z(n11407) );
  ANDN U12006 ( .B(n11435), .A(n11436), .Z(n11433) );
  XOR U12007 ( .A(n11434), .B(n11437), .Z(n11435) );
  XOR U12008 ( .A(n11416), .B(n11347), .Z(n11417) );
  XOR U12009 ( .A(n11438), .B(n11439), .Z(n11347) );
  AND U12010 ( .A(n242), .B(n11440), .Z(n11438) );
  XOR U12011 ( .A(n11441), .B(n11439), .Z(n11440) );
  XNOR U12012 ( .A(n11442), .B(n11443), .Z(n11416) );
  NAND U12013 ( .A(n11444), .B(n11445), .Z(n11443) );
  XOR U12014 ( .A(n11446), .B(n11395), .Z(n11445) );
  XOR U12015 ( .A(n11436), .B(n11437), .Z(n11395) );
  XOR U12016 ( .A(n11447), .B(n11424), .Z(n11437) );
  XOR U12017 ( .A(n11448), .B(n11449), .Z(n11424) );
  ANDN U12018 ( .B(n11450), .A(n11451), .Z(n11448) );
  XOR U12019 ( .A(n11449), .B(n11452), .Z(n11450) );
  IV U12020 ( .A(n11422), .Z(n11447) );
  XOR U12021 ( .A(n11420), .B(n11453), .Z(n11422) );
  XOR U12022 ( .A(n11454), .B(n11455), .Z(n11453) );
  ANDN U12023 ( .B(n11456), .A(n11457), .Z(n11454) );
  XOR U12024 ( .A(n11458), .B(n11455), .Z(n11456) );
  IV U12025 ( .A(n11423), .Z(n11420) );
  XOR U12026 ( .A(n11459), .B(n11460), .Z(n11423) );
  ANDN U12027 ( .B(n11461), .A(n11462), .Z(n11459) );
  XOR U12028 ( .A(n11460), .B(n11463), .Z(n11461) );
  XOR U12029 ( .A(n11464), .B(n11465), .Z(n11436) );
  XNOR U12030 ( .A(n11431), .B(n11466), .Z(n11465) );
  IV U12031 ( .A(n11434), .Z(n11466) );
  XOR U12032 ( .A(n11467), .B(n11468), .Z(n11434) );
  ANDN U12033 ( .B(n11469), .A(n11470), .Z(n11467) );
  XOR U12034 ( .A(n11468), .B(n11471), .Z(n11469) );
  XNOR U12035 ( .A(n11472), .B(n11473), .Z(n11431) );
  ANDN U12036 ( .B(n11474), .A(n11475), .Z(n11472) );
  XOR U12037 ( .A(n11473), .B(n11476), .Z(n11474) );
  IV U12038 ( .A(n11430), .Z(n11464) );
  XOR U12039 ( .A(n11428), .B(n11477), .Z(n11430) );
  XOR U12040 ( .A(n11478), .B(n11479), .Z(n11477) );
  ANDN U12041 ( .B(n11480), .A(n11481), .Z(n11478) );
  XOR U12042 ( .A(n11482), .B(n11479), .Z(n11480) );
  IV U12043 ( .A(n11432), .Z(n11428) );
  XOR U12044 ( .A(n11483), .B(n11484), .Z(n11432) );
  ANDN U12045 ( .B(n11485), .A(n11486), .Z(n11483) );
  XOR U12046 ( .A(n11487), .B(n11484), .Z(n11485) );
  IV U12047 ( .A(n11442), .Z(n11446) );
  XOR U12048 ( .A(n11442), .B(n11397), .Z(n11444) );
  XOR U12049 ( .A(n11488), .B(n11489), .Z(n11397) );
  AND U12050 ( .A(n242), .B(n11490), .Z(n11488) );
  XOR U12051 ( .A(n11491), .B(n11489), .Z(n11490) );
  NANDN U12052 ( .A(n11399), .B(n11401), .Z(n11442) );
  XOR U12053 ( .A(n11492), .B(n11493), .Z(n11401) );
  AND U12054 ( .A(n242), .B(n11494), .Z(n11492) );
  XOR U12055 ( .A(n11493), .B(n11495), .Z(n11494) );
  XNOR U12056 ( .A(n11496), .B(n11497), .Z(n242) );
  AND U12057 ( .A(n11498), .B(n11499), .Z(n11496) );
  XOR U12058 ( .A(n11497), .B(n11412), .Z(n11499) );
  XNOR U12059 ( .A(n11500), .B(n11501), .Z(n11412) );
  ANDN U12060 ( .B(n11502), .A(n11503), .Z(n11500) );
  XOR U12061 ( .A(n11501), .B(n11504), .Z(n11502) );
  XNOR U12062 ( .A(n11497), .B(n11414), .Z(n11498) );
  XOR U12063 ( .A(n11505), .B(n11506), .Z(n11414) );
  AND U12064 ( .A(n246), .B(n11507), .Z(n11505) );
  XOR U12065 ( .A(n11508), .B(n11506), .Z(n11507) );
  XNOR U12066 ( .A(n11509), .B(n11510), .Z(n11497) );
  AND U12067 ( .A(n11511), .B(n11512), .Z(n11509) );
  XNOR U12068 ( .A(n11510), .B(n11439), .Z(n11512) );
  XOR U12069 ( .A(n11503), .B(n11504), .Z(n11439) );
  XNOR U12070 ( .A(n11513), .B(n11514), .Z(n11504) );
  ANDN U12071 ( .B(n11515), .A(n11516), .Z(n11513) );
  XOR U12072 ( .A(n11517), .B(n11518), .Z(n11515) );
  XOR U12073 ( .A(n11519), .B(n11520), .Z(n11503) );
  XNOR U12074 ( .A(n11521), .B(n11522), .Z(n11520) );
  ANDN U12075 ( .B(n11523), .A(n11524), .Z(n11521) );
  XNOR U12076 ( .A(n11525), .B(n11526), .Z(n11523) );
  IV U12077 ( .A(n11501), .Z(n11519) );
  XOR U12078 ( .A(n11527), .B(n11528), .Z(n11501) );
  ANDN U12079 ( .B(n11529), .A(n11530), .Z(n11527) );
  XOR U12080 ( .A(n11528), .B(n11531), .Z(n11529) );
  XOR U12081 ( .A(n11510), .B(n11441), .Z(n11511) );
  XOR U12082 ( .A(n11532), .B(n11533), .Z(n11441) );
  AND U12083 ( .A(n246), .B(n11534), .Z(n11532) );
  XOR U12084 ( .A(n11535), .B(n11533), .Z(n11534) );
  XNOR U12085 ( .A(n11536), .B(n11537), .Z(n11510) );
  NAND U12086 ( .A(n11538), .B(n11539), .Z(n11537) );
  XOR U12087 ( .A(n11540), .B(n11489), .Z(n11539) );
  XOR U12088 ( .A(n11530), .B(n11531), .Z(n11489) );
  XOR U12089 ( .A(n11541), .B(n11518), .Z(n11531) );
  XOR U12090 ( .A(n11542), .B(n11543), .Z(n11518) );
  ANDN U12091 ( .B(n11544), .A(n11545), .Z(n11542) );
  XOR U12092 ( .A(n11543), .B(n11546), .Z(n11544) );
  IV U12093 ( .A(n11516), .Z(n11541) );
  XOR U12094 ( .A(n11514), .B(n11547), .Z(n11516) );
  XOR U12095 ( .A(n11548), .B(n11549), .Z(n11547) );
  ANDN U12096 ( .B(n11550), .A(n11551), .Z(n11548) );
  XOR U12097 ( .A(n11552), .B(n11549), .Z(n11550) );
  IV U12098 ( .A(n11517), .Z(n11514) );
  XOR U12099 ( .A(n11553), .B(n11554), .Z(n11517) );
  ANDN U12100 ( .B(n11555), .A(n11556), .Z(n11553) );
  XOR U12101 ( .A(n11554), .B(n11557), .Z(n11555) );
  XOR U12102 ( .A(n11558), .B(n11559), .Z(n11530) );
  XNOR U12103 ( .A(n11525), .B(n11560), .Z(n11559) );
  IV U12104 ( .A(n11528), .Z(n11560) );
  XOR U12105 ( .A(n11561), .B(n11562), .Z(n11528) );
  ANDN U12106 ( .B(n11563), .A(n11564), .Z(n11561) );
  XOR U12107 ( .A(n11562), .B(n11565), .Z(n11563) );
  XNOR U12108 ( .A(n11566), .B(n11567), .Z(n11525) );
  ANDN U12109 ( .B(n11568), .A(n11569), .Z(n11566) );
  XOR U12110 ( .A(n11567), .B(n11570), .Z(n11568) );
  IV U12111 ( .A(n11524), .Z(n11558) );
  XOR U12112 ( .A(n11522), .B(n11571), .Z(n11524) );
  XOR U12113 ( .A(n11572), .B(n11573), .Z(n11571) );
  ANDN U12114 ( .B(n11574), .A(n11575), .Z(n11572) );
  XOR U12115 ( .A(n11576), .B(n11573), .Z(n11574) );
  IV U12116 ( .A(n11526), .Z(n11522) );
  XOR U12117 ( .A(n11577), .B(n11578), .Z(n11526) );
  ANDN U12118 ( .B(n11579), .A(n11580), .Z(n11577) );
  XOR U12119 ( .A(n11581), .B(n11578), .Z(n11579) );
  IV U12120 ( .A(n11536), .Z(n11540) );
  XOR U12121 ( .A(n11536), .B(n11491), .Z(n11538) );
  XOR U12122 ( .A(n11582), .B(n11583), .Z(n11491) );
  AND U12123 ( .A(n246), .B(n11584), .Z(n11582) );
  XOR U12124 ( .A(n11585), .B(n11583), .Z(n11584) );
  NANDN U12125 ( .A(n11493), .B(n11495), .Z(n11536) );
  XOR U12126 ( .A(n11586), .B(n11587), .Z(n11495) );
  AND U12127 ( .A(n246), .B(n11588), .Z(n11586) );
  XOR U12128 ( .A(n11587), .B(n11589), .Z(n11588) );
  XNOR U12129 ( .A(n11590), .B(n11591), .Z(n246) );
  AND U12130 ( .A(n11592), .B(n11593), .Z(n11590) );
  XOR U12131 ( .A(n11591), .B(n11506), .Z(n11593) );
  XNOR U12132 ( .A(n11594), .B(n11595), .Z(n11506) );
  ANDN U12133 ( .B(n11596), .A(n11597), .Z(n11594) );
  XOR U12134 ( .A(n11595), .B(n11598), .Z(n11596) );
  XNOR U12135 ( .A(n11591), .B(n11508), .Z(n11592) );
  XOR U12136 ( .A(n11599), .B(n11600), .Z(n11508) );
  AND U12137 ( .A(n250), .B(n11601), .Z(n11599) );
  XOR U12138 ( .A(n11602), .B(n11600), .Z(n11601) );
  XNOR U12139 ( .A(n11603), .B(n11604), .Z(n11591) );
  AND U12140 ( .A(n11605), .B(n11606), .Z(n11603) );
  XNOR U12141 ( .A(n11604), .B(n11533), .Z(n11606) );
  XOR U12142 ( .A(n11597), .B(n11598), .Z(n11533) );
  XNOR U12143 ( .A(n11607), .B(n11608), .Z(n11598) );
  ANDN U12144 ( .B(n11609), .A(n11610), .Z(n11607) );
  XOR U12145 ( .A(n11611), .B(n11612), .Z(n11609) );
  XOR U12146 ( .A(n11613), .B(n11614), .Z(n11597) );
  XNOR U12147 ( .A(n11615), .B(n11616), .Z(n11614) );
  ANDN U12148 ( .B(n11617), .A(n11618), .Z(n11615) );
  XNOR U12149 ( .A(n11619), .B(n11620), .Z(n11617) );
  IV U12150 ( .A(n11595), .Z(n11613) );
  XOR U12151 ( .A(n11621), .B(n11622), .Z(n11595) );
  ANDN U12152 ( .B(n11623), .A(n11624), .Z(n11621) );
  XOR U12153 ( .A(n11622), .B(n11625), .Z(n11623) );
  XOR U12154 ( .A(n11604), .B(n11535), .Z(n11605) );
  XOR U12155 ( .A(n11626), .B(n11627), .Z(n11535) );
  AND U12156 ( .A(n250), .B(n11628), .Z(n11626) );
  XOR U12157 ( .A(n11629), .B(n11627), .Z(n11628) );
  XNOR U12158 ( .A(n11630), .B(n11631), .Z(n11604) );
  NAND U12159 ( .A(n11632), .B(n11633), .Z(n11631) );
  XOR U12160 ( .A(n11634), .B(n11583), .Z(n11633) );
  XOR U12161 ( .A(n11624), .B(n11625), .Z(n11583) );
  XOR U12162 ( .A(n11635), .B(n11612), .Z(n11625) );
  XOR U12163 ( .A(n11636), .B(n11637), .Z(n11612) );
  ANDN U12164 ( .B(n11638), .A(n11639), .Z(n11636) );
  XOR U12165 ( .A(n11637), .B(n11640), .Z(n11638) );
  IV U12166 ( .A(n11610), .Z(n11635) );
  XOR U12167 ( .A(n11608), .B(n11641), .Z(n11610) );
  XOR U12168 ( .A(n11642), .B(n11643), .Z(n11641) );
  ANDN U12169 ( .B(n11644), .A(n11645), .Z(n11642) );
  XOR U12170 ( .A(n11646), .B(n11643), .Z(n11644) );
  IV U12171 ( .A(n11611), .Z(n11608) );
  XOR U12172 ( .A(n11647), .B(n11648), .Z(n11611) );
  ANDN U12173 ( .B(n11649), .A(n11650), .Z(n11647) );
  XOR U12174 ( .A(n11648), .B(n11651), .Z(n11649) );
  XOR U12175 ( .A(n11652), .B(n11653), .Z(n11624) );
  XNOR U12176 ( .A(n11619), .B(n11654), .Z(n11653) );
  IV U12177 ( .A(n11622), .Z(n11654) );
  XOR U12178 ( .A(n11655), .B(n11656), .Z(n11622) );
  ANDN U12179 ( .B(n11657), .A(n11658), .Z(n11655) );
  XOR U12180 ( .A(n11656), .B(n11659), .Z(n11657) );
  XNOR U12181 ( .A(n11660), .B(n11661), .Z(n11619) );
  ANDN U12182 ( .B(n11662), .A(n11663), .Z(n11660) );
  XOR U12183 ( .A(n11661), .B(n11664), .Z(n11662) );
  IV U12184 ( .A(n11618), .Z(n11652) );
  XOR U12185 ( .A(n11616), .B(n11665), .Z(n11618) );
  XOR U12186 ( .A(n11666), .B(n11667), .Z(n11665) );
  ANDN U12187 ( .B(n11668), .A(n11669), .Z(n11666) );
  XOR U12188 ( .A(n11670), .B(n11667), .Z(n11668) );
  IV U12189 ( .A(n11620), .Z(n11616) );
  XOR U12190 ( .A(n11671), .B(n11672), .Z(n11620) );
  ANDN U12191 ( .B(n11673), .A(n11674), .Z(n11671) );
  XOR U12192 ( .A(n11675), .B(n11672), .Z(n11673) );
  IV U12193 ( .A(n11630), .Z(n11634) );
  XOR U12194 ( .A(n11630), .B(n11585), .Z(n11632) );
  XOR U12195 ( .A(n11676), .B(n11677), .Z(n11585) );
  AND U12196 ( .A(n250), .B(n11678), .Z(n11676) );
  XOR U12197 ( .A(n11679), .B(n11677), .Z(n11678) );
  NANDN U12198 ( .A(n11587), .B(n11589), .Z(n11630) );
  XOR U12199 ( .A(n11680), .B(n11681), .Z(n11589) );
  AND U12200 ( .A(n250), .B(n11682), .Z(n11680) );
  XOR U12201 ( .A(n11681), .B(n11683), .Z(n11682) );
  XNOR U12202 ( .A(n11684), .B(n11685), .Z(n250) );
  AND U12203 ( .A(n11686), .B(n11687), .Z(n11684) );
  XOR U12204 ( .A(n11685), .B(n11600), .Z(n11687) );
  XNOR U12205 ( .A(n11688), .B(n11689), .Z(n11600) );
  ANDN U12206 ( .B(n11690), .A(n11691), .Z(n11688) );
  XOR U12207 ( .A(n11689), .B(n11692), .Z(n11690) );
  XNOR U12208 ( .A(n11685), .B(n11602), .Z(n11686) );
  XOR U12209 ( .A(n11693), .B(n11694), .Z(n11602) );
  AND U12210 ( .A(n254), .B(n11695), .Z(n11693) );
  XOR U12211 ( .A(n11696), .B(n11694), .Z(n11695) );
  XNOR U12212 ( .A(n11697), .B(n11698), .Z(n11685) );
  AND U12213 ( .A(n11699), .B(n11700), .Z(n11697) );
  XNOR U12214 ( .A(n11698), .B(n11627), .Z(n11700) );
  XOR U12215 ( .A(n11691), .B(n11692), .Z(n11627) );
  XNOR U12216 ( .A(n11701), .B(n11702), .Z(n11692) );
  ANDN U12217 ( .B(n11703), .A(n11704), .Z(n11701) );
  XOR U12218 ( .A(n11705), .B(n11706), .Z(n11703) );
  XOR U12219 ( .A(n11707), .B(n11708), .Z(n11691) );
  XNOR U12220 ( .A(n11709), .B(n11710), .Z(n11708) );
  ANDN U12221 ( .B(n11711), .A(n11712), .Z(n11709) );
  XNOR U12222 ( .A(n11713), .B(n11714), .Z(n11711) );
  IV U12223 ( .A(n11689), .Z(n11707) );
  XOR U12224 ( .A(n11715), .B(n11716), .Z(n11689) );
  ANDN U12225 ( .B(n11717), .A(n11718), .Z(n11715) );
  XOR U12226 ( .A(n11716), .B(n11719), .Z(n11717) );
  XOR U12227 ( .A(n11698), .B(n11629), .Z(n11699) );
  XOR U12228 ( .A(n11720), .B(n11721), .Z(n11629) );
  AND U12229 ( .A(n254), .B(n11722), .Z(n11720) );
  XOR U12230 ( .A(n11723), .B(n11721), .Z(n11722) );
  XNOR U12231 ( .A(n11724), .B(n11725), .Z(n11698) );
  NAND U12232 ( .A(n11726), .B(n11727), .Z(n11725) );
  XOR U12233 ( .A(n11728), .B(n11677), .Z(n11727) );
  XOR U12234 ( .A(n11718), .B(n11719), .Z(n11677) );
  XOR U12235 ( .A(n11729), .B(n11706), .Z(n11719) );
  XOR U12236 ( .A(n11730), .B(n11731), .Z(n11706) );
  ANDN U12237 ( .B(n11732), .A(n11733), .Z(n11730) );
  XOR U12238 ( .A(n11731), .B(n11734), .Z(n11732) );
  IV U12239 ( .A(n11704), .Z(n11729) );
  XOR U12240 ( .A(n11702), .B(n11735), .Z(n11704) );
  XOR U12241 ( .A(n11736), .B(n11737), .Z(n11735) );
  ANDN U12242 ( .B(n11738), .A(n11739), .Z(n11736) );
  XOR U12243 ( .A(n11740), .B(n11737), .Z(n11738) );
  IV U12244 ( .A(n11705), .Z(n11702) );
  XOR U12245 ( .A(n11741), .B(n11742), .Z(n11705) );
  ANDN U12246 ( .B(n11743), .A(n11744), .Z(n11741) );
  XOR U12247 ( .A(n11742), .B(n11745), .Z(n11743) );
  XOR U12248 ( .A(n11746), .B(n11747), .Z(n11718) );
  XNOR U12249 ( .A(n11713), .B(n11748), .Z(n11747) );
  IV U12250 ( .A(n11716), .Z(n11748) );
  XOR U12251 ( .A(n11749), .B(n11750), .Z(n11716) );
  ANDN U12252 ( .B(n11751), .A(n11752), .Z(n11749) );
  XOR U12253 ( .A(n11750), .B(n11753), .Z(n11751) );
  XNOR U12254 ( .A(n11754), .B(n11755), .Z(n11713) );
  ANDN U12255 ( .B(n11756), .A(n11757), .Z(n11754) );
  XOR U12256 ( .A(n11755), .B(n11758), .Z(n11756) );
  IV U12257 ( .A(n11712), .Z(n11746) );
  XOR U12258 ( .A(n11710), .B(n11759), .Z(n11712) );
  XOR U12259 ( .A(n11760), .B(n11761), .Z(n11759) );
  ANDN U12260 ( .B(n11762), .A(n11763), .Z(n11760) );
  XOR U12261 ( .A(n11764), .B(n11761), .Z(n11762) );
  IV U12262 ( .A(n11714), .Z(n11710) );
  XOR U12263 ( .A(n11765), .B(n11766), .Z(n11714) );
  ANDN U12264 ( .B(n11767), .A(n11768), .Z(n11765) );
  XOR U12265 ( .A(n11769), .B(n11766), .Z(n11767) );
  IV U12266 ( .A(n11724), .Z(n11728) );
  XOR U12267 ( .A(n11724), .B(n11679), .Z(n11726) );
  XOR U12268 ( .A(n11770), .B(n11771), .Z(n11679) );
  AND U12269 ( .A(n254), .B(n11772), .Z(n11770) );
  XOR U12270 ( .A(n11773), .B(n11771), .Z(n11772) );
  NANDN U12271 ( .A(n11681), .B(n11683), .Z(n11724) );
  XOR U12272 ( .A(n11774), .B(n11775), .Z(n11683) );
  AND U12273 ( .A(n254), .B(n11776), .Z(n11774) );
  XOR U12274 ( .A(n11775), .B(n11777), .Z(n11776) );
  XNOR U12275 ( .A(n11778), .B(n11779), .Z(n254) );
  AND U12276 ( .A(n11780), .B(n11781), .Z(n11778) );
  XOR U12277 ( .A(n11779), .B(n11694), .Z(n11781) );
  XNOR U12278 ( .A(n11782), .B(n11783), .Z(n11694) );
  ANDN U12279 ( .B(n11784), .A(n11785), .Z(n11782) );
  XOR U12280 ( .A(n11783), .B(n11786), .Z(n11784) );
  XNOR U12281 ( .A(n11779), .B(n11696), .Z(n11780) );
  XOR U12282 ( .A(n11787), .B(n11788), .Z(n11696) );
  AND U12283 ( .A(n258), .B(n11789), .Z(n11787) );
  XOR U12284 ( .A(n11790), .B(n11788), .Z(n11789) );
  XNOR U12285 ( .A(n11791), .B(n11792), .Z(n11779) );
  AND U12286 ( .A(n11793), .B(n11794), .Z(n11791) );
  XNOR U12287 ( .A(n11792), .B(n11721), .Z(n11794) );
  XOR U12288 ( .A(n11785), .B(n11786), .Z(n11721) );
  XNOR U12289 ( .A(n11795), .B(n11796), .Z(n11786) );
  ANDN U12290 ( .B(n11797), .A(n11798), .Z(n11795) );
  XOR U12291 ( .A(n11799), .B(n11800), .Z(n11797) );
  XOR U12292 ( .A(n11801), .B(n11802), .Z(n11785) );
  XNOR U12293 ( .A(n11803), .B(n11804), .Z(n11802) );
  ANDN U12294 ( .B(n11805), .A(n11806), .Z(n11803) );
  XNOR U12295 ( .A(n11807), .B(n11808), .Z(n11805) );
  IV U12296 ( .A(n11783), .Z(n11801) );
  XOR U12297 ( .A(n11809), .B(n11810), .Z(n11783) );
  ANDN U12298 ( .B(n11811), .A(n11812), .Z(n11809) );
  XOR U12299 ( .A(n11810), .B(n11813), .Z(n11811) );
  XOR U12300 ( .A(n11792), .B(n11723), .Z(n11793) );
  XOR U12301 ( .A(n11814), .B(n11815), .Z(n11723) );
  AND U12302 ( .A(n258), .B(n11816), .Z(n11814) );
  XOR U12303 ( .A(n11817), .B(n11815), .Z(n11816) );
  XNOR U12304 ( .A(n11818), .B(n11819), .Z(n11792) );
  NAND U12305 ( .A(n11820), .B(n11821), .Z(n11819) );
  XOR U12306 ( .A(n11822), .B(n11771), .Z(n11821) );
  XOR U12307 ( .A(n11812), .B(n11813), .Z(n11771) );
  XOR U12308 ( .A(n11823), .B(n11800), .Z(n11813) );
  XOR U12309 ( .A(n11824), .B(n11825), .Z(n11800) );
  ANDN U12310 ( .B(n11826), .A(n11827), .Z(n11824) );
  XOR U12311 ( .A(n11825), .B(n11828), .Z(n11826) );
  IV U12312 ( .A(n11798), .Z(n11823) );
  XOR U12313 ( .A(n11796), .B(n11829), .Z(n11798) );
  XOR U12314 ( .A(n11830), .B(n11831), .Z(n11829) );
  ANDN U12315 ( .B(n11832), .A(n11833), .Z(n11830) );
  XOR U12316 ( .A(n11834), .B(n11831), .Z(n11832) );
  IV U12317 ( .A(n11799), .Z(n11796) );
  XOR U12318 ( .A(n11835), .B(n11836), .Z(n11799) );
  ANDN U12319 ( .B(n11837), .A(n11838), .Z(n11835) );
  XOR U12320 ( .A(n11836), .B(n11839), .Z(n11837) );
  XOR U12321 ( .A(n11840), .B(n11841), .Z(n11812) );
  XNOR U12322 ( .A(n11807), .B(n11842), .Z(n11841) );
  IV U12323 ( .A(n11810), .Z(n11842) );
  XOR U12324 ( .A(n11843), .B(n11844), .Z(n11810) );
  ANDN U12325 ( .B(n11845), .A(n11846), .Z(n11843) );
  XOR U12326 ( .A(n11844), .B(n11847), .Z(n11845) );
  XNOR U12327 ( .A(n11848), .B(n11849), .Z(n11807) );
  ANDN U12328 ( .B(n11850), .A(n11851), .Z(n11848) );
  XOR U12329 ( .A(n11849), .B(n11852), .Z(n11850) );
  IV U12330 ( .A(n11806), .Z(n11840) );
  XOR U12331 ( .A(n11804), .B(n11853), .Z(n11806) );
  XOR U12332 ( .A(n11854), .B(n11855), .Z(n11853) );
  ANDN U12333 ( .B(n11856), .A(n11857), .Z(n11854) );
  XOR U12334 ( .A(n11858), .B(n11855), .Z(n11856) );
  IV U12335 ( .A(n11808), .Z(n11804) );
  XOR U12336 ( .A(n11859), .B(n11860), .Z(n11808) );
  ANDN U12337 ( .B(n11861), .A(n11862), .Z(n11859) );
  XOR U12338 ( .A(n11863), .B(n11860), .Z(n11861) );
  IV U12339 ( .A(n11818), .Z(n11822) );
  XOR U12340 ( .A(n11818), .B(n11773), .Z(n11820) );
  XOR U12341 ( .A(n11864), .B(n11865), .Z(n11773) );
  AND U12342 ( .A(n258), .B(n11866), .Z(n11864) );
  XOR U12343 ( .A(n11867), .B(n11865), .Z(n11866) );
  NANDN U12344 ( .A(n11775), .B(n11777), .Z(n11818) );
  XOR U12345 ( .A(n11868), .B(n11869), .Z(n11777) );
  AND U12346 ( .A(n258), .B(n11870), .Z(n11868) );
  XOR U12347 ( .A(n11869), .B(n11871), .Z(n11870) );
  XNOR U12348 ( .A(n11872), .B(n11873), .Z(n258) );
  AND U12349 ( .A(n11874), .B(n11875), .Z(n11872) );
  XOR U12350 ( .A(n11873), .B(n11788), .Z(n11875) );
  XNOR U12351 ( .A(n11876), .B(n11877), .Z(n11788) );
  ANDN U12352 ( .B(n11878), .A(n11879), .Z(n11876) );
  XOR U12353 ( .A(n11877), .B(n11880), .Z(n11878) );
  XNOR U12354 ( .A(n11873), .B(n11790), .Z(n11874) );
  XOR U12355 ( .A(n11881), .B(n11882), .Z(n11790) );
  AND U12356 ( .A(n262), .B(n11883), .Z(n11881) );
  XOR U12357 ( .A(n11884), .B(n11882), .Z(n11883) );
  XNOR U12358 ( .A(n11885), .B(n11886), .Z(n11873) );
  AND U12359 ( .A(n11887), .B(n11888), .Z(n11885) );
  XNOR U12360 ( .A(n11886), .B(n11815), .Z(n11888) );
  XOR U12361 ( .A(n11879), .B(n11880), .Z(n11815) );
  XNOR U12362 ( .A(n11889), .B(n11890), .Z(n11880) );
  ANDN U12363 ( .B(n11891), .A(n11892), .Z(n11889) );
  XOR U12364 ( .A(n11893), .B(n11894), .Z(n11891) );
  XOR U12365 ( .A(n11895), .B(n11896), .Z(n11879) );
  XNOR U12366 ( .A(n11897), .B(n11898), .Z(n11896) );
  ANDN U12367 ( .B(n11899), .A(n11900), .Z(n11897) );
  XNOR U12368 ( .A(n11901), .B(n11902), .Z(n11899) );
  IV U12369 ( .A(n11877), .Z(n11895) );
  XOR U12370 ( .A(n11903), .B(n11904), .Z(n11877) );
  ANDN U12371 ( .B(n11905), .A(n11906), .Z(n11903) );
  XOR U12372 ( .A(n11904), .B(n11907), .Z(n11905) );
  XOR U12373 ( .A(n11886), .B(n11817), .Z(n11887) );
  XOR U12374 ( .A(n11908), .B(n11909), .Z(n11817) );
  AND U12375 ( .A(n262), .B(n11910), .Z(n11908) );
  XOR U12376 ( .A(n11911), .B(n11909), .Z(n11910) );
  XNOR U12377 ( .A(n11912), .B(n11913), .Z(n11886) );
  NAND U12378 ( .A(n11914), .B(n11915), .Z(n11913) );
  XOR U12379 ( .A(n11916), .B(n11865), .Z(n11915) );
  XOR U12380 ( .A(n11906), .B(n11907), .Z(n11865) );
  XOR U12381 ( .A(n11917), .B(n11894), .Z(n11907) );
  XOR U12382 ( .A(n11918), .B(n11919), .Z(n11894) );
  ANDN U12383 ( .B(n11920), .A(n11921), .Z(n11918) );
  XOR U12384 ( .A(n11919), .B(n11922), .Z(n11920) );
  IV U12385 ( .A(n11892), .Z(n11917) );
  XOR U12386 ( .A(n11890), .B(n11923), .Z(n11892) );
  XOR U12387 ( .A(n11924), .B(n11925), .Z(n11923) );
  ANDN U12388 ( .B(n11926), .A(n11927), .Z(n11924) );
  XOR U12389 ( .A(n11928), .B(n11925), .Z(n11926) );
  IV U12390 ( .A(n11893), .Z(n11890) );
  XOR U12391 ( .A(n11929), .B(n11930), .Z(n11893) );
  ANDN U12392 ( .B(n11931), .A(n11932), .Z(n11929) );
  XOR U12393 ( .A(n11930), .B(n11933), .Z(n11931) );
  XOR U12394 ( .A(n11934), .B(n11935), .Z(n11906) );
  XNOR U12395 ( .A(n11901), .B(n11936), .Z(n11935) );
  IV U12396 ( .A(n11904), .Z(n11936) );
  XOR U12397 ( .A(n11937), .B(n11938), .Z(n11904) );
  ANDN U12398 ( .B(n11939), .A(n11940), .Z(n11937) );
  XOR U12399 ( .A(n11938), .B(n11941), .Z(n11939) );
  XNOR U12400 ( .A(n11942), .B(n11943), .Z(n11901) );
  ANDN U12401 ( .B(n11944), .A(n11945), .Z(n11942) );
  XOR U12402 ( .A(n11943), .B(n11946), .Z(n11944) );
  IV U12403 ( .A(n11900), .Z(n11934) );
  XOR U12404 ( .A(n11898), .B(n11947), .Z(n11900) );
  XOR U12405 ( .A(n11948), .B(n11949), .Z(n11947) );
  ANDN U12406 ( .B(n11950), .A(n11951), .Z(n11948) );
  XOR U12407 ( .A(n11952), .B(n11949), .Z(n11950) );
  IV U12408 ( .A(n11902), .Z(n11898) );
  XOR U12409 ( .A(n11953), .B(n11954), .Z(n11902) );
  ANDN U12410 ( .B(n11955), .A(n11956), .Z(n11953) );
  XOR U12411 ( .A(n11957), .B(n11954), .Z(n11955) );
  IV U12412 ( .A(n11912), .Z(n11916) );
  XOR U12413 ( .A(n11912), .B(n11867), .Z(n11914) );
  XOR U12414 ( .A(n11958), .B(n11959), .Z(n11867) );
  AND U12415 ( .A(n262), .B(n11960), .Z(n11958) );
  XOR U12416 ( .A(n11961), .B(n11959), .Z(n11960) );
  NANDN U12417 ( .A(n11869), .B(n11871), .Z(n11912) );
  XOR U12418 ( .A(n11962), .B(n11963), .Z(n11871) );
  AND U12419 ( .A(n262), .B(n11964), .Z(n11962) );
  XOR U12420 ( .A(n11963), .B(n11965), .Z(n11964) );
  XNOR U12421 ( .A(n11966), .B(n11967), .Z(n262) );
  AND U12422 ( .A(n11968), .B(n11969), .Z(n11966) );
  XOR U12423 ( .A(n11967), .B(n11882), .Z(n11969) );
  XNOR U12424 ( .A(n11970), .B(n11971), .Z(n11882) );
  ANDN U12425 ( .B(n11972), .A(n11973), .Z(n11970) );
  XOR U12426 ( .A(n11971), .B(n11974), .Z(n11972) );
  XNOR U12427 ( .A(n11967), .B(n11884), .Z(n11968) );
  XOR U12428 ( .A(n11975), .B(n11976), .Z(n11884) );
  AND U12429 ( .A(n266), .B(n11977), .Z(n11975) );
  XOR U12430 ( .A(n11978), .B(n11976), .Z(n11977) );
  XNOR U12431 ( .A(n11979), .B(n11980), .Z(n11967) );
  AND U12432 ( .A(n11981), .B(n11982), .Z(n11979) );
  XNOR U12433 ( .A(n11980), .B(n11909), .Z(n11982) );
  XOR U12434 ( .A(n11973), .B(n11974), .Z(n11909) );
  XNOR U12435 ( .A(n11983), .B(n11984), .Z(n11974) );
  ANDN U12436 ( .B(n11985), .A(n11986), .Z(n11983) );
  XOR U12437 ( .A(n11987), .B(n11988), .Z(n11985) );
  XOR U12438 ( .A(n11989), .B(n11990), .Z(n11973) );
  XNOR U12439 ( .A(n11991), .B(n11992), .Z(n11990) );
  ANDN U12440 ( .B(n11993), .A(n11994), .Z(n11991) );
  XNOR U12441 ( .A(n11995), .B(n11996), .Z(n11993) );
  IV U12442 ( .A(n11971), .Z(n11989) );
  XOR U12443 ( .A(n11997), .B(n11998), .Z(n11971) );
  ANDN U12444 ( .B(n11999), .A(n12000), .Z(n11997) );
  XOR U12445 ( .A(n11998), .B(n12001), .Z(n11999) );
  XOR U12446 ( .A(n11980), .B(n11911), .Z(n11981) );
  XOR U12447 ( .A(n12002), .B(n12003), .Z(n11911) );
  AND U12448 ( .A(n266), .B(n12004), .Z(n12002) );
  XOR U12449 ( .A(n12005), .B(n12003), .Z(n12004) );
  XNOR U12450 ( .A(n12006), .B(n12007), .Z(n11980) );
  NAND U12451 ( .A(n12008), .B(n12009), .Z(n12007) );
  XOR U12452 ( .A(n12010), .B(n11959), .Z(n12009) );
  XOR U12453 ( .A(n12000), .B(n12001), .Z(n11959) );
  XOR U12454 ( .A(n12011), .B(n11988), .Z(n12001) );
  XOR U12455 ( .A(n12012), .B(n12013), .Z(n11988) );
  ANDN U12456 ( .B(n12014), .A(n12015), .Z(n12012) );
  XOR U12457 ( .A(n12013), .B(n12016), .Z(n12014) );
  IV U12458 ( .A(n11986), .Z(n12011) );
  XOR U12459 ( .A(n11984), .B(n12017), .Z(n11986) );
  XOR U12460 ( .A(n12018), .B(n12019), .Z(n12017) );
  ANDN U12461 ( .B(n12020), .A(n12021), .Z(n12018) );
  XOR U12462 ( .A(n12022), .B(n12019), .Z(n12020) );
  IV U12463 ( .A(n11987), .Z(n11984) );
  XOR U12464 ( .A(n12023), .B(n12024), .Z(n11987) );
  ANDN U12465 ( .B(n12025), .A(n12026), .Z(n12023) );
  XOR U12466 ( .A(n12024), .B(n12027), .Z(n12025) );
  XOR U12467 ( .A(n12028), .B(n12029), .Z(n12000) );
  XNOR U12468 ( .A(n11995), .B(n12030), .Z(n12029) );
  IV U12469 ( .A(n11998), .Z(n12030) );
  XOR U12470 ( .A(n12031), .B(n12032), .Z(n11998) );
  ANDN U12471 ( .B(n12033), .A(n12034), .Z(n12031) );
  XOR U12472 ( .A(n12032), .B(n12035), .Z(n12033) );
  XNOR U12473 ( .A(n12036), .B(n12037), .Z(n11995) );
  ANDN U12474 ( .B(n12038), .A(n12039), .Z(n12036) );
  XOR U12475 ( .A(n12037), .B(n12040), .Z(n12038) );
  IV U12476 ( .A(n11994), .Z(n12028) );
  XOR U12477 ( .A(n11992), .B(n12041), .Z(n11994) );
  XOR U12478 ( .A(n12042), .B(n12043), .Z(n12041) );
  ANDN U12479 ( .B(n12044), .A(n12045), .Z(n12042) );
  XOR U12480 ( .A(n12046), .B(n12043), .Z(n12044) );
  IV U12481 ( .A(n11996), .Z(n11992) );
  XOR U12482 ( .A(n12047), .B(n12048), .Z(n11996) );
  ANDN U12483 ( .B(n12049), .A(n12050), .Z(n12047) );
  XOR U12484 ( .A(n12051), .B(n12048), .Z(n12049) );
  IV U12485 ( .A(n12006), .Z(n12010) );
  XOR U12486 ( .A(n12006), .B(n11961), .Z(n12008) );
  XOR U12487 ( .A(n12052), .B(n12053), .Z(n11961) );
  AND U12488 ( .A(n266), .B(n12054), .Z(n12052) );
  XOR U12489 ( .A(n12055), .B(n12053), .Z(n12054) );
  NANDN U12490 ( .A(n11963), .B(n11965), .Z(n12006) );
  XOR U12491 ( .A(n12056), .B(n12057), .Z(n11965) );
  AND U12492 ( .A(n266), .B(n12058), .Z(n12056) );
  XOR U12493 ( .A(n12057), .B(n12059), .Z(n12058) );
  XNOR U12494 ( .A(n12060), .B(n12061), .Z(n266) );
  AND U12495 ( .A(n12062), .B(n12063), .Z(n12060) );
  XOR U12496 ( .A(n12061), .B(n11976), .Z(n12063) );
  XNOR U12497 ( .A(n12064), .B(n12065), .Z(n11976) );
  ANDN U12498 ( .B(n12066), .A(n12067), .Z(n12064) );
  XOR U12499 ( .A(n12065), .B(n12068), .Z(n12066) );
  XNOR U12500 ( .A(n12061), .B(n11978), .Z(n12062) );
  XOR U12501 ( .A(n12069), .B(n12070), .Z(n11978) );
  AND U12502 ( .A(n270), .B(n12071), .Z(n12069) );
  XOR U12503 ( .A(n12072), .B(n12070), .Z(n12071) );
  XNOR U12504 ( .A(n12073), .B(n12074), .Z(n12061) );
  AND U12505 ( .A(n12075), .B(n12076), .Z(n12073) );
  XNOR U12506 ( .A(n12074), .B(n12003), .Z(n12076) );
  XOR U12507 ( .A(n12067), .B(n12068), .Z(n12003) );
  XNOR U12508 ( .A(n12077), .B(n12078), .Z(n12068) );
  ANDN U12509 ( .B(n12079), .A(n12080), .Z(n12077) );
  XOR U12510 ( .A(n12081), .B(n12082), .Z(n12079) );
  XOR U12511 ( .A(n12083), .B(n12084), .Z(n12067) );
  XNOR U12512 ( .A(n12085), .B(n12086), .Z(n12084) );
  ANDN U12513 ( .B(n12087), .A(n12088), .Z(n12085) );
  XNOR U12514 ( .A(n12089), .B(n12090), .Z(n12087) );
  IV U12515 ( .A(n12065), .Z(n12083) );
  XOR U12516 ( .A(n12091), .B(n12092), .Z(n12065) );
  ANDN U12517 ( .B(n12093), .A(n12094), .Z(n12091) );
  XOR U12518 ( .A(n12092), .B(n12095), .Z(n12093) );
  XOR U12519 ( .A(n12074), .B(n12005), .Z(n12075) );
  XOR U12520 ( .A(n12096), .B(n12097), .Z(n12005) );
  AND U12521 ( .A(n270), .B(n12098), .Z(n12096) );
  XOR U12522 ( .A(n12099), .B(n12097), .Z(n12098) );
  XNOR U12523 ( .A(n12100), .B(n12101), .Z(n12074) );
  NAND U12524 ( .A(n12102), .B(n12103), .Z(n12101) );
  XOR U12525 ( .A(n12104), .B(n12053), .Z(n12103) );
  XOR U12526 ( .A(n12094), .B(n12095), .Z(n12053) );
  XOR U12527 ( .A(n12105), .B(n12082), .Z(n12095) );
  XOR U12528 ( .A(n12106), .B(n12107), .Z(n12082) );
  ANDN U12529 ( .B(n12108), .A(n12109), .Z(n12106) );
  XOR U12530 ( .A(n12107), .B(n12110), .Z(n12108) );
  IV U12531 ( .A(n12080), .Z(n12105) );
  XOR U12532 ( .A(n12078), .B(n12111), .Z(n12080) );
  XOR U12533 ( .A(n12112), .B(n12113), .Z(n12111) );
  ANDN U12534 ( .B(n12114), .A(n12115), .Z(n12112) );
  XOR U12535 ( .A(n12116), .B(n12113), .Z(n12114) );
  IV U12536 ( .A(n12081), .Z(n12078) );
  XOR U12537 ( .A(n12117), .B(n12118), .Z(n12081) );
  ANDN U12538 ( .B(n12119), .A(n12120), .Z(n12117) );
  XOR U12539 ( .A(n12118), .B(n12121), .Z(n12119) );
  XOR U12540 ( .A(n12122), .B(n12123), .Z(n12094) );
  XNOR U12541 ( .A(n12089), .B(n12124), .Z(n12123) );
  IV U12542 ( .A(n12092), .Z(n12124) );
  XOR U12543 ( .A(n12125), .B(n12126), .Z(n12092) );
  ANDN U12544 ( .B(n12127), .A(n12128), .Z(n12125) );
  XOR U12545 ( .A(n12126), .B(n12129), .Z(n12127) );
  XNOR U12546 ( .A(n12130), .B(n12131), .Z(n12089) );
  ANDN U12547 ( .B(n12132), .A(n12133), .Z(n12130) );
  XOR U12548 ( .A(n12131), .B(n12134), .Z(n12132) );
  IV U12549 ( .A(n12088), .Z(n12122) );
  XOR U12550 ( .A(n12086), .B(n12135), .Z(n12088) );
  XOR U12551 ( .A(n12136), .B(n12137), .Z(n12135) );
  ANDN U12552 ( .B(n12138), .A(n12139), .Z(n12136) );
  XOR U12553 ( .A(n12140), .B(n12137), .Z(n12138) );
  IV U12554 ( .A(n12090), .Z(n12086) );
  XOR U12555 ( .A(n12141), .B(n12142), .Z(n12090) );
  ANDN U12556 ( .B(n12143), .A(n12144), .Z(n12141) );
  XOR U12557 ( .A(n12145), .B(n12142), .Z(n12143) );
  IV U12558 ( .A(n12100), .Z(n12104) );
  XOR U12559 ( .A(n12100), .B(n12055), .Z(n12102) );
  XOR U12560 ( .A(n12146), .B(n12147), .Z(n12055) );
  AND U12561 ( .A(n270), .B(n12148), .Z(n12146) );
  XOR U12562 ( .A(n12149), .B(n12147), .Z(n12148) );
  NANDN U12563 ( .A(n12057), .B(n12059), .Z(n12100) );
  XOR U12564 ( .A(n12150), .B(n12151), .Z(n12059) );
  AND U12565 ( .A(n270), .B(n12152), .Z(n12150) );
  XOR U12566 ( .A(n12151), .B(n12153), .Z(n12152) );
  XNOR U12567 ( .A(n12154), .B(n12155), .Z(n270) );
  AND U12568 ( .A(n12156), .B(n12157), .Z(n12154) );
  XOR U12569 ( .A(n12155), .B(n12070), .Z(n12157) );
  XNOR U12570 ( .A(n12158), .B(n12159), .Z(n12070) );
  ANDN U12571 ( .B(n12160), .A(n12161), .Z(n12158) );
  XOR U12572 ( .A(n12159), .B(n12162), .Z(n12160) );
  XNOR U12573 ( .A(n12155), .B(n12072), .Z(n12156) );
  XOR U12574 ( .A(n12163), .B(n12164), .Z(n12072) );
  AND U12575 ( .A(n274), .B(n12165), .Z(n12163) );
  XOR U12576 ( .A(n12166), .B(n12164), .Z(n12165) );
  XNOR U12577 ( .A(n12167), .B(n12168), .Z(n12155) );
  AND U12578 ( .A(n12169), .B(n12170), .Z(n12167) );
  XNOR U12579 ( .A(n12168), .B(n12097), .Z(n12170) );
  XOR U12580 ( .A(n12161), .B(n12162), .Z(n12097) );
  XNOR U12581 ( .A(n12171), .B(n12172), .Z(n12162) );
  ANDN U12582 ( .B(n12173), .A(n12174), .Z(n12171) );
  XOR U12583 ( .A(n12175), .B(n12176), .Z(n12173) );
  XOR U12584 ( .A(n12177), .B(n12178), .Z(n12161) );
  XNOR U12585 ( .A(n12179), .B(n12180), .Z(n12178) );
  ANDN U12586 ( .B(n12181), .A(n12182), .Z(n12179) );
  XNOR U12587 ( .A(n12183), .B(n12184), .Z(n12181) );
  IV U12588 ( .A(n12159), .Z(n12177) );
  XOR U12589 ( .A(n12185), .B(n12186), .Z(n12159) );
  ANDN U12590 ( .B(n12187), .A(n12188), .Z(n12185) );
  XOR U12591 ( .A(n12186), .B(n12189), .Z(n12187) );
  XOR U12592 ( .A(n12168), .B(n12099), .Z(n12169) );
  XOR U12593 ( .A(n12190), .B(n12191), .Z(n12099) );
  AND U12594 ( .A(n274), .B(n12192), .Z(n12190) );
  XOR U12595 ( .A(n12193), .B(n12191), .Z(n12192) );
  XNOR U12596 ( .A(n12194), .B(n12195), .Z(n12168) );
  NAND U12597 ( .A(n12196), .B(n12197), .Z(n12195) );
  XOR U12598 ( .A(n12198), .B(n12147), .Z(n12197) );
  XOR U12599 ( .A(n12188), .B(n12189), .Z(n12147) );
  XOR U12600 ( .A(n12199), .B(n12176), .Z(n12189) );
  XOR U12601 ( .A(n12200), .B(n12201), .Z(n12176) );
  ANDN U12602 ( .B(n12202), .A(n12203), .Z(n12200) );
  XOR U12603 ( .A(n12201), .B(n12204), .Z(n12202) );
  IV U12604 ( .A(n12174), .Z(n12199) );
  XOR U12605 ( .A(n12172), .B(n12205), .Z(n12174) );
  XOR U12606 ( .A(n12206), .B(n12207), .Z(n12205) );
  ANDN U12607 ( .B(n12208), .A(n12209), .Z(n12206) );
  XOR U12608 ( .A(n12210), .B(n12207), .Z(n12208) );
  IV U12609 ( .A(n12175), .Z(n12172) );
  XOR U12610 ( .A(n12211), .B(n12212), .Z(n12175) );
  ANDN U12611 ( .B(n12213), .A(n12214), .Z(n12211) );
  XOR U12612 ( .A(n12212), .B(n12215), .Z(n12213) );
  XOR U12613 ( .A(n12216), .B(n12217), .Z(n12188) );
  XNOR U12614 ( .A(n12183), .B(n12218), .Z(n12217) );
  IV U12615 ( .A(n12186), .Z(n12218) );
  XOR U12616 ( .A(n12219), .B(n12220), .Z(n12186) );
  ANDN U12617 ( .B(n12221), .A(n12222), .Z(n12219) );
  XOR U12618 ( .A(n12220), .B(n12223), .Z(n12221) );
  XNOR U12619 ( .A(n12224), .B(n12225), .Z(n12183) );
  ANDN U12620 ( .B(n12226), .A(n12227), .Z(n12224) );
  XOR U12621 ( .A(n12225), .B(n12228), .Z(n12226) );
  IV U12622 ( .A(n12182), .Z(n12216) );
  XOR U12623 ( .A(n12180), .B(n12229), .Z(n12182) );
  XOR U12624 ( .A(n12230), .B(n12231), .Z(n12229) );
  ANDN U12625 ( .B(n12232), .A(n12233), .Z(n12230) );
  XOR U12626 ( .A(n12234), .B(n12231), .Z(n12232) );
  IV U12627 ( .A(n12184), .Z(n12180) );
  XOR U12628 ( .A(n12235), .B(n12236), .Z(n12184) );
  ANDN U12629 ( .B(n12237), .A(n12238), .Z(n12235) );
  XOR U12630 ( .A(n12239), .B(n12236), .Z(n12237) );
  IV U12631 ( .A(n12194), .Z(n12198) );
  XOR U12632 ( .A(n12194), .B(n12149), .Z(n12196) );
  XOR U12633 ( .A(n12240), .B(n12241), .Z(n12149) );
  AND U12634 ( .A(n274), .B(n12242), .Z(n12240) );
  XOR U12635 ( .A(n12243), .B(n12241), .Z(n12242) );
  NANDN U12636 ( .A(n12151), .B(n12153), .Z(n12194) );
  XOR U12637 ( .A(n12244), .B(n12245), .Z(n12153) );
  AND U12638 ( .A(n274), .B(n12246), .Z(n12244) );
  XOR U12639 ( .A(n12245), .B(n12247), .Z(n12246) );
  XNOR U12640 ( .A(n12248), .B(n12249), .Z(n274) );
  AND U12641 ( .A(n12250), .B(n12251), .Z(n12248) );
  XOR U12642 ( .A(n12249), .B(n12164), .Z(n12251) );
  XNOR U12643 ( .A(n12252), .B(n12253), .Z(n12164) );
  ANDN U12644 ( .B(n12254), .A(n12255), .Z(n12252) );
  XOR U12645 ( .A(n12253), .B(n12256), .Z(n12254) );
  XNOR U12646 ( .A(n12249), .B(n12166), .Z(n12250) );
  XOR U12647 ( .A(n12257), .B(n12258), .Z(n12166) );
  AND U12648 ( .A(n278), .B(n12259), .Z(n12257) );
  XOR U12649 ( .A(n12260), .B(n12258), .Z(n12259) );
  XNOR U12650 ( .A(n12261), .B(n12262), .Z(n12249) );
  AND U12651 ( .A(n12263), .B(n12264), .Z(n12261) );
  XNOR U12652 ( .A(n12262), .B(n12191), .Z(n12264) );
  XOR U12653 ( .A(n12255), .B(n12256), .Z(n12191) );
  XNOR U12654 ( .A(n12265), .B(n12266), .Z(n12256) );
  ANDN U12655 ( .B(n12267), .A(n12268), .Z(n12265) );
  XOR U12656 ( .A(n12269), .B(n12270), .Z(n12267) );
  XOR U12657 ( .A(n12271), .B(n12272), .Z(n12255) );
  XNOR U12658 ( .A(n12273), .B(n12274), .Z(n12272) );
  ANDN U12659 ( .B(n12275), .A(n12276), .Z(n12273) );
  XNOR U12660 ( .A(n12277), .B(n12278), .Z(n12275) );
  IV U12661 ( .A(n12253), .Z(n12271) );
  XOR U12662 ( .A(n12279), .B(n12280), .Z(n12253) );
  ANDN U12663 ( .B(n12281), .A(n12282), .Z(n12279) );
  XOR U12664 ( .A(n12280), .B(n12283), .Z(n12281) );
  XOR U12665 ( .A(n12262), .B(n12193), .Z(n12263) );
  XOR U12666 ( .A(n12284), .B(n12285), .Z(n12193) );
  AND U12667 ( .A(n278), .B(n12286), .Z(n12284) );
  XOR U12668 ( .A(n12287), .B(n12285), .Z(n12286) );
  XNOR U12669 ( .A(n12288), .B(n12289), .Z(n12262) );
  NAND U12670 ( .A(n12290), .B(n12291), .Z(n12289) );
  XOR U12671 ( .A(n12292), .B(n12241), .Z(n12291) );
  XOR U12672 ( .A(n12282), .B(n12283), .Z(n12241) );
  XOR U12673 ( .A(n12293), .B(n12270), .Z(n12283) );
  XOR U12674 ( .A(n12294), .B(n12295), .Z(n12270) );
  ANDN U12675 ( .B(n12296), .A(n12297), .Z(n12294) );
  XOR U12676 ( .A(n12295), .B(n12298), .Z(n12296) );
  IV U12677 ( .A(n12268), .Z(n12293) );
  XOR U12678 ( .A(n12266), .B(n12299), .Z(n12268) );
  XOR U12679 ( .A(n12300), .B(n12301), .Z(n12299) );
  ANDN U12680 ( .B(n12302), .A(n12303), .Z(n12300) );
  XOR U12681 ( .A(n12304), .B(n12301), .Z(n12302) );
  IV U12682 ( .A(n12269), .Z(n12266) );
  XOR U12683 ( .A(n12305), .B(n12306), .Z(n12269) );
  ANDN U12684 ( .B(n12307), .A(n12308), .Z(n12305) );
  XOR U12685 ( .A(n12306), .B(n12309), .Z(n12307) );
  XOR U12686 ( .A(n12310), .B(n12311), .Z(n12282) );
  XNOR U12687 ( .A(n12277), .B(n12312), .Z(n12311) );
  IV U12688 ( .A(n12280), .Z(n12312) );
  XOR U12689 ( .A(n12313), .B(n12314), .Z(n12280) );
  ANDN U12690 ( .B(n12315), .A(n12316), .Z(n12313) );
  XOR U12691 ( .A(n12314), .B(n12317), .Z(n12315) );
  XNOR U12692 ( .A(n12318), .B(n12319), .Z(n12277) );
  ANDN U12693 ( .B(n12320), .A(n12321), .Z(n12318) );
  XOR U12694 ( .A(n12319), .B(n12322), .Z(n12320) );
  IV U12695 ( .A(n12276), .Z(n12310) );
  XOR U12696 ( .A(n12274), .B(n12323), .Z(n12276) );
  XOR U12697 ( .A(n12324), .B(n12325), .Z(n12323) );
  ANDN U12698 ( .B(n12326), .A(n12327), .Z(n12324) );
  XOR U12699 ( .A(n12328), .B(n12325), .Z(n12326) );
  IV U12700 ( .A(n12278), .Z(n12274) );
  XOR U12701 ( .A(n12329), .B(n12330), .Z(n12278) );
  ANDN U12702 ( .B(n12331), .A(n12332), .Z(n12329) );
  XOR U12703 ( .A(n12333), .B(n12330), .Z(n12331) );
  IV U12704 ( .A(n12288), .Z(n12292) );
  XOR U12705 ( .A(n12288), .B(n12243), .Z(n12290) );
  XOR U12706 ( .A(n12334), .B(n12335), .Z(n12243) );
  AND U12707 ( .A(n278), .B(n12336), .Z(n12334) );
  XOR U12708 ( .A(n12337), .B(n12335), .Z(n12336) );
  NANDN U12709 ( .A(n12245), .B(n12247), .Z(n12288) );
  XOR U12710 ( .A(n12338), .B(n12339), .Z(n12247) );
  AND U12711 ( .A(n278), .B(n12340), .Z(n12338) );
  XOR U12712 ( .A(n12339), .B(n12341), .Z(n12340) );
  XNOR U12713 ( .A(n12342), .B(n12343), .Z(n278) );
  AND U12714 ( .A(n12344), .B(n12345), .Z(n12342) );
  XOR U12715 ( .A(n12343), .B(n12258), .Z(n12345) );
  XNOR U12716 ( .A(n12346), .B(n12347), .Z(n12258) );
  ANDN U12717 ( .B(n12348), .A(n12349), .Z(n12346) );
  XOR U12718 ( .A(n12347), .B(n12350), .Z(n12348) );
  XNOR U12719 ( .A(n12343), .B(n12260), .Z(n12344) );
  XOR U12720 ( .A(n12351), .B(n12352), .Z(n12260) );
  AND U12721 ( .A(n282), .B(n12353), .Z(n12351) );
  XOR U12722 ( .A(n12354), .B(n12352), .Z(n12353) );
  XNOR U12723 ( .A(n12355), .B(n12356), .Z(n12343) );
  AND U12724 ( .A(n12357), .B(n12358), .Z(n12355) );
  XNOR U12725 ( .A(n12356), .B(n12285), .Z(n12358) );
  XOR U12726 ( .A(n12349), .B(n12350), .Z(n12285) );
  XNOR U12727 ( .A(n12359), .B(n12360), .Z(n12350) );
  ANDN U12728 ( .B(n12361), .A(n12362), .Z(n12359) );
  XOR U12729 ( .A(n12363), .B(n12364), .Z(n12361) );
  XOR U12730 ( .A(n12365), .B(n12366), .Z(n12349) );
  XNOR U12731 ( .A(n12367), .B(n12368), .Z(n12366) );
  ANDN U12732 ( .B(n12369), .A(n12370), .Z(n12367) );
  XNOR U12733 ( .A(n12371), .B(n12372), .Z(n12369) );
  IV U12734 ( .A(n12347), .Z(n12365) );
  XOR U12735 ( .A(n12373), .B(n12374), .Z(n12347) );
  ANDN U12736 ( .B(n12375), .A(n12376), .Z(n12373) );
  XOR U12737 ( .A(n12374), .B(n12377), .Z(n12375) );
  XOR U12738 ( .A(n12356), .B(n12287), .Z(n12357) );
  XOR U12739 ( .A(n12378), .B(n12379), .Z(n12287) );
  AND U12740 ( .A(n282), .B(n12380), .Z(n12378) );
  XOR U12741 ( .A(n12381), .B(n12379), .Z(n12380) );
  XNOR U12742 ( .A(n12382), .B(n12383), .Z(n12356) );
  NAND U12743 ( .A(n12384), .B(n12385), .Z(n12383) );
  XOR U12744 ( .A(n12386), .B(n12335), .Z(n12385) );
  XOR U12745 ( .A(n12376), .B(n12377), .Z(n12335) );
  XOR U12746 ( .A(n12387), .B(n12364), .Z(n12377) );
  XOR U12747 ( .A(n12388), .B(n12389), .Z(n12364) );
  ANDN U12748 ( .B(n12390), .A(n12391), .Z(n12388) );
  XOR U12749 ( .A(n12389), .B(n12392), .Z(n12390) );
  IV U12750 ( .A(n12362), .Z(n12387) );
  XOR U12751 ( .A(n12360), .B(n12393), .Z(n12362) );
  XOR U12752 ( .A(n12394), .B(n12395), .Z(n12393) );
  ANDN U12753 ( .B(n12396), .A(n12397), .Z(n12394) );
  XOR U12754 ( .A(n12398), .B(n12395), .Z(n12396) );
  IV U12755 ( .A(n12363), .Z(n12360) );
  XOR U12756 ( .A(n12399), .B(n12400), .Z(n12363) );
  ANDN U12757 ( .B(n12401), .A(n12402), .Z(n12399) );
  XOR U12758 ( .A(n12400), .B(n12403), .Z(n12401) );
  XOR U12759 ( .A(n12404), .B(n12405), .Z(n12376) );
  XNOR U12760 ( .A(n12371), .B(n12406), .Z(n12405) );
  IV U12761 ( .A(n12374), .Z(n12406) );
  XOR U12762 ( .A(n12407), .B(n12408), .Z(n12374) );
  ANDN U12763 ( .B(n12409), .A(n12410), .Z(n12407) );
  XOR U12764 ( .A(n12408), .B(n12411), .Z(n12409) );
  XNOR U12765 ( .A(n12412), .B(n12413), .Z(n12371) );
  ANDN U12766 ( .B(n12414), .A(n12415), .Z(n12412) );
  XOR U12767 ( .A(n12413), .B(n12416), .Z(n12414) );
  IV U12768 ( .A(n12370), .Z(n12404) );
  XOR U12769 ( .A(n12368), .B(n12417), .Z(n12370) );
  XOR U12770 ( .A(n12418), .B(n12419), .Z(n12417) );
  ANDN U12771 ( .B(n12420), .A(n12421), .Z(n12418) );
  XOR U12772 ( .A(n12422), .B(n12419), .Z(n12420) );
  IV U12773 ( .A(n12372), .Z(n12368) );
  XOR U12774 ( .A(n12423), .B(n12424), .Z(n12372) );
  ANDN U12775 ( .B(n12425), .A(n12426), .Z(n12423) );
  XOR U12776 ( .A(n12427), .B(n12424), .Z(n12425) );
  IV U12777 ( .A(n12382), .Z(n12386) );
  XOR U12778 ( .A(n12382), .B(n12337), .Z(n12384) );
  XOR U12779 ( .A(n12428), .B(n12429), .Z(n12337) );
  AND U12780 ( .A(n282), .B(n12430), .Z(n12428) );
  XOR U12781 ( .A(n12431), .B(n12429), .Z(n12430) );
  NANDN U12782 ( .A(n12339), .B(n12341), .Z(n12382) );
  XOR U12783 ( .A(n12432), .B(n12433), .Z(n12341) );
  AND U12784 ( .A(n282), .B(n12434), .Z(n12432) );
  XOR U12785 ( .A(n12433), .B(n12435), .Z(n12434) );
  XNOR U12786 ( .A(n12436), .B(n12437), .Z(n282) );
  AND U12787 ( .A(n12438), .B(n12439), .Z(n12436) );
  XOR U12788 ( .A(n12437), .B(n12352), .Z(n12439) );
  XNOR U12789 ( .A(n12440), .B(n12441), .Z(n12352) );
  ANDN U12790 ( .B(n12442), .A(n12443), .Z(n12440) );
  XOR U12791 ( .A(n12441), .B(n12444), .Z(n12442) );
  XNOR U12792 ( .A(n12437), .B(n12354), .Z(n12438) );
  XOR U12793 ( .A(n12445), .B(n12446), .Z(n12354) );
  AND U12794 ( .A(n286), .B(n12447), .Z(n12445) );
  XOR U12795 ( .A(n12448), .B(n12446), .Z(n12447) );
  XNOR U12796 ( .A(n12449), .B(n12450), .Z(n12437) );
  AND U12797 ( .A(n12451), .B(n12452), .Z(n12449) );
  XNOR U12798 ( .A(n12450), .B(n12379), .Z(n12452) );
  XOR U12799 ( .A(n12443), .B(n12444), .Z(n12379) );
  XNOR U12800 ( .A(n12453), .B(n12454), .Z(n12444) );
  ANDN U12801 ( .B(n12455), .A(n12456), .Z(n12453) );
  XOR U12802 ( .A(n12457), .B(n12458), .Z(n12455) );
  XOR U12803 ( .A(n12459), .B(n12460), .Z(n12443) );
  XNOR U12804 ( .A(n12461), .B(n12462), .Z(n12460) );
  ANDN U12805 ( .B(n12463), .A(n12464), .Z(n12461) );
  XNOR U12806 ( .A(n12465), .B(n12466), .Z(n12463) );
  IV U12807 ( .A(n12441), .Z(n12459) );
  XOR U12808 ( .A(n12467), .B(n12468), .Z(n12441) );
  ANDN U12809 ( .B(n12469), .A(n12470), .Z(n12467) );
  XOR U12810 ( .A(n12468), .B(n12471), .Z(n12469) );
  XOR U12811 ( .A(n12450), .B(n12381), .Z(n12451) );
  XOR U12812 ( .A(n12472), .B(n12473), .Z(n12381) );
  AND U12813 ( .A(n286), .B(n12474), .Z(n12472) );
  XOR U12814 ( .A(n12475), .B(n12473), .Z(n12474) );
  XNOR U12815 ( .A(n12476), .B(n12477), .Z(n12450) );
  NAND U12816 ( .A(n12478), .B(n12479), .Z(n12477) );
  XOR U12817 ( .A(n12480), .B(n12429), .Z(n12479) );
  XOR U12818 ( .A(n12470), .B(n12471), .Z(n12429) );
  XOR U12819 ( .A(n12481), .B(n12458), .Z(n12471) );
  XOR U12820 ( .A(n12482), .B(n12483), .Z(n12458) );
  ANDN U12821 ( .B(n12484), .A(n12485), .Z(n12482) );
  XOR U12822 ( .A(n12483), .B(n12486), .Z(n12484) );
  IV U12823 ( .A(n12456), .Z(n12481) );
  XOR U12824 ( .A(n12454), .B(n12487), .Z(n12456) );
  XOR U12825 ( .A(n12488), .B(n12489), .Z(n12487) );
  ANDN U12826 ( .B(n12490), .A(n12491), .Z(n12488) );
  XOR U12827 ( .A(n12492), .B(n12489), .Z(n12490) );
  IV U12828 ( .A(n12457), .Z(n12454) );
  XOR U12829 ( .A(n12493), .B(n12494), .Z(n12457) );
  ANDN U12830 ( .B(n12495), .A(n12496), .Z(n12493) );
  XOR U12831 ( .A(n12494), .B(n12497), .Z(n12495) );
  XOR U12832 ( .A(n12498), .B(n12499), .Z(n12470) );
  XNOR U12833 ( .A(n12465), .B(n12500), .Z(n12499) );
  IV U12834 ( .A(n12468), .Z(n12500) );
  XOR U12835 ( .A(n12501), .B(n12502), .Z(n12468) );
  ANDN U12836 ( .B(n12503), .A(n12504), .Z(n12501) );
  XOR U12837 ( .A(n12502), .B(n12505), .Z(n12503) );
  XNOR U12838 ( .A(n12506), .B(n12507), .Z(n12465) );
  ANDN U12839 ( .B(n12508), .A(n12509), .Z(n12506) );
  XOR U12840 ( .A(n12507), .B(n12510), .Z(n12508) );
  IV U12841 ( .A(n12464), .Z(n12498) );
  XOR U12842 ( .A(n12462), .B(n12511), .Z(n12464) );
  XOR U12843 ( .A(n12512), .B(n12513), .Z(n12511) );
  ANDN U12844 ( .B(n12514), .A(n12515), .Z(n12512) );
  XOR U12845 ( .A(n12516), .B(n12513), .Z(n12514) );
  IV U12846 ( .A(n12466), .Z(n12462) );
  XOR U12847 ( .A(n12517), .B(n12518), .Z(n12466) );
  ANDN U12848 ( .B(n12519), .A(n12520), .Z(n12517) );
  XOR U12849 ( .A(n12521), .B(n12518), .Z(n12519) );
  IV U12850 ( .A(n12476), .Z(n12480) );
  XOR U12851 ( .A(n12476), .B(n12431), .Z(n12478) );
  XOR U12852 ( .A(n12522), .B(n12523), .Z(n12431) );
  AND U12853 ( .A(n286), .B(n12524), .Z(n12522) );
  XOR U12854 ( .A(n12525), .B(n12523), .Z(n12524) );
  NANDN U12855 ( .A(n12433), .B(n12435), .Z(n12476) );
  XOR U12856 ( .A(n12526), .B(n12527), .Z(n12435) );
  AND U12857 ( .A(n286), .B(n12528), .Z(n12526) );
  XOR U12858 ( .A(n12527), .B(n12529), .Z(n12528) );
  XNOR U12859 ( .A(n12530), .B(n12531), .Z(n286) );
  AND U12860 ( .A(n12532), .B(n12533), .Z(n12530) );
  XOR U12861 ( .A(n12531), .B(n12446), .Z(n12533) );
  XNOR U12862 ( .A(n12534), .B(n12535), .Z(n12446) );
  ANDN U12863 ( .B(n12536), .A(n12537), .Z(n12534) );
  XOR U12864 ( .A(n12535), .B(n12538), .Z(n12536) );
  XNOR U12865 ( .A(n12531), .B(n12448), .Z(n12532) );
  XOR U12866 ( .A(n12539), .B(n12540), .Z(n12448) );
  AND U12867 ( .A(n290), .B(n12541), .Z(n12539) );
  XOR U12868 ( .A(n12542), .B(n12540), .Z(n12541) );
  XNOR U12869 ( .A(n12543), .B(n12544), .Z(n12531) );
  AND U12870 ( .A(n12545), .B(n12546), .Z(n12543) );
  XNOR U12871 ( .A(n12544), .B(n12473), .Z(n12546) );
  XOR U12872 ( .A(n12537), .B(n12538), .Z(n12473) );
  XNOR U12873 ( .A(n12547), .B(n12548), .Z(n12538) );
  ANDN U12874 ( .B(n12549), .A(n12550), .Z(n12547) );
  XOR U12875 ( .A(n12551), .B(n12552), .Z(n12549) );
  XOR U12876 ( .A(n12553), .B(n12554), .Z(n12537) );
  XNOR U12877 ( .A(n12555), .B(n12556), .Z(n12554) );
  ANDN U12878 ( .B(n12557), .A(n12558), .Z(n12555) );
  XNOR U12879 ( .A(n12559), .B(n12560), .Z(n12557) );
  IV U12880 ( .A(n12535), .Z(n12553) );
  XOR U12881 ( .A(n12561), .B(n12562), .Z(n12535) );
  ANDN U12882 ( .B(n12563), .A(n12564), .Z(n12561) );
  XOR U12883 ( .A(n12562), .B(n12565), .Z(n12563) );
  XOR U12884 ( .A(n12544), .B(n12475), .Z(n12545) );
  XOR U12885 ( .A(n12566), .B(n12567), .Z(n12475) );
  AND U12886 ( .A(n290), .B(n12568), .Z(n12566) );
  XOR U12887 ( .A(n12569), .B(n12567), .Z(n12568) );
  XNOR U12888 ( .A(n12570), .B(n12571), .Z(n12544) );
  NAND U12889 ( .A(n12572), .B(n12573), .Z(n12571) );
  XOR U12890 ( .A(n12574), .B(n12523), .Z(n12573) );
  XOR U12891 ( .A(n12564), .B(n12565), .Z(n12523) );
  XOR U12892 ( .A(n12575), .B(n12552), .Z(n12565) );
  XOR U12893 ( .A(n12576), .B(n12577), .Z(n12552) );
  ANDN U12894 ( .B(n12578), .A(n12579), .Z(n12576) );
  XOR U12895 ( .A(n12577), .B(n12580), .Z(n12578) );
  IV U12896 ( .A(n12550), .Z(n12575) );
  XOR U12897 ( .A(n12548), .B(n12581), .Z(n12550) );
  XOR U12898 ( .A(n12582), .B(n12583), .Z(n12581) );
  ANDN U12899 ( .B(n12584), .A(n12585), .Z(n12582) );
  XOR U12900 ( .A(n12586), .B(n12583), .Z(n12584) );
  IV U12901 ( .A(n12551), .Z(n12548) );
  XOR U12902 ( .A(n12587), .B(n12588), .Z(n12551) );
  ANDN U12903 ( .B(n12589), .A(n12590), .Z(n12587) );
  XOR U12904 ( .A(n12588), .B(n12591), .Z(n12589) );
  XOR U12905 ( .A(n12592), .B(n12593), .Z(n12564) );
  XNOR U12906 ( .A(n12559), .B(n12594), .Z(n12593) );
  IV U12907 ( .A(n12562), .Z(n12594) );
  XOR U12908 ( .A(n12595), .B(n12596), .Z(n12562) );
  ANDN U12909 ( .B(n12597), .A(n12598), .Z(n12595) );
  XOR U12910 ( .A(n12596), .B(n12599), .Z(n12597) );
  XNOR U12911 ( .A(n12600), .B(n12601), .Z(n12559) );
  ANDN U12912 ( .B(n12602), .A(n12603), .Z(n12600) );
  XOR U12913 ( .A(n12601), .B(n12604), .Z(n12602) );
  IV U12914 ( .A(n12558), .Z(n12592) );
  XOR U12915 ( .A(n12556), .B(n12605), .Z(n12558) );
  XOR U12916 ( .A(n12606), .B(n12607), .Z(n12605) );
  ANDN U12917 ( .B(n12608), .A(n12609), .Z(n12606) );
  XOR U12918 ( .A(n12610), .B(n12607), .Z(n12608) );
  IV U12919 ( .A(n12560), .Z(n12556) );
  XOR U12920 ( .A(n12611), .B(n12612), .Z(n12560) );
  ANDN U12921 ( .B(n12613), .A(n12614), .Z(n12611) );
  XOR U12922 ( .A(n12615), .B(n12612), .Z(n12613) );
  IV U12923 ( .A(n12570), .Z(n12574) );
  XOR U12924 ( .A(n12570), .B(n12525), .Z(n12572) );
  XOR U12925 ( .A(n12616), .B(n12617), .Z(n12525) );
  AND U12926 ( .A(n290), .B(n12618), .Z(n12616) );
  XOR U12927 ( .A(n12619), .B(n12617), .Z(n12618) );
  NANDN U12928 ( .A(n12527), .B(n12529), .Z(n12570) );
  XOR U12929 ( .A(n12620), .B(n12621), .Z(n12529) );
  AND U12930 ( .A(n290), .B(n12622), .Z(n12620) );
  XOR U12931 ( .A(n12621), .B(n12623), .Z(n12622) );
  XNOR U12932 ( .A(n12624), .B(n12625), .Z(n290) );
  AND U12933 ( .A(n12626), .B(n12627), .Z(n12624) );
  XOR U12934 ( .A(n12625), .B(n12540), .Z(n12627) );
  XNOR U12935 ( .A(n12628), .B(n12629), .Z(n12540) );
  ANDN U12936 ( .B(n12630), .A(n12631), .Z(n12628) );
  XOR U12937 ( .A(n12629), .B(n12632), .Z(n12630) );
  XNOR U12938 ( .A(n12625), .B(n12542), .Z(n12626) );
  XOR U12939 ( .A(n12633), .B(n12634), .Z(n12542) );
  AND U12940 ( .A(n294), .B(n12635), .Z(n12633) );
  XOR U12941 ( .A(n12636), .B(n12634), .Z(n12635) );
  XNOR U12942 ( .A(n12637), .B(n12638), .Z(n12625) );
  AND U12943 ( .A(n12639), .B(n12640), .Z(n12637) );
  XNOR U12944 ( .A(n12638), .B(n12567), .Z(n12640) );
  XOR U12945 ( .A(n12631), .B(n12632), .Z(n12567) );
  XNOR U12946 ( .A(n12641), .B(n12642), .Z(n12632) );
  ANDN U12947 ( .B(n12643), .A(n12644), .Z(n12641) );
  XOR U12948 ( .A(n12645), .B(n12646), .Z(n12643) );
  XOR U12949 ( .A(n12647), .B(n12648), .Z(n12631) );
  XNOR U12950 ( .A(n12649), .B(n12650), .Z(n12648) );
  ANDN U12951 ( .B(n12651), .A(n12652), .Z(n12649) );
  XNOR U12952 ( .A(n12653), .B(n12654), .Z(n12651) );
  IV U12953 ( .A(n12629), .Z(n12647) );
  XOR U12954 ( .A(n12655), .B(n12656), .Z(n12629) );
  ANDN U12955 ( .B(n12657), .A(n12658), .Z(n12655) );
  XOR U12956 ( .A(n12656), .B(n12659), .Z(n12657) );
  XOR U12957 ( .A(n12638), .B(n12569), .Z(n12639) );
  XOR U12958 ( .A(n12660), .B(n12661), .Z(n12569) );
  AND U12959 ( .A(n294), .B(n12662), .Z(n12660) );
  XOR U12960 ( .A(n12663), .B(n12661), .Z(n12662) );
  XNOR U12961 ( .A(n12664), .B(n12665), .Z(n12638) );
  NAND U12962 ( .A(n12666), .B(n12667), .Z(n12665) );
  XOR U12963 ( .A(n12668), .B(n12617), .Z(n12667) );
  XOR U12964 ( .A(n12658), .B(n12659), .Z(n12617) );
  XOR U12965 ( .A(n12669), .B(n12646), .Z(n12659) );
  XOR U12966 ( .A(n12670), .B(n12671), .Z(n12646) );
  ANDN U12967 ( .B(n12672), .A(n12673), .Z(n12670) );
  XOR U12968 ( .A(n12671), .B(n12674), .Z(n12672) );
  IV U12969 ( .A(n12644), .Z(n12669) );
  XOR U12970 ( .A(n12642), .B(n12675), .Z(n12644) );
  XOR U12971 ( .A(n12676), .B(n12677), .Z(n12675) );
  ANDN U12972 ( .B(n12678), .A(n12679), .Z(n12676) );
  XOR U12973 ( .A(n12680), .B(n12677), .Z(n12678) );
  IV U12974 ( .A(n12645), .Z(n12642) );
  XOR U12975 ( .A(n12681), .B(n12682), .Z(n12645) );
  ANDN U12976 ( .B(n12683), .A(n12684), .Z(n12681) );
  XOR U12977 ( .A(n12682), .B(n12685), .Z(n12683) );
  XOR U12978 ( .A(n12686), .B(n12687), .Z(n12658) );
  XNOR U12979 ( .A(n12653), .B(n12688), .Z(n12687) );
  IV U12980 ( .A(n12656), .Z(n12688) );
  XOR U12981 ( .A(n12689), .B(n12690), .Z(n12656) );
  ANDN U12982 ( .B(n12691), .A(n12692), .Z(n12689) );
  XOR U12983 ( .A(n12690), .B(n12693), .Z(n12691) );
  XNOR U12984 ( .A(n12694), .B(n12695), .Z(n12653) );
  ANDN U12985 ( .B(n12696), .A(n12697), .Z(n12694) );
  XOR U12986 ( .A(n12695), .B(n12698), .Z(n12696) );
  IV U12987 ( .A(n12652), .Z(n12686) );
  XOR U12988 ( .A(n12650), .B(n12699), .Z(n12652) );
  XOR U12989 ( .A(n12700), .B(n12701), .Z(n12699) );
  ANDN U12990 ( .B(n12702), .A(n12703), .Z(n12700) );
  XOR U12991 ( .A(n12704), .B(n12701), .Z(n12702) );
  IV U12992 ( .A(n12654), .Z(n12650) );
  XOR U12993 ( .A(n12705), .B(n12706), .Z(n12654) );
  ANDN U12994 ( .B(n12707), .A(n12708), .Z(n12705) );
  XOR U12995 ( .A(n12709), .B(n12706), .Z(n12707) );
  IV U12996 ( .A(n12664), .Z(n12668) );
  XOR U12997 ( .A(n12664), .B(n12619), .Z(n12666) );
  XOR U12998 ( .A(n12710), .B(n12711), .Z(n12619) );
  AND U12999 ( .A(n294), .B(n12712), .Z(n12710) );
  XOR U13000 ( .A(n12713), .B(n12711), .Z(n12712) );
  NANDN U13001 ( .A(n12621), .B(n12623), .Z(n12664) );
  XOR U13002 ( .A(n12714), .B(n12715), .Z(n12623) );
  AND U13003 ( .A(n294), .B(n12716), .Z(n12714) );
  XOR U13004 ( .A(n12715), .B(n12717), .Z(n12716) );
  XNOR U13005 ( .A(n12718), .B(n12719), .Z(n294) );
  AND U13006 ( .A(n12720), .B(n12721), .Z(n12718) );
  XOR U13007 ( .A(n12719), .B(n12634), .Z(n12721) );
  XNOR U13008 ( .A(n12722), .B(n12723), .Z(n12634) );
  ANDN U13009 ( .B(n12724), .A(n12725), .Z(n12722) );
  XOR U13010 ( .A(n12723), .B(n12726), .Z(n12724) );
  XNOR U13011 ( .A(n12719), .B(n12636), .Z(n12720) );
  XOR U13012 ( .A(n12727), .B(n12728), .Z(n12636) );
  AND U13013 ( .A(n298), .B(n12729), .Z(n12727) );
  XOR U13014 ( .A(n12730), .B(n12728), .Z(n12729) );
  XNOR U13015 ( .A(n12731), .B(n12732), .Z(n12719) );
  AND U13016 ( .A(n12733), .B(n12734), .Z(n12731) );
  XNOR U13017 ( .A(n12732), .B(n12661), .Z(n12734) );
  XOR U13018 ( .A(n12725), .B(n12726), .Z(n12661) );
  XNOR U13019 ( .A(n12735), .B(n12736), .Z(n12726) );
  ANDN U13020 ( .B(n12737), .A(n12738), .Z(n12735) );
  XOR U13021 ( .A(n12739), .B(n12740), .Z(n12737) );
  XOR U13022 ( .A(n12741), .B(n12742), .Z(n12725) );
  XNOR U13023 ( .A(n12743), .B(n12744), .Z(n12742) );
  ANDN U13024 ( .B(n12745), .A(n12746), .Z(n12743) );
  XNOR U13025 ( .A(n12747), .B(n12748), .Z(n12745) );
  IV U13026 ( .A(n12723), .Z(n12741) );
  XOR U13027 ( .A(n12749), .B(n12750), .Z(n12723) );
  ANDN U13028 ( .B(n12751), .A(n12752), .Z(n12749) );
  XOR U13029 ( .A(n12750), .B(n12753), .Z(n12751) );
  XOR U13030 ( .A(n12732), .B(n12663), .Z(n12733) );
  XOR U13031 ( .A(n12754), .B(n12755), .Z(n12663) );
  AND U13032 ( .A(n298), .B(n12756), .Z(n12754) );
  XOR U13033 ( .A(n12757), .B(n12755), .Z(n12756) );
  XNOR U13034 ( .A(n12758), .B(n12759), .Z(n12732) );
  NAND U13035 ( .A(n12760), .B(n12761), .Z(n12759) );
  XOR U13036 ( .A(n12762), .B(n12711), .Z(n12761) );
  XOR U13037 ( .A(n12752), .B(n12753), .Z(n12711) );
  XOR U13038 ( .A(n12763), .B(n12740), .Z(n12753) );
  XOR U13039 ( .A(n12764), .B(n12765), .Z(n12740) );
  ANDN U13040 ( .B(n12766), .A(n12767), .Z(n12764) );
  XOR U13041 ( .A(n12765), .B(n12768), .Z(n12766) );
  IV U13042 ( .A(n12738), .Z(n12763) );
  XOR U13043 ( .A(n12736), .B(n12769), .Z(n12738) );
  XOR U13044 ( .A(n12770), .B(n12771), .Z(n12769) );
  ANDN U13045 ( .B(n12772), .A(n12773), .Z(n12770) );
  XOR U13046 ( .A(n12774), .B(n12771), .Z(n12772) );
  IV U13047 ( .A(n12739), .Z(n12736) );
  XOR U13048 ( .A(n12775), .B(n12776), .Z(n12739) );
  ANDN U13049 ( .B(n12777), .A(n12778), .Z(n12775) );
  XOR U13050 ( .A(n12776), .B(n12779), .Z(n12777) );
  XOR U13051 ( .A(n12780), .B(n12781), .Z(n12752) );
  XNOR U13052 ( .A(n12747), .B(n12782), .Z(n12781) );
  IV U13053 ( .A(n12750), .Z(n12782) );
  XOR U13054 ( .A(n12783), .B(n12784), .Z(n12750) );
  ANDN U13055 ( .B(n12785), .A(n12786), .Z(n12783) );
  XOR U13056 ( .A(n12784), .B(n12787), .Z(n12785) );
  XNOR U13057 ( .A(n12788), .B(n12789), .Z(n12747) );
  ANDN U13058 ( .B(n12790), .A(n12791), .Z(n12788) );
  XOR U13059 ( .A(n12789), .B(n12792), .Z(n12790) );
  IV U13060 ( .A(n12746), .Z(n12780) );
  XOR U13061 ( .A(n12744), .B(n12793), .Z(n12746) );
  XOR U13062 ( .A(n12794), .B(n12795), .Z(n12793) );
  ANDN U13063 ( .B(n12796), .A(n12797), .Z(n12794) );
  XOR U13064 ( .A(n12798), .B(n12795), .Z(n12796) );
  IV U13065 ( .A(n12748), .Z(n12744) );
  XOR U13066 ( .A(n12799), .B(n12800), .Z(n12748) );
  ANDN U13067 ( .B(n12801), .A(n12802), .Z(n12799) );
  XOR U13068 ( .A(n12803), .B(n12800), .Z(n12801) );
  IV U13069 ( .A(n12758), .Z(n12762) );
  XOR U13070 ( .A(n12758), .B(n12713), .Z(n12760) );
  XOR U13071 ( .A(n12804), .B(n12805), .Z(n12713) );
  AND U13072 ( .A(n298), .B(n12806), .Z(n12804) );
  XOR U13073 ( .A(n12807), .B(n12805), .Z(n12806) );
  NANDN U13074 ( .A(n12715), .B(n12717), .Z(n12758) );
  XOR U13075 ( .A(n12808), .B(n12809), .Z(n12717) );
  AND U13076 ( .A(n298), .B(n12810), .Z(n12808) );
  XOR U13077 ( .A(n12809), .B(n12811), .Z(n12810) );
  XNOR U13078 ( .A(n12812), .B(n12813), .Z(n298) );
  AND U13079 ( .A(n12814), .B(n12815), .Z(n12812) );
  XOR U13080 ( .A(n12813), .B(n12728), .Z(n12815) );
  XNOR U13081 ( .A(n12816), .B(n12817), .Z(n12728) );
  ANDN U13082 ( .B(n12818), .A(n12819), .Z(n12816) );
  XOR U13083 ( .A(n12817), .B(n12820), .Z(n12818) );
  XNOR U13084 ( .A(n12813), .B(n12730), .Z(n12814) );
  XOR U13085 ( .A(n12821), .B(n12822), .Z(n12730) );
  AND U13086 ( .A(n302), .B(n12823), .Z(n12821) );
  XOR U13087 ( .A(n12824), .B(n12822), .Z(n12823) );
  XNOR U13088 ( .A(n12825), .B(n12826), .Z(n12813) );
  AND U13089 ( .A(n12827), .B(n12828), .Z(n12825) );
  XNOR U13090 ( .A(n12826), .B(n12755), .Z(n12828) );
  XOR U13091 ( .A(n12819), .B(n12820), .Z(n12755) );
  XNOR U13092 ( .A(n12829), .B(n12830), .Z(n12820) );
  ANDN U13093 ( .B(n12831), .A(n12832), .Z(n12829) );
  XOR U13094 ( .A(n12833), .B(n12834), .Z(n12831) );
  XOR U13095 ( .A(n12835), .B(n12836), .Z(n12819) );
  XNOR U13096 ( .A(n12837), .B(n12838), .Z(n12836) );
  ANDN U13097 ( .B(n12839), .A(n12840), .Z(n12837) );
  XNOR U13098 ( .A(n12841), .B(n12842), .Z(n12839) );
  IV U13099 ( .A(n12817), .Z(n12835) );
  XOR U13100 ( .A(n12843), .B(n12844), .Z(n12817) );
  ANDN U13101 ( .B(n12845), .A(n12846), .Z(n12843) );
  XOR U13102 ( .A(n12844), .B(n12847), .Z(n12845) );
  XOR U13103 ( .A(n12826), .B(n12757), .Z(n12827) );
  XOR U13104 ( .A(n12848), .B(n12849), .Z(n12757) );
  AND U13105 ( .A(n302), .B(n12850), .Z(n12848) );
  XOR U13106 ( .A(n12851), .B(n12849), .Z(n12850) );
  XNOR U13107 ( .A(n12852), .B(n12853), .Z(n12826) );
  NAND U13108 ( .A(n12854), .B(n12855), .Z(n12853) );
  XOR U13109 ( .A(n12856), .B(n12805), .Z(n12855) );
  XOR U13110 ( .A(n12846), .B(n12847), .Z(n12805) );
  XOR U13111 ( .A(n12857), .B(n12834), .Z(n12847) );
  XOR U13112 ( .A(n12858), .B(n12859), .Z(n12834) );
  ANDN U13113 ( .B(n12860), .A(n12861), .Z(n12858) );
  XOR U13114 ( .A(n12859), .B(n12862), .Z(n12860) );
  IV U13115 ( .A(n12832), .Z(n12857) );
  XOR U13116 ( .A(n12830), .B(n12863), .Z(n12832) );
  XOR U13117 ( .A(n12864), .B(n12865), .Z(n12863) );
  ANDN U13118 ( .B(n12866), .A(n12867), .Z(n12864) );
  XOR U13119 ( .A(n12868), .B(n12865), .Z(n12866) );
  IV U13120 ( .A(n12833), .Z(n12830) );
  XOR U13121 ( .A(n12869), .B(n12870), .Z(n12833) );
  ANDN U13122 ( .B(n12871), .A(n12872), .Z(n12869) );
  XOR U13123 ( .A(n12870), .B(n12873), .Z(n12871) );
  XOR U13124 ( .A(n12874), .B(n12875), .Z(n12846) );
  XNOR U13125 ( .A(n12841), .B(n12876), .Z(n12875) );
  IV U13126 ( .A(n12844), .Z(n12876) );
  XOR U13127 ( .A(n12877), .B(n12878), .Z(n12844) );
  ANDN U13128 ( .B(n12879), .A(n12880), .Z(n12877) );
  XOR U13129 ( .A(n12878), .B(n12881), .Z(n12879) );
  XNOR U13130 ( .A(n12882), .B(n12883), .Z(n12841) );
  ANDN U13131 ( .B(n12884), .A(n12885), .Z(n12882) );
  XOR U13132 ( .A(n12883), .B(n12886), .Z(n12884) );
  IV U13133 ( .A(n12840), .Z(n12874) );
  XOR U13134 ( .A(n12838), .B(n12887), .Z(n12840) );
  XOR U13135 ( .A(n12888), .B(n12889), .Z(n12887) );
  ANDN U13136 ( .B(n12890), .A(n12891), .Z(n12888) );
  XOR U13137 ( .A(n12892), .B(n12889), .Z(n12890) );
  IV U13138 ( .A(n12842), .Z(n12838) );
  XOR U13139 ( .A(n12893), .B(n12894), .Z(n12842) );
  ANDN U13140 ( .B(n12895), .A(n12896), .Z(n12893) );
  XOR U13141 ( .A(n12897), .B(n12894), .Z(n12895) );
  IV U13142 ( .A(n12852), .Z(n12856) );
  XOR U13143 ( .A(n12852), .B(n12807), .Z(n12854) );
  XOR U13144 ( .A(n12898), .B(n12899), .Z(n12807) );
  AND U13145 ( .A(n302), .B(n12900), .Z(n12898) );
  XOR U13146 ( .A(n12901), .B(n12899), .Z(n12900) );
  NANDN U13147 ( .A(n12809), .B(n12811), .Z(n12852) );
  XOR U13148 ( .A(n12902), .B(n12903), .Z(n12811) );
  AND U13149 ( .A(n302), .B(n12904), .Z(n12902) );
  XOR U13150 ( .A(n12903), .B(n12905), .Z(n12904) );
  XNOR U13151 ( .A(n12906), .B(n12907), .Z(n302) );
  AND U13152 ( .A(n12908), .B(n12909), .Z(n12906) );
  XOR U13153 ( .A(n12907), .B(n12822), .Z(n12909) );
  XNOR U13154 ( .A(n12910), .B(n12911), .Z(n12822) );
  ANDN U13155 ( .B(n12912), .A(n12913), .Z(n12910) );
  XOR U13156 ( .A(n12911), .B(n12914), .Z(n12912) );
  XNOR U13157 ( .A(n12907), .B(n12824), .Z(n12908) );
  XOR U13158 ( .A(n12915), .B(n12916), .Z(n12824) );
  AND U13159 ( .A(n306), .B(n12917), .Z(n12915) );
  XOR U13160 ( .A(n12918), .B(n12916), .Z(n12917) );
  XNOR U13161 ( .A(n12919), .B(n12920), .Z(n12907) );
  AND U13162 ( .A(n12921), .B(n12922), .Z(n12919) );
  XNOR U13163 ( .A(n12920), .B(n12849), .Z(n12922) );
  XOR U13164 ( .A(n12913), .B(n12914), .Z(n12849) );
  XNOR U13165 ( .A(n12923), .B(n12924), .Z(n12914) );
  ANDN U13166 ( .B(n12925), .A(n12926), .Z(n12923) );
  XOR U13167 ( .A(n12927), .B(n12928), .Z(n12925) );
  XOR U13168 ( .A(n12929), .B(n12930), .Z(n12913) );
  XNOR U13169 ( .A(n12931), .B(n12932), .Z(n12930) );
  ANDN U13170 ( .B(n12933), .A(n12934), .Z(n12931) );
  XNOR U13171 ( .A(n12935), .B(n12936), .Z(n12933) );
  IV U13172 ( .A(n12911), .Z(n12929) );
  XOR U13173 ( .A(n12937), .B(n12938), .Z(n12911) );
  ANDN U13174 ( .B(n12939), .A(n12940), .Z(n12937) );
  XOR U13175 ( .A(n12938), .B(n12941), .Z(n12939) );
  XOR U13176 ( .A(n12920), .B(n12851), .Z(n12921) );
  XOR U13177 ( .A(n12942), .B(n12943), .Z(n12851) );
  AND U13178 ( .A(n306), .B(n12944), .Z(n12942) );
  XOR U13179 ( .A(n12945), .B(n12943), .Z(n12944) );
  XNOR U13180 ( .A(n12946), .B(n12947), .Z(n12920) );
  NAND U13181 ( .A(n12948), .B(n12949), .Z(n12947) );
  XOR U13182 ( .A(n12950), .B(n12899), .Z(n12949) );
  XOR U13183 ( .A(n12940), .B(n12941), .Z(n12899) );
  XOR U13184 ( .A(n12951), .B(n12928), .Z(n12941) );
  XOR U13185 ( .A(n12952), .B(n12953), .Z(n12928) );
  ANDN U13186 ( .B(n12954), .A(n12955), .Z(n12952) );
  XOR U13187 ( .A(n12953), .B(n12956), .Z(n12954) );
  IV U13188 ( .A(n12926), .Z(n12951) );
  XOR U13189 ( .A(n12924), .B(n12957), .Z(n12926) );
  XOR U13190 ( .A(n12958), .B(n12959), .Z(n12957) );
  ANDN U13191 ( .B(n12960), .A(n12961), .Z(n12958) );
  XOR U13192 ( .A(n12962), .B(n12959), .Z(n12960) );
  IV U13193 ( .A(n12927), .Z(n12924) );
  XOR U13194 ( .A(n12963), .B(n12964), .Z(n12927) );
  ANDN U13195 ( .B(n12965), .A(n12966), .Z(n12963) );
  XOR U13196 ( .A(n12964), .B(n12967), .Z(n12965) );
  XOR U13197 ( .A(n12968), .B(n12969), .Z(n12940) );
  XNOR U13198 ( .A(n12935), .B(n12970), .Z(n12969) );
  IV U13199 ( .A(n12938), .Z(n12970) );
  XOR U13200 ( .A(n12971), .B(n12972), .Z(n12938) );
  ANDN U13201 ( .B(n12973), .A(n12974), .Z(n12971) );
  XOR U13202 ( .A(n12972), .B(n12975), .Z(n12973) );
  XNOR U13203 ( .A(n12976), .B(n12977), .Z(n12935) );
  ANDN U13204 ( .B(n12978), .A(n12979), .Z(n12976) );
  XOR U13205 ( .A(n12977), .B(n12980), .Z(n12978) );
  IV U13206 ( .A(n12934), .Z(n12968) );
  XOR U13207 ( .A(n12932), .B(n12981), .Z(n12934) );
  XOR U13208 ( .A(n12982), .B(n12983), .Z(n12981) );
  ANDN U13209 ( .B(n12984), .A(n12985), .Z(n12982) );
  XOR U13210 ( .A(n12986), .B(n12983), .Z(n12984) );
  IV U13211 ( .A(n12936), .Z(n12932) );
  XOR U13212 ( .A(n12987), .B(n12988), .Z(n12936) );
  ANDN U13213 ( .B(n12989), .A(n12990), .Z(n12987) );
  XOR U13214 ( .A(n12991), .B(n12988), .Z(n12989) );
  IV U13215 ( .A(n12946), .Z(n12950) );
  XOR U13216 ( .A(n12946), .B(n12901), .Z(n12948) );
  XOR U13217 ( .A(n12992), .B(n12993), .Z(n12901) );
  AND U13218 ( .A(n306), .B(n12994), .Z(n12992) );
  XOR U13219 ( .A(n12995), .B(n12993), .Z(n12994) );
  NANDN U13220 ( .A(n12903), .B(n12905), .Z(n12946) );
  XOR U13221 ( .A(n12996), .B(n12997), .Z(n12905) );
  AND U13222 ( .A(n306), .B(n12998), .Z(n12996) );
  XOR U13223 ( .A(n12997), .B(n12999), .Z(n12998) );
  XNOR U13224 ( .A(n13000), .B(n13001), .Z(n306) );
  AND U13225 ( .A(n13002), .B(n13003), .Z(n13000) );
  XOR U13226 ( .A(n13001), .B(n12916), .Z(n13003) );
  XNOR U13227 ( .A(n13004), .B(n13005), .Z(n12916) );
  ANDN U13228 ( .B(n13006), .A(n13007), .Z(n13004) );
  XOR U13229 ( .A(n13005), .B(n13008), .Z(n13006) );
  XNOR U13230 ( .A(n13001), .B(n12918), .Z(n13002) );
  XOR U13231 ( .A(n13009), .B(n13010), .Z(n12918) );
  AND U13232 ( .A(n310), .B(n13011), .Z(n13009) );
  XOR U13233 ( .A(n13012), .B(n13010), .Z(n13011) );
  XNOR U13234 ( .A(n13013), .B(n13014), .Z(n13001) );
  AND U13235 ( .A(n13015), .B(n13016), .Z(n13013) );
  XNOR U13236 ( .A(n13014), .B(n12943), .Z(n13016) );
  XOR U13237 ( .A(n13007), .B(n13008), .Z(n12943) );
  XNOR U13238 ( .A(n13017), .B(n13018), .Z(n13008) );
  ANDN U13239 ( .B(n13019), .A(n13020), .Z(n13017) );
  XOR U13240 ( .A(n13021), .B(n13022), .Z(n13019) );
  XOR U13241 ( .A(n13023), .B(n13024), .Z(n13007) );
  XNOR U13242 ( .A(n13025), .B(n13026), .Z(n13024) );
  ANDN U13243 ( .B(n13027), .A(n13028), .Z(n13025) );
  XNOR U13244 ( .A(n13029), .B(n13030), .Z(n13027) );
  IV U13245 ( .A(n13005), .Z(n13023) );
  XOR U13246 ( .A(n13031), .B(n13032), .Z(n13005) );
  ANDN U13247 ( .B(n13033), .A(n13034), .Z(n13031) );
  XOR U13248 ( .A(n13032), .B(n13035), .Z(n13033) );
  XOR U13249 ( .A(n13014), .B(n12945), .Z(n13015) );
  XOR U13250 ( .A(n13036), .B(n13037), .Z(n12945) );
  AND U13251 ( .A(n310), .B(n13038), .Z(n13036) );
  XOR U13252 ( .A(n13039), .B(n13037), .Z(n13038) );
  XNOR U13253 ( .A(n13040), .B(n13041), .Z(n13014) );
  NAND U13254 ( .A(n13042), .B(n13043), .Z(n13041) );
  XOR U13255 ( .A(n13044), .B(n12993), .Z(n13043) );
  XOR U13256 ( .A(n13034), .B(n13035), .Z(n12993) );
  XOR U13257 ( .A(n13045), .B(n13022), .Z(n13035) );
  XOR U13258 ( .A(n13046), .B(n13047), .Z(n13022) );
  ANDN U13259 ( .B(n13048), .A(n13049), .Z(n13046) );
  XOR U13260 ( .A(n13047), .B(n13050), .Z(n13048) );
  IV U13261 ( .A(n13020), .Z(n13045) );
  XOR U13262 ( .A(n13018), .B(n13051), .Z(n13020) );
  XOR U13263 ( .A(n13052), .B(n13053), .Z(n13051) );
  ANDN U13264 ( .B(n13054), .A(n13055), .Z(n13052) );
  XOR U13265 ( .A(n13056), .B(n13053), .Z(n13054) );
  IV U13266 ( .A(n13021), .Z(n13018) );
  XOR U13267 ( .A(n13057), .B(n13058), .Z(n13021) );
  ANDN U13268 ( .B(n13059), .A(n13060), .Z(n13057) );
  XOR U13269 ( .A(n13058), .B(n13061), .Z(n13059) );
  XOR U13270 ( .A(n13062), .B(n13063), .Z(n13034) );
  XNOR U13271 ( .A(n13029), .B(n13064), .Z(n13063) );
  IV U13272 ( .A(n13032), .Z(n13064) );
  XOR U13273 ( .A(n13065), .B(n13066), .Z(n13032) );
  ANDN U13274 ( .B(n13067), .A(n13068), .Z(n13065) );
  XOR U13275 ( .A(n13066), .B(n13069), .Z(n13067) );
  XNOR U13276 ( .A(n13070), .B(n13071), .Z(n13029) );
  ANDN U13277 ( .B(n13072), .A(n13073), .Z(n13070) );
  XOR U13278 ( .A(n13071), .B(n13074), .Z(n13072) );
  IV U13279 ( .A(n13028), .Z(n13062) );
  XOR U13280 ( .A(n13026), .B(n13075), .Z(n13028) );
  XOR U13281 ( .A(n13076), .B(n13077), .Z(n13075) );
  ANDN U13282 ( .B(n13078), .A(n13079), .Z(n13076) );
  XOR U13283 ( .A(n13080), .B(n13077), .Z(n13078) );
  IV U13284 ( .A(n13030), .Z(n13026) );
  XOR U13285 ( .A(n13081), .B(n13082), .Z(n13030) );
  ANDN U13286 ( .B(n13083), .A(n13084), .Z(n13081) );
  XOR U13287 ( .A(n13085), .B(n13082), .Z(n13083) );
  IV U13288 ( .A(n13040), .Z(n13044) );
  XOR U13289 ( .A(n13040), .B(n12995), .Z(n13042) );
  XOR U13290 ( .A(n13086), .B(n13087), .Z(n12995) );
  AND U13291 ( .A(n310), .B(n13088), .Z(n13086) );
  XOR U13292 ( .A(n13089), .B(n13087), .Z(n13088) );
  NANDN U13293 ( .A(n12997), .B(n12999), .Z(n13040) );
  XOR U13294 ( .A(n13090), .B(n13091), .Z(n12999) );
  AND U13295 ( .A(n310), .B(n13092), .Z(n13090) );
  XOR U13296 ( .A(n13091), .B(n13093), .Z(n13092) );
  XNOR U13297 ( .A(n13094), .B(n13095), .Z(n310) );
  AND U13298 ( .A(n13096), .B(n13097), .Z(n13094) );
  XOR U13299 ( .A(n13095), .B(n13010), .Z(n13097) );
  XNOR U13300 ( .A(n13098), .B(n13099), .Z(n13010) );
  ANDN U13301 ( .B(n13100), .A(n13101), .Z(n13098) );
  XOR U13302 ( .A(n13099), .B(n13102), .Z(n13100) );
  XNOR U13303 ( .A(n13095), .B(n13012), .Z(n13096) );
  XOR U13304 ( .A(n13103), .B(n13104), .Z(n13012) );
  AND U13305 ( .A(n314), .B(n13105), .Z(n13103) );
  XOR U13306 ( .A(n13106), .B(n13104), .Z(n13105) );
  XNOR U13307 ( .A(n13107), .B(n13108), .Z(n13095) );
  AND U13308 ( .A(n13109), .B(n13110), .Z(n13107) );
  XNOR U13309 ( .A(n13108), .B(n13037), .Z(n13110) );
  XOR U13310 ( .A(n13101), .B(n13102), .Z(n13037) );
  XNOR U13311 ( .A(n13111), .B(n13112), .Z(n13102) );
  ANDN U13312 ( .B(n13113), .A(n13114), .Z(n13111) );
  XOR U13313 ( .A(n13115), .B(n13116), .Z(n13113) );
  XOR U13314 ( .A(n13117), .B(n13118), .Z(n13101) );
  XNOR U13315 ( .A(n13119), .B(n13120), .Z(n13118) );
  ANDN U13316 ( .B(n13121), .A(n13122), .Z(n13119) );
  XNOR U13317 ( .A(n13123), .B(n13124), .Z(n13121) );
  IV U13318 ( .A(n13099), .Z(n13117) );
  XOR U13319 ( .A(n13125), .B(n13126), .Z(n13099) );
  ANDN U13320 ( .B(n13127), .A(n13128), .Z(n13125) );
  XOR U13321 ( .A(n13126), .B(n13129), .Z(n13127) );
  XOR U13322 ( .A(n13108), .B(n13039), .Z(n13109) );
  XOR U13323 ( .A(n13130), .B(n13131), .Z(n13039) );
  AND U13324 ( .A(n314), .B(n13132), .Z(n13130) );
  XOR U13325 ( .A(n13133), .B(n13131), .Z(n13132) );
  XNOR U13326 ( .A(n13134), .B(n13135), .Z(n13108) );
  NAND U13327 ( .A(n13136), .B(n13137), .Z(n13135) );
  XOR U13328 ( .A(n13138), .B(n13087), .Z(n13137) );
  XOR U13329 ( .A(n13128), .B(n13129), .Z(n13087) );
  XOR U13330 ( .A(n13139), .B(n13116), .Z(n13129) );
  XOR U13331 ( .A(n13140), .B(n13141), .Z(n13116) );
  ANDN U13332 ( .B(n13142), .A(n13143), .Z(n13140) );
  XOR U13333 ( .A(n13141), .B(n13144), .Z(n13142) );
  IV U13334 ( .A(n13114), .Z(n13139) );
  XOR U13335 ( .A(n13112), .B(n13145), .Z(n13114) );
  XOR U13336 ( .A(n13146), .B(n13147), .Z(n13145) );
  ANDN U13337 ( .B(n13148), .A(n13149), .Z(n13146) );
  XOR U13338 ( .A(n13150), .B(n13147), .Z(n13148) );
  IV U13339 ( .A(n13115), .Z(n13112) );
  XOR U13340 ( .A(n13151), .B(n13152), .Z(n13115) );
  ANDN U13341 ( .B(n13153), .A(n13154), .Z(n13151) );
  XOR U13342 ( .A(n13152), .B(n13155), .Z(n13153) );
  XOR U13343 ( .A(n13156), .B(n13157), .Z(n13128) );
  XNOR U13344 ( .A(n13123), .B(n13158), .Z(n13157) );
  IV U13345 ( .A(n13126), .Z(n13158) );
  XOR U13346 ( .A(n13159), .B(n13160), .Z(n13126) );
  ANDN U13347 ( .B(n13161), .A(n13162), .Z(n13159) );
  XOR U13348 ( .A(n13160), .B(n13163), .Z(n13161) );
  XNOR U13349 ( .A(n13164), .B(n13165), .Z(n13123) );
  ANDN U13350 ( .B(n13166), .A(n13167), .Z(n13164) );
  XOR U13351 ( .A(n13165), .B(n13168), .Z(n13166) );
  IV U13352 ( .A(n13122), .Z(n13156) );
  XOR U13353 ( .A(n13120), .B(n13169), .Z(n13122) );
  XOR U13354 ( .A(n13170), .B(n13171), .Z(n13169) );
  ANDN U13355 ( .B(n13172), .A(n13173), .Z(n13170) );
  XOR U13356 ( .A(n13174), .B(n13171), .Z(n13172) );
  IV U13357 ( .A(n13124), .Z(n13120) );
  XOR U13358 ( .A(n13175), .B(n13176), .Z(n13124) );
  ANDN U13359 ( .B(n13177), .A(n13178), .Z(n13175) );
  XOR U13360 ( .A(n13179), .B(n13176), .Z(n13177) );
  IV U13361 ( .A(n13134), .Z(n13138) );
  XOR U13362 ( .A(n13134), .B(n13089), .Z(n13136) );
  XOR U13363 ( .A(n13180), .B(n13181), .Z(n13089) );
  AND U13364 ( .A(n314), .B(n13182), .Z(n13180) );
  XOR U13365 ( .A(n13183), .B(n13181), .Z(n13182) );
  NANDN U13366 ( .A(n13091), .B(n13093), .Z(n13134) );
  XOR U13367 ( .A(n13184), .B(n13185), .Z(n13093) );
  AND U13368 ( .A(n314), .B(n13186), .Z(n13184) );
  XOR U13369 ( .A(n13185), .B(n13187), .Z(n13186) );
  XNOR U13370 ( .A(n13188), .B(n13189), .Z(n314) );
  AND U13371 ( .A(n13190), .B(n13191), .Z(n13188) );
  XOR U13372 ( .A(n13189), .B(n13104), .Z(n13191) );
  XNOR U13373 ( .A(n13192), .B(n13193), .Z(n13104) );
  ANDN U13374 ( .B(n13194), .A(n13195), .Z(n13192) );
  XOR U13375 ( .A(n13193), .B(n13196), .Z(n13194) );
  XNOR U13376 ( .A(n13189), .B(n13106), .Z(n13190) );
  XOR U13377 ( .A(n13197), .B(n13198), .Z(n13106) );
  AND U13378 ( .A(n318), .B(n13199), .Z(n13197) );
  XOR U13379 ( .A(n13200), .B(n13198), .Z(n13199) );
  XNOR U13380 ( .A(n13201), .B(n13202), .Z(n13189) );
  AND U13381 ( .A(n13203), .B(n13204), .Z(n13201) );
  XNOR U13382 ( .A(n13202), .B(n13131), .Z(n13204) );
  XOR U13383 ( .A(n13195), .B(n13196), .Z(n13131) );
  XNOR U13384 ( .A(n13205), .B(n13206), .Z(n13196) );
  ANDN U13385 ( .B(n13207), .A(n13208), .Z(n13205) );
  XOR U13386 ( .A(n13209), .B(n13210), .Z(n13207) );
  XOR U13387 ( .A(n13211), .B(n13212), .Z(n13195) );
  XNOR U13388 ( .A(n13213), .B(n13214), .Z(n13212) );
  ANDN U13389 ( .B(n13215), .A(n13216), .Z(n13213) );
  XNOR U13390 ( .A(n13217), .B(n13218), .Z(n13215) );
  IV U13391 ( .A(n13193), .Z(n13211) );
  XOR U13392 ( .A(n13219), .B(n13220), .Z(n13193) );
  ANDN U13393 ( .B(n13221), .A(n13222), .Z(n13219) );
  XOR U13394 ( .A(n13220), .B(n13223), .Z(n13221) );
  XOR U13395 ( .A(n13202), .B(n13133), .Z(n13203) );
  XOR U13396 ( .A(n13224), .B(n13225), .Z(n13133) );
  AND U13397 ( .A(n318), .B(n13226), .Z(n13224) );
  XOR U13398 ( .A(n13227), .B(n13225), .Z(n13226) );
  XNOR U13399 ( .A(n13228), .B(n13229), .Z(n13202) );
  NAND U13400 ( .A(n13230), .B(n13231), .Z(n13229) );
  XOR U13401 ( .A(n13232), .B(n13181), .Z(n13231) );
  XOR U13402 ( .A(n13222), .B(n13223), .Z(n13181) );
  XOR U13403 ( .A(n13233), .B(n13210), .Z(n13223) );
  XOR U13404 ( .A(n13234), .B(n13235), .Z(n13210) );
  ANDN U13405 ( .B(n13236), .A(n13237), .Z(n13234) );
  XOR U13406 ( .A(n13235), .B(n13238), .Z(n13236) );
  IV U13407 ( .A(n13208), .Z(n13233) );
  XOR U13408 ( .A(n13206), .B(n13239), .Z(n13208) );
  XOR U13409 ( .A(n13240), .B(n13241), .Z(n13239) );
  ANDN U13410 ( .B(n13242), .A(n13243), .Z(n13240) );
  XOR U13411 ( .A(n13244), .B(n13241), .Z(n13242) );
  IV U13412 ( .A(n13209), .Z(n13206) );
  XOR U13413 ( .A(n13245), .B(n13246), .Z(n13209) );
  ANDN U13414 ( .B(n13247), .A(n13248), .Z(n13245) );
  XOR U13415 ( .A(n13246), .B(n13249), .Z(n13247) );
  XOR U13416 ( .A(n13250), .B(n13251), .Z(n13222) );
  XNOR U13417 ( .A(n13217), .B(n13252), .Z(n13251) );
  IV U13418 ( .A(n13220), .Z(n13252) );
  XOR U13419 ( .A(n13253), .B(n13254), .Z(n13220) );
  ANDN U13420 ( .B(n13255), .A(n13256), .Z(n13253) );
  XOR U13421 ( .A(n13254), .B(n13257), .Z(n13255) );
  XNOR U13422 ( .A(n13258), .B(n13259), .Z(n13217) );
  ANDN U13423 ( .B(n13260), .A(n13261), .Z(n13258) );
  XOR U13424 ( .A(n13259), .B(n13262), .Z(n13260) );
  IV U13425 ( .A(n13216), .Z(n13250) );
  XOR U13426 ( .A(n13214), .B(n13263), .Z(n13216) );
  XOR U13427 ( .A(n13264), .B(n13265), .Z(n13263) );
  ANDN U13428 ( .B(n13266), .A(n13267), .Z(n13264) );
  XOR U13429 ( .A(n13268), .B(n13265), .Z(n13266) );
  IV U13430 ( .A(n13218), .Z(n13214) );
  XOR U13431 ( .A(n13269), .B(n13270), .Z(n13218) );
  ANDN U13432 ( .B(n13271), .A(n13272), .Z(n13269) );
  XOR U13433 ( .A(n13273), .B(n13270), .Z(n13271) );
  IV U13434 ( .A(n13228), .Z(n13232) );
  XOR U13435 ( .A(n13228), .B(n13183), .Z(n13230) );
  XOR U13436 ( .A(n13274), .B(n13275), .Z(n13183) );
  AND U13437 ( .A(n318), .B(n13276), .Z(n13274) );
  XOR U13438 ( .A(n13277), .B(n13275), .Z(n13276) );
  NANDN U13439 ( .A(n13185), .B(n13187), .Z(n13228) );
  XOR U13440 ( .A(n13278), .B(n13279), .Z(n13187) );
  AND U13441 ( .A(n318), .B(n13280), .Z(n13278) );
  XOR U13442 ( .A(n13279), .B(n13281), .Z(n13280) );
  XNOR U13443 ( .A(n13282), .B(n13283), .Z(n318) );
  AND U13444 ( .A(n13284), .B(n13285), .Z(n13282) );
  XOR U13445 ( .A(n13283), .B(n13198), .Z(n13285) );
  XNOR U13446 ( .A(n13286), .B(n13287), .Z(n13198) );
  ANDN U13447 ( .B(n13288), .A(n13289), .Z(n13286) );
  XOR U13448 ( .A(n13287), .B(n13290), .Z(n13288) );
  XNOR U13449 ( .A(n13283), .B(n13200), .Z(n13284) );
  XOR U13450 ( .A(n13291), .B(n13292), .Z(n13200) );
  AND U13451 ( .A(n322), .B(n13293), .Z(n13291) );
  XOR U13452 ( .A(n13294), .B(n13292), .Z(n13293) );
  XNOR U13453 ( .A(n13295), .B(n13296), .Z(n13283) );
  AND U13454 ( .A(n13297), .B(n13298), .Z(n13295) );
  XNOR U13455 ( .A(n13296), .B(n13225), .Z(n13298) );
  XOR U13456 ( .A(n13289), .B(n13290), .Z(n13225) );
  XNOR U13457 ( .A(n13299), .B(n13300), .Z(n13290) );
  ANDN U13458 ( .B(n13301), .A(n13302), .Z(n13299) );
  XOR U13459 ( .A(n13303), .B(n13304), .Z(n13301) );
  XOR U13460 ( .A(n13305), .B(n13306), .Z(n13289) );
  XNOR U13461 ( .A(n13307), .B(n13308), .Z(n13306) );
  ANDN U13462 ( .B(n13309), .A(n13310), .Z(n13307) );
  XNOR U13463 ( .A(n13311), .B(n13312), .Z(n13309) );
  IV U13464 ( .A(n13287), .Z(n13305) );
  XOR U13465 ( .A(n13313), .B(n13314), .Z(n13287) );
  ANDN U13466 ( .B(n13315), .A(n13316), .Z(n13313) );
  XOR U13467 ( .A(n13314), .B(n13317), .Z(n13315) );
  XOR U13468 ( .A(n13296), .B(n13227), .Z(n13297) );
  XOR U13469 ( .A(n13318), .B(n13319), .Z(n13227) );
  AND U13470 ( .A(n322), .B(n13320), .Z(n13318) );
  XOR U13471 ( .A(n13321), .B(n13319), .Z(n13320) );
  XNOR U13472 ( .A(n13322), .B(n13323), .Z(n13296) );
  NAND U13473 ( .A(n13324), .B(n13325), .Z(n13323) );
  XOR U13474 ( .A(n13326), .B(n13275), .Z(n13325) );
  XOR U13475 ( .A(n13316), .B(n13317), .Z(n13275) );
  XOR U13476 ( .A(n13327), .B(n13304), .Z(n13317) );
  XOR U13477 ( .A(n13328), .B(n13329), .Z(n13304) );
  ANDN U13478 ( .B(n13330), .A(n13331), .Z(n13328) );
  XOR U13479 ( .A(n13329), .B(n13332), .Z(n13330) );
  IV U13480 ( .A(n13302), .Z(n13327) );
  XOR U13481 ( .A(n13300), .B(n13333), .Z(n13302) );
  XOR U13482 ( .A(n13334), .B(n13335), .Z(n13333) );
  ANDN U13483 ( .B(n13336), .A(n13337), .Z(n13334) );
  XOR U13484 ( .A(n13338), .B(n13335), .Z(n13336) );
  IV U13485 ( .A(n13303), .Z(n13300) );
  XOR U13486 ( .A(n13339), .B(n13340), .Z(n13303) );
  ANDN U13487 ( .B(n13341), .A(n13342), .Z(n13339) );
  XOR U13488 ( .A(n13340), .B(n13343), .Z(n13341) );
  XOR U13489 ( .A(n13344), .B(n13345), .Z(n13316) );
  XNOR U13490 ( .A(n13311), .B(n13346), .Z(n13345) );
  IV U13491 ( .A(n13314), .Z(n13346) );
  XOR U13492 ( .A(n13347), .B(n13348), .Z(n13314) );
  ANDN U13493 ( .B(n13349), .A(n13350), .Z(n13347) );
  XOR U13494 ( .A(n13348), .B(n13351), .Z(n13349) );
  XNOR U13495 ( .A(n13352), .B(n13353), .Z(n13311) );
  ANDN U13496 ( .B(n13354), .A(n13355), .Z(n13352) );
  XOR U13497 ( .A(n13353), .B(n13356), .Z(n13354) );
  IV U13498 ( .A(n13310), .Z(n13344) );
  XOR U13499 ( .A(n13308), .B(n13357), .Z(n13310) );
  XOR U13500 ( .A(n13358), .B(n13359), .Z(n13357) );
  ANDN U13501 ( .B(n13360), .A(n13361), .Z(n13358) );
  XOR U13502 ( .A(n13362), .B(n13359), .Z(n13360) );
  IV U13503 ( .A(n13312), .Z(n13308) );
  XOR U13504 ( .A(n13363), .B(n13364), .Z(n13312) );
  ANDN U13505 ( .B(n13365), .A(n13366), .Z(n13363) );
  XOR U13506 ( .A(n13367), .B(n13364), .Z(n13365) );
  IV U13507 ( .A(n13322), .Z(n13326) );
  XOR U13508 ( .A(n13322), .B(n13277), .Z(n13324) );
  XOR U13509 ( .A(n13368), .B(n13369), .Z(n13277) );
  AND U13510 ( .A(n322), .B(n13370), .Z(n13368) );
  XOR U13511 ( .A(n13371), .B(n13369), .Z(n13370) );
  NANDN U13512 ( .A(n13279), .B(n13281), .Z(n13322) );
  XOR U13513 ( .A(n13372), .B(n13373), .Z(n13281) );
  AND U13514 ( .A(n322), .B(n13374), .Z(n13372) );
  XOR U13515 ( .A(n13373), .B(n13375), .Z(n13374) );
  XNOR U13516 ( .A(n13376), .B(n13377), .Z(n322) );
  AND U13517 ( .A(n13378), .B(n13379), .Z(n13376) );
  XOR U13518 ( .A(n13377), .B(n13292), .Z(n13379) );
  XNOR U13519 ( .A(n13380), .B(n13381), .Z(n13292) );
  ANDN U13520 ( .B(n13382), .A(n13383), .Z(n13380) );
  XOR U13521 ( .A(n13381), .B(n13384), .Z(n13382) );
  XNOR U13522 ( .A(n13377), .B(n13294), .Z(n13378) );
  XOR U13523 ( .A(n13385), .B(n13386), .Z(n13294) );
  AND U13524 ( .A(n326), .B(n13387), .Z(n13385) );
  XOR U13525 ( .A(n13388), .B(n13386), .Z(n13387) );
  XNOR U13526 ( .A(n13389), .B(n13390), .Z(n13377) );
  AND U13527 ( .A(n13391), .B(n13392), .Z(n13389) );
  XNOR U13528 ( .A(n13390), .B(n13319), .Z(n13392) );
  XOR U13529 ( .A(n13383), .B(n13384), .Z(n13319) );
  XNOR U13530 ( .A(n13393), .B(n13394), .Z(n13384) );
  ANDN U13531 ( .B(n13395), .A(n13396), .Z(n13393) );
  XOR U13532 ( .A(n13397), .B(n13398), .Z(n13395) );
  XOR U13533 ( .A(n13399), .B(n13400), .Z(n13383) );
  XNOR U13534 ( .A(n13401), .B(n13402), .Z(n13400) );
  ANDN U13535 ( .B(n13403), .A(n13404), .Z(n13401) );
  XNOR U13536 ( .A(n13405), .B(n13406), .Z(n13403) );
  IV U13537 ( .A(n13381), .Z(n13399) );
  XOR U13538 ( .A(n13407), .B(n13408), .Z(n13381) );
  ANDN U13539 ( .B(n13409), .A(n13410), .Z(n13407) );
  XOR U13540 ( .A(n13408), .B(n13411), .Z(n13409) );
  XOR U13541 ( .A(n13390), .B(n13321), .Z(n13391) );
  XOR U13542 ( .A(n13412), .B(n13413), .Z(n13321) );
  AND U13543 ( .A(n326), .B(n13414), .Z(n13412) );
  XOR U13544 ( .A(n13415), .B(n13413), .Z(n13414) );
  XNOR U13545 ( .A(n13416), .B(n13417), .Z(n13390) );
  NAND U13546 ( .A(n13418), .B(n13419), .Z(n13417) );
  XOR U13547 ( .A(n13420), .B(n13369), .Z(n13419) );
  XOR U13548 ( .A(n13410), .B(n13411), .Z(n13369) );
  XOR U13549 ( .A(n13421), .B(n13398), .Z(n13411) );
  XOR U13550 ( .A(n13422), .B(n13423), .Z(n13398) );
  ANDN U13551 ( .B(n13424), .A(n13425), .Z(n13422) );
  XOR U13552 ( .A(n13423), .B(n13426), .Z(n13424) );
  IV U13553 ( .A(n13396), .Z(n13421) );
  XOR U13554 ( .A(n13394), .B(n13427), .Z(n13396) );
  XOR U13555 ( .A(n13428), .B(n13429), .Z(n13427) );
  ANDN U13556 ( .B(n13430), .A(n13431), .Z(n13428) );
  XOR U13557 ( .A(n13432), .B(n13429), .Z(n13430) );
  IV U13558 ( .A(n13397), .Z(n13394) );
  XOR U13559 ( .A(n13433), .B(n13434), .Z(n13397) );
  ANDN U13560 ( .B(n13435), .A(n13436), .Z(n13433) );
  XOR U13561 ( .A(n13434), .B(n13437), .Z(n13435) );
  XOR U13562 ( .A(n13438), .B(n13439), .Z(n13410) );
  XNOR U13563 ( .A(n13405), .B(n13440), .Z(n13439) );
  IV U13564 ( .A(n13408), .Z(n13440) );
  XOR U13565 ( .A(n13441), .B(n13442), .Z(n13408) );
  ANDN U13566 ( .B(n13443), .A(n13444), .Z(n13441) );
  XOR U13567 ( .A(n13442), .B(n13445), .Z(n13443) );
  XNOR U13568 ( .A(n13446), .B(n13447), .Z(n13405) );
  ANDN U13569 ( .B(n13448), .A(n13449), .Z(n13446) );
  XOR U13570 ( .A(n13447), .B(n13450), .Z(n13448) );
  IV U13571 ( .A(n13404), .Z(n13438) );
  XOR U13572 ( .A(n13402), .B(n13451), .Z(n13404) );
  XOR U13573 ( .A(n13452), .B(n13453), .Z(n13451) );
  ANDN U13574 ( .B(n13454), .A(n13455), .Z(n13452) );
  XOR U13575 ( .A(n13456), .B(n13453), .Z(n13454) );
  IV U13576 ( .A(n13406), .Z(n13402) );
  XOR U13577 ( .A(n13457), .B(n13458), .Z(n13406) );
  ANDN U13578 ( .B(n13459), .A(n13460), .Z(n13457) );
  XOR U13579 ( .A(n13461), .B(n13458), .Z(n13459) );
  IV U13580 ( .A(n13416), .Z(n13420) );
  XOR U13581 ( .A(n13416), .B(n13371), .Z(n13418) );
  XOR U13582 ( .A(n13462), .B(n13463), .Z(n13371) );
  AND U13583 ( .A(n326), .B(n13464), .Z(n13462) );
  XOR U13584 ( .A(n13465), .B(n13463), .Z(n13464) );
  NANDN U13585 ( .A(n13373), .B(n13375), .Z(n13416) );
  XOR U13586 ( .A(n13466), .B(n13467), .Z(n13375) );
  AND U13587 ( .A(n326), .B(n13468), .Z(n13466) );
  XOR U13588 ( .A(n13467), .B(n13469), .Z(n13468) );
  XNOR U13589 ( .A(n13470), .B(n13471), .Z(n326) );
  AND U13590 ( .A(n13472), .B(n13473), .Z(n13470) );
  XOR U13591 ( .A(n13471), .B(n13386), .Z(n13473) );
  XNOR U13592 ( .A(n13474), .B(n13475), .Z(n13386) );
  ANDN U13593 ( .B(n13476), .A(n13477), .Z(n13474) );
  XOR U13594 ( .A(n13475), .B(n13478), .Z(n13476) );
  XNOR U13595 ( .A(n13471), .B(n13388), .Z(n13472) );
  XOR U13596 ( .A(n13479), .B(n13480), .Z(n13388) );
  AND U13597 ( .A(n330), .B(n13481), .Z(n13479) );
  XOR U13598 ( .A(n13482), .B(n13480), .Z(n13481) );
  XNOR U13599 ( .A(n13483), .B(n13484), .Z(n13471) );
  AND U13600 ( .A(n13485), .B(n13486), .Z(n13483) );
  XNOR U13601 ( .A(n13484), .B(n13413), .Z(n13486) );
  XOR U13602 ( .A(n13477), .B(n13478), .Z(n13413) );
  XNOR U13603 ( .A(n13487), .B(n13488), .Z(n13478) );
  ANDN U13604 ( .B(n13489), .A(n13490), .Z(n13487) );
  XOR U13605 ( .A(n13491), .B(n13492), .Z(n13489) );
  XOR U13606 ( .A(n13493), .B(n13494), .Z(n13477) );
  XNOR U13607 ( .A(n13495), .B(n13496), .Z(n13494) );
  ANDN U13608 ( .B(n13497), .A(n13498), .Z(n13495) );
  XNOR U13609 ( .A(n13499), .B(n13500), .Z(n13497) );
  IV U13610 ( .A(n13475), .Z(n13493) );
  XOR U13611 ( .A(n13501), .B(n13502), .Z(n13475) );
  ANDN U13612 ( .B(n13503), .A(n13504), .Z(n13501) );
  XOR U13613 ( .A(n13502), .B(n13505), .Z(n13503) );
  XOR U13614 ( .A(n13484), .B(n13415), .Z(n13485) );
  XOR U13615 ( .A(n13506), .B(n13507), .Z(n13415) );
  AND U13616 ( .A(n330), .B(n13508), .Z(n13506) );
  XOR U13617 ( .A(n13509), .B(n13507), .Z(n13508) );
  XNOR U13618 ( .A(n13510), .B(n13511), .Z(n13484) );
  NAND U13619 ( .A(n13512), .B(n13513), .Z(n13511) );
  XOR U13620 ( .A(n13514), .B(n13463), .Z(n13513) );
  XOR U13621 ( .A(n13504), .B(n13505), .Z(n13463) );
  XOR U13622 ( .A(n13515), .B(n13492), .Z(n13505) );
  XOR U13623 ( .A(n13516), .B(n13517), .Z(n13492) );
  ANDN U13624 ( .B(n13518), .A(n13519), .Z(n13516) );
  XOR U13625 ( .A(n13517), .B(n13520), .Z(n13518) );
  IV U13626 ( .A(n13490), .Z(n13515) );
  XOR U13627 ( .A(n13488), .B(n13521), .Z(n13490) );
  XOR U13628 ( .A(n13522), .B(n13523), .Z(n13521) );
  ANDN U13629 ( .B(n13524), .A(n13525), .Z(n13522) );
  XOR U13630 ( .A(n13526), .B(n13523), .Z(n13524) );
  IV U13631 ( .A(n13491), .Z(n13488) );
  XOR U13632 ( .A(n13527), .B(n13528), .Z(n13491) );
  ANDN U13633 ( .B(n13529), .A(n13530), .Z(n13527) );
  XOR U13634 ( .A(n13528), .B(n13531), .Z(n13529) );
  XOR U13635 ( .A(n13532), .B(n13533), .Z(n13504) );
  XNOR U13636 ( .A(n13499), .B(n13534), .Z(n13533) );
  IV U13637 ( .A(n13502), .Z(n13534) );
  XOR U13638 ( .A(n13535), .B(n13536), .Z(n13502) );
  ANDN U13639 ( .B(n13537), .A(n13538), .Z(n13535) );
  XOR U13640 ( .A(n13536), .B(n13539), .Z(n13537) );
  XNOR U13641 ( .A(n13540), .B(n13541), .Z(n13499) );
  ANDN U13642 ( .B(n13542), .A(n13543), .Z(n13540) );
  XOR U13643 ( .A(n13541), .B(n13544), .Z(n13542) );
  IV U13644 ( .A(n13498), .Z(n13532) );
  XOR U13645 ( .A(n13496), .B(n13545), .Z(n13498) );
  XOR U13646 ( .A(n13546), .B(n13547), .Z(n13545) );
  ANDN U13647 ( .B(n13548), .A(n13549), .Z(n13546) );
  XOR U13648 ( .A(n13550), .B(n13547), .Z(n13548) );
  IV U13649 ( .A(n13500), .Z(n13496) );
  XOR U13650 ( .A(n13551), .B(n13552), .Z(n13500) );
  ANDN U13651 ( .B(n13553), .A(n13554), .Z(n13551) );
  XOR U13652 ( .A(n13555), .B(n13552), .Z(n13553) );
  IV U13653 ( .A(n13510), .Z(n13514) );
  XOR U13654 ( .A(n13510), .B(n13465), .Z(n13512) );
  XOR U13655 ( .A(n13556), .B(n13557), .Z(n13465) );
  AND U13656 ( .A(n330), .B(n13558), .Z(n13556) );
  XOR U13657 ( .A(n13559), .B(n13557), .Z(n13558) );
  NANDN U13658 ( .A(n13467), .B(n13469), .Z(n13510) );
  XOR U13659 ( .A(n13560), .B(n13561), .Z(n13469) );
  AND U13660 ( .A(n330), .B(n13562), .Z(n13560) );
  XOR U13661 ( .A(n13561), .B(n13563), .Z(n13562) );
  XNOR U13662 ( .A(n13564), .B(n13565), .Z(n330) );
  AND U13663 ( .A(n13566), .B(n13567), .Z(n13564) );
  XOR U13664 ( .A(n13565), .B(n13480), .Z(n13567) );
  XNOR U13665 ( .A(n13568), .B(n13569), .Z(n13480) );
  ANDN U13666 ( .B(n13570), .A(n13571), .Z(n13568) );
  XOR U13667 ( .A(n13569), .B(n13572), .Z(n13570) );
  XNOR U13668 ( .A(n13565), .B(n13482), .Z(n13566) );
  XOR U13669 ( .A(n13573), .B(n13574), .Z(n13482) );
  AND U13670 ( .A(n334), .B(n13575), .Z(n13573) );
  XOR U13671 ( .A(n13576), .B(n13574), .Z(n13575) );
  XNOR U13672 ( .A(n13577), .B(n13578), .Z(n13565) );
  AND U13673 ( .A(n13579), .B(n13580), .Z(n13577) );
  XNOR U13674 ( .A(n13578), .B(n13507), .Z(n13580) );
  XOR U13675 ( .A(n13571), .B(n13572), .Z(n13507) );
  XNOR U13676 ( .A(n13581), .B(n13582), .Z(n13572) );
  ANDN U13677 ( .B(n13583), .A(n13584), .Z(n13581) );
  XOR U13678 ( .A(n13585), .B(n13586), .Z(n13583) );
  XOR U13679 ( .A(n13587), .B(n13588), .Z(n13571) );
  XNOR U13680 ( .A(n13589), .B(n13590), .Z(n13588) );
  ANDN U13681 ( .B(n13591), .A(n13592), .Z(n13589) );
  XNOR U13682 ( .A(n13593), .B(n13594), .Z(n13591) );
  IV U13683 ( .A(n13569), .Z(n13587) );
  XOR U13684 ( .A(n13595), .B(n13596), .Z(n13569) );
  ANDN U13685 ( .B(n13597), .A(n13598), .Z(n13595) );
  XOR U13686 ( .A(n13596), .B(n13599), .Z(n13597) );
  XOR U13687 ( .A(n13578), .B(n13509), .Z(n13579) );
  XOR U13688 ( .A(n13600), .B(n13601), .Z(n13509) );
  AND U13689 ( .A(n334), .B(n13602), .Z(n13600) );
  XOR U13690 ( .A(n13603), .B(n13601), .Z(n13602) );
  XNOR U13691 ( .A(n13604), .B(n13605), .Z(n13578) );
  NAND U13692 ( .A(n13606), .B(n13607), .Z(n13605) );
  XOR U13693 ( .A(n13608), .B(n13557), .Z(n13607) );
  XOR U13694 ( .A(n13598), .B(n13599), .Z(n13557) );
  XOR U13695 ( .A(n13609), .B(n13586), .Z(n13599) );
  XOR U13696 ( .A(n13610), .B(n13611), .Z(n13586) );
  ANDN U13697 ( .B(n13612), .A(n13613), .Z(n13610) );
  XOR U13698 ( .A(n13611), .B(n13614), .Z(n13612) );
  IV U13699 ( .A(n13584), .Z(n13609) );
  XOR U13700 ( .A(n13582), .B(n13615), .Z(n13584) );
  XOR U13701 ( .A(n13616), .B(n13617), .Z(n13615) );
  ANDN U13702 ( .B(n13618), .A(n13619), .Z(n13616) );
  XOR U13703 ( .A(n13620), .B(n13617), .Z(n13618) );
  IV U13704 ( .A(n13585), .Z(n13582) );
  XOR U13705 ( .A(n13621), .B(n13622), .Z(n13585) );
  ANDN U13706 ( .B(n13623), .A(n13624), .Z(n13621) );
  XOR U13707 ( .A(n13622), .B(n13625), .Z(n13623) );
  XOR U13708 ( .A(n13626), .B(n13627), .Z(n13598) );
  XNOR U13709 ( .A(n13593), .B(n13628), .Z(n13627) );
  IV U13710 ( .A(n13596), .Z(n13628) );
  XOR U13711 ( .A(n13629), .B(n13630), .Z(n13596) );
  ANDN U13712 ( .B(n13631), .A(n13632), .Z(n13629) );
  XOR U13713 ( .A(n13630), .B(n13633), .Z(n13631) );
  XNOR U13714 ( .A(n13634), .B(n13635), .Z(n13593) );
  ANDN U13715 ( .B(n13636), .A(n13637), .Z(n13634) );
  XOR U13716 ( .A(n13635), .B(n13638), .Z(n13636) );
  IV U13717 ( .A(n13592), .Z(n13626) );
  XOR U13718 ( .A(n13590), .B(n13639), .Z(n13592) );
  XOR U13719 ( .A(n13640), .B(n13641), .Z(n13639) );
  ANDN U13720 ( .B(n13642), .A(n13643), .Z(n13640) );
  XOR U13721 ( .A(n13644), .B(n13641), .Z(n13642) );
  IV U13722 ( .A(n13594), .Z(n13590) );
  XOR U13723 ( .A(n13645), .B(n13646), .Z(n13594) );
  ANDN U13724 ( .B(n13647), .A(n13648), .Z(n13645) );
  XOR U13725 ( .A(n13649), .B(n13646), .Z(n13647) );
  IV U13726 ( .A(n13604), .Z(n13608) );
  XOR U13727 ( .A(n13604), .B(n13559), .Z(n13606) );
  XOR U13728 ( .A(n13650), .B(n13651), .Z(n13559) );
  AND U13729 ( .A(n334), .B(n13652), .Z(n13650) );
  XOR U13730 ( .A(n13653), .B(n13651), .Z(n13652) );
  NANDN U13731 ( .A(n13561), .B(n13563), .Z(n13604) );
  XOR U13732 ( .A(n13654), .B(n13655), .Z(n13563) );
  AND U13733 ( .A(n334), .B(n13656), .Z(n13654) );
  XOR U13734 ( .A(n13655), .B(n13657), .Z(n13656) );
  XNOR U13735 ( .A(n13658), .B(n13659), .Z(n334) );
  AND U13736 ( .A(n13660), .B(n13661), .Z(n13658) );
  XOR U13737 ( .A(n13659), .B(n13574), .Z(n13661) );
  XNOR U13738 ( .A(n13662), .B(n13663), .Z(n13574) );
  ANDN U13739 ( .B(n13664), .A(n13665), .Z(n13662) );
  XOR U13740 ( .A(n13663), .B(n13666), .Z(n13664) );
  XNOR U13741 ( .A(n13659), .B(n13576), .Z(n13660) );
  XOR U13742 ( .A(n13667), .B(n13668), .Z(n13576) );
  AND U13743 ( .A(n338), .B(n13669), .Z(n13667) );
  XOR U13744 ( .A(n13670), .B(n13668), .Z(n13669) );
  XNOR U13745 ( .A(n13671), .B(n13672), .Z(n13659) );
  AND U13746 ( .A(n13673), .B(n13674), .Z(n13671) );
  XNOR U13747 ( .A(n13672), .B(n13601), .Z(n13674) );
  XOR U13748 ( .A(n13665), .B(n13666), .Z(n13601) );
  XNOR U13749 ( .A(n13675), .B(n13676), .Z(n13666) );
  ANDN U13750 ( .B(n13677), .A(n13678), .Z(n13675) );
  XOR U13751 ( .A(n13679), .B(n13680), .Z(n13677) );
  XOR U13752 ( .A(n13681), .B(n13682), .Z(n13665) );
  XNOR U13753 ( .A(n13683), .B(n13684), .Z(n13682) );
  ANDN U13754 ( .B(n13685), .A(n13686), .Z(n13683) );
  XNOR U13755 ( .A(n13687), .B(n13688), .Z(n13685) );
  IV U13756 ( .A(n13663), .Z(n13681) );
  XOR U13757 ( .A(n13689), .B(n13690), .Z(n13663) );
  ANDN U13758 ( .B(n13691), .A(n13692), .Z(n13689) );
  XOR U13759 ( .A(n13690), .B(n13693), .Z(n13691) );
  XOR U13760 ( .A(n13672), .B(n13603), .Z(n13673) );
  XOR U13761 ( .A(n13694), .B(n13695), .Z(n13603) );
  AND U13762 ( .A(n338), .B(n13696), .Z(n13694) );
  XOR U13763 ( .A(n13697), .B(n13695), .Z(n13696) );
  XNOR U13764 ( .A(n13698), .B(n13699), .Z(n13672) );
  NAND U13765 ( .A(n13700), .B(n13701), .Z(n13699) );
  XOR U13766 ( .A(n13702), .B(n13651), .Z(n13701) );
  XOR U13767 ( .A(n13692), .B(n13693), .Z(n13651) );
  XOR U13768 ( .A(n13703), .B(n13680), .Z(n13693) );
  XOR U13769 ( .A(n13704), .B(n13705), .Z(n13680) );
  ANDN U13770 ( .B(n13706), .A(n13707), .Z(n13704) );
  XOR U13771 ( .A(n13705), .B(n13708), .Z(n13706) );
  IV U13772 ( .A(n13678), .Z(n13703) );
  XOR U13773 ( .A(n13676), .B(n13709), .Z(n13678) );
  XOR U13774 ( .A(n13710), .B(n13711), .Z(n13709) );
  ANDN U13775 ( .B(n13712), .A(n13713), .Z(n13710) );
  XOR U13776 ( .A(n13714), .B(n13711), .Z(n13712) );
  IV U13777 ( .A(n13679), .Z(n13676) );
  XOR U13778 ( .A(n13715), .B(n13716), .Z(n13679) );
  ANDN U13779 ( .B(n13717), .A(n13718), .Z(n13715) );
  XOR U13780 ( .A(n13716), .B(n13719), .Z(n13717) );
  XOR U13781 ( .A(n13720), .B(n13721), .Z(n13692) );
  XNOR U13782 ( .A(n13687), .B(n13722), .Z(n13721) );
  IV U13783 ( .A(n13690), .Z(n13722) );
  XOR U13784 ( .A(n13723), .B(n13724), .Z(n13690) );
  ANDN U13785 ( .B(n13725), .A(n13726), .Z(n13723) );
  XOR U13786 ( .A(n13724), .B(n13727), .Z(n13725) );
  XNOR U13787 ( .A(n13728), .B(n13729), .Z(n13687) );
  ANDN U13788 ( .B(n13730), .A(n13731), .Z(n13728) );
  XOR U13789 ( .A(n13729), .B(n13732), .Z(n13730) );
  IV U13790 ( .A(n13686), .Z(n13720) );
  XOR U13791 ( .A(n13684), .B(n13733), .Z(n13686) );
  XOR U13792 ( .A(n13734), .B(n13735), .Z(n13733) );
  ANDN U13793 ( .B(n13736), .A(n13737), .Z(n13734) );
  XOR U13794 ( .A(n13738), .B(n13735), .Z(n13736) );
  IV U13795 ( .A(n13688), .Z(n13684) );
  XOR U13796 ( .A(n13739), .B(n13740), .Z(n13688) );
  ANDN U13797 ( .B(n13741), .A(n13742), .Z(n13739) );
  XOR U13798 ( .A(n13743), .B(n13740), .Z(n13741) );
  IV U13799 ( .A(n13698), .Z(n13702) );
  XOR U13800 ( .A(n13698), .B(n13653), .Z(n13700) );
  XOR U13801 ( .A(n13744), .B(n13745), .Z(n13653) );
  AND U13802 ( .A(n338), .B(n13746), .Z(n13744) );
  XOR U13803 ( .A(n13747), .B(n13745), .Z(n13746) );
  NANDN U13804 ( .A(n13655), .B(n13657), .Z(n13698) );
  XOR U13805 ( .A(n13748), .B(n13749), .Z(n13657) );
  AND U13806 ( .A(n338), .B(n13750), .Z(n13748) );
  XOR U13807 ( .A(n13749), .B(n13751), .Z(n13750) );
  XNOR U13808 ( .A(n13752), .B(n13753), .Z(n338) );
  AND U13809 ( .A(n13754), .B(n13755), .Z(n13752) );
  XOR U13810 ( .A(n13753), .B(n13668), .Z(n13755) );
  XNOR U13811 ( .A(n13756), .B(n13757), .Z(n13668) );
  ANDN U13812 ( .B(n13758), .A(n13759), .Z(n13756) );
  XOR U13813 ( .A(n13757), .B(n13760), .Z(n13758) );
  XNOR U13814 ( .A(n13753), .B(n13670), .Z(n13754) );
  XOR U13815 ( .A(n13761), .B(n13762), .Z(n13670) );
  AND U13816 ( .A(n342), .B(n13763), .Z(n13761) );
  XOR U13817 ( .A(n13764), .B(n13762), .Z(n13763) );
  XNOR U13818 ( .A(n13765), .B(n13766), .Z(n13753) );
  AND U13819 ( .A(n13767), .B(n13768), .Z(n13765) );
  XNOR U13820 ( .A(n13766), .B(n13695), .Z(n13768) );
  XOR U13821 ( .A(n13759), .B(n13760), .Z(n13695) );
  XNOR U13822 ( .A(n13769), .B(n13770), .Z(n13760) );
  ANDN U13823 ( .B(n13771), .A(n13772), .Z(n13769) );
  XOR U13824 ( .A(n13773), .B(n13774), .Z(n13771) );
  XOR U13825 ( .A(n13775), .B(n13776), .Z(n13759) );
  XNOR U13826 ( .A(n13777), .B(n13778), .Z(n13776) );
  ANDN U13827 ( .B(n13779), .A(n13780), .Z(n13777) );
  XNOR U13828 ( .A(n13781), .B(n13782), .Z(n13779) );
  IV U13829 ( .A(n13757), .Z(n13775) );
  XOR U13830 ( .A(n13783), .B(n13784), .Z(n13757) );
  ANDN U13831 ( .B(n13785), .A(n13786), .Z(n13783) );
  XOR U13832 ( .A(n13784), .B(n13787), .Z(n13785) );
  XOR U13833 ( .A(n13766), .B(n13697), .Z(n13767) );
  XOR U13834 ( .A(n13788), .B(n13789), .Z(n13697) );
  AND U13835 ( .A(n342), .B(n13790), .Z(n13788) );
  XOR U13836 ( .A(n13791), .B(n13789), .Z(n13790) );
  XNOR U13837 ( .A(n13792), .B(n13793), .Z(n13766) );
  NAND U13838 ( .A(n13794), .B(n13795), .Z(n13793) );
  XOR U13839 ( .A(n13796), .B(n13745), .Z(n13795) );
  XOR U13840 ( .A(n13786), .B(n13787), .Z(n13745) );
  XOR U13841 ( .A(n13797), .B(n13774), .Z(n13787) );
  XOR U13842 ( .A(n13798), .B(n13799), .Z(n13774) );
  ANDN U13843 ( .B(n13800), .A(n13801), .Z(n13798) );
  XOR U13844 ( .A(n13799), .B(n13802), .Z(n13800) );
  IV U13845 ( .A(n13772), .Z(n13797) );
  XOR U13846 ( .A(n13770), .B(n13803), .Z(n13772) );
  XOR U13847 ( .A(n13804), .B(n13805), .Z(n13803) );
  ANDN U13848 ( .B(n13806), .A(n13807), .Z(n13804) );
  XOR U13849 ( .A(n13808), .B(n13805), .Z(n13806) );
  IV U13850 ( .A(n13773), .Z(n13770) );
  XOR U13851 ( .A(n13809), .B(n13810), .Z(n13773) );
  ANDN U13852 ( .B(n13811), .A(n13812), .Z(n13809) );
  XOR U13853 ( .A(n13810), .B(n13813), .Z(n13811) );
  XOR U13854 ( .A(n13814), .B(n13815), .Z(n13786) );
  XNOR U13855 ( .A(n13781), .B(n13816), .Z(n13815) );
  IV U13856 ( .A(n13784), .Z(n13816) );
  XOR U13857 ( .A(n13817), .B(n13818), .Z(n13784) );
  ANDN U13858 ( .B(n13819), .A(n13820), .Z(n13817) );
  XOR U13859 ( .A(n13818), .B(n13821), .Z(n13819) );
  XNOR U13860 ( .A(n13822), .B(n13823), .Z(n13781) );
  ANDN U13861 ( .B(n13824), .A(n13825), .Z(n13822) );
  XOR U13862 ( .A(n13823), .B(n13826), .Z(n13824) );
  IV U13863 ( .A(n13780), .Z(n13814) );
  XOR U13864 ( .A(n13778), .B(n13827), .Z(n13780) );
  XOR U13865 ( .A(n13828), .B(n13829), .Z(n13827) );
  ANDN U13866 ( .B(n13830), .A(n13831), .Z(n13828) );
  XOR U13867 ( .A(n13832), .B(n13829), .Z(n13830) );
  IV U13868 ( .A(n13782), .Z(n13778) );
  XOR U13869 ( .A(n13833), .B(n13834), .Z(n13782) );
  ANDN U13870 ( .B(n13835), .A(n13836), .Z(n13833) );
  XOR U13871 ( .A(n13837), .B(n13834), .Z(n13835) );
  IV U13872 ( .A(n13792), .Z(n13796) );
  XOR U13873 ( .A(n13792), .B(n13747), .Z(n13794) );
  XOR U13874 ( .A(n13838), .B(n13839), .Z(n13747) );
  AND U13875 ( .A(n342), .B(n13840), .Z(n13838) );
  XOR U13876 ( .A(n13841), .B(n13839), .Z(n13840) );
  NANDN U13877 ( .A(n13749), .B(n13751), .Z(n13792) );
  XOR U13878 ( .A(n13842), .B(n13843), .Z(n13751) );
  AND U13879 ( .A(n342), .B(n13844), .Z(n13842) );
  XOR U13880 ( .A(n13843), .B(n13845), .Z(n13844) );
  XNOR U13881 ( .A(n13846), .B(n13847), .Z(n342) );
  AND U13882 ( .A(n13848), .B(n13849), .Z(n13846) );
  XOR U13883 ( .A(n13847), .B(n13762), .Z(n13849) );
  XNOR U13884 ( .A(n13850), .B(n13851), .Z(n13762) );
  ANDN U13885 ( .B(n13852), .A(n13853), .Z(n13850) );
  XOR U13886 ( .A(n13851), .B(n13854), .Z(n13852) );
  XNOR U13887 ( .A(n13847), .B(n13764), .Z(n13848) );
  XOR U13888 ( .A(n13855), .B(n13856), .Z(n13764) );
  AND U13889 ( .A(n346), .B(n13857), .Z(n13855) );
  XOR U13890 ( .A(n13858), .B(n13856), .Z(n13857) );
  XNOR U13891 ( .A(n13859), .B(n13860), .Z(n13847) );
  AND U13892 ( .A(n13861), .B(n13862), .Z(n13859) );
  XNOR U13893 ( .A(n13860), .B(n13789), .Z(n13862) );
  XOR U13894 ( .A(n13853), .B(n13854), .Z(n13789) );
  XNOR U13895 ( .A(n13863), .B(n13864), .Z(n13854) );
  ANDN U13896 ( .B(n13865), .A(n13866), .Z(n13863) );
  XOR U13897 ( .A(n13867), .B(n13868), .Z(n13865) );
  XOR U13898 ( .A(n13869), .B(n13870), .Z(n13853) );
  XNOR U13899 ( .A(n13871), .B(n13872), .Z(n13870) );
  ANDN U13900 ( .B(n13873), .A(n13874), .Z(n13871) );
  XNOR U13901 ( .A(n13875), .B(n13876), .Z(n13873) );
  IV U13902 ( .A(n13851), .Z(n13869) );
  XOR U13903 ( .A(n13877), .B(n13878), .Z(n13851) );
  ANDN U13904 ( .B(n13879), .A(n13880), .Z(n13877) );
  XOR U13905 ( .A(n13878), .B(n13881), .Z(n13879) );
  XOR U13906 ( .A(n13860), .B(n13791), .Z(n13861) );
  XOR U13907 ( .A(n13882), .B(n13883), .Z(n13791) );
  AND U13908 ( .A(n346), .B(n13884), .Z(n13882) );
  XOR U13909 ( .A(n13885), .B(n13883), .Z(n13884) );
  XNOR U13910 ( .A(n13886), .B(n13887), .Z(n13860) );
  NAND U13911 ( .A(n13888), .B(n13889), .Z(n13887) );
  XOR U13912 ( .A(n13890), .B(n13839), .Z(n13889) );
  XOR U13913 ( .A(n13880), .B(n13881), .Z(n13839) );
  XOR U13914 ( .A(n13891), .B(n13868), .Z(n13881) );
  XOR U13915 ( .A(n13892), .B(n13893), .Z(n13868) );
  ANDN U13916 ( .B(n13894), .A(n13895), .Z(n13892) );
  XOR U13917 ( .A(n13893), .B(n13896), .Z(n13894) );
  IV U13918 ( .A(n13866), .Z(n13891) );
  XOR U13919 ( .A(n13864), .B(n13897), .Z(n13866) );
  XOR U13920 ( .A(n13898), .B(n13899), .Z(n13897) );
  ANDN U13921 ( .B(n13900), .A(n13901), .Z(n13898) );
  XOR U13922 ( .A(n13902), .B(n13899), .Z(n13900) );
  IV U13923 ( .A(n13867), .Z(n13864) );
  XOR U13924 ( .A(n13903), .B(n13904), .Z(n13867) );
  ANDN U13925 ( .B(n13905), .A(n13906), .Z(n13903) );
  XOR U13926 ( .A(n13904), .B(n13907), .Z(n13905) );
  XOR U13927 ( .A(n13908), .B(n13909), .Z(n13880) );
  XNOR U13928 ( .A(n13875), .B(n13910), .Z(n13909) );
  IV U13929 ( .A(n13878), .Z(n13910) );
  XOR U13930 ( .A(n13911), .B(n13912), .Z(n13878) );
  ANDN U13931 ( .B(n13913), .A(n13914), .Z(n13911) );
  XOR U13932 ( .A(n13912), .B(n13915), .Z(n13913) );
  XNOR U13933 ( .A(n13916), .B(n13917), .Z(n13875) );
  ANDN U13934 ( .B(n13918), .A(n13919), .Z(n13916) );
  XOR U13935 ( .A(n13917), .B(n13920), .Z(n13918) );
  IV U13936 ( .A(n13874), .Z(n13908) );
  XOR U13937 ( .A(n13872), .B(n13921), .Z(n13874) );
  XOR U13938 ( .A(n13922), .B(n13923), .Z(n13921) );
  ANDN U13939 ( .B(n13924), .A(n13925), .Z(n13922) );
  XOR U13940 ( .A(n13926), .B(n13923), .Z(n13924) );
  IV U13941 ( .A(n13876), .Z(n13872) );
  XOR U13942 ( .A(n13927), .B(n13928), .Z(n13876) );
  ANDN U13943 ( .B(n13929), .A(n13930), .Z(n13927) );
  XOR U13944 ( .A(n13931), .B(n13928), .Z(n13929) );
  IV U13945 ( .A(n13886), .Z(n13890) );
  XOR U13946 ( .A(n13886), .B(n13841), .Z(n13888) );
  XOR U13947 ( .A(n13932), .B(n13933), .Z(n13841) );
  AND U13948 ( .A(n346), .B(n13934), .Z(n13932) );
  XOR U13949 ( .A(n13935), .B(n13933), .Z(n13934) );
  NANDN U13950 ( .A(n13843), .B(n13845), .Z(n13886) );
  XOR U13951 ( .A(n13936), .B(n13937), .Z(n13845) );
  AND U13952 ( .A(n346), .B(n13938), .Z(n13936) );
  XOR U13953 ( .A(n13937), .B(n13939), .Z(n13938) );
  XNOR U13954 ( .A(n13940), .B(n13941), .Z(n346) );
  AND U13955 ( .A(n13942), .B(n13943), .Z(n13940) );
  XOR U13956 ( .A(n13941), .B(n13856), .Z(n13943) );
  XNOR U13957 ( .A(n13944), .B(n13945), .Z(n13856) );
  ANDN U13958 ( .B(n13946), .A(n13947), .Z(n13944) );
  XOR U13959 ( .A(n13945), .B(n13948), .Z(n13946) );
  XNOR U13960 ( .A(n13941), .B(n13858), .Z(n13942) );
  XOR U13961 ( .A(n13949), .B(n13950), .Z(n13858) );
  AND U13962 ( .A(n350), .B(n13951), .Z(n13949) );
  XOR U13963 ( .A(n13952), .B(n13950), .Z(n13951) );
  XNOR U13964 ( .A(n13953), .B(n13954), .Z(n13941) );
  AND U13965 ( .A(n13955), .B(n13956), .Z(n13953) );
  XNOR U13966 ( .A(n13954), .B(n13883), .Z(n13956) );
  XOR U13967 ( .A(n13947), .B(n13948), .Z(n13883) );
  XNOR U13968 ( .A(n13957), .B(n13958), .Z(n13948) );
  ANDN U13969 ( .B(n13959), .A(n13960), .Z(n13957) );
  XOR U13970 ( .A(n13961), .B(n13962), .Z(n13959) );
  XOR U13971 ( .A(n13963), .B(n13964), .Z(n13947) );
  XNOR U13972 ( .A(n13965), .B(n13966), .Z(n13964) );
  ANDN U13973 ( .B(n13967), .A(n13968), .Z(n13965) );
  XNOR U13974 ( .A(n13969), .B(n13970), .Z(n13967) );
  IV U13975 ( .A(n13945), .Z(n13963) );
  XOR U13976 ( .A(n13971), .B(n13972), .Z(n13945) );
  ANDN U13977 ( .B(n13973), .A(n13974), .Z(n13971) );
  XOR U13978 ( .A(n13972), .B(n13975), .Z(n13973) );
  XOR U13979 ( .A(n13954), .B(n13885), .Z(n13955) );
  XOR U13980 ( .A(n13976), .B(n13977), .Z(n13885) );
  AND U13981 ( .A(n350), .B(n13978), .Z(n13976) );
  XOR U13982 ( .A(n13979), .B(n13977), .Z(n13978) );
  XNOR U13983 ( .A(n13980), .B(n13981), .Z(n13954) );
  NAND U13984 ( .A(n13982), .B(n13983), .Z(n13981) );
  XOR U13985 ( .A(n13984), .B(n13933), .Z(n13983) );
  XOR U13986 ( .A(n13974), .B(n13975), .Z(n13933) );
  XOR U13987 ( .A(n13985), .B(n13962), .Z(n13975) );
  XOR U13988 ( .A(n13986), .B(n13987), .Z(n13962) );
  ANDN U13989 ( .B(n13988), .A(n13989), .Z(n13986) );
  XOR U13990 ( .A(n13987), .B(n13990), .Z(n13988) );
  IV U13991 ( .A(n13960), .Z(n13985) );
  XOR U13992 ( .A(n13958), .B(n13991), .Z(n13960) );
  XOR U13993 ( .A(n13992), .B(n13993), .Z(n13991) );
  ANDN U13994 ( .B(n13994), .A(n13995), .Z(n13992) );
  XOR U13995 ( .A(n13996), .B(n13993), .Z(n13994) );
  IV U13996 ( .A(n13961), .Z(n13958) );
  XOR U13997 ( .A(n13997), .B(n13998), .Z(n13961) );
  ANDN U13998 ( .B(n13999), .A(n14000), .Z(n13997) );
  XOR U13999 ( .A(n13998), .B(n14001), .Z(n13999) );
  XOR U14000 ( .A(n14002), .B(n14003), .Z(n13974) );
  XNOR U14001 ( .A(n13969), .B(n14004), .Z(n14003) );
  IV U14002 ( .A(n13972), .Z(n14004) );
  XOR U14003 ( .A(n14005), .B(n14006), .Z(n13972) );
  ANDN U14004 ( .B(n14007), .A(n14008), .Z(n14005) );
  XOR U14005 ( .A(n14006), .B(n14009), .Z(n14007) );
  XNOR U14006 ( .A(n14010), .B(n14011), .Z(n13969) );
  ANDN U14007 ( .B(n14012), .A(n14013), .Z(n14010) );
  XOR U14008 ( .A(n14011), .B(n14014), .Z(n14012) );
  IV U14009 ( .A(n13968), .Z(n14002) );
  XOR U14010 ( .A(n13966), .B(n14015), .Z(n13968) );
  XOR U14011 ( .A(n14016), .B(n14017), .Z(n14015) );
  ANDN U14012 ( .B(n14018), .A(n14019), .Z(n14016) );
  XOR U14013 ( .A(n14020), .B(n14017), .Z(n14018) );
  IV U14014 ( .A(n13970), .Z(n13966) );
  XOR U14015 ( .A(n14021), .B(n14022), .Z(n13970) );
  ANDN U14016 ( .B(n14023), .A(n14024), .Z(n14021) );
  XOR U14017 ( .A(n14025), .B(n14022), .Z(n14023) );
  IV U14018 ( .A(n13980), .Z(n13984) );
  XOR U14019 ( .A(n13980), .B(n13935), .Z(n13982) );
  XOR U14020 ( .A(n14026), .B(n14027), .Z(n13935) );
  AND U14021 ( .A(n350), .B(n14028), .Z(n14026) );
  XOR U14022 ( .A(n14029), .B(n14027), .Z(n14028) );
  NANDN U14023 ( .A(n13937), .B(n13939), .Z(n13980) );
  XOR U14024 ( .A(n14030), .B(n14031), .Z(n13939) );
  AND U14025 ( .A(n350), .B(n14032), .Z(n14030) );
  XOR U14026 ( .A(n14031), .B(n14033), .Z(n14032) );
  XNOR U14027 ( .A(n14034), .B(n14035), .Z(n350) );
  AND U14028 ( .A(n14036), .B(n14037), .Z(n14034) );
  XOR U14029 ( .A(n14035), .B(n13950), .Z(n14037) );
  XNOR U14030 ( .A(n14038), .B(n14039), .Z(n13950) );
  ANDN U14031 ( .B(n14040), .A(n14041), .Z(n14038) );
  XOR U14032 ( .A(n14039), .B(n14042), .Z(n14040) );
  XNOR U14033 ( .A(n14035), .B(n13952), .Z(n14036) );
  XOR U14034 ( .A(n14043), .B(n14044), .Z(n13952) );
  AND U14035 ( .A(n354), .B(n14045), .Z(n14043) );
  XOR U14036 ( .A(n14046), .B(n14044), .Z(n14045) );
  XNOR U14037 ( .A(n14047), .B(n14048), .Z(n14035) );
  AND U14038 ( .A(n14049), .B(n14050), .Z(n14047) );
  XNOR U14039 ( .A(n14048), .B(n13977), .Z(n14050) );
  XOR U14040 ( .A(n14041), .B(n14042), .Z(n13977) );
  XNOR U14041 ( .A(n14051), .B(n14052), .Z(n14042) );
  ANDN U14042 ( .B(n14053), .A(n14054), .Z(n14051) );
  XOR U14043 ( .A(n14055), .B(n14056), .Z(n14053) );
  XOR U14044 ( .A(n14057), .B(n14058), .Z(n14041) );
  XNOR U14045 ( .A(n14059), .B(n14060), .Z(n14058) );
  ANDN U14046 ( .B(n14061), .A(n14062), .Z(n14059) );
  XNOR U14047 ( .A(n14063), .B(n14064), .Z(n14061) );
  IV U14048 ( .A(n14039), .Z(n14057) );
  XOR U14049 ( .A(n14065), .B(n14066), .Z(n14039) );
  ANDN U14050 ( .B(n14067), .A(n14068), .Z(n14065) );
  XOR U14051 ( .A(n14066), .B(n14069), .Z(n14067) );
  XOR U14052 ( .A(n14048), .B(n13979), .Z(n14049) );
  XOR U14053 ( .A(n14070), .B(n14071), .Z(n13979) );
  AND U14054 ( .A(n354), .B(n14072), .Z(n14070) );
  XOR U14055 ( .A(n14073), .B(n14071), .Z(n14072) );
  XNOR U14056 ( .A(n14074), .B(n14075), .Z(n14048) );
  NAND U14057 ( .A(n14076), .B(n14077), .Z(n14075) );
  XOR U14058 ( .A(n14078), .B(n14027), .Z(n14077) );
  XOR U14059 ( .A(n14068), .B(n14069), .Z(n14027) );
  XOR U14060 ( .A(n14079), .B(n14056), .Z(n14069) );
  XOR U14061 ( .A(n14080), .B(n14081), .Z(n14056) );
  ANDN U14062 ( .B(n14082), .A(n14083), .Z(n14080) );
  XOR U14063 ( .A(n14081), .B(n14084), .Z(n14082) );
  IV U14064 ( .A(n14054), .Z(n14079) );
  XOR U14065 ( .A(n14052), .B(n14085), .Z(n14054) );
  XOR U14066 ( .A(n14086), .B(n14087), .Z(n14085) );
  ANDN U14067 ( .B(n14088), .A(n14089), .Z(n14086) );
  XOR U14068 ( .A(n14090), .B(n14087), .Z(n14088) );
  IV U14069 ( .A(n14055), .Z(n14052) );
  XOR U14070 ( .A(n14091), .B(n14092), .Z(n14055) );
  ANDN U14071 ( .B(n14093), .A(n14094), .Z(n14091) );
  XOR U14072 ( .A(n14092), .B(n14095), .Z(n14093) );
  XOR U14073 ( .A(n14096), .B(n14097), .Z(n14068) );
  XNOR U14074 ( .A(n14063), .B(n14098), .Z(n14097) );
  IV U14075 ( .A(n14066), .Z(n14098) );
  XOR U14076 ( .A(n14099), .B(n14100), .Z(n14066) );
  ANDN U14077 ( .B(n14101), .A(n14102), .Z(n14099) );
  XOR U14078 ( .A(n14100), .B(n14103), .Z(n14101) );
  XNOR U14079 ( .A(n14104), .B(n14105), .Z(n14063) );
  ANDN U14080 ( .B(n14106), .A(n14107), .Z(n14104) );
  XOR U14081 ( .A(n14105), .B(n14108), .Z(n14106) );
  IV U14082 ( .A(n14062), .Z(n14096) );
  XOR U14083 ( .A(n14060), .B(n14109), .Z(n14062) );
  XOR U14084 ( .A(n14110), .B(n14111), .Z(n14109) );
  ANDN U14085 ( .B(n14112), .A(n14113), .Z(n14110) );
  XOR U14086 ( .A(n14114), .B(n14111), .Z(n14112) );
  IV U14087 ( .A(n14064), .Z(n14060) );
  XOR U14088 ( .A(n14115), .B(n14116), .Z(n14064) );
  ANDN U14089 ( .B(n14117), .A(n14118), .Z(n14115) );
  XOR U14090 ( .A(n14119), .B(n14116), .Z(n14117) );
  IV U14091 ( .A(n14074), .Z(n14078) );
  XOR U14092 ( .A(n14074), .B(n14029), .Z(n14076) );
  XOR U14093 ( .A(n14120), .B(n14121), .Z(n14029) );
  AND U14094 ( .A(n354), .B(n14122), .Z(n14120) );
  XOR U14095 ( .A(n14123), .B(n14121), .Z(n14122) );
  NANDN U14096 ( .A(n14031), .B(n14033), .Z(n14074) );
  XOR U14097 ( .A(n14124), .B(n14125), .Z(n14033) );
  AND U14098 ( .A(n354), .B(n14126), .Z(n14124) );
  XOR U14099 ( .A(n14125), .B(n14127), .Z(n14126) );
  XNOR U14100 ( .A(n14128), .B(n14129), .Z(n354) );
  AND U14101 ( .A(n14130), .B(n14131), .Z(n14128) );
  XOR U14102 ( .A(n14129), .B(n14044), .Z(n14131) );
  XNOR U14103 ( .A(n14132), .B(n14133), .Z(n14044) );
  ANDN U14104 ( .B(n14134), .A(n14135), .Z(n14132) );
  XOR U14105 ( .A(n14133), .B(n14136), .Z(n14134) );
  XNOR U14106 ( .A(n14129), .B(n14046), .Z(n14130) );
  XOR U14107 ( .A(n14137), .B(n14138), .Z(n14046) );
  AND U14108 ( .A(n358), .B(n14139), .Z(n14137) );
  XOR U14109 ( .A(n14140), .B(n14138), .Z(n14139) );
  XNOR U14110 ( .A(n14141), .B(n14142), .Z(n14129) );
  AND U14111 ( .A(n14143), .B(n14144), .Z(n14141) );
  XNOR U14112 ( .A(n14142), .B(n14071), .Z(n14144) );
  XOR U14113 ( .A(n14135), .B(n14136), .Z(n14071) );
  XNOR U14114 ( .A(n14145), .B(n14146), .Z(n14136) );
  ANDN U14115 ( .B(n14147), .A(n14148), .Z(n14145) );
  XOR U14116 ( .A(n14149), .B(n14150), .Z(n14147) );
  XOR U14117 ( .A(n14151), .B(n14152), .Z(n14135) );
  XNOR U14118 ( .A(n14153), .B(n14154), .Z(n14152) );
  ANDN U14119 ( .B(n14155), .A(n14156), .Z(n14153) );
  XNOR U14120 ( .A(n14157), .B(n14158), .Z(n14155) );
  IV U14121 ( .A(n14133), .Z(n14151) );
  XOR U14122 ( .A(n14159), .B(n14160), .Z(n14133) );
  ANDN U14123 ( .B(n14161), .A(n14162), .Z(n14159) );
  XOR U14124 ( .A(n14160), .B(n14163), .Z(n14161) );
  XOR U14125 ( .A(n14142), .B(n14073), .Z(n14143) );
  XOR U14126 ( .A(n14164), .B(n14165), .Z(n14073) );
  AND U14127 ( .A(n358), .B(n14166), .Z(n14164) );
  XOR U14128 ( .A(n14167), .B(n14165), .Z(n14166) );
  XNOR U14129 ( .A(n14168), .B(n14169), .Z(n14142) );
  NAND U14130 ( .A(n14170), .B(n14171), .Z(n14169) );
  XOR U14131 ( .A(n14172), .B(n14121), .Z(n14171) );
  XOR U14132 ( .A(n14162), .B(n14163), .Z(n14121) );
  XOR U14133 ( .A(n14173), .B(n14150), .Z(n14163) );
  XOR U14134 ( .A(n14174), .B(n14175), .Z(n14150) );
  ANDN U14135 ( .B(n14176), .A(n14177), .Z(n14174) );
  XOR U14136 ( .A(n14175), .B(n14178), .Z(n14176) );
  IV U14137 ( .A(n14148), .Z(n14173) );
  XOR U14138 ( .A(n14146), .B(n14179), .Z(n14148) );
  XOR U14139 ( .A(n14180), .B(n14181), .Z(n14179) );
  ANDN U14140 ( .B(n14182), .A(n14183), .Z(n14180) );
  XOR U14141 ( .A(n14184), .B(n14181), .Z(n14182) );
  IV U14142 ( .A(n14149), .Z(n14146) );
  XOR U14143 ( .A(n14185), .B(n14186), .Z(n14149) );
  ANDN U14144 ( .B(n14187), .A(n14188), .Z(n14185) );
  XOR U14145 ( .A(n14186), .B(n14189), .Z(n14187) );
  XOR U14146 ( .A(n14190), .B(n14191), .Z(n14162) );
  XNOR U14147 ( .A(n14157), .B(n14192), .Z(n14191) );
  IV U14148 ( .A(n14160), .Z(n14192) );
  XOR U14149 ( .A(n14193), .B(n14194), .Z(n14160) );
  ANDN U14150 ( .B(n14195), .A(n14196), .Z(n14193) );
  XOR U14151 ( .A(n14194), .B(n14197), .Z(n14195) );
  XNOR U14152 ( .A(n14198), .B(n14199), .Z(n14157) );
  ANDN U14153 ( .B(n14200), .A(n14201), .Z(n14198) );
  XOR U14154 ( .A(n14199), .B(n14202), .Z(n14200) );
  IV U14155 ( .A(n14156), .Z(n14190) );
  XOR U14156 ( .A(n14154), .B(n14203), .Z(n14156) );
  XOR U14157 ( .A(n14204), .B(n14205), .Z(n14203) );
  ANDN U14158 ( .B(n14206), .A(n14207), .Z(n14204) );
  XOR U14159 ( .A(n14208), .B(n14205), .Z(n14206) );
  IV U14160 ( .A(n14158), .Z(n14154) );
  XOR U14161 ( .A(n14209), .B(n14210), .Z(n14158) );
  ANDN U14162 ( .B(n14211), .A(n14212), .Z(n14209) );
  XOR U14163 ( .A(n14213), .B(n14210), .Z(n14211) );
  IV U14164 ( .A(n14168), .Z(n14172) );
  XOR U14165 ( .A(n14168), .B(n14123), .Z(n14170) );
  XOR U14166 ( .A(n14214), .B(n14215), .Z(n14123) );
  AND U14167 ( .A(n358), .B(n14216), .Z(n14214) );
  XOR U14168 ( .A(n14217), .B(n14215), .Z(n14216) );
  NANDN U14169 ( .A(n14125), .B(n14127), .Z(n14168) );
  XOR U14170 ( .A(n14218), .B(n14219), .Z(n14127) );
  AND U14171 ( .A(n358), .B(n14220), .Z(n14218) );
  XOR U14172 ( .A(n14219), .B(n14221), .Z(n14220) );
  XNOR U14173 ( .A(n14222), .B(n14223), .Z(n358) );
  AND U14174 ( .A(n14224), .B(n14225), .Z(n14222) );
  XOR U14175 ( .A(n14223), .B(n14138), .Z(n14225) );
  XNOR U14176 ( .A(n14226), .B(n14227), .Z(n14138) );
  ANDN U14177 ( .B(n14228), .A(n14229), .Z(n14226) );
  XOR U14178 ( .A(n14227), .B(n14230), .Z(n14228) );
  XNOR U14179 ( .A(n14223), .B(n14140), .Z(n14224) );
  XOR U14180 ( .A(n14231), .B(n14232), .Z(n14140) );
  AND U14181 ( .A(n362), .B(n14233), .Z(n14231) );
  XOR U14182 ( .A(n14234), .B(n14232), .Z(n14233) );
  XNOR U14183 ( .A(n14235), .B(n14236), .Z(n14223) );
  AND U14184 ( .A(n14237), .B(n14238), .Z(n14235) );
  XNOR U14185 ( .A(n14236), .B(n14165), .Z(n14238) );
  XOR U14186 ( .A(n14229), .B(n14230), .Z(n14165) );
  XNOR U14187 ( .A(n14239), .B(n14240), .Z(n14230) );
  ANDN U14188 ( .B(n14241), .A(n14242), .Z(n14239) );
  XOR U14189 ( .A(n14243), .B(n14244), .Z(n14241) );
  XOR U14190 ( .A(n14245), .B(n14246), .Z(n14229) );
  XNOR U14191 ( .A(n14247), .B(n14248), .Z(n14246) );
  ANDN U14192 ( .B(n14249), .A(n14250), .Z(n14247) );
  XNOR U14193 ( .A(n14251), .B(n14252), .Z(n14249) );
  IV U14194 ( .A(n14227), .Z(n14245) );
  XOR U14195 ( .A(n14253), .B(n14254), .Z(n14227) );
  ANDN U14196 ( .B(n14255), .A(n14256), .Z(n14253) );
  XOR U14197 ( .A(n14254), .B(n14257), .Z(n14255) );
  XOR U14198 ( .A(n14236), .B(n14167), .Z(n14237) );
  XOR U14199 ( .A(n14258), .B(n14259), .Z(n14167) );
  AND U14200 ( .A(n362), .B(n14260), .Z(n14258) );
  XOR U14201 ( .A(n14261), .B(n14259), .Z(n14260) );
  XNOR U14202 ( .A(n14262), .B(n14263), .Z(n14236) );
  NAND U14203 ( .A(n14264), .B(n14265), .Z(n14263) );
  XOR U14204 ( .A(n14266), .B(n14215), .Z(n14265) );
  XOR U14205 ( .A(n14256), .B(n14257), .Z(n14215) );
  XOR U14206 ( .A(n14267), .B(n14244), .Z(n14257) );
  XOR U14207 ( .A(n14268), .B(n14269), .Z(n14244) );
  ANDN U14208 ( .B(n14270), .A(n14271), .Z(n14268) );
  XOR U14209 ( .A(n14269), .B(n14272), .Z(n14270) );
  IV U14210 ( .A(n14242), .Z(n14267) );
  XOR U14211 ( .A(n14240), .B(n14273), .Z(n14242) );
  XOR U14212 ( .A(n14274), .B(n14275), .Z(n14273) );
  ANDN U14213 ( .B(n14276), .A(n14277), .Z(n14274) );
  XOR U14214 ( .A(n14278), .B(n14275), .Z(n14276) );
  IV U14215 ( .A(n14243), .Z(n14240) );
  XOR U14216 ( .A(n14279), .B(n14280), .Z(n14243) );
  ANDN U14217 ( .B(n14281), .A(n14282), .Z(n14279) );
  XOR U14218 ( .A(n14280), .B(n14283), .Z(n14281) );
  XOR U14219 ( .A(n14284), .B(n14285), .Z(n14256) );
  XNOR U14220 ( .A(n14251), .B(n14286), .Z(n14285) );
  IV U14221 ( .A(n14254), .Z(n14286) );
  XOR U14222 ( .A(n14287), .B(n14288), .Z(n14254) );
  ANDN U14223 ( .B(n14289), .A(n14290), .Z(n14287) );
  XOR U14224 ( .A(n14288), .B(n14291), .Z(n14289) );
  XNOR U14225 ( .A(n14292), .B(n14293), .Z(n14251) );
  ANDN U14226 ( .B(n14294), .A(n14295), .Z(n14292) );
  XOR U14227 ( .A(n14293), .B(n14296), .Z(n14294) );
  IV U14228 ( .A(n14250), .Z(n14284) );
  XOR U14229 ( .A(n14248), .B(n14297), .Z(n14250) );
  XOR U14230 ( .A(n14298), .B(n14299), .Z(n14297) );
  ANDN U14231 ( .B(n14300), .A(n14301), .Z(n14298) );
  XOR U14232 ( .A(n14302), .B(n14299), .Z(n14300) );
  IV U14233 ( .A(n14252), .Z(n14248) );
  XOR U14234 ( .A(n14303), .B(n14304), .Z(n14252) );
  ANDN U14235 ( .B(n14305), .A(n14306), .Z(n14303) );
  XOR U14236 ( .A(n14307), .B(n14304), .Z(n14305) );
  IV U14237 ( .A(n14262), .Z(n14266) );
  XOR U14238 ( .A(n14262), .B(n14217), .Z(n14264) );
  XOR U14239 ( .A(n14308), .B(n14309), .Z(n14217) );
  AND U14240 ( .A(n362), .B(n14310), .Z(n14308) );
  XOR U14241 ( .A(n14311), .B(n14309), .Z(n14310) );
  NANDN U14242 ( .A(n14219), .B(n14221), .Z(n14262) );
  XOR U14243 ( .A(n14312), .B(n14313), .Z(n14221) );
  AND U14244 ( .A(n362), .B(n14314), .Z(n14312) );
  XOR U14245 ( .A(n14313), .B(n14315), .Z(n14314) );
  XNOR U14246 ( .A(n14316), .B(n14317), .Z(n362) );
  AND U14247 ( .A(n14318), .B(n14319), .Z(n14316) );
  XOR U14248 ( .A(n14317), .B(n14232), .Z(n14319) );
  XNOR U14249 ( .A(n14320), .B(n14321), .Z(n14232) );
  ANDN U14250 ( .B(n14322), .A(n14323), .Z(n14320) );
  XOR U14251 ( .A(n14321), .B(n14324), .Z(n14322) );
  XNOR U14252 ( .A(n14317), .B(n14234), .Z(n14318) );
  XOR U14253 ( .A(n14325), .B(n14326), .Z(n14234) );
  AND U14254 ( .A(n366), .B(n14327), .Z(n14325) );
  XOR U14255 ( .A(n14328), .B(n14326), .Z(n14327) );
  XNOR U14256 ( .A(n14329), .B(n14330), .Z(n14317) );
  AND U14257 ( .A(n14331), .B(n14332), .Z(n14329) );
  XNOR U14258 ( .A(n14330), .B(n14259), .Z(n14332) );
  XOR U14259 ( .A(n14323), .B(n14324), .Z(n14259) );
  XNOR U14260 ( .A(n14333), .B(n14334), .Z(n14324) );
  ANDN U14261 ( .B(n14335), .A(n14336), .Z(n14333) );
  XOR U14262 ( .A(n14337), .B(n14338), .Z(n14335) );
  XOR U14263 ( .A(n14339), .B(n14340), .Z(n14323) );
  XNOR U14264 ( .A(n14341), .B(n14342), .Z(n14340) );
  ANDN U14265 ( .B(n14343), .A(n14344), .Z(n14341) );
  XNOR U14266 ( .A(n14345), .B(n14346), .Z(n14343) );
  IV U14267 ( .A(n14321), .Z(n14339) );
  XOR U14268 ( .A(n14347), .B(n14348), .Z(n14321) );
  ANDN U14269 ( .B(n14349), .A(n14350), .Z(n14347) );
  XOR U14270 ( .A(n14348), .B(n14351), .Z(n14349) );
  XOR U14271 ( .A(n14330), .B(n14261), .Z(n14331) );
  XOR U14272 ( .A(n14352), .B(n14353), .Z(n14261) );
  AND U14273 ( .A(n366), .B(n14354), .Z(n14352) );
  XOR U14274 ( .A(n14355), .B(n14353), .Z(n14354) );
  XNOR U14275 ( .A(n14356), .B(n14357), .Z(n14330) );
  NAND U14276 ( .A(n14358), .B(n14359), .Z(n14357) );
  XOR U14277 ( .A(n14360), .B(n14309), .Z(n14359) );
  XOR U14278 ( .A(n14350), .B(n14351), .Z(n14309) );
  XOR U14279 ( .A(n14361), .B(n14338), .Z(n14351) );
  XOR U14280 ( .A(n14362), .B(n14363), .Z(n14338) );
  ANDN U14281 ( .B(n14364), .A(n14365), .Z(n14362) );
  XOR U14282 ( .A(n14363), .B(n14366), .Z(n14364) );
  IV U14283 ( .A(n14336), .Z(n14361) );
  XOR U14284 ( .A(n14334), .B(n14367), .Z(n14336) );
  XOR U14285 ( .A(n14368), .B(n14369), .Z(n14367) );
  ANDN U14286 ( .B(n14370), .A(n14371), .Z(n14368) );
  XOR U14287 ( .A(n14372), .B(n14369), .Z(n14370) );
  IV U14288 ( .A(n14337), .Z(n14334) );
  XOR U14289 ( .A(n14373), .B(n14374), .Z(n14337) );
  ANDN U14290 ( .B(n14375), .A(n14376), .Z(n14373) );
  XOR U14291 ( .A(n14374), .B(n14377), .Z(n14375) );
  XOR U14292 ( .A(n14378), .B(n14379), .Z(n14350) );
  XNOR U14293 ( .A(n14345), .B(n14380), .Z(n14379) );
  IV U14294 ( .A(n14348), .Z(n14380) );
  XOR U14295 ( .A(n14381), .B(n14382), .Z(n14348) );
  ANDN U14296 ( .B(n14383), .A(n14384), .Z(n14381) );
  XOR U14297 ( .A(n14382), .B(n14385), .Z(n14383) );
  XNOR U14298 ( .A(n14386), .B(n14387), .Z(n14345) );
  ANDN U14299 ( .B(n14388), .A(n14389), .Z(n14386) );
  XOR U14300 ( .A(n14387), .B(n14390), .Z(n14388) );
  IV U14301 ( .A(n14344), .Z(n14378) );
  XOR U14302 ( .A(n14342), .B(n14391), .Z(n14344) );
  XOR U14303 ( .A(n14392), .B(n14393), .Z(n14391) );
  ANDN U14304 ( .B(n14394), .A(n14395), .Z(n14392) );
  XOR U14305 ( .A(n14396), .B(n14393), .Z(n14394) );
  IV U14306 ( .A(n14346), .Z(n14342) );
  XOR U14307 ( .A(n14397), .B(n14398), .Z(n14346) );
  ANDN U14308 ( .B(n14399), .A(n14400), .Z(n14397) );
  XOR U14309 ( .A(n14401), .B(n14398), .Z(n14399) );
  IV U14310 ( .A(n14356), .Z(n14360) );
  XOR U14311 ( .A(n14356), .B(n14311), .Z(n14358) );
  XOR U14312 ( .A(n14402), .B(n14403), .Z(n14311) );
  AND U14313 ( .A(n366), .B(n14404), .Z(n14402) );
  XOR U14314 ( .A(n14405), .B(n14403), .Z(n14404) );
  NANDN U14315 ( .A(n14313), .B(n14315), .Z(n14356) );
  XOR U14316 ( .A(n14406), .B(n14407), .Z(n14315) );
  AND U14317 ( .A(n366), .B(n14408), .Z(n14406) );
  XOR U14318 ( .A(n14407), .B(n14409), .Z(n14408) );
  XNOR U14319 ( .A(n14410), .B(n14411), .Z(n366) );
  AND U14320 ( .A(n14412), .B(n14413), .Z(n14410) );
  XOR U14321 ( .A(n14411), .B(n14326), .Z(n14413) );
  XNOR U14322 ( .A(n14414), .B(n14415), .Z(n14326) );
  ANDN U14323 ( .B(n14416), .A(n14417), .Z(n14414) );
  XOR U14324 ( .A(n14415), .B(n14418), .Z(n14416) );
  XNOR U14325 ( .A(n14411), .B(n14328), .Z(n14412) );
  XOR U14326 ( .A(n14419), .B(n14420), .Z(n14328) );
  AND U14327 ( .A(n370), .B(n14421), .Z(n14419) );
  XOR U14328 ( .A(n14422), .B(n14420), .Z(n14421) );
  XNOR U14329 ( .A(n14423), .B(n14424), .Z(n14411) );
  AND U14330 ( .A(n14425), .B(n14426), .Z(n14423) );
  XNOR U14331 ( .A(n14424), .B(n14353), .Z(n14426) );
  XOR U14332 ( .A(n14417), .B(n14418), .Z(n14353) );
  XNOR U14333 ( .A(n14427), .B(n14428), .Z(n14418) );
  ANDN U14334 ( .B(n14429), .A(n14430), .Z(n14427) );
  XOR U14335 ( .A(n14431), .B(n14432), .Z(n14429) );
  XOR U14336 ( .A(n14433), .B(n14434), .Z(n14417) );
  XNOR U14337 ( .A(n14435), .B(n14436), .Z(n14434) );
  ANDN U14338 ( .B(n14437), .A(n14438), .Z(n14435) );
  XNOR U14339 ( .A(n14439), .B(n14440), .Z(n14437) );
  IV U14340 ( .A(n14415), .Z(n14433) );
  XOR U14341 ( .A(n14441), .B(n14442), .Z(n14415) );
  ANDN U14342 ( .B(n14443), .A(n14444), .Z(n14441) );
  XOR U14343 ( .A(n14442), .B(n14445), .Z(n14443) );
  XOR U14344 ( .A(n14424), .B(n14355), .Z(n14425) );
  XOR U14345 ( .A(n14446), .B(n14447), .Z(n14355) );
  AND U14346 ( .A(n370), .B(n14448), .Z(n14446) );
  XOR U14347 ( .A(n14449), .B(n14447), .Z(n14448) );
  XNOR U14348 ( .A(n14450), .B(n14451), .Z(n14424) );
  NAND U14349 ( .A(n14452), .B(n14453), .Z(n14451) );
  XOR U14350 ( .A(n14454), .B(n14403), .Z(n14453) );
  XOR U14351 ( .A(n14444), .B(n14445), .Z(n14403) );
  XOR U14352 ( .A(n14455), .B(n14432), .Z(n14445) );
  XOR U14353 ( .A(n14456), .B(n14457), .Z(n14432) );
  ANDN U14354 ( .B(n14458), .A(n14459), .Z(n14456) );
  XOR U14355 ( .A(n14457), .B(n14460), .Z(n14458) );
  IV U14356 ( .A(n14430), .Z(n14455) );
  XOR U14357 ( .A(n14428), .B(n14461), .Z(n14430) );
  XOR U14358 ( .A(n14462), .B(n14463), .Z(n14461) );
  ANDN U14359 ( .B(n14464), .A(n14465), .Z(n14462) );
  XOR U14360 ( .A(n14466), .B(n14463), .Z(n14464) );
  IV U14361 ( .A(n14431), .Z(n14428) );
  XOR U14362 ( .A(n14467), .B(n14468), .Z(n14431) );
  ANDN U14363 ( .B(n14469), .A(n14470), .Z(n14467) );
  XOR U14364 ( .A(n14468), .B(n14471), .Z(n14469) );
  XOR U14365 ( .A(n14472), .B(n14473), .Z(n14444) );
  XNOR U14366 ( .A(n14439), .B(n14474), .Z(n14473) );
  IV U14367 ( .A(n14442), .Z(n14474) );
  XOR U14368 ( .A(n14475), .B(n14476), .Z(n14442) );
  ANDN U14369 ( .B(n14477), .A(n14478), .Z(n14475) );
  XOR U14370 ( .A(n14476), .B(n14479), .Z(n14477) );
  XNOR U14371 ( .A(n14480), .B(n14481), .Z(n14439) );
  ANDN U14372 ( .B(n14482), .A(n14483), .Z(n14480) );
  XOR U14373 ( .A(n14481), .B(n14484), .Z(n14482) );
  IV U14374 ( .A(n14438), .Z(n14472) );
  XOR U14375 ( .A(n14436), .B(n14485), .Z(n14438) );
  XOR U14376 ( .A(n14486), .B(n14487), .Z(n14485) );
  ANDN U14377 ( .B(n14488), .A(n14489), .Z(n14486) );
  XOR U14378 ( .A(n14490), .B(n14487), .Z(n14488) );
  IV U14379 ( .A(n14440), .Z(n14436) );
  XOR U14380 ( .A(n14491), .B(n14492), .Z(n14440) );
  ANDN U14381 ( .B(n14493), .A(n14494), .Z(n14491) );
  XOR U14382 ( .A(n14495), .B(n14492), .Z(n14493) );
  IV U14383 ( .A(n14450), .Z(n14454) );
  XOR U14384 ( .A(n14450), .B(n14405), .Z(n14452) );
  XOR U14385 ( .A(n14496), .B(n14497), .Z(n14405) );
  AND U14386 ( .A(n370), .B(n14498), .Z(n14496) );
  XOR U14387 ( .A(n14499), .B(n14497), .Z(n14498) );
  NANDN U14388 ( .A(n14407), .B(n14409), .Z(n14450) );
  XOR U14389 ( .A(n14500), .B(n14501), .Z(n14409) );
  AND U14390 ( .A(n370), .B(n14502), .Z(n14500) );
  XOR U14391 ( .A(n14501), .B(n14503), .Z(n14502) );
  XNOR U14392 ( .A(n14504), .B(n14505), .Z(n370) );
  AND U14393 ( .A(n14506), .B(n14507), .Z(n14504) );
  XOR U14394 ( .A(n14505), .B(n14420), .Z(n14507) );
  XNOR U14395 ( .A(n14508), .B(n14509), .Z(n14420) );
  ANDN U14396 ( .B(n14510), .A(n14511), .Z(n14508) );
  XOR U14397 ( .A(n14509), .B(n14512), .Z(n14510) );
  XNOR U14398 ( .A(n14505), .B(n14422), .Z(n14506) );
  XOR U14399 ( .A(n14513), .B(n14514), .Z(n14422) );
  AND U14400 ( .A(n374), .B(n14515), .Z(n14513) );
  XOR U14401 ( .A(n14516), .B(n14514), .Z(n14515) );
  XNOR U14402 ( .A(n14517), .B(n14518), .Z(n14505) );
  AND U14403 ( .A(n14519), .B(n14520), .Z(n14517) );
  XNOR U14404 ( .A(n14518), .B(n14447), .Z(n14520) );
  XOR U14405 ( .A(n14511), .B(n14512), .Z(n14447) );
  XNOR U14406 ( .A(n14521), .B(n14522), .Z(n14512) );
  ANDN U14407 ( .B(n14523), .A(n14524), .Z(n14521) );
  XOR U14408 ( .A(n14525), .B(n14526), .Z(n14523) );
  XOR U14409 ( .A(n14527), .B(n14528), .Z(n14511) );
  XNOR U14410 ( .A(n14529), .B(n14530), .Z(n14528) );
  ANDN U14411 ( .B(n14531), .A(n14532), .Z(n14529) );
  XNOR U14412 ( .A(n14533), .B(n14534), .Z(n14531) );
  IV U14413 ( .A(n14509), .Z(n14527) );
  XOR U14414 ( .A(n14535), .B(n14536), .Z(n14509) );
  ANDN U14415 ( .B(n14537), .A(n14538), .Z(n14535) );
  XOR U14416 ( .A(n14536), .B(n14539), .Z(n14537) );
  XOR U14417 ( .A(n14518), .B(n14449), .Z(n14519) );
  XOR U14418 ( .A(n14540), .B(n14541), .Z(n14449) );
  AND U14419 ( .A(n374), .B(n14542), .Z(n14540) );
  XOR U14420 ( .A(n14543), .B(n14541), .Z(n14542) );
  XNOR U14421 ( .A(n14544), .B(n14545), .Z(n14518) );
  NAND U14422 ( .A(n14546), .B(n14547), .Z(n14545) );
  XOR U14423 ( .A(n14548), .B(n14497), .Z(n14547) );
  XOR U14424 ( .A(n14538), .B(n14539), .Z(n14497) );
  XOR U14425 ( .A(n14549), .B(n14526), .Z(n14539) );
  XOR U14426 ( .A(n14550), .B(n14551), .Z(n14526) );
  ANDN U14427 ( .B(n14552), .A(n14553), .Z(n14550) );
  XOR U14428 ( .A(n14551), .B(n14554), .Z(n14552) );
  IV U14429 ( .A(n14524), .Z(n14549) );
  XOR U14430 ( .A(n14522), .B(n14555), .Z(n14524) );
  XOR U14431 ( .A(n14556), .B(n14557), .Z(n14555) );
  ANDN U14432 ( .B(n14558), .A(n14559), .Z(n14556) );
  XOR U14433 ( .A(n14560), .B(n14557), .Z(n14558) );
  IV U14434 ( .A(n14525), .Z(n14522) );
  XOR U14435 ( .A(n14561), .B(n14562), .Z(n14525) );
  ANDN U14436 ( .B(n14563), .A(n14564), .Z(n14561) );
  XOR U14437 ( .A(n14562), .B(n14565), .Z(n14563) );
  XOR U14438 ( .A(n14566), .B(n14567), .Z(n14538) );
  XNOR U14439 ( .A(n14533), .B(n14568), .Z(n14567) );
  IV U14440 ( .A(n14536), .Z(n14568) );
  XOR U14441 ( .A(n14569), .B(n14570), .Z(n14536) );
  ANDN U14442 ( .B(n14571), .A(n14572), .Z(n14569) );
  XOR U14443 ( .A(n14570), .B(n14573), .Z(n14571) );
  XNOR U14444 ( .A(n14574), .B(n14575), .Z(n14533) );
  ANDN U14445 ( .B(n14576), .A(n14577), .Z(n14574) );
  XOR U14446 ( .A(n14575), .B(n14578), .Z(n14576) );
  IV U14447 ( .A(n14532), .Z(n14566) );
  XOR U14448 ( .A(n14530), .B(n14579), .Z(n14532) );
  XOR U14449 ( .A(n14580), .B(n14581), .Z(n14579) );
  ANDN U14450 ( .B(n14582), .A(n14583), .Z(n14580) );
  XOR U14451 ( .A(n14584), .B(n14581), .Z(n14582) );
  IV U14452 ( .A(n14534), .Z(n14530) );
  XOR U14453 ( .A(n14585), .B(n14586), .Z(n14534) );
  ANDN U14454 ( .B(n14587), .A(n14588), .Z(n14585) );
  XOR U14455 ( .A(n14589), .B(n14586), .Z(n14587) );
  IV U14456 ( .A(n14544), .Z(n14548) );
  XOR U14457 ( .A(n14544), .B(n14499), .Z(n14546) );
  XOR U14458 ( .A(n14590), .B(n14591), .Z(n14499) );
  AND U14459 ( .A(n374), .B(n14592), .Z(n14590) );
  XOR U14460 ( .A(n14593), .B(n14591), .Z(n14592) );
  NANDN U14461 ( .A(n14501), .B(n14503), .Z(n14544) );
  XOR U14462 ( .A(n14594), .B(n14595), .Z(n14503) );
  AND U14463 ( .A(n374), .B(n14596), .Z(n14594) );
  XOR U14464 ( .A(n14595), .B(n14597), .Z(n14596) );
  XNOR U14465 ( .A(n14598), .B(n14599), .Z(n374) );
  AND U14466 ( .A(n14600), .B(n14601), .Z(n14598) );
  XOR U14467 ( .A(n14599), .B(n14514), .Z(n14601) );
  XNOR U14468 ( .A(n14602), .B(n14603), .Z(n14514) );
  ANDN U14469 ( .B(n14604), .A(n14605), .Z(n14602) );
  XOR U14470 ( .A(n14603), .B(n14606), .Z(n14604) );
  XNOR U14471 ( .A(n14599), .B(n14516), .Z(n14600) );
  XOR U14472 ( .A(n14607), .B(n14608), .Z(n14516) );
  AND U14473 ( .A(n378), .B(n14609), .Z(n14607) );
  XOR U14474 ( .A(n14610), .B(n14608), .Z(n14609) );
  XNOR U14475 ( .A(n14611), .B(n14612), .Z(n14599) );
  AND U14476 ( .A(n14613), .B(n14614), .Z(n14611) );
  XNOR U14477 ( .A(n14612), .B(n14541), .Z(n14614) );
  XOR U14478 ( .A(n14605), .B(n14606), .Z(n14541) );
  XNOR U14479 ( .A(n14615), .B(n14616), .Z(n14606) );
  ANDN U14480 ( .B(n14617), .A(n14618), .Z(n14615) );
  XOR U14481 ( .A(n14619), .B(n14620), .Z(n14617) );
  XOR U14482 ( .A(n14621), .B(n14622), .Z(n14605) );
  XNOR U14483 ( .A(n14623), .B(n14624), .Z(n14622) );
  ANDN U14484 ( .B(n14625), .A(n14626), .Z(n14623) );
  XNOR U14485 ( .A(n14627), .B(n14628), .Z(n14625) );
  IV U14486 ( .A(n14603), .Z(n14621) );
  XOR U14487 ( .A(n14629), .B(n14630), .Z(n14603) );
  ANDN U14488 ( .B(n14631), .A(n14632), .Z(n14629) );
  XOR U14489 ( .A(n14630), .B(n14633), .Z(n14631) );
  XOR U14490 ( .A(n14612), .B(n14543), .Z(n14613) );
  XOR U14491 ( .A(n14634), .B(n14635), .Z(n14543) );
  AND U14492 ( .A(n378), .B(n14636), .Z(n14634) );
  XOR U14493 ( .A(n14637), .B(n14635), .Z(n14636) );
  XNOR U14494 ( .A(n14638), .B(n14639), .Z(n14612) );
  NAND U14495 ( .A(n14640), .B(n14641), .Z(n14639) );
  XOR U14496 ( .A(n14642), .B(n14591), .Z(n14641) );
  XOR U14497 ( .A(n14632), .B(n14633), .Z(n14591) );
  XOR U14498 ( .A(n14643), .B(n14620), .Z(n14633) );
  XOR U14499 ( .A(n14644), .B(n14645), .Z(n14620) );
  ANDN U14500 ( .B(n14646), .A(n14647), .Z(n14644) );
  XOR U14501 ( .A(n14645), .B(n14648), .Z(n14646) );
  IV U14502 ( .A(n14618), .Z(n14643) );
  XOR U14503 ( .A(n14616), .B(n14649), .Z(n14618) );
  XOR U14504 ( .A(n14650), .B(n14651), .Z(n14649) );
  ANDN U14505 ( .B(n14652), .A(n14653), .Z(n14650) );
  XOR U14506 ( .A(n14654), .B(n14651), .Z(n14652) );
  IV U14507 ( .A(n14619), .Z(n14616) );
  XOR U14508 ( .A(n14655), .B(n14656), .Z(n14619) );
  ANDN U14509 ( .B(n14657), .A(n14658), .Z(n14655) );
  XOR U14510 ( .A(n14656), .B(n14659), .Z(n14657) );
  XOR U14511 ( .A(n14660), .B(n14661), .Z(n14632) );
  XNOR U14512 ( .A(n14627), .B(n14662), .Z(n14661) );
  IV U14513 ( .A(n14630), .Z(n14662) );
  XOR U14514 ( .A(n14663), .B(n14664), .Z(n14630) );
  ANDN U14515 ( .B(n14665), .A(n14666), .Z(n14663) );
  XOR U14516 ( .A(n14664), .B(n14667), .Z(n14665) );
  XNOR U14517 ( .A(n14668), .B(n14669), .Z(n14627) );
  ANDN U14518 ( .B(n14670), .A(n14671), .Z(n14668) );
  XOR U14519 ( .A(n14669), .B(n14672), .Z(n14670) );
  IV U14520 ( .A(n14626), .Z(n14660) );
  XOR U14521 ( .A(n14624), .B(n14673), .Z(n14626) );
  XOR U14522 ( .A(n14674), .B(n14675), .Z(n14673) );
  ANDN U14523 ( .B(n14676), .A(n14677), .Z(n14674) );
  XOR U14524 ( .A(n14678), .B(n14675), .Z(n14676) );
  IV U14525 ( .A(n14628), .Z(n14624) );
  XOR U14526 ( .A(n14679), .B(n14680), .Z(n14628) );
  ANDN U14527 ( .B(n14681), .A(n14682), .Z(n14679) );
  XOR U14528 ( .A(n14683), .B(n14680), .Z(n14681) );
  IV U14529 ( .A(n14638), .Z(n14642) );
  XOR U14530 ( .A(n14638), .B(n14593), .Z(n14640) );
  XOR U14531 ( .A(n14684), .B(n14685), .Z(n14593) );
  AND U14532 ( .A(n378), .B(n14686), .Z(n14684) );
  XOR U14533 ( .A(n14687), .B(n14685), .Z(n14686) );
  NANDN U14534 ( .A(n14595), .B(n14597), .Z(n14638) );
  XOR U14535 ( .A(n14688), .B(n14689), .Z(n14597) );
  AND U14536 ( .A(n378), .B(n14690), .Z(n14688) );
  XOR U14537 ( .A(n14689), .B(n14691), .Z(n14690) );
  XNOR U14538 ( .A(n14692), .B(n14693), .Z(n378) );
  AND U14539 ( .A(n14694), .B(n14695), .Z(n14692) );
  XOR U14540 ( .A(n14693), .B(n14608), .Z(n14695) );
  XNOR U14541 ( .A(n14696), .B(n14697), .Z(n14608) );
  ANDN U14542 ( .B(n14698), .A(n14699), .Z(n14696) );
  XOR U14543 ( .A(n14697), .B(n14700), .Z(n14698) );
  XNOR U14544 ( .A(n14693), .B(n14610), .Z(n14694) );
  XOR U14545 ( .A(n14701), .B(n14702), .Z(n14610) );
  AND U14546 ( .A(n382), .B(n14703), .Z(n14701) );
  XOR U14547 ( .A(n14704), .B(n14702), .Z(n14703) );
  XNOR U14548 ( .A(n14705), .B(n14706), .Z(n14693) );
  AND U14549 ( .A(n14707), .B(n14708), .Z(n14705) );
  XNOR U14550 ( .A(n14706), .B(n14635), .Z(n14708) );
  XOR U14551 ( .A(n14699), .B(n14700), .Z(n14635) );
  XNOR U14552 ( .A(n14709), .B(n14710), .Z(n14700) );
  ANDN U14553 ( .B(n14711), .A(n14712), .Z(n14709) );
  XOR U14554 ( .A(n14713), .B(n14714), .Z(n14711) );
  XOR U14555 ( .A(n14715), .B(n14716), .Z(n14699) );
  XNOR U14556 ( .A(n14717), .B(n14718), .Z(n14716) );
  ANDN U14557 ( .B(n14719), .A(n14720), .Z(n14717) );
  XNOR U14558 ( .A(n14721), .B(n14722), .Z(n14719) );
  IV U14559 ( .A(n14697), .Z(n14715) );
  XOR U14560 ( .A(n14723), .B(n14724), .Z(n14697) );
  ANDN U14561 ( .B(n14725), .A(n14726), .Z(n14723) );
  XOR U14562 ( .A(n14724), .B(n14727), .Z(n14725) );
  XOR U14563 ( .A(n14706), .B(n14637), .Z(n14707) );
  XOR U14564 ( .A(n14728), .B(n14729), .Z(n14637) );
  AND U14565 ( .A(n382), .B(n14730), .Z(n14728) );
  XOR U14566 ( .A(n14731), .B(n14729), .Z(n14730) );
  XNOR U14567 ( .A(n14732), .B(n14733), .Z(n14706) );
  NAND U14568 ( .A(n14734), .B(n14735), .Z(n14733) );
  XOR U14569 ( .A(n14736), .B(n14685), .Z(n14735) );
  XOR U14570 ( .A(n14726), .B(n14727), .Z(n14685) );
  XOR U14571 ( .A(n14737), .B(n14714), .Z(n14727) );
  XOR U14572 ( .A(n14738), .B(n14739), .Z(n14714) );
  ANDN U14573 ( .B(n14740), .A(n14741), .Z(n14738) );
  XOR U14574 ( .A(n14739), .B(n14742), .Z(n14740) );
  IV U14575 ( .A(n14712), .Z(n14737) );
  XOR U14576 ( .A(n14710), .B(n14743), .Z(n14712) );
  XOR U14577 ( .A(n14744), .B(n14745), .Z(n14743) );
  ANDN U14578 ( .B(n14746), .A(n14747), .Z(n14744) );
  XOR U14579 ( .A(n14748), .B(n14745), .Z(n14746) );
  IV U14580 ( .A(n14713), .Z(n14710) );
  XOR U14581 ( .A(n14749), .B(n14750), .Z(n14713) );
  ANDN U14582 ( .B(n14751), .A(n14752), .Z(n14749) );
  XOR U14583 ( .A(n14750), .B(n14753), .Z(n14751) );
  XOR U14584 ( .A(n14754), .B(n14755), .Z(n14726) );
  XNOR U14585 ( .A(n14721), .B(n14756), .Z(n14755) );
  IV U14586 ( .A(n14724), .Z(n14756) );
  XOR U14587 ( .A(n14757), .B(n14758), .Z(n14724) );
  ANDN U14588 ( .B(n14759), .A(n14760), .Z(n14757) );
  XOR U14589 ( .A(n14758), .B(n14761), .Z(n14759) );
  XNOR U14590 ( .A(n14762), .B(n14763), .Z(n14721) );
  ANDN U14591 ( .B(n14764), .A(n14765), .Z(n14762) );
  XOR U14592 ( .A(n14763), .B(n14766), .Z(n14764) );
  IV U14593 ( .A(n14720), .Z(n14754) );
  XOR U14594 ( .A(n14718), .B(n14767), .Z(n14720) );
  XOR U14595 ( .A(n14768), .B(n14769), .Z(n14767) );
  ANDN U14596 ( .B(n14770), .A(n14771), .Z(n14768) );
  XOR U14597 ( .A(n14772), .B(n14769), .Z(n14770) );
  IV U14598 ( .A(n14722), .Z(n14718) );
  XOR U14599 ( .A(n14773), .B(n14774), .Z(n14722) );
  ANDN U14600 ( .B(n14775), .A(n14776), .Z(n14773) );
  XOR U14601 ( .A(n14777), .B(n14774), .Z(n14775) );
  IV U14602 ( .A(n14732), .Z(n14736) );
  XOR U14603 ( .A(n14732), .B(n14687), .Z(n14734) );
  XOR U14604 ( .A(n14778), .B(n14779), .Z(n14687) );
  AND U14605 ( .A(n382), .B(n14780), .Z(n14778) );
  XOR U14606 ( .A(n14781), .B(n14779), .Z(n14780) );
  NANDN U14607 ( .A(n14689), .B(n14691), .Z(n14732) );
  XOR U14608 ( .A(n14782), .B(n14783), .Z(n14691) );
  AND U14609 ( .A(n382), .B(n14784), .Z(n14782) );
  XOR U14610 ( .A(n14783), .B(n14785), .Z(n14784) );
  XNOR U14611 ( .A(n14786), .B(n14787), .Z(n382) );
  AND U14612 ( .A(n14788), .B(n14789), .Z(n14786) );
  XOR U14613 ( .A(n14787), .B(n14702), .Z(n14789) );
  XNOR U14614 ( .A(n14790), .B(n14791), .Z(n14702) );
  ANDN U14615 ( .B(n14792), .A(n14793), .Z(n14790) );
  XOR U14616 ( .A(n14791), .B(n14794), .Z(n14792) );
  XNOR U14617 ( .A(n14787), .B(n14704), .Z(n14788) );
  XOR U14618 ( .A(n14795), .B(n14796), .Z(n14704) );
  AND U14619 ( .A(n386), .B(n14797), .Z(n14795) );
  XOR U14620 ( .A(n14798), .B(n14796), .Z(n14797) );
  XNOR U14621 ( .A(n14799), .B(n14800), .Z(n14787) );
  AND U14622 ( .A(n14801), .B(n14802), .Z(n14799) );
  XNOR U14623 ( .A(n14800), .B(n14729), .Z(n14802) );
  XOR U14624 ( .A(n14793), .B(n14794), .Z(n14729) );
  XNOR U14625 ( .A(n14803), .B(n14804), .Z(n14794) );
  ANDN U14626 ( .B(n14805), .A(n14806), .Z(n14803) );
  XOR U14627 ( .A(n14807), .B(n14808), .Z(n14805) );
  XOR U14628 ( .A(n14809), .B(n14810), .Z(n14793) );
  XNOR U14629 ( .A(n14811), .B(n14812), .Z(n14810) );
  ANDN U14630 ( .B(n14813), .A(n14814), .Z(n14811) );
  XNOR U14631 ( .A(n14815), .B(n14816), .Z(n14813) );
  IV U14632 ( .A(n14791), .Z(n14809) );
  XOR U14633 ( .A(n14817), .B(n14818), .Z(n14791) );
  ANDN U14634 ( .B(n14819), .A(n14820), .Z(n14817) );
  XOR U14635 ( .A(n14818), .B(n14821), .Z(n14819) );
  XOR U14636 ( .A(n14800), .B(n14731), .Z(n14801) );
  XOR U14637 ( .A(n14822), .B(n14823), .Z(n14731) );
  AND U14638 ( .A(n386), .B(n14824), .Z(n14822) );
  XOR U14639 ( .A(n14825), .B(n14823), .Z(n14824) );
  XNOR U14640 ( .A(n14826), .B(n14827), .Z(n14800) );
  NAND U14641 ( .A(n14828), .B(n14829), .Z(n14827) );
  XOR U14642 ( .A(n14830), .B(n14779), .Z(n14829) );
  XOR U14643 ( .A(n14820), .B(n14821), .Z(n14779) );
  XOR U14644 ( .A(n14831), .B(n14808), .Z(n14821) );
  XOR U14645 ( .A(n14832), .B(n14833), .Z(n14808) );
  ANDN U14646 ( .B(n14834), .A(n14835), .Z(n14832) );
  XOR U14647 ( .A(n14833), .B(n14836), .Z(n14834) );
  IV U14648 ( .A(n14806), .Z(n14831) );
  XOR U14649 ( .A(n14804), .B(n14837), .Z(n14806) );
  XOR U14650 ( .A(n14838), .B(n14839), .Z(n14837) );
  ANDN U14651 ( .B(n14840), .A(n14841), .Z(n14838) );
  XOR U14652 ( .A(n14842), .B(n14839), .Z(n14840) );
  IV U14653 ( .A(n14807), .Z(n14804) );
  XOR U14654 ( .A(n14843), .B(n14844), .Z(n14807) );
  ANDN U14655 ( .B(n14845), .A(n14846), .Z(n14843) );
  XOR U14656 ( .A(n14844), .B(n14847), .Z(n14845) );
  XOR U14657 ( .A(n14848), .B(n14849), .Z(n14820) );
  XNOR U14658 ( .A(n14815), .B(n14850), .Z(n14849) );
  IV U14659 ( .A(n14818), .Z(n14850) );
  XOR U14660 ( .A(n14851), .B(n14852), .Z(n14818) );
  ANDN U14661 ( .B(n14853), .A(n14854), .Z(n14851) );
  XOR U14662 ( .A(n14852), .B(n14855), .Z(n14853) );
  XNOR U14663 ( .A(n14856), .B(n14857), .Z(n14815) );
  ANDN U14664 ( .B(n14858), .A(n14859), .Z(n14856) );
  XOR U14665 ( .A(n14857), .B(n14860), .Z(n14858) );
  IV U14666 ( .A(n14814), .Z(n14848) );
  XOR U14667 ( .A(n14812), .B(n14861), .Z(n14814) );
  XOR U14668 ( .A(n14862), .B(n14863), .Z(n14861) );
  ANDN U14669 ( .B(n14864), .A(n14865), .Z(n14862) );
  XOR U14670 ( .A(n14866), .B(n14863), .Z(n14864) );
  IV U14671 ( .A(n14816), .Z(n14812) );
  XOR U14672 ( .A(n14867), .B(n14868), .Z(n14816) );
  ANDN U14673 ( .B(n14869), .A(n14870), .Z(n14867) );
  XOR U14674 ( .A(n14871), .B(n14868), .Z(n14869) );
  IV U14675 ( .A(n14826), .Z(n14830) );
  XOR U14676 ( .A(n14826), .B(n14781), .Z(n14828) );
  XOR U14677 ( .A(n14872), .B(n14873), .Z(n14781) );
  AND U14678 ( .A(n386), .B(n14874), .Z(n14872) );
  XOR U14679 ( .A(n14875), .B(n14873), .Z(n14874) );
  NANDN U14680 ( .A(n14783), .B(n14785), .Z(n14826) );
  XOR U14681 ( .A(n14876), .B(n14877), .Z(n14785) );
  AND U14682 ( .A(n386), .B(n14878), .Z(n14876) );
  XOR U14683 ( .A(n14877), .B(n14879), .Z(n14878) );
  XNOR U14684 ( .A(n14880), .B(n14881), .Z(n386) );
  AND U14685 ( .A(n14882), .B(n14883), .Z(n14880) );
  XOR U14686 ( .A(n14881), .B(n14796), .Z(n14883) );
  XNOR U14687 ( .A(n14884), .B(n14885), .Z(n14796) );
  ANDN U14688 ( .B(n14886), .A(n14887), .Z(n14884) );
  XOR U14689 ( .A(n14885), .B(n14888), .Z(n14886) );
  XNOR U14690 ( .A(n14881), .B(n14798), .Z(n14882) );
  XOR U14691 ( .A(n14889), .B(n14890), .Z(n14798) );
  AND U14692 ( .A(n390), .B(n14891), .Z(n14889) );
  XOR U14693 ( .A(n14892), .B(n14890), .Z(n14891) );
  XNOR U14694 ( .A(n14893), .B(n14894), .Z(n14881) );
  AND U14695 ( .A(n14895), .B(n14896), .Z(n14893) );
  XNOR U14696 ( .A(n14894), .B(n14823), .Z(n14896) );
  XOR U14697 ( .A(n14887), .B(n14888), .Z(n14823) );
  XNOR U14698 ( .A(n14897), .B(n14898), .Z(n14888) );
  ANDN U14699 ( .B(n14899), .A(n14900), .Z(n14897) );
  XOR U14700 ( .A(n14901), .B(n14902), .Z(n14899) );
  XOR U14701 ( .A(n14903), .B(n14904), .Z(n14887) );
  XNOR U14702 ( .A(n14905), .B(n14906), .Z(n14904) );
  ANDN U14703 ( .B(n14907), .A(n14908), .Z(n14905) );
  XNOR U14704 ( .A(n14909), .B(n14910), .Z(n14907) );
  IV U14705 ( .A(n14885), .Z(n14903) );
  XOR U14706 ( .A(n14911), .B(n14912), .Z(n14885) );
  ANDN U14707 ( .B(n14913), .A(n14914), .Z(n14911) );
  XOR U14708 ( .A(n14912), .B(n14915), .Z(n14913) );
  XOR U14709 ( .A(n14894), .B(n14825), .Z(n14895) );
  XOR U14710 ( .A(n14916), .B(n14917), .Z(n14825) );
  AND U14711 ( .A(n390), .B(n14918), .Z(n14916) );
  XOR U14712 ( .A(n14919), .B(n14917), .Z(n14918) );
  XNOR U14713 ( .A(n14920), .B(n14921), .Z(n14894) );
  NAND U14714 ( .A(n14922), .B(n14923), .Z(n14921) );
  XOR U14715 ( .A(n14924), .B(n14873), .Z(n14923) );
  XOR U14716 ( .A(n14914), .B(n14915), .Z(n14873) );
  XOR U14717 ( .A(n14925), .B(n14902), .Z(n14915) );
  XOR U14718 ( .A(n14926), .B(n14927), .Z(n14902) );
  ANDN U14719 ( .B(n14928), .A(n14929), .Z(n14926) );
  XOR U14720 ( .A(n14927), .B(n14930), .Z(n14928) );
  IV U14721 ( .A(n14900), .Z(n14925) );
  XOR U14722 ( .A(n14898), .B(n14931), .Z(n14900) );
  XOR U14723 ( .A(n14932), .B(n14933), .Z(n14931) );
  ANDN U14724 ( .B(n14934), .A(n14935), .Z(n14932) );
  XOR U14725 ( .A(n14936), .B(n14933), .Z(n14934) );
  IV U14726 ( .A(n14901), .Z(n14898) );
  XOR U14727 ( .A(n14937), .B(n14938), .Z(n14901) );
  ANDN U14728 ( .B(n14939), .A(n14940), .Z(n14937) );
  XOR U14729 ( .A(n14938), .B(n14941), .Z(n14939) );
  XOR U14730 ( .A(n14942), .B(n14943), .Z(n14914) );
  XNOR U14731 ( .A(n14909), .B(n14944), .Z(n14943) );
  IV U14732 ( .A(n14912), .Z(n14944) );
  XOR U14733 ( .A(n14945), .B(n14946), .Z(n14912) );
  ANDN U14734 ( .B(n14947), .A(n14948), .Z(n14945) );
  XOR U14735 ( .A(n14946), .B(n14949), .Z(n14947) );
  XNOR U14736 ( .A(n14950), .B(n14951), .Z(n14909) );
  ANDN U14737 ( .B(n14952), .A(n14953), .Z(n14950) );
  XOR U14738 ( .A(n14951), .B(n14954), .Z(n14952) );
  IV U14739 ( .A(n14908), .Z(n14942) );
  XOR U14740 ( .A(n14906), .B(n14955), .Z(n14908) );
  XOR U14741 ( .A(n14956), .B(n14957), .Z(n14955) );
  ANDN U14742 ( .B(n14958), .A(n14959), .Z(n14956) );
  XOR U14743 ( .A(n14960), .B(n14957), .Z(n14958) );
  IV U14744 ( .A(n14910), .Z(n14906) );
  XOR U14745 ( .A(n14961), .B(n14962), .Z(n14910) );
  ANDN U14746 ( .B(n14963), .A(n14964), .Z(n14961) );
  XOR U14747 ( .A(n14965), .B(n14962), .Z(n14963) );
  IV U14748 ( .A(n14920), .Z(n14924) );
  XOR U14749 ( .A(n14920), .B(n14875), .Z(n14922) );
  XOR U14750 ( .A(n14966), .B(n14967), .Z(n14875) );
  AND U14751 ( .A(n390), .B(n14968), .Z(n14966) );
  XOR U14752 ( .A(n14969), .B(n14967), .Z(n14968) );
  NANDN U14753 ( .A(n14877), .B(n14879), .Z(n14920) );
  XOR U14754 ( .A(n14970), .B(n14971), .Z(n14879) );
  AND U14755 ( .A(n390), .B(n14972), .Z(n14970) );
  XOR U14756 ( .A(n14971), .B(n14973), .Z(n14972) );
  XNOR U14757 ( .A(n14974), .B(n14975), .Z(n390) );
  AND U14758 ( .A(n14976), .B(n14977), .Z(n14974) );
  XOR U14759 ( .A(n14975), .B(n14890), .Z(n14977) );
  XNOR U14760 ( .A(n14978), .B(n14979), .Z(n14890) );
  ANDN U14761 ( .B(n14980), .A(n14981), .Z(n14978) );
  XOR U14762 ( .A(n14979), .B(n14982), .Z(n14980) );
  XNOR U14763 ( .A(n14975), .B(n14892), .Z(n14976) );
  XOR U14764 ( .A(n14983), .B(n14984), .Z(n14892) );
  AND U14765 ( .A(n394), .B(n14985), .Z(n14983) );
  XOR U14766 ( .A(n14986), .B(n14984), .Z(n14985) );
  XNOR U14767 ( .A(n14987), .B(n14988), .Z(n14975) );
  AND U14768 ( .A(n14989), .B(n14990), .Z(n14987) );
  XNOR U14769 ( .A(n14988), .B(n14917), .Z(n14990) );
  XOR U14770 ( .A(n14981), .B(n14982), .Z(n14917) );
  XNOR U14771 ( .A(n14991), .B(n14992), .Z(n14982) );
  ANDN U14772 ( .B(n14993), .A(n14994), .Z(n14991) );
  XOR U14773 ( .A(n14995), .B(n14996), .Z(n14993) );
  XOR U14774 ( .A(n14997), .B(n14998), .Z(n14981) );
  XNOR U14775 ( .A(n14999), .B(n15000), .Z(n14998) );
  ANDN U14776 ( .B(n15001), .A(n15002), .Z(n14999) );
  XNOR U14777 ( .A(n15003), .B(n15004), .Z(n15001) );
  IV U14778 ( .A(n14979), .Z(n14997) );
  XOR U14779 ( .A(n15005), .B(n15006), .Z(n14979) );
  ANDN U14780 ( .B(n15007), .A(n15008), .Z(n15005) );
  XOR U14781 ( .A(n15006), .B(n15009), .Z(n15007) );
  XOR U14782 ( .A(n14988), .B(n14919), .Z(n14989) );
  XOR U14783 ( .A(n15010), .B(n15011), .Z(n14919) );
  AND U14784 ( .A(n394), .B(n15012), .Z(n15010) );
  XOR U14785 ( .A(n15013), .B(n15011), .Z(n15012) );
  XNOR U14786 ( .A(n15014), .B(n15015), .Z(n14988) );
  NAND U14787 ( .A(n15016), .B(n15017), .Z(n15015) );
  XOR U14788 ( .A(n15018), .B(n14967), .Z(n15017) );
  XOR U14789 ( .A(n15008), .B(n15009), .Z(n14967) );
  XOR U14790 ( .A(n15019), .B(n14996), .Z(n15009) );
  XOR U14791 ( .A(n15020), .B(n15021), .Z(n14996) );
  ANDN U14792 ( .B(n15022), .A(n15023), .Z(n15020) );
  XOR U14793 ( .A(n15021), .B(n15024), .Z(n15022) );
  IV U14794 ( .A(n14994), .Z(n15019) );
  XOR U14795 ( .A(n14992), .B(n15025), .Z(n14994) );
  XOR U14796 ( .A(n15026), .B(n15027), .Z(n15025) );
  ANDN U14797 ( .B(n15028), .A(n15029), .Z(n15026) );
  XOR U14798 ( .A(n15030), .B(n15027), .Z(n15028) );
  IV U14799 ( .A(n14995), .Z(n14992) );
  XOR U14800 ( .A(n15031), .B(n15032), .Z(n14995) );
  ANDN U14801 ( .B(n15033), .A(n15034), .Z(n15031) );
  XOR U14802 ( .A(n15032), .B(n15035), .Z(n15033) );
  XOR U14803 ( .A(n15036), .B(n15037), .Z(n15008) );
  XNOR U14804 ( .A(n15003), .B(n15038), .Z(n15037) );
  IV U14805 ( .A(n15006), .Z(n15038) );
  XOR U14806 ( .A(n15039), .B(n15040), .Z(n15006) );
  ANDN U14807 ( .B(n15041), .A(n15042), .Z(n15039) );
  XOR U14808 ( .A(n15040), .B(n15043), .Z(n15041) );
  XNOR U14809 ( .A(n15044), .B(n15045), .Z(n15003) );
  ANDN U14810 ( .B(n15046), .A(n15047), .Z(n15044) );
  XOR U14811 ( .A(n15045), .B(n15048), .Z(n15046) );
  IV U14812 ( .A(n15002), .Z(n15036) );
  XOR U14813 ( .A(n15000), .B(n15049), .Z(n15002) );
  XOR U14814 ( .A(n15050), .B(n15051), .Z(n15049) );
  ANDN U14815 ( .B(n15052), .A(n15053), .Z(n15050) );
  XOR U14816 ( .A(n15054), .B(n15051), .Z(n15052) );
  IV U14817 ( .A(n15004), .Z(n15000) );
  XOR U14818 ( .A(n15055), .B(n15056), .Z(n15004) );
  ANDN U14819 ( .B(n15057), .A(n15058), .Z(n15055) );
  XOR U14820 ( .A(n15059), .B(n15056), .Z(n15057) );
  IV U14821 ( .A(n15014), .Z(n15018) );
  XOR U14822 ( .A(n15014), .B(n14969), .Z(n15016) );
  XOR U14823 ( .A(n15060), .B(n15061), .Z(n14969) );
  AND U14824 ( .A(n394), .B(n15062), .Z(n15060) );
  XOR U14825 ( .A(n15063), .B(n15061), .Z(n15062) );
  NANDN U14826 ( .A(n14971), .B(n14973), .Z(n15014) );
  XOR U14827 ( .A(n15064), .B(n15065), .Z(n14973) );
  AND U14828 ( .A(n394), .B(n15066), .Z(n15064) );
  XOR U14829 ( .A(n15065), .B(n15067), .Z(n15066) );
  XNOR U14830 ( .A(n15068), .B(n15069), .Z(n394) );
  AND U14831 ( .A(n15070), .B(n15071), .Z(n15068) );
  XOR U14832 ( .A(n15069), .B(n14984), .Z(n15071) );
  XNOR U14833 ( .A(n15072), .B(n15073), .Z(n14984) );
  ANDN U14834 ( .B(n15074), .A(n15075), .Z(n15072) );
  XOR U14835 ( .A(n15073), .B(n15076), .Z(n15074) );
  XNOR U14836 ( .A(n15069), .B(n14986), .Z(n15070) );
  XOR U14837 ( .A(n15077), .B(n15078), .Z(n14986) );
  AND U14838 ( .A(n398), .B(n15079), .Z(n15077) );
  XOR U14839 ( .A(n15080), .B(n15078), .Z(n15079) );
  XNOR U14840 ( .A(n15081), .B(n15082), .Z(n15069) );
  AND U14841 ( .A(n15083), .B(n15084), .Z(n15081) );
  XNOR U14842 ( .A(n15082), .B(n15011), .Z(n15084) );
  XOR U14843 ( .A(n15075), .B(n15076), .Z(n15011) );
  XNOR U14844 ( .A(n15085), .B(n15086), .Z(n15076) );
  ANDN U14845 ( .B(n15087), .A(n15088), .Z(n15085) );
  XOR U14846 ( .A(n15089), .B(n15090), .Z(n15087) );
  XOR U14847 ( .A(n15091), .B(n15092), .Z(n15075) );
  XNOR U14848 ( .A(n15093), .B(n15094), .Z(n15092) );
  ANDN U14849 ( .B(n15095), .A(n15096), .Z(n15093) );
  XNOR U14850 ( .A(n15097), .B(n15098), .Z(n15095) );
  IV U14851 ( .A(n15073), .Z(n15091) );
  XOR U14852 ( .A(n15099), .B(n15100), .Z(n15073) );
  ANDN U14853 ( .B(n15101), .A(n15102), .Z(n15099) );
  XOR U14854 ( .A(n15100), .B(n15103), .Z(n15101) );
  XOR U14855 ( .A(n15082), .B(n15013), .Z(n15083) );
  XOR U14856 ( .A(n15104), .B(n15105), .Z(n15013) );
  AND U14857 ( .A(n398), .B(n15106), .Z(n15104) );
  XOR U14858 ( .A(n15107), .B(n15105), .Z(n15106) );
  XNOR U14859 ( .A(n15108), .B(n15109), .Z(n15082) );
  NAND U14860 ( .A(n15110), .B(n15111), .Z(n15109) );
  XOR U14861 ( .A(n15112), .B(n15061), .Z(n15111) );
  XOR U14862 ( .A(n15102), .B(n15103), .Z(n15061) );
  XOR U14863 ( .A(n15113), .B(n15090), .Z(n15103) );
  XOR U14864 ( .A(n15114), .B(n15115), .Z(n15090) );
  ANDN U14865 ( .B(n15116), .A(n15117), .Z(n15114) );
  XOR U14866 ( .A(n15115), .B(n15118), .Z(n15116) );
  IV U14867 ( .A(n15088), .Z(n15113) );
  XOR U14868 ( .A(n15086), .B(n15119), .Z(n15088) );
  XOR U14869 ( .A(n15120), .B(n15121), .Z(n15119) );
  ANDN U14870 ( .B(n15122), .A(n15123), .Z(n15120) );
  XOR U14871 ( .A(n15124), .B(n15121), .Z(n15122) );
  IV U14872 ( .A(n15089), .Z(n15086) );
  XOR U14873 ( .A(n15125), .B(n15126), .Z(n15089) );
  ANDN U14874 ( .B(n15127), .A(n15128), .Z(n15125) );
  XOR U14875 ( .A(n15126), .B(n15129), .Z(n15127) );
  XOR U14876 ( .A(n15130), .B(n15131), .Z(n15102) );
  XNOR U14877 ( .A(n15097), .B(n15132), .Z(n15131) );
  IV U14878 ( .A(n15100), .Z(n15132) );
  XOR U14879 ( .A(n15133), .B(n15134), .Z(n15100) );
  ANDN U14880 ( .B(n15135), .A(n15136), .Z(n15133) );
  XOR U14881 ( .A(n15134), .B(n15137), .Z(n15135) );
  XNOR U14882 ( .A(n15138), .B(n15139), .Z(n15097) );
  ANDN U14883 ( .B(n15140), .A(n15141), .Z(n15138) );
  XOR U14884 ( .A(n15139), .B(n15142), .Z(n15140) );
  IV U14885 ( .A(n15096), .Z(n15130) );
  XOR U14886 ( .A(n15094), .B(n15143), .Z(n15096) );
  XOR U14887 ( .A(n15144), .B(n15145), .Z(n15143) );
  ANDN U14888 ( .B(n15146), .A(n15147), .Z(n15144) );
  XOR U14889 ( .A(n15148), .B(n15145), .Z(n15146) );
  IV U14890 ( .A(n15098), .Z(n15094) );
  XOR U14891 ( .A(n15149), .B(n15150), .Z(n15098) );
  ANDN U14892 ( .B(n15151), .A(n15152), .Z(n15149) );
  XOR U14893 ( .A(n15153), .B(n15150), .Z(n15151) );
  IV U14894 ( .A(n15108), .Z(n15112) );
  XOR U14895 ( .A(n15108), .B(n15063), .Z(n15110) );
  XOR U14896 ( .A(n15154), .B(n15155), .Z(n15063) );
  AND U14897 ( .A(n398), .B(n15156), .Z(n15154) );
  XOR U14898 ( .A(n15157), .B(n15155), .Z(n15156) );
  NANDN U14899 ( .A(n15065), .B(n15067), .Z(n15108) );
  XOR U14900 ( .A(n15158), .B(n15159), .Z(n15067) );
  AND U14901 ( .A(n398), .B(n15160), .Z(n15158) );
  XOR U14902 ( .A(n15159), .B(n15161), .Z(n15160) );
  XNOR U14903 ( .A(n15162), .B(n15163), .Z(n398) );
  AND U14904 ( .A(n15164), .B(n15165), .Z(n15162) );
  XOR U14905 ( .A(n15163), .B(n15078), .Z(n15165) );
  XNOR U14906 ( .A(n15166), .B(n15167), .Z(n15078) );
  ANDN U14907 ( .B(n15168), .A(n15169), .Z(n15166) );
  XOR U14908 ( .A(n15167), .B(n15170), .Z(n15168) );
  XNOR U14909 ( .A(n15163), .B(n15080), .Z(n15164) );
  XOR U14910 ( .A(n15171), .B(n15172), .Z(n15080) );
  AND U14911 ( .A(n402), .B(n15173), .Z(n15171) );
  XOR U14912 ( .A(n15174), .B(n15172), .Z(n15173) );
  XNOR U14913 ( .A(n15175), .B(n15176), .Z(n15163) );
  AND U14914 ( .A(n15177), .B(n15178), .Z(n15175) );
  XNOR U14915 ( .A(n15176), .B(n15105), .Z(n15178) );
  XOR U14916 ( .A(n15169), .B(n15170), .Z(n15105) );
  XNOR U14917 ( .A(n15179), .B(n15180), .Z(n15170) );
  ANDN U14918 ( .B(n15181), .A(n15182), .Z(n15179) );
  XOR U14919 ( .A(n15183), .B(n15184), .Z(n15181) );
  XOR U14920 ( .A(n15185), .B(n15186), .Z(n15169) );
  XNOR U14921 ( .A(n15187), .B(n15188), .Z(n15186) );
  ANDN U14922 ( .B(n15189), .A(n15190), .Z(n15187) );
  XNOR U14923 ( .A(n15191), .B(n15192), .Z(n15189) );
  IV U14924 ( .A(n15167), .Z(n15185) );
  XOR U14925 ( .A(n15193), .B(n15194), .Z(n15167) );
  ANDN U14926 ( .B(n15195), .A(n15196), .Z(n15193) );
  XOR U14927 ( .A(n15194), .B(n15197), .Z(n15195) );
  XOR U14928 ( .A(n15176), .B(n15107), .Z(n15177) );
  XOR U14929 ( .A(n15198), .B(n15199), .Z(n15107) );
  AND U14930 ( .A(n402), .B(n15200), .Z(n15198) );
  XOR U14931 ( .A(n15201), .B(n15199), .Z(n15200) );
  XNOR U14932 ( .A(n15202), .B(n15203), .Z(n15176) );
  NAND U14933 ( .A(n15204), .B(n15205), .Z(n15203) );
  XOR U14934 ( .A(n15206), .B(n15155), .Z(n15205) );
  XOR U14935 ( .A(n15196), .B(n15197), .Z(n15155) );
  XOR U14936 ( .A(n15207), .B(n15184), .Z(n15197) );
  XOR U14937 ( .A(n15208), .B(n15209), .Z(n15184) );
  ANDN U14938 ( .B(n15210), .A(n15211), .Z(n15208) );
  XOR U14939 ( .A(n15209), .B(n15212), .Z(n15210) );
  IV U14940 ( .A(n15182), .Z(n15207) );
  XOR U14941 ( .A(n15180), .B(n15213), .Z(n15182) );
  XOR U14942 ( .A(n15214), .B(n15215), .Z(n15213) );
  ANDN U14943 ( .B(n15216), .A(n15217), .Z(n15214) );
  XOR U14944 ( .A(n15218), .B(n15215), .Z(n15216) );
  IV U14945 ( .A(n15183), .Z(n15180) );
  XOR U14946 ( .A(n15219), .B(n15220), .Z(n15183) );
  ANDN U14947 ( .B(n15221), .A(n15222), .Z(n15219) );
  XOR U14948 ( .A(n15220), .B(n15223), .Z(n15221) );
  XOR U14949 ( .A(n15224), .B(n15225), .Z(n15196) );
  XNOR U14950 ( .A(n15191), .B(n15226), .Z(n15225) );
  IV U14951 ( .A(n15194), .Z(n15226) );
  XOR U14952 ( .A(n15227), .B(n15228), .Z(n15194) );
  ANDN U14953 ( .B(n15229), .A(n15230), .Z(n15227) );
  XOR U14954 ( .A(n15228), .B(n15231), .Z(n15229) );
  XNOR U14955 ( .A(n15232), .B(n15233), .Z(n15191) );
  ANDN U14956 ( .B(n15234), .A(n15235), .Z(n15232) );
  XOR U14957 ( .A(n15233), .B(n15236), .Z(n15234) );
  IV U14958 ( .A(n15190), .Z(n15224) );
  XOR U14959 ( .A(n15188), .B(n15237), .Z(n15190) );
  XOR U14960 ( .A(n15238), .B(n15239), .Z(n15237) );
  ANDN U14961 ( .B(n15240), .A(n15241), .Z(n15238) );
  XOR U14962 ( .A(n15242), .B(n15239), .Z(n15240) );
  IV U14963 ( .A(n15192), .Z(n15188) );
  XOR U14964 ( .A(n15243), .B(n15244), .Z(n15192) );
  ANDN U14965 ( .B(n15245), .A(n15246), .Z(n15243) );
  XOR U14966 ( .A(n15247), .B(n15244), .Z(n15245) );
  IV U14967 ( .A(n15202), .Z(n15206) );
  XOR U14968 ( .A(n15202), .B(n15157), .Z(n15204) );
  XOR U14969 ( .A(n15248), .B(n15249), .Z(n15157) );
  AND U14970 ( .A(n402), .B(n15250), .Z(n15248) );
  XOR U14971 ( .A(n15251), .B(n15249), .Z(n15250) );
  NANDN U14972 ( .A(n15159), .B(n15161), .Z(n15202) );
  XOR U14973 ( .A(n15252), .B(n15253), .Z(n15161) );
  AND U14974 ( .A(n402), .B(n15254), .Z(n15252) );
  XOR U14975 ( .A(n15253), .B(n15255), .Z(n15254) );
  XNOR U14976 ( .A(n15256), .B(n15257), .Z(n402) );
  AND U14977 ( .A(n15258), .B(n15259), .Z(n15256) );
  XOR U14978 ( .A(n15257), .B(n15172), .Z(n15259) );
  XNOR U14979 ( .A(n15260), .B(n15261), .Z(n15172) );
  ANDN U14980 ( .B(n15262), .A(n15263), .Z(n15260) );
  XOR U14981 ( .A(n15261), .B(n15264), .Z(n15262) );
  XNOR U14982 ( .A(n15257), .B(n15174), .Z(n15258) );
  XOR U14983 ( .A(n15265), .B(n15266), .Z(n15174) );
  AND U14984 ( .A(n406), .B(n15267), .Z(n15265) );
  XOR U14985 ( .A(n15268), .B(n15266), .Z(n15267) );
  XNOR U14986 ( .A(n15269), .B(n15270), .Z(n15257) );
  AND U14987 ( .A(n15271), .B(n15272), .Z(n15269) );
  XNOR U14988 ( .A(n15270), .B(n15199), .Z(n15272) );
  XOR U14989 ( .A(n15263), .B(n15264), .Z(n15199) );
  XNOR U14990 ( .A(n15273), .B(n15274), .Z(n15264) );
  ANDN U14991 ( .B(n15275), .A(n15276), .Z(n15273) );
  XOR U14992 ( .A(n15277), .B(n15278), .Z(n15275) );
  XOR U14993 ( .A(n15279), .B(n15280), .Z(n15263) );
  XNOR U14994 ( .A(n15281), .B(n15282), .Z(n15280) );
  ANDN U14995 ( .B(n15283), .A(n15284), .Z(n15281) );
  XNOR U14996 ( .A(n15285), .B(n15286), .Z(n15283) );
  IV U14997 ( .A(n15261), .Z(n15279) );
  XOR U14998 ( .A(n15287), .B(n15288), .Z(n15261) );
  ANDN U14999 ( .B(n15289), .A(n15290), .Z(n15287) );
  XOR U15000 ( .A(n15288), .B(n15291), .Z(n15289) );
  XOR U15001 ( .A(n15270), .B(n15201), .Z(n15271) );
  XOR U15002 ( .A(n15292), .B(n15293), .Z(n15201) );
  AND U15003 ( .A(n406), .B(n15294), .Z(n15292) );
  XOR U15004 ( .A(n15295), .B(n15293), .Z(n15294) );
  XNOR U15005 ( .A(n15296), .B(n15297), .Z(n15270) );
  NAND U15006 ( .A(n15298), .B(n15299), .Z(n15297) );
  XOR U15007 ( .A(n15300), .B(n15249), .Z(n15299) );
  XOR U15008 ( .A(n15290), .B(n15291), .Z(n15249) );
  XOR U15009 ( .A(n15301), .B(n15278), .Z(n15291) );
  XOR U15010 ( .A(n15302), .B(n15303), .Z(n15278) );
  ANDN U15011 ( .B(n15304), .A(n15305), .Z(n15302) );
  XOR U15012 ( .A(n15303), .B(n15306), .Z(n15304) );
  IV U15013 ( .A(n15276), .Z(n15301) );
  XOR U15014 ( .A(n15274), .B(n15307), .Z(n15276) );
  XOR U15015 ( .A(n15308), .B(n15309), .Z(n15307) );
  ANDN U15016 ( .B(n15310), .A(n15311), .Z(n15308) );
  XOR U15017 ( .A(n15312), .B(n15309), .Z(n15310) );
  IV U15018 ( .A(n15277), .Z(n15274) );
  XOR U15019 ( .A(n15313), .B(n15314), .Z(n15277) );
  ANDN U15020 ( .B(n15315), .A(n15316), .Z(n15313) );
  XOR U15021 ( .A(n15314), .B(n15317), .Z(n15315) );
  XOR U15022 ( .A(n15318), .B(n15319), .Z(n15290) );
  XNOR U15023 ( .A(n15285), .B(n15320), .Z(n15319) );
  IV U15024 ( .A(n15288), .Z(n15320) );
  XOR U15025 ( .A(n15321), .B(n15322), .Z(n15288) );
  ANDN U15026 ( .B(n15323), .A(n15324), .Z(n15321) );
  XOR U15027 ( .A(n15322), .B(n15325), .Z(n15323) );
  XNOR U15028 ( .A(n15326), .B(n15327), .Z(n15285) );
  ANDN U15029 ( .B(n15328), .A(n15329), .Z(n15326) );
  XOR U15030 ( .A(n15327), .B(n15330), .Z(n15328) );
  IV U15031 ( .A(n15284), .Z(n15318) );
  XOR U15032 ( .A(n15282), .B(n15331), .Z(n15284) );
  XOR U15033 ( .A(n15332), .B(n15333), .Z(n15331) );
  ANDN U15034 ( .B(n15334), .A(n15335), .Z(n15332) );
  XOR U15035 ( .A(n15336), .B(n15333), .Z(n15334) );
  IV U15036 ( .A(n15286), .Z(n15282) );
  XOR U15037 ( .A(n15337), .B(n15338), .Z(n15286) );
  ANDN U15038 ( .B(n15339), .A(n15340), .Z(n15337) );
  XOR U15039 ( .A(n15341), .B(n15338), .Z(n15339) );
  IV U15040 ( .A(n15296), .Z(n15300) );
  XOR U15041 ( .A(n15296), .B(n15251), .Z(n15298) );
  XOR U15042 ( .A(n15342), .B(n15343), .Z(n15251) );
  AND U15043 ( .A(n406), .B(n15344), .Z(n15342) );
  XOR U15044 ( .A(n15345), .B(n15343), .Z(n15344) );
  NANDN U15045 ( .A(n15253), .B(n15255), .Z(n15296) );
  XOR U15046 ( .A(n15346), .B(n15347), .Z(n15255) );
  AND U15047 ( .A(n406), .B(n15348), .Z(n15346) );
  XOR U15048 ( .A(n15347), .B(n15349), .Z(n15348) );
  XNOR U15049 ( .A(n15350), .B(n15351), .Z(n406) );
  AND U15050 ( .A(n15352), .B(n15353), .Z(n15350) );
  XOR U15051 ( .A(n15351), .B(n15266), .Z(n15353) );
  XNOR U15052 ( .A(n15354), .B(n15355), .Z(n15266) );
  ANDN U15053 ( .B(n15356), .A(n15357), .Z(n15354) );
  XOR U15054 ( .A(n15355), .B(n15358), .Z(n15356) );
  XNOR U15055 ( .A(n15351), .B(n15268), .Z(n15352) );
  XOR U15056 ( .A(n15359), .B(n15360), .Z(n15268) );
  AND U15057 ( .A(n410), .B(n15361), .Z(n15359) );
  XOR U15058 ( .A(n15362), .B(n15360), .Z(n15361) );
  XNOR U15059 ( .A(n15363), .B(n15364), .Z(n15351) );
  AND U15060 ( .A(n15365), .B(n15366), .Z(n15363) );
  XNOR U15061 ( .A(n15364), .B(n15293), .Z(n15366) );
  XOR U15062 ( .A(n15357), .B(n15358), .Z(n15293) );
  XNOR U15063 ( .A(n15367), .B(n15368), .Z(n15358) );
  ANDN U15064 ( .B(n15369), .A(n15370), .Z(n15367) );
  XOR U15065 ( .A(n15371), .B(n15372), .Z(n15369) );
  XOR U15066 ( .A(n15373), .B(n15374), .Z(n15357) );
  XNOR U15067 ( .A(n15375), .B(n15376), .Z(n15374) );
  ANDN U15068 ( .B(n15377), .A(n15378), .Z(n15375) );
  XNOR U15069 ( .A(n15379), .B(n15380), .Z(n15377) );
  IV U15070 ( .A(n15355), .Z(n15373) );
  XOR U15071 ( .A(n15381), .B(n15382), .Z(n15355) );
  ANDN U15072 ( .B(n15383), .A(n15384), .Z(n15381) );
  XOR U15073 ( .A(n15382), .B(n15385), .Z(n15383) );
  XOR U15074 ( .A(n15364), .B(n15295), .Z(n15365) );
  XOR U15075 ( .A(n15386), .B(n15387), .Z(n15295) );
  AND U15076 ( .A(n410), .B(n15388), .Z(n15386) );
  XOR U15077 ( .A(n15389), .B(n15387), .Z(n15388) );
  XNOR U15078 ( .A(n15390), .B(n15391), .Z(n15364) );
  NAND U15079 ( .A(n15392), .B(n15393), .Z(n15391) );
  XOR U15080 ( .A(n15394), .B(n15343), .Z(n15393) );
  XOR U15081 ( .A(n15384), .B(n15385), .Z(n15343) );
  XOR U15082 ( .A(n15395), .B(n15372), .Z(n15385) );
  XOR U15083 ( .A(n15396), .B(n15397), .Z(n15372) );
  ANDN U15084 ( .B(n15398), .A(n15399), .Z(n15396) );
  XOR U15085 ( .A(n15397), .B(n15400), .Z(n15398) );
  IV U15086 ( .A(n15370), .Z(n15395) );
  XOR U15087 ( .A(n15368), .B(n15401), .Z(n15370) );
  XOR U15088 ( .A(n15402), .B(n15403), .Z(n15401) );
  ANDN U15089 ( .B(n15404), .A(n15405), .Z(n15402) );
  XOR U15090 ( .A(n15406), .B(n15403), .Z(n15404) );
  IV U15091 ( .A(n15371), .Z(n15368) );
  XOR U15092 ( .A(n15407), .B(n15408), .Z(n15371) );
  ANDN U15093 ( .B(n15409), .A(n15410), .Z(n15407) );
  XOR U15094 ( .A(n15408), .B(n15411), .Z(n15409) );
  XOR U15095 ( .A(n15412), .B(n15413), .Z(n15384) );
  XNOR U15096 ( .A(n15379), .B(n15414), .Z(n15413) );
  IV U15097 ( .A(n15382), .Z(n15414) );
  XOR U15098 ( .A(n15415), .B(n15416), .Z(n15382) );
  ANDN U15099 ( .B(n15417), .A(n15418), .Z(n15415) );
  XOR U15100 ( .A(n15416), .B(n15419), .Z(n15417) );
  XNOR U15101 ( .A(n15420), .B(n15421), .Z(n15379) );
  ANDN U15102 ( .B(n15422), .A(n15423), .Z(n15420) );
  XOR U15103 ( .A(n15421), .B(n15424), .Z(n15422) );
  IV U15104 ( .A(n15378), .Z(n15412) );
  XOR U15105 ( .A(n15376), .B(n15425), .Z(n15378) );
  XOR U15106 ( .A(n15426), .B(n15427), .Z(n15425) );
  ANDN U15107 ( .B(n15428), .A(n15429), .Z(n15426) );
  XOR U15108 ( .A(n15430), .B(n15427), .Z(n15428) );
  IV U15109 ( .A(n15380), .Z(n15376) );
  XOR U15110 ( .A(n15431), .B(n15432), .Z(n15380) );
  ANDN U15111 ( .B(n15433), .A(n15434), .Z(n15431) );
  XOR U15112 ( .A(n15435), .B(n15432), .Z(n15433) );
  IV U15113 ( .A(n15390), .Z(n15394) );
  XOR U15114 ( .A(n15390), .B(n15345), .Z(n15392) );
  XOR U15115 ( .A(n15436), .B(n15437), .Z(n15345) );
  AND U15116 ( .A(n410), .B(n15438), .Z(n15436) );
  XOR U15117 ( .A(n15439), .B(n15437), .Z(n15438) );
  NANDN U15118 ( .A(n15347), .B(n15349), .Z(n15390) );
  XOR U15119 ( .A(n15440), .B(n15441), .Z(n15349) );
  AND U15120 ( .A(n410), .B(n15442), .Z(n15440) );
  XOR U15121 ( .A(n15441), .B(n15443), .Z(n15442) );
  XNOR U15122 ( .A(n15444), .B(n15445), .Z(n410) );
  AND U15123 ( .A(n15446), .B(n15447), .Z(n15444) );
  XOR U15124 ( .A(n15445), .B(n15360), .Z(n15447) );
  XNOR U15125 ( .A(n15448), .B(n15449), .Z(n15360) );
  ANDN U15126 ( .B(n15450), .A(n15451), .Z(n15448) );
  XOR U15127 ( .A(n15449), .B(n15452), .Z(n15450) );
  XNOR U15128 ( .A(n15445), .B(n15362), .Z(n15446) );
  XOR U15129 ( .A(n15453), .B(n15454), .Z(n15362) );
  AND U15130 ( .A(n414), .B(n15455), .Z(n15453) );
  XOR U15131 ( .A(n15456), .B(n15454), .Z(n15455) );
  XNOR U15132 ( .A(n15457), .B(n15458), .Z(n15445) );
  AND U15133 ( .A(n15459), .B(n15460), .Z(n15457) );
  XNOR U15134 ( .A(n15458), .B(n15387), .Z(n15460) );
  XOR U15135 ( .A(n15451), .B(n15452), .Z(n15387) );
  XNOR U15136 ( .A(n15461), .B(n15462), .Z(n15452) );
  ANDN U15137 ( .B(n15463), .A(n15464), .Z(n15461) );
  XOR U15138 ( .A(n15465), .B(n15466), .Z(n15463) );
  XOR U15139 ( .A(n15467), .B(n15468), .Z(n15451) );
  XNOR U15140 ( .A(n15469), .B(n15470), .Z(n15468) );
  ANDN U15141 ( .B(n15471), .A(n15472), .Z(n15469) );
  XNOR U15142 ( .A(n15473), .B(n15474), .Z(n15471) );
  IV U15143 ( .A(n15449), .Z(n15467) );
  XOR U15144 ( .A(n15475), .B(n15476), .Z(n15449) );
  ANDN U15145 ( .B(n15477), .A(n15478), .Z(n15475) );
  XOR U15146 ( .A(n15476), .B(n15479), .Z(n15477) );
  XOR U15147 ( .A(n15458), .B(n15389), .Z(n15459) );
  XOR U15148 ( .A(n15480), .B(n15481), .Z(n15389) );
  AND U15149 ( .A(n414), .B(n15482), .Z(n15480) );
  XOR U15150 ( .A(n15483), .B(n15481), .Z(n15482) );
  XNOR U15151 ( .A(n15484), .B(n15485), .Z(n15458) );
  NAND U15152 ( .A(n15486), .B(n15487), .Z(n15485) );
  XOR U15153 ( .A(n15488), .B(n15437), .Z(n15487) );
  XOR U15154 ( .A(n15478), .B(n15479), .Z(n15437) );
  XOR U15155 ( .A(n15489), .B(n15466), .Z(n15479) );
  XOR U15156 ( .A(n15490), .B(n15491), .Z(n15466) );
  ANDN U15157 ( .B(n15492), .A(n15493), .Z(n15490) );
  XOR U15158 ( .A(n15491), .B(n15494), .Z(n15492) );
  IV U15159 ( .A(n15464), .Z(n15489) );
  XOR U15160 ( .A(n15462), .B(n15495), .Z(n15464) );
  XOR U15161 ( .A(n15496), .B(n15497), .Z(n15495) );
  ANDN U15162 ( .B(n15498), .A(n15499), .Z(n15496) );
  XOR U15163 ( .A(n15500), .B(n15497), .Z(n15498) );
  IV U15164 ( .A(n15465), .Z(n15462) );
  XOR U15165 ( .A(n15501), .B(n15502), .Z(n15465) );
  ANDN U15166 ( .B(n15503), .A(n15504), .Z(n15501) );
  XOR U15167 ( .A(n15502), .B(n15505), .Z(n15503) );
  XOR U15168 ( .A(n15506), .B(n15507), .Z(n15478) );
  XNOR U15169 ( .A(n15473), .B(n15508), .Z(n15507) );
  IV U15170 ( .A(n15476), .Z(n15508) );
  XOR U15171 ( .A(n15509), .B(n15510), .Z(n15476) );
  ANDN U15172 ( .B(n15511), .A(n15512), .Z(n15509) );
  XOR U15173 ( .A(n15510), .B(n15513), .Z(n15511) );
  XNOR U15174 ( .A(n15514), .B(n15515), .Z(n15473) );
  ANDN U15175 ( .B(n15516), .A(n15517), .Z(n15514) );
  XOR U15176 ( .A(n15515), .B(n15518), .Z(n15516) );
  IV U15177 ( .A(n15472), .Z(n15506) );
  XOR U15178 ( .A(n15470), .B(n15519), .Z(n15472) );
  XOR U15179 ( .A(n15520), .B(n15521), .Z(n15519) );
  ANDN U15180 ( .B(n15522), .A(n15523), .Z(n15520) );
  XOR U15181 ( .A(n15524), .B(n15521), .Z(n15522) );
  IV U15182 ( .A(n15474), .Z(n15470) );
  XOR U15183 ( .A(n15525), .B(n15526), .Z(n15474) );
  ANDN U15184 ( .B(n15527), .A(n15528), .Z(n15525) );
  XOR U15185 ( .A(n15529), .B(n15526), .Z(n15527) );
  IV U15186 ( .A(n15484), .Z(n15488) );
  XOR U15187 ( .A(n15484), .B(n15439), .Z(n15486) );
  XOR U15188 ( .A(n15530), .B(n15531), .Z(n15439) );
  AND U15189 ( .A(n414), .B(n15532), .Z(n15530) );
  XOR U15190 ( .A(n15533), .B(n15531), .Z(n15532) );
  NANDN U15191 ( .A(n15441), .B(n15443), .Z(n15484) );
  XOR U15192 ( .A(n15534), .B(n15535), .Z(n15443) );
  AND U15193 ( .A(n414), .B(n15536), .Z(n15534) );
  XOR U15194 ( .A(n15535), .B(n15537), .Z(n15536) );
  XNOR U15195 ( .A(n15538), .B(n15539), .Z(n414) );
  AND U15196 ( .A(n15540), .B(n15541), .Z(n15538) );
  XOR U15197 ( .A(n15539), .B(n15454), .Z(n15541) );
  XNOR U15198 ( .A(n15542), .B(n15543), .Z(n15454) );
  ANDN U15199 ( .B(n15544), .A(n15545), .Z(n15542) );
  XOR U15200 ( .A(n15543), .B(n15546), .Z(n15544) );
  XNOR U15201 ( .A(n15539), .B(n15456), .Z(n15540) );
  XOR U15202 ( .A(n15547), .B(n15548), .Z(n15456) );
  AND U15203 ( .A(n418), .B(n15549), .Z(n15547) );
  XOR U15204 ( .A(n15550), .B(n15548), .Z(n15549) );
  XNOR U15205 ( .A(n15551), .B(n15552), .Z(n15539) );
  AND U15206 ( .A(n15553), .B(n15554), .Z(n15551) );
  XNOR U15207 ( .A(n15552), .B(n15481), .Z(n15554) );
  XOR U15208 ( .A(n15545), .B(n15546), .Z(n15481) );
  XNOR U15209 ( .A(n15555), .B(n15556), .Z(n15546) );
  ANDN U15210 ( .B(n15557), .A(n15558), .Z(n15555) );
  XOR U15211 ( .A(n15559), .B(n15560), .Z(n15557) );
  XOR U15212 ( .A(n15561), .B(n15562), .Z(n15545) );
  XNOR U15213 ( .A(n15563), .B(n15564), .Z(n15562) );
  ANDN U15214 ( .B(n15565), .A(n15566), .Z(n15563) );
  XNOR U15215 ( .A(n15567), .B(n15568), .Z(n15565) );
  IV U15216 ( .A(n15543), .Z(n15561) );
  XOR U15217 ( .A(n15569), .B(n15570), .Z(n15543) );
  ANDN U15218 ( .B(n15571), .A(n15572), .Z(n15569) );
  XOR U15219 ( .A(n15570), .B(n15573), .Z(n15571) );
  XOR U15220 ( .A(n15552), .B(n15483), .Z(n15553) );
  XOR U15221 ( .A(n15574), .B(n15575), .Z(n15483) );
  AND U15222 ( .A(n418), .B(n15576), .Z(n15574) );
  XOR U15223 ( .A(n15577), .B(n15575), .Z(n15576) );
  XNOR U15224 ( .A(n15578), .B(n15579), .Z(n15552) );
  NAND U15225 ( .A(n15580), .B(n15581), .Z(n15579) );
  XOR U15226 ( .A(n15582), .B(n15531), .Z(n15581) );
  XOR U15227 ( .A(n15572), .B(n15573), .Z(n15531) );
  XOR U15228 ( .A(n15583), .B(n15560), .Z(n15573) );
  XOR U15229 ( .A(n15584), .B(n15585), .Z(n15560) );
  ANDN U15230 ( .B(n15586), .A(n15587), .Z(n15584) );
  XOR U15231 ( .A(n15585), .B(n15588), .Z(n15586) );
  IV U15232 ( .A(n15558), .Z(n15583) );
  XOR U15233 ( .A(n15556), .B(n15589), .Z(n15558) );
  XOR U15234 ( .A(n15590), .B(n15591), .Z(n15589) );
  ANDN U15235 ( .B(n15592), .A(n15593), .Z(n15590) );
  XOR U15236 ( .A(n15594), .B(n15591), .Z(n15592) );
  IV U15237 ( .A(n15559), .Z(n15556) );
  XOR U15238 ( .A(n15595), .B(n15596), .Z(n15559) );
  ANDN U15239 ( .B(n15597), .A(n15598), .Z(n15595) );
  XOR U15240 ( .A(n15596), .B(n15599), .Z(n15597) );
  XOR U15241 ( .A(n15600), .B(n15601), .Z(n15572) );
  XNOR U15242 ( .A(n15567), .B(n15602), .Z(n15601) );
  IV U15243 ( .A(n15570), .Z(n15602) );
  XOR U15244 ( .A(n15603), .B(n15604), .Z(n15570) );
  ANDN U15245 ( .B(n15605), .A(n15606), .Z(n15603) );
  XOR U15246 ( .A(n15604), .B(n15607), .Z(n15605) );
  XNOR U15247 ( .A(n15608), .B(n15609), .Z(n15567) );
  ANDN U15248 ( .B(n15610), .A(n15611), .Z(n15608) );
  XOR U15249 ( .A(n15609), .B(n15612), .Z(n15610) );
  IV U15250 ( .A(n15566), .Z(n15600) );
  XOR U15251 ( .A(n15564), .B(n15613), .Z(n15566) );
  XOR U15252 ( .A(n15614), .B(n15615), .Z(n15613) );
  ANDN U15253 ( .B(n15616), .A(n15617), .Z(n15614) );
  XOR U15254 ( .A(n15618), .B(n15615), .Z(n15616) );
  IV U15255 ( .A(n15568), .Z(n15564) );
  XOR U15256 ( .A(n15619), .B(n15620), .Z(n15568) );
  ANDN U15257 ( .B(n15621), .A(n15622), .Z(n15619) );
  XOR U15258 ( .A(n15623), .B(n15620), .Z(n15621) );
  IV U15259 ( .A(n15578), .Z(n15582) );
  XOR U15260 ( .A(n15578), .B(n15533), .Z(n15580) );
  XOR U15261 ( .A(n15624), .B(n15625), .Z(n15533) );
  AND U15262 ( .A(n418), .B(n15626), .Z(n15624) );
  XOR U15263 ( .A(n15627), .B(n15625), .Z(n15626) );
  NANDN U15264 ( .A(n15535), .B(n15537), .Z(n15578) );
  XOR U15265 ( .A(n15628), .B(n15629), .Z(n15537) );
  AND U15266 ( .A(n418), .B(n15630), .Z(n15628) );
  XOR U15267 ( .A(n15629), .B(n15631), .Z(n15630) );
  XNOR U15268 ( .A(n15632), .B(n15633), .Z(n418) );
  AND U15269 ( .A(n15634), .B(n15635), .Z(n15632) );
  XOR U15270 ( .A(n15633), .B(n15548), .Z(n15635) );
  XNOR U15271 ( .A(n15636), .B(n15637), .Z(n15548) );
  ANDN U15272 ( .B(n15638), .A(n15639), .Z(n15636) );
  XOR U15273 ( .A(n15637), .B(n15640), .Z(n15638) );
  XNOR U15274 ( .A(n15633), .B(n15550), .Z(n15634) );
  XOR U15275 ( .A(n15641), .B(n15642), .Z(n15550) );
  AND U15276 ( .A(n422), .B(n15643), .Z(n15641) );
  XOR U15277 ( .A(n15644), .B(n15642), .Z(n15643) );
  XNOR U15278 ( .A(n15645), .B(n15646), .Z(n15633) );
  AND U15279 ( .A(n15647), .B(n15648), .Z(n15645) );
  XNOR U15280 ( .A(n15646), .B(n15575), .Z(n15648) );
  XOR U15281 ( .A(n15639), .B(n15640), .Z(n15575) );
  XNOR U15282 ( .A(n15649), .B(n15650), .Z(n15640) );
  ANDN U15283 ( .B(n15651), .A(n15652), .Z(n15649) );
  XOR U15284 ( .A(n15653), .B(n15654), .Z(n15651) );
  XOR U15285 ( .A(n15655), .B(n15656), .Z(n15639) );
  XNOR U15286 ( .A(n15657), .B(n15658), .Z(n15656) );
  ANDN U15287 ( .B(n15659), .A(n15660), .Z(n15657) );
  XNOR U15288 ( .A(n15661), .B(n15662), .Z(n15659) );
  IV U15289 ( .A(n15637), .Z(n15655) );
  XOR U15290 ( .A(n15663), .B(n15664), .Z(n15637) );
  ANDN U15291 ( .B(n15665), .A(n15666), .Z(n15663) );
  XOR U15292 ( .A(n15664), .B(n15667), .Z(n15665) );
  XOR U15293 ( .A(n15646), .B(n15577), .Z(n15647) );
  XOR U15294 ( .A(n15668), .B(n15669), .Z(n15577) );
  AND U15295 ( .A(n422), .B(n15670), .Z(n15668) );
  XOR U15296 ( .A(n15671), .B(n15669), .Z(n15670) );
  XNOR U15297 ( .A(n15672), .B(n15673), .Z(n15646) );
  NAND U15298 ( .A(n15674), .B(n15675), .Z(n15673) );
  XOR U15299 ( .A(n15676), .B(n15625), .Z(n15675) );
  XOR U15300 ( .A(n15666), .B(n15667), .Z(n15625) );
  XOR U15301 ( .A(n15677), .B(n15654), .Z(n15667) );
  XOR U15302 ( .A(n15678), .B(n15679), .Z(n15654) );
  ANDN U15303 ( .B(n15680), .A(n15681), .Z(n15678) );
  XOR U15304 ( .A(n15679), .B(n15682), .Z(n15680) );
  IV U15305 ( .A(n15652), .Z(n15677) );
  XOR U15306 ( .A(n15650), .B(n15683), .Z(n15652) );
  XOR U15307 ( .A(n15684), .B(n15685), .Z(n15683) );
  ANDN U15308 ( .B(n15686), .A(n15687), .Z(n15684) );
  XOR U15309 ( .A(n15688), .B(n15685), .Z(n15686) );
  IV U15310 ( .A(n15653), .Z(n15650) );
  XOR U15311 ( .A(n15689), .B(n15690), .Z(n15653) );
  ANDN U15312 ( .B(n15691), .A(n15692), .Z(n15689) );
  XOR U15313 ( .A(n15690), .B(n15693), .Z(n15691) );
  XOR U15314 ( .A(n15694), .B(n15695), .Z(n15666) );
  XNOR U15315 ( .A(n15661), .B(n15696), .Z(n15695) );
  IV U15316 ( .A(n15664), .Z(n15696) );
  XOR U15317 ( .A(n15697), .B(n15698), .Z(n15664) );
  ANDN U15318 ( .B(n15699), .A(n15700), .Z(n15697) );
  XOR U15319 ( .A(n15698), .B(n15701), .Z(n15699) );
  XNOR U15320 ( .A(n15702), .B(n15703), .Z(n15661) );
  ANDN U15321 ( .B(n15704), .A(n15705), .Z(n15702) );
  XOR U15322 ( .A(n15703), .B(n15706), .Z(n15704) );
  IV U15323 ( .A(n15660), .Z(n15694) );
  XOR U15324 ( .A(n15658), .B(n15707), .Z(n15660) );
  XOR U15325 ( .A(n15708), .B(n15709), .Z(n15707) );
  ANDN U15326 ( .B(n15710), .A(n15711), .Z(n15708) );
  XOR U15327 ( .A(n15712), .B(n15709), .Z(n15710) );
  IV U15328 ( .A(n15662), .Z(n15658) );
  XOR U15329 ( .A(n15713), .B(n15714), .Z(n15662) );
  ANDN U15330 ( .B(n15715), .A(n15716), .Z(n15713) );
  XOR U15331 ( .A(n15717), .B(n15714), .Z(n15715) );
  IV U15332 ( .A(n15672), .Z(n15676) );
  XOR U15333 ( .A(n15672), .B(n15627), .Z(n15674) );
  XOR U15334 ( .A(n15718), .B(n15719), .Z(n15627) );
  AND U15335 ( .A(n422), .B(n15720), .Z(n15718) );
  XOR U15336 ( .A(n15721), .B(n15719), .Z(n15720) );
  NANDN U15337 ( .A(n15629), .B(n15631), .Z(n15672) );
  XOR U15338 ( .A(n15722), .B(n15723), .Z(n15631) );
  AND U15339 ( .A(n422), .B(n15724), .Z(n15722) );
  XOR U15340 ( .A(n15723), .B(n15725), .Z(n15724) );
  XNOR U15341 ( .A(n15726), .B(n15727), .Z(n422) );
  AND U15342 ( .A(n15728), .B(n15729), .Z(n15726) );
  XOR U15343 ( .A(n15727), .B(n15642), .Z(n15729) );
  XNOR U15344 ( .A(n15730), .B(n15731), .Z(n15642) );
  ANDN U15345 ( .B(n15732), .A(n15733), .Z(n15730) );
  XOR U15346 ( .A(n15731), .B(n15734), .Z(n15732) );
  XNOR U15347 ( .A(n15727), .B(n15644), .Z(n15728) );
  XOR U15348 ( .A(n15735), .B(n15736), .Z(n15644) );
  AND U15349 ( .A(n426), .B(n15737), .Z(n15735) );
  XOR U15350 ( .A(n15738), .B(n15736), .Z(n15737) );
  XNOR U15351 ( .A(n15739), .B(n15740), .Z(n15727) );
  AND U15352 ( .A(n15741), .B(n15742), .Z(n15739) );
  XNOR U15353 ( .A(n15740), .B(n15669), .Z(n15742) );
  XOR U15354 ( .A(n15733), .B(n15734), .Z(n15669) );
  XNOR U15355 ( .A(n15743), .B(n15744), .Z(n15734) );
  ANDN U15356 ( .B(n15745), .A(n15746), .Z(n15743) );
  XOR U15357 ( .A(n15747), .B(n15748), .Z(n15745) );
  XOR U15358 ( .A(n15749), .B(n15750), .Z(n15733) );
  XNOR U15359 ( .A(n15751), .B(n15752), .Z(n15750) );
  ANDN U15360 ( .B(n15753), .A(n15754), .Z(n15751) );
  XNOR U15361 ( .A(n15755), .B(n15756), .Z(n15753) );
  IV U15362 ( .A(n15731), .Z(n15749) );
  XOR U15363 ( .A(n15757), .B(n15758), .Z(n15731) );
  ANDN U15364 ( .B(n15759), .A(n15760), .Z(n15757) );
  XOR U15365 ( .A(n15758), .B(n15761), .Z(n15759) );
  XOR U15366 ( .A(n15740), .B(n15671), .Z(n15741) );
  XOR U15367 ( .A(n15762), .B(n15763), .Z(n15671) );
  AND U15368 ( .A(n426), .B(n15764), .Z(n15762) );
  XOR U15369 ( .A(n15765), .B(n15763), .Z(n15764) );
  XNOR U15370 ( .A(n15766), .B(n15767), .Z(n15740) );
  NAND U15371 ( .A(n15768), .B(n15769), .Z(n15767) );
  XOR U15372 ( .A(n15770), .B(n15719), .Z(n15769) );
  XOR U15373 ( .A(n15760), .B(n15761), .Z(n15719) );
  XOR U15374 ( .A(n15771), .B(n15748), .Z(n15761) );
  XOR U15375 ( .A(n15772), .B(n15773), .Z(n15748) );
  ANDN U15376 ( .B(n15774), .A(n15775), .Z(n15772) );
  XOR U15377 ( .A(n15773), .B(n15776), .Z(n15774) );
  IV U15378 ( .A(n15746), .Z(n15771) );
  XOR U15379 ( .A(n15744), .B(n15777), .Z(n15746) );
  XOR U15380 ( .A(n15778), .B(n15779), .Z(n15777) );
  ANDN U15381 ( .B(n15780), .A(n15781), .Z(n15778) );
  XOR U15382 ( .A(n15782), .B(n15779), .Z(n15780) );
  IV U15383 ( .A(n15747), .Z(n15744) );
  XOR U15384 ( .A(n15783), .B(n15784), .Z(n15747) );
  ANDN U15385 ( .B(n15785), .A(n15786), .Z(n15783) );
  XOR U15386 ( .A(n15784), .B(n15787), .Z(n15785) );
  XOR U15387 ( .A(n15788), .B(n15789), .Z(n15760) );
  XNOR U15388 ( .A(n15755), .B(n15790), .Z(n15789) );
  IV U15389 ( .A(n15758), .Z(n15790) );
  XOR U15390 ( .A(n15791), .B(n15792), .Z(n15758) );
  ANDN U15391 ( .B(n15793), .A(n15794), .Z(n15791) );
  XOR U15392 ( .A(n15792), .B(n15795), .Z(n15793) );
  XNOR U15393 ( .A(n15796), .B(n15797), .Z(n15755) );
  ANDN U15394 ( .B(n15798), .A(n15799), .Z(n15796) );
  XOR U15395 ( .A(n15797), .B(n15800), .Z(n15798) );
  IV U15396 ( .A(n15754), .Z(n15788) );
  XOR U15397 ( .A(n15752), .B(n15801), .Z(n15754) );
  XOR U15398 ( .A(n15802), .B(n15803), .Z(n15801) );
  ANDN U15399 ( .B(n15804), .A(n15805), .Z(n15802) );
  XOR U15400 ( .A(n15806), .B(n15803), .Z(n15804) );
  IV U15401 ( .A(n15756), .Z(n15752) );
  XOR U15402 ( .A(n15807), .B(n15808), .Z(n15756) );
  ANDN U15403 ( .B(n15809), .A(n15810), .Z(n15807) );
  XOR U15404 ( .A(n15811), .B(n15808), .Z(n15809) );
  IV U15405 ( .A(n15766), .Z(n15770) );
  XOR U15406 ( .A(n15766), .B(n15721), .Z(n15768) );
  XOR U15407 ( .A(n15812), .B(n15813), .Z(n15721) );
  AND U15408 ( .A(n426), .B(n15814), .Z(n15812) );
  XOR U15409 ( .A(n15815), .B(n15813), .Z(n15814) );
  NANDN U15410 ( .A(n15723), .B(n15725), .Z(n15766) );
  XOR U15411 ( .A(n15816), .B(n15817), .Z(n15725) );
  AND U15412 ( .A(n426), .B(n15818), .Z(n15816) );
  XOR U15413 ( .A(n15817), .B(n15819), .Z(n15818) );
  XNOR U15414 ( .A(n15820), .B(n15821), .Z(n426) );
  AND U15415 ( .A(n15822), .B(n15823), .Z(n15820) );
  XOR U15416 ( .A(n15821), .B(n15736), .Z(n15823) );
  XNOR U15417 ( .A(n15824), .B(n15825), .Z(n15736) );
  ANDN U15418 ( .B(n15826), .A(n15827), .Z(n15824) );
  XOR U15419 ( .A(n15825), .B(n15828), .Z(n15826) );
  XNOR U15420 ( .A(n15821), .B(n15738), .Z(n15822) );
  XOR U15421 ( .A(n15829), .B(n15830), .Z(n15738) );
  AND U15422 ( .A(n430), .B(n15831), .Z(n15829) );
  XOR U15423 ( .A(n15832), .B(n15830), .Z(n15831) );
  XNOR U15424 ( .A(n15833), .B(n15834), .Z(n15821) );
  AND U15425 ( .A(n15835), .B(n15836), .Z(n15833) );
  XNOR U15426 ( .A(n15834), .B(n15763), .Z(n15836) );
  XOR U15427 ( .A(n15827), .B(n15828), .Z(n15763) );
  XNOR U15428 ( .A(n15837), .B(n15838), .Z(n15828) );
  ANDN U15429 ( .B(n15839), .A(n15840), .Z(n15837) );
  XOR U15430 ( .A(n15841), .B(n15842), .Z(n15839) );
  XOR U15431 ( .A(n15843), .B(n15844), .Z(n15827) );
  XNOR U15432 ( .A(n15845), .B(n15846), .Z(n15844) );
  ANDN U15433 ( .B(n15847), .A(n15848), .Z(n15845) );
  XNOR U15434 ( .A(n15849), .B(n15850), .Z(n15847) );
  IV U15435 ( .A(n15825), .Z(n15843) );
  XOR U15436 ( .A(n15851), .B(n15852), .Z(n15825) );
  ANDN U15437 ( .B(n15853), .A(n15854), .Z(n15851) );
  XOR U15438 ( .A(n15852), .B(n15855), .Z(n15853) );
  XOR U15439 ( .A(n15834), .B(n15765), .Z(n15835) );
  XOR U15440 ( .A(n15856), .B(n15857), .Z(n15765) );
  AND U15441 ( .A(n430), .B(n15858), .Z(n15856) );
  XOR U15442 ( .A(n15859), .B(n15857), .Z(n15858) );
  XNOR U15443 ( .A(n15860), .B(n15861), .Z(n15834) );
  NAND U15444 ( .A(n15862), .B(n15863), .Z(n15861) );
  XOR U15445 ( .A(n15864), .B(n15813), .Z(n15863) );
  XOR U15446 ( .A(n15854), .B(n15855), .Z(n15813) );
  XOR U15447 ( .A(n15865), .B(n15842), .Z(n15855) );
  XOR U15448 ( .A(n15866), .B(n15867), .Z(n15842) );
  ANDN U15449 ( .B(n15868), .A(n15869), .Z(n15866) );
  XOR U15450 ( .A(n15867), .B(n15870), .Z(n15868) );
  IV U15451 ( .A(n15840), .Z(n15865) );
  XOR U15452 ( .A(n15838), .B(n15871), .Z(n15840) );
  XOR U15453 ( .A(n15872), .B(n15873), .Z(n15871) );
  ANDN U15454 ( .B(n15874), .A(n15875), .Z(n15872) );
  XOR U15455 ( .A(n15876), .B(n15873), .Z(n15874) );
  IV U15456 ( .A(n15841), .Z(n15838) );
  XOR U15457 ( .A(n15877), .B(n15878), .Z(n15841) );
  ANDN U15458 ( .B(n15879), .A(n15880), .Z(n15877) );
  XOR U15459 ( .A(n15878), .B(n15881), .Z(n15879) );
  XOR U15460 ( .A(n15882), .B(n15883), .Z(n15854) );
  XNOR U15461 ( .A(n15849), .B(n15884), .Z(n15883) );
  IV U15462 ( .A(n15852), .Z(n15884) );
  XOR U15463 ( .A(n15885), .B(n15886), .Z(n15852) );
  ANDN U15464 ( .B(n15887), .A(n15888), .Z(n15885) );
  XOR U15465 ( .A(n15886), .B(n15889), .Z(n15887) );
  XNOR U15466 ( .A(n15890), .B(n15891), .Z(n15849) );
  ANDN U15467 ( .B(n15892), .A(n15893), .Z(n15890) );
  XOR U15468 ( .A(n15891), .B(n15894), .Z(n15892) );
  IV U15469 ( .A(n15848), .Z(n15882) );
  XOR U15470 ( .A(n15846), .B(n15895), .Z(n15848) );
  XOR U15471 ( .A(n15896), .B(n15897), .Z(n15895) );
  ANDN U15472 ( .B(n15898), .A(n15899), .Z(n15896) );
  XOR U15473 ( .A(n15900), .B(n15897), .Z(n15898) );
  IV U15474 ( .A(n15850), .Z(n15846) );
  XOR U15475 ( .A(n15901), .B(n15902), .Z(n15850) );
  ANDN U15476 ( .B(n15903), .A(n15904), .Z(n15901) );
  XOR U15477 ( .A(n15905), .B(n15902), .Z(n15903) );
  IV U15478 ( .A(n15860), .Z(n15864) );
  XOR U15479 ( .A(n15860), .B(n15815), .Z(n15862) );
  XOR U15480 ( .A(n15906), .B(n15907), .Z(n15815) );
  AND U15481 ( .A(n430), .B(n15908), .Z(n15906) );
  XOR U15482 ( .A(n15909), .B(n15907), .Z(n15908) );
  NANDN U15483 ( .A(n15817), .B(n15819), .Z(n15860) );
  XOR U15484 ( .A(n15910), .B(n15911), .Z(n15819) );
  AND U15485 ( .A(n430), .B(n15912), .Z(n15910) );
  XOR U15486 ( .A(n15911), .B(n15913), .Z(n15912) );
  XNOR U15487 ( .A(n15914), .B(n15915), .Z(n430) );
  AND U15488 ( .A(n15916), .B(n15917), .Z(n15914) );
  XOR U15489 ( .A(n15915), .B(n15830), .Z(n15917) );
  XNOR U15490 ( .A(n15918), .B(n15919), .Z(n15830) );
  ANDN U15491 ( .B(n15920), .A(n15921), .Z(n15918) );
  XOR U15492 ( .A(n15919), .B(n15922), .Z(n15920) );
  XNOR U15493 ( .A(n15915), .B(n15832), .Z(n15916) );
  XOR U15494 ( .A(n15923), .B(n15924), .Z(n15832) );
  AND U15495 ( .A(n434), .B(n15925), .Z(n15923) );
  XOR U15496 ( .A(n15926), .B(n15924), .Z(n15925) );
  XNOR U15497 ( .A(n15927), .B(n15928), .Z(n15915) );
  AND U15498 ( .A(n15929), .B(n15930), .Z(n15927) );
  XNOR U15499 ( .A(n15928), .B(n15857), .Z(n15930) );
  XOR U15500 ( .A(n15921), .B(n15922), .Z(n15857) );
  XNOR U15501 ( .A(n15931), .B(n15932), .Z(n15922) );
  ANDN U15502 ( .B(n15933), .A(n15934), .Z(n15931) );
  XOR U15503 ( .A(n15935), .B(n15936), .Z(n15933) );
  XOR U15504 ( .A(n15937), .B(n15938), .Z(n15921) );
  XNOR U15505 ( .A(n15939), .B(n15940), .Z(n15938) );
  ANDN U15506 ( .B(n15941), .A(n15942), .Z(n15939) );
  XNOR U15507 ( .A(n15943), .B(n15944), .Z(n15941) );
  IV U15508 ( .A(n15919), .Z(n15937) );
  XOR U15509 ( .A(n15945), .B(n15946), .Z(n15919) );
  ANDN U15510 ( .B(n15947), .A(n15948), .Z(n15945) );
  XOR U15511 ( .A(n15946), .B(n15949), .Z(n15947) );
  XOR U15512 ( .A(n15928), .B(n15859), .Z(n15929) );
  XOR U15513 ( .A(n15950), .B(n15951), .Z(n15859) );
  AND U15514 ( .A(n434), .B(n15952), .Z(n15950) );
  XOR U15515 ( .A(n15953), .B(n15951), .Z(n15952) );
  XNOR U15516 ( .A(n15954), .B(n15955), .Z(n15928) );
  NAND U15517 ( .A(n15956), .B(n15957), .Z(n15955) );
  XOR U15518 ( .A(n15958), .B(n15907), .Z(n15957) );
  XOR U15519 ( .A(n15948), .B(n15949), .Z(n15907) );
  XOR U15520 ( .A(n15959), .B(n15936), .Z(n15949) );
  XOR U15521 ( .A(n15960), .B(n15961), .Z(n15936) );
  ANDN U15522 ( .B(n15962), .A(n15963), .Z(n15960) );
  XOR U15523 ( .A(n15961), .B(n15964), .Z(n15962) );
  IV U15524 ( .A(n15934), .Z(n15959) );
  XOR U15525 ( .A(n15932), .B(n15965), .Z(n15934) );
  XOR U15526 ( .A(n15966), .B(n15967), .Z(n15965) );
  ANDN U15527 ( .B(n15968), .A(n15969), .Z(n15966) );
  XOR U15528 ( .A(n15970), .B(n15967), .Z(n15968) );
  IV U15529 ( .A(n15935), .Z(n15932) );
  XOR U15530 ( .A(n15971), .B(n15972), .Z(n15935) );
  ANDN U15531 ( .B(n15973), .A(n15974), .Z(n15971) );
  XOR U15532 ( .A(n15972), .B(n15975), .Z(n15973) );
  XOR U15533 ( .A(n15976), .B(n15977), .Z(n15948) );
  XNOR U15534 ( .A(n15943), .B(n15978), .Z(n15977) );
  IV U15535 ( .A(n15946), .Z(n15978) );
  XOR U15536 ( .A(n15979), .B(n15980), .Z(n15946) );
  ANDN U15537 ( .B(n15981), .A(n15982), .Z(n15979) );
  XOR U15538 ( .A(n15980), .B(n15983), .Z(n15981) );
  XNOR U15539 ( .A(n15984), .B(n15985), .Z(n15943) );
  ANDN U15540 ( .B(n15986), .A(n15987), .Z(n15984) );
  XOR U15541 ( .A(n15985), .B(n15988), .Z(n15986) );
  IV U15542 ( .A(n15942), .Z(n15976) );
  XOR U15543 ( .A(n15940), .B(n15989), .Z(n15942) );
  XOR U15544 ( .A(n15990), .B(n15991), .Z(n15989) );
  ANDN U15545 ( .B(n15992), .A(n15993), .Z(n15990) );
  XOR U15546 ( .A(n15994), .B(n15991), .Z(n15992) );
  IV U15547 ( .A(n15944), .Z(n15940) );
  XOR U15548 ( .A(n15995), .B(n15996), .Z(n15944) );
  ANDN U15549 ( .B(n15997), .A(n15998), .Z(n15995) );
  XOR U15550 ( .A(n15999), .B(n15996), .Z(n15997) );
  IV U15551 ( .A(n15954), .Z(n15958) );
  XOR U15552 ( .A(n15954), .B(n15909), .Z(n15956) );
  XOR U15553 ( .A(n16000), .B(n16001), .Z(n15909) );
  AND U15554 ( .A(n434), .B(n16002), .Z(n16000) );
  XOR U15555 ( .A(n16003), .B(n16001), .Z(n16002) );
  NANDN U15556 ( .A(n15911), .B(n15913), .Z(n15954) );
  XOR U15557 ( .A(n16004), .B(n16005), .Z(n15913) );
  AND U15558 ( .A(n434), .B(n16006), .Z(n16004) );
  XOR U15559 ( .A(n16005), .B(n16007), .Z(n16006) );
  XNOR U15560 ( .A(n16008), .B(n16009), .Z(n434) );
  AND U15561 ( .A(n16010), .B(n16011), .Z(n16008) );
  XOR U15562 ( .A(n16009), .B(n15924), .Z(n16011) );
  XNOR U15563 ( .A(n16012), .B(n16013), .Z(n15924) );
  ANDN U15564 ( .B(n16014), .A(n16015), .Z(n16012) );
  XOR U15565 ( .A(n16013), .B(n16016), .Z(n16014) );
  XNOR U15566 ( .A(n16009), .B(n15926), .Z(n16010) );
  XOR U15567 ( .A(n16017), .B(n16018), .Z(n15926) );
  AND U15568 ( .A(n438), .B(n16019), .Z(n16017) );
  XOR U15569 ( .A(n16020), .B(n16018), .Z(n16019) );
  XNOR U15570 ( .A(n16021), .B(n16022), .Z(n16009) );
  AND U15571 ( .A(n16023), .B(n16024), .Z(n16021) );
  XNOR U15572 ( .A(n16022), .B(n15951), .Z(n16024) );
  XOR U15573 ( .A(n16015), .B(n16016), .Z(n15951) );
  XNOR U15574 ( .A(n16025), .B(n16026), .Z(n16016) );
  ANDN U15575 ( .B(n16027), .A(n16028), .Z(n16025) );
  XOR U15576 ( .A(n16029), .B(n16030), .Z(n16027) );
  XOR U15577 ( .A(n16031), .B(n16032), .Z(n16015) );
  XNOR U15578 ( .A(n16033), .B(n16034), .Z(n16032) );
  ANDN U15579 ( .B(n16035), .A(n16036), .Z(n16033) );
  XNOR U15580 ( .A(n16037), .B(n16038), .Z(n16035) );
  IV U15581 ( .A(n16013), .Z(n16031) );
  XOR U15582 ( .A(n16039), .B(n16040), .Z(n16013) );
  ANDN U15583 ( .B(n16041), .A(n16042), .Z(n16039) );
  XOR U15584 ( .A(n16040), .B(n16043), .Z(n16041) );
  XOR U15585 ( .A(n16022), .B(n15953), .Z(n16023) );
  XOR U15586 ( .A(n16044), .B(n16045), .Z(n15953) );
  AND U15587 ( .A(n438), .B(n16046), .Z(n16044) );
  XOR U15588 ( .A(n16047), .B(n16045), .Z(n16046) );
  XNOR U15589 ( .A(n16048), .B(n16049), .Z(n16022) );
  NAND U15590 ( .A(n16050), .B(n16051), .Z(n16049) );
  XOR U15591 ( .A(n16052), .B(n16001), .Z(n16051) );
  XOR U15592 ( .A(n16042), .B(n16043), .Z(n16001) );
  XOR U15593 ( .A(n16053), .B(n16030), .Z(n16043) );
  XOR U15594 ( .A(n16054), .B(n16055), .Z(n16030) );
  ANDN U15595 ( .B(n16056), .A(n16057), .Z(n16054) );
  XOR U15596 ( .A(n16055), .B(n16058), .Z(n16056) );
  IV U15597 ( .A(n16028), .Z(n16053) );
  XOR U15598 ( .A(n16026), .B(n16059), .Z(n16028) );
  XOR U15599 ( .A(n16060), .B(n16061), .Z(n16059) );
  ANDN U15600 ( .B(n16062), .A(n16063), .Z(n16060) );
  XOR U15601 ( .A(n16064), .B(n16061), .Z(n16062) );
  IV U15602 ( .A(n16029), .Z(n16026) );
  XOR U15603 ( .A(n16065), .B(n16066), .Z(n16029) );
  ANDN U15604 ( .B(n16067), .A(n16068), .Z(n16065) );
  XOR U15605 ( .A(n16066), .B(n16069), .Z(n16067) );
  XOR U15606 ( .A(n16070), .B(n16071), .Z(n16042) );
  XNOR U15607 ( .A(n16037), .B(n16072), .Z(n16071) );
  IV U15608 ( .A(n16040), .Z(n16072) );
  XOR U15609 ( .A(n16073), .B(n16074), .Z(n16040) );
  ANDN U15610 ( .B(n16075), .A(n16076), .Z(n16073) );
  XOR U15611 ( .A(n16074), .B(n16077), .Z(n16075) );
  XNOR U15612 ( .A(n16078), .B(n16079), .Z(n16037) );
  ANDN U15613 ( .B(n16080), .A(n16081), .Z(n16078) );
  XOR U15614 ( .A(n16079), .B(n16082), .Z(n16080) );
  IV U15615 ( .A(n16036), .Z(n16070) );
  XOR U15616 ( .A(n16034), .B(n16083), .Z(n16036) );
  XOR U15617 ( .A(n16084), .B(n16085), .Z(n16083) );
  ANDN U15618 ( .B(n16086), .A(n16087), .Z(n16084) );
  XOR U15619 ( .A(n16088), .B(n16085), .Z(n16086) );
  IV U15620 ( .A(n16038), .Z(n16034) );
  XOR U15621 ( .A(n16089), .B(n16090), .Z(n16038) );
  ANDN U15622 ( .B(n16091), .A(n16092), .Z(n16089) );
  XOR U15623 ( .A(n16093), .B(n16090), .Z(n16091) );
  IV U15624 ( .A(n16048), .Z(n16052) );
  XOR U15625 ( .A(n16048), .B(n16003), .Z(n16050) );
  XOR U15626 ( .A(n16094), .B(n16095), .Z(n16003) );
  AND U15627 ( .A(n438), .B(n16096), .Z(n16094) );
  XOR U15628 ( .A(n16097), .B(n16095), .Z(n16096) );
  NANDN U15629 ( .A(n16005), .B(n16007), .Z(n16048) );
  XOR U15630 ( .A(n16098), .B(n16099), .Z(n16007) );
  AND U15631 ( .A(n438), .B(n16100), .Z(n16098) );
  XOR U15632 ( .A(n16099), .B(n16101), .Z(n16100) );
  XNOR U15633 ( .A(n16102), .B(n16103), .Z(n438) );
  AND U15634 ( .A(n16104), .B(n16105), .Z(n16102) );
  XOR U15635 ( .A(n16103), .B(n16018), .Z(n16105) );
  XNOR U15636 ( .A(n16106), .B(n16107), .Z(n16018) );
  ANDN U15637 ( .B(n16108), .A(n16109), .Z(n16106) );
  XOR U15638 ( .A(n16107), .B(n16110), .Z(n16108) );
  XNOR U15639 ( .A(n16103), .B(n16020), .Z(n16104) );
  XOR U15640 ( .A(n16111), .B(n16112), .Z(n16020) );
  AND U15641 ( .A(n442), .B(n16113), .Z(n16111) );
  XOR U15642 ( .A(n16114), .B(n16112), .Z(n16113) );
  XNOR U15643 ( .A(n16115), .B(n16116), .Z(n16103) );
  AND U15644 ( .A(n16117), .B(n16118), .Z(n16115) );
  XNOR U15645 ( .A(n16116), .B(n16045), .Z(n16118) );
  XOR U15646 ( .A(n16109), .B(n16110), .Z(n16045) );
  XNOR U15647 ( .A(n16119), .B(n16120), .Z(n16110) );
  ANDN U15648 ( .B(n16121), .A(n16122), .Z(n16119) );
  XOR U15649 ( .A(n16123), .B(n16124), .Z(n16121) );
  XOR U15650 ( .A(n16125), .B(n16126), .Z(n16109) );
  XNOR U15651 ( .A(n16127), .B(n16128), .Z(n16126) );
  ANDN U15652 ( .B(n16129), .A(n16130), .Z(n16127) );
  XNOR U15653 ( .A(n16131), .B(n16132), .Z(n16129) );
  IV U15654 ( .A(n16107), .Z(n16125) );
  XOR U15655 ( .A(n16133), .B(n16134), .Z(n16107) );
  ANDN U15656 ( .B(n16135), .A(n16136), .Z(n16133) );
  XOR U15657 ( .A(n16134), .B(n16137), .Z(n16135) );
  XOR U15658 ( .A(n16116), .B(n16047), .Z(n16117) );
  XOR U15659 ( .A(n16138), .B(n16139), .Z(n16047) );
  AND U15660 ( .A(n442), .B(n16140), .Z(n16138) );
  XOR U15661 ( .A(n16141), .B(n16139), .Z(n16140) );
  XNOR U15662 ( .A(n16142), .B(n16143), .Z(n16116) );
  NAND U15663 ( .A(n16144), .B(n16145), .Z(n16143) );
  XOR U15664 ( .A(n16146), .B(n16095), .Z(n16145) );
  XOR U15665 ( .A(n16136), .B(n16137), .Z(n16095) );
  XOR U15666 ( .A(n16147), .B(n16124), .Z(n16137) );
  XOR U15667 ( .A(n16148), .B(n16149), .Z(n16124) );
  ANDN U15668 ( .B(n16150), .A(n16151), .Z(n16148) );
  XOR U15669 ( .A(n16149), .B(n16152), .Z(n16150) );
  IV U15670 ( .A(n16122), .Z(n16147) );
  XOR U15671 ( .A(n16120), .B(n16153), .Z(n16122) );
  XOR U15672 ( .A(n16154), .B(n16155), .Z(n16153) );
  ANDN U15673 ( .B(n16156), .A(n16157), .Z(n16154) );
  XOR U15674 ( .A(n16158), .B(n16155), .Z(n16156) );
  IV U15675 ( .A(n16123), .Z(n16120) );
  XOR U15676 ( .A(n16159), .B(n16160), .Z(n16123) );
  ANDN U15677 ( .B(n16161), .A(n16162), .Z(n16159) );
  XOR U15678 ( .A(n16160), .B(n16163), .Z(n16161) );
  XOR U15679 ( .A(n16164), .B(n16165), .Z(n16136) );
  XNOR U15680 ( .A(n16131), .B(n16166), .Z(n16165) );
  IV U15681 ( .A(n16134), .Z(n16166) );
  XOR U15682 ( .A(n16167), .B(n16168), .Z(n16134) );
  ANDN U15683 ( .B(n16169), .A(n16170), .Z(n16167) );
  XOR U15684 ( .A(n16168), .B(n16171), .Z(n16169) );
  XNOR U15685 ( .A(n16172), .B(n16173), .Z(n16131) );
  ANDN U15686 ( .B(n16174), .A(n16175), .Z(n16172) );
  XOR U15687 ( .A(n16173), .B(n16176), .Z(n16174) );
  IV U15688 ( .A(n16130), .Z(n16164) );
  XOR U15689 ( .A(n16128), .B(n16177), .Z(n16130) );
  XOR U15690 ( .A(n16178), .B(n16179), .Z(n16177) );
  ANDN U15691 ( .B(n16180), .A(n16181), .Z(n16178) );
  XOR U15692 ( .A(n16182), .B(n16179), .Z(n16180) );
  IV U15693 ( .A(n16132), .Z(n16128) );
  XOR U15694 ( .A(n16183), .B(n16184), .Z(n16132) );
  ANDN U15695 ( .B(n16185), .A(n16186), .Z(n16183) );
  XOR U15696 ( .A(n16187), .B(n16184), .Z(n16185) );
  IV U15697 ( .A(n16142), .Z(n16146) );
  XOR U15698 ( .A(n16142), .B(n16097), .Z(n16144) );
  XOR U15699 ( .A(n16188), .B(n16189), .Z(n16097) );
  AND U15700 ( .A(n442), .B(n16190), .Z(n16188) );
  XOR U15701 ( .A(n16191), .B(n16189), .Z(n16190) );
  NANDN U15702 ( .A(n16099), .B(n16101), .Z(n16142) );
  XOR U15703 ( .A(n16192), .B(n16193), .Z(n16101) );
  AND U15704 ( .A(n442), .B(n16194), .Z(n16192) );
  XOR U15705 ( .A(n16193), .B(n16195), .Z(n16194) );
  XNOR U15706 ( .A(n16196), .B(n16197), .Z(n442) );
  AND U15707 ( .A(n16198), .B(n16199), .Z(n16196) );
  XOR U15708 ( .A(n16197), .B(n16112), .Z(n16199) );
  XNOR U15709 ( .A(n16200), .B(n16201), .Z(n16112) );
  ANDN U15710 ( .B(n16202), .A(n16203), .Z(n16200) );
  XOR U15711 ( .A(n16201), .B(n16204), .Z(n16202) );
  XNOR U15712 ( .A(n16197), .B(n16114), .Z(n16198) );
  XOR U15713 ( .A(n16205), .B(n16206), .Z(n16114) );
  AND U15714 ( .A(n446), .B(n16207), .Z(n16205) );
  XOR U15715 ( .A(n16208), .B(n16206), .Z(n16207) );
  XNOR U15716 ( .A(n16209), .B(n16210), .Z(n16197) );
  AND U15717 ( .A(n16211), .B(n16212), .Z(n16209) );
  XNOR U15718 ( .A(n16210), .B(n16139), .Z(n16212) );
  XOR U15719 ( .A(n16203), .B(n16204), .Z(n16139) );
  XNOR U15720 ( .A(n16213), .B(n16214), .Z(n16204) );
  ANDN U15721 ( .B(n16215), .A(n16216), .Z(n16213) );
  XOR U15722 ( .A(n16217), .B(n16218), .Z(n16215) );
  XOR U15723 ( .A(n16219), .B(n16220), .Z(n16203) );
  XNOR U15724 ( .A(n16221), .B(n16222), .Z(n16220) );
  ANDN U15725 ( .B(n16223), .A(n16224), .Z(n16221) );
  XNOR U15726 ( .A(n16225), .B(n16226), .Z(n16223) );
  IV U15727 ( .A(n16201), .Z(n16219) );
  XOR U15728 ( .A(n16227), .B(n16228), .Z(n16201) );
  ANDN U15729 ( .B(n16229), .A(n16230), .Z(n16227) );
  XOR U15730 ( .A(n16228), .B(n16231), .Z(n16229) );
  XOR U15731 ( .A(n16210), .B(n16141), .Z(n16211) );
  XOR U15732 ( .A(n16232), .B(n16233), .Z(n16141) );
  AND U15733 ( .A(n446), .B(n16234), .Z(n16232) );
  XOR U15734 ( .A(n16235), .B(n16233), .Z(n16234) );
  XNOR U15735 ( .A(n16236), .B(n16237), .Z(n16210) );
  NAND U15736 ( .A(n16238), .B(n16239), .Z(n16237) );
  XOR U15737 ( .A(n16240), .B(n16189), .Z(n16239) );
  XOR U15738 ( .A(n16230), .B(n16231), .Z(n16189) );
  XOR U15739 ( .A(n16241), .B(n16218), .Z(n16231) );
  XOR U15740 ( .A(n16242), .B(n16243), .Z(n16218) );
  ANDN U15741 ( .B(n16244), .A(n16245), .Z(n16242) );
  XOR U15742 ( .A(n16243), .B(n16246), .Z(n16244) );
  IV U15743 ( .A(n16216), .Z(n16241) );
  XOR U15744 ( .A(n16214), .B(n16247), .Z(n16216) );
  XOR U15745 ( .A(n16248), .B(n16249), .Z(n16247) );
  ANDN U15746 ( .B(n16250), .A(n16251), .Z(n16248) );
  XOR U15747 ( .A(n16252), .B(n16249), .Z(n16250) );
  IV U15748 ( .A(n16217), .Z(n16214) );
  XOR U15749 ( .A(n16253), .B(n16254), .Z(n16217) );
  ANDN U15750 ( .B(n16255), .A(n16256), .Z(n16253) );
  XOR U15751 ( .A(n16254), .B(n16257), .Z(n16255) );
  XOR U15752 ( .A(n16258), .B(n16259), .Z(n16230) );
  XNOR U15753 ( .A(n16225), .B(n16260), .Z(n16259) );
  IV U15754 ( .A(n16228), .Z(n16260) );
  XOR U15755 ( .A(n16261), .B(n16262), .Z(n16228) );
  ANDN U15756 ( .B(n16263), .A(n16264), .Z(n16261) );
  XOR U15757 ( .A(n16262), .B(n16265), .Z(n16263) );
  XNOR U15758 ( .A(n16266), .B(n16267), .Z(n16225) );
  ANDN U15759 ( .B(n16268), .A(n16269), .Z(n16266) );
  XOR U15760 ( .A(n16267), .B(n16270), .Z(n16268) );
  IV U15761 ( .A(n16224), .Z(n16258) );
  XOR U15762 ( .A(n16222), .B(n16271), .Z(n16224) );
  XOR U15763 ( .A(n16272), .B(n16273), .Z(n16271) );
  ANDN U15764 ( .B(n16274), .A(n16275), .Z(n16272) );
  XOR U15765 ( .A(n16276), .B(n16273), .Z(n16274) );
  IV U15766 ( .A(n16226), .Z(n16222) );
  XOR U15767 ( .A(n16277), .B(n16278), .Z(n16226) );
  ANDN U15768 ( .B(n16279), .A(n16280), .Z(n16277) );
  XOR U15769 ( .A(n16281), .B(n16278), .Z(n16279) );
  IV U15770 ( .A(n16236), .Z(n16240) );
  XOR U15771 ( .A(n16236), .B(n16191), .Z(n16238) );
  XOR U15772 ( .A(n16282), .B(n16283), .Z(n16191) );
  AND U15773 ( .A(n446), .B(n16284), .Z(n16282) );
  XOR U15774 ( .A(n16285), .B(n16283), .Z(n16284) );
  NANDN U15775 ( .A(n16193), .B(n16195), .Z(n16236) );
  XOR U15776 ( .A(n16286), .B(n16287), .Z(n16195) );
  AND U15777 ( .A(n446), .B(n16288), .Z(n16286) );
  XOR U15778 ( .A(n16287), .B(n16289), .Z(n16288) );
  XNOR U15779 ( .A(n16290), .B(n16291), .Z(n446) );
  AND U15780 ( .A(n16292), .B(n16293), .Z(n16290) );
  XOR U15781 ( .A(n16291), .B(n16206), .Z(n16293) );
  XNOR U15782 ( .A(n16294), .B(n16295), .Z(n16206) );
  ANDN U15783 ( .B(n16296), .A(n16297), .Z(n16294) );
  XOR U15784 ( .A(n16295), .B(n16298), .Z(n16296) );
  XNOR U15785 ( .A(n16291), .B(n16208), .Z(n16292) );
  XOR U15786 ( .A(n16299), .B(n16300), .Z(n16208) );
  AND U15787 ( .A(n450), .B(n16301), .Z(n16299) );
  XOR U15788 ( .A(n16302), .B(n16300), .Z(n16301) );
  XNOR U15789 ( .A(n16303), .B(n16304), .Z(n16291) );
  AND U15790 ( .A(n16305), .B(n16306), .Z(n16303) );
  XNOR U15791 ( .A(n16304), .B(n16233), .Z(n16306) );
  XOR U15792 ( .A(n16297), .B(n16298), .Z(n16233) );
  XNOR U15793 ( .A(n16307), .B(n16308), .Z(n16298) );
  ANDN U15794 ( .B(n16309), .A(n16310), .Z(n16307) );
  XOR U15795 ( .A(n16311), .B(n16312), .Z(n16309) );
  XOR U15796 ( .A(n16313), .B(n16314), .Z(n16297) );
  XNOR U15797 ( .A(n16315), .B(n16316), .Z(n16314) );
  ANDN U15798 ( .B(n16317), .A(n16318), .Z(n16315) );
  XNOR U15799 ( .A(n16319), .B(n16320), .Z(n16317) );
  IV U15800 ( .A(n16295), .Z(n16313) );
  XOR U15801 ( .A(n16321), .B(n16322), .Z(n16295) );
  ANDN U15802 ( .B(n16323), .A(n16324), .Z(n16321) );
  XOR U15803 ( .A(n16322), .B(n16325), .Z(n16323) );
  XOR U15804 ( .A(n16304), .B(n16235), .Z(n16305) );
  XOR U15805 ( .A(n16326), .B(n16327), .Z(n16235) );
  AND U15806 ( .A(n450), .B(n16328), .Z(n16326) );
  XOR U15807 ( .A(n16329), .B(n16327), .Z(n16328) );
  XNOR U15808 ( .A(n16330), .B(n16331), .Z(n16304) );
  NAND U15809 ( .A(n16332), .B(n16333), .Z(n16331) );
  XOR U15810 ( .A(n16334), .B(n16283), .Z(n16333) );
  XOR U15811 ( .A(n16324), .B(n16325), .Z(n16283) );
  XOR U15812 ( .A(n16335), .B(n16312), .Z(n16325) );
  XOR U15813 ( .A(n16336), .B(n16337), .Z(n16312) );
  ANDN U15814 ( .B(n16338), .A(n16339), .Z(n16336) );
  XOR U15815 ( .A(n16337), .B(n16340), .Z(n16338) );
  IV U15816 ( .A(n16310), .Z(n16335) );
  XOR U15817 ( .A(n16308), .B(n16341), .Z(n16310) );
  XOR U15818 ( .A(n16342), .B(n16343), .Z(n16341) );
  ANDN U15819 ( .B(n16344), .A(n16345), .Z(n16342) );
  XOR U15820 ( .A(n16346), .B(n16343), .Z(n16344) );
  IV U15821 ( .A(n16311), .Z(n16308) );
  XOR U15822 ( .A(n16347), .B(n16348), .Z(n16311) );
  ANDN U15823 ( .B(n16349), .A(n16350), .Z(n16347) );
  XOR U15824 ( .A(n16348), .B(n16351), .Z(n16349) );
  XOR U15825 ( .A(n16352), .B(n16353), .Z(n16324) );
  XNOR U15826 ( .A(n16319), .B(n16354), .Z(n16353) );
  IV U15827 ( .A(n16322), .Z(n16354) );
  XOR U15828 ( .A(n16355), .B(n16356), .Z(n16322) );
  ANDN U15829 ( .B(n16357), .A(n16358), .Z(n16355) );
  XOR U15830 ( .A(n16356), .B(n16359), .Z(n16357) );
  XNOR U15831 ( .A(n16360), .B(n16361), .Z(n16319) );
  ANDN U15832 ( .B(n16362), .A(n16363), .Z(n16360) );
  XOR U15833 ( .A(n16361), .B(n16364), .Z(n16362) );
  IV U15834 ( .A(n16318), .Z(n16352) );
  XOR U15835 ( .A(n16316), .B(n16365), .Z(n16318) );
  XOR U15836 ( .A(n16366), .B(n16367), .Z(n16365) );
  ANDN U15837 ( .B(n16368), .A(n16369), .Z(n16366) );
  XOR U15838 ( .A(n16370), .B(n16367), .Z(n16368) );
  IV U15839 ( .A(n16320), .Z(n16316) );
  XOR U15840 ( .A(n16371), .B(n16372), .Z(n16320) );
  ANDN U15841 ( .B(n16373), .A(n16374), .Z(n16371) );
  XOR U15842 ( .A(n16375), .B(n16372), .Z(n16373) );
  IV U15843 ( .A(n16330), .Z(n16334) );
  XOR U15844 ( .A(n16330), .B(n16285), .Z(n16332) );
  XOR U15845 ( .A(n16376), .B(n16377), .Z(n16285) );
  AND U15846 ( .A(n450), .B(n16378), .Z(n16376) );
  XOR U15847 ( .A(n16379), .B(n16377), .Z(n16378) );
  NANDN U15848 ( .A(n16287), .B(n16289), .Z(n16330) );
  XOR U15849 ( .A(n16380), .B(n16381), .Z(n16289) );
  AND U15850 ( .A(n450), .B(n16382), .Z(n16380) );
  XOR U15851 ( .A(n16381), .B(n16383), .Z(n16382) );
  XNOR U15852 ( .A(n16384), .B(n16385), .Z(n450) );
  AND U15853 ( .A(n16386), .B(n16387), .Z(n16384) );
  XOR U15854 ( .A(n16385), .B(n16300), .Z(n16387) );
  XNOR U15855 ( .A(n16388), .B(n16389), .Z(n16300) );
  ANDN U15856 ( .B(n16390), .A(n16391), .Z(n16388) );
  XOR U15857 ( .A(n16389), .B(n16392), .Z(n16390) );
  XNOR U15858 ( .A(n16385), .B(n16302), .Z(n16386) );
  XOR U15859 ( .A(n16393), .B(n16394), .Z(n16302) );
  AND U15860 ( .A(n454), .B(n16395), .Z(n16393) );
  XOR U15861 ( .A(n16396), .B(n16394), .Z(n16395) );
  XNOR U15862 ( .A(n16397), .B(n16398), .Z(n16385) );
  AND U15863 ( .A(n16399), .B(n16400), .Z(n16397) );
  XNOR U15864 ( .A(n16398), .B(n16327), .Z(n16400) );
  XOR U15865 ( .A(n16391), .B(n16392), .Z(n16327) );
  XNOR U15866 ( .A(n16401), .B(n16402), .Z(n16392) );
  ANDN U15867 ( .B(n16403), .A(n16404), .Z(n16401) );
  XOR U15868 ( .A(n16405), .B(n16406), .Z(n16403) );
  XOR U15869 ( .A(n16407), .B(n16408), .Z(n16391) );
  XNOR U15870 ( .A(n16409), .B(n16410), .Z(n16408) );
  ANDN U15871 ( .B(n16411), .A(n16412), .Z(n16409) );
  XNOR U15872 ( .A(n16413), .B(n16414), .Z(n16411) );
  IV U15873 ( .A(n16389), .Z(n16407) );
  XOR U15874 ( .A(n16415), .B(n16416), .Z(n16389) );
  ANDN U15875 ( .B(n16417), .A(n16418), .Z(n16415) );
  XOR U15876 ( .A(n16416), .B(n16419), .Z(n16417) );
  XOR U15877 ( .A(n16398), .B(n16329), .Z(n16399) );
  XOR U15878 ( .A(n16420), .B(n16421), .Z(n16329) );
  AND U15879 ( .A(n454), .B(n16422), .Z(n16420) );
  XOR U15880 ( .A(n16423), .B(n16421), .Z(n16422) );
  XNOR U15881 ( .A(n16424), .B(n16425), .Z(n16398) );
  NAND U15882 ( .A(n16426), .B(n16427), .Z(n16425) );
  XOR U15883 ( .A(n16428), .B(n16377), .Z(n16427) );
  XOR U15884 ( .A(n16418), .B(n16419), .Z(n16377) );
  XOR U15885 ( .A(n16429), .B(n16406), .Z(n16419) );
  XOR U15886 ( .A(n16430), .B(n16431), .Z(n16406) );
  ANDN U15887 ( .B(n16432), .A(n16433), .Z(n16430) );
  XOR U15888 ( .A(n16431), .B(n16434), .Z(n16432) );
  IV U15889 ( .A(n16404), .Z(n16429) );
  XOR U15890 ( .A(n16402), .B(n16435), .Z(n16404) );
  XOR U15891 ( .A(n16436), .B(n16437), .Z(n16435) );
  ANDN U15892 ( .B(n16438), .A(n16439), .Z(n16436) );
  XOR U15893 ( .A(n16440), .B(n16437), .Z(n16438) );
  IV U15894 ( .A(n16405), .Z(n16402) );
  XOR U15895 ( .A(n16441), .B(n16442), .Z(n16405) );
  ANDN U15896 ( .B(n16443), .A(n16444), .Z(n16441) );
  XOR U15897 ( .A(n16442), .B(n16445), .Z(n16443) );
  XOR U15898 ( .A(n16446), .B(n16447), .Z(n16418) );
  XNOR U15899 ( .A(n16413), .B(n16448), .Z(n16447) );
  IV U15900 ( .A(n16416), .Z(n16448) );
  XOR U15901 ( .A(n16449), .B(n16450), .Z(n16416) );
  ANDN U15902 ( .B(n16451), .A(n16452), .Z(n16449) );
  XOR U15903 ( .A(n16450), .B(n16453), .Z(n16451) );
  XNOR U15904 ( .A(n16454), .B(n16455), .Z(n16413) );
  ANDN U15905 ( .B(n16456), .A(n16457), .Z(n16454) );
  XOR U15906 ( .A(n16455), .B(n16458), .Z(n16456) );
  IV U15907 ( .A(n16412), .Z(n16446) );
  XOR U15908 ( .A(n16410), .B(n16459), .Z(n16412) );
  XOR U15909 ( .A(n16460), .B(n16461), .Z(n16459) );
  ANDN U15910 ( .B(n16462), .A(n16463), .Z(n16460) );
  XOR U15911 ( .A(n16464), .B(n16461), .Z(n16462) );
  IV U15912 ( .A(n16414), .Z(n16410) );
  XOR U15913 ( .A(n16465), .B(n16466), .Z(n16414) );
  ANDN U15914 ( .B(n16467), .A(n16468), .Z(n16465) );
  XOR U15915 ( .A(n16469), .B(n16466), .Z(n16467) );
  IV U15916 ( .A(n16424), .Z(n16428) );
  XOR U15917 ( .A(n16424), .B(n16379), .Z(n16426) );
  XOR U15918 ( .A(n16470), .B(n16471), .Z(n16379) );
  AND U15919 ( .A(n454), .B(n16472), .Z(n16470) );
  XOR U15920 ( .A(n16473), .B(n16471), .Z(n16472) );
  NANDN U15921 ( .A(n16381), .B(n16383), .Z(n16424) );
  XOR U15922 ( .A(n16474), .B(n16475), .Z(n16383) );
  AND U15923 ( .A(n454), .B(n16476), .Z(n16474) );
  XOR U15924 ( .A(n16475), .B(n16477), .Z(n16476) );
  XNOR U15925 ( .A(n16478), .B(n16479), .Z(n454) );
  AND U15926 ( .A(n16480), .B(n16481), .Z(n16478) );
  XOR U15927 ( .A(n16479), .B(n16394), .Z(n16481) );
  XNOR U15928 ( .A(n16482), .B(n16483), .Z(n16394) );
  ANDN U15929 ( .B(n16484), .A(n16485), .Z(n16482) );
  XOR U15930 ( .A(n16483), .B(n16486), .Z(n16484) );
  XNOR U15931 ( .A(n16479), .B(n16396), .Z(n16480) );
  XOR U15932 ( .A(n16487), .B(n16488), .Z(n16396) );
  AND U15933 ( .A(n458), .B(n16489), .Z(n16487) );
  XOR U15934 ( .A(n16490), .B(n16488), .Z(n16489) );
  XNOR U15935 ( .A(n16491), .B(n16492), .Z(n16479) );
  AND U15936 ( .A(n16493), .B(n16494), .Z(n16491) );
  XNOR U15937 ( .A(n16492), .B(n16421), .Z(n16494) );
  XOR U15938 ( .A(n16485), .B(n16486), .Z(n16421) );
  XNOR U15939 ( .A(n16495), .B(n16496), .Z(n16486) );
  ANDN U15940 ( .B(n16497), .A(n16498), .Z(n16495) );
  XOR U15941 ( .A(n16499), .B(n16500), .Z(n16497) );
  XOR U15942 ( .A(n16501), .B(n16502), .Z(n16485) );
  XNOR U15943 ( .A(n16503), .B(n16504), .Z(n16502) );
  ANDN U15944 ( .B(n16505), .A(n16506), .Z(n16503) );
  XNOR U15945 ( .A(n16507), .B(n16508), .Z(n16505) );
  IV U15946 ( .A(n16483), .Z(n16501) );
  XOR U15947 ( .A(n16509), .B(n16510), .Z(n16483) );
  ANDN U15948 ( .B(n16511), .A(n16512), .Z(n16509) );
  XOR U15949 ( .A(n16510), .B(n16513), .Z(n16511) );
  XOR U15950 ( .A(n16492), .B(n16423), .Z(n16493) );
  XOR U15951 ( .A(n16514), .B(n16515), .Z(n16423) );
  AND U15952 ( .A(n458), .B(n16516), .Z(n16514) );
  XOR U15953 ( .A(n16517), .B(n16515), .Z(n16516) );
  XNOR U15954 ( .A(n16518), .B(n16519), .Z(n16492) );
  NAND U15955 ( .A(n16520), .B(n16521), .Z(n16519) );
  XOR U15956 ( .A(n16522), .B(n16471), .Z(n16521) );
  XOR U15957 ( .A(n16512), .B(n16513), .Z(n16471) );
  XOR U15958 ( .A(n16523), .B(n16500), .Z(n16513) );
  XOR U15959 ( .A(n16524), .B(n16525), .Z(n16500) );
  ANDN U15960 ( .B(n16526), .A(n16527), .Z(n16524) );
  XOR U15961 ( .A(n16525), .B(n16528), .Z(n16526) );
  IV U15962 ( .A(n16498), .Z(n16523) );
  XOR U15963 ( .A(n16496), .B(n16529), .Z(n16498) );
  XOR U15964 ( .A(n16530), .B(n16531), .Z(n16529) );
  ANDN U15965 ( .B(n16532), .A(n16533), .Z(n16530) );
  XOR U15966 ( .A(n16534), .B(n16531), .Z(n16532) );
  IV U15967 ( .A(n16499), .Z(n16496) );
  XOR U15968 ( .A(n16535), .B(n16536), .Z(n16499) );
  ANDN U15969 ( .B(n16537), .A(n16538), .Z(n16535) );
  XOR U15970 ( .A(n16536), .B(n16539), .Z(n16537) );
  XOR U15971 ( .A(n16540), .B(n16541), .Z(n16512) );
  XNOR U15972 ( .A(n16507), .B(n16542), .Z(n16541) );
  IV U15973 ( .A(n16510), .Z(n16542) );
  XOR U15974 ( .A(n16543), .B(n16544), .Z(n16510) );
  ANDN U15975 ( .B(n16545), .A(n16546), .Z(n16543) );
  XOR U15976 ( .A(n16544), .B(n16547), .Z(n16545) );
  XNOR U15977 ( .A(n16548), .B(n16549), .Z(n16507) );
  ANDN U15978 ( .B(n16550), .A(n16551), .Z(n16548) );
  XOR U15979 ( .A(n16549), .B(n16552), .Z(n16550) );
  IV U15980 ( .A(n16506), .Z(n16540) );
  XOR U15981 ( .A(n16504), .B(n16553), .Z(n16506) );
  XOR U15982 ( .A(n16554), .B(n16555), .Z(n16553) );
  ANDN U15983 ( .B(n16556), .A(n16557), .Z(n16554) );
  XOR U15984 ( .A(n16558), .B(n16555), .Z(n16556) );
  IV U15985 ( .A(n16508), .Z(n16504) );
  XOR U15986 ( .A(n16559), .B(n16560), .Z(n16508) );
  ANDN U15987 ( .B(n16561), .A(n16562), .Z(n16559) );
  XOR U15988 ( .A(n16563), .B(n16560), .Z(n16561) );
  IV U15989 ( .A(n16518), .Z(n16522) );
  XOR U15990 ( .A(n16518), .B(n16473), .Z(n16520) );
  XOR U15991 ( .A(n16564), .B(n16565), .Z(n16473) );
  AND U15992 ( .A(n458), .B(n16566), .Z(n16564) );
  XOR U15993 ( .A(n16567), .B(n16565), .Z(n16566) );
  NANDN U15994 ( .A(n16475), .B(n16477), .Z(n16518) );
  XOR U15995 ( .A(n16568), .B(n16569), .Z(n16477) );
  AND U15996 ( .A(n458), .B(n16570), .Z(n16568) );
  XOR U15997 ( .A(n16569), .B(n16571), .Z(n16570) );
  XNOR U15998 ( .A(n16572), .B(n16573), .Z(n458) );
  AND U15999 ( .A(n16574), .B(n16575), .Z(n16572) );
  XOR U16000 ( .A(n16573), .B(n16488), .Z(n16575) );
  XNOR U16001 ( .A(n16576), .B(n16577), .Z(n16488) );
  ANDN U16002 ( .B(n16578), .A(n16579), .Z(n16576) );
  XOR U16003 ( .A(n16577), .B(n16580), .Z(n16578) );
  XNOR U16004 ( .A(n16573), .B(n16490), .Z(n16574) );
  XOR U16005 ( .A(n16581), .B(n16582), .Z(n16490) );
  AND U16006 ( .A(n462), .B(n16583), .Z(n16581) );
  XOR U16007 ( .A(n16584), .B(n16582), .Z(n16583) );
  XNOR U16008 ( .A(n16585), .B(n16586), .Z(n16573) );
  AND U16009 ( .A(n16587), .B(n16588), .Z(n16585) );
  XNOR U16010 ( .A(n16586), .B(n16515), .Z(n16588) );
  XOR U16011 ( .A(n16579), .B(n16580), .Z(n16515) );
  XNOR U16012 ( .A(n16589), .B(n16590), .Z(n16580) );
  ANDN U16013 ( .B(n16591), .A(n16592), .Z(n16589) );
  XOR U16014 ( .A(n16593), .B(n16594), .Z(n16591) );
  XOR U16015 ( .A(n16595), .B(n16596), .Z(n16579) );
  XNOR U16016 ( .A(n16597), .B(n16598), .Z(n16596) );
  ANDN U16017 ( .B(n16599), .A(n16600), .Z(n16597) );
  XNOR U16018 ( .A(n16601), .B(n16602), .Z(n16599) );
  IV U16019 ( .A(n16577), .Z(n16595) );
  XOR U16020 ( .A(n16603), .B(n16604), .Z(n16577) );
  ANDN U16021 ( .B(n16605), .A(n16606), .Z(n16603) );
  XOR U16022 ( .A(n16604), .B(n16607), .Z(n16605) );
  XOR U16023 ( .A(n16586), .B(n16517), .Z(n16587) );
  XOR U16024 ( .A(n16608), .B(n16609), .Z(n16517) );
  AND U16025 ( .A(n462), .B(n16610), .Z(n16608) );
  XOR U16026 ( .A(n16611), .B(n16609), .Z(n16610) );
  XNOR U16027 ( .A(n16612), .B(n16613), .Z(n16586) );
  NAND U16028 ( .A(n16614), .B(n16615), .Z(n16613) );
  XOR U16029 ( .A(n16616), .B(n16565), .Z(n16615) );
  XOR U16030 ( .A(n16606), .B(n16607), .Z(n16565) );
  XOR U16031 ( .A(n16617), .B(n16594), .Z(n16607) );
  XOR U16032 ( .A(n16618), .B(n16619), .Z(n16594) );
  ANDN U16033 ( .B(n16620), .A(n16621), .Z(n16618) );
  XOR U16034 ( .A(n16619), .B(n16622), .Z(n16620) );
  IV U16035 ( .A(n16592), .Z(n16617) );
  XOR U16036 ( .A(n16590), .B(n16623), .Z(n16592) );
  XOR U16037 ( .A(n16624), .B(n16625), .Z(n16623) );
  ANDN U16038 ( .B(n16626), .A(n16627), .Z(n16624) );
  XOR U16039 ( .A(n16628), .B(n16625), .Z(n16626) );
  IV U16040 ( .A(n16593), .Z(n16590) );
  XOR U16041 ( .A(n16629), .B(n16630), .Z(n16593) );
  ANDN U16042 ( .B(n16631), .A(n16632), .Z(n16629) );
  XOR U16043 ( .A(n16630), .B(n16633), .Z(n16631) );
  XOR U16044 ( .A(n16634), .B(n16635), .Z(n16606) );
  XNOR U16045 ( .A(n16601), .B(n16636), .Z(n16635) );
  IV U16046 ( .A(n16604), .Z(n16636) );
  XOR U16047 ( .A(n16637), .B(n16638), .Z(n16604) );
  ANDN U16048 ( .B(n16639), .A(n16640), .Z(n16637) );
  XOR U16049 ( .A(n16638), .B(n16641), .Z(n16639) );
  XNOR U16050 ( .A(n16642), .B(n16643), .Z(n16601) );
  ANDN U16051 ( .B(n16644), .A(n16645), .Z(n16642) );
  XOR U16052 ( .A(n16643), .B(n16646), .Z(n16644) );
  IV U16053 ( .A(n16600), .Z(n16634) );
  XOR U16054 ( .A(n16598), .B(n16647), .Z(n16600) );
  XOR U16055 ( .A(n16648), .B(n16649), .Z(n16647) );
  ANDN U16056 ( .B(n16650), .A(n16651), .Z(n16648) );
  XOR U16057 ( .A(n16652), .B(n16649), .Z(n16650) );
  IV U16058 ( .A(n16602), .Z(n16598) );
  XOR U16059 ( .A(n16653), .B(n16654), .Z(n16602) );
  ANDN U16060 ( .B(n16655), .A(n16656), .Z(n16653) );
  XOR U16061 ( .A(n16657), .B(n16654), .Z(n16655) );
  IV U16062 ( .A(n16612), .Z(n16616) );
  XOR U16063 ( .A(n16612), .B(n16567), .Z(n16614) );
  XOR U16064 ( .A(n16658), .B(n16659), .Z(n16567) );
  AND U16065 ( .A(n462), .B(n16660), .Z(n16658) );
  XOR U16066 ( .A(n16661), .B(n16659), .Z(n16660) );
  NANDN U16067 ( .A(n16569), .B(n16571), .Z(n16612) );
  XOR U16068 ( .A(n16662), .B(n16663), .Z(n16571) );
  AND U16069 ( .A(n462), .B(n16664), .Z(n16662) );
  XOR U16070 ( .A(n16663), .B(n16665), .Z(n16664) );
  XNOR U16071 ( .A(n16666), .B(n16667), .Z(n462) );
  AND U16072 ( .A(n16668), .B(n16669), .Z(n16666) );
  XOR U16073 ( .A(n16667), .B(n16582), .Z(n16669) );
  XNOR U16074 ( .A(n16670), .B(n16671), .Z(n16582) );
  ANDN U16075 ( .B(n16672), .A(n16673), .Z(n16670) );
  XOR U16076 ( .A(n16671), .B(n16674), .Z(n16672) );
  XNOR U16077 ( .A(n16667), .B(n16584), .Z(n16668) );
  XOR U16078 ( .A(n16675), .B(n16676), .Z(n16584) );
  AND U16079 ( .A(n466), .B(n16677), .Z(n16675) );
  XOR U16080 ( .A(n16678), .B(n16676), .Z(n16677) );
  XNOR U16081 ( .A(n16679), .B(n16680), .Z(n16667) );
  AND U16082 ( .A(n16681), .B(n16682), .Z(n16679) );
  XNOR U16083 ( .A(n16680), .B(n16609), .Z(n16682) );
  XOR U16084 ( .A(n16673), .B(n16674), .Z(n16609) );
  XNOR U16085 ( .A(n16683), .B(n16684), .Z(n16674) );
  ANDN U16086 ( .B(n16685), .A(n16686), .Z(n16683) );
  XOR U16087 ( .A(n16687), .B(n16688), .Z(n16685) );
  XOR U16088 ( .A(n16689), .B(n16690), .Z(n16673) );
  XNOR U16089 ( .A(n16691), .B(n16692), .Z(n16690) );
  ANDN U16090 ( .B(n16693), .A(n16694), .Z(n16691) );
  XNOR U16091 ( .A(n16695), .B(n16696), .Z(n16693) );
  IV U16092 ( .A(n16671), .Z(n16689) );
  XOR U16093 ( .A(n16697), .B(n16698), .Z(n16671) );
  ANDN U16094 ( .B(n16699), .A(n16700), .Z(n16697) );
  XOR U16095 ( .A(n16698), .B(n16701), .Z(n16699) );
  XOR U16096 ( .A(n16680), .B(n16611), .Z(n16681) );
  XOR U16097 ( .A(n16702), .B(n16703), .Z(n16611) );
  AND U16098 ( .A(n466), .B(n16704), .Z(n16702) );
  XOR U16099 ( .A(n16705), .B(n16703), .Z(n16704) );
  XNOR U16100 ( .A(n16706), .B(n16707), .Z(n16680) );
  NAND U16101 ( .A(n16708), .B(n16709), .Z(n16707) );
  XOR U16102 ( .A(n16710), .B(n16659), .Z(n16709) );
  XOR U16103 ( .A(n16700), .B(n16701), .Z(n16659) );
  XOR U16104 ( .A(n16711), .B(n16688), .Z(n16701) );
  XOR U16105 ( .A(n16712), .B(n16713), .Z(n16688) );
  ANDN U16106 ( .B(n16714), .A(n16715), .Z(n16712) );
  XOR U16107 ( .A(n16713), .B(n16716), .Z(n16714) );
  IV U16108 ( .A(n16686), .Z(n16711) );
  XOR U16109 ( .A(n16684), .B(n16717), .Z(n16686) );
  XOR U16110 ( .A(n16718), .B(n16719), .Z(n16717) );
  ANDN U16111 ( .B(n16720), .A(n16721), .Z(n16718) );
  XOR U16112 ( .A(n16722), .B(n16719), .Z(n16720) );
  IV U16113 ( .A(n16687), .Z(n16684) );
  XOR U16114 ( .A(n16723), .B(n16724), .Z(n16687) );
  ANDN U16115 ( .B(n16725), .A(n16726), .Z(n16723) );
  XOR U16116 ( .A(n16724), .B(n16727), .Z(n16725) );
  XOR U16117 ( .A(n16728), .B(n16729), .Z(n16700) );
  XNOR U16118 ( .A(n16695), .B(n16730), .Z(n16729) );
  IV U16119 ( .A(n16698), .Z(n16730) );
  XOR U16120 ( .A(n16731), .B(n16732), .Z(n16698) );
  ANDN U16121 ( .B(n16733), .A(n16734), .Z(n16731) );
  XOR U16122 ( .A(n16732), .B(n16735), .Z(n16733) );
  XNOR U16123 ( .A(n16736), .B(n16737), .Z(n16695) );
  ANDN U16124 ( .B(n16738), .A(n16739), .Z(n16736) );
  XOR U16125 ( .A(n16737), .B(n16740), .Z(n16738) );
  IV U16126 ( .A(n16694), .Z(n16728) );
  XOR U16127 ( .A(n16692), .B(n16741), .Z(n16694) );
  XOR U16128 ( .A(n16742), .B(n16743), .Z(n16741) );
  ANDN U16129 ( .B(n16744), .A(n16745), .Z(n16742) );
  XOR U16130 ( .A(n16746), .B(n16743), .Z(n16744) );
  IV U16131 ( .A(n16696), .Z(n16692) );
  XOR U16132 ( .A(n16747), .B(n16748), .Z(n16696) );
  ANDN U16133 ( .B(n16749), .A(n16750), .Z(n16747) );
  XOR U16134 ( .A(n16751), .B(n16748), .Z(n16749) );
  IV U16135 ( .A(n16706), .Z(n16710) );
  XOR U16136 ( .A(n16706), .B(n16661), .Z(n16708) );
  XOR U16137 ( .A(n16752), .B(n16753), .Z(n16661) );
  AND U16138 ( .A(n466), .B(n16754), .Z(n16752) );
  XOR U16139 ( .A(n16755), .B(n16753), .Z(n16754) );
  NANDN U16140 ( .A(n16663), .B(n16665), .Z(n16706) );
  XOR U16141 ( .A(n16756), .B(n16757), .Z(n16665) );
  AND U16142 ( .A(n466), .B(n16758), .Z(n16756) );
  XOR U16143 ( .A(n16757), .B(n16759), .Z(n16758) );
  XNOR U16144 ( .A(n16760), .B(n16761), .Z(n466) );
  AND U16145 ( .A(n16762), .B(n16763), .Z(n16760) );
  XOR U16146 ( .A(n16761), .B(n16676), .Z(n16763) );
  XNOR U16147 ( .A(n16764), .B(n16765), .Z(n16676) );
  ANDN U16148 ( .B(n16766), .A(n16767), .Z(n16764) );
  XOR U16149 ( .A(n16765), .B(n16768), .Z(n16766) );
  XNOR U16150 ( .A(n16761), .B(n16678), .Z(n16762) );
  XOR U16151 ( .A(n16769), .B(n16770), .Z(n16678) );
  AND U16152 ( .A(n470), .B(n16771), .Z(n16769) );
  XOR U16153 ( .A(n16772), .B(n16770), .Z(n16771) );
  XNOR U16154 ( .A(n16773), .B(n16774), .Z(n16761) );
  AND U16155 ( .A(n16775), .B(n16776), .Z(n16773) );
  XNOR U16156 ( .A(n16774), .B(n16703), .Z(n16776) );
  XOR U16157 ( .A(n16767), .B(n16768), .Z(n16703) );
  XNOR U16158 ( .A(n16777), .B(n16778), .Z(n16768) );
  ANDN U16159 ( .B(n16779), .A(n16780), .Z(n16777) );
  XOR U16160 ( .A(n16781), .B(n16782), .Z(n16779) );
  XOR U16161 ( .A(n16783), .B(n16784), .Z(n16767) );
  XNOR U16162 ( .A(n16785), .B(n16786), .Z(n16784) );
  ANDN U16163 ( .B(n16787), .A(n16788), .Z(n16785) );
  XNOR U16164 ( .A(n16789), .B(n16790), .Z(n16787) );
  IV U16165 ( .A(n16765), .Z(n16783) );
  XOR U16166 ( .A(n16791), .B(n16792), .Z(n16765) );
  ANDN U16167 ( .B(n16793), .A(n16794), .Z(n16791) );
  XOR U16168 ( .A(n16792), .B(n16795), .Z(n16793) );
  XOR U16169 ( .A(n16774), .B(n16705), .Z(n16775) );
  XOR U16170 ( .A(n16796), .B(n16797), .Z(n16705) );
  AND U16171 ( .A(n470), .B(n16798), .Z(n16796) );
  XOR U16172 ( .A(n16799), .B(n16797), .Z(n16798) );
  XNOR U16173 ( .A(n16800), .B(n16801), .Z(n16774) );
  NAND U16174 ( .A(n16802), .B(n16803), .Z(n16801) );
  XOR U16175 ( .A(n16804), .B(n16753), .Z(n16803) );
  XOR U16176 ( .A(n16794), .B(n16795), .Z(n16753) );
  XOR U16177 ( .A(n16805), .B(n16782), .Z(n16795) );
  XOR U16178 ( .A(n16806), .B(n16807), .Z(n16782) );
  ANDN U16179 ( .B(n16808), .A(n16809), .Z(n16806) );
  XOR U16180 ( .A(n16807), .B(n16810), .Z(n16808) );
  IV U16181 ( .A(n16780), .Z(n16805) );
  XOR U16182 ( .A(n16778), .B(n16811), .Z(n16780) );
  XOR U16183 ( .A(n16812), .B(n16813), .Z(n16811) );
  ANDN U16184 ( .B(n16814), .A(n16815), .Z(n16812) );
  XOR U16185 ( .A(n16816), .B(n16813), .Z(n16814) );
  IV U16186 ( .A(n16781), .Z(n16778) );
  XOR U16187 ( .A(n16817), .B(n16818), .Z(n16781) );
  ANDN U16188 ( .B(n16819), .A(n16820), .Z(n16817) );
  XOR U16189 ( .A(n16818), .B(n16821), .Z(n16819) );
  XOR U16190 ( .A(n16822), .B(n16823), .Z(n16794) );
  XNOR U16191 ( .A(n16789), .B(n16824), .Z(n16823) );
  IV U16192 ( .A(n16792), .Z(n16824) );
  XOR U16193 ( .A(n16825), .B(n16826), .Z(n16792) );
  ANDN U16194 ( .B(n16827), .A(n16828), .Z(n16825) );
  XOR U16195 ( .A(n16826), .B(n16829), .Z(n16827) );
  XNOR U16196 ( .A(n16830), .B(n16831), .Z(n16789) );
  ANDN U16197 ( .B(n16832), .A(n16833), .Z(n16830) );
  XOR U16198 ( .A(n16831), .B(n16834), .Z(n16832) );
  IV U16199 ( .A(n16788), .Z(n16822) );
  XOR U16200 ( .A(n16786), .B(n16835), .Z(n16788) );
  XOR U16201 ( .A(n16836), .B(n16837), .Z(n16835) );
  ANDN U16202 ( .B(n16838), .A(n16839), .Z(n16836) );
  XOR U16203 ( .A(n16840), .B(n16837), .Z(n16838) );
  IV U16204 ( .A(n16790), .Z(n16786) );
  XOR U16205 ( .A(n16841), .B(n16842), .Z(n16790) );
  ANDN U16206 ( .B(n16843), .A(n16844), .Z(n16841) );
  XOR U16207 ( .A(n16845), .B(n16842), .Z(n16843) );
  IV U16208 ( .A(n16800), .Z(n16804) );
  XOR U16209 ( .A(n16800), .B(n16755), .Z(n16802) );
  XOR U16210 ( .A(n16846), .B(n16847), .Z(n16755) );
  AND U16211 ( .A(n470), .B(n16848), .Z(n16846) );
  XOR U16212 ( .A(n16849), .B(n16847), .Z(n16848) );
  NANDN U16213 ( .A(n16757), .B(n16759), .Z(n16800) );
  XOR U16214 ( .A(n16850), .B(n16851), .Z(n16759) );
  AND U16215 ( .A(n470), .B(n16852), .Z(n16850) );
  XOR U16216 ( .A(n16851), .B(n16853), .Z(n16852) );
  XNOR U16217 ( .A(n16854), .B(n16855), .Z(n470) );
  AND U16218 ( .A(n16856), .B(n16857), .Z(n16854) );
  XOR U16219 ( .A(n16855), .B(n16770), .Z(n16857) );
  XNOR U16220 ( .A(n16858), .B(n16859), .Z(n16770) );
  ANDN U16221 ( .B(n16860), .A(n16861), .Z(n16858) );
  XOR U16222 ( .A(n16859), .B(n16862), .Z(n16860) );
  XNOR U16223 ( .A(n16855), .B(n16772), .Z(n16856) );
  XOR U16224 ( .A(n16863), .B(n16864), .Z(n16772) );
  AND U16225 ( .A(n474), .B(n16865), .Z(n16863) );
  XOR U16226 ( .A(n16866), .B(n16864), .Z(n16865) );
  XNOR U16227 ( .A(n16867), .B(n16868), .Z(n16855) );
  AND U16228 ( .A(n16869), .B(n16870), .Z(n16867) );
  XNOR U16229 ( .A(n16868), .B(n16797), .Z(n16870) );
  XOR U16230 ( .A(n16861), .B(n16862), .Z(n16797) );
  XNOR U16231 ( .A(n16871), .B(n16872), .Z(n16862) );
  ANDN U16232 ( .B(n16873), .A(n16874), .Z(n16871) );
  XOR U16233 ( .A(n16875), .B(n16876), .Z(n16873) );
  XOR U16234 ( .A(n16877), .B(n16878), .Z(n16861) );
  XNOR U16235 ( .A(n16879), .B(n16880), .Z(n16878) );
  ANDN U16236 ( .B(n16881), .A(n16882), .Z(n16879) );
  XNOR U16237 ( .A(n16883), .B(n16884), .Z(n16881) );
  IV U16238 ( .A(n16859), .Z(n16877) );
  XOR U16239 ( .A(n16885), .B(n16886), .Z(n16859) );
  ANDN U16240 ( .B(n16887), .A(n16888), .Z(n16885) );
  XOR U16241 ( .A(n16886), .B(n16889), .Z(n16887) );
  XOR U16242 ( .A(n16868), .B(n16799), .Z(n16869) );
  XOR U16243 ( .A(n16890), .B(n16891), .Z(n16799) );
  AND U16244 ( .A(n474), .B(n16892), .Z(n16890) );
  XOR U16245 ( .A(n16893), .B(n16891), .Z(n16892) );
  XNOR U16246 ( .A(n16894), .B(n16895), .Z(n16868) );
  NAND U16247 ( .A(n16896), .B(n16897), .Z(n16895) );
  XOR U16248 ( .A(n16898), .B(n16847), .Z(n16897) );
  XOR U16249 ( .A(n16888), .B(n16889), .Z(n16847) );
  XOR U16250 ( .A(n16899), .B(n16876), .Z(n16889) );
  XOR U16251 ( .A(n16900), .B(n16901), .Z(n16876) );
  ANDN U16252 ( .B(n16902), .A(n16903), .Z(n16900) );
  XOR U16253 ( .A(n16901), .B(n16904), .Z(n16902) );
  IV U16254 ( .A(n16874), .Z(n16899) );
  XOR U16255 ( .A(n16872), .B(n16905), .Z(n16874) );
  XOR U16256 ( .A(n16906), .B(n16907), .Z(n16905) );
  ANDN U16257 ( .B(n16908), .A(n16909), .Z(n16906) );
  XOR U16258 ( .A(n16910), .B(n16907), .Z(n16908) );
  IV U16259 ( .A(n16875), .Z(n16872) );
  XOR U16260 ( .A(n16911), .B(n16912), .Z(n16875) );
  ANDN U16261 ( .B(n16913), .A(n16914), .Z(n16911) );
  XOR U16262 ( .A(n16912), .B(n16915), .Z(n16913) );
  XOR U16263 ( .A(n16916), .B(n16917), .Z(n16888) );
  XNOR U16264 ( .A(n16883), .B(n16918), .Z(n16917) );
  IV U16265 ( .A(n16886), .Z(n16918) );
  XOR U16266 ( .A(n16919), .B(n16920), .Z(n16886) );
  ANDN U16267 ( .B(n16921), .A(n16922), .Z(n16919) );
  XOR U16268 ( .A(n16920), .B(n16923), .Z(n16921) );
  XNOR U16269 ( .A(n16924), .B(n16925), .Z(n16883) );
  ANDN U16270 ( .B(n16926), .A(n16927), .Z(n16924) );
  XOR U16271 ( .A(n16925), .B(n16928), .Z(n16926) );
  IV U16272 ( .A(n16882), .Z(n16916) );
  XOR U16273 ( .A(n16880), .B(n16929), .Z(n16882) );
  XOR U16274 ( .A(n16930), .B(n16931), .Z(n16929) );
  ANDN U16275 ( .B(n16932), .A(n16933), .Z(n16930) );
  XOR U16276 ( .A(n16934), .B(n16931), .Z(n16932) );
  IV U16277 ( .A(n16884), .Z(n16880) );
  XOR U16278 ( .A(n16935), .B(n16936), .Z(n16884) );
  ANDN U16279 ( .B(n16937), .A(n16938), .Z(n16935) );
  XOR U16280 ( .A(n16939), .B(n16936), .Z(n16937) );
  IV U16281 ( .A(n16894), .Z(n16898) );
  XOR U16282 ( .A(n16894), .B(n16849), .Z(n16896) );
  XOR U16283 ( .A(n16940), .B(n16941), .Z(n16849) );
  AND U16284 ( .A(n474), .B(n16942), .Z(n16940) );
  XOR U16285 ( .A(n16943), .B(n16941), .Z(n16942) );
  NANDN U16286 ( .A(n16851), .B(n16853), .Z(n16894) );
  XOR U16287 ( .A(n16944), .B(n16945), .Z(n16853) );
  AND U16288 ( .A(n474), .B(n16946), .Z(n16944) );
  XOR U16289 ( .A(n16945), .B(n16947), .Z(n16946) );
  XNOR U16290 ( .A(n16948), .B(n16949), .Z(n474) );
  AND U16291 ( .A(n16950), .B(n16951), .Z(n16948) );
  XOR U16292 ( .A(n16949), .B(n16864), .Z(n16951) );
  XNOR U16293 ( .A(n16952), .B(n16953), .Z(n16864) );
  ANDN U16294 ( .B(n16954), .A(n16955), .Z(n16952) );
  XOR U16295 ( .A(n16953), .B(n16956), .Z(n16954) );
  XNOR U16296 ( .A(n16949), .B(n16866), .Z(n16950) );
  XOR U16297 ( .A(n16957), .B(n16958), .Z(n16866) );
  AND U16298 ( .A(n478), .B(n16959), .Z(n16957) );
  XOR U16299 ( .A(n16960), .B(n16958), .Z(n16959) );
  XNOR U16300 ( .A(n16961), .B(n16962), .Z(n16949) );
  AND U16301 ( .A(n16963), .B(n16964), .Z(n16961) );
  XNOR U16302 ( .A(n16962), .B(n16891), .Z(n16964) );
  XOR U16303 ( .A(n16955), .B(n16956), .Z(n16891) );
  XNOR U16304 ( .A(n16965), .B(n16966), .Z(n16956) );
  ANDN U16305 ( .B(n16967), .A(n16968), .Z(n16965) );
  XOR U16306 ( .A(n16969), .B(n16970), .Z(n16967) );
  XOR U16307 ( .A(n16971), .B(n16972), .Z(n16955) );
  XNOR U16308 ( .A(n16973), .B(n16974), .Z(n16972) );
  ANDN U16309 ( .B(n16975), .A(n16976), .Z(n16973) );
  XNOR U16310 ( .A(n16977), .B(n16978), .Z(n16975) );
  IV U16311 ( .A(n16953), .Z(n16971) );
  XOR U16312 ( .A(n16979), .B(n16980), .Z(n16953) );
  ANDN U16313 ( .B(n16981), .A(n16982), .Z(n16979) );
  XOR U16314 ( .A(n16980), .B(n16983), .Z(n16981) );
  XOR U16315 ( .A(n16962), .B(n16893), .Z(n16963) );
  XOR U16316 ( .A(n16984), .B(n16985), .Z(n16893) );
  AND U16317 ( .A(n478), .B(n16986), .Z(n16984) );
  XOR U16318 ( .A(n16987), .B(n16985), .Z(n16986) );
  XNOR U16319 ( .A(n16988), .B(n16989), .Z(n16962) );
  NAND U16320 ( .A(n16990), .B(n16991), .Z(n16989) );
  XOR U16321 ( .A(n16992), .B(n16941), .Z(n16991) );
  XOR U16322 ( .A(n16982), .B(n16983), .Z(n16941) );
  XOR U16323 ( .A(n16993), .B(n16970), .Z(n16983) );
  XOR U16324 ( .A(n16994), .B(n16995), .Z(n16970) );
  ANDN U16325 ( .B(n16996), .A(n16997), .Z(n16994) );
  XOR U16326 ( .A(n16995), .B(n16998), .Z(n16996) );
  IV U16327 ( .A(n16968), .Z(n16993) );
  XOR U16328 ( .A(n16966), .B(n16999), .Z(n16968) );
  XOR U16329 ( .A(n17000), .B(n17001), .Z(n16999) );
  ANDN U16330 ( .B(n17002), .A(n17003), .Z(n17000) );
  XOR U16331 ( .A(n17004), .B(n17001), .Z(n17002) );
  IV U16332 ( .A(n16969), .Z(n16966) );
  XOR U16333 ( .A(n17005), .B(n17006), .Z(n16969) );
  ANDN U16334 ( .B(n17007), .A(n17008), .Z(n17005) );
  XOR U16335 ( .A(n17006), .B(n17009), .Z(n17007) );
  XOR U16336 ( .A(n17010), .B(n17011), .Z(n16982) );
  XNOR U16337 ( .A(n16977), .B(n17012), .Z(n17011) );
  IV U16338 ( .A(n16980), .Z(n17012) );
  XOR U16339 ( .A(n17013), .B(n17014), .Z(n16980) );
  ANDN U16340 ( .B(n17015), .A(n17016), .Z(n17013) );
  XOR U16341 ( .A(n17014), .B(n17017), .Z(n17015) );
  XNOR U16342 ( .A(n17018), .B(n17019), .Z(n16977) );
  ANDN U16343 ( .B(n17020), .A(n17021), .Z(n17018) );
  XOR U16344 ( .A(n17019), .B(n17022), .Z(n17020) );
  IV U16345 ( .A(n16976), .Z(n17010) );
  XOR U16346 ( .A(n16974), .B(n17023), .Z(n16976) );
  XOR U16347 ( .A(n17024), .B(n17025), .Z(n17023) );
  ANDN U16348 ( .B(n17026), .A(n17027), .Z(n17024) );
  XOR U16349 ( .A(n17028), .B(n17025), .Z(n17026) );
  IV U16350 ( .A(n16978), .Z(n16974) );
  XOR U16351 ( .A(n17029), .B(n17030), .Z(n16978) );
  ANDN U16352 ( .B(n17031), .A(n17032), .Z(n17029) );
  XOR U16353 ( .A(n17033), .B(n17030), .Z(n17031) );
  IV U16354 ( .A(n16988), .Z(n16992) );
  XOR U16355 ( .A(n16988), .B(n16943), .Z(n16990) );
  XOR U16356 ( .A(n17034), .B(n17035), .Z(n16943) );
  AND U16357 ( .A(n478), .B(n17036), .Z(n17034) );
  XOR U16358 ( .A(n17037), .B(n17035), .Z(n17036) );
  NANDN U16359 ( .A(n16945), .B(n16947), .Z(n16988) );
  XOR U16360 ( .A(n17038), .B(n17039), .Z(n16947) );
  AND U16361 ( .A(n478), .B(n17040), .Z(n17038) );
  XOR U16362 ( .A(n17039), .B(n17041), .Z(n17040) );
  XNOR U16363 ( .A(n17042), .B(n17043), .Z(n478) );
  AND U16364 ( .A(n17044), .B(n17045), .Z(n17042) );
  XOR U16365 ( .A(n17043), .B(n16958), .Z(n17045) );
  XNOR U16366 ( .A(n17046), .B(n17047), .Z(n16958) );
  ANDN U16367 ( .B(n17048), .A(n17049), .Z(n17046) );
  XOR U16368 ( .A(n17047), .B(n17050), .Z(n17048) );
  XNOR U16369 ( .A(n17043), .B(n16960), .Z(n17044) );
  XOR U16370 ( .A(n17051), .B(n17052), .Z(n16960) );
  AND U16371 ( .A(n482), .B(n17053), .Z(n17051) );
  XOR U16372 ( .A(n17054), .B(n17052), .Z(n17053) );
  XNOR U16373 ( .A(n17055), .B(n17056), .Z(n17043) );
  AND U16374 ( .A(n17057), .B(n17058), .Z(n17055) );
  XNOR U16375 ( .A(n17056), .B(n16985), .Z(n17058) );
  XOR U16376 ( .A(n17049), .B(n17050), .Z(n16985) );
  XNOR U16377 ( .A(n17059), .B(n17060), .Z(n17050) );
  ANDN U16378 ( .B(n17061), .A(n17062), .Z(n17059) );
  XOR U16379 ( .A(n17063), .B(n17064), .Z(n17061) );
  XOR U16380 ( .A(n17065), .B(n17066), .Z(n17049) );
  XNOR U16381 ( .A(n17067), .B(n17068), .Z(n17066) );
  ANDN U16382 ( .B(n17069), .A(n17070), .Z(n17067) );
  XNOR U16383 ( .A(n17071), .B(n17072), .Z(n17069) );
  IV U16384 ( .A(n17047), .Z(n17065) );
  XOR U16385 ( .A(n17073), .B(n17074), .Z(n17047) );
  ANDN U16386 ( .B(n17075), .A(n17076), .Z(n17073) );
  XOR U16387 ( .A(n17074), .B(n17077), .Z(n17075) );
  XOR U16388 ( .A(n17056), .B(n16987), .Z(n17057) );
  XOR U16389 ( .A(n17078), .B(n17079), .Z(n16987) );
  AND U16390 ( .A(n482), .B(n17080), .Z(n17078) );
  XOR U16391 ( .A(n17081), .B(n17079), .Z(n17080) );
  XNOR U16392 ( .A(n17082), .B(n17083), .Z(n17056) );
  NAND U16393 ( .A(n17084), .B(n17085), .Z(n17083) );
  XOR U16394 ( .A(n17086), .B(n17035), .Z(n17085) );
  XOR U16395 ( .A(n17076), .B(n17077), .Z(n17035) );
  XOR U16396 ( .A(n17087), .B(n17064), .Z(n17077) );
  XOR U16397 ( .A(n17088), .B(n17089), .Z(n17064) );
  ANDN U16398 ( .B(n17090), .A(n17091), .Z(n17088) );
  XOR U16399 ( .A(n17089), .B(n17092), .Z(n17090) );
  IV U16400 ( .A(n17062), .Z(n17087) );
  XOR U16401 ( .A(n17060), .B(n17093), .Z(n17062) );
  XOR U16402 ( .A(n17094), .B(n17095), .Z(n17093) );
  ANDN U16403 ( .B(n17096), .A(n17097), .Z(n17094) );
  XOR U16404 ( .A(n17098), .B(n17095), .Z(n17096) );
  IV U16405 ( .A(n17063), .Z(n17060) );
  XOR U16406 ( .A(n17099), .B(n17100), .Z(n17063) );
  ANDN U16407 ( .B(n17101), .A(n17102), .Z(n17099) );
  XOR U16408 ( .A(n17100), .B(n17103), .Z(n17101) );
  XOR U16409 ( .A(n17104), .B(n17105), .Z(n17076) );
  XNOR U16410 ( .A(n17071), .B(n17106), .Z(n17105) );
  IV U16411 ( .A(n17074), .Z(n17106) );
  XOR U16412 ( .A(n17107), .B(n17108), .Z(n17074) );
  ANDN U16413 ( .B(n17109), .A(n17110), .Z(n17107) );
  XOR U16414 ( .A(n17108), .B(n17111), .Z(n17109) );
  XNOR U16415 ( .A(n17112), .B(n17113), .Z(n17071) );
  ANDN U16416 ( .B(n17114), .A(n17115), .Z(n17112) );
  XOR U16417 ( .A(n17113), .B(n17116), .Z(n17114) );
  IV U16418 ( .A(n17070), .Z(n17104) );
  XOR U16419 ( .A(n17068), .B(n17117), .Z(n17070) );
  XOR U16420 ( .A(n17118), .B(n17119), .Z(n17117) );
  ANDN U16421 ( .B(n17120), .A(n17121), .Z(n17118) );
  XOR U16422 ( .A(n17122), .B(n17119), .Z(n17120) );
  IV U16423 ( .A(n17072), .Z(n17068) );
  XOR U16424 ( .A(n17123), .B(n17124), .Z(n17072) );
  ANDN U16425 ( .B(n17125), .A(n17126), .Z(n17123) );
  XOR U16426 ( .A(n17127), .B(n17124), .Z(n17125) );
  IV U16427 ( .A(n17082), .Z(n17086) );
  XOR U16428 ( .A(n17082), .B(n17037), .Z(n17084) );
  XOR U16429 ( .A(n17128), .B(n17129), .Z(n17037) );
  AND U16430 ( .A(n482), .B(n17130), .Z(n17128) );
  XOR U16431 ( .A(n17131), .B(n17129), .Z(n17130) );
  NANDN U16432 ( .A(n17039), .B(n17041), .Z(n17082) );
  XOR U16433 ( .A(n17132), .B(n17133), .Z(n17041) );
  AND U16434 ( .A(n482), .B(n17134), .Z(n17132) );
  XOR U16435 ( .A(n17133), .B(n17135), .Z(n17134) );
  XNOR U16436 ( .A(n17136), .B(n17137), .Z(n482) );
  AND U16437 ( .A(n17138), .B(n17139), .Z(n17136) );
  XOR U16438 ( .A(n17137), .B(n17052), .Z(n17139) );
  XNOR U16439 ( .A(n17140), .B(n17141), .Z(n17052) );
  ANDN U16440 ( .B(n17142), .A(n17143), .Z(n17140) );
  XOR U16441 ( .A(n17141), .B(n17144), .Z(n17142) );
  XNOR U16442 ( .A(n17137), .B(n17054), .Z(n17138) );
  XOR U16443 ( .A(n17145), .B(n17146), .Z(n17054) );
  AND U16444 ( .A(n486), .B(n17147), .Z(n17145) );
  XOR U16445 ( .A(n17148), .B(n17146), .Z(n17147) );
  XNOR U16446 ( .A(n17149), .B(n17150), .Z(n17137) );
  AND U16447 ( .A(n17151), .B(n17152), .Z(n17149) );
  XNOR U16448 ( .A(n17150), .B(n17079), .Z(n17152) );
  XOR U16449 ( .A(n17143), .B(n17144), .Z(n17079) );
  XNOR U16450 ( .A(n17153), .B(n17154), .Z(n17144) );
  ANDN U16451 ( .B(n17155), .A(n17156), .Z(n17153) );
  XOR U16452 ( .A(n17157), .B(n17158), .Z(n17155) );
  XOR U16453 ( .A(n17159), .B(n17160), .Z(n17143) );
  XNOR U16454 ( .A(n17161), .B(n17162), .Z(n17160) );
  ANDN U16455 ( .B(n17163), .A(n17164), .Z(n17161) );
  XNOR U16456 ( .A(n17165), .B(n17166), .Z(n17163) );
  IV U16457 ( .A(n17141), .Z(n17159) );
  XOR U16458 ( .A(n17167), .B(n17168), .Z(n17141) );
  ANDN U16459 ( .B(n17169), .A(n17170), .Z(n17167) );
  XOR U16460 ( .A(n17168), .B(n17171), .Z(n17169) );
  XOR U16461 ( .A(n17150), .B(n17081), .Z(n17151) );
  XOR U16462 ( .A(n17172), .B(n17173), .Z(n17081) );
  AND U16463 ( .A(n486), .B(n17174), .Z(n17172) );
  XOR U16464 ( .A(n17175), .B(n17173), .Z(n17174) );
  XNOR U16465 ( .A(n17176), .B(n17177), .Z(n17150) );
  NAND U16466 ( .A(n17178), .B(n17179), .Z(n17177) );
  XOR U16467 ( .A(n17180), .B(n17129), .Z(n17179) );
  XOR U16468 ( .A(n17170), .B(n17171), .Z(n17129) );
  XOR U16469 ( .A(n17181), .B(n17158), .Z(n17171) );
  XOR U16470 ( .A(n17182), .B(n17183), .Z(n17158) );
  ANDN U16471 ( .B(n17184), .A(n17185), .Z(n17182) );
  XOR U16472 ( .A(n17183), .B(n17186), .Z(n17184) );
  IV U16473 ( .A(n17156), .Z(n17181) );
  XOR U16474 ( .A(n17154), .B(n17187), .Z(n17156) );
  XOR U16475 ( .A(n17188), .B(n17189), .Z(n17187) );
  ANDN U16476 ( .B(n17190), .A(n17191), .Z(n17188) );
  XOR U16477 ( .A(n17192), .B(n17189), .Z(n17190) );
  IV U16478 ( .A(n17157), .Z(n17154) );
  XOR U16479 ( .A(n17193), .B(n17194), .Z(n17157) );
  ANDN U16480 ( .B(n17195), .A(n17196), .Z(n17193) );
  XOR U16481 ( .A(n17194), .B(n17197), .Z(n17195) );
  XOR U16482 ( .A(n17198), .B(n17199), .Z(n17170) );
  XNOR U16483 ( .A(n17165), .B(n17200), .Z(n17199) );
  IV U16484 ( .A(n17168), .Z(n17200) );
  XOR U16485 ( .A(n17201), .B(n17202), .Z(n17168) );
  ANDN U16486 ( .B(n17203), .A(n17204), .Z(n17201) );
  XOR U16487 ( .A(n17202), .B(n17205), .Z(n17203) );
  XNOR U16488 ( .A(n17206), .B(n17207), .Z(n17165) );
  ANDN U16489 ( .B(n17208), .A(n17209), .Z(n17206) );
  XOR U16490 ( .A(n17207), .B(n17210), .Z(n17208) );
  IV U16491 ( .A(n17164), .Z(n17198) );
  XOR U16492 ( .A(n17162), .B(n17211), .Z(n17164) );
  XOR U16493 ( .A(n17212), .B(n17213), .Z(n17211) );
  ANDN U16494 ( .B(n17214), .A(n17215), .Z(n17212) );
  XOR U16495 ( .A(n17216), .B(n17213), .Z(n17214) );
  IV U16496 ( .A(n17166), .Z(n17162) );
  XOR U16497 ( .A(n17217), .B(n17218), .Z(n17166) );
  ANDN U16498 ( .B(n17219), .A(n17220), .Z(n17217) );
  XOR U16499 ( .A(n17221), .B(n17218), .Z(n17219) );
  IV U16500 ( .A(n17176), .Z(n17180) );
  XOR U16501 ( .A(n17176), .B(n17131), .Z(n17178) );
  XOR U16502 ( .A(n17222), .B(n17223), .Z(n17131) );
  AND U16503 ( .A(n486), .B(n17224), .Z(n17222) );
  XOR U16504 ( .A(n17225), .B(n17223), .Z(n17224) );
  NANDN U16505 ( .A(n17133), .B(n17135), .Z(n17176) );
  XOR U16506 ( .A(n17226), .B(n17227), .Z(n17135) );
  AND U16507 ( .A(n486), .B(n17228), .Z(n17226) );
  XOR U16508 ( .A(n17227), .B(n17229), .Z(n17228) );
  XNOR U16509 ( .A(n17230), .B(n17231), .Z(n486) );
  AND U16510 ( .A(n17232), .B(n17233), .Z(n17230) );
  XOR U16511 ( .A(n17231), .B(n17146), .Z(n17233) );
  XNOR U16512 ( .A(n17234), .B(n17235), .Z(n17146) );
  ANDN U16513 ( .B(n17236), .A(n17237), .Z(n17234) );
  XOR U16514 ( .A(n17235), .B(n17238), .Z(n17236) );
  XNOR U16515 ( .A(n17231), .B(n17148), .Z(n17232) );
  XOR U16516 ( .A(n17239), .B(n17240), .Z(n17148) );
  AND U16517 ( .A(n490), .B(n17241), .Z(n17239) );
  XOR U16518 ( .A(n17242), .B(n17240), .Z(n17241) );
  XNOR U16519 ( .A(n17243), .B(n17244), .Z(n17231) );
  AND U16520 ( .A(n17245), .B(n17246), .Z(n17243) );
  XNOR U16521 ( .A(n17244), .B(n17173), .Z(n17246) );
  XOR U16522 ( .A(n17237), .B(n17238), .Z(n17173) );
  XNOR U16523 ( .A(n17247), .B(n17248), .Z(n17238) );
  ANDN U16524 ( .B(n17249), .A(n17250), .Z(n17247) );
  XOR U16525 ( .A(n17251), .B(n17252), .Z(n17249) );
  XOR U16526 ( .A(n17253), .B(n17254), .Z(n17237) );
  XNOR U16527 ( .A(n17255), .B(n17256), .Z(n17254) );
  ANDN U16528 ( .B(n17257), .A(n17258), .Z(n17255) );
  XNOR U16529 ( .A(n17259), .B(n17260), .Z(n17257) );
  IV U16530 ( .A(n17235), .Z(n17253) );
  XOR U16531 ( .A(n17261), .B(n17262), .Z(n17235) );
  ANDN U16532 ( .B(n17263), .A(n17264), .Z(n17261) );
  XOR U16533 ( .A(n17262), .B(n17265), .Z(n17263) );
  XOR U16534 ( .A(n17244), .B(n17175), .Z(n17245) );
  XOR U16535 ( .A(n17266), .B(n17267), .Z(n17175) );
  AND U16536 ( .A(n490), .B(n17268), .Z(n17266) );
  XOR U16537 ( .A(n17269), .B(n17267), .Z(n17268) );
  XNOR U16538 ( .A(n17270), .B(n17271), .Z(n17244) );
  NAND U16539 ( .A(n17272), .B(n17273), .Z(n17271) );
  XOR U16540 ( .A(n17274), .B(n17223), .Z(n17273) );
  XOR U16541 ( .A(n17264), .B(n17265), .Z(n17223) );
  XOR U16542 ( .A(n17275), .B(n17252), .Z(n17265) );
  XOR U16543 ( .A(n17276), .B(n17277), .Z(n17252) );
  ANDN U16544 ( .B(n17278), .A(n17279), .Z(n17276) );
  XOR U16545 ( .A(n17277), .B(n17280), .Z(n17278) );
  IV U16546 ( .A(n17250), .Z(n17275) );
  XOR U16547 ( .A(n17248), .B(n17281), .Z(n17250) );
  XOR U16548 ( .A(n17282), .B(n17283), .Z(n17281) );
  ANDN U16549 ( .B(n17284), .A(n17285), .Z(n17282) );
  XOR U16550 ( .A(n17286), .B(n17283), .Z(n17284) );
  IV U16551 ( .A(n17251), .Z(n17248) );
  XOR U16552 ( .A(n17287), .B(n17288), .Z(n17251) );
  ANDN U16553 ( .B(n17289), .A(n17290), .Z(n17287) );
  XOR U16554 ( .A(n17288), .B(n17291), .Z(n17289) );
  XOR U16555 ( .A(n17292), .B(n17293), .Z(n17264) );
  XNOR U16556 ( .A(n17259), .B(n17294), .Z(n17293) );
  IV U16557 ( .A(n17262), .Z(n17294) );
  XOR U16558 ( .A(n17295), .B(n17296), .Z(n17262) );
  ANDN U16559 ( .B(n17297), .A(n17298), .Z(n17295) );
  XOR U16560 ( .A(n17296), .B(n17299), .Z(n17297) );
  XNOR U16561 ( .A(n17300), .B(n17301), .Z(n17259) );
  ANDN U16562 ( .B(n17302), .A(n17303), .Z(n17300) );
  XOR U16563 ( .A(n17301), .B(n17304), .Z(n17302) );
  IV U16564 ( .A(n17258), .Z(n17292) );
  XOR U16565 ( .A(n17256), .B(n17305), .Z(n17258) );
  XOR U16566 ( .A(n17306), .B(n17307), .Z(n17305) );
  ANDN U16567 ( .B(n17308), .A(n17309), .Z(n17306) );
  XOR U16568 ( .A(n17310), .B(n17307), .Z(n17308) );
  IV U16569 ( .A(n17260), .Z(n17256) );
  XOR U16570 ( .A(n17311), .B(n17312), .Z(n17260) );
  ANDN U16571 ( .B(n17313), .A(n17314), .Z(n17311) );
  XOR U16572 ( .A(n17315), .B(n17312), .Z(n17313) );
  IV U16573 ( .A(n17270), .Z(n17274) );
  XOR U16574 ( .A(n17270), .B(n17225), .Z(n17272) );
  XOR U16575 ( .A(n17316), .B(n17317), .Z(n17225) );
  AND U16576 ( .A(n490), .B(n17318), .Z(n17316) );
  XOR U16577 ( .A(n17319), .B(n17317), .Z(n17318) );
  NANDN U16578 ( .A(n17227), .B(n17229), .Z(n17270) );
  XOR U16579 ( .A(n17320), .B(n17321), .Z(n17229) );
  AND U16580 ( .A(n490), .B(n17322), .Z(n17320) );
  XOR U16581 ( .A(n17321), .B(n17323), .Z(n17322) );
  XNOR U16582 ( .A(n17324), .B(n17325), .Z(n490) );
  AND U16583 ( .A(n17326), .B(n17327), .Z(n17324) );
  XOR U16584 ( .A(n17325), .B(n17240), .Z(n17327) );
  XNOR U16585 ( .A(n17328), .B(n17329), .Z(n17240) );
  ANDN U16586 ( .B(n17330), .A(n17331), .Z(n17328) );
  XOR U16587 ( .A(n17329), .B(n17332), .Z(n17330) );
  XNOR U16588 ( .A(n17325), .B(n17242), .Z(n17326) );
  XOR U16589 ( .A(n17333), .B(n17334), .Z(n17242) );
  AND U16590 ( .A(n494), .B(n17335), .Z(n17333) );
  XOR U16591 ( .A(n17336), .B(n17334), .Z(n17335) );
  XNOR U16592 ( .A(n17337), .B(n17338), .Z(n17325) );
  AND U16593 ( .A(n17339), .B(n17340), .Z(n17337) );
  XNOR U16594 ( .A(n17338), .B(n17267), .Z(n17340) );
  XOR U16595 ( .A(n17331), .B(n17332), .Z(n17267) );
  XNOR U16596 ( .A(n17341), .B(n17342), .Z(n17332) );
  ANDN U16597 ( .B(n17343), .A(n17344), .Z(n17341) );
  XOR U16598 ( .A(n17345), .B(n17346), .Z(n17343) );
  XOR U16599 ( .A(n17347), .B(n17348), .Z(n17331) );
  XNOR U16600 ( .A(n17349), .B(n17350), .Z(n17348) );
  ANDN U16601 ( .B(n17351), .A(n17352), .Z(n17349) );
  XNOR U16602 ( .A(n17353), .B(n17354), .Z(n17351) );
  IV U16603 ( .A(n17329), .Z(n17347) );
  XOR U16604 ( .A(n17355), .B(n17356), .Z(n17329) );
  ANDN U16605 ( .B(n17357), .A(n17358), .Z(n17355) );
  XOR U16606 ( .A(n17356), .B(n17359), .Z(n17357) );
  XOR U16607 ( .A(n17338), .B(n17269), .Z(n17339) );
  XOR U16608 ( .A(n17360), .B(n17361), .Z(n17269) );
  AND U16609 ( .A(n494), .B(n17362), .Z(n17360) );
  XOR U16610 ( .A(n17363), .B(n17361), .Z(n17362) );
  XNOR U16611 ( .A(n17364), .B(n17365), .Z(n17338) );
  NAND U16612 ( .A(n17366), .B(n17367), .Z(n17365) );
  XOR U16613 ( .A(n17368), .B(n17317), .Z(n17367) );
  XOR U16614 ( .A(n17358), .B(n17359), .Z(n17317) );
  XOR U16615 ( .A(n17369), .B(n17346), .Z(n17359) );
  XOR U16616 ( .A(n17370), .B(n17371), .Z(n17346) );
  ANDN U16617 ( .B(n17372), .A(n17373), .Z(n17370) );
  XOR U16618 ( .A(n17371), .B(n17374), .Z(n17372) );
  IV U16619 ( .A(n17344), .Z(n17369) );
  XOR U16620 ( .A(n17342), .B(n17375), .Z(n17344) );
  XOR U16621 ( .A(n17376), .B(n17377), .Z(n17375) );
  ANDN U16622 ( .B(n17378), .A(n17379), .Z(n17376) );
  XOR U16623 ( .A(n17380), .B(n17377), .Z(n17378) );
  IV U16624 ( .A(n17345), .Z(n17342) );
  XOR U16625 ( .A(n17381), .B(n17382), .Z(n17345) );
  ANDN U16626 ( .B(n17383), .A(n17384), .Z(n17381) );
  XOR U16627 ( .A(n17382), .B(n17385), .Z(n17383) );
  XOR U16628 ( .A(n17386), .B(n17387), .Z(n17358) );
  XNOR U16629 ( .A(n17353), .B(n17388), .Z(n17387) );
  IV U16630 ( .A(n17356), .Z(n17388) );
  XOR U16631 ( .A(n17389), .B(n17390), .Z(n17356) );
  ANDN U16632 ( .B(n17391), .A(n17392), .Z(n17389) );
  XOR U16633 ( .A(n17390), .B(n17393), .Z(n17391) );
  XNOR U16634 ( .A(n17394), .B(n17395), .Z(n17353) );
  ANDN U16635 ( .B(n17396), .A(n17397), .Z(n17394) );
  XOR U16636 ( .A(n17395), .B(n17398), .Z(n17396) );
  IV U16637 ( .A(n17352), .Z(n17386) );
  XOR U16638 ( .A(n17350), .B(n17399), .Z(n17352) );
  XOR U16639 ( .A(n17400), .B(n17401), .Z(n17399) );
  ANDN U16640 ( .B(n17402), .A(n17403), .Z(n17400) );
  XOR U16641 ( .A(n17404), .B(n17401), .Z(n17402) );
  IV U16642 ( .A(n17354), .Z(n17350) );
  XOR U16643 ( .A(n17405), .B(n17406), .Z(n17354) );
  ANDN U16644 ( .B(n17407), .A(n17408), .Z(n17405) );
  XOR U16645 ( .A(n17409), .B(n17406), .Z(n17407) );
  IV U16646 ( .A(n17364), .Z(n17368) );
  XOR U16647 ( .A(n17364), .B(n17319), .Z(n17366) );
  XOR U16648 ( .A(n17410), .B(n17411), .Z(n17319) );
  AND U16649 ( .A(n494), .B(n17412), .Z(n17410) );
  XOR U16650 ( .A(n17413), .B(n17411), .Z(n17412) );
  NANDN U16651 ( .A(n17321), .B(n17323), .Z(n17364) );
  XOR U16652 ( .A(n17414), .B(n17415), .Z(n17323) );
  AND U16653 ( .A(n494), .B(n17416), .Z(n17414) );
  XOR U16654 ( .A(n17415), .B(n17417), .Z(n17416) );
  XNOR U16655 ( .A(n17418), .B(n17419), .Z(n494) );
  AND U16656 ( .A(n17420), .B(n17421), .Z(n17418) );
  XOR U16657 ( .A(n17419), .B(n17334), .Z(n17421) );
  XNOR U16658 ( .A(n17422), .B(n17423), .Z(n17334) );
  ANDN U16659 ( .B(n17424), .A(n17425), .Z(n17422) );
  XOR U16660 ( .A(n17423), .B(n17426), .Z(n17424) );
  XNOR U16661 ( .A(n17419), .B(n17336), .Z(n17420) );
  XOR U16662 ( .A(n17427), .B(n17428), .Z(n17336) );
  AND U16663 ( .A(n498), .B(n17429), .Z(n17427) );
  XOR U16664 ( .A(n17430), .B(n17428), .Z(n17429) );
  XNOR U16665 ( .A(n17431), .B(n17432), .Z(n17419) );
  AND U16666 ( .A(n17433), .B(n17434), .Z(n17431) );
  XNOR U16667 ( .A(n17432), .B(n17361), .Z(n17434) );
  XOR U16668 ( .A(n17425), .B(n17426), .Z(n17361) );
  XNOR U16669 ( .A(n17435), .B(n17436), .Z(n17426) );
  ANDN U16670 ( .B(n17437), .A(n17438), .Z(n17435) );
  XOR U16671 ( .A(n17439), .B(n17440), .Z(n17437) );
  XOR U16672 ( .A(n17441), .B(n17442), .Z(n17425) );
  XNOR U16673 ( .A(n17443), .B(n17444), .Z(n17442) );
  ANDN U16674 ( .B(n17445), .A(n17446), .Z(n17443) );
  XNOR U16675 ( .A(n17447), .B(n17448), .Z(n17445) );
  IV U16676 ( .A(n17423), .Z(n17441) );
  XOR U16677 ( .A(n17449), .B(n17450), .Z(n17423) );
  ANDN U16678 ( .B(n17451), .A(n17452), .Z(n17449) );
  XOR U16679 ( .A(n17450), .B(n17453), .Z(n17451) );
  XOR U16680 ( .A(n17432), .B(n17363), .Z(n17433) );
  XOR U16681 ( .A(n17454), .B(n17455), .Z(n17363) );
  AND U16682 ( .A(n498), .B(n17456), .Z(n17454) );
  XOR U16683 ( .A(n17457), .B(n17455), .Z(n17456) );
  XNOR U16684 ( .A(n17458), .B(n17459), .Z(n17432) );
  NAND U16685 ( .A(n17460), .B(n17461), .Z(n17459) );
  XOR U16686 ( .A(n17462), .B(n17411), .Z(n17461) );
  XOR U16687 ( .A(n17452), .B(n17453), .Z(n17411) );
  XOR U16688 ( .A(n17463), .B(n17440), .Z(n17453) );
  XOR U16689 ( .A(n17464), .B(n17465), .Z(n17440) );
  ANDN U16690 ( .B(n17466), .A(n17467), .Z(n17464) );
  XOR U16691 ( .A(n17465), .B(n17468), .Z(n17466) );
  IV U16692 ( .A(n17438), .Z(n17463) );
  XOR U16693 ( .A(n17436), .B(n17469), .Z(n17438) );
  XOR U16694 ( .A(n17470), .B(n17471), .Z(n17469) );
  ANDN U16695 ( .B(n17472), .A(n17473), .Z(n17470) );
  XOR U16696 ( .A(n17474), .B(n17471), .Z(n17472) );
  IV U16697 ( .A(n17439), .Z(n17436) );
  XOR U16698 ( .A(n17475), .B(n17476), .Z(n17439) );
  ANDN U16699 ( .B(n17477), .A(n17478), .Z(n17475) );
  XOR U16700 ( .A(n17476), .B(n17479), .Z(n17477) );
  XOR U16701 ( .A(n17480), .B(n17481), .Z(n17452) );
  XNOR U16702 ( .A(n17447), .B(n17482), .Z(n17481) );
  IV U16703 ( .A(n17450), .Z(n17482) );
  XOR U16704 ( .A(n17483), .B(n17484), .Z(n17450) );
  ANDN U16705 ( .B(n17485), .A(n17486), .Z(n17483) );
  XOR U16706 ( .A(n17484), .B(n17487), .Z(n17485) );
  XNOR U16707 ( .A(n17488), .B(n17489), .Z(n17447) );
  ANDN U16708 ( .B(n17490), .A(n17491), .Z(n17488) );
  XOR U16709 ( .A(n17489), .B(n17492), .Z(n17490) );
  IV U16710 ( .A(n17446), .Z(n17480) );
  XOR U16711 ( .A(n17444), .B(n17493), .Z(n17446) );
  XOR U16712 ( .A(n17494), .B(n17495), .Z(n17493) );
  ANDN U16713 ( .B(n17496), .A(n17497), .Z(n17494) );
  XOR U16714 ( .A(n17498), .B(n17495), .Z(n17496) );
  IV U16715 ( .A(n17448), .Z(n17444) );
  XOR U16716 ( .A(n17499), .B(n17500), .Z(n17448) );
  ANDN U16717 ( .B(n17501), .A(n17502), .Z(n17499) );
  XOR U16718 ( .A(n17503), .B(n17500), .Z(n17501) );
  IV U16719 ( .A(n17458), .Z(n17462) );
  XOR U16720 ( .A(n17458), .B(n17413), .Z(n17460) );
  XOR U16721 ( .A(n17504), .B(n17505), .Z(n17413) );
  AND U16722 ( .A(n498), .B(n17506), .Z(n17504) );
  XOR U16723 ( .A(n17507), .B(n17505), .Z(n17506) );
  NANDN U16724 ( .A(n17415), .B(n17417), .Z(n17458) );
  XOR U16725 ( .A(n17508), .B(n17509), .Z(n17417) );
  AND U16726 ( .A(n498), .B(n17510), .Z(n17508) );
  XOR U16727 ( .A(n17509), .B(n17511), .Z(n17510) );
  XNOR U16728 ( .A(n17512), .B(n17513), .Z(n498) );
  AND U16729 ( .A(n17514), .B(n17515), .Z(n17512) );
  XOR U16730 ( .A(n17513), .B(n17428), .Z(n17515) );
  XNOR U16731 ( .A(n17516), .B(n17517), .Z(n17428) );
  ANDN U16732 ( .B(n17518), .A(n17519), .Z(n17516) );
  XOR U16733 ( .A(n17517), .B(n17520), .Z(n17518) );
  XNOR U16734 ( .A(n17513), .B(n17430), .Z(n17514) );
  XOR U16735 ( .A(n17521), .B(n17522), .Z(n17430) );
  AND U16736 ( .A(n502), .B(n17523), .Z(n17521) );
  XOR U16737 ( .A(n17524), .B(n17522), .Z(n17523) );
  XNOR U16738 ( .A(n17525), .B(n17526), .Z(n17513) );
  AND U16739 ( .A(n17527), .B(n17528), .Z(n17525) );
  XNOR U16740 ( .A(n17526), .B(n17455), .Z(n17528) );
  XOR U16741 ( .A(n17519), .B(n17520), .Z(n17455) );
  XNOR U16742 ( .A(n17529), .B(n17530), .Z(n17520) );
  ANDN U16743 ( .B(n17531), .A(n17532), .Z(n17529) );
  XOR U16744 ( .A(n17533), .B(n17534), .Z(n17531) );
  XOR U16745 ( .A(n17535), .B(n17536), .Z(n17519) );
  XNOR U16746 ( .A(n17537), .B(n17538), .Z(n17536) );
  ANDN U16747 ( .B(n17539), .A(n17540), .Z(n17537) );
  XNOR U16748 ( .A(n17541), .B(n17542), .Z(n17539) );
  IV U16749 ( .A(n17517), .Z(n17535) );
  XOR U16750 ( .A(n17543), .B(n17544), .Z(n17517) );
  ANDN U16751 ( .B(n17545), .A(n17546), .Z(n17543) );
  XOR U16752 ( .A(n17544), .B(n17547), .Z(n17545) );
  XOR U16753 ( .A(n17526), .B(n17457), .Z(n17527) );
  XOR U16754 ( .A(n17548), .B(n17549), .Z(n17457) );
  AND U16755 ( .A(n502), .B(n17550), .Z(n17548) );
  XOR U16756 ( .A(n17551), .B(n17549), .Z(n17550) );
  XNOR U16757 ( .A(n17552), .B(n17553), .Z(n17526) );
  NAND U16758 ( .A(n17554), .B(n17555), .Z(n17553) );
  XOR U16759 ( .A(n17556), .B(n17505), .Z(n17555) );
  XOR U16760 ( .A(n17546), .B(n17547), .Z(n17505) );
  XOR U16761 ( .A(n17557), .B(n17534), .Z(n17547) );
  XOR U16762 ( .A(n17558), .B(n17559), .Z(n17534) );
  ANDN U16763 ( .B(n17560), .A(n17561), .Z(n17558) );
  XOR U16764 ( .A(n17559), .B(n17562), .Z(n17560) );
  IV U16765 ( .A(n17532), .Z(n17557) );
  XOR U16766 ( .A(n17530), .B(n17563), .Z(n17532) );
  XOR U16767 ( .A(n17564), .B(n17565), .Z(n17563) );
  ANDN U16768 ( .B(n17566), .A(n17567), .Z(n17564) );
  XOR U16769 ( .A(n17568), .B(n17565), .Z(n17566) );
  IV U16770 ( .A(n17533), .Z(n17530) );
  XOR U16771 ( .A(n17569), .B(n17570), .Z(n17533) );
  ANDN U16772 ( .B(n17571), .A(n17572), .Z(n17569) );
  XOR U16773 ( .A(n17570), .B(n17573), .Z(n17571) );
  XOR U16774 ( .A(n17574), .B(n17575), .Z(n17546) );
  XNOR U16775 ( .A(n17541), .B(n17576), .Z(n17575) );
  IV U16776 ( .A(n17544), .Z(n17576) );
  XOR U16777 ( .A(n17577), .B(n17578), .Z(n17544) );
  ANDN U16778 ( .B(n17579), .A(n17580), .Z(n17577) );
  XOR U16779 ( .A(n17578), .B(n17581), .Z(n17579) );
  XNOR U16780 ( .A(n17582), .B(n17583), .Z(n17541) );
  ANDN U16781 ( .B(n17584), .A(n17585), .Z(n17582) );
  XOR U16782 ( .A(n17583), .B(n17586), .Z(n17584) );
  IV U16783 ( .A(n17540), .Z(n17574) );
  XOR U16784 ( .A(n17538), .B(n17587), .Z(n17540) );
  XOR U16785 ( .A(n17588), .B(n17589), .Z(n17587) );
  ANDN U16786 ( .B(n17590), .A(n17591), .Z(n17588) );
  XOR U16787 ( .A(n17592), .B(n17589), .Z(n17590) );
  IV U16788 ( .A(n17542), .Z(n17538) );
  XOR U16789 ( .A(n17593), .B(n17594), .Z(n17542) );
  ANDN U16790 ( .B(n17595), .A(n17596), .Z(n17593) );
  XOR U16791 ( .A(n17597), .B(n17594), .Z(n17595) );
  IV U16792 ( .A(n17552), .Z(n17556) );
  XOR U16793 ( .A(n17552), .B(n17507), .Z(n17554) );
  XOR U16794 ( .A(n17598), .B(n17599), .Z(n17507) );
  AND U16795 ( .A(n502), .B(n17600), .Z(n17598) );
  XOR U16796 ( .A(n17601), .B(n17599), .Z(n17600) );
  NANDN U16797 ( .A(n17509), .B(n17511), .Z(n17552) );
  XOR U16798 ( .A(n17602), .B(n17603), .Z(n17511) );
  AND U16799 ( .A(n502), .B(n17604), .Z(n17602) );
  XOR U16800 ( .A(n17603), .B(n17605), .Z(n17604) );
  XNOR U16801 ( .A(n17606), .B(n17607), .Z(n502) );
  AND U16802 ( .A(n17608), .B(n17609), .Z(n17606) );
  XOR U16803 ( .A(n17607), .B(n17522), .Z(n17609) );
  XNOR U16804 ( .A(n17610), .B(n17611), .Z(n17522) );
  ANDN U16805 ( .B(n17612), .A(n17613), .Z(n17610) );
  XOR U16806 ( .A(n17611), .B(n17614), .Z(n17612) );
  XNOR U16807 ( .A(n17607), .B(n17524), .Z(n17608) );
  XOR U16808 ( .A(n17615), .B(n17616), .Z(n17524) );
  AND U16809 ( .A(n506), .B(n17617), .Z(n17615) );
  XOR U16810 ( .A(n17618), .B(n17616), .Z(n17617) );
  XNOR U16811 ( .A(n17619), .B(n17620), .Z(n17607) );
  AND U16812 ( .A(n17621), .B(n17622), .Z(n17619) );
  XNOR U16813 ( .A(n17620), .B(n17549), .Z(n17622) );
  XOR U16814 ( .A(n17613), .B(n17614), .Z(n17549) );
  XNOR U16815 ( .A(n17623), .B(n17624), .Z(n17614) );
  ANDN U16816 ( .B(n17625), .A(n17626), .Z(n17623) );
  XOR U16817 ( .A(n17627), .B(n17628), .Z(n17625) );
  XOR U16818 ( .A(n17629), .B(n17630), .Z(n17613) );
  XNOR U16819 ( .A(n17631), .B(n17632), .Z(n17630) );
  ANDN U16820 ( .B(n17633), .A(n17634), .Z(n17631) );
  XNOR U16821 ( .A(n17635), .B(n17636), .Z(n17633) );
  IV U16822 ( .A(n17611), .Z(n17629) );
  XOR U16823 ( .A(n17637), .B(n17638), .Z(n17611) );
  ANDN U16824 ( .B(n17639), .A(n17640), .Z(n17637) );
  XOR U16825 ( .A(n17638), .B(n17641), .Z(n17639) );
  XOR U16826 ( .A(n17620), .B(n17551), .Z(n17621) );
  XOR U16827 ( .A(n17642), .B(n17643), .Z(n17551) );
  AND U16828 ( .A(n506), .B(n17644), .Z(n17642) );
  XNOR U16829 ( .A(n17645), .B(n17643), .Z(n17644) );
  XNOR U16830 ( .A(n17646), .B(n17647), .Z(n17620) );
  NAND U16831 ( .A(n17648), .B(n17649), .Z(n17647) );
  XOR U16832 ( .A(n17650), .B(n17599), .Z(n17649) );
  XOR U16833 ( .A(n17640), .B(n17641), .Z(n17599) );
  XOR U16834 ( .A(n17651), .B(n17628), .Z(n17641) );
  XOR U16835 ( .A(n17652), .B(n17653), .Z(n17628) );
  ANDN U16836 ( .B(n17654), .A(n17655), .Z(n17652) );
  XOR U16837 ( .A(n17653), .B(n17656), .Z(n17654) );
  IV U16838 ( .A(n17626), .Z(n17651) );
  XOR U16839 ( .A(n17624), .B(n17657), .Z(n17626) );
  XOR U16840 ( .A(n17658), .B(n17659), .Z(n17657) );
  ANDN U16841 ( .B(n17660), .A(n17661), .Z(n17658) );
  XOR U16842 ( .A(n17662), .B(n17659), .Z(n17660) );
  IV U16843 ( .A(n17627), .Z(n17624) );
  XOR U16844 ( .A(n17663), .B(n17664), .Z(n17627) );
  ANDN U16845 ( .B(n17665), .A(n17666), .Z(n17663) );
  XOR U16846 ( .A(n17664), .B(n17667), .Z(n17665) );
  XOR U16847 ( .A(n17668), .B(n17669), .Z(n17640) );
  XNOR U16848 ( .A(n17635), .B(n17670), .Z(n17669) );
  IV U16849 ( .A(n17638), .Z(n17670) );
  XOR U16850 ( .A(n17671), .B(n17672), .Z(n17638) );
  ANDN U16851 ( .B(n17673), .A(n17674), .Z(n17671) );
  XOR U16852 ( .A(n17672), .B(n17675), .Z(n17673) );
  XNOR U16853 ( .A(n17676), .B(n17677), .Z(n17635) );
  ANDN U16854 ( .B(n17678), .A(n17679), .Z(n17676) );
  XOR U16855 ( .A(n17677), .B(n17680), .Z(n17678) );
  IV U16856 ( .A(n17634), .Z(n17668) );
  XOR U16857 ( .A(n17632), .B(n17681), .Z(n17634) );
  XOR U16858 ( .A(n17682), .B(n17683), .Z(n17681) );
  ANDN U16859 ( .B(n17684), .A(n17685), .Z(n17682) );
  XOR U16860 ( .A(n17686), .B(n17683), .Z(n17684) );
  IV U16861 ( .A(n17636), .Z(n17632) );
  XOR U16862 ( .A(n17687), .B(n17688), .Z(n17636) );
  ANDN U16863 ( .B(n17689), .A(n17690), .Z(n17687) );
  XOR U16864 ( .A(n17691), .B(n17688), .Z(n17689) );
  IV U16865 ( .A(n17646), .Z(n17650) );
  XOR U16866 ( .A(n17646), .B(n17601), .Z(n17648) );
  XOR U16867 ( .A(n17692), .B(n17693), .Z(n17601) );
  AND U16868 ( .A(n506), .B(n17694), .Z(n17692) );
  XNOR U16869 ( .A(n17695), .B(n17693), .Z(n17694) );
  NANDN U16870 ( .A(n17603), .B(n17605), .Z(n17646) );
  XOR U16871 ( .A(n17696), .B(n17697), .Z(n17605) );
  AND U16872 ( .A(n506), .B(n17698), .Z(n17696) );
  XOR U16873 ( .A(n17697), .B(n17699), .Z(n17698) );
  XNOR U16874 ( .A(n17700), .B(n17701), .Z(n506) );
  AND U16875 ( .A(n17702), .B(n17703), .Z(n17700) );
  XOR U16876 ( .A(n17701), .B(n17616), .Z(n17703) );
  XNOR U16877 ( .A(n17704), .B(n17705), .Z(n17616) );
  ANDN U16878 ( .B(n17706), .A(n17707), .Z(n17704) );
  XOR U16879 ( .A(n17705), .B(n17708), .Z(n17706) );
  XNOR U16880 ( .A(n17701), .B(n17618), .Z(n17702) );
  XNOR U16881 ( .A(n17709), .B(n17710), .Z(n17618) );
  ANDN U16882 ( .B(n17711), .A(n17712), .Z(n17709) );
  XOR U16883 ( .A(n17710), .B(n17713), .Z(n17711) );
  XNOR U16884 ( .A(n17714), .B(n17715), .Z(n17701) );
  AND U16885 ( .A(n17716), .B(n17717), .Z(n17714) );
  XNOR U16886 ( .A(n17715), .B(n17643), .Z(n17717) );
  XOR U16887 ( .A(n17707), .B(n17708), .Z(n17643) );
  XNOR U16888 ( .A(n17718), .B(n17719), .Z(n17708) );
  ANDN U16889 ( .B(n17720), .A(n17721), .Z(n17718) );
  XOR U16890 ( .A(n17722), .B(n17723), .Z(n17720) );
  XOR U16891 ( .A(n17724), .B(n17725), .Z(n17707) );
  XNOR U16892 ( .A(n17726), .B(n17727), .Z(n17725) );
  ANDN U16893 ( .B(n17728), .A(n17729), .Z(n17726) );
  XNOR U16894 ( .A(n17730), .B(n17731), .Z(n17728) );
  IV U16895 ( .A(n17705), .Z(n17724) );
  XOR U16896 ( .A(n17732), .B(n17733), .Z(n17705) );
  ANDN U16897 ( .B(n17734), .A(n17735), .Z(n17732) );
  XOR U16898 ( .A(n17733), .B(n17736), .Z(n17734) );
  XNOR U16899 ( .A(n17715), .B(n17645), .Z(n17716) );
  XOR U16900 ( .A(n17737), .B(n17713), .Z(n17645) );
  XNOR U16901 ( .A(n17738), .B(n17739), .Z(n17713) );
  ANDN U16902 ( .B(n17740), .A(n17741), .Z(n17738) );
  XOR U16903 ( .A(n17742), .B(n17743), .Z(n17740) );
  IV U16904 ( .A(n17712), .Z(n17737) );
  XOR U16905 ( .A(n17744), .B(n17745), .Z(n17712) );
  XNOR U16906 ( .A(n17746), .B(n17747), .Z(n17745) );
  ANDN U16907 ( .B(n17748), .A(n17749), .Z(n17746) );
  XNOR U16908 ( .A(n17750), .B(n17751), .Z(n17748) );
  IV U16909 ( .A(n17710), .Z(n17744) );
  XOR U16910 ( .A(n17752), .B(n17753), .Z(n17710) );
  ANDN U16911 ( .B(n17754), .A(n17755), .Z(n17752) );
  XOR U16912 ( .A(n17753), .B(n17756), .Z(n17754) );
  XNOR U16913 ( .A(n17757), .B(n17758), .Z(n17715) );
  NAND U16914 ( .A(n17759), .B(n17760), .Z(n17758) );
  XOR U16915 ( .A(n17761), .B(n17693), .Z(n17760) );
  XOR U16916 ( .A(n17735), .B(n17736), .Z(n17693) );
  XOR U16917 ( .A(n17762), .B(n17723), .Z(n17736) );
  XOR U16918 ( .A(n17763), .B(n17764), .Z(n17723) );
  ANDN U16919 ( .B(n17765), .A(n17766), .Z(n17763) );
  XOR U16920 ( .A(n17764), .B(n17767), .Z(n17765) );
  IV U16921 ( .A(n17721), .Z(n17762) );
  XOR U16922 ( .A(n17719), .B(n17768), .Z(n17721) );
  XOR U16923 ( .A(n17769), .B(n17770), .Z(n17768) );
  ANDN U16924 ( .B(n17771), .A(n17772), .Z(n17769) );
  XOR U16925 ( .A(n17773), .B(n17770), .Z(n17771) );
  IV U16926 ( .A(n17722), .Z(n17719) );
  XOR U16927 ( .A(n17774), .B(n17775), .Z(n17722) );
  ANDN U16928 ( .B(n17776), .A(n17777), .Z(n17774) );
  XOR U16929 ( .A(n17775), .B(n17778), .Z(n17776) );
  XOR U16930 ( .A(n17779), .B(n17780), .Z(n17735) );
  XNOR U16931 ( .A(n17730), .B(n17781), .Z(n17780) );
  IV U16932 ( .A(n17733), .Z(n17781) );
  XOR U16933 ( .A(n17782), .B(n17783), .Z(n17733) );
  ANDN U16934 ( .B(n17784), .A(n17785), .Z(n17782) );
  XOR U16935 ( .A(n17783), .B(n17786), .Z(n17784) );
  XNOR U16936 ( .A(n17787), .B(n17788), .Z(n17730) );
  ANDN U16937 ( .B(n17789), .A(n17790), .Z(n17787) );
  XOR U16938 ( .A(n17788), .B(n17791), .Z(n17789) );
  IV U16939 ( .A(n17729), .Z(n17779) );
  XOR U16940 ( .A(n17727), .B(n17792), .Z(n17729) );
  XOR U16941 ( .A(n17793), .B(n17794), .Z(n17792) );
  ANDN U16942 ( .B(n17795), .A(n17796), .Z(n17793) );
  XOR U16943 ( .A(n17797), .B(n17794), .Z(n17795) );
  IV U16944 ( .A(n17731), .Z(n17727) );
  XOR U16945 ( .A(n17798), .B(n17799), .Z(n17731) );
  ANDN U16946 ( .B(n17800), .A(n17801), .Z(n17798) );
  XOR U16947 ( .A(n17802), .B(n17799), .Z(n17800) );
  IV U16948 ( .A(n17757), .Z(n17761) );
  XNOR U16949 ( .A(n17757), .B(n17695), .Z(n17759) );
  XOR U16950 ( .A(n17803), .B(n17756), .Z(n17695) );
  XOR U16951 ( .A(n17804), .B(n17743), .Z(n17756) );
  XOR U16952 ( .A(n17805), .B(n17806), .Z(n17743) );
  ANDN U16953 ( .B(n17807), .A(n17808), .Z(n17805) );
  XOR U16954 ( .A(n17806), .B(n17809), .Z(n17807) );
  IV U16955 ( .A(n17741), .Z(n17804) );
  XOR U16956 ( .A(n17739), .B(n17810), .Z(n17741) );
  XOR U16957 ( .A(n17811), .B(n17812), .Z(n17810) );
  ANDN U16958 ( .B(n17813), .A(n17814), .Z(n17811) );
  XOR U16959 ( .A(n17815), .B(n17812), .Z(n17813) );
  IV U16960 ( .A(n17742), .Z(n17739) );
  XOR U16961 ( .A(n17816), .B(n17817), .Z(n17742) );
  ANDN U16962 ( .B(n17818), .A(n17819), .Z(n17816) );
  XOR U16963 ( .A(n17817), .B(n17820), .Z(n17818) );
  IV U16964 ( .A(n17755), .Z(n17803) );
  XOR U16965 ( .A(n17821), .B(n17822), .Z(n17755) );
  XNOR U16966 ( .A(n17750), .B(n17823), .Z(n17822) );
  IV U16967 ( .A(n17753), .Z(n17823) );
  XNOR U16968 ( .A(n17824), .B(n17825), .Z(n17753) );
  ANDN U16969 ( .B(n17826), .A(n17827), .Z(n17824) );
  XNOR U16970 ( .A(n17825), .B(n17828), .Z(n17826) );
  XNOR U16971 ( .A(n17829), .B(n17830), .Z(n17750) );
  ANDN U16972 ( .B(n17831), .A(n17832), .Z(n17829) );
  XOR U16973 ( .A(n17830), .B(n17833), .Z(n17831) );
  IV U16974 ( .A(n17749), .Z(n17821) );
  XOR U16975 ( .A(n17747), .B(n17834), .Z(n17749) );
  XOR U16976 ( .A(n17835), .B(n17836), .Z(n17834) );
  ANDN U16977 ( .B(n17837), .A(n17838), .Z(n17835) );
  XOR U16978 ( .A(n17839), .B(n17836), .Z(n17837) );
  IV U16979 ( .A(n17751), .Z(n17747) );
  XOR U16980 ( .A(n17840), .B(n17841), .Z(n17751) );
  ANDN U16981 ( .B(n17842), .A(n17843), .Z(n17840) );
  XOR U16982 ( .A(n17844), .B(n17841), .Z(n17842) );
  NANDN U16983 ( .A(n17697), .B(n17699), .Z(n17757) );
  XOR U16984 ( .A(n17845), .B(n17828), .Z(n17699) );
  XOR U16985 ( .A(n17846), .B(n17820), .Z(n17828) );
  XOR U16986 ( .A(n17847), .B(n17809), .Z(n17820) );
  XNOR U16987 ( .A(q[14]), .B(DB[14]), .Z(n17809) );
  IV U16988 ( .A(n17808), .Z(n17847) );
  XNOR U16989 ( .A(n17806), .B(n17848), .Z(n17808) );
  XNOR U16990 ( .A(q[13]), .B(DB[13]), .Z(n17848) );
  XNOR U16991 ( .A(q[12]), .B(DB[12]), .Z(n17806) );
  IV U16992 ( .A(n17819), .Z(n17846) );
  XOR U16993 ( .A(n17849), .B(n17850), .Z(n17819) );
  XNOR U16994 ( .A(n17815), .B(n17817), .Z(n17850) );
  XNOR U16995 ( .A(q[8]), .B(DB[8]), .Z(n17817) );
  XNOR U16996 ( .A(q[11]), .B(DB[11]), .Z(n17815) );
  IV U16997 ( .A(n17814), .Z(n17849) );
  XNOR U16998 ( .A(n17812), .B(n17851), .Z(n17814) );
  XNOR U16999 ( .A(q[10]), .B(DB[10]), .Z(n17851) );
  XNOR U17000 ( .A(q[9]), .B(DB[9]), .Z(n17812) );
  IV U17001 ( .A(n17827), .Z(n17845) );
  XOR U17002 ( .A(n17852), .B(n17853), .Z(n17827) );
  XOR U17003 ( .A(n17825), .B(n17844), .Z(n17853) );
  XOR U17004 ( .A(n17854), .B(n17833), .Z(n17844) );
  XNOR U17005 ( .A(q[7]), .B(DB[7]), .Z(n17833) );
  IV U17006 ( .A(n17832), .Z(n17854) );
  XNOR U17007 ( .A(n17830), .B(n17855), .Z(n17832) );
  XNOR U17008 ( .A(q[6]), .B(DB[6]), .Z(n17855) );
  XNOR U17009 ( .A(q[5]), .B(DB[5]), .Z(n17830) );
  XOR U17010 ( .A(q[0]), .B(DB[0]), .Z(n17825) );
  IV U17011 ( .A(n17843), .Z(n17852) );
  XOR U17012 ( .A(n17856), .B(n17857), .Z(n17843) );
  XNOR U17013 ( .A(n17839), .B(n17841), .Z(n17857) );
  XNOR U17014 ( .A(q[1]), .B(DB[1]), .Z(n17841) );
  XNOR U17015 ( .A(q[4]), .B(DB[4]), .Z(n17839) );
  IV U17016 ( .A(n17838), .Z(n17856) );
  XNOR U17017 ( .A(n17836), .B(n17858), .Z(n17838) );
  XNOR U17018 ( .A(q[3]), .B(DB[3]), .Z(n17858) );
  XNOR U17019 ( .A(q[2]), .B(DB[2]), .Z(n17836) );
  XOR U17020 ( .A(n17859), .B(n17786), .Z(n17697) );
  XOR U17021 ( .A(n17860), .B(n17778), .Z(n17786) );
  XOR U17022 ( .A(n17861), .B(n17767), .Z(n17778) );
  XNOR U17023 ( .A(q[14]), .B(DB[29]), .Z(n17767) );
  IV U17024 ( .A(n17766), .Z(n17861) );
  XNOR U17025 ( .A(n17764), .B(n17862), .Z(n17766) );
  XNOR U17026 ( .A(q[13]), .B(DB[28]), .Z(n17862) );
  XNOR U17027 ( .A(q[12]), .B(DB[27]), .Z(n17764) );
  IV U17028 ( .A(n17777), .Z(n17860) );
  XOR U17029 ( .A(n17863), .B(n17864), .Z(n17777) );
  XNOR U17030 ( .A(n17773), .B(n17775), .Z(n17864) );
  XNOR U17031 ( .A(q[8]), .B(DB[23]), .Z(n17775) );
  XNOR U17032 ( .A(q[11]), .B(DB[26]), .Z(n17773) );
  IV U17033 ( .A(n17772), .Z(n17863) );
  XNOR U17034 ( .A(n17770), .B(n17865), .Z(n17772) );
  XNOR U17035 ( .A(q[10]), .B(DB[25]), .Z(n17865) );
  XNOR U17036 ( .A(q[9]), .B(DB[24]), .Z(n17770) );
  IV U17037 ( .A(n17785), .Z(n17859) );
  XOR U17038 ( .A(n17866), .B(n17867), .Z(n17785) );
  XNOR U17039 ( .A(n17802), .B(n17783), .Z(n17867) );
  XNOR U17040 ( .A(q[0]), .B(DB[15]), .Z(n17783) );
  XOR U17041 ( .A(n17868), .B(n17791), .Z(n17802) );
  XNOR U17042 ( .A(q[7]), .B(DB[22]), .Z(n17791) );
  IV U17043 ( .A(n17790), .Z(n17868) );
  XNOR U17044 ( .A(n17788), .B(n17869), .Z(n17790) );
  XNOR U17045 ( .A(q[6]), .B(DB[21]), .Z(n17869) );
  XNOR U17046 ( .A(q[5]), .B(DB[20]), .Z(n17788) );
  IV U17047 ( .A(n17801), .Z(n17866) );
  XOR U17048 ( .A(n17870), .B(n17871), .Z(n17801) );
  XNOR U17049 ( .A(n17797), .B(n17799), .Z(n17871) );
  XNOR U17050 ( .A(q[1]), .B(DB[16]), .Z(n17799) );
  XNOR U17051 ( .A(q[4]), .B(DB[19]), .Z(n17797) );
  IV U17052 ( .A(n17796), .Z(n17870) );
  XNOR U17053 ( .A(n17794), .B(n17872), .Z(n17796) );
  XNOR U17054 ( .A(q[3]), .B(DB[18]), .Z(n17872) );
  XNOR U17055 ( .A(q[2]), .B(DB[17]), .Z(n17794) );
  XOR U17056 ( .A(n17873), .B(n17675), .Z(n17603) );
  XOR U17057 ( .A(n17874), .B(n17667), .Z(n17675) );
  XOR U17058 ( .A(n17875), .B(n17656), .Z(n17667) );
  XNOR U17059 ( .A(q[14]), .B(DB[44]), .Z(n17656) );
  IV U17060 ( .A(n17655), .Z(n17875) );
  XNOR U17061 ( .A(n17653), .B(n17876), .Z(n17655) );
  XNOR U17062 ( .A(q[13]), .B(DB[43]), .Z(n17876) );
  XNOR U17063 ( .A(q[12]), .B(DB[42]), .Z(n17653) );
  IV U17064 ( .A(n17666), .Z(n17874) );
  XOR U17065 ( .A(n17877), .B(n17878), .Z(n17666) );
  XNOR U17066 ( .A(n17662), .B(n17664), .Z(n17878) );
  XNOR U17067 ( .A(q[8]), .B(DB[38]), .Z(n17664) );
  XNOR U17068 ( .A(q[11]), .B(DB[41]), .Z(n17662) );
  IV U17069 ( .A(n17661), .Z(n17877) );
  XNOR U17070 ( .A(n17659), .B(n17879), .Z(n17661) );
  XNOR U17071 ( .A(q[10]), .B(DB[40]), .Z(n17879) );
  XNOR U17072 ( .A(q[9]), .B(DB[39]), .Z(n17659) );
  IV U17073 ( .A(n17674), .Z(n17873) );
  XOR U17074 ( .A(n17880), .B(n17881), .Z(n17674) );
  XNOR U17075 ( .A(n17691), .B(n17672), .Z(n17881) );
  XNOR U17076 ( .A(q[0]), .B(DB[30]), .Z(n17672) );
  XOR U17077 ( .A(n17882), .B(n17680), .Z(n17691) );
  XNOR U17078 ( .A(q[7]), .B(DB[37]), .Z(n17680) );
  IV U17079 ( .A(n17679), .Z(n17882) );
  XNOR U17080 ( .A(n17677), .B(n17883), .Z(n17679) );
  XNOR U17081 ( .A(q[6]), .B(DB[36]), .Z(n17883) );
  XNOR U17082 ( .A(q[5]), .B(DB[35]), .Z(n17677) );
  IV U17083 ( .A(n17690), .Z(n17880) );
  XOR U17084 ( .A(n17884), .B(n17885), .Z(n17690) );
  XNOR U17085 ( .A(n17686), .B(n17688), .Z(n17885) );
  XNOR U17086 ( .A(q[1]), .B(DB[31]), .Z(n17688) );
  XNOR U17087 ( .A(q[4]), .B(DB[34]), .Z(n17686) );
  IV U17088 ( .A(n17685), .Z(n17884) );
  XNOR U17089 ( .A(n17683), .B(n17886), .Z(n17685) );
  XNOR U17090 ( .A(q[3]), .B(DB[33]), .Z(n17886) );
  XNOR U17091 ( .A(q[2]), .B(DB[32]), .Z(n17683) );
  XOR U17092 ( .A(n17887), .B(n17581), .Z(n17509) );
  XOR U17093 ( .A(n17888), .B(n17573), .Z(n17581) );
  XOR U17094 ( .A(n17889), .B(n17562), .Z(n17573) );
  XNOR U17095 ( .A(q[14]), .B(DB[59]), .Z(n17562) );
  IV U17096 ( .A(n17561), .Z(n17889) );
  XNOR U17097 ( .A(n17559), .B(n17890), .Z(n17561) );
  XNOR U17098 ( .A(q[13]), .B(DB[58]), .Z(n17890) );
  XNOR U17099 ( .A(q[12]), .B(DB[57]), .Z(n17559) );
  IV U17100 ( .A(n17572), .Z(n17888) );
  XOR U17101 ( .A(n17891), .B(n17892), .Z(n17572) );
  XNOR U17102 ( .A(n17568), .B(n17570), .Z(n17892) );
  XNOR U17103 ( .A(q[8]), .B(DB[53]), .Z(n17570) );
  XNOR U17104 ( .A(q[11]), .B(DB[56]), .Z(n17568) );
  IV U17105 ( .A(n17567), .Z(n17891) );
  XNOR U17106 ( .A(n17565), .B(n17893), .Z(n17567) );
  XNOR U17107 ( .A(q[10]), .B(DB[55]), .Z(n17893) );
  XNOR U17108 ( .A(q[9]), .B(DB[54]), .Z(n17565) );
  IV U17109 ( .A(n17580), .Z(n17887) );
  XOR U17110 ( .A(n17894), .B(n17895), .Z(n17580) );
  XNOR U17111 ( .A(n17597), .B(n17578), .Z(n17895) );
  XNOR U17112 ( .A(q[0]), .B(DB[45]), .Z(n17578) );
  XOR U17113 ( .A(n17896), .B(n17586), .Z(n17597) );
  XNOR U17114 ( .A(q[7]), .B(DB[52]), .Z(n17586) );
  IV U17115 ( .A(n17585), .Z(n17896) );
  XNOR U17116 ( .A(n17583), .B(n17897), .Z(n17585) );
  XNOR U17117 ( .A(q[6]), .B(DB[51]), .Z(n17897) );
  XNOR U17118 ( .A(q[5]), .B(DB[50]), .Z(n17583) );
  IV U17119 ( .A(n17596), .Z(n17894) );
  XOR U17120 ( .A(n17898), .B(n17899), .Z(n17596) );
  XNOR U17121 ( .A(n17592), .B(n17594), .Z(n17899) );
  XNOR U17122 ( .A(q[1]), .B(DB[46]), .Z(n17594) );
  XNOR U17123 ( .A(q[4]), .B(DB[49]), .Z(n17592) );
  IV U17124 ( .A(n17591), .Z(n17898) );
  XNOR U17125 ( .A(n17589), .B(n17900), .Z(n17591) );
  XNOR U17126 ( .A(q[3]), .B(DB[48]), .Z(n17900) );
  XNOR U17127 ( .A(q[2]), .B(DB[47]), .Z(n17589) );
  XOR U17128 ( .A(n17901), .B(n17487), .Z(n17415) );
  XOR U17129 ( .A(n17902), .B(n17479), .Z(n17487) );
  XOR U17130 ( .A(n17903), .B(n17468), .Z(n17479) );
  XNOR U17131 ( .A(q[14]), .B(DB[74]), .Z(n17468) );
  IV U17132 ( .A(n17467), .Z(n17903) );
  XNOR U17133 ( .A(n17465), .B(n17904), .Z(n17467) );
  XNOR U17134 ( .A(q[13]), .B(DB[73]), .Z(n17904) );
  XNOR U17135 ( .A(q[12]), .B(DB[72]), .Z(n17465) );
  IV U17136 ( .A(n17478), .Z(n17902) );
  XOR U17137 ( .A(n17905), .B(n17906), .Z(n17478) );
  XNOR U17138 ( .A(n17474), .B(n17476), .Z(n17906) );
  XNOR U17139 ( .A(q[8]), .B(DB[68]), .Z(n17476) );
  XNOR U17140 ( .A(q[11]), .B(DB[71]), .Z(n17474) );
  IV U17141 ( .A(n17473), .Z(n17905) );
  XNOR U17142 ( .A(n17471), .B(n17907), .Z(n17473) );
  XNOR U17143 ( .A(q[10]), .B(DB[70]), .Z(n17907) );
  XNOR U17144 ( .A(q[9]), .B(DB[69]), .Z(n17471) );
  IV U17145 ( .A(n17486), .Z(n17901) );
  XOR U17146 ( .A(n17908), .B(n17909), .Z(n17486) );
  XNOR U17147 ( .A(n17503), .B(n17484), .Z(n17909) );
  XNOR U17148 ( .A(q[0]), .B(DB[60]), .Z(n17484) );
  XOR U17149 ( .A(n17910), .B(n17492), .Z(n17503) );
  XNOR U17150 ( .A(q[7]), .B(DB[67]), .Z(n17492) );
  IV U17151 ( .A(n17491), .Z(n17910) );
  XNOR U17152 ( .A(n17489), .B(n17911), .Z(n17491) );
  XNOR U17153 ( .A(q[6]), .B(DB[66]), .Z(n17911) );
  XNOR U17154 ( .A(q[5]), .B(DB[65]), .Z(n17489) );
  IV U17155 ( .A(n17502), .Z(n17908) );
  XOR U17156 ( .A(n17912), .B(n17913), .Z(n17502) );
  XNOR U17157 ( .A(n17498), .B(n17500), .Z(n17913) );
  XNOR U17158 ( .A(q[1]), .B(DB[61]), .Z(n17500) );
  XNOR U17159 ( .A(q[4]), .B(DB[64]), .Z(n17498) );
  IV U17160 ( .A(n17497), .Z(n17912) );
  XNOR U17161 ( .A(n17495), .B(n17914), .Z(n17497) );
  XNOR U17162 ( .A(q[3]), .B(DB[63]), .Z(n17914) );
  XNOR U17163 ( .A(q[2]), .B(DB[62]), .Z(n17495) );
  XOR U17164 ( .A(n17915), .B(n17393), .Z(n17321) );
  XOR U17165 ( .A(n17916), .B(n17385), .Z(n17393) );
  XOR U17166 ( .A(n17917), .B(n17374), .Z(n17385) );
  XNOR U17167 ( .A(q[14]), .B(DB[89]), .Z(n17374) );
  IV U17168 ( .A(n17373), .Z(n17917) );
  XNOR U17169 ( .A(n17371), .B(n17918), .Z(n17373) );
  XNOR U17170 ( .A(q[13]), .B(DB[88]), .Z(n17918) );
  XNOR U17171 ( .A(q[12]), .B(DB[87]), .Z(n17371) );
  IV U17172 ( .A(n17384), .Z(n17916) );
  XOR U17173 ( .A(n17919), .B(n17920), .Z(n17384) );
  XNOR U17174 ( .A(n17380), .B(n17382), .Z(n17920) );
  XNOR U17175 ( .A(q[8]), .B(DB[83]), .Z(n17382) );
  XNOR U17176 ( .A(q[11]), .B(DB[86]), .Z(n17380) );
  IV U17177 ( .A(n17379), .Z(n17919) );
  XNOR U17178 ( .A(n17377), .B(n17921), .Z(n17379) );
  XNOR U17179 ( .A(q[10]), .B(DB[85]), .Z(n17921) );
  XNOR U17180 ( .A(q[9]), .B(DB[84]), .Z(n17377) );
  IV U17181 ( .A(n17392), .Z(n17915) );
  XOR U17182 ( .A(n17922), .B(n17923), .Z(n17392) );
  XNOR U17183 ( .A(n17409), .B(n17390), .Z(n17923) );
  XNOR U17184 ( .A(q[0]), .B(DB[75]), .Z(n17390) );
  XOR U17185 ( .A(n17924), .B(n17398), .Z(n17409) );
  XNOR U17186 ( .A(q[7]), .B(DB[82]), .Z(n17398) );
  IV U17187 ( .A(n17397), .Z(n17924) );
  XNOR U17188 ( .A(n17395), .B(n17925), .Z(n17397) );
  XNOR U17189 ( .A(q[6]), .B(DB[81]), .Z(n17925) );
  XNOR U17190 ( .A(q[5]), .B(DB[80]), .Z(n17395) );
  IV U17191 ( .A(n17408), .Z(n17922) );
  XOR U17192 ( .A(n17926), .B(n17927), .Z(n17408) );
  XNOR U17193 ( .A(n17404), .B(n17406), .Z(n17927) );
  XNOR U17194 ( .A(q[1]), .B(DB[76]), .Z(n17406) );
  XNOR U17195 ( .A(q[4]), .B(DB[79]), .Z(n17404) );
  IV U17196 ( .A(n17403), .Z(n17926) );
  XNOR U17197 ( .A(n17401), .B(n17928), .Z(n17403) );
  XNOR U17198 ( .A(q[3]), .B(DB[78]), .Z(n17928) );
  XNOR U17199 ( .A(q[2]), .B(DB[77]), .Z(n17401) );
  XOR U17200 ( .A(n17929), .B(n17299), .Z(n17227) );
  XOR U17201 ( .A(n17930), .B(n17291), .Z(n17299) );
  XOR U17202 ( .A(n17931), .B(n17280), .Z(n17291) );
  XNOR U17203 ( .A(q[14]), .B(DB[104]), .Z(n17280) );
  IV U17204 ( .A(n17279), .Z(n17931) );
  XNOR U17205 ( .A(n17277), .B(n17932), .Z(n17279) );
  XNOR U17206 ( .A(q[13]), .B(DB[103]), .Z(n17932) );
  XNOR U17207 ( .A(q[12]), .B(DB[102]), .Z(n17277) );
  IV U17208 ( .A(n17290), .Z(n17930) );
  XOR U17209 ( .A(n17933), .B(n17934), .Z(n17290) );
  XNOR U17210 ( .A(n17286), .B(n17288), .Z(n17934) );
  XNOR U17211 ( .A(q[8]), .B(DB[98]), .Z(n17288) );
  XNOR U17212 ( .A(q[11]), .B(DB[101]), .Z(n17286) );
  IV U17213 ( .A(n17285), .Z(n17933) );
  XNOR U17214 ( .A(n17283), .B(n17935), .Z(n17285) );
  XNOR U17215 ( .A(q[10]), .B(DB[100]), .Z(n17935) );
  XNOR U17216 ( .A(q[9]), .B(DB[99]), .Z(n17283) );
  IV U17217 ( .A(n17298), .Z(n17929) );
  XOR U17218 ( .A(n17936), .B(n17937), .Z(n17298) );
  XNOR U17219 ( .A(n17315), .B(n17296), .Z(n17937) );
  XNOR U17220 ( .A(q[0]), .B(DB[90]), .Z(n17296) );
  XOR U17221 ( .A(n17938), .B(n17304), .Z(n17315) );
  XNOR U17222 ( .A(q[7]), .B(DB[97]), .Z(n17304) );
  IV U17223 ( .A(n17303), .Z(n17938) );
  XNOR U17224 ( .A(n17301), .B(n17939), .Z(n17303) );
  XNOR U17225 ( .A(q[6]), .B(DB[96]), .Z(n17939) );
  XNOR U17226 ( .A(q[5]), .B(DB[95]), .Z(n17301) );
  IV U17227 ( .A(n17314), .Z(n17936) );
  XOR U17228 ( .A(n17940), .B(n17941), .Z(n17314) );
  XNOR U17229 ( .A(n17310), .B(n17312), .Z(n17941) );
  XNOR U17230 ( .A(q[1]), .B(DB[91]), .Z(n17312) );
  XNOR U17231 ( .A(q[4]), .B(DB[94]), .Z(n17310) );
  IV U17232 ( .A(n17309), .Z(n17940) );
  XNOR U17233 ( .A(n17307), .B(n17942), .Z(n17309) );
  XNOR U17234 ( .A(q[3]), .B(DB[93]), .Z(n17942) );
  XNOR U17235 ( .A(q[2]), .B(DB[92]), .Z(n17307) );
  XOR U17236 ( .A(n17943), .B(n17205), .Z(n17133) );
  XOR U17237 ( .A(n17944), .B(n17197), .Z(n17205) );
  XOR U17238 ( .A(n17945), .B(n17186), .Z(n17197) );
  XNOR U17239 ( .A(q[14]), .B(DB[119]), .Z(n17186) );
  IV U17240 ( .A(n17185), .Z(n17945) );
  XNOR U17241 ( .A(n17183), .B(n17946), .Z(n17185) );
  XNOR U17242 ( .A(q[13]), .B(DB[118]), .Z(n17946) );
  XNOR U17243 ( .A(q[12]), .B(DB[117]), .Z(n17183) );
  IV U17244 ( .A(n17196), .Z(n17944) );
  XOR U17245 ( .A(n17947), .B(n17948), .Z(n17196) );
  XNOR U17246 ( .A(n17192), .B(n17194), .Z(n17948) );
  XNOR U17247 ( .A(q[8]), .B(DB[113]), .Z(n17194) );
  XNOR U17248 ( .A(q[11]), .B(DB[116]), .Z(n17192) );
  IV U17249 ( .A(n17191), .Z(n17947) );
  XNOR U17250 ( .A(n17189), .B(n17949), .Z(n17191) );
  XNOR U17251 ( .A(q[10]), .B(DB[115]), .Z(n17949) );
  XNOR U17252 ( .A(q[9]), .B(DB[114]), .Z(n17189) );
  IV U17253 ( .A(n17204), .Z(n17943) );
  XOR U17254 ( .A(n17950), .B(n17951), .Z(n17204) );
  XNOR U17255 ( .A(n17221), .B(n17202), .Z(n17951) );
  XNOR U17256 ( .A(q[0]), .B(DB[105]), .Z(n17202) );
  XOR U17257 ( .A(n17952), .B(n17210), .Z(n17221) );
  XNOR U17258 ( .A(q[7]), .B(DB[112]), .Z(n17210) );
  IV U17259 ( .A(n17209), .Z(n17952) );
  XNOR U17260 ( .A(n17207), .B(n17953), .Z(n17209) );
  XNOR U17261 ( .A(q[6]), .B(DB[111]), .Z(n17953) );
  XNOR U17262 ( .A(q[5]), .B(DB[110]), .Z(n17207) );
  IV U17263 ( .A(n17220), .Z(n17950) );
  XOR U17264 ( .A(n17954), .B(n17955), .Z(n17220) );
  XNOR U17265 ( .A(n17216), .B(n17218), .Z(n17955) );
  XNOR U17266 ( .A(q[1]), .B(DB[106]), .Z(n17218) );
  XNOR U17267 ( .A(q[4]), .B(DB[109]), .Z(n17216) );
  IV U17268 ( .A(n17215), .Z(n17954) );
  XNOR U17269 ( .A(n17213), .B(n17956), .Z(n17215) );
  XNOR U17270 ( .A(q[3]), .B(DB[108]), .Z(n17956) );
  XNOR U17271 ( .A(q[2]), .B(DB[107]), .Z(n17213) );
  XOR U17272 ( .A(n17957), .B(n17111), .Z(n17039) );
  XOR U17273 ( .A(n17958), .B(n17103), .Z(n17111) );
  XOR U17274 ( .A(n17959), .B(n17092), .Z(n17103) );
  XNOR U17275 ( .A(q[14]), .B(DB[134]), .Z(n17092) );
  IV U17276 ( .A(n17091), .Z(n17959) );
  XNOR U17277 ( .A(n17089), .B(n17960), .Z(n17091) );
  XNOR U17278 ( .A(q[13]), .B(DB[133]), .Z(n17960) );
  XNOR U17279 ( .A(q[12]), .B(DB[132]), .Z(n17089) );
  IV U17280 ( .A(n17102), .Z(n17958) );
  XOR U17281 ( .A(n17961), .B(n17962), .Z(n17102) );
  XNOR U17282 ( .A(n17098), .B(n17100), .Z(n17962) );
  XNOR U17283 ( .A(q[8]), .B(DB[128]), .Z(n17100) );
  XNOR U17284 ( .A(q[11]), .B(DB[131]), .Z(n17098) );
  IV U17285 ( .A(n17097), .Z(n17961) );
  XNOR U17286 ( .A(n17095), .B(n17963), .Z(n17097) );
  XNOR U17287 ( .A(q[10]), .B(DB[130]), .Z(n17963) );
  XNOR U17288 ( .A(q[9]), .B(DB[129]), .Z(n17095) );
  IV U17289 ( .A(n17110), .Z(n17957) );
  XOR U17290 ( .A(n17964), .B(n17965), .Z(n17110) );
  XNOR U17291 ( .A(n17127), .B(n17108), .Z(n17965) );
  XNOR U17292 ( .A(q[0]), .B(DB[120]), .Z(n17108) );
  XOR U17293 ( .A(n17966), .B(n17116), .Z(n17127) );
  XNOR U17294 ( .A(q[7]), .B(DB[127]), .Z(n17116) );
  IV U17295 ( .A(n17115), .Z(n17966) );
  XNOR U17296 ( .A(n17113), .B(n17967), .Z(n17115) );
  XNOR U17297 ( .A(q[6]), .B(DB[126]), .Z(n17967) );
  XNOR U17298 ( .A(q[5]), .B(DB[125]), .Z(n17113) );
  IV U17299 ( .A(n17126), .Z(n17964) );
  XOR U17300 ( .A(n17968), .B(n17969), .Z(n17126) );
  XNOR U17301 ( .A(n17122), .B(n17124), .Z(n17969) );
  XNOR U17302 ( .A(q[1]), .B(DB[121]), .Z(n17124) );
  XNOR U17303 ( .A(q[4]), .B(DB[124]), .Z(n17122) );
  IV U17304 ( .A(n17121), .Z(n17968) );
  XNOR U17305 ( .A(n17119), .B(n17970), .Z(n17121) );
  XNOR U17306 ( .A(q[3]), .B(DB[123]), .Z(n17970) );
  XNOR U17307 ( .A(q[2]), .B(DB[122]), .Z(n17119) );
  XOR U17308 ( .A(n17971), .B(n17017), .Z(n16945) );
  XOR U17309 ( .A(n17972), .B(n17009), .Z(n17017) );
  XOR U17310 ( .A(n17973), .B(n16998), .Z(n17009) );
  XNOR U17311 ( .A(q[14]), .B(DB[149]), .Z(n16998) );
  IV U17312 ( .A(n16997), .Z(n17973) );
  XNOR U17313 ( .A(n16995), .B(n17974), .Z(n16997) );
  XNOR U17314 ( .A(q[13]), .B(DB[148]), .Z(n17974) );
  XNOR U17315 ( .A(q[12]), .B(DB[147]), .Z(n16995) );
  IV U17316 ( .A(n17008), .Z(n17972) );
  XOR U17317 ( .A(n17975), .B(n17976), .Z(n17008) );
  XNOR U17318 ( .A(n17004), .B(n17006), .Z(n17976) );
  XNOR U17319 ( .A(q[8]), .B(DB[143]), .Z(n17006) );
  XNOR U17320 ( .A(q[11]), .B(DB[146]), .Z(n17004) );
  IV U17321 ( .A(n17003), .Z(n17975) );
  XNOR U17322 ( .A(n17001), .B(n17977), .Z(n17003) );
  XNOR U17323 ( .A(q[10]), .B(DB[145]), .Z(n17977) );
  XNOR U17324 ( .A(q[9]), .B(DB[144]), .Z(n17001) );
  IV U17325 ( .A(n17016), .Z(n17971) );
  XOR U17326 ( .A(n17978), .B(n17979), .Z(n17016) );
  XNOR U17327 ( .A(n17033), .B(n17014), .Z(n17979) );
  XNOR U17328 ( .A(q[0]), .B(DB[135]), .Z(n17014) );
  XOR U17329 ( .A(n17980), .B(n17022), .Z(n17033) );
  XNOR U17330 ( .A(q[7]), .B(DB[142]), .Z(n17022) );
  IV U17331 ( .A(n17021), .Z(n17980) );
  XNOR U17332 ( .A(n17019), .B(n17981), .Z(n17021) );
  XNOR U17333 ( .A(q[6]), .B(DB[141]), .Z(n17981) );
  XNOR U17334 ( .A(q[5]), .B(DB[140]), .Z(n17019) );
  IV U17335 ( .A(n17032), .Z(n17978) );
  XOR U17336 ( .A(n17982), .B(n17983), .Z(n17032) );
  XNOR U17337 ( .A(n17028), .B(n17030), .Z(n17983) );
  XNOR U17338 ( .A(q[1]), .B(DB[136]), .Z(n17030) );
  XNOR U17339 ( .A(q[4]), .B(DB[139]), .Z(n17028) );
  IV U17340 ( .A(n17027), .Z(n17982) );
  XNOR U17341 ( .A(n17025), .B(n17984), .Z(n17027) );
  XNOR U17342 ( .A(q[3]), .B(DB[138]), .Z(n17984) );
  XNOR U17343 ( .A(q[2]), .B(DB[137]), .Z(n17025) );
  XOR U17344 ( .A(n17985), .B(n16923), .Z(n16851) );
  XOR U17345 ( .A(n17986), .B(n16915), .Z(n16923) );
  XOR U17346 ( .A(n17987), .B(n16904), .Z(n16915) );
  XNOR U17347 ( .A(q[14]), .B(DB[164]), .Z(n16904) );
  IV U17348 ( .A(n16903), .Z(n17987) );
  XNOR U17349 ( .A(n16901), .B(n17988), .Z(n16903) );
  XNOR U17350 ( .A(q[13]), .B(DB[163]), .Z(n17988) );
  XNOR U17351 ( .A(q[12]), .B(DB[162]), .Z(n16901) );
  IV U17352 ( .A(n16914), .Z(n17986) );
  XOR U17353 ( .A(n17989), .B(n17990), .Z(n16914) );
  XNOR U17354 ( .A(n16910), .B(n16912), .Z(n17990) );
  XNOR U17355 ( .A(q[8]), .B(DB[158]), .Z(n16912) );
  XNOR U17356 ( .A(q[11]), .B(DB[161]), .Z(n16910) );
  IV U17357 ( .A(n16909), .Z(n17989) );
  XNOR U17358 ( .A(n16907), .B(n17991), .Z(n16909) );
  XNOR U17359 ( .A(q[10]), .B(DB[160]), .Z(n17991) );
  XNOR U17360 ( .A(q[9]), .B(DB[159]), .Z(n16907) );
  IV U17361 ( .A(n16922), .Z(n17985) );
  XOR U17362 ( .A(n17992), .B(n17993), .Z(n16922) );
  XNOR U17363 ( .A(n16939), .B(n16920), .Z(n17993) );
  XNOR U17364 ( .A(q[0]), .B(DB[150]), .Z(n16920) );
  XOR U17365 ( .A(n17994), .B(n16928), .Z(n16939) );
  XNOR U17366 ( .A(q[7]), .B(DB[157]), .Z(n16928) );
  IV U17367 ( .A(n16927), .Z(n17994) );
  XNOR U17368 ( .A(n16925), .B(n17995), .Z(n16927) );
  XNOR U17369 ( .A(q[6]), .B(DB[156]), .Z(n17995) );
  XNOR U17370 ( .A(q[5]), .B(DB[155]), .Z(n16925) );
  IV U17371 ( .A(n16938), .Z(n17992) );
  XOR U17372 ( .A(n17996), .B(n17997), .Z(n16938) );
  XNOR U17373 ( .A(n16934), .B(n16936), .Z(n17997) );
  XNOR U17374 ( .A(q[1]), .B(DB[151]), .Z(n16936) );
  XNOR U17375 ( .A(q[4]), .B(DB[154]), .Z(n16934) );
  IV U17376 ( .A(n16933), .Z(n17996) );
  XNOR U17377 ( .A(n16931), .B(n17998), .Z(n16933) );
  XNOR U17378 ( .A(q[3]), .B(DB[153]), .Z(n17998) );
  XNOR U17379 ( .A(q[2]), .B(DB[152]), .Z(n16931) );
  XOR U17380 ( .A(n17999), .B(n16829), .Z(n16757) );
  XOR U17381 ( .A(n18000), .B(n16821), .Z(n16829) );
  XOR U17382 ( .A(n18001), .B(n16810), .Z(n16821) );
  XNOR U17383 ( .A(q[14]), .B(DB[179]), .Z(n16810) );
  IV U17384 ( .A(n16809), .Z(n18001) );
  XNOR U17385 ( .A(n16807), .B(n18002), .Z(n16809) );
  XNOR U17386 ( .A(q[13]), .B(DB[178]), .Z(n18002) );
  XNOR U17387 ( .A(q[12]), .B(DB[177]), .Z(n16807) );
  IV U17388 ( .A(n16820), .Z(n18000) );
  XOR U17389 ( .A(n18003), .B(n18004), .Z(n16820) );
  XNOR U17390 ( .A(n16816), .B(n16818), .Z(n18004) );
  XNOR U17391 ( .A(q[8]), .B(DB[173]), .Z(n16818) );
  XNOR U17392 ( .A(q[11]), .B(DB[176]), .Z(n16816) );
  IV U17393 ( .A(n16815), .Z(n18003) );
  XNOR U17394 ( .A(n16813), .B(n18005), .Z(n16815) );
  XNOR U17395 ( .A(q[10]), .B(DB[175]), .Z(n18005) );
  XNOR U17396 ( .A(q[9]), .B(DB[174]), .Z(n16813) );
  IV U17397 ( .A(n16828), .Z(n17999) );
  XOR U17398 ( .A(n18006), .B(n18007), .Z(n16828) );
  XNOR U17399 ( .A(n16845), .B(n16826), .Z(n18007) );
  XNOR U17400 ( .A(q[0]), .B(DB[165]), .Z(n16826) );
  XOR U17401 ( .A(n18008), .B(n16834), .Z(n16845) );
  XNOR U17402 ( .A(q[7]), .B(DB[172]), .Z(n16834) );
  IV U17403 ( .A(n16833), .Z(n18008) );
  XNOR U17404 ( .A(n16831), .B(n18009), .Z(n16833) );
  XNOR U17405 ( .A(q[6]), .B(DB[171]), .Z(n18009) );
  XNOR U17406 ( .A(q[5]), .B(DB[170]), .Z(n16831) );
  IV U17407 ( .A(n16844), .Z(n18006) );
  XOR U17408 ( .A(n18010), .B(n18011), .Z(n16844) );
  XNOR U17409 ( .A(n16840), .B(n16842), .Z(n18011) );
  XNOR U17410 ( .A(q[1]), .B(DB[166]), .Z(n16842) );
  XNOR U17411 ( .A(q[4]), .B(DB[169]), .Z(n16840) );
  IV U17412 ( .A(n16839), .Z(n18010) );
  XNOR U17413 ( .A(n16837), .B(n18012), .Z(n16839) );
  XNOR U17414 ( .A(q[3]), .B(DB[168]), .Z(n18012) );
  XNOR U17415 ( .A(q[2]), .B(DB[167]), .Z(n16837) );
  XOR U17416 ( .A(n18013), .B(n16735), .Z(n16663) );
  XOR U17417 ( .A(n18014), .B(n16727), .Z(n16735) );
  XOR U17418 ( .A(n18015), .B(n16716), .Z(n16727) );
  XNOR U17419 ( .A(q[14]), .B(DB[194]), .Z(n16716) );
  IV U17420 ( .A(n16715), .Z(n18015) );
  XNOR U17421 ( .A(n16713), .B(n18016), .Z(n16715) );
  XNOR U17422 ( .A(q[13]), .B(DB[193]), .Z(n18016) );
  XNOR U17423 ( .A(q[12]), .B(DB[192]), .Z(n16713) );
  IV U17424 ( .A(n16726), .Z(n18014) );
  XOR U17425 ( .A(n18017), .B(n18018), .Z(n16726) );
  XNOR U17426 ( .A(n16722), .B(n16724), .Z(n18018) );
  XNOR U17427 ( .A(q[8]), .B(DB[188]), .Z(n16724) );
  XNOR U17428 ( .A(q[11]), .B(DB[191]), .Z(n16722) );
  IV U17429 ( .A(n16721), .Z(n18017) );
  XNOR U17430 ( .A(n16719), .B(n18019), .Z(n16721) );
  XNOR U17431 ( .A(q[10]), .B(DB[190]), .Z(n18019) );
  XNOR U17432 ( .A(q[9]), .B(DB[189]), .Z(n16719) );
  IV U17433 ( .A(n16734), .Z(n18013) );
  XOR U17434 ( .A(n18020), .B(n18021), .Z(n16734) );
  XNOR U17435 ( .A(n16751), .B(n16732), .Z(n18021) );
  XNOR U17436 ( .A(q[0]), .B(DB[180]), .Z(n16732) );
  XOR U17437 ( .A(n18022), .B(n16740), .Z(n16751) );
  XNOR U17438 ( .A(q[7]), .B(DB[187]), .Z(n16740) );
  IV U17439 ( .A(n16739), .Z(n18022) );
  XNOR U17440 ( .A(n16737), .B(n18023), .Z(n16739) );
  XNOR U17441 ( .A(q[6]), .B(DB[186]), .Z(n18023) );
  XNOR U17442 ( .A(q[5]), .B(DB[185]), .Z(n16737) );
  IV U17443 ( .A(n16750), .Z(n18020) );
  XOR U17444 ( .A(n18024), .B(n18025), .Z(n16750) );
  XNOR U17445 ( .A(n16746), .B(n16748), .Z(n18025) );
  XNOR U17446 ( .A(q[1]), .B(DB[181]), .Z(n16748) );
  XNOR U17447 ( .A(q[4]), .B(DB[184]), .Z(n16746) );
  IV U17448 ( .A(n16745), .Z(n18024) );
  XNOR U17449 ( .A(n16743), .B(n18026), .Z(n16745) );
  XNOR U17450 ( .A(q[3]), .B(DB[183]), .Z(n18026) );
  XNOR U17451 ( .A(q[2]), .B(DB[182]), .Z(n16743) );
  XOR U17452 ( .A(n18027), .B(n16641), .Z(n16569) );
  XOR U17453 ( .A(n18028), .B(n16633), .Z(n16641) );
  XOR U17454 ( .A(n18029), .B(n16622), .Z(n16633) );
  XNOR U17455 ( .A(q[14]), .B(DB[209]), .Z(n16622) );
  IV U17456 ( .A(n16621), .Z(n18029) );
  XNOR U17457 ( .A(n16619), .B(n18030), .Z(n16621) );
  XNOR U17458 ( .A(q[13]), .B(DB[208]), .Z(n18030) );
  XNOR U17459 ( .A(q[12]), .B(DB[207]), .Z(n16619) );
  IV U17460 ( .A(n16632), .Z(n18028) );
  XOR U17461 ( .A(n18031), .B(n18032), .Z(n16632) );
  XNOR U17462 ( .A(n16628), .B(n16630), .Z(n18032) );
  XNOR U17463 ( .A(q[8]), .B(DB[203]), .Z(n16630) );
  XNOR U17464 ( .A(q[11]), .B(DB[206]), .Z(n16628) );
  IV U17465 ( .A(n16627), .Z(n18031) );
  XNOR U17466 ( .A(n16625), .B(n18033), .Z(n16627) );
  XNOR U17467 ( .A(q[10]), .B(DB[205]), .Z(n18033) );
  XNOR U17468 ( .A(q[9]), .B(DB[204]), .Z(n16625) );
  IV U17469 ( .A(n16640), .Z(n18027) );
  XOR U17470 ( .A(n18034), .B(n18035), .Z(n16640) );
  XNOR U17471 ( .A(n16657), .B(n16638), .Z(n18035) );
  XNOR U17472 ( .A(q[0]), .B(DB[195]), .Z(n16638) );
  XOR U17473 ( .A(n18036), .B(n16646), .Z(n16657) );
  XNOR U17474 ( .A(q[7]), .B(DB[202]), .Z(n16646) );
  IV U17475 ( .A(n16645), .Z(n18036) );
  XNOR U17476 ( .A(n16643), .B(n18037), .Z(n16645) );
  XNOR U17477 ( .A(q[6]), .B(DB[201]), .Z(n18037) );
  XNOR U17478 ( .A(q[5]), .B(DB[200]), .Z(n16643) );
  IV U17479 ( .A(n16656), .Z(n18034) );
  XOR U17480 ( .A(n18038), .B(n18039), .Z(n16656) );
  XNOR U17481 ( .A(n16652), .B(n16654), .Z(n18039) );
  XNOR U17482 ( .A(q[1]), .B(DB[196]), .Z(n16654) );
  XNOR U17483 ( .A(q[4]), .B(DB[199]), .Z(n16652) );
  IV U17484 ( .A(n16651), .Z(n18038) );
  XNOR U17485 ( .A(n16649), .B(n18040), .Z(n16651) );
  XNOR U17486 ( .A(q[3]), .B(DB[198]), .Z(n18040) );
  XNOR U17487 ( .A(q[2]), .B(DB[197]), .Z(n16649) );
  XOR U17488 ( .A(n18041), .B(n16547), .Z(n16475) );
  XOR U17489 ( .A(n18042), .B(n16539), .Z(n16547) );
  XOR U17490 ( .A(n18043), .B(n16528), .Z(n16539) );
  XNOR U17491 ( .A(q[14]), .B(DB[224]), .Z(n16528) );
  IV U17492 ( .A(n16527), .Z(n18043) );
  XNOR U17493 ( .A(n16525), .B(n18044), .Z(n16527) );
  XNOR U17494 ( .A(q[13]), .B(DB[223]), .Z(n18044) );
  XNOR U17495 ( .A(q[12]), .B(DB[222]), .Z(n16525) );
  IV U17496 ( .A(n16538), .Z(n18042) );
  XOR U17497 ( .A(n18045), .B(n18046), .Z(n16538) );
  XNOR U17498 ( .A(n16534), .B(n16536), .Z(n18046) );
  XNOR U17499 ( .A(q[8]), .B(DB[218]), .Z(n16536) );
  XNOR U17500 ( .A(q[11]), .B(DB[221]), .Z(n16534) );
  IV U17501 ( .A(n16533), .Z(n18045) );
  XNOR U17502 ( .A(n16531), .B(n18047), .Z(n16533) );
  XNOR U17503 ( .A(q[10]), .B(DB[220]), .Z(n18047) );
  XNOR U17504 ( .A(q[9]), .B(DB[219]), .Z(n16531) );
  IV U17505 ( .A(n16546), .Z(n18041) );
  XOR U17506 ( .A(n18048), .B(n18049), .Z(n16546) );
  XNOR U17507 ( .A(n16563), .B(n16544), .Z(n18049) );
  XNOR U17508 ( .A(q[0]), .B(DB[210]), .Z(n16544) );
  XOR U17509 ( .A(n18050), .B(n16552), .Z(n16563) );
  XNOR U17510 ( .A(q[7]), .B(DB[217]), .Z(n16552) );
  IV U17511 ( .A(n16551), .Z(n18050) );
  XNOR U17512 ( .A(n16549), .B(n18051), .Z(n16551) );
  XNOR U17513 ( .A(q[6]), .B(DB[216]), .Z(n18051) );
  XNOR U17514 ( .A(q[5]), .B(DB[215]), .Z(n16549) );
  IV U17515 ( .A(n16562), .Z(n18048) );
  XOR U17516 ( .A(n18052), .B(n18053), .Z(n16562) );
  XNOR U17517 ( .A(n16558), .B(n16560), .Z(n18053) );
  XNOR U17518 ( .A(q[1]), .B(DB[211]), .Z(n16560) );
  XNOR U17519 ( .A(q[4]), .B(DB[214]), .Z(n16558) );
  IV U17520 ( .A(n16557), .Z(n18052) );
  XNOR U17521 ( .A(n16555), .B(n18054), .Z(n16557) );
  XNOR U17522 ( .A(q[3]), .B(DB[213]), .Z(n18054) );
  XNOR U17523 ( .A(q[2]), .B(DB[212]), .Z(n16555) );
  XOR U17524 ( .A(n18055), .B(n16453), .Z(n16381) );
  XOR U17525 ( .A(n18056), .B(n16445), .Z(n16453) );
  XOR U17526 ( .A(n18057), .B(n16434), .Z(n16445) );
  XNOR U17527 ( .A(q[14]), .B(DB[239]), .Z(n16434) );
  IV U17528 ( .A(n16433), .Z(n18057) );
  XNOR U17529 ( .A(n16431), .B(n18058), .Z(n16433) );
  XNOR U17530 ( .A(q[13]), .B(DB[238]), .Z(n18058) );
  XNOR U17531 ( .A(q[12]), .B(DB[237]), .Z(n16431) );
  IV U17532 ( .A(n16444), .Z(n18056) );
  XOR U17533 ( .A(n18059), .B(n18060), .Z(n16444) );
  XNOR U17534 ( .A(n16440), .B(n16442), .Z(n18060) );
  XNOR U17535 ( .A(q[8]), .B(DB[233]), .Z(n16442) );
  XNOR U17536 ( .A(q[11]), .B(DB[236]), .Z(n16440) );
  IV U17537 ( .A(n16439), .Z(n18059) );
  XNOR U17538 ( .A(n16437), .B(n18061), .Z(n16439) );
  XNOR U17539 ( .A(q[10]), .B(DB[235]), .Z(n18061) );
  XNOR U17540 ( .A(q[9]), .B(DB[234]), .Z(n16437) );
  IV U17541 ( .A(n16452), .Z(n18055) );
  XOR U17542 ( .A(n18062), .B(n18063), .Z(n16452) );
  XNOR U17543 ( .A(n16469), .B(n16450), .Z(n18063) );
  XNOR U17544 ( .A(q[0]), .B(DB[225]), .Z(n16450) );
  XOR U17545 ( .A(n18064), .B(n16458), .Z(n16469) );
  XNOR U17546 ( .A(q[7]), .B(DB[232]), .Z(n16458) );
  IV U17547 ( .A(n16457), .Z(n18064) );
  XNOR U17548 ( .A(n16455), .B(n18065), .Z(n16457) );
  XNOR U17549 ( .A(q[6]), .B(DB[231]), .Z(n18065) );
  XNOR U17550 ( .A(q[5]), .B(DB[230]), .Z(n16455) );
  IV U17551 ( .A(n16468), .Z(n18062) );
  XOR U17552 ( .A(n18066), .B(n18067), .Z(n16468) );
  XNOR U17553 ( .A(n16464), .B(n16466), .Z(n18067) );
  XNOR U17554 ( .A(q[1]), .B(DB[226]), .Z(n16466) );
  XNOR U17555 ( .A(q[4]), .B(DB[229]), .Z(n16464) );
  IV U17556 ( .A(n16463), .Z(n18066) );
  XNOR U17557 ( .A(n16461), .B(n18068), .Z(n16463) );
  XNOR U17558 ( .A(q[3]), .B(DB[228]), .Z(n18068) );
  XNOR U17559 ( .A(q[2]), .B(DB[227]), .Z(n16461) );
  XOR U17560 ( .A(n18069), .B(n16359), .Z(n16287) );
  XOR U17561 ( .A(n18070), .B(n16351), .Z(n16359) );
  XOR U17562 ( .A(n18071), .B(n16340), .Z(n16351) );
  XNOR U17563 ( .A(q[14]), .B(DB[254]), .Z(n16340) );
  IV U17564 ( .A(n16339), .Z(n18071) );
  XNOR U17565 ( .A(n16337), .B(n18072), .Z(n16339) );
  XNOR U17566 ( .A(q[13]), .B(DB[253]), .Z(n18072) );
  XNOR U17567 ( .A(q[12]), .B(DB[252]), .Z(n16337) );
  IV U17568 ( .A(n16350), .Z(n18070) );
  XOR U17569 ( .A(n18073), .B(n18074), .Z(n16350) );
  XNOR U17570 ( .A(n16346), .B(n16348), .Z(n18074) );
  XNOR U17571 ( .A(q[8]), .B(DB[248]), .Z(n16348) );
  XNOR U17572 ( .A(q[11]), .B(DB[251]), .Z(n16346) );
  IV U17573 ( .A(n16345), .Z(n18073) );
  XNOR U17574 ( .A(n16343), .B(n18075), .Z(n16345) );
  XNOR U17575 ( .A(q[10]), .B(DB[250]), .Z(n18075) );
  XNOR U17576 ( .A(q[9]), .B(DB[249]), .Z(n16343) );
  IV U17577 ( .A(n16358), .Z(n18069) );
  XOR U17578 ( .A(n18076), .B(n18077), .Z(n16358) );
  XNOR U17579 ( .A(n16375), .B(n16356), .Z(n18077) );
  XNOR U17580 ( .A(q[0]), .B(DB[240]), .Z(n16356) );
  XOR U17581 ( .A(n18078), .B(n16364), .Z(n16375) );
  XNOR U17582 ( .A(q[7]), .B(DB[247]), .Z(n16364) );
  IV U17583 ( .A(n16363), .Z(n18078) );
  XNOR U17584 ( .A(n16361), .B(n18079), .Z(n16363) );
  XNOR U17585 ( .A(q[6]), .B(DB[246]), .Z(n18079) );
  XNOR U17586 ( .A(q[5]), .B(DB[245]), .Z(n16361) );
  IV U17587 ( .A(n16374), .Z(n18076) );
  XOR U17588 ( .A(n18080), .B(n18081), .Z(n16374) );
  XNOR U17589 ( .A(n16370), .B(n16372), .Z(n18081) );
  XNOR U17590 ( .A(q[1]), .B(DB[241]), .Z(n16372) );
  XNOR U17591 ( .A(q[4]), .B(DB[244]), .Z(n16370) );
  IV U17592 ( .A(n16369), .Z(n18080) );
  XNOR U17593 ( .A(n16367), .B(n18082), .Z(n16369) );
  XNOR U17594 ( .A(q[3]), .B(DB[243]), .Z(n18082) );
  XNOR U17595 ( .A(q[2]), .B(DB[242]), .Z(n16367) );
  XOR U17596 ( .A(n18083), .B(n16265), .Z(n16193) );
  XOR U17597 ( .A(n18084), .B(n16257), .Z(n16265) );
  XOR U17598 ( .A(n18085), .B(n16246), .Z(n16257) );
  XNOR U17599 ( .A(q[14]), .B(DB[269]), .Z(n16246) );
  IV U17600 ( .A(n16245), .Z(n18085) );
  XNOR U17601 ( .A(n16243), .B(n18086), .Z(n16245) );
  XNOR U17602 ( .A(q[13]), .B(DB[268]), .Z(n18086) );
  XNOR U17603 ( .A(q[12]), .B(DB[267]), .Z(n16243) );
  IV U17604 ( .A(n16256), .Z(n18084) );
  XOR U17605 ( .A(n18087), .B(n18088), .Z(n16256) );
  XNOR U17606 ( .A(n16252), .B(n16254), .Z(n18088) );
  XNOR U17607 ( .A(q[8]), .B(DB[263]), .Z(n16254) );
  XNOR U17608 ( .A(q[11]), .B(DB[266]), .Z(n16252) );
  IV U17609 ( .A(n16251), .Z(n18087) );
  XNOR U17610 ( .A(n16249), .B(n18089), .Z(n16251) );
  XNOR U17611 ( .A(q[10]), .B(DB[265]), .Z(n18089) );
  XNOR U17612 ( .A(q[9]), .B(DB[264]), .Z(n16249) );
  IV U17613 ( .A(n16264), .Z(n18083) );
  XOR U17614 ( .A(n18090), .B(n18091), .Z(n16264) );
  XNOR U17615 ( .A(n16281), .B(n16262), .Z(n18091) );
  XNOR U17616 ( .A(q[0]), .B(DB[255]), .Z(n16262) );
  XOR U17617 ( .A(n18092), .B(n16270), .Z(n16281) );
  XNOR U17618 ( .A(q[7]), .B(DB[262]), .Z(n16270) );
  IV U17619 ( .A(n16269), .Z(n18092) );
  XNOR U17620 ( .A(n16267), .B(n18093), .Z(n16269) );
  XNOR U17621 ( .A(q[6]), .B(DB[261]), .Z(n18093) );
  XNOR U17622 ( .A(q[5]), .B(DB[260]), .Z(n16267) );
  IV U17623 ( .A(n16280), .Z(n18090) );
  XOR U17624 ( .A(n18094), .B(n18095), .Z(n16280) );
  XNOR U17625 ( .A(n16276), .B(n16278), .Z(n18095) );
  XNOR U17626 ( .A(q[1]), .B(DB[256]), .Z(n16278) );
  XNOR U17627 ( .A(q[4]), .B(DB[259]), .Z(n16276) );
  IV U17628 ( .A(n16275), .Z(n18094) );
  XNOR U17629 ( .A(n16273), .B(n18096), .Z(n16275) );
  XNOR U17630 ( .A(q[3]), .B(DB[258]), .Z(n18096) );
  XNOR U17631 ( .A(q[2]), .B(DB[257]), .Z(n16273) );
  XOR U17632 ( .A(n18097), .B(n16171), .Z(n16099) );
  XOR U17633 ( .A(n18098), .B(n16163), .Z(n16171) );
  XOR U17634 ( .A(n18099), .B(n16152), .Z(n16163) );
  XNOR U17635 ( .A(q[14]), .B(DB[284]), .Z(n16152) );
  IV U17636 ( .A(n16151), .Z(n18099) );
  XNOR U17637 ( .A(n16149), .B(n18100), .Z(n16151) );
  XNOR U17638 ( .A(q[13]), .B(DB[283]), .Z(n18100) );
  XNOR U17639 ( .A(q[12]), .B(DB[282]), .Z(n16149) );
  IV U17640 ( .A(n16162), .Z(n18098) );
  XOR U17641 ( .A(n18101), .B(n18102), .Z(n16162) );
  XNOR U17642 ( .A(n16158), .B(n16160), .Z(n18102) );
  XNOR U17643 ( .A(q[8]), .B(DB[278]), .Z(n16160) );
  XNOR U17644 ( .A(q[11]), .B(DB[281]), .Z(n16158) );
  IV U17645 ( .A(n16157), .Z(n18101) );
  XNOR U17646 ( .A(n16155), .B(n18103), .Z(n16157) );
  XNOR U17647 ( .A(q[10]), .B(DB[280]), .Z(n18103) );
  XNOR U17648 ( .A(q[9]), .B(DB[279]), .Z(n16155) );
  IV U17649 ( .A(n16170), .Z(n18097) );
  XOR U17650 ( .A(n18104), .B(n18105), .Z(n16170) );
  XNOR U17651 ( .A(n16187), .B(n16168), .Z(n18105) );
  XNOR U17652 ( .A(q[0]), .B(DB[270]), .Z(n16168) );
  XOR U17653 ( .A(n18106), .B(n16176), .Z(n16187) );
  XNOR U17654 ( .A(q[7]), .B(DB[277]), .Z(n16176) );
  IV U17655 ( .A(n16175), .Z(n18106) );
  XNOR U17656 ( .A(n16173), .B(n18107), .Z(n16175) );
  XNOR U17657 ( .A(q[6]), .B(DB[276]), .Z(n18107) );
  XNOR U17658 ( .A(q[5]), .B(DB[275]), .Z(n16173) );
  IV U17659 ( .A(n16186), .Z(n18104) );
  XOR U17660 ( .A(n18108), .B(n18109), .Z(n16186) );
  XNOR U17661 ( .A(n16182), .B(n16184), .Z(n18109) );
  XNOR U17662 ( .A(q[1]), .B(DB[271]), .Z(n16184) );
  XNOR U17663 ( .A(q[4]), .B(DB[274]), .Z(n16182) );
  IV U17664 ( .A(n16181), .Z(n18108) );
  XNOR U17665 ( .A(n16179), .B(n18110), .Z(n16181) );
  XNOR U17666 ( .A(q[3]), .B(DB[273]), .Z(n18110) );
  XNOR U17667 ( .A(q[2]), .B(DB[272]), .Z(n16179) );
  XOR U17668 ( .A(n18111), .B(n16077), .Z(n16005) );
  XOR U17669 ( .A(n18112), .B(n16069), .Z(n16077) );
  XOR U17670 ( .A(n18113), .B(n16058), .Z(n16069) );
  XNOR U17671 ( .A(q[14]), .B(DB[299]), .Z(n16058) );
  IV U17672 ( .A(n16057), .Z(n18113) );
  XNOR U17673 ( .A(n16055), .B(n18114), .Z(n16057) );
  XNOR U17674 ( .A(q[13]), .B(DB[298]), .Z(n18114) );
  XNOR U17675 ( .A(q[12]), .B(DB[297]), .Z(n16055) );
  IV U17676 ( .A(n16068), .Z(n18112) );
  XOR U17677 ( .A(n18115), .B(n18116), .Z(n16068) );
  XNOR U17678 ( .A(n16064), .B(n16066), .Z(n18116) );
  XNOR U17679 ( .A(q[8]), .B(DB[293]), .Z(n16066) );
  XNOR U17680 ( .A(q[11]), .B(DB[296]), .Z(n16064) );
  IV U17681 ( .A(n16063), .Z(n18115) );
  XNOR U17682 ( .A(n16061), .B(n18117), .Z(n16063) );
  XNOR U17683 ( .A(q[10]), .B(DB[295]), .Z(n18117) );
  XNOR U17684 ( .A(q[9]), .B(DB[294]), .Z(n16061) );
  IV U17685 ( .A(n16076), .Z(n18111) );
  XOR U17686 ( .A(n18118), .B(n18119), .Z(n16076) );
  XNOR U17687 ( .A(n16093), .B(n16074), .Z(n18119) );
  XNOR U17688 ( .A(q[0]), .B(DB[285]), .Z(n16074) );
  XOR U17689 ( .A(n18120), .B(n16082), .Z(n16093) );
  XNOR U17690 ( .A(q[7]), .B(DB[292]), .Z(n16082) );
  IV U17691 ( .A(n16081), .Z(n18120) );
  XNOR U17692 ( .A(n16079), .B(n18121), .Z(n16081) );
  XNOR U17693 ( .A(q[6]), .B(DB[291]), .Z(n18121) );
  XNOR U17694 ( .A(q[5]), .B(DB[290]), .Z(n16079) );
  IV U17695 ( .A(n16092), .Z(n18118) );
  XOR U17696 ( .A(n18122), .B(n18123), .Z(n16092) );
  XNOR U17697 ( .A(n16088), .B(n16090), .Z(n18123) );
  XNOR U17698 ( .A(q[1]), .B(DB[286]), .Z(n16090) );
  XNOR U17699 ( .A(q[4]), .B(DB[289]), .Z(n16088) );
  IV U17700 ( .A(n16087), .Z(n18122) );
  XNOR U17701 ( .A(n16085), .B(n18124), .Z(n16087) );
  XNOR U17702 ( .A(q[3]), .B(DB[288]), .Z(n18124) );
  XNOR U17703 ( .A(q[2]), .B(DB[287]), .Z(n16085) );
  XOR U17704 ( .A(n18125), .B(n15983), .Z(n15911) );
  XOR U17705 ( .A(n18126), .B(n15975), .Z(n15983) );
  XOR U17706 ( .A(n18127), .B(n15964), .Z(n15975) );
  XNOR U17707 ( .A(q[14]), .B(DB[314]), .Z(n15964) );
  IV U17708 ( .A(n15963), .Z(n18127) );
  XNOR U17709 ( .A(n15961), .B(n18128), .Z(n15963) );
  XNOR U17710 ( .A(q[13]), .B(DB[313]), .Z(n18128) );
  XNOR U17711 ( .A(q[12]), .B(DB[312]), .Z(n15961) );
  IV U17712 ( .A(n15974), .Z(n18126) );
  XOR U17713 ( .A(n18129), .B(n18130), .Z(n15974) );
  XNOR U17714 ( .A(n15970), .B(n15972), .Z(n18130) );
  XNOR U17715 ( .A(q[8]), .B(DB[308]), .Z(n15972) );
  XNOR U17716 ( .A(q[11]), .B(DB[311]), .Z(n15970) );
  IV U17717 ( .A(n15969), .Z(n18129) );
  XNOR U17718 ( .A(n15967), .B(n18131), .Z(n15969) );
  XNOR U17719 ( .A(q[10]), .B(DB[310]), .Z(n18131) );
  XNOR U17720 ( .A(q[9]), .B(DB[309]), .Z(n15967) );
  IV U17721 ( .A(n15982), .Z(n18125) );
  XOR U17722 ( .A(n18132), .B(n18133), .Z(n15982) );
  XNOR U17723 ( .A(n15999), .B(n15980), .Z(n18133) );
  XNOR U17724 ( .A(q[0]), .B(DB[300]), .Z(n15980) );
  XOR U17725 ( .A(n18134), .B(n15988), .Z(n15999) );
  XNOR U17726 ( .A(q[7]), .B(DB[307]), .Z(n15988) );
  IV U17727 ( .A(n15987), .Z(n18134) );
  XNOR U17728 ( .A(n15985), .B(n18135), .Z(n15987) );
  XNOR U17729 ( .A(q[6]), .B(DB[306]), .Z(n18135) );
  XNOR U17730 ( .A(q[5]), .B(DB[305]), .Z(n15985) );
  IV U17731 ( .A(n15998), .Z(n18132) );
  XOR U17732 ( .A(n18136), .B(n18137), .Z(n15998) );
  XNOR U17733 ( .A(n15994), .B(n15996), .Z(n18137) );
  XNOR U17734 ( .A(q[1]), .B(DB[301]), .Z(n15996) );
  XNOR U17735 ( .A(q[4]), .B(DB[304]), .Z(n15994) );
  IV U17736 ( .A(n15993), .Z(n18136) );
  XNOR U17737 ( .A(n15991), .B(n18138), .Z(n15993) );
  XNOR U17738 ( .A(q[3]), .B(DB[303]), .Z(n18138) );
  XNOR U17739 ( .A(q[2]), .B(DB[302]), .Z(n15991) );
  XOR U17740 ( .A(n18139), .B(n15889), .Z(n15817) );
  XOR U17741 ( .A(n18140), .B(n15881), .Z(n15889) );
  XOR U17742 ( .A(n18141), .B(n15870), .Z(n15881) );
  XNOR U17743 ( .A(q[14]), .B(DB[329]), .Z(n15870) );
  IV U17744 ( .A(n15869), .Z(n18141) );
  XNOR U17745 ( .A(n15867), .B(n18142), .Z(n15869) );
  XNOR U17746 ( .A(q[13]), .B(DB[328]), .Z(n18142) );
  XNOR U17747 ( .A(q[12]), .B(DB[327]), .Z(n15867) );
  IV U17748 ( .A(n15880), .Z(n18140) );
  XOR U17749 ( .A(n18143), .B(n18144), .Z(n15880) );
  XNOR U17750 ( .A(n15876), .B(n15878), .Z(n18144) );
  XNOR U17751 ( .A(q[8]), .B(DB[323]), .Z(n15878) );
  XNOR U17752 ( .A(q[11]), .B(DB[326]), .Z(n15876) );
  IV U17753 ( .A(n15875), .Z(n18143) );
  XNOR U17754 ( .A(n15873), .B(n18145), .Z(n15875) );
  XNOR U17755 ( .A(q[10]), .B(DB[325]), .Z(n18145) );
  XNOR U17756 ( .A(q[9]), .B(DB[324]), .Z(n15873) );
  IV U17757 ( .A(n15888), .Z(n18139) );
  XOR U17758 ( .A(n18146), .B(n18147), .Z(n15888) );
  XNOR U17759 ( .A(n15905), .B(n15886), .Z(n18147) );
  XNOR U17760 ( .A(q[0]), .B(DB[315]), .Z(n15886) );
  XOR U17761 ( .A(n18148), .B(n15894), .Z(n15905) );
  XNOR U17762 ( .A(q[7]), .B(DB[322]), .Z(n15894) );
  IV U17763 ( .A(n15893), .Z(n18148) );
  XNOR U17764 ( .A(n15891), .B(n18149), .Z(n15893) );
  XNOR U17765 ( .A(q[6]), .B(DB[321]), .Z(n18149) );
  XNOR U17766 ( .A(q[5]), .B(DB[320]), .Z(n15891) );
  IV U17767 ( .A(n15904), .Z(n18146) );
  XOR U17768 ( .A(n18150), .B(n18151), .Z(n15904) );
  XNOR U17769 ( .A(n15900), .B(n15902), .Z(n18151) );
  XNOR U17770 ( .A(q[1]), .B(DB[316]), .Z(n15902) );
  XNOR U17771 ( .A(q[4]), .B(DB[319]), .Z(n15900) );
  IV U17772 ( .A(n15899), .Z(n18150) );
  XNOR U17773 ( .A(n15897), .B(n18152), .Z(n15899) );
  XNOR U17774 ( .A(q[3]), .B(DB[318]), .Z(n18152) );
  XNOR U17775 ( .A(q[2]), .B(DB[317]), .Z(n15897) );
  XOR U17776 ( .A(n18153), .B(n15795), .Z(n15723) );
  XOR U17777 ( .A(n18154), .B(n15787), .Z(n15795) );
  XOR U17778 ( .A(n18155), .B(n15776), .Z(n15787) );
  XNOR U17779 ( .A(q[14]), .B(DB[344]), .Z(n15776) );
  IV U17780 ( .A(n15775), .Z(n18155) );
  XNOR U17781 ( .A(n15773), .B(n18156), .Z(n15775) );
  XNOR U17782 ( .A(q[13]), .B(DB[343]), .Z(n18156) );
  XNOR U17783 ( .A(q[12]), .B(DB[342]), .Z(n15773) );
  IV U17784 ( .A(n15786), .Z(n18154) );
  XOR U17785 ( .A(n18157), .B(n18158), .Z(n15786) );
  XNOR U17786 ( .A(n15782), .B(n15784), .Z(n18158) );
  XNOR U17787 ( .A(q[8]), .B(DB[338]), .Z(n15784) );
  XNOR U17788 ( .A(q[11]), .B(DB[341]), .Z(n15782) );
  IV U17789 ( .A(n15781), .Z(n18157) );
  XNOR U17790 ( .A(n15779), .B(n18159), .Z(n15781) );
  XNOR U17791 ( .A(q[10]), .B(DB[340]), .Z(n18159) );
  XNOR U17792 ( .A(q[9]), .B(DB[339]), .Z(n15779) );
  IV U17793 ( .A(n15794), .Z(n18153) );
  XOR U17794 ( .A(n18160), .B(n18161), .Z(n15794) );
  XNOR U17795 ( .A(n15811), .B(n15792), .Z(n18161) );
  XNOR U17796 ( .A(q[0]), .B(DB[330]), .Z(n15792) );
  XOR U17797 ( .A(n18162), .B(n15800), .Z(n15811) );
  XNOR U17798 ( .A(q[7]), .B(DB[337]), .Z(n15800) );
  IV U17799 ( .A(n15799), .Z(n18162) );
  XNOR U17800 ( .A(n15797), .B(n18163), .Z(n15799) );
  XNOR U17801 ( .A(q[6]), .B(DB[336]), .Z(n18163) );
  XNOR U17802 ( .A(q[5]), .B(DB[335]), .Z(n15797) );
  IV U17803 ( .A(n15810), .Z(n18160) );
  XOR U17804 ( .A(n18164), .B(n18165), .Z(n15810) );
  XNOR U17805 ( .A(n15806), .B(n15808), .Z(n18165) );
  XNOR U17806 ( .A(q[1]), .B(DB[331]), .Z(n15808) );
  XNOR U17807 ( .A(q[4]), .B(DB[334]), .Z(n15806) );
  IV U17808 ( .A(n15805), .Z(n18164) );
  XNOR U17809 ( .A(n15803), .B(n18166), .Z(n15805) );
  XNOR U17810 ( .A(q[3]), .B(DB[333]), .Z(n18166) );
  XNOR U17811 ( .A(q[2]), .B(DB[332]), .Z(n15803) );
  XOR U17812 ( .A(n18167), .B(n15701), .Z(n15629) );
  XOR U17813 ( .A(n18168), .B(n15693), .Z(n15701) );
  XOR U17814 ( .A(n18169), .B(n15682), .Z(n15693) );
  XNOR U17815 ( .A(q[14]), .B(DB[359]), .Z(n15682) );
  IV U17816 ( .A(n15681), .Z(n18169) );
  XNOR U17817 ( .A(n15679), .B(n18170), .Z(n15681) );
  XNOR U17818 ( .A(q[13]), .B(DB[358]), .Z(n18170) );
  XNOR U17819 ( .A(q[12]), .B(DB[357]), .Z(n15679) );
  IV U17820 ( .A(n15692), .Z(n18168) );
  XOR U17821 ( .A(n18171), .B(n18172), .Z(n15692) );
  XNOR U17822 ( .A(n15688), .B(n15690), .Z(n18172) );
  XNOR U17823 ( .A(q[8]), .B(DB[353]), .Z(n15690) );
  XNOR U17824 ( .A(q[11]), .B(DB[356]), .Z(n15688) );
  IV U17825 ( .A(n15687), .Z(n18171) );
  XNOR U17826 ( .A(n15685), .B(n18173), .Z(n15687) );
  XNOR U17827 ( .A(q[10]), .B(DB[355]), .Z(n18173) );
  XNOR U17828 ( .A(q[9]), .B(DB[354]), .Z(n15685) );
  IV U17829 ( .A(n15700), .Z(n18167) );
  XOR U17830 ( .A(n18174), .B(n18175), .Z(n15700) );
  XNOR U17831 ( .A(n15717), .B(n15698), .Z(n18175) );
  XNOR U17832 ( .A(q[0]), .B(DB[345]), .Z(n15698) );
  XOR U17833 ( .A(n18176), .B(n15706), .Z(n15717) );
  XNOR U17834 ( .A(q[7]), .B(DB[352]), .Z(n15706) );
  IV U17835 ( .A(n15705), .Z(n18176) );
  XNOR U17836 ( .A(n15703), .B(n18177), .Z(n15705) );
  XNOR U17837 ( .A(q[6]), .B(DB[351]), .Z(n18177) );
  XNOR U17838 ( .A(q[5]), .B(DB[350]), .Z(n15703) );
  IV U17839 ( .A(n15716), .Z(n18174) );
  XOR U17840 ( .A(n18178), .B(n18179), .Z(n15716) );
  XNOR U17841 ( .A(n15712), .B(n15714), .Z(n18179) );
  XNOR U17842 ( .A(q[1]), .B(DB[346]), .Z(n15714) );
  XNOR U17843 ( .A(q[4]), .B(DB[349]), .Z(n15712) );
  IV U17844 ( .A(n15711), .Z(n18178) );
  XNOR U17845 ( .A(n15709), .B(n18180), .Z(n15711) );
  XNOR U17846 ( .A(q[3]), .B(DB[348]), .Z(n18180) );
  XNOR U17847 ( .A(q[2]), .B(DB[347]), .Z(n15709) );
  XOR U17848 ( .A(n18181), .B(n15607), .Z(n15535) );
  XOR U17849 ( .A(n18182), .B(n15599), .Z(n15607) );
  XOR U17850 ( .A(n18183), .B(n15588), .Z(n15599) );
  XNOR U17851 ( .A(q[14]), .B(DB[374]), .Z(n15588) );
  IV U17852 ( .A(n15587), .Z(n18183) );
  XNOR U17853 ( .A(n15585), .B(n18184), .Z(n15587) );
  XNOR U17854 ( .A(q[13]), .B(DB[373]), .Z(n18184) );
  XNOR U17855 ( .A(q[12]), .B(DB[372]), .Z(n15585) );
  IV U17856 ( .A(n15598), .Z(n18182) );
  XOR U17857 ( .A(n18185), .B(n18186), .Z(n15598) );
  XNOR U17858 ( .A(n15594), .B(n15596), .Z(n18186) );
  XNOR U17859 ( .A(q[8]), .B(DB[368]), .Z(n15596) );
  XNOR U17860 ( .A(q[11]), .B(DB[371]), .Z(n15594) );
  IV U17861 ( .A(n15593), .Z(n18185) );
  XNOR U17862 ( .A(n15591), .B(n18187), .Z(n15593) );
  XNOR U17863 ( .A(q[10]), .B(DB[370]), .Z(n18187) );
  XNOR U17864 ( .A(q[9]), .B(DB[369]), .Z(n15591) );
  IV U17865 ( .A(n15606), .Z(n18181) );
  XOR U17866 ( .A(n18188), .B(n18189), .Z(n15606) );
  XNOR U17867 ( .A(n15623), .B(n15604), .Z(n18189) );
  XNOR U17868 ( .A(q[0]), .B(DB[360]), .Z(n15604) );
  XOR U17869 ( .A(n18190), .B(n15612), .Z(n15623) );
  XNOR U17870 ( .A(q[7]), .B(DB[367]), .Z(n15612) );
  IV U17871 ( .A(n15611), .Z(n18190) );
  XNOR U17872 ( .A(n15609), .B(n18191), .Z(n15611) );
  XNOR U17873 ( .A(q[6]), .B(DB[366]), .Z(n18191) );
  XNOR U17874 ( .A(q[5]), .B(DB[365]), .Z(n15609) );
  IV U17875 ( .A(n15622), .Z(n18188) );
  XOR U17876 ( .A(n18192), .B(n18193), .Z(n15622) );
  XNOR U17877 ( .A(n15618), .B(n15620), .Z(n18193) );
  XNOR U17878 ( .A(q[1]), .B(DB[361]), .Z(n15620) );
  XNOR U17879 ( .A(q[4]), .B(DB[364]), .Z(n15618) );
  IV U17880 ( .A(n15617), .Z(n18192) );
  XNOR U17881 ( .A(n15615), .B(n18194), .Z(n15617) );
  XNOR U17882 ( .A(q[3]), .B(DB[363]), .Z(n18194) );
  XNOR U17883 ( .A(q[2]), .B(DB[362]), .Z(n15615) );
  XOR U17884 ( .A(n18195), .B(n15513), .Z(n15441) );
  XOR U17885 ( .A(n18196), .B(n15505), .Z(n15513) );
  XOR U17886 ( .A(n18197), .B(n15494), .Z(n15505) );
  XNOR U17887 ( .A(q[14]), .B(DB[389]), .Z(n15494) );
  IV U17888 ( .A(n15493), .Z(n18197) );
  XNOR U17889 ( .A(n15491), .B(n18198), .Z(n15493) );
  XNOR U17890 ( .A(q[13]), .B(DB[388]), .Z(n18198) );
  XNOR U17891 ( .A(q[12]), .B(DB[387]), .Z(n15491) );
  IV U17892 ( .A(n15504), .Z(n18196) );
  XOR U17893 ( .A(n18199), .B(n18200), .Z(n15504) );
  XNOR U17894 ( .A(n15500), .B(n15502), .Z(n18200) );
  XNOR U17895 ( .A(q[8]), .B(DB[383]), .Z(n15502) );
  XNOR U17896 ( .A(q[11]), .B(DB[386]), .Z(n15500) );
  IV U17897 ( .A(n15499), .Z(n18199) );
  XNOR U17898 ( .A(n15497), .B(n18201), .Z(n15499) );
  XNOR U17899 ( .A(q[10]), .B(DB[385]), .Z(n18201) );
  XNOR U17900 ( .A(q[9]), .B(DB[384]), .Z(n15497) );
  IV U17901 ( .A(n15512), .Z(n18195) );
  XOR U17902 ( .A(n18202), .B(n18203), .Z(n15512) );
  XNOR U17903 ( .A(n15529), .B(n15510), .Z(n18203) );
  XNOR U17904 ( .A(q[0]), .B(DB[375]), .Z(n15510) );
  XOR U17905 ( .A(n18204), .B(n15518), .Z(n15529) );
  XNOR U17906 ( .A(q[7]), .B(DB[382]), .Z(n15518) );
  IV U17907 ( .A(n15517), .Z(n18204) );
  XNOR U17908 ( .A(n15515), .B(n18205), .Z(n15517) );
  XNOR U17909 ( .A(q[6]), .B(DB[381]), .Z(n18205) );
  XNOR U17910 ( .A(q[5]), .B(DB[380]), .Z(n15515) );
  IV U17911 ( .A(n15528), .Z(n18202) );
  XOR U17912 ( .A(n18206), .B(n18207), .Z(n15528) );
  XNOR U17913 ( .A(n15524), .B(n15526), .Z(n18207) );
  XNOR U17914 ( .A(q[1]), .B(DB[376]), .Z(n15526) );
  XNOR U17915 ( .A(q[4]), .B(DB[379]), .Z(n15524) );
  IV U17916 ( .A(n15523), .Z(n18206) );
  XNOR U17917 ( .A(n15521), .B(n18208), .Z(n15523) );
  XNOR U17918 ( .A(q[3]), .B(DB[378]), .Z(n18208) );
  XNOR U17919 ( .A(q[2]), .B(DB[377]), .Z(n15521) );
  XOR U17920 ( .A(n18209), .B(n15419), .Z(n15347) );
  XOR U17921 ( .A(n18210), .B(n15411), .Z(n15419) );
  XOR U17922 ( .A(n18211), .B(n15400), .Z(n15411) );
  XNOR U17923 ( .A(q[14]), .B(DB[404]), .Z(n15400) );
  IV U17924 ( .A(n15399), .Z(n18211) );
  XNOR U17925 ( .A(n15397), .B(n18212), .Z(n15399) );
  XNOR U17926 ( .A(q[13]), .B(DB[403]), .Z(n18212) );
  XNOR U17927 ( .A(q[12]), .B(DB[402]), .Z(n15397) );
  IV U17928 ( .A(n15410), .Z(n18210) );
  XOR U17929 ( .A(n18213), .B(n18214), .Z(n15410) );
  XNOR U17930 ( .A(n15406), .B(n15408), .Z(n18214) );
  XNOR U17931 ( .A(q[8]), .B(DB[398]), .Z(n15408) );
  XNOR U17932 ( .A(q[11]), .B(DB[401]), .Z(n15406) );
  IV U17933 ( .A(n15405), .Z(n18213) );
  XNOR U17934 ( .A(n15403), .B(n18215), .Z(n15405) );
  XNOR U17935 ( .A(q[10]), .B(DB[400]), .Z(n18215) );
  XNOR U17936 ( .A(q[9]), .B(DB[399]), .Z(n15403) );
  IV U17937 ( .A(n15418), .Z(n18209) );
  XOR U17938 ( .A(n18216), .B(n18217), .Z(n15418) );
  XNOR U17939 ( .A(n15435), .B(n15416), .Z(n18217) );
  XNOR U17940 ( .A(q[0]), .B(DB[390]), .Z(n15416) );
  XOR U17941 ( .A(n18218), .B(n15424), .Z(n15435) );
  XNOR U17942 ( .A(q[7]), .B(DB[397]), .Z(n15424) );
  IV U17943 ( .A(n15423), .Z(n18218) );
  XNOR U17944 ( .A(n15421), .B(n18219), .Z(n15423) );
  XNOR U17945 ( .A(q[6]), .B(DB[396]), .Z(n18219) );
  XNOR U17946 ( .A(q[5]), .B(DB[395]), .Z(n15421) );
  IV U17947 ( .A(n15434), .Z(n18216) );
  XOR U17948 ( .A(n18220), .B(n18221), .Z(n15434) );
  XNOR U17949 ( .A(n15430), .B(n15432), .Z(n18221) );
  XNOR U17950 ( .A(q[1]), .B(DB[391]), .Z(n15432) );
  XNOR U17951 ( .A(q[4]), .B(DB[394]), .Z(n15430) );
  IV U17952 ( .A(n15429), .Z(n18220) );
  XNOR U17953 ( .A(n15427), .B(n18222), .Z(n15429) );
  XNOR U17954 ( .A(q[3]), .B(DB[393]), .Z(n18222) );
  XNOR U17955 ( .A(q[2]), .B(DB[392]), .Z(n15427) );
  XOR U17956 ( .A(n18223), .B(n15325), .Z(n15253) );
  XOR U17957 ( .A(n18224), .B(n15317), .Z(n15325) );
  XOR U17958 ( .A(n18225), .B(n15306), .Z(n15317) );
  XNOR U17959 ( .A(q[14]), .B(DB[419]), .Z(n15306) );
  IV U17960 ( .A(n15305), .Z(n18225) );
  XNOR U17961 ( .A(n15303), .B(n18226), .Z(n15305) );
  XNOR U17962 ( .A(q[13]), .B(DB[418]), .Z(n18226) );
  XNOR U17963 ( .A(q[12]), .B(DB[417]), .Z(n15303) );
  IV U17964 ( .A(n15316), .Z(n18224) );
  XOR U17965 ( .A(n18227), .B(n18228), .Z(n15316) );
  XNOR U17966 ( .A(n15312), .B(n15314), .Z(n18228) );
  XNOR U17967 ( .A(q[8]), .B(DB[413]), .Z(n15314) );
  XNOR U17968 ( .A(q[11]), .B(DB[416]), .Z(n15312) );
  IV U17969 ( .A(n15311), .Z(n18227) );
  XNOR U17970 ( .A(n15309), .B(n18229), .Z(n15311) );
  XNOR U17971 ( .A(q[10]), .B(DB[415]), .Z(n18229) );
  XNOR U17972 ( .A(q[9]), .B(DB[414]), .Z(n15309) );
  IV U17973 ( .A(n15324), .Z(n18223) );
  XOR U17974 ( .A(n18230), .B(n18231), .Z(n15324) );
  XNOR U17975 ( .A(n15341), .B(n15322), .Z(n18231) );
  XNOR U17976 ( .A(q[0]), .B(DB[405]), .Z(n15322) );
  XOR U17977 ( .A(n18232), .B(n15330), .Z(n15341) );
  XNOR U17978 ( .A(q[7]), .B(DB[412]), .Z(n15330) );
  IV U17979 ( .A(n15329), .Z(n18232) );
  XNOR U17980 ( .A(n15327), .B(n18233), .Z(n15329) );
  XNOR U17981 ( .A(q[6]), .B(DB[411]), .Z(n18233) );
  XNOR U17982 ( .A(q[5]), .B(DB[410]), .Z(n15327) );
  IV U17983 ( .A(n15340), .Z(n18230) );
  XOR U17984 ( .A(n18234), .B(n18235), .Z(n15340) );
  XNOR U17985 ( .A(n15336), .B(n15338), .Z(n18235) );
  XNOR U17986 ( .A(q[1]), .B(DB[406]), .Z(n15338) );
  XNOR U17987 ( .A(q[4]), .B(DB[409]), .Z(n15336) );
  IV U17988 ( .A(n15335), .Z(n18234) );
  XNOR U17989 ( .A(n15333), .B(n18236), .Z(n15335) );
  XNOR U17990 ( .A(q[3]), .B(DB[408]), .Z(n18236) );
  XNOR U17991 ( .A(q[2]), .B(DB[407]), .Z(n15333) );
  XOR U17992 ( .A(n18237), .B(n15231), .Z(n15159) );
  XOR U17993 ( .A(n18238), .B(n15223), .Z(n15231) );
  XOR U17994 ( .A(n18239), .B(n15212), .Z(n15223) );
  XNOR U17995 ( .A(q[14]), .B(DB[434]), .Z(n15212) );
  IV U17996 ( .A(n15211), .Z(n18239) );
  XNOR U17997 ( .A(n15209), .B(n18240), .Z(n15211) );
  XNOR U17998 ( .A(q[13]), .B(DB[433]), .Z(n18240) );
  XNOR U17999 ( .A(q[12]), .B(DB[432]), .Z(n15209) );
  IV U18000 ( .A(n15222), .Z(n18238) );
  XOR U18001 ( .A(n18241), .B(n18242), .Z(n15222) );
  XNOR U18002 ( .A(n15218), .B(n15220), .Z(n18242) );
  XNOR U18003 ( .A(q[8]), .B(DB[428]), .Z(n15220) );
  XNOR U18004 ( .A(q[11]), .B(DB[431]), .Z(n15218) );
  IV U18005 ( .A(n15217), .Z(n18241) );
  XNOR U18006 ( .A(n15215), .B(n18243), .Z(n15217) );
  XNOR U18007 ( .A(q[10]), .B(DB[430]), .Z(n18243) );
  XNOR U18008 ( .A(q[9]), .B(DB[429]), .Z(n15215) );
  IV U18009 ( .A(n15230), .Z(n18237) );
  XOR U18010 ( .A(n18244), .B(n18245), .Z(n15230) );
  XNOR U18011 ( .A(n15247), .B(n15228), .Z(n18245) );
  XNOR U18012 ( .A(q[0]), .B(DB[420]), .Z(n15228) );
  XOR U18013 ( .A(n18246), .B(n15236), .Z(n15247) );
  XNOR U18014 ( .A(q[7]), .B(DB[427]), .Z(n15236) );
  IV U18015 ( .A(n15235), .Z(n18246) );
  XNOR U18016 ( .A(n15233), .B(n18247), .Z(n15235) );
  XNOR U18017 ( .A(q[6]), .B(DB[426]), .Z(n18247) );
  XNOR U18018 ( .A(q[5]), .B(DB[425]), .Z(n15233) );
  IV U18019 ( .A(n15246), .Z(n18244) );
  XOR U18020 ( .A(n18248), .B(n18249), .Z(n15246) );
  XNOR U18021 ( .A(n15242), .B(n15244), .Z(n18249) );
  XNOR U18022 ( .A(q[1]), .B(DB[421]), .Z(n15244) );
  XNOR U18023 ( .A(q[4]), .B(DB[424]), .Z(n15242) );
  IV U18024 ( .A(n15241), .Z(n18248) );
  XNOR U18025 ( .A(n15239), .B(n18250), .Z(n15241) );
  XNOR U18026 ( .A(q[3]), .B(DB[423]), .Z(n18250) );
  XNOR U18027 ( .A(q[2]), .B(DB[422]), .Z(n15239) );
  XOR U18028 ( .A(n18251), .B(n15137), .Z(n15065) );
  XOR U18029 ( .A(n18252), .B(n15129), .Z(n15137) );
  XOR U18030 ( .A(n18253), .B(n15118), .Z(n15129) );
  XNOR U18031 ( .A(q[14]), .B(DB[449]), .Z(n15118) );
  IV U18032 ( .A(n15117), .Z(n18253) );
  XNOR U18033 ( .A(n15115), .B(n18254), .Z(n15117) );
  XNOR U18034 ( .A(q[13]), .B(DB[448]), .Z(n18254) );
  XNOR U18035 ( .A(q[12]), .B(DB[447]), .Z(n15115) );
  IV U18036 ( .A(n15128), .Z(n18252) );
  XOR U18037 ( .A(n18255), .B(n18256), .Z(n15128) );
  XNOR U18038 ( .A(n15124), .B(n15126), .Z(n18256) );
  XNOR U18039 ( .A(q[8]), .B(DB[443]), .Z(n15126) );
  XNOR U18040 ( .A(q[11]), .B(DB[446]), .Z(n15124) );
  IV U18041 ( .A(n15123), .Z(n18255) );
  XNOR U18042 ( .A(n15121), .B(n18257), .Z(n15123) );
  XNOR U18043 ( .A(q[10]), .B(DB[445]), .Z(n18257) );
  XNOR U18044 ( .A(q[9]), .B(DB[444]), .Z(n15121) );
  IV U18045 ( .A(n15136), .Z(n18251) );
  XOR U18046 ( .A(n18258), .B(n18259), .Z(n15136) );
  XNOR U18047 ( .A(n15153), .B(n15134), .Z(n18259) );
  XNOR U18048 ( .A(q[0]), .B(DB[435]), .Z(n15134) );
  XOR U18049 ( .A(n18260), .B(n15142), .Z(n15153) );
  XNOR U18050 ( .A(q[7]), .B(DB[442]), .Z(n15142) );
  IV U18051 ( .A(n15141), .Z(n18260) );
  XNOR U18052 ( .A(n15139), .B(n18261), .Z(n15141) );
  XNOR U18053 ( .A(q[6]), .B(DB[441]), .Z(n18261) );
  XNOR U18054 ( .A(q[5]), .B(DB[440]), .Z(n15139) );
  IV U18055 ( .A(n15152), .Z(n18258) );
  XOR U18056 ( .A(n18262), .B(n18263), .Z(n15152) );
  XNOR U18057 ( .A(n15148), .B(n15150), .Z(n18263) );
  XNOR U18058 ( .A(q[1]), .B(DB[436]), .Z(n15150) );
  XNOR U18059 ( .A(q[4]), .B(DB[439]), .Z(n15148) );
  IV U18060 ( .A(n15147), .Z(n18262) );
  XNOR U18061 ( .A(n15145), .B(n18264), .Z(n15147) );
  XNOR U18062 ( .A(q[3]), .B(DB[438]), .Z(n18264) );
  XNOR U18063 ( .A(q[2]), .B(DB[437]), .Z(n15145) );
  XOR U18064 ( .A(n18265), .B(n15043), .Z(n14971) );
  XOR U18065 ( .A(n18266), .B(n15035), .Z(n15043) );
  XOR U18066 ( .A(n18267), .B(n15024), .Z(n15035) );
  XNOR U18067 ( .A(q[14]), .B(DB[464]), .Z(n15024) );
  IV U18068 ( .A(n15023), .Z(n18267) );
  XNOR U18069 ( .A(n15021), .B(n18268), .Z(n15023) );
  XNOR U18070 ( .A(q[13]), .B(DB[463]), .Z(n18268) );
  XNOR U18071 ( .A(q[12]), .B(DB[462]), .Z(n15021) );
  IV U18072 ( .A(n15034), .Z(n18266) );
  XOR U18073 ( .A(n18269), .B(n18270), .Z(n15034) );
  XNOR U18074 ( .A(n15030), .B(n15032), .Z(n18270) );
  XNOR U18075 ( .A(q[8]), .B(DB[458]), .Z(n15032) );
  XNOR U18076 ( .A(q[11]), .B(DB[461]), .Z(n15030) );
  IV U18077 ( .A(n15029), .Z(n18269) );
  XNOR U18078 ( .A(n15027), .B(n18271), .Z(n15029) );
  XNOR U18079 ( .A(q[10]), .B(DB[460]), .Z(n18271) );
  XNOR U18080 ( .A(q[9]), .B(DB[459]), .Z(n15027) );
  IV U18081 ( .A(n15042), .Z(n18265) );
  XOR U18082 ( .A(n18272), .B(n18273), .Z(n15042) );
  XNOR U18083 ( .A(n15059), .B(n15040), .Z(n18273) );
  XNOR U18084 ( .A(q[0]), .B(DB[450]), .Z(n15040) );
  XOR U18085 ( .A(n18274), .B(n15048), .Z(n15059) );
  XNOR U18086 ( .A(q[7]), .B(DB[457]), .Z(n15048) );
  IV U18087 ( .A(n15047), .Z(n18274) );
  XNOR U18088 ( .A(n15045), .B(n18275), .Z(n15047) );
  XNOR U18089 ( .A(q[6]), .B(DB[456]), .Z(n18275) );
  XNOR U18090 ( .A(q[5]), .B(DB[455]), .Z(n15045) );
  IV U18091 ( .A(n15058), .Z(n18272) );
  XOR U18092 ( .A(n18276), .B(n18277), .Z(n15058) );
  XNOR U18093 ( .A(n15054), .B(n15056), .Z(n18277) );
  XNOR U18094 ( .A(q[1]), .B(DB[451]), .Z(n15056) );
  XNOR U18095 ( .A(q[4]), .B(DB[454]), .Z(n15054) );
  IV U18096 ( .A(n15053), .Z(n18276) );
  XNOR U18097 ( .A(n15051), .B(n18278), .Z(n15053) );
  XNOR U18098 ( .A(q[3]), .B(DB[453]), .Z(n18278) );
  XNOR U18099 ( .A(q[2]), .B(DB[452]), .Z(n15051) );
  XOR U18100 ( .A(n18279), .B(n14949), .Z(n14877) );
  XOR U18101 ( .A(n18280), .B(n14941), .Z(n14949) );
  XOR U18102 ( .A(n18281), .B(n14930), .Z(n14941) );
  XNOR U18103 ( .A(q[14]), .B(DB[479]), .Z(n14930) );
  IV U18104 ( .A(n14929), .Z(n18281) );
  XNOR U18105 ( .A(n14927), .B(n18282), .Z(n14929) );
  XNOR U18106 ( .A(q[13]), .B(DB[478]), .Z(n18282) );
  XNOR U18107 ( .A(q[12]), .B(DB[477]), .Z(n14927) );
  IV U18108 ( .A(n14940), .Z(n18280) );
  XOR U18109 ( .A(n18283), .B(n18284), .Z(n14940) );
  XNOR U18110 ( .A(n14936), .B(n14938), .Z(n18284) );
  XNOR U18111 ( .A(q[8]), .B(DB[473]), .Z(n14938) );
  XNOR U18112 ( .A(q[11]), .B(DB[476]), .Z(n14936) );
  IV U18113 ( .A(n14935), .Z(n18283) );
  XNOR U18114 ( .A(n14933), .B(n18285), .Z(n14935) );
  XNOR U18115 ( .A(q[10]), .B(DB[475]), .Z(n18285) );
  XNOR U18116 ( .A(q[9]), .B(DB[474]), .Z(n14933) );
  IV U18117 ( .A(n14948), .Z(n18279) );
  XOR U18118 ( .A(n18286), .B(n18287), .Z(n14948) );
  XNOR U18119 ( .A(n14965), .B(n14946), .Z(n18287) );
  XNOR U18120 ( .A(q[0]), .B(DB[465]), .Z(n14946) );
  XOR U18121 ( .A(n18288), .B(n14954), .Z(n14965) );
  XNOR U18122 ( .A(q[7]), .B(DB[472]), .Z(n14954) );
  IV U18123 ( .A(n14953), .Z(n18288) );
  XNOR U18124 ( .A(n14951), .B(n18289), .Z(n14953) );
  XNOR U18125 ( .A(q[6]), .B(DB[471]), .Z(n18289) );
  XNOR U18126 ( .A(q[5]), .B(DB[470]), .Z(n14951) );
  IV U18127 ( .A(n14964), .Z(n18286) );
  XOR U18128 ( .A(n18290), .B(n18291), .Z(n14964) );
  XNOR U18129 ( .A(n14960), .B(n14962), .Z(n18291) );
  XNOR U18130 ( .A(q[1]), .B(DB[466]), .Z(n14962) );
  XNOR U18131 ( .A(q[4]), .B(DB[469]), .Z(n14960) );
  IV U18132 ( .A(n14959), .Z(n18290) );
  XNOR U18133 ( .A(n14957), .B(n18292), .Z(n14959) );
  XNOR U18134 ( .A(q[3]), .B(DB[468]), .Z(n18292) );
  XNOR U18135 ( .A(q[2]), .B(DB[467]), .Z(n14957) );
  XOR U18136 ( .A(n18293), .B(n14855), .Z(n14783) );
  XOR U18137 ( .A(n18294), .B(n14847), .Z(n14855) );
  XOR U18138 ( .A(n18295), .B(n14836), .Z(n14847) );
  XNOR U18139 ( .A(q[14]), .B(DB[494]), .Z(n14836) );
  IV U18140 ( .A(n14835), .Z(n18295) );
  XNOR U18141 ( .A(n14833), .B(n18296), .Z(n14835) );
  XNOR U18142 ( .A(q[13]), .B(DB[493]), .Z(n18296) );
  XNOR U18143 ( .A(q[12]), .B(DB[492]), .Z(n14833) );
  IV U18144 ( .A(n14846), .Z(n18294) );
  XOR U18145 ( .A(n18297), .B(n18298), .Z(n14846) );
  XNOR U18146 ( .A(n14842), .B(n14844), .Z(n18298) );
  XNOR U18147 ( .A(q[8]), .B(DB[488]), .Z(n14844) );
  XNOR U18148 ( .A(q[11]), .B(DB[491]), .Z(n14842) );
  IV U18149 ( .A(n14841), .Z(n18297) );
  XNOR U18150 ( .A(n14839), .B(n18299), .Z(n14841) );
  XNOR U18151 ( .A(q[10]), .B(DB[490]), .Z(n18299) );
  XNOR U18152 ( .A(q[9]), .B(DB[489]), .Z(n14839) );
  IV U18153 ( .A(n14854), .Z(n18293) );
  XOR U18154 ( .A(n18300), .B(n18301), .Z(n14854) );
  XNOR U18155 ( .A(n14871), .B(n14852), .Z(n18301) );
  XNOR U18156 ( .A(q[0]), .B(DB[480]), .Z(n14852) );
  XOR U18157 ( .A(n18302), .B(n14860), .Z(n14871) );
  XNOR U18158 ( .A(q[7]), .B(DB[487]), .Z(n14860) );
  IV U18159 ( .A(n14859), .Z(n18302) );
  XNOR U18160 ( .A(n14857), .B(n18303), .Z(n14859) );
  XNOR U18161 ( .A(q[6]), .B(DB[486]), .Z(n18303) );
  XNOR U18162 ( .A(q[5]), .B(DB[485]), .Z(n14857) );
  IV U18163 ( .A(n14870), .Z(n18300) );
  XOR U18164 ( .A(n18304), .B(n18305), .Z(n14870) );
  XNOR U18165 ( .A(n14866), .B(n14868), .Z(n18305) );
  XNOR U18166 ( .A(q[1]), .B(DB[481]), .Z(n14868) );
  XNOR U18167 ( .A(q[4]), .B(DB[484]), .Z(n14866) );
  IV U18168 ( .A(n14865), .Z(n18304) );
  XNOR U18169 ( .A(n14863), .B(n18306), .Z(n14865) );
  XNOR U18170 ( .A(q[3]), .B(DB[483]), .Z(n18306) );
  XNOR U18171 ( .A(q[2]), .B(DB[482]), .Z(n14863) );
  XOR U18172 ( .A(n18307), .B(n14761), .Z(n14689) );
  XOR U18173 ( .A(n18308), .B(n14753), .Z(n14761) );
  XOR U18174 ( .A(n18309), .B(n14742), .Z(n14753) );
  XNOR U18175 ( .A(q[14]), .B(DB[509]), .Z(n14742) );
  IV U18176 ( .A(n14741), .Z(n18309) );
  XNOR U18177 ( .A(n14739), .B(n18310), .Z(n14741) );
  XNOR U18178 ( .A(q[13]), .B(DB[508]), .Z(n18310) );
  XNOR U18179 ( .A(q[12]), .B(DB[507]), .Z(n14739) );
  IV U18180 ( .A(n14752), .Z(n18308) );
  XOR U18181 ( .A(n18311), .B(n18312), .Z(n14752) );
  XNOR U18182 ( .A(n14748), .B(n14750), .Z(n18312) );
  XNOR U18183 ( .A(q[8]), .B(DB[503]), .Z(n14750) );
  XNOR U18184 ( .A(q[11]), .B(DB[506]), .Z(n14748) );
  IV U18185 ( .A(n14747), .Z(n18311) );
  XNOR U18186 ( .A(n14745), .B(n18313), .Z(n14747) );
  XNOR U18187 ( .A(q[10]), .B(DB[505]), .Z(n18313) );
  XNOR U18188 ( .A(q[9]), .B(DB[504]), .Z(n14745) );
  IV U18189 ( .A(n14760), .Z(n18307) );
  XOR U18190 ( .A(n18314), .B(n18315), .Z(n14760) );
  XNOR U18191 ( .A(n14777), .B(n14758), .Z(n18315) );
  XNOR U18192 ( .A(q[0]), .B(DB[495]), .Z(n14758) );
  XOR U18193 ( .A(n18316), .B(n14766), .Z(n14777) );
  XNOR U18194 ( .A(q[7]), .B(DB[502]), .Z(n14766) );
  IV U18195 ( .A(n14765), .Z(n18316) );
  XNOR U18196 ( .A(n14763), .B(n18317), .Z(n14765) );
  XNOR U18197 ( .A(q[6]), .B(DB[501]), .Z(n18317) );
  XNOR U18198 ( .A(q[5]), .B(DB[500]), .Z(n14763) );
  IV U18199 ( .A(n14776), .Z(n18314) );
  XOR U18200 ( .A(n18318), .B(n18319), .Z(n14776) );
  XNOR U18201 ( .A(n14772), .B(n14774), .Z(n18319) );
  XNOR U18202 ( .A(q[1]), .B(DB[496]), .Z(n14774) );
  XNOR U18203 ( .A(q[4]), .B(DB[499]), .Z(n14772) );
  IV U18204 ( .A(n14771), .Z(n18318) );
  XNOR U18205 ( .A(n14769), .B(n18320), .Z(n14771) );
  XNOR U18206 ( .A(q[3]), .B(DB[498]), .Z(n18320) );
  XNOR U18207 ( .A(q[2]), .B(DB[497]), .Z(n14769) );
  XOR U18208 ( .A(n18321), .B(n14667), .Z(n14595) );
  XOR U18209 ( .A(n18322), .B(n14659), .Z(n14667) );
  XOR U18210 ( .A(n18323), .B(n14648), .Z(n14659) );
  XNOR U18211 ( .A(q[14]), .B(DB[524]), .Z(n14648) );
  IV U18212 ( .A(n14647), .Z(n18323) );
  XNOR U18213 ( .A(n14645), .B(n18324), .Z(n14647) );
  XNOR U18214 ( .A(q[13]), .B(DB[523]), .Z(n18324) );
  XNOR U18215 ( .A(q[12]), .B(DB[522]), .Z(n14645) );
  IV U18216 ( .A(n14658), .Z(n18322) );
  XOR U18217 ( .A(n18325), .B(n18326), .Z(n14658) );
  XNOR U18218 ( .A(n14654), .B(n14656), .Z(n18326) );
  XNOR U18219 ( .A(q[8]), .B(DB[518]), .Z(n14656) );
  XNOR U18220 ( .A(q[11]), .B(DB[521]), .Z(n14654) );
  IV U18221 ( .A(n14653), .Z(n18325) );
  XNOR U18222 ( .A(n14651), .B(n18327), .Z(n14653) );
  XNOR U18223 ( .A(q[10]), .B(DB[520]), .Z(n18327) );
  XNOR U18224 ( .A(q[9]), .B(DB[519]), .Z(n14651) );
  IV U18225 ( .A(n14666), .Z(n18321) );
  XOR U18226 ( .A(n18328), .B(n18329), .Z(n14666) );
  XNOR U18227 ( .A(n14683), .B(n14664), .Z(n18329) );
  XNOR U18228 ( .A(q[0]), .B(DB[510]), .Z(n14664) );
  XOR U18229 ( .A(n18330), .B(n14672), .Z(n14683) );
  XNOR U18230 ( .A(q[7]), .B(DB[517]), .Z(n14672) );
  IV U18231 ( .A(n14671), .Z(n18330) );
  XNOR U18232 ( .A(n14669), .B(n18331), .Z(n14671) );
  XNOR U18233 ( .A(q[6]), .B(DB[516]), .Z(n18331) );
  XNOR U18234 ( .A(q[5]), .B(DB[515]), .Z(n14669) );
  IV U18235 ( .A(n14682), .Z(n18328) );
  XOR U18236 ( .A(n18332), .B(n18333), .Z(n14682) );
  XNOR U18237 ( .A(n14678), .B(n14680), .Z(n18333) );
  XNOR U18238 ( .A(q[1]), .B(DB[511]), .Z(n14680) );
  XNOR U18239 ( .A(q[4]), .B(DB[514]), .Z(n14678) );
  IV U18240 ( .A(n14677), .Z(n18332) );
  XNOR U18241 ( .A(n14675), .B(n18334), .Z(n14677) );
  XNOR U18242 ( .A(q[3]), .B(DB[513]), .Z(n18334) );
  XNOR U18243 ( .A(q[2]), .B(DB[512]), .Z(n14675) );
  XOR U18244 ( .A(n18335), .B(n14573), .Z(n14501) );
  XOR U18245 ( .A(n18336), .B(n14565), .Z(n14573) );
  XOR U18246 ( .A(n18337), .B(n14554), .Z(n14565) );
  XNOR U18247 ( .A(q[14]), .B(DB[539]), .Z(n14554) );
  IV U18248 ( .A(n14553), .Z(n18337) );
  XNOR U18249 ( .A(n14551), .B(n18338), .Z(n14553) );
  XNOR U18250 ( .A(q[13]), .B(DB[538]), .Z(n18338) );
  XNOR U18251 ( .A(q[12]), .B(DB[537]), .Z(n14551) );
  IV U18252 ( .A(n14564), .Z(n18336) );
  XOR U18253 ( .A(n18339), .B(n18340), .Z(n14564) );
  XNOR U18254 ( .A(n14560), .B(n14562), .Z(n18340) );
  XNOR U18255 ( .A(q[8]), .B(DB[533]), .Z(n14562) );
  XNOR U18256 ( .A(q[11]), .B(DB[536]), .Z(n14560) );
  IV U18257 ( .A(n14559), .Z(n18339) );
  XNOR U18258 ( .A(n14557), .B(n18341), .Z(n14559) );
  XNOR U18259 ( .A(q[10]), .B(DB[535]), .Z(n18341) );
  XNOR U18260 ( .A(q[9]), .B(DB[534]), .Z(n14557) );
  IV U18261 ( .A(n14572), .Z(n18335) );
  XOR U18262 ( .A(n18342), .B(n18343), .Z(n14572) );
  XNOR U18263 ( .A(n14589), .B(n14570), .Z(n18343) );
  XNOR U18264 ( .A(q[0]), .B(DB[525]), .Z(n14570) );
  XOR U18265 ( .A(n18344), .B(n14578), .Z(n14589) );
  XNOR U18266 ( .A(q[7]), .B(DB[532]), .Z(n14578) );
  IV U18267 ( .A(n14577), .Z(n18344) );
  XNOR U18268 ( .A(n14575), .B(n18345), .Z(n14577) );
  XNOR U18269 ( .A(q[6]), .B(DB[531]), .Z(n18345) );
  XNOR U18270 ( .A(q[5]), .B(DB[530]), .Z(n14575) );
  IV U18271 ( .A(n14588), .Z(n18342) );
  XOR U18272 ( .A(n18346), .B(n18347), .Z(n14588) );
  XNOR U18273 ( .A(n14584), .B(n14586), .Z(n18347) );
  XNOR U18274 ( .A(q[1]), .B(DB[526]), .Z(n14586) );
  XNOR U18275 ( .A(q[4]), .B(DB[529]), .Z(n14584) );
  IV U18276 ( .A(n14583), .Z(n18346) );
  XNOR U18277 ( .A(n14581), .B(n18348), .Z(n14583) );
  XNOR U18278 ( .A(q[3]), .B(DB[528]), .Z(n18348) );
  XNOR U18279 ( .A(q[2]), .B(DB[527]), .Z(n14581) );
  XOR U18280 ( .A(n18349), .B(n14479), .Z(n14407) );
  XOR U18281 ( .A(n18350), .B(n14471), .Z(n14479) );
  XOR U18282 ( .A(n18351), .B(n14460), .Z(n14471) );
  XNOR U18283 ( .A(q[14]), .B(DB[554]), .Z(n14460) );
  IV U18284 ( .A(n14459), .Z(n18351) );
  XNOR U18285 ( .A(n14457), .B(n18352), .Z(n14459) );
  XNOR U18286 ( .A(q[13]), .B(DB[553]), .Z(n18352) );
  XNOR U18287 ( .A(q[12]), .B(DB[552]), .Z(n14457) );
  IV U18288 ( .A(n14470), .Z(n18350) );
  XOR U18289 ( .A(n18353), .B(n18354), .Z(n14470) );
  XNOR U18290 ( .A(n14466), .B(n14468), .Z(n18354) );
  XNOR U18291 ( .A(q[8]), .B(DB[548]), .Z(n14468) );
  XNOR U18292 ( .A(q[11]), .B(DB[551]), .Z(n14466) );
  IV U18293 ( .A(n14465), .Z(n18353) );
  XNOR U18294 ( .A(n14463), .B(n18355), .Z(n14465) );
  XNOR U18295 ( .A(q[10]), .B(DB[550]), .Z(n18355) );
  XNOR U18296 ( .A(q[9]), .B(DB[549]), .Z(n14463) );
  IV U18297 ( .A(n14478), .Z(n18349) );
  XOR U18298 ( .A(n18356), .B(n18357), .Z(n14478) );
  XNOR U18299 ( .A(n14495), .B(n14476), .Z(n18357) );
  XNOR U18300 ( .A(q[0]), .B(DB[540]), .Z(n14476) );
  XOR U18301 ( .A(n18358), .B(n14484), .Z(n14495) );
  XNOR U18302 ( .A(q[7]), .B(DB[547]), .Z(n14484) );
  IV U18303 ( .A(n14483), .Z(n18358) );
  XNOR U18304 ( .A(n14481), .B(n18359), .Z(n14483) );
  XNOR U18305 ( .A(q[6]), .B(DB[546]), .Z(n18359) );
  XNOR U18306 ( .A(q[5]), .B(DB[545]), .Z(n14481) );
  IV U18307 ( .A(n14494), .Z(n18356) );
  XOR U18308 ( .A(n18360), .B(n18361), .Z(n14494) );
  XNOR U18309 ( .A(n14490), .B(n14492), .Z(n18361) );
  XNOR U18310 ( .A(q[1]), .B(DB[541]), .Z(n14492) );
  XNOR U18311 ( .A(q[4]), .B(DB[544]), .Z(n14490) );
  IV U18312 ( .A(n14489), .Z(n18360) );
  XNOR U18313 ( .A(n14487), .B(n18362), .Z(n14489) );
  XNOR U18314 ( .A(q[3]), .B(DB[543]), .Z(n18362) );
  XNOR U18315 ( .A(q[2]), .B(DB[542]), .Z(n14487) );
  XOR U18316 ( .A(n18363), .B(n14385), .Z(n14313) );
  XOR U18317 ( .A(n18364), .B(n14377), .Z(n14385) );
  XOR U18318 ( .A(n18365), .B(n14366), .Z(n14377) );
  XNOR U18319 ( .A(q[14]), .B(DB[569]), .Z(n14366) );
  IV U18320 ( .A(n14365), .Z(n18365) );
  XNOR U18321 ( .A(n14363), .B(n18366), .Z(n14365) );
  XNOR U18322 ( .A(q[13]), .B(DB[568]), .Z(n18366) );
  XNOR U18323 ( .A(q[12]), .B(DB[567]), .Z(n14363) );
  IV U18324 ( .A(n14376), .Z(n18364) );
  XOR U18325 ( .A(n18367), .B(n18368), .Z(n14376) );
  XNOR U18326 ( .A(n14372), .B(n14374), .Z(n18368) );
  XNOR U18327 ( .A(q[8]), .B(DB[563]), .Z(n14374) );
  XNOR U18328 ( .A(q[11]), .B(DB[566]), .Z(n14372) );
  IV U18329 ( .A(n14371), .Z(n18367) );
  XNOR U18330 ( .A(n14369), .B(n18369), .Z(n14371) );
  XNOR U18331 ( .A(q[10]), .B(DB[565]), .Z(n18369) );
  XNOR U18332 ( .A(q[9]), .B(DB[564]), .Z(n14369) );
  IV U18333 ( .A(n14384), .Z(n18363) );
  XOR U18334 ( .A(n18370), .B(n18371), .Z(n14384) );
  XNOR U18335 ( .A(n14401), .B(n14382), .Z(n18371) );
  XNOR U18336 ( .A(q[0]), .B(DB[555]), .Z(n14382) );
  XOR U18337 ( .A(n18372), .B(n14390), .Z(n14401) );
  XNOR U18338 ( .A(q[7]), .B(DB[562]), .Z(n14390) );
  IV U18339 ( .A(n14389), .Z(n18372) );
  XNOR U18340 ( .A(n14387), .B(n18373), .Z(n14389) );
  XNOR U18341 ( .A(q[6]), .B(DB[561]), .Z(n18373) );
  XNOR U18342 ( .A(q[5]), .B(DB[560]), .Z(n14387) );
  IV U18343 ( .A(n14400), .Z(n18370) );
  XOR U18344 ( .A(n18374), .B(n18375), .Z(n14400) );
  XNOR U18345 ( .A(n14396), .B(n14398), .Z(n18375) );
  XNOR U18346 ( .A(q[1]), .B(DB[556]), .Z(n14398) );
  XNOR U18347 ( .A(q[4]), .B(DB[559]), .Z(n14396) );
  IV U18348 ( .A(n14395), .Z(n18374) );
  XNOR U18349 ( .A(n14393), .B(n18376), .Z(n14395) );
  XNOR U18350 ( .A(q[3]), .B(DB[558]), .Z(n18376) );
  XNOR U18351 ( .A(q[2]), .B(DB[557]), .Z(n14393) );
  XOR U18352 ( .A(n18377), .B(n14291), .Z(n14219) );
  XOR U18353 ( .A(n18378), .B(n14283), .Z(n14291) );
  XOR U18354 ( .A(n18379), .B(n14272), .Z(n14283) );
  XNOR U18355 ( .A(q[14]), .B(DB[584]), .Z(n14272) );
  IV U18356 ( .A(n14271), .Z(n18379) );
  XNOR U18357 ( .A(n14269), .B(n18380), .Z(n14271) );
  XNOR U18358 ( .A(q[13]), .B(DB[583]), .Z(n18380) );
  XNOR U18359 ( .A(q[12]), .B(DB[582]), .Z(n14269) );
  IV U18360 ( .A(n14282), .Z(n18378) );
  XOR U18361 ( .A(n18381), .B(n18382), .Z(n14282) );
  XNOR U18362 ( .A(n14278), .B(n14280), .Z(n18382) );
  XNOR U18363 ( .A(q[8]), .B(DB[578]), .Z(n14280) );
  XNOR U18364 ( .A(q[11]), .B(DB[581]), .Z(n14278) );
  IV U18365 ( .A(n14277), .Z(n18381) );
  XNOR U18366 ( .A(n14275), .B(n18383), .Z(n14277) );
  XNOR U18367 ( .A(q[10]), .B(DB[580]), .Z(n18383) );
  XNOR U18368 ( .A(q[9]), .B(DB[579]), .Z(n14275) );
  IV U18369 ( .A(n14290), .Z(n18377) );
  XOR U18370 ( .A(n18384), .B(n18385), .Z(n14290) );
  XNOR U18371 ( .A(n14307), .B(n14288), .Z(n18385) );
  XNOR U18372 ( .A(q[0]), .B(DB[570]), .Z(n14288) );
  XOR U18373 ( .A(n18386), .B(n14296), .Z(n14307) );
  XNOR U18374 ( .A(q[7]), .B(DB[577]), .Z(n14296) );
  IV U18375 ( .A(n14295), .Z(n18386) );
  XNOR U18376 ( .A(n14293), .B(n18387), .Z(n14295) );
  XNOR U18377 ( .A(q[6]), .B(DB[576]), .Z(n18387) );
  XNOR U18378 ( .A(q[5]), .B(DB[575]), .Z(n14293) );
  IV U18379 ( .A(n14306), .Z(n18384) );
  XOR U18380 ( .A(n18388), .B(n18389), .Z(n14306) );
  XNOR U18381 ( .A(n14302), .B(n14304), .Z(n18389) );
  XNOR U18382 ( .A(q[1]), .B(DB[571]), .Z(n14304) );
  XNOR U18383 ( .A(q[4]), .B(DB[574]), .Z(n14302) );
  IV U18384 ( .A(n14301), .Z(n18388) );
  XNOR U18385 ( .A(n14299), .B(n18390), .Z(n14301) );
  XNOR U18386 ( .A(q[3]), .B(DB[573]), .Z(n18390) );
  XNOR U18387 ( .A(q[2]), .B(DB[572]), .Z(n14299) );
  XOR U18388 ( .A(n18391), .B(n14197), .Z(n14125) );
  XOR U18389 ( .A(n18392), .B(n14189), .Z(n14197) );
  XOR U18390 ( .A(n18393), .B(n14178), .Z(n14189) );
  XNOR U18391 ( .A(q[14]), .B(DB[599]), .Z(n14178) );
  IV U18392 ( .A(n14177), .Z(n18393) );
  XNOR U18393 ( .A(n14175), .B(n18394), .Z(n14177) );
  XNOR U18394 ( .A(q[13]), .B(DB[598]), .Z(n18394) );
  XNOR U18395 ( .A(q[12]), .B(DB[597]), .Z(n14175) );
  IV U18396 ( .A(n14188), .Z(n18392) );
  XOR U18397 ( .A(n18395), .B(n18396), .Z(n14188) );
  XNOR U18398 ( .A(n14184), .B(n14186), .Z(n18396) );
  XNOR U18399 ( .A(q[8]), .B(DB[593]), .Z(n14186) );
  XNOR U18400 ( .A(q[11]), .B(DB[596]), .Z(n14184) );
  IV U18401 ( .A(n14183), .Z(n18395) );
  XNOR U18402 ( .A(n14181), .B(n18397), .Z(n14183) );
  XNOR U18403 ( .A(q[10]), .B(DB[595]), .Z(n18397) );
  XNOR U18404 ( .A(q[9]), .B(DB[594]), .Z(n14181) );
  IV U18405 ( .A(n14196), .Z(n18391) );
  XOR U18406 ( .A(n18398), .B(n18399), .Z(n14196) );
  XNOR U18407 ( .A(n14213), .B(n14194), .Z(n18399) );
  XNOR U18408 ( .A(q[0]), .B(DB[585]), .Z(n14194) );
  XOR U18409 ( .A(n18400), .B(n14202), .Z(n14213) );
  XNOR U18410 ( .A(q[7]), .B(DB[592]), .Z(n14202) );
  IV U18411 ( .A(n14201), .Z(n18400) );
  XNOR U18412 ( .A(n14199), .B(n18401), .Z(n14201) );
  XNOR U18413 ( .A(q[6]), .B(DB[591]), .Z(n18401) );
  XNOR U18414 ( .A(q[5]), .B(DB[590]), .Z(n14199) );
  IV U18415 ( .A(n14212), .Z(n18398) );
  XOR U18416 ( .A(n18402), .B(n18403), .Z(n14212) );
  XNOR U18417 ( .A(n14208), .B(n14210), .Z(n18403) );
  XNOR U18418 ( .A(q[1]), .B(DB[586]), .Z(n14210) );
  XNOR U18419 ( .A(q[4]), .B(DB[589]), .Z(n14208) );
  IV U18420 ( .A(n14207), .Z(n18402) );
  XNOR U18421 ( .A(n14205), .B(n18404), .Z(n14207) );
  XNOR U18422 ( .A(q[3]), .B(DB[588]), .Z(n18404) );
  XNOR U18423 ( .A(q[2]), .B(DB[587]), .Z(n14205) );
  XOR U18424 ( .A(n18405), .B(n14103), .Z(n14031) );
  XOR U18425 ( .A(n18406), .B(n14095), .Z(n14103) );
  XOR U18426 ( .A(n18407), .B(n14084), .Z(n14095) );
  XNOR U18427 ( .A(q[14]), .B(DB[614]), .Z(n14084) );
  IV U18428 ( .A(n14083), .Z(n18407) );
  XNOR U18429 ( .A(n14081), .B(n18408), .Z(n14083) );
  XNOR U18430 ( .A(q[13]), .B(DB[613]), .Z(n18408) );
  XNOR U18431 ( .A(q[12]), .B(DB[612]), .Z(n14081) );
  IV U18432 ( .A(n14094), .Z(n18406) );
  XOR U18433 ( .A(n18409), .B(n18410), .Z(n14094) );
  XNOR U18434 ( .A(n14090), .B(n14092), .Z(n18410) );
  XNOR U18435 ( .A(q[8]), .B(DB[608]), .Z(n14092) );
  XNOR U18436 ( .A(q[11]), .B(DB[611]), .Z(n14090) );
  IV U18437 ( .A(n14089), .Z(n18409) );
  XNOR U18438 ( .A(n14087), .B(n18411), .Z(n14089) );
  XNOR U18439 ( .A(q[10]), .B(DB[610]), .Z(n18411) );
  XNOR U18440 ( .A(q[9]), .B(DB[609]), .Z(n14087) );
  IV U18441 ( .A(n14102), .Z(n18405) );
  XOR U18442 ( .A(n18412), .B(n18413), .Z(n14102) );
  XNOR U18443 ( .A(n14119), .B(n14100), .Z(n18413) );
  XNOR U18444 ( .A(q[0]), .B(DB[600]), .Z(n14100) );
  XOR U18445 ( .A(n18414), .B(n14108), .Z(n14119) );
  XNOR U18446 ( .A(q[7]), .B(DB[607]), .Z(n14108) );
  IV U18447 ( .A(n14107), .Z(n18414) );
  XNOR U18448 ( .A(n14105), .B(n18415), .Z(n14107) );
  XNOR U18449 ( .A(q[6]), .B(DB[606]), .Z(n18415) );
  XNOR U18450 ( .A(q[5]), .B(DB[605]), .Z(n14105) );
  IV U18451 ( .A(n14118), .Z(n18412) );
  XOR U18452 ( .A(n18416), .B(n18417), .Z(n14118) );
  XNOR U18453 ( .A(n14114), .B(n14116), .Z(n18417) );
  XNOR U18454 ( .A(q[1]), .B(DB[601]), .Z(n14116) );
  XNOR U18455 ( .A(q[4]), .B(DB[604]), .Z(n14114) );
  IV U18456 ( .A(n14113), .Z(n18416) );
  XNOR U18457 ( .A(n14111), .B(n18418), .Z(n14113) );
  XNOR U18458 ( .A(q[3]), .B(DB[603]), .Z(n18418) );
  XNOR U18459 ( .A(q[2]), .B(DB[602]), .Z(n14111) );
  XOR U18460 ( .A(n18419), .B(n14009), .Z(n13937) );
  XOR U18461 ( .A(n18420), .B(n14001), .Z(n14009) );
  XOR U18462 ( .A(n18421), .B(n13990), .Z(n14001) );
  XNOR U18463 ( .A(q[14]), .B(DB[629]), .Z(n13990) );
  IV U18464 ( .A(n13989), .Z(n18421) );
  XNOR U18465 ( .A(n13987), .B(n18422), .Z(n13989) );
  XNOR U18466 ( .A(q[13]), .B(DB[628]), .Z(n18422) );
  XNOR U18467 ( .A(q[12]), .B(DB[627]), .Z(n13987) );
  IV U18468 ( .A(n14000), .Z(n18420) );
  XOR U18469 ( .A(n18423), .B(n18424), .Z(n14000) );
  XNOR U18470 ( .A(n13996), .B(n13998), .Z(n18424) );
  XNOR U18471 ( .A(q[8]), .B(DB[623]), .Z(n13998) );
  XNOR U18472 ( .A(q[11]), .B(DB[626]), .Z(n13996) );
  IV U18473 ( .A(n13995), .Z(n18423) );
  XNOR U18474 ( .A(n13993), .B(n18425), .Z(n13995) );
  XNOR U18475 ( .A(q[10]), .B(DB[625]), .Z(n18425) );
  XNOR U18476 ( .A(q[9]), .B(DB[624]), .Z(n13993) );
  IV U18477 ( .A(n14008), .Z(n18419) );
  XOR U18478 ( .A(n18426), .B(n18427), .Z(n14008) );
  XNOR U18479 ( .A(n14025), .B(n14006), .Z(n18427) );
  XNOR U18480 ( .A(q[0]), .B(DB[615]), .Z(n14006) );
  XOR U18481 ( .A(n18428), .B(n14014), .Z(n14025) );
  XNOR U18482 ( .A(q[7]), .B(DB[622]), .Z(n14014) );
  IV U18483 ( .A(n14013), .Z(n18428) );
  XNOR U18484 ( .A(n14011), .B(n18429), .Z(n14013) );
  XNOR U18485 ( .A(q[6]), .B(DB[621]), .Z(n18429) );
  XNOR U18486 ( .A(q[5]), .B(DB[620]), .Z(n14011) );
  IV U18487 ( .A(n14024), .Z(n18426) );
  XOR U18488 ( .A(n18430), .B(n18431), .Z(n14024) );
  XNOR U18489 ( .A(n14020), .B(n14022), .Z(n18431) );
  XNOR U18490 ( .A(q[1]), .B(DB[616]), .Z(n14022) );
  XNOR U18491 ( .A(q[4]), .B(DB[619]), .Z(n14020) );
  IV U18492 ( .A(n14019), .Z(n18430) );
  XNOR U18493 ( .A(n14017), .B(n18432), .Z(n14019) );
  XNOR U18494 ( .A(q[3]), .B(DB[618]), .Z(n18432) );
  XNOR U18495 ( .A(q[2]), .B(DB[617]), .Z(n14017) );
  XOR U18496 ( .A(n18433), .B(n13915), .Z(n13843) );
  XOR U18497 ( .A(n18434), .B(n13907), .Z(n13915) );
  XOR U18498 ( .A(n18435), .B(n13896), .Z(n13907) );
  XNOR U18499 ( .A(q[14]), .B(DB[644]), .Z(n13896) );
  IV U18500 ( .A(n13895), .Z(n18435) );
  XNOR U18501 ( .A(n13893), .B(n18436), .Z(n13895) );
  XNOR U18502 ( .A(q[13]), .B(DB[643]), .Z(n18436) );
  XNOR U18503 ( .A(q[12]), .B(DB[642]), .Z(n13893) );
  IV U18504 ( .A(n13906), .Z(n18434) );
  XOR U18505 ( .A(n18437), .B(n18438), .Z(n13906) );
  XNOR U18506 ( .A(n13902), .B(n13904), .Z(n18438) );
  XNOR U18507 ( .A(q[8]), .B(DB[638]), .Z(n13904) );
  XNOR U18508 ( .A(q[11]), .B(DB[641]), .Z(n13902) );
  IV U18509 ( .A(n13901), .Z(n18437) );
  XNOR U18510 ( .A(n13899), .B(n18439), .Z(n13901) );
  XNOR U18511 ( .A(q[10]), .B(DB[640]), .Z(n18439) );
  XNOR U18512 ( .A(q[9]), .B(DB[639]), .Z(n13899) );
  IV U18513 ( .A(n13914), .Z(n18433) );
  XOR U18514 ( .A(n18440), .B(n18441), .Z(n13914) );
  XNOR U18515 ( .A(n13931), .B(n13912), .Z(n18441) );
  XNOR U18516 ( .A(q[0]), .B(DB[630]), .Z(n13912) );
  XOR U18517 ( .A(n18442), .B(n13920), .Z(n13931) );
  XNOR U18518 ( .A(q[7]), .B(DB[637]), .Z(n13920) );
  IV U18519 ( .A(n13919), .Z(n18442) );
  XNOR U18520 ( .A(n13917), .B(n18443), .Z(n13919) );
  XNOR U18521 ( .A(q[6]), .B(DB[636]), .Z(n18443) );
  XNOR U18522 ( .A(q[5]), .B(DB[635]), .Z(n13917) );
  IV U18523 ( .A(n13930), .Z(n18440) );
  XOR U18524 ( .A(n18444), .B(n18445), .Z(n13930) );
  XNOR U18525 ( .A(n13926), .B(n13928), .Z(n18445) );
  XNOR U18526 ( .A(q[1]), .B(DB[631]), .Z(n13928) );
  XNOR U18527 ( .A(q[4]), .B(DB[634]), .Z(n13926) );
  IV U18528 ( .A(n13925), .Z(n18444) );
  XNOR U18529 ( .A(n13923), .B(n18446), .Z(n13925) );
  XNOR U18530 ( .A(q[3]), .B(DB[633]), .Z(n18446) );
  XNOR U18531 ( .A(q[2]), .B(DB[632]), .Z(n13923) );
  XOR U18532 ( .A(n18447), .B(n13821), .Z(n13749) );
  XOR U18533 ( .A(n18448), .B(n13813), .Z(n13821) );
  XOR U18534 ( .A(n18449), .B(n13802), .Z(n13813) );
  XNOR U18535 ( .A(q[14]), .B(DB[659]), .Z(n13802) );
  IV U18536 ( .A(n13801), .Z(n18449) );
  XNOR U18537 ( .A(n13799), .B(n18450), .Z(n13801) );
  XNOR U18538 ( .A(q[13]), .B(DB[658]), .Z(n18450) );
  XNOR U18539 ( .A(q[12]), .B(DB[657]), .Z(n13799) );
  IV U18540 ( .A(n13812), .Z(n18448) );
  XOR U18541 ( .A(n18451), .B(n18452), .Z(n13812) );
  XNOR U18542 ( .A(n13808), .B(n13810), .Z(n18452) );
  XNOR U18543 ( .A(q[8]), .B(DB[653]), .Z(n13810) );
  XNOR U18544 ( .A(q[11]), .B(DB[656]), .Z(n13808) );
  IV U18545 ( .A(n13807), .Z(n18451) );
  XNOR U18546 ( .A(n13805), .B(n18453), .Z(n13807) );
  XNOR U18547 ( .A(q[10]), .B(DB[655]), .Z(n18453) );
  XNOR U18548 ( .A(q[9]), .B(DB[654]), .Z(n13805) );
  IV U18549 ( .A(n13820), .Z(n18447) );
  XOR U18550 ( .A(n18454), .B(n18455), .Z(n13820) );
  XNOR U18551 ( .A(n13837), .B(n13818), .Z(n18455) );
  XNOR U18552 ( .A(q[0]), .B(DB[645]), .Z(n13818) );
  XOR U18553 ( .A(n18456), .B(n13826), .Z(n13837) );
  XNOR U18554 ( .A(q[7]), .B(DB[652]), .Z(n13826) );
  IV U18555 ( .A(n13825), .Z(n18456) );
  XNOR U18556 ( .A(n13823), .B(n18457), .Z(n13825) );
  XNOR U18557 ( .A(q[6]), .B(DB[651]), .Z(n18457) );
  XNOR U18558 ( .A(q[5]), .B(DB[650]), .Z(n13823) );
  IV U18559 ( .A(n13836), .Z(n18454) );
  XOR U18560 ( .A(n18458), .B(n18459), .Z(n13836) );
  XNOR U18561 ( .A(n13832), .B(n13834), .Z(n18459) );
  XNOR U18562 ( .A(q[1]), .B(DB[646]), .Z(n13834) );
  XNOR U18563 ( .A(q[4]), .B(DB[649]), .Z(n13832) );
  IV U18564 ( .A(n13831), .Z(n18458) );
  XNOR U18565 ( .A(n13829), .B(n18460), .Z(n13831) );
  XNOR U18566 ( .A(q[3]), .B(DB[648]), .Z(n18460) );
  XNOR U18567 ( .A(q[2]), .B(DB[647]), .Z(n13829) );
  XOR U18568 ( .A(n18461), .B(n13727), .Z(n13655) );
  XOR U18569 ( .A(n18462), .B(n13719), .Z(n13727) );
  XOR U18570 ( .A(n18463), .B(n13708), .Z(n13719) );
  XNOR U18571 ( .A(q[14]), .B(DB[674]), .Z(n13708) );
  IV U18572 ( .A(n13707), .Z(n18463) );
  XNOR U18573 ( .A(n13705), .B(n18464), .Z(n13707) );
  XNOR U18574 ( .A(q[13]), .B(DB[673]), .Z(n18464) );
  XNOR U18575 ( .A(q[12]), .B(DB[672]), .Z(n13705) );
  IV U18576 ( .A(n13718), .Z(n18462) );
  XOR U18577 ( .A(n18465), .B(n18466), .Z(n13718) );
  XNOR U18578 ( .A(n13714), .B(n13716), .Z(n18466) );
  XNOR U18579 ( .A(q[8]), .B(DB[668]), .Z(n13716) );
  XNOR U18580 ( .A(q[11]), .B(DB[671]), .Z(n13714) );
  IV U18581 ( .A(n13713), .Z(n18465) );
  XNOR U18582 ( .A(n13711), .B(n18467), .Z(n13713) );
  XNOR U18583 ( .A(q[10]), .B(DB[670]), .Z(n18467) );
  XNOR U18584 ( .A(q[9]), .B(DB[669]), .Z(n13711) );
  IV U18585 ( .A(n13726), .Z(n18461) );
  XOR U18586 ( .A(n18468), .B(n18469), .Z(n13726) );
  XNOR U18587 ( .A(n13743), .B(n13724), .Z(n18469) );
  XNOR U18588 ( .A(q[0]), .B(DB[660]), .Z(n13724) );
  XOR U18589 ( .A(n18470), .B(n13732), .Z(n13743) );
  XNOR U18590 ( .A(q[7]), .B(DB[667]), .Z(n13732) );
  IV U18591 ( .A(n13731), .Z(n18470) );
  XNOR U18592 ( .A(n13729), .B(n18471), .Z(n13731) );
  XNOR U18593 ( .A(q[6]), .B(DB[666]), .Z(n18471) );
  XNOR U18594 ( .A(q[5]), .B(DB[665]), .Z(n13729) );
  IV U18595 ( .A(n13742), .Z(n18468) );
  XOR U18596 ( .A(n18472), .B(n18473), .Z(n13742) );
  XNOR U18597 ( .A(n13738), .B(n13740), .Z(n18473) );
  XNOR U18598 ( .A(q[1]), .B(DB[661]), .Z(n13740) );
  XNOR U18599 ( .A(q[4]), .B(DB[664]), .Z(n13738) );
  IV U18600 ( .A(n13737), .Z(n18472) );
  XNOR U18601 ( .A(n13735), .B(n18474), .Z(n13737) );
  XNOR U18602 ( .A(q[3]), .B(DB[663]), .Z(n18474) );
  XNOR U18603 ( .A(q[2]), .B(DB[662]), .Z(n13735) );
  XOR U18604 ( .A(n18475), .B(n13633), .Z(n13561) );
  XOR U18605 ( .A(n18476), .B(n13625), .Z(n13633) );
  XOR U18606 ( .A(n18477), .B(n13614), .Z(n13625) );
  XNOR U18607 ( .A(q[14]), .B(DB[689]), .Z(n13614) );
  IV U18608 ( .A(n13613), .Z(n18477) );
  XNOR U18609 ( .A(n13611), .B(n18478), .Z(n13613) );
  XNOR U18610 ( .A(q[13]), .B(DB[688]), .Z(n18478) );
  XNOR U18611 ( .A(q[12]), .B(DB[687]), .Z(n13611) );
  IV U18612 ( .A(n13624), .Z(n18476) );
  XOR U18613 ( .A(n18479), .B(n18480), .Z(n13624) );
  XNOR U18614 ( .A(n13620), .B(n13622), .Z(n18480) );
  XNOR U18615 ( .A(q[8]), .B(DB[683]), .Z(n13622) );
  XNOR U18616 ( .A(q[11]), .B(DB[686]), .Z(n13620) );
  IV U18617 ( .A(n13619), .Z(n18479) );
  XNOR U18618 ( .A(n13617), .B(n18481), .Z(n13619) );
  XNOR U18619 ( .A(q[10]), .B(DB[685]), .Z(n18481) );
  XNOR U18620 ( .A(q[9]), .B(DB[684]), .Z(n13617) );
  IV U18621 ( .A(n13632), .Z(n18475) );
  XOR U18622 ( .A(n18482), .B(n18483), .Z(n13632) );
  XNOR U18623 ( .A(n13649), .B(n13630), .Z(n18483) );
  XNOR U18624 ( .A(q[0]), .B(DB[675]), .Z(n13630) );
  XOR U18625 ( .A(n18484), .B(n13638), .Z(n13649) );
  XNOR U18626 ( .A(q[7]), .B(DB[682]), .Z(n13638) );
  IV U18627 ( .A(n13637), .Z(n18484) );
  XNOR U18628 ( .A(n13635), .B(n18485), .Z(n13637) );
  XNOR U18629 ( .A(q[6]), .B(DB[681]), .Z(n18485) );
  XNOR U18630 ( .A(q[5]), .B(DB[680]), .Z(n13635) );
  IV U18631 ( .A(n13648), .Z(n18482) );
  XOR U18632 ( .A(n18486), .B(n18487), .Z(n13648) );
  XNOR U18633 ( .A(n13644), .B(n13646), .Z(n18487) );
  XNOR U18634 ( .A(q[1]), .B(DB[676]), .Z(n13646) );
  XNOR U18635 ( .A(q[4]), .B(DB[679]), .Z(n13644) );
  IV U18636 ( .A(n13643), .Z(n18486) );
  XNOR U18637 ( .A(n13641), .B(n18488), .Z(n13643) );
  XNOR U18638 ( .A(q[3]), .B(DB[678]), .Z(n18488) );
  XNOR U18639 ( .A(q[2]), .B(DB[677]), .Z(n13641) );
  XOR U18640 ( .A(n18489), .B(n13539), .Z(n13467) );
  XOR U18641 ( .A(n18490), .B(n13531), .Z(n13539) );
  XOR U18642 ( .A(n18491), .B(n13520), .Z(n13531) );
  XNOR U18643 ( .A(q[14]), .B(DB[704]), .Z(n13520) );
  IV U18644 ( .A(n13519), .Z(n18491) );
  XNOR U18645 ( .A(n13517), .B(n18492), .Z(n13519) );
  XNOR U18646 ( .A(q[13]), .B(DB[703]), .Z(n18492) );
  XNOR U18647 ( .A(q[12]), .B(DB[702]), .Z(n13517) );
  IV U18648 ( .A(n13530), .Z(n18490) );
  XOR U18649 ( .A(n18493), .B(n18494), .Z(n13530) );
  XNOR U18650 ( .A(n13526), .B(n13528), .Z(n18494) );
  XNOR U18651 ( .A(q[8]), .B(DB[698]), .Z(n13528) );
  XNOR U18652 ( .A(q[11]), .B(DB[701]), .Z(n13526) );
  IV U18653 ( .A(n13525), .Z(n18493) );
  XNOR U18654 ( .A(n13523), .B(n18495), .Z(n13525) );
  XNOR U18655 ( .A(q[10]), .B(DB[700]), .Z(n18495) );
  XNOR U18656 ( .A(q[9]), .B(DB[699]), .Z(n13523) );
  IV U18657 ( .A(n13538), .Z(n18489) );
  XOR U18658 ( .A(n18496), .B(n18497), .Z(n13538) );
  XNOR U18659 ( .A(n13555), .B(n13536), .Z(n18497) );
  XNOR U18660 ( .A(q[0]), .B(DB[690]), .Z(n13536) );
  XOR U18661 ( .A(n18498), .B(n13544), .Z(n13555) );
  XNOR U18662 ( .A(q[7]), .B(DB[697]), .Z(n13544) );
  IV U18663 ( .A(n13543), .Z(n18498) );
  XNOR U18664 ( .A(n13541), .B(n18499), .Z(n13543) );
  XNOR U18665 ( .A(q[6]), .B(DB[696]), .Z(n18499) );
  XNOR U18666 ( .A(q[5]), .B(DB[695]), .Z(n13541) );
  IV U18667 ( .A(n13554), .Z(n18496) );
  XOR U18668 ( .A(n18500), .B(n18501), .Z(n13554) );
  XNOR U18669 ( .A(n13550), .B(n13552), .Z(n18501) );
  XNOR U18670 ( .A(q[1]), .B(DB[691]), .Z(n13552) );
  XNOR U18671 ( .A(q[4]), .B(DB[694]), .Z(n13550) );
  IV U18672 ( .A(n13549), .Z(n18500) );
  XNOR U18673 ( .A(n13547), .B(n18502), .Z(n13549) );
  XNOR U18674 ( .A(q[3]), .B(DB[693]), .Z(n18502) );
  XNOR U18675 ( .A(q[2]), .B(DB[692]), .Z(n13547) );
  XOR U18676 ( .A(n18503), .B(n13445), .Z(n13373) );
  XOR U18677 ( .A(n18504), .B(n13437), .Z(n13445) );
  XOR U18678 ( .A(n18505), .B(n13426), .Z(n13437) );
  XNOR U18679 ( .A(q[14]), .B(DB[719]), .Z(n13426) );
  IV U18680 ( .A(n13425), .Z(n18505) );
  XNOR U18681 ( .A(n13423), .B(n18506), .Z(n13425) );
  XNOR U18682 ( .A(q[13]), .B(DB[718]), .Z(n18506) );
  XNOR U18683 ( .A(q[12]), .B(DB[717]), .Z(n13423) );
  IV U18684 ( .A(n13436), .Z(n18504) );
  XOR U18685 ( .A(n18507), .B(n18508), .Z(n13436) );
  XNOR U18686 ( .A(n13432), .B(n13434), .Z(n18508) );
  XNOR U18687 ( .A(q[8]), .B(DB[713]), .Z(n13434) );
  XNOR U18688 ( .A(q[11]), .B(DB[716]), .Z(n13432) );
  IV U18689 ( .A(n13431), .Z(n18507) );
  XNOR U18690 ( .A(n13429), .B(n18509), .Z(n13431) );
  XNOR U18691 ( .A(q[10]), .B(DB[715]), .Z(n18509) );
  XNOR U18692 ( .A(q[9]), .B(DB[714]), .Z(n13429) );
  IV U18693 ( .A(n13444), .Z(n18503) );
  XOR U18694 ( .A(n18510), .B(n18511), .Z(n13444) );
  XNOR U18695 ( .A(n13461), .B(n13442), .Z(n18511) );
  XNOR U18696 ( .A(q[0]), .B(DB[705]), .Z(n13442) );
  XOR U18697 ( .A(n18512), .B(n13450), .Z(n13461) );
  XNOR U18698 ( .A(q[7]), .B(DB[712]), .Z(n13450) );
  IV U18699 ( .A(n13449), .Z(n18512) );
  XNOR U18700 ( .A(n13447), .B(n18513), .Z(n13449) );
  XNOR U18701 ( .A(q[6]), .B(DB[711]), .Z(n18513) );
  XNOR U18702 ( .A(q[5]), .B(DB[710]), .Z(n13447) );
  IV U18703 ( .A(n13460), .Z(n18510) );
  XOR U18704 ( .A(n18514), .B(n18515), .Z(n13460) );
  XNOR U18705 ( .A(n13456), .B(n13458), .Z(n18515) );
  XNOR U18706 ( .A(q[1]), .B(DB[706]), .Z(n13458) );
  XNOR U18707 ( .A(q[4]), .B(DB[709]), .Z(n13456) );
  IV U18708 ( .A(n13455), .Z(n18514) );
  XNOR U18709 ( .A(n13453), .B(n18516), .Z(n13455) );
  XNOR U18710 ( .A(q[3]), .B(DB[708]), .Z(n18516) );
  XNOR U18711 ( .A(q[2]), .B(DB[707]), .Z(n13453) );
  XOR U18712 ( .A(n18517), .B(n13351), .Z(n13279) );
  XOR U18713 ( .A(n18518), .B(n13343), .Z(n13351) );
  XOR U18714 ( .A(n18519), .B(n13332), .Z(n13343) );
  XNOR U18715 ( .A(q[14]), .B(DB[734]), .Z(n13332) );
  IV U18716 ( .A(n13331), .Z(n18519) );
  XNOR U18717 ( .A(n13329), .B(n18520), .Z(n13331) );
  XNOR U18718 ( .A(q[13]), .B(DB[733]), .Z(n18520) );
  XNOR U18719 ( .A(q[12]), .B(DB[732]), .Z(n13329) );
  IV U18720 ( .A(n13342), .Z(n18518) );
  XOR U18721 ( .A(n18521), .B(n18522), .Z(n13342) );
  XNOR U18722 ( .A(n13338), .B(n13340), .Z(n18522) );
  XNOR U18723 ( .A(q[8]), .B(DB[728]), .Z(n13340) );
  XNOR U18724 ( .A(q[11]), .B(DB[731]), .Z(n13338) );
  IV U18725 ( .A(n13337), .Z(n18521) );
  XNOR U18726 ( .A(n13335), .B(n18523), .Z(n13337) );
  XNOR U18727 ( .A(q[10]), .B(DB[730]), .Z(n18523) );
  XNOR U18728 ( .A(q[9]), .B(DB[729]), .Z(n13335) );
  IV U18729 ( .A(n13350), .Z(n18517) );
  XOR U18730 ( .A(n18524), .B(n18525), .Z(n13350) );
  XNOR U18731 ( .A(n13367), .B(n13348), .Z(n18525) );
  XNOR U18732 ( .A(q[0]), .B(DB[720]), .Z(n13348) );
  XOR U18733 ( .A(n18526), .B(n13356), .Z(n13367) );
  XNOR U18734 ( .A(q[7]), .B(DB[727]), .Z(n13356) );
  IV U18735 ( .A(n13355), .Z(n18526) );
  XNOR U18736 ( .A(n13353), .B(n18527), .Z(n13355) );
  XNOR U18737 ( .A(q[6]), .B(DB[726]), .Z(n18527) );
  XNOR U18738 ( .A(q[5]), .B(DB[725]), .Z(n13353) );
  IV U18739 ( .A(n13366), .Z(n18524) );
  XOR U18740 ( .A(n18528), .B(n18529), .Z(n13366) );
  XNOR U18741 ( .A(n13362), .B(n13364), .Z(n18529) );
  XNOR U18742 ( .A(q[1]), .B(DB[721]), .Z(n13364) );
  XNOR U18743 ( .A(q[4]), .B(DB[724]), .Z(n13362) );
  IV U18744 ( .A(n13361), .Z(n18528) );
  XNOR U18745 ( .A(n13359), .B(n18530), .Z(n13361) );
  XNOR U18746 ( .A(q[3]), .B(DB[723]), .Z(n18530) );
  XNOR U18747 ( .A(q[2]), .B(DB[722]), .Z(n13359) );
  XOR U18748 ( .A(n18531), .B(n13257), .Z(n13185) );
  XOR U18749 ( .A(n18532), .B(n13249), .Z(n13257) );
  XOR U18750 ( .A(n18533), .B(n13238), .Z(n13249) );
  XNOR U18751 ( .A(q[14]), .B(DB[749]), .Z(n13238) );
  IV U18752 ( .A(n13237), .Z(n18533) );
  XNOR U18753 ( .A(n13235), .B(n18534), .Z(n13237) );
  XNOR U18754 ( .A(q[13]), .B(DB[748]), .Z(n18534) );
  XNOR U18755 ( .A(q[12]), .B(DB[747]), .Z(n13235) );
  IV U18756 ( .A(n13248), .Z(n18532) );
  XOR U18757 ( .A(n18535), .B(n18536), .Z(n13248) );
  XNOR U18758 ( .A(n13244), .B(n13246), .Z(n18536) );
  XNOR U18759 ( .A(q[8]), .B(DB[743]), .Z(n13246) );
  XNOR U18760 ( .A(q[11]), .B(DB[746]), .Z(n13244) );
  IV U18761 ( .A(n13243), .Z(n18535) );
  XNOR U18762 ( .A(n13241), .B(n18537), .Z(n13243) );
  XNOR U18763 ( .A(q[10]), .B(DB[745]), .Z(n18537) );
  XNOR U18764 ( .A(q[9]), .B(DB[744]), .Z(n13241) );
  IV U18765 ( .A(n13256), .Z(n18531) );
  XOR U18766 ( .A(n18538), .B(n18539), .Z(n13256) );
  XNOR U18767 ( .A(n13273), .B(n13254), .Z(n18539) );
  XNOR U18768 ( .A(q[0]), .B(DB[735]), .Z(n13254) );
  XOR U18769 ( .A(n18540), .B(n13262), .Z(n13273) );
  XNOR U18770 ( .A(q[7]), .B(DB[742]), .Z(n13262) );
  IV U18771 ( .A(n13261), .Z(n18540) );
  XNOR U18772 ( .A(n13259), .B(n18541), .Z(n13261) );
  XNOR U18773 ( .A(q[6]), .B(DB[741]), .Z(n18541) );
  XNOR U18774 ( .A(q[5]), .B(DB[740]), .Z(n13259) );
  IV U18775 ( .A(n13272), .Z(n18538) );
  XOR U18776 ( .A(n18542), .B(n18543), .Z(n13272) );
  XNOR U18777 ( .A(n13268), .B(n13270), .Z(n18543) );
  XNOR U18778 ( .A(q[1]), .B(DB[736]), .Z(n13270) );
  XNOR U18779 ( .A(q[4]), .B(DB[739]), .Z(n13268) );
  IV U18780 ( .A(n13267), .Z(n18542) );
  XNOR U18781 ( .A(n13265), .B(n18544), .Z(n13267) );
  XNOR U18782 ( .A(q[3]), .B(DB[738]), .Z(n18544) );
  XNOR U18783 ( .A(q[2]), .B(DB[737]), .Z(n13265) );
  XOR U18784 ( .A(n18545), .B(n13163), .Z(n13091) );
  XOR U18785 ( .A(n18546), .B(n13155), .Z(n13163) );
  XOR U18786 ( .A(n18547), .B(n13144), .Z(n13155) );
  XNOR U18787 ( .A(q[14]), .B(DB[764]), .Z(n13144) );
  IV U18788 ( .A(n13143), .Z(n18547) );
  XNOR U18789 ( .A(n13141), .B(n18548), .Z(n13143) );
  XNOR U18790 ( .A(q[13]), .B(DB[763]), .Z(n18548) );
  XNOR U18791 ( .A(q[12]), .B(DB[762]), .Z(n13141) );
  IV U18792 ( .A(n13154), .Z(n18546) );
  XOR U18793 ( .A(n18549), .B(n18550), .Z(n13154) );
  XNOR U18794 ( .A(n13150), .B(n13152), .Z(n18550) );
  XNOR U18795 ( .A(q[8]), .B(DB[758]), .Z(n13152) );
  XNOR U18796 ( .A(q[11]), .B(DB[761]), .Z(n13150) );
  IV U18797 ( .A(n13149), .Z(n18549) );
  XNOR U18798 ( .A(n13147), .B(n18551), .Z(n13149) );
  XNOR U18799 ( .A(q[10]), .B(DB[760]), .Z(n18551) );
  XNOR U18800 ( .A(q[9]), .B(DB[759]), .Z(n13147) );
  IV U18801 ( .A(n13162), .Z(n18545) );
  XOR U18802 ( .A(n18552), .B(n18553), .Z(n13162) );
  XNOR U18803 ( .A(n13179), .B(n13160), .Z(n18553) );
  XNOR U18804 ( .A(q[0]), .B(DB[750]), .Z(n13160) );
  XOR U18805 ( .A(n18554), .B(n13168), .Z(n13179) );
  XNOR U18806 ( .A(q[7]), .B(DB[757]), .Z(n13168) );
  IV U18807 ( .A(n13167), .Z(n18554) );
  XNOR U18808 ( .A(n13165), .B(n18555), .Z(n13167) );
  XNOR U18809 ( .A(q[6]), .B(DB[756]), .Z(n18555) );
  XNOR U18810 ( .A(q[5]), .B(DB[755]), .Z(n13165) );
  IV U18811 ( .A(n13178), .Z(n18552) );
  XOR U18812 ( .A(n18556), .B(n18557), .Z(n13178) );
  XNOR U18813 ( .A(n13174), .B(n13176), .Z(n18557) );
  XNOR U18814 ( .A(q[1]), .B(DB[751]), .Z(n13176) );
  XNOR U18815 ( .A(q[4]), .B(DB[754]), .Z(n13174) );
  IV U18816 ( .A(n13173), .Z(n18556) );
  XNOR U18817 ( .A(n13171), .B(n18558), .Z(n13173) );
  XNOR U18818 ( .A(q[3]), .B(DB[753]), .Z(n18558) );
  XNOR U18819 ( .A(q[2]), .B(DB[752]), .Z(n13171) );
  XOR U18820 ( .A(n18559), .B(n13069), .Z(n12997) );
  XOR U18821 ( .A(n18560), .B(n13061), .Z(n13069) );
  XOR U18822 ( .A(n18561), .B(n13050), .Z(n13061) );
  XNOR U18823 ( .A(q[14]), .B(DB[779]), .Z(n13050) );
  IV U18824 ( .A(n13049), .Z(n18561) );
  XNOR U18825 ( .A(n13047), .B(n18562), .Z(n13049) );
  XNOR U18826 ( .A(q[13]), .B(DB[778]), .Z(n18562) );
  XNOR U18827 ( .A(q[12]), .B(DB[777]), .Z(n13047) );
  IV U18828 ( .A(n13060), .Z(n18560) );
  XOR U18829 ( .A(n18563), .B(n18564), .Z(n13060) );
  XNOR U18830 ( .A(n13056), .B(n13058), .Z(n18564) );
  XNOR U18831 ( .A(q[8]), .B(DB[773]), .Z(n13058) );
  XNOR U18832 ( .A(q[11]), .B(DB[776]), .Z(n13056) );
  IV U18833 ( .A(n13055), .Z(n18563) );
  XNOR U18834 ( .A(n13053), .B(n18565), .Z(n13055) );
  XNOR U18835 ( .A(q[10]), .B(DB[775]), .Z(n18565) );
  XNOR U18836 ( .A(q[9]), .B(DB[774]), .Z(n13053) );
  IV U18837 ( .A(n13068), .Z(n18559) );
  XOR U18838 ( .A(n18566), .B(n18567), .Z(n13068) );
  XNOR U18839 ( .A(n13085), .B(n13066), .Z(n18567) );
  XNOR U18840 ( .A(q[0]), .B(DB[765]), .Z(n13066) );
  XOR U18841 ( .A(n18568), .B(n13074), .Z(n13085) );
  XNOR U18842 ( .A(q[7]), .B(DB[772]), .Z(n13074) );
  IV U18843 ( .A(n13073), .Z(n18568) );
  XNOR U18844 ( .A(n13071), .B(n18569), .Z(n13073) );
  XNOR U18845 ( .A(q[6]), .B(DB[771]), .Z(n18569) );
  XNOR U18846 ( .A(q[5]), .B(DB[770]), .Z(n13071) );
  IV U18847 ( .A(n13084), .Z(n18566) );
  XOR U18848 ( .A(n18570), .B(n18571), .Z(n13084) );
  XNOR U18849 ( .A(n13080), .B(n13082), .Z(n18571) );
  XNOR U18850 ( .A(q[1]), .B(DB[766]), .Z(n13082) );
  XNOR U18851 ( .A(q[4]), .B(DB[769]), .Z(n13080) );
  IV U18852 ( .A(n13079), .Z(n18570) );
  XNOR U18853 ( .A(n13077), .B(n18572), .Z(n13079) );
  XNOR U18854 ( .A(q[3]), .B(DB[768]), .Z(n18572) );
  XNOR U18855 ( .A(q[2]), .B(DB[767]), .Z(n13077) );
  XOR U18856 ( .A(n18573), .B(n12975), .Z(n12903) );
  XOR U18857 ( .A(n18574), .B(n12967), .Z(n12975) );
  XOR U18858 ( .A(n18575), .B(n12956), .Z(n12967) );
  XNOR U18859 ( .A(q[14]), .B(DB[794]), .Z(n12956) );
  IV U18860 ( .A(n12955), .Z(n18575) );
  XNOR U18861 ( .A(n12953), .B(n18576), .Z(n12955) );
  XNOR U18862 ( .A(q[13]), .B(DB[793]), .Z(n18576) );
  XNOR U18863 ( .A(q[12]), .B(DB[792]), .Z(n12953) );
  IV U18864 ( .A(n12966), .Z(n18574) );
  XOR U18865 ( .A(n18577), .B(n18578), .Z(n12966) );
  XNOR U18866 ( .A(n12962), .B(n12964), .Z(n18578) );
  XNOR U18867 ( .A(q[8]), .B(DB[788]), .Z(n12964) );
  XNOR U18868 ( .A(q[11]), .B(DB[791]), .Z(n12962) );
  IV U18869 ( .A(n12961), .Z(n18577) );
  XNOR U18870 ( .A(n12959), .B(n18579), .Z(n12961) );
  XNOR U18871 ( .A(q[10]), .B(DB[790]), .Z(n18579) );
  XNOR U18872 ( .A(q[9]), .B(DB[789]), .Z(n12959) );
  IV U18873 ( .A(n12974), .Z(n18573) );
  XOR U18874 ( .A(n18580), .B(n18581), .Z(n12974) );
  XNOR U18875 ( .A(n12991), .B(n12972), .Z(n18581) );
  XNOR U18876 ( .A(q[0]), .B(DB[780]), .Z(n12972) );
  XOR U18877 ( .A(n18582), .B(n12980), .Z(n12991) );
  XNOR U18878 ( .A(q[7]), .B(DB[787]), .Z(n12980) );
  IV U18879 ( .A(n12979), .Z(n18582) );
  XNOR U18880 ( .A(n12977), .B(n18583), .Z(n12979) );
  XNOR U18881 ( .A(q[6]), .B(DB[786]), .Z(n18583) );
  XNOR U18882 ( .A(q[5]), .B(DB[785]), .Z(n12977) );
  IV U18883 ( .A(n12990), .Z(n18580) );
  XOR U18884 ( .A(n18584), .B(n18585), .Z(n12990) );
  XNOR U18885 ( .A(n12986), .B(n12988), .Z(n18585) );
  XNOR U18886 ( .A(q[1]), .B(DB[781]), .Z(n12988) );
  XNOR U18887 ( .A(q[4]), .B(DB[784]), .Z(n12986) );
  IV U18888 ( .A(n12985), .Z(n18584) );
  XNOR U18889 ( .A(n12983), .B(n18586), .Z(n12985) );
  XNOR U18890 ( .A(q[3]), .B(DB[783]), .Z(n18586) );
  XNOR U18891 ( .A(q[2]), .B(DB[782]), .Z(n12983) );
  XOR U18892 ( .A(n18587), .B(n12881), .Z(n12809) );
  XOR U18893 ( .A(n18588), .B(n12873), .Z(n12881) );
  XOR U18894 ( .A(n18589), .B(n12862), .Z(n12873) );
  XNOR U18895 ( .A(q[14]), .B(DB[809]), .Z(n12862) );
  IV U18896 ( .A(n12861), .Z(n18589) );
  XNOR U18897 ( .A(n12859), .B(n18590), .Z(n12861) );
  XNOR U18898 ( .A(q[13]), .B(DB[808]), .Z(n18590) );
  XNOR U18899 ( .A(q[12]), .B(DB[807]), .Z(n12859) );
  IV U18900 ( .A(n12872), .Z(n18588) );
  XOR U18901 ( .A(n18591), .B(n18592), .Z(n12872) );
  XNOR U18902 ( .A(n12868), .B(n12870), .Z(n18592) );
  XNOR U18903 ( .A(q[8]), .B(DB[803]), .Z(n12870) );
  XNOR U18904 ( .A(q[11]), .B(DB[806]), .Z(n12868) );
  IV U18905 ( .A(n12867), .Z(n18591) );
  XNOR U18906 ( .A(n12865), .B(n18593), .Z(n12867) );
  XNOR U18907 ( .A(q[10]), .B(DB[805]), .Z(n18593) );
  XNOR U18908 ( .A(q[9]), .B(DB[804]), .Z(n12865) );
  IV U18909 ( .A(n12880), .Z(n18587) );
  XOR U18910 ( .A(n18594), .B(n18595), .Z(n12880) );
  XNOR U18911 ( .A(n12897), .B(n12878), .Z(n18595) );
  XNOR U18912 ( .A(q[0]), .B(DB[795]), .Z(n12878) );
  XOR U18913 ( .A(n18596), .B(n12886), .Z(n12897) );
  XNOR U18914 ( .A(q[7]), .B(DB[802]), .Z(n12886) );
  IV U18915 ( .A(n12885), .Z(n18596) );
  XNOR U18916 ( .A(n12883), .B(n18597), .Z(n12885) );
  XNOR U18917 ( .A(q[6]), .B(DB[801]), .Z(n18597) );
  XNOR U18918 ( .A(q[5]), .B(DB[800]), .Z(n12883) );
  IV U18919 ( .A(n12896), .Z(n18594) );
  XOR U18920 ( .A(n18598), .B(n18599), .Z(n12896) );
  XNOR U18921 ( .A(n12892), .B(n12894), .Z(n18599) );
  XNOR U18922 ( .A(q[1]), .B(DB[796]), .Z(n12894) );
  XNOR U18923 ( .A(q[4]), .B(DB[799]), .Z(n12892) );
  IV U18924 ( .A(n12891), .Z(n18598) );
  XNOR U18925 ( .A(n12889), .B(n18600), .Z(n12891) );
  XNOR U18926 ( .A(q[3]), .B(DB[798]), .Z(n18600) );
  XNOR U18927 ( .A(q[2]), .B(DB[797]), .Z(n12889) );
  XOR U18928 ( .A(n18601), .B(n12787), .Z(n12715) );
  XOR U18929 ( .A(n18602), .B(n12779), .Z(n12787) );
  XOR U18930 ( .A(n18603), .B(n12768), .Z(n12779) );
  XNOR U18931 ( .A(q[14]), .B(DB[824]), .Z(n12768) );
  IV U18932 ( .A(n12767), .Z(n18603) );
  XNOR U18933 ( .A(n12765), .B(n18604), .Z(n12767) );
  XNOR U18934 ( .A(q[13]), .B(DB[823]), .Z(n18604) );
  XNOR U18935 ( .A(q[12]), .B(DB[822]), .Z(n12765) );
  IV U18936 ( .A(n12778), .Z(n18602) );
  XOR U18937 ( .A(n18605), .B(n18606), .Z(n12778) );
  XNOR U18938 ( .A(n12774), .B(n12776), .Z(n18606) );
  XNOR U18939 ( .A(q[8]), .B(DB[818]), .Z(n12776) );
  XNOR U18940 ( .A(q[11]), .B(DB[821]), .Z(n12774) );
  IV U18941 ( .A(n12773), .Z(n18605) );
  XNOR U18942 ( .A(n12771), .B(n18607), .Z(n12773) );
  XNOR U18943 ( .A(q[10]), .B(DB[820]), .Z(n18607) );
  XNOR U18944 ( .A(q[9]), .B(DB[819]), .Z(n12771) );
  IV U18945 ( .A(n12786), .Z(n18601) );
  XOR U18946 ( .A(n18608), .B(n18609), .Z(n12786) );
  XNOR U18947 ( .A(n12803), .B(n12784), .Z(n18609) );
  XNOR U18948 ( .A(q[0]), .B(DB[810]), .Z(n12784) );
  XOR U18949 ( .A(n18610), .B(n12792), .Z(n12803) );
  XNOR U18950 ( .A(q[7]), .B(DB[817]), .Z(n12792) );
  IV U18951 ( .A(n12791), .Z(n18610) );
  XNOR U18952 ( .A(n12789), .B(n18611), .Z(n12791) );
  XNOR U18953 ( .A(q[6]), .B(DB[816]), .Z(n18611) );
  XNOR U18954 ( .A(q[5]), .B(DB[815]), .Z(n12789) );
  IV U18955 ( .A(n12802), .Z(n18608) );
  XOR U18956 ( .A(n18612), .B(n18613), .Z(n12802) );
  XNOR U18957 ( .A(n12798), .B(n12800), .Z(n18613) );
  XNOR U18958 ( .A(q[1]), .B(DB[811]), .Z(n12800) );
  XNOR U18959 ( .A(q[4]), .B(DB[814]), .Z(n12798) );
  IV U18960 ( .A(n12797), .Z(n18612) );
  XNOR U18961 ( .A(n12795), .B(n18614), .Z(n12797) );
  XNOR U18962 ( .A(q[3]), .B(DB[813]), .Z(n18614) );
  XNOR U18963 ( .A(q[2]), .B(DB[812]), .Z(n12795) );
  XOR U18964 ( .A(n18615), .B(n12693), .Z(n12621) );
  XOR U18965 ( .A(n18616), .B(n12685), .Z(n12693) );
  XOR U18966 ( .A(n18617), .B(n12674), .Z(n12685) );
  XNOR U18967 ( .A(q[14]), .B(DB[839]), .Z(n12674) );
  IV U18968 ( .A(n12673), .Z(n18617) );
  XNOR U18969 ( .A(n12671), .B(n18618), .Z(n12673) );
  XNOR U18970 ( .A(q[13]), .B(DB[838]), .Z(n18618) );
  XNOR U18971 ( .A(q[12]), .B(DB[837]), .Z(n12671) );
  IV U18972 ( .A(n12684), .Z(n18616) );
  XOR U18973 ( .A(n18619), .B(n18620), .Z(n12684) );
  XNOR U18974 ( .A(n12680), .B(n12682), .Z(n18620) );
  XNOR U18975 ( .A(q[8]), .B(DB[833]), .Z(n12682) );
  XNOR U18976 ( .A(q[11]), .B(DB[836]), .Z(n12680) );
  IV U18977 ( .A(n12679), .Z(n18619) );
  XNOR U18978 ( .A(n12677), .B(n18621), .Z(n12679) );
  XNOR U18979 ( .A(q[10]), .B(DB[835]), .Z(n18621) );
  XNOR U18980 ( .A(q[9]), .B(DB[834]), .Z(n12677) );
  IV U18981 ( .A(n12692), .Z(n18615) );
  XOR U18982 ( .A(n18622), .B(n18623), .Z(n12692) );
  XNOR U18983 ( .A(n12709), .B(n12690), .Z(n18623) );
  XNOR U18984 ( .A(q[0]), .B(DB[825]), .Z(n12690) );
  XOR U18985 ( .A(n18624), .B(n12698), .Z(n12709) );
  XNOR U18986 ( .A(q[7]), .B(DB[832]), .Z(n12698) );
  IV U18987 ( .A(n12697), .Z(n18624) );
  XNOR U18988 ( .A(n12695), .B(n18625), .Z(n12697) );
  XNOR U18989 ( .A(q[6]), .B(DB[831]), .Z(n18625) );
  XNOR U18990 ( .A(q[5]), .B(DB[830]), .Z(n12695) );
  IV U18991 ( .A(n12708), .Z(n18622) );
  XOR U18992 ( .A(n18626), .B(n18627), .Z(n12708) );
  XNOR U18993 ( .A(n12704), .B(n12706), .Z(n18627) );
  XNOR U18994 ( .A(q[1]), .B(DB[826]), .Z(n12706) );
  XNOR U18995 ( .A(q[4]), .B(DB[829]), .Z(n12704) );
  IV U18996 ( .A(n12703), .Z(n18626) );
  XNOR U18997 ( .A(n12701), .B(n18628), .Z(n12703) );
  XNOR U18998 ( .A(q[3]), .B(DB[828]), .Z(n18628) );
  XNOR U18999 ( .A(q[2]), .B(DB[827]), .Z(n12701) );
  XOR U19000 ( .A(n18629), .B(n12599), .Z(n12527) );
  XOR U19001 ( .A(n18630), .B(n12591), .Z(n12599) );
  XOR U19002 ( .A(n18631), .B(n12580), .Z(n12591) );
  XNOR U19003 ( .A(q[14]), .B(DB[854]), .Z(n12580) );
  IV U19004 ( .A(n12579), .Z(n18631) );
  XNOR U19005 ( .A(n12577), .B(n18632), .Z(n12579) );
  XNOR U19006 ( .A(q[13]), .B(DB[853]), .Z(n18632) );
  XNOR U19007 ( .A(q[12]), .B(DB[852]), .Z(n12577) );
  IV U19008 ( .A(n12590), .Z(n18630) );
  XOR U19009 ( .A(n18633), .B(n18634), .Z(n12590) );
  XNOR U19010 ( .A(n12586), .B(n12588), .Z(n18634) );
  XNOR U19011 ( .A(q[8]), .B(DB[848]), .Z(n12588) );
  XNOR U19012 ( .A(q[11]), .B(DB[851]), .Z(n12586) );
  IV U19013 ( .A(n12585), .Z(n18633) );
  XNOR U19014 ( .A(n12583), .B(n18635), .Z(n12585) );
  XNOR U19015 ( .A(q[10]), .B(DB[850]), .Z(n18635) );
  XNOR U19016 ( .A(q[9]), .B(DB[849]), .Z(n12583) );
  IV U19017 ( .A(n12598), .Z(n18629) );
  XOR U19018 ( .A(n18636), .B(n18637), .Z(n12598) );
  XNOR U19019 ( .A(n12615), .B(n12596), .Z(n18637) );
  XNOR U19020 ( .A(q[0]), .B(DB[840]), .Z(n12596) );
  XOR U19021 ( .A(n18638), .B(n12604), .Z(n12615) );
  XNOR U19022 ( .A(q[7]), .B(DB[847]), .Z(n12604) );
  IV U19023 ( .A(n12603), .Z(n18638) );
  XNOR U19024 ( .A(n12601), .B(n18639), .Z(n12603) );
  XNOR U19025 ( .A(q[6]), .B(DB[846]), .Z(n18639) );
  XNOR U19026 ( .A(q[5]), .B(DB[845]), .Z(n12601) );
  IV U19027 ( .A(n12614), .Z(n18636) );
  XOR U19028 ( .A(n18640), .B(n18641), .Z(n12614) );
  XNOR U19029 ( .A(n12610), .B(n12612), .Z(n18641) );
  XNOR U19030 ( .A(q[1]), .B(DB[841]), .Z(n12612) );
  XNOR U19031 ( .A(q[4]), .B(DB[844]), .Z(n12610) );
  IV U19032 ( .A(n12609), .Z(n18640) );
  XNOR U19033 ( .A(n12607), .B(n18642), .Z(n12609) );
  XNOR U19034 ( .A(q[3]), .B(DB[843]), .Z(n18642) );
  XNOR U19035 ( .A(q[2]), .B(DB[842]), .Z(n12607) );
  XOR U19036 ( .A(n18643), .B(n12505), .Z(n12433) );
  XOR U19037 ( .A(n18644), .B(n12497), .Z(n12505) );
  XOR U19038 ( .A(n18645), .B(n12486), .Z(n12497) );
  XNOR U19039 ( .A(q[14]), .B(DB[869]), .Z(n12486) );
  IV U19040 ( .A(n12485), .Z(n18645) );
  XNOR U19041 ( .A(n12483), .B(n18646), .Z(n12485) );
  XNOR U19042 ( .A(q[13]), .B(DB[868]), .Z(n18646) );
  XNOR U19043 ( .A(q[12]), .B(DB[867]), .Z(n12483) );
  IV U19044 ( .A(n12496), .Z(n18644) );
  XOR U19045 ( .A(n18647), .B(n18648), .Z(n12496) );
  XNOR U19046 ( .A(n12492), .B(n12494), .Z(n18648) );
  XNOR U19047 ( .A(q[8]), .B(DB[863]), .Z(n12494) );
  XNOR U19048 ( .A(q[11]), .B(DB[866]), .Z(n12492) );
  IV U19049 ( .A(n12491), .Z(n18647) );
  XNOR U19050 ( .A(n12489), .B(n18649), .Z(n12491) );
  XNOR U19051 ( .A(q[10]), .B(DB[865]), .Z(n18649) );
  XNOR U19052 ( .A(q[9]), .B(DB[864]), .Z(n12489) );
  IV U19053 ( .A(n12504), .Z(n18643) );
  XOR U19054 ( .A(n18650), .B(n18651), .Z(n12504) );
  XNOR U19055 ( .A(n12521), .B(n12502), .Z(n18651) );
  XNOR U19056 ( .A(q[0]), .B(DB[855]), .Z(n12502) );
  XOR U19057 ( .A(n18652), .B(n12510), .Z(n12521) );
  XNOR U19058 ( .A(q[7]), .B(DB[862]), .Z(n12510) );
  IV U19059 ( .A(n12509), .Z(n18652) );
  XNOR U19060 ( .A(n12507), .B(n18653), .Z(n12509) );
  XNOR U19061 ( .A(q[6]), .B(DB[861]), .Z(n18653) );
  XNOR U19062 ( .A(q[5]), .B(DB[860]), .Z(n12507) );
  IV U19063 ( .A(n12520), .Z(n18650) );
  XOR U19064 ( .A(n18654), .B(n18655), .Z(n12520) );
  XNOR U19065 ( .A(n12516), .B(n12518), .Z(n18655) );
  XNOR U19066 ( .A(q[1]), .B(DB[856]), .Z(n12518) );
  XNOR U19067 ( .A(q[4]), .B(DB[859]), .Z(n12516) );
  IV U19068 ( .A(n12515), .Z(n18654) );
  XNOR U19069 ( .A(n12513), .B(n18656), .Z(n12515) );
  XNOR U19070 ( .A(q[3]), .B(DB[858]), .Z(n18656) );
  XNOR U19071 ( .A(q[2]), .B(DB[857]), .Z(n12513) );
  XOR U19072 ( .A(n18657), .B(n12411), .Z(n12339) );
  XOR U19073 ( .A(n18658), .B(n12403), .Z(n12411) );
  XOR U19074 ( .A(n18659), .B(n12392), .Z(n12403) );
  XNOR U19075 ( .A(q[14]), .B(DB[884]), .Z(n12392) );
  IV U19076 ( .A(n12391), .Z(n18659) );
  XNOR U19077 ( .A(n12389), .B(n18660), .Z(n12391) );
  XNOR U19078 ( .A(q[13]), .B(DB[883]), .Z(n18660) );
  XNOR U19079 ( .A(q[12]), .B(DB[882]), .Z(n12389) );
  IV U19080 ( .A(n12402), .Z(n18658) );
  XOR U19081 ( .A(n18661), .B(n18662), .Z(n12402) );
  XNOR U19082 ( .A(n12398), .B(n12400), .Z(n18662) );
  XNOR U19083 ( .A(q[8]), .B(DB[878]), .Z(n12400) );
  XNOR U19084 ( .A(q[11]), .B(DB[881]), .Z(n12398) );
  IV U19085 ( .A(n12397), .Z(n18661) );
  XNOR U19086 ( .A(n12395), .B(n18663), .Z(n12397) );
  XNOR U19087 ( .A(q[10]), .B(DB[880]), .Z(n18663) );
  XNOR U19088 ( .A(q[9]), .B(DB[879]), .Z(n12395) );
  IV U19089 ( .A(n12410), .Z(n18657) );
  XOR U19090 ( .A(n18664), .B(n18665), .Z(n12410) );
  XNOR U19091 ( .A(n12427), .B(n12408), .Z(n18665) );
  XNOR U19092 ( .A(q[0]), .B(DB[870]), .Z(n12408) );
  XOR U19093 ( .A(n18666), .B(n12416), .Z(n12427) );
  XNOR U19094 ( .A(q[7]), .B(DB[877]), .Z(n12416) );
  IV U19095 ( .A(n12415), .Z(n18666) );
  XNOR U19096 ( .A(n12413), .B(n18667), .Z(n12415) );
  XNOR U19097 ( .A(q[6]), .B(DB[876]), .Z(n18667) );
  XNOR U19098 ( .A(q[5]), .B(DB[875]), .Z(n12413) );
  IV U19099 ( .A(n12426), .Z(n18664) );
  XOR U19100 ( .A(n18668), .B(n18669), .Z(n12426) );
  XNOR U19101 ( .A(n12422), .B(n12424), .Z(n18669) );
  XNOR U19102 ( .A(q[1]), .B(DB[871]), .Z(n12424) );
  XNOR U19103 ( .A(q[4]), .B(DB[874]), .Z(n12422) );
  IV U19104 ( .A(n12421), .Z(n18668) );
  XNOR U19105 ( .A(n12419), .B(n18670), .Z(n12421) );
  XNOR U19106 ( .A(q[3]), .B(DB[873]), .Z(n18670) );
  XNOR U19107 ( .A(q[2]), .B(DB[872]), .Z(n12419) );
  XOR U19108 ( .A(n18671), .B(n12317), .Z(n12245) );
  XOR U19109 ( .A(n18672), .B(n12309), .Z(n12317) );
  XOR U19110 ( .A(n18673), .B(n12298), .Z(n12309) );
  XNOR U19111 ( .A(q[14]), .B(DB[899]), .Z(n12298) );
  IV U19112 ( .A(n12297), .Z(n18673) );
  XNOR U19113 ( .A(n12295), .B(n18674), .Z(n12297) );
  XNOR U19114 ( .A(q[13]), .B(DB[898]), .Z(n18674) );
  XNOR U19115 ( .A(q[12]), .B(DB[897]), .Z(n12295) );
  IV U19116 ( .A(n12308), .Z(n18672) );
  XOR U19117 ( .A(n18675), .B(n18676), .Z(n12308) );
  XNOR U19118 ( .A(n12304), .B(n12306), .Z(n18676) );
  XNOR U19119 ( .A(q[8]), .B(DB[893]), .Z(n12306) );
  XNOR U19120 ( .A(q[11]), .B(DB[896]), .Z(n12304) );
  IV U19121 ( .A(n12303), .Z(n18675) );
  XNOR U19122 ( .A(n12301), .B(n18677), .Z(n12303) );
  XNOR U19123 ( .A(q[10]), .B(DB[895]), .Z(n18677) );
  XNOR U19124 ( .A(q[9]), .B(DB[894]), .Z(n12301) );
  IV U19125 ( .A(n12316), .Z(n18671) );
  XOR U19126 ( .A(n18678), .B(n18679), .Z(n12316) );
  XNOR U19127 ( .A(n12333), .B(n12314), .Z(n18679) );
  XNOR U19128 ( .A(q[0]), .B(DB[885]), .Z(n12314) );
  XOR U19129 ( .A(n18680), .B(n12322), .Z(n12333) );
  XNOR U19130 ( .A(q[7]), .B(DB[892]), .Z(n12322) );
  IV U19131 ( .A(n12321), .Z(n18680) );
  XNOR U19132 ( .A(n12319), .B(n18681), .Z(n12321) );
  XNOR U19133 ( .A(q[6]), .B(DB[891]), .Z(n18681) );
  XNOR U19134 ( .A(q[5]), .B(DB[890]), .Z(n12319) );
  IV U19135 ( .A(n12332), .Z(n18678) );
  XOR U19136 ( .A(n18682), .B(n18683), .Z(n12332) );
  XNOR U19137 ( .A(n12328), .B(n12330), .Z(n18683) );
  XNOR U19138 ( .A(q[1]), .B(DB[886]), .Z(n12330) );
  XNOR U19139 ( .A(q[4]), .B(DB[889]), .Z(n12328) );
  IV U19140 ( .A(n12327), .Z(n18682) );
  XNOR U19141 ( .A(n12325), .B(n18684), .Z(n12327) );
  XNOR U19142 ( .A(q[3]), .B(DB[888]), .Z(n18684) );
  XNOR U19143 ( .A(q[2]), .B(DB[887]), .Z(n12325) );
  XOR U19144 ( .A(n18685), .B(n12223), .Z(n12151) );
  XOR U19145 ( .A(n18686), .B(n12215), .Z(n12223) );
  XOR U19146 ( .A(n18687), .B(n12204), .Z(n12215) );
  XNOR U19147 ( .A(q[14]), .B(DB[914]), .Z(n12204) );
  IV U19148 ( .A(n12203), .Z(n18687) );
  XNOR U19149 ( .A(n12201), .B(n18688), .Z(n12203) );
  XNOR U19150 ( .A(q[13]), .B(DB[913]), .Z(n18688) );
  XNOR U19151 ( .A(q[12]), .B(DB[912]), .Z(n12201) );
  IV U19152 ( .A(n12214), .Z(n18686) );
  XOR U19153 ( .A(n18689), .B(n18690), .Z(n12214) );
  XNOR U19154 ( .A(n12210), .B(n12212), .Z(n18690) );
  XNOR U19155 ( .A(q[8]), .B(DB[908]), .Z(n12212) );
  XNOR U19156 ( .A(q[11]), .B(DB[911]), .Z(n12210) );
  IV U19157 ( .A(n12209), .Z(n18689) );
  XNOR U19158 ( .A(n12207), .B(n18691), .Z(n12209) );
  XNOR U19159 ( .A(q[10]), .B(DB[910]), .Z(n18691) );
  XNOR U19160 ( .A(q[9]), .B(DB[909]), .Z(n12207) );
  IV U19161 ( .A(n12222), .Z(n18685) );
  XOR U19162 ( .A(n18692), .B(n18693), .Z(n12222) );
  XNOR U19163 ( .A(n12239), .B(n12220), .Z(n18693) );
  XNOR U19164 ( .A(q[0]), .B(DB[900]), .Z(n12220) );
  XOR U19165 ( .A(n18694), .B(n12228), .Z(n12239) );
  XNOR U19166 ( .A(q[7]), .B(DB[907]), .Z(n12228) );
  IV U19167 ( .A(n12227), .Z(n18694) );
  XNOR U19168 ( .A(n12225), .B(n18695), .Z(n12227) );
  XNOR U19169 ( .A(q[6]), .B(DB[906]), .Z(n18695) );
  XNOR U19170 ( .A(q[5]), .B(DB[905]), .Z(n12225) );
  IV U19171 ( .A(n12238), .Z(n18692) );
  XOR U19172 ( .A(n18696), .B(n18697), .Z(n12238) );
  XNOR U19173 ( .A(n12234), .B(n12236), .Z(n18697) );
  XNOR U19174 ( .A(q[1]), .B(DB[901]), .Z(n12236) );
  XNOR U19175 ( .A(q[4]), .B(DB[904]), .Z(n12234) );
  IV U19176 ( .A(n12233), .Z(n18696) );
  XNOR U19177 ( .A(n12231), .B(n18698), .Z(n12233) );
  XNOR U19178 ( .A(q[3]), .B(DB[903]), .Z(n18698) );
  XNOR U19179 ( .A(q[2]), .B(DB[902]), .Z(n12231) );
  XOR U19180 ( .A(n18699), .B(n12129), .Z(n12057) );
  XOR U19181 ( .A(n18700), .B(n12121), .Z(n12129) );
  XOR U19182 ( .A(n18701), .B(n12110), .Z(n12121) );
  XNOR U19183 ( .A(q[14]), .B(DB[929]), .Z(n12110) );
  IV U19184 ( .A(n12109), .Z(n18701) );
  XNOR U19185 ( .A(n12107), .B(n18702), .Z(n12109) );
  XNOR U19186 ( .A(q[13]), .B(DB[928]), .Z(n18702) );
  XNOR U19187 ( .A(q[12]), .B(DB[927]), .Z(n12107) );
  IV U19188 ( .A(n12120), .Z(n18700) );
  XOR U19189 ( .A(n18703), .B(n18704), .Z(n12120) );
  XNOR U19190 ( .A(n12116), .B(n12118), .Z(n18704) );
  XNOR U19191 ( .A(q[8]), .B(DB[923]), .Z(n12118) );
  XNOR U19192 ( .A(q[11]), .B(DB[926]), .Z(n12116) );
  IV U19193 ( .A(n12115), .Z(n18703) );
  XNOR U19194 ( .A(n12113), .B(n18705), .Z(n12115) );
  XNOR U19195 ( .A(q[10]), .B(DB[925]), .Z(n18705) );
  XNOR U19196 ( .A(q[9]), .B(DB[924]), .Z(n12113) );
  IV U19197 ( .A(n12128), .Z(n18699) );
  XOR U19198 ( .A(n18706), .B(n18707), .Z(n12128) );
  XNOR U19199 ( .A(n12145), .B(n12126), .Z(n18707) );
  XNOR U19200 ( .A(q[0]), .B(DB[915]), .Z(n12126) );
  XOR U19201 ( .A(n18708), .B(n12134), .Z(n12145) );
  XNOR U19202 ( .A(q[7]), .B(DB[922]), .Z(n12134) );
  IV U19203 ( .A(n12133), .Z(n18708) );
  XNOR U19204 ( .A(n12131), .B(n18709), .Z(n12133) );
  XNOR U19205 ( .A(q[6]), .B(DB[921]), .Z(n18709) );
  XNOR U19206 ( .A(q[5]), .B(DB[920]), .Z(n12131) );
  IV U19207 ( .A(n12144), .Z(n18706) );
  XOR U19208 ( .A(n18710), .B(n18711), .Z(n12144) );
  XNOR U19209 ( .A(n12140), .B(n12142), .Z(n18711) );
  XNOR U19210 ( .A(q[1]), .B(DB[916]), .Z(n12142) );
  XNOR U19211 ( .A(q[4]), .B(DB[919]), .Z(n12140) );
  IV U19212 ( .A(n12139), .Z(n18710) );
  XNOR U19213 ( .A(n12137), .B(n18712), .Z(n12139) );
  XNOR U19214 ( .A(q[3]), .B(DB[918]), .Z(n18712) );
  XNOR U19215 ( .A(q[2]), .B(DB[917]), .Z(n12137) );
  XOR U19216 ( .A(n18713), .B(n12035), .Z(n11963) );
  XOR U19217 ( .A(n18714), .B(n12027), .Z(n12035) );
  XOR U19218 ( .A(n18715), .B(n12016), .Z(n12027) );
  XNOR U19219 ( .A(q[14]), .B(DB[944]), .Z(n12016) );
  IV U19220 ( .A(n12015), .Z(n18715) );
  XNOR U19221 ( .A(n12013), .B(n18716), .Z(n12015) );
  XNOR U19222 ( .A(q[13]), .B(DB[943]), .Z(n18716) );
  XNOR U19223 ( .A(q[12]), .B(DB[942]), .Z(n12013) );
  IV U19224 ( .A(n12026), .Z(n18714) );
  XOR U19225 ( .A(n18717), .B(n18718), .Z(n12026) );
  XNOR U19226 ( .A(n12022), .B(n12024), .Z(n18718) );
  XNOR U19227 ( .A(q[8]), .B(DB[938]), .Z(n12024) );
  XNOR U19228 ( .A(q[11]), .B(DB[941]), .Z(n12022) );
  IV U19229 ( .A(n12021), .Z(n18717) );
  XNOR U19230 ( .A(n12019), .B(n18719), .Z(n12021) );
  XNOR U19231 ( .A(q[10]), .B(DB[940]), .Z(n18719) );
  XNOR U19232 ( .A(q[9]), .B(DB[939]), .Z(n12019) );
  IV U19233 ( .A(n12034), .Z(n18713) );
  XOR U19234 ( .A(n18720), .B(n18721), .Z(n12034) );
  XNOR U19235 ( .A(n12051), .B(n12032), .Z(n18721) );
  XNOR U19236 ( .A(q[0]), .B(DB[930]), .Z(n12032) );
  XOR U19237 ( .A(n18722), .B(n12040), .Z(n12051) );
  XNOR U19238 ( .A(q[7]), .B(DB[937]), .Z(n12040) );
  IV U19239 ( .A(n12039), .Z(n18722) );
  XNOR U19240 ( .A(n12037), .B(n18723), .Z(n12039) );
  XNOR U19241 ( .A(q[6]), .B(DB[936]), .Z(n18723) );
  XNOR U19242 ( .A(q[5]), .B(DB[935]), .Z(n12037) );
  IV U19243 ( .A(n12050), .Z(n18720) );
  XOR U19244 ( .A(n18724), .B(n18725), .Z(n12050) );
  XNOR U19245 ( .A(n12046), .B(n12048), .Z(n18725) );
  XNOR U19246 ( .A(q[1]), .B(DB[931]), .Z(n12048) );
  XNOR U19247 ( .A(q[4]), .B(DB[934]), .Z(n12046) );
  IV U19248 ( .A(n12045), .Z(n18724) );
  XNOR U19249 ( .A(n12043), .B(n18726), .Z(n12045) );
  XNOR U19250 ( .A(q[3]), .B(DB[933]), .Z(n18726) );
  XNOR U19251 ( .A(q[2]), .B(DB[932]), .Z(n12043) );
  XOR U19252 ( .A(n18727), .B(n11941), .Z(n11869) );
  XOR U19253 ( .A(n18728), .B(n11933), .Z(n11941) );
  XOR U19254 ( .A(n18729), .B(n11922), .Z(n11933) );
  XNOR U19255 ( .A(q[14]), .B(DB[959]), .Z(n11922) );
  IV U19256 ( .A(n11921), .Z(n18729) );
  XNOR U19257 ( .A(n11919), .B(n18730), .Z(n11921) );
  XNOR U19258 ( .A(q[13]), .B(DB[958]), .Z(n18730) );
  XNOR U19259 ( .A(q[12]), .B(DB[957]), .Z(n11919) );
  IV U19260 ( .A(n11932), .Z(n18728) );
  XOR U19261 ( .A(n18731), .B(n18732), .Z(n11932) );
  XNOR U19262 ( .A(n11928), .B(n11930), .Z(n18732) );
  XNOR U19263 ( .A(q[8]), .B(DB[953]), .Z(n11930) );
  XNOR U19264 ( .A(q[11]), .B(DB[956]), .Z(n11928) );
  IV U19265 ( .A(n11927), .Z(n18731) );
  XNOR U19266 ( .A(n11925), .B(n18733), .Z(n11927) );
  XNOR U19267 ( .A(q[10]), .B(DB[955]), .Z(n18733) );
  XNOR U19268 ( .A(q[9]), .B(DB[954]), .Z(n11925) );
  IV U19269 ( .A(n11940), .Z(n18727) );
  XOR U19270 ( .A(n18734), .B(n18735), .Z(n11940) );
  XNOR U19271 ( .A(n11957), .B(n11938), .Z(n18735) );
  XNOR U19272 ( .A(q[0]), .B(DB[945]), .Z(n11938) );
  XOR U19273 ( .A(n18736), .B(n11946), .Z(n11957) );
  XNOR U19274 ( .A(q[7]), .B(DB[952]), .Z(n11946) );
  IV U19275 ( .A(n11945), .Z(n18736) );
  XNOR U19276 ( .A(n11943), .B(n18737), .Z(n11945) );
  XNOR U19277 ( .A(q[6]), .B(DB[951]), .Z(n18737) );
  XNOR U19278 ( .A(q[5]), .B(DB[950]), .Z(n11943) );
  IV U19279 ( .A(n11956), .Z(n18734) );
  XOR U19280 ( .A(n18738), .B(n18739), .Z(n11956) );
  XNOR U19281 ( .A(n11952), .B(n11954), .Z(n18739) );
  XNOR U19282 ( .A(q[1]), .B(DB[946]), .Z(n11954) );
  XNOR U19283 ( .A(q[4]), .B(DB[949]), .Z(n11952) );
  IV U19284 ( .A(n11951), .Z(n18738) );
  XNOR U19285 ( .A(n11949), .B(n18740), .Z(n11951) );
  XNOR U19286 ( .A(q[3]), .B(DB[948]), .Z(n18740) );
  XNOR U19287 ( .A(q[2]), .B(DB[947]), .Z(n11949) );
  XOR U19288 ( .A(n18741), .B(n11847), .Z(n11775) );
  XOR U19289 ( .A(n18742), .B(n11839), .Z(n11847) );
  XOR U19290 ( .A(n18743), .B(n11828), .Z(n11839) );
  XNOR U19291 ( .A(q[14]), .B(DB[974]), .Z(n11828) );
  IV U19292 ( .A(n11827), .Z(n18743) );
  XNOR U19293 ( .A(n11825), .B(n18744), .Z(n11827) );
  XNOR U19294 ( .A(q[13]), .B(DB[973]), .Z(n18744) );
  XNOR U19295 ( .A(q[12]), .B(DB[972]), .Z(n11825) );
  IV U19296 ( .A(n11838), .Z(n18742) );
  XOR U19297 ( .A(n18745), .B(n18746), .Z(n11838) );
  XNOR U19298 ( .A(n11834), .B(n11836), .Z(n18746) );
  XNOR U19299 ( .A(q[8]), .B(DB[968]), .Z(n11836) );
  XNOR U19300 ( .A(q[11]), .B(DB[971]), .Z(n11834) );
  IV U19301 ( .A(n11833), .Z(n18745) );
  XNOR U19302 ( .A(n11831), .B(n18747), .Z(n11833) );
  XNOR U19303 ( .A(q[10]), .B(DB[970]), .Z(n18747) );
  XNOR U19304 ( .A(q[9]), .B(DB[969]), .Z(n11831) );
  IV U19305 ( .A(n11846), .Z(n18741) );
  XOR U19306 ( .A(n18748), .B(n18749), .Z(n11846) );
  XNOR U19307 ( .A(n11863), .B(n11844), .Z(n18749) );
  XNOR U19308 ( .A(q[0]), .B(DB[960]), .Z(n11844) );
  XOR U19309 ( .A(n18750), .B(n11852), .Z(n11863) );
  XNOR U19310 ( .A(q[7]), .B(DB[967]), .Z(n11852) );
  IV U19311 ( .A(n11851), .Z(n18750) );
  XNOR U19312 ( .A(n11849), .B(n18751), .Z(n11851) );
  XNOR U19313 ( .A(q[6]), .B(DB[966]), .Z(n18751) );
  XNOR U19314 ( .A(q[5]), .B(DB[965]), .Z(n11849) );
  IV U19315 ( .A(n11862), .Z(n18748) );
  XOR U19316 ( .A(n18752), .B(n18753), .Z(n11862) );
  XNOR U19317 ( .A(n11858), .B(n11860), .Z(n18753) );
  XNOR U19318 ( .A(q[1]), .B(DB[961]), .Z(n11860) );
  XNOR U19319 ( .A(q[4]), .B(DB[964]), .Z(n11858) );
  IV U19320 ( .A(n11857), .Z(n18752) );
  XNOR U19321 ( .A(n11855), .B(n18754), .Z(n11857) );
  XNOR U19322 ( .A(q[3]), .B(DB[963]), .Z(n18754) );
  XNOR U19323 ( .A(q[2]), .B(DB[962]), .Z(n11855) );
  XOR U19324 ( .A(n18755), .B(n11753), .Z(n11681) );
  XOR U19325 ( .A(n18756), .B(n11745), .Z(n11753) );
  XOR U19326 ( .A(n18757), .B(n11734), .Z(n11745) );
  XNOR U19327 ( .A(q[14]), .B(DB[989]), .Z(n11734) );
  IV U19328 ( .A(n11733), .Z(n18757) );
  XNOR U19329 ( .A(n11731), .B(n18758), .Z(n11733) );
  XNOR U19330 ( .A(q[13]), .B(DB[988]), .Z(n18758) );
  XNOR U19331 ( .A(q[12]), .B(DB[987]), .Z(n11731) );
  IV U19332 ( .A(n11744), .Z(n18756) );
  XOR U19333 ( .A(n18759), .B(n18760), .Z(n11744) );
  XNOR U19334 ( .A(n11740), .B(n11742), .Z(n18760) );
  XNOR U19335 ( .A(q[8]), .B(DB[983]), .Z(n11742) );
  XNOR U19336 ( .A(q[11]), .B(DB[986]), .Z(n11740) );
  IV U19337 ( .A(n11739), .Z(n18759) );
  XNOR U19338 ( .A(n11737), .B(n18761), .Z(n11739) );
  XNOR U19339 ( .A(q[10]), .B(DB[985]), .Z(n18761) );
  XNOR U19340 ( .A(q[9]), .B(DB[984]), .Z(n11737) );
  IV U19341 ( .A(n11752), .Z(n18755) );
  XOR U19342 ( .A(n18762), .B(n18763), .Z(n11752) );
  XNOR U19343 ( .A(n11769), .B(n11750), .Z(n18763) );
  XNOR U19344 ( .A(q[0]), .B(DB[975]), .Z(n11750) );
  XOR U19345 ( .A(n18764), .B(n11758), .Z(n11769) );
  XNOR U19346 ( .A(q[7]), .B(DB[982]), .Z(n11758) );
  IV U19347 ( .A(n11757), .Z(n18764) );
  XNOR U19348 ( .A(n11755), .B(n18765), .Z(n11757) );
  XNOR U19349 ( .A(q[6]), .B(DB[981]), .Z(n18765) );
  XNOR U19350 ( .A(q[5]), .B(DB[980]), .Z(n11755) );
  IV U19351 ( .A(n11768), .Z(n18762) );
  XOR U19352 ( .A(n18766), .B(n18767), .Z(n11768) );
  XNOR U19353 ( .A(n11764), .B(n11766), .Z(n18767) );
  XNOR U19354 ( .A(q[1]), .B(DB[976]), .Z(n11766) );
  XNOR U19355 ( .A(q[4]), .B(DB[979]), .Z(n11764) );
  IV U19356 ( .A(n11763), .Z(n18766) );
  XNOR U19357 ( .A(n11761), .B(n18768), .Z(n11763) );
  XNOR U19358 ( .A(q[3]), .B(DB[978]), .Z(n18768) );
  XNOR U19359 ( .A(q[2]), .B(DB[977]), .Z(n11761) );
  XOR U19360 ( .A(n18769), .B(n11659), .Z(n11587) );
  XOR U19361 ( .A(n18770), .B(n11651), .Z(n11659) );
  XOR U19362 ( .A(n18771), .B(n11640), .Z(n11651) );
  XNOR U19363 ( .A(q[14]), .B(DB[1004]), .Z(n11640) );
  IV U19364 ( .A(n11639), .Z(n18771) );
  XNOR U19365 ( .A(n11637), .B(n18772), .Z(n11639) );
  XNOR U19366 ( .A(q[13]), .B(DB[1003]), .Z(n18772) );
  XNOR U19367 ( .A(q[12]), .B(DB[1002]), .Z(n11637) );
  IV U19368 ( .A(n11650), .Z(n18770) );
  XOR U19369 ( .A(n18773), .B(n18774), .Z(n11650) );
  XNOR U19370 ( .A(n11646), .B(n11648), .Z(n18774) );
  XNOR U19371 ( .A(q[8]), .B(DB[998]), .Z(n11648) );
  XNOR U19372 ( .A(q[11]), .B(DB[1001]), .Z(n11646) );
  IV U19373 ( .A(n11645), .Z(n18773) );
  XNOR U19374 ( .A(n11643), .B(n18775), .Z(n11645) );
  XNOR U19375 ( .A(q[10]), .B(DB[1000]), .Z(n18775) );
  XNOR U19376 ( .A(q[9]), .B(DB[999]), .Z(n11643) );
  IV U19377 ( .A(n11658), .Z(n18769) );
  XOR U19378 ( .A(n18776), .B(n18777), .Z(n11658) );
  XNOR U19379 ( .A(n11675), .B(n11656), .Z(n18777) );
  XNOR U19380 ( .A(q[0]), .B(DB[990]), .Z(n11656) );
  XOR U19381 ( .A(n18778), .B(n11664), .Z(n11675) );
  XNOR U19382 ( .A(q[7]), .B(DB[997]), .Z(n11664) );
  IV U19383 ( .A(n11663), .Z(n18778) );
  XNOR U19384 ( .A(n11661), .B(n18779), .Z(n11663) );
  XNOR U19385 ( .A(q[6]), .B(DB[996]), .Z(n18779) );
  XNOR U19386 ( .A(q[5]), .B(DB[995]), .Z(n11661) );
  IV U19387 ( .A(n11674), .Z(n18776) );
  XOR U19388 ( .A(n18780), .B(n18781), .Z(n11674) );
  XNOR U19389 ( .A(n11670), .B(n11672), .Z(n18781) );
  XNOR U19390 ( .A(q[1]), .B(DB[991]), .Z(n11672) );
  XNOR U19391 ( .A(q[4]), .B(DB[994]), .Z(n11670) );
  IV U19392 ( .A(n11669), .Z(n18780) );
  XNOR U19393 ( .A(n11667), .B(n18782), .Z(n11669) );
  XNOR U19394 ( .A(q[3]), .B(DB[993]), .Z(n18782) );
  XNOR U19395 ( .A(q[2]), .B(DB[992]), .Z(n11667) );
  XOR U19396 ( .A(n18783), .B(n11565), .Z(n11493) );
  XOR U19397 ( .A(n18784), .B(n11557), .Z(n11565) );
  XOR U19398 ( .A(n18785), .B(n11546), .Z(n11557) );
  XNOR U19399 ( .A(q[14]), .B(DB[1019]), .Z(n11546) );
  IV U19400 ( .A(n11545), .Z(n18785) );
  XNOR U19401 ( .A(n11543), .B(n18786), .Z(n11545) );
  XNOR U19402 ( .A(q[13]), .B(DB[1018]), .Z(n18786) );
  XNOR U19403 ( .A(q[12]), .B(DB[1017]), .Z(n11543) );
  IV U19404 ( .A(n11556), .Z(n18784) );
  XOR U19405 ( .A(n18787), .B(n18788), .Z(n11556) );
  XNOR U19406 ( .A(n11552), .B(n11554), .Z(n18788) );
  XNOR U19407 ( .A(q[8]), .B(DB[1013]), .Z(n11554) );
  XNOR U19408 ( .A(q[11]), .B(DB[1016]), .Z(n11552) );
  IV U19409 ( .A(n11551), .Z(n18787) );
  XNOR U19410 ( .A(n11549), .B(n18789), .Z(n11551) );
  XNOR U19411 ( .A(q[10]), .B(DB[1015]), .Z(n18789) );
  XNOR U19412 ( .A(q[9]), .B(DB[1014]), .Z(n11549) );
  IV U19413 ( .A(n11564), .Z(n18783) );
  XOR U19414 ( .A(n18790), .B(n18791), .Z(n11564) );
  XNOR U19415 ( .A(n11581), .B(n11562), .Z(n18791) );
  XNOR U19416 ( .A(q[0]), .B(DB[1005]), .Z(n11562) );
  XOR U19417 ( .A(n18792), .B(n11570), .Z(n11581) );
  XNOR U19418 ( .A(q[7]), .B(DB[1012]), .Z(n11570) );
  IV U19419 ( .A(n11569), .Z(n18792) );
  XNOR U19420 ( .A(n11567), .B(n18793), .Z(n11569) );
  XNOR U19421 ( .A(q[6]), .B(DB[1011]), .Z(n18793) );
  XNOR U19422 ( .A(q[5]), .B(DB[1010]), .Z(n11567) );
  IV U19423 ( .A(n11580), .Z(n18790) );
  XOR U19424 ( .A(n18794), .B(n18795), .Z(n11580) );
  XNOR U19425 ( .A(n11576), .B(n11578), .Z(n18795) );
  XNOR U19426 ( .A(q[1]), .B(DB[1006]), .Z(n11578) );
  XNOR U19427 ( .A(q[4]), .B(DB[1009]), .Z(n11576) );
  IV U19428 ( .A(n11575), .Z(n18794) );
  XNOR U19429 ( .A(n11573), .B(n18796), .Z(n11575) );
  XNOR U19430 ( .A(q[3]), .B(DB[1008]), .Z(n18796) );
  XNOR U19431 ( .A(q[2]), .B(DB[1007]), .Z(n11573) );
  XOR U19432 ( .A(n18797), .B(n11471), .Z(n11399) );
  XOR U19433 ( .A(n18798), .B(n11463), .Z(n11471) );
  XOR U19434 ( .A(n18799), .B(n11452), .Z(n11463) );
  XNOR U19435 ( .A(q[14]), .B(DB[1034]), .Z(n11452) );
  IV U19436 ( .A(n11451), .Z(n18799) );
  XNOR U19437 ( .A(n11449), .B(n18800), .Z(n11451) );
  XNOR U19438 ( .A(q[13]), .B(DB[1033]), .Z(n18800) );
  XNOR U19439 ( .A(q[12]), .B(DB[1032]), .Z(n11449) );
  IV U19440 ( .A(n11462), .Z(n18798) );
  XOR U19441 ( .A(n18801), .B(n18802), .Z(n11462) );
  XNOR U19442 ( .A(n11458), .B(n11460), .Z(n18802) );
  XNOR U19443 ( .A(q[8]), .B(DB[1028]), .Z(n11460) );
  XNOR U19444 ( .A(q[11]), .B(DB[1031]), .Z(n11458) );
  IV U19445 ( .A(n11457), .Z(n18801) );
  XNOR U19446 ( .A(n11455), .B(n18803), .Z(n11457) );
  XNOR U19447 ( .A(q[10]), .B(DB[1030]), .Z(n18803) );
  XNOR U19448 ( .A(q[9]), .B(DB[1029]), .Z(n11455) );
  IV U19449 ( .A(n11470), .Z(n18797) );
  XOR U19450 ( .A(n18804), .B(n18805), .Z(n11470) );
  XNOR U19451 ( .A(n11487), .B(n11468), .Z(n18805) );
  XNOR U19452 ( .A(q[0]), .B(DB[1020]), .Z(n11468) );
  XOR U19453 ( .A(n18806), .B(n11476), .Z(n11487) );
  XNOR U19454 ( .A(q[7]), .B(DB[1027]), .Z(n11476) );
  IV U19455 ( .A(n11475), .Z(n18806) );
  XNOR U19456 ( .A(n11473), .B(n18807), .Z(n11475) );
  XNOR U19457 ( .A(q[6]), .B(DB[1026]), .Z(n18807) );
  XNOR U19458 ( .A(q[5]), .B(DB[1025]), .Z(n11473) );
  IV U19459 ( .A(n11486), .Z(n18804) );
  XOR U19460 ( .A(n18808), .B(n18809), .Z(n11486) );
  XNOR U19461 ( .A(n11482), .B(n11484), .Z(n18809) );
  XNOR U19462 ( .A(q[1]), .B(DB[1021]), .Z(n11484) );
  XNOR U19463 ( .A(q[4]), .B(DB[1024]), .Z(n11482) );
  IV U19464 ( .A(n11481), .Z(n18808) );
  XNOR U19465 ( .A(n11479), .B(n18810), .Z(n11481) );
  XNOR U19466 ( .A(q[3]), .B(DB[1023]), .Z(n18810) );
  XNOR U19467 ( .A(q[2]), .B(DB[1022]), .Z(n11479) );
  XOR U19468 ( .A(n18811), .B(n11377), .Z(n11305) );
  XOR U19469 ( .A(n18812), .B(n11369), .Z(n11377) );
  XOR U19470 ( .A(n18813), .B(n11358), .Z(n11369) );
  XNOR U19471 ( .A(q[14]), .B(DB[1049]), .Z(n11358) );
  IV U19472 ( .A(n11357), .Z(n18813) );
  XNOR U19473 ( .A(n11355), .B(n18814), .Z(n11357) );
  XNOR U19474 ( .A(q[13]), .B(DB[1048]), .Z(n18814) );
  XNOR U19475 ( .A(q[12]), .B(DB[1047]), .Z(n11355) );
  IV U19476 ( .A(n11368), .Z(n18812) );
  XOR U19477 ( .A(n18815), .B(n18816), .Z(n11368) );
  XNOR U19478 ( .A(n11364), .B(n11366), .Z(n18816) );
  XNOR U19479 ( .A(q[8]), .B(DB[1043]), .Z(n11366) );
  XNOR U19480 ( .A(q[11]), .B(DB[1046]), .Z(n11364) );
  IV U19481 ( .A(n11363), .Z(n18815) );
  XNOR U19482 ( .A(n11361), .B(n18817), .Z(n11363) );
  XNOR U19483 ( .A(q[10]), .B(DB[1045]), .Z(n18817) );
  XNOR U19484 ( .A(q[9]), .B(DB[1044]), .Z(n11361) );
  IV U19485 ( .A(n11376), .Z(n18811) );
  XOR U19486 ( .A(n18818), .B(n18819), .Z(n11376) );
  XNOR U19487 ( .A(n11393), .B(n11374), .Z(n18819) );
  XNOR U19488 ( .A(q[0]), .B(DB[1035]), .Z(n11374) );
  XOR U19489 ( .A(n18820), .B(n11382), .Z(n11393) );
  XNOR U19490 ( .A(q[7]), .B(DB[1042]), .Z(n11382) );
  IV U19491 ( .A(n11381), .Z(n18820) );
  XNOR U19492 ( .A(n11379), .B(n18821), .Z(n11381) );
  XNOR U19493 ( .A(q[6]), .B(DB[1041]), .Z(n18821) );
  XNOR U19494 ( .A(q[5]), .B(DB[1040]), .Z(n11379) );
  IV U19495 ( .A(n11392), .Z(n18818) );
  XOR U19496 ( .A(n18822), .B(n18823), .Z(n11392) );
  XNOR U19497 ( .A(n11388), .B(n11390), .Z(n18823) );
  XNOR U19498 ( .A(q[1]), .B(DB[1036]), .Z(n11390) );
  XNOR U19499 ( .A(q[4]), .B(DB[1039]), .Z(n11388) );
  IV U19500 ( .A(n11387), .Z(n18822) );
  XNOR U19501 ( .A(n11385), .B(n18824), .Z(n11387) );
  XNOR U19502 ( .A(q[3]), .B(DB[1038]), .Z(n18824) );
  XNOR U19503 ( .A(q[2]), .B(DB[1037]), .Z(n11385) );
  XOR U19504 ( .A(n18825), .B(n11283), .Z(n11211) );
  XOR U19505 ( .A(n18826), .B(n11275), .Z(n11283) );
  XOR U19506 ( .A(n18827), .B(n11264), .Z(n11275) );
  XNOR U19507 ( .A(q[14]), .B(DB[1064]), .Z(n11264) );
  IV U19508 ( .A(n11263), .Z(n18827) );
  XNOR U19509 ( .A(n11261), .B(n18828), .Z(n11263) );
  XNOR U19510 ( .A(q[13]), .B(DB[1063]), .Z(n18828) );
  XNOR U19511 ( .A(q[12]), .B(DB[1062]), .Z(n11261) );
  IV U19512 ( .A(n11274), .Z(n18826) );
  XOR U19513 ( .A(n18829), .B(n18830), .Z(n11274) );
  XNOR U19514 ( .A(n11270), .B(n11272), .Z(n18830) );
  XNOR U19515 ( .A(q[8]), .B(DB[1058]), .Z(n11272) );
  XNOR U19516 ( .A(q[11]), .B(DB[1061]), .Z(n11270) );
  IV U19517 ( .A(n11269), .Z(n18829) );
  XNOR U19518 ( .A(n11267), .B(n18831), .Z(n11269) );
  XNOR U19519 ( .A(q[10]), .B(DB[1060]), .Z(n18831) );
  XNOR U19520 ( .A(q[9]), .B(DB[1059]), .Z(n11267) );
  IV U19521 ( .A(n11282), .Z(n18825) );
  XOR U19522 ( .A(n18832), .B(n18833), .Z(n11282) );
  XNOR U19523 ( .A(n11299), .B(n11280), .Z(n18833) );
  XNOR U19524 ( .A(q[0]), .B(DB[1050]), .Z(n11280) );
  XOR U19525 ( .A(n18834), .B(n11288), .Z(n11299) );
  XNOR U19526 ( .A(q[7]), .B(DB[1057]), .Z(n11288) );
  IV U19527 ( .A(n11287), .Z(n18834) );
  XNOR U19528 ( .A(n11285), .B(n18835), .Z(n11287) );
  XNOR U19529 ( .A(q[6]), .B(DB[1056]), .Z(n18835) );
  XNOR U19530 ( .A(q[5]), .B(DB[1055]), .Z(n11285) );
  IV U19531 ( .A(n11298), .Z(n18832) );
  XOR U19532 ( .A(n18836), .B(n18837), .Z(n11298) );
  XNOR U19533 ( .A(n11294), .B(n11296), .Z(n18837) );
  XNOR U19534 ( .A(q[1]), .B(DB[1051]), .Z(n11296) );
  XNOR U19535 ( .A(q[4]), .B(DB[1054]), .Z(n11294) );
  IV U19536 ( .A(n11293), .Z(n18836) );
  XNOR U19537 ( .A(n11291), .B(n18838), .Z(n11293) );
  XNOR U19538 ( .A(q[3]), .B(DB[1053]), .Z(n18838) );
  XNOR U19539 ( .A(q[2]), .B(DB[1052]), .Z(n11291) );
  XOR U19540 ( .A(n18839), .B(n11189), .Z(n11117) );
  XOR U19541 ( .A(n18840), .B(n11181), .Z(n11189) );
  XOR U19542 ( .A(n18841), .B(n11170), .Z(n11181) );
  XNOR U19543 ( .A(q[14]), .B(DB[1079]), .Z(n11170) );
  IV U19544 ( .A(n11169), .Z(n18841) );
  XNOR U19545 ( .A(n11167), .B(n18842), .Z(n11169) );
  XNOR U19546 ( .A(q[13]), .B(DB[1078]), .Z(n18842) );
  XNOR U19547 ( .A(q[12]), .B(DB[1077]), .Z(n11167) );
  IV U19548 ( .A(n11180), .Z(n18840) );
  XOR U19549 ( .A(n18843), .B(n18844), .Z(n11180) );
  XNOR U19550 ( .A(n11176), .B(n11178), .Z(n18844) );
  XNOR U19551 ( .A(q[8]), .B(DB[1073]), .Z(n11178) );
  XNOR U19552 ( .A(q[11]), .B(DB[1076]), .Z(n11176) );
  IV U19553 ( .A(n11175), .Z(n18843) );
  XNOR U19554 ( .A(n11173), .B(n18845), .Z(n11175) );
  XNOR U19555 ( .A(q[10]), .B(DB[1075]), .Z(n18845) );
  XNOR U19556 ( .A(q[9]), .B(DB[1074]), .Z(n11173) );
  IV U19557 ( .A(n11188), .Z(n18839) );
  XOR U19558 ( .A(n18846), .B(n18847), .Z(n11188) );
  XNOR U19559 ( .A(n11205), .B(n11186), .Z(n18847) );
  XNOR U19560 ( .A(q[0]), .B(DB[1065]), .Z(n11186) );
  XOR U19561 ( .A(n18848), .B(n11194), .Z(n11205) );
  XNOR U19562 ( .A(q[7]), .B(DB[1072]), .Z(n11194) );
  IV U19563 ( .A(n11193), .Z(n18848) );
  XNOR U19564 ( .A(n11191), .B(n18849), .Z(n11193) );
  XNOR U19565 ( .A(q[6]), .B(DB[1071]), .Z(n18849) );
  XNOR U19566 ( .A(q[5]), .B(DB[1070]), .Z(n11191) );
  IV U19567 ( .A(n11204), .Z(n18846) );
  XOR U19568 ( .A(n18850), .B(n18851), .Z(n11204) );
  XNOR U19569 ( .A(n11200), .B(n11202), .Z(n18851) );
  XNOR U19570 ( .A(q[1]), .B(DB[1066]), .Z(n11202) );
  XNOR U19571 ( .A(q[4]), .B(DB[1069]), .Z(n11200) );
  IV U19572 ( .A(n11199), .Z(n18850) );
  XNOR U19573 ( .A(n11197), .B(n18852), .Z(n11199) );
  XNOR U19574 ( .A(q[3]), .B(DB[1068]), .Z(n18852) );
  XNOR U19575 ( .A(q[2]), .B(DB[1067]), .Z(n11197) );
  XOR U19576 ( .A(n18853), .B(n11095), .Z(n11023) );
  XOR U19577 ( .A(n18854), .B(n11087), .Z(n11095) );
  XOR U19578 ( .A(n18855), .B(n11076), .Z(n11087) );
  XNOR U19579 ( .A(q[14]), .B(DB[1094]), .Z(n11076) );
  IV U19580 ( .A(n11075), .Z(n18855) );
  XNOR U19581 ( .A(n11073), .B(n18856), .Z(n11075) );
  XNOR U19582 ( .A(q[13]), .B(DB[1093]), .Z(n18856) );
  XNOR U19583 ( .A(q[12]), .B(DB[1092]), .Z(n11073) );
  IV U19584 ( .A(n11086), .Z(n18854) );
  XOR U19585 ( .A(n18857), .B(n18858), .Z(n11086) );
  XNOR U19586 ( .A(n11082), .B(n11084), .Z(n18858) );
  XNOR U19587 ( .A(q[8]), .B(DB[1088]), .Z(n11084) );
  XNOR U19588 ( .A(q[11]), .B(DB[1091]), .Z(n11082) );
  IV U19589 ( .A(n11081), .Z(n18857) );
  XNOR U19590 ( .A(n11079), .B(n18859), .Z(n11081) );
  XNOR U19591 ( .A(q[10]), .B(DB[1090]), .Z(n18859) );
  XNOR U19592 ( .A(q[9]), .B(DB[1089]), .Z(n11079) );
  IV U19593 ( .A(n11094), .Z(n18853) );
  XOR U19594 ( .A(n18860), .B(n18861), .Z(n11094) );
  XNOR U19595 ( .A(n11111), .B(n11092), .Z(n18861) );
  XNOR U19596 ( .A(q[0]), .B(DB[1080]), .Z(n11092) );
  XOR U19597 ( .A(n18862), .B(n11100), .Z(n11111) );
  XNOR U19598 ( .A(q[7]), .B(DB[1087]), .Z(n11100) );
  IV U19599 ( .A(n11099), .Z(n18862) );
  XNOR U19600 ( .A(n11097), .B(n18863), .Z(n11099) );
  XNOR U19601 ( .A(q[6]), .B(DB[1086]), .Z(n18863) );
  XNOR U19602 ( .A(q[5]), .B(DB[1085]), .Z(n11097) );
  IV U19603 ( .A(n11110), .Z(n18860) );
  XOR U19604 ( .A(n18864), .B(n18865), .Z(n11110) );
  XNOR U19605 ( .A(n11106), .B(n11108), .Z(n18865) );
  XNOR U19606 ( .A(q[1]), .B(DB[1081]), .Z(n11108) );
  XNOR U19607 ( .A(q[4]), .B(DB[1084]), .Z(n11106) );
  IV U19608 ( .A(n11105), .Z(n18864) );
  XNOR U19609 ( .A(n11103), .B(n18866), .Z(n11105) );
  XNOR U19610 ( .A(q[3]), .B(DB[1083]), .Z(n18866) );
  XNOR U19611 ( .A(q[2]), .B(DB[1082]), .Z(n11103) );
  XOR U19612 ( .A(n18867), .B(n11001), .Z(n10929) );
  XOR U19613 ( .A(n18868), .B(n10993), .Z(n11001) );
  XOR U19614 ( .A(n18869), .B(n10982), .Z(n10993) );
  XNOR U19615 ( .A(q[14]), .B(DB[1109]), .Z(n10982) );
  IV U19616 ( .A(n10981), .Z(n18869) );
  XNOR U19617 ( .A(n10979), .B(n18870), .Z(n10981) );
  XNOR U19618 ( .A(q[13]), .B(DB[1108]), .Z(n18870) );
  XNOR U19619 ( .A(q[12]), .B(DB[1107]), .Z(n10979) );
  IV U19620 ( .A(n10992), .Z(n18868) );
  XOR U19621 ( .A(n18871), .B(n18872), .Z(n10992) );
  XNOR U19622 ( .A(n10988), .B(n10990), .Z(n18872) );
  XNOR U19623 ( .A(q[8]), .B(DB[1103]), .Z(n10990) );
  XNOR U19624 ( .A(q[11]), .B(DB[1106]), .Z(n10988) );
  IV U19625 ( .A(n10987), .Z(n18871) );
  XNOR U19626 ( .A(n10985), .B(n18873), .Z(n10987) );
  XNOR U19627 ( .A(q[10]), .B(DB[1105]), .Z(n18873) );
  XNOR U19628 ( .A(q[9]), .B(DB[1104]), .Z(n10985) );
  IV U19629 ( .A(n11000), .Z(n18867) );
  XOR U19630 ( .A(n18874), .B(n18875), .Z(n11000) );
  XNOR U19631 ( .A(n11017), .B(n10998), .Z(n18875) );
  XNOR U19632 ( .A(q[0]), .B(DB[1095]), .Z(n10998) );
  XOR U19633 ( .A(n18876), .B(n11006), .Z(n11017) );
  XNOR U19634 ( .A(q[7]), .B(DB[1102]), .Z(n11006) );
  IV U19635 ( .A(n11005), .Z(n18876) );
  XNOR U19636 ( .A(n11003), .B(n18877), .Z(n11005) );
  XNOR U19637 ( .A(q[6]), .B(DB[1101]), .Z(n18877) );
  XNOR U19638 ( .A(q[5]), .B(DB[1100]), .Z(n11003) );
  IV U19639 ( .A(n11016), .Z(n18874) );
  XOR U19640 ( .A(n18878), .B(n18879), .Z(n11016) );
  XNOR U19641 ( .A(n11012), .B(n11014), .Z(n18879) );
  XNOR U19642 ( .A(q[1]), .B(DB[1096]), .Z(n11014) );
  XNOR U19643 ( .A(q[4]), .B(DB[1099]), .Z(n11012) );
  IV U19644 ( .A(n11011), .Z(n18878) );
  XNOR U19645 ( .A(n11009), .B(n18880), .Z(n11011) );
  XNOR U19646 ( .A(q[3]), .B(DB[1098]), .Z(n18880) );
  XNOR U19647 ( .A(q[2]), .B(DB[1097]), .Z(n11009) );
  XOR U19648 ( .A(n18881), .B(n10907), .Z(n10835) );
  XOR U19649 ( .A(n18882), .B(n10899), .Z(n10907) );
  XOR U19650 ( .A(n18883), .B(n10888), .Z(n10899) );
  XNOR U19651 ( .A(q[14]), .B(DB[1124]), .Z(n10888) );
  IV U19652 ( .A(n10887), .Z(n18883) );
  XNOR U19653 ( .A(n10885), .B(n18884), .Z(n10887) );
  XNOR U19654 ( .A(q[13]), .B(DB[1123]), .Z(n18884) );
  XNOR U19655 ( .A(q[12]), .B(DB[1122]), .Z(n10885) );
  IV U19656 ( .A(n10898), .Z(n18882) );
  XOR U19657 ( .A(n18885), .B(n18886), .Z(n10898) );
  XNOR U19658 ( .A(n10894), .B(n10896), .Z(n18886) );
  XNOR U19659 ( .A(q[8]), .B(DB[1118]), .Z(n10896) );
  XNOR U19660 ( .A(q[11]), .B(DB[1121]), .Z(n10894) );
  IV U19661 ( .A(n10893), .Z(n18885) );
  XNOR U19662 ( .A(n10891), .B(n18887), .Z(n10893) );
  XNOR U19663 ( .A(q[10]), .B(DB[1120]), .Z(n18887) );
  XNOR U19664 ( .A(q[9]), .B(DB[1119]), .Z(n10891) );
  IV U19665 ( .A(n10906), .Z(n18881) );
  XOR U19666 ( .A(n18888), .B(n18889), .Z(n10906) );
  XNOR U19667 ( .A(n10923), .B(n10904), .Z(n18889) );
  XNOR U19668 ( .A(q[0]), .B(DB[1110]), .Z(n10904) );
  XOR U19669 ( .A(n18890), .B(n10912), .Z(n10923) );
  XNOR U19670 ( .A(q[7]), .B(DB[1117]), .Z(n10912) );
  IV U19671 ( .A(n10911), .Z(n18890) );
  XNOR U19672 ( .A(n10909), .B(n18891), .Z(n10911) );
  XNOR U19673 ( .A(q[6]), .B(DB[1116]), .Z(n18891) );
  XNOR U19674 ( .A(q[5]), .B(DB[1115]), .Z(n10909) );
  IV U19675 ( .A(n10922), .Z(n18888) );
  XOR U19676 ( .A(n18892), .B(n18893), .Z(n10922) );
  XNOR U19677 ( .A(n10918), .B(n10920), .Z(n18893) );
  XNOR U19678 ( .A(q[1]), .B(DB[1111]), .Z(n10920) );
  XNOR U19679 ( .A(q[4]), .B(DB[1114]), .Z(n10918) );
  IV U19680 ( .A(n10917), .Z(n18892) );
  XNOR U19681 ( .A(n10915), .B(n18894), .Z(n10917) );
  XNOR U19682 ( .A(q[3]), .B(DB[1113]), .Z(n18894) );
  XNOR U19683 ( .A(q[2]), .B(DB[1112]), .Z(n10915) );
  XOR U19684 ( .A(n18895), .B(n10813), .Z(n10741) );
  XOR U19685 ( .A(n18896), .B(n10805), .Z(n10813) );
  XOR U19686 ( .A(n18897), .B(n10794), .Z(n10805) );
  XNOR U19687 ( .A(q[14]), .B(DB[1139]), .Z(n10794) );
  IV U19688 ( .A(n10793), .Z(n18897) );
  XNOR U19689 ( .A(n10791), .B(n18898), .Z(n10793) );
  XNOR U19690 ( .A(q[13]), .B(DB[1138]), .Z(n18898) );
  XNOR U19691 ( .A(q[12]), .B(DB[1137]), .Z(n10791) );
  IV U19692 ( .A(n10804), .Z(n18896) );
  XOR U19693 ( .A(n18899), .B(n18900), .Z(n10804) );
  XNOR U19694 ( .A(n10800), .B(n10802), .Z(n18900) );
  XNOR U19695 ( .A(q[8]), .B(DB[1133]), .Z(n10802) );
  XNOR U19696 ( .A(q[11]), .B(DB[1136]), .Z(n10800) );
  IV U19697 ( .A(n10799), .Z(n18899) );
  XNOR U19698 ( .A(n10797), .B(n18901), .Z(n10799) );
  XNOR U19699 ( .A(q[10]), .B(DB[1135]), .Z(n18901) );
  XNOR U19700 ( .A(q[9]), .B(DB[1134]), .Z(n10797) );
  IV U19701 ( .A(n10812), .Z(n18895) );
  XOR U19702 ( .A(n18902), .B(n18903), .Z(n10812) );
  XNOR U19703 ( .A(n10829), .B(n10810), .Z(n18903) );
  XNOR U19704 ( .A(q[0]), .B(DB[1125]), .Z(n10810) );
  XOR U19705 ( .A(n18904), .B(n10818), .Z(n10829) );
  XNOR U19706 ( .A(q[7]), .B(DB[1132]), .Z(n10818) );
  IV U19707 ( .A(n10817), .Z(n18904) );
  XNOR U19708 ( .A(n10815), .B(n18905), .Z(n10817) );
  XNOR U19709 ( .A(q[6]), .B(DB[1131]), .Z(n18905) );
  XNOR U19710 ( .A(q[5]), .B(DB[1130]), .Z(n10815) );
  IV U19711 ( .A(n10828), .Z(n18902) );
  XOR U19712 ( .A(n18906), .B(n18907), .Z(n10828) );
  XNOR U19713 ( .A(n10824), .B(n10826), .Z(n18907) );
  XNOR U19714 ( .A(q[1]), .B(DB[1126]), .Z(n10826) );
  XNOR U19715 ( .A(q[4]), .B(DB[1129]), .Z(n10824) );
  IV U19716 ( .A(n10823), .Z(n18906) );
  XNOR U19717 ( .A(n10821), .B(n18908), .Z(n10823) );
  XNOR U19718 ( .A(q[3]), .B(DB[1128]), .Z(n18908) );
  XNOR U19719 ( .A(q[2]), .B(DB[1127]), .Z(n10821) );
  XOR U19720 ( .A(n18909), .B(n10719), .Z(n10647) );
  XOR U19721 ( .A(n18910), .B(n10711), .Z(n10719) );
  XOR U19722 ( .A(n18911), .B(n10700), .Z(n10711) );
  XNOR U19723 ( .A(q[14]), .B(DB[1154]), .Z(n10700) );
  IV U19724 ( .A(n10699), .Z(n18911) );
  XNOR U19725 ( .A(n10697), .B(n18912), .Z(n10699) );
  XNOR U19726 ( .A(q[13]), .B(DB[1153]), .Z(n18912) );
  XNOR U19727 ( .A(q[12]), .B(DB[1152]), .Z(n10697) );
  IV U19728 ( .A(n10710), .Z(n18910) );
  XOR U19729 ( .A(n18913), .B(n18914), .Z(n10710) );
  XNOR U19730 ( .A(n10706), .B(n10708), .Z(n18914) );
  XNOR U19731 ( .A(q[8]), .B(DB[1148]), .Z(n10708) );
  XNOR U19732 ( .A(q[11]), .B(DB[1151]), .Z(n10706) );
  IV U19733 ( .A(n10705), .Z(n18913) );
  XNOR U19734 ( .A(n10703), .B(n18915), .Z(n10705) );
  XNOR U19735 ( .A(q[10]), .B(DB[1150]), .Z(n18915) );
  XNOR U19736 ( .A(q[9]), .B(DB[1149]), .Z(n10703) );
  IV U19737 ( .A(n10718), .Z(n18909) );
  XOR U19738 ( .A(n18916), .B(n18917), .Z(n10718) );
  XNOR U19739 ( .A(n10735), .B(n10716), .Z(n18917) );
  XNOR U19740 ( .A(q[0]), .B(DB[1140]), .Z(n10716) );
  XOR U19741 ( .A(n18918), .B(n10724), .Z(n10735) );
  XNOR U19742 ( .A(q[7]), .B(DB[1147]), .Z(n10724) );
  IV U19743 ( .A(n10723), .Z(n18918) );
  XNOR U19744 ( .A(n10721), .B(n18919), .Z(n10723) );
  XNOR U19745 ( .A(q[6]), .B(DB[1146]), .Z(n18919) );
  XNOR U19746 ( .A(q[5]), .B(DB[1145]), .Z(n10721) );
  IV U19747 ( .A(n10734), .Z(n18916) );
  XOR U19748 ( .A(n18920), .B(n18921), .Z(n10734) );
  XNOR U19749 ( .A(n10730), .B(n10732), .Z(n18921) );
  XNOR U19750 ( .A(q[1]), .B(DB[1141]), .Z(n10732) );
  XNOR U19751 ( .A(q[4]), .B(DB[1144]), .Z(n10730) );
  IV U19752 ( .A(n10729), .Z(n18920) );
  XNOR U19753 ( .A(n10727), .B(n18922), .Z(n10729) );
  XNOR U19754 ( .A(q[3]), .B(DB[1143]), .Z(n18922) );
  XNOR U19755 ( .A(q[2]), .B(DB[1142]), .Z(n10727) );
  XOR U19756 ( .A(n18923), .B(n10625), .Z(n10553) );
  XOR U19757 ( .A(n18924), .B(n10617), .Z(n10625) );
  XOR U19758 ( .A(n18925), .B(n10606), .Z(n10617) );
  XNOR U19759 ( .A(q[14]), .B(DB[1169]), .Z(n10606) );
  IV U19760 ( .A(n10605), .Z(n18925) );
  XNOR U19761 ( .A(n10603), .B(n18926), .Z(n10605) );
  XNOR U19762 ( .A(q[13]), .B(DB[1168]), .Z(n18926) );
  XNOR U19763 ( .A(q[12]), .B(DB[1167]), .Z(n10603) );
  IV U19764 ( .A(n10616), .Z(n18924) );
  XOR U19765 ( .A(n18927), .B(n18928), .Z(n10616) );
  XNOR U19766 ( .A(n10612), .B(n10614), .Z(n18928) );
  XNOR U19767 ( .A(q[8]), .B(DB[1163]), .Z(n10614) );
  XNOR U19768 ( .A(q[11]), .B(DB[1166]), .Z(n10612) );
  IV U19769 ( .A(n10611), .Z(n18927) );
  XNOR U19770 ( .A(n10609), .B(n18929), .Z(n10611) );
  XNOR U19771 ( .A(q[10]), .B(DB[1165]), .Z(n18929) );
  XNOR U19772 ( .A(q[9]), .B(DB[1164]), .Z(n10609) );
  IV U19773 ( .A(n10624), .Z(n18923) );
  XOR U19774 ( .A(n18930), .B(n18931), .Z(n10624) );
  XNOR U19775 ( .A(n10641), .B(n10622), .Z(n18931) );
  XNOR U19776 ( .A(q[0]), .B(DB[1155]), .Z(n10622) );
  XOR U19777 ( .A(n18932), .B(n10630), .Z(n10641) );
  XNOR U19778 ( .A(q[7]), .B(DB[1162]), .Z(n10630) );
  IV U19779 ( .A(n10629), .Z(n18932) );
  XNOR U19780 ( .A(n10627), .B(n18933), .Z(n10629) );
  XNOR U19781 ( .A(q[6]), .B(DB[1161]), .Z(n18933) );
  XNOR U19782 ( .A(q[5]), .B(DB[1160]), .Z(n10627) );
  IV U19783 ( .A(n10640), .Z(n18930) );
  XOR U19784 ( .A(n18934), .B(n18935), .Z(n10640) );
  XNOR U19785 ( .A(n10636), .B(n10638), .Z(n18935) );
  XNOR U19786 ( .A(q[1]), .B(DB[1156]), .Z(n10638) );
  XNOR U19787 ( .A(q[4]), .B(DB[1159]), .Z(n10636) );
  IV U19788 ( .A(n10635), .Z(n18934) );
  XNOR U19789 ( .A(n10633), .B(n18936), .Z(n10635) );
  XNOR U19790 ( .A(q[3]), .B(DB[1158]), .Z(n18936) );
  XNOR U19791 ( .A(q[2]), .B(DB[1157]), .Z(n10633) );
  XOR U19792 ( .A(n18937), .B(n10531), .Z(n10459) );
  XOR U19793 ( .A(n18938), .B(n10523), .Z(n10531) );
  XOR U19794 ( .A(n18939), .B(n10512), .Z(n10523) );
  XNOR U19795 ( .A(q[14]), .B(DB[1184]), .Z(n10512) );
  IV U19796 ( .A(n10511), .Z(n18939) );
  XNOR U19797 ( .A(n10509), .B(n18940), .Z(n10511) );
  XNOR U19798 ( .A(q[13]), .B(DB[1183]), .Z(n18940) );
  XNOR U19799 ( .A(q[12]), .B(DB[1182]), .Z(n10509) );
  IV U19800 ( .A(n10522), .Z(n18938) );
  XOR U19801 ( .A(n18941), .B(n18942), .Z(n10522) );
  XNOR U19802 ( .A(n10518), .B(n10520), .Z(n18942) );
  XNOR U19803 ( .A(q[8]), .B(DB[1178]), .Z(n10520) );
  XNOR U19804 ( .A(q[11]), .B(DB[1181]), .Z(n10518) );
  IV U19805 ( .A(n10517), .Z(n18941) );
  XNOR U19806 ( .A(n10515), .B(n18943), .Z(n10517) );
  XNOR U19807 ( .A(q[10]), .B(DB[1180]), .Z(n18943) );
  XNOR U19808 ( .A(q[9]), .B(DB[1179]), .Z(n10515) );
  IV U19809 ( .A(n10530), .Z(n18937) );
  XOR U19810 ( .A(n18944), .B(n18945), .Z(n10530) );
  XNOR U19811 ( .A(n10547), .B(n10528), .Z(n18945) );
  XNOR U19812 ( .A(q[0]), .B(DB[1170]), .Z(n10528) );
  XOR U19813 ( .A(n18946), .B(n10536), .Z(n10547) );
  XNOR U19814 ( .A(q[7]), .B(DB[1177]), .Z(n10536) );
  IV U19815 ( .A(n10535), .Z(n18946) );
  XNOR U19816 ( .A(n10533), .B(n18947), .Z(n10535) );
  XNOR U19817 ( .A(q[6]), .B(DB[1176]), .Z(n18947) );
  XNOR U19818 ( .A(q[5]), .B(DB[1175]), .Z(n10533) );
  IV U19819 ( .A(n10546), .Z(n18944) );
  XOR U19820 ( .A(n18948), .B(n18949), .Z(n10546) );
  XNOR U19821 ( .A(n10542), .B(n10544), .Z(n18949) );
  XNOR U19822 ( .A(q[1]), .B(DB[1171]), .Z(n10544) );
  XNOR U19823 ( .A(q[4]), .B(DB[1174]), .Z(n10542) );
  IV U19824 ( .A(n10541), .Z(n18948) );
  XNOR U19825 ( .A(n10539), .B(n18950), .Z(n10541) );
  XNOR U19826 ( .A(q[3]), .B(DB[1173]), .Z(n18950) );
  XNOR U19827 ( .A(q[2]), .B(DB[1172]), .Z(n10539) );
  XOR U19828 ( .A(n18951), .B(n10437), .Z(n10365) );
  XOR U19829 ( .A(n18952), .B(n10429), .Z(n10437) );
  XOR U19830 ( .A(n18953), .B(n10418), .Z(n10429) );
  XNOR U19831 ( .A(q[14]), .B(DB[1199]), .Z(n10418) );
  IV U19832 ( .A(n10417), .Z(n18953) );
  XNOR U19833 ( .A(n10415), .B(n18954), .Z(n10417) );
  XNOR U19834 ( .A(q[13]), .B(DB[1198]), .Z(n18954) );
  XNOR U19835 ( .A(q[12]), .B(DB[1197]), .Z(n10415) );
  IV U19836 ( .A(n10428), .Z(n18952) );
  XOR U19837 ( .A(n18955), .B(n18956), .Z(n10428) );
  XNOR U19838 ( .A(n10424), .B(n10426), .Z(n18956) );
  XNOR U19839 ( .A(q[8]), .B(DB[1193]), .Z(n10426) );
  XNOR U19840 ( .A(q[11]), .B(DB[1196]), .Z(n10424) );
  IV U19841 ( .A(n10423), .Z(n18955) );
  XNOR U19842 ( .A(n10421), .B(n18957), .Z(n10423) );
  XNOR U19843 ( .A(q[10]), .B(DB[1195]), .Z(n18957) );
  XNOR U19844 ( .A(q[9]), .B(DB[1194]), .Z(n10421) );
  IV U19845 ( .A(n10436), .Z(n18951) );
  XOR U19846 ( .A(n18958), .B(n18959), .Z(n10436) );
  XNOR U19847 ( .A(n10453), .B(n10434), .Z(n18959) );
  XNOR U19848 ( .A(q[0]), .B(DB[1185]), .Z(n10434) );
  XOR U19849 ( .A(n18960), .B(n10442), .Z(n10453) );
  XNOR U19850 ( .A(q[7]), .B(DB[1192]), .Z(n10442) );
  IV U19851 ( .A(n10441), .Z(n18960) );
  XNOR U19852 ( .A(n10439), .B(n18961), .Z(n10441) );
  XNOR U19853 ( .A(q[6]), .B(DB[1191]), .Z(n18961) );
  XNOR U19854 ( .A(q[5]), .B(DB[1190]), .Z(n10439) );
  IV U19855 ( .A(n10452), .Z(n18958) );
  XOR U19856 ( .A(n18962), .B(n18963), .Z(n10452) );
  XNOR U19857 ( .A(n10448), .B(n10450), .Z(n18963) );
  XNOR U19858 ( .A(q[1]), .B(DB[1186]), .Z(n10450) );
  XNOR U19859 ( .A(q[4]), .B(DB[1189]), .Z(n10448) );
  IV U19860 ( .A(n10447), .Z(n18962) );
  XNOR U19861 ( .A(n10445), .B(n18964), .Z(n10447) );
  XNOR U19862 ( .A(q[3]), .B(DB[1188]), .Z(n18964) );
  XNOR U19863 ( .A(q[2]), .B(DB[1187]), .Z(n10445) );
  XOR U19864 ( .A(n18965), .B(n10343), .Z(n10271) );
  XOR U19865 ( .A(n18966), .B(n10335), .Z(n10343) );
  XOR U19866 ( .A(n18967), .B(n10324), .Z(n10335) );
  XNOR U19867 ( .A(q[14]), .B(DB[1214]), .Z(n10324) );
  IV U19868 ( .A(n10323), .Z(n18967) );
  XNOR U19869 ( .A(n10321), .B(n18968), .Z(n10323) );
  XNOR U19870 ( .A(q[13]), .B(DB[1213]), .Z(n18968) );
  XNOR U19871 ( .A(q[12]), .B(DB[1212]), .Z(n10321) );
  IV U19872 ( .A(n10334), .Z(n18966) );
  XOR U19873 ( .A(n18969), .B(n18970), .Z(n10334) );
  XNOR U19874 ( .A(n10330), .B(n10332), .Z(n18970) );
  XNOR U19875 ( .A(q[8]), .B(DB[1208]), .Z(n10332) );
  XNOR U19876 ( .A(q[11]), .B(DB[1211]), .Z(n10330) );
  IV U19877 ( .A(n10329), .Z(n18969) );
  XNOR U19878 ( .A(n10327), .B(n18971), .Z(n10329) );
  XNOR U19879 ( .A(q[10]), .B(DB[1210]), .Z(n18971) );
  XNOR U19880 ( .A(q[9]), .B(DB[1209]), .Z(n10327) );
  IV U19881 ( .A(n10342), .Z(n18965) );
  XOR U19882 ( .A(n18972), .B(n18973), .Z(n10342) );
  XNOR U19883 ( .A(n10359), .B(n10340), .Z(n18973) );
  XNOR U19884 ( .A(q[0]), .B(DB[1200]), .Z(n10340) );
  XOR U19885 ( .A(n18974), .B(n10348), .Z(n10359) );
  XNOR U19886 ( .A(q[7]), .B(DB[1207]), .Z(n10348) );
  IV U19887 ( .A(n10347), .Z(n18974) );
  XNOR U19888 ( .A(n10345), .B(n18975), .Z(n10347) );
  XNOR U19889 ( .A(q[6]), .B(DB[1206]), .Z(n18975) );
  XNOR U19890 ( .A(q[5]), .B(DB[1205]), .Z(n10345) );
  IV U19891 ( .A(n10358), .Z(n18972) );
  XOR U19892 ( .A(n18976), .B(n18977), .Z(n10358) );
  XNOR U19893 ( .A(n10354), .B(n10356), .Z(n18977) );
  XNOR U19894 ( .A(q[1]), .B(DB[1201]), .Z(n10356) );
  XNOR U19895 ( .A(q[4]), .B(DB[1204]), .Z(n10354) );
  IV U19896 ( .A(n10353), .Z(n18976) );
  XNOR U19897 ( .A(n10351), .B(n18978), .Z(n10353) );
  XNOR U19898 ( .A(q[3]), .B(DB[1203]), .Z(n18978) );
  XNOR U19899 ( .A(q[2]), .B(DB[1202]), .Z(n10351) );
  XOR U19900 ( .A(n18979), .B(n10249), .Z(n10177) );
  XOR U19901 ( .A(n18980), .B(n10241), .Z(n10249) );
  XOR U19902 ( .A(n18981), .B(n10230), .Z(n10241) );
  XNOR U19903 ( .A(q[14]), .B(DB[1229]), .Z(n10230) );
  IV U19904 ( .A(n10229), .Z(n18981) );
  XNOR U19905 ( .A(n10227), .B(n18982), .Z(n10229) );
  XNOR U19906 ( .A(q[13]), .B(DB[1228]), .Z(n18982) );
  XNOR U19907 ( .A(q[12]), .B(DB[1227]), .Z(n10227) );
  IV U19908 ( .A(n10240), .Z(n18980) );
  XOR U19909 ( .A(n18983), .B(n18984), .Z(n10240) );
  XNOR U19910 ( .A(n10236), .B(n10238), .Z(n18984) );
  XNOR U19911 ( .A(q[8]), .B(DB[1223]), .Z(n10238) );
  XNOR U19912 ( .A(q[11]), .B(DB[1226]), .Z(n10236) );
  IV U19913 ( .A(n10235), .Z(n18983) );
  XNOR U19914 ( .A(n10233), .B(n18985), .Z(n10235) );
  XNOR U19915 ( .A(q[10]), .B(DB[1225]), .Z(n18985) );
  XNOR U19916 ( .A(q[9]), .B(DB[1224]), .Z(n10233) );
  IV U19917 ( .A(n10248), .Z(n18979) );
  XOR U19918 ( .A(n18986), .B(n18987), .Z(n10248) );
  XNOR U19919 ( .A(n10265), .B(n10246), .Z(n18987) );
  XNOR U19920 ( .A(q[0]), .B(DB[1215]), .Z(n10246) );
  XOR U19921 ( .A(n18988), .B(n10254), .Z(n10265) );
  XNOR U19922 ( .A(q[7]), .B(DB[1222]), .Z(n10254) );
  IV U19923 ( .A(n10253), .Z(n18988) );
  XNOR U19924 ( .A(n10251), .B(n18989), .Z(n10253) );
  XNOR U19925 ( .A(q[6]), .B(DB[1221]), .Z(n18989) );
  XNOR U19926 ( .A(q[5]), .B(DB[1220]), .Z(n10251) );
  IV U19927 ( .A(n10264), .Z(n18986) );
  XOR U19928 ( .A(n18990), .B(n18991), .Z(n10264) );
  XNOR U19929 ( .A(n10260), .B(n10262), .Z(n18991) );
  XNOR U19930 ( .A(q[1]), .B(DB[1216]), .Z(n10262) );
  XNOR U19931 ( .A(q[4]), .B(DB[1219]), .Z(n10260) );
  IV U19932 ( .A(n10259), .Z(n18990) );
  XNOR U19933 ( .A(n10257), .B(n18992), .Z(n10259) );
  XNOR U19934 ( .A(q[3]), .B(DB[1218]), .Z(n18992) );
  XNOR U19935 ( .A(q[2]), .B(DB[1217]), .Z(n10257) );
  XOR U19936 ( .A(n18993), .B(n10155), .Z(n10083) );
  XOR U19937 ( .A(n18994), .B(n10147), .Z(n10155) );
  XOR U19938 ( .A(n18995), .B(n10136), .Z(n10147) );
  XNOR U19939 ( .A(q[14]), .B(DB[1244]), .Z(n10136) );
  IV U19940 ( .A(n10135), .Z(n18995) );
  XNOR U19941 ( .A(n10133), .B(n18996), .Z(n10135) );
  XNOR U19942 ( .A(q[13]), .B(DB[1243]), .Z(n18996) );
  XNOR U19943 ( .A(q[12]), .B(DB[1242]), .Z(n10133) );
  IV U19944 ( .A(n10146), .Z(n18994) );
  XOR U19945 ( .A(n18997), .B(n18998), .Z(n10146) );
  XNOR U19946 ( .A(n10142), .B(n10144), .Z(n18998) );
  XNOR U19947 ( .A(q[8]), .B(DB[1238]), .Z(n10144) );
  XNOR U19948 ( .A(q[11]), .B(DB[1241]), .Z(n10142) );
  IV U19949 ( .A(n10141), .Z(n18997) );
  XNOR U19950 ( .A(n10139), .B(n18999), .Z(n10141) );
  XNOR U19951 ( .A(q[10]), .B(DB[1240]), .Z(n18999) );
  XNOR U19952 ( .A(q[9]), .B(DB[1239]), .Z(n10139) );
  IV U19953 ( .A(n10154), .Z(n18993) );
  XOR U19954 ( .A(n19000), .B(n19001), .Z(n10154) );
  XNOR U19955 ( .A(n10171), .B(n10152), .Z(n19001) );
  XNOR U19956 ( .A(q[0]), .B(DB[1230]), .Z(n10152) );
  XOR U19957 ( .A(n19002), .B(n10160), .Z(n10171) );
  XNOR U19958 ( .A(q[7]), .B(DB[1237]), .Z(n10160) );
  IV U19959 ( .A(n10159), .Z(n19002) );
  XNOR U19960 ( .A(n10157), .B(n19003), .Z(n10159) );
  XNOR U19961 ( .A(q[6]), .B(DB[1236]), .Z(n19003) );
  XNOR U19962 ( .A(q[5]), .B(DB[1235]), .Z(n10157) );
  IV U19963 ( .A(n10170), .Z(n19000) );
  XOR U19964 ( .A(n19004), .B(n19005), .Z(n10170) );
  XNOR U19965 ( .A(n10166), .B(n10168), .Z(n19005) );
  XNOR U19966 ( .A(q[1]), .B(DB[1231]), .Z(n10168) );
  XNOR U19967 ( .A(q[4]), .B(DB[1234]), .Z(n10166) );
  IV U19968 ( .A(n10165), .Z(n19004) );
  XNOR U19969 ( .A(n10163), .B(n19006), .Z(n10165) );
  XNOR U19970 ( .A(q[3]), .B(DB[1233]), .Z(n19006) );
  XNOR U19971 ( .A(q[2]), .B(DB[1232]), .Z(n10163) );
  XOR U19972 ( .A(n19007), .B(n10061), .Z(n9989) );
  XOR U19973 ( .A(n19008), .B(n10053), .Z(n10061) );
  XOR U19974 ( .A(n19009), .B(n10042), .Z(n10053) );
  XNOR U19975 ( .A(q[14]), .B(DB[1259]), .Z(n10042) );
  IV U19976 ( .A(n10041), .Z(n19009) );
  XNOR U19977 ( .A(n10039), .B(n19010), .Z(n10041) );
  XNOR U19978 ( .A(q[13]), .B(DB[1258]), .Z(n19010) );
  XNOR U19979 ( .A(q[12]), .B(DB[1257]), .Z(n10039) );
  IV U19980 ( .A(n10052), .Z(n19008) );
  XOR U19981 ( .A(n19011), .B(n19012), .Z(n10052) );
  XNOR U19982 ( .A(n10048), .B(n10050), .Z(n19012) );
  XNOR U19983 ( .A(q[8]), .B(DB[1253]), .Z(n10050) );
  XNOR U19984 ( .A(q[11]), .B(DB[1256]), .Z(n10048) );
  IV U19985 ( .A(n10047), .Z(n19011) );
  XNOR U19986 ( .A(n10045), .B(n19013), .Z(n10047) );
  XNOR U19987 ( .A(q[10]), .B(DB[1255]), .Z(n19013) );
  XNOR U19988 ( .A(q[9]), .B(DB[1254]), .Z(n10045) );
  IV U19989 ( .A(n10060), .Z(n19007) );
  XOR U19990 ( .A(n19014), .B(n19015), .Z(n10060) );
  XNOR U19991 ( .A(n10077), .B(n10058), .Z(n19015) );
  XNOR U19992 ( .A(q[0]), .B(DB[1245]), .Z(n10058) );
  XOR U19993 ( .A(n19016), .B(n10066), .Z(n10077) );
  XNOR U19994 ( .A(q[7]), .B(DB[1252]), .Z(n10066) );
  IV U19995 ( .A(n10065), .Z(n19016) );
  XNOR U19996 ( .A(n10063), .B(n19017), .Z(n10065) );
  XNOR U19997 ( .A(q[6]), .B(DB[1251]), .Z(n19017) );
  XNOR U19998 ( .A(q[5]), .B(DB[1250]), .Z(n10063) );
  IV U19999 ( .A(n10076), .Z(n19014) );
  XOR U20000 ( .A(n19018), .B(n19019), .Z(n10076) );
  XNOR U20001 ( .A(n10072), .B(n10074), .Z(n19019) );
  XNOR U20002 ( .A(q[1]), .B(DB[1246]), .Z(n10074) );
  XNOR U20003 ( .A(q[4]), .B(DB[1249]), .Z(n10072) );
  IV U20004 ( .A(n10071), .Z(n19018) );
  XNOR U20005 ( .A(n10069), .B(n19020), .Z(n10071) );
  XNOR U20006 ( .A(q[3]), .B(DB[1248]), .Z(n19020) );
  XNOR U20007 ( .A(q[2]), .B(DB[1247]), .Z(n10069) );
  XOR U20008 ( .A(n19021), .B(n9967), .Z(n9895) );
  XOR U20009 ( .A(n19022), .B(n9959), .Z(n9967) );
  XOR U20010 ( .A(n19023), .B(n9948), .Z(n9959) );
  XNOR U20011 ( .A(q[14]), .B(DB[1274]), .Z(n9948) );
  IV U20012 ( .A(n9947), .Z(n19023) );
  XNOR U20013 ( .A(n9945), .B(n19024), .Z(n9947) );
  XNOR U20014 ( .A(q[13]), .B(DB[1273]), .Z(n19024) );
  XNOR U20015 ( .A(q[12]), .B(DB[1272]), .Z(n9945) );
  IV U20016 ( .A(n9958), .Z(n19022) );
  XOR U20017 ( .A(n19025), .B(n19026), .Z(n9958) );
  XNOR U20018 ( .A(n9954), .B(n9956), .Z(n19026) );
  XNOR U20019 ( .A(q[8]), .B(DB[1268]), .Z(n9956) );
  XNOR U20020 ( .A(q[11]), .B(DB[1271]), .Z(n9954) );
  IV U20021 ( .A(n9953), .Z(n19025) );
  XNOR U20022 ( .A(n9951), .B(n19027), .Z(n9953) );
  XNOR U20023 ( .A(q[10]), .B(DB[1270]), .Z(n19027) );
  XNOR U20024 ( .A(q[9]), .B(DB[1269]), .Z(n9951) );
  IV U20025 ( .A(n9966), .Z(n19021) );
  XOR U20026 ( .A(n19028), .B(n19029), .Z(n9966) );
  XNOR U20027 ( .A(n9983), .B(n9964), .Z(n19029) );
  XNOR U20028 ( .A(q[0]), .B(DB[1260]), .Z(n9964) );
  XOR U20029 ( .A(n19030), .B(n9972), .Z(n9983) );
  XNOR U20030 ( .A(q[7]), .B(DB[1267]), .Z(n9972) );
  IV U20031 ( .A(n9971), .Z(n19030) );
  XNOR U20032 ( .A(n9969), .B(n19031), .Z(n9971) );
  XNOR U20033 ( .A(q[6]), .B(DB[1266]), .Z(n19031) );
  XNOR U20034 ( .A(q[5]), .B(DB[1265]), .Z(n9969) );
  IV U20035 ( .A(n9982), .Z(n19028) );
  XOR U20036 ( .A(n19032), .B(n19033), .Z(n9982) );
  XNOR U20037 ( .A(n9978), .B(n9980), .Z(n19033) );
  XNOR U20038 ( .A(q[1]), .B(DB[1261]), .Z(n9980) );
  XNOR U20039 ( .A(q[4]), .B(DB[1264]), .Z(n9978) );
  IV U20040 ( .A(n9977), .Z(n19032) );
  XNOR U20041 ( .A(n9975), .B(n19034), .Z(n9977) );
  XNOR U20042 ( .A(q[3]), .B(DB[1263]), .Z(n19034) );
  XNOR U20043 ( .A(q[2]), .B(DB[1262]), .Z(n9975) );
  XOR U20044 ( .A(n19035), .B(n9873), .Z(n9801) );
  XOR U20045 ( .A(n19036), .B(n9865), .Z(n9873) );
  XOR U20046 ( .A(n19037), .B(n9854), .Z(n9865) );
  XNOR U20047 ( .A(q[14]), .B(DB[1289]), .Z(n9854) );
  IV U20048 ( .A(n9853), .Z(n19037) );
  XNOR U20049 ( .A(n9851), .B(n19038), .Z(n9853) );
  XNOR U20050 ( .A(q[13]), .B(DB[1288]), .Z(n19038) );
  XNOR U20051 ( .A(q[12]), .B(DB[1287]), .Z(n9851) );
  IV U20052 ( .A(n9864), .Z(n19036) );
  XOR U20053 ( .A(n19039), .B(n19040), .Z(n9864) );
  XNOR U20054 ( .A(n9860), .B(n9862), .Z(n19040) );
  XNOR U20055 ( .A(q[8]), .B(DB[1283]), .Z(n9862) );
  XNOR U20056 ( .A(q[11]), .B(DB[1286]), .Z(n9860) );
  IV U20057 ( .A(n9859), .Z(n19039) );
  XNOR U20058 ( .A(n9857), .B(n19041), .Z(n9859) );
  XNOR U20059 ( .A(q[10]), .B(DB[1285]), .Z(n19041) );
  XNOR U20060 ( .A(q[9]), .B(DB[1284]), .Z(n9857) );
  IV U20061 ( .A(n9872), .Z(n19035) );
  XOR U20062 ( .A(n19042), .B(n19043), .Z(n9872) );
  XNOR U20063 ( .A(n9889), .B(n9870), .Z(n19043) );
  XNOR U20064 ( .A(q[0]), .B(DB[1275]), .Z(n9870) );
  XOR U20065 ( .A(n19044), .B(n9878), .Z(n9889) );
  XNOR U20066 ( .A(q[7]), .B(DB[1282]), .Z(n9878) );
  IV U20067 ( .A(n9877), .Z(n19044) );
  XNOR U20068 ( .A(n9875), .B(n19045), .Z(n9877) );
  XNOR U20069 ( .A(q[6]), .B(DB[1281]), .Z(n19045) );
  XNOR U20070 ( .A(q[5]), .B(DB[1280]), .Z(n9875) );
  IV U20071 ( .A(n9888), .Z(n19042) );
  XOR U20072 ( .A(n19046), .B(n19047), .Z(n9888) );
  XNOR U20073 ( .A(n9884), .B(n9886), .Z(n19047) );
  XNOR U20074 ( .A(q[1]), .B(DB[1276]), .Z(n9886) );
  XNOR U20075 ( .A(q[4]), .B(DB[1279]), .Z(n9884) );
  IV U20076 ( .A(n9883), .Z(n19046) );
  XNOR U20077 ( .A(n9881), .B(n19048), .Z(n9883) );
  XNOR U20078 ( .A(q[3]), .B(DB[1278]), .Z(n19048) );
  XNOR U20079 ( .A(q[2]), .B(DB[1277]), .Z(n9881) );
  XOR U20080 ( .A(n19049), .B(n9779), .Z(n9707) );
  XOR U20081 ( .A(n19050), .B(n9771), .Z(n9779) );
  XOR U20082 ( .A(n19051), .B(n9760), .Z(n9771) );
  XNOR U20083 ( .A(q[14]), .B(DB[1304]), .Z(n9760) );
  IV U20084 ( .A(n9759), .Z(n19051) );
  XNOR U20085 ( .A(n9757), .B(n19052), .Z(n9759) );
  XNOR U20086 ( .A(q[13]), .B(DB[1303]), .Z(n19052) );
  XNOR U20087 ( .A(q[12]), .B(DB[1302]), .Z(n9757) );
  IV U20088 ( .A(n9770), .Z(n19050) );
  XOR U20089 ( .A(n19053), .B(n19054), .Z(n9770) );
  XNOR U20090 ( .A(n9766), .B(n9768), .Z(n19054) );
  XNOR U20091 ( .A(q[8]), .B(DB[1298]), .Z(n9768) );
  XNOR U20092 ( .A(q[11]), .B(DB[1301]), .Z(n9766) );
  IV U20093 ( .A(n9765), .Z(n19053) );
  XNOR U20094 ( .A(n9763), .B(n19055), .Z(n9765) );
  XNOR U20095 ( .A(q[10]), .B(DB[1300]), .Z(n19055) );
  XNOR U20096 ( .A(q[9]), .B(DB[1299]), .Z(n9763) );
  IV U20097 ( .A(n9778), .Z(n19049) );
  XOR U20098 ( .A(n19056), .B(n19057), .Z(n9778) );
  XNOR U20099 ( .A(n9795), .B(n9776), .Z(n19057) );
  XNOR U20100 ( .A(q[0]), .B(DB[1290]), .Z(n9776) );
  XOR U20101 ( .A(n19058), .B(n9784), .Z(n9795) );
  XNOR U20102 ( .A(q[7]), .B(DB[1297]), .Z(n9784) );
  IV U20103 ( .A(n9783), .Z(n19058) );
  XNOR U20104 ( .A(n9781), .B(n19059), .Z(n9783) );
  XNOR U20105 ( .A(q[6]), .B(DB[1296]), .Z(n19059) );
  XNOR U20106 ( .A(q[5]), .B(DB[1295]), .Z(n9781) );
  IV U20107 ( .A(n9794), .Z(n19056) );
  XOR U20108 ( .A(n19060), .B(n19061), .Z(n9794) );
  XNOR U20109 ( .A(n9790), .B(n9792), .Z(n19061) );
  XNOR U20110 ( .A(q[1]), .B(DB[1291]), .Z(n9792) );
  XNOR U20111 ( .A(q[4]), .B(DB[1294]), .Z(n9790) );
  IV U20112 ( .A(n9789), .Z(n19060) );
  XNOR U20113 ( .A(n9787), .B(n19062), .Z(n9789) );
  XNOR U20114 ( .A(q[3]), .B(DB[1293]), .Z(n19062) );
  XNOR U20115 ( .A(q[2]), .B(DB[1292]), .Z(n9787) );
  XOR U20116 ( .A(n19063), .B(n9685), .Z(n9613) );
  XOR U20117 ( .A(n19064), .B(n9677), .Z(n9685) );
  XOR U20118 ( .A(n19065), .B(n9666), .Z(n9677) );
  XNOR U20119 ( .A(q[14]), .B(DB[1319]), .Z(n9666) );
  IV U20120 ( .A(n9665), .Z(n19065) );
  XNOR U20121 ( .A(n9663), .B(n19066), .Z(n9665) );
  XNOR U20122 ( .A(q[13]), .B(DB[1318]), .Z(n19066) );
  XNOR U20123 ( .A(q[12]), .B(DB[1317]), .Z(n9663) );
  IV U20124 ( .A(n9676), .Z(n19064) );
  XOR U20125 ( .A(n19067), .B(n19068), .Z(n9676) );
  XNOR U20126 ( .A(n9672), .B(n9674), .Z(n19068) );
  XNOR U20127 ( .A(q[8]), .B(DB[1313]), .Z(n9674) );
  XNOR U20128 ( .A(q[11]), .B(DB[1316]), .Z(n9672) );
  IV U20129 ( .A(n9671), .Z(n19067) );
  XNOR U20130 ( .A(n9669), .B(n19069), .Z(n9671) );
  XNOR U20131 ( .A(q[10]), .B(DB[1315]), .Z(n19069) );
  XNOR U20132 ( .A(q[9]), .B(DB[1314]), .Z(n9669) );
  IV U20133 ( .A(n9684), .Z(n19063) );
  XOR U20134 ( .A(n19070), .B(n19071), .Z(n9684) );
  XNOR U20135 ( .A(n9701), .B(n9682), .Z(n19071) );
  XNOR U20136 ( .A(q[0]), .B(DB[1305]), .Z(n9682) );
  XOR U20137 ( .A(n19072), .B(n9690), .Z(n9701) );
  XNOR U20138 ( .A(q[7]), .B(DB[1312]), .Z(n9690) );
  IV U20139 ( .A(n9689), .Z(n19072) );
  XNOR U20140 ( .A(n9687), .B(n19073), .Z(n9689) );
  XNOR U20141 ( .A(q[6]), .B(DB[1311]), .Z(n19073) );
  XNOR U20142 ( .A(q[5]), .B(DB[1310]), .Z(n9687) );
  IV U20143 ( .A(n9700), .Z(n19070) );
  XOR U20144 ( .A(n19074), .B(n19075), .Z(n9700) );
  XNOR U20145 ( .A(n9696), .B(n9698), .Z(n19075) );
  XNOR U20146 ( .A(q[1]), .B(DB[1306]), .Z(n9698) );
  XNOR U20147 ( .A(q[4]), .B(DB[1309]), .Z(n9696) );
  IV U20148 ( .A(n9695), .Z(n19074) );
  XNOR U20149 ( .A(n9693), .B(n19076), .Z(n9695) );
  XNOR U20150 ( .A(q[3]), .B(DB[1308]), .Z(n19076) );
  XNOR U20151 ( .A(q[2]), .B(DB[1307]), .Z(n9693) );
  XOR U20152 ( .A(n19077), .B(n9591), .Z(n9519) );
  XOR U20153 ( .A(n19078), .B(n9583), .Z(n9591) );
  XOR U20154 ( .A(n19079), .B(n9572), .Z(n9583) );
  XNOR U20155 ( .A(q[14]), .B(DB[1334]), .Z(n9572) );
  IV U20156 ( .A(n9571), .Z(n19079) );
  XNOR U20157 ( .A(n9569), .B(n19080), .Z(n9571) );
  XNOR U20158 ( .A(q[13]), .B(DB[1333]), .Z(n19080) );
  XNOR U20159 ( .A(q[12]), .B(DB[1332]), .Z(n9569) );
  IV U20160 ( .A(n9582), .Z(n19078) );
  XOR U20161 ( .A(n19081), .B(n19082), .Z(n9582) );
  XNOR U20162 ( .A(n9578), .B(n9580), .Z(n19082) );
  XNOR U20163 ( .A(q[8]), .B(DB[1328]), .Z(n9580) );
  XNOR U20164 ( .A(q[11]), .B(DB[1331]), .Z(n9578) );
  IV U20165 ( .A(n9577), .Z(n19081) );
  XNOR U20166 ( .A(n9575), .B(n19083), .Z(n9577) );
  XNOR U20167 ( .A(q[10]), .B(DB[1330]), .Z(n19083) );
  XNOR U20168 ( .A(q[9]), .B(DB[1329]), .Z(n9575) );
  IV U20169 ( .A(n9590), .Z(n19077) );
  XOR U20170 ( .A(n19084), .B(n19085), .Z(n9590) );
  XNOR U20171 ( .A(n9607), .B(n9588), .Z(n19085) );
  XNOR U20172 ( .A(q[0]), .B(DB[1320]), .Z(n9588) );
  XOR U20173 ( .A(n19086), .B(n9596), .Z(n9607) );
  XNOR U20174 ( .A(q[7]), .B(DB[1327]), .Z(n9596) );
  IV U20175 ( .A(n9595), .Z(n19086) );
  XNOR U20176 ( .A(n9593), .B(n19087), .Z(n9595) );
  XNOR U20177 ( .A(q[6]), .B(DB[1326]), .Z(n19087) );
  XNOR U20178 ( .A(q[5]), .B(DB[1325]), .Z(n9593) );
  IV U20179 ( .A(n9606), .Z(n19084) );
  XOR U20180 ( .A(n19088), .B(n19089), .Z(n9606) );
  XNOR U20181 ( .A(n9602), .B(n9604), .Z(n19089) );
  XNOR U20182 ( .A(q[1]), .B(DB[1321]), .Z(n9604) );
  XNOR U20183 ( .A(q[4]), .B(DB[1324]), .Z(n9602) );
  IV U20184 ( .A(n9601), .Z(n19088) );
  XNOR U20185 ( .A(n9599), .B(n19090), .Z(n9601) );
  XNOR U20186 ( .A(q[3]), .B(DB[1323]), .Z(n19090) );
  XNOR U20187 ( .A(q[2]), .B(DB[1322]), .Z(n9599) );
  XOR U20188 ( .A(n19091), .B(n9497), .Z(n9425) );
  XOR U20189 ( .A(n19092), .B(n9489), .Z(n9497) );
  XOR U20190 ( .A(n19093), .B(n9478), .Z(n9489) );
  XNOR U20191 ( .A(q[14]), .B(DB[1349]), .Z(n9478) );
  IV U20192 ( .A(n9477), .Z(n19093) );
  XNOR U20193 ( .A(n9475), .B(n19094), .Z(n9477) );
  XNOR U20194 ( .A(q[13]), .B(DB[1348]), .Z(n19094) );
  XNOR U20195 ( .A(q[12]), .B(DB[1347]), .Z(n9475) );
  IV U20196 ( .A(n9488), .Z(n19092) );
  XOR U20197 ( .A(n19095), .B(n19096), .Z(n9488) );
  XNOR U20198 ( .A(n9484), .B(n9486), .Z(n19096) );
  XNOR U20199 ( .A(q[8]), .B(DB[1343]), .Z(n9486) );
  XNOR U20200 ( .A(q[11]), .B(DB[1346]), .Z(n9484) );
  IV U20201 ( .A(n9483), .Z(n19095) );
  XNOR U20202 ( .A(n9481), .B(n19097), .Z(n9483) );
  XNOR U20203 ( .A(q[10]), .B(DB[1345]), .Z(n19097) );
  XNOR U20204 ( .A(q[9]), .B(DB[1344]), .Z(n9481) );
  IV U20205 ( .A(n9496), .Z(n19091) );
  XOR U20206 ( .A(n19098), .B(n19099), .Z(n9496) );
  XNOR U20207 ( .A(n9513), .B(n9494), .Z(n19099) );
  XNOR U20208 ( .A(q[0]), .B(DB[1335]), .Z(n9494) );
  XOR U20209 ( .A(n19100), .B(n9502), .Z(n9513) );
  XNOR U20210 ( .A(q[7]), .B(DB[1342]), .Z(n9502) );
  IV U20211 ( .A(n9501), .Z(n19100) );
  XNOR U20212 ( .A(n9499), .B(n19101), .Z(n9501) );
  XNOR U20213 ( .A(q[6]), .B(DB[1341]), .Z(n19101) );
  XNOR U20214 ( .A(q[5]), .B(DB[1340]), .Z(n9499) );
  IV U20215 ( .A(n9512), .Z(n19098) );
  XOR U20216 ( .A(n19102), .B(n19103), .Z(n9512) );
  XNOR U20217 ( .A(n9508), .B(n9510), .Z(n19103) );
  XNOR U20218 ( .A(q[1]), .B(DB[1336]), .Z(n9510) );
  XNOR U20219 ( .A(q[4]), .B(DB[1339]), .Z(n9508) );
  IV U20220 ( .A(n9507), .Z(n19102) );
  XNOR U20221 ( .A(n9505), .B(n19104), .Z(n9507) );
  XNOR U20222 ( .A(q[3]), .B(DB[1338]), .Z(n19104) );
  XNOR U20223 ( .A(q[2]), .B(DB[1337]), .Z(n9505) );
  XOR U20224 ( .A(n19105), .B(n9403), .Z(n9331) );
  XOR U20225 ( .A(n19106), .B(n9395), .Z(n9403) );
  XOR U20226 ( .A(n19107), .B(n9384), .Z(n9395) );
  XNOR U20227 ( .A(q[14]), .B(DB[1364]), .Z(n9384) );
  IV U20228 ( .A(n9383), .Z(n19107) );
  XNOR U20229 ( .A(n9381), .B(n19108), .Z(n9383) );
  XNOR U20230 ( .A(q[13]), .B(DB[1363]), .Z(n19108) );
  XNOR U20231 ( .A(q[12]), .B(DB[1362]), .Z(n9381) );
  IV U20232 ( .A(n9394), .Z(n19106) );
  XOR U20233 ( .A(n19109), .B(n19110), .Z(n9394) );
  XNOR U20234 ( .A(n9390), .B(n9392), .Z(n19110) );
  XNOR U20235 ( .A(q[8]), .B(DB[1358]), .Z(n9392) );
  XNOR U20236 ( .A(q[11]), .B(DB[1361]), .Z(n9390) );
  IV U20237 ( .A(n9389), .Z(n19109) );
  XNOR U20238 ( .A(n9387), .B(n19111), .Z(n9389) );
  XNOR U20239 ( .A(q[10]), .B(DB[1360]), .Z(n19111) );
  XNOR U20240 ( .A(q[9]), .B(DB[1359]), .Z(n9387) );
  IV U20241 ( .A(n9402), .Z(n19105) );
  XOR U20242 ( .A(n19112), .B(n19113), .Z(n9402) );
  XNOR U20243 ( .A(n9419), .B(n9400), .Z(n19113) );
  XNOR U20244 ( .A(q[0]), .B(DB[1350]), .Z(n9400) );
  XOR U20245 ( .A(n19114), .B(n9408), .Z(n9419) );
  XNOR U20246 ( .A(q[7]), .B(DB[1357]), .Z(n9408) );
  IV U20247 ( .A(n9407), .Z(n19114) );
  XNOR U20248 ( .A(n9405), .B(n19115), .Z(n9407) );
  XNOR U20249 ( .A(q[6]), .B(DB[1356]), .Z(n19115) );
  XNOR U20250 ( .A(q[5]), .B(DB[1355]), .Z(n9405) );
  IV U20251 ( .A(n9418), .Z(n19112) );
  XOR U20252 ( .A(n19116), .B(n19117), .Z(n9418) );
  XNOR U20253 ( .A(n9414), .B(n9416), .Z(n19117) );
  XNOR U20254 ( .A(q[1]), .B(DB[1351]), .Z(n9416) );
  XNOR U20255 ( .A(q[4]), .B(DB[1354]), .Z(n9414) );
  IV U20256 ( .A(n9413), .Z(n19116) );
  XNOR U20257 ( .A(n9411), .B(n19118), .Z(n9413) );
  XNOR U20258 ( .A(q[3]), .B(DB[1353]), .Z(n19118) );
  XNOR U20259 ( .A(q[2]), .B(DB[1352]), .Z(n9411) );
  XOR U20260 ( .A(n19119), .B(n9309), .Z(n9237) );
  XOR U20261 ( .A(n19120), .B(n9301), .Z(n9309) );
  XOR U20262 ( .A(n19121), .B(n9290), .Z(n9301) );
  XNOR U20263 ( .A(q[14]), .B(DB[1379]), .Z(n9290) );
  IV U20264 ( .A(n9289), .Z(n19121) );
  XNOR U20265 ( .A(n9287), .B(n19122), .Z(n9289) );
  XNOR U20266 ( .A(q[13]), .B(DB[1378]), .Z(n19122) );
  XNOR U20267 ( .A(q[12]), .B(DB[1377]), .Z(n9287) );
  IV U20268 ( .A(n9300), .Z(n19120) );
  XOR U20269 ( .A(n19123), .B(n19124), .Z(n9300) );
  XNOR U20270 ( .A(n9296), .B(n9298), .Z(n19124) );
  XNOR U20271 ( .A(q[8]), .B(DB[1373]), .Z(n9298) );
  XNOR U20272 ( .A(q[11]), .B(DB[1376]), .Z(n9296) );
  IV U20273 ( .A(n9295), .Z(n19123) );
  XNOR U20274 ( .A(n9293), .B(n19125), .Z(n9295) );
  XNOR U20275 ( .A(q[10]), .B(DB[1375]), .Z(n19125) );
  XNOR U20276 ( .A(q[9]), .B(DB[1374]), .Z(n9293) );
  IV U20277 ( .A(n9308), .Z(n19119) );
  XOR U20278 ( .A(n19126), .B(n19127), .Z(n9308) );
  XNOR U20279 ( .A(n9325), .B(n9306), .Z(n19127) );
  XNOR U20280 ( .A(q[0]), .B(DB[1365]), .Z(n9306) );
  XOR U20281 ( .A(n19128), .B(n9314), .Z(n9325) );
  XNOR U20282 ( .A(q[7]), .B(DB[1372]), .Z(n9314) );
  IV U20283 ( .A(n9313), .Z(n19128) );
  XNOR U20284 ( .A(n9311), .B(n19129), .Z(n9313) );
  XNOR U20285 ( .A(q[6]), .B(DB[1371]), .Z(n19129) );
  XNOR U20286 ( .A(q[5]), .B(DB[1370]), .Z(n9311) );
  IV U20287 ( .A(n9324), .Z(n19126) );
  XOR U20288 ( .A(n19130), .B(n19131), .Z(n9324) );
  XNOR U20289 ( .A(n9320), .B(n9322), .Z(n19131) );
  XNOR U20290 ( .A(q[1]), .B(DB[1366]), .Z(n9322) );
  XNOR U20291 ( .A(q[4]), .B(DB[1369]), .Z(n9320) );
  IV U20292 ( .A(n9319), .Z(n19130) );
  XNOR U20293 ( .A(n9317), .B(n19132), .Z(n9319) );
  XNOR U20294 ( .A(q[3]), .B(DB[1368]), .Z(n19132) );
  XNOR U20295 ( .A(q[2]), .B(DB[1367]), .Z(n9317) );
  XOR U20296 ( .A(n19133), .B(n9215), .Z(n9143) );
  XOR U20297 ( .A(n19134), .B(n9207), .Z(n9215) );
  XOR U20298 ( .A(n19135), .B(n9196), .Z(n9207) );
  XNOR U20299 ( .A(q[14]), .B(DB[1394]), .Z(n9196) );
  IV U20300 ( .A(n9195), .Z(n19135) );
  XNOR U20301 ( .A(n9193), .B(n19136), .Z(n9195) );
  XNOR U20302 ( .A(q[13]), .B(DB[1393]), .Z(n19136) );
  XNOR U20303 ( .A(q[12]), .B(DB[1392]), .Z(n9193) );
  IV U20304 ( .A(n9206), .Z(n19134) );
  XOR U20305 ( .A(n19137), .B(n19138), .Z(n9206) );
  XNOR U20306 ( .A(n9202), .B(n9204), .Z(n19138) );
  XNOR U20307 ( .A(q[8]), .B(DB[1388]), .Z(n9204) );
  XNOR U20308 ( .A(q[11]), .B(DB[1391]), .Z(n9202) );
  IV U20309 ( .A(n9201), .Z(n19137) );
  XNOR U20310 ( .A(n9199), .B(n19139), .Z(n9201) );
  XNOR U20311 ( .A(q[10]), .B(DB[1390]), .Z(n19139) );
  XNOR U20312 ( .A(q[9]), .B(DB[1389]), .Z(n9199) );
  IV U20313 ( .A(n9214), .Z(n19133) );
  XOR U20314 ( .A(n19140), .B(n19141), .Z(n9214) );
  XNOR U20315 ( .A(n9231), .B(n9212), .Z(n19141) );
  XNOR U20316 ( .A(q[0]), .B(DB[1380]), .Z(n9212) );
  XOR U20317 ( .A(n19142), .B(n9220), .Z(n9231) );
  XNOR U20318 ( .A(q[7]), .B(DB[1387]), .Z(n9220) );
  IV U20319 ( .A(n9219), .Z(n19142) );
  XNOR U20320 ( .A(n9217), .B(n19143), .Z(n9219) );
  XNOR U20321 ( .A(q[6]), .B(DB[1386]), .Z(n19143) );
  XNOR U20322 ( .A(q[5]), .B(DB[1385]), .Z(n9217) );
  IV U20323 ( .A(n9230), .Z(n19140) );
  XOR U20324 ( .A(n19144), .B(n19145), .Z(n9230) );
  XNOR U20325 ( .A(n9226), .B(n9228), .Z(n19145) );
  XNOR U20326 ( .A(q[1]), .B(DB[1381]), .Z(n9228) );
  XNOR U20327 ( .A(q[4]), .B(DB[1384]), .Z(n9226) );
  IV U20328 ( .A(n9225), .Z(n19144) );
  XNOR U20329 ( .A(n9223), .B(n19146), .Z(n9225) );
  XNOR U20330 ( .A(q[3]), .B(DB[1383]), .Z(n19146) );
  XNOR U20331 ( .A(q[2]), .B(DB[1382]), .Z(n9223) );
  XOR U20332 ( .A(n19147), .B(n9121), .Z(n9049) );
  XOR U20333 ( .A(n19148), .B(n9113), .Z(n9121) );
  XOR U20334 ( .A(n19149), .B(n9102), .Z(n9113) );
  XNOR U20335 ( .A(q[14]), .B(DB[1409]), .Z(n9102) );
  IV U20336 ( .A(n9101), .Z(n19149) );
  XNOR U20337 ( .A(n9099), .B(n19150), .Z(n9101) );
  XNOR U20338 ( .A(q[13]), .B(DB[1408]), .Z(n19150) );
  XNOR U20339 ( .A(q[12]), .B(DB[1407]), .Z(n9099) );
  IV U20340 ( .A(n9112), .Z(n19148) );
  XOR U20341 ( .A(n19151), .B(n19152), .Z(n9112) );
  XNOR U20342 ( .A(n9108), .B(n9110), .Z(n19152) );
  XNOR U20343 ( .A(q[8]), .B(DB[1403]), .Z(n9110) );
  XNOR U20344 ( .A(q[11]), .B(DB[1406]), .Z(n9108) );
  IV U20345 ( .A(n9107), .Z(n19151) );
  XNOR U20346 ( .A(n9105), .B(n19153), .Z(n9107) );
  XNOR U20347 ( .A(q[10]), .B(DB[1405]), .Z(n19153) );
  XNOR U20348 ( .A(q[9]), .B(DB[1404]), .Z(n9105) );
  IV U20349 ( .A(n9120), .Z(n19147) );
  XOR U20350 ( .A(n19154), .B(n19155), .Z(n9120) );
  XNOR U20351 ( .A(n9137), .B(n9118), .Z(n19155) );
  XNOR U20352 ( .A(q[0]), .B(DB[1395]), .Z(n9118) );
  XOR U20353 ( .A(n19156), .B(n9126), .Z(n9137) );
  XNOR U20354 ( .A(q[7]), .B(DB[1402]), .Z(n9126) );
  IV U20355 ( .A(n9125), .Z(n19156) );
  XNOR U20356 ( .A(n9123), .B(n19157), .Z(n9125) );
  XNOR U20357 ( .A(q[6]), .B(DB[1401]), .Z(n19157) );
  XNOR U20358 ( .A(q[5]), .B(DB[1400]), .Z(n9123) );
  IV U20359 ( .A(n9136), .Z(n19154) );
  XOR U20360 ( .A(n19158), .B(n19159), .Z(n9136) );
  XNOR U20361 ( .A(n9132), .B(n9134), .Z(n19159) );
  XNOR U20362 ( .A(q[1]), .B(DB[1396]), .Z(n9134) );
  XNOR U20363 ( .A(q[4]), .B(DB[1399]), .Z(n9132) );
  IV U20364 ( .A(n9131), .Z(n19158) );
  XNOR U20365 ( .A(n9129), .B(n19160), .Z(n9131) );
  XNOR U20366 ( .A(q[3]), .B(DB[1398]), .Z(n19160) );
  XNOR U20367 ( .A(q[2]), .B(DB[1397]), .Z(n9129) );
  XOR U20368 ( .A(n19161), .B(n9027), .Z(n8955) );
  XOR U20369 ( .A(n19162), .B(n9019), .Z(n9027) );
  XOR U20370 ( .A(n19163), .B(n9008), .Z(n9019) );
  XNOR U20371 ( .A(q[14]), .B(DB[1424]), .Z(n9008) );
  IV U20372 ( .A(n9007), .Z(n19163) );
  XNOR U20373 ( .A(n9005), .B(n19164), .Z(n9007) );
  XNOR U20374 ( .A(q[13]), .B(DB[1423]), .Z(n19164) );
  XNOR U20375 ( .A(q[12]), .B(DB[1422]), .Z(n9005) );
  IV U20376 ( .A(n9018), .Z(n19162) );
  XOR U20377 ( .A(n19165), .B(n19166), .Z(n9018) );
  XNOR U20378 ( .A(n9014), .B(n9016), .Z(n19166) );
  XNOR U20379 ( .A(q[8]), .B(DB[1418]), .Z(n9016) );
  XNOR U20380 ( .A(q[11]), .B(DB[1421]), .Z(n9014) );
  IV U20381 ( .A(n9013), .Z(n19165) );
  XNOR U20382 ( .A(n9011), .B(n19167), .Z(n9013) );
  XNOR U20383 ( .A(q[10]), .B(DB[1420]), .Z(n19167) );
  XNOR U20384 ( .A(q[9]), .B(DB[1419]), .Z(n9011) );
  IV U20385 ( .A(n9026), .Z(n19161) );
  XOR U20386 ( .A(n19168), .B(n19169), .Z(n9026) );
  XNOR U20387 ( .A(n9043), .B(n9024), .Z(n19169) );
  XNOR U20388 ( .A(q[0]), .B(DB[1410]), .Z(n9024) );
  XOR U20389 ( .A(n19170), .B(n9032), .Z(n9043) );
  XNOR U20390 ( .A(q[7]), .B(DB[1417]), .Z(n9032) );
  IV U20391 ( .A(n9031), .Z(n19170) );
  XNOR U20392 ( .A(n9029), .B(n19171), .Z(n9031) );
  XNOR U20393 ( .A(q[6]), .B(DB[1416]), .Z(n19171) );
  XNOR U20394 ( .A(q[5]), .B(DB[1415]), .Z(n9029) );
  IV U20395 ( .A(n9042), .Z(n19168) );
  XOR U20396 ( .A(n19172), .B(n19173), .Z(n9042) );
  XNOR U20397 ( .A(n9038), .B(n9040), .Z(n19173) );
  XNOR U20398 ( .A(q[1]), .B(DB[1411]), .Z(n9040) );
  XNOR U20399 ( .A(q[4]), .B(DB[1414]), .Z(n9038) );
  IV U20400 ( .A(n9037), .Z(n19172) );
  XNOR U20401 ( .A(n9035), .B(n19174), .Z(n9037) );
  XNOR U20402 ( .A(q[3]), .B(DB[1413]), .Z(n19174) );
  XNOR U20403 ( .A(q[2]), .B(DB[1412]), .Z(n9035) );
  XOR U20404 ( .A(n19175), .B(n8933), .Z(n8861) );
  XOR U20405 ( .A(n19176), .B(n8925), .Z(n8933) );
  XOR U20406 ( .A(n19177), .B(n8914), .Z(n8925) );
  XNOR U20407 ( .A(q[14]), .B(DB[1439]), .Z(n8914) );
  IV U20408 ( .A(n8913), .Z(n19177) );
  XNOR U20409 ( .A(n8911), .B(n19178), .Z(n8913) );
  XNOR U20410 ( .A(q[13]), .B(DB[1438]), .Z(n19178) );
  XNOR U20411 ( .A(q[12]), .B(DB[1437]), .Z(n8911) );
  IV U20412 ( .A(n8924), .Z(n19176) );
  XOR U20413 ( .A(n19179), .B(n19180), .Z(n8924) );
  XNOR U20414 ( .A(n8920), .B(n8922), .Z(n19180) );
  XNOR U20415 ( .A(q[8]), .B(DB[1433]), .Z(n8922) );
  XNOR U20416 ( .A(q[11]), .B(DB[1436]), .Z(n8920) );
  IV U20417 ( .A(n8919), .Z(n19179) );
  XNOR U20418 ( .A(n8917), .B(n19181), .Z(n8919) );
  XNOR U20419 ( .A(q[10]), .B(DB[1435]), .Z(n19181) );
  XNOR U20420 ( .A(q[9]), .B(DB[1434]), .Z(n8917) );
  IV U20421 ( .A(n8932), .Z(n19175) );
  XOR U20422 ( .A(n19182), .B(n19183), .Z(n8932) );
  XNOR U20423 ( .A(n8949), .B(n8930), .Z(n19183) );
  XNOR U20424 ( .A(q[0]), .B(DB[1425]), .Z(n8930) );
  XOR U20425 ( .A(n19184), .B(n8938), .Z(n8949) );
  XNOR U20426 ( .A(q[7]), .B(DB[1432]), .Z(n8938) );
  IV U20427 ( .A(n8937), .Z(n19184) );
  XNOR U20428 ( .A(n8935), .B(n19185), .Z(n8937) );
  XNOR U20429 ( .A(q[6]), .B(DB[1431]), .Z(n19185) );
  XNOR U20430 ( .A(q[5]), .B(DB[1430]), .Z(n8935) );
  IV U20431 ( .A(n8948), .Z(n19182) );
  XOR U20432 ( .A(n19186), .B(n19187), .Z(n8948) );
  XNOR U20433 ( .A(n8944), .B(n8946), .Z(n19187) );
  XNOR U20434 ( .A(q[1]), .B(DB[1426]), .Z(n8946) );
  XNOR U20435 ( .A(q[4]), .B(DB[1429]), .Z(n8944) );
  IV U20436 ( .A(n8943), .Z(n19186) );
  XNOR U20437 ( .A(n8941), .B(n19188), .Z(n8943) );
  XNOR U20438 ( .A(q[3]), .B(DB[1428]), .Z(n19188) );
  XNOR U20439 ( .A(q[2]), .B(DB[1427]), .Z(n8941) );
  XOR U20440 ( .A(n19189), .B(n8839), .Z(n8767) );
  XOR U20441 ( .A(n19190), .B(n8831), .Z(n8839) );
  XOR U20442 ( .A(n19191), .B(n8820), .Z(n8831) );
  XNOR U20443 ( .A(q[14]), .B(DB[1454]), .Z(n8820) );
  IV U20444 ( .A(n8819), .Z(n19191) );
  XNOR U20445 ( .A(n8817), .B(n19192), .Z(n8819) );
  XNOR U20446 ( .A(q[13]), .B(DB[1453]), .Z(n19192) );
  XNOR U20447 ( .A(q[12]), .B(DB[1452]), .Z(n8817) );
  IV U20448 ( .A(n8830), .Z(n19190) );
  XOR U20449 ( .A(n19193), .B(n19194), .Z(n8830) );
  XNOR U20450 ( .A(n8826), .B(n8828), .Z(n19194) );
  XNOR U20451 ( .A(q[8]), .B(DB[1448]), .Z(n8828) );
  XNOR U20452 ( .A(q[11]), .B(DB[1451]), .Z(n8826) );
  IV U20453 ( .A(n8825), .Z(n19193) );
  XNOR U20454 ( .A(n8823), .B(n19195), .Z(n8825) );
  XNOR U20455 ( .A(q[10]), .B(DB[1450]), .Z(n19195) );
  XNOR U20456 ( .A(q[9]), .B(DB[1449]), .Z(n8823) );
  IV U20457 ( .A(n8838), .Z(n19189) );
  XOR U20458 ( .A(n19196), .B(n19197), .Z(n8838) );
  XNOR U20459 ( .A(n8855), .B(n8836), .Z(n19197) );
  XNOR U20460 ( .A(q[0]), .B(DB[1440]), .Z(n8836) );
  XOR U20461 ( .A(n19198), .B(n8844), .Z(n8855) );
  XNOR U20462 ( .A(q[7]), .B(DB[1447]), .Z(n8844) );
  IV U20463 ( .A(n8843), .Z(n19198) );
  XNOR U20464 ( .A(n8841), .B(n19199), .Z(n8843) );
  XNOR U20465 ( .A(q[6]), .B(DB[1446]), .Z(n19199) );
  XNOR U20466 ( .A(q[5]), .B(DB[1445]), .Z(n8841) );
  IV U20467 ( .A(n8854), .Z(n19196) );
  XOR U20468 ( .A(n19200), .B(n19201), .Z(n8854) );
  XNOR U20469 ( .A(n8850), .B(n8852), .Z(n19201) );
  XNOR U20470 ( .A(q[1]), .B(DB[1441]), .Z(n8852) );
  XNOR U20471 ( .A(q[4]), .B(DB[1444]), .Z(n8850) );
  IV U20472 ( .A(n8849), .Z(n19200) );
  XNOR U20473 ( .A(n8847), .B(n19202), .Z(n8849) );
  XNOR U20474 ( .A(q[3]), .B(DB[1443]), .Z(n19202) );
  XNOR U20475 ( .A(q[2]), .B(DB[1442]), .Z(n8847) );
  XOR U20476 ( .A(n19203), .B(n8745), .Z(n8673) );
  XOR U20477 ( .A(n19204), .B(n8737), .Z(n8745) );
  XOR U20478 ( .A(n19205), .B(n8726), .Z(n8737) );
  XNOR U20479 ( .A(q[14]), .B(DB[1469]), .Z(n8726) );
  IV U20480 ( .A(n8725), .Z(n19205) );
  XNOR U20481 ( .A(n8723), .B(n19206), .Z(n8725) );
  XNOR U20482 ( .A(q[13]), .B(DB[1468]), .Z(n19206) );
  XNOR U20483 ( .A(q[12]), .B(DB[1467]), .Z(n8723) );
  IV U20484 ( .A(n8736), .Z(n19204) );
  XOR U20485 ( .A(n19207), .B(n19208), .Z(n8736) );
  XNOR U20486 ( .A(n8732), .B(n8734), .Z(n19208) );
  XNOR U20487 ( .A(q[8]), .B(DB[1463]), .Z(n8734) );
  XNOR U20488 ( .A(q[11]), .B(DB[1466]), .Z(n8732) );
  IV U20489 ( .A(n8731), .Z(n19207) );
  XNOR U20490 ( .A(n8729), .B(n19209), .Z(n8731) );
  XNOR U20491 ( .A(q[10]), .B(DB[1465]), .Z(n19209) );
  XNOR U20492 ( .A(q[9]), .B(DB[1464]), .Z(n8729) );
  IV U20493 ( .A(n8744), .Z(n19203) );
  XOR U20494 ( .A(n19210), .B(n19211), .Z(n8744) );
  XNOR U20495 ( .A(n8761), .B(n8742), .Z(n19211) );
  XNOR U20496 ( .A(q[0]), .B(DB[1455]), .Z(n8742) );
  XOR U20497 ( .A(n19212), .B(n8750), .Z(n8761) );
  XNOR U20498 ( .A(q[7]), .B(DB[1462]), .Z(n8750) );
  IV U20499 ( .A(n8749), .Z(n19212) );
  XNOR U20500 ( .A(n8747), .B(n19213), .Z(n8749) );
  XNOR U20501 ( .A(q[6]), .B(DB[1461]), .Z(n19213) );
  XNOR U20502 ( .A(q[5]), .B(DB[1460]), .Z(n8747) );
  IV U20503 ( .A(n8760), .Z(n19210) );
  XOR U20504 ( .A(n19214), .B(n19215), .Z(n8760) );
  XNOR U20505 ( .A(n8756), .B(n8758), .Z(n19215) );
  XNOR U20506 ( .A(q[1]), .B(DB[1456]), .Z(n8758) );
  XNOR U20507 ( .A(q[4]), .B(DB[1459]), .Z(n8756) );
  IV U20508 ( .A(n8755), .Z(n19214) );
  XNOR U20509 ( .A(n8753), .B(n19216), .Z(n8755) );
  XNOR U20510 ( .A(q[3]), .B(DB[1458]), .Z(n19216) );
  XNOR U20511 ( .A(q[2]), .B(DB[1457]), .Z(n8753) );
  XOR U20512 ( .A(n19217), .B(n8651), .Z(n8579) );
  XOR U20513 ( .A(n19218), .B(n8643), .Z(n8651) );
  XOR U20514 ( .A(n19219), .B(n8632), .Z(n8643) );
  XNOR U20515 ( .A(q[14]), .B(DB[1484]), .Z(n8632) );
  IV U20516 ( .A(n8631), .Z(n19219) );
  XNOR U20517 ( .A(n8629), .B(n19220), .Z(n8631) );
  XNOR U20518 ( .A(q[13]), .B(DB[1483]), .Z(n19220) );
  XNOR U20519 ( .A(q[12]), .B(DB[1482]), .Z(n8629) );
  IV U20520 ( .A(n8642), .Z(n19218) );
  XOR U20521 ( .A(n19221), .B(n19222), .Z(n8642) );
  XNOR U20522 ( .A(n8638), .B(n8640), .Z(n19222) );
  XNOR U20523 ( .A(q[8]), .B(DB[1478]), .Z(n8640) );
  XNOR U20524 ( .A(q[11]), .B(DB[1481]), .Z(n8638) );
  IV U20525 ( .A(n8637), .Z(n19221) );
  XNOR U20526 ( .A(n8635), .B(n19223), .Z(n8637) );
  XNOR U20527 ( .A(q[10]), .B(DB[1480]), .Z(n19223) );
  XNOR U20528 ( .A(q[9]), .B(DB[1479]), .Z(n8635) );
  IV U20529 ( .A(n8650), .Z(n19217) );
  XOR U20530 ( .A(n19224), .B(n19225), .Z(n8650) );
  XNOR U20531 ( .A(n8667), .B(n8648), .Z(n19225) );
  XNOR U20532 ( .A(q[0]), .B(DB[1470]), .Z(n8648) );
  XOR U20533 ( .A(n19226), .B(n8656), .Z(n8667) );
  XNOR U20534 ( .A(q[7]), .B(DB[1477]), .Z(n8656) );
  IV U20535 ( .A(n8655), .Z(n19226) );
  XNOR U20536 ( .A(n8653), .B(n19227), .Z(n8655) );
  XNOR U20537 ( .A(q[6]), .B(DB[1476]), .Z(n19227) );
  XNOR U20538 ( .A(q[5]), .B(DB[1475]), .Z(n8653) );
  IV U20539 ( .A(n8666), .Z(n19224) );
  XOR U20540 ( .A(n19228), .B(n19229), .Z(n8666) );
  XNOR U20541 ( .A(n8662), .B(n8664), .Z(n19229) );
  XNOR U20542 ( .A(q[1]), .B(DB[1471]), .Z(n8664) );
  XNOR U20543 ( .A(q[4]), .B(DB[1474]), .Z(n8662) );
  IV U20544 ( .A(n8661), .Z(n19228) );
  XNOR U20545 ( .A(n8659), .B(n19230), .Z(n8661) );
  XNOR U20546 ( .A(q[3]), .B(DB[1473]), .Z(n19230) );
  XNOR U20547 ( .A(q[2]), .B(DB[1472]), .Z(n8659) );
  XOR U20548 ( .A(n19231), .B(n8557), .Z(n8485) );
  XOR U20549 ( .A(n19232), .B(n8549), .Z(n8557) );
  XOR U20550 ( .A(n19233), .B(n8538), .Z(n8549) );
  XNOR U20551 ( .A(q[14]), .B(DB[1499]), .Z(n8538) );
  IV U20552 ( .A(n8537), .Z(n19233) );
  XNOR U20553 ( .A(n8535), .B(n19234), .Z(n8537) );
  XNOR U20554 ( .A(q[13]), .B(DB[1498]), .Z(n19234) );
  XNOR U20555 ( .A(q[12]), .B(DB[1497]), .Z(n8535) );
  IV U20556 ( .A(n8548), .Z(n19232) );
  XOR U20557 ( .A(n19235), .B(n19236), .Z(n8548) );
  XNOR U20558 ( .A(n8544), .B(n8546), .Z(n19236) );
  XNOR U20559 ( .A(q[8]), .B(DB[1493]), .Z(n8546) );
  XNOR U20560 ( .A(q[11]), .B(DB[1496]), .Z(n8544) );
  IV U20561 ( .A(n8543), .Z(n19235) );
  XNOR U20562 ( .A(n8541), .B(n19237), .Z(n8543) );
  XNOR U20563 ( .A(q[10]), .B(DB[1495]), .Z(n19237) );
  XNOR U20564 ( .A(q[9]), .B(DB[1494]), .Z(n8541) );
  IV U20565 ( .A(n8556), .Z(n19231) );
  XOR U20566 ( .A(n19238), .B(n19239), .Z(n8556) );
  XNOR U20567 ( .A(n8573), .B(n8554), .Z(n19239) );
  XNOR U20568 ( .A(q[0]), .B(DB[1485]), .Z(n8554) );
  XOR U20569 ( .A(n19240), .B(n8562), .Z(n8573) );
  XNOR U20570 ( .A(q[7]), .B(DB[1492]), .Z(n8562) );
  IV U20571 ( .A(n8561), .Z(n19240) );
  XNOR U20572 ( .A(n8559), .B(n19241), .Z(n8561) );
  XNOR U20573 ( .A(q[6]), .B(DB[1491]), .Z(n19241) );
  XNOR U20574 ( .A(q[5]), .B(DB[1490]), .Z(n8559) );
  IV U20575 ( .A(n8572), .Z(n19238) );
  XOR U20576 ( .A(n19242), .B(n19243), .Z(n8572) );
  XNOR U20577 ( .A(n8568), .B(n8570), .Z(n19243) );
  XNOR U20578 ( .A(q[1]), .B(DB[1486]), .Z(n8570) );
  XNOR U20579 ( .A(q[4]), .B(DB[1489]), .Z(n8568) );
  IV U20580 ( .A(n8567), .Z(n19242) );
  XNOR U20581 ( .A(n8565), .B(n19244), .Z(n8567) );
  XNOR U20582 ( .A(q[3]), .B(DB[1488]), .Z(n19244) );
  XNOR U20583 ( .A(q[2]), .B(DB[1487]), .Z(n8565) );
  XOR U20584 ( .A(n19245), .B(n8463), .Z(n8391) );
  XOR U20585 ( .A(n19246), .B(n8455), .Z(n8463) );
  XOR U20586 ( .A(n19247), .B(n8444), .Z(n8455) );
  XNOR U20587 ( .A(q[14]), .B(DB[1514]), .Z(n8444) );
  IV U20588 ( .A(n8443), .Z(n19247) );
  XNOR U20589 ( .A(n8441), .B(n19248), .Z(n8443) );
  XNOR U20590 ( .A(q[13]), .B(DB[1513]), .Z(n19248) );
  XNOR U20591 ( .A(q[12]), .B(DB[1512]), .Z(n8441) );
  IV U20592 ( .A(n8454), .Z(n19246) );
  XOR U20593 ( .A(n19249), .B(n19250), .Z(n8454) );
  XNOR U20594 ( .A(n8450), .B(n8452), .Z(n19250) );
  XNOR U20595 ( .A(q[8]), .B(DB[1508]), .Z(n8452) );
  XNOR U20596 ( .A(q[11]), .B(DB[1511]), .Z(n8450) );
  IV U20597 ( .A(n8449), .Z(n19249) );
  XNOR U20598 ( .A(n8447), .B(n19251), .Z(n8449) );
  XNOR U20599 ( .A(q[10]), .B(DB[1510]), .Z(n19251) );
  XNOR U20600 ( .A(q[9]), .B(DB[1509]), .Z(n8447) );
  IV U20601 ( .A(n8462), .Z(n19245) );
  XOR U20602 ( .A(n19252), .B(n19253), .Z(n8462) );
  XNOR U20603 ( .A(n8479), .B(n8460), .Z(n19253) );
  XNOR U20604 ( .A(q[0]), .B(DB[1500]), .Z(n8460) );
  XOR U20605 ( .A(n19254), .B(n8468), .Z(n8479) );
  XNOR U20606 ( .A(q[7]), .B(DB[1507]), .Z(n8468) );
  IV U20607 ( .A(n8467), .Z(n19254) );
  XNOR U20608 ( .A(n8465), .B(n19255), .Z(n8467) );
  XNOR U20609 ( .A(q[6]), .B(DB[1506]), .Z(n19255) );
  XNOR U20610 ( .A(q[5]), .B(DB[1505]), .Z(n8465) );
  IV U20611 ( .A(n8478), .Z(n19252) );
  XOR U20612 ( .A(n19256), .B(n19257), .Z(n8478) );
  XNOR U20613 ( .A(n8474), .B(n8476), .Z(n19257) );
  XNOR U20614 ( .A(q[1]), .B(DB[1501]), .Z(n8476) );
  XNOR U20615 ( .A(q[4]), .B(DB[1504]), .Z(n8474) );
  IV U20616 ( .A(n8473), .Z(n19256) );
  XNOR U20617 ( .A(n8471), .B(n19258), .Z(n8473) );
  XNOR U20618 ( .A(q[3]), .B(DB[1503]), .Z(n19258) );
  XNOR U20619 ( .A(q[2]), .B(DB[1502]), .Z(n8471) );
  XOR U20620 ( .A(n19259), .B(n8369), .Z(n8297) );
  XOR U20621 ( .A(n19260), .B(n8361), .Z(n8369) );
  XOR U20622 ( .A(n19261), .B(n8350), .Z(n8361) );
  XNOR U20623 ( .A(q[14]), .B(DB[1529]), .Z(n8350) );
  IV U20624 ( .A(n8349), .Z(n19261) );
  XNOR U20625 ( .A(n8347), .B(n19262), .Z(n8349) );
  XNOR U20626 ( .A(q[13]), .B(DB[1528]), .Z(n19262) );
  XNOR U20627 ( .A(q[12]), .B(DB[1527]), .Z(n8347) );
  IV U20628 ( .A(n8360), .Z(n19260) );
  XOR U20629 ( .A(n19263), .B(n19264), .Z(n8360) );
  XNOR U20630 ( .A(n8356), .B(n8358), .Z(n19264) );
  XNOR U20631 ( .A(q[8]), .B(DB[1523]), .Z(n8358) );
  XNOR U20632 ( .A(q[11]), .B(DB[1526]), .Z(n8356) );
  IV U20633 ( .A(n8355), .Z(n19263) );
  XNOR U20634 ( .A(n8353), .B(n19265), .Z(n8355) );
  XNOR U20635 ( .A(q[10]), .B(DB[1525]), .Z(n19265) );
  XNOR U20636 ( .A(q[9]), .B(DB[1524]), .Z(n8353) );
  IV U20637 ( .A(n8368), .Z(n19259) );
  XOR U20638 ( .A(n19266), .B(n19267), .Z(n8368) );
  XNOR U20639 ( .A(n8385), .B(n8366), .Z(n19267) );
  XNOR U20640 ( .A(q[0]), .B(DB[1515]), .Z(n8366) );
  XOR U20641 ( .A(n19268), .B(n8374), .Z(n8385) );
  XNOR U20642 ( .A(q[7]), .B(DB[1522]), .Z(n8374) );
  IV U20643 ( .A(n8373), .Z(n19268) );
  XNOR U20644 ( .A(n8371), .B(n19269), .Z(n8373) );
  XNOR U20645 ( .A(q[6]), .B(DB[1521]), .Z(n19269) );
  XNOR U20646 ( .A(q[5]), .B(DB[1520]), .Z(n8371) );
  IV U20647 ( .A(n8384), .Z(n19266) );
  XOR U20648 ( .A(n19270), .B(n19271), .Z(n8384) );
  XNOR U20649 ( .A(n8380), .B(n8382), .Z(n19271) );
  XNOR U20650 ( .A(q[1]), .B(DB[1516]), .Z(n8382) );
  XNOR U20651 ( .A(q[4]), .B(DB[1519]), .Z(n8380) );
  IV U20652 ( .A(n8379), .Z(n19270) );
  XNOR U20653 ( .A(n8377), .B(n19272), .Z(n8379) );
  XNOR U20654 ( .A(q[3]), .B(DB[1518]), .Z(n19272) );
  XNOR U20655 ( .A(q[2]), .B(DB[1517]), .Z(n8377) );
  XOR U20656 ( .A(n19273), .B(n8275), .Z(n8203) );
  XOR U20657 ( .A(n19274), .B(n8267), .Z(n8275) );
  XOR U20658 ( .A(n19275), .B(n8256), .Z(n8267) );
  XNOR U20659 ( .A(q[14]), .B(DB[1544]), .Z(n8256) );
  IV U20660 ( .A(n8255), .Z(n19275) );
  XNOR U20661 ( .A(n8253), .B(n19276), .Z(n8255) );
  XNOR U20662 ( .A(q[13]), .B(DB[1543]), .Z(n19276) );
  XNOR U20663 ( .A(q[12]), .B(DB[1542]), .Z(n8253) );
  IV U20664 ( .A(n8266), .Z(n19274) );
  XOR U20665 ( .A(n19277), .B(n19278), .Z(n8266) );
  XNOR U20666 ( .A(n8262), .B(n8264), .Z(n19278) );
  XNOR U20667 ( .A(q[8]), .B(DB[1538]), .Z(n8264) );
  XNOR U20668 ( .A(q[11]), .B(DB[1541]), .Z(n8262) );
  IV U20669 ( .A(n8261), .Z(n19277) );
  XNOR U20670 ( .A(n8259), .B(n19279), .Z(n8261) );
  XNOR U20671 ( .A(q[10]), .B(DB[1540]), .Z(n19279) );
  XNOR U20672 ( .A(q[9]), .B(DB[1539]), .Z(n8259) );
  IV U20673 ( .A(n8274), .Z(n19273) );
  XOR U20674 ( .A(n19280), .B(n19281), .Z(n8274) );
  XNOR U20675 ( .A(n8291), .B(n8272), .Z(n19281) );
  XNOR U20676 ( .A(q[0]), .B(DB[1530]), .Z(n8272) );
  XOR U20677 ( .A(n19282), .B(n8280), .Z(n8291) );
  XNOR U20678 ( .A(q[7]), .B(DB[1537]), .Z(n8280) );
  IV U20679 ( .A(n8279), .Z(n19282) );
  XNOR U20680 ( .A(n8277), .B(n19283), .Z(n8279) );
  XNOR U20681 ( .A(q[6]), .B(DB[1536]), .Z(n19283) );
  XNOR U20682 ( .A(q[5]), .B(DB[1535]), .Z(n8277) );
  IV U20683 ( .A(n8290), .Z(n19280) );
  XOR U20684 ( .A(n19284), .B(n19285), .Z(n8290) );
  XNOR U20685 ( .A(n8286), .B(n8288), .Z(n19285) );
  XNOR U20686 ( .A(q[1]), .B(DB[1531]), .Z(n8288) );
  XNOR U20687 ( .A(q[4]), .B(DB[1534]), .Z(n8286) );
  IV U20688 ( .A(n8285), .Z(n19284) );
  XNOR U20689 ( .A(n8283), .B(n19286), .Z(n8285) );
  XNOR U20690 ( .A(q[3]), .B(DB[1533]), .Z(n19286) );
  XNOR U20691 ( .A(q[2]), .B(DB[1532]), .Z(n8283) );
  XOR U20692 ( .A(n19287), .B(n8181), .Z(n8109) );
  XOR U20693 ( .A(n19288), .B(n8173), .Z(n8181) );
  XOR U20694 ( .A(n19289), .B(n8162), .Z(n8173) );
  XNOR U20695 ( .A(q[14]), .B(DB[1559]), .Z(n8162) );
  IV U20696 ( .A(n8161), .Z(n19289) );
  XNOR U20697 ( .A(n8159), .B(n19290), .Z(n8161) );
  XNOR U20698 ( .A(q[13]), .B(DB[1558]), .Z(n19290) );
  XNOR U20699 ( .A(q[12]), .B(DB[1557]), .Z(n8159) );
  IV U20700 ( .A(n8172), .Z(n19288) );
  XOR U20701 ( .A(n19291), .B(n19292), .Z(n8172) );
  XNOR U20702 ( .A(n8168), .B(n8170), .Z(n19292) );
  XNOR U20703 ( .A(q[8]), .B(DB[1553]), .Z(n8170) );
  XNOR U20704 ( .A(q[11]), .B(DB[1556]), .Z(n8168) );
  IV U20705 ( .A(n8167), .Z(n19291) );
  XNOR U20706 ( .A(n8165), .B(n19293), .Z(n8167) );
  XNOR U20707 ( .A(q[10]), .B(DB[1555]), .Z(n19293) );
  XNOR U20708 ( .A(q[9]), .B(DB[1554]), .Z(n8165) );
  IV U20709 ( .A(n8180), .Z(n19287) );
  XOR U20710 ( .A(n19294), .B(n19295), .Z(n8180) );
  XNOR U20711 ( .A(n8197), .B(n8178), .Z(n19295) );
  XNOR U20712 ( .A(q[0]), .B(DB[1545]), .Z(n8178) );
  XOR U20713 ( .A(n19296), .B(n8186), .Z(n8197) );
  XNOR U20714 ( .A(q[7]), .B(DB[1552]), .Z(n8186) );
  IV U20715 ( .A(n8185), .Z(n19296) );
  XNOR U20716 ( .A(n8183), .B(n19297), .Z(n8185) );
  XNOR U20717 ( .A(q[6]), .B(DB[1551]), .Z(n19297) );
  XNOR U20718 ( .A(q[5]), .B(DB[1550]), .Z(n8183) );
  IV U20719 ( .A(n8196), .Z(n19294) );
  XOR U20720 ( .A(n19298), .B(n19299), .Z(n8196) );
  XNOR U20721 ( .A(n8192), .B(n8194), .Z(n19299) );
  XNOR U20722 ( .A(q[1]), .B(DB[1546]), .Z(n8194) );
  XNOR U20723 ( .A(q[4]), .B(DB[1549]), .Z(n8192) );
  IV U20724 ( .A(n8191), .Z(n19298) );
  XNOR U20725 ( .A(n8189), .B(n19300), .Z(n8191) );
  XNOR U20726 ( .A(q[3]), .B(DB[1548]), .Z(n19300) );
  XNOR U20727 ( .A(q[2]), .B(DB[1547]), .Z(n8189) );
  XOR U20728 ( .A(n19301), .B(n8087), .Z(n8015) );
  XOR U20729 ( .A(n19302), .B(n8079), .Z(n8087) );
  XOR U20730 ( .A(n19303), .B(n8068), .Z(n8079) );
  XNOR U20731 ( .A(q[14]), .B(DB[1574]), .Z(n8068) );
  IV U20732 ( .A(n8067), .Z(n19303) );
  XNOR U20733 ( .A(n8065), .B(n19304), .Z(n8067) );
  XNOR U20734 ( .A(q[13]), .B(DB[1573]), .Z(n19304) );
  XNOR U20735 ( .A(q[12]), .B(DB[1572]), .Z(n8065) );
  IV U20736 ( .A(n8078), .Z(n19302) );
  XOR U20737 ( .A(n19305), .B(n19306), .Z(n8078) );
  XNOR U20738 ( .A(n8074), .B(n8076), .Z(n19306) );
  XNOR U20739 ( .A(q[8]), .B(DB[1568]), .Z(n8076) );
  XNOR U20740 ( .A(q[11]), .B(DB[1571]), .Z(n8074) );
  IV U20741 ( .A(n8073), .Z(n19305) );
  XNOR U20742 ( .A(n8071), .B(n19307), .Z(n8073) );
  XNOR U20743 ( .A(q[10]), .B(DB[1570]), .Z(n19307) );
  XNOR U20744 ( .A(q[9]), .B(DB[1569]), .Z(n8071) );
  IV U20745 ( .A(n8086), .Z(n19301) );
  XOR U20746 ( .A(n19308), .B(n19309), .Z(n8086) );
  XNOR U20747 ( .A(n8103), .B(n8084), .Z(n19309) );
  XNOR U20748 ( .A(q[0]), .B(DB[1560]), .Z(n8084) );
  XOR U20749 ( .A(n19310), .B(n8092), .Z(n8103) );
  XNOR U20750 ( .A(q[7]), .B(DB[1567]), .Z(n8092) );
  IV U20751 ( .A(n8091), .Z(n19310) );
  XNOR U20752 ( .A(n8089), .B(n19311), .Z(n8091) );
  XNOR U20753 ( .A(q[6]), .B(DB[1566]), .Z(n19311) );
  XNOR U20754 ( .A(q[5]), .B(DB[1565]), .Z(n8089) );
  IV U20755 ( .A(n8102), .Z(n19308) );
  XOR U20756 ( .A(n19312), .B(n19313), .Z(n8102) );
  XNOR U20757 ( .A(n8098), .B(n8100), .Z(n19313) );
  XNOR U20758 ( .A(q[1]), .B(DB[1561]), .Z(n8100) );
  XNOR U20759 ( .A(q[4]), .B(DB[1564]), .Z(n8098) );
  IV U20760 ( .A(n8097), .Z(n19312) );
  XNOR U20761 ( .A(n8095), .B(n19314), .Z(n8097) );
  XNOR U20762 ( .A(q[3]), .B(DB[1563]), .Z(n19314) );
  XNOR U20763 ( .A(q[2]), .B(DB[1562]), .Z(n8095) );
  XOR U20764 ( .A(n19315), .B(n7993), .Z(n7921) );
  XOR U20765 ( .A(n19316), .B(n7985), .Z(n7993) );
  XOR U20766 ( .A(n19317), .B(n7974), .Z(n7985) );
  XNOR U20767 ( .A(q[14]), .B(DB[1589]), .Z(n7974) );
  IV U20768 ( .A(n7973), .Z(n19317) );
  XNOR U20769 ( .A(n7971), .B(n19318), .Z(n7973) );
  XNOR U20770 ( .A(q[13]), .B(DB[1588]), .Z(n19318) );
  XNOR U20771 ( .A(q[12]), .B(DB[1587]), .Z(n7971) );
  IV U20772 ( .A(n7984), .Z(n19316) );
  XOR U20773 ( .A(n19319), .B(n19320), .Z(n7984) );
  XNOR U20774 ( .A(n7980), .B(n7982), .Z(n19320) );
  XNOR U20775 ( .A(q[8]), .B(DB[1583]), .Z(n7982) );
  XNOR U20776 ( .A(q[11]), .B(DB[1586]), .Z(n7980) );
  IV U20777 ( .A(n7979), .Z(n19319) );
  XNOR U20778 ( .A(n7977), .B(n19321), .Z(n7979) );
  XNOR U20779 ( .A(q[10]), .B(DB[1585]), .Z(n19321) );
  XNOR U20780 ( .A(q[9]), .B(DB[1584]), .Z(n7977) );
  IV U20781 ( .A(n7992), .Z(n19315) );
  XOR U20782 ( .A(n19322), .B(n19323), .Z(n7992) );
  XNOR U20783 ( .A(n8009), .B(n7990), .Z(n19323) );
  XNOR U20784 ( .A(q[0]), .B(DB[1575]), .Z(n7990) );
  XOR U20785 ( .A(n19324), .B(n7998), .Z(n8009) );
  XNOR U20786 ( .A(q[7]), .B(DB[1582]), .Z(n7998) );
  IV U20787 ( .A(n7997), .Z(n19324) );
  XNOR U20788 ( .A(n7995), .B(n19325), .Z(n7997) );
  XNOR U20789 ( .A(q[6]), .B(DB[1581]), .Z(n19325) );
  XNOR U20790 ( .A(q[5]), .B(DB[1580]), .Z(n7995) );
  IV U20791 ( .A(n8008), .Z(n19322) );
  XOR U20792 ( .A(n19326), .B(n19327), .Z(n8008) );
  XNOR U20793 ( .A(n8004), .B(n8006), .Z(n19327) );
  XNOR U20794 ( .A(q[1]), .B(DB[1576]), .Z(n8006) );
  XNOR U20795 ( .A(q[4]), .B(DB[1579]), .Z(n8004) );
  IV U20796 ( .A(n8003), .Z(n19326) );
  XNOR U20797 ( .A(n8001), .B(n19328), .Z(n8003) );
  XNOR U20798 ( .A(q[3]), .B(DB[1578]), .Z(n19328) );
  XNOR U20799 ( .A(q[2]), .B(DB[1577]), .Z(n8001) );
  XOR U20800 ( .A(n19329), .B(n7899), .Z(n7827) );
  XOR U20801 ( .A(n19330), .B(n7891), .Z(n7899) );
  XOR U20802 ( .A(n19331), .B(n7880), .Z(n7891) );
  XNOR U20803 ( .A(q[14]), .B(DB[1604]), .Z(n7880) );
  IV U20804 ( .A(n7879), .Z(n19331) );
  XNOR U20805 ( .A(n7877), .B(n19332), .Z(n7879) );
  XNOR U20806 ( .A(q[13]), .B(DB[1603]), .Z(n19332) );
  XNOR U20807 ( .A(q[12]), .B(DB[1602]), .Z(n7877) );
  IV U20808 ( .A(n7890), .Z(n19330) );
  XOR U20809 ( .A(n19333), .B(n19334), .Z(n7890) );
  XNOR U20810 ( .A(n7886), .B(n7888), .Z(n19334) );
  XNOR U20811 ( .A(q[8]), .B(DB[1598]), .Z(n7888) );
  XNOR U20812 ( .A(q[11]), .B(DB[1601]), .Z(n7886) );
  IV U20813 ( .A(n7885), .Z(n19333) );
  XNOR U20814 ( .A(n7883), .B(n19335), .Z(n7885) );
  XNOR U20815 ( .A(q[10]), .B(DB[1600]), .Z(n19335) );
  XNOR U20816 ( .A(q[9]), .B(DB[1599]), .Z(n7883) );
  IV U20817 ( .A(n7898), .Z(n19329) );
  XOR U20818 ( .A(n19336), .B(n19337), .Z(n7898) );
  XNOR U20819 ( .A(n7915), .B(n7896), .Z(n19337) );
  XNOR U20820 ( .A(q[0]), .B(DB[1590]), .Z(n7896) );
  XOR U20821 ( .A(n19338), .B(n7904), .Z(n7915) );
  XNOR U20822 ( .A(q[7]), .B(DB[1597]), .Z(n7904) );
  IV U20823 ( .A(n7903), .Z(n19338) );
  XNOR U20824 ( .A(n7901), .B(n19339), .Z(n7903) );
  XNOR U20825 ( .A(q[6]), .B(DB[1596]), .Z(n19339) );
  XNOR U20826 ( .A(q[5]), .B(DB[1595]), .Z(n7901) );
  IV U20827 ( .A(n7914), .Z(n19336) );
  XOR U20828 ( .A(n19340), .B(n19341), .Z(n7914) );
  XNOR U20829 ( .A(n7910), .B(n7912), .Z(n19341) );
  XNOR U20830 ( .A(q[1]), .B(DB[1591]), .Z(n7912) );
  XNOR U20831 ( .A(q[4]), .B(DB[1594]), .Z(n7910) );
  IV U20832 ( .A(n7909), .Z(n19340) );
  XNOR U20833 ( .A(n7907), .B(n19342), .Z(n7909) );
  XNOR U20834 ( .A(q[3]), .B(DB[1593]), .Z(n19342) );
  XNOR U20835 ( .A(q[2]), .B(DB[1592]), .Z(n7907) );
  XOR U20836 ( .A(n19343), .B(n7805), .Z(n7733) );
  XOR U20837 ( .A(n19344), .B(n7797), .Z(n7805) );
  XOR U20838 ( .A(n19345), .B(n7786), .Z(n7797) );
  XNOR U20839 ( .A(q[14]), .B(DB[1619]), .Z(n7786) );
  IV U20840 ( .A(n7785), .Z(n19345) );
  XNOR U20841 ( .A(n7783), .B(n19346), .Z(n7785) );
  XNOR U20842 ( .A(q[13]), .B(DB[1618]), .Z(n19346) );
  XNOR U20843 ( .A(q[12]), .B(DB[1617]), .Z(n7783) );
  IV U20844 ( .A(n7796), .Z(n19344) );
  XOR U20845 ( .A(n19347), .B(n19348), .Z(n7796) );
  XNOR U20846 ( .A(n7792), .B(n7794), .Z(n19348) );
  XNOR U20847 ( .A(q[8]), .B(DB[1613]), .Z(n7794) );
  XNOR U20848 ( .A(q[11]), .B(DB[1616]), .Z(n7792) );
  IV U20849 ( .A(n7791), .Z(n19347) );
  XNOR U20850 ( .A(n7789), .B(n19349), .Z(n7791) );
  XNOR U20851 ( .A(q[10]), .B(DB[1615]), .Z(n19349) );
  XNOR U20852 ( .A(q[9]), .B(DB[1614]), .Z(n7789) );
  IV U20853 ( .A(n7804), .Z(n19343) );
  XOR U20854 ( .A(n19350), .B(n19351), .Z(n7804) );
  XNOR U20855 ( .A(n7821), .B(n7802), .Z(n19351) );
  XNOR U20856 ( .A(q[0]), .B(DB[1605]), .Z(n7802) );
  XOR U20857 ( .A(n19352), .B(n7810), .Z(n7821) );
  XNOR U20858 ( .A(q[7]), .B(DB[1612]), .Z(n7810) );
  IV U20859 ( .A(n7809), .Z(n19352) );
  XNOR U20860 ( .A(n7807), .B(n19353), .Z(n7809) );
  XNOR U20861 ( .A(q[6]), .B(DB[1611]), .Z(n19353) );
  XNOR U20862 ( .A(q[5]), .B(DB[1610]), .Z(n7807) );
  IV U20863 ( .A(n7820), .Z(n19350) );
  XOR U20864 ( .A(n19354), .B(n19355), .Z(n7820) );
  XNOR U20865 ( .A(n7816), .B(n7818), .Z(n19355) );
  XNOR U20866 ( .A(q[1]), .B(DB[1606]), .Z(n7818) );
  XNOR U20867 ( .A(q[4]), .B(DB[1609]), .Z(n7816) );
  IV U20868 ( .A(n7815), .Z(n19354) );
  XNOR U20869 ( .A(n7813), .B(n19356), .Z(n7815) );
  XNOR U20870 ( .A(q[3]), .B(DB[1608]), .Z(n19356) );
  XNOR U20871 ( .A(q[2]), .B(DB[1607]), .Z(n7813) );
  XOR U20872 ( .A(n19357), .B(n7711), .Z(n7639) );
  XOR U20873 ( .A(n19358), .B(n7703), .Z(n7711) );
  XOR U20874 ( .A(n19359), .B(n7692), .Z(n7703) );
  XNOR U20875 ( .A(q[14]), .B(DB[1634]), .Z(n7692) );
  IV U20876 ( .A(n7691), .Z(n19359) );
  XNOR U20877 ( .A(n7689), .B(n19360), .Z(n7691) );
  XNOR U20878 ( .A(q[13]), .B(DB[1633]), .Z(n19360) );
  XNOR U20879 ( .A(q[12]), .B(DB[1632]), .Z(n7689) );
  IV U20880 ( .A(n7702), .Z(n19358) );
  XOR U20881 ( .A(n19361), .B(n19362), .Z(n7702) );
  XNOR U20882 ( .A(n7698), .B(n7700), .Z(n19362) );
  XNOR U20883 ( .A(q[8]), .B(DB[1628]), .Z(n7700) );
  XNOR U20884 ( .A(q[11]), .B(DB[1631]), .Z(n7698) );
  IV U20885 ( .A(n7697), .Z(n19361) );
  XNOR U20886 ( .A(n7695), .B(n19363), .Z(n7697) );
  XNOR U20887 ( .A(q[10]), .B(DB[1630]), .Z(n19363) );
  XNOR U20888 ( .A(q[9]), .B(DB[1629]), .Z(n7695) );
  IV U20889 ( .A(n7710), .Z(n19357) );
  XOR U20890 ( .A(n19364), .B(n19365), .Z(n7710) );
  XNOR U20891 ( .A(n7727), .B(n7708), .Z(n19365) );
  XNOR U20892 ( .A(q[0]), .B(DB[1620]), .Z(n7708) );
  XOR U20893 ( .A(n19366), .B(n7716), .Z(n7727) );
  XNOR U20894 ( .A(q[7]), .B(DB[1627]), .Z(n7716) );
  IV U20895 ( .A(n7715), .Z(n19366) );
  XNOR U20896 ( .A(n7713), .B(n19367), .Z(n7715) );
  XNOR U20897 ( .A(q[6]), .B(DB[1626]), .Z(n19367) );
  XNOR U20898 ( .A(q[5]), .B(DB[1625]), .Z(n7713) );
  IV U20899 ( .A(n7726), .Z(n19364) );
  XOR U20900 ( .A(n19368), .B(n19369), .Z(n7726) );
  XNOR U20901 ( .A(n7722), .B(n7724), .Z(n19369) );
  XNOR U20902 ( .A(q[1]), .B(DB[1621]), .Z(n7724) );
  XNOR U20903 ( .A(q[4]), .B(DB[1624]), .Z(n7722) );
  IV U20904 ( .A(n7721), .Z(n19368) );
  XNOR U20905 ( .A(n7719), .B(n19370), .Z(n7721) );
  XNOR U20906 ( .A(q[3]), .B(DB[1623]), .Z(n19370) );
  XNOR U20907 ( .A(q[2]), .B(DB[1622]), .Z(n7719) );
  XOR U20908 ( .A(n19371), .B(n7617), .Z(n7545) );
  XOR U20909 ( .A(n19372), .B(n7609), .Z(n7617) );
  XOR U20910 ( .A(n19373), .B(n7598), .Z(n7609) );
  XNOR U20911 ( .A(q[14]), .B(DB[1649]), .Z(n7598) );
  IV U20912 ( .A(n7597), .Z(n19373) );
  XNOR U20913 ( .A(n7595), .B(n19374), .Z(n7597) );
  XNOR U20914 ( .A(q[13]), .B(DB[1648]), .Z(n19374) );
  XNOR U20915 ( .A(q[12]), .B(DB[1647]), .Z(n7595) );
  IV U20916 ( .A(n7608), .Z(n19372) );
  XOR U20917 ( .A(n19375), .B(n19376), .Z(n7608) );
  XNOR U20918 ( .A(n7604), .B(n7606), .Z(n19376) );
  XNOR U20919 ( .A(q[8]), .B(DB[1643]), .Z(n7606) );
  XNOR U20920 ( .A(q[11]), .B(DB[1646]), .Z(n7604) );
  IV U20921 ( .A(n7603), .Z(n19375) );
  XNOR U20922 ( .A(n7601), .B(n19377), .Z(n7603) );
  XNOR U20923 ( .A(q[10]), .B(DB[1645]), .Z(n19377) );
  XNOR U20924 ( .A(q[9]), .B(DB[1644]), .Z(n7601) );
  IV U20925 ( .A(n7616), .Z(n19371) );
  XOR U20926 ( .A(n19378), .B(n19379), .Z(n7616) );
  XNOR U20927 ( .A(n7633), .B(n7614), .Z(n19379) );
  XNOR U20928 ( .A(q[0]), .B(DB[1635]), .Z(n7614) );
  XOR U20929 ( .A(n19380), .B(n7622), .Z(n7633) );
  XNOR U20930 ( .A(q[7]), .B(DB[1642]), .Z(n7622) );
  IV U20931 ( .A(n7621), .Z(n19380) );
  XNOR U20932 ( .A(n7619), .B(n19381), .Z(n7621) );
  XNOR U20933 ( .A(q[6]), .B(DB[1641]), .Z(n19381) );
  XNOR U20934 ( .A(q[5]), .B(DB[1640]), .Z(n7619) );
  IV U20935 ( .A(n7632), .Z(n19378) );
  XOR U20936 ( .A(n19382), .B(n19383), .Z(n7632) );
  XNOR U20937 ( .A(n7628), .B(n7630), .Z(n19383) );
  XNOR U20938 ( .A(q[1]), .B(DB[1636]), .Z(n7630) );
  XNOR U20939 ( .A(q[4]), .B(DB[1639]), .Z(n7628) );
  IV U20940 ( .A(n7627), .Z(n19382) );
  XNOR U20941 ( .A(n7625), .B(n19384), .Z(n7627) );
  XNOR U20942 ( .A(q[3]), .B(DB[1638]), .Z(n19384) );
  XNOR U20943 ( .A(q[2]), .B(DB[1637]), .Z(n7625) );
  XOR U20944 ( .A(n19385), .B(n7523), .Z(n7451) );
  XOR U20945 ( .A(n19386), .B(n7515), .Z(n7523) );
  XOR U20946 ( .A(n19387), .B(n7504), .Z(n7515) );
  XNOR U20947 ( .A(q[14]), .B(DB[1664]), .Z(n7504) );
  IV U20948 ( .A(n7503), .Z(n19387) );
  XNOR U20949 ( .A(n7501), .B(n19388), .Z(n7503) );
  XNOR U20950 ( .A(q[13]), .B(DB[1663]), .Z(n19388) );
  XNOR U20951 ( .A(q[12]), .B(DB[1662]), .Z(n7501) );
  IV U20952 ( .A(n7514), .Z(n19386) );
  XOR U20953 ( .A(n19389), .B(n19390), .Z(n7514) );
  XNOR U20954 ( .A(n7510), .B(n7512), .Z(n19390) );
  XNOR U20955 ( .A(q[8]), .B(DB[1658]), .Z(n7512) );
  XNOR U20956 ( .A(q[11]), .B(DB[1661]), .Z(n7510) );
  IV U20957 ( .A(n7509), .Z(n19389) );
  XNOR U20958 ( .A(n7507), .B(n19391), .Z(n7509) );
  XNOR U20959 ( .A(q[10]), .B(DB[1660]), .Z(n19391) );
  XNOR U20960 ( .A(q[9]), .B(DB[1659]), .Z(n7507) );
  IV U20961 ( .A(n7522), .Z(n19385) );
  XOR U20962 ( .A(n19392), .B(n19393), .Z(n7522) );
  XNOR U20963 ( .A(n7539), .B(n7520), .Z(n19393) );
  XNOR U20964 ( .A(q[0]), .B(DB[1650]), .Z(n7520) );
  XOR U20965 ( .A(n19394), .B(n7528), .Z(n7539) );
  XNOR U20966 ( .A(q[7]), .B(DB[1657]), .Z(n7528) );
  IV U20967 ( .A(n7527), .Z(n19394) );
  XNOR U20968 ( .A(n7525), .B(n19395), .Z(n7527) );
  XNOR U20969 ( .A(q[6]), .B(DB[1656]), .Z(n19395) );
  XNOR U20970 ( .A(q[5]), .B(DB[1655]), .Z(n7525) );
  IV U20971 ( .A(n7538), .Z(n19392) );
  XOR U20972 ( .A(n19396), .B(n19397), .Z(n7538) );
  XNOR U20973 ( .A(n7534), .B(n7536), .Z(n19397) );
  XNOR U20974 ( .A(q[1]), .B(DB[1651]), .Z(n7536) );
  XNOR U20975 ( .A(q[4]), .B(DB[1654]), .Z(n7534) );
  IV U20976 ( .A(n7533), .Z(n19396) );
  XNOR U20977 ( .A(n7531), .B(n19398), .Z(n7533) );
  XNOR U20978 ( .A(q[3]), .B(DB[1653]), .Z(n19398) );
  XNOR U20979 ( .A(q[2]), .B(DB[1652]), .Z(n7531) );
  XOR U20980 ( .A(n19399), .B(n7429), .Z(n7357) );
  XOR U20981 ( .A(n19400), .B(n7421), .Z(n7429) );
  XOR U20982 ( .A(n19401), .B(n7410), .Z(n7421) );
  XNOR U20983 ( .A(q[14]), .B(DB[1679]), .Z(n7410) );
  IV U20984 ( .A(n7409), .Z(n19401) );
  XNOR U20985 ( .A(n7407), .B(n19402), .Z(n7409) );
  XNOR U20986 ( .A(q[13]), .B(DB[1678]), .Z(n19402) );
  XNOR U20987 ( .A(q[12]), .B(DB[1677]), .Z(n7407) );
  IV U20988 ( .A(n7420), .Z(n19400) );
  XOR U20989 ( .A(n19403), .B(n19404), .Z(n7420) );
  XNOR U20990 ( .A(n7416), .B(n7418), .Z(n19404) );
  XNOR U20991 ( .A(q[8]), .B(DB[1673]), .Z(n7418) );
  XNOR U20992 ( .A(q[11]), .B(DB[1676]), .Z(n7416) );
  IV U20993 ( .A(n7415), .Z(n19403) );
  XNOR U20994 ( .A(n7413), .B(n19405), .Z(n7415) );
  XNOR U20995 ( .A(q[10]), .B(DB[1675]), .Z(n19405) );
  XNOR U20996 ( .A(q[9]), .B(DB[1674]), .Z(n7413) );
  IV U20997 ( .A(n7428), .Z(n19399) );
  XOR U20998 ( .A(n19406), .B(n19407), .Z(n7428) );
  XNOR U20999 ( .A(n7445), .B(n7426), .Z(n19407) );
  XNOR U21000 ( .A(q[0]), .B(DB[1665]), .Z(n7426) );
  XOR U21001 ( .A(n19408), .B(n7434), .Z(n7445) );
  XNOR U21002 ( .A(q[7]), .B(DB[1672]), .Z(n7434) );
  IV U21003 ( .A(n7433), .Z(n19408) );
  XNOR U21004 ( .A(n7431), .B(n19409), .Z(n7433) );
  XNOR U21005 ( .A(q[6]), .B(DB[1671]), .Z(n19409) );
  XNOR U21006 ( .A(q[5]), .B(DB[1670]), .Z(n7431) );
  IV U21007 ( .A(n7444), .Z(n19406) );
  XOR U21008 ( .A(n19410), .B(n19411), .Z(n7444) );
  XNOR U21009 ( .A(n7440), .B(n7442), .Z(n19411) );
  XNOR U21010 ( .A(q[1]), .B(DB[1666]), .Z(n7442) );
  XNOR U21011 ( .A(q[4]), .B(DB[1669]), .Z(n7440) );
  IV U21012 ( .A(n7439), .Z(n19410) );
  XNOR U21013 ( .A(n7437), .B(n19412), .Z(n7439) );
  XNOR U21014 ( .A(q[3]), .B(DB[1668]), .Z(n19412) );
  XNOR U21015 ( .A(q[2]), .B(DB[1667]), .Z(n7437) );
  XOR U21016 ( .A(n19413), .B(n7335), .Z(n7263) );
  XOR U21017 ( .A(n19414), .B(n7327), .Z(n7335) );
  XOR U21018 ( .A(n19415), .B(n7316), .Z(n7327) );
  XNOR U21019 ( .A(q[14]), .B(DB[1694]), .Z(n7316) );
  IV U21020 ( .A(n7315), .Z(n19415) );
  XNOR U21021 ( .A(n7313), .B(n19416), .Z(n7315) );
  XNOR U21022 ( .A(q[13]), .B(DB[1693]), .Z(n19416) );
  XNOR U21023 ( .A(q[12]), .B(DB[1692]), .Z(n7313) );
  IV U21024 ( .A(n7326), .Z(n19414) );
  XOR U21025 ( .A(n19417), .B(n19418), .Z(n7326) );
  XNOR U21026 ( .A(n7322), .B(n7324), .Z(n19418) );
  XNOR U21027 ( .A(q[8]), .B(DB[1688]), .Z(n7324) );
  XNOR U21028 ( .A(q[11]), .B(DB[1691]), .Z(n7322) );
  IV U21029 ( .A(n7321), .Z(n19417) );
  XNOR U21030 ( .A(n7319), .B(n19419), .Z(n7321) );
  XNOR U21031 ( .A(q[10]), .B(DB[1690]), .Z(n19419) );
  XNOR U21032 ( .A(q[9]), .B(DB[1689]), .Z(n7319) );
  IV U21033 ( .A(n7334), .Z(n19413) );
  XOR U21034 ( .A(n19420), .B(n19421), .Z(n7334) );
  XNOR U21035 ( .A(n7351), .B(n7332), .Z(n19421) );
  XNOR U21036 ( .A(q[0]), .B(DB[1680]), .Z(n7332) );
  XOR U21037 ( .A(n19422), .B(n7340), .Z(n7351) );
  XNOR U21038 ( .A(q[7]), .B(DB[1687]), .Z(n7340) );
  IV U21039 ( .A(n7339), .Z(n19422) );
  XNOR U21040 ( .A(n7337), .B(n19423), .Z(n7339) );
  XNOR U21041 ( .A(q[6]), .B(DB[1686]), .Z(n19423) );
  XNOR U21042 ( .A(q[5]), .B(DB[1685]), .Z(n7337) );
  IV U21043 ( .A(n7350), .Z(n19420) );
  XOR U21044 ( .A(n19424), .B(n19425), .Z(n7350) );
  XNOR U21045 ( .A(n7346), .B(n7348), .Z(n19425) );
  XNOR U21046 ( .A(q[1]), .B(DB[1681]), .Z(n7348) );
  XNOR U21047 ( .A(q[4]), .B(DB[1684]), .Z(n7346) );
  IV U21048 ( .A(n7345), .Z(n19424) );
  XNOR U21049 ( .A(n7343), .B(n19426), .Z(n7345) );
  XNOR U21050 ( .A(q[3]), .B(DB[1683]), .Z(n19426) );
  XNOR U21051 ( .A(q[2]), .B(DB[1682]), .Z(n7343) );
  XOR U21052 ( .A(n19427), .B(n7241), .Z(n7169) );
  XOR U21053 ( .A(n19428), .B(n7233), .Z(n7241) );
  XOR U21054 ( .A(n19429), .B(n7222), .Z(n7233) );
  XNOR U21055 ( .A(q[14]), .B(DB[1709]), .Z(n7222) );
  IV U21056 ( .A(n7221), .Z(n19429) );
  XNOR U21057 ( .A(n7219), .B(n19430), .Z(n7221) );
  XNOR U21058 ( .A(q[13]), .B(DB[1708]), .Z(n19430) );
  XNOR U21059 ( .A(q[12]), .B(DB[1707]), .Z(n7219) );
  IV U21060 ( .A(n7232), .Z(n19428) );
  XOR U21061 ( .A(n19431), .B(n19432), .Z(n7232) );
  XNOR U21062 ( .A(n7228), .B(n7230), .Z(n19432) );
  XNOR U21063 ( .A(q[8]), .B(DB[1703]), .Z(n7230) );
  XNOR U21064 ( .A(q[11]), .B(DB[1706]), .Z(n7228) );
  IV U21065 ( .A(n7227), .Z(n19431) );
  XNOR U21066 ( .A(n7225), .B(n19433), .Z(n7227) );
  XNOR U21067 ( .A(q[10]), .B(DB[1705]), .Z(n19433) );
  XNOR U21068 ( .A(q[9]), .B(DB[1704]), .Z(n7225) );
  IV U21069 ( .A(n7240), .Z(n19427) );
  XOR U21070 ( .A(n19434), .B(n19435), .Z(n7240) );
  XNOR U21071 ( .A(n7257), .B(n7238), .Z(n19435) );
  XNOR U21072 ( .A(q[0]), .B(DB[1695]), .Z(n7238) );
  XOR U21073 ( .A(n19436), .B(n7246), .Z(n7257) );
  XNOR U21074 ( .A(q[7]), .B(DB[1702]), .Z(n7246) );
  IV U21075 ( .A(n7245), .Z(n19436) );
  XNOR U21076 ( .A(n7243), .B(n19437), .Z(n7245) );
  XNOR U21077 ( .A(q[6]), .B(DB[1701]), .Z(n19437) );
  XNOR U21078 ( .A(q[5]), .B(DB[1700]), .Z(n7243) );
  IV U21079 ( .A(n7256), .Z(n19434) );
  XOR U21080 ( .A(n19438), .B(n19439), .Z(n7256) );
  XNOR U21081 ( .A(n7252), .B(n7254), .Z(n19439) );
  XNOR U21082 ( .A(q[1]), .B(DB[1696]), .Z(n7254) );
  XNOR U21083 ( .A(q[4]), .B(DB[1699]), .Z(n7252) );
  IV U21084 ( .A(n7251), .Z(n19438) );
  XNOR U21085 ( .A(n7249), .B(n19440), .Z(n7251) );
  XNOR U21086 ( .A(q[3]), .B(DB[1698]), .Z(n19440) );
  XNOR U21087 ( .A(q[2]), .B(DB[1697]), .Z(n7249) );
  XOR U21088 ( .A(n19441), .B(n7147), .Z(n7075) );
  XOR U21089 ( .A(n19442), .B(n7139), .Z(n7147) );
  XOR U21090 ( .A(n19443), .B(n7128), .Z(n7139) );
  XNOR U21091 ( .A(q[14]), .B(DB[1724]), .Z(n7128) );
  IV U21092 ( .A(n7127), .Z(n19443) );
  XNOR U21093 ( .A(n7125), .B(n19444), .Z(n7127) );
  XNOR U21094 ( .A(q[13]), .B(DB[1723]), .Z(n19444) );
  XNOR U21095 ( .A(q[12]), .B(DB[1722]), .Z(n7125) );
  IV U21096 ( .A(n7138), .Z(n19442) );
  XOR U21097 ( .A(n19445), .B(n19446), .Z(n7138) );
  XNOR U21098 ( .A(n7134), .B(n7136), .Z(n19446) );
  XNOR U21099 ( .A(q[8]), .B(DB[1718]), .Z(n7136) );
  XNOR U21100 ( .A(q[11]), .B(DB[1721]), .Z(n7134) );
  IV U21101 ( .A(n7133), .Z(n19445) );
  XNOR U21102 ( .A(n7131), .B(n19447), .Z(n7133) );
  XNOR U21103 ( .A(q[10]), .B(DB[1720]), .Z(n19447) );
  XNOR U21104 ( .A(q[9]), .B(DB[1719]), .Z(n7131) );
  IV U21105 ( .A(n7146), .Z(n19441) );
  XOR U21106 ( .A(n19448), .B(n19449), .Z(n7146) );
  XNOR U21107 ( .A(n7163), .B(n7144), .Z(n19449) );
  XNOR U21108 ( .A(q[0]), .B(DB[1710]), .Z(n7144) );
  XOR U21109 ( .A(n19450), .B(n7152), .Z(n7163) );
  XNOR U21110 ( .A(q[7]), .B(DB[1717]), .Z(n7152) );
  IV U21111 ( .A(n7151), .Z(n19450) );
  XNOR U21112 ( .A(n7149), .B(n19451), .Z(n7151) );
  XNOR U21113 ( .A(q[6]), .B(DB[1716]), .Z(n19451) );
  XNOR U21114 ( .A(q[5]), .B(DB[1715]), .Z(n7149) );
  IV U21115 ( .A(n7162), .Z(n19448) );
  XOR U21116 ( .A(n19452), .B(n19453), .Z(n7162) );
  XNOR U21117 ( .A(n7158), .B(n7160), .Z(n19453) );
  XNOR U21118 ( .A(q[1]), .B(DB[1711]), .Z(n7160) );
  XNOR U21119 ( .A(q[4]), .B(DB[1714]), .Z(n7158) );
  IV U21120 ( .A(n7157), .Z(n19452) );
  XNOR U21121 ( .A(n7155), .B(n19454), .Z(n7157) );
  XNOR U21122 ( .A(q[3]), .B(DB[1713]), .Z(n19454) );
  XNOR U21123 ( .A(q[2]), .B(DB[1712]), .Z(n7155) );
  XOR U21124 ( .A(n19455), .B(n7053), .Z(n6981) );
  XOR U21125 ( .A(n19456), .B(n7045), .Z(n7053) );
  XOR U21126 ( .A(n19457), .B(n7034), .Z(n7045) );
  XNOR U21127 ( .A(q[14]), .B(DB[1739]), .Z(n7034) );
  IV U21128 ( .A(n7033), .Z(n19457) );
  XNOR U21129 ( .A(n7031), .B(n19458), .Z(n7033) );
  XNOR U21130 ( .A(q[13]), .B(DB[1738]), .Z(n19458) );
  XNOR U21131 ( .A(q[12]), .B(DB[1737]), .Z(n7031) );
  IV U21132 ( .A(n7044), .Z(n19456) );
  XOR U21133 ( .A(n19459), .B(n19460), .Z(n7044) );
  XNOR U21134 ( .A(n7040), .B(n7042), .Z(n19460) );
  XNOR U21135 ( .A(q[8]), .B(DB[1733]), .Z(n7042) );
  XNOR U21136 ( .A(q[11]), .B(DB[1736]), .Z(n7040) );
  IV U21137 ( .A(n7039), .Z(n19459) );
  XNOR U21138 ( .A(n7037), .B(n19461), .Z(n7039) );
  XNOR U21139 ( .A(q[10]), .B(DB[1735]), .Z(n19461) );
  XNOR U21140 ( .A(q[9]), .B(DB[1734]), .Z(n7037) );
  IV U21141 ( .A(n7052), .Z(n19455) );
  XOR U21142 ( .A(n19462), .B(n19463), .Z(n7052) );
  XNOR U21143 ( .A(n7069), .B(n7050), .Z(n19463) );
  XNOR U21144 ( .A(q[0]), .B(DB[1725]), .Z(n7050) );
  XOR U21145 ( .A(n19464), .B(n7058), .Z(n7069) );
  XNOR U21146 ( .A(q[7]), .B(DB[1732]), .Z(n7058) );
  IV U21147 ( .A(n7057), .Z(n19464) );
  XNOR U21148 ( .A(n7055), .B(n19465), .Z(n7057) );
  XNOR U21149 ( .A(q[6]), .B(DB[1731]), .Z(n19465) );
  XNOR U21150 ( .A(q[5]), .B(DB[1730]), .Z(n7055) );
  IV U21151 ( .A(n7068), .Z(n19462) );
  XOR U21152 ( .A(n19466), .B(n19467), .Z(n7068) );
  XNOR U21153 ( .A(n7064), .B(n7066), .Z(n19467) );
  XNOR U21154 ( .A(q[1]), .B(DB[1726]), .Z(n7066) );
  XNOR U21155 ( .A(q[4]), .B(DB[1729]), .Z(n7064) );
  IV U21156 ( .A(n7063), .Z(n19466) );
  XNOR U21157 ( .A(n7061), .B(n19468), .Z(n7063) );
  XNOR U21158 ( .A(q[3]), .B(DB[1728]), .Z(n19468) );
  XNOR U21159 ( .A(q[2]), .B(DB[1727]), .Z(n7061) );
  XOR U21160 ( .A(n19469), .B(n6959), .Z(n6887) );
  XOR U21161 ( .A(n19470), .B(n6951), .Z(n6959) );
  XOR U21162 ( .A(n19471), .B(n6940), .Z(n6951) );
  XNOR U21163 ( .A(q[14]), .B(DB[1754]), .Z(n6940) );
  IV U21164 ( .A(n6939), .Z(n19471) );
  XNOR U21165 ( .A(n6937), .B(n19472), .Z(n6939) );
  XNOR U21166 ( .A(q[13]), .B(DB[1753]), .Z(n19472) );
  XNOR U21167 ( .A(q[12]), .B(DB[1752]), .Z(n6937) );
  IV U21168 ( .A(n6950), .Z(n19470) );
  XOR U21169 ( .A(n19473), .B(n19474), .Z(n6950) );
  XNOR U21170 ( .A(n6946), .B(n6948), .Z(n19474) );
  XNOR U21171 ( .A(q[8]), .B(DB[1748]), .Z(n6948) );
  XNOR U21172 ( .A(q[11]), .B(DB[1751]), .Z(n6946) );
  IV U21173 ( .A(n6945), .Z(n19473) );
  XNOR U21174 ( .A(n6943), .B(n19475), .Z(n6945) );
  XNOR U21175 ( .A(q[10]), .B(DB[1750]), .Z(n19475) );
  XNOR U21176 ( .A(q[9]), .B(DB[1749]), .Z(n6943) );
  IV U21177 ( .A(n6958), .Z(n19469) );
  XOR U21178 ( .A(n19476), .B(n19477), .Z(n6958) );
  XNOR U21179 ( .A(n6975), .B(n6956), .Z(n19477) );
  XNOR U21180 ( .A(q[0]), .B(DB[1740]), .Z(n6956) );
  XOR U21181 ( .A(n19478), .B(n6964), .Z(n6975) );
  XNOR U21182 ( .A(q[7]), .B(DB[1747]), .Z(n6964) );
  IV U21183 ( .A(n6963), .Z(n19478) );
  XNOR U21184 ( .A(n6961), .B(n19479), .Z(n6963) );
  XNOR U21185 ( .A(q[6]), .B(DB[1746]), .Z(n19479) );
  XNOR U21186 ( .A(q[5]), .B(DB[1745]), .Z(n6961) );
  IV U21187 ( .A(n6974), .Z(n19476) );
  XOR U21188 ( .A(n19480), .B(n19481), .Z(n6974) );
  XNOR U21189 ( .A(n6970), .B(n6972), .Z(n19481) );
  XNOR U21190 ( .A(q[1]), .B(DB[1741]), .Z(n6972) );
  XNOR U21191 ( .A(q[4]), .B(DB[1744]), .Z(n6970) );
  IV U21192 ( .A(n6969), .Z(n19480) );
  XNOR U21193 ( .A(n6967), .B(n19482), .Z(n6969) );
  XNOR U21194 ( .A(q[3]), .B(DB[1743]), .Z(n19482) );
  XNOR U21195 ( .A(q[2]), .B(DB[1742]), .Z(n6967) );
  XOR U21196 ( .A(n19483), .B(n6865), .Z(n6793) );
  XOR U21197 ( .A(n19484), .B(n6857), .Z(n6865) );
  XOR U21198 ( .A(n19485), .B(n6846), .Z(n6857) );
  XNOR U21199 ( .A(q[14]), .B(DB[1769]), .Z(n6846) );
  IV U21200 ( .A(n6845), .Z(n19485) );
  XNOR U21201 ( .A(n6843), .B(n19486), .Z(n6845) );
  XNOR U21202 ( .A(q[13]), .B(DB[1768]), .Z(n19486) );
  XNOR U21203 ( .A(q[12]), .B(DB[1767]), .Z(n6843) );
  IV U21204 ( .A(n6856), .Z(n19484) );
  XOR U21205 ( .A(n19487), .B(n19488), .Z(n6856) );
  XNOR U21206 ( .A(n6852), .B(n6854), .Z(n19488) );
  XNOR U21207 ( .A(q[8]), .B(DB[1763]), .Z(n6854) );
  XNOR U21208 ( .A(q[11]), .B(DB[1766]), .Z(n6852) );
  IV U21209 ( .A(n6851), .Z(n19487) );
  XNOR U21210 ( .A(n6849), .B(n19489), .Z(n6851) );
  XNOR U21211 ( .A(q[10]), .B(DB[1765]), .Z(n19489) );
  XNOR U21212 ( .A(q[9]), .B(DB[1764]), .Z(n6849) );
  IV U21213 ( .A(n6864), .Z(n19483) );
  XOR U21214 ( .A(n19490), .B(n19491), .Z(n6864) );
  XNOR U21215 ( .A(n6881), .B(n6862), .Z(n19491) );
  XNOR U21216 ( .A(q[0]), .B(DB[1755]), .Z(n6862) );
  XOR U21217 ( .A(n19492), .B(n6870), .Z(n6881) );
  XNOR U21218 ( .A(q[7]), .B(DB[1762]), .Z(n6870) );
  IV U21219 ( .A(n6869), .Z(n19492) );
  XNOR U21220 ( .A(n6867), .B(n19493), .Z(n6869) );
  XNOR U21221 ( .A(q[6]), .B(DB[1761]), .Z(n19493) );
  XNOR U21222 ( .A(q[5]), .B(DB[1760]), .Z(n6867) );
  IV U21223 ( .A(n6880), .Z(n19490) );
  XOR U21224 ( .A(n19494), .B(n19495), .Z(n6880) );
  XNOR U21225 ( .A(n6876), .B(n6878), .Z(n19495) );
  XNOR U21226 ( .A(q[1]), .B(DB[1756]), .Z(n6878) );
  XNOR U21227 ( .A(q[4]), .B(DB[1759]), .Z(n6876) );
  IV U21228 ( .A(n6875), .Z(n19494) );
  XNOR U21229 ( .A(n6873), .B(n19496), .Z(n6875) );
  XNOR U21230 ( .A(q[3]), .B(DB[1758]), .Z(n19496) );
  XNOR U21231 ( .A(q[2]), .B(DB[1757]), .Z(n6873) );
  XOR U21232 ( .A(n19497), .B(n6771), .Z(n6699) );
  XOR U21233 ( .A(n19498), .B(n6763), .Z(n6771) );
  XOR U21234 ( .A(n19499), .B(n6752), .Z(n6763) );
  XNOR U21235 ( .A(q[14]), .B(DB[1784]), .Z(n6752) );
  IV U21236 ( .A(n6751), .Z(n19499) );
  XNOR U21237 ( .A(n6749), .B(n19500), .Z(n6751) );
  XNOR U21238 ( .A(q[13]), .B(DB[1783]), .Z(n19500) );
  XNOR U21239 ( .A(q[12]), .B(DB[1782]), .Z(n6749) );
  IV U21240 ( .A(n6762), .Z(n19498) );
  XOR U21241 ( .A(n19501), .B(n19502), .Z(n6762) );
  XNOR U21242 ( .A(n6758), .B(n6760), .Z(n19502) );
  XNOR U21243 ( .A(q[8]), .B(DB[1778]), .Z(n6760) );
  XNOR U21244 ( .A(q[11]), .B(DB[1781]), .Z(n6758) );
  IV U21245 ( .A(n6757), .Z(n19501) );
  XNOR U21246 ( .A(n6755), .B(n19503), .Z(n6757) );
  XNOR U21247 ( .A(q[10]), .B(DB[1780]), .Z(n19503) );
  XNOR U21248 ( .A(q[9]), .B(DB[1779]), .Z(n6755) );
  IV U21249 ( .A(n6770), .Z(n19497) );
  XOR U21250 ( .A(n19504), .B(n19505), .Z(n6770) );
  XNOR U21251 ( .A(n6787), .B(n6768), .Z(n19505) );
  XNOR U21252 ( .A(q[0]), .B(DB[1770]), .Z(n6768) );
  XOR U21253 ( .A(n19506), .B(n6776), .Z(n6787) );
  XNOR U21254 ( .A(q[7]), .B(DB[1777]), .Z(n6776) );
  IV U21255 ( .A(n6775), .Z(n19506) );
  XNOR U21256 ( .A(n6773), .B(n19507), .Z(n6775) );
  XNOR U21257 ( .A(q[6]), .B(DB[1776]), .Z(n19507) );
  XNOR U21258 ( .A(q[5]), .B(DB[1775]), .Z(n6773) );
  IV U21259 ( .A(n6786), .Z(n19504) );
  XOR U21260 ( .A(n19508), .B(n19509), .Z(n6786) );
  XNOR U21261 ( .A(n6782), .B(n6784), .Z(n19509) );
  XNOR U21262 ( .A(q[1]), .B(DB[1771]), .Z(n6784) );
  XNOR U21263 ( .A(q[4]), .B(DB[1774]), .Z(n6782) );
  IV U21264 ( .A(n6781), .Z(n19508) );
  XNOR U21265 ( .A(n6779), .B(n19510), .Z(n6781) );
  XNOR U21266 ( .A(q[3]), .B(DB[1773]), .Z(n19510) );
  XNOR U21267 ( .A(q[2]), .B(DB[1772]), .Z(n6779) );
  XOR U21268 ( .A(n19511), .B(n6677), .Z(n6605) );
  XOR U21269 ( .A(n19512), .B(n6669), .Z(n6677) );
  XOR U21270 ( .A(n19513), .B(n6658), .Z(n6669) );
  XNOR U21271 ( .A(q[14]), .B(DB[1799]), .Z(n6658) );
  IV U21272 ( .A(n6657), .Z(n19513) );
  XNOR U21273 ( .A(n6655), .B(n19514), .Z(n6657) );
  XNOR U21274 ( .A(q[13]), .B(DB[1798]), .Z(n19514) );
  XNOR U21275 ( .A(q[12]), .B(DB[1797]), .Z(n6655) );
  IV U21276 ( .A(n6668), .Z(n19512) );
  XOR U21277 ( .A(n19515), .B(n19516), .Z(n6668) );
  XNOR U21278 ( .A(n6664), .B(n6666), .Z(n19516) );
  XNOR U21279 ( .A(q[8]), .B(DB[1793]), .Z(n6666) );
  XNOR U21280 ( .A(q[11]), .B(DB[1796]), .Z(n6664) );
  IV U21281 ( .A(n6663), .Z(n19515) );
  XNOR U21282 ( .A(n6661), .B(n19517), .Z(n6663) );
  XNOR U21283 ( .A(q[10]), .B(DB[1795]), .Z(n19517) );
  XNOR U21284 ( .A(q[9]), .B(DB[1794]), .Z(n6661) );
  IV U21285 ( .A(n6676), .Z(n19511) );
  XOR U21286 ( .A(n19518), .B(n19519), .Z(n6676) );
  XNOR U21287 ( .A(n6693), .B(n6674), .Z(n19519) );
  XNOR U21288 ( .A(q[0]), .B(DB[1785]), .Z(n6674) );
  XOR U21289 ( .A(n19520), .B(n6682), .Z(n6693) );
  XNOR U21290 ( .A(q[7]), .B(DB[1792]), .Z(n6682) );
  IV U21291 ( .A(n6681), .Z(n19520) );
  XNOR U21292 ( .A(n6679), .B(n19521), .Z(n6681) );
  XNOR U21293 ( .A(q[6]), .B(DB[1791]), .Z(n19521) );
  XNOR U21294 ( .A(q[5]), .B(DB[1790]), .Z(n6679) );
  IV U21295 ( .A(n6692), .Z(n19518) );
  XOR U21296 ( .A(n19522), .B(n19523), .Z(n6692) );
  XNOR U21297 ( .A(n6688), .B(n6690), .Z(n19523) );
  XNOR U21298 ( .A(q[1]), .B(DB[1786]), .Z(n6690) );
  XNOR U21299 ( .A(q[4]), .B(DB[1789]), .Z(n6688) );
  IV U21300 ( .A(n6687), .Z(n19522) );
  XNOR U21301 ( .A(n6685), .B(n19524), .Z(n6687) );
  XNOR U21302 ( .A(q[3]), .B(DB[1788]), .Z(n19524) );
  XNOR U21303 ( .A(q[2]), .B(DB[1787]), .Z(n6685) );
  XOR U21304 ( .A(n19525), .B(n6583), .Z(n6511) );
  XOR U21305 ( .A(n19526), .B(n6575), .Z(n6583) );
  XOR U21306 ( .A(n19527), .B(n6564), .Z(n6575) );
  XNOR U21307 ( .A(q[14]), .B(DB[1814]), .Z(n6564) );
  IV U21308 ( .A(n6563), .Z(n19527) );
  XNOR U21309 ( .A(n6561), .B(n19528), .Z(n6563) );
  XNOR U21310 ( .A(q[13]), .B(DB[1813]), .Z(n19528) );
  XNOR U21311 ( .A(q[12]), .B(DB[1812]), .Z(n6561) );
  IV U21312 ( .A(n6574), .Z(n19526) );
  XOR U21313 ( .A(n19529), .B(n19530), .Z(n6574) );
  XNOR U21314 ( .A(n6570), .B(n6572), .Z(n19530) );
  XNOR U21315 ( .A(q[8]), .B(DB[1808]), .Z(n6572) );
  XNOR U21316 ( .A(q[11]), .B(DB[1811]), .Z(n6570) );
  IV U21317 ( .A(n6569), .Z(n19529) );
  XNOR U21318 ( .A(n6567), .B(n19531), .Z(n6569) );
  XNOR U21319 ( .A(q[10]), .B(DB[1810]), .Z(n19531) );
  XNOR U21320 ( .A(q[9]), .B(DB[1809]), .Z(n6567) );
  IV U21321 ( .A(n6582), .Z(n19525) );
  XOR U21322 ( .A(n19532), .B(n19533), .Z(n6582) );
  XNOR U21323 ( .A(n6599), .B(n6580), .Z(n19533) );
  XNOR U21324 ( .A(q[0]), .B(DB[1800]), .Z(n6580) );
  XOR U21325 ( .A(n19534), .B(n6588), .Z(n6599) );
  XNOR U21326 ( .A(q[7]), .B(DB[1807]), .Z(n6588) );
  IV U21327 ( .A(n6587), .Z(n19534) );
  XNOR U21328 ( .A(n6585), .B(n19535), .Z(n6587) );
  XNOR U21329 ( .A(q[6]), .B(DB[1806]), .Z(n19535) );
  XNOR U21330 ( .A(q[5]), .B(DB[1805]), .Z(n6585) );
  IV U21331 ( .A(n6598), .Z(n19532) );
  XOR U21332 ( .A(n19536), .B(n19537), .Z(n6598) );
  XNOR U21333 ( .A(n6594), .B(n6596), .Z(n19537) );
  XNOR U21334 ( .A(q[1]), .B(DB[1801]), .Z(n6596) );
  XNOR U21335 ( .A(q[4]), .B(DB[1804]), .Z(n6594) );
  IV U21336 ( .A(n6593), .Z(n19536) );
  XNOR U21337 ( .A(n6591), .B(n19538), .Z(n6593) );
  XNOR U21338 ( .A(q[3]), .B(DB[1803]), .Z(n19538) );
  XNOR U21339 ( .A(q[2]), .B(DB[1802]), .Z(n6591) );
  XOR U21340 ( .A(n19539), .B(n6489), .Z(n6417) );
  XOR U21341 ( .A(n19540), .B(n6481), .Z(n6489) );
  XOR U21342 ( .A(n19541), .B(n6470), .Z(n6481) );
  XNOR U21343 ( .A(q[14]), .B(DB[1829]), .Z(n6470) );
  IV U21344 ( .A(n6469), .Z(n19541) );
  XNOR U21345 ( .A(n6467), .B(n19542), .Z(n6469) );
  XNOR U21346 ( .A(q[13]), .B(DB[1828]), .Z(n19542) );
  XNOR U21347 ( .A(q[12]), .B(DB[1827]), .Z(n6467) );
  IV U21348 ( .A(n6480), .Z(n19540) );
  XOR U21349 ( .A(n19543), .B(n19544), .Z(n6480) );
  XNOR U21350 ( .A(n6476), .B(n6478), .Z(n19544) );
  XNOR U21351 ( .A(q[8]), .B(DB[1823]), .Z(n6478) );
  XNOR U21352 ( .A(q[11]), .B(DB[1826]), .Z(n6476) );
  IV U21353 ( .A(n6475), .Z(n19543) );
  XNOR U21354 ( .A(n6473), .B(n19545), .Z(n6475) );
  XNOR U21355 ( .A(q[10]), .B(DB[1825]), .Z(n19545) );
  XNOR U21356 ( .A(q[9]), .B(DB[1824]), .Z(n6473) );
  IV U21357 ( .A(n6488), .Z(n19539) );
  XOR U21358 ( .A(n19546), .B(n19547), .Z(n6488) );
  XNOR U21359 ( .A(n6505), .B(n6486), .Z(n19547) );
  XNOR U21360 ( .A(q[0]), .B(DB[1815]), .Z(n6486) );
  XOR U21361 ( .A(n19548), .B(n6494), .Z(n6505) );
  XNOR U21362 ( .A(q[7]), .B(DB[1822]), .Z(n6494) );
  IV U21363 ( .A(n6493), .Z(n19548) );
  XNOR U21364 ( .A(n6491), .B(n19549), .Z(n6493) );
  XNOR U21365 ( .A(q[6]), .B(DB[1821]), .Z(n19549) );
  XNOR U21366 ( .A(q[5]), .B(DB[1820]), .Z(n6491) );
  IV U21367 ( .A(n6504), .Z(n19546) );
  XOR U21368 ( .A(n19550), .B(n19551), .Z(n6504) );
  XNOR U21369 ( .A(n6500), .B(n6502), .Z(n19551) );
  XNOR U21370 ( .A(q[1]), .B(DB[1816]), .Z(n6502) );
  XNOR U21371 ( .A(q[4]), .B(DB[1819]), .Z(n6500) );
  IV U21372 ( .A(n6499), .Z(n19550) );
  XNOR U21373 ( .A(n6497), .B(n19552), .Z(n6499) );
  XNOR U21374 ( .A(q[3]), .B(DB[1818]), .Z(n19552) );
  XNOR U21375 ( .A(q[2]), .B(DB[1817]), .Z(n6497) );
  XOR U21376 ( .A(n19553), .B(n6395), .Z(n6323) );
  XOR U21377 ( .A(n19554), .B(n6387), .Z(n6395) );
  XOR U21378 ( .A(n19555), .B(n6376), .Z(n6387) );
  XNOR U21379 ( .A(q[14]), .B(DB[1844]), .Z(n6376) );
  IV U21380 ( .A(n6375), .Z(n19555) );
  XNOR U21381 ( .A(n6373), .B(n19556), .Z(n6375) );
  XNOR U21382 ( .A(q[13]), .B(DB[1843]), .Z(n19556) );
  XNOR U21383 ( .A(q[12]), .B(DB[1842]), .Z(n6373) );
  IV U21384 ( .A(n6386), .Z(n19554) );
  XOR U21385 ( .A(n19557), .B(n19558), .Z(n6386) );
  XNOR U21386 ( .A(n6382), .B(n6384), .Z(n19558) );
  XNOR U21387 ( .A(q[8]), .B(DB[1838]), .Z(n6384) );
  XNOR U21388 ( .A(q[11]), .B(DB[1841]), .Z(n6382) );
  IV U21389 ( .A(n6381), .Z(n19557) );
  XNOR U21390 ( .A(n6379), .B(n19559), .Z(n6381) );
  XNOR U21391 ( .A(q[10]), .B(DB[1840]), .Z(n19559) );
  XNOR U21392 ( .A(q[9]), .B(DB[1839]), .Z(n6379) );
  IV U21393 ( .A(n6394), .Z(n19553) );
  XOR U21394 ( .A(n19560), .B(n19561), .Z(n6394) );
  XNOR U21395 ( .A(n6411), .B(n6392), .Z(n19561) );
  XNOR U21396 ( .A(q[0]), .B(DB[1830]), .Z(n6392) );
  XOR U21397 ( .A(n19562), .B(n6400), .Z(n6411) );
  XNOR U21398 ( .A(q[7]), .B(DB[1837]), .Z(n6400) );
  IV U21399 ( .A(n6399), .Z(n19562) );
  XNOR U21400 ( .A(n6397), .B(n19563), .Z(n6399) );
  XNOR U21401 ( .A(q[6]), .B(DB[1836]), .Z(n19563) );
  XNOR U21402 ( .A(q[5]), .B(DB[1835]), .Z(n6397) );
  IV U21403 ( .A(n6410), .Z(n19560) );
  XOR U21404 ( .A(n19564), .B(n19565), .Z(n6410) );
  XNOR U21405 ( .A(n6406), .B(n6408), .Z(n19565) );
  XNOR U21406 ( .A(q[1]), .B(DB[1831]), .Z(n6408) );
  XNOR U21407 ( .A(q[4]), .B(DB[1834]), .Z(n6406) );
  IV U21408 ( .A(n6405), .Z(n19564) );
  XNOR U21409 ( .A(n6403), .B(n19566), .Z(n6405) );
  XNOR U21410 ( .A(q[3]), .B(DB[1833]), .Z(n19566) );
  XNOR U21411 ( .A(q[2]), .B(DB[1832]), .Z(n6403) );
  XOR U21412 ( .A(n19567), .B(n6301), .Z(n6229) );
  XOR U21413 ( .A(n19568), .B(n6293), .Z(n6301) );
  XOR U21414 ( .A(n19569), .B(n6282), .Z(n6293) );
  XNOR U21415 ( .A(q[14]), .B(DB[1859]), .Z(n6282) );
  IV U21416 ( .A(n6281), .Z(n19569) );
  XNOR U21417 ( .A(n6279), .B(n19570), .Z(n6281) );
  XNOR U21418 ( .A(q[13]), .B(DB[1858]), .Z(n19570) );
  XNOR U21419 ( .A(q[12]), .B(DB[1857]), .Z(n6279) );
  IV U21420 ( .A(n6292), .Z(n19568) );
  XOR U21421 ( .A(n19571), .B(n19572), .Z(n6292) );
  XNOR U21422 ( .A(n6288), .B(n6290), .Z(n19572) );
  XNOR U21423 ( .A(q[8]), .B(DB[1853]), .Z(n6290) );
  XNOR U21424 ( .A(q[11]), .B(DB[1856]), .Z(n6288) );
  IV U21425 ( .A(n6287), .Z(n19571) );
  XNOR U21426 ( .A(n6285), .B(n19573), .Z(n6287) );
  XNOR U21427 ( .A(q[10]), .B(DB[1855]), .Z(n19573) );
  XNOR U21428 ( .A(q[9]), .B(DB[1854]), .Z(n6285) );
  IV U21429 ( .A(n6300), .Z(n19567) );
  XOR U21430 ( .A(n19574), .B(n19575), .Z(n6300) );
  XNOR U21431 ( .A(n6317), .B(n6298), .Z(n19575) );
  XNOR U21432 ( .A(q[0]), .B(DB[1845]), .Z(n6298) );
  XOR U21433 ( .A(n19576), .B(n6306), .Z(n6317) );
  XNOR U21434 ( .A(q[7]), .B(DB[1852]), .Z(n6306) );
  IV U21435 ( .A(n6305), .Z(n19576) );
  XNOR U21436 ( .A(n6303), .B(n19577), .Z(n6305) );
  XNOR U21437 ( .A(q[6]), .B(DB[1851]), .Z(n19577) );
  XNOR U21438 ( .A(q[5]), .B(DB[1850]), .Z(n6303) );
  IV U21439 ( .A(n6316), .Z(n19574) );
  XOR U21440 ( .A(n19578), .B(n19579), .Z(n6316) );
  XNOR U21441 ( .A(n6312), .B(n6314), .Z(n19579) );
  XNOR U21442 ( .A(q[1]), .B(DB[1846]), .Z(n6314) );
  XNOR U21443 ( .A(q[4]), .B(DB[1849]), .Z(n6312) );
  IV U21444 ( .A(n6311), .Z(n19578) );
  XNOR U21445 ( .A(n6309), .B(n19580), .Z(n6311) );
  XNOR U21446 ( .A(q[3]), .B(DB[1848]), .Z(n19580) );
  XNOR U21447 ( .A(q[2]), .B(DB[1847]), .Z(n6309) );
  XOR U21448 ( .A(n19581), .B(n6207), .Z(n6135) );
  XOR U21449 ( .A(n19582), .B(n6199), .Z(n6207) );
  XOR U21450 ( .A(n19583), .B(n6188), .Z(n6199) );
  XNOR U21451 ( .A(q[14]), .B(DB[1874]), .Z(n6188) );
  IV U21452 ( .A(n6187), .Z(n19583) );
  XNOR U21453 ( .A(n6185), .B(n19584), .Z(n6187) );
  XNOR U21454 ( .A(q[13]), .B(DB[1873]), .Z(n19584) );
  XNOR U21455 ( .A(q[12]), .B(DB[1872]), .Z(n6185) );
  IV U21456 ( .A(n6198), .Z(n19582) );
  XOR U21457 ( .A(n19585), .B(n19586), .Z(n6198) );
  XNOR U21458 ( .A(n6194), .B(n6196), .Z(n19586) );
  XNOR U21459 ( .A(q[8]), .B(DB[1868]), .Z(n6196) );
  XNOR U21460 ( .A(q[11]), .B(DB[1871]), .Z(n6194) );
  IV U21461 ( .A(n6193), .Z(n19585) );
  XNOR U21462 ( .A(n6191), .B(n19587), .Z(n6193) );
  XNOR U21463 ( .A(q[10]), .B(DB[1870]), .Z(n19587) );
  XNOR U21464 ( .A(q[9]), .B(DB[1869]), .Z(n6191) );
  IV U21465 ( .A(n6206), .Z(n19581) );
  XOR U21466 ( .A(n19588), .B(n19589), .Z(n6206) );
  XNOR U21467 ( .A(n6223), .B(n6204), .Z(n19589) );
  XNOR U21468 ( .A(q[0]), .B(DB[1860]), .Z(n6204) );
  XOR U21469 ( .A(n19590), .B(n6212), .Z(n6223) );
  XNOR U21470 ( .A(q[7]), .B(DB[1867]), .Z(n6212) );
  IV U21471 ( .A(n6211), .Z(n19590) );
  XNOR U21472 ( .A(n6209), .B(n19591), .Z(n6211) );
  XNOR U21473 ( .A(q[6]), .B(DB[1866]), .Z(n19591) );
  XNOR U21474 ( .A(q[5]), .B(DB[1865]), .Z(n6209) );
  IV U21475 ( .A(n6222), .Z(n19588) );
  XOR U21476 ( .A(n19592), .B(n19593), .Z(n6222) );
  XNOR U21477 ( .A(n6218), .B(n6220), .Z(n19593) );
  XNOR U21478 ( .A(q[1]), .B(DB[1861]), .Z(n6220) );
  XNOR U21479 ( .A(q[4]), .B(DB[1864]), .Z(n6218) );
  IV U21480 ( .A(n6217), .Z(n19592) );
  XNOR U21481 ( .A(n6215), .B(n19594), .Z(n6217) );
  XNOR U21482 ( .A(q[3]), .B(DB[1863]), .Z(n19594) );
  XNOR U21483 ( .A(q[2]), .B(DB[1862]), .Z(n6215) );
  XOR U21484 ( .A(n19595), .B(n6113), .Z(n6041) );
  XOR U21485 ( .A(n19596), .B(n6105), .Z(n6113) );
  XOR U21486 ( .A(n19597), .B(n6094), .Z(n6105) );
  XNOR U21487 ( .A(q[14]), .B(DB[1889]), .Z(n6094) );
  IV U21488 ( .A(n6093), .Z(n19597) );
  XNOR U21489 ( .A(n6091), .B(n19598), .Z(n6093) );
  XNOR U21490 ( .A(q[13]), .B(DB[1888]), .Z(n19598) );
  XNOR U21491 ( .A(q[12]), .B(DB[1887]), .Z(n6091) );
  IV U21492 ( .A(n6104), .Z(n19596) );
  XOR U21493 ( .A(n19599), .B(n19600), .Z(n6104) );
  XNOR U21494 ( .A(n6100), .B(n6102), .Z(n19600) );
  XNOR U21495 ( .A(q[8]), .B(DB[1883]), .Z(n6102) );
  XNOR U21496 ( .A(q[11]), .B(DB[1886]), .Z(n6100) );
  IV U21497 ( .A(n6099), .Z(n19599) );
  XNOR U21498 ( .A(n6097), .B(n19601), .Z(n6099) );
  XNOR U21499 ( .A(q[10]), .B(DB[1885]), .Z(n19601) );
  XNOR U21500 ( .A(q[9]), .B(DB[1884]), .Z(n6097) );
  IV U21501 ( .A(n6112), .Z(n19595) );
  XOR U21502 ( .A(n19602), .B(n19603), .Z(n6112) );
  XNOR U21503 ( .A(n6129), .B(n6110), .Z(n19603) );
  XNOR U21504 ( .A(q[0]), .B(DB[1875]), .Z(n6110) );
  XOR U21505 ( .A(n19604), .B(n6118), .Z(n6129) );
  XNOR U21506 ( .A(q[7]), .B(DB[1882]), .Z(n6118) );
  IV U21507 ( .A(n6117), .Z(n19604) );
  XNOR U21508 ( .A(n6115), .B(n19605), .Z(n6117) );
  XNOR U21509 ( .A(q[6]), .B(DB[1881]), .Z(n19605) );
  XNOR U21510 ( .A(q[5]), .B(DB[1880]), .Z(n6115) );
  IV U21511 ( .A(n6128), .Z(n19602) );
  XOR U21512 ( .A(n19606), .B(n19607), .Z(n6128) );
  XNOR U21513 ( .A(n6124), .B(n6126), .Z(n19607) );
  XNOR U21514 ( .A(q[1]), .B(DB[1876]), .Z(n6126) );
  XNOR U21515 ( .A(q[4]), .B(DB[1879]), .Z(n6124) );
  IV U21516 ( .A(n6123), .Z(n19606) );
  XNOR U21517 ( .A(n6121), .B(n19608), .Z(n6123) );
  XNOR U21518 ( .A(q[3]), .B(DB[1878]), .Z(n19608) );
  XNOR U21519 ( .A(q[2]), .B(DB[1877]), .Z(n6121) );
  XOR U21520 ( .A(n19609), .B(n6019), .Z(n5945) );
  XOR U21521 ( .A(n19610), .B(n6011), .Z(n6019) );
  XOR U21522 ( .A(n19611), .B(n6000), .Z(n6011) );
  XNOR U21523 ( .A(q[14]), .B(DB[1904]), .Z(n6000) );
  IV U21524 ( .A(n5999), .Z(n19611) );
  XNOR U21525 ( .A(n5997), .B(n19612), .Z(n5999) );
  XNOR U21526 ( .A(q[13]), .B(DB[1903]), .Z(n19612) );
  XOR U21527 ( .A(q[12]), .B(n4313), .Z(n5997) );
  IV U21528 ( .A(DB[1902]), .Z(n4313) );
  IV U21529 ( .A(n6010), .Z(n19610) );
  XOR U21530 ( .A(n19613), .B(n19614), .Z(n6010) );
  XNOR U21531 ( .A(n6006), .B(n6008), .Z(n19614) );
  XNOR U21532 ( .A(q[8]), .B(DB[1898]), .Z(n6008) );
  XOR U21533 ( .A(q[11]), .B(n4695), .Z(n6006) );
  IV U21534 ( .A(DB[1901]), .Z(n4695) );
  IV U21535 ( .A(n6005), .Z(n19613) );
  XNOR U21536 ( .A(n6003), .B(n19615), .Z(n6005) );
  XNOR U21537 ( .A(q[10]), .B(DB[1900]), .Z(n19615) );
  XNOR U21538 ( .A(q[9]), .B(DB[1899]), .Z(n6003) );
  IV U21539 ( .A(n6018), .Z(n19609) );
  XOR U21540 ( .A(n19616), .B(n19617), .Z(n6018) );
  XNOR U21541 ( .A(n6035), .B(n6016), .Z(n19617) );
  XNOR U21542 ( .A(q[0]), .B(DB[1890]), .Z(n6016) );
  XOR U21543 ( .A(n19618), .B(n6024), .Z(n6035) );
  XNOR U21544 ( .A(q[7]), .B(DB[1897]), .Z(n6024) );
  IV U21545 ( .A(n6023), .Z(n19618) );
  XNOR U21546 ( .A(n6021), .B(n19619), .Z(n6023) );
  XNOR U21547 ( .A(q[6]), .B(DB[1896]), .Z(n19619) );
  XNOR U21548 ( .A(q[5]), .B(DB[1895]), .Z(n6021) );
  IV U21549 ( .A(n6034), .Z(n19616) );
  XOR U21550 ( .A(n19620), .B(n19621), .Z(n6034) );
  XNOR U21551 ( .A(n6030), .B(n6032), .Z(n19621) );
  XNOR U21552 ( .A(q[1]), .B(DB[1891]), .Z(n6032) );
  XNOR U21553 ( .A(q[4]), .B(DB[1894]), .Z(n6030) );
  IV U21554 ( .A(n6029), .Z(n19620) );
  XNOR U21555 ( .A(n6027), .B(n19622), .Z(n6029) );
  XNOR U21556 ( .A(q[3]), .B(DB[1893]), .Z(n19622) );
  XNOR U21557 ( .A(q[2]), .B(DB[1892]), .Z(n6027) );
endmodule

