

    module a23_gc_main_CODE_MEM_SIZE32_G_MEM_SIZE8_E_MEM_SIZE8_OUT_MEM_SIZE8_STACK_MEM_SIZE8 ( 
        clk, rst, p_init, g_init, e_init, o, terminate );
  input [1023:0] p_init;
  input [255:0] g_init;
  input [255:0] e_init;
  output [255:0] o;
  input clk, rst;
  output terminate;
  wire   m_write_en, \u_a23_core/status_bits_flags_wen ,
         \u_a23_core/reg_bank_wen[14] , \u_a23_core/reg_bank_wen[13] ,
         \u_a23_core/reg_bank_wen[12] , \u_a23_core/reg_bank_wen[11] ,
         \u_a23_core/reg_bank_wen[10] , \u_a23_core/reg_bank_wen[9] ,
         \u_a23_core/reg_bank_wen[8] , \u_a23_core/reg_bank_wen[7] ,
         \u_a23_core/reg_bank_wen[6] , \u_a23_core/reg_bank_wen[5] ,
         \u_a23_core/reg_bank_wen[4] , \u_a23_core/reg_bank_wen[3] ,
         \u_a23_core/reg_bank_wen[2] , \u_a23_core/reg_bank_wen[1] ,
         \u_a23_core/reg_bank_wen[0] , \u_a23_core/pc_wen ,
         \u_a23_core/write_data_wen , \u_a23_core/reg_write_sel[1] ,
         \u_a23_core/reg_write_sel[0] , \u_a23_core/status_bits_sel[2] ,
         \u_a23_core/status_bits_sel[0] , \u_a23_core/byte_enable_sel[0] ,
         \u_a23_core/pc_sel[1] , \u_a23_core/pc_sel[0] ,
         \u_a23_core/address_sel[3] , \u_a23_core/address_sel[2] ,
         \u_a23_core/address_sel[1] , \u_a23_core/address_sel[0] ,
         \u_a23_core/multiply_function[1] , \u_a23_core/multiply_function[0] ,
         \u_a23_core/alu_function[8] , \u_a23_core/alu_function[7] ,
         \u_a23_core/alu_function[6] , \u_a23_core/alu_function[5] ,
         \u_a23_core/alu_function[4] , \u_a23_core/alu_function[3] ,
         \u_a23_core/alu_function[2] , \u_a23_core/alu_function[1] ,
         \u_a23_core/alu_function[0] , \u_a23_core/use_carry_in ,
         \u_a23_core/barrel_shift_function[1] ,
         \u_a23_core/barrel_shift_function[0] ,
         \u_a23_core/barrel_shift_data_sel[1] ,
         \u_a23_core/barrel_shift_data_sel[0] ,
         \u_a23_core/barrel_shift_amount_sel[1] ,
         \u_a23_core/barrel_shift_amount_sel[0] , \u_a23_core/rn_sel_nxt[3] ,
         \u_a23_core/rn_sel_nxt[2] , \u_a23_core/rn_sel_nxt[1] ,
         \u_a23_core/rn_sel_nxt[0] , \u_a23_core/rds_sel_nxt[3] ,
         \u_a23_core/rds_sel_nxt[2] , \u_a23_core/rds_sel_nxt[1] ,
         \u_a23_core/rds_sel_nxt[0] , \u_a23_core/rm_sel_nxt[3] ,
         \u_a23_core/rm_sel_nxt[2] , \u_a23_core/rm_sel_nxt[1] ,
         \u_a23_core/rm_sel_nxt[0] , \u_a23_core/rn_sel[3] ,
         \u_a23_core/rn_sel[2] , \u_a23_core/rn_sel[1] ,
         \u_a23_core/rn_sel[0] , \u_a23_core/rds_sel[3] ,
         \u_a23_core/rds_sel[2] , \u_a23_core/rds_sel[1] ,
         \u_a23_core/rds_sel[0] , \u_a23_core/rm_sel[3] ,
         \u_a23_core/rm_sel[2] , \u_a23_core/rm_sel[1] ,
         \u_a23_core/rm_sel[0] , \u_a23_core/condition[3] ,
         \u_a23_core/condition[2] , \u_a23_core/condition[1] ,
         \u_a23_core/condition[0] , \u_a23_core/shift_imm_zero ,
         \u_a23_core/imm_shift_amount[4] , \u_a23_core/imm_shift_amount[3] ,
         \u_a23_core/imm_shift_amount[2] , \u_a23_core/imm_shift_amount[1] ,
         \u_a23_core/imm_shift_amount[0] , \u_a23_core/imm32[31] ,
         \u_a23_core/imm32[30] , \u_a23_core/imm32[29] ,
         \u_a23_core/imm32[28] , \u_a23_core/imm32[27] ,
         \u_a23_core/imm32[26] , \u_a23_core/imm32[25] ,
         \u_a23_core/imm32[24] , \u_a23_core/imm32[23] ,
         \u_a23_core/imm32[22] , \u_a23_core/imm32[21] ,
         \u_a23_core/imm32[20] , \u_a23_core/imm32[19] ,
         \u_a23_core/imm32[18] , \u_a23_core/imm32[17] ,
         \u_a23_core/imm32[16] , \u_a23_core/imm32[15] ,
         \u_a23_core/imm32[14] , \u_a23_core/imm32[13] ,
         \u_a23_core/imm32[12] , \u_a23_core/imm32[11] ,
         \u_a23_core/imm32[10] , \u_a23_core/imm32[9] , \u_a23_core/imm32[8] ,
         \u_a23_core/imm32[7] , \u_a23_core/imm32[6] , \u_a23_core/imm32[5] ,
         \u_a23_core/imm32[4] , \u_a23_core/imm32[3] , \u_a23_core/imm32[2] ,
         \u_a23_core/imm32[1] , \u_a23_core/imm32[0] ,
         \u_a23_core/multiply_done , \u_a23_core/read_data_alignment[4] ,
         \u_a23_core/read_data_alignment[3] , \u_a23_core/read_data_s2[31] ,
         \u_a23_core/read_data_s2[30] , \u_a23_core/read_data_s2[29] ,
         \u_a23_core/read_data_s2[28] , \u_a23_core/read_data_s2[27] ,
         \u_a23_core/read_data_s2[26] , \u_a23_core/read_data_s2[25] ,
         \u_a23_core/read_data_s2[24] , \u_a23_core/read_data_s2[23] ,
         \u_a23_core/read_data_s2[22] , \u_a23_core/read_data_s2[21] ,
         \u_a23_core/read_data_s2[20] , \u_a23_core/read_data_s2[19] ,
         \u_a23_core/read_data_s2[18] , \u_a23_core/read_data_s2[17] ,
         \u_a23_core/read_data_s2[16] , \u_a23_core/read_data_s2[15] ,
         \u_a23_core/read_data_s2[14] , \u_a23_core/read_data_s2[13] ,
         \u_a23_core/read_data_s2[12] , \u_a23_core/read_data_s2[11] ,
         \u_a23_core/read_data_s2[10] , \u_a23_core/read_data_s2[9] ,
         \u_a23_core/read_data_s2[8] , \u_a23_core/read_data_s2[7] ,
         \u_a23_core/read_data_s2[6] , \u_a23_core/read_data_s2[5] ,
         \u_a23_core/read_data_s2[4] , \u_a23_core/read_data_s2[3] ,
         \u_a23_core/read_data_s2[2] , \u_a23_core/read_data_s2[1] ,
         \u_a23_core/read_data_s2[0] , \u_a23_core/read_data[31] ,
         \u_a23_core/read_data[30] , \u_a23_core/read_data[29] ,
         \u_a23_core/read_data[28] , \u_a23_core/read_data[27] ,
         \u_a23_core/read_data[26] , \u_a23_core/read_data[25] ,
         \u_a23_core/read_data[24] , \u_a23_core/read_data[23] ,
         \u_a23_core/read_data[22] , \u_a23_core/read_data[21] ,
         \u_a23_core/read_data[20] , \u_a23_core/read_data[19] ,
         \u_a23_core/read_data[18] , \u_a23_core/read_data[17] ,
         \u_a23_core/read_data[16] , \u_a23_core/read_data[15] ,
         \u_a23_core/read_data[14] , \u_a23_core/read_data[13] ,
         \u_a23_core/read_data[12] , \u_a23_core/read_data[11] ,
         \u_a23_core/read_data[10] , \u_a23_core/read_data[9] ,
         \u_a23_core/read_data[8] , \u_a23_core/read_data[7] ,
         \u_a23_core/read_data[6] , \u_a23_core/read_data[5] ,
         \u_a23_core/read_data[4] , \u_a23_core/read_data[3] ,
         \u_a23_core/read_data[2] , \u_a23_core/read_data[1] ,
         \u_a23_core/read_data[0] , \u_a23_core/execute_address_nxt[0] ,
         \u_a23_core/execute_address_nxt[1] ,
         \u_a23_core/execute_address_nxt[2] ,
         \u_a23_core/execute_address_nxt[3] ,
         \u_a23_core/execute_address_nxt[4] ,
         \u_a23_core/execute_address_nxt[5] ,
         \u_a23_core/execute_address_nxt[6] ,
         \u_a23_core/execute_address_nxt[7] ,
         \u_a23_core/execute_address_nxt[8] ,
         \u_a23_core/execute_address_nxt[9] ,
         \u_a23_core/execute_address_nxt[10] ,
         \u_a23_core/execute_address_nxt[11] ,
         \u_a23_core/execute_address_nxt[12] ,
         \u_a23_core/execute_address_nxt[13] ,
         \u_a23_core/execute_address_nxt[14] ,
         \u_a23_core/execute_address_nxt[15] ,
         \u_a23_core/execute_address_nxt[16] ,
         \u_a23_core/execute_address_nxt[17] ,
         \u_a23_core/execute_address_nxt[18] ,
         \u_a23_core/execute_address_nxt[19] ,
         \u_a23_core/execute_address_nxt[20] ,
         \u_a23_core/execute_address_nxt[21] ,
         \u_a23_core/execute_address_nxt[22] ,
         \u_a23_core/execute_address_nxt[23] ,
         \u_a23_core/execute_address_nxt[24] ,
         \u_a23_core/execute_address_nxt[25] ,
         \u_a23_core/execute_address_nxt[26] ,
         \u_a23_core/execute_address_nxt[27] ,
         \u_a23_core/execute_address_nxt[28] ,
         \u_a23_core/execute_address_nxt[29] ,
         \u_a23_core/execute_address_nxt[30] ,
         \u_a23_core/execute_address_nxt[31] , \u_a23_core/execute_address[1] ,
         \u_a23_mem/n23820 , \u_a23_mem/n23819 , \u_a23_mem/n23812 ,
         \u_a23_mem/n23805 , \u_a23_mem/n23804 , \u_a23_mem/n23797 ,
         \u_a23_mem/n23790 , \u_a23_mem/n23789 , \u_a23_mem/n23782 ,
         \u_a23_mem/n23775 , \u_a23_mem/n23774 , \u_a23_mem/n23767 ,
         \u_a23_mem/n23760 , \u_a23_mem/n23759 , \u_a23_mem/n23752 ,
         \u_a23_mem/n23745 , \u_a23_mem/n23744 , \u_a23_mem/n23737 ,
         \u_a23_mem/n23730 , \u_a23_mem/n23729 , \u_a23_mem/n23722 ,
         \u_a23_mem/n23715 , \u_a23_mem/n23714 , \u_a23_mem/n23707 ,
         \u_a23_mem/n23700 , \u_a23_mem/n23699 , \u_a23_mem/n23692 ,
         \u_a23_mem/n23685 , \u_a23_mem/n23684 , \u_a23_mem/n23677 ,
         \u_a23_mem/n23670 , \u_a23_mem/n23669 , \u_a23_mem/n23662 ,
         \u_a23_mem/n23655 , \u_a23_mem/n23654 , \u_a23_mem/n23647 ,
         \u_a23_mem/n23640 , \u_a23_mem/n23639 , \u_a23_mem/n23632 ,
         \u_a23_mem/n23625 , \u_a23_mem/n23624 , \u_a23_mem/n23617 ,
         \u_a23_mem/n23610 , \u_a23_mem/n23609 , \u_a23_mem/n23602 ,
         \u_a23_mem/n23595 , \u_a23_mem/n23594 , \u_a23_mem/n23587 ,
         \u_a23_mem/n23580 , \u_a23_mem/n23579 , \u_a23_mem/n23572 ,
         \u_a23_mem/n23565 , \u_a23_mem/n23564 , \u_a23_mem/n23557 ,
         \u_a23_mem/n23550 , \u_a23_mem/n23549 , \u_a23_mem/n23542 ,
         \u_a23_mem/n23535 , \u_a23_mem/n23534 , \u_a23_mem/n23527 ,
         \u_a23_mem/n23520 , \u_a23_mem/n23519 , \u_a23_mem/n23512 ,
         \u_a23_mem/n23505 , \u_a23_mem/n23504 , \u_a23_mem/n23497 ,
         \u_a23_mem/n23490 , \u_a23_mem/n23489 , \u_a23_mem/n23482 ,
         \u_a23_mem/n23475 , \u_a23_mem/n23474 , \u_a23_mem/n23467 ,
         \u_a23_mem/n23460 , \u_a23_mem/n23459 , \u_a23_mem/n23452 ,
         \u_a23_mem/n23445 , \u_a23_mem/n23444 , \u_a23_mem/n23437 ,
         \u_a23_mem/n23430 , \u_a23_mem/n23429 , \u_a23_mem/n23422 ,
         \u_a23_mem/n23415 , \u_a23_mem/n23414 , \u_a23_mem/n23407 ,
         \u_a23_mem/n23400 , \u_a23_mem/n23399 , \u_a23_mem/n23392 ,
         \u_a23_mem/n23385 , \u_a23_mem/n23384 , \u_a23_mem/n23377 ,
         \u_a23_mem/n23370 , \u_a23_mem/n23369 , \u_a23_mem/n23362 ,
         \u_a23_mem/n23355 , \u_a23_mem/n23354 , \u_a23_mem/n23347 ,
         \u_a23_mem/n23340 , \u_a23_mem/n23339 , \u_a23_mem/n23332 ,
         \u_a23_mem/n23325 , \u_a23_mem/n23324 , \u_a23_mem/n23317 ,
         \u_a23_mem/n23310 , \u_a23_mem/n23309 , \u_a23_mem/n23302 ,
         \u_a23_mem/n23295 , \u_a23_mem/n23294 , \u_a23_mem/n23287 ,
         \u_a23_mem/n23280 , \u_a23_mem/n23279 , \u_a23_mem/n23272 ,
         \u_a23_mem/n23265 , \u_a23_mem/n23264 , \u_a23_mem/n23257 ,
         \u_a23_mem/n23250 , \u_a23_mem/n23249 , \u_a23_mem/n23242 ,
         \u_a23_mem/n23235 , \u_a23_mem/n23234 , \u_a23_mem/n23227 ,
         \u_a23_mem/n23220 , \u_a23_mem/n23219 , \u_a23_mem/n23212 ,
         \u_a23_mem/n23205 , \u_a23_mem/n23204 , \u_a23_mem/n23197 ,
         \u_a23_mem/n23190 , \u_a23_mem/n23189 , \u_a23_mem/n23182 ,
         \u_a23_mem/n23175 , \u_a23_mem/n23174 , \u_a23_mem/n23167 ,
         \u_a23_mem/n23160 , \u_a23_mem/n23159 , \u_a23_mem/n23152 ,
         \u_a23_mem/n23145 , \u_a23_mem/n23144 , \u_a23_mem/n23137 ,
         \u_a23_mem/n23130 , \u_a23_mem/n23129 , \u_a23_mem/n23122 ,
         \u_a23_mem/n23115 , \u_a23_mem/n23114 , \u_a23_mem/n23107 ,
         \u_a23_mem/n23100 , \u_a23_mem/n23099 , \u_a23_mem/n23092 ,
         \u_a23_mem/n23085 , \u_a23_mem/n23084 , \u_a23_mem/n23077 ,
         \u_a23_mem/n23070 , \u_a23_mem/n23069 , \u_a23_mem/n23062 ,
         \u_a23_mem/n23055 , \u_a23_mem/n23054 , \u_a23_mem/n23047 ,
         \u_a23_mem/n23040 , \u_a23_mem/n23039 , \u_a23_mem/n23032 ,
         \u_a23_mem/n23025 , \u_a23_mem/n23024 , \u_a23_mem/n23017 ,
         \u_a23_mem/n23010 , \u_a23_mem/n23009 , \u_a23_mem/n23002 ,
         \u_a23_mem/n22995 , \u_a23_mem/n22994 , \u_a23_mem/n22987 ,
         \u_a23_mem/n22980 , \u_a23_mem/n22979 , \u_a23_mem/n22972 ,
         \u_a23_mem/n22965 , \u_a23_mem/n22964 , \u_a23_mem/n22957 ,
         \u_a23_mem/n22950 , \u_a23_mem/n22949 , \u_a23_mem/n22942 ,
         \u_a23_mem/n22935 , \u_a23_mem/n22934 , \u_a23_mem/n22927 ,
         \u_a23_mem/n22920 , \u_a23_mem/n22919 , \u_a23_mem/n22912 ,
         \u_a23_mem/n22905 , \u_a23_mem/n22904 , \u_a23_mem/n22897 ,
         \u_a23_mem/n22890 , \u_a23_mem/n22889 , \u_a23_mem/n22882 ,
         \u_a23_mem/n22875 , \u_a23_mem/n22874 , \u_a23_mem/n22867 ,
         \u_a23_mem/n22860 , \u_a23_mem/n22859 , \u_a23_mem/n22858 ,
         \u_a23_mem/n22857 , \u_a23_mem/n22850 , \u_a23_mem/n22843 ,
         \u_a23_mem/n22842 , \u_a23_mem/n22835 , \u_a23_mem/n22828 ,
         \u_a23_mem/n22827 , \u_a23_mem/n22826 , \u_a23_mem/n22819 ,
         \u_a23_mem/n22812 , \u_a23_mem/n22811 , \u_a23_mem/n22804 ,
         \u_a23_mem/n22797 , \u_a23_mem/n22796 , \u_a23_mem/n22795 ,
         \u_a23_mem/n22794 , \u_a23_mem/n22787 , \u_a23_mem/n22780 ,
         \u_a23_mem/n22779 , \u_a23_mem/n22772 , \u_a23_mem/n22765 ,
         \u_a23_mem/n22764 , \u_a23_mem/n22763 , \u_a23_mem/n22756 ,
         \u_a23_mem/n22749 , \u_a23_mem/n22748 , \u_a23_mem/n22741 ,
         \u_a23_mem/n22734 , \u_a23_mem/n22733 , \u_a23_mem/n22732 ,
         \u_a23_mem/n22731 , \u_a23_mem/n22724 , \u_a23_mem/n22717 ,
         \u_a23_mem/n22716 , \u_a23_mem/n22709 , \u_a23_mem/n22702 ,
         \u_a23_mem/n22701 , \u_a23_mem/n22700 , \u_a23_mem/n22693 ,
         \u_a23_mem/n22686 , \u_a23_mem/n22685 , \u_a23_mem/n22678 ,
         \u_a23_mem/n22671 , \u_a23_mem/n22670 , \u_a23_mem/n22669 ,
         \u_a23_mem/n22668 , \u_a23_mem/n22661 , \u_a23_mem/n22654 ,
         \u_a23_mem/n22653 , \u_a23_mem/n22646 , \u_a23_mem/n22639 ,
         \u_a23_mem/n22638 , \u_a23_mem/n22637 , \u_a23_mem/n22630 ,
         \u_a23_mem/n22623 , \u_a23_mem/n22622 , \u_a23_mem/n22615 ,
         \u_a23_mem/n22608 , \u_a23_mem/n22607 , \u_a23_mem/n22606 ,
         \u_a23_mem/n22605 , \u_a23_mem/n22598 , \u_a23_mem/n22591 ,
         \u_a23_mem/n22590 , \u_a23_mem/n22583 , \u_a23_mem/n22576 ,
         \u_a23_mem/n22575 , \u_a23_mem/n22574 , \u_a23_mem/n22567 ,
         \u_a23_mem/n22560 , \u_a23_mem/n22559 , \u_a23_mem/n22552 ,
         \u_a23_mem/n22545 , \u_a23_mem/n22544 , \u_a23_mem/n22543 ,
         \u_a23_mem/n22542 , \u_a23_mem/n22535 , \u_a23_mem/n22528 ,
         \u_a23_mem/n22527 , \u_a23_mem/n22520 , \u_a23_mem/n22513 ,
         \u_a23_mem/n22512 , \u_a23_mem/n22511 , \u_a23_mem/n22504 ,
         \u_a23_mem/n22497 , \u_a23_mem/n22496 , \u_a23_mem/n22489 ,
         \u_a23_mem/n22482 , \u_a23_mem/n22481 , \u_a23_mem/n22480 ,
         \u_a23_mem/n22479 , \u_a23_mem/n22472 , \u_a23_mem/n22465 ,
         \u_a23_mem/n22464 , \u_a23_mem/n22457 , \u_a23_mem/n22450 ,
         \u_a23_mem/n22449 , \u_a23_mem/n22448 , \u_a23_mem/n22441 ,
         \u_a23_mem/n22434 , \u_a23_mem/n22433 , \u_a23_mem/n22426 ,
         \u_a23_mem/n22419 , \u_a23_mem/n22418 , \u_a23_mem/n22417 ,
         \u_a23_mem/n22416 , \u_a23_mem/n22409 , \u_a23_mem/n22402 ,
         \u_a23_mem/n22401 , \u_a23_mem/n22394 , \u_a23_mem/n22387 ,
         \u_a23_mem/n22386 , \u_a23_mem/n22385 , \u_a23_mem/n22378 ,
         \u_a23_mem/n22371 , \u_a23_mem/n22370 , \u_a23_mem/n22363 ,
         \u_a23_mem/n22356 , \u_a23_mem/n22355 , \u_a23_mem/n22354 ,
         \u_a23_mem/n22353 , \u_a23_mem/n22346 , \u_a23_mem/n22339 ,
         \u_a23_mem/n22338 , \u_a23_mem/n22331 , \u_a23_mem/n22324 ,
         \u_a23_mem/n22323 , \u_a23_mem/n22322 , \u_a23_mem/n22315 ,
         \u_a23_mem/n22308 , \u_a23_mem/n22307 , \u_a23_mem/n22300 ,
         \u_a23_mem/n22293 , \u_a23_mem/n22292 , \u_a23_mem/n22291 ,
         \u_a23_mem/n22290 , \u_a23_mem/n22283 , \u_a23_mem/n22276 ,
         \u_a23_mem/n22275 , \u_a23_mem/n22268 , \u_a23_mem/n22261 ,
         \u_a23_mem/n22260 , \u_a23_mem/n22259 , \u_a23_mem/n22252 ,
         \u_a23_mem/n22245 , \u_a23_mem/n22244 , \u_a23_mem/n22237 ,
         \u_a23_mem/n22230 , \u_a23_mem/n22229 , \u_a23_mem/n22228 ,
         \u_a23_mem/n22227 , \u_a23_mem/n22220 , \u_a23_mem/n22213 ,
         \u_a23_mem/n22212 , \u_a23_mem/n22205 , \u_a23_mem/n22198 ,
         \u_a23_mem/n22197 , \u_a23_mem/n22196 , \u_a23_mem/n22189 ,
         \u_a23_mem/n22182 , \u_a23_mem/n22181 , \u_a23_mem/n22174 ,
         \u_a23_mem/n22167 , \u_a23_mem/n22166 , \u_a23_mem/n22165 ,
         \u_a23_mem/n22164 , \u_a23_mem/n22157 , \u_a23_mem/n22150 ,
         \u_a23_mem/n22149 , \u_a23_mem/n22142 , \u_a23_mem/n22135 ,
         \u_a23_mem/n22134 , \u_a23_mem/n22133 , \u_a23_mem/n22126 ,
         \u_a23_mem/n22119 , \u_a23_mem/n22118 , \u_a23_mem/n22111 ,
         \u_a23_mem/n22104 , \u_a23_mem/n22103 , \u_a23_mem/n22102 ,
         \u_a23_mem/n22101 , \u_a23_mem/n22094 , \u_a23_mem/n22087 ,
         \u_a23_mem/n22086 , \u_a23_mem/n22079 , \u_a23_mem/n22072 ,
         \u_a23_mem/n22071 , \u_a23_mem/n22070 , \u_a23_mem/n22063 ,
         \u_a23_mem/n22056 , \u_a23_mem/n22055 , \u_a23_mem/n22048 ,
         \u_a23_mem/n22041 , \u_a23_mem/n22040 , \u_a23_mem/n22039 ,
         \u_a23_mem/n22038 , \u_a23_mem/n22031 , \u_a23_mem/n22024 ,
         \u_a23_mem/n22023 , \u_a23_mem/n22016 , \u_a23_mem/n22009 ,
         \u_a23_mem/n22008 , \u_a23_mem/n22007 , \u_a23_mem/n22000 ,
         \u_a23_mem/n21993 , \u_a23_mem/n21992 , \u_a23_mem/n21985 ,
         \u_a23_mem/n21978 , \u_a23_mem/n21977 , \u_a23_mem/n21976 ,
         \u_a23_mem/n21975 , \u_a23_mem/n21968 , \u_a23_mem/n21961 ,
         \u_a23_mem/n21960 , \u_a23_mem/n21953 , \u_a23_mem/n21946 ,
         \u_a23_mem/n21945 , \u_a23_mem/n21944 , \u_a23_mem/n21937 ,
         \u_a23_mem/n21930 , \u_a23_mem/n21929 , \u_a23_mem/n21922 ,
         \u_a23_mem/n21915 , \u_a23_mem/n21914 , \u_a23_mem/n21913 ,
         \u_a23_mem/n21912 , \u_a23_mem/n21905 , \u_a23_mem/n21898 ,
         \u_a23_mem/n21897 , \u_a23_mem/n21890 , \u_a23_mem/n21883 ,
         \u_a23_mem/n21882 , \u_a23_mem/n21881 , \u_a23_mem/n21874 ,
         \u_a23_mem/n21867 , \u_a23_mem/n21866 , \u_a23_mem/n21859 ,
         \u_a23_mem/n21731 , \u_a23_mem/n21730 , \u_a23_mem/n21729 ,
         \u_a23_mem/n21728 , \u_a23_mem/n21727 , \u_a23_mem/n21726 ,
         \u_a23_mem/n21725 , \u_a23_mem/n21724 , \u_a23_mem/n21723 ,
         \u_a23_mem/n21722 , \u_a23_mem/n21721 , \u_a23_mem/n21720 ,
         \u_a23_mem/n21719 , \u_a23_mem/n21718 , \u_a23_mem/n21716 ,
         \u_a23_mem/n21715 , \u_a23_mem/n21714 , \u_a23_mem/n21713 ,
         \u_a23_mem/n21712 , \u_a23_mem/n21711 , \u_a23_mem/n21710 ,
         \u_a23_mem/n21702 , \u_a23_mem/n21701 , \u_a23_mem/n21700 ,
         \u_a23_mem/n21699 , \u_a23_mem/n21698 , \u_a23_mem/n21697 ,
         \u_a23_mem/n21696 , \u_a23_mem/n21695 , \u_a23_mem/n21694 ,
         \u_a23_mem/n21693 , \u_a23_mem/n21692 , \u_a23_mem/n21691 ,
         \u_a23_mem/n21690 , \u_a23_mem/n21689 , \u_a23_mem/n21687 ,
         \u_a23_mem/n21686 , \u_a23_mem/n21685 , \u_a23_mem/n21684 ,
         \u_a23_mem/n21683 , \u_a23_mem/n21682 , \u_a23_mem/n21681 ,
         \u_a23_mem/n21673 , \u_a23_mem/n21672 , \u_a23_mem/n21671 ,
         \u_a23_mem/n21670 , \u_a23_mem/n21669 , \u_a23_mem/n21668 ,
         \u_a23_mem/n21667 , \u_a23_mem/n21666 , \u_a23_mem/n21665 ,
         \u_a23_mem/n21664 , \u_a23_mem/n21663 , \u_a23_mem/n21662 ,
         \u_a23_mem/n21661 , \u_a23_mem/n21660 , \u_a23_mem/n21658 ,
         \u_a23_mem/n21657 , \u_a23_mem/n21656 , \u_a23_mem/n21655 ,
         \u_a23_mem/n21654 , \u_a23_mem/n21653 , \u_a23_mem/n21652 ,
         \u_a23_mem/n21644 , \u_a23_mem/n21643 , \u_a23_mem/n21642 ,
         \u_a23_mem/n21641 , \u_a23_mem/n21640 , \u_a23_mem/n21639 ,
         \u_a23_mem/n21638 , \u_a23_mem/n21637 , \u_a23_mem/n21636 ,
         \u_a23_mem/n21635 , \u_a23_mem/n21634 , \u_a23_mem/n21633 ,
         \u_a23_mem/n21632 , \u_a23_mem/n21631 , \u_a23_mem/n21629 ,
         \u_a23_mem/n21628 , \u_a23_mem/n21627 , \u_a23_mem/n21626 ,
         \u_a23_mem/n21625 , \u_a23_mem/n21624 , \u_a23_mem/n21623 ,
         \u_a23_mem/n21615 , \u_a23_mem/n21614 , \u_a23_mem/n21613 ,
         \u_a23_mem/n21612 , \u_a23_mem/n21611 , \u_a23_mem/n21610 ,
         \u_a23_mem/n21609 , \u_a23_mem/n21608 , \u_a23_mem/n21607 ,
         \u_a23_mem/n21606 , \u_a23_mem/n21605 , \u_a23_mem/n21604 ,
         \u_a23_mem/n21603 , \u_a23_mem/n21602 , \u_a23_mem/n21600 ,
         \u_a23_mem/n21599 , \u_a23_mem/n21598 , \u_a23_mem/n21597 ,
         \u_a23_mem/n21596 , \u_a23_mem/n21595 , \u_a23_mem/n21594 ,
         \u_a23_mem/n21586 , \u_a23_mem/n21585 , \u_a23_mem/n21584 ,
         \u_a23_mem/n21583 , \u_a23_mem/n21582 , \u_a23_mem/n21581 ,
         \u_a23_mem/n21580 , \u_a23_mem/n21579 , \u_a23_mem/n21578 ,
         \u_a23_mem/n21577 , \u_a23_mem/n21576 , \u_a23_mem/n21575 ,
         \u_a23_mem/n21574 , \u_a23_mem/n21573 , \u_a23_mem/n21571 ,
         \u_a23_mem/n21570 , \u_a23_mem/n21569 , \u_a23_mem/n21568 ,
         \u_a23_mem/n21567 , \u_a23_mem/n21566 , \u_a23_mem/n21565 ,
         \u_a23_mem/n21557 , \u_a23_mem/n21556 , \u_a23_mem/n21555 ,
         \u_a23_mem/n21554 , \u_a23_mem/n21553 , \u_a23_mem/n21552 ,
         \u_a23_mem/n21551 , \u_a23_mem/n21550 , \u_a23_mem/n21549 ,
         \u_a23_mem/n21548 , \u_a23_mem/n21547 , \u_a23_mem/n21546 ,
         \u_a23_mem/n21545 , \u_a23_mem/n21544 , \u_a23_mem/n21542 ,
         \u_a23_mem/n21541 , \u_a23_mem/n21540 , \u_a23_mem/n21539 ,
         \u_a23_mem/n21538 , \u_a23_mem/n21537 , \u_a23_mem/n21536 ,
         \u_a23_mem/n21528 , \u_a23_mem/n21527 , \u_a23_mem/n21526 ,
         \u_a23_mem/n21525 , \u_a23_mem/n21524 , \u_a23_mem/n21523 ,
         \u_a23_mem/n21522 , \u_a23_mem/n21521 , \u_a23_mem/n21520 ,
         \u_a23_mem/n21519 , \u_a23_mem/n21518 , \u_a23_mem/n21517 ,
         \u_a23_mem/n21516 , \u_a23_mem/n21515 , \u_a23_mem/n21513 ,
         \u_a23_mem/n21512 , \u_a23_mem/n21511 , \u_a23_mem/n21510 ,
         \u_a23_mem/n21509 , \u_a23_mem/n21508 , \u_a23_mem/n21507 ,
         \u_a23_mem/n21475 , \u_a23_mem/n21474 , \u_a23_mem/n21473 ,
         \u_a23_mem/n21472 , \u_a23_mem/n21471 , \u_a23_mem/n21470 ,
         \u_a23_mem/n21469 , \u_a23_mem/n21468 , \u_a23_mem/n21467 ,
         \u_a23_mem/n21466 , \u_a23_mem/n21465 , \u_a23_mem/n21464 ,
         \u_a23_mem/n21463 , \u_a23_mem/n21462 , \u_a23_mem/n21460 ,
         \u_a23_mem/n21459 , \u_a23_mem/n21458 , \u_a23_mem/n21457 ,
         \u_a23_mem/n21456 , \u_a23_mem/n21455 , \u_a23_mem/n21454 ,
         \u_a23_mem/n21446 , \u_a23_mem/n21445 , \u_a23_mem/n21444 ,
         \u_a23_mem/n21443 , \u_a23_mem/n21442 , \u_a23_mem/n21441 ,
         \u_a23_mem/n21440 , \u_a23_mem/n21439 , \u_a23_mem/n21438 ,
         \u_a23_mem/n21437 , \u_a23_mem/n21436 , \u_a23_mem/n21435 ,
         \u_a23_mem/n21434 , \u_a23_mem/n21433 , \u_a23_mem/n21431 ,
         \u_a23_mem/n21430 , \u_a23_mem/n21429 , \u_a23_mem/n21428 ,
         \u_a23_mem/n21427 , \u_a23_mem/n21426 , \u_a23_mem/n21425 ,
         \u_a23_mem/n21417 , \u_a23_mem/n21416 , \u_a23_mem/n21415 ,
         \u_a23_mem/n21414 , \u_a23_mem/n21413 , \u_a23_mem/n21412 ,
         \u_a23_mem/n21411 , \u_a23_mem/n21410 , \u_a23_mem/n21409 ,
         \u_a23_mem/n21408 , \u_a23_mem/n21407 , \u_a23_mem/n21406 ,
         \u_a23_mem/n21405 , \u_a23_mem/n21404 , \u_a23_mem/n21402 ,
         \u_a23_mem/n21401 , \u_a23_mem/n21400 , \u_a23_mem/n21399 ,
         \u_a23_mem/n21398 , \u_a23_mem/n21397 , \u_a23_mem/n21396 ,
         \u_a23_mem/n21388 , \u_a23_mem/n21387 , \u_a23_mem/n21386 ,
         \u_a23_mem/n21385 , \u_a23_mem/n21384 , \u_a23_mem/n21383 ,
         \u_a23_mem/n21382 , \u_a23_mem/n21381 , \u_a23_mem/n21380 ,
         \u_a23_mem/n21379 , \u_a23_mem/n21378 , \u_a23_mem/n21377 ,
         \u_a23_mem/n21376 , \u_a23_mem/n21375 , \u_a23_mem/n21373 ,
         \u_a23_mem/n21372 , \u_a23_mem/n21371 , \u_a23_mem/n21370 ,
         \u_a23_mem/n21369 , \u_a23_mem/n21368 , \u_a23_mem/n21367 ,
         \u_a23_mem/n21359 , \u_a23_mem/n21358 , \u_a23_mem/n21357 ,
         \u_a23_mem/n21356 , \u_a23_mem/n21355 , \u_a23_mem/n21354 ,
         \u_a23_mem/n21353 , \u_a23_mem/n21352 , \u_a23_mem/n21351 ,
         \u_a23_mem/n21350 , \u_a23_mem/n21349 , \u_a23_mem/n21348 ,
         \u_a23_mem/n21347 , \u_a23_mem/n21346 , \u_a23_mem/n21344 ,
         \u_a23_mem/n21343 , \u_a23_mem/n21342 , \u_a23_mem/n21341 ,
         \u_a23_mem/n21340 , \u_a23_mem/n21339 , \u_a23_mem/n21338 ,
         \u_a23_mem/n21330 , \u_a23_mem/n21329 , \u_a23_mem/n21328 ,
         \u_a23_mem/n21327 , \u_a23_mem/n21326 , \u_a23_mem/n21325 ,
         \u_a23_mem/n21324 , \u_a23_mem/n21323 , \u_a23_mem/n21322 ,
         \u_a23_mem/n21321 , \u_a23_mem/n21320 , \u_a23_mem/n21319 ,
         \u_a23_mem/n21318 , \u_a23_mem/n21317 , \u_a23_mem/n21315 ,
         \u_a23_mem/n21314 , \u_a23_mem/n21313 , \u_a23_mem/n21312 ,
         \u_a23_mem/n21311 , \u_a23_mem/n21310 , \u_a23_mem/n21309 ,
         \u_a23_mem/n21301 , \u_a23_mem/n21300 , \u_a23_mem/n21299 ,
         \u_a23_mem/n21298 , \u_a23_mem/n21297 , \u_a23_mem/n21296 ,
         \u_a23_mem/n21295 , \u_a23_mem/n21294 , \u_a23_mem/n21293 ,
         \u_a23_mem/n21292 , \u_a23_mem/n21291 , \u_a23_mem/n21290 ,
         \u_a23_mem/n21289 , \u_a23_mem/n21288 , \u_a23_mem/n21286 ,
         \u_a23_mem/n21285 , \u_a23_mem/n21284 , \u_a23_mem/n21283 ,
         \u_a23_mem/n21282 , \u_a23_mem/n21281 , \u_a23_mem/n21280 ,
         \u_a23_mem/n21272 , \u_a23_mem/n21271 , \u_a23_mem/n21270 ,
         \u_a23_mem/n21269 , \u_a23_mem/n21268 , \u_a23_mem/n21267 ,
         \u_a23_mem/n21266 , \u_a23_mem/n21265 , \u_a23_mem/n21264 ,
         \u_a23_mem/n21263 , \u_a23_mem/n21262 , \u_a23_mem/n21261 ,
         \u_a23_mem/n21260 , \u_a23_mem/n21259 , \u_a23_mem/n21257 ,
         \u_a23_mem/n21256 , \u_a23_mem/n21255 , \u_a23_mem/n21254 ,
         \u_a23_mem/n21253 , \u_a23_mem/n21252 , \u_a23_mem/n21251 ,
         \u_a23_mem/n21219 , \u_a23_mem/n21218 , \u_a23_mem/n21217 ,
         \u_a23_mem/n21216 , \u_a23_mem/n21215 , \u_a23_mem/n21214 ,
         \u_a23_mem/n21213 , \u_a23_mem/n21212 , \u_a23_mem/n21211 ,
         \u_a23_mem/n21210 , \u_a23_mem/n21209 , \u_a23_mem/n21208 ,
         \u_a23_mem/n21207 , \u_a23_mem/n21206 , \u_a23_mem/n21204 ,
         \u_a23_mem/n21203 , \u_a23_mem/n21202 , \u_a23_mem/n21201 ,
         \u_a23_mem/n21200 , \u_a23_mem/n21199 , \u_a23_mem/n21198 ,
         \u_a23_mem/n21190 , \u_a23_mem/n21189 , \u_a23_mem/n21188 ,
         \u_a23_mem/n21187 , \u_a23_mem/n21186 , \u_a23_mem/n21185 ,
         \u_a23_mem/n21184 , \u_a23_mem/n21183 , \u_a23_mem/n21182 ,
         \u_a23_mem/n21181 , \u_a23_mem/n21180 , \u_a23_mem/n21179 ,
         \u_a23_mem/n21178 , \u_a23_mem/n21177 , \u_a23_mem/n21175 ,
         \u_a23_mem/n21174 , \u_a23_mem/n21173 , \u_a23_mem/n21172 ,
         \u_a23_mem/n21171 , \u_a23_mem/n21170 , \u_a23_mem/n21169 ,
         \u_a23_mem/n21161 , \u_a23_mem/n21160 , \u_a23_mem/n21159 ,
         \u_a23_mem/n21158 , \u_a23_mem/n21157 , \u_a23_mem/n21156 ,
         \u_a23_mem/n21155 , \u_a23_mem/n21154 , \u_a23_mem/n21153 ,
         \u_a23_mem/n21152 , \u_a23_mem/n21151 , \u_a23_mem/n21150 ,
         \u_a23_mem/n21149 , \u_a23_mem/n21148 , \u_a23_mem/n21146 ,
         \u_a23_mem/n21145 , \u_a23_mem/n21144 , \u_a23_mem/n21143 ,
         \u_a23_mem/n21142 , \u_a23_mem/n21141 , \u_a23_mem/n21140 ,
         \u_a23_mem/n21132 , \u_a23_mem/n21131 , \u_a23_mem/n21130 ,
         \u_a23_mem/n21129 , \u_a23_mem/n21128 , \u_a23_mem/n21127 ,
         \u_a23_mem/n21126 , \u_a23_mem/n21125 , \u_a23_mem/n21124 ,
         \u_a23_mem/n21123 , \u_a23_mem/n21122 , \u_a23_mem/n21121 ,
         \u_a23_mem/n21120 , \u_a23_mem/n21119 , \u_a23_mem/n21117 ,
         \u_a23_mem/n21116 , \u_a23_mem/n21115 , \u_a23_mem/n21114 ,
         \u_a23_mem/n21113 , \u_a23_mem/n21112 , \u_a23_mem/n21111 ,
         \u_a23_mem/n21103 , \u_a23_mem/n21102 , \u_a23_mem/n21101 ,
         \u_a23_mem/n21100 , \u_a23_mem/n21099 , \u_a23_mem/n21098 ,
         \u_a23_mem/n21097 , \u_a23_mem/n21096 , \u_a23_mem/n21095 ,
         \u_a23_mem/n21094 , \u_a23_mem/n21093 , \u_a23_mem/n21092 ,
         \u_a23_mem/n21091 , \u_a23_mem/n21090 , \u_a23_mem/n21088 ,
         \u_a23_mem/n21087 , \u_a23_mem/n21086 , \u_a23_mem/n21085 ,
         \u_a23_mem/n21084 , \u_a23_mem/n21083 , \u_a23_mem/n21082 ,
         \u_a23_mem/n21074 , \u_a23_mem/n21073 , \u_a23_mem/n21072 ,
         \u_a23_mem/n21071 , \u_a23_mem/n21070 , \u_a23_mem/n21069 ,
         \u_a23_mem/n21068 , \u_a23_mem/n21067 , \u_a23_mem/n21066 ,
         \u_a23_mem/n21065 , \u_a23_mem/n21064 , \u_a23_mem/n21063 ,
         \u_a23_mem/n21062 , \u_a23_mem/n21061 , \u_a23_mem/n21059 ,
         \u_a23_mem/n21058 , \u_a23_mem/n21057 , \u_a23_mem/n21056 ,
         \u_a23_mem/n21055 , \u_a23_mem/n21054 , \u_a23_mem/n21053 ,
         \u_a23_mem/n21045 , \u_a23_mem/n21044 , \u_a23_mem/n21043 ,
         \u_a23_mem/n21042 , \u_a23_mem/n21041 , \u_a23_mem/n21040 ,
         \u_a23_mem/n21039 , \u_a23_mem/n21038 , \u_a23_mem/n21037 ,
         \u_a23_mem/n21036 , \u_a23_mem/n21035 , \u_a23_mem/n21034 ,
         \u_a23_mem/n21033 , \u_a23_mem/n21032 , \u_a23_mem/n21030 ,
         \u_a23_mem/n21029 , \u_a23_mem/n21028 , \u_a23_mem/n21027 ,
         \u_a23_mem/n21026 , \u_a23_mem/n21025 , \u_a23_mem/n21024 ,
         \u_a23_mem/n21016 , \u_a23_mem/n21015 , \u_a23_mem/n21014 ,
         \u_a23_mem/n21013 , \u_a23_mem/n21012 , \u_a23_mem/n21011 ,
         \u_a23_mem/n21010 , \u_a23_mem/n21009 , \u_a23_mem/n21008 ,
         \u_a23_mem/n21007 , \u_a23_mem/n21006 , \u_a23_mem/n21005 ,
         \u_a23_mem/n21004 , \u_a23_mem/n21003 , \u_a23_mem/n21001 ,
         \u_a23_mem/n21000 , \u_a23_mem/n20999 , \u_a23_mem/n20998 ,
         \u_a23_mem/n20997 , \u_a23_mem/n20996 , \u_a23_mem/n20995 ,
         \u_a23_mem/n20963 , \u_a23_mem/n20962 , \u_a23_mem/n20961 ,
         \u_a23_mem/n20960 , \u_a23_mem/n20959 , \u_a23_mem/n20958 ,
         \u_a23_mem/n20957 , \u_a23_mem/n20956 , \u_a23_mem/n20955 ,
         \u_a23_mem/n20954 , \u_a23_mem/n20953 , \u_a23_mem/n20952 ,
         \u_a23_mem/n20951 , \u_a23_mem/n20950 , \u_a23_mem/n20948 ,
         \u_a23_mem/n20947 , \u_a23_mem/n20946 , \u_a23_mem/n20945 ,
         \u_a23_mem/n20944 , \u_a23_mem/n20943 , \u_a23_mem/n20942 ,
         \u_a23_mem/n20934 , \u_a23_mem/n20933 , \u_a23_mem/n20932 ,
         \u_a23_mem/n20931 , \u_a23_mem/n20930 , \u_a23_mem/n20929 ,
         \u_a23_mem/n20928 , \u_a23_mem/n20927 , \u_a23_mem/n20926 ,
         \u_a23_mem/n20925 , \u_a23_mem/n20924 , \u_a23_mem/n20923 ,
         \u_a23_mem/n20922 , \u_a23_mem/n20921 , \u_a23_mem/n20919 ,
         \u_a23_mem/n20918 , \u_a23_mem/n20917 , \u_a23_mem/n20916 ,
         \u_a23_mem/n20915 , \u_a23_mem/n20914 , \u_a23_mem/n20913 ,
         \u_a23_mem/n20905 , \u_a23_mem/n20904 , \u_a23_mem/n20903 ,
         \u_a23_mem/n20902 , \u_a23_mem/n20901 , \u_a23_mem/n20900 ,
         \u_a23_mem/n20899 , \u_a23_mem/n20898 , \u_a23_mem/n20897 ,
         \u_a23_mem/n20896 , \u_a23_mem/n20895 , \u_a23_mem/n20894 ,
         \u_a23_mem/n20893 , \u_a23_mem/n20892 , \u_a23_mem/n20890 ,
         \u_a23_mem/n20889 , \u_a23_mem/n20888 , \u_a23_mem/n20887 ,
         \u_a23_mem/n20886 , \u_a23_mem/n20885 , \u_a23_mem/n20884 ,
         \u_a23_mem/n20876 , \u_a23_mem/n20875 , \u_a23_mem/n20874 ,
         \u_a23_mem/n20873 , \u_a23_mem/n20872 , \u_a23_mem/n20871 ,
         \u_a23_mem/n20870 , \u_a23_mem/n20869 , \u_a23_mem/n20868 ,
         \u_a23_mem/n20867 , \u_a23_mem/n20866 , \u_a23_mem/n20865 ,
         \u_a23_mem/n20864 , \u_a23_mem/n20863 , \u_a23_mem/n20861 ,
         \u_a23_mem/n20860 , \u_a23_mem/n20859 , \u_a23_mem/n20858 ,
         \u_a23_mem/n20857 , \u_a23_mem/n20856 , \u_a23_mem/n20855 ,
         \u_a23_mem/n20847 , \u_a23_mem/n20846 , \u_a23_mem/n20845 ,
         \u_a23_mem/n20844 , \u_a23_mem/n20843 , \u_a23_mem/n20842 ,
         \u_a23_mem/n20841 , \u_a23_mem/n20840 , \u_a23_mem/n20839 ,
         \u_a23_mem/n20838 , \u_a23_mem/n20837 , \u_a23_mem/n20836 ,
         \u_a23_mem/n20835 , \u_a23_mem/n20834 , \u_a23_mem/n20832 ,
         \u_a23_mem/n20831 , \u_a23_mem/n20830 , \u_a23_mem/n20829 ,
         \u_a23_mem/n20828 , \u_a23_mem/n20827 , \u_a23_mem/n20826 ,
         \u_a23_mem/n20818 , \u_a23_mem/n20817 , \u_a23_mem/n20816 ,
         \u_a23_mem/n20815 , \u_a23_mem/n20814 , \u_a23_mem/n20813 ,
         \u_a23_mem/n20812 , \u_a23_mem/n20811 , \u_a23_mem/n20810 ,
         \u_a23_mem/n20809 , \u_a23_mem/n20808 , \u_a23_mem/n20807 ,
         \u_a23_mem/n20806 , \u_a23_mem/n20805 , \u_a23_mem/n20803 ,
         \u_a23_mem/n20802 , \u_a23_mem/n20801 , \u_a23_mem/n20800 ,
         \u_a23_mem/n20799 , \u_a23_mem/n20798 , \u_a23_mem/n20797 ,
         \u_a23_mem/n20789 , \u_a23_mem/n20788 , \u_a23_mem/n20787 ,
         \u_a23_mem/n20786 , \u_a23_mem/n20785 , \u_a23_mem/n20784 ,
         \u_a23_mem/n20783 , \u_a23_mem/n20782 , \u_a23_mem/n20781 ,
         \u_a23_mem/n20780 , \u_a23_mem/n20779 , \u_a23_mem/n20778 ,
         \u_a23_mem/n20777 , \u_a23_mem/n20776 , \u_a23_mem/n20774 ,
         \u_a23_mem/n20773 , \u_a23_mem/n20772 , \u_a23_mem/n20771 ,
         \u_a23_mem/n20770 , \u_a23_mem/n20769 , \u_a23_mem/n20768 ,
         \u_a23_mem/n20760 , \u_a23_mem/n20759 , \u_a23_mem/n20758 ,
         \u_a23_mem/n20757 , \u_a23_mem/n20756 , \u_a23_mem/n20755 ,
         \u_a23_mem/n20754 , \u_a23_mem/n20753 , \u_a23_mem/n20752 ,
         \u_a23_mem/n20751 , \u_a23_mem/n20750 , \u_a23_mem/n20749 ,
         \u_a23_mem/n20748 , \u_a23_mem/n20747 , \u_a23_mem/n20745 ,
         \u_a23_mem/n20744 , \u_a23_mem/n20743 , \u_a23_mem/n20742 ,
         \u_a23_mem/n20741 , \u_a23_mem/n20740 , \u_a23_mem/n20739 ,
         \u_a23_mem/n20651 , \u_a23_mem/n20650 , \u_a23_mem/n20649 ,
         \u_a23_mem/n20648 , \u_a23_mem/n20647 , \u_a23_mem/n20646 ,
         \u_a23_mem/n20645 , \u_a23_mem/n20644 , \u_a23_mem/n20643 ,
         \u_a23_mem/n20642 , \u_a23_mem/n20641 , \u_a23_mem/n20640 ,
         \u_a23_mem/n20639 , \u_a23_mem/n20638 , \u_a23_mem/n20637 ,
         \u_a23_mem/n20636 , \u_a23_mem/n20635 , \u_a23_mem/n20634 ,
         \u_a23_mem/n20633 , \u_a23_mem/n20632 , \u_a23_mem/n20631 ,
         \u_a23_mem/n20630 , \u_a23_mem/n20629 , \u_a23_mem/n20628 ,
         \u_a23_mem/n20627 , \u_a23_mem/n20626 , \u_a23_mem/n20625 ,
         \u_a23_mem/n20624 , \u_a23_mem/n20623 , \u_a23_mem/n20622 ,
         \u_a23_mem/n20621 , \u_a23_mem/n20620 , \u_a23_mem/n20619 ,
         \u_a23_mem/n20618 , \u_a23_mem/n20617 , \u_a23_mem/n20616 ,
         \u_a23_mem/n20615 , \u_a23_mem/n20614 , \u_a23_mem/n20613 ,
         \u_a23_mem/n20612 , \u_a23_mem/n20611 , \u_a23_mem/n20610 ,
         \u_a23_mem/n20609 , \u_a23_mem/n20608 , \u_a23_mem/n20607 ,
         \u_a23_mem/n20606 , \u_a23_mem/n20605 , \u_a23_mem/n20604 ,
         \u_a23_mem/n20603 , \u_a23_mem/n20602 , \u_a23_mem/n20601 ,
         \u_a23_mem/n20600 , \u_a23_mem/n20599 , \u_a23_mem/n20598 ,
         \u_a23_mem/n20597 , \u_a23_mem/n20596 , \u_a23_mem/n20595 ,
         \u_a23_mem/n20594 , \u_a23_mem/n20593 , \u_a23_mem/n20592 ,
         \u_a23_mem/n20591 , \u_a23_mem/n20590 , \u_a23_mem/n20588 ,
         \u_a23_mem/n20587 , \u_a23_mem/n20586 , \u_a23_mem/n20585 ,
         \u_a23_mem/n20584 , \u_a23_mem/n20583 , \u_a23_mem/n20582 ,
         \u_a23_mem/n20581 , \u_a23_mem/n20580 , \u_a23_mem/n20579 ,
         \u_a23_mem/n20578 , \u_a23_mem/n20577 , \u_a23_mem/n20576 ,
         \u_a23_mem/n20575 , \u_a23_mem/n20574 , \u_a23_mem/n20573 ,
         \u_a23_mem/n20572 , \u_a23_mem/n20571 , \u_a23_mem/n20570 ,
         \u_a23_mem/n20569 , \u_a23_mem/n20568 , \u_a23_mem/n20567 ,
         \u_a23_mem/n20566 , \u_a23_mem/n20565 , \u_a23_mem/n20564 ,
         \u_a23_mem/n20563 , \u_a23_mem/n20562 , \u_a23_mem/n20561 ,
         \u_a23_mem/n20560 , \u_a23_mem/n20559 , \u_a23_mem/n20558 ,
         \u_a23_mem/n20526 , \u_a23_mem/n20525 , \u_a23_mem/n20524 ,
         \u_a23_mem/n20523 , \u_a23_mem/n20522 , \u_a23_mem/n20521 ,
         \u_a23_mem/n20520 , \u_a23_mem/n20519 , \u_a23_mem/n20518 ,
         \u_a23_mem/n20517 , \u_a23_mem/n20516 , \u_a23_mem/n20515 ,
         \u_a23_mem/n20514 , \u_a23_mem/n20513 , \u_a23_mem/n20512 ,
         \u_a23_mem/n20511 , \u_a23_mem/n20510 , \u_a23_mem/n20509 ,
         \u_a23_mem/n20508 , \u_a23_mem/n20507 , \u_a23_mem/n20506 ,
         \u_a23_mem/n20505 , \u_a23_mem/n20504 , \u_a23_mem/n20503 ,
         \u_a23_mem/n20502 , \u_a23_mem/n20501 , \u_a23_mem/n20500 ,
         \u_a23_mem/n20499 , \u_a23_mem/n20498 , \u_a23_mem/n20497 ,
         \u_a23_mem/n20496 , \u_a23_mem/n20495 , \u_a23_mem/n20494 ,
         \u_a23_mem/n20493 , \u_a23_mem/n20492 , \u_a23_mem/n20491 ,
         \u_a23_mem/n20490 , \u_a23_mem/n20489 , \u_a23_mem/n20488 ,
         \u_a23_mem/n20487 , \u_a23_mem/n20486 , \u_a23_mem/n20485 ,
         \u_a23_mem/n20484 , \u_a23_mem/n20483 , \u_a23_mem/n20482 ,
         \u_a23_mem/n20481 , \u_a23_mem/n20480 , \u_a23_mem/n20479 ,
         \u_a23_mem/n20478 , \u_a23_mem/n20477 , \u_a23_mem/n20476 ,
         \u_a23_mem/n20475 , \u_a23_mem/n20474 , \u_a23_mem/n20473 ,
         \u_a23_mem/n20472 , \u_a23_mem/n20471 , \u_a23_mem/n20470 ,
         \u_a23_mem/n20469 , \u_a23_mem/n20468 , \u_a23_mem/n20467 ,
         \u_a23_mem/n20466 , \u_a23_mem/n20465 , \u_a23_mem/n20463 ,
         \u_a23_mem/n20462 , \u_a23_mem/n20461 , \u_a23_mem/n20460 ,
         \u_a23_mem/n20459 , \u_a23_mem/n20458 , \u_a23_mem/n20457 ,
         \u_a23_mem/n20456 , \u_a23_mem/n20455 , \u_a23_mem/n20454 ,
         \u_a23_mem/n20453 , \u_a23_mem/n20452 , \u_a23_mem/n20451 ,
         \u_a23_mem/n20450 , \u_a23_mem/n20449 , \u_a23_mem/n20448 ,
         \u_a23_mem/n20447 , \u_a23_mem/n20446 , \u_a23_mem/n20445 ,
         \u_a23_mem/n20444 , \u_a23_mem/n20443 , \u_a23_mem/n20442 ,
         \u_a23_mem/n20441 , \u_a23_mem/n20440 , \u_a23_mem/n20439 ,
         \u_a23_mem/n20438 , \u_a23_mem/n20437 , \u_a23_mem/n20436 ,
         \u_a23_mem/n20435 , \u_a23_mem/n20434 , \u_a23_mem/n20433 ,
         \u_a23_mem/n20401 , \u_a23_mem/n20400 , \u_a23_mem/n20399 ,
         \u_a23_mem/n20398 , \u_a23_mem/n20397 , \u_a23_mem/n20396 ,
         \u_a23_mem/n20395 , \u_a23_mem/n20394 , \u_a23_mem/n20393 ,
         \u_a23_mem/n20392 , \u_a23_mem/n20391 , \u_a23_mem/n20390 ,
         \u_a23_mem/n20389 , \u_a23_mem/n20388 , \u_a23_mem/n20387 ,
         \u_a23_mem/n20386 , \u_a23_mem/n20385 , \u_a23_mem/n20384 ,
         \u_a23_mem/n20383 , \u_a23_mem/n20382 , \u_a23_mem/n20381 ,
         \u_a23_mem/n20380 , \u_a23_mem/n20379 , \u_a23_mem/n20378 ,
         \u_a23_mem/n20377 , \u_a23_mem/n20376 , \u_a23_mem/n20375 ,
         \u_a23_mem/n20374 , \u_a23_mem/n20373 , \u_a23_mem/n20372 ,
         \u_a23_mem/n20371 , \u_a23_mem/n20370 , \u_a23_mem/n20369 ,
         \u_a23_mem/n20368 , \u_a23_mem/n20367 , \u_a23_mem/n20366 ,
         \u_a23_mem/n20365 , \u_a23_mem/n20364 , \u_a23_mem/n20363 ,
         \u_a23_mem/n20362 , \u_a23_mem/n20361 , \u_a23_mem/n20360 ,
         \u_a23_mem/n20359 , \u_a23_mem/n20358 , \u_a23_mem/n20357 ,
         \u_a23_mem/n20356 , \u_a23_mem/n20355 , \u_a23_mem/n20354 ,
         \u_a23_mem/n20353 , \u_a23_mem/n20352 , \u_a23_mem/n20351 ,
         \u_a23_mem/n20350 , \u_a23_mem/n20349 , \u_a23_mem/n20348 ,
         \u_a23_mem/n20347 , \u_a23_mem/n20346 , \u_a23_mem/n20345 ,
         \u_a23_mem/n20344 , \u_a23_mem/n20343 , \u_a23_mem/n20342 ,
         \u_a23_mem/n20341 , \u_a23_mem/n20340 , \u_a23_mem/n20338 ,
         \u_a23_mem/n20337 , \u_a23_mem/n20336 , \u_a23_mem/n20335 ,
         \u_a23_mem/n20334 , \u_a23_mem/n20333 , \u_a23_mem/n20332 ,
         \u_a23_mem/n20331 , \u_a23_mem/n20330 , \u_a23_mem/n20329 ,
         \u_a23_mem/n20328 , \u_a23_mem/n20327 , \u_a23_mem/n20326 ,
         \u_a23_mem/n20325 , \u_a23_mem/n20324 , \u_a23_mem/n20323 ,
         \u_a23_mem/n20322 , \u_a23_mem/n20321 , \u_a23_mem/n20320 ,
         \u_a23_mem/n20319 , \u_a23_mem/n20318 , \u_a23_mem/n20317 ,
         \u_a23_mem/n20316 , \u_a23_mem/n20315 , \u_a23_mem/n20314 ,
         \u_a23_mem/n20313 , \u_a23_mem/n20312 , \u_a23_mem/n20311 ,
         \u_a23_mem/n20310 , \u_a23_mem/n20309 , \u_a23_mem/n20308 ,
         \u_a23_mem/n20276 , \u_a23_mem/n20275 , \u_a23_mem/n20274 ,
         \u_a23_mem/n20273 , \u_a23_mem/n20272 , \u_a23_mem/n20271 ,
         \u_a23_mem/n20270 , \u_a23_mem/n20269 , \u_a23_mem/n20268 ,
         \u_a23_mem/n20267 , \u_a23_mem/n20266 , \u_a23_mem/n20265 ,
         \u_a23_mem/n20264 , \u_a23_mem/n20263 , \u_a23_mem/n20262 ,
         \u_a23_mem/n20261 , \u_a23_mem/n20260 , \u_a23_mem/n20259 ,
         \u_a23_mem/n20258 , \u_a23_mem/n20257 , \u_a23_mem/n20256 ,
         \u_a23_mem/n20255 , \u_a23_mem/n20254 , \u_a23_mem/n20253 ,
         \u_a23_mem/n20252 , \u_a23_mem/n20251 , \u_a23_mem/n20250 ,
         \u_a23_mem/n20249 , \u_a23_mem/n20248 , \u_a23_mem/n20247 ,
         \u_a23_mem/n20246 , \u_a23_mem/n20245 , \u_a23_mem/n20244 ,
         \u_a23_mem/n20243 , \u_a23_mem/n20242 , \u_a23_mem/n20241 ,
         \u_a23_mem/n20240 , \u_a23_mem/n20239 , \u_a23_mem/n20238 ,
         \u_a23_mem/n20237 , \u_a23_mem/n20236 , \u_a23_mem/n20235 ,
         \u_a23_mem/n20234 , \u_a23_mem/n20233 , \u_a23_mem/n20232 ,
         \u_a23_mem/n20231 , \u_a23_mem/n20230 , \u_a23_mem/n20229 ,
         \u_a23_mem/n20228 , \u_a23_mem/n20227 , \u_a23_mem/n20226 ,
         \u_a23_mem/n20225 , \u_a23_mem/n20224 , \u_a23_mem/n20223 ,
         \u_a23_mem/n20222 , \u_a23_mem/n20221 , \u_a23_mem/n20220 ,
         \u_a23_mem/n20219 , \u_a23_mem/n20218 , \u_a23_mem/n20217 ,
         \u_a23_mem/n20216 , \u_a23_mem/n20215 , \u_a23_mem/n20213 ,
         \u_a23_mem/n20212 , \u_a23_mem/n20211 , \u_a23_mem/n20210 ,
         \u_a23_mem/n20209 , \u_a23_mem/n20208 , \u_a23_mem/n20207 ,
         \u_a23_mem/n20206 , \u_a23_mem/n20205 , \u_a23_mem/n20204 ,
         \u_a23_mem/n20203 , \u_a23_mem/n20202 , \u_a23_mem/n20201 ,
         \u_a23_mem/n20200 , \u_a23_mem/n20199 , \u_a23_mem/n20198 ,
         \u_a23_mem/n20197 , \u_a23_mem/n20196 , \u_a23_mem/n20195 ,
         \u_a23_mem/n20194 , \u_a23_mem/n20193 , \u_a23_mem/n20192 ,
         \u_a23_mem/n20191 , \u_a23_mem/n20190 , \u_a23_mem/n20189 ,
         \u_a23_mem/n20188 , \u_a23_mem/n20187 , \u_a23_mem/n20186 ,
         \u_a23_mem/n20185 , \u_a23_mem/n20184 , \u_a23_mem/n20183 ,
         \u_a23_mem/n20151 , \u_a23_mem/n20150 , \u_a23_mem/n20149 ,
         \u_a23_mem/n20148 , \u_a23_mem/n20147 , \u_a23_mem/n20146 ,
         \u_a23_mem/n20145 , \u_a23_mem/n20144 , \u_a23_mem/n20143 ,
         \u_a23_mem/n20142 , \u_a23_mem/n20141 , \u_a23_mem/n20140 ,
         \u_a23_mem/n20139 , \u_a23_mem/n20138 , \u_a23_mem/n20137 ,
         \u_a23_mem/n20136 , \u_a23_mem/n20135 , \u_a23_mem/n20134 ,
         \u_a23_mem/n20133 , \u_a23_mem/n20132 , \u_a23_mem/n20131 ,
         \u_a23_mem/n20130 , \u_a23_mem/n20129 , \u_a23_mem/n20128 ,
         \u_a23_mem/n20127 , \u_a23_mem/n20126 , \u_a23_mem/n20125 ,
         \u_a23_mem/n20124 , \u_a23_mem/n20123 , \u_a23_mem/n20122 ,
         \u_a23_mem/n20121 , \u_a23_mem/n20120 , \u_a23_mem/n20119 ,
         \u_a23_mem/n20118 , \u_a23_mem/n20117 , \u_a23_mem/n20116 ,
         \u_a23_mem/n20115 , \u_a23_mem/n20114 , \u_a23_mem/n20113 ,
         \u_a23_mem/n20112 , \u_a23_mem/n20111 , \u_a23_mem/n20110 ,
         \u_a23_mem/n20109 , \u_a23_mem/n20108 , \u_a23_mem/n20107 ,
         \u_a23_mem/n20106 , \u_a23_mem/n20105 , \u_a23_mem/n20104 ,
         \u_a23_mem/n20103 , \u_a23_mem/n20102 , \u_a23_mem/n20101 ,
         \u_a23_mem/n20100 , \u_a23_mem/n20099 , \u_a23_mem/n20098 ,
         \u_a23_mem/n20097 , \u_a23_mem/n20096 , \u_a23_mem/n20095 ,
         \u_a23_mem/n20094 , \u_a23_mem/n20093 , \u_a23_mem/n20092 ,
         \u_a23_mem/n20091 , \u_a23_mem/n20090 , \u_a23_mem/n20088 ,
         \u_a23_mem/n20087 , \u_a23_mem/n20086 , \u_a23_mem/n20085 ,
         \u_a23_mem/n20084 , \u_a23_mem/n20083 , \u_a23_mem/n20082 ,
         \u_a23_mem/n20081 , \u_a23_mem/n20080 , \u_a23_mem/n20079 ,
         \u_a23_mem/n20078 , \u_a23_mem/n20077 , \u_a23_mem/n20076 ,
         \u_a23_mem/n20075 , \u_a23_mem/n20074 , \u_a23_mem/n20073 ,
         \u_a23_mem/n20072 , \u_a23_mem/n20071 , \u_a23_mem/n20070 ,
         \u_a23_mem/n20069 , \u_a23_mem/n20068 , \u_a23_mem/n20067 ,
         \u_a23_mem/n20066 , \u_a23_mem/n20065 , \u_a23_mem/n20064 ,
         \u_a23_mem/n20063 , \u_a23_mem/n20062 , \u_a23_mem/n20061 ,
         \u_a23_mem/n20060 , \u_a23_mem/n20059 , \u_a23_mem/n20058 ,
         \u_a23_mem/n20026 , \u_a23_mem/n20025 , \u_a23_mem/n20024 ,
         \u_a23_mem/n20023 , \u_a23_mem/n20022 , \u_a23_mem/n20021 ,
         \u_a23_mem/n20020 , \u_a23_mem/n20019 , \u_a23_mem/n20018 ,
         \u_a23_mem/n20017 , \u_a23_mem/n20016 , \u_a23_mem/n20015 ,
         \u_a23_mem/n20014 , \u_a23_mem/n20013 , \u_a23_mem/n20012 ,
         \u_a23_mem/n20011 , \u_a23_mem/n20010 , \u_a23_mem/n20009 ,
         \u_a23_mem/n20008 , \u_a23_mem/n20007 , \u_a23_mem/n20006 ,
         \u_a23_mem/n20005 , \u_a23_mem/n20004 , \u_a23_mem/n20003 ,
         \u_a23_mem/n20002 , \u_a23_mem/n20001 , \u_a23_mem/n20000 ,
         \u_a23_mem/n19999 , \u_a23_mem/n19998 , \u_a23_mem/n19997 ,
         \u_a23_mem/n19996 , \u_a23_mem/n19995 , \u_a23_mem/n19994 ,
         \u_a23_mem/n19993 , \u_a23_mem/n19992 , \u_a23_mem/n19991 ,
         \u_a23_mem/n19990 , \u_a23_mem/n19989 , \u_a23_mem/n19988 ,
         \u_a23_mem/n19987 , \u_a23_mem/n19986 , \u_a23_mem/n19985 ,
         \u_a23_mem/n19984 , \u_a23_mem/n19983 , \u_a23_mem/n19982 ,
         \u_a23_mem/n19981 , \u_a23_mem/n19980 , \u_a23_mem/n19979 ,
         \u_a23_mem/n19978 , \u_a23_mem/n19977 , \u_a23_mem/n19976 ,
         \u_a23_mem/n19975 , \u_a23_mem/n19974 , \u_a23_mem/n19973 ,
         \u_a23_mem/n19972 , \u_a23_mem/n19971 , \u_a23_mem/n19970 ,
         \u_a23_mem/n19969 , \u_a23_mem/n19968 , \u_a23_mem/n19967 ,
         \u_a23_mem/n19966 , \u_a23_mem/n19965 , \u_a23_mem/n19963 ,
         \u_a23_mem/n19962 , \u_a23_mem/n19961 , \u_a23_mem/n19960 ,
         \u_a23_mem/n19959 , \u_a23_mem/n19958 , \u_a23_mem/n19957 ,
         \u_a23_mem/n19956 , \u_a23_mem/n19955 , \u_a23_mem/n19954 ,
         \u_a23_mem/n19953 , \u_a23_mem/n19952 , \u_a23_mem/n19951 ,
         \u_a23_mem/n19950 , \u_a23_mem/n19949 , \u_a23_mem/n19948 ,
         \u_a23_mem/n19947 , \u_a23_mem/n19946 , \u_a23_mem/n19945 ,
         \u_a23_mem/n19944 , \u_a23_mem/n19943 , \u_a23_mem/n19942 ,
         \u_a23_mem/n19941 , \u_a23_mem/n19940 , \u_a23_mem/n19939 ,
         \u_a23_mem/n19938 , \u_a23_mem/n19937 , \u_a23_mem/n19936 ,
         \u_a23_mem/n19935 , \u_a23_mem/n19934 , \u_a23_mem/n19933 ,
         \u_a23_mem/n19901 , \u_a23_mem/n19900 , \u_a23_mem/n19899 ,
         \u_a23_mem/n19898 , \u_a23_mem/n19897 , \u_a23_mem/n19896 ,
         \u_a23_mem/n19895 , \u_a23_mem/n19894 , \u_a23_mem/n19893 ,
         \u_a23_mem/n19892 , \u_a23_mem/n19891 , \u_a23_mem/n19890 ,
         \u_a23_mem/n19889 , \u_a23_mem/n19888 , \u_a23_mem/n19887 ,
         \u_a23_mem/n19886 , \u_a23_mem/n19885 , \u_a23_mem/n19884 ,
         \u_a23_mem/n19883 , \u_a23_mem/n19882 , \u_a23_mem/n19881 ,
         \u_a23_mem/n19880 , \u_a23_mem/n19879 , \u_a23_mem/n19878 ,
         \u_a23_mem/n19877 , \u_a23_mem/n19876 , \u_a23_mem/n19875 ,
         \u_a23_mem/n19874 , \u_a23_mem/n19873 , \u_a23_mem/n19872 ,
         \u_a23_mem/n19871 , \u_a23_mem/n19870 , \u_a23_mem/n19869 ,
         \u_a23_mem/n19868 , \u_a23_mem/n19867 , \u_a23_mem/n19866 ,
         \u_a23_mem/n19865 , \u_a23_mem/n19864 , \u_a23_mem/n19863 ,
         \u_a23_mem/n19862 , \u_a23_mem/n19861 , \u_a23_mem/n19860 ,
         \u_a23_mem/n19859 , \u_a23_mem/n19858 , \u_a23_mem/n19857 ,
         \u_a23_mem/n19856 , \u_a23_mem/n19855 , \u_a23_mem/n19854 ,
         \u_a23_mem/n19853 , \u_a23_mem/n19852 , \u_a23_mem/n19851 ,
         \u_a23_mem/n19850 , \u_a23_mem/n19849 , \u_a23_mem/n19848 ,
         \u_a23_mem/n19847 , \u_a23_mem/n19846 , \u_a23_mem/n19845 ,
         \u_a23_mem/n19844 , \u_a23_mem/n19843 , \u_a23_mem/n19842 ,
         \u_a23_mem/n19841 , \u_a23_mem/n19840 , \u_a23_mem/n19838 ,
         \u_a23_mem/n19837 , \u_a23_mem/n19836 , \u_a23_mem/n19835 ,
         \u_a23_mem/n19834 , \u_a23_mem/n19833 , \u_a23_mem/n19832 ,
         \u_a23_mem/n19831 , \u_a23_mem/n19830 , \u_a23_mem/n19829 ,
         \u_a23_mem/n19828 , \u_a23_mem/n19827 , \u_a23_mem/n19826 ,
         \u_a23_mem/n19825 , \u_a23_mem/n19824 , \u_a23_mem/n19823 ,
         \u_a23_mem/n19822 , \u_a23_mem/n19821 , \u_a23_mem/n19820 ,
         \u_a23_mem/n19819 , \u_a23_mem/n19818 , \u_a23_mem/n19817 ,
         \u_a23_mem/n19816 , \u_a23_mem/n19815 , \u_a23_mem/n19814 ,
         \u_a23_mem/n19813 , \u_a23_mem/n19812 , \u_a23_mem/n19811 ,
         \u_a23_mem/n19810 , \u_a23_mem/n19809 , \u_a23_mem/n19808 ,
         \u_a23_mem/n19776 , \u_a23_mem/n19775 , \u_a23_mem/n19774 ,
         \u_a23_mem/n19773 , \u_a23_mem/n19772 , \u_a23_mem/n19771 ,
         \u_a23_mem/n19770 , \u_a23_mem/n19769 , \u_a23_mem/n19768 ,
         \u_a23_mem/n19767 , \u_a23_mem/n19766 , \u_a23_mem/n19765 ,
         \u_a23_mem/n19764 , \u_a23_mem/n19763 , \u_a23_mem/n19762 ,
         \u_a23_mem/n19761 , \u_a23_mem/n19760 , \u_a23_mem/n19759 ,
         \u_a23_mem/n19758 , \u_a23_mem/n19757 , \u_a23_mem/n19756 ,
         \u_a23_mem/n19755 , \u_a23_mem/n19754 , \u_a23_mem/n19753 ,
         \u_a23_mem/n19752 , \u_a23_mem/n19751 , \u_a23_mem/n19750 ,
         \u_a23_mem/n19749 , \u_a23_mem/n19748 , \u_a23_mem/n19747 ,
         \u_a23_mem/n19746 , \u_a23_mem/n19745 , \u_a23_mem/n19744 ,
         \u_a23_mem/n19743 , \u_a23_mem/n19742 , \u_a23_mem/n19741 ,
         \u_a23_mem/n19740 , \u_a23_mem/n19739 , \u_a23_mem/n19738 ,
         \u_a23_mem/n19737 , \u_a23_mem/n19736 , \u_a23_mem/n19735 ,
         \u_a23_mem/n19734 , \u_a23_mem/n19733 , \u_a23_mem/n19732 ,
         \u_a23_mem/n19731 , \u_a23_mem/n19730 , \u_a23_mem/n19729 ,
         \u_a23_mem/n19728 , \u_a23_mem/n19727 , \u_a23_mem/n19726 ,
         \u_a23_mem/n19725 , \u_a23_mem/n19724 , \u_a23_mem/n19723 ,
         \u_a23_mem/n19722 , \u_a23_mem/n19721 , \u_a23_mem/n19720 ,
         \u_a23_mem/n19719 , \u_a23_mem/n19718 , \u_a23_mem/n19717 ,
         \u_a23_mem/n19716 , \u_a23_mem/n19715 , \u_a23_mem/n19713 ,
         \u_a23_mem/n19712 , \u_a23_mem/n19711 , \u_a23_mem/n19710 ,
         \u_a23_mem/n19709 , \u_a23_mem/n19708 , \u_a23_mem/n19707 ,
         \u_a23_mem/n19706 , \u_a23_mem/n19705 , \u_a23_mem/n19704 ,
         \u_a23_mem/n19703 , \u_a23_mem/n19702 , \u_a23_mem/n19701 ,
         \u_a23_mem/n19700 , \u_a23_mem/n19699 , \u_a23_mem/n19698 ,
         \u_a23_mem/n19697 , \u_a23_mem/n19696 , \u_a23_mem/n19695 ,
         \u_a23_mem/n19694 , \u_a23_mem/n19693 , \u_a23_mem/n19692 ,
         \u_a23_mem/n19691 , \u_a23_mem/n19690 , \u_a23_mem/n19689 ,
         \u_a23_mem/n19688 , \u_a23_mem/n19687 , \u_a23_mem/n19686 ,
         \u_a23_mem/n19685 , \u_a23_mem/n19684 , \u_a23_mem/n19683 ,
         \u_a23_mem/n19652 , \u_a23_mem/n19651 , \u_a23_mem/n19650 ,
         \u_a23_mem/n19649 , \u_a23_mem/n19648 , \u_a23_mem/n19647 ,
         \u_a23_mem/n19646 , \u_a23_mem/n19645 , \u_a23_mem/n19644 ,
         \u_a23_mem/n19643 , \u_a23_mem/n19642 , \u_a23_mem/n19641 ,
         \u_a23_mem/n19640 , \u_a23_mem/n19639 , \u_a23_mem/n19638 ,
         \u_a23_mem/n19637 , \u_a23_mem/n19636 , \u_a23_mem/n19635 ,
         \u_a23_mem/n19634 , \u_a23_mem/n19633 , \u_a23_mem/n19632 ,
         \u_a23_mem/n19631 , \u_a23_mem/n19630 , \u_a23_mem/n19629 ,
         \u_a23_mem/n19628 , \u_a23_mem/n19627 , \u_a23_mem/n19626 ,
         \u_a23_mem/n19625 , \u_a23_mem/n19624 , \u_a23_mem/n19623 ,
         \u_a23_mem/n19622 , \u_a23_mem/n19621 , \u_a23_mem/n19620 ,
         \u_a23_mem/n19619 , \u_a23_mem/n19618 , \u_a23_mem/n19617 ,
         \u_a23_mem/n19616 , \u_a23_mem/n19615 , \u_a23_mem/n19614 ,
         \u_a23_mem/n19613 , \u_a23_mem/n19612 , \u_a23_mem/n19611 ,
         \u_a23_mem/n19610 , \u_a23_mem/n19609 , \u_a23_mem/n19608 ,
         \u_a23_mem/n19607 , \u_a23_mem/n19606 , \u_a23_mem/n19605 ,
         \u_a23_mem/n19604 , \u_a23_mem/n19603 , \u_a23_mem/n19602 ,
         \u_a23_mem/n19601 , \u_a23_mem/n19600 , \u_a23_mem/n19599 ,
         \u_a23_mem/n19598 , \u_a23_mem/n19597 , \u_a23_mem/n19596 ,
         \u_a23_mem/n19595 , \u_a23_mem/n19594 , \u_a23_mem/n19593 ,
         \u_a23_mem/n19592 , \u_a23_mem/n19591 , \u_a23_mem/n19590 ,
         \u_a23_mem/n19589 , \u_a23_mem/n19588 , \u_a23_mem/n19587 ,
         \u_a23_mem/n19586 , \u_a23_mem/n19585 , \u_a23_mem/n19584 ,
         \u_a23_mem/n19583 , \u_a23_mem/n19582 , \u_a23_mem/n19581 ,
         \u_a23_mem/n19580 , \u_a23_mem/n19579 , \u_a23_mem/n19578 ,
         \u_a23_mem/n19577 , \u_a23_mem/n19576 , \u_a23_mem/n19575 ,
         \u_a23_mem/n19574 , \u_a23_mem/n19573 , \u_a23_mem/n19572 ,
         \u_a23_mem/n19571 , \u_a23_mem/n19570 , \u_a23_mem/n19569 ,
         \u_a23_mem/n19568 , \u_a23_mem/n19567 , \u_a23_mem/n19566 ,
         \u_a23_mem/n19565 , \u_a23_mem/n19564 , \u_a23_mem/n19563 ,
         \u_a23_mem/n19562 , \u_a23_mem/n19561 , \u_a23_mem/n19560 ,
         \u_a23_mem/n19559 , \u_a23_mem/n19558 , \u_a23_mem/n19557 ,
         \u_a23_mem/n19556 , \u_a23_mem/n19555 , \u_a23_mem/n19554 ,
         \u_a23_mem/n19553 , \u_a23_mem/n19552 , \u_a23_mem/n19551 ,
         \u_a23_mem/n19550 , \u_a23_mem/n19549 , \u_a23_mem/n19548 ,
         \u_a23_mem/n19547 , \u_a23_mem/n19546 , \u_a23_mem/n19545 ,
         \u_a23_mem/n19544 , \u_a23_mem/n19543 , \u_a23_mem/n19542 ,
         \u_a23_mem/n19541 , \u_a23_mem/n19540 , \u_a23_mem/n19539 ,
         \u_a23_mem/n19538 , \u_a23_mem/n19537 , \u_a23_mem/n19536 ,
         \u_a23_mem/n19535 , \u_a23_mem/n19534 , \u_a23_mem/n19533 ,
         \u_a23_mem/n19532 , \u_a23_mem/n19531 , \u_a23_mem/n19530 ,
         \u_a23_mem/n19529 , \u_a23_mem/n19528 , \u_a23_mem/n19527 ,
         \u_a23_mem/n19526 , \u_a23_mem/n19525 , \u_a23_mem/n19524 ,
         \u_a23_mem/n19523 , \u_a23_mem/n19522 , \u_a23_mem/n19521 ,
         \u_a23_mem/n19520 , \u_a23_mem/n19519 , \u_a23_mem/n19518 ,
         \u_a23_mem/n19517 , \u_a23_mem/n19516 , \u_a23_mem/n19515 ,
         \u_a23_mem/n19514 , \u_a23_mem/n19513 , \u_a23_mem/n19512 ,
         \u_a23_mem/n19511 , \u_a23_mem/n19510 , \u_a23_mem/n19509 ,
         \u_a23_mem/n19508 , \u_a23_mem/n19507 , \u_a23_mem/n19506 ,
         \u_a23_mem/n19505 , \u_a23_mem/n19504 , \u_a23_mem/n19503 ,
         \u_a23_mem/n19502 , \u_a23_mem/n19501 , \u_a23_mem/n19500 ,
         \u_a23_mem/n19499 , \u_a23_mem/n19498 , \u_a23_mem/n19497 ,
         \u_a23_mem/n19496 , \u_a23_mem/n19495 , \u_a23_mem/n19494 ,
         \u_a23_mem/n19493 , \u_a23_mem/n19492 , \u_a23_mem/n19491 ,
         \u_a23_mem/n19490 , \u_a23_mem/n19489 , \u_a23_mem/n19488 ,
         \u_a23_mem/n19487 , \u_a23_mem/n19486 , \u_a23_mem/n19485 ,
         \u_a23_mem/n19484 , \u_a23_mem/n19483 , \u_a23_mem/n19482 ,
         \u_a23_mem/n19481 , \u_a23_mem/n19480 , \u_a23_mem/n19479 ,
         \u_a23_mem/n19478 , \u_a23_mem/n19477 , \u_a23_mem/n19476 ,
         \u_a23_mem/n19475 , \u_a23_mem/n19474 , \u_a23_mem/n19473 ,
         \u_a23_mem/n19472 , \u_a23_mem/n19471 , \u_a23_mem/n19470 ,
         \u_a23_mem/n19469 , \u_a23_mem/n19468 , \u_a23_mem/n19467 ,
         \u_a23_mem/n19466 , \u_a23_mem/n19465 , \u_a23_mem/n19464 ,
         \u_a23_mem/n19463 , \u_a23_mem/n19462 , \u_a23_mem/n19461 ,
         \u_a23_mem/n19460 , \u_a23_mem/n19459 , \u_a23_mem/n19458 ,
         \u_a23_mem/n19457 , \u_a23_mem/n19456 , \u_a23_mem/n19455 ,
         \u_a23_mem/n19454 , \u_a23_mem/n19453 , \u_a23_mem/n19452 ,
         \u_a23_mem/n19451 , \u_a23_mem/n19450 , \u_a23_mem/n19449 ,
         \u_a23_mem/n19448 , \u_a23_mem/n19447 , \u_a23_mem/n19446 ,
         \u_a23_mem/n19445 , \u_a23_mem/n19444 , \u_a23_mem/n19443 ,
         \u_a23_mem/n19442 , \u_a23_mem/n19441 , \u_a23_mem/n19440 ,
         \u_a23_mem/n19439 , \u_a23_mem/n19438 , \u_a23_mem/n19437 ,
         \u_a23_mem/n19436 , \u_a23_mem/n19435 , \u_a23_mem/n19434 ,
         \u_a23_mem/n19433 , \u_a23_mem/n19432 , \u_a23_mem/n19431 ,
         \u_a23_mem/n19430 , \u_a23_mem/n19429 , \u_a23_mem/n19428 ,
         \u_a23_mem/n19427 , \u_a23_mem/n19426 , \u_a23_mem/n19425 ,
         \u_a23_mem/n19424 , \u_a23_mem/n19423 , \u_a23_mem/n19422 ,
         \u_a23_mem/n19421 , \u_a23_mem/n19420 , \u_a23_mem/n19419 ,
         \u_a23_mem/n19418 , \u_a23_mem/n19417 , \u_a23_mem/n19416 ,
         \u_a23_mem/n19415 , \u_a23_mem/n19414 , \u_a23_mem/n19413 ,
         \u_a23_mem/n19412 , \u_a23_mem/n19411 , \u_a23_mem/n19410 ,
         \u_a23_mem/n19409 , \u_a23_mem/n19408 , \u_a23_mem/n19407 ,
         \u_a23_mem/n19406 , \u_a23_mem/n19405 , \u_a23_mem/n19404 ,
         \u_a23_mem/n19403 , \u_a23_mem/n19402 , \u_a23_mem/n19401 ,
         \u_a23_mem/n19400 , \u_a23_mem/n19399 , \u_a23_mem/n19398 ,
         \u_a23_mem/n19397 , \u_a23_mem/n19396 , \u_a23_mem/n19395 ,
         \u_a23_mem/n19394 , \u_a23_mem/n19393 , \u_a23_mem/n19392 ,
         \u_a23_mem/n19391 , \u_a23_mem/n19390 , \u_a23_mem/n19389 ,
         \u_a23_mem/n19388 , \u_a23_mem/n19387 , \u_a23_mem/n19386 ,
         \u_a23_mem/n19385 , \u_a23_mem/n19384 , \u_a23_mem/n19383 ,
         \u_a23_mem/n19382 , \u_a23_mem/n19381 , \u_a23_mem/n19380 ,
         \u_a23_mem/n19379 , \u_a23_mem/n19378 , \u_a23_mem/n19377 ,
         \u_a23_mem/n19376 , \u_a23_mem/n19375 , \u_a23_mem/n19374 ,
         \u_a23_mem/n19373 , \u_a23_mem/n19372 , \u_a23_mem/n19371 ,
         \u_a23_mem/n19370 , \u_a23_mem/n19369 , \u_a23_mem/n19368 ,
         \u_a23_mem/n19367 , \u_a23_mem/n19366 , \u_a23_mem/n19365 ,
         \u_a23_mem/n19364 , \u_a23_mem/n19363 , \u_a23_mem/n19362 ,
         \u_a23_mem/n19361 , \u_a23_mem/n19360 , \u_a23_mem/n19359 ,
         \u_a23_mem/n19358 , \u_a23_mem/n19357 , \u_a23_mem/n19356 ,
         \u_a23_mem/n19355 , \u_a23_mem/n19354 , \u_a23_mem/n19353 ,
         \u_a23_mem/n19352 , \u_a23_mem/n19351 , \u_a23_mem/n19350 ,
         \u_a23_mem/n19349 , \u_a23_mem/n19348 , \u_a23_mem/n19347 ,
         \u_a23_mem/n19346 , \u_a23_mem/n19345 , \u_a23_mem/n19344 ,
         \u_a23_mem/n19343 , \u_a23_mem/n19342 , \u_a23_mem/n19341 ,
         \u_a23_mem/n19340 , \u_a23_mem/n19339 , \u_a23_mem/n19338 ,
         \u_a23_mem/n19337 , \u_a23_mem/n19336 , \u_a23_mem/n19335 ,
         \u_a23_mem/n19334 , \u_a23_mem/n19333 , \u_a23_mem/n19332 ,
         \u_a23_mem/n19331 , \u_a23_mem/n19330 , \u_a23_mem/n19329 ,
         \u_a23_mem/n19328 , \u_a23_mem/n19327 , \u_a23_mem/n19326 ,
         \u_a23_mem/n19325 , \u_a23_mem/n19324 , \u_a23_mem/n19323 ,
         \u_a23_mem/n19322 , \u_a23_mem/n19321 , \u_a23_mem/n19320 ,
         \u_a23_mem/n19319 , \u_a23_mem/n19318 , \u_a23_mem/n19317 ,
         \u_a23_mem/n19316 , \u_a23_mem/n19315 , \u_a23_mem/n19314 ,
         \u_a23_mem/n19313 , \u_a23_mem/n19312 , \u_a23_mem/n19311 ,
         \u_a23_mem/n19310 , \u_a23_mem/n19309 , \u_a23_mem/n19308 ,
         \u_a23_mem/n19307 , \u_a23_mem/n19306 , \u_a23_mem/n19305 ,
         \u_a23_mem/n19304 , \u_a23_mem/n19303 , \u_a23_mem/n19302 ,
         \u_a23_mem/n19301 , \u_a23_mem/n19300 , \u_a23_mem/n19299 ,
         \u_a23_mem/n19298 , \u_a23_mem/n19297 , \u_a23_mem/n19296 ,
         \u_a23_mem/n19295 , \u_a23_mem/n19294 , \u_a23_mem/n19293 ,
         \u_a23_mem/n19292 , \u_a23_mem/n19291 , \u_a23_mem/n19290 ,
         \u_a23_mem/n19289 , \u_a23_mem/n19288 , \u_a23_mem/n19287 ,
         \u_a23_mem/n19286 , \u_a23_mem/n19285 , \u_a23_mem/n19284 ,
         \u_a23_mem/n19283 , \u_a23_mem/n19282 , \u_a23_mem/n19281 ,
         \u_a23_mem/n19280 , \u_a23_mem/n19279 , \u_a23_mem/n19278 ,
         \u_a23_mem/n19277 , \u_a23_mem/n19276 , \u_a23_mem/n19275 ,
         \u_a23_mem/n19274 , \u_a23_mem/n19273 , \u_a23_mem/n19272 ,
         \u_a23_mem/n19271 , \u_a23_mem/n19270 , \u_a23_mem/n19269 ,
         \u_a23_mem/n19268 , \u_a23_mem/n19267 , \u_a23_mem/n19266 ,
         \u_a23_mem/n19265 , \u_a23_mem/n19264 , \u_a23_mem/n19263 ,
         \u_a23_mem/n19262 , \u_a23_mem/n19261 , \u_a23_mem/n19260 ,
         \u_a23_mem/n19259 , \u_a23_mem/n19258 , \u_a23_mem/n19257 ,
         \u_a23_mem/n19256 , \u_a23_mem/n19255 , \u_a23_mem/n19254 ,
         \u_a23_mem/n19253 , \u_a23_mem/n19252 , \u_a23_mem/n19251 ,
         \u_a23_mem/n19250 , \u_a23_mem/n19249 , \u_a23_mem/n19248 ,
         \u_a23_mem/n19247 , \u_a23_mem/n19246 , \u_a23_mem/n19245 ,
         \u_a23_mem/n19244 , \u_a23_mem/n19243 , \u_a23_mem/n19242 ,
         \u_a23_mem/n19241 , \u_a23_mem/n19240 , \u_a23_mem/n19239 ,
         \u_a23_mem/n19238 , \u_a23_mem/n19237 , \u_a23_mem/n19236 ,
         \u_a23_mem/n19235 , \u_a23_mem/n19234 , \u_a23_mem/n19233 ,
         \u_a23_mem/n19232 , \u_a23_mem/n19231 , \u_a23_mem/n19230 ,
         \u_a23_mem/n19229 , \u_a23_mem/n19228 , \u_a23_mem/n19227 ,
         \u_a23_mem/n19226 , \u_a23_mem/n19225 , \u_a23_mem/n19224 ,
         \u_a23_mem/n19223 , \u_a23_mem/n19222 , \u_a23_mem/n19221 ,
         \u_a23_mem/n19220 , \u_a23_mem/n19219 , \u_a23_mem/n19218 ,
         \u_a23_mem/n19217 , \u_a23_mem/n19216 , \u_a23_mem/n19215 ,
         \u_a23_mem/n19214 , \u_a23_mem/n19213 , \u_a23_mem/n19212 ,
         \u_a23_mem/n19211 , \u_a23_mem/n19210 , \u_a23_mem/n19209 ,
         \u_a23_mem/n19208 , \u_a23_mem/n19207 , \u_a23_mem/n19206 ,
         \u_a23_mem/n19205 , \u_a23_mem/n19204 , \u_a23_mem/n19203 ,
         \u_a23_mem/n19202 , \u_a23_mem/n19201 , \u_a23_mem/n19200 ,
         \u_a23_mem/n19199 , \u_a23_mem/n19198 , \u_a23_mem/n19197 ,
         \u_a23_mem/n19196 , \u_a23_mem/n19195 , \u_a23_mem/n19194 ,
         \u_a23_mem/n19193 , \u_a23_mem/n19192 , \u_a23_mem/n19191 ,
         \u_a23_mem/n19190 , \u_a23_mem/n19189 , \u_a23_mem/n19188 ,
         \u_a23_mem/n19187 , \u_a23_mem/n19186 , \u_a23_mem/n19185 ,
         \u_a23_mem/n19184 , \u_a23_mem/n19183 , \u_a23_mem/n19182 ,
         \u_a23_mem/n19181 , \u_a23_mem/n19180 , \u_a23_mem/n19179 ,
         \u_a23_mem/n19178 , \u_a23_mem/n19177 , \u_a23_mem/n19176 ,
         \u_a23_mem/n19175 , \u_a23_mem/n19174 , \u_a23_mem/n19173 ,
         \u_a23_mem/n19172 , \u_a23_mem/n19171 , \u_a23_mem/n19170 ,
         \u_a23_mem/n19169 , \u_a23_mem/n19168 , \u_a23_mem/n19167 ,
         \u_a23_mem/n19166 , \u_a23_mem/n19165 , \u_a23_mem/n19164 ,
         \u_a23_mem/n19163 , \u_a23_mem/n19162 , \u_a23_mem/n19161 ,
         \u_a23_mem/n19160 , \u_a23_mem/n19159 , \u_a23_mem/n19158 ,
         \u_a23_mem/n19157 , \u_a23_mem/n19156 , \u_a23_mem/n19155 ,
         \u_a23_mem/n19154 , \u_a23_mem/n19153 , \u_a23_mem/n19152 ,
         \u_a23_mem/n19151 , \u_a23_mem/n19150 , \u_a23_mem/n19149 ,
         \u_a23_mem/n19148 , \u_a23_mem/n19147 , \u_a23_mem/n19146 ,
         \u_a23_mem/n19145 , \u_a23_mem/n19144 , \u_a23_mem/n19143 ,
         \u_a23_mem/n19142 , \u_a23_mem/n19141 , \u_a23_mem/n19140 ,
         \u_a23_mem/n19139 , \u_a23_mem/n19138 , \u_a23_mem/n19137 ,
         \u_a23_mem/n19136 , \u_a23_mem/n19135 , \u_a23_mem/n19134 ,
         \u_a23_mem/n19133 , \u_a23_mem/n19132 , \u_a23_mem/n19131 ,
         \u_a23_mem/n19130 , \u_a23_mem/n19129 , \u_a23_mem/n19128 ,
         \u_a23_mem/n19127 , \u_a23_mem/n19126 , \u_a23_mem/n19125 ,
         \u_a23_mem/n19124 , \u_a23_mem/n19123 , \u_a23_mem/n19122 ,
         \u_a23_mem/n19121 , \u_a23_mem/n19120 , \u_a23_mem/n19119 ,
         \u_a23_mem/n19118 , \u_a23_mem/n19117 , \u_a23_mem/n19116 ,
         \u_a23_mem/n19115 , \u_a23_mem/n19114 , \u_a23_mem/n19113 ,
         \u_a23_mem/n19112 , \u_a23_mem/n19111 , \u_a23_mem/n19110 ,
         \u_a23_mem/n19109 , \u_a23_mem/n19108 , \u_a23_mem/n19107 ,
         \u_a23_mem/n19106 , \u_a23_mem/n19105 , \u_a23_mem/n19104 ,
         \u_a23_mem/n19103 , \u_a23_mem/n19102 , \u_a23_mem/n19101 ,
         \u_a23_mem/n19100 , \u_a23_mem/n19099 , \u_a23_mem/n19098 ,
         \u_a23_mem/n19097 , \u_a23_mem/n19096 , \u_a23_mem/n19095 ,
         \u_a23_mem/n19094 , \u_a23_mem/n19093 , \u_a23_mem/n19092 ,
         \u_a23_mem/n19091 , \u_a23_mem/n19090 , \u_a23_mem/n19089 ,
         \u_a23_mem/n19088 , \u_a23_mem/n19087 , \u_a23_mem/n19086 ,
         \u_a23_mem/n19085 , \u_a23_mem/n19084 , \u_a23_mem/n19083 ,
         \u_a23_mem/n19082 , \u_a23_mem/n19081 , \u_a23_mem/n19080 ,
         \u_a23_mem/n19079 , \u_a23_mem/n19078 , \u_a23_mem/n19077 ,
         \u_a23_mem/n19076 , \u_a23_mem/n19075 , \u_a23_mem/n19074 ,
         \u_a23_mem/n19073 , \u_a23_mem/n19072 , \u_a23_mem/n19071 ,
         \u_a23_mem/n19070 , \u_a23_mem/n19069 , \u_a23_mem/n19068 ,
         \u_a23_mem/n19067 , \u_a23_mem/n19066 , \u_a23_mem/n19065 ,
         \u_a23_mem/n19064 , \u_a23_mem/n19063 , \u_a23_mem/n19062 ,
         \u_a23_mem/n19061 , \u_a23_mem/n19060 , \u_a23_mem/n19059 ,
         \u_a23_mem/n19058 , \u_a23_mem/n19057 , \u_a23_mem/n19056 ,
         \u_a23_mem/n19055 , \u_a23_mem/n19054 , \u_a23_mem/n19053 ,
         \u_a23_mem/n19052 , \u_a23_mem/n19051 , \u_a23_mem/n19050 ,
         \u_a23_mem/n19049 , \u_a23_mem/n19048 , \u_a23_mem/n19047 ,
         \u_a23_mem/n19046 , \u_a23_mem/n19045 , \u_a23_mem/n19044 ,
         \u_a23_mem/n19043 , \u_a23_mem/n19042 , \u_a23_mem/n19041 ,
         \u_a23_mem/n19040 , \u_a23_mem/n19039 , \u_a23_mem/n19038 ,
         \u_a23_mem/n19037 , \u_a23_mem/n19036 , \u_a23_mem/n19035 ,
         \u_a23_mem/n19034 , \u_a23_mem/n19033 , \u_a23_mem/n19032 ,
         \u_a23_mem/n19031 , \u_a23_mem/n19030 , \u_a23_mem/n19029 ,
         \u_a23_mem/n19028 , \u_a23_mem/n19027 , \u_a23_mem/n19026 ,
         \u_a23_mem/n19025 , \u_a23_mem/n19024 , \u_a23_mem/n19023 ,
         \u_a23_mem/n19022 , \u_a23_mem/n19021 , \u_a23_mem/n19020 ,
         \u_a23_mem/n19019 , \u_a23_mem/n19018 , \u_a23_mem/n19017 ,
         \u_a23_mem/n19016 , \u_a23_mem/n19015 , \u_a23_mem/n19014 ,
         \u_a23_mem/n19013 , \u_a23_mem/n19012 , \u_a23_mem/n19011 ,
         \u_a23_mem/n19010 , \u_a23_mem/n19009 , \u_a23_mem/n19008 ,
         \u_a23_mem/n19007 , \u_a23_mem/n19006 , \u_a23_mem/n19005 ,
         \u_a23_mem/n19004 , \u_a23_mem/n19003 , \u_a23_mem/n19002 ,
         \u_a23_mem/n19001 , \u_a23_mem/n19000 , \u_a23_mem/n18999 ,
         \u_a23_mem/n18998 , \u_a23_mem/n18997 , \u_a23_mem/n18996 ,
         \u_a23_mem/n18995 , \u_a23_mem/n18994 , \u_a23_mem/n18993 ,
         \u_a23_mem/n18992 , \u_a23_mem/n18991 , \u_a23_mem/n18990 ,
         \u_a23_mem/n18989 , \u_a23_mem/n18988 , \u_a23_mem/n18987 ,
         \u_a23_mem/n18986 , \u_a23_mem/n18985 , \u_a23_mem/n18984 ,
         \u_a23_mem/n18983 , \u_a23_mem/n18982 , \u_a23_mem/n18981 ,
         \u_a23_mem/n18980 , \u_a23_mem/n18979 , \u_a23_mem/n18978 ,
         \u_a23_mem/n18977 , \u_a23_mem/n18976 , \u_a23_mem/n18975 ,
         \u_a23_mem/n18974 , \u_a23_mem/n18973 , \u_a23_mem/n18972 ,
         \u_a23_mem/n18971 , \u_a23_mem/n18970 , \u_a23_mem/n18969 ,
         \u_a23_mem/n18968 , \u_a23_mem/n18967 , \u_a23_mem/n18966 ,
         \u_a23_mem/n18965 , \u_a23_mem/n18964 , \u_a23_mem/n18963 ,
         \u_a23_mem/n18962 , \u_a23_mem/n18961 , \u_a23_mem/n18960 ,
         \u_a23_mem/n18959 , \u_a23_mem/n18958 , \u_a23_mem/n18957 ,
         \u_a23_mem/n18956 , \u_a23_mem/n18955 , \u_a23_mem/n18954 ,
         \u_a23_mem/n18953 , \u_a23_mem/n18952 , \u_a23_mem/n18951 ,
         \u_a23_mem/n18950 , \u_a23_mem/n18949 , \u_a23_mem/n18948 ,
         \u_a23_mem/n18947 , \u_a23_mem/n18946 , \u_a23_mem/n18945 ,
         \u_a23_mem/n18944 , \u_a23_mem/n18943 , \u_a23_mem/n18942 ,
         \u_a23_mem/n18941 , \u_a23_mem/n18940 , \u_a23_mem/n18939 ,
         \u_a23_mem/n18938 , \u_a23_mem/n18937 , \u_a23_mem/n18936 ,
         \u_a23_mem/n18935 , \u_a23_mem/n18934 , \u_a23_mem/n18933 ,
         \u_a23_mem/n18932 , \u_a23_mem/n18931 , \u_a23_mem/n18930 ,
         \u_a23_mem/n18929 , \u_a23_mem/n18928 , \u_a23_mem/n18927 ,
         \u_a23_mem/n18926 , \u_a23_mem/n18925 , \u_a23_mem/n18924 ,
         \u_a23_mem/n18923 , \u_a23_mem/n18922 , \u_a23_mem/n18921 ,
         \u_a23_mem/n18920 , \u_a23_mem/n18919 , \u_a23_mem/n18918 ,
         \u_a23_mem/n18917 , \u_a23_mem/n18916 , \u_a23_mem/n18915 ,
         \u_a23_mem/n18914 , \u_a23_mem/n18913 , \u_a23_mem/n18912 ,
         \u_a23_mem/n18911 , \u_a23_mem/n18910 , \u_a23_mem/n18909 ,
         \u_a23_mem/n18908 , \u_a23_mem/n18907 , \u_a23_mem/n18906 ,
         \u_a23_mem/n18905 , \u_a23_mem/n18904 , \u_a23_mem/n18903 ,
         \u_a23_mem/n18902 , \u_a23_mem/n18901 , \u_a23_mem/n18900 ,
         \u_a23_mem/n18899 , \u_a23_mem/n18898 , \u_a23_mem/n18897 ,
         \u_a23_mem/n18896 , \u_a23_mem/n18895 , \u_a23_mem/n18894 ,
         \u_a23_mem/n18893 , \u_a23_mem/n18892 , \u_a23_mem/n18891 ,
         \u_a23_mem/n18890 , \u_a23_mem/n18889 , \u_a23_mem/n18888 ,
         \u_a23_mem/n18887 , \u_a23_mem/n18886 , \u_a23_mem/n18885 ,
         \u_a23_mem/n18884 , \u_a23_mem/n18883 , \u_a23_mem/n18882 ,
         \u_a23_mem/n18881 , \u_a23_mem/n18880 , \u_a23_mem/n18879 ,
         \u_a23_mem/n18878 , \u_a23_mem/n18877 , \u_a23_mem/n18876 ,
         \u_a23_mem/n18875 , \u_a23_mem/n18874 , \u_a23_mem/n18873 ,
         \u_a23_mem/n18872 , \u_a23_mem/n18871 , \u_a23_mem/n18870 ,
         \u_a23_mem/n18869 , \u_a23_mem/n18868 , \u_a23_mem/n18867 ,
         \u_a23_mem/n18866 , \u_a23_mem/n18865 , \u_a23_mem/n18864 ,
         \u_a23_mem/n18863 , \u_a23_mem/n18862 , \u_a23_mem/n18861 ,
         \u_a23_mem/n18860 , \u_a23_mem/n18859 , \u_a23_mem/n18858 ,
         \u_a23_mem/n18857 , \u_a23_mem/n18856 , \u_a23_mem/n18855 ,
         \u_a23_mem/n18854 , \u_a23_mem/n18853 , \u_a23_mem/n18852 ,
         \u_a23_mem/n18851 , \u_a23_mem/n18850 , \u_a23_mem/n18849 ,
         \u_a23_mem/n18848 , \u_a23_mem/n18847 , \u_a23_mem/n18846 ,
         \u_a23_mem/n18845 , \u_a23_mem/n18844 , \u_a23_mem/n18843 ,
         \u_a23_mem/n18842 , \u_a23_mem/n18841 , \u_a23_mem/n18840 ,
         \u_a23_mem/n18839 , \u_a23_mem/n18838 , \u_a23_mem/n18837 ,
         \u_a23_mem/n18836 , \u_a23_mem/n18835 , \u_a23_mem/n18834 ,
         \u_a23_mem/n18833 , \u_a23_mem/n18832 , \u_a23_mem/n18831 ,
         \u_a23_mem/n18830 , \u_a23_mem/n18829 , \u_a23_mem/n18828 ,
         \u_a23_mem/n18827 , \u_a23_mem/n18826 , \u_a23_mem/n18825 ,
         \u_a23_mem/n18824 , \u_a23_mem/n18823 , \u_a23_mem/n18822 ,
         \u_a23_mem/n18821 , \u_a23_mem/n18820 , \u_a23_mem/n18819 ,
         \u_a23_mem/n18818 , \u_a23_mem/n18817 , \u_a23_mem/n18816 ,
         \u_a23_mem/n18815 , \u_a23_mem/n18814 , \u_a23_mem/n18813 ,
         \u_a23_mem/n18812 , \u_a23_mem/n18811 , \u_a23_mem/n18810 ,
         \u_a23_mem/n18809 , \u_a23_mem/n18808 , \u_a23_mem/n18807 ,
         \u_a23_mem/n18806 , \u_a23_mem/n18805 , \u_a23_mem/n18804 ,
         \u_a23_mem/n18803 , \u_a23_mem/n18802 , \u_a23_mem/n18801 ,
         \u_a23_mem/n18800 , \u_a23_mem/n18799 , \u_a23_mem/n18798 ,
         \u_a23_mem/n18797 , \u_a23_mem/n18796 , \u_a23_mem/n18795 ,
         \u_a23_mem/n18794 , \u_a23_mem/n18793 , \u_a23_mem/n18792 ,
         \u_a23_mem/n18791 , \u_a23_mem/n18790 , \u_a23_mem/n18789 ,
         \u_a23_mem/n18788 , \u_a23_mem/n18787 , \u_a23_mem/n18786 ,
         \u_a23_mem/n18785 , \u_a23_mem/n18784 , \u_a23_mem/n18783 ,
         \u_a23_mem/n18782 , \u_a23_mem/n18781 , \u_a23_mem/n18780 ,
         \u_a23_mem/n18779 , \u_a23_mem/n18778 , \u_a23_mem/n18777 ,
         \u_a23_mem/n18776 , \u_a23_mem/n18775 , \u_a23_mem/n18774 ,
         \u_a23_mem/n18773 , \u_a23_mem/n18772 , \u_a23_mem/n18771 ,
         \u_a23_mem/n18770 , \u_a23_mem/n18769 , \u_a23_mem/n18768 ,
         \u_a23_mem/n18767 , \u_a23_mem/n18766 , \u_a23_mem/n18765 ,
         \u_a23_mem/n18764 , \u_a23_mem/n18763 , \u_a23_mem/n18762 ,
         \u_a23_mem/n18761 , \u_a23_mem/n18760 , \u_a23_mem/n18759 ,
         \u_a23_mem/n18758 , \u_a23_mem/n18757 , \u_a23_mem/n18756 ,
         \u_a23_mem/n18755 , \u_a23_mem/n18754 , \u_a23_mem/n18753 ,
         \u_a23_mem/n18752 , \u_a23_mem/n18751 , \u_a23_mem/n18750 ,
         \u_a23_mem/n18749 , \u_a23_mem/n18748 , \u_a23_mem/n18747 ,
         \u_a23_mem/n18746 , \u_a23_mem/n18745 , \u_a23_mem/n18744 ,
         \u_a23_mem/n18743 , \u_a23_mem/n18742 , \u_a23_mem/n18741 ,
         \u_a23_mem/n18740 , \u_a23_mem/n18739 , \u_a23_mem/n18738 ,
         \u_a23_mem/n18737 , \u_a23_mem/n18736 , \u_a23_mem/n18735 ,
         \u_a23_mem/n18734 , \u_a23_mem/n18733 , \u_a23_mem/n18732 ,
         \u_a23_mem/n18731 , \u_a23_mem/n18730 , \u_a23_mem/n18729 ,
         \u_a23_mem/n18728 , \u_a23_mem/n18727 , \u_a23_mem/n18726 ,
         \u_a23_mem/n18725 , \u_a23_mem/n18724 , \u_a23_mem/n18723 ,
         \u_a23_mem/n18722 , \u_a23_mem/n18721 , \u_a23_mem/n18720 ,
         \u_a23_mem/n18719 , \u_a23_mem/n18718 , \u_a23_mem/n18717 ,
         \u_a23_mem/n18716 , \u_a23_mem/n18715 , \u_a23_mem/n18714 ,
         \u_a23_mem/n18713 , \u_a23_mem/n18712 , \u_a23_mem/n18711 ,
         \u_a23_mem/n18710 , \u_a23_mem/n18709 , \u_a23_mem/n18708 ,
         \u_a23_mem/n18707 , \u_a23_mem/n18706 , \u_a23_mem/n18705 ,
         \u_a23_mem/n18704 , \u_a23_mem/n18703 , \u_a23_mem/n18702 ,
         \u_a23_mem/n18701 , \u_a23_mem/n18700 , \u_a23_mem/n18699 ,
         \u_a23_mem/n18698 , \u_a23_mem/n18697 , \u_a23_mem/n18696 ,
         \u_a23_mem/n18695 , \u_a23_mem/n18694 , \u_a23_mem/n18693 ,
         \u_a23_mem/n18692 , \u_a23_mem/n18691 , \u_a23_mem/n18690 ,
         \u_a23_mem/n18689 , \u_a23_mem/n18688 , \u_a23_mem/n18687 ,
         \u_a23_mem/n18686 , \u_a23_mem/n18685 , \u_a23_mem/n18684 ,
         \u_a23_mem/n18683 , \u_a23_mem/n18682 , \u_a23_mem/n18681 ,
         \u_a23_mem/n18680 , \u_a23_mem/n18679 , \u_a23_mem/n18678 ,
         \u_a23_mem/n18677 , \u_a23_mem/n18676 , \u_a23_mem/n18675 ,
         \u_a23_mem/n18674 , \u_a23_mem/n18673 , \u_a23_mem/n18672 ,
         \u_a23_mem/n18671 , \u_a23_mem/n18670 , \u_a23_mem/n18669 ,
         \u_a23_mem/n18668 , \u_a23_mem/n18667 , \u_a23_mem/n18666 ,
         \u_a23_mem/n18665 , \u_a23_mem/n18664 , \u_a23_mem/n18663 ,
         \u_a23_mem/n18662 , \u_a23_mem/n18661 , \u_a23_mem/n18660 ,
         \u_a23_mem/n18659 , \u_a23_mem/n18658 , \u_a23_mem/n18657 ,
         \u_a23_mem/n18656 , \u_a23_mem/n18655 , \u_a23_mem/n18654 ,
         \u_a23_mem/n18653 , \u_a23_mem/n18652 , \u_a23_mem/n18651 ,
         \u_a23_mem/n18650 , \u_a23_mem/n18649 , \u_a23_mem/n18648 ,
         \u_a23_mem/n18647 , \u_a23_mem/n18646 , \u_a23_mem/n18645 ,
         \u_a23_mem/n18644 , \u_a23_mem/n18643 , \u_a23_mem/n18642 ,
         \u_a23_mem/n18641 , \u_a23_mem/n18640 , \u_a23_mem/n18639 ,
         \u_a23_mem/n18638 , \u_a23_mem/n18637 , \u_a23_mem/n18636 ,
         \u_a23_mem/n18635 , \u_a23_mem/n18634 , \u_a23_mem/n18633 ,
         \u_a23_mem/n18632 , \u_a23_mem/n18631 , \u_a23_mem/n18630 ,
         \u_a23_mem/n18629 , \u_a23_mem/n18628 , \u_a23_mem/n18627 ,
         \u_a23_mem/n18626 , \u_a23_mem/n18625 , \u_a23_mem/n18624 ,
         \u_a23_mem/n18623 , \u_a23_mem/n18622 , \u_a23_mem/n18621 ,
         \u_a23_mem/n18620 , \u_a23_mem/n18619 , \u_a23_mem/n18618 ,
         \u_a23_mem/n18617 , \u_a23_mem/n18616 , \u_a23_mem/n18615 ,
         \u_a23_mem/n18614 , \u_a23_mem/n18613 , \u_a23_mem/n18612 ,
         \u_a23_mem/n18611 , \u_a23_mem/n18610 , \u_a23_mem/n18609 ,
         \u_a23_mem/n18608 , \u_a23_mem/n18607 , \u_a23_mem/n18606 ,
         \u_a23_mem/n18605 , \u_a23_mem/n18604 , \u_a23_mem/n18603 ,
         \u_a23_mem/n18602 , \u_a23_mem/n18601 , \u_a23_mem/n18600 ,
         \u_a23_mem/n18599 , \u_a23_mem/n18598 , \u_a23_mem/n18597 ,
         \u_a23_mem/n18596 , \u_a23_mem/n18595 , \u_a23_mem/n18594 ,
         \u_a23_mem/n18593 , \u_a23_mem/n18592 , \u_a23_mem/n18591 ,
         \u_a23_mem/n18590 , \u_a23_mem/n18589 , \u_a23_mem/n18588 ,
         \u_a23_mem/n18587 , \u_a23_mem/n18586 , \u_a23_mem/n18585 ,
         \u_a23_mem/n18584 , \u_a23_mem/n18583 , \u_a23_mem/n18582 ,
         \u_a23_mem/n18581 , \u_a23_mem/n18580 , \u_a23_mem/n18579 ,
         \u_a23_mem/n18578 , \u_a23_mem/n18577 , \u_a23_mem/n18576 ,
         \u_a23_mem/n18575 , \u_a23_mem/n18574 , \u_a23_mem/n18573 ,
         \u_a23_mem/n18572 , \u_a23_mem/n18571 , \u_a23_mem/n18570 ,
         \u_a23_mem/n18569 , \u_a23_mem/n18568 , \u_a23_mem/n18567 ,
         \u_a23_mem/n18566 , \u_a23_mem/n18565 , \u_a23_mem/n18564 ,
         \u_a23_mem/n18563 , \u_a23_mem/n18562 , \u_a23_mem/n18561 ,
         \u_a23_mem/n18560 , \u_a23_mem/n18559 , \u_a23_mem/n18558 ,
         \u_a23_mem/n18557 , \u_a23_mem/n18556 , \u_a23_mem/n18555 ,
         \u_a23_mem/n18554 , \u_a23_mem/n18553 , \u_a23_mem/n18552 ,
         \u_a23_mem/n18551 , \u_a23_mem/n18550 , \u_a23_mem/n18549 ,
         \u_a23_mem/n18548 , \u_a23_mem/n18547 , \u_a23_mem/n18546 ,
         \u_a23_mem/n18545 , \u_a23_mem/n18544 , \u_a23_mem/n18543 ,
         \u_a23_mem/n18542 , \u_a23_mem/n18541 , \u_a23_mem/n18540 ,
         \u_a23_mem/n18539 , \u_a23_mem/n18538 , \u_a23_mem/n18537 ,
         \u_a23_mem/n18536 , \u_a23_mem/n18535 , \u_a23_mem/n18534 ,
         \u_a23_mem/n18533 , \u_a23_mem/n18532 , \u_a23_mem/n18531 ,
         \u_a23_mem/n18530 , \u_a23_mem/n18529 , \u_a23_mem/n18528 ,
         \u_a23_mem/n18527 , \u_a23_mem/n18526 , \u_a23_mem/n18525 ,
         \u_a23_mem/n18524 , \u_a23_mem/n18523 , \u_a23_mem/n18522 ,
         \u_a23_mem/n18521 , \u_a23_mem/n18520 , \u_a23_mem/n18519 ,
         \u_a23_mem/n18518 , \u_a23_mem/n18517 , \u_a23_mem/n18516 ,
         \u_a23_mem/n18515 , \u_a23_mem/n18514 , \u_a23_mem/n18513 ,
         \u_a23_mem/n18512 , \u_a23_mem/n18511 , \u_a23_mem/n18510 ,
         \u_a23_mem/n18509 , \u_a23_mem/n18508 , \u_a23_mem/n18507 ,
         \u_a23_mem/n18506 , \u_a23_mem/n18505 , \u_a23_mem/n18504 ,
         \u_a23_mem/n18503 , \u_a23_mem/n18502 , \u_a23_mem/n18501 ,
         \u_a23_mem/n18500 , \u_a23_mem/n18499 , \u_a23_mem/n18498 ,
         \u_a23_mem/n18497 , \u_a23_mem/n18496 , \u_a23_mem/n18495 ,
         \u_a23_mem/n18494 , \u_a23_mem/n18493 , \u_a23_mem/n18492 ,
         \u_a23_mem/n18491 , \u_a23_mem/n18490 , \u_a23_mem/n18489 ,
         \u_a23_mem/n18488 , \u_a23_mem/n18487 , \u_a23_mem/n18486 ,
         \u_a23_mem/n18485 , \u_a23_mem/n18484 , \u_a23_mem/n18483 ,
         \u_a23_mem/n18482 , \u_a23_mem/n18481 , \u_a23_mem/n18480 ,
         \u_a23_mem/n18479 , \u_a23_mem/n18478 , \u_a23_mem/n18477 ,
         \u_a23_mem/n18476 , \u_a23_mem/n18475 , \u_a23_mem/n18474 ,
         \u_a23_mem/n18473 , \u_a23_mem/n18472 , \u_a23_mem/n18471 ,
         \u_a23_mem/n18470 , \u_a23_mem/n18469 , \u_a23_mem/n18468 ,
         \u_a23_mem/n18467 , \u_a23_mem/n18466 , \u_a23_mem/n18465 ,
         \u_a23_mem/n18464 , \u_a23_mem/n18463 , \u_a23_mem/n18462 ,
         \u_a23_mem/n18461 , \u_a23_mem/n18460 , \u_a23_mem/n18459 ,
         \u_a23_mem/n18458 , \u_a23_mem/n18457 , \u_a23_mem/n18456 ,
         \u_a23_mem/n18455 , \u_a23_mem/n18454 , \u_a23_mem/n18453 ,
         \u_a23_mem/n18452 , \u_a23_mem/n18451 , \u_a23_mem/n18450 ,
         \u_a23_mem/n18449 , \u_a23_mem/n18448 , \u_a23_mem/n18447 ,
         \u_a23_mem/n18446 , \u_a23_mem/n18445 , \u_a23_mem/n18444 ,
         \u_a23_mem/n18443 , \u_a23_mem/n18442 , \u_a23_mem/n18441 ,
         \u_a23_mem/n18440 , \u_a23_mem/n18439 , \u_a23_mem/n18438 ,
         \u_a23_mem/n18437 , \u_a23_mem/n18436 , \u_a23_mem/n18435 ,
         \u_a23_mem/n18434 , \u_a23_mem/n18433 , \u_a23_mem/n18432 ,
         \u_a23_mem/n18431 , \u_a23_mem/n18430 , \u_a23_mem/n18429 ,
         \u_a23_mem/n18428 , \u_a23_mem/n18427 , \u_a23_mem/n18426 ,
         \u_a23_mem/n18425 , \u_a23_mem/n18424 , \u_a23_mem/n18423 ,
         \u_a23_mem/n18422 , \u_a23_mem/n18421 , \u_a23_mem/n18420 ,
         \u_a23_mem/n18419 , \u_a23_mem/n18418 , \u_a23_mem/n18417 ,
         \u_a23_mem/n18416 , \u_a23_mem/n18415 , \u_a23_mem/n18414 ,
         \u_a23_mem/n18413 , \u_a23_mem/n18412 , \u_a23_mem/n18411 ,
         \u_a23_mem/n18410 , \u_a23_mem/n18409 , \u_a23_mem/n18408 ,
         \u_a23_mem/n18407 , \u_a23_mem/n18406 , \u_a23_mem/n18405 ,
         \u_a23_mem/n18404 , \u_a23_mem/n18403 , \u_a23_mem/n18402 ,
         \u_a23_mem/n18401 , \u_a23_mem/n18400 , \u_a23_mem/n18399 ,
         \u_a23_mem/n18398 , \u_a23_mem/n18397 , \u_a23_mem/n18396 ,
         \u_a23_mem/n18395 , \u_a23_mem/n18394 , \u_a23_mem/n18393 ,
         \u_a23_mem/n18392 , \u_a23_mem/n18391 , \u_a23_mem/n18390 ,
         \u_a23_mem/n18389 , \u_a23_mem/n18388 , \u_a23_mem/n18387 ,
         \u_a23_mem/n18386 , \u_a23_mem/n18385 , \u_a23_mem/n18384 ,
         \u_a23_mem/n18383 , \u_a23_mem/n18382 , \u_a23_mem/n18381 ,
         \u_a23_mem/n18380 , \u_a23_mem/n18379 , \u_a23_mem/n18378 ,
         \u_a23_mem/n18377 , \u_a23_mem/n18376 , \u_a23_mem/n18375 ,
         \u_a23_mem/n18374 , \u_a23_mem/n18373 , \u_a23_mem/n18372 ,
         \u_a23_mem/n18371 , \u_a23_mem/n18370 , \u_a23_mem/n18369 ,
         \u_a23_mem/n18368 , \u_a23_mem/n18367 , \u_a23_mem/n18366 ,
         \u_a23_mem/n18365 , \u_a23_mem/n18364 , \u_a23_mem/n18363 ,
         \u_a23_mem/n18362 , \u_a23_mem/n18361 , \u_a23_mem/n18360 ,
         \u_a23_mem/n18359 , \u_a23_mem/n18358 , \u_a23_mem/n18357 ,
         \u_a23_mem/n18356 , \u_a23_mem/n18355 , \u_a23_mem/n18354 ,
         \u_a23_mem/n18353 , \u_a23_mem/n18352 , \u_a23_mem/n18351 ,
         \u_a23_mem/n18350 , \u_a23_mem/n18349 , \u_a23_mem/n18348 ,
         \u_a23_mem/n18347 , \u_a23_mem/n18346 , \u_a23_mem/n18345 ,
         \u_a23_mem/n18344 , \u_a23_mem/n18343 , \u_a23_mem/n18342 ,
         \u_a23_mem/n18341 , \u_a23_mem/n18340 , \u_a23_mem/n18339 ,
         \u_a23_mem/n18338 , \u_a23_mem/n18337 , \u_a23_mem/n18336 ,
         \u_a23_mem/n18335 , \u_a23_mem/n18334 , \u_a23_mem/n18333 ,
         \u_a23_mem/n18332 , \u_a23_mem/n18331 , \u_a23_mem/n18330 ,
         \u_a23_mem/n18329 , \u_a23_mem/n18328 , \u_a23_mem/n18327 ,
         \u_a23_mem/n18326 , \u_a23_mem/n18325 , \u_a23_mem/n18324 ,
         \u_a23_mem/n18323 , \u_a23_mem/n18322 , \u_a23_mem/n18321 ,
         \u_a23_mem/n18320 , \u_a23_mem/n18319 , \u_a23_mem/n18318 ,
         \u_a23_mem/n18317 , \u_a23_mem/n18316 , \u_a23_mem/n18315 ,
         \u_a23_mem/n18314 , \u_a23_mem/n18313 , \u_a23_mem/n18312 ,
         \u_a23_mem/n18311 , \u_a23_mem/n18310 , \u_a23_mem/n18309 ,
         \u_a23_mem/n18308 , \u_a23_mem/n18307 , \u_a23_mem/n18306 ,
         \u_a23_mem/n18305 , \u_a23_mem/n18304 , \u_a23_mem/n18303 ,
         \u_a23_mem/n18302 , \u_a23_mem/n18301 , \u_a23_mem/n18300 ,
         \u_a23_mem/n18299 , \u_a23_mem/n18298 , \u_a23_mem/n18297 ,
         \u_a23_mem/n18296 , \u_a23_mem/n18295 , \u_a23_mem/n18294 ,
         \u_a23_mem/n18293 , \u_a23_mem/n18292 , \u_a23_mem/n18291 ,
         \u_a23_mem/n18290 , \u_a23_mem/n18289 , \u_a23_mem/n18288 ,
         \u_a23_mem/n18287 , \u_a23_mem/n18286 , \u_a23_mem/n18285 ,
         \u_a23_mem/n18284 , \u_a23_mem/n18283 , \u_a23_mem/n18282 ,
         \u_a23_mem/n18281 , \u_a23_mem/n18280 , \u_a23_mem/n18279 ,
         \u_a23_mem/n18278 , \u_a23_mem/n18277 , \u_a23_mem/n18276 ,
         \u_a23_mem/n18275 , \u_a23_mem/n18274 , \u_a23_mem/n18273 ,
         \u_a23_mem/n18272 , \u_a23_mem/n18271 , \u_a23_mem/n18270 ,
         \u_a23_mem/n18269 , \u_a23_mem/n18268 , \u_a23_mem/n18267 ,
         \u_a23_mem/n18266 , \u_a23_mem/n18265 , \u_a23_mem/n18264 ,
         \u_a23_mem/n18263 , \u_a23_mem/n18262 , \u_a23_mem/n18261 ,
         \u_a23_mem/n18260 , \u_a23_mem/n18259 , \u_a23_mem/n18258 ,
         \u_a23_mem/n18257 , \u_a23_mem/n18256 , \u_a23_mem/n18255 ,
         \u_a23_mem/n18254 , \u_a23_mem/n18253 , \u_a23_mem/n18252 ,
         \u_a23_mem/n18251 , \u_a23_mem/n18250 , \u_a23_mem/n18249 ,
         \u_a23_mem/n18248 , \u_a23_mem/n18247 , \u_a23_mem/n18246 ,
         \u_a23_mem/n18245 , \u_a23_mem/n18244 , \u_a23_mem/n18243 ,
         \u_a23_mem/n18242 , \u_a23_mem/n18241 , \u_a23_mem/n18240 ,
         \u_a23_mem/n18239 , \u_a23_mem/n18238 , \u_a23_mem/n18237 ,
         \u_a23_mem/n18236 , \u_a23_mem/n18235 , \u_a23_mem/n18234 ,
         \u_a23_mem/n18233 , \u_a23_mem/n18232 , \u_a23_mem/n18231 ,
         \u_a23_mem/n18230 , \u_a23_mem/n18229 , \u_a23_mem/n18228 ,
         \u_a23_mem/n18227 , \u_a23_mem/n18226 , \u_a23_mem/n18225 ,
         \u_a23_mem/n18224 , \u_a23_mem/n18223 , \u_a23_mem/n18222 ,
         \u_a23_mem/n18221 , \u_a23_mem/n18220 , \u_a23_mem/n18219 ,
         \u_a23_mem/n18218 , \u_a23_mem/n18217 , \u_a23_mem/n18216 ,
         \u_a23_mem/n18215 , \u_a23_mem/n18214 , \u_a23_mem/n18213 ,
         \u_a23_mem/n18212 , \u_a23_mem/n18211 , \u_a23_mem/n18210 ,
         \u_a23_mem/n18209 , \u_a23_mem/n18208 , \u_a23_mem/n18207 ,
         \u_a23_mem/n18206 , \u_a23_mem/n18205 , \u_a23_mem/n18204 ,
         \u_a23_mem/n18203 , \u_a23_mem/n18202 , \u_a23_mem/n18201 ,
         \u_a23_mem/n18200 , \u_a23_mem/n18199 , \u_a23_mem/n18198 ,
         \u_a23_mem/n18197 , \u_a23_mem/n18196 , \u_a23_mem/n18195 ,
         \u_a23_mem/n18194 , \u_a23_mem/n18193 , \u_a23_mem/n18192 ,
         \u_a23_mem/n18191 , \u_a23_mem/n18190 , \u_a23_mem/n18189 ,
         \u_a23_mem/n18188 , \u_a23_mem/n18187 , \u_a23_mem/n18186 ,
         \u_a23_mem/n18185 , \u_a23_mem/n18184 , \u_a23_mem/n18183 ,
         \u_a23_mem/n18182 , \u_a23_mem/n18181 , \u_a23_mem/n18180 ,
         \u_a23_mem/n18179 , \u_a23_mem/n18178 , \u_a23_mem/n18177 ,
         \u_a23_mem/n18176 , \u_a23_mem/n18175 , \u_a23_mem/n18174 ,
         \u_a23_mem/n18173 , \u_a23_mem/n18172 , \u_a23_mem/n18171 ,
         \u_a23_mem/n18170 , \u_a23_mem/n18169 , \u_a23_mem/n18168 ,
         \u_a23_mem/n18167 , \u_a23_mem/n18166 , \u_a23_mem/n18165 ,
         \u_a23_mem/n18164 , \u_a23_mem/n18163 , \u_a23_mem/n18162 ,
         \u_a23_mem/n18161 , \u_a23_mem/n18160 , \u_a23_mem/n18159 ,
         \u_a23_mem/n18158 , \u_a23_mem/n18157 , \u_a23_mem/n18156 ,
         \u_a23_mem/n18155 , \u_a23_mem/n18154 , \u_a23_mem/n18153 ,
         \u_a23_mem/n18152 , \u_a23_mem/n18151 , \u_a23_mem/n18150 ,
         \u_a23_mem/n18149 , \u_a23_mem/n18148 , \u_a23_mem/n18147 ,
         \u_a23_mem/n18146 , \u_a23_mem/n18145 , \u_a23_mem/n18144 ,
         \u_a23_mem/n18143 , \u_a23_mem/n18142 , \u_a23_mem/n18141 ,
         \u_a23_mem/n18140 , \u_a23_mem/n18139 , \u_a23_mem/n18138 ,
         \u_a23_mem/n18137 , \u_a23_mem/n18136 , \u_a23_mem/n18135 ,
         \u_a23_mem/n18134 , \u_a23_mem/n18133 , \u_a23_mem/n18132 ,
         \u_a23_mem/n18131 , \u_a23_mem/n18130 , \u_a23_mem/n18129 ,
         \u_a23_mem/n18128 , \u_a23_mem/n18127 , \u_a23_mem/n18126 ,
         \u_a23_mem/n18125 , \u_a23_mem/n18124 , \u_a23_mem/n18123 ,
         \u_a23_mem/n18122 , \u_a23_mem/n18121 , \u_a23_mem/n18120 ,
         \u_a23_mem/n18119 , \u_a23_mem/n18118 , \u_a23_mem/n18117 ,
         \u_a23_mem/N1974 , \u_a23_mem/N1973 , \u_a23_mem/N1972 ,
         \u_a23_mem/N1971 , \u_a23_mem/N1970 , \u_a23_mem/N1969 ,
         \u_a23_mem/N1968 , \u_a23_mem/N1967 , \u_a23_mem/stack_mem[0][0] ,
         \u_a23_mem/stack_mem[0][1] , \u_a23_mem/stack_mem[0][2] ,
         \u_a23_mem/stack_mem[0][3] , \u_a23_mem/stack_mem[0][4] ,
         \u_a23_mem/stack_mem[0][5] , \u_a23_mem/stack_mem[0][6] ,
         \u_a23_mem/stack_mem[0][7] , \u_a23_mem/stack_mem[1][0] ,
         \u_a23_mem/stack_mem[1][1] , \u_a23_mem/stack_mem[1][2] ,
         \u_a23_mem/stack_mem[1][3] , \u_a23_mem/stack_mem[1][4] ,
         \u_a23_mem/stack_mem[1][5] , \u_a23_mem/stack_mem[1][6] ,
         \u_a23_mem/stack_mem[1][7] , \u_a23_mem/stack_mem[2][0] ,
         \u_a23_mem/stack_mem[2][1] , \u_a23_mem/stack_mem[2][2] ,
         \u_a23_mem/stack_mem[2][3] , \u_a23_mem/stack_mem[2][4] ,
         \u_a23_mem/stack_mem[2][5] , \u_a23_mem/stack_mem[2][6] ,
         \u_a23_mem/stack_mem[2][7] , \u_a23_mem/stack_mem[3][0] ,
         \u_a23_mem/stack_mem[3][1] , \u_a23_mem/stack_mem[3][2] ,
         \u_a23_mem/stack_mem[3][3] , \u_a23_mem/stack_mem[3][4] ,
         \u_a23_mem/stack_mem[3][5] , \u_a23_mem/stack_mem[3][6] ,
         \u_a23_mem/stack_mem[3][7] , \u_a23_mem/stack_mem[4][0] ,
         \u_a23_mem/stack_mem[4][1] , \u_a23_mem/stack_mem[4][2] ,
         \u_a23_mem/stack_mem[4][3] , \u_a23_mem/stack_mem[4][4] ,
         \u_a23_mem/stack_mem[4][5] , \u_a23_mem/stack_mem[4][6] ,
         \u_a23_mem/stack_mem[4][7] , \u_a23_mem/stack_mem[5][0] ,
         \u_a23_mem/stack_mem[5][1] , \u_a23_mem/stack_mem[5][2] ,
         \u_a23_mem/stack_mem[5][3] , \u_a23_mem/stack_mem[5][4] ,
         \u_a23_mem/stack_mem[5][5] , \u_a23_mem/stack_mem[5][6] ,
         \u_a23_mem/stack_mem[5][7] , \u_a23_mem/stack_mem[6][0] ,
         \u_a23_mem/stack_mem[6][1] , \u_a23_mem/stack_mem[6][2] ,
         \u_a23_mem/stack_mem[6][3] , \u_a23_mem/stack_mem[6][4] ,
         \u_a23_mem/stack_mem[6][5] , \u_a23_mem/stack_mem[6][6] ,
         \u_a23_mem/stack_mem[6][7] , \u_a23_mem/stack_mem[7][0] ,
         \u_a23_mem/stack_mem[7][1] , \u_a23_mem/stack_mem[7][2] ,
         \u_a23_mem/stack_mem[7][3] , \u_a23_mem/stack_mem[7][4] ,
         \u_a23_mem/stack_mem[7][5] , \u_a23_mem/stack_mem[7][6] ,
         \u_a23_mem/stack_mem[7][7] , \u_a23_mem/stack_mem[8][0] ,
         \u_a23_mem/stack_mem[8][1] , \u_a23_mem/stack_mem[8][2] ,
         \u_a23_mem/stack_mem[8][3] , \u_a23_mem/stack_mem[8][4] ,
         \u_a23_mem/stack_mem[8][5] , \u_a23_mem/stack_mem[8][6] ,
         \u_a23_mem/stack_mem[8][7] , \u_a23_mem/stack_mem[9][0] ,
         \u_a23_mem/stack_mem[9][1] , \u_a23_mem/stack_mem[9][2] ,
         \u_a23_mem/stack_mem[9][3] , \u_a23_mem/stack_mem[9][4] ,
         \u_a23_mem/stack_mem[9][5] , \u_a23_mem/stack_mem[9][6] ,
         \u_a23_mem/stack_mem[9][7] , \u_a23_mem/stack_mem[10][0] ,
         \u_a23_mem/stack_mem[10][1] , \u_a23_mem/stack_mem[10][2] ,
         \u_a23_mem/stack_mem[10][3] , \u_a23_mem/stack_mem[10][4] ,
         \u_a23_mem/stack_mem[10][5] , \u_a23_mem/stack_mem[10][6] ,
         \u_a23_mem/stack_mem[10][7] , \u_a23_mem/stack_mem[11][0] ,
         \u_a23_mem/stack_mem[11][1] , \u_a23_mem/stack_mem[11][2] ,
         \u_a23_mem/stack_mem[11][3] , \u_a23_mem/stack_mem[11][4] ,
         \u_a23_mem/stack_mem[11][5] , \u_a23_mem/stack_mem[11][6] ,
         \u_a23_mem/stack_mem[11][7] , \u_a23_mem/stack_mem[12][0] ,
         \u_a23_mem/stack_mem[12][1] , \u_a23_mem/stack_mem[12][2] ,
         \u_a23_mem/stack_mem[12][3] , \u_a23_mem/stack_mem[12][4] ,
         \u_a23_mem/stack_mem[12][5] , \u_a23_mem/stack_mem[12][6] ,
         \u_a23_mem/stack_mem[12][7] , \u_a23_mem/stack_mem[13][0] ,
         \u_a23_mem/stack_mem[13][1] , \u_a23_mem/stack_mem[13][2] ,
         \u_a23_mem/stack_mem[13][3] , \u_a23_mem/stack_mem[13][4] ,
         \u_a23_mem/stack_mem[13][5] , \u_a23_mem/stack_mem[13][6] ,
         \u_a23_mem/stack_mem[13][7] , \u_a23_mem/stack_mem[14][0] ,
         \u_a23_mem/stack_mem[14][1] , \u_a23_mem/stack_mem[14][2] ,
         \u_a23_mem/stack_mem[14][3] , \u_a23_mem/stack_mem[14][4] ,
         \u_a23_mem/stack_mem[14][5] , \u_a23_mem/stack_mem[14][6] ,
         \u_a23_mem/stack_mem[14][7] , \u_a23_mem/stack_mem[15][0] ,
         \u_a23_mem/stack_mem[15][1] , \u_a23_mem/stack_mem[15][2] ,
         \u_a23_mem/stack_mem[15][3] , \u_a23_mem/stack_mem[15][4] ,
         \u_a23_mem/stack_mem[15][5] , \u_a23_mem/stack_mem[15][6] ,
         \u_a23_mem/stack_mem[15][7] , \u_a23_mem/stack_mem[16][0] ,
         \u_a23_mem/stack_mem[16][1] , \u_a23_mem/stack_mem[16][2] ,
         \u_a23_mem/stack_mem[16][3] , \u_a23_mem/stack_mem[16][4] ,
         \u_a23_mem/stack_mem[16][5] , \u_a23_mem/stack_mem[16][6] ,
         \u_a23_mem/stack_mem[16][7] , \u_a23_mem/stack_mem[17][0] ,
         \u_a23_mem/stack_mem[17][1] , \u_a23_mem/stack_mem[17][2] ,
         \u_a23_mem/stack_mem[17][3] , \u_a23_mem/stack_mem[17][4] ,
         \u_a23_mem/stack_mem[17][5] , \u_a23_mem/stack_mem[17][6] ,
         \u_a23_mem/stack_mem[17][7] , \u_a23_mem/stack_mem[18][0] ,
         \u_a23_mem/stack_mem[18][1] , \u_a23_mem/stack_mem[18][2] ,
         \u_a23_mem/stack_mem[18][3] , \u_a23_mem/stack_mem[18][4] ,
         \u_a23_mem/stack_mem[18][5] , \u_a23_mem/stack_mem[18][6] ,
         \u_a23_mem/stack_mem[18][7] , \u_a23_mem/stack_mem[19][0] ,
         \u_a23_mem/stack_mem[19][1] , \u_a23_mem/stack_mem[19][2] ,
         \u_a23_mem/stack_mem[19][3] , \u_a23_mem/stack_mem[19][4] ,
         \u_a23_mem/stack_mem[19][5] , \u_a23_mem/stack_mem[19][6] ,
         \u_a23_mem/stack_mem[19][7] , \u_a23_mem/stack_mem[20][0] ,
         \u_a23_mem/stack_mem[20][1] , \u_a23_mem/stack_mem[20][2] ,
         \u_a23_mem/stack_mem[20][3] , \u_a23_mem/stack_mem[20][4] ,
         \u_a23_mem/stack_mem[20][5] , \u_a23_mem/stack_mem[20][6] ,
         \u_a23_mem/stack_mem[20][7] , \u_a23_mem/stack_mem[21][0] ,
         \u_a23_mem/stack_mem[21][1] , \u_a23_mem/stack_mem[21][2] ,
         \u_a23_mem/stack_mem[21][3] , \u_a23_mem/stack_mem[21][4] ,
         \u_a23_mem/stack_mem[21][5] , \u_a23_mem/stack_mem[21][6] ,
         \u_a23_mem/stack_mem[21][7] , \u_a23_mem/stack_mem[22][0] ,
         \u_a23_mem/stack_mem[22][1] , \u_a23_mem/stack_mem[22][2] ,
         \u_a23_mem/stack_mem[22][3] , \u_a23_mem/stack_mem[22][4] ,
         \u_a23_mem/stack_mem[22][5] , \u_a23_mem/stack_mem[22][6] ,
         \u_a23_mem/stack_mem[22][7] , \u_a23_mem/stack_mem[23][0] ,
         \u_a23_mem/stack_mem[23][1] , \u_a23_mem/stack_mem[23][2] ,
         \u_a23_mem/stack_mem[23][3] , \u_a23_mem/stack_mem[23][4] ,
         \u_a23_mem/stack_mem[23][5] , \u_a23_mem/stack_mem[23][6] ,
         \u_a23_mem/stack_mem[23][7] , \u_a23_mem/stack_mem[24][0] ,
         \u_a23_mem/stack_mem[24][1] , \u_a23_mem/stack_mem[24][2] ,
         \u_a23_mem/stack_mem[24][3] , \u_a23_mem/stack_mem[24][4] ,
         \u_a23_mem/stack_mem[24][5] , \u_a23_mem/stack_mem[24][6] ,
         \u_a23_mem/stack_mem[24][7] , \u_a23_mem/stack_mem[25][0] ,
         \u_a23_mem/stack_mem[25][1] , \u_a23_mem/stack_mem[25][2] ,
         \u_a23_mem/stack_mem[25][3] , \u_a23_mem/stack_mem[25][4] ,
         \u_a23_mem/stack_mem[25][5] , \u_a23_mem/stack_mem[25][6] ,
         \u_a23_mem/stack_mem[25][7] , \u_a23_mem/stack_mem[26][0] ,
         \u_a23_mem/stack_mem[26][1] , \u_a23_mem/stack_mem[26][2] ,
         \u_a23_mem/stack_mem[26][3] , \u_a23_mem/stack_mem[26][4] ,
         \u_a23_mem/stack_mem[26][5] , \u_a23_mem/stack_mem[26][6] ,
         \u_a23_mem/stack_mem[26][7] , \u_a23_mem/stack_mem[27][0] ,
         \u_a23_mem/stack_mem[27][1] , \u_a23_mem/stack_mem[27][2] ,
         \u_a23_mem/stack_mem[27][3] , \u_a23_mem/stack_mem[27][4] ,
         \u_a23_mem/stack_mem[27][5] , \u_a23_mem/stack_mem[27][6] ,
         \u_a23_mem/stack_mem[27][7] , \u_a23_mem/stack_mem[28][0] ,
         \u_a23_mem/stack_mem[28][1] , \u_a23_mem/stack_mem[28][2] ,
         \u_a23_mem/stack_mem[28][3] , \u_a23_mem/stack_mem[28][4] ,
         \u_a23_mem/stack_mem[28][5] , \u_a23_mem/stack_mem[28][6] ,
         \u_a23_mem/stack_mem[28][7] , \u_a23_mem/stack_mem[29][0] ,
         \u_a23_mem/stack_mem[29][1] , \u_a23_mem/stack_mem[29][2] ,
         \u_a23_mem/stack_mem[29][3] , \u_a23_mem/stack_mem[29][4] ,
         \u_a23_mem/stack_mem[29][5] , \u_a23_mem/stack_mem[29][6] ,
         \u_a23_mem/stack_mem[29][7] , \u_a23_mem/stack_mem[30][0] ,
         \u_a23_mem/stack_mem[30][1] , \u_a23_mem/stack_mem[30][2] ,
         \u_a23_mem/stack_mem[30][3] , \u_a23_mem/stack_mem[30][4] ,
         \u_a23_mem/stack_mem[30][5] , \u_a23_mem/stack_mem[30][6] ,
         \u_a23_mem/stack_mem[30][7] , \u_a23_mem/stack_mem[31][0] ,
         \u_a23_mem/stack_mem[31][1] , \u_a23_mem/stack_mem[31][2] ,
         \u_a23_mem/stack_mem[31][3] , \u_a23_mem/stack_mem[31][4] ,
         \u_a23_mem/stack_mem[31][5] , \u_a23_mem/stack_mem[31][6] ,
         \u_a23_mem/stack_mem[31][7] , \u_a23_mem/N1942 , \u_a23_mem/N1941 ,
         \u_a23_mem/N1940 , \u_a23_mem/N1939 , \u_a23_mem/N1938 ,
         \u_a23_mem/N1937 , \u_a23_mem/N1936 , \u_a23_mem/N1935 ,
         \u_a23_mem/N1910 , \u_a23_mem/N1909 , \u_a23_mem/N1908 ,
         \u_a23_mem/N1907 , \u_a23_mem/N1906 , \u_a23_mem/N1905 ,
         \u_a23_mem/N1904 , \u_a23_mem/N1903 , \u_a23_mem/e_mem[0][0] ,
         \u_a23_mem/e_mem[0][1] , \u_a23_mem/e_mem[0][2] ,
         \u_a23_mem/e_mem[0][3] , \u_a23_mem/e_mem[0][4] ,
         \u_a23_mem/e_mem[0][5] , \u_a23_mem/e_mem[0][6] ,
         \u_a23_mem/e_mem[0][7] , \u_a23_mem/e_mem[1][0] ,
         \u_a23_mem/e_mem[1][1] , \u_a23_mem/e_mem[1][2] ,
         \u_a23_mem/e_mem[1][3] , \u_a23_mem/e_mem[1][4] ,
         \u_a23_mem/e_mem[1][5] , \u_a23_mem/e_mem[1][6] ,
         \u_a23_mem/e_mem[1][7] , \u_a23_mem/e_mem[2][0] ,
         \u_a23_mem/e_mem[2][1] , \u_a23_mem/e_mem[2][2] ,
         \u_a23_mem/e_mem[2][3] , \u_a23_mem/e_mem[2][4] ,
         \u_a23_mem/e_mem[2][5] , \u_a23_mem/e_mem[2][6] ,
         \u_a23_mem/e_mem[2][7] , \u_a23_mem/e_mem[3][0] ,
         \u_a23_mem/e_mem[3][1] , \u_a23_mem/e_mem[3][2] ,
         \u_a23_mem/e_mem[3][3] , \u_a23_mem/e_mem[3][4] ,
         \u_a23_mem/e_mem[3][5] , \u_a23_mem/e_mem[3][6] ,
         \u_a23_mem/e_mem[3][7] , \u_a23_mem/e_mem[4][0] ,
         \u_a23_mem/e_mem[4][1] , \u_a23_mem/e_mem[4][2] ,
         \u_a23_mem/e_mem[4][3] , \u_a23_mem/e_mem[4][4] ,
         \u_a23_mem/e_mem[4][5] , \u_a23_mem/e_mem[4][6] ,
         \u_a23_mem/e_mem[4][7] , \u_a23_mem/e_mem[5][0] ,
         \u_a23_mem/e_mem[5][1] , \u_a23_mem/e_mem[5][2] ,
         \u_a23_mem/e_mem[5][3] , \u_a23_mem/e_mem[5][4] ,
         \u_a23_mem/e_mem[5][5] , \u_a23_mem/e_mem[5][6] ,
         \u_a23_mem/e_mem[5][7] , \u_a23_mem/e_mem[6][0] ,
         \u_a23_mem/e_mem[6][1] , \u_a23_mem/e_mem[6][2] ,
         \u_a23_mem/e_mem[6][3] , \u_a23_mem/e_mem[6][4] ,
         \u_a23_mem/e_mem[6][5] , \u_a23_mem/e_mem[6][6] ,
         \u_a23_mem/e_mem[6][7] , \u_a23_mem/e_mem[7][0] ,
         \u_a23_mem/e_mem[7][1] , \u_a23_mem/e_mem[7][2] ,
         \u_a23_mem/e_mem[7][3] , \u_a23_mem/e_mem[7][4] ,
         \u_a23_mem/e_mem[7][5] , \u_a23_mem/e_mem[7][6] ,
         \u_a23_mem/e_mem[7][7] , \u_a23_mem/e_mem[8][0] ,
         \u_a23_mem/e_mem[8][1] , \u_a23_mem/e_mem[8][2] ,
         \u_a23_mem/e_mem[8][3] , \u_a23_mem/e_mem[8][4] ,
         \u_a23_mem/e_mem[8][5] , \u_a23_mem/e_mem[8][6] ,
         \u_a23_mem/e_mem[8][7] , \u_a23_mem/e_mem[9][0] ,
         \u_a23_mem/e_mem[9][1] , \u_a23_mem/e_mem[9][2] ,
         \u_a23_mem/e_mem[9][3] , \u_a23_mem/e_mem[9][4] ,
         \u_a23_mem/e_mem[9][5] , \u_a23_mem/e_mem[9][6] ,
         \u_a23_mem/e_mem[9][7] , \u_a23_mem/e_mem[10][0] ,
         \u_a23_mem/e_mem[10][1] , \u_a23_mem/e_mem[10][2] ,
         \u_a23_mem/e_mem[10][3] , \u_a23_mem/e_mem[10][4] ,
         \u_a23_mem/e_mem[10][5] , \u_a23_mem/e_mem[10][6] ,
         \u_a23_mem/e_mem[10][7] , \u_a23_mem/e_mem[11][0] ,
         \u_a23_mem/e_mem[11][1] , \u_a23_mem/e_mem[11][2] ,
         \u_a23_mem/e_mem[11][3] , \u_a23_mem/e_mem[11][4] ,
         \u_a23_mem/e_mem[11][5] , \u_a23_mem/e_mem[11][6] ,
         \u_a23_mem/e_mem[11][7] , \u_a23_mem/e_mem[12][0] ,
         \u_a23_mem/e_mem[12][1] , \u_a23_mem/e_mem[12][2] ,
         \u_a23_mem/e_mem[12][3] , \u_a23_mem/e_mem[12][4] ,
         \u_a23_mem/e_mem[12][5] , \u_a23_mem/e_mem[12][6] ,
         \u_a23_mem/e_mem[12][7] , \u_a23_mem/e_mem[13][0] ,
         \u_a23_mem/e_mem[13][1] , \u_a23_mem/e_mem[13][2] ,
         \u_a23_mem/e_mem[13][3] , \u_a23_mem/e_mem[13][4] ,
         \u_a23_mem/e_mem[13][5] , \u_a23_mem/e_mem[13][6] ,
         \u_a23_mem/e_mem[13][7] , \u_a23_mem/e_mem[14][0] ,
         \u_a23_mem/e_mem[14][1] , \u_a23_mem/e_mem[14][2] ,
         \u_a23_mem/e_mem[14][3] , \u_a23_mem/e_mem[14][4] ,
         \u_a23_mem/e_mem[14][5] , \u_a23_mem/e_mem[14][6] ,
         \u_a23_mem/e_mem[14][7] , \u_a23_mem/e_mem[15][0] ,
         \u_a23_mem/e_mem[15][1] , \u_a23_mem/e_mem[15][2] ,
         \u_a23_mem/e_mem[15][3] , \u_a23_mem/e_mem[15][4] ,
         \u_a23_mem/e_mem[15][5] , \u_a23_mem/e_mem[15][6] ,
         \u_a23_mem/e_mem[15][7] , \u_a23_mem/e_mem[16][0] ,
         \u_a23_mem/e_mem[16][1] , \u_a23_mem/e_mem[16][2] ,
         \u_a23_mem/e_mem[16][3] , \u_a23_mem/e_mem[16][4] ,
         \u_a23_mem/e_mem[16][5] , \u_a23_mem/e_mem[16][6] ,
         \u_a23_mem/e_mem[16][7] , \u_a23_mem/e_mem[17][0] ,
         \u_a23_mem/e_mem[17][1] , \u_a23_mem/e_mem[17][2] ,
         \u_a23_mem/e_mem[17][3] , \u_a23_mem/e_mem[17][4] ,
         \u_a23_mem/e_mem[17][5] , \u_a23_mem/e_mem[17][6] ,
         \u_a23_mem/e_mem[17][7] , \u_a23_mem/e_mem[18][0] ,
         \u_a23_mem/e_mem[18][1] , \u_a23_mem/e_mem[18][2] ,
         \u_a23_mem/e_mem[18][3] , \u_a23_mem/e_mem[18][4] ,
         \u_a23_mem/e_mem[18][5] , \u_a23_mem/e_mem[18][6] ,
         \u_a23_mem/e_mem[18][7] , \u_a23_mem/e_mem[19][0] ,
         \u_a23_mem/e_mem[19][1] , \u_a23_mem/e_mem[19][2] ,
         \u_a23_mem/e_mem[19][3] , \u_a23_mem/e_mem[19][4] ,
         \u_a23_mem/e_mem[19][5] , \u_a23_mem/e_mem[19][6] ,
         \u_a23_mem/e_mem[19][7] , \u_a23_mem/e_mem[20][0] ,
         \u_a23_mem/e_mem[20][1] , \u_a23_mem/e_mem[20][2] ,
         \u_a23_mem/e_mem[20][3] , \u_a23_mem/e_mem[20][4] ,
         \u_a23_mem/e_mem[20][5] , \u_a23_mem/e_mem[20][6] ,
         \u_a23_mem/e_mem[20][7] , \u_a23_mem/e_mem[21][0] ,
         \u_a23_mem/e_mem[21][1] , \u_a23_mem/e_mem[21][2] ,
         \u_a23_mem/e_mem[21][3] , \u_a23_mem/e_mem[21][4] ,
         \u_a23_mem/e_mem[21][5] , \u_a23_mem/e_mem[21][6] ,
         \u_a23_mem/e_mem[21][7] , \u_a23_mem/e_mem[22][0] ,
         \u_a23_mem/e_mem[22][1] , \u_a23_mem/e_mem[22][2] ,
         \u_a23_mem/e_mem[22][3] , \u_a23_mem/e_mem[22][4] ,
         \u_a23_mem/e_mem[22][5] , \u_a23_mem/e_mem[22][6] ,
         \u_a23_mem/e_mem[22][7] , \u_a23_mem/e_mem[23][0] ,
         \u_a23_mem/e_mem[23][1] , \u_a23_mem/e_mem[23][2] ,
         \u_a23_mem/e_mem[23][3] , \u_a23_mem/e_mem[23][4] ,
         \u_a23_mem/e_mem[23][5] , \u_a23_mem/e_mem[23][6] ,
         \u_a23_mem/e_mem[23][7] , \u_a23_mem/e_mem[24][0] ,
         \u_a23_mem/e_mem[24][1] , \u_a23_mem/e_mem[24][2] ,
         \u_a23_mem/e_mem[24][3] , \u_a23_mem/e_mem[24][4] ,
         \u_a23_mem/e_mem[24][5] , \u_a23_mem/e_mem[24][6] ,
         \u_a23_mem/e_mem[24][7] , \u_a23_mem/e_mem[25][0] ,
         \u_a23_mem/e_mem[25][1] , \u_a23_mem/e_mem[25][2] ,
         \u_a23_mem/e_mem[25][3] , \u_a23_mem/e_mem[25][4] ,
         \u_a23_mem/e_mem[25][5] , \u_a23_mem/e_mem[25][6] ,
         \u_a23_mem/e_mem[25][7] , \u_a23_mem/e_mem[26][0] ,
         \u_a23_mem/e_mem[26][1] , \u_a23_mem/e_mem[26][2] ,
         \u_a23_mem/e_mem[26][3] , \u_a23_mem/e_mem[26][4] ,
         \u_a23_mem/e_mem[26][5] , \u_a23_mem/e_mem[26][6] ,
         \u_a23_mem/e_mem[26][7] , \u_a23_mem/e_mem[27][0] ,
         \u_a23_mem/e_mem[27][1] , \u_a23_mem/e_mem[27][2] ,
         \u_a23_mem/e_mem[27][3] , \u_a23_mem/e_mem[27][4] ,
         \u_a23_mem/e_mem[27][5] , \u_a23_mem/e_mem[27][6] ,
         \u_a23_mem/e_mem[27][7] , \u_a23_mem/e_mem[28][0] ,
         \u_a23_mem/e_mem[28][1] , \u_a23_mem/e_mem[28][2] ,
         \u_a23_mem/e_mem[28][3] , \u_a23_mem/e_mem[28][4] ,
         \u_a23_mem/e_mem[28][5] , \u_a23_mem/e_mem[28][6] ,
         \u_a23_mem/e_mem[28][7] , \u_a23_mem/e_mem[29][0] ,
         \u_a23_mem/e_mem[29][1] , \u_a23_mem/e_mem[29][2] ,
         \u_a23_mem/e_mem[29][3] , \u_a23_mem/e_mem[29][4] ,
         \u_a23_mem/e_mem[29][5] , \u_a23_mem/e_mem[29][6] ,
         \u_a23_mem/e_mem[29][7] , \u_a23_mem/e_mem[30][0] ,
         \u_a23_mem/e_mem[30][1] , \u_a23_mem/e_mem[30][2] ,
         \u_a23_mem/e_mem[30][3] , \u_a23_mem/e_mem[30][4] ,
         \u_a23_mem/e_mem[30][5] , \u_a23_mem/e_mem[30][6] ,
         \u_a23_mem/e_mem[30][7] , \u_a23_mem/e_mem[31][0] ,
         \u_a23_mem/e_mem[31][1] , \u_a23_mem/e_mem[31][2] ,
         \u_a23_mem/e_mem[31][3] , \u_a23_mem/e_mem[31][4] ,
         \u_a23_mem/e_mem[31][5] , \u_a23_mem/e_mem[31][6] ,
         \u_a23_mem/e_mem[31][7] , \u_a23_mem/N1878 , \u_a23_mem/N1877 ,
         \u_a23_mem/N1876 , \u_a23_mem/N1875 , \u_a23_mem/N1874 ,
         \u_a23_mem/N1873 , \u_a23_mem/N1872 , \u_a23_mem/N1871 ,
         \u_a23_mem/g_mem[0][0] , \u_a23_mem/g_mem[0][1] ,
         \u_a23_mem/g_mem[0][2] , \u_a23_mem/g_mem[0][3] ,
         \u_a23_mem/g_mem[0][4] , \u_a23_mem/g_mem[0][5] ,
         \u_a23_mem/g_mem[0][6] , \u_a23_mem/g_mem[0][7] ,
         \u_a23_mem/g_mem[1][0] , \u_a23_mem/g_mem[1][1] ,
         \u_a23_mem/g_mem[1][2] , \u_a23_mem/g_mem[1][3] ,
         \u_a23_mem/g_mem[1][4] , \u_a23_mem/g_mem[1][5] ,
         \u_a23_mem/g_mem[1][6] , \u_a23_mem/g_mem[1][7] ,
         \u_a23_mem/g_mem[2][0] , \u_a23_mem/g_mem[2][1] ,
         \u_a23_mem/g_mem[2][2] , \u_a23_mem/g_mem[2][3] ,
         \u_a23_mem/g_mem[2][4] , \u_a23_mem/g_mem[2][5] ,
         \u_a23_mem/g_mem[2][6] , \u_a23_mem/g_mem[2][7] ,
         \u_a23_mem/g_mem[3][0] , \u_a23_mem/g_mem[3][1] ,
         \u_a23_mem/g_mem[3][2] , \u_a23_mem/g_mem[3][3] ,
         \u_a23_mem/g_mem[3][4] , \u_a23_mem/g_mem[3][5] ,
         \u_a23_mem/g_mem[3][6] , \u_a23_mem/g_mem[3][7] ,
         \u_a23_mem/g_mem[4][0] , \u_a23_mem/g_mem[4][1] ,
         \u_a23_mem/g_mem[4][2] , \u_a23_mem/g_mem[4][3] ,
         \u_a23_mem/g_mem[4][4] , \u_a23_mem/g_mem[4][5] ,
         \u_a23_mem/g_mem[4][6] , \u_a23_mem/g_mem[4][7] ,
         \u_a23_mem/g_mem[5][0] , \u_a23_mem/g_mem[5][1] ,
         \u_a23_mem/g_mem[5][2] , \u_a23_mem/g_mem[5][3] ,
         \u_a23_mem/g_mem[5][4] , \u_a23_mem/g_mem[5][5] ,
         \u_a23_mem/g_mem[5][6] , \u_a23_mem/g_mem[5][7] ,
         \u_a23_mem/g_mem[6][0] , \u_a23_mem/g_mem[6][1] ,
         \u_a23_mem/g_mem[6][2] , \u_a23_mem/g_mem[6][3] ,
         \u_a23_mem/g_mem[6][4] , \u_a23_mem/g_mem[6][5] ,
         \u_a23_mem/g_mem[6][6] , \u_a23_mem/g_mem[6][7] ,
         \u_a23_mem/g_mem[7][0] , \u_a23_mem/g_mem[7][1] ,
         \u_a23_mem/g_mem[7][2] , \u_a23_mem/g_mem[7][3] ,
         \u_a23_mem/g_mem[7][4] , \u_a23_mem/g_mem[7][5] ,
         \u_a23_mem/g_mem[7][6] , \u_a23_mem/g_mem[7][7] ,
         \u_a23_mem/g_mem[8][0] , \u_a23_mem/g_mem[8][1] ,
         \u_a23_mem/g_mem[8][2] , \u_a23_mem/g_mem[8][3] ,
         \u_a23_mem/g_mem[8][4] , \u_a23_mem/g_mem[8][5] ,
         \u_a23_mem/g_mem[8][6] , \u_a23_mem/g_mem[8][7] ,
         \u_a23_mem/g_mem[9][0] , \u_a23_mem/g_mem[9][1] ,
         \u_a23_mem/g_mem[9][2] , \u_a23_mem/g_mem[9][3] ,
         \u_a23_mem/g_mem[9][4] , \u_a23_mem/g_mem[9][5] ,
         \u_a23_mem/g_mem[9][6] , \u_a23_mem/g_mem[9][7] ,
         \u_a23_mem/g_mem[10][0] , \u_a23_mem/g_mem[10][1] ,
         \u_a23_mem/g_mem[10][2] , \u_a23_mem/g_mem[10][3] ,
         \u_a23_mem/g_mem[10][4] , \u_a23_mem/g_mem[10][5] ,
         \u_a23_mem/g_mem[10][6] , \u_a23_mem/g_mem[10][7] ,
         \u_a23_mem/g_mem[11][0] , \u_a23_mem/g_mem[11][1] ,
         \u_a23_mem/g_mem[11][2] , \u_a23_mem/g_mem[11][3] ,
         \u_a23_mem/g_mem[11][4] , \u_a23_mem/g_mem[11][5] ,
         \u_a23_mem/g_mem[11][6] , \u_a23_mem/g_mem[11][7] ,
         \u_a23_mem/g_mem[12][0] , \u_a23_mem/g_mem[12][1] ,
         \u_a23_mem/g_mem[12][2] , \u_a23_mem/g_mem[12][3] ,
         \u_a23_mem/g_mem[12][4] , \u_a23_mem/g_mem[12][5] ,
         \u_a23_mem/g_mem[12][6] , \u_a23_mem/g_mem[12][7] ,
         \u_a23_mem/g_mem[13][0] , \u_a23_mem/g_mem[13][1] ,
         \u_a23_mem/g_mem[13][2] , \u_a23_mem/g_mem[13][3] ,
         \u_a23_mem/g_mem[13][4] , \u_a23_mem/g_mem[13][5] ,
         \u_a23_mem/g_mem[13][6] , \u_a23_mem/g_mem[13][7] ,
         \u_a23_mem/g_mem[14][0] , \u_a23_mem/g_mem[14][1] ,
         \u_a23_mem/g_mem[14][2] , \u_a23_mem/g_mem[14][3] ,
         \u_a23_mem/g_mem[14][4] , \u_a23_mem/g_mem[14][5] ,
         \u_a23_mem/g_mem[14][6] , \u_a23_mem/g_mem[14][7] ,
         \u_a23_mem/g_mem[15][0] , \u_a23_mem/g_mem[15][1] ,
         \u_a23_mem/g_mem[15][2] , \u_a23_mem/g_mem[15][3] ,
         \u_a23_mem/g_mem[15][4] , \u_a23_mem/g_mem[15][5] ,
         \u_a23_mem/g_mem[15][6] , \u_a23_mem/g_mem[15][7] ,
         \u_a23_mem/g_mem[16][0] , \u_a23_mem/g_mem[16][1] ,
         \u_a23_mem/g_mem[16][2] , \u_a23_mem/g_mem[16][3] ,
         \u_a23_mem/g_mem[16][4] , \u_a23_mem/g_mem[16][5] ,
         \u_a23_mem/g_mem[16][6] , \u_a23_mem/g_mem[16][7] ,
         \u_a23_mem/g_mem[17][0] , \u_a23_mem/g_mem[17][1] ,
         \u_a23_mem/g_mem[17][2] , \u_a23_mem/g_mem[17][3] ,
         \u_a23_mem/g_mem[17][4] , \u_a23_mem/g_mem[17][5] ,
         \u_a23_mem/g_mem[17][6] , \u_a23_mem/g_mem[17][7] ,
         \u_a23_mem/g_mem[18][0] , \u_a23_mem/g_mem[18][1] ,
         \u_a23_mem/g_mem[18][2] , \u_a23_mem/g_mem[18][3] ,
         \u_a23_mem/g_mem[18][4] , \u_a23_mem/g_mem[18][5] ,
         \u_a23_mem/g_mem[18][6] , \u_a23_mem/g_mem[18][7] ,
         \u_a23_mem/g_mem[19][0] , \u_a23_mem/g_mem[19][1] ,
         \u_a23_mem/g_mem[19][2] , \u_a23_mem/g_mem[19][3] ,
         \u_a23_mem/g_mem[19][4] , \u_a23_mem/g_mem[19][5] ,
         \u_a23_mem/g_mem[19][6] , \u_a23_mem/g_mem[19][7] ,
         \u_a23_mem/g_mem[20][0] , \u_a23_mem/g_mem[20][1] ,
         \u_a23_mem/g_mem[20][2] , \u_a23_mem/g_mem[20][3] ,
         \u_a23_mem/g_mem[20][4] , \u_a23_mem/g_mem[20][5] ,
         \u_a23_mem/g_mem[20][6] , \u_a23_mem/g_mem[20][7] ,
         \u_a23_mem/g_mem[21][0] , \u_a23_mem/g_mem[21][1] ,
         \u_a23_mem/g_mem[21][2] , \u_a23_mem/g_mem[21][3] ,
         \u_a23_mem/g_mem[21][4] , \u_a23_mem/g_mem[21][5] ,
         \u_a23_mem/g_mem[21][6] , \u_a23_mem/g_mem[21][7] ,
         \u_a23_mem/g_mem[22][0] , \u_a23_mem/g_mem[22][1] ,
         \u_a23_mem/g_mem[22][2] , \u_a23_mem/g_mem[22][3] ,
         \u_a23_mem/g_mem[22][4] , \u_a23_mem/g_mem[22][5] ,
         \u_a23_mem/g_mem[22][6] , \u_a23_mem/g_mem[22][7] ,
         \u_a23_mem/g_mem[23][0] , \u_a23_mem/g_mem[23][1] ,
         \u_a23_mem/g_mem[23][2] , \u_a23_mem/g_mem[23][3] ,
         \u_a23_mem/g_mem[23][4] , \u_a23_mem/g_mem[23][5] ,
         \u_a23_mem/g_mem[23][6] , \u_a23_mem/g_mem[23][7] ,
         \u_a23_mem/g_mem[24][0] , \u_a23_mem/g_mem[24][1] ,
         \u_a23_mem/g_mem[24][2] , \u_a23_mem/g_mem[24][3] ,
         \u_a23_mem/g_mem[24][4] , \u_a23_mem/g_mem[24][5] ,
         \u_a23_mem/g_mem[24][6] , \u_a23_mem/g_mem[24][7] ,
         \u_a23_mem/g_mem[25][0] , \u_a23_mem/g_mem[25][1] ,
         \u_a23_mem/g_mem[25][2] , \u_a23_mem/g_mem[25][3] ,
         \u_a23_mem/g_mem[25][4] , \u_a23_mem/g_mem[25][5] ,
         \u_a23_mem/g_mem[25][6] , \u_a23_mem/g_mem[25][7] ,
         \u_a23_mem/g_mem[26][0] , \u_a23_mem/g_mem[26][1] ,
         \u_a23_mem/g_mem[26][2] , \u_a23_mem/g_mem[26][3] ,
         \u_a23_mem/g_mem[26][4] , \u_a23_mem/g_mem[26][5] ,
         \u_a23_mem/g_mem[26][6] , \u_a23_mem/g_mem[26][7] ,
         \u_a23_mem/g_mem[27][0] , \u_a23_mem/g_mem[27][1] ,
         \u_a23_mem/g_mem[27][2] , \u_a23_mem/g_mem[27][3] ,
         \u_a23_mem/g_mem[27][4] , \u_a23_mem/g_mem[27][5] ,
         \u_a23_mem/g_mem[27][6] , \u_a23_mem/g_mem[27][7] ,
         \u_a23_mem/g_mem[28][0] , \u_a23_mem/g_mem[28][1] ,
         \u_a23_mem/g_mem[28][2] , \u_a23_mem/g_mem[28][3] ,
         \u_a23_mem/g_mem[28][4] , \u_a23_mem/g_mem[28][5] ,
         \u_a23_mem/g_mem[28][6] , \u_a23_mem/g_mem[28][7] ,
         \u_a23_mem/g_mem[29][0] , \u_a23_mem/g_mem[29][1] ,
         \u_a23_mem/g_mem[29][2] , \u_a23_mem/g_mem[29][3] ,
         \u_a23_mem/g_mem[29][4] , \u_a23_mem/g_mem[29][5] ,
         \u_a23_mem/g_mem[29][6] , \u_a23_mem/g_mem[29][7] ,
         \u_a23_mem/g_mem[30][0] , \u_a23_mem/g_mem[30][1] ,
         \u_a23_mem/g_mem[30][2] , \u_a23_mem/g_mem[30][3] ,
         \u_a23_mem/g_mem[30][4] , \u_a23_mem/g_mem[30][5] ,
         \u_a23_mem/g_mem[30][6] , \u_a23_mem/g_mem[30][7] ,
         \u_a23_mem/g_mem[31][0] , \u_a23_mem/g_mem[31][1] ,
         \u_a23_mem/g_mem[31][2] , \u_a23_mem/g_mem[31][3] ,
         \u_a23_mem/g_mem[31][4] , \u_a23_mem/g_mem[31][5] ,
         \u_a23_mem/g_mem[31][6] , \u_a23_mem/g_mem[31][7] , \u_a23_mem/N1846 ,
         \u_a23_mem/N1845 , \u_a23_mem/N1844 , \u_a23_mem/N1843 ,
         \u_a23_mem/N1842 , \u_a23_mem/N1841 , \u_a23_mem/N1840 ,
         \u_a23_mem/N1839 , \u_a23_mem/p_mem[0][0] , \u_a23_mem/p_mem[0][1] ,
         \u_a23_mem/p_mem[0][2] , \u_a23_mem/p_mem[0][3] ,
         \u_a23_mem/p_mem[0][4] , \u_a23_mem/p_mem[0][5] ,
         \u_a23_mem/p_mem[0][6] , \u_a23_mem/p_mem[0][7] ,
         \u_a23_mem/p_mem[1][0] , \u_a23_mem/p_mem[1][1] ,
         \u_a23_mem/p_mem[1][2] , \u_a23_mem/p_mem[1][3] ,
         \u_a23_mem/p_mem[1][4] , \u_a23_mem/p_mem[1][5] ,
         \u_a23_mem/p_mem[1][6] , \u_a23_mem/p_mem[1][7] ,
         \u_a23_mem/p_mem[2][0] , \u_a23_mem/p_mem[2][1] ,
         \u_a23_mem/p_mem[2][2] , \u_a23_mem/p_mem[2][3] ,
         \u_a23_mem/p_mem[2][4] , \u_a23_mem/p_mem[2][5] ,
         \u_a23_mem/p_mem[2][6] , \u_a23_mem/p_mem[2][7] ,
         \u_a23_mem/p_mem[3][0] , \u_a23_mem/p_mem[3][1] ,
         \u_a23_mem/p_mem[3][2] , \u_a23_mem/p_mem[3][3] ,
         \u_a23_mem/p_mem[3][4] , \u_a23_mem/p_mem[3][5] ,
         \u_a23_mem/p_mem[3][6] , \u_a23_mem/p_mem[3][7] ,
         \u_a23_mem/p_mem[4][0] , \u_a23_mem/p_mem[4][1] ,
         \u_a23_mem/p_mem[4][2] , \u_a23_mem/p_mem[4][3] ,
         \u_a23_mem/p_mem[4][4] , \u_a23_mem/p_mem[4][5] ,
         \u_a23_mem/p_mem[4][6] , \u_a23_mem/p_mem[4][7] ,
         \u_a23_mem/p_mem[5][0] , \u_a23_mem/p_mem[5][1] ,
         \u_a23_mem/p_mem[5][2] , \u_a23_mem/p_mem[5][3] ,
         \u_a23_mem/p_mem[5][4] , \u_a23_mem/p_mem[5][5] ,
         \u_a23_mem/p_mem[5][6] , \u_a23_mem/p_mem[5][7] ,
         \u_a23_mem/p_mem[6][0] , \u_a23_mem/p_mem[6][1] ,
         \u_a23_mem/p_mem[6][2] , \u_a23_mem/p_mem[6][3] ,
         \u_a23_mem/p_mem[6][4] , \u_a23_mem/p_mem[6][5] ,
         \u_a23_mem/p_mem[6][6] , \u_a23_mem/p_mem[6][7] ,
         \u_a23_mem/p_mem[7][0] , \u_a23_mem/p_mem[7][1] ,
         \u_a23_mem/p_mem[7][2] , \u_a23_mem/p_mem[7][3] ,
         \u_a23_mem/p_mem[7][4] , \u_a23_mem/p_mem[7][5] ,
         \u_a23_mem/p_mem[7][6] , \u_a23_mem/p_mem[7][7] ,
         \u_a23_mem/p_mem[8][0] , \u_a23_mem/p_mem[8][1] ,
         \u_a23_mem/p_mem[8][2] , \u_a23_mem/p_mem[8][3] ,
         \u_a23_mem/p_mem[8][4] , \u_a23_mem/p_mem[8][5] ,
         \u_a23_mem/p_mem[8][6] , \u_a23_mem/p_mem[8][7] ,
         \u_a23_mem/p_mem[9][0] , \u_a23_mem/p_mem[9][1] ,
         \u_a23_mem/p_mem[9][2] , \u_a23_mem/p_mem[9][3] ,
         \u_a23_mem/p_mem[9][4] , \u_a23_mem/p_mem[9][5] ,
         \u_a23_mem/p_mem[9][6] , \u_a23_mem/p_mem[9][7] ,
         \u_a23_mem/p_mem[10][0] , \u_a23_mem/p_mem[10][1] ,
         \u_a23_mem/p_mem[10][2] , \u_a23_mem/p_mem[10][3] ,
         \u_a23_mem/p_mem[10][4] , \u_a23_mem/p_mem[10][5] ,
         \u_a23_mem/p_mem[10][6] , \u_a23_mem/p_mem[10][7] ,
         \u_a23_mem/p_mem[11][0] , \u_a23_mem/p_mem[11][1] ,
         \u_a23_mem/p_mem[11][2] , \u_a23_mem/p_mem[11][3] ,
         \u_a23_mem/p_mem[11][4] , \u_a23_mem/p_mem[11][5] ,
         \u_a23_mem/p_mem[11][6] , \u_a23_mem/p_mem[11][7] ,
         \u_a23_mem/p_mem[12][0] , \u_a23_mem/p_mem[12][1] ,
         \u_a23_mem/p_mem[12][2] , \u_a23_mem/p_mem[12][3] ,
         \u_a23_mem/p_mem[12][4] , \u_a23_mem/p_mem[12][5] ,
         \u_a23_mem/p_mem[12][6] , \u_a23_mem/p_mem[12][7] ,
         \u_a23_mem/p_mem[13][0] , \u_a23_mem/p_mem[13][1] ,
         \u_a23_mem/p_mem[13][2] , \u_a23_mem/p_mem[13][3] ,
         \u_a23_mem/p_mem[13][4] , \u_a23_mem/p_mem[13][5] ,
         \u_a23_mem/p_mem[13][6] , \u_a23_mem/p_mem[13][7] ,
         \u_a23_mem/p_mem[14][0] , \u_a23_mem/p_mem[14][1] ,
         \u_a23_mem/p_mem[14][2] , \u_a23_mem/p_mem[14][3] ,
         \u_a23_mem/p_mem[14][4] , \u_a23_mem/p_mem[14][5] ,
         \u_a23_mem/p_mem[14][6] , \u_a23_mem/p_mem[14][7] ,
         \u_a23_mem/p_mem[15][0] , \u_a23_mem/p_mem[15][1] ,
         \u_a23_mem/p_mem[15][2] , \u_a23_mem/p_mem[15][3] ,
         \u_a23_mem/p_mem[15][4] , \u_a23_mem/p_mem[15][5] ,
         \u_a23_mem/p_mem[15][6] , \u_a23_mem/p_mem[15][7] ,
         \u_a23_mem/p_mem[16][0] , \u_a23_mem/p_mem[16][1] ,
         \u_a23_mem/p_mem[16][2] , \u_a23_mem/p_mem[16][3] ,
         \u_a23_mem/p_mem[16][4] , \u_a23_mem/p_mem[16][5] ,
         \u_a23_mem/p_mem[16][6] , \u_a23_mem/p_mem[16][7] ,
         \u_a23_mem/p_mem[17][0] , \u_a23_mem/p_mem[17][1] ,
         \u_a23_mem/p_mem[17][2] , \u_a23_mem/p_mem[17][3] ,
         \u_a23_mem/p_mem[17][4] , \u_a23_mem/p_mem[17][5] ,
         \u_a23_mem/p_mem[17][6] , \u_a23_mem/p_mem[17][7] ,
         \u_a23_mem/p_mem[18][0] , \u_a23_mem/p_mem[18][1] ,
         \u_a23_mem/p_mem[18][2] , \u_a23_mem/p_mem[18][3] ,
         \u_a23_mem/p_mem[18][4] , \u_a23_mem/p_mem[18][5] ,
         \u_a23_mem/p_mem[18][6] , \u_a23_mem/p_mem[18][7] ,
         \u_a23_mem/p_mem[19][0] , \u_a23_mem/p_mem[19][1] ,
         \u_a23_mem/p_mem[19][2] , \u_a23_mem/p_mem[19][3] ,
         \u_a23_mem/p_mem[19][4] , \u_a23_mem/p_mem[19][5] ,
         \u_a23_mem/p_mem[19][6] , \u_a23_mem/p_mem[19][7] ,
         \u_a23_mem/p_mem[20][0] , \u_a23_mem/p_mem[20][1] ,
         \u_a23_mem/p_mem[20][2] , \u_a23_mem/p_mem[20][3] ,
         \u_a23_mem/p_mem[20][4] , \u_a23_mem/p_mem[20][5] ,
         \u_a23_mem/p_mem[20][6] , \u_a23_mem/p_mem[20][7] ,
         \u_a23_mem/p_mem[21][0] , \u_a23_mem/p_mem[21][1] ,
         \u_a23_mem/p_mem[21][2] , \u_a23_mem/p_mem[21][3] ,
         \u_a23_mem/p_mem[21][4] , \u_a23_mem/p_mem[21][5] ,
         \u_a23_mem/p_mem[21][6] , \u_a23_mem/p_mem[21][7] ,
         \u_a23_mem/p_mem[22][0] , \u_a23_mem/p_mem[22][1] ,
         \u_a23_mem/p_mem[22][2] , \u_a23_mem/p_mem[22][3] ,
         \u_a23_mem/p_mem[22][4] , \u_a23_mem/p_mem[22][5] ,
         \u_a23_mem/p_mem[22][6] , \u_a23_mem/p_mem[22][7] ,
         \u_a23_mem/p_mem[23][0] , \u_a23_mem/p_mem[23][1] ,
         \u_a23_mem/p_mem[23][2] , \u_a23_mem/p_mem[23][3] ,
         \u_a23_mem/p_mem[23][4] , \u_a23_mem/p_mem[23][5] ,
         \u_a23_mem/p_mem[23][6] , \u_a23_mem/p_mem[23][7] ,
         \u_a23_mem/p_mem[24][0] , \u_a23_mem/p_mem[24][1] ,
         \u_a23_mem/p_mem[24][2] , \u_a23_mem/p_mem[24][3] ,
         \u_a23_mem/p_mem[24][4] , \u_a23_mem/p_mem[24][5] ,
         \u_a23_mem/p_mem[24][6] , \u_a23_mem/p_mem[24][7] ,
         \u_a23_mem/p_mem[25][0] , \u_a23_mem/p_mem[25][1] ,
         \u_a23_mem/p_mem[25][2] , \u_a23_mem/p_mem[25][3] ,
         \u_a23_mem/p_mem[25][4] , \u_a23_mem/p_mem[25][5] ,
         \u_a23_mem/p_mem[25][6] , \u_a23_mem/p_mem[25][7] ,
         \u_a23_mem/p_mem[26][0] , \u_a23_mem/p_mem[26][1] ,
         \u_a23_mem/p_mem[26][2] , \u_a23_mem/p_mem[26][3] ,
         \u_a23_mem/p_mem[26][4] , \u_a23_mem/p_mem[26][5] ,
         \u_a23_mem/p_mem[26][6] , \u_a23_mem/p_mem[26][7] ,
         \u_a23_mem/p_mem[27][0] , \u_a23_mem/p_mem[27][1] ,
         \u_a23_mem/p_mem[27][2] , \u_a23_mem/p_mem[27][3] ,
         \u_a23_mem/p_mem[27][4] , \u_a23_mem/p_mem[27][5] ,
         \u_a23_mem/p_mem[27][6] , \u_a23_mem/p_mem[27][7] ,
         \u_a23_mem/p_mem[28][0] , \u_a23_mem/p_mem[28][1] ,
         \u_a23_mem/p_mem[28][2] , \u_a23_mem/p_mem[28][3] ,
         \u_a23_mem/p_mem[28][4] , \u_a23_mem/p_mem[28][5] ,
         \u_a23_mem/p_mem[28][6] , \u_a23_mem/p_mem[28][7] ,
         \u_a23_mem/p_mem[29][0] , \u_a23_mem/p_mem[29][1] ,
         \u_a23_mem/p_mem[29][2] , \u_a23_mem/p_mem[29][3] ,
         \u_a23_mem/p_mem[29][4] , \u_a23_mem/p_mem[29][5] ,
         \u_a23_mem/p_mem[29][6] , \u_a23_mem/p_mem[29][7] ,
         \u_a23_mem/p_mem[30][0] , \u_a23_mem/p_mem[30][1] ,
         \u_a23_mem/p_mem[30][2] , \u_a23_mem/p_mem[30][3] ,
         \u_a23_mem/p_mem[30][4] , \u_a23_mem/p_mem[30][5] ,
         \u_a23_mem/p_mem[30][6] , \u_a23_mem/p_mem[30][7] ,
         \u_a23_mem/p_mem[31][0] , \u_a23_mem/p_mem[31][1] ,
         \u_a23_mem/p_mem[31][2] , \u_a23_mem/p_mem[31][3] ,
         \u_a23_mem/p_mem[31][4] , \u_a23_mem/p_mem[31][5] ,
         \u_a23_mem/p_mem[31][6] , \u_a23_mem/p_mem[31][7] ,
         \u_a23_mem/p_mem[32][0] , \u_a23_mem/p_mem[32][1] ,
         \u_a23_mem/p_mem[32][2] , \u_a23_mem/p_mem[32][3] ,
         \u_a23_mem/p_mem[32][4] , \u_a23_mem/p_mem[32][5] ,
         \u_a23_mem/p_mem[32][6] , \u_a23_mem/p_mem[32][7] ,
         \u_a23_mem/p_mem[33][0] , \u_a23_mem/p_mem[33][1] ,
         \u_a23_mem/p_mem[33][2] , \u_a23_mem/p_mem[33][3] ,
         \u_a23_mem/p_mem[33][4] , \u_a23_mem/p_mem[33][5] ,
         \u_a23_mem/p_mem[33][6] , \u_a23_mem/p_mem[33][7] ,
         \u_a23_mem/p_mem[34][0] , \u_a23_mem/p_mem[34][1] ,
         \u_a23_mem/p_mem[34][2] , \u_a23_mem/p_mem[34][3] ,
         \u_a23_mem/p_mem[34][4] , \u_a23_mem/p_mem[34][5] ,
         \u_a23_mem/p_mem[34][6] , \u_a23_mem/p_mem[34][7] ,
         \u_a23_mem/p_mem[35][0] , \u_a23_mem/p_mem[35][1] ,
         \u_a23_mem/p_mem[35][2] , \u_a23_mem/p_mem[35][3] ,
         \u_a23_mem/p_mem[35][4] , \u_a23_mem/p_mem[35][5] ,
         \u_a23_mem/p_mem[35][6] , \u_a23_mem/p_mem[35][7] ,
         \u_a23_mem/p_mem[36][0] , \u_a23_mem/p_mem[36][1] ,
         \u_a23_mem/p_mem[36][2] , \u_a23_mem/p_mem[36][3] ,
         \u_a23_mem/p_mem[36][4] , \u_a23_mem/p_mem[36][5] ,
         \u_a23_mem/p_mem[36][6] , \u_a23_mem/p_mem[36][7] ,
         \u_a23_mem/p_mem[37][0] , \u_a23_mem/p_mem[37][1] ,
         \u_a23_mem/p_mem[37][2] , \u_a23_mem/p_mem[37][3] ,
         \u_a23_mem/p_mem[37][4] , \u_a23_mem/p_mem[37][5] ,
         \u_a23_mem/p_mem[37][6] , \u_a23_mem/p_mem[37][7] ,
         \u_a23_mem/p_mem[38][0] , \u_a23_mem/p_mem[38][1] ,
         \u_a23_mem/p_mem[38][2] , \u_a23_mem/p_mem[38][3] ,
         \u_a23_mem/p_mem[38][4] , \u_a23_mem/p_mem[38][5] ,
         \u_a23_mem/p_mem[38][6] , \u_a23_mem/p_mem[38][7] ,
         \u_a23_mem/p_mem[39][0] , \u_a23_mem/p_mem[39][1] ,
         \u_a23_mem/p_mem[39][2] , \u_a23_mem/p_mem[39][3] ,
         \u_a23_mem/p_mem[39][4] , \u_a23_mem/p_mem[39][5] ,
         \u_a23_mem/p_mem[39][6] , \u_a23_mem/p_mem[39][7] ,
         \u_a23_mem/p_mem[40][0] , \u_a23_mem/p_mem[40][1] ,
         \u_a23_mem/p_mem[40][2] , \u_a23_mem/p_mem[40][3] ,
         \u_a23_mem/p_mem[40][4] , \u_a23_mem/p_mem[40][5] ,
         \u_a23_mem/p_mem[40][6] , \u_a23_mem/p_mem[40][7] ,
         \u_a23_mem/p_mem[41][0] , \u_a23_mem/p_mem[41][1] ,
         \u_a23_mem/p_mem[41][2] , \u_a23_mem/p_mem[41][3] ,
         \u_a23_mem/p_mem[41][4] , \u_a23_mem/p_mem[41][5] ,
         \u_a23_mem/p_mem[41][6] , \u_a23_mem/p_mem[41][7] ,
         \u_a23_mem/p_mem[42][0] , \u_a23_mem/p_mem[42][1] ,
         \u_a23_mem/p_mem[42][2] , \u_a23_mem/p_mem[42][3] ,
         \u_a23_mem/p_mem[42][4] , \u_a23_mem/p_mem[42][5] ,
         \u_a23_mem/p_mem[42][6] , \u_a23_mem/p_mem[42][7] ,
         \u_a23_mem/p_mem[43][0] , \u_a23_mem/p_mem[43][1] ,
         \u_a23_mem/p_mem[43][2] , \u_a23_mem/p_mem[43][3] ,
         \u_a23_mem/p_mem[43][4] , \u_a23_mem/p_mem[43][5] ,
         \u_a23_mem/p_mem[43][6] , \u_a23_mem/p_mem[43][7] ,
         \u_a23_mem/p_mem[44][0] , \u_a23_mem/p_mem[44][1] ,
         \u_a23_mem/p_mem[44][2] , \u_a23_mem/p_mem[44][3] ,
         \u_a23_mem/p_mem[44][4] , \u_a23_mem/p_mem[44][5] ,
         \u_a23_mem/p_mem[44][6] , \u_a23_mem/p_mem[44][7] ,
         \u_a23_mem/p_mem[45][0] , \u_a23_mem/p_mem[45][1] ,
         \u_a23_mem/p_mem[45][2] , \u_a23_mem/p_mem[45][3] ,
         \u_a23_mem/p_mem[45][4] , \u_a23_mem/p_mem[45][5] ,
         \u_a23_mem/p_mem[45][6] , \u_a23_mem/p_mem[45][7] ,
         \u_a23_mem/p_mem[46][0] , \u_a23_mem/p_mem[46][1] ,
         \u_a23_mem/p_mem[46][2] , \u_a23_mem/p_mem[46][3] ,
         \u_a23_mem/p_mem[46][4] , \u_a23_mem/p_mem[46][5] ,
         \u_a23_mem/p_mem[46][6] , \u_a23_mem/p_mem[46][7] ,
         \u_a23_mem/p_mem[47][0] , \u_a23_mem/p_mem[47][1] ,
         \u_a23_mem/p_mem[47][2] , \u_a23_mem/p_mem[47][3] ,
         \u_a23_mem/p_mem[47][4] , \u_a23_mem/p_mem[47][5] ,
         \u_a23_mem/p_mem[47][6] , \u_a23_mem/p_mem[47][7] ,
         \u_a23_mem/p_mem[48][0] , \u_a23_mem/p_mem[48][1] ,
         \u_a23_mem/p_mem[48][2] , \u_a23_mem/p_mem[48][3] ,
         \u_a23_mem/p_mem[48][4] , \u_a23_mem/p_mem[48][5] ,
         \u_a23_mem/p_mem[48][6] , \u_a23_mem/p_mem[48][7] ,
         \u_a23_mem/p_mem[49][0] , \u_a23_mem/p_mem[49][1] ,
         \u_a23_mem/p_mem[49][2] , \u_a23_mem/p_mem[49][3] ,
         \u_a23_mem/p_mem[49][4] , \u_a23_mem/p_mem[49][5] ,
         \u_a23_mem/p_mem[49][6] , \u_a23_mem/p_mem[49][7] ,
         \u_a23_mem/p_mem[50][0] , \u_a23_mem/p_mem[50][1] ,
         \u_a23_mem/p_mem[50][2] , \u_a23_mem/p_mem[50][3] ,
         \u_a23_mem/p_mem[50][4] , \u_a23_mem/p_mem[50][5] ,
         \u_a23_mem/p_mem[50][6] , \u_a23_mem/p_mem[50][7] ,
         \u_a23_mem/p_mem[51][0] , \u_a23_mem/p_mem[51][1] ,
         \u_a23_mem/p_mem[51][2] , \u_a23_mem/p_mem[51][3] ,
         \u_a23_mem/p_mem[51][4] , \u_a23_mem/p_mem[51][5] ,
         \u_a23_mem/p_mem[51][6] , \u_a23_mem/p_mem[51][7] ,
         \u_a23_mem/p_mem[52][0] , \u_a23_mem/p_mem[52][1] ,
         \u_a23_mem/p_mem[52][2] , \u_a23_mem/p_mem[52][3] ,
         \u_a23_mem/p_mem[52][4] , \u_a23_mem/p_mem[52][5] ,
         \u_a23_mem/p_mem[52][6] , \u_a23_mem/p_mem[52][7] ,
         \u_a23_mem/p_mem[53][0] , \u_a23_mem/p_mem[53][1] ,
         \u_a23_mem/p_mem[53][2] , \u_a23_mem/p_mem[53][3] ,
         \u_a23_mem/p_mem[53][4] , \u_a23_mem/p_mem[53][5] ,
         \u_a23_mem/p_mem[53][6] , \u_a23_mem/p_mem[53][7] ,
         \u_a23_mem/p_mem[54][0] , \u_a23_mem/p_mem[54][1] ,
         \u_a23_mem/p_mem[54][2] , \u_a23_mem/p_mem[54][3] ,
         \u_a23_mem/p_mem[54][4] , \u_a23_mem/p_mem[54][5] ,
         \u_a23_mem/p_mem[54][6] , \u_a23_mem/p_mem[54][7] ,
         \u_a23_mem/p_mem[55][0] , \u_a23_mem/p_mem[55][1] ,
         \u_a23_mem/p_mem[55][2] , \u_a23_mem/p_mem[55][3] ,
         \u_a23_mem/p_mem[55][4] , \u_a23_mem/p_mem[55][5] ,
         \u_a23_mem/p_mem[55][6] , \u_a23_mem/p_mem[55][7] ,
         \u_a23_mem/p_mem[56][0] , \u_a23_mem/p_mem[56][1] ,
         \u_a23_mem/p_mem[56][2] , \u_a23_mem/p_mem[56][3] ,
         \u_a23_mem/p_mem[56][4] , \u_a23_mem/p_mem[56][5] ,
         \u_a23_mem/p_mem[56][6] , \u_a23_mem/p_mem[56][7] ,
         \u_a23_mem/p_mem[57][0] , \u_a23_mem/p_mem[57][1] ,
         \u_a23_mem/p_mem[57][2] , \u_a23_mem/p_mem[57][3] ,
         \u_a23_mem/p_mem[57][4] , \u_a23_mem/p_mem[57][5] ,
         \u_a23_mem/p_mem[57][6] , \u_a23_mem/p_mem[57][7] ,
         \u_a23_mem/p_mem[58][0] , \u_a23_mem/p_mem[58][1] ,
         \u_a23_mem/p_mem[58][2] , \u_a23_mem/p_mem[58][3] ,
         \u_a23_mem/p_mem[58][4] , \u_a23_mem/p_mem[58][5] ,
         \u_a23_mem/p_mem[58][6] , \u_a23_mem/p_mem[58][7] ,
         \u_a23_mem/p_mem[59][0] , \u_a23_mem/p_mem[59][1] ,
         \u_a23_mem/p_mem[59][2] , \u_a23_mem/p_mem[59][3] ,
         \u_a23_mem/p_mem[59][4] , \u_a23_mem/p_mem[59][5] ,
         \u_a23_mem/p_mem[59][6] , \u_a23_mem/p_mem[59][7] ,
         \u_a23_mem/p_mem[60][0] , \u_a23_mem/p_mem[60][1] ,
         \u_a23_mem/p_mem[60][2] , \u_a23_mem/p_mem[60][3] ,
         \u_a23_mem/p_mem[60][4] , \u_a23_mem/p_mem[60][5] ,
         \u_a23_mem/p_mem[60][6] , \u_a23_mem/p_mem[60][7] ,
         \u_a23_mem/p_mem[61][0] , \u_a23_mem/p_mem[61][1] ,
         \u_a23_mem/p_mem[61][2] , \u_a23_mem/p_mem[61][3] ,
         \u_a23_mem/p_mem[61][4] , \u_a23_mem/p_mem[61][5] ,
         \u_a23_mem/p_mem[61][6] , \u_a23_mem/p_mem[61][7] ,
         \u_a23_mem/p_mem[62][0] , \u_a23_mem/p_mem[62][1] ,
         \u_a23_mem/p_mem[62][2] , \u_a23_mem/p_mem[62][3] ,
         \u_a23_mem/p_mem[62][4] , \u_a23_mem/p_mem[62][5] ,
         \u_a23_mem/p_mem[62][6] , \u_a23_mem/p_mem[62][7] ,
         \u_a23_mem/p_mem[63][0] , \u_a23_mem/p_mem[63][1] ,
         \u_a23_mem/p_mem[63][2] , \u_a23_mem/p_mem[63][3] ,
         \u_a23_mem/p_mem[63][4] , \u_a23_mem/p_mem[63][5] ,
         \u_a23_mem/p_mem[63][6] , \u_a23_mem/p_mem[63][7] ,
         \u_a23_mem/p_mem[64][0] , \u_a23_mem/p_mem[64][1] ,
         \u_a23_mem/p_mem[64][2] , \u_a23_mem/p_mem[64][3] ,
         \u_a23_mem/p_mem[64][4] , \u_a23_mem/p_mem[64][5] ,
         \u_a23_mem/p_mem[64][6] , \u_a23_mem/p_mem[64][7] ,
         \u_a23_mem/p_mem[65][0] , \u_a23_mem/p_mem[65][1] ,
         \u_a23_mem/p_mem[65][2] , \u_a23_mem/p_mem[65][3] ,
         \u_a23_mem/p_mem[65][4] , \u_a23_mem/p_mem[65][5] ,
         \u_a23_mem/p_mem[65][6] , \u_a23_mem/p_mem[65][7] ,
         \u_a23_mem/p_mem[66][0] , \u_a23_mem/p_mem[66][1] ,
         \u_a23_mem/p_mem[66][2] , \u_a23_mem/p_mem[66][3] ,
         \u_a23_mem/p_mem[66][4] , \u_a23_mem/p_mem[66][5] ,
         \u_a23_mem/p_mem[66][6] , \u_a23_mem/p_mem[66][7] ,
         \u_a23_mem/p_mem[67][0] , \u_a23_mem/p_mem[67][1] ,
         \u_a23_mem/p_mem[67][2] , \u_a23_mem/p_mem[67][3] ,
         \u_a23_mem/p_mem[67][4] , \u_a23_mem/p_mem[67][5] ,
         \u_a23_mem/p_mem[67][6] , \u_a23_mem/p_mem[67][7] ,
         \u_a23_mem/p_mem[68][0] , \u_a23_mem/p_mem[68][1] ,
         \u_a23_mem/p_mem[68][2] , \u_a23_mem/p_mem[68][3] ,
         \u_a23_mem/p_mem[68][4] , \u_a23_mem/p_mem[68][5] ,
         \u_a23_mem/p_mem[68][6] , \u_a23_mem/p_mem[68][7] ,
         \u_a23_mem/p_mem[69][0] , \u_a23_mem/p_mem[69][1] ,
         \u_a23_mem/p_mem[69][2] , \u_a23_mem/p_mem[69][3] ,
         \u_a23_mem/p_mem[69][4] , \u_a23_mem/p_mem[69][5] ,
         \u_a23_mem/p_mem[69][6] , \u_a23_mem/p_mem[69][7] ,
         \u_a23_mem/p_mem[70][0] , \u_a23_mem/p_mem[70][1] ,
         \u_a23_mem/p_mem[70][2] , \u_a23_mem/p_mem[70][3] ,
         \u_a23_mem/p_mem[70][4] , \u_a23_mem/p_mem[70][5] ,
         \u_a23_mem/p_mem[70][6] , \u_a23_mem/p_mem[70][7] ,
         \u_a23_mem/p_mem[71][0] , \u_a23_mem/p_mem[71][1] ,
         \u_a23_mem/p_mem[71][2] , \u_a23_mem/p_mem[71][3] ,
         \u_a23_mem/p_mem[71][4] , \u_a23_mem/p_mem[71][5] ,
         \u_a23_mem/p_mem[71][6] , \u_a23_mem/p_mem[71][7] ,
         \u_a23_mem/p_mem[72][0] , \u_a23_mem/p_mem[72][1] ,
         \u_a23_mem/p_mem[72][2] , \u_a23_mem/p_mem[72][3] ,
         \u_a23_mem/p_mem[72][4] , \u_a23_mem/p_mem[72][5] ,
         \u_a23_mem/p_mem[72][6] , \u_a23_mem/p_mem[72][7] ,
         \u_a23_mem/p_mem[73][0] , \u_a23_mem/p_mem[73][1] ,
         \u_a23_mem/p_mem[73][2] , \u_a23_mem/p_mem[73][3] ,
         \u_a23_mem/p_mem[73][4] , \u_a23_mem/p_mem[73][5] ,
         \u_a23_mem/p_mem[73][6] , \u_a23_mem/p_mem[73][7] ,
         \u_a23_mem/p_mem[74][0] , \u_a23_mem/p_mem[74][1] ,
         \u_a23_mem/p_mem[74][2] , \u_a23_mem/p_mem[74][3] ,
         \u_a23_mem/p_mem[74][4] , \u_a23_mem/p_mem[74][5] ,
         \u_a23_mem/p_mem[74][6] , \u_a23_mem/p_mem[74][7] ,
         \u_a23_mem/p_mem[75][0] , \u_a23_mem/p_mem[75][1] ,
         \u_a23_mem/p_mem[75][2] , \u_a23_mem/p_mem[75][3] ,
         \u_a23_mem/p_mem[75][4] , \u_a23_mem/p_mem[75][5] ,
         \u_a23_mem/p_mem[75][6] , \u_a23_mem/p_mem[75][7] ,
         \u_a23_mem/p_mem[76][0] , \u_a23_mem/p_mem[76][1] ,
         \u_a23_mem/p_mem[76][2] , \u_a23_mem/p_mem[76][3] ,
         \u_a23_mem/p_mem[76][4] , \u_a23_mem/p_mem[76][5] ,
         \u_a23_mem/p_mem[76][6] , \u_a23_mem/p_mem[76][7] ,
         \u_a23_mem/p_mem[77][0] , \u_a23_mem/p_mem[77][1] ,
         \u_a23_mem/p_mem[77][2] , \u_a23_mem/p_mem[77][3] ,
         \u_a23_mem/p_mem[77][4] , \u_a23_mem/p_mem[77][5] ,
         \u_a23_mem/p_mem[77][6] , \u_a23_mem/p_mem[77][7] ,
         \u_a23_mem/p_mem[78][0] , \u_a23_mem/p_mem[78][1] ,
         \u_a23_mem/p_mem[78][2] , \u_a23_mem/p_mem[78][3] ,
         \u_a23_mem/p_mem[78][4] , \u_a23_mem/p_mem[78][5] ,
         \u_a23_mem/p_mem[78][6] , \u_a23_mem/p_mem[78][7] ,
         \u_a23_mem/p_mem[79][0] , \u_a23_mem/p_mem[79][1] ,
         \u_a23_mem/p_mem[79][2] , \u_a23_mem/p_mem[79][3] ,
         \u_a23_mem/p_mem[79][4] , \u_a23_mem/p_mem[79][5] ,
         \u_a23_mem/p_mem[79][6] , \u_a23_mem/p_mem[79][7] ,
         \u_a23_mem/p_mem[80][0] , \u_a23_mem/p_mem[80][1] ,
         \u_a23_mem/p_mem[80][2] , \u_a23_mem/p_mem[80][3] ,
         \u_a23_mem/p_mem[80][4] , \u_a23_mem/p_mem[80][5] ,
         \u_a23_mem/p_mem[80][6] , \u_a23_mem/p_mem[80][7] ,
         \u_a23_mem/p_mem[81][0] , \u_a23_mem/p_mem[81][1] ,
         \u_a23_mem/p_mem[81][2] , \u_a23_mem/p_mem[81][3] ,
         \u_a23_mem/p_mem[81][4] , \u_a23_mem/p_mem[81][5] ,
         \u_a23_mem/p_mem[81][6] , \u_a23_mem/p_mem[81][7] ,
         \u_a23_mem/p_mem[82][0] , \u_a23_mem/p_mem[82][1] ,
         \u_a23_mem/p_mem[82][2] , \u_a23_mem/p_mem[82][3] ,
         \u_a23_mem/p_mem[82][4] , \u_a23_mem/p_mem[82][5] ,
         \u_a23_mem/p_mem[82][6] , \u_a23_mem/p_mem[82][7] ,
         \u_a23_mem/p_mem[83][0] , \u_a23_mem/p_mem[83][1] ,
         \u_a23_mem/p_mem[83][2] , \u_a23_mem/p_mem[83][3] ,
         \u_a23_mem/p_mem[83][4] , \u_a23_mem/p_mem[83][5] ,
         \u_a23_mem/p_mem[83][6] , \u_a23_mem/p_mem[83][7] ,
         \u_a23_mem/p_mem[84][0] , \u_a23_mem/p_mem[84][1] ,
         \u_a23_mem/p_mem[84][2] , \u_a23_mem/p_mem[84][3] ,
         \u_a23_mem/p_mem[84][4] , \u_a23_mem/p_mem[84][5] ,
         \u_a23_mem/p_mem[84][6] , \u_a23_mem/p_mem[84][7] ,
         \u_a23_mem/p_mem[85][0] , \u_a23_mem/p_mem[85][1] ,
         \u_a23_mem/p_mem[85][2] , \u_a23_mem/p_mem[85][3] ,
         \u_a23_mem/p_mem[85][4] , \u_a23_mem/p_mem[85][5] ,
         \u_a23_mem/p_mem[85][6] , \u_a23_mem/p_mem[85][7] ,
         \u_a23_mem/p_mem[86][0] , \u_a23_mem/p_mem[86][1] ,
         \u_a23_mem/p_mem[86][2] , \u_a23_mem/p_mem[86][3] ,
         \u_a23_mem/p_mem[86][4] , \u_a23_mem/p_mem[86][5] ,
         \u_a23_mem/p_mem[86][6] , \u_a23_mem/p_mem[86][7] ,
         \u_a23_mem/p_mem[87][0] , \u_a23_mem/p_mem[87][1] ,
         \u_a23_mem/p_mem[87][2] , \u_a23_mem/p_mem[87][3] ,
         \u_a23_mem/p_mem[87][4] , \u_a23_mem/p_mem[87][5] ,
         \u_a23_mem/p_mem[87][6] , \u_a23_mem/p_mem[87][7] ,
         \u_a23_mem/p_mem[88][0] , \u_a23_mem/p_mem[88][1] ,
         \u_a23_mem/p_mem[88][2] , \u_a23_mem/p_mem[88][3] ,
         \u_a23_mem/p_mem[88][4] , \u_a23_mem/p_mem[88][5] ,
         \u_a23_mem/p_mem[88][6] , \u_a23_mem/p_mem[88][7] ,
         \u_a23_mem/p_mem[89][0] , \u_a23_mem/p_mem[89][1] ,
         \u_a23_mem/p_mem[89][2] , \u_a23_mem/p_mem[89][3] ,
         \u_a23_mem/p_mem[89][4] , \u_a23_mem/p_mem[89][5] ,
         \u_a23_mem/p_mem[89][6] , \u_a23_mem/p_mem[89][7] ,
         \u_a23_mem/p_mem[90][0] , \u_a23_mem/p_mem[90][1] ,
         \u_a23_mem/p_mem[90][2] , \u_a23_mem/p_mem[90][3] ,
         \u_a23_mem/p_mem[90][4] , \u_a23_mem/p_mem[90][5] ,
         \u_a23_mem/p_mem[90][6] , \u_a23_mem/p_mem[90][7] ,
         \u_a23_mem/p_mem[91][0] , \u_a23_mem/p_mem[91][1] ,
         \u_a23_mem/p_mem[91][2] , \u_a23_mem/p_mem[91][3] ,
         \u_a23_mem/p_mem[91][4] , \u_a23_mem/p_mem[91][5] ,
         \u_a23_mem/p_mem[91][6] , \u_a23_mem/p_mem[91][7] ,
         \u_a23_mem/p_mem[92][0] , \u_a23_mem/p_mem[92][1] ,
         \u_a23_mem/p_mem[92][2] , \u_a23_mem/p_mem[92][3] ,
         \u_a23_mem/p_mem[92][4] , \u_a23_mem/p_mem[92][5] ,
         \u_a23_mem/p_mem[92][6] , \u_a23_mem/p_mem[92][7] ,
         \u_a23_mem/p_mem[93][0] , \u_a23_mem/p_mem[93][1] ,
         \u_a23_mem/p_mem[93][2] , \u_a23_mem/p_mem[93][3] ,
         \u_a23_mem/p_mem[93][4] , \u_a23_mem/p_mem[93][5] ,
         \u_a23_mem/p_mem[93][6] , \u_a23_mem/p_mem[93][7] ,
         \u_a23_mem/p_mem[94][0] , \u_a23_mem/p_mem[94][1] ,
         \u_a23_mem/p_mem[94][2] , \u_a23_mem/p_mem[94][3] ,
         \u_a23_mem/p_mem[94][4] , \u_a23_mem/p_mem[94][5] ,
         \u_a23_mem/p_mem[94][6] , \u_a23_mem/p_mem[94][7] ,
         \u_a23_mem/p_mem[95][0] , \u_a23_mem/p_mem[95][1] ,
         \u_a23_mem/p_mem[95][2] , \u_a23_mem/p_mem[95][3] ,
         \u_a23_mem/p_mem[95][4] , \u_a23_mem/p_mem[95][5] ,
         \u_a23_mem/p_mem[95][6] , \u_a23_mem/p_mem[95][7] ,
         \u_a23_mem/p_mem[96][0] , \u_a23_mem/p_mem[96][1] ,
         \u_a23_mem/p_mem[96][2] , \u_a23_mem/p_mem[96][3] ,
         \u_a23_mem/p_mem[96][4] , \u_a23_mem/p_mem[96][5] ,
         \u_a23_mem/p_mem[96][6] , \u_a23_mem/p_mem[96][7] ,
         \u_a23_mem/p_mem[97][0] , \u_a23_mem/p_mem[97][1] ,
         \u_a23_mem/p_mem[97][2] , \u_a23_mem/p_mem[97][3] ,
         \u_a23_mem/p_mem[97][4] , \u_a23_mem/p_mem[97][5] ,
         \u_a23_mem/p_mem[97][6] , \u_a23_mem/p_mem[97][7] ,
         \u_a23_mem/p_mem[98][0] , \u_a23_mem/p_mem[98][1] ,
         \u_a23_mem/p_mem[98][2] , \u_a23_mem/p_mem[98][3] ,
         \u_a23_mem/p_mem[98][4] , \u_a23_mem/p_mem[98][5] ,
         \u_a23_mem/p_mem[98][6] , \u_a23_mem/p_mem[98][7] ,
         \u_a23_mem/p_mem[99][0] , \u_a23_mem/p_mem[99][1] ,
         \u_a23_mem/p_mem[99][2] , \u_a23_mem/p_mem[99][3] ,
         \u_a23_mem/p_mem[99][4] , \u_a23_mem/p_mem[99][5] ,
         \u_a23_mem/p_mem[99][6] , \u_a23_mem/p_mem[99][7] ,
         \u_a23_mem/p_mem[100][0] , \u_a23_mem/p_mem[100][1] ,
         \u_a23_mem/p_mem[100][2] , \u_a23_mem/p_mem[100][3] ,
         \u_a23_mem/p_mem[100][4] , \u_a23_mem/p_mem[100][5] ,
         \u_a23_mem/p_mem[100][6] , \u_a23_mem/p_mem[100][7] ,
         \u_a23_mem/p_mem[101][0] , \u_a23_mem/p_mem[101][1] ,
         \u_a23_mem/p_mem[101][2] , \u_a23_mem/p_mem[101][3] ,
         \u_a23_mem/p_mem[101][4] , \u_a23_mem/p_mem[101][5] ,
         \u_a23_mem/p_mem[101][6] , \u_a23_mem/p_mem[101][7] ,
         \u_a23_mem/p_mem[102][0] , \u_a23_mem/p_mem[102][1] ,
         \u_a23_mem/p_mem[102][2] , \u_a23_mem/p_mem[102][3] ,
         \u_a23_mem/p_mem[102][4] , \u_a23_mem/p_mem[102][5] ,
         \u_a23_mem/p_mem[102][6] , \u_a23_mem/p_mem[102][7] ,
         \u_a23_mem/p_mem[103][0] , \u_a23_mem/p_mem[103][1] ,
         \u_a23_mem/p_mem[103][2] , \u_a23_mem/p_mem[103][3] ,
         \u_a23_mem/p_mem[103][4] , \u_a23_mem/p_mem[103][5] ,
         \u_a23_mem/p_mem[103][6] , \u_a23_mem/p_mem[103][7] ,
         \u_a23_mem/p_mem[104][0] , \u_a23_mem/p_mem[104][1] ,
         \u_a23_mem/p_mem[104][2] , \u_a23_mem/p_mem[104][3] ,
         \u_a23_mem/p_mem[104][4] , \u_a23_mem/p_mem[104][5] ,
         \u_a23_mem/p_mem[104][6] , \u_a23_mem/p_mem[104][7] ,
         \u_a23_mem/p_mem[105][0] , \u_a23_mem/p_mem[105][1] ,
         \u_a23_mem/p_mem[105][2] , \u_a23_mem/p_mem[105][3] ,
         \u_a23_mem/p_mem[105][4] , \u_a23_mem/p_mem[105][5] ,
         \u_a23_mem/p_mem[105][6] , \u_a23_mem/p_mem[105][7] ,
         \u_a23_mem/p_mem[106][0] , \u_a23_mem/p_mem[106][1] ,
         \u_a23_mem/p_mem[106][2] , \u_a23_mem/p_mem[106][3] ,
         \u_a23_mem/p_mem[106][4] , \u_a23_mem/p_mem[106][5] ,
         \u_a23_mem/p_mem[106][6] , \u_a23_mem/p_mem[106][7] ,
         \u_a23_mem/p_mem[107][0] , \u_a23_mem/p_mem[107][1] ,
         \u_a23_mem/p_mem[107][2] , \u_a23_mem/p_mem[107][3] ,
         \u_a23_mem/p_mem[107][4] , \u_a23_mem/p_mem[107][5] ,
         \u_a23_mem/p_mem[107][6] , \u_a23_mem/p_mem[107][7] ,
         \u_a23_mem/p_mem[108][0] , \u_a23_mem/p_mem[108][1] ,
         \u_a23_mem/p_mem[108][2] , \u_a23_mem/p_mem[108][3] ,
         \u_a23_mem/p_mem[108][4] , \u_a23_mem/p_mem[108][5] ,
         \u_a23_mem/p_mem[108][6] , \u_a23_mem/p_mem[108][7] ,
         \u_a23_mem/p_mem[109][0] , \u_a23_mem/p_mem[109][1] ,
         \u_a23_mem/p_mem[109][2] , \u_a23_mem/p_mem[109][3] ,
         \u_a23_mem/p_mem[109][4] , \u_a23_mem/p_mem[109][5] ,
         \u_a23_mem/p_mem[109][6] , \u_a23_mem/p_mem[109][7] ,
         \u_a23_mem/p_mem[110][0] , \u_a23_mem/p_mem[110][1] ,
         \u_a23_mem/p_mem[110][2] , \u_a23_mem/p_mem[110][3] ,
         \u_a23_mem/p_mem[110][4] , \u_a23_mem/p_mem[110][5] ,
         \u_a23_mem/p_mem[110][6] , \u_a23_mem/p_mem[110][7] ,
         \u_a23_mem/p_mem[111][0] , \u_a23_mem/p_mem[111][1] ,
         \u_a23_mem/p_mem[111][2] , \u_a23_mem/p_mem[111][3] ,
         \u_a23_mem/p_mem[111][4] , \u_a23_mem/p_mem[111][5] ,
         \u_a23_mem/p_mem[111][6] , \u_a23_mem/p_mem[111][7] ,
         \u_a23_mem/p_mem[112][0] , \u_a23_mem/p_mem[112][1] ,
         \u_a23_mem/p_mem[112][2] , \u_a23_mem/p_mem[112][3] ,
         \u_a23_mem/p_mem[112][4] , \u_a23_mem/p_mem[112][5] ,
         \u_a23_mem/p_mem[112][6] , \u_a23_mem/p_mem[112][7] ,
         \u_a23_mem/p_mem[113][0] , \u_a23_mem/p_mem[113][1] ,
         \u_a23_mem/p_mem[113][2] , \u_a23_mem/p_mem[113][3] ,
         \u_a23_mem/p_mem[113][4] , \u_a23_mem/p_mem[113][5] ,
         \u_a23_mem/p_mem[113][6] , \u_a23_mem/p_mem[113][7] ,
         \u_a23_mem/p_mem[114][0] , \u_a23_mem/p_mem[114][1] ,
         \u_a23_mem/p_mem[114][2] , \u_a23_mem/p_mem[114][3] ,
         \u_a23_mem/p_mem[114][4] , \u_a23_mem/p_mem[114][5] ,
         \u_a23_mem/p_mem[114][6] , \u_a23_mem/p_mem[114][7] ,
         \u_a23_mem/p_mem[115][0] , \u_a23_mem/p_mem[115][1] ,
         \u_a23_mem/p_mem[115][2] , \u_a23_mem/p_mem[115][3] ,
         \u_a23_mem/p_mem[115][4] , \u_a23_mem/p_mem[115][5] ,
         \u_a23_mem/p_mem[115][6] , \u_a23_mem/p_mem[115][7] ,
         \u_a23_mem/p_mem[116][0] , \u_a23_mem/p_mem[116][1] ,
         \u_a23_mem/p_mem[116][2] , \u_a23_mem/p_mem[116][3] ,
         \u_a23_mem/p_mem[116][4] , \u_a23_mem/p_mem[116][5] ,
         \u_a23_mem/p_mem[116][6] , \u_a23_mem/p_mem[116][7] ,
         \u_a23_mem/p_mem[117][0] , \u_a23_mem/p_mem[117][1] ,
         \u_a23_mem/p_mem[117][2] , \u_a23_mem/p_mem[117][3] ,
         \u_a23_mem/p_mem[117][4] , \u_a23_mem/p_mem[117][5] ,
         \u_a23_mem/p_mem[117][6] , \u_a23_mem/p_mem[117][7] ,
         \u_a23_mem/p_mem[118][0] , \u_a23_mem/p_mem[118][1] ,
         \u_a23_mem/p_mem[118][2] , \u_a23_mem/p_mem[118][3] ,
         \u_a23_mem/p_mem[118][4] , \u_a23_mem/p_mem[118][5] ,
         \u_a23_mem/p_mem[118][6] , \u_a23_mem/p_mem[118][7] ,
         \u_a23_mem/p_mem[119][0] , \u_a23_mem/p_mem[119][1] ,
         \u_a23_mem/p_mem[119][2] , \u_a23_mem/p_mem[119][3] ,
         \u_a23_mem/p_mem[119][4] , \u_a23_mem/p_mem[119][5] ,
         \u_a23_mem/p_mem[119][6] , \u_a23_mem/p_mem[119][7] ,
         \u_a23_mem/p_mem[120][0] , \u_a23_mem/p_mem[120][1] ,
         \u_a23_mem/p_mem[120][2] , \u_a23_mem/p_mem[120][3] ,
         \u_a23_mem/p_mem[120][4] , \u_a23_mem/p_mem[120][5] ,
         \u_a23_mem/p_mem[120][6] , \u_a23_mem/p_mem[120][7] ,
         \u_a23_mem/p_mem[121][0] , \u_a23_mem/p_mem[121][1] ,
         \u_a23_mem/p_mem[121][2] , \u_a23_mem/p_mem[121][3] ,
         \u_a23_mem/p_mem[121][4] , \u_a23_mem/p_mem[121][5] ,
         \u_a23_mem/p_mem[121][6] , \u_a23_mem/p_mem[121][7] ,
         \u_a23_mem/p_mem[122][0] , \u_a23_mem/p_mem[122][1] ,
         \u_a23_mem/p_mem[122][2] , \u_a23_mem/p_mem[122][3] ,
         \u_a23_mem/p_mem[122][4] , \u_a23_mem/p_mem[122][5] ,
         \u_a23_mem/p_mem[122][6] , \u_a23_mem/p_mem[122][7] ,
         \u_a23_mem/p_mem[123][0] , \u_a23_mem/p_mem[123][1] ,
         \u_a23_mem/p_mem[123][2] , \u_a23_mem/p_mem[123][3] ,
         \u_a23_mem/p_mem[123][4] , \u_a23_mem/p_mem[123][5] ,
         \u_a23_mem/p_mem[123][6] , \u_a23_mem/p_mem[123][7] ,
         \u_a23_mem/p_mem[124][0] , \u_a23_mem/p_mem[124][1] ,
         \u_a23_mem/p_mem[124][2] , \u_a23_mem/p_mem[124][3] ,
         \u_a23_mem/p_mem[124][4] , \u_a23_mem/p_mem[124][5] ,
         \u_a23_mem/p_mem[124][6] , \u_a23_mem/p_mem[124][7] ,
         \u_a23_mem/p_mem[125][0] , \u_a23_mem/p_mem[125][1] ,
         \u_a23_mem/p_mem[125][2] , \u_a23_mem/p_mem[125][3] ,
         \u_a23_mem/p_mem[125][4] , \u_a23_mem/p_mem[125][5] ,
         \u_a23_mem/p_mem[125][6] , \u_a23_mem/p_mem[125][7] ,
         \u_a23_mem/p_mem[126][0] , \u_a23_mem/p_mem[126][1] ,
         \u_a23_mem/p_mem[126][2] , \u_a23_mem/p_mem[126][3] ,
         \u_a23_mem/p_mem[126][4] , \u_a23_mem/p_mem[126][5] ,
         \u_a23_mem/p_mem[126][6] , \u_a23_mem/p_mem[126][7] ,
         \u_a23_mem/p_mem[127][0] , \u_a23_mem/p_mem[127][1] ,
         \u_a23_mem/p_mem[127][2] , \u_a23_mem/p_mem[127][3] ,
         \u_a23_mem/p_mem[127][4] , \u_a23_mem/p_mem[127][5] ,
         \u_a23_mem/p_mem[127][6] , \u_a23_mem/p_mem[127][7] ,
         \u_a23_core/u_decode/n1511 , \u_a23_core/u_decode/n1510 ,
         \u_a23_core/u_decode/n1509 , \u_a23_core/u_decode/n1508 ,
         \u_a23_core/u_decode/n1507 , \u_a23_core/u_decode/n1506 ,
         \u_a23_core/u_decode/n1505 , \u_a23_core/u_decode/n1504 ,
         \u_a23_core/u_decode/n1503 , \u_a23_core/u_decode/n1502 ,
         \u_a23_core/u_decode/n1501 , \u_a23_core/u_decode/n1500 ,
         \u_a23_core/u_decode/n1499 , \u_a23_core/u_decode/n1498 ,
         \u_a23_core/u_decode/n1495 , \u_a23_core/u_decode/n1494 ,
         \u_a23_core/u_decode/n1493 , \u_a23_core/u_decode/n1492 ,
         \u_a23_core/u_decode/n1491 , \u_a23_core/u_decode/n1490 ,
         \u_a23_core/u_decode/n1489 , \u_a23_core/u_decode/n1488 ,
         \u_a23_core/u_decode/n1487 , \u_a23_core/u_decode/n1486 ,
         \u_a23_core/u_decode/n1485 , \u_a23_core/u_decode/n1484 ,
         \u_a23_core/u_decode/n1483 , \u_a23_core/u_decode/n1482 ,
         \u_a23_core/u_decode/n1481 , \u_a23_core/u_decode/n1480 ,
         \u_a23_core/u_decode/n1479 , \u_a23_core/u_decode/n1478 ,
         \u_a23_core/u_decode/n1477 , \u_a23_core/u_decode/n1476 ,
         \u_a23_core/u_decode/n1475 , \u_a23_core/u_decode/n1474 ,
         \u_a23_core/u_decode/n1473 , \u_a23_core/u_decode/n1472 ,
         \u_a23_core/u_decode/n1471 , \u_a23_core/u_decode/n1470 ,
         \u_a23_core/u_decode/n1469 , \u_a23_core/u_decode/n1468 ,
         \u_a23_core/u_decode/n1467 , \u_a23_core/u_decode/n1466 ,
         \u_a23_core/u_decode/n1465 , \u_a23_core/u_decode/n1464 ,
         \u_a23_core/u_decode/n1463 , \u_a23_core/u_decode/n1462 ,
         \u_a23_core/u_decode/n1461 , \u_a23_core/u_decode/n1460 ,
         \u_a23_core/u_decode/n1459 , \u_a23_core/u_decode/n1458 ,
         \u_a23_core/u_decode/n1457 , \u_a23_core/u_decode/n1456 ,
         \u_a23_core/u_decode/n1455 , \u_a23_core/u_decode/n1454 ,
         \u_a23_core/u_decode/n1453 , \u_a23_core/u_decode/n1452 ,
         \u_a23_core/u_decode/n1451 , \u_a23_core/u_decode/n1450 ,
         \u_a23_core/u_decode/n1449 , \u_a23_core/u_decode/n1448 ,
         \u_a23_core/u_decode/n1447 , \u_a23_core/u_decode/n1446 ,
         \u_a23_core/u_decode/n1445 , \u_a23_core/u_decode/n1444 ,
         \u_a23_core/u_decode/n1443 , \u_a23_core/u_decode/n1442 ,
         \u_a23_core/u_decode/n1441 , \u_a23_core/u_decode/n1440 ,
         \u_a23_core/u_decode/n1439 , \u_a23_core/u_decode/n1438 ,
         \u_a23_core/u_decode/n1437 , \u_a23_core/u_decode/n1436 ,
         \u_a23_core/u_decode/n1435 , \u_a23_core/u_decode/n1434 ,
         \u_a23_core/u_decode/n1433 , \u_a23_core/u_decode/n1431 ,
         \u_a23_core/u_decode/n1429 , \u_a23_core/u_decode/n1427 ,
         \u_a23_core/u_decode/N1089 , \u_a23_core/u_decode/mtrans_reg_d1[3] ,
         \u_a23_core/u_decode/mtrans_reg_d1[2] ,
         \u_a23_core/u_decode/mtrans_reg_d1[1] ,
         \u_a23_core/u_decode/mtrans_reg_d1[0] ,
         \u_a23_core/u_decode/control_state_nxt[4] ,
         \u_a23_core/u_decode/control_state_nxt[3] ,
         \u_a23_core/u_decode/control_state_nxt[2] ,
         \u_a23_core/u_decode/control_state_nxt[1] ,
         \u_a23_core/u_decode/control_state_nxt[0] ,
         \u_a23_core/u_decode/status_bits_flags_wen_nxt ,
         \u_a23_core/u_decode/write_data_wen_nxt ,
         \u_a23_core/u_decode/reg_write_sel_nxt[0] ,
         \u_a23_core/u_decode/status_bits_sel_nxt_0 ,
         \u_a23_core/u_decode/status_bits_sel_nxt[2] ,
         \u_a23_core/u_decode/byte_enable_sel_nxt[0] ,
         \u_a23_core/u_decode/address_sel_nxt[2] ,
         \u_a23_core/u_decode/address_sel_nxt[1] ,
         \u_a23_core/u_decode/address_sel_nxt[0] ,
         \u_a23_core/u_decode/use_carry_in_nxt ,
         \u_a23_core/u_decode/barrel_shift_function_nxt[1] ,
         \u_a23_core/u_decode/barrel_shift_function_nxt[0] ,
         \u_a23_core/u_decode/barrel_shift_data_sel_nxt[1] ,
         \u_a23_core/u_decode/barrel_shift_data_sel_nxt[0] ,
         \u_a23_core/u_decode/mtrans_reg_d2[0] ,
         \u_a23_core/u_decode/mtrans_reg_d2[1] ,
         \u_a23_core/u_decode/mtrans_reg_d2[2] ,
         \u_a23_core/u_decode/mtrans_reg_d2[3] ,
         \u_a23_core/u_decode/mtrans_num_registers[0] ,
         \u_a23_core/u_decode/mtrans_num_registers[1] ,
         \u_a23_core/u_decode/mtrans_num_registers[2] ,
         \u_a23_core/u_decode/mtrans_num_registers[3] ,
         \u_a23_core/u_decode/mtrans_num_registers[4] ,
         \u_a23_core/u_decode/N550 , \u_a23_core/u_decode/N549 ,
         \u_a23_core/u_decode/N548 , \u_a23_core/u_decode/N547 ,
         \u_a23_core/u_decode/N544 , \u_a23_core/u_decode/N543 ,
         \u_a23_core/u_decode/N542 , \u_a23_core/u_decode/N539 ,
         \u_a23_core/u_decode/N538 , \u_a23_core/u_decode/N537 ,
         \u_a23_core/u_decode/N533 , \u_a23_core/u_decode/N532 ,
         \u_a23_core/u_decode/N528 , \u_a23_core/u_decode/N527 ,
         \u_a23_core/u_decode/N524 , \u_a23_core/u_decode/N523 ,
         \u_a23_core/u_decode/N521 , \u_a23_core/u_decode/N520 ,
         \u_a23_core/u_decode/N519 , \u_a23_core/u_decode/N518 ,
         \u_a23_core/u_decode/N384 , \u_a23_core/u_decode/N348 ,
         \u_a23_core/u_decode/N319 , \u_a23_core/u_decode/N298 ,
         \u_a23_core/u_decode/alu_function_nxt[0] ,
         \u_a23_core/u_decode/alu_function_nxt[1] ,
         \u_a23_core/u_decode/alu_function_nxt[2] ,
         \u_a23_core/u_decode/alu_function_nxt[3] ,
         \u_a23_core/u_decode/alu_function_nxt[4] ,
         \u_a23_core/u_decode/alu_function_nxt[5] ,
         \u_a23_core/u_decode/alu_function_nxt[6] ,
         \u_a23_core/u_decode/alu_function_nxt[7] ,
         \u_a23_core/u_decode/alu_function_nxt[8] ,
         \u_a23_core/u_decode/shift_imm_zero_nxt ,
         \u_a23_core/u_decode/barrel_shift_amount_sel_nxt[0] ,
         \u_a23_core/u_decode/barrel_shift_amount_sel_nxt[1] ,
         \u_a23_core/u_decode/imm32_nxt[31] ,
         \u_a23_core/u_decode/imm32_nxt[30] ,
         \u_a23_core/u_decode/imm32_nxt[29] ,
         \u_a23_core/u_decode/imm32_nxt[28] ,
         \u_a23_core/u_decode/imm32_nxt[27] ,
         \u_a23_core/u_decode/imm32_nxt[26] ,
         \u_a23_core/u_decode/imm32_nxt[25] ,
         \u_a23_core/u_decode/imm32_nxt[24] ,
         \u_a23_core/u_decode/imm32_nxt[23] ,
         \u_a23_core/u_decode/imm32_nxt[22] ,
         \u_a23_core/u_decode/imm32_nxt[21] ,
         \u_a23_core/u_decode/imm32_nxt[20] ,
         \u_a23_core/u_decode/imm32_nxt[19] ,
         \u_a23_core/u_decode/imm32_nxt[18] ,
         \u_a23_core/u_decode/imm32_nxt[17] ,
         \u_a23_core/u_decode/imm32_nxt[16] ,
         \u_a23_core/u_decode/imm32_nxt[15] ,
         \u_a23_core/u_decode/imm32_nxt[14] ,
         \u_a23_core/u_decode/imm32_nxt[13] ,
         \u_a23_core/u_decode/imm32_nxt[12] ,
         \u_a23_core/u_decode/imm32_nxt[11] ,
         \u_a23_core/u_decode/imm32_nxt[10] ,
         \u_a23_core/u_decode/imm32_nxt[9] ,
         \u_a23_core/u_decode/imm32_nxt[8] ,
         \u_a23_core/u_decode/imm32_nxt[7] ,
         \u_a23_core/u_decode/imm32_nxt[6] ,
         \u_a23_core/u_decode/imm32_nxt[5] ,
         \u_a23_core/u_decode/imm32_nxt[4] ,
         \u_a23_core/u_decode/imm32_nxt[3] ,
         \u_a23_core/u_decode/imm32_nxt[2] ,
         \u_a23_core/u_decode/imm32_nxt[1] ,
         \u_a23_core/u_decode/imm32_nxt[0] ,
         \u_a23_core/u_decode/pc_sel_nxt[0] ,
         \u_a23_core/u_decode/pc_sel_nxt[1] , \u_a23_core/u_decode/pc_wen_nxt ,
         \u_a23_core/u_decode/pre_fetch_instruction[0] ,
         \u_a23_core/u_decode/pre_fetch_instruction[1] ,
         \u_a23_core/u_decode/pre_fetch_instruction[2] ,
         \u_a23_core/u_decode/pre_fetch_instruction[3] ,
         \u_a23_core/u_decode/pre_fetch_instruction[4] ,
         \u_a23_core/u_decode/pre_fetch_instruction[5] ,
         \u_a23_core/u_decode/pre_fetch_instruction[6] ,
         \u_a23_core/u_decode/pre_fetch_instruction[7] ,
         \u_a23_core/u_decode/pre_fetch_instruction[8] ,
         \u_a23_core/u_decode/pre_fetch_instruction[9] ,
         \u_a23_core/u_decode/pre_fetch_instruction[10] ,
         \u_a23_core/u_decode/pre_fetch_instruction[11] ,
         \u_a23_core/u_decode/pre_fetch_instruction[12] ,
         \u_a23_core/u_decode/pre_fetch_instruction[13] ,
         \u_a23_core/u_decode/pre_fetch_instruction[14] ,
         \u_a23_core/u_decode/pre_fetch_instruction[15] ,
         \u_a23_core/u_decode/pre_fetch_instruction[16] ,
         \u_a23_core/u_decode/pre_fetch_instruction[17] ,
         \u_a23_core/u_decode/pre_fetch_instruction[18] ,
         \u_a23_core/u_decode/pre_fetch_instruction[19] ,
         \u_a23_core/u_decode/pre_fetch_instruction[20] ,
         \u_a23_core/u_decode/pre_fetch_instruction[21] ,
         \u_a23_core/u_decode/pre_fetch_instruction[22] ,
         \u_a23_core/u_decode/pre_fetch_instruction[23] ,
         \u_a23_core/u_decode/pre_fetch_instruction[24] ,
         \u_a23_core/u_decode/pre_fetch_instruction[25] ,
         \u_a23_core/u_decode/pre_fetch_instruction[26] ,
         \u_a23_core/u_decode/pre_fetch_instruction[27] ,
         \u_a23_core/u_decode/pre_fetch_instruction[28] ,
         \u_a23_core/u_decode/pre_fetch_instruction[29] ,
         \u_a23_core/u_decode/pre_fetch_instruction[30] ,
         \u_a23_core/u_decode/pre_fetch_instruction[31] ,
         \u_a23_core/u_decode/saved_current_instruction[0] ,
         \u_a23_core/u_decode/saved_current_instruction[1] ,
         \u_a23_core/u_decode/saved_current_instruction[2] ,
         \u_a23_core/u_decode/saved_current_instruction[3] ,
         \u_a23_core/u_decode/saved_current_instruction[4] ,
         \u_a23_core/u_decode/saved_current_instruction[5] ,
         \u_a23_core/u_decode/saved_current_instruction[6] ,
         \u_a23_core/u_decode/saved_current_instruction[7] ,
         \u_a23_core/u_decode/saved_current_instruction[8] ,
         \u_a23_core/u_decode/saved_current_instruction[9] ,
         \u_a23_core/u_decode/saved_current_instruction[10] ,
         \u_a23_core/u_decode/saved_current_instruction[11] ,
         \u_a23_core/u_decode/saved_current_instruction[12] ,
         \u_a23_core/u_decode/saved_current_instruction[13] ,
         \u_a23_core/u_decode/saved_current_instruction[14] ,
         \u_a23_core/u_decode/saved_current_instruction[15] ,
         \u_a23_core/u_decode/saved_current_instruction[16] ,
         \u_a23_core/u_decode/saved_current_instruction[17] ,
         \u_a23_core/u_decode/saved_current_instruction[18] ,
         \u_a23_core/u_decode/saved_current_instruction[19] ,
         \u_a23_core/u_decode/saved_current_instruction[20] ,
         \u_a23_core/u_decode/saved_current_instruction[21] ,
         \u_a23_core/u_decode/saved_current_instruction[22] ,
         \u_a23_core/u_decode/saved_current_instruction[23] ,
         \u_a23_core/u_decode/saved_current_instruction[24] ,
         \u_a23_core/u_decode/saved_current_instruction[25] ,
         \u_a23_core/u_decode/saved_current_instruction[26] ,
         \u_a23_core/u_decode/saved_current_instruction[27] ,
         \u_a23_core/u_decode/instruction[4] ,
         \u_a23_core/u_decode/instruction[5] ,
         \u_a23_core/u_decode/instruction[6] ,
         \u_a23_core/u_decode/instruction[7] ,
         \u_a23_core/u_decode/instruction[8] ,
         \u_a23_core/u_decode/instruction[9] ,
         \u_a23_core/u_decode/instruction[10] ,
         \u_a23_core/u_decode/instruction[11] ,
         \u_a23_core/u_decode/control_state[0] ,
         \u_a23_core/u_decode/control_state[1] ,
         \u_a23_core/u_decode/control_state[2] ,
         \u_a23_core/u_decode/control_state[3] ,
         \u_a23_core/u_decode/control_state[4] , \u_a23_core/u_execute/n1076 ,
         \u_a23_core/u_execute/n1075 , \u_a23_core/u_execute/n1074 ,
         \u_a23_core/u_execute/n1073 , \u_a23_core/u_execute/write_enable_nxt ,
         \u_a23_core/u_execute/write_data_nxt[2] ,
         \u_a23_core/u_execute/write_data_nxt[3] ,
         \u_a23_core/u_execute/write_data_nxt[4] ,
         \u_a23_core/u_execute/write_data_nxt[5] ,
         \u_a23_core/u_execute/write_data_nxt[6] ,
         \u_a23_core/u_execute/write_data_nxt[7] ,
         \u_a23_core/u_execute/write_data_nxt[8] ,
         \u_a23_core/u_execute/write_data_nxt[9] ,
         \u_a23_core/u_execute/write_data_nxt[10] ,
         \u_a23_core/u_execute/write_data_nxt[11] ,
         \u_a23_core/u_execute/write_data_nxt[12] ,
         \u_a23_core/u_execute/write_data_nxt[13] ,
         \u_a23_core/u_execute/write_data_nxt[14] ,
         \u_a23_core/u_execute/write_data_nxt[15] ,
         \u_a23_core/u_execute/write_data_nxt[16] ,
         \u_a23_core/u_execute/write_data_nxt[17] ,
         \u_a23_core/u_execute/write_data_nxt[18] ,
         \u_a23_core/u_execute/write_data_nxt[19] ,
         \u_a23_core/u_execute/write_data_nxt[20] ,
         \u_a23_core/u_execute/write_data_nxt[21] ,
         \u_a23_core/u_execute/write_data_nxt[22] ,
         \u_a23_core/u_execute/write_data_nxt[23] ,
         \u_a23_core/u_execute/write_data_nxt[24] ,
         \u_a23_core/u_execute/write_data_nxt[25] ,
         \u_a23_core/u_execute/write_data_nxt[26] ,
         \u_a23_core/u_execute/write_data_nxt[27] ,
         \u_a23_core/u_execute/write_data_nxt[28] ,
         \u_a23_core/u_execute/write_data_nxt[29] ,
         \u_a23_core/u_execute/write_data_nxt[30] ,
         \u_a23_core/u_execute/write_data_nxt[31] ,
         \u_a23_core/u_execute/byte_enable_nxt[3] ,
         \u_a23_core/u_execute/byte_enable_nxt[2] ,
         \u_a23_core/u_execute/byte_enable_nxt[1] ,
         \u_a23_core/u_execute/byte_enable_nxt[0] ,
         \u_a23_core/u_execute/multiply_out[31] ,
         \u_a23_core/u_execute/multiply_out[30] ,
         \u_a23_core/u_execute/multiply_out[29] ,
         \u_a23_core/u_execute/multiply_out[28] ,
         \u_a23_core/u_execute/multiply_out[27] ,
         \u_a23_core/u_execute/multiply_out[26] ,
         \u_a23_core/u_execute/multiply_out[25] ,
         \u_a23_core/u_execute/multiply_out[24] ,
         \u_a23_core/u_execute/multiply_out[23] ,
         \u_a23_core/u_execute/multiply_out[22] ,
         \u_a23_core/u_execute/multiply_out[21] ,
         \u_a23_core/u_execute/multiply_out[20] ,
         \u_a23_core/u_execute/multiply_out[19] ,
         \u_a23_core/u_execute/multiply_out[18] ,
         \u_a23_core/u_execute/multiply_out[17] ,
         \u_a23_core/u_execute/multiply_out[16] ,
         \u_a23_core/u_execute/multiply_out[15] ,
         \u_a23_core/u_execute/multiply_out[14] ,
         \u_a23_core/u_execute/multiply_out[13] ,
         \u_a23_core/u_execute/multiply_out[12] ,
         \u_a23_core/u_execute/multiply_out[11] ,
         \u_a23_core/u_execute/multiply_out[10] ,
         \u_a23_core/u_execute/multiply_out[9] ,
         \u_a23_core/u_execute/multiply_out[8] ,
         \u_a23_core/u_execute/multiply_out[7] ,
         \u_a23_core/u_execute/multiply_out[6] ,
         \u_a23_core/u_execute/multiply_out[5] ,
         \u_a23_core/u_execute/multiply_out[4] ,
         \u_a23_core/u_execute/multiply_out[3] ,
         \u_a23_core/u_execute/multiply_out[2] ,
         \u_a23_core/u_execute/multiply_out[1] ,
         \u_a23_core/u_execute/multiply_out[0] ,
         \u_a23_core/u_execute/save_int_pc_m4[28] ,
         \u_a23_core/u_execute/save_int_pc_m4[29] ,
         \u_a23_core/u_execute/save_int_pc_m4[30] ,
         \u_a23_core/u_execute/save_int_pc_m4[31] ,
         \u_a23_core/u_execute/alu_out_pc_filtered[2] ,
         \u_a23_core/u_execute/alu_out_pc_filtered[3] ,
         \u_a23_core/u_execute/alu_out_pc_filtered[4] ,
         \u_a23_core/u_execute/alu_out_pc_filtered[5] ,
         \u_a23_core/u_execute/alu_out_pc_filtered[6] ,
         \u_a23_core/u_execute/alu_out_pc_filtered[7] ,
         \u_a23_core/u_execute/alu_out_pc_filtered[8] ,
         \u_a23_core/u_execute/alu_out_pc_filtered[9] ,
         \u_a23_core/u_execute/alu_out_pc_filtered[10] ,
         \u_a23_core/u_execute/alu_out_pc_filtered[11] ,
         \u_a23_core/u_execute/alu_out_pc_filtered[12] ,
         \u_a23_core/u_execute/alu_out_pc_filtered[13] ,
         \u_a23_core/u_execute/alu_out_pc_filtered[14] ,
         \u_a23_core/u_execute/alu_out_pc_filtered[15] ,
         \u_a23_core/u_execute/alu_out_pc_filtered[16] ,
         \u_a23_core/u_execute/alu_out_pc_filtered[17] ,
         \u_a23_core/u_execute/alu_out_pc_filtered[18] ,
         \u_a23_core/u_execute/alu_out_pc_filtered[19] ,
         \u_a23_core/u_execute/alu_out_pc_filtered[20] ,
         \u_a23_core/u_execute/alu_out_pc_filtered[21] ,
         \u_a23_core/u_execute/alu_out_pc_filtered[22] ,
         \u_a23_core/u_execute/alu_out_pc_filtered[23] ,
         \u_a23_core/u_execute/alu_out_pc_filtered[24] ,
         \u_a23_core/u_execute/alu_out_pc_filtered[25] ,
         \u_a23_core/u_execute/rs[0] , \u_a23_core/u_execute/rs[1] ,
         \u_a23_core/u_execute/rs[2] , \u_a23_core/u_execute/rs[3] ,
         \u_a23_core/u_execute/rs[4] , \u_a23_core/u_execute/rs[5] ,
         \u_a23_core/u_execute/rs[6] , \u_a23_core/u_execute/rs[7] ,
         \u_a23_core/u_execute/rs[8] , \u_a23_core/u_execute/rs[9] ,
         \u_a23_core/u_execute/rs[10] , \u_a23_core/u_execute/rs[11] ,
         \u_a23_core/u_execute/rs[12] , \u_a23_core/u_execute/rs[13] ,
         \u_a23_core/u_execute/rs[14] , \u_a23_core/u_execute/rs[15] ,
         \u_a23_core/u_execute/rs[16] , \u_a23_core/u_execute/rs[17] ,
         \u_a23_core/u_execute/rs[18] , \u_a23_core/u_execute/rs[19] ,
         \u_a23_core/u_execute/rs[20] , \u_a23_core/u_execute/rs[21] ,
         \u_a23_core/u_execute/rs[22] , \u_a23_core/u_execute/rs[23] ,
         \u_a23_core/u_execute/rs[24] , \u_a23_core/u_execute/rs[25] ,
         \u_a23_core/u_execute/rs[26] , \u_a23_core/u_execute/rs[27] ,
         \u_a23_core/u_execute/rs[28] , \u_a23_core/u_execute/rs[29] ,
         \u_a23_core/u_execute/rs[30] , \u_a23_core/u_execute/rs[31] ,
         \u_a23_core/u_execute/rn_plus4[31] ,
         \u_a23_core/u_execute/rn_plus4[30] ,
         \u_a23_core/u_execute/rn_plus4[29] ,
         \u_a23_core/u_execute/rn_plus4[28] ,
         \u_a23_core/u_execute/rn_plus4[27] ,
         \u_a23_core/u_execute/rn_plus4[26] ,
         \u_a23_core/u_execute/rn_plus4[25] ,
         \u_a23_core/u_execute/rn_plus4[24] ,
         \u_a23_core/u_execute/rn_plus4[23] ,
         \u_a23_core/u_execute/rn_plus4[22] ,
         \u_a23_core/u_execute/rn_plus4[21] ,
         \u_a23_core/u_execute/rn_plus4[20] ,
         \u_a23_core/u_execute/rn_plus4[19] ,
         \u_a23_core/u_execute/rn_plus4[18] ,
         \u_a23_core/u_execute/rn_plus4[17] ,
         \u_a23_core/u_execute/rn_plus4[16] ,
         \u_a23_core/u_execute/rn_plus4[15] ,
         \u_a23_core/u_execute/rn_plus4[14] ,
         \u_a23_core/u_execute/rn_plus4[13] ,
         \u_a23_core/u_execute/rn_plus4[12] ,
         \u_a23_core/u_execute/rn_plus4[11] ,
         \u_a23_core/u_execute/rn_plus4[10] ,
         \u_a23_core/u_execute/rn_plus4[9] ,
         \u_a23_core/u_execute/rn_plus4[8] ,
         \u_a23_core/u_execute/rn_plus4[7] ,
         \u_a23_core/u_execute/rn_plus4[6] ,
         \u_a23_core/u_execute/rn_plus4[5] ,
         \u_a23_core/u_execute/rn_plus4[4] ,
         \u_a23_core/u_execute/rn_plus4[3] , \u_a23_core/u_execute/rn[2] ,
         \u_a23_core/u_execute/rn[3] , \u_a23_core/u_execute/rn[4] ,
         \u_a23_core/u_execute/rn[5] , \u_a23_core/u_execute/rn[6] ,
         \u_a23_core/u_execute/rn[7] , \u_a23_core/u_execute/rn[8] ,
         \u_a23_core/u_execute/rn[9] , \u_a23_core/u_execute/rn[10] ,
         \u_a23_core/u_execute/rn[11] , \u_a23_core/u_execute/rn[12] ,
         \u_a23_core/u_execute/rn[13] , \u_a23_core/u_execute/rn[14] ,
         \u_a23_core/u_execute/rn[15] , \u_a23_core/u_execute/rn[16] ,
         \u_a23_core/u_execute/rn[17] , \u_a23_core/u_execute/rn[18] ,
         \u_a23_core/u_execute/rn[19] , \u_a23_core/u_execute/rn[20] ,
         \u_a23_core/u_execute/rn[21] , \u_a23_core/u_execute/rn[22] ,
         \u_a23_core/u_execute/rn[23] , \u_a23_core/u_execute/rn[24] ,
         \u_a23_core/u_execute/rn[25] , \u_a23_core/u_execute/rn[26] ,
         \u_a23_core/u_execute/rn[27] , \u_a23_core/u_execute/rn[28] ,
         \u_a23_core/u_execute/rn[29] , \u_a23_core/u_execute/rn[30] ,
         \u_a23_core/u_execute/rn[31] , \u_a23_core/u_execute/alu_plus4[31] ,
         \u_a23_core/u_execute/alu_plus4[30] ,
         \u_a23_core/u_execute/alu_plus4[29] ,
         \u_a23_core/u_execute/alu_plus4[28] ,
         \u_a23_core/u_execute/alu_plus4[27] ,
         \u_a23_core/u_execute/alu_plus4[26] ,
         \u_a23_core/u_execute/alu_plus4[25] ,
         \u_a23_core/u_execute/alu_plus4[24] ,
         \u_a23_core/u_execute/alu_plus4[23] ,
         \u_a23_core/u_execute/alu_plus4[22] ,
         \u_a23_core/u_execute/alu_plus4[21] ,
         \u_a23_core/u_execute/alu_plus4[20] ,
         \u_a23_core/u_execute/alu_plus4[19] ,
         \u_a23_core/u_execute/alu_plus4[18] ,
         \u_a23_core/u_execute/alu_plus4[17] ,
         \u_a23_core/u_execute/alu_plus4[16] ,
         \u_a23_core/u_execute/alu_plus4[15] ,
         \u_a23_core/u_execute/alu_plus4[14] ,
         \u_a23_core/u_execute/alu_plus4[13] ,
         \u_a23_core/u_execute/alu_plus4[12] ,
         \u_a23_core/u_execute/alu_plus4[11] ,
         \u_a23_core/u_execute/alu_plus4[10] ,
         \u_a23_core/u_execute/alu_plus4[9] ,
         \u_a23_core/u_execute/alu_plus4[8] ,
         \u_a23_core/u_execute/alu_plus4[7] ,
         \u_a23_core/u_execute/alu_plus4[6] ,
         \u_a23_core/u_execute/alu_plus4[5] ,
         \u_a23_core/u_execute/alu_plus4[4] ,
         \u_a23_core/u_execute/alu_plus4[3] ,
         \u_a23_core/u_execute/address_plus4[31] ,
         \u_a23_core/u_execute/address_plus4[30] ,
         \u_a23_core/u_execute/address_plus4[29] ,
         \u_a23_core/u_execute/address_plus4[28] ,
         \u_a23_core/u_execute/address_plus4[27] ,
         \u_a23_core/u_execute/address_plus4[26] ,
         \u_a23_core/u_execute/address_plus4[25] ,
         \u_a23_core/u_execute/address_plus4[24] ,
         \u_a23_core/u_execute/address_plus4[23] ,
         \u_a23_core/u_execute/address_plus4[22] ,
         \u_a23_core/u_execute/address_plus4[21] ,
         \u_a23_core/u_execute/address_plus4[20] ,
         \u_a23_core/u_execute/address_plus4[19] ,
         \u_a23_core/u_execute/address_plus4[18] ,
         \u_a23_core/u_execute/address_plus4[17] ,
         \u_a23_core/u_execute/address_plus4[16] ,
         \u_a23_core/u_execute/address_plus4[15] ,
         \u_a23_core/u_execute/address_plus4[14] ,
         \u_a23_core/u_execute/address_plus4[13] ,
         \u_a23_core/u_execute/address_plus4[12] ,
         \u_a23_core/u_execute/address_plus4[11] ,
         \u_a23_core/u_execute/address_plus4[10] ,
         \u_a23_core/u_execute/address_plus4[9] ,
         \u_a23_core/u_execute/address_plus4[8] ,
         \u_a23_core/u_execute/address_plus4[7] ,
         \u_a23_core/u_execute/address_plus4[6] ,
         \u_a23_core/u_execute/address_plus4[5] ,
         \u_a23_core/u_execute/address_plus4[4] ,
         \u_a23_core/u_execute/address_plus4[3] ,
         \u_a23_core/u_execute/address_plus4[0] ,
         \u_a23_core/u_execute/pc_minus4[3] ,
         \u_a23_core/u_execute/pc_minus4[4] ,
         \u_a23_core/u_execute/pc_minus4[5] ,
         \u_a23_core/u_execute/pc_minus4[6] ,
         \u_a23_core/u_execute/pc_minus4[7] ,
         \u_a23_core/u_execute/pc_minus4[8] ,
         \u_a23_core/u_execute/pc_minus4[9] ,
         \u_a23_core/u_execute/pc_minus4[10] ,
         \u_a23_core/u_execute/pc_minus4[11] ,
         \u_a23_core/u_execute/pc_minus4[12] ,
         \u_a23_core/u_execute/pc_minus4[13] ,
         \u_a23_core/u_execute/pc_minus4[14] ,
         \u_a23_core/u_execute/pc_minus4[15] ,
         \u_a23_core/u_execute/pc_minus4[16] ,
         \u_a23_core/u_execute/pc_minus4[17] ,
         \u_a23_core/u_execute/pc_minus4[18] ,
         \u_a23_core/u_execute/pc_minus4[19] ,
         \u_a23_core/u_execute/pc_minus4[20] ,
         \u_a23_core/u_execute/pc_minus4[21] ,
         \u_a23_core/u_execute/pc_minus4[22] ,
         \u_a23_core/u_execute/pc_minus4[23] ,
         \u_a23_core/u_execute/pc_minus4[24] ,
         \u_a23_core/u_execute/pc_minus4[25] ,
         \u_a23_core/u_execute/pc_plus4[3] ,
         \u_a23_core/u_execute/pc_plus4[4] ,
         \u_a23_core/u_execute/pc_plus4[5] ,
         \u_a23_core/u_execute/pc_plus4[6] ,
         \u_a23_core/u_execute/pc_plus4[7] ,
         \u_a23_core/u_execute/pc_plus4[8] ,
         \u_a23_core/u_execute/pc_plus4[9] ,
         \u_a23_core/u_execute/pc_plus4[10] ,
         \u_a23_core/u_execute/pc_plus4[11] ,
         \u_a23_core/u_execute/pc_plus4[12] ,
         \u_a23_core/u_execute/pc_plus4[13] ,
         \u_a23_core/u_execute/pc_plus4[14] ,
         \u_a23_core/u_execute/pc_plus4[15] ,
         \u_a23_core/u_execute/pc_plus4[16] ,
         \u_a23_core/u_execute/pc_plus4[17] ,
         \u_a23_core/u_execute/pc_plus4[18] ,
         \u_a23_core/u_execute/pc_plus4[19] ,
         \u_a23_core/u_execute/pc_plus4[20] ,
         \u_a23_core/u_execute/pc_plus4[21] ,
         \u_a23_core/u_execute/pc_plus4[22] ,
         \u_a23_core/u_execute/pc_plus4[23] ,
         \u_a23_core/u_execute/pc_plus4[24] ,
         \u_a23_core/u_execute/pc_plus4[25] ,
         \u_a23_core/u_execute/pc_plus4[26] , \u_a23_core/u_execute/pc[2] ,
         \u_a23_core/u_execute/pc[3] , \u_a23_core/u_execute/pc[4] ,
         \u_a23_core/u_execute/pc[5] , \u_a23_core/u_execute/pc[6] ,
         \u_a23_core/u_execute/pc[7] , \u_a23_core/u_execute/pc[8] ,
         \u_a23_core/u_execute/pc[9] , \u_a23_core/u_execute/pc[10] ,
         \u_a23_core/u_execute/pc[11] , \u_a23_core/u_execute/pc[12] ,
         \u_a23_core/u_execute/pc[13] , \u_a23_core/u_execute/pc[14] ,
         \u_a23_core/u_execute/pc[15] , \u_a23_core/u_execute/pc[16] ,
         \u_a23_core/u_execute/pc[17] , \u_a23_core/u_execute/pc[18] ,
         \u_a23_core/u_execute/pc[19] , \u_a23_core/u_execute/pc[20] ,
         \u_a23_core/u_execute/pc[21] , \u_a23_core/u_execute/pc[22] ,
         \u_a23_core/u_execute/pc[23] , \u_a23_core/u_execute/pc[24] ,
         \u_a23_core/u_execute/pc[25] , \u_a23_core/u_execute/alu_out[26] ,
         \u_a23_core/u_execute/alu_out[27] ,
         \u_a23_core/u_execute/alu_out[28] ,
         \u_a23_core/u_execute/alu_out[29] ,
         \u_a23_core/u_execute/alu_out[30] ,
         \u_a23_core/u_execute/alu_out[31] ,
         \u_a23_core/u_execute/u_alu/fadder_out[0] ,
         \u_a23_core/u_execute/u_alu/fadder_out[1] ,
         \u_a23_core/u_execute/u_alu/fadder_out[2] ,
         \u_a23_core/u_execute/u_alu/fadder_out[3] ,
         \u_a23_core/u_execute/u_alu/fadder_out[4] ,
         \u_a23_core/u_execute/u_alu/fadder_out[5] ,
         \u_a23_core/u_execute/u_alu/fadder_out[6] ,
         \u_a23_core/u_execute/u_alu/fadder_out[7] ,
         \u_a23_core/u_execute/u_alu/fadder_out[8] ,
         \u_a23_core/u_execute/u_alu/fadder_out[9] ,
         \u_a23_core/u_execute/u_alu/fadder_out[10] ,
         \u_a23_core/u_execute/u_alu/fadder_out[11] ,
         \u_a23_core/u_execute/u_alu/fadder_out[12] ,
         \u_a23_core/u_execute/u_alu/fadder_out[13] ,
         \u_a23_core/u_execute/u_alu/fadder_out[14] ,
         \u_a23_core/u_execute/u_alu/fadder_out[15] ,
         \u_a23_core/u_execute/u_alu/fadder_out[16] ,
         \u_a23_core/u_execute/u_alu/fadder_out[17] ,
         \u_a23_core/u_execute/u_alu/fadder_out[18] ,
         \u_a23_core/u_execute/u_alu/fadder_out[19] ,
         \u_a23_core/u_execute/u_alu/fadder_out[20] ,
         \u_a23_core/u_execute/u_alu/fadder_out[21] ,
         \u_a23_core/u_execute/u_alu/fadder_out[22] ,
         \u_a23_core/u_execute/u_alu/fadder_out[23] ,
         \u_a23_core/u_execute/u_alu/fadder_out[24] ,
         \u_a23_core/u_execute/u_alu/fadder_out[25] ,
         \u_a23_core/u_execute/u_alu/fadder_out[26] ,
         \u_a23_core/u_execute/u_alu/fadder_out[27] ,
         \u_a23_core/u_execute/u_alu/fadder_out[28] ,
         \u_a23_core/u_execute/u_alu/fadder_out[29] ,
         \u_a23_core/u_execute/u_alu/fadder_out[30] ,
         \u_a23_core/u_execute/u_alu/fadder_out[31] ,
         \u_a23_core/u_execute/u_alu/fadder_out[32] ,
         \u_a23_core/u_execute/u_alu/carry_in ,
         \u_a23_core/u_execute/u_alu/b_not[0] ,
         \u_a23_core/u_execute/u_alu/b_not[1] ,
         \u_a23_core/u_execute/u_alu/b_not[2] ,
         \u_a23_core/u_execute/u_alu/b_not[3] ,
         \u_a23_core/u_execute/u_alu/b_not[4] ,
         \u_a23_core/u_execute/u_alu/b_not[5] ,
         \u_a23_core/u_execute/u_alu/b_not[6] ,
         \u_a23_core/u_execute/u_alu/b_not[7] ,
         \u_a23_core/u_execute/u_alu/b_not[8] ,
         \u_a23_core/u_execute/u_alu/b_not[9] ,
         \u_a23_core/u_execute/u_alu/b_not[10] ,
         \u_a23_core/u_execute/u_alu/b_not[11] ,
         \u_a23_core/u_execute/u_alu/b_not[12] ,
         \u_a23_core/u_execute/u_alu/b_not[13] ,
         \u_a23_core/u_execute/u_alu/b_not[14] ,
         \u_a23_core/u_execute/u_alu/b_not[15] ,
         \u_a23_core/u_execute/u_alu/b_not[16] ,
         \u_a23_core/u_execute/u_alu/b_not[17] ,
         \u_a23_core/u_execute/u_alu/b_not[18] ,
         \u_a23_core/u_execute/u_alu/b_not[19] ,
         \u_a23_core/u_execute/u_alu/b_not[20] ,
         \u_a23_core/u_execute/u_alu/b_not[21] ,
         \u_a23_core/u_execute/u_alu/b_not[22] ,
         \u_a23_core/u_execute/u_alu/b_not[23] ,
         \u_a23_core/u_execute/u_alu/b_not[24] ,
         \u_a23_core/u_execute/u_alu/b_not[25] ,
         \u_a23_core/u_execute/u_alu/b_not[26] ,
         \u_a23_core/u_execute/u_alu/b_not[27] ,
         \u_a23_core/u_execute/u_alu/b_not[28] ,
         \u_a23_core/u_execute/u_alu/b_not[29] ,
         \u_a23_core/u_execute/u_alu/b_not[30] ,
         \u_a23_core/u_execute/u_alu/b_not[31] ,
         \u_a23_core/u_execute/u_alu/a[0] , \u_a23_core/u_execute/u_alu/a[1] ,
         \u_a23_core/u_execute/u_alu/a[2] , \u_a23_core/u_execute/u_alu/a[3] ,
         \u_a23_core/u_execute/u_alu/a[4] , \u_a23_core/u_execute/u_alu/a[5] ,
         \u_a23_core/u_execute/u_alu/a[6] , \u_a23_core/u_execute/u_alu/a[7] ,
         \u_a23_core/u_execute/u_alu/a[8] , \u_a23_core/u_execute/u_alu/a[9] ,
         \u_a23_core/u_execute/u_alu/a[10] ,
         \u_a23_core/u_execute/u_alu/a[11] ,
         \u_a23_core/u_execute/u_alu/a[12] ,
         \u_a23_core/u_execute/u_alu/a[13] ,
         \u_a23_core/u_execute/u_alu/a[14] ,
         \u_a23_core/u_execute/u_alu/a[15] ,
         \u_a23_core/u_execute/u_alu/a[16] ,
         \u_a23_core/u_execute/u_alu/a[17] ,
         \u_a23_core/u_execute/u_alu/a[18] ,
         \u_a23_core/u_execute/u_alu/a[19] ,
         \u_a23_core/u_execute/u_alu/a[20] ,
         \u_a23_core/u_execute/u_alu/a[21] ,
         \u_a23_core/u_execute/u_alu/a[22] ,
         \u_a23_core/u_execute/u_alu/a[23] ,
         \u_a23_core/u_execute/u_alu/a[24] ,
         \u_a23_core/u_execute/u_alu/a[25] ,
         \u_a23_core/u_execute/u_alu/a[26] ,
         \u_a23_core/u_execute/u_alu/a[27] ,
         \u_a23_core/u_execute/u_alu/a[28] ,
         \u_a23_core/u_execute/u_alu/a[29] ,
         \u_a23_core/u_execute/u_alu/a[30] ,
         \u_a23_core/u_execute/u_alu/a[31] ,
         \u_a23_core/u_execute/u_multiply/n611 ,
         \u_a23_core/u_execute/u_multiply/n610 ,
         \u_a23_core/u_execute/u_multiply/n609 ,
         \u_a23_core/u_execute/u_multiply/n608 ,
         \u_a23_core/u_execute/u_multiply/n607 ,
         \u_a23_core/u_execute/u_multiply/n606 ,
         \u_a23_core/u_execute/u_multiply/n605 ,
         \u_a23_core/u_execute/u_multiply/n604 ,
         \u_a23_core/u_execute/u_multiply/n603 ,
         \u_a23_core/u_execute/u_multiply/n602 ,
         \u_a23_core/u_execute/u_multiply/n601 ,
         \u_a23_core/u_execute/u_multiply/n600 ,
         \u_a23_core/u_execute/u_multiply/n599 ,
         \u_a23_core/u_execute/u_multiply/n598 ,
         \u_a23_core/u_execute/u_multiply/n597 ,
         \u_a23_core/u_execute/u_multiply/n596 ,
         \u_a23_core/u_execute/u_multiply/n595 ,
         \u_a23_core/u_execute/u_multiply/n594 ,
         \u_a23_core/u_execute/u_multiply/n593 ,
         \u_a23_core/u_execute/u_multiply/n592 ,
         \u_a23_core/u_execute/u_multiply/n591 ,
         \u_a23_core/u_execute/u_multiply/n590 ,
         \u_a23_core/u_execute/u_multiply/n589 ,
         \u_a23_core/u_execute/u_multiply/n588 ,
         \u_a23_core/u_execute/u_multiply/n587 ,
         \u_a23_core/u_execute/u_multiply/n586 ,
         \u_a23_core/u_execute/u_multiply/n585 ,
         \u_a23_core/u_execute/u_multiply/n584 ,
         \u_a23_core/u_execute/u_multiply/n583 ,
         \u_a23_core/u_execute/u_multiply/n582 ,
         \u_a23_core/u_execute/u_multiply/n581 ,
         \u_a23_core/u_execute/u_multiply/n580 ,
         \u_a23_core/u_execute/u_multiply/n579 ,
         \u_a23_core/u_execute/u_multiply/n578 ,
         \u_a23_core/u_execute/u_multiply/n577 ,
         \u_a23_core/u_execute/u_multiply/n576 ,
         \u_a23_core/u_execute/u_multiply/n575 ,
         \u_a23_core/u_execute/u_multiply/n574 ,
         \u_a23_core/u_execute/u_multiply/n573 ,
         \u_a23_core/u_execute/u_multiply/n572 ,
         \u_a23_core/u_execute/u_multiply/n571 ,
         \u_a23_core/u_execute/u_multiply/n570 ,
         \u_a23_core/u_execute/u_multiply/n569 ,
         \u_a23_core/u_execute/u_multiply/n568 ,
         \u_a23_core/u_execute/u_multiply/n567 ,
         \u_a23_core/u_execute/u_multiply/n566 ,
         \u_a23_core/u_execute/u_multiply/n565 ,
         \u_a23_core/u_execute/u_multiply/n564 ,
         \u_a23_core/u_execute/u_multiply/n563 ,
         \u_a23_core/u_execute/u_multiply/n562 ,
         \u_a23_core/u_execute/u_multiply/n561 ,
         \u_a23_core/u_execute/u_multiply/n560 ,
         \u_a23_core/u_execute/u_multiply/n559 ,
         \u_a23_core/u_execute/u_multiply/n558 ,
         \u_a23_core/u_execute/u_multiply/n557 ,
         \u_a23_core/u_execute/u_multiply/n556 ,
         \u_a23_core/u_execute/u_multiply/n555 ,
         \u_a23_core/u_execute/u_multiply/n554 ,
         \u_a23_core/u_execute/u_multiply/n553 ,
         \u_a23_core/u_execute/u_multiply/n552 ,
         \u_a23_core/u_execute/u_multiply/n551 ,
         \u_a23_core/u_execute/u_multiply/n550 ,
         \u_a23_core/u_execute/u_multiply/n549 ,
         \u_a23_core/u_execute/u_multiply/n548 ,
         \u_a23_core/u_execute/u_multiply/n547 ,
         \u_a23_core/u_execute/u_multiply/n546 ,
         \u_a23_core/u_execute/u_multiply/n545 ,
         \u_a23_core/u_execute/u_multiply/n544 ,
         \u_a23_core/u_execute/u_multiply/n543 ,
         \u_a23_core/u_execute/u_multiply/n509 ,
         \u_a23_core/u_execute/u_multiply/n507 ,
         \u_a23_core/u_execute/u_multiply/n505 ,
         \u_a23_core/u_execute/u_multiply/n503 ,
         \u_a23_core/u_execute/u_multiply/n501 ,
         \u_a23_core/u_execute/u_multiply/n499 ,
         \u_a23_core/u_execute/u_multiply/N58 ,
         \u_a23_core/u_execute/u_multiply/N57 ,
         \u_a23_core/u_execute/u_multiply/N56 ,
         \u_a23_core/u_execute/u_multiply/N55 ,
         \u_a23_core/u_execute/u_multiply/count[0] ,
         \u_a23_core/u_execute/u_multiply/count[1] ,
         \u_a23_core/u_execute/u_multiply/count[2] ,
         \u_a23_core/u_execute/u_multiply/count[3] ,
         \u_a23_core/u_execute/u_multiply/count[4] ,
         \u_a23_core/u_execute/u_multiply/count[5] ,
         \u_a23_core/u_execute/u_multiply/sum_acc1[31] ,
         \u_a23_core/u_execute/u_multiply/sum_acc1[30] ,
         \u_a23_core/u_execute/u_multiply/sum_acc1[29] ,
         \u_a23_core/u_execute/u_multiply/sum_acc1[28] ,
         \u_a23_core/u_execute/u_multiply/sum_acc1[27] ,
         \u_a23_core/u_execute/u_multiply/sum_acc1[26] ,
         \u_a23_core/u_execute/u_multiply/sum_acc1[25] ,
         \u_a23_core/u_execute/u_multiply/sum_acc1[24] ,
         \u_a23_core/u_execute/u_multiply/sum_acc1[23] ,
         \u_a23_core/u_execute/u_multiply/sum_acc1[22] ,
         \u_a23_core/u_execute/u_multiply/sum_acc1[21] ,
         \u_a23_core/u_execute/u_multiply/sum_acc1[20] ,
         \u_a23_core/u_execute/u_multiply/sum_acc1[19] ,
         \u_a23_core/u_execute/u_multiply/sum_acc1[18] ,
         \u_a23_core/u_execute/u_multiply/sum_acc1[17] ,
         \u_a23_core/u_execute/u_multiply/sum_acc1[16] ,
         \u_a23_core/u_execute/u_multiply/sum_acc1[15] ,
         \u_a23_core/u_execute/u_multiply/sum_acc1[14] ,
         \u_a23_core/u_execute/u_multiply/sum_acc1[13] ,
         \u_a23_core/u_execute/u_multiply/sum_acc1[12] ,
         \u_a23_core/u_execute/u_multiply/sum_acc1[11] ,
         \u_a23_core/u_execute/u_multiply/sum_acc1[10] ,
         \u_a23_core/u_execute/u_multiply/sum_acc1[9] ,
         \u_a23_core/u_execute/u_multiply/sum_acc1[8] ,
         \u_a23_core/u_execute/u_multiply/sum_acc1[7] ,
         \u_a23_core/u_execute/u_multiply/sum_acc1[6] ,
         \u_a23_core/u_execute/u_multiply/sum_acc1[5] ,
         \u_a23_core/u_execute/u_multiply/sum_acc1[4] ,
         \u_a23_core/u_execute/u_multiply/sum_acc1[3] ,
         \u_a23_core/u_execute/u_multiply/sum_acc1[2] ,
         \u_a23_core/u_execute/u_multiply/sum_acc1[1] ,
         \u_a23_core/u_execute/u_multiply/sum_acc1[0] ,
         \u_a23_core/u_execute/u_multiply/sum[33] ,
         \u_a23_core/u_execute/u_multiply/sum[32] ,
         \u_a23_core/u_execute/u_multiply/sum[31] ,
         \u_a23_core/u_execute/u_multiply/sum[30] ,
         \u_a23_core/u_execute/u_multiply/sum[29] ,
         \u_a23_core/u_execute/u_multiply/sum[28] ,
         \u_a23_core/u_execute/u_multiply/sum[27] ,
         \u_a23_core/u_execute/u_multiply/sum[26] ,
         \u_a23_core/u_execute/u_multiply/sum[25] ,
         \u_a23_core/u_execute/u_multiply/sum[24] ,
         \u_a23_core/u_execute/u_multiply/sum[23] ,
         \u_a23_core/u_execute/u_multiply/sum[22] ,
         \u_a23_core/u_execute/u_multiply/sum[21] ,
         \u_a23_core/u_execute/u_multiply/sum[20] ,
         \u_a23_core/u_execute/u_multiply/sum[19] ,
         \u_a23_core/u_execute/u_multiply/sum[18] ,
         \u_a23_core/u_execute/u_multiply/sum[17] ,
         \u_a23_core/u_execute/u_multiply/sum[16] ,
         \u_a23_core/u_execute/u_multiply/sum[15] ,
         \u_a23_core/u_execute/u_multiply/sum[14] ,
         \u_a23_core/u_execute/u_multiply/sum[13] ,
         \u_a23_core/u_execute/u_multiply/sum[12] ,
         \u_a23_core/u_execute/u_multiply/sum[11] ,
         \u_a23_core/u_execute/u_multiply/sum[10] ,
         \u_a23_core/u_execute/u_multiply/sum[9] ,
         \u_a23_core/u_execute/u_multiply/sum[8] ,
         \u_a23_core/u_execute/u_multiply/sum[7] ,
         \u_a23_core/u_execute/u_multiply/sum[6] ,
         \u_a23_core/u_execute/u_multiply/sum[5] ,
         \u_a23_core/u_execute/u_multiply/sum[4] ,
         \u_a23_core/u_execute/u_multiply/sum[3] ,
         \u_a23_core/u_execute/u_multiply/sum[2] ,
         \u_a23_core/u_execute/u_multiply/sum[1] ,
         \u_a23_core/u_execute/u_multiply/sum[0] ,
         \u_a23_core/u_execute/u_multiply/sum34_b[33] ,
         \u_a23_core/u_execute/u_multiply/sum34_b[31] ,
         \u_a23_core/u_execute/u_multiply/sum34_b[30] ,
         \u_a23_core/u_execute/u_multiply/sum34_b[29] ,
         \u_a23_core/u_execute/u_multiply/sum34_b[28] ,
         \u_a23_core/u_execute/u_multiply/sum34_b[27] ,
         \u_a23_core/u_execute/u_multiply/sum34_b[26] ,
         \u_a23_core/u_execute/u_multiply/sum34_b[25] ,
         \u_a23_core/u_execute/u_multiply/sum34_b[24] ,
         \u_a23_core/u_execute/u_multiply/sum34_b[23] ,
         \u_a23_core/u_execute/u_multiply/sum34_b[22] ,
         \u_a23_core/u_execute/u_multiply/sum34_b[21] ,
         \u_a23_core/u_execute/u_multiply/sum34_b[20] ,
         \u_a23_core/u_execute/u_multiply/sum34_b[19] ,
         \u_a23_core/u_execute/u_multiply/sum34_b[18] ,
         \u_a23_core/u_execute/u_multiply/sum34_b[17] ,
         \u_a23_core/u_execute/u_multiply/sum34_b[16] ,
         \u_a23_core/u_execute/u_multiply/sum34_b[15] ,
         \u_a23_core/u_execute/u_multiply/sum34_b[14] ,
         \u_a23_core/u_execute/u_multiply/sum34_b[13] ,
         \u_a23_core/u_execute/u_multiply/sum34_b[12] ,
         \u_a23_core/u_execute/u_multiply/sum34_b[11] ,
         \u_a23_core/u_execute/u_multiply/sum34_b[10] ,
         \u_a23_core/u_execute/u_multiply/sum34_b[9] ,
         \u_a23_core/u_execute/u_multiply/sum34_b[8] ,
         \u_a23_core/u_execute/u_multiply/sum34_b[7] ,
         \u_a23_core/u_execute/u_multiply/sum34_b[6] ,
         \u_a23_core/u_execute/u_multiply/sum34_b[5] ,
         \u_a23_core/u_execute/u_multiply/sum34_b[4] ,
         \u_a23_core/u_execute/u_multiply/sum34_b[3] ,
         \u_a23_core/u_execute/u_multiply/sum34_b[2] ,
         \u_a23_core/u_execute/u_multiply/sum34_b[1] ,
         \u_a23_core/u_execute/u_multiply/sum34_b[0] ,
         \u_a23_core/u_execute/u_multiply/product_0 ,
         \u_a23_core/u_execute/u_multiply/product[33] ,
         \u_a23_core/u_execute/u_multiply/product[34] ,
         \u_a23_core/u_execute/u_multiply/product[35] ,
         \u_a23_core/u_execute/u_multiply/product[36] ,
         \u_a23_core/u_execute/u_multiply/product[37] ,
         \u_a23_core/u_execute/u_multiply/product[38] ,
         \u_a23_core/u_execute/u_multiply/product[39] ,
         \u_a23_core/u_execute/u_multiply/product[40] ,
         \u_a23_core/u_execute/u_multiply/product[41] ,
         \u_a23_core/u_execute/u_multiply/product[42] ,
         \u_a23_core/u_execute/u_multiply/product[43] ,
         \u_a23_core/u_execute/u_multiply/product[44] ,
         \u_a23_core/u_execute/u_multiply/product[45] ,
         \u_a23_core/u_execute/u_multiply/product[46] ,
         \u_a23_core/u_execute/u_multiply/product[47] ,
         \u_a23_core/u_execute/u_multiply/product[48] ,
         \u_a23_core/u_execute/u_multiply/product[49] ,
         \u_a23_core/u_execute/u_multiply/product[50] ,
         \u_a23_core/u_execute/u_multiply/product[51] ,
         \u_a23_core/u_execute/u_multiply/product[52] ,
         \u_a23_core/u_execute/u_multiply/product[53] ,
         \u_a23_core/u_execute/u_multiply/product[54] ,
         \u_a23_core/u_execute/u_multiply/product[55] ,
         \u_a23_core/u_execute/u_multiply/product[56] ,
         \u_a23_core/u_execute/u_multiply/product[57] ,
         \u_a23_core/u_execute/u_multiply/product[58] ,
         \u_a23_core/u_execute/u_multiply/product[59] ,
         \u_a23_core/u_execute/u_multiply/product[60] ,
         \u_a23_core/u_execute/u_multiply/product[61] ,
         \u_a23_core/u_execute/u_multiply/product[62] ,
         \u_a23_core/u_execute/u_multiply/product[63] ,
         \u_a23_core/u_execute/u_multiply/product[64] ,
         \u_a23_core/u_execute/u_multiply/product[65] ,
         \u_a23_core/u_execute/u_multiply/product[66] ,
         \u_a23_core/u_execute/u_multiply/product[67] ,
         \u_a23_core/u_execute/u_multiply/multiplier_bar[31] ,
         \u_a23_core/u_execute/u_multiply/multiplier_bar[30] ,
         \u_a23_core/u_execute/u_multiply/multiplier_bar[29] ,
         \u_a23_core/u_execute/u_multiply/multiplier_bar[28] ,
         \u_a23_core/u_execute/u_multiply/multiplier_bar[27] ,
         \u_a23_core/u_execute/u_multiply/multiplier_bar[26] ,
         \u_a23_core/u_execute/u_multiply/multiplier_bar[25] ,
         \u_a23_core/u_execute/u_multiply/multiplier_bar[24] ,
         \u_a23_core/u_execute/u_multiply/multiplier_bar[23] ,
         \u_a23_core/u_execute/u_multiply/multiplier_bar[22] ,
         \u_a23_core/u_execute/u_multiply/multiplier_bar[21] ,
         \u_a23_core/u_execute/u_multiply/multiplier_bar[20] ,
         \u_a23_core/u_execute/u_multiply/multiplier_bar[19] ,
         \u_a23_core/u_execute/u_multiply/multiplier_bar[18] ,
         \u_a23_core/u_execute/u_multiply/multiplier_bar[17] ,
         \u_a23_core/u_execute/u_multiply/multiplier_bar[16] ,
         \u_a23_core/u_execute/u_multiply/multiplier_bar[15] ,
         \u_a23_core/u_execute/u_multiply/multiplier_bar[14] ,
         \u_a23_core/u_execute/u_multiply/multiplier_bar[13] ,
         \u_a23_core/u_execute/u_multiply/multiplier_bar[12] ,
         \u_a23_core/u_execute/u_multiply/multiplier_bar[11] ,
         \u_a23_core/u_execute/u_multiply/multiplier_bar[10] ,
         \u_a23_core/u_execute/u_multiply/multiplier_bar[9] ,
         \u_a23_core/u_execute/u_multiply/multiplier_bar[8] ,
         \u_a23_core/u_execute/u_multiply/multiplier_bar[7] ,
         \u_a23_core/u_execute/u_multiply/multiplier_bar[6] ,
         \u_a23_core/u_execute/u_multiply/multiplier_bar[5] ,
         \u_a23_core/u_execute/u_multiply/multiplier_bar[4] ,
         \u_a23_core/u_execute/u_multiply/multiplier_bar[3] ,
         \u_a23_core/u_execute/u_multiply/multiplier_bar[2] ,
         \u_a23_core/u_execute/u_multiply/multiplier_bar[1] ,
         \u_a23_core/u_execute/u_register_bank/n4981 ,
         \u_a23_core/u_execute/u_register_bank/n4979 ,
         \u_a23_core/u_execute/u_register_bank/n4977 ,
         \u_a23_core/u_execute/u_register_bank/n4975 ,
         \u_a23_core/u_execute/u_register_bank/n4973 ,
         \u_a23_core/u_execute/u_register_bank/n4971 ,
         \u_a23_core/u_execute/u_register_bank/n4969 ,
         \u_a23_core/u_execute/u_register_bank/n4967 ,
         \u_a23_core/u_execute/u_register_bank/n4965 ,
         \u_a23_core/u_execute/u_register_bank/n4963 ,
         \u_a23_core/u_execute/u_register_bank/n4961 ,
         \u_a23_core/u_execute/u_register_bank/n4959 ,
         \u_a23_core/u_execute/u_register_bank/n4957 ,
         \u_a23_core/u_execute/u_register_bank/n4955 ,
         \u_a23_core/u_execute/u_register_bank/n4953 ,
         \u_a23_core/u_execute/u_register_bank/n4951 ,
         \u_a23_core/u_execute/u_register_bank/n4949 ,
         \u_a23_core/u_execute/u_register_bank/n4947 ,
         \u_a23_core/u_execute/u_register_bank/n4945 ,
         \u_a23_core/u_execute/u_register_bank/n4943 ,
         \u_a23_core/u_execute/u_register_bank/n4941 ,
         \u_a23_core/u_execute/u_register_bank/n4939 ,
         \u_a23_core/u_execute/u_register_bank/n4937 ,
         \u_a23_core/u_execute/u_register_bank/n4935 ,
         \u_a23_core/u_execute/u_register_bank/n4933 ,
         \u_a23_core/u_execute/u_register_bank/n4931 ,
         \u_a23_core/u_execute/u_register_bank/n4929 ,
         \u_a23_core/u_execute/u_register_bank/n4927 ,
         \u_a23_core/u_execute/u_register_bank/n4925 ,
         \u_a23_core/u_execute/u_register_bank/n4923 ,
         \u_a23_core/u_execute/u_register_bank/n4921 ,
         \u_a23_core/u_execute/u_register_bank/n4919 ,
         \u_a23_core/u_execute/u_register_bank/n4917 ,
         \u_a23_core/u_execute/u_register_bank/n4915 ,
         \u_a23_core/u_execute/u_register_bank/n4913 ,
         \u_a23_core/u_execute/u_register_bank/n4911 ,
         \u_a23_core/u_execute/u_register_bank/n4909 ,
         \u_a23_core/u_execute/u_register_bank/n4907 ,
         \u_a23_core/u_execute/u_register_bank/n4905 ,
         \u_a23_core/u_execute/u_register_bank/n4903 ,
         \u_a23_core/u_execute/u_register_bank/n4901 ,
         \u_a23_core/u_execute/u_register_bank/n4899 ,
         \u_a23_core/u_execute/u_register_bank/n4897 ,
         \u_a23_core/u_execute/u_register_bank/n4895 ,
         \u_a23_core/u_execute/u_register_bank/n4893 ,
         \u_a23_core/u_execute/u_register_bank/n4891 ,
         \u_a23_core/u_execute/u_register_bank/n4889 ,
         \u_a23_core/u_execute/u_register_bank/n4887 ,
         \u_a23_core/u_execute/u_register_bank/n4885 ,
         \u_a23_core/u_execute/u_register_bank/n4883 ,
         \u_a23_core/u_execute/u_register_bank/n4881 ,
         \u_a23_core/u_execute/u_register_bank/n4879 ,
         \u_a23_core/u_execute/u_register_bank/n4877 ,
         \u_a23_core/u_execute/u_register_bank/n4875 ,
         \u_a23_core/u_execute/u_register_bank/n4873 ,
         \u_a23_core/u_execute/u_register_bank/n4871 ,
         \u_a23_core/u_execute/u_register_bank/n4869 ,
         \u_a23_core/u_execute/u_register_bank/n4867 ,
         \u_a23_core/u_execute/u_register_bank/n4865 ,
         \u_a23_core/u_execute/u_register_bank/n4863 ,
         \u_a23_core/u_execute/u_register_bank/n4861 ,
         \u_a23_core/u_execute/u_register_bank/n4859 ,
         \u_a23_core/u_execute/u_register_bank/n4857 ,
         \u_a23_core/u_execute/u_register_bank/n4855 ,
         \u_a23_core/u_execute/u_register_bank/n4853 ,
         \u_a23_core/u_execute/u_register_bank/n4851 ,
         \u_a23_core/u_execute/u_register_bank/n4849 ,
         \u_a23_core/u_execute/u_register_bank/n4847 ,
         \u_a23_core/u_execute/u_register_bank/n4845 ,
         \u_a23_core/u_execute/u_register_bank/n4843 ,
         \u_a23_core/u_execute/u_register_bank/n4841 ,
         \u_a23_core/u_execute/u_register_bank/n4839 ,
         \u_a23_core/u_execute/u_register_bank/n4837 ,
         \u_a23_core/u_execute/u_register_bank/n4835 ,
         \u_a23_core/u_execute/u_register_bank/n4833 ,
         \u_a23_core/u_execute/u_register_bank/n4831 ,
         \u_a23_core/u_execute/u_register_bank/n4829 ,
         \u_a23_core/u_execute/u_register_bank/n4827 ,
         \u_a23_core/u_execute/u_register_bank/n4825 ,
         \u_a23_core/u_execute/u_register_bank/n4823 ,
         \u_a23_core/u_execute/u_register_bank/n4821 ,
         \u_a23_core/u_execute/u_register_bank/n4819 ,
         \u_a23_core/u_execute/u_register_bank/n4817 ,
         \u_a23_core/u_execute/u_register_bank/n4815 ,
         \u_a23_core/u_execute/u_register_bank/n4813 ,
         \u_a23_core/u_execute/u_register_bank/n4811 ,
         \u_a23_core/u_execute/u_register_bank/n4809 ,
         \u_a23_core/u_execute/u_register_bank/n4807 ,
         \u_a23_core/u_execute/u_register_bank/n4805 ,
         \u_a23_core/u_execute/u_register_bank/n4803 ,
         \u_a23_core/u_execute/u_register_bank/n4801 ,
         \u_a23_core/u_execute/u_register_bank/n4799 ,
         \u_a23_core/u_execute/u_register_bank/n4797 ,
         \u_a23_core/u_execute/u_register_bank/n4795 ,
         \u_a23_core/u_execute/u_register_bank/n4793 ,
         \u_a23_core/u_execute/u_register_bank/n4791 ,
         \u_a23_core/u_execute/u_register_bank/n4789 ,
         \u_a23_core/u_execute/u_register_bank/n4787 ,
         \u_a23_core/u_execute/u_register_bank/n4785 ,
         \u_a23_core/u_execute/u_register_bank/n4783 ,
         \u_a23_core/u_execute/u_register_bank/n4781 ,
         \u_a23_core/u_execute/u_register_bank/n4779 ,
         \u_a23_core/u_execute/u_register_bank/n4777 ,
         \u_a23_core/u_execute/u_register_bank/n4775 ,
         \u_a23_core/u_execute/u_register_bank/n4773 ,
         \u_a23_core/u_execute/u_register_bank/n4771 ,
         \u_a23_core/u_execute/u_register_bank/n4769 ,
         \u_a23_core/u_execute/u_register_bank/n4767 ,
         \u_a23_core/u_execute/u_register_bank/n4765 ,
         \u_a23_core/u_execute/u_register_bank/n4763 ,
         \u_a23_core/u_execute/u_register_bank/n4761 ,
         \u_a23_core/u_execute/u_register_bank/n4759 ,
         \u_a23_core/u_execute/u_register_bank/n4757 ,
         \u_a23_core/u_execute/u_register_bank/n4755 ,
         \u_a23_core/u_execute/u_register_bank/n4753 ,
         \u_a23_core/u_execute/u_register_bank/n4751 ,
         \u_a23_core/u_execute/u_register_bank/n4749 ,
         \u_a23_core/u_execute/u_register_bank/n4747 ,
         \u_a23_core/u_execute/u_register_bank/n4745 ,
         \u_a23_core/u_execute/u_register_bank/n4743 ,
         \u_a23_core/u_execute/u_register_bank/n4741 ,
         \u_a23_core/u_execute/u_register_bank/n4739 ,
         \u_a23_core/u_execute/u_register_bank/n4737 ,
         \u_a23_core/u_execute/u_register_bank/n4735 ,
         \u_a23_core/u_execute/u_register_bank/n4733 ,
         \u_a23_core/u_execute/u_register_bank/n4731 ,
         \u_a23_core/u_execute/u_register_bank/n4729 ,
         \u_a23_core/u_execute/u_register_bank/n4727 ,
         \u_a23_core/u_execute/u_register_bank/n4725 ,
         \u_a23_core/u_execute/u_register_bank/n4723 ,
         \u_a23_core/u_execute/u_register_bank/n4721 ,
         \u_a23_core/u_execute/u_register_bank/n4719 ,
         \u_a23_core/u_execute/u_register_bank/n4717 ,
         \u_a23_core/u_execute/u_register_bank/n4715 ,
         \u_a23_core/u_execute/u_register_bank/n4713 ,
         \u_a23_core/u_execute/u_register_bank/n4711 ,
         \u_a23_core/u_execute/u_register_bank/n4709 ,
         \u_a23_core/u_execute/u_register_bank/n4707 ,
         \u_a23_core/u_execute/u_register_bank/n4705 ,
         \u_a23_core/u_execute/u_register_bank/n4703 ,
         \u_a23_core/u_execute/u_register_bank/n4701 ,
         \u_a23_core/u_execute/u_register_bank/n4699 ,
         \u_a23_core/u_execute/u_register_bank/n4697 ,
         \u_a23_core/u_execute/u_register_bank/n4695 ,
         \u_a23_core/u_execute/u_register_bank/n4693 ,
         \u_a23_core/u_execute/u_register_bank/n4691 ,
         \u_a23_core/u_execute/u_register_bank/n4689 ,
         \u_a23_core/u_execute/u_register_bank/n4687 ,
         \u_a23_core/u_execute/u_register_bank/n4685 ,
         \u_a23_core/u_execute/u_register_bank/n4683 ,
         \u_a23_core/u_execute/u_register_bank/n4681 ,
         \u_a23_core/u_execute/u_register_bank/n4679 ,
         \u_a23_core/u_execute/u_register_bank/n4677 ,
         \u_a23_core/u_execute/u_register_bank/n4675 ,
         \u_a23_core/u_execute/u_register_bank/n4673 ,
         \u_a23_core/u_execute/u_register_bank/n4671 ,
         \u_a23_core/u_execute/u_register_bank/n4669 ,
         \u_a23_core/u_execute/u_register_bank/n4667 ,
         \u_a23_core/u_execute/u_register_bank/n4665 ,
         \u_a23_core/u_execute/u_register_bank/n4663 ,
         \u_a23_core/u_execute/u_register_bank/n4661 ,
         \u_a23_core/u_execute/u_register_bank/n4659 ,
         \u_a23_core/u_execute/u_register_bank/n4657 ,
         \u_a23_core/u_execute/u_register_bank/n4655 ,
         \u_a23_core/u_execute/u_register_bank/n4653 ,
         \u_a23_core/u_execute/u_register_bank/n4651 ,
         \u_a23_core/u_execute/u_register_bank/n4649 ,
         \u_a23_core/u_execute/u_register_bank/n4647 ,
         \u_a23_core/u_execute/u_register_bank/n4645 ,
         \u_a23_core/u_execute/u_register_bank/n4643 ,
         \u_a23_core/u_execute/u_register_bank/n4641 ,
         \u_a23_core/u_execute/u_register_bank/n4639 ,
         \u_a23_core/u_execute/u_register_bank/n4637 ,
         \u_a23_core/u_execute/u_register_bank/n4635 ,
         \u_a23_core/u_execute/u_register_bank/n4633 ,
         \u_a23_core/u_execute/u_register_bank/n4631 ,
         \u_a23_core/u_execute/u_register_bank/n4629 ,
         \u_a23_core/u_execute/u_register_bank/n4627 ,
         \u_a23_core/u_execute/u_register_bank/n4625 ,
         \u_a23_core/u_execute/u_register_bank/n4623 ,
         \u_a23_core/u_execute/u_register_bank/n4621 ,
         \u_a23_core/u_execute/u_register_bank/n4619 ,
         \u_a23_core/u_execute/u_register_bank/n4617 ,
         \u_a23_core/u_execute/u_register_bank/n4615 ,
         \u_a23_core/u_execute/u_register_bank/n4613 ,
         \u_a23_core/u_execute/u_register_bank/n4611 ,
         \u_a23_core/u_execute/u_register_bank/n4609 ,
         \u_a23_core/u_execute/u_register_bank/n4607 ,
         \u_a23_core/u_execute/u_register_bank/n4605 ,
         \u_a23_core/u_execute/u_register_bank/n4603 ,
         \u_a23_core/u_execute/u_register_bank/n4601 ,
         \u_a23_core/u_execute/u_register_bank/n4599 ,
         \u_a23_core/u_execute/u_register_bank/n4597 ,
         \u_a23_core/u_execute/u_register_bank/n4595 ,
         \u_a23_core/u_execute/u_register_bank/n4593 ,
         \u_a23_core/u_execute/u_register_bank/n4591 ,
         \u_a23_core/u_execute/u_register_bank/n4589 ,
         \u_a23_core/u_execute/u_register_bank/n4587 ,
         \u_a23_core/u_execute/u_register_bank/n4585 ,
         \u_a23_core/u_execute/u_register_bank/n4583 ,
         \u_a23_core/u_execute/u_register_bank/n4581 ,
         \u_a23_core/u_execute/u_register_bank/n4579 ,
         \u_a23_core/u_execute/u_register_bank/n4577 ,
         \u_a23_core/u_execute/u_register_bank/n4575 ,
         \u_a23_core/u_execute/u_register_bank/n4573 ,
         \u_a23_core/u_execute/u_register_bank/n4571 ,
         \u_a23_core/u_execute/u_register_bank/n4569 ,
         \u_a23_core/u_execute/u_register_bank/n4567 ,
         \u_a23_core/u_execute/u_register_bank/n4565 ,
         \u_a23_core/u_execute/u_register_bank/n4563 ,
         \u_a23_core/u_execute/u_register_bank/n4561 ,
         \u_a23_core/u_execute/u_register_bank/n4559 ,
         \u_a23_core/u_execute/u_register_bank/n4557 ,
         \u_a23_core/u_execute/u_register_bank/n4555 ,
         \u_a23_core/u_execute/u_register_bank/n4553 ,
         \u_a23_core/u_execute/u_register_bank/n4551 ,
         \u_a23_core/u_execute/u_register_bank/n4549 ,
         \u_a23_core/u_execute/u_register_bank/n4547 ,
         \u_a23_core/u_execute/u_register_bank/n4545 ,
         \u_a23_core/u_execute/u_register_bank/n4543 ,
         \u_a23_core/u_execute/u_register_bank/n4541 ,
         \u_a23_core/u_execute/u_register_bank/n4539 ,
         \u_a23_core/u_execute/u_register_bank/n4537 ,
         \u_a23_core/u_execute/u_register_bank/n4535 ,
         \u_a23_core/u_execute/u_register_bank/n4533 ,
         \u_a23_core/u_execute/u_register_bank/n4531 ,
         \u_a23_core/u_execute/u_register_bank/n4529 ,
         \u_a23_core/u_execute/u_register_bank/n4527 ,
         \u_a23_core/u_execute/u_register_bank/n4525 ,
         \u_a23_core/u_execute/u_register_bank/n4523 ,
         \u_a23_core/u_execute/u_register_bank/n4521 ,
         \u_a23_core/u_execute/u_register_bank/n4519 ,
         \u_a23_core/u_execute/u_register_bank/n4517 ,
         \u_a23_core/u_execute/u_register_bank/n4515 ,
         \u_a23_core/u_execute/u_register_bank/n4513 ,
         \u_a23_core/u_execute/u_register_bank/n4511 ,
         \u_a23_core/u_execute/u_register_bank/n4509 ,
         \u_a23_core/u_execute/u_register_bank/n4507 ,
         \u_a23_core/u_execute/u_register_bank/n4505 ,
         \u_a23_core/u_execute/u_register_bank/n4503 ,
         \u_a23_core/u_execute/u_register_bank/n4501 ,
         \u_a23_core/u_execute/u_register_bank/n4499 ,
         \u_a23_core/u_execute/u_register_bank/n4497 ,
         \u_a23_core/u_execute/u_register_bank/n4495 ,
         \u_a23_core/u_execute/u_register_bank/n4493 ,
         \u_a23_core/u_execute/u_register_bank/n4491 ,
         \u_a23_core/u_execute/u_register_bank/n4489 ,
         \u_a23_core/u_execute/u_register_bank/n4487 ,
         \u_a23_core/u_execute/u_register_bank/n4485 ,
         \u_a23_core/u_execute/u_register_bank/n4483 ,
         \u_a23_core/u_execute/u_register_bank/n4481 ,
         \u_a23_core/u_execute/u_register_bank/n4479 ,
         \u_a23_core/u_execute/u_register_bank/n4477 ,
         \u_a23_core/u_execute/u_register_bank/n4475 ,
         \u_a23_core/u_execute/u_register_bank/n4473 ,
         \u_a23_core/u_execute/u_register_bank/n4471 ,
         \u_a23_core/u_execute/u_register_bank/n4469 ,
         \u_a23_core/u_execute/u_register_bank/n4467 ,
         \u_a23_core/u_execute/u_register_bank/n4465 ,
         \u_a23_core/u_execute/u_register_bank/n4463 ,
         \u_a23_core/u_execute/u_register_bank/n4461 ,
         \u_a23_core/u_execute/u_register_bank/n4459 ,
         \u_a23_core/u_execute/u_register_bank/n4457 ,
         \u_a23_core/u_execute/u_register_bank/n4455 ,
         \u_a23_core/u_execute/u_register_bank/n4453 ,
         \u_a23_core/u_execute/u_register_bank/n4451 ,
         \u_a23_core/u_execute/u_register_bank/n4449 ,
         \u_a23_core/u_execute/u_register_bank/n4447 ,
         \u_a23_core/u_execute/u_register_bank/n4445 ,
         \u_a23_core/u_execute/u_register_bank/n4443 ,
         \u_a23_core/u_execute/u_register_bank/n4441 ,
         \u_a23_core/u_execute/u_register_bank/n4439 ,
         \u_a23_core/u_execute/u_register_bank/n4437 ,
         \u_a23_core/u_execute/u_register_bank/n4435 ,
         \u_a23_core/u_execute/u_register_bank/n4433 ,
         \u_a23_core/u_execute/u_register_bank/n4431 ,
         \u_a23_core/u_execute/u_register_bank/n4429 ,
         \u_a23_core/u_execute/u_register_bank/n4427 ,
         \u_a23_core/u_execute/u_register_bank/n4425 ,
         \u_a23_core/u_execute/u_register_bank/n4423 ,
         \u_a23_core/u_execute/u_register_bank/n4421 ,
         \u_a23_core/u_execute/u_register_bank/n4419 ,
         \u_a23_core/u_execute/u_register_bank/n4417 ,
         \u_a23_core/u_execute/u_register_bank/n4415 ,
         \u_a23_core/u_execute/u_register_bank/n4413 ,
         \u_a23_core/u_execute/u_register_bank/n4411 ,
         \u_a23_core/u_execute/u_register_bank/n4409 ,
         \u_a23_core/u_execute/u_register_bank/n4407 ,
         \u_a23_core/u_execute/u_register_bank/n4405 ,
         \u_a23_core/u_execute/u_register_bank/n4403 ,
         \u_a23_core/u_execute/u_register_bank/n4401 ,
         \u_a23_core/u_execute/u_register_bank/n4399 ,
         \u_a23_core/u_execute/u_register_bank/n4397 ,
         \u_a23_core/u_execute/u_register_bank/n4395 ,
         \u_a23_core/u_execute/u_register_bank/n4393 ,
         \u_a23_core/u_execute/u_register_bank/n4391 ,
         \u_a23_core/u_execute/u_register_bank/n4389 ,
         \u_a23_core/u_execute/u_register_bank/n4387 ,
         \u_a23_core/u_execute/u_register_bank/n4385 ,
         \u_a23_core/u_execute/u_register_bank/n4383 ,
         \u_a23_core/u_execute/u_register_bank/n4381 ,
         \u_a23_core/u_execute/u_register_bank/n4379 ,
         \u_a23_core/u_execute/u_register_bank/n4377 ,
         \u_a23_core/u_execute/u_register_bank/n4375 ,
         \u_a23_core/u_execute/u_register_bank/n4373 ,
         \u_a23_core/u_execute/u_register_bank/n4371 ,
         \u_a23_core/u_execute/u_register_bank/n4369 ,
         \u_a23_core/u_execute/u_register_bank/n4367 ,
         \u_a23_core/u_execute/u_register_bank/n4365 ,
         \u_a23_core/u_execute/u_register_bank/n4363 ,
         \u_a23_core/u_execute/u_register_bank/n4361 ,
         \u_a23_core/u_execute/u_register_bank/n4359 ,
         \u_a23_core/u_execute/u_register_bank/n4357 ,
         \u_a23_core/u_execute/u_register_bank/n4355 ,
         \u_a23_core/u_execute/u_register_bank/n4353 ,
         \u_a23_core/u_execute/u_register_bank/n4351 ,
         \u_a23_core/u_execute/u_register_bank/n4349 ,
         \u_a23_core/u_execute/u_register_bank/n4347 ,
         \u_a23_core/u_execute/u_register_bank/n4345 ,
         \u_a23_core/u_execute/u_register_bank/n4343 ,
         \u_a23_core/u_execute/u_register_bank/n4341 ,
         \u_a23_core/u_execute/u_register_bank/n4339 ,
         \u_a23_core/u_execute/u_register_bank/n4337 ,
         \u_a23_core/u_execute/u_register_bank/n4335 ,
         \u_a23_core/u_execute/u_register_bank/n4333 ,
         \u_a23_core/u_execute/u_register_bank/n4331 ,
         \u_a23_core/u_execute/u_register_bank/n4329 ,
         \u_a23_core/u_execute/u_register_bank/n4327 ,
         \u_a23_core/u_execute/u_register_bank/n4325 ,
         \u_a23_core/u_execute/u_register_bank/n4323 ,
         \u_a23_core/u_execute/u_register_bank/n4321 ,
         \u_a23_core/u_execute/u_register_bank/n4319 ,
         \u_a23_core/u_execute/u_register_bank/n4317 ,
         \u_a23_core/u_execute/u_register_bank/n4315 ,
         \u_a23_core/u_execute/u_register_bank/n4313 ,
         \u_a23_core/u_execute/u_register_bank/n4311 ,
         \u_a23_core/u_execute/u_register_bank/n4309 ,
         \u_a23_core/u_execute/u_register_bank/n4307 ,
         \u_a23_core/u_execute/u_register_bank/n4305 ,
         \u_a23_core/u_execute/u_register_bank/n4303 ,
         \u_a23_core/u_execute/u_register_bank/n4301 ,
         \u_a23_core/u_execute/u_register_bank/n4299 ,
         \u_a23_core/u_execute/u_register_bank/n4297 ,
         \u_a23_core/u_execute/u_register_bank/n4295 ,
         \u_a23_core/u_execute/u_register_bank/n4293 ,
         \u_a23_core/u_execute/u_register_bank/n4291 ,
         \u_a23_core/u_execute/u_register_bank/n4289 ,
         \u_a23_core/u_execute/u_register_bank/n4287 ,
         \u_a23_core/u_execute/u_register_bank/n4285 ,
         \u_a23_core/u_execute/u_register_bank/n4283 ,
         \u_a23_core/u_execute/u_register_bank/n4281 ,
         \u_a23_core/u_execute/u_register_bank/n4279 ,
         \u_a23_core/u_execute/u_register_bank/n4277 ,
         \u_a23_core/u_execute/u_register_bank/n4275 ,
         \u_a23_core/u_execute/u_register_bank/n4273 ,
         \u_a23_core/u_execute/u_register_bank/n4271 ,
         \u_a23_core/u_execute/u_register_bank/n4269 ,
         \u_a23_core/u_execute/u_register_bank/n4267 ,
         \u_a23_core/u_execute/u_register_bank/n4265 ,
         \u_a23_core/u_execute/u_register_bank/n4263 ,
         \u_a23_core/u_execute/u_register_bank/n4261 ,
         \u_a23_core/u_execute/u_register_bank/n4259 ,
         \u_a23_core/u_execute/u_register_bank/n4257 ,
         \u_a23_core/u_execute/u_register_bank/n4255 ,
         \u_a23_core/u_execute/u_register_bank/n4253 ,
         \u_a23_core/u_execute/u_register_bank/n4251 ,
         \u_a23_core/u_execute/u_register_bank/n4249 ,
         \u_a23_core/u_execute/u_register_bank/n4247 ,
         \u_a23_core/u_execute/u_register_bank/n4245 ,
         \u_a23_core/u_execute/u_register_bank/n4243 ,
         \u_a23_core/u_execute/u_register_bank/n4241 ,
         \u_a23_core/u_execute/u_register_bank/n4239 ,
         \u_a23_core/u_execute/u_register_bank/n4237 ,
         \u_a23_core/u_execute/u_register_bank/n4235 ,
         \u_a23_core/u_execute/u_register_bank/n4233 ,
         \u_a23_core/u_execute/u_register_bank/n4231 ,
         \u_a23_core/u_execute/u_register_bank/n4229 ,
         \u_a23_core/u_execute/u_register_bank/n4227 ,
         \u_a23_core/u_execute/u_register_bank/n4225 ,
         \u_a23_core/u_execute/u_register_bank/n4223 ,
         \u_a23_core/u_execute/u_register_bank/n4221 ,
         \u_a23_core/u_execute/u_register_bank/n4219 ,
         \u_a23_core/u_execute/u_register_bank/n4217 ,
         \u_a23_core/u_execute/u_register_bank/n4215 ,
         \u_a23_core/u_execute/u_register_bank/n4213 ,
         \u_a23_core/u_execute/u_register_bank/n4211 ,
         \u_a23_core/u_execute/u_register_bank/n4209 ,
         \u_a23_core/u_execute/u_register_bank/n4207 ,
         \u_a23_core/u_execute/u_register_bank/n4205 ,
         \u_a23_core/u_execute/u_register_bank/n4203 ,
         \u_a23_core/u_execute/u_register_bank/n4201 ,
         \u_a23_core/u_execute/u_register_bank/n4199 ,
         \u_a23_core/u_execute/u_register_bank/n4197 ,
         \u_a23_core/u_execute/u_register_bank/n4195 ,
         \u_a23_core/u_execute/u_register_bank/n4193 ,
         \u_a23_core/u_execute/u_register_bank/n4191 ,
         \u_a23_core/u_execute/u_register_bank/n4189 ,
         \u_a23_core/u_execute/u_register_bank/n4187 ,
         \u_a23_core/u_execute/u_register_bank/n4185 ,
         \u_a23_core/u_execute/u_register_bank/n4183 ,
         \u_a23_core/u_execute/u_register_bank/n4181 ,
         \u_a23_core/u_execute/u_register_bank/n4179 ,
         \u_a23_core/u_execute/u_register_bank/n4177 ,
         \u_a23_core/u_execute/u_register_bank/n4175 ,
         \u_a23_core/u_execute/u_register_bank/n4173 ,
         \u_a23_core/u_execute/u_register_bank/n4171 ,
         \u_a23_core/u_execute/u_register_bank/n4169 ,
         \u_a23_core/u_execute/u_register_bank/n4167 ,
         \u_a23_core/u_execute/u_register_bank/n4165 ,
         \u_a23_core/u_execute/u_register_bank/n4163 ,
         \u_a23_core/u_execute/u_register_bank/n4161 ,
         \u_a23_core/u_execute/u_register_bank/n4159 ,
         \u_a23_core/u_execute/u_register_bank/n4157 ,
         \u_a23_core/u_execute/u_register_bank/n4155 ,
         \u_a23_core/u_execute/u_register_bank/n4153 ,
         \u_a23_core/u_execute/u_register_bank/n4151 ,
         \u_a23_core/u_execute/u_register_bank/n4149 ,
         \u_a23_core/u_execute/u_register_bank/n4147 ,
         \u_a23_core/u_execute/u_register_bank/n4145 ,
         \u_a23_core/u_execute/u_register_bank/n4143 ,
         \u_a23_core/u_execute/u_register_bank/n4141 ,
         \u_a23_core/u_execute/u_register_bank/n4139 ,
         \u_a23_core/u_execute/u_register_bank/n4137 ,
         \u_a23_core/u_execute/u_register_bank/n4135 ,
         \u_a23_core/u_execute/u_register_bank/n4133 ,
         \u_a23_core/u_execute/u_register_bank/n4131 ,
         \u_a23_core/u_execute/u_register_bank/n4129 ,
         \u_a23_core/u_execute/u_register_bank/n4127 ,
         \u_a23_core/u_execute/u_register_bank/n4125 ,
         \u_a23_core/u_execute/u_register_bank/n4123 ,
         \u_a23_core/u_execute/u_register_bank/n4121 ,
         \u_a23_core/u_execute/u_register_bank/n4119 ,
         \u_a23_core/u_execute/u_register_bank/n4117 ,
         \u_a23_core/u_execute/u_register_bank/n4115 ,
         \u_a23_core/u_execute/u_register_bank/n4113 ,
         \u_a23_core/u_execute/u_register_bank/n4111 ,
         \u_a23_core/u_execute/u_register_bank/n4109 ,
         \u_a23_core/u_execute/u_register_bank/n4107 ,
         \u_a23_core/u_execute/u_register_bank/n4105 ,
         \u_a23_core/u_execute/u_register_bank/n4103 ,
         \u_a23_core/u_execute/u_register_bank/n4101 ,
         \u_a23_core/u_execute/u_register_bank/n4099 ,
         \u_a23_core/u_execute/u_register_bank/n4097 ,
         \u_a23_core/u_execute/u_register_bank/n4095 ,
         \u_a23_core/u_execute/u_register_bank/n4093 ,
         \u_a23_core/u_execute/u_register_bank/n4091 ,
         \u_a23_core/u_execute/u_register_bank/n4089 ,
         \u_a23_core/u_execute/u_register_bank/n4087 ,
         \u_a23_core/u_execute/u_register_bank/n4085 ,
         \u_a23_core/u_execute/u_register_bank/n4083 ,
         \u_a23_core/u_execute/u_register_bank/n4081 ,
         \u_a23_core/u_execute/u_register_bank/n4079 ,
         \u_a23_core/u_execute/u_register_bank/n4077 ,
         \u_a23_core/u_execute/u_register_bank/n4075 ,
         \u_a23_core/u_execute/u_register_bank/n4073 ,
         \u_a23_core/u_execute/u_register_bank/n4071 ,
         \u_a23_core/u_execute/u_register_bank/n4069 ,
         \u_a23_core/u_execute/u_register_bank/n4067 ,
         \u_a23_core/u_execute/u_register_bank/n4065 ,
         \u_a23_core/u_execute/u_register_bank/n4063 ,
         \u_a23_core/u_execute/u_register_bank/n4061 ,
         \u_a23_core/u_execute/u_register_bank/n4059 ,
         \u_a23_core/u_execute/u_register_bank/n4057 ,
         \u_a23_core/u_execute/u_register_bank/n4055 ,
         \u_a23_core/u_execute/u_register_bank/n4053 ,
         \u_a23_core/u_execute/u_register_bank/n4051 ,
         \u_a23_core/u_execute/u_register_bank/n4049 ,
         \u_a23_core/u_execute/u_register_bank/n4047 ,
         \u_a23_core/u_execute/u_register_bank/n4045 ,
         \u_a23_core/u_execute/u_register_bank/n4043 ,
         \u_a23_core/u_execute/u_register_bank/n4041 ,
         \u_a23_core/u_execute/u_register_bank/n4039 ,
         \u_a23_core/u_execute/u_register_bank/n4037 ,
         \u_a23_core/u_execute/u_register_bank/n4035 ,
         \u_a23_core/u_execute/u_register_bank/n4033 ,
         \u_a23_core/u_execute/u_register_bank/n4031 ,
         \u_a23_core/u_execute/u_register_bank/n4029 ,
         \u_a23_core/u_execute/u_register_bank/n4027 ,
         \u_a23_core/u_execute/u_register_bank/n4025 ,
         \u_a23_core/u_execute/u_register_bank/n4023 ,
         \u_a23_core/u_execute/u_register_bank/n4021 ,
         \u_a23_core/u_execute/u_register_bank/n4019 ,
         \u_a23_core/u_execute/u_register_bank/n4017 ,
         \u_a23_core/u_execute/u_register_bank/n4015 ,
         \u_a23_core/u_execute/u_register_bank/n4013 ,
         \u_a23_core/u_execute/u_register_bank/n4011 ,
         \u_a23_core/u_execute/u_register_bank/n4009 ,
         \u_a23_core/u_execute/u_register_bank/n4007 ,
         \u_a23_core/u_execute/u_register_bank/n4005 ,
         \u_a23_core/u_execute/u_register_bank/n4003 ,
         \u_a23_core/u_execute/u_register_bank/n4001 ,
         \u_a23_core/u_execute/u_register_bank/n3999 ,
         \u_a23_core/u_execute/u_register_bank/n3997 ,
         \u_a23_core/u_execute/u_register_bank/n3995 ,
         \u_a23_core/u_execute/u_register_bank/n3993 ,
         \u_a23_core/u_execute/u_register_bank/n3991 ,
         \u_a23_core/u_execute/u_register_bank/n3989 ,
         \u_a23_core/u_execute/u_register_bank/n3987 ,
         \u_a23_core/u_execute/u_register_bank/n3985 ,
         \u_a23_core/u_execute/u_register_bank/n3983 ,
         \u_a23_core/u_execute/u_register_bank/n3981 ,
         \u_a23_core/u_execute/u_register_bank/n3979 ,
         \u_a23_core/u_execute/u_register_bank/n3977 ,
         \u_a23_core/u_execute/u_register_bank/n3975 ,
         \u_a23_core/u_execute/u_register_bank/r14[0] ,
         \u_a23_core/u_execute/u_register_bank/r14[1] ,
         \u_a23_core/u_execute/u_register_bank/r14[2] ,
         \u_a23_core/u_execute/u_register_bank/r14[3] ,
         \u_a23_core/u_execute/u_register_bank/r14[4] ,
         \u_a23_core/u_execute/u_register_bank/r14[5] ,
         \u_a23_core/u_execute/u_register_bank/r14[6] ,
         \u_a23_core/u_execute/u_register_bank/r14[7] ,
         \u_a23_core/u_execute/u_register_bank/r14[8] ,
         \u_a23_core/u_execute/u_register_bank/r14[9] ,
         \u_a23_core/u_execute/u_register_bank/r14[10] ,
         \u_a23_core/u_execute/u_register_bank/r14[11] ,
         \u_a23_core/u_execute/u_register_bank/r14[12] ,
         \u_a23_core/u_execute/u_register_bank/r14[13] ,
         \u_a23_core/u_execute/u_register_bank/r14[14] ,
         \u_a23_core/u_execute/u_register_bank/r14[15] ,
         \u_a23_core/u_execute/u_register_bank/r14[16] ,
         \u_a23_core/u_execute/u_register_bank/r14[17] ,
         \u_a23_core/u_execute/u_register_bank/r14[18] ,
         \u_a23_core/u_execute/u_register_bank/r14[19] ,
         \u_a23_core/u_execute/u_register_bank/r14[20] ,
         \u_a23_core/u_execute/u_register_bank/r14[21] ,
         \u_a23_core/u_execute/u_register_bank/r14[22] ,
         \u_a23_core/u_execute/u_register_bank/r14[23] ,
         \u_a23_core/u_execute/u_register_bank/r14[24] ,
         \u_a23_core/u_execute/u_register_bank/r14[25] ,
         \u_a23_core/u_execute/u_register_bank/r14[26] ,
         \u_a23_core/u_execute/u_register_bank/r14[27] ,
         \u_a23_core/u_execute/u_register_bank/r14[28] ,
         \u_a23_core/u_execute/u_register_bank/r14[29] ,
         \u_a23_core/u_execute/u_register_bank/r14[30] ,
         \u_a23_core/u_execute/u_register_bank/r14[31] ,
         \u_a23_core/u_execute/u_register_bank/r13[0] ,
         \u_a23_core/u_execute/u_register_bank/r13[1] ,
         \u_a23_core/u_execute/u_register_bank/r13[2] ,
         \u_a23_core/u_execute/u_register_bank/r13[3] ,
         \u_a23_core/u_execute/u_register_bank/r13[4] ,
         \u_a23_core/u_execute/u_register_bank/r13[5] ,
         \u_a23_core/u_execute/u_register_bank/r13[6] ,
         \u_a23_core/u_execute/u_register_bank/r13[7] ,
         \u_a23_core/u_execute/u_register_bank/r13[8] ,
         \u_a23_core/u_execute/u_register_bank/r13[9] ,
         \u_a23_core/u_execute/u_register_bank/r13[10] ,
         \u_a23_core/u_execute/u_register_bank/r13[11] ,
         \u_a23_core/u_execute/u_register_bank/r13[12] ,
         \u_a23_core/u_execute/u_register_bank/r13[13] ,
         \u_a23_core/u_execute/u_register_bank/r13[14] ,
         \u_a23_core/u_execute/u_register_bank/r13[15] ,
         \u_a23_core/u_execute/u_register_bank/r13[16] ,
         \u_a23_core/u_execute/u_register_bank/r13[17] ,
         \u_a23_core/u_execute/u_register_bank/r13[18] ,
         \u_a23_core/u_execute/u_register_bank/r13[19] ,
         \u_a23_core/u_execute/u_register_bank/r13[20] ,
         \u_a23_core/u_execute/u_register_bank/r13[21] ,
         \u_a23_core/u_execute/u_register_bank/r13[22] ,
         \u_a23_core/u_execute/u_register_bank/r13[23] ,
         \u_a23_core/u_execute/u_register_bank/r13[24] ,
         \u_a23_core/u_execute/u_register_bank/r13[25] ,
         \u_a23_core/u_execute/u_register_bank/r13[26] ,
         \u_a23_core/u_execute/u_register_bank/r13[27] ,
         \u_a23_core/u_execute/u_register_bank/r13[28] ,
         \u_a23_core/u_execute/u_register_bank/r13[29] ,
         \u_a23_core/u_execute/u_register_bank/r13[30] ,
         \u_a23_core/u_execute/u_register_bank/r13[31] ,
         \u_a23_core/u_execute/u_register_bank/r12[0] ,
         \u_a23_core/u_execute/u_register_bank/r12[1] ,
         \u_a23_core/u_execute/u_register_bank/r12[2] ,
         \u_a23_core/u_execute/u_register_bank/r12[3] ,
         \u_a23_core/u_execute/u_register_bank/r12[4] ,
         \u_a23_core/u_execute/u_register_bank/r12[5] ,
         \u_a23_core/u_execute/u_register_bank/r12[6] ,
         \u_a23_core/u_execute/u_register_bank/r12[7] ,
         \u_a23_core/u_execute/u_register_bank/r12[8] ,
         \u_a23_core/u_execute/u_register_bank/r12[9] ,
         \u_a23_core/u_execute/u_register_bank/r12[10] ,
         \u_a23_core/u_execute/u_register_bank/r12[11] ,
         \u_a23_core/u_execute/u_register_bank/r12[12] ,
         \u_a23_core/u_execute/u_register_bank/r12[13] ,
         \u_a23_core/u_execute/u_register_bank/r12[14] ,
         \u_a23_core/u_execute/u_register_bank/r12[15] ,
         \u_a23_core/u_execute/u_register_bank/r12[16] ,
         \u_a23_core/u_execute/u_register_bank/r12[17] ,
         \u_a23_core/u_execute/u_register_bank/r12[18] ,
         \u_a23_core/u_execute/u_register_bank/r12[19] ,
         \u_a23_core/u_execute/u_register_bank/r12[20] ,
         \u_a23_core/u_execute/u_register_bank/r12[21] ,
         \u_a23_core/u_execute/u_register_bank/r12[22] ,
         \u_a23_core/u_execute/u_register_bank/r12[23] ,
         \u_a23_core/u_execute/u_register_bank/r12[24] ,
         \u_a23_core/u_execute/u_register_bank/r12[25] ,
         \u_a23_core/u_execute/u_register_bank/r12[26] ,
         \u_a23_core/u_execute/u_register_bank/r12[27] ,
         \u_a23_core/u_execute/u_register_bank/r12[28] ,
         \u_a23_core/u_execute/u_register_bank/r12[29] ,
         \u_a23_core/u_execute/u_register_bank/r12[30] ,
         \u_a23_core/u_execute/u_register_bank/r12[31] ,
         \u_a23_core/u_execute/u_register_bank/r11[0] ,
         \u_a23_core/u_execute/u_register_bank/r11[1] ,
         \u_a23_core/u_execute/u_register_bank/r11[2] ,
         \u_a23_core/u_execute/u_register_bank/r11[3] ,
         \u_a23_core/u_execute/u_register_bank/r11[4] ,
         \u_a23_core/u_execute/u_register_bank/r11[5] ,
         \u_a23_core/u_execute/u_register_bank/r11[6] ,
         \u_a23_core/u_execute/u_register_bank/r11[7] ,
         \u_a23_core/u_execute/u_register_bank/r11[8] ,
         \u_a23_core/u_execute/u_register_bank/r11[9] ,
         \u_a23_core/u_execute/u_register_bank/r11[10] ,
         \u_a23_core/u_execute/u_register_bank/r11[11] ,
         \u_a23_core/u_execute/u_register_bank/r11[12] ,
         \u_a23_core/u_execute/u_register_bank/r11[13] ,
         \u_a23_core/u_execute/u_register_bank/r11[14] ,
         \u_a23_core/u_execute/u_register_bank/r11[15] ,
         \u_a23_core/u_execute/u_register_bank/r11[16] ,
         \u_a23_core/u_execute/u_register_bank/r11[17] ,
         \u_a23_core/u_execute/u_register_bank/r11[18] ,
         \u_a23_core/u_execute/u_register_bank/r11[19] ,
         \u_a23_core/u_execute/u_register_bank/r11[20] ,
         \u_a23_core/u_execute/u_register_bank/r11[21] ,
         \u_a23_core/u_execute/u_register_bank/r11[22] ,
         \u_a23_core/u_execute/u_register_bank/r11[23] ,
         \u_a23_core/u_execute/u_register_bank/r11[24] ,
         \u_a23_core/u_execute/u_register_bank/r11[25] ,
         \u_a23_core/u_execute/u_register_bank/r11[26] ,
         \u_a23_core/u_execute/u_register_bank/r11[27] ,
         \u_a23_core/u_execute/u_register_bank/r11[28] ,
         \u_a23_core/u_execute/u_register_bank/r11[29] ,
         \u_a23_core/u_execute/u_register_bank/r11[30] ,
         \u_a23_core/u_execute/u_register_bank/r11[31] ,
         \u_a23_core/u_execute/u_register_bank/r10[0] ,
         \u_a23_core/u_execute/u_register_bank/r10[1] ,
         \u_a23_core/u_execute/u_register_bank/r10[2] ,
         \u_a23_core/u_execute/u_register_bank/r10[3] ,
         \u_a23_core/u_execute/u_register_bank/r10[4] ,
         \u_a23_core/u_execute/u_register_bank/r10[5] ,
         \u_a23_core/u_execute/u_register_bank/r10[6] ,
         \u_a23_core/u_execute/u_register_bank/r10[7] ,
         \u_a23_core/u_execute/u_register_bank/r10[8] ,
         \u_a23_core/u_execute/u_register_bank/r10[9] ,
         \u_a23_core/u_execute/u_register_bank/r10[10] ,
         \u_a23_core/u_execute/u_register_bank/r10[11] ,
         \u_a23_core/u_execute/u_register_bank/r10[12] ,
         \u_a23_core/u_execute/u_register_bank/r10[13] ,
         \u_a23_core/u_execute/u_register_bank/r10[14] ,
         \u_a23_core/u_execute/u_register_bank/r10[15] ,
         \u_a23_core/u_execute/u_register_bank/r10[16] ,
         \u_a23_core/u_execute/u_register_bank/r10[17] ,
         \u_a23_core/u_execute/u_register_bank/r10[18] ,
         \u_a23_core/u_execute/u_register_bank/r10[19] ,
         \u_a23_core/u_execute/u_register_bank/r10[20] ,
         \u_a23_core/u_execute/u_register_bank/r10[21] ,
         \u_a23_core/u_execute/u_register_bank/r10[22] ,
         \u_a23_core/u_execute/u_register_bank/r10[23] ,
         \u_a23_core/u_execute/u_register_bank/r10[24] ,
         \u_a23_core/u_execute/u_register_bank/r10[25] ,
         \u_a23_core/u_execute/u_register_bank/r10[26] ,
         \u_a23_core/u_execute/u_register_bank/r10[27] ,
         \u_a23_core/u_execute/u_register_bank/r10[28] ,
         \u_a23_core/u_execute/u_register_bank/r10[29] ,
         \u_a23_core/u_execute/u_register_bank/r10[30] ,
         \u_a23_core/u_execute/u_register_bank/r10[31] ,
         \u_a23_core/u_execute/u_register_bank/r9[0] ,
         \u_a23_core/u_execute/u_register_bank/r9[1] ,
         \u_a23_core/u_execute/u_register_bank/r9[2] ,
         \u_a23_core/u_execute/u_register_bank/r9[3] ,
         \u_a23_core/u_execute/u_register_bank/r9[4] ,
         \u_a23_core/u_execute/u_register_bank/r9[5] ,
         \u_a23_core/u_execute/u_register_bank/r9[6] ,
         \u_a23_core/u_execute/u_register_bank/r9[7] ,
         \u_a23_core/u_execute/u_register_bank/r9[8] ,
         \u_a23_core/u_execute/u_register_bank/r9[9] ,
         \u_a23_core/u_execute/u_register_bank/r9[10] ,
         \u_a23_core/u_execute/u_register_bank/r9[11] ,
         \u_a23_core/u_execute/u_register_bank/r9[12] ,
         \u_a23_core/u_execute/u_register_bank/r9[13] ,
         \u_a23_core/u_execute/u_register_bank/r9[14] ,
         \u_a23_core/u_execute/u_register_bank/r9[15] ,
         \u_a23_core/u_execute/u_register_bank/r9[16] ,
         \u_a23_core/u_execute/u_register_bank/r9[17] ,
         \u_a23_core/u_execute/u_register_bank/r9[18] ,
         \u_a23_core/u_execute/u_register_bank/r9[19] ,
         \u_a23_core/u_execute/u_register_bank/r9[20] ,
         \u_a23_core/u_execute/u_register_bank/r9[21] ,
         \u_a23_core/u_execute/u_register_bank/r9[22] ,
         \u_a23_core/u_execute/u_register_bank/r9[23] ,
         \u_a23_core/u_execute/u_register_bank/r9[24] ,
         \u_a23_core/u_execute/u_register_bank/r9[25] ,
         \u_a23_core/u_execute/u_register_bank/r9[26] ,
         \u_a23_core/u_execute/u_register_bank/r9[27] ,
         \u_a23_core/u_execute/u_register_bank/r9[28] ,
         \u_a23_core/u_execute/u_register_bank/r9[29] ,
         \u_a23_core/u_execute/u_register_bank/r9[30] ,
         \u_a23_core/u_execute/u_register_bank/r9[31] ,
         \u_a23_core/u_execute/u_register_bank/r8[0] ,
         \u_a23_core/u_execute/u_register_bank/r8[1] ,
         \u_a23_core/u_execute/u_register_bank/r8[2] ,
         \u_a23_core/u_execute/u_register_bank/r8[3] ,
         \u_a23_core/u_execute/u_register_bank/r8[4] ,
         \u_a23_core/u_execute/u_register_bank/r8[5] ,
         \u_a23_core/u_execute/u_register_bank/r8[6] ,
         \u_a23_core/u_execute/u_register_bank/r8[7] ,
         \u_a23_core/u_execute/u_register_bank/r8[8] ,
         \u_a23_core/u_execute/u_register_bank/r8[9] ,
         \u_a23_core/u_execute/u_register_bank/r8[10] ,
         \u_a23_core/u_execute/u_register_bank/r8[11] ,
         \u_a23_core/u_execute/u_register_bank/r8[12] ,
         \u_a23_core/u_execute/u_register_bank/r8[13] ,
         \u_a23_core/u_execute/u_register_bank/r8[14] ,
         \u_a23_core/u_execute/u_register_bank/r8[15] ,
         \u_a23_core/u_execute/u_register_bank/r8[16] ,
         \u_a23_core/u_execute/u_register_bank/r8[17] ,
         \u_a23_core/u_execute/u_register_bank/r8[18] ,
         \u_a23_core/u_execute/u_register_bank/r8[19] ,
         \u_a23_core/u_execute/u_register_bank/r8[20] ,
         \u_a23_core/u_execute/u_register_bank/r8[21] ,
         \u_a23_core/u_execute/u_register_bank/r8[22] ,
         \u_a23_core/u_execute/u_register_bank/r8[23] ,
         \u_a23_core/u_execute/u_register_bank/r8[24] ,
         \u_a23_core/u_execute/u_register_bank/r8[25] ,
         \u_a23_core/u_execute/u_register_bank/r8[26] ,
         \u_a23_core/u_execute/u_register_bank/r8[27] ,
         \u_a23_core/u_execute/u_register_bank/r8[28] ,
         \u_a23_core/u_execute/u_register_bank/r8[29] ,
         \u_a23_core/u_execute/u_register_bank/r8[30] ,
         \u_a23_core/u_execute/u_register_bank/r8[31] ,
         \u_a23_core/u_execute/u_register_bank/r7[0] ,
         \u_a23_core/u_execute/u_register_bank/r7[1] ,
         \u_a23_core/u_execute/u_register_bank/r7[2] ,
         \u_a23_core/u_execute/u_register_bank/r7[3] ,
         \u_a23_core/u_execute/u_register_bank/r7[4] ,
         \u_a23_core/u_execute/u_register_bank/r7[5] ,
         \u_a23_core/u_execute/u_register_bank/r7[6] ,
         \u_a23_core/u_execute/u_register_bank/r7[7] ,
         \u_a23_core/u_execute/u_register_bank/r7[8] ,
         \u_a23_core/u_execute/u_register_bank/r7[9] ,
         \u_a23_core/u_execute/u_register_bank/r7[10] ,
         \u_a23_core/u_execute/u_register_bank/r7[11] ,
         \u_a23_core/u_execute/u_register_bank/r7[12] ,
         \u_a23_core/u_execute/u_register_bank/r7[13] ,
         \u_a23_core/u_execute/u_register_bank/r7[14] ,
         \u_a23_core/u_execute/u_register_bank/r7[15] ,
         \u_a23_core/u_execute/u_register_bank/r7[16] ,
         \u_a23_core/u_execute/u_register_bank/r7[17] ,
         \u_a23_core/u_execute/u_register_bank/r7[18] ,
         \u_a23_core/u_execute/u_register_bank/r7[19] ,
         \u_a23_core/u_execute/u_register_bank/r7[20] ,
         \u_a23_core/u_execute/u_register_bank/r7[21] ,
         \u_a23_core/u_execute/u_register_bank/r7[22] ,
         \u_a23_core/u_execute/u_register_bank/r7[23] ,
         \u_a23_core/u_execute/u_register_bank/r7[24] ,
         \u_a23_core/u_execute/u_register_bank/r7[25] ,
         \u_a23_core/u_execute/u_register_bank/r7[26] ,
         \u_a23_core/u_execute/u_register_bank/r7[27] ,
         \u_a23_core/u_execute/u_register_bank/r7[28] ,
         \u_a23_core/u_execute/u_register_bank/r7[29] ,
         \u_a23_core/u_execute/u_register_bank/r7[30] ,
         \u_a23_core/u_execute/u_register_bank/r7[31] ,
         \u_a23_core/u_execute/u_register_bank/r6[0] ,
         \u_a23_core/u_execute/u_register_bank/r6[1] ,
         \u_a23_core/u_execute/u_register_bank/r6[2] ,
         \u_a23_core/u_execute/u_register_bank/r6[3] ,
         \u_a23_core/u_execute/u_register_bank/r6[4] ,
         \u_a23_core/u_execute/u_register_bank/r6[5] ,
         \u_a23_core/u_execute/u_register_bank/r6[6] ,
         \u_a23_core/u_execute/u_register_bank/r6[7] ,
         \u_a23_core/u_execute/u_register_bank/r6[8] ,
         \u_a23_core/u_execute/u_register_bank/r6[9] ,
         \u_a23_core/u_execute/u_register_bank/r6[10] ,
         \u_a23_core/u_execute/u_register_bank/r6[11] ,
         \u_a23_core/u_execute/u_register_bank/r6[12] ,
         \u_a23_core/u_execute/u_register_bank/r6[13] ,
         \u_a23_core/u_execute/u_register_bank/r6[14] ,
         \u_a23_core/u_execute/u_register_bank/r6[15] ,
         \u_a23_core/u_execute/u_register_bank/r6[16] ,
         \u_a23_core/u_execute/u_register_bank/r6[17] ,
         \u_a23_core/u_execute/u_register_bank/r6[18] ,
         \u_a23_core/u_execute/u_register_bank/r6[19] ,
         \u_a23_core/u_execute/u_register_bank/r6[20] ,
         \u_a23_core/u_execute/u_register_bank/r6[21] ,
         \u_a23_core/u_execute/u_register_bank/r6[22] ,
         \u_a23_core/u_execute/u_register_bank/r6[23] ,
         \u_a23_core/u_execute/u_register_bank/r6[24] ,
         \u_a23_core/u_execute/u_register_bank/r6[25] ,
         \u_a23_core/u_execute/u_register_bank/r6[26] ,
         \u_a23_core/u_execute/u_register_bank/r6[27] ,
         \u_a23_core/u_execute/u_register_bank/r6[28] ,
         \u_a23_core/u_execute/u_register_bank/r6[29] ,
         \u_a23_core/u_execute/u_register_bank/r6[30] ,
         \u_a23_core/u_execute/u_register_bank/r6[31] ,
         \u_a23_core/u_execute/u_register_bank/r5[0] ,
         \u_a23_core/u_execute/u_register_bank/r5[1] ,
         \u_a23_core/u_execute/u_register_bank/r5[2] ,
         \u_a23_core/u_execute/u_register_bank/r5[3] ,
         \u_a23_core/u_execute/u_register_bank/r5[4] ,
         \u_a23_core/u_execute/u_register_bank/r5[5] ,
         \u_a23_core/u_execute/u_register_bank/r5[6] ,
         \u_a23_core/u_execute/u_register_bank/r5[7] ,
         \u_a23_core/u_execute/u_register_bank/r5[8] ,
         \u_a23_core/u_execute/u_register_bank/r5[9] ,
         \u_a23_core/u_execute/u_register_bank/r5[10] ,
         \u_a23_core/u_execute/u_register_bank/r5[11] ,
         \u_a23_core/u_execute/u_register_bank/r5[12] ,
         \u_a23_core/u_execute/u_register_bank/r5[13] ,
         \u_a23_core/u_execute/u_register_bank/r5[14] ,
         \u_a23_core/u_execute/u_register_bank/r5[15] ,
         \u_a23_core/u_execute/u_register_bank/r5[16] ,
         \u_a23_core/u_execute/u_register_bank/r5[17] ,
         \u_a23_core/u_execute/u_register_bank/r5[18] ,
         \u_a23_core/u_execute/u_register_bank/r5[19] ,
         \u_a23_core/u_execute/u_register_bank/r5[20] ,
         \u_a23_core/u_execute/u_register_bank/r5[21] ,
         \u_a23_core/u_execute/u_register_bank/r5[22] ,
         \u_a23_core/u_execute/u_register_bank/r5[23] ,
         \u_a23_core/u_execute/u_register_bank/r5[24] ,
         \u_a23_core/u_execute/u_register_bank/r5[25] ,
         \u_a23_core/u_execute/u_register_bank/r5[26] ,
         \u_a23_core/u_execute/u_register_bank/r5[27] ,
         \u_a23_core/u_execute/u_register_bank/r5[28] ,
         \u_a23_core/u_execute/u_register_bank/r5[29] ,
         \u_a23_core/u_execute/u_register_bank/r5[30] ,
         \u_a23_core/u_execute/u_register_bank/r5[31] ,
         \u_a23_core/u_execute/u_register_bank/r4[0] ,
         \u_a23_core/u_execute/u_register_bank/r4[1] ,
         \u_a23_core/u_execute/u_register_bank/r4[2] ,
         \u_a23_core/u_execute/u_register_bank/r4[3] ,
         \u_a23_core/u_execute/u_register_bank/r4[4] ,
         \u_a23_core/u_execute/u_register_bank/r4[5] ,
         \u_a23_core/u_execute/u_register_bank/r4[6] ,
         \u_a23_core/u_execute/u_register_bank/r4[7] ,
         \u_a23_core/u_execute/u_register_bank/r4[8] ,
         \u_a23_core/u_execute/u_register_bank/r4[9] ,
         \u_a23_core/u_execute/u_register_bank/r4[10] ,
         \u_a23_core/u_execute/u_register_bank/r4[11] ,
         \u_a23_core/u_execute/u_register_bank/r4[12] ,
         \u_a23_core/u_execute/u_register_bank/r4[13] ,
         \u_a23_core/u_execute/u_register_bank/r4[14] ,
         \u_a23_core/u_execute/u_register_bank/r4[15] ,
         \u_a23_core/u_execute/u_register_bank/r4[16] ,
         \u_a23_core/u_execute/u_register_bank/r4[17] ,
         \u_a23_core/u_execute/u_register_bank/r4[18] ,
         \u_a23_core/u_execute/u_register_bank/r4[19] ,
         \u_a23_core/u_execute/u_register_bank/r4[20] ,
         \u_a23_core/u_execute/u_register_bank/r4[21] ,
         \u_a23_core/u_execute/u_register_bank/r4[22] ,
         \u_a23_core/u_execute/u_register_bank/r4[23] ,
         \u_a23_core/u_execute/u_register_bank/r4[24] ,
         \u_a23_core/u_execute/u_register_bank/r4[25] ,
         \u_a23_core/u_execute/u_register_bank/r4[26] ,
         \u_a23_core/u_execute/u_register_bank/r4[27] ,
         \u_a23_core/u_execute/u_register_bank/r4[28] ,
         \u_a23_core/u_execute/u_register_bank/r4[29] ,
         \u_a23_core/u_execute/u_register_bank/r4[30] ,
         \u_a23_core/u_execute/u_register_bank/r4[31] ,
         \u_a23_core/u_execute/u_register_bank/r3[0] ,
         \u_a23_core/u_execute/u_register_bank/r3[1] ,
         \u_a23_core/u_execute/u_register_bank/r3[2] ,
         \u_a23_core/u_execute/u_register_bank/r3[3] ,
         \u_a23_core/u_execute/u_register_bank/r3[4] ,
         \u_a23_core/u_execute/u_register_bank/r3[5] ,
         \u_a23_core/u_execute/u_register_bank/r3[6] ,
         \u_a23_core/u_execute/u_register_bank/r3[7] ,
         \u_a23_core/u_execute/u_register_bank/r3[8] ,
         \u_a23_core/u_execute/u_register_bank/r3[9] ,
         \u_a23_core/u_execute/u_register_bank/r3[10] ,
         \u_a23_core/u_execute/u_register_bank/r3[11] ,
         \u_a23_core/u_execute/u_register_bank/r3[12] ,
         \u_a23_core/u_execute/u_register_bank/r3[13] ,
         \u_a23_core/u_execute/u_register_bank/r3[14] ,
         \u_a23_core/u_execute/u_register_bank/r3[15] ,
         \u_a23_core/u_execute/u_register_bank/r3[16] ,
         \u_a23_core/u_execute/u_register_bank/r3[17] ,
         \u_a23_core/u_execute/u_register_bank/r3[18] ,
         \u_a23_core/u_execute/u_register_bank/r3[19] ,
         \u_a23_core/u_execute/u_register_bank/r3[20] ,
         \u_a23_core/u_execute/u_register_bank/r3[21] ,
         \u_a23_core/u_execute/u_register_bank/r3[22] ,
         \u_a23_core/u_execute/u_register_bank/r3[23] ,
         \u_a23_core/u_execute/u_register_bank/r3[24] ,
         \u_a23_core/u_execute/u_register_bank/r3[25] ,
         \u_a23_core/u_execute/u_register_bank/r3[26] ,
         \u_a23_core/u_execute/u_register_bank/r3[27] ,
         \u_a23_core/u_execute/u_register_bank/r3[28] ,
         \u_a23_core/u_execute/u_register_bank/r3[29] ,
         \u_a23_core/u_execute/u_register_bank/r3[30] ,
         \u_a23_core/u_execute/u_register_bank/r3[31] ,
         \u_a23_core/u_execute/u_register_bank/r2[0] ,
         \u_a23_core/u_execute/u_register_bank/r2[1] ,
         \u_a23_core/u_execute/u_register_bank/r2[2] ,
         \u_a23_core/u_execute/u_register_bank/r2[3] ,
         \u_a23_core/u_execute/u_register_bank/r2[4] ,
         \u_a23_core/u_execute/u_register_bank/r2[5] ,
         \u_a23_core/u_execute/u_register_bank/r2[6] ,
         \u_a23_core/u_execute/u_register_bank/r2[7] ,
         \u_a23_core/u_execute/u_register_bank/r2[8] ,
         \u_a23_core/u_execute/u_register_bank/r2[9] ,
         \u_a23_core/u_execute/u_register_bank/r2[10] ,
         \u_a23_core/u_execute/u_register_bank/r2[11] ,
         \u_a23_core/u_execute/u_register_bank/r2[12] ,
         \u_a23_core/u_execute/u_register_bank/r2[13] ,
         \u_a23_core/u_execute/u_register_bank/r2[14] ,
         \u_a23_core/u_execute/u_register_bank/r2[15] ,
         \u_a23_core/u_execute/u_register_bank/r2[16] ,
         \u_a23_core/u_execute/u_register_bank/r2[17] ,
         \u_a23_core/u_execute/u_register_bank/r2[18] ,
         \u_a23_core/u_execute/u_register_bank/r2[19] ,
         \u_a23_core/u_execute/u_register_bank/r2[20] ,
         \u_a23_core/u_execute/u_register_bank/r2[21] ,
         \u_a23_core/u_execute/u_register_bank/r2[22] ,
         \u_a23_core/u_execute/u_register_bank/r2[23] ,
         \u_a23_core/u_execute/u_register_bank/r2[24] ,
         \u_a23_core/u_execute/u_register_bank/r2[25] ,
         \u_a23_core/u_execute/u_register_bank/r2[26] ,
         \u_a23_core/u_execute/u_register_bank/r2[27] ,
         \u_a23_core/u_execute/u_register_bank/r2[28] ,
         \u_a23_core/u_execute/u_register_bank/r2[29] ,
         \u_a23_core/u_execute/u_register_bank/r2[30] ,
         \u_a23_core/u_execute/u_register_bank/r2[31] ,
         \u_a23_core/u_execute/u_register_bank/r1[0] ,
         \u_a23_core/u_execute/u_register_bank/r1[1] ,
         \u_a23_core/u_execute/u_register_bank/r1[2] ,
         \u_a23_core/u_execute/u_register_bank/r1[3] ,
         \u_a23_core/u_execute/u_register_bank/r1[4] ,
         \u_a23_core/u_execute/u_register_bank/r1[5] ,
         \u_a23_core/u_execute/u_register_bank/r1[6] ,
         \u_a23_core/u_execute/u_register_bank/r1[7] ,
         \u_a23_core/u_execute/u_register_bank/r1[8] ,
         \u_a23_core/u_execute/u_register_bank/r1[9] ,
         \u_a23_core/u_execute/u_register_bank/r1[10] ,
         \u_a23_core/u_execute/u_register_bank/r1[11] ,
         \u_a23_core/u_execute/u_register_bank/r1[12] ,
         \u_a23_core/u_execute/u_register_bank/r1[13] ,
         \u_a23_core/u_execute/u_register_bank/r1[14] ,
         \u_a23_core/u_execute/u_register_bank/r1[15] ,
         \u_a23_core/u_execute/u_register_bank/r1[16] ,
         \u_a23_core/u_execute/u_register_bank/r1[17] ,
         \u_a23_core/u_execute/u_register_bank/r1[18] ,
         \u_a23_core/u_execute/u_register_bank/r1[19] ,
         \u_a23_core/u_execute/u_register_bank/r1[20] ,
         \u_a23_core/u_execute/u_register_bank/r1[21] ,
         \u_a23_core/u_execute/u_register_bank/r1[22] ,
         \u_a23_core/u_execute/u_register_bank/r1[23] ,
         \u_a23_core/u_execute/u_register_bank/r1[24] ,
         \u_a23_core/u_execute/u_register_bank/r1[25] ,
         \u_a23_core/u_execute/u_register_bank/r1[26] ,
         \u_a23_core/u_execute/u_register_bank/r1[27] ,
         \u_a23_core/u_execute/u_register_bank/r1[28] ,
         \u_a23_core/u_execute/u_register_bank/r1[29] ,
         \u_a23_core/u_execute/u_register_bank/r1[30] ,
         \u_a23_core/u_execute/u_register_bank/r1[31] ,
         \u_a23_core/u_execute/u_register_bank/r0[0] ,
         \u_a23_core/u_execute/u_register_bank/r0[1] ,
         \u_a23_core/u_execute/u_register_bank/r0[2] ,
         \u_a23_core/u_execute/u_register_bank/r0[3] ,
         \u_a23_core/u_execute/u_register_bank/r0[4] ,
         \u_a23_core/u_execute/u_register_bank/r0[5] ,
         \u_a23_core/u_execute/u_register_bank/r0[6] ,
         \u_a23_core/u_execute/u_register_bank/r0[7] ,
         \u_a23_core/u_execute/u_register_bank/r0[8] ,
         \u_a23_core/u_execute/u_register_bank/r0[9] ,
         \u_a23_core/u_execute/u_register_bank/r0[10] ,
         \u_a23_core/u_execute/u_register_bank/r0[11] ,
         \u_a23_core/u_execute/u_register_bank/r0[12] ,
         \u_a23_core/u_execute/u_register_bank/r0[13] ,
         \u_a23_core/u_execute/u_register_bank/r0[14] ,
         \u_a23_core/u_execute/u_register_bank/r0[15] ,
         \u_a23_core/u_execute/u_register_bank/r0[16] ,
         \u_a23_core/u_execute/u_register_bank/r0[17] ,
         \u_a23_core/u_execute/u_register_bank/r0[18] ,
         \u_a23_core/u_execute/u_register_bank/r0[19] ,
         \u_a23_core/u_execute/u_register_bank/r0[20] ,
         \u_a23_core/u_execute/u_register_bank/r0[21] ,
         \u_a23_core/u_execute/u_register_bank/r0[22] ,
         \u_a23_core/u_execute/u_register_bank/r0[23] ,
         \u_a23_core/u_execute/u_register_bank/r0[24] ,
         \u_a23_core/u_execute/u_register_bank/r0[25] ,
         \u_a23_core/u_execute/u_register_bank/r0[26] ,
         \u_a23_core/u_execute/u_register_bank/r0[27] ,
         \u_a23_core/u_execute/u_register_bank/r0[28] ,
         \u_a23_core/u_execute/u_register_bank/r0[29] ,
         \u_a23_core/u_execute/u_register_bank/r0[30] ,
         \u_a23_core/u_execute/u_register_bank/r0[31] ,
         \u_a23_core/u_execute/u_multiply/add_90/carry[32] ,
         \u_a23_core/u_execute/u_multiply/add_90/carry[31] ,
         \u_a23_core/u_execute/u_multiply/add_90/carry[30] ,
         \u_a23_core/u_execute/u_multiply/add_90/carry[29] ,
         \u_a23_core/u_execute/u_multiply/add_90/carry[28] ,
         \u_a23_core/u_execute/u_multiply/add_90/carry[27] ,
         \u_a23_core/u_execute/u_multiply/add_90/carry[26] ,
         \u_a23_core/u_execute/u_multiply/add_90/carry[25] ,
         \u_a23_core/u_execute/u_multiply/add_90/carry[24] ,
         \u_a23_core/u_execute/u_multiply/add_90/carry[23] ,
         \u_a23_core/u_execute/u_multiply/add_90/carry[22] ,
         \u_a23_core/u_execute/u_multiply/add_90/carry[21] ,
         \u_a23_core/u_execute/u_multiply/add_90/carry[20] ,
         \u_a23_core/u_execute/u_multiply/add_90/carry[19] ,
         \u_a23_core/u_execute/u_multiply/add_90/carry[18] ,
         \u_a23_core/u_execute/u_multiply/add_90/carry[17] ,
         \u_a23_core/u_execute/u_multiply/add_90/carry[16] ,
         \u_a23_core/u_execute/u_multiply/add_90/carry[15] ,
         \u_a23_core/u_execute/u_multiply/add_90/carry[14] ,
         \u_a23_core/u_execute/u_multiply/add_90/carry[13] ,
         \u_a23_core/u_execute/u_multiply/add_90/carry[12] ,
         \u_a23_core/u_execute/u_multiply/add_90/carry[11] ,
         \u_a23_core/u_execute/u_multiply/add_90/carry[10] ,
         \u_a23_core/u_execute/u_multiply/add_90/carry[9] ,
         \u_a23_core/u_execute/u_multiply/add_90/carry[8] ,
         \u_a23_core/u_execute/u_multiply/add_90/carry[7] ,
         \u_a23_core/u_execute/u_multiply/add_90/carry[6] ,
         \u_a23_core/u_execute/u_multiply/add_90/carry[5] ,
         \u_a23_core/u_execute/u_multiply/add_90/carry[4] ,
         \u_a23_core/u_execute/u_multiply/add_90/carry[3] ,
         \u_a23_core/u_execute/u_multiply/add_90/carry[2] ,
         \u_a23_core/u_execute/u_multiply/add_100/carry[33] ,
         \u_a23_core/u_execute/u_multiply/add_100/carry[32] ,
         \u_a23_core/u_execute/u_multiply/add_100/carry[31] ,
         \u_a23_core/u_execute/u_multiply/add_100/carry[30] ,
         \u_a23_core/u_execute/u_multiply/add_100/carry[29] ,
         \u_a23_core/u_execute/u_multiply/add_100/carry[28] ,
         \u_a23_core/u_execute/u_multiply/add_100/carry[27] ,
         \u_a23_core/u_execute/u_multiply/add_100/carry[26] ,
         \u_a23_core/u_execute/u_multiply/add_100/carry[25] ,
         \u_a23_core/u_execute/u_multiply/add_100/carry[24] ,
         \u_a23_core/u_execute/u_multiply/add_100/carry[23] ,
         \u_a23_core/u_execute/u_multiply/add_100/carry[22] ,
         \u_a23_core/u_execute/u_multiply/add_100/carry[21] ,
         \u_a23_core/u_execute/u_multiply/add_100/carry[20] ,
         \u_a23_core/u_execute/u_multiply/add_100/carry[19] ,
         \u_a23_core/u_execute/u_multiply/add_100/carry[18] ,
         \u_a23_core/u_execute/u_multiply/add_100/carry[17] ,
         \u_a23_core/u_execute/u_multiply/add_100/carry[16] ,
         \u_a23_core/u_execute/u_multiply/add_100/carry[15] ,
         \u_a23_core/u_execute/u_multiply/add_100/carry[14] ,
         \u_a23_core/u_execute/u_multiply/add_100/carry[13] ,
         \u_a23_core/u_execute/u_multiply/add_100/carry[12] ,
         \u_a23_core/u_execute/u_multiply/add_100/carry[11] ,
         \u_a23_core/u_execute/u_multiply/add_100/carry[10] ,
         \u_a23_core/u_execute/u_multiply/add_100/carry[9] ,
         \u_a23_core/u_execute/u_multiply/add_100/carry[8] ,
         \u_a23_core/u_execute/u_multiply/add_100/carry[7] ,
         \u_a23_core/u_execute/u_multiply/add_100/carry[6] ,
         \u_a23_core/u_execute/u_multiply/add_100/carry[5] ,
         \u_a23_core/u_execute/u_multiply/add_100/carry[4] ,
         \u_a23_core/u_execute/u_multiply/add_100/carry[3] ,
         \u_a23_core/u_execute/u_multiply/add_100/carry[2] ,
         \u_a23_core/u_execute/u_multiply/add_100/carry[1] ,
         \u_a23_core/u_execute/u_multiply/add_105/carry[31] ,
         \u_a23_core/u_execute/u_multiply/add_105/carry[30] ,
         \u_a23_core/u_execute/u_multiply/add_105/carry[29] ,
         \u_a23_core/u_execute/u_multiply/add_105/carry[28] ,
         \u_a23_core/u_execute/u_multiply/add_105/carry[27] ,
         \u_a23_core/u_execute/u_multiply/add_105/carry[26] ,
         \u_a23_core/u_execute/u_multiply/add_105/carry[25] ,
         \u_a23_core/u_execute/u_multiply/add_105/carry[24] ,
         \u_a23_core/u_execute/u_multiply/add_105/carry[23] ,
         \u_a23_core/u_execute/u_multiply/add_105/carry[22] ,
         \u_a23_core/u_execute/u_multiply/add_105/carry[21] ,
         \u_a23_core/u_execute/u_multiply/add_105/carry[20] ,
         \u_a23_core/u_execute/u_multiply/add_105/carry[19] ,
         \u_a23_core/u_execute/u_multiply/add_105/carry[18] ,
         \u_a23_core/u_execute/u_multiply/add_105/carry[17] ,
         \u_a23_core/u_execute/u_multiply/add_105/carry[16] ,
         \u_a23_core/u_execute/u_multiply/add_105/carry[15] ,
         \u_a23_core/u_execute/u_multiply/add_105/carry[14] ,
         \u_a23_core/u_execute/u_multiply/add_105/carry[13] ,
         \u_a23_core/u_execute/u_multiply/add_105/carry[12] ,
         \u_a23_core/u_execute/u_multiply/add_105/carry[11] ,
         \u_a23_core/u_execute/u_multiply/add_105/carry[10] ,
         \u_a23_core/u_execute/u_multiply/add_105/carry[9] ,
         \u_a23_core/u_execute/u_multiply/add_105/carry[8] ,
         \u_a23_core/u_execute/u_multiply/add_105/carry[7] ,
         \u_a23_core/u_execute/u_multiply/add_105/carry[6] ,
         \u_a23_core/u_execute/u_multiply/add_105/carry[5] ,
         \u_a23_core/u_execute/u_multiply/add_105/carry[4] ,
         \u_a23_core/u_execute/u_multiply/add_105/carry[3] ,
         \u_a23_core/u_execute/u_multiply/add_105/carry[2] ,
         \u_a23_core/u_execute/u_multiply/add_105/carry[1] ,
         \u_a23_core/u_execute/u_multiply/add_139/carry[5] ,
         \u_a23_core/u_execute/u_multiply/add_139/carry[4] ,
         \u_a23_core/u_execute/u_multiply/add_139/carry[3] ,
         \u_a23_core/u_execute/u_multiply/add_139/carry[2] ,
         \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[31] ,
         \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[30] ,
         \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[29] ,
         \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[28] ,
         \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[27] ,
         \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[26] ,
         \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[25] ,
         \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[24] ,
         \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[23] ,
         \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[22] ,
         \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[21] ,
         \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[20] ,
         \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[19] ,
         \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[18] ,
         \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[17] ,
         \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[16] ,
         \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[15] ,
         \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[14] ,
         \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[13] ,
         \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[12] ,
         \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[11] ,
         \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[10] ,
         \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[9] ,
         \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[8] ,
         \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[7] ,
         \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[6] ,
         \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[5] ,
         \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[4] ,
         \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[3] ,
         \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[2] ,
         \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[1] ,
         \u_a23_core/u_execute/add_165/carry[25] ,
         \u_a23_core/u_execute/add_165/carry[24] ,
         \u_a23_core/u_execute/add_165/carry[23] ,
         \u_a23_core/u_execute/add_165/carry[22] ,
         \u_a23_core/u_execute/add_165/carry[21] ,
         \u_a23_core/u_execute/add_165/carry[20] ,
         \u_a23_core/u_execute/add_165/carry[19] ,
         \u_a23_core/u_execute/add_165/carry[18] ,
         \u_a23_core/u_execute/add_165/carry[17] ,
         \u_a23_core/u_execute/add_165/carry[16] ,
         \u_a23_core/u_execute/add_165/carry[15] ,
         \u_a23_core/u_execute/add_165/carry[14] ,
         \u_a23_core/u_execute/add_165/carry[13] ,
         \u_a23_core/u_execute/add_165/carry[12] ,
         \u_a23_core/u_execute/add_165/carry[11] ,
         \u_a23_core/u_execute/add_165/carry[10] ,
         \u_a23_core/u_execute/add_165/carry[9] ,
         \u_a23_core/u_execute/add_165/carry[8] ,
         \u_a23_core/u_execute/add_165/carry[7] ,
         \u_a23_core/u_execute/add_165/carry[6] ,
         \u_a23_core/u_execute/add_165/carry[5] ,
         \u_a23_core/u_execute/add_165/carry[4] ,
         \u_a23_core/u_execute/sub_166/carry[26] ,
         \u_a23_core/u_execute/sub_166/carry[25] ,
         \u_a23_core/u_execute/sub_166/carry[24] ,
         \u_a23_core/u_execute/sub_166/carry[23] ,
         \u_a23_core/u_execute/sub_166/carry[22] ,
         \u_a23_core/u_execute/sub_166/carry[21] ,
         \u_a23_core/u_execute/sub_166/carry[20] ,
         \u_a23_core/u_execute/sub_166/carry[19] ,
         \u_a23_core/u_execute/sub_166/carry[18] ,
         \u_a23_core/u_execute/sub_166/carry[17] ,
         \u_a23_core/u_execute/sub_166/carry[16] ,
         \u_a23_core/u_execute/sub_166/carry[15] ,
         \u_a23_core/u_execute/sub_166/carry[14] ,
         \u_a23_core/u_execute/sub_166/carry[13] ,
         \u_a23_core/u_execute/sub_166/carry[12] ,
         \u_a23_core/u_execute/sub_166/carry[11] ,
         \u_a23_core/u_execute/sub_166/carry[10] ,
         \u_a23_core/u_execute/sub_166/carry[9] ,
         \u_a23_core/u_execute/sub_166/carry[8] ,
         \u_a23_core/u_execute/sub_166/carry[7] ,
         \u_a23_core/u_execute/sub_166/carry[6] ,
         \u_a23_core/u_execute/sub_166/carry[5] ,
         \u_a23_core/u_execute/sub_166/carry[4] ,
         \u_a23_core/u_execute/add_167/carry[31] ,
         \u_a23_core/u_execute/add_167/carry[30] ,
         \u_a23_core/u_execute/add_167/carry[29] ,
         \u_a23_core/u_execute/add_167/carry[28] ,
         \u_a23_core/u_execute/add_167/carry[27] ,
         \u_a23_core/u_execute/add_167/carry[26] ,
         \u_a23_core/u_execute/add_167/carry[25] ,
         \u_a23_core/u_execute/add_167/carry[24] ,
         \u_a23_core/u_execute/add_167/carry[23] ,
         \u_a23_core/u_execute/add_167/carry[22] ,
         \u_a23_core/u_execute/add_167/carry[21] ,
         \u_a23_core/u_execute/add_167/carry[20] ,
         \u_a23_core/u_execute/add_167/carry[19] ,
         \u_a23_core/u_execute/add_167/carry[18] ,
         \u_a23_core/u_execute/add_167/carry[17] ,
         \u_a23_core/u_execute/add_167/carry[16] ,
         \u_a23_core/u_execute/add_167/carry[15] ,
         \u_a23_core/u_execute/add_167/carry[14] ,
         \u_a23_core/u_execute/add_167/carry[13] ,
         \u_a23_core/u_execute/add_167/carry[12] ,
         \u_a23_core/u_execute/add_167/carry[11] ,
         \u_a23_core/u_execute/add_167/carry[10] ,
         \u_a23_core/u_execute/add_167/carry[9] ,
         \u_a23_core/u_execute/add_167/carry[8] ,
         \u_a23_core/u_execute/add_167/carry[7] ,
         \u_a23_core/u_execute/add_167/carry[6] ,
         \u_a23_core/u_execute/add_167/carry[5] ,
         \u_a23_core/u_execute/add_167/carry[4] ,
         \u_a23_core/u_execute/add_168/carry[31] ,
         \u_a23_core/u_execute/add_168/carry[30] ,
         \u_a23_core/u_execute/add_168/carry[29] ,
         \u_a23_core/u_execute/add_168/carry[28] ,
         \u_a23_core/u_execute/add_168/carry[27] ,
         \u_a23_core/u_execute/add_168/carry[26] ,
         \u_a23_core/u_execute/add_168/carry[25] ,
         \u_a23_core/u_execute/add_168/carry[24] ,
         \u_a23_core/u_execute/add_168/carry[23] ,
         \u_a23_core/u_execute/add_168/carry[22] ,
         \u_a23_core/u_execute/add_168/carry[21] ,
         \u_a23_core/u_execute/add_168/carry[20] ,
         \u_a23_core/u_execute/add_168/carry[19] ,
         \u_a23_core/u_execute/add_168/carry[18] ,
         \u_a23_core/u_execute/add_168/carry[17] ,
         \u_a23_core/u_execute/add_168/carry[16] ,
         \u_a23_core/u_execute/add_168/carry[15] ,
         \u_a23_core/u_execute/add_168/carry[14] ,
         \u_a23_core/u_execute/add_168/carry[13] ,
         \u_a23_core/u_execute/add_168/carry[12] ,
         \u_a23_core/u_execute/add_168/carry[11] ,
         \u_a23_core/u_execute/add_168/carry[10] ,
         \u_a23_core/u_execute/add_168/carry[9] ,
         \u_a23_core/u_execute/add_168/carry[8] ,
         \u_a23_core/u_execute/add_168/carry[7] ,
         \u_a23_core/u_execute/add_168/carry[6] ,
         \u_a23_core/u_execute/add_168/carry[5] ,
         \u_a23_core/u_execute/add_168/carry[4] ,
         \u_a23_core/u_execute/add_169/carry[31] ,
         \u_a23_core/u_execute/add_169/carry[30] ,
         \u_a23_core/u_execute/add_169/carry[29] ,
         \u_a23_core/u_execute/add_169/carry[28] ,
         \u_a23_core/u_execute/add_169/carry[27] ,
         \u_a23_core/u_execute/add_169/carry[26] ,
         \u_a23_core/u_execute/add_169/carry[25] ,
         \u_a23_core/u_execute/add_169/carry[24] ,
         \u_a23_core/u_execute/add_169/carry[23] ,
         \u_a23_core/u_execute/add_169/carry[22] ,
         \u_a23_core/u_execute/add_169/carry[21] ,
         \u_a23_core/u_execute/add_169/carry[20] ,
         \u_a23_core/u_execute/add_169/carry[19] ,
         \u_a23_core/u_execute/add_169/carry[18] ,
         \u_a23_core/u_execute/add_169/carry[17] ,
         \u_a23_core/u_execute/add_169/carry[16] ,
         \u_a23_core/u_execute/add_169/carry[15] ,
         \u_a23_core/u_execute/add_169/carry[14] ,
         \u_a23_core/u_execute/add_169/carry[13] ,
         \u_a23_core/u_execute/add_169/carry[12] ,
         \u_a23_core/u_execute/add_169/carry[11] ,
         \u_a23_core/u_execute/add_169/carry[10] ,
         \u_a23_core/u_execute/add_169/carry[9] ,
         \u_a23_core/u_execute/add_169/carry[8] ,
         \u_a23_core/u_execute/add_169/carry[7] ,
         \u_a23_core/u_execute/add_169/carry[6] ,
         \u_a23_core/u_execute/add_169/carry[5] ,
         \u_a23_core/u_execute/add_169/carry[4] ,
         \u_a23_core/u_decode/add_9_root_add_415_15/carry[1] ,
         \u_a23_core/u_decode/add_8_root_add_415_15/carry[1] ,
         \u_a23_core/u_decode/add_7_root_add_415_15/carry[2] ,
         \u_a23_core/u_decode/add_7_root_add_415_15/carry[1] ,
         \u_a23_core/u_decode/add_6_root_add_415_15/carry[3] ,
         \u_a23_core/u_decode/add_6_root_add_415_15/carry[2] ,
         \u_a23_core/u_decode/add_6_root_add_415_15/carry[1] , n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
         n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
         n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
         n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
         n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
         n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
         n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
         n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547,
         n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555,
         n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563,
         n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
         n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579,
         n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
         n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595,
         n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603,
         n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611,
         n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619,
         n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627,
         n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635,
         n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
         n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651,
         n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659,
         n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667,
         n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675,
         n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683,
         n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691,
         n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699,
         n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707,
         n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715,
         n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723,
         n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731,
         n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739,
         n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747,
         n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755,
         n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763,
         n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771,
         n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779,
         n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787,
         n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795,
         n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803,
         n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811,
         n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819,
         n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827,
         n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835,
         n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843,
         n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851,
         n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859,
         n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867,
         n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
         n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883,
         n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891,
         n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899,
         n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907,
         n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915,
         n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923,
         n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931,
         n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939,
         n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
         n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955,
         n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963,
         n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971,
         n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
         n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987,
         n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995,
         n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003,
         n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011,
         n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019,
         n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027,
         n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035,
         n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043,
         n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051,
         n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059,
         n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067,
         n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075,
         n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083,
         n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
         n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099,
         n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107,
         n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115,
         n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123,
         n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131,
         n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139,
         n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147,
         n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155,
         n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163,
         n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171,
         n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179,
         n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187,
         n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195,
         n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203,
         n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211,
         n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219,
         n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227,
         n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235,
         n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243,
         n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251,
         n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259,
         n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267,
         n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275,
         n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283,
         n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291,
         n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299,
         n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307,
         n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315,
         n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323,
         n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331,
         n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339,
         n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347,
         n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355,
         n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363,
         n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371,
         n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379,
         n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387,
         n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395,
         n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403,
         n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411,
         n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419,
         n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427,
         n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435,
         n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443,
         n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451,
         n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459,
         n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467,
         n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475,
         n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483,
         n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491,
         n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499,
         n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507,
         n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515,
         n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523,
         n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531,
         n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539,
         n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547,
         n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555,
         n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563,
         n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571,
         n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579,
         n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587,
         n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595,
         n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603,
         n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611,
         n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619,
         n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627,
         n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635,
         n16636, n16637;
  wire   [31:0] m_address;
  wire   [31:0] m_write;
  wire   [3:0] m_byte_enable;

  MUX \u_a23_mem/U23985  ( .IN0(\u_a23_mem/n23820 ), .IN1(\u_a23_mem/n23805 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/N1871 ) );
  MUX \u_a23_mem/U23984  ( .IN0(\u_a23_mem/n23819 ), .IN1(\u_a23_mem/n23812 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23820 ) );
  MUX \u_a23_mem/U23983  ( .IN0(\u_a23_mem/g_mem[0][7] ), .IN1(
        \u_a23_mem/g_mem[4][7] ), .SEL(m_address[2]), .F(\u_a23_mem/n23819 )
         );
  MUX \u_a23_mem/U23976  ( .IN0(\u_a23_mem/g_mem[8][7] ), .IN1(
        \u_a23_mem/g_mem[12][7] ), .SEL(m_address[2]), .F(\u_a23_mem/n23812 )
         );
  MUX \u_a23_mem/U23969  ( .IN0(\u_a23_mem/n23804 ), .IN1(\u_a23_mem/n23797 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23805 ) );
  MUX \u_a23_mem/U23968  ( .IN0(\u_a23_mem/g_mem[16][7] ), .IN1(
        \u_a23_mem/g_mem[20][7] ), .SEL(m_address[2]), .F(\u_a23_mem/n23804 )
         );
  MUX \u_a23_mem/U23961  ( .IN0(\u_a23_mem/g_mem[24][7] ), .IN1(
        \u_a23_mem/g_mem[28][7] ), .SEL(m_address[2]), .F(\u_a23_mem/n23797 )
         );
  MUX \u_a23_mem/U23954  ( .IN0(\u_a23_mem/n23790 ), .IN1(\u_a23_mem/n23775 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/N1872 ) );
  MUX \u_a23_mem/U23953  ( .IN0(\u_a23_mem/n23789 ), .IN1(\u_a23_mem/n23782 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23790 ) );
  MUX \u_a23_mem/U23952  ( .IN0(\u_a23_mem/g_mem[0][6] ), .IN1(
        \u_a23_mem/g_mem[4][6] ), .SEL(m_address[2]), .F(\u_a23_mem/n23789 )
         );
  MUX \u_a23_mem/U23945  ( .IN0(\u_a23_mem/g_mem[8][6] ), .IN1(
        \u_a23_mem/g_mem[12][6] ), .SEL(m_address[2]), .F(\u_a23_mem/n23782 )
         );
  MUX \u_a23_mem/U23938  ( .IN0(\u_a23_mem/n23774 ), .IN1(\u_a23_mem/n23767 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23775 ) );
  MUX \u_a23_mem/U23937  ( .IN0(\u_a23_mem/g_mem[16][6] ), .IN1(
        \u_a23_mem/g_mem[20][6] ), .SEL(m_address[2]), .F(\u_a23_mem/n23774 )
         );
  MUX \u_a23_mem/U23930  ( .IN0(\u_a23_mem/g_mem[24][6] ), .IN1(
        \u_a23_mem/g_mem[28][6] ), .SEL(m_address[2]), .F(\u_a23_mem/n23767 )
         );
  MUX \u_a23_mem/U23923  ( .IN0(\u_a23_mem/n23760 ), .IN1(\u_a23_mem/n23745 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/N1873 ) );
  MUX \u_a23_mem/U23922  ( .IN0(\u_a23_mem/n23759 ), .IN1(\u_a23_mem/n23752 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23760 ) );
  MUX \u_a23_mem/U23921  ( .IN0(\u_a23_mem/g_mem[0][5] ), .IN1(
        \u_a23_mem/g_mem[4][5] ), .SEL(m_address[2]), .F(\u_a23_mem/n23759 )
         );
  MUX \u_a23_mem/U23914  ( .IN0(\u_a23_mem/g_mem[8][5] ), .IN1(
        \u_a23_mem/g_mem[12][5] ), .SEL(m_address[2]), .F(\u_a23_mem/n23752 )
         );
  MUX \u_a23_mem/U23907  ( .IN0(\u_a23_mem/n23744 ), .IN1(\u_a23_mem/n23737 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23745 ) );
  MUX \u_a23_mem/U23906  ( .IN0(\u_a23_mem/g_mem[16][5] ), .IN1(
        \u_a23_mem/g_mem[20][5] ), .SEL(m_address[2]), .F(\u_a23_mem/n23744 )
         );
  MUX \u_a23_mem/U23899  ( .IN0(\u_a23_mem/g_mem[24][5] ), .IN1(
        \u_a23_mem/g_mem[28][5] ), .SEL(m_address[2]), .F(\u_a23_mem/n23737 )
         );
  MUX \u_a23_mem/U23892  ( .IN0(\u_a23_mem/n23730 ), .IN1(\u_a23_mem/n23715 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/N1874 ) );
  MUX \u_a23_mem/U23891  ( .IN0(\u_a23_mem/n23729 ), .IN1(\u_a23_mem/n23722 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23730 ) );
  MUX \u_a23_mem/U23890  ( .IN0(\u_a23_mem/g_mem[0][4] ), .IN1(
        \u_a23_mem/g_mem[4][4] ), .SEL(m_address[2]), .F(\u_a23_mem/n23729 )
         );
  MUX \u_a23_mem/U23883  ( .IN0(\u_a23_mem/g_mem[8][4] ), .IN1(
        \u_a23_mem/g_mem[12][4] ), .SEL(m_address[2]), .F(\u_a23_mem/n23722 )
         );
  MUX \u_a23_mem/U23876  ( .IN0(\u_a23_mem/n23714 ), .IN1(\u_a23_mem/n23707 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23715 ) );
  MUX \u_a23_mem/U23875  ( .IN0(\u_a23_mem/g_mem[16][4] ), .IN1(
        \u_a23_mem/g_mem[20][4] ), .SEL(m_address[2]), .F(\u_a23_mem/n23714 )
         );
  MUX \u_a23_mem/U23868  ( .IN0(\u_a23_mem/g_mem[24][4] ), .IN1(
        \u_a23_mem/g_mem[28][4] ), .SEL(m_address[2]), .F(\u_a23_mem/n23707 )
         );
  MUX \u_a23_mem/U23861  ( .IN0(\u_a23_mem/n23700 ), .IN1(\u_a23_mem/n23685 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/N1875 ) );
  MUX \u_a23_mem/U23860  ( .IN0(\u_a23_mem/n23699 ), .IN1(\u_a23_mem/n23692 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23700 ) );
  MUX \u_a23_mem/U23859  ( .IN0(\u_a23_mem/g_mem[0][3] ), .IN1(
        \u_a23_mem/g_mem[4][3] ), .SEL(m_address[2]), .F(\u_a23_mem/n23699 )
         );
  MUX \u_a23_mem/U23852  ( .IN0(\u_a23_mem/g_mem[8][3] ), .IN1(
        \u_a23_mem/g_mem[12][3] ), .SEL(m_address[2]), .F(\u_a23_mem/n23692 )
         );
  MUX \u_a23_mem/U23845  ( .IN0(\u_a23_mem/n23684 ), .IN1(\u_a23_mem/n23677 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23685 ) );
  MUX \u_a23_mem/U23844  ( .IN0(\u_a23_mem/g_mem[16][3] ), .IN1(
        \u_a23_mem/g_mem[20][3] ), .SEL(m_address[2]), .F(\u_a23_mem/n23684 )
         );
  MUX \u_a23_mem/U23837  ( .IN0(\u_a23_mem/g_mem[24][3] ), .IN1(
        \u_a23_mem/g_mem[28][3] ), .SEL(m_address[2]), .F(\u_a23_mem/n23677 )
         );
  MUX \u_a23_mem/U23830  ( .IN0(\u_a23_mem/n23670 ), .IN1(\u_a23_mem/n23655 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/N1876 ) );
  MUX \u_a23_mem/U23829  ( .IN0(\u_a23_mem/n23669 ), .IN1(\u_a23_mem/n23662 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23670 ) );
  MUX \u_a23_mem/U23828  ( .IN0(\u_a23_mem/g_mem[0][2] ), .IN1(
        \u_a23_mem/g_mem[4][2] ), .SEL(m_address[2]), .F(\u_a23_mem/n23669 )
         );
  MUX \u_a23_mem/U23821  ( .IN0(\u_a23_mem/g_mem[8][2] ), .IN1(
        \u_a23_mem/g_mem[12][2] ), .SEL(m_address[2]), .F(\u_a23_mem/n23662 )
         );
  MUX \u_a23_mem/U23814  ( .IN0(\u_a23_mem/n23654 ), .IN1(\u_a23_mem/n23647 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23655 ) );
  MUX \u_a23_mem/U23813  ( .IN0(\u_a23_mem/g_mem[16][2] ), .IN1(
        \u_a23_mem/g_mem[20][2] ), .SEL(m_address[2]), .F(\u_a23_mem/n23654 )
         );
  MUX \u_a23_mem/U23806  ( .IN0(\u_a23_mem/g_mem[24][2] ), .IN1(
        \u_a23_mem/g_mem[28][2] ), .SEL(m_address[2]), .F(\u_a23_mem/n23647 )
         );
  MUX \u_a23_mem/U23799  ( .IN0(\u_a23_mem/n23640 ), .IN1(\u_a23_mem/n23625 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/N1877 ) );
  MUX \u_a23_mem/U23798  ( .IN0(\u_a23_mem/n23639 ), .IN1(\u_a23_mem/n23632 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23640 ) );
  MUX \u_a23_mem/U23797  ( .IN0(\u_a23_mem/g_mem[0][1] ), .IN1(
        \u_a23_mem/g_mem[4][1] ), .SEL(m_address[2]), .F(\u_a23_mem/n23639 )
         );
  MUX \u_a23_mem/U23790  ( .IN0(\u_a23_mem/g_mem[8][1] ), .IN1(
        \u_a23_mem/g_mem[12][1] ), .SEL(m_address[2]), .F(\u_a23_mem/n23632 )
         );
  MUX \u_a23_mem/U23783  ( .IN0(\u_a23_mem/n23624 ), .IN1(\u_a23_mem/n23617 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23625 ) );
  MUX \u_a23_mem/U23782  ( .IN0(\u_a23_mem/g_mem[16][1] ), .IN1(
        \u_a23_mem/g_mem[20][1] ), .SEL(m_address[2]), .F(\u_a23_mem/n23624 )
         );
  MUX \u_a23_mem/U23775  ( .IN0(\u_a23_mem/g_mem[24][1] ), .IN1(
        \u_a23_mem/g_mem[28][1] ), .SEL(m_address[2]), .F(\u_a23_mem/n23617 )
         );
  MUX \u_a23_mem/U23768  ( .IN0(\u_a23_mem/n23610 ), .IN1(\u_a23_mem/n23595 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/N1878 ) );
  MUX \u_a23_mem/U23767  ( .IN0(\u_a23_mem/n23609 ), .IN1(\u_a23_mem/n23602 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23610 ) );
  MUX \u_a23_mem/U23766  ( .IN0(\u_a23_mem/g_mem[0][0] ), .IN1(
        \u_a23_mem/g_mem[4][0] ), .SEL(m_address[2]), .F(\u_a23_mem/n23609 )
         );
  MUX \u_a23_mem/U23759  ( .IN0(\u_a23_mem/g_mem[8][0] ), .IN1(
        \u_a23_mem/g_mem[12][0] ), .SEL(m_address[2]), .F(\u_a23_mem/n23602 )
         );
  MUX \u_a23_mem/U23752  ( .IN0(\u_a23_mem/n23594 ), .IN1(\u_a23_mem/n23587 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23595 ) );
  MUX \u_a23_mem/U23751  ( .IN0(\u_a23_mem/g_mem[16][0] ), .IN1(
        \u_a23_mem/g_mem[20][0] ), .SEL(m_address[2]), .F(\u_a23_mem/n23594 )
         );
  MUX \u_a23_mem/U23744  ( .IN0(\u_a23_mem/g_mem[24][0] ), .IN1(
        \u_a23_mem/g_mem[28][0] ), .SEL(m_address[2]), .F(\u_a23_mem/n23587 )
         );
  MUX \u_a23_mem/U23737  ( .IN0(\u_a23_mem/n23580 ), .IN1(\u_a23_mem/n23565 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/N1903 ) );
  MUX \u_a23_mem/U23736  ( .IN0(\u_a23_mem/n23579 ), .IN1(\u_a23_mem/n23572 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23580 ) );
  MUX \u_a23_mem/U23735  ( .IN0(\u_a23_mem/e_mem[0][7] ), .IN1(
        \u_a23_mem/e_mem[4][7] ), .SEL(m_address[2]), .F(\u_a23_mem/n23579 )
         );
  MUX \u_a23_mem/U23728  ( .IN0(\u_a23_mem/e_mem[8][7] ), .IN1(
        \u_a23_mem/e_mem[12][7] ), .SEL(m_address[2]), .F(\u_a23_mem/n23572 )
         );
  MUX \u_a23_mem/U23721  ( .IN0(\u_a23_mem/n23564 ), .IN1(\u_a23_mem/n23557 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23565 ) );
  MUX \u_a23_mem/U23720  ( .IN0(\u_a23_mem/e_mem[16][7] ), .IN1(
        \u_a23_mem/e_mem[20][7] ), .SEL(m_address[2]), .F(\u_a23_mem/n23564 )
         );
  MUX \u_a23_mem/U23713  ( .IN0(\u_a23_mem/e_mem[24][7] ), .IN1(
        \u_a23_mem/e_mem[28][7] ), .SEL(m_address[2]), .F(\u_a23_mem/n23557 )
         );
  MUX \u_a23_mem/U23706  ( .IN0(\u_a23_mem/n23550 ), .IN1(\u_a23_mem/n23535 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/N1904 ) );
  MUX \u_a23_mem/U23705  ( .IN0(\u_a23_mem/n23549 ), .IN1(\u_a23_mem/n23542 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23550 ) );
  MUX \u_a23_mem/U23704  ( .IN0(\u_a23_mem/e_mem[0][6] ), .IN1(
        \u_a23_mem/e_mem[4][6] ), .SEL(m_address[2]), .F(\u_a23_mem/n23549 )
         );
  MUX \u_a23_mem/U23697  ( .IN0(\u_a23_mem/e_mem[8][6] ), .IN1(
        \u_a23_mem/e_mem[12][6] ), .SEL(m_address[2]), .F(\u_a23_mem/n23542 )
         );
  MUX \u_a23_mem/U23690  ( .IN0(\u_a23_mem/n23534 ), .IN1(\u_a23_mem/n23527 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23535 ) );
  MUX \u_a23_mem/U23689  ( .IN0(\u_a23_mem/e_mem[16][6] ), .IN1(
        \u_a23_mem/e_mem[20][6] ), .SEL(m_address[2]), .F(\u_a23_mem/n23534 )
         );
  MUX \u_a23_mem/U23682  ( .IN0(\u_a23_mem/e_mem[24][6] ), .IN1(
        \u_a23_mem/e_mem[28][6] ), .SEL(m_address[2]), .F(\u_a23_mem/n23527 )
         );
  MUX \u_a23_mem/U23675  ( .IN0(\u_a23_mem/n23520 ), .IN1(\u_a23_mem/n23505 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/N1905 ) );
  MUX \u_a23_mem/U23674  ( .IN0(\u_a23_mem/n23519 ), .IN1(\u_a23_mem/n23512 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23520 ) );
  MUX \u_a23_mem/U23673  ( .IN0(\u_a23_mem/e_mem[0][5] ), .IN1(
        \u_a23_mem/e_mem[4][5] ), .SEL(m_address[2]), .F(\u_a23_mem/n23519 )
         );
  MUX \u_a23_mem/U23666  ( .IN0(\u_a23_mem/e_mem[8][5] ), .IN1(
        \u_a23_mem/e_mem[12][5] ), .SEL(m_address[2]), .F(\u_a23_mem/n23512 )
         );
  MUX \u_a23_mem/U23659  ( .IN0(\u_a23_mem/n23504 ), .IN1(\u_a23_mem/n23497 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23505 ) );
  MUX \u_a23_mem/U23658  ( .IN0(\u_a23_mem/e_mem[16][5] ), .IN1(
        \u_a23_mem/e_mem[20][5] ), .SEL(m_address[2]), .F(\u_a23_mem/n23504 )
         );
  MUX \u_a23_mem/U23651  ( .IN0(\u_a23_mem/e_mem[24][5] ), .IN1(
        \u_a23_mem/e_mem[28][5] ), .SEL(m_address[2]), .F(\u_a23_mem/n23497 )
         );
  MUX \u_a23_mem/U23644  ( .IN0(\u_a23_mem/n23490 ), .IN1(\u_a23_mem/n23475 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/N1906 ) );
  MUX \u_a23_mem/U23643  ( .IN0(\u_a23_mem/n23489 ), .IN1(\u_a23_mem/n23482 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23490 ) );
  MUX \u_a23_mem/U23642  ( .IN0(\u_a23_mem/e_mem[0][4] ), .IN1(
        \u_a23_mem/e_mem[4][4] ), .SEL(m_address[2]), .F(\u_a23_mem/n23489 )
         );
  MUX \u_a23_mem/U23635  ( .IN0(\u_a23_mem/e_mem[8][4] ), .IN1(
        \u_a23_mem/e_mem[12][4] ), .SEL(m_address[2]), .F(\u_a23_mem/n23482 )
         );
  MUX \u_a23_mem/U23628  ( .IN0(\u_a23_mem/n23474 ), .IN1(\u_a23_mem/n23467 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23475 ) );
  MUX \u_a23_mem/U23627  ( .IN0(\u_a23_mem/e_mem[16][4] ), .IN1(
        \u_a23_mem/e_mem[20][4] ), .SEL(m_address[2]), .F(\u_a23_mem/n23474 )
         );
  MUX \u_a23_mem/U23620  ( .IN0(\u_a23_mem/e_mem[24][4] ), .IN1(
        \u_a23_mem/e_mem[28][4] ), .SEL(m_address[2]), .F(\u_a23_mem/n23467 )
         );
  MUX \u_a23_mem/U23613  ( .IN0(\u_a23_mem/n23460 ), .IN1(\u_a23_mem/n23445 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/N1907 ) );
  MUX \u_a23_mem/U23612  ( .IN0(\u_a23_mem/n23459 ), .IN1(\u_a23_mem/n23452 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23460 ) );
  MUX \u_a23_mem/U23611  ( .IN0(\u_a23_mem/e_mem[0][3] ), .IN1(
        \u_a23_mem/e_mem[4][3] ), .SEL(m_address[2]), .F(\u_a23_mem/n23459 )
         );
  MUX \u_a23_mem/U23604  ( .IN0(\u_a23_mem/e_mem[8][3] ), .IN1(
        \u_a23_mem/e_mem[12][3] ), .SEL(m_address[2]), .F(\u_a23_mem/n23452 )
         );
  MUX \u_a23_mem/U23597  ( .IN0(\u_a23_mem/n23444 ), .IN1(\u_a23_mem/n23437 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23445 ) );
  MUX \u_a23_mem/U23596  ( .IN0(\u_a23_mem/e_mem[16][3] ), .IN1(
        \u_a23_mem/e_mem[20][3] ), .SEL(m_address[2]), .F(\u_a23_mem/n23444 )
         );
  MUX \u_a23_mem/U23589  ( .IN0(\u_a23_mem/e_mem[24][3] ), .IN1(
        \u_a23_mem/e_mem[28][3] ), .SEL(m_address[2]), .F(\u_a23_mem/n23437 )
         );
  MUX \u_a23_mem/U23582  ( .IN0(\u_a23_mem/n23430 ), .IN1(\u_a23_mem/n23415 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/N1908 ) );
  MUX \u_a23_mem/U23581  ( .IN0(\u_a23_mem/n23429 ), .IN1(\u_a23_mem/n23422 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23430 ) );
  MUX \u_a23_mem/U23580  ( .IN0(\u_a23_mem/e_mem[0][2] ), .IN1(
        \u_a23_mem/e_mem[4][2] ), .SEL(m_address[2]), .F(\u_a23_mem/n23429 )
         );
  MUX \u_a23_mem/U23573  ( .IN0(\u_a23_mem/e_mem[8][2] ), .IN1(
        \u_a23_mem/e_mem[12][2] ), .SEL(m_address[2]), .F(\u_a23_mem/n23422 )
         );
  MUX \u_a23_mem/U23566  ( .IN0(\u_a23_mem/n23414 ), .IN1(\u_a23_mem/n23407 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23415 ) );
  MUX \u_a23_mem/U23565  ( .IN0(\u_a23_mem/e_mem[16][2] ), .IN1(
        \u_a23_mem/e_mem[20][2] ), .SEL(m_address[2]), .F(\u_a23_mem/n23414 )
         );
  MUX \u_a23_mem/U23558  ( .IN0(\u_a23_mem/e_mem[24][2] ), .IN1(
        \u_a23_mem/e_mem[28][2] ), .SEL(m_address[2]), .F(\u_a23_mem/n23407 )
         );
  MUX \u_a23_mem/U23551  ( .IN0(\u_a23_mem/n23400 ), .IN1(\u_a23_mem/n23385 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/N1909 ) );
  MUX \u_a23_mem/U23550  ( .IN0(\u_a23_mem/n23399 ), .IN1(\u_a23_mem/n23392 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23400 ) );
  MUX \u_a23_mem/U23549  ( .IN0(\u_a23_mem/e_mem[0][1] ), .IN1(
        \u_a23_mem/e_mem[4][1] ), .SEL(m_address[2]), .F(\u_a23_mem/n23399 )
         );
  MUX \u_a23_mem/U23542  ( .IN0(\u_a23_mem/e_mem[8][1] ), .IN1(
        \u_a23_mem/e_mem[12][1] ), .SEL(m_address[2]), .F(\u_a23_mem/n23392 )
         );
  MUX \u_a23_mem/U23535  ( .IN0(\u_a23_mem/n23384 ), .IN1(\u_a23_mem/n23377 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23385 ) );
  MUX \u_a23_mem/U23534  ( .IN0(\u_a23_mem/e_mem[16][1] ), .IN1(
        \u_a23_mem/e_mem[20][1] ), .SEL(m_address[2]), .F(\u_a23_mem/n23384 )
         );
  MUX \u_a23_mem/U23527  ( .IN0(\u_a23_mem/e_mem[24][1] ), .IN1(
        \u_a23_mem/e_mem[28][1] ), .SEL(m_address[2]), .F(\u_a23_mem/n23377 )
         );
  MUX \u_a23_mem/U23520  ( .IN0(\u_a23_mem/n23370 ), .IN1(\u_a23_mem/n23355 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/N1910 ) );
  MUX \u_a23_mem/U23519  ( .IN0(\u_a23_mem/n23369 ), .IN1(\u_a23_mem/n23362 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23370 ) );
  MUX \u_a23_mem/U23518  ( .IN0(\u_a23_mem/e_mem[0][0] ), .IN1(
        \u_a23_mem/e_mem[4][0] ), .SEL(m_address[2]), .F(\u_a23_mem/n23369 )
         );
  MUX \u_a23_mem/U23511  ( .IN0(\u_a23_mem/e_mem[8][0] ), .IN1(
        \u_a23_mem/e_mem[12][0] ), .SEL(m_address[2]), .F(\u_a23_mem/n23362 )
         );
  MUX \u_a23_mem/U23504  ( .IN0(\u_a23_mem/n23354 ), .IN1(\u_a23_mem/n23347 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23355 ) );
  MUX \u_a23_mem/U23503  ( .IN0(\u_a23_mem/e_mem[16][0] ), .IN1(
        \u_a23_mem/e_mem[20][0] ), .SEL(m_address[2]), .F(\u_a23_mem/n23354 )
         );
  MUX \u_a23_mem/U23496  ( .IN0(\u_a23_mem/e_mem[24][0] ), .IN1(
        \u_a23_mem/e_mem[28][0] ), .SEL(m_address[2]), .F(\u_a23_mem/n23347 )
         );
  MUX \u_a23_mem/U23489  ( .IN0(\u_a23_mem/n23340 ), .IN1(\u_a23_mem/n23325 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/N1935 ) );
  MUX \u_a23_mem/U23488  ( .IN0(\u_a23_mem/n23339 ), .IN1(\u_a23_mem/n23332 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23340 ) );
  MUX \u_a23_mem/U23487  ( .IN0(o[7]), .IN1(o[39]), .SEL(m_address[2]), .F(
        \u_a23_mem/n23339 ) );
  MUX \u_a23_mem/U23480  ( .IN0(o[71]), .IN1(o[103]), .SEL(m_address[2]), .F(
        \u_a23_mem/n23332 ) );
  MUX \u_a23_mem/U23473  ( .IN0(\u_a23_mem/n23324 ), .IN1(\u_a23_mem/n23317 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23325 ) );
  MUX \u_a23_mem/U23472  ( .IN0(o[135]), .IN1(o[167]), .SEL(m_address[2]), .F(
        \u_a23_mem/n23324 ) );
  MUX \u_a23_mem/U23465  ( .IN0(o[199]), .IN1(o[231]), .SEL(m_address[2]), .F(
        \u_a23_mem/n23317 ) );
  MUX \u_a23_mem/U23458  ( .IN0(\u_a23_mem/n23310 ), .IN1(\u_a23_mem/n23295 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/N1936 ) );
  MUX \u_a23_mem/U23457  ( .IN0(\u_a23_mem/n23309 ), .IN1(\u_a23_mem/n23302 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23310 ) );
  MUX \u_a23_mem/U23456  ( .IN0(o[6]), .IN1(o[38]), .SEL(m_address[2]), .F(
        \u_a23_mem/n23309 ) );
  MUX \u_a23_mem/U23449  ( .IN0(o[70]), .IN1(o[102]), .SEL(m_address[2]), .F(
        \u_a23_mem/n23302 ) );
  MUX \u_a23_mem/U23442  ( .IN0(\u_a23_mem/n23294 ), .IN1(\u_a23_mem/n23287 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23295 ) );
  MUX \u_a23_mem/U23441  ( .IN0(o[134]), .IN1(o[166]), .SEL(m_address[2]), .F(
        \u_a23_mem/n23294 ) );
  MUX \u_a23_mem/U23434  ( .IN0(o[198]), .IN1(o[230]), .SEL(m_address[2]), .F(
        \u_a23_mem/n23287 ) );
  MUX \u_a23_mem/U23427  ( .IN0(\u_a23_mem/n23280 ), .IN1(\u_a23_mem/n23265 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/N1937 ) );
  MUX \u_a23_mem/U23426  ( .IN0(\u_a23_mem/n23279 ), .IN1(\u_a23_mem/n23272 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23280 ) );
  MUX \u_a23_mem/U23425  ( .IN0(o[5]), .IN1(o[37]), .SEL(m_address[2]), .F(
        \u_a23_mem/n23279 ) );
  MUX \u_a23_mem/U23418  ( .IN0(o[69]), .IN1(o[101]), .SEL(m_address[2]), .F(
        \u_a23_mem/n23272 ) );
  MUX \u_a23_mem/U23411  ( .IN0(\u_a23_mem/n23264 ), .IN1(\u_a23_mem/n23257 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23265 ) );
  MUX \u_a23_mem/U23410  ( .IN0(o[133]), .IN1(o[165]), .SEL(m_address[2]), .F(
        \u_a23_mem/n23264 ) );
  MUX \u_a23_mem/U23403  ( .IN0(o[197]), .IN1(o[229]), .SEL(m_address[2]), .F(
        \u_a23_mem/n23257 ) );
  MUX \u_a23_mem/U23396  ( .IN0(\u_a23_mem/n23250 ), .IN1(\u_a23_mem/n23235 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/N1938 ) );
  MUX \u_a23_mem/U23395  ( .IN0(\u_a23_mem/n23249 ), .IN1(\u_a23_mem/n23242 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23250 ) );
  MUX \u_a23_mem/U23394  ( .IN0(o[4]), .IN1(o[36]), .SEL(m_address[2]), .F(
        \u_a23_mem/n23249 ) );
  MUX \u_a23_mem/U23387  ( .IN0(o[68]), .IN1(o[100]), .SEL(m_address[2]), .F(
        \u_a23_mem/n23242 ) );
  MUX \u_a23_mem/U23380  ( .IN0(\u_a23_mem/n23234 ), .IN1(\u_a23_mem/n23227 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23235 ) );
  MUX \u_a23_mem/U23379  ( .IN0(o[132]), .IN1(o[164]), .SEL(m_address[2]), .F(
        \u_a23_mem/n23234 ) );
  MUX \u_a23_mem/U23372  ( .IN0(o[196]), .IN1(o[228]), .SEL(m_address[2]), .F(
        \u_a23_mem/n23227 ) );
  MUX \u_a23_mem/U23365  ( .IN0(\u_a23_mem/n23220 ), .IN1(\u_a23_mem/n23205 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/N1939 ) );
  MUX \u_a23_mem/U23364  ( .IN0(\u_a23_mem/n23219 ), .IN1(\u_a23_mem/n23212 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23220 ) );
  MUX \u_a23_mem/U23363  ( .IN0(o[3]), .IN1(o[35]), .SEL(m_address[2]), .F(
        \u_a23_mem/n23219 ) );
  MUX \u_a23_mem/U23356  ( .IN0(o[67]), .IN1(o[99]), .SEL(m_address[2]), .F(
        \u_a23_mem/n23212 ) );
  MUX \u_a23_mem/U23349  ( .IN0(\u_a23_mem/n23204 ), .IN1(\u_a23_mem/n23197 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23205 ) );
  MUX \u_a23_mem/U23348  ( .IN0(o[131]), .IN1(o[163]), .SEL(m_address[2]), .F(
        \u_a23_mem/n23204 ) );
  MUX \u_a23_mem/U23341  ( .IN0(o[195]), .IN1(o[227]), .SEL(m_address[2]), .F(
        \u_a23_mem/n23197 ) );
  MUX \u_a23_mem/U23334  ( .IN0(\u_a23_mem/n23190 ), .IN1(\u_a23_mem/n23175 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/N1940 ) );
  MUX \u_a23_mem/U23333  ( .IN0(\u_a23_mem/n23189 ), .IN1(\u_a23_mem/n23182 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23190 ) );
  MUX \u_a23_mem/U23332  ( .IN0(o[2]), .IN1(o[34]), .SEL(m_address[2]), .F(
        \u_a23_mem/n23189 ) );
  MUX \u_a23_mem/U23325  ( .IN0(o[66]), .IN1(o[98]), .SEL(m_address[2]), .F(
        \u_a23_mem/n23182 ) );
  MUX \u_a23_mem/U23318  ( .IN0(\u_a23_mem/n23174 ), .IN1(\u_a23_mem/n23167 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23175 ) );
  MUX \u_a23_mem/U23317  ( .IN0(o[130]), .IN1(o[162]), .SEL(m_address[2]), .F(
        \u_a23_mem/n23174 ) );
  MUX \u_a23_mem/U23310  ( .IN0(o[194]), .IN1(o[226]), .SEL(m_address[2]), .F(
        \u_a23_mem/n23167 ) );
  MUX \u_a23_mem/U23303  ( .IN0(\u_a23_mem/n23160 ), .IN1(\u_a23_mem/n23145 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/N1941 ) );
  MUX \u_a23_mem/U23302  ( .IN0(\u_a23_mem/n23159 ), .IN1(\u_a23_mem/n23152 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23160 ) );
  MUX \u_a23_mem/U23301  ( .IN0(o[1]), .IN1(o[33]), .SEL(m_address[2]), .F(
        \u_a23_mem/n23159 ) );
  MUX \u_a23_mem/U23294  ( .IN0(o[65]), .IN1(o[97]), .SEL(m_address[2]), .F(
        \u_a23_mem/n23152 ) );
  MUX \u_a23_mem/U23287  ( .IN0(\u_a23_mem/n23144 ), .IN1(\u_a23_mem/n23137 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23145 ) );
  MUX \u_a23_mem/U23286  ( .IN0(o[129]), .IN1(o[161]), .SEL(m_address[2]), .F(
        \u_a23_mem/n23144 ) );
  MUX \u_a23_mem/U23279  ( .IN0(o[193]), .IN1(o[225]), .SEL(m_address[2]), .F(
        \u_a23_mem/n23137 ) );
  MUX \u_a23_mem/U23272  ( .IN0(\u_a23_mem/n23130 ), .IN1(\u_a23_mem/n23115 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/N1942 ) );
  MUX \u_a23_mem/U23271  ( .IN0(\u_a23_mem/n23129 ), .IN1(\u_a23_mem/n23122 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23130 ) );
  MUX \u_a23_mem/U23270  ( .IN0(o[0]), .IN1(o[32]), .SEL(m_address[2]), .F(
        \u_a23_mem/n23129 ) );
  MUX \u_a23_mem/U23263  ( .IN0(o[64]), .IN1(o[96]), .SEL(m_address[2]), .F(
        \u_a23_mem/n23122 ) );
  MUX \u_a23_mem/U23256  ( .IN0(\u_a23_mem/n23114 ), .IN1(\u_a23_mem/n23107 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23115 ) );
  MUX \u_a23_mem/U23255  ( .IN0(o[128]), .IN1(o[160]), .SEL(m_address[2]), .F(
        \u_a23_mem/n23114 ) );
  MUX \u_a23_mem/U23248  ( .IN0(o[192]), .IN1(o[224]), .SEL(m_address[2]), .F(
        \u_a23_mem/n23107 ) );
  MUX \u_a23_mem/U23241  ( .IN0(\u_a23_mem/n23100 ), .IN1(\u_a23_mem/n23085 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/N1967 ) );
  MUX \u_a23_mem/U23240  ( .IN0(\u_a23_mem/n23099 ), .IN1(\u_a23_mem/n23092 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23100 ) );
  MUX \u_a23_mem/U23239  ( .IN0(\u_a23_mem/stack_mem[0][7] ), .IN1(
        \u_a23_mem/stack_mem[4][7] ), .SEL(m_address[2]), .F(
        \u_a23_mem/n23099 ) );
  MUX \u_a23_mem/U23232  ( .IN0(\u_a23_mem/stack_mem[8][7] ), .IN1(
        \u_a23_mem/stack_mem[12][7] ), .SEL(m_address[2]), .F(
        \u_a23_mem/n23092 ) );
  MUX \u_a23_mem/U23225  ( .IN0(\u_a23_mem/n23084 ), .IN1(\u_a23_mem/n23077 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23085 ) );
  MUX \u_a23_mem/U23224  ( .IN0(\u_a23_mem/stack_mem[16][7] ), .IN1(
        \u_a23_mem/stack_mem[20][7] ), .SEL(m_address[2]), .F(
        \u_a23_mem/n23084 ) );
  MUX \u_a23_mem/U23217  ( .IN0(\u_a23_mem/stack_mem[24][7] ), .IN1(
        \u_a23_mem/stack_mem[28][7] ), .SEL(m_address[2]), .F(
        \u_a23_mem/n23077 ) );
  MUX \u_a23_mem/U23210  ( .IN0(\u_a23_mem/n23070 ), .IN1(\u_a23_mem/n23055 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/N1968 ) );
  MUX \u_a23_mem/U23209  ( .IN0(\u_a23_mem/n23069 ), .IN1(\u_a23_mem/n23062 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23070 ) );
  MUX \u_a23_mem/U23208  ( .IN0(\u_a23_mem/stack_mem[0][6] ), .IN1(
        \u_a23_mem/stack_mem[4][6] ), .SEL(m_address[2]), .F(
        \u_a23_mem/n23069 ) );
  MUX \u_a23_mem/U23201  ( .IN0(\u_a23_mem/stack_mem[8][6] ), .IN1(
        \u_a23_mem/stack_mem[12][6] ), .SEL(m_address[2]), .F(
        \u_a23_mem/n23062 ) );
  MUX \u_a23_mem/U23194  ( .IN0(\u_a23_mem/n23054 ), .IN1(\u_a23_mem/n23047 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23055 ) );
  MUX \u_a23_mem/U23193  ( .IN0(\u_a23_mem/stack_mem[16][6] ), .IN1(
        \u_a23_mem/stack_mem[20][6] ), .SEL(m_address[2]), .F(
        \u_a23_mem/n23054 ) );
  MUX \u_a23_mem/U23186  ( .IN0(\u_a23_mem/stack_mem[24][6] ), .IN1(
        \u_a23_mem/stack_mem[28][6] ), .SEL(m_address[2]), .F(
        \u_a23_mem/n23047 ) );
  MUX \u_a23_mem/U23179  ( .IN0(\u_a23_mem/n23040 ), .IN1(\u_a23_mem/n23025 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/N1969 ) );
  MUX \u_a23_mem/U23178  ( .IN0(\u_a23_mem/n23039 ), .IN1(\u_a23_mem/n23032 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23040 ) );
  MUX \u_a23_mem/U23177  ( .IN0(\u_a23_mem/stack_mem[0][5] ), .IN1(
        \u_a23_mem/stack_mem[4][5] ), .SEL(m_address[2]), .F(
        \u_a23_mem/n23039 ) );
  MUX \u_a23_mem/U23170  ( .IN0(\u_a23_mem/stack_mem[8][5] ), .IN1(
        \u_a23_mem/stack_mem[12][5] ), .SEL(m_address[2]), .F(
        \u_a23_mem/n23032 ) );
  MUX \u_a23_mem/U23163  ( .IN0(\u_a23_mem/n23024 ), .IN1(\u_a23_mem/n23017 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23025 ) );
  MUX \u_a23_mem/U23162  ( .IN0(\u_a23_mem/stack_mem[16][5] ), .IN1(
        \u_a23_mem/stack_mem[20][5] ), .SEL(m_address[2]), .F(
        \u_a23_mem/n23024 ) );
  MUX \u_a23_mem/U23155  ( .IN0(\u_a23_mem/stack_mem[24][5] ), .IN1(
        \u_a23_mem/stack_mem[28][5] ), .SEL(m_address[2]), .F(
        \u_a23_mem/n23017 ) );
  MUX \u_a23_mem/U23148  ( .IN0(\u_a23_mem/n23010 ), .IN1(\u_a23_mem/n22995 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/N1970 ) );
  MUX \u_a23_mem/U23147  ( .IN0(\u_a23_mem/n23009 ), .IN1(\u_a23_mem/n23002 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n23010 ) );
  MUX \u_a23_mem/U23146  ( .IN0(\u_a23_mem/stack_mem[0][4] ), .IN1(
        \u_a23_mem/stack_mem[4][4] ), .SEL(m_address[2]), .F(
        \u_a23_mem/n23009 ) );
  MUX \u_a23_mem/U23139  ( .IN0(\u_a23_mem/stack_mem[8][4] ), .IN1(
        \u_a23_mem/stack_mem[12][4] ), .SEL(m_address[2]), .F(
        \u_a23_mem/n23002 ) );
  MUX \u_a23_mem/U23132  ( .IN0(\u_a23_mem/n22994 ), .IN1(\u_a23_mem/n22987 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22995 ) );
  MUX \u_a23_mem/U23131  ( .IN0(\u_a23_mem/stack_mem[16][4] ), .IN1(
        \u_a23_mem/stack_mem[20][4] ), .SEL(m_address[2]), .F(
        \u_a23_mem/n22994 ) );
  MUX \u_a23_mem/U23124  ( .IN0(\u_a23_mem/stack_mem[24][4] ), .IN1(
        \u_a23_mem/stack_mem[28][4] ), .SEL(m_address[2]), .F(
        \u_a23_mem/n22987 ) );
  MUX \u_a23_mem/U23117  ( .IN0(\u_a23_mem/n22980 ), .IN1(\u_a23_mem/n22965 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/N1971 ) );
  MUX \u_a23_mem/U23116  ( .IN0(\u_a23_mem/n22979 ), .IN1(\u_a23_mem/n22972 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22980 ) );
  MUX \u_a23_mem/U23115  ( .IN0(\u_a23_mem/stack_mem[0][3] ), .IN1(
        \u_a23_mem/stack_mem[4][3] ), .SEL(m_address[2]), .F(
        \u_a23_mem/n22979 ) );
  MUX \u_a23_mem/U23108  ( .IN0(\u_a23_mem/stack_mem[8][3] ), .IN1(
        \u_a23_mem/stack_mem[12][3] ), .SEL(m_address[2]), .F(
        \u_a23_mem/n22972 ) );
  MUX \u_a23_mem/U23101  ( .IN0(\u_a23_mem/n22964 ), .IN1(\u_a23_mem/n22957 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22965 ) );
  MUX \u_a23_mem/U23100  ( .IN0(\u_a23_mem/stack_mem[16][3] ), .IN1(
        \u_a23_mem/stack_mem[20][3] ), .SEL(m_address[2]), .F(
        \u_a23_mem/n22964 ) );
  MUX \u_a23_mem/U23093  ( .IN0(\u_a23_mem/stack_mem[24][3] ), .IN1(
        \u_a23_mem/stack_mem[28][3] ), .SEL(m_address[2]), .F(
        \u_a23_mem/n22957 ) );
  MUX \u_a23_mem/U23086  ( .IN0(\u_a23_mem/n22950 ), .IN1(\u_a23_mem/n22935 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/N1972 ) );
  MUX \u_a23_mem/U23085  ( .IN0(\u_a23_mem/n22949 ), .IN1(\u_a23_mem/n22942 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22950 ) );
  MUX \u_a23_mem/U23084  ( .IN0(\u_a23_mem/stack_mem[0][2] ), .IN1(
        \u_a23_mem/stack_mem[4][2] ), .SEL(m_address[2]), .F(
        \u_a23_mem/n22949 ) );
  MUX \u_a23_mem/U23077  ( .IN0(\u_a23_mem/stack_mem[8][2] ), .IN1(
        \u_a23_mem/stack_mem[12][2] ), .SEL(m_address[2]), .F(
        \u_a23_mem/n22942 ) );
  MUX \u_a23_mem/U23070  ( .IN0(\u_a23_mem/n22934 ), .IN1(\u_a23_mem/n22927 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22935 ) );
  MUX \u_a23_mem/U23069  ( .IN0(\u_a23_mem/stack_mem[16][2] ), .IN1(
        \u_a23_mem/stack_mem[20][2] ), .SEL(m_address[2]), .F(
        \u_a23_mem/n22934 ) );
  MUX \u_a23_mem/U23062  ( .IN0(\u_a23_mem/stack_mem[24][2] ), .IN1(
        \u_a23_mem/stack_mem[28][2] ), .SEL(m_address[2]), .F(
        \u_a23_mem/n22927 ) );
  MUX \u_a23_mem/U23055  ( .IN0(\u_a23_mem/n22920 ), .IN1(\u_a23_mem/n22905 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/N1973 ) );
  MUX \u_a23_mem/U23054  ( .IN0(\u_a23_mem/n22919 ), .IN1(\u_a23_mem/n22912 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22920 ) );
  MUX \u_a23_mem/U23053  ( .IN0(\u_a23_mem/stack_mem[0][1] ), .IN1(
        \u_a23_mem/stack_mem[4][1] ), .SEL(m_address[2]), .F(
        \u_a23_mem/n22919 ) );
  MUX \u_a23_mem/U23046  ( .IN0(\u_a23_mem/stack_mem[8][1] ), .IN1(
        \u_a23_mem/stack_mem[12][1] ), .SEL(m_address[2]), .F(
        \u_a23_mem/n22912 ) );
  MUX \u_a23_mem/U23039  ( .IN0(\u_a23_mem/n22904 ), .IN1(\u_a23_mem/n22897 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22905 ) );
  MUX \u_a23_mem/U23038  ( .IN0(\u_a23_mem/stack_mem[16][1] ), .IN1(
        \u_a23_mem/stack_mem[20][1] ), .SEL(m_address[2]), .F(
        \u_a23_mem/n22904 ) );
  MUX \u_a23_mem/U23031  ( .IN0(\u_a23_mem/stack_mem[24][1] ), .IN1(
        \u_a23_mem/stack_mem[28][1] ), .SEL(m_address[2]), .F(
        \u_a23_mem/n22897 ) );
  MUX \u_a23_mem/U23024  ( .IN0(\u_a23_mem/n22890 ), .IN1(\u_a23_mem/n22875 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/N1974 ) );
  MUX \u_a23_mem/U23023  ( .IN0(\u_a23_mem/n22889 ), .IN1(\u_a23_mem/n22882 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22890 ) );
  MUX \u_a23_mem/U23022  ( .IN0(\u_a23_mem/stack_mem[0][0] ), .IN1(
        \u_a23_mem/stack_mem[4][0] ), .SEL(m_address[2]), .F(
        \u_a23_mem/n22889 ) );
  MUX \u_a23_mem/U23015  ( .IN0(\u_a23_mem/stack_mem[8][0] ), .IN1(
        \u_a23_mem/stack_mem[12][0] ), .SEL(m_address[2]), .F(
        \u_a23_mem/n22882 ) );
  MUX \u_a23_mem/U23008  ( .IN0(\u_a23_mem/n22874 ), .IN1(\u_a23_mem/n22867 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22875 ) );
  MUX \u_a23_mem/U23007  ( .IN0(\u_a23_mem/stack_mem[16][0] ), .IN1(
        \u_a23_mem/stack_mem[20][0] ), .SEL(m_address[2]), .F(
        \u_a23_mem/n22874 ) );
  MUX \u_a23_mem/U23000  ( .IN0(\u_a23_mem/stack_mem[24][0] ), .IN1(
        \u_a23_mem/stack_mem[28][0] ), .SEL(m_address[2]), .F(
        \u_a23_mem/n22867 ) );
  MUX \u_a23_mem/U22993  ( .IN0(\u_a23_mem/n22860 ), .IN1(\u_a23_mem/n22797 ), 
        .SEL(m_address[6]), .F(\u_a23_mem/N1839 ) );
  MUX \u_a23_mem/U22992  ( .IN0(\u_a23_mem/n22859 ), .IN1(\u_a23_mem/n22828 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n22860 ) );
  MUX \u_a23_mem/U22991  ( .IN0(\u_a23_mem/n22858 ), .IN1(\u_a23_mem/n22843 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n22859 ) );
  MUX \u_a23_mem/U22990  ( .IN0(\u_a23_mem/n22857 ), .IN1(\u_a23_mem/n22850 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22858 ) );
  MUX \u_a23_mem/U22989  ( .IN0(\u_a23_mem/p_mem[0][7] ), .IN1(
        \u_a23_mem/p_mem[4][7] ), .SEL(m_address[2]), .F(\u_a23_mem/n22857 )
         );
  MUX \u_a23_mem/U22982  ( .IN0(\u_a23_mem/p_mem[8][7] ), .IN1(
        \u_a23_mem/p_mem[12][7] ), .SEL(m_address[2]), .F(\u_a23_mem/n22850 )
         );
  MUX \u_a23_mem/U22975  ( .IN0(\u_a23_mem/n22842 ), .IN1(\u_a23_mem/n22835 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22843 ) );
  MUX \u_a23_mem/U22974  ( .IN0(\u_a23_mem/p_mem[16][7] ), .IN1(
        \u_a23_mem/p_mem[20][7] ), .SEL(m_address[2]), .F(\u_a23_mem/n22842 )
         );
  MUX \u_a23_mem/U22967  ( .IN0(\u_a23_mem/p_mem[24][7] ), .IN1(
        \u_a23_mem/p_mem[28][7] ), .SEL(m_address[2]), .F(\u_a23_mem/n22835 )
         );
  MUX \u_a23_mem/U22960  ( .IN0(\u_a23_mem/n22827 ), .IN1(\u_a23_mem/n22812 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n22828 ) );
  MUX \u_a23_mem/U22959  ( .IN0(\u_a23_mem/n22826 ), .IN1(\u_a23_mem/n22819 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22827 ) );
  MUX \u_a23_mem/U22958  ( .IN0(\u_a23_mem/p_mem[32][7] ), .IN1(
        \u_a23_mem/p_mem[36][7] ), .SEL(m_address[2]), .F(\u_a23_mem/n22826 )
         );
  MUX \u_a23_mem/U22951  ( .IN0(\u_a23_mem/p_mem[40][7] ), .IN1(
        \u_a23_mem/p_mem[44][7] ), .SEL(m_address[2]), .F(\u_a23_mem/n22819 )
         );
  MUX \u_a23_mem/U22944  ( .IN0(\u_a23_mem/n22811 ), .IN1(\u_a23_mem/n22804 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22812 ) );
  MUX \u_a23_mem/U22943  ( .IN0(\u_a23_mem/p_mem[48][7] ), .IN1(
        \u_a23_mem/p_mem[52][7] ), .SEL(m_address[2]), .F(\u_a23_mem/n22811 )
         );
  MUX \u_a23_mem/U22936  ( .IN0(\u_a23_mem/p_mem[56][7] ), .IN1(
        \u_a23_mem/p_mem[60][7] ), .SEL(m_address[2]), .F(\u_a23_mem/n22804 )
         );
  MUX \u_a23_mem/U22929  ( .IN0(\u_a23_mem/n22796 ), .IN1(\u_a23_mem/n22765 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n22797 ) );
  MUX \u_a23_mem/U22928  ( .IN0(\u_a23_mem/n22795 ), .IN1(\u_a23_mem/n22780 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n22796 ) );
  MUX \u_a23_mem/U22927  ( .IN0(\u_a23_mem/n22794 ), .IN1(\u_a23_mem/n22787 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22795 ) );
  MUX \u_a23_mem/U22926  ( .IN0(\u_a23_mem/p_mem[64][7] ), .IN1(
        \u_a23_mem/p_mem[68][7] ), .SEL(m_address[2]), .F(\u_a23_mem/n22794 )
         );
  MUX \u_a23_mem/U22919  ( .IN0(\u_a23_mem/p_mem[72][7] ), .IN1(
        \u_a23_mem/p_mem[76][7] ), .SEL(m_address[2]), .F(\u_a23_mem/n22787 )
         );
  MUX \u_a23_mem/U22912  ( .IN0(\u_a23_mem/n22779 ), .IN1(\u_a23_mem/n22772 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22780 ) );
  MUX \u_a23_mem/U22911  ( .IN0(\u_a23_mem/p_mem[80][7] ), .IN1(
        \u_a23_mem/p_mem[84][7] ), .SEL(m_address[2]), .F(\u_a23_mem/n22779 )
         );
  MUX \u_a23_mem/U22904  ( .IN0(\u_a23_mem/p_mem[88][7] ), .IN1(
        \u_a23_mem/p_mem[92][7] ), .SEL(m_address[2]), .F(\u_a23_mem/n22772 )
         );
  MUX \u_a23_mem/U22897  ( .IN0(\u_a23_mem/n22764 ), .IN1(\u_a23_mem/n22749 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n22765 ) );
  MUX \u_a23_mem/U22896  ( .IN0(\u_a23_mem/n22763 ), .IN1(\u_a23_mem/n22756 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22764 ) );
  MUX \u_a23_mem/U22895  ( .IN0(\u_a23_mem/p_mem[96][7] ), .IN1(
        \u_a23_mem/p_mem[100][7] ), .SEL(m_address[2]), .F(\u_a23_mem/n22763 )
         );
  MUX \u_a23_mem/U22888  ( .IN0(\u_a23_mem/p_mem[104][7] ), .IN1(
        \u_a23_mem/p_mem[108][7] ), .SEL(m_address[2]), .F(\u_a23_mem/n22756 )
         );
  MUX \u_a23_mem/U22881  ( .IN0(\u_a23_mem/n22748 ), .IN1(\u_a23_mem/n22741 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22749 ) );
  MUX \u_a23_mem/U22880  ( .IN0(\u_a23_mem/p_mem[112][7] ), .IN1(
        \u_a23_mem/p_mem[116][7] ), .SEL(m_address[2]), .F(\u_a23_mem/n22748 )
         );
  MUX \u_a23_mem/U22873  ( .IN0(\u_a23_mem/p_mem[120][7] ), .IN1(
        \u_a23_mem/p_mem[124][7] ), .SEL(m_address[2]), .F(\u_a23_mem/n22741 )
         );
  MUX \u_a23_mem/U22866  ( .IN0(\u_a23_mem/n22734 ), .IN1(\u_a23_mem/n22671 ), 
        .SEL(m_address[6]), .F(\u_a23_mem/N1840 ) );
  MUX \u_a23_mem/U22865  ( .IN0(\u_a23_mem/n22733 ), .IN1(\u_a23_mem/n22702 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n22734 ) );
  MUX \u_a23_mem/U22864  ( .IN0(\u_a23_mem/n22732 ), .IN1(\u_a23_mem/n22717 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n22733 ) );
  MUX \u_a23_mem/U22863  ( .IN0(\u_a23_mem/n22731 ), .IN1(\u_a23_mem/n22724 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22732 ) );
  MUX \u_a23_mem/U22862  ( .IN0(\u_a23_mem/p_mem[0][6] ), .IN1(
        \u_a23_mem/p_mem[4][6] ), .SEL(m_address[2]), .F(\u_a23_mem/n22731 )
         );
  MUX \u_a23_mem/U22855  ( .IN0(\u_a23_mem/p_mem[8][6] ), .IN1(
        \u_a23_mem/p_mem[12][6] ), .SEL(m_address[2]), .F(\u_a23_mem/n22724 )
         );
  MUX \u_a23_mem/U22848  ( .IN0(\u_a23_mem/n22716 ), .IN1(\u_a23_mem/n22709 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22717 ) );
  MUX \u_a23_mem/U22847  ( .IN0(\u_a23_mem/p_mem[16][6] ), .IN1(
        \u_a23_mem/p_mem[20][6] ), .SEL(m_address[2]), .F(\u_a23_mem/n22716 )
         );
  MUX \u_a23_mem/U22840  ( .IN0(\u_a23_mem/p_mem[24][6] ), .IN1(
        \u_a23_mem/p_mem[28][6] ), .SEL(m_address[2]), .F(\u_a23_mem/n22709 )
         );
  MUX \u_a23_mem/U22833  ( .IN0(\u_a23_mem/n22701 ), .IN1(\u_a23_mem/n22686 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n22702 ) );
  MUX \u_a23_mem/U22832  ( .IN0(\u_a23_mem/n22700 ), .IN1(\u_a23_mem/n22693 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22701 ) );
  MUX \u_a23_mem/U22831  ( .IN0(\u_a23_mem/p_mem[32][6] ), .IN1(
        \u_a23_mem/p_mem[36][6] ), .SEL(m_address[2]), .F(\u_a23_mem/n22700 )
         );
  MUX \u_a23_mem/U22824  ( .IN0(\u_a23_mem/p_mem[40][6] ), .IN1(
        \u_a23_mem/p_mem[44][6] ), .SEL(m_address[2]), .F(\u_a23_mem/n22693 )
         );
  MUX \u_a23_mem/U22817  ( .IN0(\u_a23_mem/n22685 ), .IN1(\u_a23_mem/n22678 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22686 ) );
  MUX \u_a23_mem/U22816  ( .IN0(\u_a23_mem/p_mem[48][6] ), .IN1(
        \u_a23_mem/p_mem[52][6] ), .SEL(m_address[2]), .F(\u_a23_mem/n22685 )
         );
  MUX \u_a23_mem/U22809  ( .IN0(\u_a23_mem/p_mem[56][6] ), .IN1(
        \u_a23_mem/p_mem[60][6] ), .SEL(m_address[2]), .F(\u_a23_mem/n22678 )
         );
  MUX \u_a23_mem/U22802  ( .IN0(\u_a23_mem/n22670 ), .IN1(\u_a23_mem/n22639 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n22671 ) );
  MUX \u_a23_mem/U22801  ( .IN0(\u_a23_mem/n22669 ), .IN1(\u_a23_mem/n22654 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n22670 ) );
  MUX \u_a23_mem/U22800  ( .IN0(\u_a23_mem/n22668 ), .IN1(\u_a23_mem/n22661 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22669 ) );
  MUX \u_a23_mem/U22799  ( .IN0(\u_a23_mem/p_mem[64][6] ), .IN1(
        \u_a23_mem/p_mem[68][6] ), .SEL(m_address[2]), .F(\u_a23_mem/n22668 )
         );
  MUX \u_a23_mem/U22792  ( .IN0(\u_a23_mem/p_mem[72][6] ), .IN1(
        \u_a23_mem/p_mem[76][6] ), .SEL(m_address[2]), .F(\u_a23_mem/n22661 )
         );
  MUX \u_a23_mem/U22785  ( .IN0(\u_a23_mem/n22653 ), .IN1(\u_a23_mem/n22646 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22654 ) );
  MUX \u_a23_mem/U22784  ( .IN0(\u_a23_mem/p_mem[80][6] ), .IN1(
        \u_a23_mem/p_mem[84][6] ), .SEL(m_address[2]), .F(\u_a23_mem/n22653 )
         );
  MUX \u_a23_mem/U22777  ( .IN0(\u_a23_mem/p_mem[88][6] ), .IN1(
        \u_a23_mem/p_mem[92][6] ), .SEL(m_address[2]), .F(\u_a23_mem/n22646 )
         );
  MUX \u_a23_mem/U22770  ( .IN0(\u_a23_mem/n22638 ), .IN1(\u_a23_mem/n22623 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n22639 ) );
  MUX \u_a23_mem/U22769  ( .IN0(\u_a23_mem/n22637 ), .IN1(\u_a23_mem/n22630 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22638 ) );
  MUX \u_a23_mem/U22768  ( .IN0(\u_a23_mem/p_mem[96][6] ), .IN1(
        \u_a23_mem/p_mem[100][6] ), .SEL(m_address[2]), .F(\u_a23_mem/n22637 )
         );
  MUX \u_a23_mem/U22761  ( .IN0(\u_a23_mem/p_mem[104][6] ), .IN1(
        \u_a23_mem/p_mem[108][6] ), .SEL(m_address[2]), .F(\u_a23_mem/n22630 )
         );
  MUX \u_a23_mem/U22754  ( .IN0(\u_a23_mem/n22622 ), .IN1(\u_a23_mem/n22615 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22623 ) );
  MUX \u_a23_mem/U22753  ( .IN0(\u_a23_mem/p_mem[112][6] ), .IN1(
        \u_a23_mem/p_mem[116][6] ), .SEL(m_address[2]), .F(\u_a23_mem/n22622 )
         );
  MUX \u_a23_mem/U22746  ( .IN0(\u_a23_mem/p_mem[120][6] ), .IN1(
        \u_a23_mem/p_mem[124][6] ), .SEL(m_address[2]), .F(\u_a23_mem/n22615 )
         );
  MUX \u_a23_mem/U22739  ( .IN0(\u_a23_mem/n22608 ), .IN1(\u_a23_mem/n22545 ), 
        .SEL(m_address[6]), .F(\u_a23_mem/N1841 ) );
  MUX \u_a23_mem/U22738  ( .IN0(\u_a23_mem/n22607 ), .IN1(\u_a23_mem/n22576 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n22608 ) );
  MUX \u_a23_mem/U22737  ( .IN0(\u_a23_mem/n22606 ), .IN1(\u_a23_mem/n22591 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n22607 ) );
  MUX \u_a23_mem/U22736  ( .IN0(\u_a23_mem/n22605 ), .IN1(\u_a23_mem/n22598 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22606 ) );
  MUX \u_a23_mem/U22735  ( .IN0(\u_a23_mem/p_mem[0][5] ), .IN1(
        \u_a23_mem/p_mem[4][5] ), .SEL(m_address[2]), .F(\u_a23_mem/n22605 )
         );
  MUX \u_a23_mem/U22728  ( .IN0(\u_a23_mem/p_mem[8][5] ), .IN1(
        \u_a23_mem/p_mem[12][5] ), .SEL(m_address[2]), .F(\u_a23_mem/n22598 )
         );
  MUX \u_a23_mem/U22721  ( .IN0(\u_a23_mem/n22590 ), .IN1(\u_a23_mem/n22583 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22591 ) );
  MUX \u_a23_mem/U22720  ( .IN0(\u_a23_mem/p_mem[16][5] ), .IN1(
        \u_a23_mem/p_mem[20][5] ), .SEL(m_address[2]), .F(\u_a23_mem/n22590 )
         );
  MUX \u_a23_mem/U22713  ( .IN0(\u_a23_mem/p_mem[24][5] ), .IN1(
        \u_a23_mem/p_mem[28][5] ), .SEL(m_address[2]), .F(\u_a23_mem/n22583 )
         );
  MUX \u_a23_mem/U22706  ( .IN0(\u_a23_mem/n22575 ), .IN1(\u_a23_mem/n22560 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n22576 ) );
  MUX \u_a23_mem/U22705  ( .IN0(\u_a23_mem/n22574 ), .IN1(\u_a23_mem/n22567 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22575 ) );
  MUX \u_a23_mem/U22704  ( .IN0(\u_a23_mem/p_mem[32][5] ), .IN1(
        \u_a23_mem/p_mem[36][5] ), .SEL(m_address[2]), .F(\u_a23_mem/n22574 )
         );
  MUX \u_a23_mem/U22697  ( .IN0(\u_a23_mem/p_mem[40][5] ), .IN1(
        \u_a23_mem/p_mem[44][5] ), .SEL(m_address[2]), .F(\u_a23_mem/n22567 )
         );
  MUX \u_a23_mem/U22690  ( .IN0(\u_a23_mem/n22559 ), .IN1(\u_a23_mem/n22552 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22560 ) );
  MUX \u_a23_mem/U22689  ( .IN0(\u_a23_mem/p_mem[48][5] ), .IN1(
        \u_a23_mem/p_mem[52][5] ), .SEL(m_address[2]), .F(\u_a23_mem/n22559 )
         );
  MUX \u_a23_mem/U22682  ( .IN0(\u_a23_mem/p_mem[56][5] ), .IN1(
        \u_a23_mem/p_mem[60][5] ), .SEL(m_address[2]), .F(\u_a23_mem/n22552 )
         );
  MUX \u_a23_mem/U22675  ( .IN0(\u_a23_mem/n22544 ), .IN1(\u_a23_mem/n22513 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n22545 ) );
  MUX \u_a23_mem/U22674  ( .IN0(\u_a23_mem/n22543 ), .IN1(\u_a23_mem/n22528 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n22544 ) );
  MUX \u_a23_mem/U22673  ( .IN0(\u_a23_mem/n22542 ), .IN1(\u_a23_mem/n22535 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22543 ) );
  MUX \u_a23_mem/U22672  ( .IN0(\u_a23_mem/p_mem[64][5] ), .IN1(
        \u_a23_mem/p_mem[68][5] ), .SEL(m_address[2]), .F(\u_a23_mem/n22542 )
         );
  MUX \u_a23_mem/U22665  ( .IN0(\u_a23_mem/p_mem[72][5] ), .IN1(
        \u_a23_mem/p_mem[76][5] ), .SEL(m_address[2]), .F(\u_a23_mem/n22535 )
         );
  MUX \u_a23_mem/U22658  ( .IN0(\u_a23_mem/n22527 ), .IN1(\u_a23_mem/n22520 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22528 ) );
  MUX \u_a23_mem/U22657  ( .IN0(\u_a23_mem/p_mem[80][5] ), .IN1(
        \u_a23_mem/p_mem[84][5] ), .SEL(m_address[2]), .F(\u_a23_mem/n22527 )
         );
  MUX \u_a23_mem/U22650  ( .IN0(\u_a23_mem/p_mem[88][5] ), .IN1(
        \u_a23_mem/p_mem[92][5] ), .SEL(m_address[2]), .F(\u_a23_mem/n22520 )
         );
  MUX \u_a23_mem/U22643  ( .IN0(\u_a23_mem/n22512 ), .IN1(\u_a23_mem/n22497 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n22513 ) );
  MUX \u_a23_mem/U22642  ( .IN0(\u_a23_mem/n22511 ), .IN1(\u_a23_mem/n22504 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22512 ) );
  MUX \u_a23_mem/U22641  ( .IN0(\u_a23_mem/p_mem[96][5] ), .IN1(
        \u_a23_mem/p_mem[100][5] ), .SEL(m_address[2]), .F(\u_a23_mem/n22511 )
         );
  MUX \u_a23_mem/U22634  ( .IN0(\u_a23_mem/p_mem[104][5] ), .IN1(
        \u_a23_mem/p_mem[108][5] ), .SEL(m_address[2]), .F(\u_a23_mem/n22504 )
         );
  MUX \u_a23_mem/U22627  ( .IN0(\u_a23_mem/n22496 ), .IN1(\u_a23_mem/n22489 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22497 ) );
  MUX \u_a23_mem/U22626  ( .IN0(\u_a23_mem/p_mem[112][5] ), .IN1(
        \u_a23_mem/p_mem[116][5] ), .SEL(m_address[2]), .F(\u_a23_mem/n22496 )
         );
  MUX \u_a23_mem/U22619  ( .IN0(\u_a23_mem/p_mem[120][5] ), .IN1(
        \u_a23_mem/p_mem[124][5] ), .SEL(m_address[2]), .F(\u_a23_mem/n22489 )
         );
  MUX \u_a23_mem/U22612  ( .IN0(\u_a23_mem/n22482 ), .IN1(\u_a23_mem/n22419 ), 
        .SEL(m_address[6]), .F(\u_a23_mem/N1842 ) );
  MUX \u_a23_mem/U22611  ( .IN0(\u_a23_mem/n22481 ), .IN1(\u_a23_mem/n22450 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n22482 ) );
  MUX \u_a23_mem/U22610  ( .IN0(\u_a23_mem/n22480 ), .IN1(\u_a23_mem/n22465 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n22481 ) );
  MUX \u_a23_mem/U22609  ( .IN0(\u_a23_mem/n22479 ), .IN1(\u_a23_mem/n22472 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22480 ) );
  MUX \u_a23_mem/U22608  ( .IN0(\u_a23_mem/p_mem[0][4] ), .IN1(
        \u_a23_mem/p_mem[4][4] ), .SEL(m_address[2]), .F(\u_a23_mem/n22479 )
         );
  MUX \u_a23_mem/U22601  ( .IN0(\u_a23_mem/p_mem[8][4] ), .IN1(
        \u_a23_mem/p_mem[12][4] ), .SEL(m_address[2]), .F(\u_a23_mem/n22472 )
         );
  MUX \u_a23_mem/U22594  ( .IN0(\u_a23_mem/n22464 ), .IN1(\u_a23_mem/n22457 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22465 ) );
  MUX \u_a23_mem/U22593  ( .IN0(\u_a23_mem/p_mem[16][4] ), .IN1(
        \u_a23_mem/p_mem[20][4] ), .SEL(m_address[2]), .F(\u_a23_mem/n22464 )
         );
  MUX \u_a23_mem/U22586  ( .IN0(\u_a23_mem/p_mem[24][4] ), .IN1(
        \u_a23_mem/p_mem[28][4] ), .SEL(m_address[2]), .F(\u_a23_mem/n22457 )
         );
  MUX \u_a23_mem/U22579  ( .IN0(\u_a23_mem/n22449 ), .IN1(\u_a23_mem/n22434 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n22450 ) );
  MUX \u_a23_mem/U22578  ( .IN0(\u_a23_mem/n22448 ), .IN1(\u_a23_mem/n22441 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22449 ) );
  MUX \u_a23_mem/U22577  ( .IN0(\u_a23_mem/p_mem[32][4] ), .IN1(
        \u_a23_mem/p_mem[36][4] ), .SEL(m_address[2]), .F(\u_a23_mem/n22448 )
         );
  MUX \u_a23_mem/U22570  ( .IN0(\u_a23_mem/p_mem[40][4] ), .IN1(
        \u_a23_mem/p_mem[44][4] ), .SEL(m_address[2]), .F(\u_a23_mem/n22441 )
         );
  MUX \u_a23_mem/U22563  ( .IN0(\u_a23_mem/n22433 ), .IN1(\u_a23_mem/n22426 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22434 ) );
  MUX \u_a23_mem/U22562  ( .IN0(\u_a23_mem/p_mem[48][4] ), .IN1(
        \u_a23_mem/p_mem[52][4] ), .SEL(m_address[2]), .F(\u_a23_mem/n22433 )
         );
  MUX \u_a23_mem/U22555  ( .IN0(\u_a23_mem/p_mem[56][4] ), .IN1(
        \u_a23_mem/p_mem[60][4] ), .SEL(m_address[2]), .F(\u_a23_mem/n22426 )
         );
  MUX \u_a23_mem/U22548  ( .IN0(\u_a23_mem/n22418 ), .IN1(\u_a23_mem/n22387 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n22419 ) );
  MUX \u_a23_mem/U22547  ( .IN0(\u_a23_mem/n22417 ), .IN1(\u_a23_mem/n22402 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n22418 ) );
  MUX \u_a23_mem/U22546  ( .IN0(\u_a23_mem/n22416 ), .IN1(\u_a23_mem/n22409 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22417 ) );
  MUX \u_a23_mem/U22545  ( .IN0(\u_a23_mem/p_mem[64][4] ), .IN1(
        \u_a23_mem/p_mem[68][4] ), .SEL(m_address[2]), .F(\u_a23_mem/n22416 )
         );
  MUX \u_a23_mem/U22538  ( .IN0(\u_a23_mem/p_mem[72][4] ), .IN1(
        \u_a23_mem/p_mem[76][4] ), .SEL(m_address[2]), .F(\u_a23_mem/n22409 )
         );
  MUX \u_a23_mem/U22531  ( .IN0(\u_a23_mem/n22401 ), .IN1(\u_a23_mem/n22394 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22402 ) );
  MUX \u_a23_mem/U22530  ( .IN0(\u_a23_mem/p_mem[80][4] ), .IN1(
        \u_a23_mem/p_mem[84][4] ), .SEL(m_address[2]), .F(\u_a23_mem/n22401 )
         );
  MUX \u_a23_mem/U22523  ( .IN0(\u_a23_mem/p_mem[88][4] ), .IN1(
        \u_a23_mem/p_mem[92][4] ), .SEL(m_address[2]), .F(\u_a23_mem/n22394 )
         );
  MUX \u_a23_mem/U22516  ( .IN0(\u_a23_mem/n22386 ), .IN1(\u_a23_mem/n22371 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n22387 ) );
  MUX \u_a23_mem/U22515  ( .IN0(\u_a23_mem/n22385 ), .IN1(\u_a23_mem/n22378 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22386 ) );
  MUX \u_a23_mem/U22514  ( .IN0(\u_a23_mem/p_mem[96][4] ), .IN1(
        \u_a23_mem/p_mem[100][4] ), .SEL(m_address[2]), .F(\u_a23_mem/n22385 )
         );
  MUX \u_a23_mem/U22507  ( .IN0(\u_a23_mem/p_mem[104][4] ), .IN1(
        \u_a23_mem/p_mem[108][4] ), .SEL(m_address[2]), .F(\u_a23_mem/n22378 )
         );
  MUX \u_a23_mem/U22500  ( .IN0(\u_a23_mem/n22370 ), .IN1(\u_a23_mem/n22363 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22371 ) );
  MUX \u_a23_mem/U22499  ( .IN0(\u_a23_mem/p_mem[112][4] ), .IN1(
        \u_a23_mem/p_mem[116][4] ), .SEL(m_address[2]), .F(\u_a23_mem/n22370 )
         );
  MUX \u_a23_mem/U22492  ( .IN0(\u_a23_mem/p_mem[120][4] ), .IN1(
        \u_a23_mem/p_mem[124][4] ), .SEL(m_address[2]), .F(\u_a23_mem/n22363 )
         );
  MUX \u_a23_mem/U22485  ( .IN0(\u_a23_mem/n22356 ), .IN1(\u_a23_mem/n22293 ), 
        .SEL(m_address[6]), .F(\u_a23_mem/N1843 ) );
  MUX \u_a23_mem/U22484  ( .IN0(\u_a23_mem/n22355 ), .IN1(\u_a23_mem/n22324 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n22356 ) );
  MUX \u_a23_mem/U22483  ( .IN0(\u_a23_mem/n22354 ), .IN1(\u_a23_mem/n22339 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n22355 ) );
  MUX \u_a23_mem/U22482  ( .IN0(\u_a23_mem/n22353 ), .IN1(\u_a23_mem/n22346 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22354 ) );
  MUX \u_a23_mem/U22481  ( .IN0(\u_a23_mem/p_mem[0][3] ), .IN1(
        \u_a23_mem/p_mem[4][3] ), .SEL(m_address[2]), .F(\u_a23_mem/n22353 )
         );
  MUX \u_a23_mem/U22474  ( .IN0(\u_a23_mem/p_mem[8][3] ), .IN1(
        \u_a23_mem/p_mem[12][3] ), .SEL(m_address[2]), .F(\u_a23_mem/n22346 )
         );
  MUX \u_a23_mem/U22467  ( .IN0(\u_a23_mem/n22338 ), .IN1(\u_a23_mem/n22331 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22339 ) );
  MUX \u_a23_mem/U22466  ( .IN0(\u_a23_mem/p_mem[16][3] ), .IN1(
        \u_a23_mem/p_mem[20][3] ), .SEL(m_address[2]), .F(\u_a23_mem/n22338 )
         );
  MUX \u_a23_mem/U22459  ( .IN0(\u_a23_mem/p_mem[24][3] ), .IN1(
        \u_a23_mem/p_mem[28][3] ), .SEL(m_address[2]), .F(\u_a23_mem/n22331 )
         );
  MUX \u_a23_mem/U22452  ( .IN0(\u_a23_mem/n22323 ), .IN1(\u_a23_mem/n22308 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n22324 ) );
  MUX \u_a23_mem/U22451  ( .IN0(\u_a23_mem/n22322 ), .IN1(\u_a23_mem/n22315 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22323 ) );
  MUX \u_a23_mem/U22450  ( .IN0(\u_a23_mem/p_mem[32][3] ), .IN1(
        \u_a23_mem/p_mem[36][3] ), .SEL(m_address[2]), .F(\u_a23_mem/n22322 )
         );
  MUX \u_a23_mem/U22443  ( .IN0(\u_a23_mem/p_mem[40][3] ), .IN1(
        \u_a23_mem/p_mem[44][3] ), .SEL(m_address[2]), .F(\u_a23_mem/n22315 )
         );
  MUX \u_a23_mem/U22436  ( .IN0(\u_a23_mem/n22307 ), .IN1(\u_a23_mem/n22300 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22308 ) );
  MUX \u_a23_mem/U22435  ( .IN0(\u_a23_mem/p_mem[48][3] ), .IN1(
        \u_a23_mem/p_mem[52][3] ), .SEL(m_address[2]), .F(\u_a23_mem/n22307 )
         );
  MUX \u_a23_mem/U22428  ( .IN0(\u_a23_mem/p_mem[56][3] ), .IN1(
        \u_a23_mem/p_mem[60][3] ), .SEL(m_address[2]), .F(\u_a23_mem/n22300 )
         );
  MUX \u_a23_mem/U22421  ( .IN0(\u_a23_mem/n22292 ), .IN1(\u_a23_mem/n22261 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n22293 ) );
  MUX \u_a23_mem/U22420  ( .IN0(\u_a23_mem/n22291 ), .IN1(\u_a23_mem/n22276 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n22292 ) );
  MUX \u_a23_mem/U22419  ( .IN0(\u_a23_mem/n22290 ), .IN1(\u_a23_mem/n22283 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22291 ) );
  MUX \u_a23_mem/U22418  ( .IN0(\u_a23_mem/p_mem[64][3] ), .IN1(
        \u_a23_mem/p_mem[68][3] ), .SEL(m_address[2]), .F(\u_a23_mem/n22290 )
         );
  MUX \u_a23_mem/U22411  ( .IN0(\u_a23_mem/p_mem[72][3] ), .IN1(
        \u_a23_mem/p_mem[76][3] ), .SEL(m_address[2]), .F(\u_a23_mem/n22283 )
         );
  MUX \u_a23_mem/U22404  ( .IN0(\u_a23_mem/n22275 ), .IN1(\u_a23_mem/n22268 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22276 ) );
  MUX \u_a23_mem/U22403  ( .IN0(\u_a23_mem/p_mem[80][3] ), .IN1(
        \u_a23_mem/p_mem[84][3] ), .SEL(m_address[2]), .F(\u_a23_mem/n22275 )
         );
  MUX \u_a23_mem/U22396  ( .IN0(\u_a23_mem/p_mem[88][3] ), .IN1(
        \u_a23_mem/p_mem[92][3] ), .SEL(m_address[2]), .F(\u_a23_mem/n22268 )
         );
  MUX \u_a23_mem/U22389  ( .IN0(\u_a23_mem/n22260 ), .IN1(\u_a23_mem/n22245 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n22261 ) );
  MUX \u_a23_mem/U22388  ( .IN0(\u_a23_mem/n22259 ), .IN1(\u_a23_mem/n22252 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22260 ) );
  MUX \u_a23_mem/U22387  ( .IN0(\u_a23_mem/p_mem[96][3] ), .IN1(
        \u_a23_mem/p_mem[100][3] ), .SEL(m_address[2]), .F(\u_a23_mem/n22259 )
         );
  MUX \u_a23_mem/U22380  ( .IN0(\u_a23_mem/p_mem[104][3] ), .IN1(
        \u_a23_mem/p_mem[108][3] ), .SEL(m_address[2]), .F(\u_a23_mem/n22252 )
         );
  MUX \u_a23_mem/U22373  ( .IN0(\u_a23_mem/n22244 ), .IN1(\u_a23_mem/n22237 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22245 ) );
  MUX \u_a23_mem/U22372  ( .IN0(\u_a23_mem/p_mem[112][3] ), .IN1(
        \u_a23_mem/p_mem[116][3] ), .SEL(m_address[2]), .F(\u_a23_mem/n22244 )
         );
  MUX \u_a23_mem/U22365  ( .IN0(\u_a23_mem/p_mem[120][3] ), .IN1(
        \u_a23_mem/p_mem[124][3] ), .SEL(m_address[2]), .F(\u_a23_mem/n22237 )
         );
  MUX \u_a23_mem/U22358  ( .IN0(\u_a23_mem/n22230 ), .IN1(\u_a23_mem/n22167 ), 
        .SEL(m_address[6]), .F(\u_a23_mem/N1844 ) );
  MUX \u_a23_mem/U22357  ( .IN0(\u_a23_mem/n22229 ), .IN1(\u_a23_mem/n22198 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n22230 ) );
  MUX \u_a23_mem/U22356  ( .IN0(\u_a23_mem/n22228 ), .IN1(\u_a23_mem/n22213 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n22229 ) );
  MUX \u_a23_mem/U22355  ( .IN0(\u_a23_mem/n22227 ), .IN1(\u_a23_mem/n22220 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22228 ) );
  MUX \u_a23_mem/U22354  ( .IN0(\u_a23_mem/p_mem[0][2] ), .IN1(
        \u_a23_mem/p_mem[4][2] ), .SEL(m_address[2]), .F(\u_a23_mem/n22227 )
         );
  MUX \u_a23_mem/U22347  ( .IN0(\u_a23_mem/p_mem[8][2] ), .IN1(
        \u_a23_mem/p_mem[12][2] ), .SEL(m_address[2]), .F(\u_a23_mem/n22220 )
         );
  MUX \u_a23_mem/U22340  ( .IN0(\u_a23_mem/n22212 ), .IN1(\u_a23_mem/n22205 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22213 ) );
  MUX \u_a23_mem/U22339  ( .IN0(\u_a23_mem/p_mem[16][2] ), .IN1(
        \u_a23_mem/p_mem[20][2] ), .SEL(m_address[2]), .F(\u_a23_mem/n22212 )
         );
  MUX \u_a23_mem/U22332  ( .IN0(\u_a23_mem/p_mem[24][2] ), .IN1(
        \u_a23_mem/p_mem[28][2] ), .SEL(m_address[2]), .F(\u_a23_mem/n22205 )
         );
  MUX \u_a23_mem/U22325  ( .IN0(\u_a23_mem/n22197 ), .IN1(\u_a23_mem/n22182 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n22198 ) );
  MUX \u_a23_mem/U22324  ( .IN0(\u_a23_mem/n22196 ), .IN1(\u_a23_mem/n22189 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22197 ) );
  MUX \u_a23_mem/U22323  ( .IN0(\u_a23_mem/p_mem[32][2] ), .IN1(
        \u_a23_mem/p_mem[36][2] ), .SEL(m_address[2]), .F(\u_a23_mem/n22196 )
         );
  MUX \u_a23_mem/U22316  ( .IN0(\u_a23_mem/p_mem[40][2] ), .IN1(
        \u_a23_mem/p_mem[44][2] ), .SEL(m_address[2]), .F(\u_a23_mem/n22189 )
         );
  MUX \u_a23_mem/U22309  ( .IN0(\u_a23_mem/n22181 ), .IN1(\u_a23_mem/n22174 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22182 ) );
  MUX \u_a23_mem/U22308  ( .IN0(\u_a23_mem/p_mem[48][2] ), .IN1(
        \u_a23_mem/p_mem[52][2] ), .SEL(m_address[2]), .F(\u_a23_mem/n22181 )
         );
  MUX \u_a23_mem/U22301  ( .IN0(\u_a23_mem/p_mem[56][2] ), .IN1(
        \u_a23_mem/p_mem[60][2] ), .SEL(m_address[2]), .F(\u_a23_mem/n22174 )
         );
  MUX \u_a23_mem/U22294  ( .IN0(\u_a23_mem/n22166 ), .IN1(\u_a23_mem/n22135 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n22167 ) );
  MUX \u_a23_mem/U22293  ( .IN0(\u_a23_mem/n22165 ), .IN1(\u_a23_mem/n22150 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n22166 ) );
  MUX \u_a23_mem/U22292  ( .IN0(\u_a23_mem/n22164 ), .IN1(\u_a23_mem/n22157 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22165 ) );
  MUX \u_a23_mem/U22291  ( .IN0(\u_a23_mem/p_mem[64][2] ), .IN1(
        \u_a23_mem/p_mem[68][2] ), .SEL(m_address[2]), .F(\u_a23_mem/n22164 )
         );
  MUX \u_a23_mem/U22284  ( .IN0(\u_a23_mem/p_mem[72][2] ), .IN1(
        \u_a23_mem/p_mem[76][2] ), .SEL(m_address[2]), .F(\u_a23_mem/n22157 )
         );
  MUX \u_a23_mem/U22277  ( .IN0(\u_a23_mem/n22149 ), .IN1(\u_a23_mem/n22142 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22150 ) );
  MUX \u_a23_mem/U22276  ( .IN0(\u_a23_mem/p_mem[80][2] ), .IN1(
        \u_a23_mem/p_mem[84][2] ), .SEL(m_address[2]), .F(\u_a23_mem/n22149 )
         );
  MUX \u_a23_mem/U22269  ( .IN0(\u_a23_mem/p_mem[88][2] ), .IN1(
        \u_a23_mem/p_mem[92][2] ), .SEL(m_address[2]), .F(\u_a23_mem/n22142 )
         );
  MUX \u_a23_mem/U22262  ( .IN0(\u_a23_mem/n22134 ), .IN1(\u_a23_mem/n22119 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n22135 ) );
  MUX \u_a23_mem/U22261  ( .IN0(\u_a23_mem/n22133 ), .IN1(\u_a23_mem/n22126 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22134 ) );
  MUX \u_a23_mem/U22260  ( .IN0(\u_a23_mem/p_mem[96][2] ), .IN1(
        \u_a23_mem/p_mem[100][2] ), .SEL(m_address[2]), .F(\u_a23_mem/n22133 )
         );
  MUX \u_a23_mem/U22253  ( .IN0(\u_a23_mem/p_mem[104][2] ), .IN1(
        \u_a23_mem/p_mem[108][2] ), .SEL(m_address[2]), .F(\u_a23_mem/n22126 )
         );
  MUX \u_a23_mem/U22246  ( .IN0(\u_a23_mem/n22118 ), .IN1(\u_a23_mem/n22111 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22119 ) );
  MUX \u_a23_mem/U22245  ( .IN0(\u_a23_mem/p_mem[112][2] ), .IN1(
        \u_a23_mem/p_mem[116][2] ), .SEL(m_address[2]), .F(\u_a23_mem/n22118 )
         );
  MUX \u_a23_mem/U22238  ( .IN0(\u_a23_mem/p_mem[120][2] ), .IN1(
        \u_a23_mem/p_mem[124][2] ), .SEL(m_address[2]), .F(\u_a23_mem/n22111 )
         );
  MUX \u_a23_mem/U22231  ( .IN0(\u_a23_mem/n22104 ), .IN1(\u_a23_mem/n22041 ), 
        .SEL(m_address[6]), .F(\u_a23_mem/N1845 ) );
  MUX \u_a23_mem/U22230  ( .IN0(\u_a23_mem/n22103 ), .IN1(\u_a23_mem/n22072 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n22104 ) );
  MUX \u_a23_mem/U22229  ( .IN0(\u_a23_mem/n22102 ), .IN1(\u_a23_mem/n22087 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n22103 ) );
  MUX \u_a23_mem/U22228  ( .IN0(\u_a23_mem/n22101 ), .IN1(\u_a23_mem/n22094 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22102 ) );
  MUX \u_a23_mem/U22227  ( .IN0(\u_a23_mem/p_mem[0][1] ), .IN1(
        \u_a23_mem/p_mem[4][1] ), .SEL(m_address[2]), .F(\u_a23_mem/n22101 )
         );
  MUX \u_a23_mem/U22220  ( .IN0(\u_a23_mem/p_mem[8][1] ), .IN1(
        \u_a23_mem/p_mem[12][1] ), .SEL(m_address[2]), .F(\u_a23_mem/n22094 )
         );
  MUX \u_a23_mem/U22213  ( .IN0(\u_a23_mem/n22086 ), .IN1(\u_a23_mem/n22079 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22087 ) );
  MUX \u_a23_mem/U22212  ( .IN0(\u_a23_mem/p_mem[16][1] ), .IN1(
        \u_a23_mem/p_mem[20][1] ), .SEL(m_address[2]), .F(\u_a23_mem/n22086 )
         );
  MUX \u_a23_mem/U22205  ( .IN0(\u_a23_mem/p_mem[24][1] ), .IN1(
        \u_a23_mem/p_mem[28][1] ), .SEL(m_address[2]), .F(\u_a23_mem/n22079 )
         );
  MUX \u_a23_mem/U22198  ( .IN0(\u_a23_mem/n22071 ), .IN1(\u_a23_mem/n22056 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n22072 ) );
  MUX \u_a23_mem/U22197  ( .IN0(\u_a23_mem/n22070 ), .IN1(\u_a23_mem/n22063 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22071 ) );
  MUX \u_a23_mem/U22196  ( .IN0(\u_a23_mem/p_mem[32][1] ), .IN1(
        \u_a23_mem/p_mem[36][1] ), .SEL(m_address[2]), .F(\u_a23_mem/n22070 )
         );
  MUX \u_a23_mem/U22189  ( .IN0(\u_a23_mem/p_mem[40][1] ), .IN1(
        \u_a23_mem/p_mem[44][1] ), .SEL(m_address[2]), .F(\u_a23_mem/n22063 )
         );
  MUX \u_a23_mem/U22182  ( .IN0(\u_a23_mem/n22055 ), .IN1(\u_a23_mem/n22048 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22056 ) );
  MUX \u_a23_mem/U22181  ( .IN0(\u_a23_mem/p_mem[48][1] ), .IN1(
        \u_a23_mem/p_mem[52][1] ), .SEL(m_address[2]), .F(\u_a23_mem/n22055 )
         );
  MUX \u_a23_mem/U22174  ( .IN0(\u_a23_mem/p_mem[56][1] ), .IN1(
        \u_a23_mem/p_mem[60][1] ), .SEL(m_address[2]), .F(\u_a23_mem/n22048 )
         );
  MUX \u_a23_mem/U22167  ( .IN0(\u_a23_mem/n22040 ), .IN1(\u_a23_mem/n22009 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n22041 ) );
  MUX \u_a23_mem/U22166  ( .IN0(\u_a23_mem/n22039 ), .IN1(\u_a23_mem/n22024 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n22040 ) );
  MUX \u_a23_mem/U22165  ( .IN0(\u_a23_mem/n22038 ), .IN1(\u_a23_mem/n22031 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22039 ) );
  MUX \u_a23_mem/U22164  ( .IN0(\u_a23_mem/p_mem[64][1] ), .IN1(
        \u_a23_mem/p_mem[68][1] ), .SEL(m_address[2]), .F(\u_a23_mem/n22038 )
         );
  MUX \u_a23_mem/U22157  ( .IN0(\u_a23_mem/p_mem[72][1] ), .IN1(
        \u_a23_mem/p_mem[76][1] ), .SEL(m_address[2]), .F(\u_a23_mem/n22031 )
         );
  MUX \u_a23_mem/U22150  ( .IN0(\u_a23_mem/n22023 ), .IN1(\u_a23_mem/n22016 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22024 ) );
  MUX \u_a23_mem/U22149  ( .IN0(\u_a23_mem/p_mem[80][1] ), .IN1(
        \u_a23_mem/p_mem[84][1] ), .SEL(m_address[2]), .F(\u_a23_mem/n22023 )
         );
  MUX \u_a23_mem/U22142  ( .IN0(\u_a23_mem/p_mem[88][1] ), .IN1(
        \u_a23_mem/p_mem[92][1] ), .SEL(m_address[2]), .F(\u_a23_mem/n22016 )
         );
  MUX \u_a23_mem/U22135  ( .IN0(\u_a23_mem/n22008 ), .IN1(\u_a23_mem/n21993 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n22009 ) );
  MUX \u_a23_mem/U22134  ( .IN0(\u_a23_mem/n22007 ), .IN1(\u_a23_mem/n22000 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n22008 ) );
  MUX \u_a23_mem/U22133  ( .IN0(\u_a23_mem/p_mem[96][1] ), .IN1(
        \u_a23_mem/p_mem[100][1] ), .SEL(m_address[2]), .F(\u_a23_mem/n22007 )
         );
  MUX \u_a23_mem/U22126  ( .IN0(\u_a23_mem/p_mem[104][1] ), .IN1(
        \u_a23_mem/p_mem[108][1] ), .SEL(m_address[2]), .F(\u_a23_mem/n22000 )
         );
  MUX \u_a23_mem/U22119  ( .IN0(\u_a23_mem/n21992 ), .IN1(\u_a23_mem/n21985 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21993 ) );
  MUX \u_a23_mem/U22118  ( .IN0(\u_a23_mem/p_mem[112][1] ), .IN1(
        \u_a23_mem/p_mem[116][1] ), .SEL(m_address[2]), .F(\u_a23_mem/n21992 )
         );
  MUX \u_a23_mem/U22111  ( .IN0(\u_a23_mem/p_mem[120][1] ), .IN1(
        \u_a23_mem/p_mem[124][1] ), .SEL(m_address[2]), .F(\u_a23_mem/n21985 )
         );
  MUX \u_a23_mem/U22104  ( .IN0(\u_a23_mem/n21978 ), .IN1(\u_a23_mem/n21915 ), 
        .SEL(m_address[6]), .F(\u_a23_mem/N1846 ) );
  MUX \u_a23_mem/U22103  ( .IN0(\u_a23_mem/n21977 ), .IN1(\u_a23_mem/n21946 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n21978 ) );
  MUX \u_a23_mem/U22102  ( .IN0(\u_a23_mem/n21976 ), .IN1(\u_a23_mem/n21961 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n21977 ) );
  MUX \u_a23_mem/U22101  ( .IN0(\u_a23_mem/n21975 ), .IN1(\u_a23_mem/n21968 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21976 ) );
  MUX \u_a23_mem/U22100  ( .IN0(\u_a23_mem/p_mem[0][0] ), .IN1(
        \u_a23_mem/p_mem[4][0] ), .SEL(m_address[2]), .F(\u_a23_mem/n21975 )
         );
  MUX \u_a23_mem/U22093  ( .IN0(\u_a23_mem/p_mem[8][0] ), .IN1(
        \u_a23_mem/p_mem[12][0] ), .SEL(m_address[2]), .F(\u_a23_mem/n21968 )
         );
  MUX \u_a23_mem/U22086  ( .IN0(\u_a23_mem/n21960 ), .IN1(\u_a23_mem/n21953 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21961 ) );
  MUX \u_a23_mem/U22085  ( .IN0(\u_a23_mem/p_mem[16][0] ), .IN1(
        \u_a23_mem/p_mem[20][0] ), .SEL(m_address[2]), .F(\u_a23_mem/n21960 )
         );
  MUX \u_a23_mem/U22078  ( .IN0(\u_a23_mem/p_mem[24][0] ), .IN1(
        \u_a23_mem/p_mem[28][0] ), .SEL(m_address[2]), .F(\u_a23_mem/n21953 )
         );
  MUX \u_a23_mem/U22071  ( .IN0(\u_a23_mem/n21945 ), .IN1(\u_a23_mem/n21930 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n21946 ) );
  MUX \u_a23_mem/U22070  ( .IN0(\u_a23_mem/n21944 ), .IN1(\u_a23_mem/n21937 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21945 ) );
  MUX \u_a23_mem/U22069  ( .IN0(\u_a23_mem/p_mem[32][0] ), .IN1(
        \u_a23_mem/p_mem[36][0] ), .SEL(m_address[2]), .F(\u_a23_mem/n21944 )
         );
  MUX \u_a23_mem/U22062  ( .IN0(\u_a23_mem/p_mem[40][0] ), .IN1(
        \u_a23_mem/p_mem[44][0] ), .SEL(m_address[2]), .F(\u_a23_mem/n21937 )
         );
  MUX \u_a23_mem/U22055  ( .IN0(\u_a23_mem/n21929 ), .IN1(\u_a23_mem/n21922 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21930 ) );
  MUX \u_a23_mem/U22054  ( .IN0(\u_a23_mem/p_mem[48][0] ), .IN1(
        \u_a23_mem/p_mem[52][0] ), .SEL(m_address[2]), .F(\u_a23_mem/n21929 )
         );
  MUX \u_a23_mem/U22047  ( .IN0(\u_a23_mem/p_mem[56][0] ), .IN1(
        \u_a23_mem/p_mem[60][0] ), .SEL(m_address[2]), .F(\u_a23_mem/n21922 )
         );
  MUX \u_a23_mem/U22040  ( .IN0(\u_a23_mem/n21914 ), .IN1(\u_a23_mem/n21883 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n21915 ) );
  MUX \u_a23_mem/U22039  ( .IN0(\u_a23_mem/n21913 ), .IN1(\u_a23_mem/n21898 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n21914 ) );
  MUX \u_a23_mem/U22038  ( .IN0(\u_a23_mem/n21912 ), .IN1(\u_a23_mem/n21905 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21913 ) );
  MUX \u_a23_mem/U22037  ( .IN0(\u_a23_mem/p_mem[64][0] ), .IN1(
        \u_a23_mem/p_mem[68][0] ), .SEL(m_address[2]), .F(\u_a23_mem/n21912 )
         );
  MUX \u_a23_mem/U22030  ( .IN0(\u_a23_mem/p_mem[72][0] ), .IN1(
        \u_a23_mem/p_mem[76][0] ), .SEL(m_address[2]), .F(\u_a23_mem/n21905 )
         );
  MUX \u_a23_mem/U22023  ( .IN0(\u_a23_mem/n21897 ), .IN1(\u_a23_mem/n21890 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21898 ) );
  MUX \u_a23_mem/U22022  ( .IN0(\u_a23_mem/p_mem[80][0] ), .IN1(
        \u_a23_mem/p_mem[84][0] ), .SEL(m_address[2]), .F(\u_a23_mem/n21897 )
         );
  MUX \u_a23_mem/U22015  ( .IN0(\u_a23_mem/p_mem[88][0] ), .IN1(
        \u_a23_mem/p_mem[92][0] ), .SEL(m_address[2]), .F(\u_a23_mem/n21890 )
         );
  MUX \u_a23_mem/U22008  ( .IN0(\u_a23_mem/n21882 ), .IN1(\u_a23_mem/n21867 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n21883 ) );
  MUX \u_a23_mem/U22007  ( .IN0(\u_a23_mem/n21881 ), .IN1(\u_a23_mem/n21874 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21882 ) );
  MUX \u_a23_mem/U22006  ( .IN0(\u_a23_mem/p_mem[96][0] ), .IN1(
        \u_a23_mem/p_mem[100][0] ), .SEL(m_address[2]), .F(\u_a23_mem/n21881 )
         );
  MUX \u_a23_mem/U21999  ( .IN0(\u_a23_mem/p_mem[104][0] ), .IN1(
        \u_a23_mem/p_mem[108][0] ), .SEL(m_address[2]), .F(\u_a23_mem/n21874 )
         );
  MUX \u_a23_mem/U21992  ( .IN0(\u_a23_mem/n21866 ), .IN1(\u_a23_mem/n21859 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21867 ) );
  MUX \u_a23_mem/U21991  ( .IN0(\u_a23_mem/p_mem[112][0] ), .IN1(
        \u_a23_mem/p_mem[116][0] ), .SEL(m_address[2]), .F(\u_a23_mem/n21866 )
         );
  MUX \u_a23_mem/U21984  ( .IN0(\u_a23_mem/p_mem[120][0] ), .IN1(
        \u_a23_mem/p_mem[124][0] ), .SEL(m_address[2]), .F(\u_a23_mem/n21859 )
         );
  MUX \u_a23_mem/U21839  ( .IN0(\u_a23_mem/n21730 ), .IN1(\u_a23_mem/n21727 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21731 ) );
  MUX \u_a23_mem/U21838  ( .IN0(\u_a23_mem/n21729 ), .IN1(\u_a23_mem/n21728 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21730 ) );
  MUX \u_a23_mem/U21837  ( .IN0(\u_a23_mem/g_mem[1][7] ), .IN1(
        \u_a23_mem/g_mem[17][7] ), .SEL(m_address[4]), .F(\u_a23_mem/n21729 )
         );
  MUX \u_a23_mem/U21836  ( .IN0(\u_a23_mem/g_mem[9][7] ), .IN1(
        \u_a23_mem/g_mem[25][7] ), .SEL(m_address[4]), .F(\u_a23_mem/n21728 )
         );
  MUX \u_a23_mem/U21835  ( .IN0(\u_a23_mem/n21726 ), .IN1(\u_a23_mem/n21725 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21727 ) );
  MUX \u_a23_mem/U21834  ( .IN0(\u_a23_mem/g_mem[5][7] ), .IN1(
        \u_a23_mem/g_mem[21][7] ), .SEL(m_address[4]), .F(\u_a23_mem/n21726 )
         );
  MUX \u_a23_mem/U21833  ( .IN0(\u_a23_mem/g_mem[13][7] ), .IN1(
        \u_a23_mem/g_mem[29][7] ), .SEL(m_address[4]), .F(\u_a23_mem/n21725 )
         );
  MUX \u_a23_mem/U21832  ( .IN0(\u_a23_mem/n21723 ), .IN1(\u_a23_mem/n21720 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21724 ) );
  MUX \u_a23_mem/U21831  ( .IN0(\u_a23_mem/n21722 ), .IN1(\u_a23_mem/n21721 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21723 ) );
  MUX \u_a23_mem/U21830  ( .IN0(\u_a23_mem/g_mem[3][7] ), .IN1(
        \u_a23_mem/g_mem[19][7] ), .SEL(m_address[4]), .F(\u_a23_mem/n21722 )
         );
  MUX \u_a23_mem/U21829  ( .IN0(\u_a23_mem/g_mem[11][7] ), .IN1(
        \u_a23_mem/g_mem[27][7] ), .SEL(m_address[4]), .F(\u_a23_mem/n21721 )
         );
  MUX \u_a23_mem/U21828  ( .IN0(\u_a23_mem/n21719 ), .IN1(\u_a23_mem/n21718 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21720 ) );
  MUX \u_a23_mem/U21827  ( .IN0(\u_a23_mem/g_mem[7][7] ), .IN1(
        \u_a23_mem/g_mem[23][7] ), .SEL(m_address[4]), .F(\u_a23_mem/n21719 )
         );
  MUX \u_a23_mem/U21826  ( .IN0(\u_a23_mem/g_mem[15][7] ), .IN1(
        \u_a23_mem/g_mem[31][7] ), .SEL(m_address[4]), .F(\u_a23_mem/n21718 )
         );
  MUX \u_a23_mem/U21824  ( .IN0(\u_a23_mem/n21715 ), .IN1(\u_a23_mem/n21712 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21716 ) );
  MUX \u_a23_mem/U21823  ( .IN0(\u_a23_mem/n21714 ), .IN1(\u_a23_mem/n21713 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21715 ) );
  MUX \u_a23_mem/U21822  ( .IN0(\u_a23_mem/g_mem[2][7] ), .IN1(
        \u_a23_mem/g_mem[18][7] ), .SEL(m_address[4]), .F(\u_a23_mem/n21714 )
         );
  MUX \u_a23_mem/U21821  ( .IN0(\u_a23_mem/g_mem[10][7] ), .IN1(
        \u_a23_mem/g_mem[26][7] ), .SEL(m_address[4]), .F(\u_a23_mem/n21713 )
         );
  MUX \u_a23_mem/U21820  ( .IN0(\u_a23_mem/n21711 ), .IN1(\u_a23_mem/n21710 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21712 ) );
  MUX \u_a23_mem/U21819  ( .IN0(\u_a23_mem/g_mem[6][7] ), .IN1(
        \u_a23_mem/g_mem[22][7] ), .SEL(m_address[4]), .F(\u_a23_mem/n21711 )
         );
  MUX \u_a23_mem/U21818  ( .IN0(\u_a23_mem/g_mem[14][7] ), .IN1(
        \u_a23_mem/g_mem[30][7] ), .SEL(m_address[4]), .F(\u_a23_mem/n21710 )
         );
  MUX \u_a23_mem/U21809  ( .IN0(\u_a23_mem/n21701 ), .IN1(\u_a23_mem/n21698 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21702 ) );
  MUX \u_a23_mem/U21808  ( .IN0(\u_a23_mem/n21700 ), .IN1(\u_a23_mem/n21699 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21701 ) );
  MUX \u_a23_mem/U21807  ( .IN0(\u_a23_mem/g_mem[1][6] ), .IN1(
        \u_a23_mem/g_mem[17][6] ), .SEL(m_address[4]), .F(\u_a23_mem/n21700 )
         );
  MUX \u_a23_mem/U21806  ( .IN0(\u_a23_mem/g_mem[9][6] ), .IN1(
        \u_a23_mem/g_mem[25][6] ), .SEL(m_address[4]), .F(\u_a23_mem/n21699 )
         );
  MUX \u_a23_mem/U21805  ( .IN0(\u_a23_mem/n21697 ), .IN1(\u_a23_mem/n21696 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21698 ) );
  MUX \u_a23_mem/U21804  ( .IN0(\u_a23_mem/g_mem[5][6] ), .IN1(
        \u_a23_mem/g_mem[21][6] ), .SEL(m_address[4]), .F(\u_a23_mem/n21697 )
         );
  MUX \u_a23_mem/U21803  ( .IN0(\u_a23_mem/g_mem[13][6] ), .IN1(
        \u_a23_mem/g_mem[29][6] ), .SEL(m_address[4]), .F(\u_a23_mem/n21696 )
         );
  MUX \u_a23_mem/U21802  ( .IN0(\u_a23_mem/n21694 ), .IN1(\u_a23_mem/n21691 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21695 ) );
  MUX \u_a23_mem/U21801  ( .IN0(\u_a23_mem/n21693 ), .IN1(\u_a23_mem/n21692 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21694 ) );
  MUX \u_a23_mem/U21800  ( .IN0(\u_a23_mem/g_mem[3][6] ), .IN1(
        \u_a23_mem/g_mem[19][6] ), .SEL(m_address[4]), .F(\u_a23_mem/n21693 )
         );
  MUX \u_a23_mem/U21799  ( .IN0(\u_a23_mem/g_mem[11][6] ), .IN1(
        \u_a23_mem/g_mem[27][6] ), .SEL(m_address[4]), .F(\u_a23_mem/n21692 )
         );
  MUX \u_a23_mem/U21798  ( .IN0(\u_a23_mem/n21690 ), .IN1(\u_a23_mem/n21689 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21691 ) );
  MUX \u_a23_mem/U21797  ( .IN0(\u_a23_mem/g_mem[7][6] ), .IN1(
        \u_a23_mem/g_mem[23][6] ), .SEL(m_address[4]), .F(\u_a23_mem/n21690 )
         );
  MUX \u_a23_mem/U21796  ( .IN0(\u_a23_mem/g_mem[15][6] ), .IN1(
        \u_a23_mem/g_mem[31][6] ), .SEL(m_address[4]), .F(\u_a23_mem/n21689 )
         );
  MUX \u_a23_mem/U21794  ( .IN0(\u_a23_mem/n21686 ), .IN1(\u_a23_mem/n21683 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21687 ) );
  MUX \u_a23_mem/U21793  ( .IN0(\u_a23_mem/n21685 ), .IN1(\u_a23_mem/n21684 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21686 ) );
  MUX \u_a23_mem/U21792  ( .IN0(\u_a23_mem/g_mem[2][6] ), .IN1(
        \u_a23_mem/g_mem[18][6] ), .SEL(m_address[4]), .F(\u_a23_mem/n21685 )
         );
  MUX \u_a23_mem/U21791  ( .IN0(\u_a23_mem/g_mem[10][6] ), .IN1(
        \u_a23_mem/g_mem[26][6] ), .SEL(m_address[4]), .F(\u_a23_mem/n21684 )
         );
  MUX \u_a23_mem/U21790  ( .IN0(\u_a23_mem/n21682 ), .IN1(\u_a23_mem/n21681 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21683 ) );
  MUX \u_a23_mem/U21789  ( .IN0(\u_a23_mem/g_mem[6][6] ), .IN1(
        \u_a23_mem/g_mem[22][6] ), .SEL(m_address[4]), .F(\u_a23_mem/n21682 )
         );
  MUX \u_a23_mem/U21788  ( .IN0(\u_a23_mem/g_mem[14][6] ), .IN1(
        \u_a23_mem/g_mem[30][6] ), .SEL(m_address[4]), .F(\u_a23_mem/n21681 )
         );
  MUX \u_a23_mem/U21779  ( .IN0(\u_a23_mem/n21672 ), .IN1(\u_a23_mem/n21669 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21673 ) );
  MUX \u_a23_mem/U21778  ( .IN0(\u_a23_mem/n21671 ), .IN1(\u_a23_mem/n21670 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21672 ) );
  MUX \u_a23_mem/U21777  ( .IN0(\u_a23_mem/g_mem[1][5] ), .IN1(
        \u_a23_mem/g_mem[17][5] ), .SEL(m_address[4]), .F(\u_a23_mem/n21671 )
         );
  MUX \u_a23_mem/U21776  ( .IN0(\u_a23_mem/g_mem[9][5] ), .IN1(
        \u_a23_mem/g_mem[25][5] ), .SEL(m_address[4]), .F(\u_a23_mem/n21670 )
         );
  MUX \u_a23_mem/U21775  ( .IN0(\u_a23_mem/n21668 ), .IN1(\u_a23_mem/n21667 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21669 ) );
  MUX \u_a23_mem/U21774  ( .IN0(\u_a23_mem/g_mem[5][5] ), .IN1(
        \u_a23_mem/g_mem[21][5] ), .SEL(m_address[4]), .F(\u_a23_mem/n21668 )
         );
  MUX \u_a23_mem/U21773  ( .IN0(\u_a23_mem/g_mem[13][5] ), .IN1(
        \u_a23_mem/g_mem[29][5] ), .SEL(m_address[4]), .F(\u_a23_mem/n21667 )
         );
  MUX \u_a23_mem/U21772  ( .IN0(\u_a23_mem/n21665 ), .IN1(\u_a23_mem/n21662 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21666 ) );
  MUX \u_a23_mem/U21771  ( .IN0(\u_a23_mem/n21664 ), .IN1(\u_a23_mem/n21663 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21665 ) );
  MUX \u_a23_mem/U21770  ( .IN0(\u_a23_mem/g_mem[3][5] ), .IN1(
        \u_a23_mem/g_mem[19][5] ), .SEL(m_address[4]), .F(\u_a23_mem/n21664 )
         );
  MUX \u_a23_mem/U21769  ( .IN0(\u_a23_mem/g_mem[11][5] ), .IN1(
        \u_a23_mem/g_mem[27][5] ), .SEL(m_address[4]), .F(\u_a23_mem/n21663 )
         );
  MUX \u_a23_mem/U21768  ( .IN0(\u_a23_mem/n21661 ), .IN1(\u_a23_mem/n21660 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21662 ) );
  MUX \u_a23_mem/U21767  ( .IN0(\u_a23_mem/g_mem[7][5] ), .IN1(
        \u_a23_mem/g_mem[23][5] ), .SEL(m_address[4]), .F(\u_a23_mem/n21661 )
         );
  MUX \u_a23_mem/U21766  ( .IN0(\u_a23_mem/g_mem[15][5] ), .IN1(
        \u_a23_mem/g_mem[31][5] ), .SEL(m_address[4]), .F(\u_a23_mem/n21660 )
         );
  MUX \u_a23_mem/U21764  ( .IN0(\u_a23_mem/n21657 ), .IN1(\u_a23_mem/n21654 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21658 ) );
  MUX \u_a23_mem/U21763  ( .IN0(\u_a23_mem/n21656 ), .IN1(\u_a23_mem/n21655 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21657 ) );
  MUX \u_a23_mem/U21762  ( .IN0(\u_a23_mem/g_mem[2][5] ), .IN1(
        \u_a23_mem/g_mem[18][5] ), .SEL(m_address[4]), .F(\u_a23_mem/n21656 )
         );
  MUX \u_a23_mem/U21761  ( .IN0(\u_a23_mem/g_mem[10][5] ), .IN1(
        \u_a23_mem/g_mem[26][5] ), .SEL(m_address[4]), .F(\u_a23_mem/n21655 )
         );
  MUX \u_a23_mem/U21760  ( .IN0(\u_a23_mem/n21653 ), .IN1(\u_a23_mem/n21652 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21654 ) );
  MUX \u_a23_mem/U21759  ( .IN0(\u_a23_mem/g_mem[6][5] ), .IN1(
        \u_a23_mem/g_mem[22][5] ), .SEL(m_address[4]), .F(\u_a23_mem/n21653 )
         );
  MUX \u_a23_mem/U21758  ( .IN0(\u_a23_mem/g_mem[14][5] ), .IN1(
        \u_a23_mem/g_mem[30][5] ), .SEL(m_address[4]), .F(\u_a23_mem/n21652 )
         );
  MUX \u_a23_mem/U21749  ( .IN0(\u_a23_mem/n21643 ), .IN1(\u_a23_mem/n21640 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21644 ) );
  MUX \u_a23_mem/U21748  ( .IN0(\u_a23_mem/n21642 ), .IN1(\u_a23_mem/n21641 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21643 ) );
  MUX \u_a23_mem/U21747  ( .IN0(\u_a23_mem/g_mem[1][4] ), .IN1(
        \u_a23_mem/g_mem[17][4] ), .SEL(m_address[4]), .F(\u_a23_mem/n21642 )
         );
  MUX \u_a23_mem/U21746  ( .IN0(\u_a23_mem/g_mem[9][4] ), .IN1(
        \u_a23_mem/g_mem[25][4] ), .SEL(m_address[4]), .F(\u_a23_mem/n21641 )
         );
  MUX \u_a23_mem/U21745  ( .IN0(\u_a23_mem/n21639 ), .IN1(\u_a23_mem/n21638 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21640 ) );
  MUX \u_a23_mem/U21744  ( .IN0(\u_a23_mem/g_mem[5][4] ), .IN1(
        \u_a23_mem/g_mem[21][4] ), .SEL(m_address[4]), .F(\u_a23_mem/n21639 )
         );
  MUX \u_a23_mem/U21743  ( .IN0(\u_a23_mem/g_mem[13][4] ), .IN1(
        \u_a23_mem/g_mem[29][4] ), .SEL(m_address[4]), .F(\u_a23_mem/n21638 )
         );
  MUX \u_a23_mem/U21742  ( .IN0(\u_a23_mem/n21636 ), .IN1(\u_a23_mem/n21633 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21637 ) );
  MUX \u_a23_mem/U21741  ( .IN0(\u_a23_mem/n21635 ), .IN1(\u_a23_mem/n21634 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21636 ) );
  MUX \u_a23_mem/U21740  ( .IN0(\u_a23_mem/g_mem[3][4] ), .IN1(
        \u_a23_mem/g_mem[19][4] ), .SEL(m_address[4]), .F(\u_a23_mem/n21635 )
         );
  MUX \u_a23_mem/U21739  ( .IN0(\u_a23_mem/g_mem[11][4] ), .IN1(
        \u_a23_mem/g_mem[27][4] ), .SEL(m_address[4]), .F(\u_a23_mem/n21634 )
         );
  MUX \u_a23_mem/U21738  ( .IN0(\u_a23_mem/n21632 ), .IN1(\u_a23_mem/n21631 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21633 ) );
  MUX \u_a23_mem/U21737  ( .IN0(\u_a23_mem/g_mem[7][4] ), .IN1(
        \u_a23_mem/g_mem[23][4] ), .SEL(m_address[4]), .F(\u_a23_mem/n21632 )
         );
  MUX \u_a23_mem/U21736  ( .IN0(\u_a23_mem/g_mem[15][4] ), .IN1(
        \u_a23_mem/g_mem[31][4] ), .SEL(m_address[4]), .F(\u_a23_mem/n21631 )
         );
  MUX \u_a23_mem/U21734  ( .IN0(\u_a23_mem/n21628 ), .IN1(\u_a23_mem/n21625 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21629 ) );
  MUX \u_a23_mem/U21733  ( .IN0(\u_a23_mem/n21627 ), .IN1(\u_a23_mem/n21626 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21628 ) );
  MUX \u_a23_mem/U21732  ( .IN0(\u_a23_mem/g_mem[2][4] ), .IN1(
        \u_a23_mem/g_mem[18][4] ), .SEL(m_address[4]), .F(\u_a23_mem/n21627 )
         );
  MUX \u_a23_mem/U21731  ( .IN0(\u_a23_mem/g_mem[10][4] ), .IN1(
        \u_a23_mem/g_mem[26][4] ), .SEL(m_address[4]), .F(\u_a23_mem/n21626 )
         );
  MUX \u_a23_mem/U21730  ( .IN0(\u_a23_mem/n21624 ), .IN1(\u_a23_mem/n21623 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21625 ) );
  MUX \u_a23_mem/U21729  ( .IN0(\u_a23_mem/g_mem[6][4] ), .IN1(
        \u_a23_mem/g_mem[22][4] ), .SEL(m_address[4]), .F(\u_a23_mem/n21624 )
         );
  MUX \u_a23_mem/U21728  ( .IN0(\u_a23_mem/g_mem[14][4] ), .IN1(
        \u_a23_mem/g_mem[30][4] ), .SEL(m_address[4]), .F(\u_a23_mem/n21623 )
         );
  MUX \u_a23_mem/U21719  ( .IN0(\u_a23_mem/n21614 ), .IN1(\u_a23_mem/n21611 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21615 ) );
  MUX \u_a23_mem/U21718  ( .IN0(\u_a23_mem/n21613 ), .IN1(\u_a23_mem/n21612 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21614 ) );
  MUX \u_a23_mem/U21717  ( .IN0(\u_a23_mem/g_mem[1][3] ), .IN1(
        \u_a23_mem/g_mem[17][3] ), .SEL(m_address[4]), .F(\u_a23_mem/n21613 )
         );
  MUX \u_a23_mem/U21716  ( .IN0(\u_a23_mem/g_mem[9][3] ), .IN1(
        \u_a23_mem/g_mem[25][3] ), .SEL(m_address[4]), .F(\u_a23_mem/n21612 )
         );
  MUX \u_a23_mem/U21715  ( .IN0(\u_a23_mem/n21610 ), .IN1(\u_a23_mem/n21609 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21611 ) );
  MUX \u_a23_mem/U21714  ( .IN0(\u_a23_mem/g_mem[5][3] ), .IN1(
        \u_a23_mem/g_mem[21][3] ), .SEL(m_address[4]), .F(\u_a23_mem/n21610 )
         );
  MUX \u_a23_mem/U21713  ( .IN0(\u_a23_mem/g_mem[13][3] ), .IN1(
        \u_a23_mem/g_mem[29][3] ), .SEL(m_address[4]), .F(\u_a23_mem/n21609 )
         );
  MUX \u_a23_mem/U21712  ( .IN0(\u_a23_mem/n21607 ), .IN1(\u_a23_mem/n21604 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21608 ) );
  MUX \u_a23_mem/U21711  ( .IN0(\u_a23_mem/n21606 ), .IN1(\u_a23_mem/n21605 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21607 ) );
  MUX \u_a23_mem/U21710  ( .IN0(\u_a23_mem/g_mem[3][3] ), .IN1(
        \u_a23_mem/g_mem[19][3] ), .SEL(m_address[4]), .F(\u_a23_mem/n21606 )
         );
  MUX \u_a23_mem/U21709  ( .IN0(\u_a23_mem/g_mem[11][3] ), .IN1(
        \u_a23_mem/g_mem[27][3] ), .SEL(m_address[4]), .F(\u_a23_mem/n21605 )
         );
  MUX \u_a23_mem/U21708  ( .IN0(\u_a23_mem/n21603 ), .IN1(\u_a23_mem/n21602 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21604 ) );
  MUX \u_a23_mem/U21707  ( .IN0(\u_a23_mem/g_mem[7][3] ), .IN1(
        \u_a23_mem/g_mem[23][3] ), .SEL(m_address[4]), .F(\u_a23_mem/n21603 )
         );
  MUX \u_a23_mem/U21706  ( .IN0(\u_a23_mem/g_mem[15][3] ), .IN1(
        \u_a23_mem/g_mem[31][3] ), .SEL(m_address[4]), .F(\u_a23_mem/n21602 )
         );
  MUX \u_a23_mem/U21704  ( .IN0(\u_a23_mem/n21599 ), .IN1(\u_a23_mem/n21596 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21600 ) );
  MUX \u_a23_mem/U21703  ( .IN0(\u_a23_mem/n21598 ), .IN1(\u_a23_mem/n21597 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21599 ) );
  MUX \u_a23_mem/U21702  ( .IN0(\u_a23_mem/g_mem[2][3] ), .IN1(
        \u_a23_mem/g_mem[18][3] ), .SEL(m_address[4]), .F(\u_a23_mem/n21598 )
         );
  MUX \u_a23_mem/U21701  ( .IN0(\u_a23_mem/g_mem[10][3] ), .IN1(
        \u_a23_mem/g_mem[26][3] ), .SEL(m_address[4]), .F(\u_a23_mem/n21597 )
         );
  MUX \u_a23_mem/U21700  ( .IN0(\u_a23_mem/n21595 ), .IN1(\u_a23_mem/n21594 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21596 ) );
  MUX \u_a23_mem/U21699  ( .IN0(\u_a23_mem/g_mem[6][3] ), .IN1(
        \u_a23_mem/g_mem[22][3] ), .SEL(m_address[4]), .F(\u_a23_mem/n21595 )
         );
  MUX \u_a23_mem/U21698  ( .IN0(\u_a23_mem/g_mem[14][3] ), .IN1(
        \u_a23_mem/g_mem[30][3] ), .SEL(m_address[4]), .F(\u_a23_mem/n21594 )
         );
  MUX \u_a23_mem/U21689  ( .IN0(\u_a23_mem/n21585 ), .IN1(\u_a23_mem/n21582 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21586 ) );
  MUX \u_a23_mem/U21688  ( .IN0(\u_a23_mem/n21584 ), .IN1(\u_a23_mem/n21583 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21585 ) );
  MUX \u_a23_mem/U21687  ( .IN0(\u_a23_mem/g_mem[1][2] ), .IN1(
        \u_a23_mem/g_mem[17][2] ), .SEL(m_address[4]), .F(\u_a23_mem/n21584 )
         );
  MUX \u_a23_mem/U21686  ( .IN0(\u_a23_mem/g_mem[9][2] ), .IN1(
        \u_a23_mem/g_mem[25][2] ), .SEL(m_address[4]), .F(\u_a23_mem/n21583 )
         );
  MUX \u_a23_mem/U21685  ( .IN0(\u_a23_mem/n21581 ), .IN1(\u_a23_mem/n21580 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21582 ) );
  MUX \u_a23_mem/U21684  ( .IN0(\u_a23_mem/g_mem[5][2] ), .IN1(
        \u_a23_mem/g_mem[21][2] ), .SEL(m_address[4]), .F(\u_a23_mem/n21581 )
         );
  MUX \u_a23_mem/U21683  ( .IN0(\u_a23_mem/g_mem[13][2] ), .IN1(
        \u_a23_mem/g_mem[29][2] ), .SEL(m_address[4]), .F(\u_a23_mem/n21580 )
         );
  MUX \u_a23_mem/U21682  ( .IN0(\u_a23_mem/n21578 ), .IN1(\u_a23_mem/n21575 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21579 ) );
  MUX \u_a23_mem/U21681  ( .IN0(\u_a23_mem/n21577 ), .IN1(\u_a23_mem/n21576 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21578 ) );
  MUX \u_a23_mem/U21680  ( .IN0(\u_a23_mem/g_mem[3][2] ), .IN1(
        \u_a23_mem/g_mem[19][2] ), .SEL(m_address[4]), .F(\u_a23_mem/n21577 )
         );
  MUX \u_a23_mem/U21679  ( .IN0(\u_a23_mem/g_mem[11][2] ), .IN1(
        \u_a23_mem/g_mem[27][2] ), .SEL(m_address[4]), .F(\u_a23_mem/n21576 )
         );
  MUX \u_a23_mem/U21678  ( .IN0(\u_a23_mem/n21574 ), .IN1(\u_a23_mem/n21573 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21575 ) );
  MUX \u_a23_mem/U21677  ( .IN0(\u_a23_mem/g_mem[7][2] ), .IN1(
        \u_a23_mem/g_mem[23][2] ), .SEL(m_address[4]), .F(\u_a23_mem/n21574 )
         );
  MUX \u_a23_mem/U21676  ( .IN0(\u_a23_mem/g_mem[15][2] ), .IN1(
        \u_a23_mem/g_mem[31][2] ), .SEL(m_address[4]), .F(\u_a23_mem/n21573 )
         );
  MUX \u_a23_mem/U21674  ( .IN0(\u_a23_mem/n21570 ), .IN1(\u_a23_mem/n21567 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21571 ) );
  MUX \u_a23_mem/U21673  ( .IN0(\u_a23_mem/n21569 ), .IN1(\u_a23_mem/n21568 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21570 ) );
  MUX \u_a23_mem/U21672  ( .IN0(\u_a23_mem/g_mem[2][2] ), .IN1(
        \u_a23_mem/g_mem[18][2] ), .SEL(m_address[4]), .F(\u_a23_mem/n21569 )
         );
  MUX \u_a23_mem/U21671  ( .IN0(\u_a23_mem/g_mem[10][2] ), .IN1(
        \u_a23_mem/g_mem[26][2] ), .SEL(m_address[4]), .F(\u_a23_mem/n21568 )
         );
  MUX \u_a23_mem/U21670  ( .IN0(\u_a23_mem/n21566 ), .IN1(\u_a23_mem/n21565 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21567 ) );
  MUX \u_a23_mem/U21669  ( .IN0(\u_a23_mem/g_mem[6][2] ), .IN1(
        \u_a23_mem/g_mem[22][2] ), .SEL(m_address[4]), .F(\u_a23_mem/n21566 )
         );
  MUX \u_a23_mem/U21668  ( .IN0(\u_a23_mem/g_mem[14][2] ), .IN1(
        \u_a23_mem/g_mem[30][2] ), .SEL(m_address[4]), .F(\u_a23_mem/n21565 )
         );
  MUX \u_a23_mem/U21659  ( .IN0(\u_a23_mem/n21556 ), .IN1(\u_a23_mem/n21553 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21557 ) );
  MUX \u_a23_mem/U21658  ( .IN0(\u_a23_mem/n21555 ), .IN1(\u_a23_mem/n21554 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21556 ) );
  MUX \u_a23_mem/U21657  ( .IN0(\u_a23_mem/g_mem[1][1] ), .IN1(
        \u_a23_mem/g_mem[17][1] ), .SEL(m_address[4]), .F(\u_a23_mem/n21555 )
         );
  MUX \u_a23_mem/U21656  ( .IN0(\u_a23_mem/g_mem[9][1] ), .IN1(
        \u_a23_mem/g_mem[25][1] ), .SEL(m_address[4]), .F(\u_a23_mem/n21554 )
         );
  MUX \u_a23_mem/U21655  ( .IN0(\u_a23_mem/n21552 ), .IN1(\u_a23_mem/n21551 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21553 ) );
  MUX \u_a23_mem/U21654  ( .IN0(\u_a23_mem/g_mem[5][1] ), .IN1(
        \u_a23_mem/g_mem[21][1] ), .SEL(m_address[4]), .F(\u_a23_mem/n21552 )
         );
  MUX \u_a23_mem/U21653  ( .IN0(\u_a23_mem/g_mem[13][1] ), .IN1(
        \u_a23_mem/g_mem[29][1] ), .SEL(m_address[4]), .F(\u_a23_mem/n21551 )
         );
  MUX \u_a23_mem/U21652  ( .IN0(\u_a23_mem/n21549 ), .IN1(\u_a23_mem/n21546 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21550 ) );
  MUX \u_a23_mem/U21651  ( .IN0(\u_a23_mem/n21548 ), .IN1(\u_a23_mem/n21547 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21549 ) );
  MUX \u_a23_mem/U21650  ( .IN0(\u_a23_mem/g_mem[3][1] ), .IN1(
        \u_a23_mem/g_mem[19][1] ), .SEL(m_address[4]), .F(\u_a23_mem/n21548 )
         );
  MUX \u_a23_mem/U21649  ( .IN0(\u_a23_mem/g_mem[11][1] ), .IN1(
        \u_a23_mem/g_mem[27][1] ), .SEL(m_address[4]), .F(\u_a23_mem/n21547 )
         );
  MUX \u_a23_mem/U21648  ( .IN0(\u_a23_mem/n21545 ), .IN1(\u_a23_mem/n21544 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21546 ) );
  MUX \u_a23_mem/U21647  ( .IN0(\u_a23_mem/g_mem[7][1] ), .IN1(
        \u_a23_mem/g_mem[23][1] ), .SEL(m_address[4]), .F(\u_a23_mem/n21545 )
         );
  MUX \u_a23_mem/U21646  ( .IN0(\u_a23_mem/g_mem[15][1] ), .IN1(
        \u_a23_mem/g_mem[31][1] ), .SEL(m_address[4]), .F(\u_a23_mem/n21544 )
         );
  MUX \u_a23_mem/U21644  ( .IN0(\u_a23_mem/n21541 ), .IN1(\u_a23_mem/n21538 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21542 ) );
  MUX \u_a23_mem/U21643  ( .IN0(\u_a23_mem/n21540 ), .IN1(\u_a23_mem/n21539 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21541 ) );
  MUX \u_a23_mem/U21642  ( .IN0(\u_a23_mem/g_mem[2][1] ), .IN1(
        \u_a23_mem/g_mem[18][1] ), .SEL(m_address[4]), .F(\u_a23_mem/n21540 )
         );
  MUX \u_a23_mem/U21641  ( .IN0(\u_a23_mem/g_mem[10][1] ), .IN1(
        \u_a23_mem/g_mem[26][1] ), .SEL(m_address[4]), .F(\u_a23_mem/n21539 )
         );
  MUX \u_a23_mem/U21640  ( .IN0(\u_a23_mem/n21537 ), .IN1(\u_a23_mem/n21536 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21538 ) );
  MUX \u_a23_mem/U21639  ( .IN0(\u_a23_mem/g_mem[6][1] ), .IN1(
        \u_a23_mem/g_mem[22][1] ), .SEL(m_address[4]), .F(\u_a23_mem/n21537 )
         );
  MUX \u_a23_mem/U21638  ( .IN0(\u_a23_mem/g_mem[14][1] ), .IN1(
        \u_a23_mem/g_mem[30][1] ), .SEL(m_address[4]), .F(\u_a23_mem/n21536 )
         );
  MUX \u_a23_mem/U21629  ( .IN0(\u_a23_mem/n21527 ), .IN1(\u_a23_mem/n21524 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21528 ) );
  MUX \u_a23_mem/U21628  ( .IN0(\u_a23_mem/n21526 ), .IN1(\u_a23_mem/n21525 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21527 ) );
  MUX \u_a23_mem/U21627  ( .IN0(\u_a23_mem/g_mem[1][0] ), .IN1(
        \u_a23_mem/g_mem[17][0] ), .SEL(m_address[4]), .F(\u_a23_mem/n21526 )
         );
  MUX \u_a23_mem/U21626  ( .IN0(\u_a23_mem/g_mem[9][0] ), .IN1(
        \u_a23_mem/g_mem[25][0] ), .SEL(m_address[4]), .F(\u_a23_mem/n21525 )
         );
  MUX \u_a23_mem/U21625  ( .IN0(\u_a23_mem/n21523 ), .IN1(\u_a23_mem/n21522 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21524 ) );
  MUX \u_a23_mem/U21624  ( .IN0(\u_a23_mem/g_mem[5][0] ), .IN1(
        \u_a23_mem/g_mem[21][0] ), .SEL(m_address[4]), .F(\u_a23_mem/n21523 )
         );
  MUX \u_a23_mem/U21623  ( .IN0(\u_a23_mem/g_mem[13][0] ), .IN1(
        \u_a23_mem/g_mem[29][0] ), .SEL(m_address[4]), .F(\u_a23_mem/n21522 )
         );
  MUX \u_a23_mem/U21622  ( .IN0(\u_a23_mem/n21520 ), .IN1(\u_a23_mem/n21517 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21521 ) );
  MUX \u_a23_mem/U21621  ( .IN0(\u_a23_mem/n21519 ), .IN1(\u_a23_mem/n21518 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21520 ) );
  MUX \u_a23_mem/U21620  ( .IN0(\u_a23_mem/g_mem[3][0] ), .IN1(
        \u_a23_mem/g_mem[19][0] ), .SEL(m_address[4]), .F(\u_a23_mem/n21519 )
         );
  MUX \u_a23_mem/U21619  ( .IN0(\u_a23_mem/g_mem[11][0] ), .IN1(
        \u_a23_mem/g_mem[27][0] ), .SEL(m_address[4]), .F(\u_a23_mem/n21518 )
         );
  MUX \u_a23_mem/U21618  ( .IN0(\u_a23_mem/n21516 ), .IN1(\u_a23_mem/n21515 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21517 ) );
  MUX \u_a23_mem/U21617  ( .IN0(\u_a23_mem/g_mem[7][0] ), .IN1(
        \u_a23_mem/g_mem[23][0] ), .SEL(m_address[4]), .F(\u_a23_mem/n21516 )
         );
  MUX \u_a23_mem/U21616  ( .IN0(\u_a23_mem/g_mem[15][0] ), .IN1(
        \u_a23_mem/g_mem[31][0] ), .SEL(m_address[4]), .F(\u_a23_mem/n21515 )
         );
  MUX \u_a23_mem/U21614  ( .IN0(\u_a23_mem/n21512 ), .IN1(\u_a23_mem/n21509 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21513 ) );
  MUX \u_a23_mem/U21613  ( .IN0(\u_a23_mem/n21511 ), .IN1(\u_a23_mem/n21510 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21512 ) );
  MUX \u_a23_mem/U21612  ( .IN0(\u_a23_mem/g_mem[2][0] ), .IN1(
        \u_a23_mem/g_mem[18][0] ), .SEL(m_address[4]), .F(\u_a23_mem/n21511 )
         );
  MUX \u_a23_mem/U21611  ( .IN0(\u_a23_mem/g_mem[10][0] ), .IN1(
        \u_a23_mem/g_mem[26][0] ), .SEL(m_address[4]), .F(\u_a23_mem/n21510 )
         );
  MUX \u_a23_mem/U21610  ( .IN0(\u_a23_mem/n21508 ), .IN1(\u_a23_mem/n21507 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21509 ) );
  MUX \u_a23_mem/U21609  ( .IN0(\u_a23_mem/g_mem[6][0] ), .IN1(
        \u_a23_mem/g_mem[22][0] ), .SEL(m_address[4]), .F(\u_a23_mem/n21508 )
         );
  MUX \u_a23_mem/U21608  ( .IN0(\u_a23_mem/g_mem[14][0] ), .IN1(
        \u_a23_mem/g_mem[30][0] ), .SEL(m_address[4]), .F(\u_a23_mem/n21507 )
         );
  MUX \u_a23_mem/U21559  ( .IN0(\u_a23_mem/n21474 ), .IN1(\u_a23_mem/n21471 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21475 ) );
  MUX \u_a23_mem/U21558  ( .IN0(\u_a23_mem/n21473 ), .IN1(\u_a23_mem/n21472 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21474 ) );
  MUX \u_a23_mem/U21557  ( .IN0(\u_a23_mem/e_mem[1][7] ), .IN1(
        \u_a23_mem/e_mem[17][7] ), .SEL(m_address[4]), .F(\u_a23_mem/n21473 )
         );
  MUX \u_a23_mem/U21556  ( .IN0(\u_a23_mem/e_mem[9][7] ), .IN1(
        \u_a23_mem/e_mem[25][7] ), .SEL(m_address[4]), .F(\u_a23_mem/n21472 )
         );
  MUX \u_a23_mem/U21555  ( .IN0(\u_a23_mem/n21470 ), .IN1(\u_a23_mem/n21469 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21471 ) );
  MUX \u_a23_mem/U21554  ( .IN0(\u_a23_mem/e_mem[5][7] ), .IN1(
        \u_a23_mem/e_mem[21][7] ), .SEL(m_address[4]), .F(\u_a23_mem/n21470 )
         );
  MUX \u_a23_mem/U21553  ( .IN0(\u_a23_mem/e_mem[13][7] ), .IN1(
        \u_a23_mem/e_mem[29][7] ), .SEL(m_address[4]), .F(\u_a23_mem/n21469 )
         );
  MUX \u_a23_mem/U21552  ( .IN0(\u_a23_mem/n21467 ), .IN1(\u_a23_mem/n21464 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21468 ) );
  MUX \u_a23_mem/U21551  ( .IN0(\u_a23_mem/n21466 ), .IN1(\u_a23_mem/n21465 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21467 ) );
  MUX \u_a23_mem/U21550  ( .IN0(\u_a23_mem/e_mem[3][7] ), .IN1(
        \u_a23_mem/e_mem[19][7] ), .SEL(m_address[4]), .F(\u_a23_mem/n21466 )
         );
  MUX \u_a23_mem/U21549  ( .IN0(\u_a23_mem/e_mem[11][7] ), .IN1(
        \u_a23_mem/e_mem[27][7] ), .SEL(m_address[4]), .F(\u_a23_mem/n21465 )
         );
  MUX \u_a23_mem/U21548  ( .IN0(\u_a23_mem/n21463 ), .IN1(\u_a23_mem/n21462 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21464 ) );
  MUX \u_a23_mem/U21547  ( .IN0(\u_a23_mem/e_mem[7][7] ), .IN1(
        \u_a23_mem/e_mem[23][7] ), .SEL(m_address[4]), .F(\u_a23_mem/n21463 )
         );
  MUX \u_a23_mem/U21546  ( .IN0(\u_a23_mem/e_mem[15][7] ), .IN1(
        \u_a23_mem/e_mem[31][7] ), .SEL(m_address[4]), .F(\u_a23_mem/n21462 )
         );
  MUX \u_a23_mem/U21544  ( .IN0(\u_a23_mem/n21459 ), .IN1(\u_a23_mem/n21456 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21460 ) );
  MUX \u_a23_mem/U21543  ( .IN0(\u_a23_mem/n21458 ), .IN1(\u_a23_mem/n21457 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21459 ) );
  MUX \u_a23_mem/U21542  ( .IN0(\u_a23_mem/e_mem[2][7] ), .IN1(
        \u_a23_mem/e_mem[18][7] ), .SEL(m_address[4]), .F(\u_a23_mem/n21458 )
         );
  MUX \u_a23_mem/U21541  ( .IN0(\u_a23_mem/e_mem[10][7] ), .IN1(
        \u_a23_mem/e_mem[26][7] ), .SEL(m_address[4]), .F(\u_a23_mem/n21457 )
         );
  MUX \u_a23_mem/U21540  ( .IN0(\u_a23_mem/n21455 ), .IN1(\u_a23_mem/n21454 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21456 ) );
  MUX \u_a23_mem/U21539  ( .IN0(\u_a23_mem/e_mem[6][7] ), .IN1(
        \u_a23_mem/e_mem[22][7] ), .SEL(m_address[4]), .F(\u_a23_mem/n21455 )
         );
  MUX \u_a23_mem/U21538  ( .IN0(\u_a23_mem/e_mem[14][7] ), .IN1(
        \u_a23_mem/e_mem[30][7] ), .SEL(m_address[4]), .F(\u_a23_mem/n21454 )
         );
  MUX \u_a23_mem/U21529  ( .IN0(\u_a23_mem/n21445 ), .IN1(\u_a23_mem/n21442 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21446 ) );
  MUX \u_a23_mem/U21528  ( .IN0(\u_a23_mem/n21444 ), .IN1(\u_a23_mem/n21443 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21445 ) );
  MUX \u_a23_mem/U21527  ( .IN0(\u_a23_mem/e_mem[1][6] ), .IN1(
        \u_a23_mem/e_mem[17][6] ), .SEL(m_address[4]), .F(\u_a23_mem/n21444 )
         );
  MUX \u_a23_mem/U21526  ( .IN0(\u_a23_mem/e_mem[9][6] ), .IN1(
        \u_a23_mem/e_mem[25][6] ), .SEL(m_address[4]), .F(\u_a23_mem/n21443 )
         );
  MUX \u_a23_mem/U21525  ( .IN0(\u_a23_mem/n21441 ), .IN1(\u_a23_mem/n21440 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21442 ) );
  MUX \u_a23_mem/U21524  ( .IN0(\u_a23_mem/e_mem[5][6] ), .IN1(
        \u_a23_mem/e_mem[21][6] ), .SEL(m_address[4]), .F(\u_a23_mem/n21441 )
         );
  MUX \u_a23_mem/U21523  ( .IN0(\u_a23_mem/e_mem[13][6] ), .IN1(
        \u_a23_mem/e_mem[29][6] ), .SEL(m_address[4]), .F(\u_a23_mem/n21440 )
         );
  MUX \u_a23_mem/U21522  ( .IN0(\u_a23_mem/n21438 ), .IN1(\u_a23_mem/n21435 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21439 ) );
  MUX \u_a23_mem/U21521  ( .IN0(\u_a23_mem/n21437 ), .IN1(\u_a23_mem/n21436 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21438 ) );
  MUX \u_a23_mem/U21520  ( .IN0(\u_a23_mem/e_mem[3][6] ), .IN1(
        \u_a23_mem/e_mem[19][6] ), .SEL(m_address[4]), .F(\u_a23_mem/n21437 )
         );
  MUX \u_a23_mem/U21519  ( .IN0(\u_a23_mem/e_mem[11][6] ), .IN1(
        \u_a23_mem/e_mem[27][6] ), .SEL(m_address[4]), .F(\u_a23_mem/n21436 )
         );
  MUX \u_a23_mem/U21518  ( .IN0(\u_a23_mem/n21434 ), .IN1(\u_a23_mem/n21433 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21435 ) );
  MUX \u_a23_mem/U21517  ( .IN0(\u_a23_mem/e_mem[7][6] ), .IN1(
        \u_a23_mem/e_mem[23][6] ), .SEL(m_address[4]), .F(\u_a23_mem/n21434 )
         );
  MUX \u_a23_mem/U21516  ( .IN0(\u_a23_mem/e_mem[15][6] ), .IN1(
        \u_a23_mem/e_mem[31][6] ), .SEL(m_address[4]), .F(\u_a23_mem/n21433 )
         );
  MUX \u_a23_mem/U21514  ( .IN0(\u_a23_mem/n21430 ), .IN1(\u_a23_mem/n21427 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21431 ) );
  MUX \u_a23_mem/U21513  ( .IN0(\u_a23_mem/n21429 ), .IN1(\u_a23_mem/n21428 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21430 ) );
  MUX \u_a23_mem/U21512  ( .IN0(\u_a23_mem/e_mem[2][6] ), .IN1(
        \u_a23_mem/e_mem[18][6] ), .SEL(m_address[4]), .F(\u_a23_mem/n21429 )
         );
  MUX \u_a23_mem/U21511  ( .IN0(\u_a23_mem/e_mem[10][6] ), .IN1(
        \u_a23_mem/e_mem[26][6] ), .SEL(m_address[4]), .F(\u_a23_mem/n21428 )
         );
  MUX \u_a23_mem/U21510  ( .IN0(\u_a23_mem/n21426 ), .IN1(\u_a23_mem/n21425 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21427 ) );
  MUX \u_a23_mem/U21509  ( .IN0(\u_a23_mem/e_mem[6][6] ), .IN1(
        \u_a23_mem/e_mem[22][6] ), .SEL(m_address[4]), .F(\u_a23_mem/n21426 )
         );
  MUX \u_a23_mem/U21508  ( .IN0(\u_a23_mem/e_mem[14][6] ), .IN1(
        \u_a23_mem/e_mem[30][6] ), .SEL(m_address[4]), .F(\u_a23_mem/n21425 )
         );
  MUX \u_a23_mem/U21499  ( .IN0(\u_a23_mem/n21416 ), .IN1(\u_a23_mem/n21413 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21417 ) );
  MUX \u_a23_mem/U21498  ( .IN0(\u_a23_mem/n21415 ), .IN1(\u_a23_mem/n21414 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21416 ) );
  MUX \u_a23_mem/U21497  ( .IN0(\u_a23_mem/e_mem[1][5] ), .IN1(
        \u_a23_mem/e_mem[17][5] ), .SEL(m_address[4]), .F(\u_a23_mem/n21415 )
         );
  MUX \u_a23_mem/U21496  ( .IN0(\u_a23_mem/e_mem[9][5] ), .IN1(
        \u_a23_mem/e_mem[25][5] ), .SEL(m_address[4]), .F(\u_a23_mem/n21414 )
         );
  MUX \u_a23_mem/U21495  ( .IN0(\u_a23_mem/n21412 ), .IN1(\u_a23_mem/n21411 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21413 ) );
  MUX \u_a23_mem/U21494  ( .IN0(\u_a23_mem/e_mem[5][5] ), .IN1(
        \u_a23_mem/e_mem[21][5] ), .SEL(m_address[4]), .F(\u_a23_mem/n21412 )
         );
  MUX \u_a23_mem/U21493  ( .IN0(\u_a23_mem/e_mem[13][5] ), .IN1(
        \u_a23_mem/e_mem[29][5] ), .SEL(m_address[4]), .F(\u_a23_mem/n21411 )
         );
  MUX \u_a23_mem/U21492  ( .IN0(\u_a23_mem/n21409 ), .IN1(\u_a23_mem/n21406 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21410 ) );
  MUX \u_a23_mem/U21491  ( .IN0(\u_a23_mem/n21408 ), .IN1(\u_a23_mem/n21407 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21409 ) );
  MUX \u_a23_mem/U21490  ( .IN0(\u_a23_mem/e_mem[3][5] ), .IN1(
        \u_a23_mem/e_mem[19][5] ), .SEL(m_address[4]), .F(\u_a23_mem/n21408 )
         );
  MUX \u_a23_mem/U21489  ( .IN0(\u_a23_mem/e_mem[11][5] ), .IN1(
        \u_a23_mem/e_mem[27][5] ), .SEL(m_address[4]), .F(\u_a23_mem/n21407 )
         );
  MUX \u_a23_mem/U21488  ( .IN0(\u_a23_mem/n21405 ), .IN1(\u_a23_mem/n21404 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21406 ) );
  MUX \u_a23_mem/U21487  ( .IN0(\u_a23_mem/e_mem[7][5] ), .IN1(
        \u_a23_mem/e_mem[23][5] ), .SEL(m_address[4]), .F(\u_a23_mem/n21405 )
         );
  MUX \u_a23_mem/U21486  ( .IN0(\u_a23_mem/e_mem[15][5] ), .IN1(
        \u_a23_mem/e_mem[31][5] ), .SEL(m_address[4]), .F(\u_a23_mem/n21404 )
         );
  MUX \u_a23_mem/U21484  ( .IN0(\u_a23_mem/n21401 ), .IN1(\u_a23_mem/n21398 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21402 ) );
  MUX \u_a23_mem/U21483  ( .IN0(\u_a23_mem/n21400 ), .IN1(\u_a23_mem/n21399 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21401 ) );
  MUX \u_a23_mem/U21482  ( .IN0(\u_a23_mem/e_mem[2][5] ), .IN1(
        \u_a23_mem/e_mem[18][5] ), .SEL(m_address[4]), .F(\u_a23_mem/n21400 )
         );
  MUX \u_a23_mem/U21481  ( .IN0(\u_a23_mem/e_mem[10][5] ), .IN1(
        \u_a23_mem/e_mem[26][5] ), .SEL(m_address[4]), .F(\u_a23_mem/n21399 )
         );
  MUX \u_a23_mem/U21480  ( .IN0(\u_a23_mem/n21397 ), .IN1(\u_a23_mem/n21396 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21398 ) );
  MUX \u_a23_mem/U21479  ( .IN0(\u_a23_mem/e_mem[6][5] ), .IN1(
        \u_a23_mem/e_mem[22][5] ), .SEL(m_address[4]), .F(\u_a23_mem/n21397 )
         );
  MUX \u_a23_mem/U21478  ( .IN0(\u_a23_mem/e_mem[14][5] ), .IN1(
        \u_a23_mem/e_mem[30][5] ), .SEL(m_address[4]), .F(\u_a23_mem/n21396 )
         );
  MUX \u_a23_mem/U21469  ( .IN0(\u_a23_mem/n21387 ), .IN1(\u_a23_mem/n21384 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21388 ) );
  MUX \u_a23_mem/U21468  ( .IN0(\u_a23_mem/n21386 ), .IN1(\u_a23_mem/n21385 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21387 ) );
  MUX \u_a23_mem/U21467  ( .IN0(\u_a23_mem/e_mem[1][4] ), .IN1(
        \u_a23_mem/e_mem[17][4] ), .SEL(m_address[4]), .F(\u_a23_mem/n21386 )
         );
  MUX \u_a23_mem/U21466  ( .IN0(\u_a23_mem/e_mem[9][4] ), .IN1(
        \u_a23_mem/e_mem[25][4] ), .SEL(m_address[4]), .F(\u_a23_mem/n21385 )
         );
  MUX \u_a23_mem/U21465  ( .IN0(\u_a23_mem/n21383 ), .IN1(\u_a23_mem/n21382 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21384 ) );
  MUX \u_a23_mem/U21464  ( .IN0(\u_a23_mem/e_mem[5][4] ), .IN1(
        \u_a23_mem/e_mem[21][4] ), .SEL(m_address[4]), .F(\u_a23_mem/n21383 )
         );
  MUX \u_a23_mem/U21463  ( .IN0(\u_a23_mem/e_mem[13][4] ), .IN1(
        \u_a23_mem/e_mem[29][4] ), .SEL(m_address[4]), .F(\u_a23_mem/n21382 )
         );
  MUX \u_a23_mem/U21462  ( .IN0(\u_a23_mem/n21380 ), .IN1(\u_a23_mem/n21377 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21381 ) );
  MUX \u_a23_mem/U21461  ( .IN0(\u_a23_mem/n21379 ), .IN1(\u_a23_mem/n21378 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21380 ) );
  MUX \u_a23_mem/U21460  ( .IN0(\u_a23_mem/e_mem[3][4] ), .IN1(
        \u_a23_mem/e_mem[19][4] ), .SEL(m_address[4]), .F(\u_a23_mem/n21379 )
         );
  MUX \u_a23_mem/U21459  ( .IN0(\u_a23_mem/e_mem[11][4] ), .IN1(
        \u_a23_mem/e_mem[27][4] ), .SEL(m_address[4]), .F(\u_a23_mem/n21378 )
         );
  MUX \u_a23_mem/U21458  ( .IN0(\u_a23_mem/n21376 ), .IN1(\u_a23_mem/n21375 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21377 ) );
  MUX \u_a23_mem/U21457  ( .IN0(\u_a23_mem/e_mem[7][4] ), .IN1(
        \u_a23_mem/e_mem[23][4] ), .SEL(m_address[4]), .F(\u_a23_mem/n21376 )
         );
  MUX \u_a23_mem/U21456  ( .IN0(\u_a23_mem/e_mem[15][4] ), .IN1(
        \u_a23_mem/e_mem[31][4] ), .SEL(m_address[4]), .F(\u_a23_mem/n21375 )
         );
  MUX \u_a23_mem/U21454  ( .IN0(\u_a23_mem/n21372 ), .IN1(\u_a23_mem/n21369 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21373 ) );
  MUX \u_a23_mem/U21453  ( .IN0(\u_a23_mem/n21371 ), .IN1(\u_a23_mem/n21370 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21372 ) );
  MUX \u_a23_mem/U21452  ( .IN0(\u_a23_mem/e_mem[2][4] ), .IN1(
        \u_a23_mem/e_mem[18][4] ), .SEL(m_address[4]), .F(\u_a23_mem/n21371 )
         );
  MUX \u_a23_mem/U21451  ( .IN0(\u_a23_mem/e_mem[10][4] ), .IN1(
        \u_a23_mem/e_mem[26][4] ), .SEL(m_address[4]), .F(\u_a23_mem/n21370 )
         );
  MUX \u_a23_mem/U21450  ( .IN0(\u_a23_mem/n21368 ), .IN1(\u_a23_mem/n21367 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21369 ) );
  MUX \u_a23_mem/U21449  ( .IN0(\u_a23_mem/e_mem[6][4] ), .IN1(
        \u_a23_mem/e_mem[22][4] ), .SEL(m_address[4]), .F(\u_a23_mem/n21368 )
         );
  MUX \u_a23_mem/U21448  ( .IN0(\u_a23_mem/e_mem[14][4] ), .IN1(
        \u_a23_mem/e_mem[30][4] ), .SEL(m_address[4]), .F(\u_a23_mem/n21367 )
         );
  MUX \u_a23_mem/U21439  ( .IN0(\u_a23_mem/n21358 ), .IN1(\u_a23_mem/n21355 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21359 ) );
  MUX \u_a23_mem/U21438  ( .IN0(\u_a23_mem/n21357 ), .IN1(\u_a23_mem/n21356 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21358 ) );
  MUX \u_a23_mem/U21437  ( .IN0(\u_a23_mem/e_mem[1][3] ), .IN1(
        \u_a23_mem/e_mem[17][3] ), .SEL(m_address[4]), .F(\u_a23_mem/n21357 )
         );
  MUX \u_a23_mem/U21436  ( .IN0(\u_a23_mem/e_mem[9][3] ), .IN1(
        \u_a23_mem/e_mem[25][3] ), .SEL(m_address[4]), .F(\u_a23_mem/n21356 )
         );
  MUX \u_a23_mem/U21435  ( .IN0(\u_a23_mem/n21354 ), .IN1(\u_a23_mem/n21353 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21355 ) );
  MUX \u_a23_mem/U21434  ( .IN0(\u_a23_mem/e_mem[5][3] ), .IN1(
        \u_a23_mem/e_mem[21][3] ), .SEL(m_address[4]), .F(\u_a23_mem/n21354 )
         );
  MUX \u_a23_mem/U21433  ( .IN0(\u_a23_mem/e_mem[13][3] ), .IN1(
        \u_a23_mem/e_mem[29][3] ), .SEL(m_address[4]), .F(\u_a23_mem/n21353 )
         );
  MUX \u_a23_mem/U21432  ( .IN0(\u_a23_mem/n21351 ), .IN1(\u_a23_mem/n21348 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21352 ) );
  MUX \u_a23_mem/U21431  ( .IN0(\u_a23_mem/n21350 ), .IN1(\u_a23_mem/n21349 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21351 ) );
  MUX \u_a23_mem/U21430  ( .IN0(\u_a23_mem/e_mem[3][3] ), .IN1(
        \u_a23_mem/e_mem[19][3] ), .SEL(m_address[4]), .F(\u_a23_mem/n21350 )
         );
  MUX \u_a23_mem/U21429  ( .IN0(\u_a23_mem/e_mem[11][3] ), .IN1(
        \u_a23_mem/e_mem[27][3] ), .SEL(m_address[4]), .F(\u_a23_mem/n21349 )
         );
  MUX \u_a23_mem/U21428  ( .IN0(\u_a23_mem/n21347 ), .IN1(\u_a23_mem/n21346 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21348 ) );
  MUX \u_a23_mem/U21427  ( .IN0(\u_a23_mem/e_mem[7][3] ), .IN1(
        \u_a23_mem/e_mem[23][3] ), .SEL(m_address[4]), .F(\u_a23_mem/n21347 )
         );
  MUX \u_a23_mem/U21426  ( .IN0(\u_a23_mem/e_mem[15][3] ), .IN1(
        \u_a23_mem/e_mem[31][3] ), .SEL(m_address[4]), .F(\u_a23_mem/n21346 )
         );
  MUX \u_a23_mem/U21424  ( .IN0(\u_a23_mem/n21343 ), .IN1(\u_a23_mem/n21340 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21344 ) );
  MUX \u_a23_mem/U21423  ( .IN0(\u_a23_mem/n21342 ), .IN1(\u_a23_mem/n21341 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21343 ) );
  MUX \u_a23_mem/U21422  ( .IN0(\u_a23_mem/e_mem[2][3] ), .IN1(
        \u_a23_mem/e_mem[18][3] ), .SEL(m_address[4]), .F(\u_a23_mem/n21342 )
         );
  MUX \u_a23_mem/U21421  ( .IN0(\u_a23_mem/e_mem[10][3] ), .IN1(
        \u_a23_mem/e_mem[26][3] ), .SEL(m_address[4]), .F(\u_a23_mem/n21341 )
         );
  MUX \u_a23_mem/U21420  ( .IN0(\u_a23_mem/n21339 ), .IN1(\u_a23_mem/n21338 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21340 ) );
  MUX \u_a23_mem/U21419  ( .IN0(\u_a23_mem/e_mem[6][3] ), .IN1(
        \u_a23_mem/e_mem[22][3] ), .SEL(m_address[4]), .F(\u_a23_mem/n21339 )
         );
  MUX \u_a23_mem/U21418  ( .IN0(\u_a23_mem/e_mem[14][3] ), .IN1(
        \u_a23_mem/e_mem[30][3] ), .SEL(m_address[4]), .F(\u_a23_mem/n21338 )
         );
  MUX \u_a23_mem/U21409  ( .IN0(\u_a23_mem/n21329 ), .IN1(\u_a23_mem/n21326 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21330 ) );
  MUX \u_a23_mem/U21408  ( .IN0(\u_a23_mem/n21328 ), .IN1(\u_a23_mem/n21327 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21329 ) );
  MUX \u_a23_mem/U21407  ( .IN0(\u_a23_mem/e_mem[1][2] ), .IN1(
        \u_a23_mem/e_mem[17][2] ), .SEL(m_address[4]), .F(\u_a23_mem/n21328 )
         );
  MUX \u_a23_mem/U21406  ( .IN0(\u_a23_mem/e_mem[9][2] ), .IN1(
        \u_a23_mem/e_mem[25][2] ), .SEL(m_address[4]), .F(\u_a23_mem/n21327 )
         );
  MUX \u_a23_mem/U21405  ( .IN0(\u_a23_mem/n21325 ), .IN1(\u_a23_mem/n21324 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21326 ) );
  MUX \u_a23_mem/U21404  ( .IN0(\u_a23_mem/e_mem[5][2] ), .IN1(
        \u_a23_mem/e_mem[21][2] ), .SEL(m_address[4]), .F(\u_a23_mem/n21325 )
         );
  MUX \u_a23_mem/U21403  ( .IN0(\u_a23_mem/e_mem[13][2] ), .IN1(
        \u_a23_mem/e_mem[29][2] ), .SEL(m_address[4]), .F(\u_a23_mem/n21324 )
         );
  MUX \u_a23_mem/U21402  ( .IN0(\u_a23_mem/n21322 ), .IN1(\u_a23_mem/n21319 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21323 ) );
  MUX \u_a23_mem/U21401  ( .IN0(\u_a23_mem/n21321 ), .IN1(\u_a23_mem/n21320 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21322 ) );
  MUX \u_a23_mem/U21400  ( .IN0(\u_a23_mem/e_mem[3][2] ), .IN1(
        \u_a23_mem/e_mem[19][2] ), .SEL(m_address[4]), .F(\u_a23_mem/n21321 )
         );
  MUX \u_a23_mem/U21399  ( .IN0(\u_a23_mem/e_mem[11][2] ), .IN1(
        \u_a23_mem/e_mem[27][2] ), .SEL(m_address[4]), .F(\u_a23_mem/n21320 )
         );
  MUX \u_a23_mem/U21398  ( .IN0(\u_a23_mem/n21318 ), .IN1(\u_a23_mem/n21317 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21319 ) );
  MUX \u_a23_mem/U21397  ( .IN0(\u_a23_mem/e_mem[7][2] ), .IN1(
        \u_a23_mem/e_mem[23][2] ), .SEL(m_address[4]), .F(\u_a23_mem/n21318 )
         );
  MUX \u_a23_mem/U21396  ( .IN0(\u_a23_mem/e_mem[15][2] ), .IN1(
        \u_a23_mem/e_mem[31][2] ), .SEL(m_address[4]), .F(\u_a23_mem/n21317 )
         );
  MUX \u_a23_mem/U21394  ( .IN0(\u_a23_mem/n21314 ), .IN1(\u_a23_mem/n21311 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21315 ) );
  MUX \u_a23_mem/U21393  ( .IN0(\u_a23_mem/n21313 ), .IN1(\u_a23_mem/n21312 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21314 ) );
  MUX \u_a23_mem/U21392  ( .IN0(\u_a23_mem/e_mem[2][2] ), .IN1(
        \u_a23_mem/e_mem[18][2] ), .SEL(m_address[4]), .F(\u_a23_mem/n21313 )
         );
  MUX \u_a23_mem/U21391  ( .IN0(\u_a23_mem/e_mem[10][2] ), .IN1(
        \u_a23_mem/e_mem[26][2] ), .SEL(m_address[4]), .F(\u_a23_mem/n21312 )
         );
  MUX \u_a23_mem/U21390  ( .IN0(\u_a23_mem/n21310 ), .IN1(\u_a23_mem/n21309 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21311 ) );
  MUX \u_a23_mem/U21389  ( .IN0(\u_a23_mem/e_mem[6][2] ), .IN1(
        \u_a23_mem/e_mem[22][2] ), .SEL(m_address[4]), .F(\u_a23_mem/n21310 )
         );
  MUX \u_a23_mem/U21388  ( .IN0(\u_a23_mem/e_mem[14][2] ), .IN1(
        \u_a23_mem/e_mem[30][2] ), .SEL(m_address[4]), .F(\u_a23_mem/n21309 )
         );
  MUX \u_a23_mem/U21379  ( .IN0(\u_a23_mem/n21300 ), .IN1(\u_a23_mem/n21297 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21301 ) );
  MUX \u_a23_mem/U21378  ( .IN0(\u_a23_mem/n21299 ), .IN1(\u_a23_mem/n21298 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21300 ) );
  MUX \u_a23_mem/U21377  ( .IN0(\u_a23_mem/e_mem[1][1] ), .IN1(
        \u_a23_mem/e_mem[17][1] ), .SEL(m_address[4]), .F(\u_a23_mem/n21299 )
         );
  MUX \u_a23_mem/U21376  ( .IN0(\u_a23_mem/e_mem[9][1] ), .IN1(
        \u_a23_mem/e_mem[25][1] ), .SEL(m_address[4]), .F(\u_a23_mem/n21298 )
         );
  MUX \u_a23_mem/U21375  ( .IN0(\u_a23_mem/n21296 ), .IN1(\u_a23_mem/n21295 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21297 ) );
  MUX \u_a23_mem/U21374  ( .IN0(\u_a23_mem/e_mem[5][1] ), .IN1(
        \u_a23_mem/e_mem[21][1] ), .SEL(m_address[4]), .F(\u_a23_mem/n21296 )
         );
  MUX \u_a23_mem/U21373  ( .IN0(\u_a23_mem/e_mem[13][1] ), .IN1(
        \u_a23_mem/e_mem[29][1] ), .SEL(m_address[4]), .F(\u_a23_mem/n21295 )
         );
  MUX \u_a23_mem/U21372  ( .IN0(\u_a23_mem/n21293 ), .IN1(\u_a23_mem/n21290 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21294 ) );
  MUX \u_a23_mem/U21371  ( .IN0(\u_a23_mem/n21292 ), .IN1(\u_a23_mem/n21291 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21293 ) );
  MUX \u_a23_mem/U21370  ( .IN0(\u_a23_mem/e_mem[3][1] ), .IN1(
        \u_a23_mem/e_mem[19][1] ), .SEL(m_address[4]), .F(\u_a23_mem/n21292 )
         );
  MUX \u_a23_mem/U21369  ( .IN0(\u_a23_mem/e_mem[11][1] ), .IN1(
        \u_a23_mem/e_mem[27][1] ), .SEL(m_address[4]), .F(\u_a23_mem/n21291 )
         );
  MUX \u_a23_mem/U21368  ( .IN0(\u_a23_mem/n21289 ), .IN1(\u_a23_mem/n21288 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21290 ) );
  MUX \u_a23_mem/U21367  ( .IN0(\u_a23_mem/e_mem[7][1] ), .IN1(
        \u_a23_mem/e_mem[23][1] ), .SEL(m_address[4]), .F(\u_a23_mem/n21289 )
         );
  MUX \u_a23_mem/U21366  ( .IN0(\u_a23_mem/e_mem[15][1] ), .IN1(
        \u_a23_mem/e_mem[31][1] ), .SEL(m_address[4]), .F(\u_a23_mem/n21288 )
         );
  MUX \u_a23_mem/U21364  ( .IN0(\u_a23_mem/n21285 ), .IN1(\u_a23_mem/n21282 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21286 ) );
  MUX \u_a23_mem/U21363  ( .IN0(\u_a23_mem/n21284 ), .IN1(\u_a23_mem/n21283 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21285 ) );
  MUX \u_a23_mem/U21362  ( .IN0(\u_a23_mem/e_mem[2][1] ), .IN1(
        \u_a23_mem/e_mem[18][1] ), .SEL(m_address[4]), .F(\u_a23_mem/n21284 )
         );
  MUX \u_a23_mem/U21361  ( .IN0(\u_a23_mem/e_mem[10][1] ), .IN1(
        \u_a23_mem/e_mem[26][1] ), .SEL(m_address[4]), .F(\u_a23_mem/n21283 )
         );
  MUX \u_a23_mem/U21360  ( .IN0(\u_a23_mem/n21281 ), .IN1(\u_a23_mem/n21280 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21282 ) );
  MUX \u_a23_mem/U21359  ( .IN0(\u_a23_mem/e_mem[6][1] ), .IN1(
        \u_a23_mem/e_mem[22][1] ), .SEL(m_address[4]), .F(\u_a23_mem/n21281 )
         );
  MUX \u_a23_mem/U21358  ( .IN0(\u_a23_mem/e_mem[14][1] ), .IN1(
        \u_a23_mem/e_mem[30][1] ), .SEL(m_address[4]), .F(\u_a23_mem/n21280 )
         );
  MUX \u_a23_mem/U21349  ( .IN0(\u_a23_mem/n21271 ), .IN1(\u_a23_mem/n21268 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21272 ) );
  MUX \u_a23_mem/U21348  ( .IN0(\u_a23_mem/n21270 ), .IN1(\u_a23_mem/n21269 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21271 ) );
  MUX \u_a23_mem/U21347  ( .IN0(\u_a23_mem/e_mem[1][0] ), .IN1(
        \u_a23_mem/e_mem[17][0] ), .SEL(m_address[4]), .F(\u_a23_mem/n21270 )
         );
  MUX \u_a23_mem/U21346  ( .IN0(\u_a23_mem/e_mem[9][0] ), .IN1(
        \u_a23_mem/e_mem[25][0] ), .SEL(m_address[4]), .F(\u_a23_mem/n21269 )
         );
  MUX \u_a23_mem/U21345  ( .IN0(\u_a23_mem/n21267 ), .IN1(\u_a23_mem/n21266 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21268 ) );
  MUX \u_a23_mem/U21344  ( .IN0(\u_a23_mem/e_mem[5][0] ), .IN1(
        \u_a23_mem/e_mem[21][0] ), .SEL(m_address[4]), .F(\u_a23_mem/n21267 )
         );
  MUX \u_a23_mem/U21343  ( .IN0(\u_a23_mem/e_mem[13][0] ), .IN1(
        \u_a23_mem/e_mem[29][0] ), .SEL(m_address[4]), .F(\u_a23_mem/n21266 )
         );
  MUX \u_a23_mem/U21342  ( .IN0(\u_a23_mem/n21264 ), .IN1(\u_a23_mem/n21261 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21265 ) );
  MUX \u_a23_mem/U21341  ( .IN0(\u_a23_mem/n21263 ), .IN1(\u_a23_mem/n21262 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21264 ) );
  MUX \u_a23_mem/U21340  ( .IN0(\u_a23_mem/e_mem[3][0] ), .IN1(
        \u_a23_mem/e_mem[19][0] ), .SEL(m_address[4]), .F(\u_a23_mem/n21263 )
         );
  MUX \u_a23_mem/U21339  ( .IN0(\u_a23_mem/e_mem[11][0] ), .IN1(
        \u_a23_mem/e_mem[27][0] ), .SEL(m_address[4]), .F(\u_a23_mem/n21262 )
         );
  MUX \u_a23_mem/U21338  ( .IN0(\u_a23_mem/n21260 ), .IN1(\u_a23_mem/n21259 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21261 ) );
  MUX \u_a23_mem/U21337  ( .IN0(\u_a23_mem/e_mem[7][0] ), .IN1(
        \u_a23_mem/e_mem[23][0] ), .SEL(m_address[4]), .F(\u_a23_mem/n21260 )
         );
  MUX \u_a23_mem/U21336  ( .IN0(\u_a23_mem/e_mem[15][0] ), .IN1(
        \u_a23_mem/e_mem[31][0] ), .SEL(m_address[4]), .F(\u_a23_mem/n21259 )
         );
  MUX \u_a23_mem/U21334  ( .IN0(\u_a23_mem/n21256 ), .IN1(\u_a23_mem/n21253 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21257 ) );
  MUX \u_a23_mem/U21333  ( .IN0(\u_a23_mem/n21255 ), .IN1(\u_a23_mem/n21254 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21256 ) );
  MUX \u_a23_mem/U21332  ( .IN0(\u_a23_mem/e_mem[2][0] ), .IN1(
        \u_a23_mem/e_mem[18][0] ), .SEL(m_address[4]), .F(\u_a23_mem/n21255 )
         );
  MUX \u_a23_mem/U21331  ( .IN0(\u_a23_mem/e_mem[10][0] ), .IN1(
        \u_a23_mem/e_mem[26][0] ), .SEL(m_address[4]), .F(\u_a23_mem/n21254 )
         );
  MUX \u_a23_mem/U21330  ( .IN0(\u_a23_mem/n21252 ), .IN1(\u_a23_mem/n21251 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21253 ) );
  MUX \u_a23_mem/U21329  ( .IN0(\u_a23_mem/e_mem[6][0] ), .IN1(
        \u_a23_mem/e_mem[22][0] ), .SEL(m_address[4]), .F(\u_a23_mem/n21252 )
         );
  MUX \u_a23_mem/U21328  ( .IN0(\u_a23_mem/e_mem[14][0] ), .IN1(
        \u_a23_mem/e_mem[30][0] ), .SEL(m_address[4]), .F(\u_a23_mem/n21251 )
         );
  MUX \u_a23_mem/U21279  ( .IN0(\u_a23_mem/n21218 ), .IN1(\u_a23_mem/n21215 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21219 ) );
  MUX \u_a23_mem/U21278  ( .IN0(\u_a23_mem/n21217 ), .IN1(\u_a23_mem/n21216 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21218 ) );
  MUX \u_a23_mem/U21277  ( .IN0(o[15]), .IN1(o[143]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21217 ) );
  MUX \u_a23_mem/U21276  ( .IN0(o[79]), .IN1(o[207]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21216 ) );
  MUX \u_a23_mem/U21275  ( .IN0(\u_a23_mem/n21214 ), .IN1(\u_a23_mem/n21213 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21215 ) );
  MUX \u_a23_mem/U21274  ( .IN0(o[47]), .IN1(o[175]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21214 ) );
  MUX \u_a23_mem/U21273  ( .IN0(o[111]), .IN1(o[239]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21213 ) );
  MUX \u_a23_mem/U21272  ( .IN0(\u_a23_mem/n21211 ), .IN1(\u_a23_mem/n21208 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21212 ) );
  MUX \u_a23_mem/U21271  ( .IN0(\u_a23_mem/n21210 ), .IN1(\u_a23_mem/n21209 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21211 ) );
  MUX \u_a23_mem/U21270  ( .IN0(o[31]), .IN1(o[159]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21210 ) );
  MUX \u_a23_mem/U21269  ( .IN0(o[95]), .IN1(o[223]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21209 ) );
  MUX \u_a23_mem/U21268  ( .IN0(\u_a23_mem/n21207 ), .IN1(\u_a23_mem/n21206 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21208 ) );
  MUX \u_a23_mem/U21267  ( .IN0(o[63]), .IN1(o[191]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21207 ) );
  MUX \u_a23_mem/U21266  ( .IN0(o[127]), .IN1(o[255]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21206 ) );
  MUX \u_a23_mem/U21264  ( .IN0(\u_a23_mem/n21203 ), .IN1(\u_a23_mem/n21200 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21204 ) );
  MUX \u_a23_mem/U21263  ( .IN0(\u_a23_mem/n21202 ), .IN1(\u_a23_mem/n21201 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21203 ) );
  MUX \u_a23_mem/U21262  ( .IN0(o[23]), .IN1(o[151]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21202 ) );
  MUX \u_a23_mem/U21261  ( .IN0(o[87]), .IN1(o[215]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21201 ) );
  MUX \u_a23_mem/U21260  ( .IN0(\u_a23_mem/n21199 ), .IN1(\u_a23_mem/n21198 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21200 ) );
  MUX \u_a23_mem/U21259  ( .IN0(o[55]), .IN1(o[183]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21199 ) );
  MUX \u_a23_mem/U21258  ( .IN0(o[119]), .IN1(o[247]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21198 ) );
  MUX \u_a23_mem/U21249  ( .IN0(\u_a23_mem/n21189 ), .IN1(\u_a23_mem/n21186 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21190 ) );
  MUX \u_a23_mem/U21248  ( .IN0(\u_a23_mem/n21188 ), .IN1(\u_a23_mem/n21187 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21189 ) );
  MUX \u_a23_mem/U21247  ( .IN0(o[14]), .IN1(o[142]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21188 ) );
  MUX \u_a23_mem/U21246  ( .IN0(o[78]), .IN1(o[206]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21187 ) );
  MUX \u_a23_mem/U21245  ( .IN0(\u_a23_mem/n21185 ), .IN1(\u_a23_mem/n21184 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21186 ) );
  MUX \u_a23_mem/U21244  ( .IN0(o[46]), .IN1(o[174]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21185 ) );
  MUX \u_a23_mem/U21243  ( .IN0(o[110]), .IN1(o[238]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21184 ) );
  MUX \u_a23_mem/U21242  ( .IN0(\u_a23_mem/n21182 ), .IN1(\u_a23_mem/n21179 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21183 ) );
  MUX \u_a23_mem/U21241  ( .IN0(\u_a23_mem/n21181 ), .IN1(\u_a23_mem/n21180 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21182 ) );
  MUX \u_a23_mem/U21240  ( .IN0(o[30]), .IN1(o[158]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21181 ) );
  MUX \u_a23_mem/U21239  ( .IN0(o[94]), .IN1(o[222]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21180 ) );
  MUX \u_a23_mem/U21238  ( .IN0(\u_a23_mem/n21178 ), .IN1(\u_a23_mem/n21177 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21179 ) );
  MUX \u_a23_mem/U21237  ( .IN0(o[62]), .IN1(o[190]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21178 ) );
  MUX \u_a23_mem/U21236  ( .IN0(o[126]), .IN1(o[254]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21177 ) );
  MUX \u_a23_mem/U21234  ( .IN0(\u_a23_mem/n21174 ), .IN1(\u_a23_mem/n21171 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21175 ) );
  MUX \u_a23_mem/U21233  ( .IN0(\u_a23_mem/n21173 ), .IN1(\u_a23_mem/n21172 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21174 ) );
  MUX \u_a23_mem/U21232  ( .IN0(o[22]), .IN1(o[150]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21173 ) );
  MUX \u_a23_mem/U21231  ( .IN0(o[86]), .IN1(o[214]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21172 ) );
  MUX \u_a23_mem/U21230  ( .IN0(\u_a23_mem/n21170 ), .IN1(\u_a23_mem/n21169 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21171 ) );
  MUX \u_a23_mem/U21229  ( .IN0(o[54]), .IN1(o[182]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21170 ) );
  MUX \u_a23_mem/U21228  ( .IN0(o[118]), .IN1(o[246]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21169 ) );
  MUX \u_a23_mem/U21219  ( .IN0(\u_a23_mem/n21160 ), .IN1(\u_a23_mem/n21157 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21161 ) );
  MUX \u_a23_mem/U21218  ( .IN0(\u_a23_mem/n21159 ), .IN1(\u_a23_mem/n21158 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21160 ) );
  MUX \u_a23_mem/U21217  ( .IN0(o[13]), .IN1(o[141]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21159 ) );
  MUX \u_a23_mem/U21216  ( .IN0(o[77]), .IN1(o[205]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21158 ) );
  MUX \u_a23_mem/U21215  ( .IN0(\u_a23_mem/n21156 ), .IN1(\u_a23_mem/n21155 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21157 ) );
  MUX \u_a23_mem/U21214  ( .IN0(o[45]), .IN1(o[173]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21156 ) );
  MUX \u_a23_mem/U21213  ( .IN0(o[109]), .IN1(o[237]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21155 ) );
  MUX \u_a23_mem/U21212  ( .IN0(\u_a23_mem/n21153 ), .IN1(\u_a23_mem/n21150 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21154 ) );
  MUX \u_a23_mem/U21211  ( .IN0(\u_a23_mem/n21152 ), .IN1(\u_a23_mem/n21151 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21153 ) );
  MUX \u_a23_mem/U21210  ( .IN0(o[29]), .IN1(o[157]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21152 ) );
  MUX \u_a23_mem/U21209  ( .IN0(o[93]), .IN1(o[221]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21151 ) );
  MUX \u_a23_mem/U21208  ( .IN0(\u_a23_mem/n21149 ), .IN1(\u_a23_mem/n21148 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21150 ) );
  MUX \u_a23_mem/U21207  ( .IN0(o[61]), .IN1(o[189]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21149 ) );
  MUX \u_a23_mem/U21206  ( .IN0(o[125]), .IN1(o[253]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21148 ) );
  MUX \u_a23_mem/U21204  ( .IN0(\u_a23_mem/n21145 ), .IN1(\u_a23_mem/n21142 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21146 ) );
  MUX \u_a23_mem/U21203  ( .IN0(\u_a23_mem/n21144 ), .IN1(\u_a23_mem/n21143 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21145 ) );
  MUX \u_a23_mem/U21202  ( .IN0(o[21]), .IN1(o[149]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21144 ) );
  MUX \u_a23_mem/U21201  ( .IN0(o[85]), .IN1(o[213]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21143 ) );
  MUX \u_a23_mem/U21200  ( .IN0(\u_a23_mem/n21141 ), .IN1(\u_a23_mem/n21140 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21142 ) );
  MUX \u_a23_mem/U21199  ( .IN0(o[53]), .IN1(o[181]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21141 ) );
  MUX \u_a23_mem/U21198  ( .IN0(o[117]), .IN1(o[245]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21140 ) );
  MUX \u_a23_mem/U21189  ( .IN0(\u_a23_mem/n21131 ), .IN1(\u_a23_mem/n21128 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21132 ) );
  MUX \u_a23_mem/U21188  ( .IN0(\u_a23_mem/n21130 ), .IN1(\u_a23_mem/n21129 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21131 ) );
  MUX \u_a23_mem/U21187  ( .IN0(o[12]), .IN1(o[140]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21130 ) );
  MUX \u_a23_mem/U21186  ( .IN0(o[76]), .IN1(o[204]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21129 ) );
  MUX \u_a23_mem/U21185  ( .IN0(\u_a23_mem/n21127 ), .IN1(\u_a23_mem/n21126 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21128 ) );
  MUX \u_a23_mem/U21184  ( .IN0(o[44]), .IN1(o[172]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21127 ) );
  MUX \u_a23_mem/U21183  ( .IN0(o[108]), .IN1(o[236]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21126 ) );
  MUX \u_a23_mem/U21182  ( .IN0(\u_a23_mem/n21124 ), .IN1(\u_a23_mem/n21121 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21125 ) );
  MUX \u_a23_mem/U21181  ( .IN0(\u_a23_mem/n21123 ), .IN1(\u_a23_mem/n21122 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21124 ) );
  MUX \u_a23_mem/U21180  ( .IN0(o[28]), .IN1(o[156]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21123 ) );
  MUX \u_a23_mem/U21179  ( .IN0(o[92]), .IN1(o[220]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21122 ) );
  MUX \u_a23_mem/U21178  ( .IN0(\u_a23_mem/n21120 ), .IN1(\u_a23_mem/n21119 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21121 ) );
  MUX \u_a23_mem/U21177  ( .IN0(o[60]), .IN1(o[188]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21120 ) );
  MUX \u_a23_mem/U21176  ( .IN0(o[124]), .IN1(o[252]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21119 ) );
  MUX \u_a23_mem/U21174  ( .IN0(\u_a23_mem/n21116 ), .IN1(\u_a23_mem/n21113 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21117 ) );
  MUX \u_a23_mem/U21173  ( .IN0(\u_a23_mem/n21115 ), .IN1(\u_a23_mem/n21114 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21116 ) );
  MUX \u_a23_mem/U21172  ( .IN0(o[20]), .IN1(o[148]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21115 ) );
  MUX \u_a23_mem/U21171  ( .IN0(o[84]), .IN1(o[212]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21114 ) );
  MUX \u_a23_mem/U21170  ( .IN0(\u_a23_mem/n21112 ), .IN1(\u_a23_mem/n21111 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21113 ) );
  MUX \u_a23_mem/U21169  ( .IN0(o[52]), .IN1(o[180]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21112 ) );
  MUX \u_a23_mem/U21168  ( .IN0(o[116]), .IN1(o[244]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21111 ) );
  MUX \u_a23_mem/U21159  ( .IN0(\u_a23_mem/n21102 ), .IN1(\u_a23_mem/n21099 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21103 ) );
  MUX \u_a23_mem/U21158  ( .IN0(\u_a23_mem/n21101 ), .IN1(\u_a23_mem/n21100 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21102 ) );
  MUX \u_a23_mem/U21157  ( .IN0(o[11]), .IN1(o[139]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21101 ) );
  MUX \u_a23_mem/U21156  ( .IN0(o[75]), .IN1(o[203]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21100 ) );
  MUX \u_a23_mem/U21155  ( .IN0(\u_a23_mem/n21098 ), .IN1(\u_a23_mem/n21097 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21099 ) );
  MUX \u_a23_mem/U21154  ( .IN0(o[43]), .IN1(o[171]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21098 ) );
  MUX \u_a23_mem/U21153  ( .IN0(o[107]), .IN1(o[235]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21097 ) );
  MUX \u_a23_mem/U21152  ( .IN0(\u_a23_mem/n21095 ), .IN1(\u_a23_mem/n21092 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21096 ) );
  MUX \u_a23_mem/U21151  ( .IN0(\u_a23_mem/n21094 ), .IN1(\u_a23_mem/n21093 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21095 ) );
  MUX \u_a23_mem/U21150  ( .IN0(o[27]), .IN1(o[155]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21094 ) );
  MUX \u_a23_mem/U21149  ( .IN0(o[91]), .IN1(o[219]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21093 ) );
  MUX \u_a23_mem/U21148  ( .IN0(\u_a23_mem/n21091 ), .IN1(\u_a23_mem/n21090 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21092 ) );
  MUX \u_a23_mem/U21147  ( .IN0(o[59]), .IN1(o[187]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21091 ) );
  MUX \u_a23_mem/U21146  ( .IN0(o[123]), .IN1(o[251]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21090 ) );
  MUX \u_a23_mem/U21144  ( .IN0(\u_a23_mem/n21087 ), .IN1(\u_a23_mem/n21084 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21088 ) );
  MUX \u_a23_mem/U21143  ( .IN0(\u_a23_mem/n21086 ), .IN1(\u_a23_mem/n21085 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21087 ) );
  MUX \u_a23_mem/U21142  ( .IN0(o[19]), .IN1(o[147]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21086 ) );
  MUX \u_a23_mem/U21141  ( .IN0(o[83]), .IN1(o[211]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21085 ) );
  MUX \u_a23_mem/U21140  ( .IN0(\u_a23_mem/n21083 ), .IN1(\u_a23_mem/n21082 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21084 ) );
  MUX \u_a23_mem/U21139  ( .IN0(o[51]), .IN1(o[179]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21083 ) );
  MUX \u_a23_mem/U21138  ( .IN0(o[115]), .IN1(o[243]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21082 ) );
  MUX \u_a23_mem/U21129  ( .IN0(\u_a23_mem/n21073 ), .IN1(\u_a23_mem/n21070 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21074 ) );
  MUX \u_a23_mem/U21128  ( .IN0(\u_a23_mem/n21072 ), .IN1(\u_a23_mem/n21071 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21073 ) );
  MUX \u_a23_mem/U21127  ( .IN0(o[10]), .IN1(o[138]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21072 ) );
  MUX \u_a23_mem/U21126  ( .IN0(o[74]), .IN1(o[202]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21071 ) );
  MUX \u_a23_mem/U21125  ( .IN0(\u_a23_mem/n21069 ), .IN1(\u_a23_mem/n21068 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21070 ) );
  MUX \u_a23_mem/U21124  ( .IN0(o[42]), .IN1(o[170]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21069 ) );
  MUX \u_a23_mem/U21123  ( .IN0(o[106]), .IN1(o[234]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21068 ) );
  MUX \u_a23_mem/U21122  ( .IN0(\u_a23_mem/n21066 ), .IN1(\u_a23_mem/n21063 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21067 ) );
  MUX \u_a23_mem/U21121  ( .IN0(\u_a23_mem/n21065 ), .IN1(\u_a23_mem/n21064 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21066 ) );
  MUX \u_a23_mem/U21120  ( .IN0(o[26]), .IN1(o[154]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21065 ) );
  MUX \u_a23_mem/U21119  ( .IN0(o[90]), .IN1(o[218]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21064 ) );
  MUX \u_a23_mem/U21118  ( .IN0(\u_a23_mem/n21062 ), .IN1(\u_a23_mem/n21061 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21063 ) );
  MUX \u_a23_mem/U21117  ( .IN0(o[58]), .IN1(o[186]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21062 ) );
  MUX \u_a23_mem/U21116  ( .IN0(o[122]), .IN1(o[250]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21061 ) );
  MUX \u_a23_mem/U21114  ( .IN0(\u_a23_mem/n21058 ), .IN1(\u_a23_mem/n21055 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21059 ) );
  MUX \u_a23_mem/U21113  ( .IN0(\u_a23_mem/n21057 ), .IN1(\u_a23_mem/n21056 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21058 ) );
  MUX \u_a23_mem/U21112  ( .IN0(o[18]), .IN1(o[146]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21057 ) );
  MUX \u_a23_mem/U21111  ( .IN0(o[82]), .IN1(o[210]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21056 ) );
  MUX \u_a23_mem/U21110  ( .IN0(\u_a23_mem/n21054 ), .IN1(\u_a23_mem/n21053 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21055 ) );
  MUX \u_a23_mem/U21109  ( .IN0(o[50]), .IN1(o[178]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21054 ) );
  MUX \u_a23_mem/U21108  ( .IN0(o[114]), .IN1(o[242]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21053 ) );
  MUX \u_a23_mem/U21099  ( .IN0(\u_a23_mem/n21044 ), .IN1(\u_a23_mem/n21041 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21045 ) );
  MUX \u_a23_mem/U21098  ( .IN0(\u_a23_mem/n21043 ), .IN1(\u_a23_mem/n21042 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21044 ) );
  MUX \u_a23_mem/U21097  ( .IN0(o[9]), .IN1(o[137]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21043 ) );
  MUX \u_a23_mem/U21096  ( .IN0(o[73]), .IN1(o[201]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21042 ) );
  MUX \u_a23_mem/U21095  ( .IN0(\u_a23_mem/n21040 ), .IN1(\u_a23_mem/n21039 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21041 ) );
  MUX \u_a23_mem/U21094  ( .IN0(o[41]), .IN1(o[169]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21040 ) );
  MUX \u_a23_mem/U21093  ( .IN0(o[105]), .IN1(o[233]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21039 ) );
  MUX \u_a23_mem/U21092  ( .IN0(\u_a23_mem/n21037 ), .IN1(\u_a23_mem/n21034 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21038 ) );
  MUX \u_a23_mem/U21091  ( .IN0(\u_a23_mem/n21036 ), .IN1(\u_a23_mem/n21035 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21037 ) );
  MUX \u_a23_mem/U21090  ( .IN0(o[25]), .IN1(o[153]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21036 ) );
  MUX \u_a23_mem/U21089  ( .IN0(o[89]), .IN1(o[217]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21035 ) );
  MUX \u_a23_mem/U21088  ( .IN0(\u_a23_mem/n21033 ), .IN1(\u_a23_mem/n21032 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21034 ) );
  MUX \u_a23_mem/U21087  ( .IN0(o[57]), .IN1(o[185]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21033 ) );
  MUX \u_a23_mem/U21086  ( .IN0(o[121]), .IN1(o[249]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21032 ) );
  MUX \u_a23_mem/U21084  ( .IN0(\u_a23_mem/n21029 ), .IN1(\u_a23_mem/n21026 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21030 ) );
  MUX \u_a23_mem/U21083  ( .IN0(\u_a23_mem/n21028 ), .IN1(\u_a23_mem/n21027 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21029 ) );
  MUX \u_a23_mem/U21082  ( .IN0(o[17]), .IN1(o[145]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21028 ) );
  MUX \u_a23_mem/U21081  ( .IN0(o[81]), .IN1(o[209]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21027 ) );
  MUX \u_a23_mem/U21080  ( .IN0(\u_a23_mem/n21025 ), .IN1(\u_a23_mem/n21024 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21026 ) );
  MUX \u_a23_mem/U21079  ( .IN0(o[49]), .IN1(o[177]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21025 ) );
  MUX \u_a23_mem/U21078  ( .IN0(o[113]), .IN1(o[241]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21024 ) );
  MUX \u_a23_mem/U21069  ( .IN0(\u_a23_mem/n21015 ), .IN1(\u_a23_mem/n21012 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21016 ) );
  MUX \u_a23_mem/U21068  ( .IN0(\u_a23_mem/n21014 ), .IN1(\u_a23_mem/n21013 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21015 ) );
  MUX \u_a23_mem/U21067  ( .IN0(o[8]), .IN1(o[136]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21014 ) );
  MUX \u_a23_mem/U21066  ( .IN0(o[72]), .IN1(o[200]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21013 ) );
  MUX \u_a23_mem/U21065  ( .IN0(\u_a23_mem/n21011 ), .IN1(\u_a23_mem/n21010 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21012 ) );
  MUX \u_a23_mem/U21064  ( .IN0(o[40]), .IN1(o[168]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21011 ) );
  MUX \u_a23_mem/U21063  ( .IN0(o[104]), .IN1(o[232]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21010 ) );
  MUX \u_a23_mem/U21062  ( .IN0(\u_a23_mem/n21008 ), .IN1(\u_a23_mem/n21005 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21009 ) );
  MUX \u_a23_mem/U21061  ( .IN0(\u_a23_mem/n21007 ), .IN1(\u_a23_mem/n21006 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21008 ) );
  MUX \u_a23_mem/U21060  ( .IN0(o[24]), .IN1(o[152]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21007 ) );
  MUX \u_a23_mem/U21059  ( .IN0(o[88]), .IN1(o[216]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21006 ) );
  MUX \u_a23_mem/U21058  ( .IN0(\u_a23_mem/n21004 ), .IN1(\u_a23_mem/n21003 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21005 ) );
  MUX \u_a23_mem/U21057  ( .IN0(o[56]), .IN1(o[184]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21004 ) );
  MUX \u_a23_mem/U21056  ( .IN0(o[120]), .IN1(o[248]), .SEL(m_address[4]), .F(
        \u_a23_mem/n21003 ) );
  MUX \u_a23_mem/U21054  ( .IN0(\u_a23_mem/n21000 ), .IN1(\u_a23_mem/n20997 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n21001 ) );
  MUX \u_a23_mem/U21053  ( .IN0(\u_a23_mem/n20999 ), .IN1(\u_a23_mem/n20998 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n21000 ) );
  MUX \u_a23_mem/U21052  ( .IN0(o[16]), .IN1(o[144]), .SEL(m_address[4]), .F(
        \u_a23_mem/n20999 ) );
  MUX \u_a23_mem/U21051  ( .IN0(o[80]), .IN1(o[208]), .SEL(m_address[4]), .F(
        \u_a23_mem/n20998 ) );
  MUX \u_a23_mem/U21050  ( .IN0(\u_a23_mem/n20996 ), .IN1(\u_a23_mem/n20995 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20997 ) );
  MUX \u_a23_mem/U21049  ( .IN0(o[48]), .IN1(o[176]), .SEL(m_address[4]), .F(
        \u_a23_mem/n20996 ) );
  MUX \u_a23_mem/U21048  ( .IN0(o[112]), .IN1(o[240]), .SEL(m_address[4]), .F(
        \u_a23_mem/n20995 ) );
  MUX \u_a23_mem/U20999  ( .IN0(\u_a23_mem/n20962 ), .IN1(\u_a23_mem/n20959 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20963 ) );
  MUX \u_a23_mem/U20998  ( .IN0(\u_a23_mem/n20961 ), .IN1(\u_a23_mem/n20960 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20962 ) );
  MUX \u_a23_mem/U20997  ( .IN0(\u_a23_mem/stack_mem[1][7] ), .IN1(
        \u_a23_mem/stack_mem[17][7] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20961 ) );
  MUX \u_a23_mem/U20996  ( .IN0(\u_a23_mem/stack_mem[9][7] ), .IN1(
        \u_a23_mem/stack_mem[25][7] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20960 ) );
  MUX \u_a23_mem/U20995  ( .IN0(\u_a23_mem/n20958 ), .IN1(\u_a23_mem/n20957 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20959 ) );
  MUX \u_a23_mem/U20994  ( .IN0(\u_a23_mem/stack_mem[5][7] ), .IN1(
        \u_a23_mem/stack_mem[21][7] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20958 ) );
  MUX \u_a23_mem/U20993  ( .IN0(\u_a23_mem/stack_mem[13][7] ), .IN1(
        \u_a23_mem/stack_mem[29][7] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20957 ) );
  MUX \u_a23_mem/U20992  ( .IN0(\u_a23_mem/n20955 ), .IN1(\u_a23_mem/n20952 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20956 ) );
  MUX \u_a23_mem/U20991  ( .IN0(\u_a23_mem/n20954 ), .IN1(\u_a23_mem/n20953 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20955 ) );
  MUX \u_a23_mem/U20990  ( .IN0(\u_a23_mem/stack_mem[3][7] ), .IN1(
        \u_a23_mem/stack_mem[19][7] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20954 ) );
  MUX \u_a23_mem/U20989  ( .IN0(\u_a23_mem/stack_mem[11][7] ), .IN1(
        \u_a23_mem/stack_mem[27][7] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20953 ) );
  MUX \u_a23_mem/U20988  ( .IN0(\u_a23_mem/n20951 ), .IN1(\u_a23_mem/n20950 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20952 ) );
  MUX \u_a23_mem/U20987  ( .IN0(\u_a23_mem/stack_mem[7][7] ), .IN1(
        \u_a23_mem/stack_mem[23][7] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20951 ) );
  MUX \u_a23_mem/U20986  ( .IN0(\u_a23_mem/stack_mem[15][7] ), .IN1(
        \u_a23_mem/stack_mem[31][7] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20950 ) );
  MUX \u_a23_mem/U20984  ( .IN0(\u_a23_mem/n20947 ), .IN1(\u_a23_mem/n20944 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20948 ) );
  MUX \u_a23_mem/U20983  ( .IN0(\u_a23_mem/n20946 ), .IN1(\u_a23_mem/n20945 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20947 ) );
  MUX \u_a23_mem/U20982  ( .IN0(\u_a23_mem/stack_mem[2][7] ), .IN1(
        \u_a23_mem/stack_mem[18][7] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20946 ) );
  MUX \u_a23_mem/U20981  ( .IN0(\u_a23_mem/stack_mem[10][7] ), .IN1(
        \u_a23_mem/stack_mem[26][7] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20945 ) );
  MUX \u_a23_mem/U20980  ( .IN0(\u_a23_mem/n20943 ), .IN1(\u_a23_mem/n20942 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20944 ) );
  MUX \u_a23_mem/U20979  ( .IN0(\u_a23_mem/stack_mem[6][7] ), .IN1(
        \u_a23_mem/stack_mem[22][7] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20943 ) );
  MUX \u_a23_mem/U20978  ( .IN0(\u_a23_mem/stack_mem[14][7] ), .IN1(
        \u_a23_mem/stack_mem[30][7] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20942 ) );
  MUX \u_a23_mem/U20969  ( .IN0(\u_a23_mem/n20933 ), .IN1(\u_a23_mem/n20930 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20934 ) );
  MUX \u_a23_mem/U20968  ( .IN0(\u_a23_mem/n20932 ), .IN1(\u_a23_mem/n20931 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20933 ) );
  MUX \u_a23_mem/U20967  ( .IN0(\u_a23_mem/stack_mem[1][6] ), .IN1(
        \u_a23_mem/stack_mem[17][6] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20932 ) );
  MUX \u_a23_mem/U20966  ( .IN0(\u_a23_mem/stack_mem[9][6] ), .IN1(
        \u_a23_mem/stack_mem[25][6] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20931 ) );
  MUX \u_a23_mem/U20965  ( .IN0(\u_a23_mem/n20929 ), .IN1(\u_a23_mem/n20928 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20930 ) );
  MUX \u_a23_mem/U20964  ( .IN0(\u_a23_mem/stack_mem[5][6] ), .IN1(
        \u_a23_mem/stack_mem[21][6] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20929 ) );
  MUX \u_a23_mem/U20963  ( .IN0(\u_a23_mem/stack_mem[13][6] ), .IN1(
        \u_a23_mem/stack_mem[29][6] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20928 ) );
  MUX \u_a23_mem/U20962  ( .IN0(\u_a23_mem/n20926 ), .IN1(\u_a23_mem/n20923 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20927 ) );
  MUX \u_a23_mem/U20961  ( .IN0(\u_a23_mem/n20925 ), .IN1(\u_a23_mem/n20924 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20926 ) );
  MUX \u_a23_mem/U20960  ( .IN0(\u_a23_mem/stack_mem[3][6] ), .IN1(
        \u_a23_mem/stack_mem[19][6] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20925 ) );
  MUX \u_a23_mem/U20959  ( .IN0(\u_a23_mem/stack_mem[11][6] ), .IN1(
        \u_a23_mem/stack_mem[27][6] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20924 ) );
  MUX \u_a23_mem/U20958  ( .IN0(\u_a23_mem/n20922 ), .IN1(\u_a23_mem/n20921 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20923 ) );
  MUX \u_a23_mem/U20957  ( .IN0(\u_a23_mem/stack_mem[7][6] ), .IN1(
        \u_a23_mem/stack_mem[23][6] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20922 ) );
  MUX \u_a23_mem/U20956  ( .IN0(\u_a23_mem/stack_mem[15][6] ), .IN1(
        \u_a23_mem/stack_mem[31][6] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20921 ) );
  MUX \u_a23_mem/U20954  ( .IN0(\u_a23_mem/n20918 ), .IN1(\u_a23_mem/n20915 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20919 ) );
  MUX \u_a23_mem/U20953  ( .IN0(\u_a23_mem/n20917 ), .IN1(\u_a23_mem/n20916 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20918 ) );
  MUX \u_a23_mem/U20952  ( .IN0(\u_a23_mem/stack_mem[2][6] ), .IN1(
        \u_a23_mem/stack_mem[18][6] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20917 ) );
  MUX \u_a23_mem/U20951  ( .IN0(\u_a23_mem/stack_mem[10][6] ), .IN1(
        \u_a23_mem/stack_mem[26][6] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20916 ) );
  MUX \u_a23_mem/U20950  ( .IN0(\u_a23_mem/n20914 ), .IN1(\u_a23_mem/n20913 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20915 ) );
  MUX \u_a23_mem/U20949  ( .IN0(\u_a23_mem/stack_mem[6][6] ), .IN1(
        \u_a23_mem/stack_mem[22][6] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20914 ) );
  MUX \u_a23_mem/U20948  ( .IN0(\u_a23_mem/stack_mem[14][6] ), .IN1(
        \u_a23_mem/stack_mem[30][6] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20913 ) );
  MUX \u_a23_mem/U20939  ( .IN0(\u_a23_mem/n20904 ), .IN1(\u_a23_mem/n20901 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20905 ) );
  MUX \u_a23_mem/U20938  ( .IN0(\u_a23_mem/n20903 ), .IN1(\u_a23_mem/n20902 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20904 ) );
  MUX \u_a23_mem/U20937  ( .IN0(\u_a23_mem/stack_mem[1][5] ), .IN1(
        \u_a23_mem/stack_mem[17][5] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20903 ) );
  MUX \u_a23_mem/U20936  ( .IN0(\u_a23_mem/stack_mem[9][5] ), .IN1(
        \u_a23_mem/stack_mem[25][5] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20902 ) );
  MUX \u_a23_mem/U20935  ( .IN0(\u_a23_mem/n20900 ), .IN1(\u_a23_mem/n20899 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20901 ) );
  MUX \u_a23_mem/U20934  ( .IN0(\u_a23_mem/stack_mem[5][5] ), .IN1(
        \u_a23_mem/stack_mem[21][5] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20900 ) );
  MUX \u_a23_mem/U20933  ( .IN0(\u_a23_mem/stack_mem[13][5] ), .IN1(
        \u_a23_mem/stack_mem[29][5] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20899 ) );
  MUX \u_a23_mem/U20932  ( .IN0(\u_a23_mem/n20897 ), .IN1(\u_a23_mem/n20894 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20898 ) );
  MUX \u_a23_mem/U20931  ( .IN0(\u_a23_mem/n20896 ), .IN1(\u_a23_mem/n20895 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20897 ) );
  MUX \u_a23_mem/U20930  ( .IN0(\u_a23_mem/stack_mem[3][5] ), .IN1(
        \u_a23_mem/stack_mem[19][5] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20896 ) );
  MUX \u_a23_mem/U20929  ( .IN0(\u_a23_mem/stack_mem[11][5] ), .IN1(
        \u_a23_mem/stack_mem[27][5] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20895 ) );
  MUX \u_a23_mem/U20928  ( .IN0(\u_a23_mem/n20893 ), .IN1(\u_a23_mem/n20892 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20894 ) );
  MUX \u_a23_mem/U20927  ( .IN0(\u_a23_mem/stack_mem[7][5] ), .IN1(
        \u_a23_mem/stack_mem[23][5] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20893 ) );
  MUX \u_a23_mem/U20926  ( .IN0(\u_a23_mem/stack_mem[15][5] ), .IN1(
        \u_a23_mem/stack_mem[31][5] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20892 ) );
  MUX \u_a23_mem/U20924  ( .IN0(\u_a23_mem/n20889 ), .IN1(\u_a23_mem/n20886 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20890 ) );
  MUX \u_a23_mem/U20923  ( .IN0(\u_a23_mem/n20888 ), .IN1(\u_a23_mem/n20887 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20889 ) );
  MUX \u_a23_mem/U20922  ( .IN0(\u_a23_mem/stack_mem[2][5] ), .IN1(
        \u_a23_mem/stack_mem[18][5] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20888 ) );
  MUX \u_a23_mem/U20921  ( .IN0(\u_a23_mem/stack_mem[10][5] ), .IN1(
        \u_a23_mem/stack_mem[26][5] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20887 ) );
  MUX \u_a23_mem/U20920  ( .IN0(\u_a23_mem/n20885 ), .IN1(\u_a23_mem/n20884 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20886 ) );
  MUX \u_a23_mem/U20919  ( .IN0(\u_a23_mem/stack_mem[6][5] ), .IN1(
        \u_a23_mem/stack_mem[22][5] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20885 ) );
  MUX \u_a23_mem/U20918  ( .IN0(\u_a23_mem/stack_mem[14][5] ), .IN1(
        \u_a23_mem/stack_mem[30][5] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20884 ) );
  MUX \u_a23_mem/U20909  ( .IN0(\u_a23_mem/n20875 ), .IN1(\u_a23_mem/n20872 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20876 ) );
  MUX \u_a23_mem/U20908  ( .IN0(\u_a23_mem/n20874 ), .IN1(\u_a23_mem/n20873 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20875 ) );
  MUX \u_a23_mem/U20907  ( .IN0(\u_a23_mem/stack_mem[1][4] ), .IN1(
        \u_a23_mem/stack_mem[17][4] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20874 ) );
  MUX \u_a23_mem/U20906  ( .IN0(\u_a23_mem/stack_mem[9][4] ), .IN1(
        \u_a23_mem/stack_mem[25][4] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20873 ) );
  MUX \u_a23_mem/U20905  ( .IN0(\u_a23_mem/n20871 ), .IN1(\u_a23_mem/n20870 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20872 ) );
  MUX \u_a23_mem/U20904  ( .IN0(\u_a23_mem/stack_mem[5][4] ), .IN1(
        \u_a23_mem/stack_mem[21][4] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20871 ) );
  MUX \u_a23_mem/U20903  ( .IN0(\u_a23_mem/stack_mem[13][4] ), .IN1(
        \u_a23_mem/stack_mem[29][4] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20870 ) );
  MUX \u_a23_mem/U20902  ( .IN0(\u_a23_mem/n20868 ), .IN1(\u_a23_mem/n20865 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20869 ) );
  MUX \u_a23_mem/U20901  ( .IN0(\u_a23_mem/n20867 ), .IN1(\u_a23_mem/n20866 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20868 ) );
  MUX \u_a23_mem/U20900  ( .IN0(\u_a23_mem/stack_mem[3][4] ), .IN1(
        \u_a23_mem/stack_mem[19][4] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20867 ) );
  MUX \u_a23_mem/U20899  ( .IN0(\u_a23_mem/stack_mem[11][4] ), .IN1(
        \u_a23_mem/stack_mem[27][4] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20866 ) );
  MUX \u_a23_mem/U20898  ( .IN0(\u_a23_mem/n20864 ), .IN1(\u_a23_mem/n20863 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20865 ) );
  MUX \u_a23_mem/U20897  ( .IN0(\u_a23_mem/stack_mem[7][4] ), .IN1(
        \u_a23_mem/stack_mem[23][4] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20864 ) );
  MUX \u_a23_mem/U20896  ( .IN0(\u_a23_mem/stack_mem[15][4] ), .IN1(
        \u_a23_mem/stack_mem[31][4] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20863 ) );
  MUX \u_a23_mem/U20894  ( .IN0(\u_a23_mem/n20860 ), .IN1(\u_a23_mem/n20857 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20861 ) );
  MUX \u_a23_mem/U20893  ( .IN0(\u_a23_mem/n20859 ), .IN1(\u_a23_mem/n20858 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20860 ) );
  MUX \u_a23_mem/U20892  ( .IN0(\u_a23_mem/stack_mem[2][4] ), .IN1(
        \u_a23_mem/stack_mem[18][4] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20859 ) );
  MUX \u_a23_mem/U20891  ( .IN0(\u_a23_mem/stack_mem[10][4] ), .IN1(
        \u_a23_mem/stack_mem[26][4] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20858 ) );
  MUX \u_a23_mem/U20890  ( .IN0(\u_a23_mem/n20856 ), .IN1(\u_a23_mem/n20855 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20857 ) );
  MUX \u_a23_mem/U20889  ( .IN0(\u_a23_mem/stack_mem[6][4] ), .IN1(
        \u_a23_mem/stack_mem[22][4] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20856 ) );
  MUX \u_a23_mem/U20888  ( .IN0(\u_a23_mem/stack_mem[14][4] ), .IN1(
        \u_a23_mem/stack_mem[30][4] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20855 ) );
  MUX \u_a23_mem/U20879  ( .IN0(\u_a23_mem/n20846 ), .IN1(\u_a23_mem/n20843 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20847 ) );
  MUX \u_a23_mem/U20878  ( .IN0(\u_a23_mem/n20845 ), .IN1(\u_a23_mem/n20844 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20846 ) );
  MUX \u_a23_mem/U20877  ( .IN0(\u_a23_mem/stack_mem[1][3] ), .IN1(
        \u_a23_mem/stack_mem[17][3] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20845 ) );
  MUX \u_a23_mem/U20876  ( .IN0(\u_a23_mem/stack_mem[9][3] ), .IN1(
        \u_a23_mem/stack_mem[25][3] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20844 ) );
  MUX \u_a23_mem/U20875  ( .IN0(\u_a23_mem/n20842 ), .IN1(\u_a23_mem/n20841 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20843 ) );
  MUX \u_a23_mem/U20874  ( .IN0(\u_a23_mem/stack_mem[5][3] ), .IN1(
        \u_a23_mem/stack_mem[21][3] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20842 ) );
  MUX \u_a23_mem/U20873  ( .IN0(\u_a23_mem/stack_mem[13][3] ), .IN1(
        \u_a23_mem/stack_mem[29][3] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20841 ) );
  MUX \u_a23_mem/U20872  ( .IN0(\u_a23_mem/n20839 ), .IN1(\u_a23_mem/n20836 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20840 ) );
  MUX \u_a23_mem/U20871  ( .IN0(\u_a23_mem/n20838 ), .IN1(\u_a23_mem/n20837 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20839 ) );
  MUX \u_a23_mem/U20870  ( .IN0(\u_a23_mem/stack_mem[3][3] ), .IN1(
        \u_a23_mem/stack_mem[19][3] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20838 ) );
  MUX \u_a23_mem/U20869  ( .IN0(\u_a23_mem/stack_mem[11][3] ), .IN1(
        \u_a23_mem/stack_mem[27][3] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20837 ) );
  MUX \u_a23_mem/U20868  ( .IN0(\u_a23_mem/n20835 ), .IN1(\u_a23_mem/n20834 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20836 ) );
  MUX \u_a23_mem/U20867  ( .IN0(\u_a23_mem/stack_mem[7][3] ), .IN1(
        \u_a23_mem/stack_mem[23][3] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20835 ) );
  MUX \u_a23_mem/U20866  ( .IN0(\u_a23_mem/stack_mem[15][3] ), .IN1(
        \u_a23_mem/stack_mem[31][3] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20834 ) );
  MUX \u_a23_mem/U20864  ( .IN0(\u_a23_mem/n20831 ), .IN1(\u_a23_mem/n20828 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20832 ) );
  MUX \u_a23_mem/U20863  ( .IN0(\u_a23_mem/n20830 ), .IN1(\u_a23_mem/n20829 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20831 ) );
  MUX \u_a23_mem/U20862  ( .IN0(\u_a23_mem/stack_mem[2][3] ), .IN1(
        \u_a23_mem/stack_mem[18][3] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20830 ) );
  MUX \u_a23_mem/U20861  ( .IN0(\u_a23_mem/stack_mem[10][3] ), .IN1(
        \u_a23_mem/stack_mem[26][3] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20829 ) );
  MUX \u_a23_mem/U20860  ( .IN0(\u_a23_mem/n20827 ), .IN1(\u_a23_mem/n20826 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20828 ) );
  MUX \u_a23_mem/U20859  ( .IN0(\u_a23_mem/stack_mem[6][3] ), .IN1(
        \u_a23_mem/stack_mem[22][3] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20827 ) );
  MUX \u_a23_mem/U20858  ( .IN0(\u_a23_mem/stack_mem[14][3] ), .IN1(
        \u_a23_mem/stack_mem[30][3] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20826 ) );
  MUX \u_a23_mem/U20849  ( .IN0(\u_a23_mem/n20817 ), .IN1(\u_a23_mem/n20814 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20818 ) );
  MUX \u_a23_mem/U20848  ( .IN0(\u_a23_mem/n20816 ), .IN1(\u_a23_mem/n20815 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20817 ) );
  MUX \u_a23_mem/U20847  ( .IN0(\u_a23_mem/stack_mem[1][2] ), .IN1(
        \u_a23_mem/stack_mem[17][2] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20816 ) );
  MUX \u_a23_mem/U20846  ( .IN0(\u_a23_mem/stack_mem[9][2] ), .IN1(
        \u_a23_mem/stack_mem[25][2] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20815 ) );
  MUX \u_a23_mem/U20845  ( .IN0(\u_a23_mem/n20813 ), .IN1(\u_a23_mem/n20812 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20814 ) );
  MUX \u_a23_mem/U20844  ( .IN0(\u_a23_mem/stack_mem[5][2] ), .IN1(
        \u_a23_mem/stack_mem[21][2] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20813 ) );
  MUX \u_a23_mem/U20843  ( .IN0(\u_a23_mem/stack_mem[13][2] ), .IN1(
        \u_a23_mem/stack_mem[29][2] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20812 ) );
  MUX \u_a23_mem/U20842  ( .IN0(\u_a23_mem/n20810 ), .IN1(\u_a23_mem/n20807 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20811 ) );
  MUX \u_a23_mem/U20841  ( .IN0(\u_a23_mem/n20809 ), .IN1(\u_a23_mem/n20808 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20810 ) );
  MUX \u_a23_mem/U20840  ( .IN0(\u_a23_mem/stack_mem[3][2] ), .IN1(
        \u_a23_mem/stack_mem[19][2] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20809 ) );
  MUX \u_a23_mem/U20839  ( .IN0(\u_a23_mem/stack_mem[11][2] ), .IN1(
        \u_a23_mem/stack_mem[27][2] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20808 ) );
  MUX \u_a23_mem/U20838  ( .IN0(\u_a23_mem/n20806 ), .IN1(\u_a23_mem/n20805 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20807 ) );
  MUX \u_a23_mem/U20837  ( .IN0(\u_a23_mem/stack_mem[7][2] ), .IN1(
        \u_a23_mem/stack_mem[23][2] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20806 ) );
  MUX \u_a23_mem/U20836  ( .IN0(\u_a23_mem/stack_mem[15][2] ), .IN1(
        \u_a23_mem/stack_mem[31][2] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20805 ) );
  MUX \u_a23_mem/U20834  ( .IN0(\u_a23_mem/n20802 ), .IN1(\u_a23_mem/n20799 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20803 ) );
  MUX \u_a23_mem/U20833  ( .IN0(\u_a23_mem/n20801 ), .IN1(\u_a23_mem/n20800 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20802 ) );
  MUX \u_a23_mem/U20832  ( .IN0(\u_a23_mem/stack_mem[2][2] ), .IN1(
        \u_a23_mem/stack_mem[18][2] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20801 ) );
  MUX \u_a23_mem/U20831  ( .IN0(\u_a23_mem/stack_mem[10][2] ), .IN1(
        \u_a23_mem/stack_mem[26][2] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20800 ) );
  MUX \u_a23_mem/U20830  ( .IN0(\u_a23_mem/n20798 ), .IN1(\u_a23_mem/n20797 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20799 ) );
  MUX \u_a23_mem/U20829  ( .IN0(\u_a23_mem/stack_mem[6][2] ), .IN1(
        \u_a23_mem/stack_mem[22][2] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20798 ) );
  MUX \u_a23_mem/U20828  ( .IN0(\u_a23_mem/stack_mem[14][2] ), .IN1(
        \u_a23_mem/stack_mem[30][2] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20797 ) );
  MUX \u_a23_mem/U20819  ( .IN0(\u_a23_mem/n20788 ), .IN1(\u_a23_mem/n20785 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20789 ) );
  MUX \u_a23_mem/U20818  ( .IN0(\u_a23_mem/n20787 ), .IN1(\u_a23_mem/n20786 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20788 ) );
  MUX \u_a23_mem/U20817  ( .IN0(\u_a23_mem/stack_mem[1][1] ), .IN1(
        \u_a23_mem/stack_mem[17][1] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20787 ) );
  MUX \u_a23_mem/U20816  ( .IN0(\u_a23_mem/stack_mem[9][1] ), .IN1(
        \u_a23_mem/stack_mem[25][1] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20786 ) );
  MUX \u_a23_mem/U20815  ( .IN0(\u_a23_mem/n20784 ), .IN1(\u_a23_mem/n20783 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20785 ) );
  MUX \u_a23_mem/U20814  ( .IN0(\u_a23_mem/stack_mem[5][1] ), .IN1(
        \u_a23_mem/stack_mem[21][1] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20784 ) );
  MUX \u_a23_mem/U20813  ( .IN0(\u_a23_mem/stack_mem[13][1] ), .IN1(
        \u_a23_mem/stack_mem[29][1] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20783 ) );
  MUX \u_a23_mem/U20812  ( .IN0(\u_a23_mem/n20781 ), .IN1(\u_a23_mem/n20778 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20782 ) );
  MUX \u_a23_mem/U20811  ( .IN0(\u_a23_mem/n20780 ), .IN1(\u_a23_mem/n20779 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20781 ) );
  MUX \u_a23_mem/U20810  ( .IN0(\u_a23_mem/stack_mem[3][1] ), .IN1(
        \u_a23_mem/stack_mem[19][1] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20780 ) );
  MUX \u_a23_mem/U20809  ( .IN0(\u_a23_mem/stack_mem[11][1] ), .IN1(
        \u_a23_mem/stack_mem[27][1] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20779 ) );
  MUX \u_a23_mem/U20808  ( .IN0(\u_a23_mem/n20777 ), .IN1(\u_a23_mem/n20776 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20778 ) );
  MUX \u_a23_mem/U20807  ( .IN0(\u_a23_mem/stack_mem[7][1] ), .IN1(
        \u_a23_mem/stack_mem[23][1] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20777 ) );
  MUX \u_a23_mem/U20806  ( .IN0(\u_a23_mem/stack_mem[15][1] ), .IN1(
        \u_a23_mem/stack_mem[31][1] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20776 ) );
  MUX \u_a23_mem/U20804  ( .IN0(\u_a23_mem/n20773 ), .IN1(\u_a23_mem/n20770 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20774 ) );
  MUX \u_a23_mem/U20803  ( .IN0(\u_a23_mem/n20772 ), .IN1(\u_a23_mem/n20771 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20773 ) );
  MUX \u_a23_mem/U20802  ( .IN0(\u_a23_mem/stack_mem[2][1] ), .IN1(
        \u_a23_mem/stack_mem[18][1] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20772 ) );
  MUX \u_a23_mem/U20801  ( .IN0(\u_a23_mem/stack_mem[10][1] ), .IN1(
        \u_a23_mem/stack_mem[26][1] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20771 ) );
  MUX \u_a23_mem/U20800  ( .IN0(\u_a23_mem/n20769 ), .IN1(\u_a23_mem/n20768 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20770 ) );
  MUX \u_a23_mem/U20799  ( .IN0(\u_a23_mem/stack_mem[6][1] ), .IN1(
        \u_a23_mem/stack_mem[22][1] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20769 ) );
  MUX \u_a23_mem/U20798  ( .IN0(\u_a23_mem/stack_mem[14][1] ), .IN1(
        \u_a23_mem/stack_mem[30][1] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20768 ) );
  MUX \u_a23_mem/U20789  ( .IN0(\u_a23_mem/n20759 ), .IN1(\u_a23_mem/n20756 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20760 ) );
  MUX \u_a23_mem/U20788  ( .IN0(\u_a23_mem/n20758 ), .IN1(\u_a23_mem/n20757 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20759 ) );
  MUX \u_a23_mem/U20787  ( .IN0(\u_a23_mem/stack_mem[1][0] ), .IN1(
        \u_a23_mem/stack_mem[17][0] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20758 ) );
  MUX \u_a23_mem/U20786  ( .IN0(\u_a23_mem/stack_mem[9][0] ), .IN1(
        \u_a23_mem/stack_mem[25][0] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20757 ) );
  MUX \u_a23_mem/U20785  ( .IN0(\u_a23_mem/n20755 ), .IN1(\u_a23_mem/n20754 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20756 ) );
  MUX \u_a23_mem/U20784  ( .IN0(\u_a23_mem/stack_mem[5][0] ), .IN1(
        \u_a23_mem/stack_mem[21][0] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20755 ) );
  MUX \u_a23_mem/U20783  ( .IN0(\u_a23_mem/stack_mem[13][0] ), .IN1(
        \u_a23_mem/stack_mem[29][0] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20754 ) );
  MUX \u_a23_mem/U20782  ( .IN0(\u_a23_mem/n20752 ), .IN1(\u_a23_mem/n20749 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20753 ) );
  MUX \u_a23_mem/U20781  ( .IN0(\u_a23_mem/n20751 ), .IN1(\u_a23_mem/n20750 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20752 ) );
  MUX \u_a23_mem/U20780  ( .IN0(\u_a23_mem/stack_mem[3][0] ), .IN1(
        \u_a23_mem/stack_mem[19][0] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20751 ) );
  MUX \u_a23_mem/U20779  ( .IN0(\u_a23_mem/stack_mem[11][0] ), .IN1(
        \u_a23_mem/stack_mem[27][0] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20750 ) );
  MUX \u_a23_mem/U20778  ( .IN0(\u_a23_mem/n20748 ), .IN1(\u_a23_mem/n20747 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20749 ) );
  MUX \u_a23_mem/U20777  ( .IN0(\u_a23_mem/stack_mem[7][0] ), .IN1(
        \u_a23_mem/stack_mem[23][0] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20748 ) );
  MUX \u_a23_mem/U20776  ( .IN0(\u_a23_mem/stack_mem[15][0] ), .IN1(
        \u_a23_mem/stack_mem[31][0] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20747 ) );
  MUX \u_a23_mem/U20774  ( .IN0(\u_a23_mem/n20744 ), .IN1(\u_a23_mem/n20741 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20745 ) );
  MUX \u_a23_mem/U20773  ( .IN0(\u_a23_mem/n20743 ), .IN1(\u_a23_mem/n20742 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20744 ) );
  MUX \u_a23_mem/U20772  ( .IN0(\u_a23_mem/stack_mem[2][0] ), .IN1(
        \u_a23_mem/stack_mem[18][0] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20743 ) );
  MUX \u_a23_mem/U20771  ( .IN0(\u_a23_mem/stack_mem[10][0] ), .IN1(
        \u_a23_mem/stack_mem[26][0] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20742 ) );
  MUX \u_a23_mem/U20770  ( .IN0(\u_a23_mem/n20740 ), .IN1(\u_a23_mem/n20739 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20741 ) );
  MUX \u_a23_mem/U20769  ( .IN0(\u_a23_mem/stack_mem[6][0] ), .IN1(
        \u_a23_mem/stack_mem[22][0] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20740 ) );
  MUX \u_a23_mem/U20768  ( .IN0(\u_a23_mem/stack_mem[14][0] ), .IN1(
        \u_a23_mem/stack_mem[30][0] ), .SEL(m_address[4]), .F(
        \u_a23_mem/n20739 ) );
  MUX \u_a23_mem/U20663  ( .IN0(\u_a23_mem/n20650 ), .IN1(\u_a23_mem/n20635 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20651 ) );
  MUX \u_a23_mem/U20662  ( .IN0(\u_a23_mem/n20649 ), .IN1(\u_a23_mem/n20642 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20650 ) );
  MUX \u_a23_mem/U20661  ( .IN0(\u_a23_mem/n20648 ), .IN1(\u_a23_mem/n20645 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20649 ) );
  MUX \u_a23_mem/U20660  ( .IN0(\u_a23_mem/n20647 ), .IN1(\u_a23_mem/n20646 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20648 ) );
  MUX \u_a23_mem/U20659  ( .IN0(\u_a23_mem/p_mem[1][7] ), .IN1(
        \u_a23_mem/p_mem[65][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20647 )
         );
  MUX \u_a23_mem/U20658  ( .IN0(\u_a23_mem/p_mem[33][7] ), .IN1(
        \u_a23_mem/p_mem[97][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20646 )
         );
  MUX \u_a23_mem/U20657  ( .IN0(\u_a23_mem/n20644 ), .IN1(\u_a23_mem/n20643 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20645 ) );
  MUX \u_a23_mem/U20656  ( .IN0(\u_a23_mem/p_mem[17][7] ), .IN1(
        \u_a23_mem/p_mem[81][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20644 )
         );
  MUX \u_a23_mem/U20655  ( .IN0(\u_a23_mem/p_mem[49][7] ), .IN1(
        \u_a23_mem/p_mem[113][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20643 )
         );
  MUX \u_a23_mem/U20654  ( .IN0(\u_a23_mem/n20641 ), .IN1(\u_a23_mem/n20638 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20642 ) );
  MUX \u_a23_mem/U20653  ( .IN0(\u_a23_mem/n20640 ), .IN1(\u_a23_mem/n20639 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20641 ) );
  MUX \u_a23_mem/U20652  ( .IN0(\u_a23_mem/p_mem[9][7] ), .IN1(
        \u_a23_mem/p_mem[73][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20640 )
         );
  MUX \u_a23_mem/U20651  ( .IN0(\u_a23_mem/p_mem[41][7] ), .IN1(
        \u_a23_mem/p_mem[105][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20639 )
         );
  MUX \u_a23_mem/U20650  ( .IN0(\u_a23_mem/n20637 ), .IN1(\u_a23_mem/n20636 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20638 ) );
  MUX \u_a23_mem/U20649  ( .IN0(\u_a23_mem/p_mem[25][7] ), .IN1(
        \u_a23_mem/p_mem[89][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20637 )
         );
  MUX \u_a23_mem/U20648  ( .IN0(\u_a23_mem/p_mem[57][7] ), .IN1(
        \u_a23_mem/p_mem[121][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20636 )
         );
  MUX \u_a23_mem/U20647  ( .IN0(\u_a23_mem/n20634 ), .IN1(\u_a23_mem/n20627 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20635 ) );
  MUX \u_a23_mem/U20646  ( .IN0(\u_a23_mem/n20633 ), .IN1(\u_a23_mem/n20630 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20634 ) );
  MUX \u_a23_mem/U20645  ( .IN0(\u_a23_mem/n20632 ), .IN1(\u_a23_mem/n20631 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20633 ) );
  MUX \u_a23_mem/U20644  ( .IN0(\u_a23_mem/p_mem[5][7] ), .IN1(
        \u_a23_mem/p_mem[69][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20632 )
         );
  MUX \u_a23_mem/U20643  ( .IN0(\u_a23_mem/p_mem[37][7] ), .IN1(
        \u_a23_mem/p_mem[101][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20631 )
         );
  MUX \u_a23_mem/U20642  ( .IN0(\u_a23_mem/n20629 ), .IN1(\u_a23_mem/n20628 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20630 ) );
  MUX \u_a23_mem/U20641  ( .IN0(\u_a23_mem/p_mem[21][7] ), .IN1(
        \u_a23_mem/p_mem[85][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20629 )
         );
  MUX \u_a23_mem/U20640  ( .IN0(\u_a23_mem/p_mem[53][7] ), .IN1(
        \u_a23_mem/p_mem[117][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20628 )
         );
  MUX \u_a23_mem/U20639  ( .IN0(\u_a23_mem/n20626 ), .IN1(\u_a23_mem/n20623 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20627 ) );
  MUX \u_a23_mem/U20638  ( .IN0(\u_a23_mem/n20625 ), .IN1(\u_a23_mem/n20624 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20626 ) );
  MUX \u_a23_mem/U20637  ( .IN0(\u_a23_mem/p_mem[13][7] ), .IN1(
        \u_a23_mem/p_mem[77][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20625 )
         );
  MUX \u_a23_mem/U20636  ( .IN0(\u_a23_mem/p_mem[45][7] ), .IN1(
        \u_a23_mem/p_mem[109][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20624 )
         );
  MUX \u_a23_mem/U20635  ( .IN0(\u_a23_mem/n20622 ), .IN1(\u_a23_mem/n20621 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20623 ) );
  MUX \u_a23_mem/U20634  ( .IN0(\u_a23_mem/p_mem[29][7] ), .IN1(
        \u_a23_mem/p_mem[93][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20622 )
         );
  MUX \u_a23_mem/U20633  ( .IN0(\u_a23_mem/p_mem[61][7] ), .IN1(
        \u_a23_mem/p_mem[125][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20621 )
         );
  MUX \u_a23_mem/U20632  ( .IN0(\u_a23_mem/n20619 ), .IN1(\u_a23_mem/n20604 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20620 ) );
  MUX \u_a23_mem/U20631  ( .IN0(\u_a23_mem/n20618 ), .IN1(\u_a23_mem/n20611 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20619 ) );
  MUX \u_a23_mem/U20630  ( .IN0(\u_a23_mem/n20617 ), .IN1(\u_a23_mem/n20614 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20618 ) );
  MUX \u_a23_mem/U20629  ( .IN0(\u_a23_mem/n20616 ), .IN1(\u_a23_mem/n20615 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20617 ) );
  MUX \u_a23_mem/U20628  ( .IN0(\u_a23_mem/p_mem[3][7] ), .IN1(
        \u_a23_mem/p_mem[67][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20616 )
         );
  MUX \u_a23_mem/U20627  ( .IN0(\u_a23_mem/p_mem[35][7] ), .IN1(
        \u_a23_mem/p_mem[99][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20615 )
         );
  MUX \u_a23_mem/U20626  ( .IN0(\u_a23_mem/n20613 ), .IN1(\u_a23_mem/n20612 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20614 ) );
  MUX \u_a23_mem/U20625  ( .IN0(\u_a23_mem/p_mem[19][7] ), .IN1(
        \u_a23_mem/p_mem[83][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20613 )
         );
  MUX \u_a23_mem/U20624  ( .IN0(\u_a23_mem/p_mem[51][7] ), .IN1(
        \u_a23_mem/p_mem[115][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20612 )
         );
  MUX \u_a23_mem/U20623  ( .IN0(\u_a23_mem/n20610 ), .IN1(\u_a23_mem/n20607 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20611 ) );
  MUX \u_a23_mem/U20622  ( .IN0(\u_a23_mem/n20609 ), .IN1(\u_a23_mem/n20608 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20610 ) );
  MUX \u_a23_mem/U20621  ( .IN0(\u_a23_mem/p_mem[11][7] ), .IN1(
        \u_a23_mem/p_mem[75][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20609 )
         );
  MUX \u_a23_mem/U20620  ( .IN0(\u_a23_mem/p_mem[43][7] ), .IN1(
        \u_a23_mem/p_mem[107][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20608 )
         );
  MUX \u_a23_mem/U20619  ( .IN0(\u_a23_mem/n20606 ), .IN1(\u_a23_mem/n20605 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20607 ) );
  MUX \u_a23_mem/U20618  ( .IN0(\u_a23_mem/p_mem[27][7] ), .IN1(
        \u_a23_mem/p_mem[91][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20606 )
         );
  MUX \u_a23_mem/U20617  ( .IN0(\u_a23_mem/p_mem[59][7] ), .IN1(
        \u_a23_mem/p_mem[123][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20605 )
         );
  MUX \u_a23_mem/U20616  ( .IN0(\u_a23_mem/n20603 ), .IN1(\u_a23_mem/n20596 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20604 ) );
  MUX \u_a23_mem/U20615  ( .IN0(\u_a23_mem/n20602 ), .IN1(\u_a23_mem/n20599 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20603 ) );
  MUX \u_a23_mem/U20614  ( .IN0(\u_a23_mem/n20601 ), .IN1(\u_a23_mem/n20600 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20602 ) );
  MUX \u_a23_mem/U20613  ( .IN0(\u_a23_mem/p_mem[7][7] ), .IN1(
        \u_a23_mem/p_mem[71][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20601 )
         );
  MUX \u_a23_mem/U20612  ( .IN0(\u_a23_mem/p_mem[39][7] ), .IN1(
        \u_a23_mem/p_mem[103][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20600 )
         );
  MUX \u_a23_mem/U20611  ( .IN0(\u_a23_mem/n20598 ), .IN1(\u_a23_mem/n20597 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20599 ) );
  MUX \u_a23_mem/U20610  ( .IN0(\u_a23_mem/p_mem[23][7] ), .IN1(
        \u_a23_mem/p_mem[87][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20598 )
         );
  MUX \u_a23_mem/U20609  ( .IN0(\u_a23_mem/p_mem[55][7] ), .IN1(
        \u_a23_mem/p_mem[119][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20597 )
         );
  MUX \u_a23_mem/U20608  ( .IN0(\u_a23_mem/n20595 ), .IN1(\u_a23_mem/n20592 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20596 ) );
  MUX \u_a23_mem/U20607  ( .IN0(\u_a23_mem/n20594 ), .IN1(\u_a23_mem/n20593 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20595 ) );
  MUX \u_a23_mem/U20606  ( .IN0(\u_a23_mem/p_mem[15][7] ), .IN1(
        \u_a23_mem/p_mem[79][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20594 )
         );
  MUX \u_a23_mem/U20605  ( .IN0(\u_a23_mem/p_mem[47][7] ), .IN1(
        \u_a23_mem/p_mem[111][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20593 )
         );
  MUX \u_a23_mem/U20604  ( .IN0(\u_a23_mem/n20591 ), .IN1(\u_a23_mem/n20590 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20592 ) );
  MUX \u_a23_mem/U20603  ( .IN0(\u_a23_mem/p_mem[31][7] ), .IN1(
        \u_a23_mem/p_mem[95][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20591 )
         );
  MUX \u_a23_mem/U20602  ( .IN0(\u_a23_mem/p_mem[63][7] ), .IN1(
        \u_a23_mem/p_mem[127][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20590 )
         );
  MUX \u_a23_mem/U20600  ( .IN0(\u_a23_mem/n20587 ), .IN1(\u_a23_mem/n20572 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20588 ) );
  MUX \u_a23_mem/U20599  ( .IN0(\u_a23_mem/n20586 ), .IN1(\u_a23_mem/n20579 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20587 ) );
  MUX \u_a23_mem/U20598  ( .IN0(\u_a23_mem/n20585 ), .IN1(\u_a23_mem/n20582 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20586 ) );
  MUX \u_a23_mem/U20597  ( .IN0(\u_a23_mem/n20584 ), .IN1(\u_a23_mem/n20583 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20585 ) );
  MUX \u_a23_mem/U20596  ( .IN0(\u_a23_mem/p_mem[2][7] ), .IN1(
        \u_a23_mem/p_mem[66][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20584 )
         );
  MUX \u_a23_mem/U20595  ( .IN0(\u_a23_mem/p_mem[34][7] ), .IN1(
        \u_a23_mem/p_mem[98][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20583 )
         );
  MUX \u_a23_mem/U20594  ( .IN0(\u_a23_mem/n20581 ), .IN1(\u_a23_mem/n20580 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20582 ) );
  MUX \u_a23_mem/U20593  ( .IN0(\u_a23_mem/p_mem[18][7] ), .IN1(
        \u_a23_mem/p_mem[82][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20581 )
         );
  MUX \u_a23_mem/U20592  ( .IN0(\u_a23_mem/p_mem[50][7] ), .IN1(
        \u_a23_mem/p_mem[114][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20580 )
         );
  MUX \u_a23_mem/U20591  ( .IN0(\u_a23_mem/n20578 ), .IN1(\u_a23_mem/n20575 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20579 ) );
  MUX \u_a23_mem/U20590  ( .IN0(\u_a23_mem/n20577 ), .IN1(\u_a23_mem/n20576 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20578 ) );
  MUX \u_a23_mem/U20589  ( .IN0(\u_a23_mem/p_mem[10][7] ), .IN1(
        \u_a23_mem/p_mem[74][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20577 )
         );
  MUX \u_a23_mem/U20588  ( .IN0(\u_a23_mem/p_mem[42][7] ), .IN1(
        \u_a23_mem/p_mem[106][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20576 )
         );
  MUX \u_a23_mem/U20587  ( .IN0(\u_a23_mem/n20574 ), .IN1(\u_a23_mem/n20573 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20575 ) );
  MUX \u_a23_mem/U20586  ( .IN0(\u_a23_mem/p_mem[26][7] ), .IN1(
        \u_a23_mem/p_mem[90][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20574 )
         );
  MUX \u_a23_mem/U20585  ( .IN0(\u_a23_mem/p_mem[58][7] ), .IN1(
        \u_a23_mem/p_mem[122][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20573 )
         );
  MUX \u_a23_mem/U20584  ( .IN0(\u_a23_mem/n20571 ), .IN1(\u_a23_mem/n20564 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20572 ) );
  MUX \u_a23_mem/U20583  ( .IN0(\u_a23_mem/n20570 ), .IN1(\u_a23_mem/n20567 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20571 ) );
  MUX \u_a23_mem/U20582  ( .IN0(\u_a23_mem/n20569 ), .IN1(\u_a23_mem/n20568 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20570 ) );
  MUX \u_a23_mem/U20581  ( .IN0(\u_a23_mem/p_mem[6][7] ), .IN1(
        \u_a23_mem/p_mem[70][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20569 )
         );
  MUX \u_a23_mem/U20580  ( .IN0(\u_a23_mem/p_mem[38][7] ), .IN1(
        \u_a23_mem/p_mem[102][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20568 )
         );
  MUX \u_a23_mem/U20579  ( .IN0(\u_a23_mem/n20566 ), .IN1(\u_a23_mem/n20565 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20567 ) );
  MUX \u_a23_mem/U20578  ( .IN0(\u_a23_mem/p_mem[22][7] ), .IN1(
        \u_a23_mem/p_mem[86][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20566 )
         );
  MUX \u_a23_mem/U20577  ( .IN0(\u_a23_mem/p_mem[54][7] ), .IN1(
        \u_a23_mem/p_mem[118][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20565 )
         );
  MUX \u_a23_mem/U20576  ( .IN0(\u_a23_mem/n20563 ), .IN1(\u_a23_mem/n20560 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20564 ) );
  MUX \u_a23_mem/U20575  ( .IN0(\u_a23_mem/n20562 ), .IN1(\u_a23_mem/n20561 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20563 ) );
  MUX \u_a23_mem/U20574  ( .IN0(\u_a23_mem/p_mem[14][7] ), .IN1(
        \u_a23_mem/p_mem[78][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20562 )
         );
  MUX \u_a23_mem/U20573  ( .IN0(\u_a23_mem/p_mem[46][7] ), .IN1(
        \u_a23_mem/p_mem[110][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20561 )
         );
  MUX \u_a23_mem/U20572  ( .IN0(\u_a23_mem/n20559 ), .IN1(\u_a23_mem/n20558 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20560 ) );
  MUX \u_a23_mem/U20571  ( .IN0(\u_a23_mem/p_mem[30][7] ), .IN1(
        \u_a23_mem/p_mem[94][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20559 )
         );
  MUX \u_a23_mem/U20570  ( .IN0(\u_a23_mem/p_mem[62][7] ), .IN1(
        \u_a23_mem/p_mem[126][7] ), .SEL(m_address[6]), .F(\u_a23_mem/n20558 )
         );
  MUX \u_a23_mem/U20537  ( .IN0(\u_a23_mem/n20525 ), .IN1(\u_a23_mem/n20510 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20526 ) );
  MUX \u_a23_mem/U20536  ( .IN0(\u_a23_mem/n20524 ), .IN1(\u_a23_mem/n20517 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20525 ) );
  MUX \u_a23_mem/U20535  ( .IN0(\u_a23_mem/n20523 ), .IN1(\u_a23_mem/n20520 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20524 ) );
  MUX \u_a23_mem/U20534  ( .IN0(\u_a23_mem/n20522 ), .IN1(\u_a23_mem/n20521 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20523 ) );
  MUX \u_a23_mem/U20533  ( .IN0(\u_a23_mem/p_mem[1][6] ), .IN1(
        \u_a23_mem/p_mem[65][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20522 )
         );
  MUX \u_a23_mem/U20532  ( .IN0(\u_a23_mem/p_mem[33][6] ), .IN1(
        \u_a23_mem/p_mem[97][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20521 )
         );
  MUX \u_a23_mem/U20531  ( .IN0(\u_a23_mem/n20519 ), .IN1(\u_a23_mem/n20518 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20520 ) );
  MUX \u_a23_mem/U20530  ( .IN0(\u_a23_mem/p_mem[17][6] ), .IN1(
        \u_a23_mem/p_mem[81][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20519 )
         );
  MUX \u_a23_mem/U20529  ( .IN0(\u_a23_mem/p_mem[49][6] ), .IN1(
        \u_a23_mem/p_mem[113][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20518 )
         );
  MUX \u_a23_mem/U20528  ( .IN0(\u_a23_mem/n20516 ), .IN1(\u_a23_mem/n20513 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20517 ) );
  MUX \u_a23_mem/U20527  ( .IN0(\u_a23_mem/n20515 ), .IN1(\u_a23_mem/n20514 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20516 ) );
  MUX \u_a23_mem/U20526  ( .IN0(\u_a23_mem/p_mem[9][6] ), .IN1(
        \u_a23_mem/p_mem[73][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20515 )
         );
  MUX \u_a23_mem/U20525  ( .IN0(\u_a23_mem/p_mem[41][6] ), .IN1(
        \u_a23_mem/p_mem[105][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20514 )
         );
  MUX \u_a23_mem/U20524  ( .IN0(\u_a23_mem/n20512 ), .IN1(\u_a23_mem/n20511 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20513 ) );
  MUX \u_a23_mem/U20523  ( .IN0(\u_a23_mem/p_mem[25][6] ), .IN1(
        \u_a23_mem/p_mem[89][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20512 )
         );
  MUX \u_a23_mem/U20522  ( .IN0(\u_a23_mem/p_mem[57][6] ), .IN1(
        \u_a23_mem/p_mem[121][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20511 )
         );
  MUX \u_a23_mem/U20521  ( .IN0(\u_a23_mem/n20509 ), .IN1(\u_a23_mem/n20502 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20510 ) );
  MUX \u_a23_mem/U20520  ( .IN0(\u_a23_mem/n20508 ), .IN1(\u_a23_mem/n20505 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20509 ) );
  MUX \u_a23_mem/U20519  ( .IN0(\u_a23_mem/n20507 ), .IN1(\u_a23_mem/n20506 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20508 ) );
  MUX \u_a23_mem/U20518  ( .IN0(\u_a23_mem/p_mem[5][6] ), .IN1(
        \u_a23_mem/p_mem[69][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20507 )
         );
  MUX \u_a23_mem/U20517  ( .IN0(\u_a23_mem/p_mem[37][6] ), .IN1(
        \u_a23_mem/p_mem[101][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20506 )
         );
  MUX \u_a23_mem/U20516  ( .IN0(\u_a23_mem/n20504 ), .IN1(\u_a23_mem/n20503 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20505 ) );
  MUX \u_a23_mem/U20515  ( .IN0(\u_a23_mem/p_mem[21][6] ), .IN1(
        \u_a23_mem/p_mem[85][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20504 )
         );
  MUX \u_a23_mem/U20514  ( .IN0(\u_a23_mem/p_mem[53][6] ), .IN1(
        \u_a23_mem/p_mem[117][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20503 )
         );
  MUX \u_a23_mem/U20513  ( .IN0(\u_a23_mem/n20501 ), .IN1(\u_a23_mem/n20498 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20502 ) );
  MUX \u_a23_mem/U20512  ( .IN0(\u_a23_mem/n20500 ), .IN1(\u_a23_mem/n20499 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20501 ) );
  MUX \u_a23_mem/U20511  ( .IN0(\u_a23_mem/p_mem[13][6] ), .IN1(
        \u_a23_mem/p_mem[77][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20500 )
         );
  MUX \u_a23_mem/U20510  ( .IN0(\u_a23_mem/p_mem[45][6] ), .IN1(
        \u_a23_mem/p_mem[109][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20499 )
         );
  MUX \u_a23_mem/U20509  ( .IN0(\u_a23_mem/n20497 ), .IN1(\u_a23_mem/n20496 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20498 ) );
  MUX \u_a23_mem/U20508  ( .IN0(\u_a23_mem/p_mem[29][6] ), .IN1(
        \u_a23_mem/p_mem[93][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20497 )
         );
  MUX \u_a23_mem/U20507  ( .IN0(\u_a23_mem/p_mem[61][6] ), .IN1(
        \u_a23_mem/p_mem[125][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20496 )
         );
  MUX \u_a23_mem/U20506  ( .IN0(\u_a23_mem/n20494 ), .IN1(\u_a23_mem/n20479 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20495 ) );
  MUX \u_a23_mem/U20505  ( .IN0(\u_a23_mem/n20493 ), .IN1(\u_a23_mem/n20486 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20494 ) );
  MUX \u_a23_mem/U20504  ( .IN0(\u_a23_mem/n20492 ), .IN1(\u_a23_mem/n20489 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20493 ) );
  MUX \u_a23_mem/U20503  ( .IN0(\u_a23_mem/n20491 ), .IN1(\u_a23_mem/n20490 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20492 ) );
  MUX \u_a23_mem/U20502  ( .IN0(\u_a23_mem/p_mem[3][6] ), .IN1(
        \u_a23_mem/p_mem[67][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20491 )
         );
  MUX \u_a23_mem/U20501  ( .IN0(\u_a23_mem/p_mem[35][6] ), .IN1(
        \u_a23_mem/p_mem[99][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20490 )
         );
  MUX \u_a23_mem/U20500  ( .IN0(\u_a23_mem/n20488 ), .IN1(\u_a23_mem/n20487 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20489 ) );
  MUX \u_a23_mem/U20499  ( .IN0(\u_a23_mem/p_mem[19][6] ), .IN1(
        \u_a23_mem/p_mem[83][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20488 )
         );
  MUX \u_a23_mem/U20498  ( .IN0(\u_a23_mem/p_mem[51][6] ), .IN1(
        \u_a23_mem/p_mem[115][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20487 )
         );
  MUX \u_a23_mem/U20497  ( .IN0(\u_a23_mem/n20485 ), .IN1(\u_a23_mem/n20482 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20486 ) );
  MUX \u_a23_mem/U20496  ( .IN0(\u_a23_mem/n20484 ), .IN1(\u_a23_mem/n20483 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20485 ) );
  MUX \u_a23_mem/U20495  ( .IN0(\u_a23_mem/p_mem[11][6] ), .IN1(
        \u_a23_mem/p_mem[75][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20484 )
         );
  MUX \u_a23_mem/U20494  ( .IN0(\u_a23_mem/p_mem[43][6] ), .IN1(
        \u_a23_mem/p_mem[107][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20483 )
         );
  MUX \u_a23_mem/U20493  ( .IN0(\u_a23_mem/n20481 ), .IN1(\u_a23_mem/n20480 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20482 ) );
  MUX \u_a23_mem/U20492  ( .IN0(\u_a23_mem/p_mem[27][6] ), .IN1(
        \u_a23_mem/p_mem[91][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20481 )
         );
  MUX \u_a23_mem/U20491  ( .IN0(\u_a23_mem/p_mem[59][6] ), .IN1(
        \u_a23_mem/p_mem[123][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20480 )
         );
  MUX \u_a23_mem/U20490  ( .IN0(\u_a23_mem/n20478 ), .IN1(\u_a23_mem/n20471 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20479 ) );
  MUX \u_a23_mem/U20489  ( .IN0(\u_a23_mem/n20477 ), .IN1(\u_a23_mem/n20474 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20478 ) );
  MUX \u_a23_mem/U20488  ( .IN0(\u_a23_mem/n20476 ), .IN1(\u_a23_mem/n20475 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20477 ) );
  MUX \u_a23_mem/U20487  ( .IN0(\u_a23_mem/p_mem[7][6] ), .IN1(
        \u_a23_mem/p_mem[71][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20476 )
         );
  MUX \u_a23_mem/U20486  ( .IN0(\u_a23_mem/p_mem[39][6] ), .IN1(
        \u_a23_mem/p_mem[103][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20475 )
         );
  MUX \u_a23_mem/U20485  ( .IN0(\u_a23_mem/n20473 ), .IN1(\u_a23_mem/n20472 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20474 ) );
  MUX \u_a23_mem/U20484  ( .IN0(\u_a23_mem/p_mem[23][6] ), .IN1(
        \u_a23_mem/p_mem[87][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20473 )
         );
  MUX \u_a23_mem/U20483  ( .IN0(\u_a23_mem/p_mem[55][6] ), .IN1(
        \u_a23_mem/p_mem[119][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20472 )
         );
  MUX \u_a23_mem/U20482  ( .IN0(\u_a23_mem/n20470 ), .IN1(\u_a23_mem/n20467 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20471 ) );
  MUX \u_a23_mem/U20481  ( .IN0(\u_a23_mem/n20469 ), .IN1(\u_a23_mem/n20468 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20470 ) );
  MUX \u_a23_mem/U20480  ( .IN0(\u_a23_mem/p_mem[15][6] ), .IN1(
        \u_a23_mem/p_mem[79][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20469 )
         );
  MUX \u_a23_mem/U20479  ( .IN0(\u_a23_mem/p_mem[47][6] ), .IN1(
        \u_a23_mem/p_mem[111][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20468 )
         );
  MUX \u_a23_mem/U20478  ( .IN0(\u_a23_mem/n20466 ), .IN1(\u_a23_mem/n20465 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20467 ) );
  MUX \u_a23_mem/U20477  ( .IN0(\u_a23_mem/p_mem[31][6] ), .IN1(
        \u_a23_mem/p_mem[95][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20466 )
         );
  MUX \u_a23_mem/U20476  ( .IN0(\u_a23_mem/p_mem[63][6] ), .IN1(
        \u_a23_mem/p_mem[127][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20465 )
         );
  MUX \u_a23_mem/U20474  ( .IN0(\u_a23_mem/n20462 ), .IN1(\u_a23_mem/n20447 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20463 ) );
  MUX \u_a23_mem/U20473  ( .IN0(\u_a23_mem/n20461 ), .IN1(\u_a23_mem/n20454 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20462 ) );
  MUX \u_a23_mem/U20472  ( .IN0(\u_a23_mem/n20460 ), .IN1(\u_a23_mem/n20457 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20461 ) );
  MUX \u_a23_mem/U20471  ( .IN0(\u_a23_mem/n20459 ), .IN1(\u_a23_mem/n20458 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20460 ) );
  MUX \u_a23_mem/U20470  ( .IN0(\u_a23_mem/p_mem[2][6] ), .IN1(
        \u_a23_mem/p_mem[66][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20459 )
         );
  MUX \u_a23_mem/U20469  ( .IN0(\u_a23_mem/p_mem[34][6] ), .IN1(
        \u_a23_mem/p_mem[98][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20458 )
         );
  MUX \u_a23_mem/U20468  ( .IN0(\u_a23_mem/n20456 ), .IN1(\u_a23_mem/n20455 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20457 ) );
  MUX \u_a23_mem/U20467  ( .IN0(\u_a23_mem/p_mem[18][6] ), .IN1(
        \u_a23_mem/p_mem[82][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20456 )
         );
  MUX \u_a23_mem/U20466  ( .IN0(\u_a23_mem/p_mem[50][6] ), .IN1(
        \u_a23_mem/p_mem[114][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20455 )
         );
  MUX \u_a23_mem/U20465  ( .IN0(\u_a23_mem/n20453 ), .IN1(\u_a23_mem/n20450 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20454 ) );
  MUX \u_a23_mem/U20464  ( .IN0(\u_a23_mem/n20452 ), .IN1(\u_a23_mem/n20451 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20453 ) );
  MUX \u_a23_mem/U20463  ( .IN0(\u_a23_mem/p_mem[10][6] ), .IN1(
        \u_a23_mem/p_mem[74][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20452 )
         );
  MUX \u_a23_mem/U20462  ( .IN0(\u_a23_mem/p_mem[42][6] ), .IN1(
        \u_a23_mem/p_mem[106][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20451 )
         );
  MUX \u_a23_mem/U20461  ( .IN0(\u_a23_mem/n20449 ), .IN1(\u_a23_mem/n20448 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20450 ) );
  MUX \u_a23_mem/U20460  ( .IN0(\u_a23_mem/p_mem[26][6] ), .IN1(
        \u_a23_mem/p_mem[90][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20449 )
         );
  MUX \u_a23_mem/U20459  ( .IN0(\u_a23_mem/p_mem[58][6] ), .IN1(
        \u_a23_mem/p_mem[122][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20448 )
         );
  MUX \u_a23_mem/U20458  ( .IN0(\u_a23_mem/n20446 ), .IN1(\u_a23_mem/n20439 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20447 ) );
  MUX \u_a23_mem/U20457  ( .IN0(\u_a23_mem/n20445 ), .IN1(\u_a23_mem/n20442 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20446 ) );
  MUX \u_a23_mem/U20456  ( .IN0(\u_a23_mem/n20444 ), .IN1(\u_a23_mem/n20443 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20445 ) );
  MUX \u_a23_mem/U20455  ( .IN0(\u_a23_mem/p_mem[6][6] ), .IN1(
        \u_a23_mem/p_mem[70][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20444 )
         );
  MUX \u_a23_mem/U20454  ( .IN0(\u_a23_mem/p_mem[38][6] ), .IN1(
        \u_a23_mem/p_mem[102][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20443 )
         );
  MUX \u_a23_mem/U20453  ( .IN0(\u_a23_mem/n20441 ), .IN1(\u_a23_mem/n20440 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20442 ) );
  MUX \u_a23_mem/U20452  ( .IN0(\u_a23_mem/p_mem[22][6] ), .IN1(
        \u_a23_mem/p_mem[86][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20441 )
         );
  MUX \u_a23_mem/U20451  ( .IN0(\u_a23_mem/p_mem[54][6] ), .IN1(
        \u_a23_mem/p_mem[118][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20440 )
         );
  MUX \u_a23_mem/U20450  ( .IN0(\u_a23_mem/n20438 ), .IN1(\u_a23_mem/n20435 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20439 ) );
  MUX \u_a23_mem/U20449  ( .IN0(\u_a23_mem/n20437 ), .IN1(\u_a23_mem/n20436 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20438 ) );
  MUX \u_a23_mem/U20448  ( .IN0(\u_a23_mem/p_mem[14][6] ), .IN1(
        \u_a23_mem/p_mem[78][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20437 )
         );
  MUX \u_a23_mem/U20447  ( .IN0(\u_a23_mem/p_mem[46][6] ), .IN1(
        \u_a23_mem/p_mem[110][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20436 )
         );
  MUX \u_a23_mem/U20446  ( .IN0(\u_a23_mem/n20434 ), .IN1(\u_a23_mem/n20433 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20435 ) );
  MUX \u_a23_mem/U20445  ( .IN0(\u_a23_mem/p_mem[30][6] ), .IN1(
        \u_a23_mem/p_mem[94][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20434 )
         );
  MUX \u_a23_mem/U20444  ( .IN0(\u_a23_mem/p_mem[62][6] ), .IN1(
        \u_a23_mem/p_mem[126][6] ), .SEL(m_address[6]), .F(\u_a23_mem/n20433 )
         );
  MUX \u_a23_mem/U20411  ( .IN0(\u_a23_mem/n20400 ), .IN1(\u_a23_mem/n20385 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20401 ) );
  MUX \u_a23_mem/U20410  ( .IN0(\u_a23_mem/n20399 ), .IN1(\u_a23_mem/n20392 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20400 ) );
  MUX \u_a23_mem/U20409  ( .IN0(\u_a23_mem/n20398 ), .IN1(\u_a23_mem/n20395 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20399 ) );
  MUX \u_a23_mem/U20408  ( .IN0(\u_a23_mem/n20397 ), .IN1(\u_a23_mem/n20396 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20398 ) );
  MUX \u_a23_mem/U20407  ( .IN0(\u_a23_mem/p_mem[1][5] ), .IN1(
        \u_a23_mem/p_mem[65][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20397 )
         );
  MUX \u_a23_mem/U20406  ( .IN0(\u_a23_mem/p_mem[33][5] ), .IN1(
        \u_a23_mem/p_mem[97][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20396 )
         );
  MUX \u_a23_mem/U20405  ( .IN0(\u_a23_mem/n20394 ), .IN1(\u_a23_mem/n20393 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20395 ) );
  MUX \u_a23_mem/U20404  ( .IN0(\u_a23_mem/p_mem[17][5] ), .IN1(
        \u_a23_mem/p_mem[81][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20394 )
         );
  MUX \u_a23_mem/U20403  ( .IN0(\u_a23_mem/p_mem[49][5] ), .IN1(
        \u_a23_mem/p_mem[113][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20393 )
         );
  MUX \u_a23_mem/U20402  ( .IN0(\u_a23_mem/n20391 ), .IN1(\u_a23_mem/n20388 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20392 ) );
  MUX \u_a23_mem/U20401  ( .IN0(\u_a23_mem/n20390 ), .IN1(\u_a23_mem/n20389 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20391 ) );
  MUX \u_a23_mem/U20400  ( .IN0(\u_a23_mem/p_mem[9][5] ), .IN1(
        \u_a23_mem/p_mem[73][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20390 )
         );
  MUX \u_a23_mem/U20399  ( .IN0(\u_a23_mem/p_mem[41][5] ), .IN1(
        \u_a23_mem/p_mem[105][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20389 )
         );
  MUX \u_a23_mem/U20398  ( .IN0(\u_a23_mem/n20387 ), .IN1(\u_a23_mem/n20386 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20388 ) );
  MUX \u_a23_mem/U20397  ( .IN0(\u_a23_mem/p_mem[25][5] ), .IN1(
        \u_a23_mem/p_mem[89][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20387 )
         );
  MUX \u_a23_mem/U20396  ( .IN0(\u_a23_mem/p_mem[57][5] ), .IN1(
        \u_a23_mem/p_mem[121][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20386 )
         );
  MUX \u_a23_mem/U20395  ( .IN0(\u_a23_mem/n20384 ), .IN1(\u_a23_mem/n20377 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20385 ) );
  MUX \u_a23_mem/U20394  ( .IN0(\u_a23_mem/n20383 ), .IN1(\u_a23_mem/n20380 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20384 ) );
  MUX \u_a23_mem/U20393  ( .IN0(\u_a23_mem/n20382 ), .IN1(\u_a23_mem/n20381 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20383 ) );
  MUX \u_a23_mem/U20392  ( .IN0(\u_a23_mem/p_mem[5][5] ), .IN1(
        \u_a23_mem/p_mem[69][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20382 )
         );
  MUX \u_a23_mem/U20391  ( .IN0(\u_a23_mem/p_mem[37][5] ), .IN1(
        \u_a23_mem/p_mem[101][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20381 )
         );
  MUX \u_a23_mem/U20390  ( .IN0(\u_a23_mem/n20379 ), .IN1(\u_a23_mem/n20378 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20380 ) );
  MUX \u_a23_mem/U20389  ( .IN0(\u_a23_mem/p_mem[21][5] ), .IN1(
        \u_a23_mem/p_mem[85][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20379 )
         );
  MUX \u_a23_mem/U20388  ( .IN0(\u_a23_mem/p_mem[53][5] ), .IN1(
        \u_a23_mem/p_mem[117][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20378 )
         );
  MUX \u_a23_mem/U20387  ( .IN0(\u_a23_mem/n20376 ), .IN1(\u_a23_mem/n20373 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20377 ) );
  MUX \u_a23_mem/U20386  ( .IN0(\u_a23_mem/n20375 ), .IN1(\u_a23_mem/n20374 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20376 ) );
  MUX \u_a23_mem/U20385  ( .IN0(\u_a23_mem/p_mem[13][5] ), .IN1(
        \u_a23_mem/p_mem[77][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20375 )
         );
  MUX \u_a23_mem/U20384  ( .IN0(\u_a23_mem/p_mem[45][5] ), .IN1(
        \u_a23_mem/p_mem[109][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20374 )
         );
  MUX \u_a23_mem/U20383  ( .IN0(\u_a23_mem/n20372 ), .IN1(\u_a23_mem/n20371 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20373 ) );
  MUX \u_a23_mem/U20382  ( .IN0(\u_a23_mem/p_mem[29][5] ), .IN1(
        \u_a23_mem/p_mem[93][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20372 )
         );
  MUX \u_a23_mem/U20381  ( .IN0(\u_a23_mem/p_mem[61][5] ), .IN1(
        \u_a23_mem/p_mem[125][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20371 )
         );
  MUX \u_a23_mem/U20380  ( .IN0(\u_a23_mem/n20369 ), .IN1(\u_a23_mem/n20354 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20370 ) );
  MUX \u_a23_mem/U20379  ( .IN0(\u_a23_mem/n20368 ), .IN1(\u_a23_mem/n20361 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20369 ) );
  MUX \u_a23_mem/U20378  ( .IN0(\u_a23_mem/n20367 ), .IN1(\u_a23_mem/n20364 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20368 ) );
  MUX \u_a23_mem/U20377  ( .IN0(\u_a23_mem/n20366 ), .IN1(\u_a23_mem/n20365 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20367 ) );
  MUX \u_a23_mem/U20376  ( .IN0(\u_a23_mem/p_mem[3][5] ), .IN1(
        \u_a23_mem/p_mem[67][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20366 )
         );
  MUX \u_a23_mem/U20375  ( .IN0(\u_a23_mem/p_mem[35][5] ), .IN1(
        \u_a23_mem/p_mem[99][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20365 )
         );
  MUX \u_a23_mem/U20374  ( .IN0(\u_a23_mem/n20363 ), .IN1(\u_a23_mem/n20362 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20364 ) );
  MUX \u_a23_mem/U20373  ( .IN0(\u_a23_mem/p_mem[19][5] ), .IN1(
        \u_a23_mem/p_mem[83][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20363 )
         );
  MUX \u_a23_mem/U20372  ( .IN0(\u_a23_mem/p_mem[51][5] ), .IN1(
        \u_a23_mem/p_mem[115][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20362 )
         );
  MUX \u_a23_mem/U20371  ( .IN0(\u_a23_mem/n20360 ), .IN1(\u_a23_mem/n20357 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20361 ) );
  MUX \u_a23_mem/U20370  ( .IN0(\u_a23_mem/n20359 ), .IN1(\u_a23_mem/n20358 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20360 ) );
  MUX \u_a23_mem/U20369  ( .IN0(\u_a23_mem/p_mem[11][5] ), .IN1(
        \u_a23_mem/p_mem[75][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20359 )
         );
  MUX \u_a23_mem/U20368  ( .IN0(\u_a23_mem/p_mem[43][5] ), .IN1(
        \u_a23_mem/p_mem[107][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20358 )
         );
  MUX \u_a23_mem/U20367  ( .IN0(\u_a23_mem/n20356 ), .IN1(\u_a23_mem/n20355 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20357 ) );
  MUX \u_a23_mem/U20366  ( .IN0(\u_a23_mem/p_mem[27][5] ), .IN1(
        \u_a23_mem/p_mem[91][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20356 )
         );
  MUX \u_a23_mem/U20365  ( .IN0(\u_a23_mem/p_mem[59][5] ), .IN1(
        \u_a23_mem/p_mem[123][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20355 )
         );
  MUX \u_a23_mem/U20364  ( .IN0(\u_a23_mem/n20353 ), .IN1(\u_a23_mem/n20346 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20354 ) );
  MUX \u_a23_mem/U20363  ( .IN0(\u_a23_mem/n20352 ), .IN1(\u_a23_mem/n20349 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20353 ) );
  MUX \u_a23_mem/U20362  ( .IN0(\u_a23_mem/n20351 ), .IN1(\u_a23_mem/n20350 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20352 ) );
  MUX \u_a23_mem/U20361  ( .IN0(\u_a23_mem/p_mem[7][5] ), .IN1(
        \u_a23_mem/p_mem[71][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20351 )
         );
  MUX \u_a23_mem/U20360  ( .IN0(\u_a23_mem/p_mem[39][5] ), .IN1(
        \u_a23_mem/p_mem[103][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20350 )
         );
  MUX \u_a23_mem/U20359  ( .IN0(\u_a23_mem/n20348 ), .IN1(\u_a23_mem/n20347 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20349 ) );
  MUX \u_a23_mem/U20358  ( .IN0(\u_a23_mem/p_mem[23][5] ), .IN1(
        \u_a23_mem/p_mem[87][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20348 )
         );
  MUX \u_a23_mem/U20357  ( .IN0(\u_a23_mem/p_mem[55][5] ), .IN1(
        \u_a23_mem/p_mem[119][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20347 )
         );
  MUX \u_a23_mem/U20356  ( .IN0(\u_a23_mem/n20345 ), .IN1(\u_a23_mem/n20342 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20346 ) );
  MUX \u_a23_mem/U20355  ( .IN0(\u_a23_mem/n20344 ), .IN1(\u_a23_mem/n20343 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20345 ) );
  MUX \u_a23_mem/U20354  ( .IN0(\u_a23_mem/p_mem[15][5] ), .IN1(
        \u_a23_mem/p_mem[79][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20344 )
         );
  MUX \u_a23_mem/U20353  ( .IN0(\u_a23_mem/p_mem[47][5] ), .IN1(
        \u_a23_mem/p_mem[111][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20343 )
         );
  MUX \u_a23_mem/U20352  ( .IN0(\u_a23_mem/n20341 ), .IN1(\u_a23_mem/n20340 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20342 ) );
  MUX \u_a23_mem/U20351  ( .IN0(\u_a23_mem/p_mem[31][5] ), .IN1(
        \u_a23_mem/p_mem[95][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20341 )
         );
  MUX \u_a23_mem/U20350  ( .IN0(\u_a23_mem/p_mem[63][5] ), .IN1(
        \u_a23_mem/p_mem[127][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20340 )
         );
  MUX \u_a23_mem/U20348  ( .IN0(\u_a23_mem/n20337 ), .IN1(\u_a23_mem/n20322 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20338 ) );
  MUX \u_a23_mem/U20347  ( .IN0(\u_a23_mem/n20336 ), .IN1(\u_a23_mem/n20329 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20337 ) );
  MUX \u_a23_mem/U20346  ( .IN0(\u_a23_mem/n20335 ), .IN1(\u_a23_mem/n20332 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20336 ) );
  MUX \u_a23_mem/U20345  ( .IN0(\u_a23_mem/n20334 ), .IN1(\u_a23_mem/n20333 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20335 ) );
  MUX \u_a23_mem/U20344  ( .IN0(\u_a23_mem/p_mem[2][5] ), .IN1(
        \u_a23_mem/p_mem[66][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20334 )
         );
  MUX \u_a23_mem/U20343  ( .IN0(\u_a23_mem/p_mem[34][5] ), .IN1(
        \u_a23_mem/p_mem[98][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20333 )
         );
  MUX \u_a23_mem/U20342  ( .IN0(\u_a23_mem/n20331 ), .IN1(\u_a23_mem/n20330 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20332 ) );
  MUX \u_a23_mem/U20341  ( .IN0(\u_a23_mem/p_mem[18][5] ), .IN1(
        \u_a23_mem/p_mem[82][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20331 )
         );
  MUX \u_a23_mem/U20340  ( .IN0(\u_a23_mem/p_mem[50][5] ), .IN1(
        \u_a23_mem/p_mem[114][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20330 )
         );
  MUX \u_a23_mem/U20339  ( .IN0(\u_a23_mem/n20328 ), .IN1(\u_a23_mem/n20325 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20329 ) );
  MUX \u_a23_mem/U20338  ( .IN0(\u_a23_mem/n20327 ), .IN1(\u_a23_mem/n20326 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20328 ) );
  MUX \u_a23_mem/U20337  ( .IN0(\u_a23_mem/p_mem[10][5] ), .IN1(
        \u_a23_mem/p_mem[74][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20327 )
         );
  MUX \u_a23_mem/U20336  ( .IN0(\u_a23_mem/p_mem[42][5] ), .IN1(
        \u_a23_mem/p_mem[106][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20326 )
         );
  MUX \u_a23_mem/U20335  ( .IN0(\u_a23_mem/n20324 ), .IN1(\u_a23_mem/n20323 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20325 ) );
  MUX \u_a23_mem/U20334  ( .IN0(\u_a23_mem/p_mem[26][5] ), .IN1(
        \u_a23_mem/p_mem[90][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20324 )
         );
  MUX \u_a23_mem/U20333  ( .IN0(\u_a23_mem/p_mem[58][5] ), .IN1(
        \u_a23_mem/p_mem[122][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20323 )
         );
  MUX \u_a23_mem/U20332  ( .IN0(\u_a23_mem/n20321 ), .IN1(\u_a23_mem/n20314 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20322 ) );
  MUX \u_a23_mem/U20331  ( .IN0(\u_a23_mem/n20320 ), .IN1(\u_a23_mem/n20317 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20321 ) );
  MUX \u_a23_mem/U20330  ( .IN0(\u_a23_mem/n20319 ), .IN1(\u_a23_mem/n20318 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20320 ) );
  MUX \u_a23_mem/U20329  ( .IN0(\u_a23_mem/p_mem[6][5] ), .IN1(
        \u_a23_mem/p_mem[70][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20319 )
         );
  MUX \u_a23_mem/U20328  ( .IN0(\u_a23_mem/p_mem[38][5] ), .IN1(
        \u_a23_mem/p_mem[102][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20318 )
         );
  MUX \u_a23_mem/U20327  ( .IN0(\u_a23_mem/n20316 ), .IN1(\u_a23_mem/n20315 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20317 ) );
  MUX \u_a23_mem/U20326  ( .IN0(\u_a23_mem/p_mem[22][5] ), .IN1(
        \u_a23_mem/p_mem[86][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20316 )
         );
  MUX \u_a23_mem/U20325  ( .IN0(\u_a23_mem/p_mem[54][5] ), .IN1(
        \u_a23_mem/p_mem[118][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20315 )
         );
  MUX \u_a23_mem/U20324  ( .IN0(\u_a23_mem/n20313 ), .IN1(\u_a23_mem/n20310 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20314 ) );
  MUX \u_a23_mem/U20323  ( .IN0(\u_a23_mem/n20312 ), .IN1(\u_a23_mem/n20311 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20313 ) );
  MUX \u_a23_mem/U20322  ( .IN0(\u_a23_mem/p_mem[14][5] ), .IN1(
        \u_a23_mem/p_mem[78][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20312 )
         );
  MUX \u_a23_mem/U20321  ( .IN0(\u_a23_mem/p_mem[46][5] ), .IN1(
        \u_a23_mem/p_mem[110][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20311 )
         );
  MUX \u_a23_mem/U20320  ( .IN0(\u_a23_mem/n20309 ), .IN1(\u_a23_mem/n20308 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20310 ) );
  MUX \u_a23_mem/U20319  ( .IN0(\u_a23_mem/p_mem[30][5] ), .IN1(
        \u_a23_mem/p_mem[94][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20309 )
         );
  MUX \u_a23_mem/U20318  ( .IN0(\u_a23_mem/p_mem[62][5] ), .IN1(
        \u_a23_mem/p_mem[126][5] ), .SEL(m_address[6]), .F(\u_a23_mem/n20308 )
         );
  MUX \u_a23_mem/U20285  ( .IN0(\u_a23_mem/n20275 ), .IN1(\u_a23_mem/n20260 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20276 ) );
  MUX \u_a23_mem/U20284  ( .IN0(\u_a23_mem/n20274 ), .IN1(\u_a23_mem/n20267 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20275 ) );
  MUX \u_a23_mem/U20283  ( .IN0(\u_a23_mem/n20273 ), .IN1(\u_a23_mem/n20270 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20274 ) );
  MUX \u_a23_mem/U20282  ( .IN0(\u_a23_mem/n20272 ), .IN1(\u_a23_mem/n20271 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20273 ) );
  MUX \u_a23_mem/U20281  ( .IN0(\u_a23_mem/p_mem[1][4] ), .IN1(
        \u_a23_mem/p_mem[65][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20272 )
         );
  MUX \u_a23_mem/U20280  ( .IN0(\u_a23_mem/p_mem[33][4] ), .IN1(
        \u_a23_mem/p_mem[97][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20271 )
         );
  MUX \u_a23_mem/U20279  ( .IN0(\u_a23_mem/n20269 ), .IN1(\u_a23_mem/n20268 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20270 ) );
  MUX \u_a23_mem/U20278  ( .IN0(\u_a23_mem/p_mem[17][4] ), .IN1(
        \u_a23_mem/p_mem[81][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20269 )
         );
  MUX \u_a23_mem/U20277  ( .IN0(\u_a23_mem/p_mem[49][4] ), .IN1(
        \u_a23_mem/p_mem[113][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20268 )
         );
  MUX \u_a23_mem/U20276  ( .IN0(\u_a23_mem/n20266 ), .IN1(\u_a23_mem/n20263 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20267 ) );
  MUX \u_a23_mem/U20275  ( .IN0(\u_a23_mem/n20265 ), .IN1(\u_a23_mem/n20264 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20266 ) );
  MUX \u_a23_mem/U20274  ( .IN0(\u_a23_mem/p_mem[9][4] ), .IN1(
        \u_a23_mem/p_mem[73][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20265 )
         );
  MUX \u_a23_mem/U20273  ( .IN0(\u_a23_mem/p_mem[41][4] ), .IN1(
        \u_a23_mem/p_mem[105][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20264 )
         );
  MUX \u_a23_mem/U20272  ( .IN0(\u_a23_mem/n20262 ), .IN1(\u_a23_mem/n20261 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20263 ) );
  MUX \u_a23_mem/U20271  ( .IN0(\u_a23_mem/p_mem[25][4] ), .IN1(
        \u_a23_mem/p_mem[89][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20262 )
         );
  MUX \u_a23_mem/U20270  ( .IN0(\u_a23_mem/p_mem[57][4] ), .IN1(
        \u_a23_mem/p_mem[121][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20261 )
         );
  MUX \u_a23_mem/U20269  ( .IN0(\u_a23_mem/n20259 ), .IN1(\u_a23_mem/n20252 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20260 ) );
  MUX \u_a23_mem/U20268  ( .IN0(\u_a23_mem/n20258 ), .IN1(\u_a23_mem/n20255 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20259 ) );
  MUX \u_a23_mem/U20267  ( .IN0(\u_a23_mem/n20257 ), .IN1(\u_a23_mem/n20256 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20258 ) );
  MUX \u_a23_mem/U20266  ( .IN0(\u_a23_mem/p_mem[5][4] ), .IN1(
        \u_a23_mem/p_mem[69][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20257 )
         );
  MUX \u_a23_mem/U20265  ( .IN0(\u_a23_mem/p_mem[37][4] ), .IN1(
        \u_a23_mem/p_mem[101][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20256 )
         );
  MUX \u_a23_mem/U20264  ( .IN0(\u_a23_mem/n20254 ), .IN1(\u_a23_mem/n20253 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20255 ) );
  MUX \u_a23_mem/U20263  ( .IN0(\u_a23_mem/p_mem[21][4] ), .IN1(
        \u_a23_mem/p_mem[85][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20254 )
         );
  MUX \u_a23_mem/U20262  ( .IN0(\u_a23_mem/p_mem[53][4] ), .IN1(
        \u_a23_mem/p_mem[117][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20253 )
         );
  MUX \u_a23_mem/U20261  ( .IN0(\u_a23_mem/n20251 ), .IN1(\u_a23_mem/n20248 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20252 ) );
  MUX \u_a23_mem/U20260  ( .IN0(\u_a23_mem/n20250 ), .IN1(\u_a23_mem/n20249 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20251 ) );
  MUX \u_a23_mem/U20259  ( .IN0(\u_a23_mem/p_mem[13][4] ), .IN1(
        \u_a23_mem/p_mem[77][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20250 )
         );
  MUX \u_a23_mem/U20258  ( .IN0(\u_a23_mem/p_mem[45][4] ), .IN1(
        \u_a23_mem/p_mem[109][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20249 )
         );
  MUX \u_a23_mem/U20257  ( .IN0(\u_a23_mem/n20247 ), .IN1(\u_a23_mem/n20246 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20248 ) );
  MUX \u_a23_mem/U20256  ( .IN0(\u_a23_mem/p_mem[29][4] ), .IN1(
        \u_a23_mem/p_mem[93][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20247 )
         );
  MUX \u_a23_mem/U20255  ( .IN0(\u_a23_mem/p_mem[61][4] ), .IN1(
        \u_a23_mem/p_mem[125][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20246 )
         );
  MUX \u_a23_mem/U20254  ( .IN0(\u_a23_mem/n20244 ), .IN1(\u_a23_mem/n20229 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20245 ) );
  MUX \u_a23_mem/U20253  ( .IN0(\u_a23_mem/n20243 ), .IN1(\u_a23_mem/n20236 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20244 ) );
  MUX \u_a23_mem/U20252  ( .IN0(\u_a23_mem/n20242 ), .IN1(\u_a23_mem/n20239 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20243 ) );
  MUX \u_a23_mem/U20251  ( .IN0(\u_a23_mem/n20241 ), .IN1(\u_a23_mem/n20240 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20242 ) );
  MUX \u_a23_mem/U20250  ( .IN0(\u_a23_mem/p_mem[3][4] ), .IN1(
        \u_a23_mem/p_mem[67][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20241 )
         );
  MUX \u_a23_mem/U20249  ( .IN0(\u_a23_mem/p_mem[35][4] ), .IN1(
        \u_a23_mem/p_mem[99][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20240 )
         );
  MUX \u_a23_mem/U20248  ( .IN0(\u_a23_mem/n20238 ), .IN1(\u_a23_mem/n20237 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20239 ) );
  MUX \u_a23_mem/U20247  ( .IN0(\u_a23_mem/p_mem[19][4] ), .IN1(
        \u_a23_mem/p_mem[83][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20238 )
         );
  MUX \u_a23_mem/U20246  ( .IN0(\u_a23_mem/p_mem[51][4] ), .IN1(
        \u_a23_mem/p_mem[115][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20237 )
         );
  MUX \u_a23_mem/U20245  ( .IN0(\u_a23_mem/n20235 ), .IN1(\u_a23_mem/n20232 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20236 ) );
  MUX \u_a23_mem/U20244  ( .IN0(\u_a23_mem/n20234 ), .IN1(\u_a23_mem/n20233 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20235 ) );
  MUX \u_a23_mem/U20243  ( .IN0(\u_a23_mem/p_mem[11][4] ), .IN1(
        \u_a23_mem/p_mem[75][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20234 )
         );
  MUX \u_a23_mem/U20242  ( .IN0(\u_a23_mem/p_mem[43][4] ), .IN1(
        \u_a23_mem/p_mem[107][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20233 )
         );
  MUX \u_a23_mem/U20241  ( .IN0(\u_a23_mem/n20231 ), .IN1(\u_a23_mem/n20230 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20232 ) );
  MUX \u_a23_mem/U20240  ( .IN0(\u_a23_mem/p_mem[27][4] ), .IN1(
        \u_a23_mem/p_mem[91][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20231 )
         );
  MUX \u_a23_mem/U20239  ( .IN0(\u_a23_mem/p_mem[59][4] ), .IN1(
        \u_a23_mem/p_mem[123][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20230 )
         );
  MUX \u_a23_mem/U20238  ( .IN0(\u_a23_mem/n20228 ), .IN1(\u_a23_mem/n20221 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20229 ) );
  MUX \u_a23_mem/U20237  ( .IN0(\u_a23_mem/n20227 ), .IN1(\u_a23_mem/n20224 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20228 ) );
  MUX \u_a23_mem/U20236  ( .IN0(\u_a23_mem/n20226 ), .IN1(\u_a23_mem/n20225 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20227 ) );
  MUX \u_a23_mem/U20235  ( .IN0(\u_a23_mem/p_mem[7][4] ), .IN1(
        \u_a23_mem/p_mem[71][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20226 )
         );
  MUX \u_a23_mem/U20234  ( .IN0(\u_a23_mem/p_mem[39][4] ), .IN1(
        \u_a23_mem/p_mem[103][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20225 )
         );
  MUX \u_a23_mem/U20233  ( .IN0(\u_a23_mem/n20223 ), .IN1(\u_a23_mem/n20222 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20224 ) );
  MUX \u_a23_mem/U20232  ( .IN0(\u_a23_mem/p_mem[23][4] ), .IN1(
        \u_a23_mem/p_mem[87][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20223 )
         );
  MUX \u_a23_mem/U20231  ( .IN0(\u_a23_mem/p_mem[55][4] ), .IN1(
        \u_a23_mem/p_mem[119][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20222 )
         );
  MUX \u_a23_mem/U20230  ( .IN0(\u_a23_mem/n20220 ), .IN1(\u_a23_mem/n20217 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20221 ) );
  MUX \u_a23_mem/U20229  ( .IN0(\u_a23_mem/n20219 ), .IN1(\u_a23_mem/n20218 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20220 ) );
  MUX \u_a23_mem/U20228  ( .IN0(\u_a23_mem/p_mem[15][4] ), .IN1(
        \u_a23_mem/p_mem[79][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20219 )
         );
  MUX \u_a23_mem/U20227  ( .IN0(\u_a23_mem/p_mem[47][4] ), .IN1(
        \u_a23_mem/p_mem[111][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20218 )
         );
  MUX \u_a23_mem/U20226  ( .IN0(\u_a23_mem/n20216 ), .IN1(\u_a23_mem/n20215 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20217 ) );
  MUX \u_a23_mem/U20225  ( .IN0(\u_a23_mem/p_mem[31][4] ), .IN1(
        \u_a23_mem/p_mem[95][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20216 )
         );
  MUX \u_a23_mem/U20224  ( .IN0(\u_a23_mem/p_mem[63][4] ), .IN1(
        \u_a23_mem/p_mem[127][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20215 )
         );
  MUX \u_a23_mem/U20222  ( .IN0(\u_a23_mem/n20212 ), .IN1(\u_a23_mem/n20197 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20213 ) );
  MUX \u_a23_mem/U20221  ( .IN0(\u_a23_mem/n20211 ), .IN1(\u_a23_mem/n20204 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20212 ) );
  MUX \u_a23_mem/U20220  ( .IN0(\u_a23_mem/n20210 ), .IN1(\u_a23_mem/n20207 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20211 ) );
  MUX \u_a23_mem/U20219  ( .IN0(\u_a23_mem/n20209 ), .IN1(\u_a23_mem/n20208 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20210 ) );
  MUX \u_a23_mem/U20218  ( .IN0(\u_a23_mem/p_mem[2][4] ), .IN1(
        \u_a23_mem/p_mem[66][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20209 )
         );
  MUX \u_a23_mem/U20217  ( .IN0(\u_a23_mem/p_mem[34][4] ), .IN1(
        \u_a23_mem/p_mem[98][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20208 )
         );
  MUX \u_a23_mem/U20216  ( .IN0(\u_a23_mem/n20206 ), .IN1(\u_a23_mem/n20205 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20207 ) );
  MUX \u_a23_mem/U20215  ( .IN0(\u_a23_mem/p_mem[18][4] ), .IN1(
        \u_a23_mem/p_mem[82][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20206 )
         );
  MUX \u_a23_mem/U20214  ( .IN0(\u_a23_mem/p_mem[50][4] ), .IN1(
        \u_a23_mem/p_mem[114][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20205 )
         );
  MUX \u_a23_mem/U20213  ( .IN0(\u_a23_mem/n20203 ), .IN1(\u_a23_mem/n20200 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20204 ) );
  MUX \u_a23_mem/U20212  ( .IN0(\u_a23_mem/n20202 ), .IN1(\u_a23_mem/n20201 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20203 ) );
  MUX \u_a23_mem/U20211  ( .IN0(\u_a23_mem/p_mem[10][4] ), .IN1(
        \u_a23_mem/p_mem[74][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20202 )
         );
  MUX \u_a23_mem/U20210  ( .IN0(\u_a23_mem/p_mem[42][4] ), .IN1(
        \u_a23_mem/p_mem[106][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20201 )
         );
  MUX \u_a23_mem/U20209  ( .IN0(\u_a23_mem/n20199 ), .IN1(\u_a23_mem/n20198 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20200 ) );
  MUX \u_a23_mem/U20208  ( .IN0(\u_a23_mem/p_mem[26][4] ), .IN1(
        \u_a23_mem/p_mem[90][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20199 )
         );
  MUX \u_a23_mem/U20207  ( .IN0(\u_a23_mem/p_mem[58][4] ), .IN1(
        \u_a23_mem/p_mem[122][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20198 )
         );
  MUX \u_a23_mem/U20206  ( .IN0(\u_a23_mem/n20196 ), .IN1(\u_a23_mem/n20189 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20197 ) );
  MUX \u_a23_mem/U20205  ( .IN0(\u_a23_mem/n20195 ), .IN1(\u_a23_mem/n20192 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20196 ) );
  MUX \u_a23_mem/U20204  ( .IN0(\u_a23_mem/n20194 ), .IN1(\u_a23_mem/n20193 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20195 ) );
  MUX \u_a23_mem/U20203  ( .IN0(\u_a23_mem/p_mem[6][4] ), .IN1(
        \u_a23_mem/p_mem[70][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20194 )
         );
  MUX \u_a23_mem/U20202  ( .IN0(\u_a23_mem/p_mem[38][4] ), .IN1(
        \u_a23_mem/p_mem[102][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20193 )
         );
  MUX \u_a23_mem/U20201  ( .IN0(\u_a23_mem/n20191 ), .IN1(\u_a23_mem/n20190 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20192 ) );
  MUX \u_a23_mem/U20200  ( .IN0(\u_a23_mem/p_mem[22][4] ), .IN1(
        \u_a23_mem/p_mem[86][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20191 )
         );
  MUX \u_a23_mem/U20199  ( .IN0(\u_a23_mem/p_mem[54][4] ), .IN1(
        \u_a23_mem/p_mem[118][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20190 )
         );
  MUX \u_a23_mem/U20198  ( .IN0(\u_a23_mem/n20188 ), .IN1(\u_a23_mem/n20185 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20189 ) );
  MUX \u_a23_mem/U20197  ( .IN0(\u_a23_mem/n20187 ), .IN1(\u_a23_mem/n20186 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20188 ) );
  MUX \u_a23_mem/U20196  ( .IN0(\u_a23_mem/p_mem[14][4] ), .IN1(
        \u_a23_mem/p_mem[78][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20187 )
         );
  MUX \u_a23_mem/U20195  ( .IN0(\u_a23_mem/p_mem[46][4] ), .IN1(
        \u_a23_mem/p_mem[110][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20186 )
         );
  MUX \u_a23_mem/U20194  ( .IN0(\u_a23_mem/n20184 ), .IN1(\u_a23_mem/n20183 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20185 ) );
  MUX \u_a23_mem/U20193  ( .IN0(\u_a23_mem/p_mem[30][4] ), .IN1(
        \u_a23_mem/p_mem[94][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20184 )
         );
  MUX \u_a23_mem/U20192  ( .IN0(\u_a23_mem/p_mem[62][4] ), .IN1(
        \u_a23_mem/p_mem[126][4] ), .SEL(m_address[6]), .F(\u_a23_mem/n20183 )
         );
  MUX \u_a23_mem/U20159  ( .IN0(\u_a23_mem/n20150 ), .IN1(\u_a23_mem/n20135 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20151 ) );
  MUX \u_a23_mem/U20158  ( .IN0(\u_a23_mem/n20149 ), .IN1(\u_a23_mem/n20142 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20150 ) );
  MUX \u_a23_mem/U20157  ( .IN0(\u_a23_mem/n20148 ), .IN1(\u_a23_mem/n20145 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20149 ) );
  MUX \u_a23_mem/U20156  ( .IN0(\u_a23_mem/n20147 ), .IN1(\u_a23_mem/n20146 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20148 ) );
  MUX \u_a23_mem/U20155  ( .IN0(\u_a23_mem/p_mem[1][3] ), .IN1(
        \u_a23_mem/p_mem[65][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20147 )
         );
  MUX \u_a23_mem/U20154  ( .IN0(\u_a23_mem/p_mem[33][3] ), .IN1(
        \u_a23_mem/p_mem[97][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20146 )
         );
  MUX \u_a23_mem/U20153  ( .IN0(\u_a23_mem/n20144 ), .IN1(\u_a23_mem/n20143 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20145 ) );
  MUX \u_a23_mem/U20152  ( .IN0(\u_a23_mem/p_mem[17][3] ), .IN1(
        \u_a23_mem/p_mem[81][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20144 )
         );
  MUX \u_a23_mem/U20151  ( .IN0(\u_a23_mem/p_mem[49][3] ), .IN1(
        \u_a23_mem/p_mem[113][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20143 )
         );
  MUX \u_a23_mem/U20150  ( .IN0(\u_a23_mem/n20141 ), .IN1(\u_a23_mem/n20138 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20142 ) );
  MUX \u_a23_mem/U20149  ( .IN0(\u_a23_mem/n20140 ), .IN1(\u_a23_mem/n20139 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20141 ) );
  MUX \u_a23_mem/U20148  ( .IN0(\u_a23_mem/p_mem[9][3] ), .IN1(
        \u_a23_mem/p_mem[73][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20140 )
         );
  MUX \u_a23_mem/U20147  ( .IN0(\u_a23_mem/p_mem[41][3] ), .IN1(
        \u_a23_mem/p_mem[105][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20139 )
         );
  MUX \u_a23_mem/U20146  ( .IN0(\u_a23_mem/n20137 ), .IN1(\u_a23_mem/n20136 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20138 ) );
  MUX \u_a23_mem/U20145  ( .IN0(\u_a23_mem/p_mem[25][3] ), .IN1(
        \u_a23_mem/p_mem[89][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20137 )
         );
  MUX \u_a23_mem/U20144  ( .IN0(\u_a23_mem/p_mem[57][3] ), .IN1(
        \u_a23_mem/p_mem[121][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20136 )
         );
  MUX \u_a23_mem/U20143  ( .IN0(\u_a23_mem/n20134 ), .IN1(\u_a23_mem/n20127 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20135 ) );
  MUX \u_a23_mem/U20142  ( .IN0(\u_a23_mem/n20133 ), .IN1(\u_a23_mem/n20130 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20134 ) );
  MUX \u_a23_mem/U20141  ( .IN0(\u_a23_mem/n20132 ), .IN1(\u_a23_mem/n20131 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20133 ) );
  MUX \u_a23_mem/U20140  ( .IN0(\u_a23_mem/p_mem[5][3] ), .IN1(
        \u_a23_mem/p_mem[69][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20132 )
         );
  MUX \u_a23_mem/U20139  ( .IN0(\u_a23_mem/p_mem[37][3] ), .IN1(
        \u_a23_mem/p_mem[101][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20131 )
         );
  MUX \u_a23_mem/U20138  ( .IN0(\u_a23_mem/n20129 ), .IN1(\u_a23_mem/n20128 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20130 ) );
  MUX \u_a23_mem/U20137  ( .IN0(\u_a23_mem/p_mem[21][3] ), .IN1(
        \u_a23_mem/p_mem[85][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20129 )
         );
  MUX \u_a23_mem/U20136  ( .IN0(\u_a23_mem/p_mem[53][3] ), .IN1(
        \u_a23_mem/p_mem[117][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20128 )
         );
  MUX \u_a23_mem/U20135  ( .IN0(\u_a23_mem/n20126 ), .IN1(\u_a23_mem/n20123 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20127 ) );
  MUX \u_a23_mem/U20134  ( .IN0(\u_a23_mem/n20125 ), .IN1(\u_a23_mem/n20124 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20126 ) );
  MUX \u_a23_mem/U20133  ( .IN0(\u_a23_mem/p_mem[13][3] ), .IN1(
        \u_a23_mem/p_mem[77][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20125 )
         );
  MUX \u_a23_mem/U20132  ( .IN0(\u_a23_mem/p_mem[45][3] ), .IN1(
        \u_a23_mem/p_mem[109][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20124 )
         );
  MUX \u_a23_mem/U20131  ( .IN0(\u_a23_mem/n20122 ), .IN1(\u_a23_mem/n20121 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20123 ) );
  MUX \u_a23_mem/U20130  ( .IN0(\u_a23_mem/p_mem[29][3] ), .IN1(
        \u_a23_mem/p_mem[93][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20122 )
         );
  MUX \u_a23_mem/U20129  ( .IN0(\u_a23_mem/p_mem[61][3] ), .IN1(
        \u_a23_mem/p_mem[125][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20121 )
         );
  MUX \u_a23_mem/U20128  ( .IN0(\u_a23_mem/n20119 ), .IN1(\u_a23_mem/n20104 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20120 ) );
  MUX \u_a23_mem/U20127  ( .IN0(\u_a23_mem/n20118 ), .IN1(\u_a23_mem/n20111 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20119 ) );
  MUX \u_a23_mem/U20126  ( .IN0(\u_a23_mem/n20117 ), .IN1(\u_a23_mem/n20114 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20118 ) );
  MUX \u_a23_mem/U20125  ( .IN0(\u_a23_mem/n20116 ), .IN1(\u_a23_mem/n20115 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20117 ) );
  MUX \u_a23_mem/U20124  ( .IN0(\u_a23_mem/p_mem[3][3] ), .IN1(
        \u_a23_mem/p_mem[67][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20116 )
         );
  MUX \u_a23_mem/U20123  ( .IN0(\u_a23_mem/p_mem[35][3] ), .IN1(
        \u_a23_mem/p_mem[99][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20115 )
         );
  MUX \u_a23_mem/U20122  ( .IN0(\u_a23_mem/n20113 ), .IN1(\u_a23_mem/n20112 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20114 ) );
  MUX \u_a23_mem/U20121  ( .IN0(\u_a23_mem/p_mem[19][3] ), .IN1(
        \u_a23_mem/p_mem[83][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20113 )
         );
  MUX \u_a23_mem/U20120  ( .IN0(\u_a23_mem/p_mem[51][3] ), .IN1(
        \u_a23_mem/p_mem[115][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20112 )
         );
  MUX \u_a23_mem/U20119  ( .IN0(\u_a23_mem/n20110 ), .IN1(\u_a23_mem/n20107 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20111 ) );
  MUX \u_a23_mem/U20118  ( .IN0(\u_a23_mem/n20109 ), .IN1(\u_a23_mem/n20108 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20110 ) );
  MUX \u_a23_mem/U20117  ( .IN0(\u_a23_mem/p_mem[11][3] ), .IN1(
        \u_a23_mem/p_mem[75][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20109 )
         );
  MUX \u_a23_mem/U20116  ( .IN0(\u_a23_mem/p_mem[43][3] ), .IN1(
        \u_a23_mem/p_mem[107][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20108 )
         );
  MUX \u_a23_mem/U20115  ( .IN0(\u_a23_mem/n20106 ), .IN1(\u_a23_mem/n20105 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20107 ) );
  MUX \u_a23_mem/U20114  ( .IN0(\u_a23_mem/p_mem[27][3] ), .IN1(
        \u_a23_mem/p_mem[91][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20106 )
         );
  MUX \u_a23_mem/U20113  ( .IN0(\u_a23_mem/p_mem[59][3] ), .IN1(
        \u_a23_mem/p_mem[123][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20105 )
         );
  MUX \u_a23_mem/U20112  ( .IN0(\u_a23_mem/n20103 ), .IN1(\u_a23_mem/n20096 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20104 ) );
  MUX \u_a23_mem/U20111  ( .IN0(\u_a23_mem/n20102 ), .IN1(\u_a23_mem/n20099 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20103 ) );
  MUX \u_a23_mem/U20110  ( .IN0(\u_a23_mem/n20101 ), .IN1(\u_a23_mem/n20100 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20102 ) );
  MUX \u_a23_mem/U20109  ( .IN0(\u_a23_mem/p_mem[7][3] ), .IN1(
        \u_a23_mem/p_mem[71][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20101 )
         );
  MUX \u_a23_mem/U20108  ( .IN0(\u_a23_mem/p_mem[39][3] ), .IN1(
        \u_a23_mem/p_mem[103][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20100 )
         );
  MUX \u_a23_mem/U20107  ( .IN0(\u_a23_mem/n20098 ), .IN1(\u_a23_mem/n20097 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20099 ) );
  MUX \u_a23_mem/U20106  ( .IN0(\u_a23_mem/p_mem[23][3] ), .IN1(
        \u_a23_mem/p_mem[87][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20098 )
         );
  MUX \u_a23_mem/U20105  ( .IN0(\u_a23_mem/p_mem[55][3] ), .IN1(
        \u_a23_mem/p_mem[119][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20097 )
         );
  MUX \u_a23_mem/U20104  ( .IN0(\u_a23_mem/n20095 ), .IN1(\u_a23_mem/n20092 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20096 ) );
  MUX \u_a23_mem/U20103  ( .IN0(\u_a23_mem/n20094 ), .IN1(\u_a23_mem/n20093 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20095 ) );
  MUX \u_a23_mem/U20102  ( .IN0(\u_a23_mem/p_mem[15][3] ), .IN1(
        \u_a23_mem/p_mem[79][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20094 )
         );
  MUX \u_a23_mem/U20101  ( .IN0(\u_a23_mem/p_mem[47][3] ), .IN1(
        \u_a23_mem/p_mem[111][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20093 )
         );
  MUX \u_a23_mem/U20100  ( .IN0(\u_a23_mem/n20091 ), .IN1(\u_a23_mem/n20090 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20092 ) );
  MUX \u_a23_mem/U20099  ( .IN0(\u_a23_mem/p_mem[31][3] ), .IN1(
        \u_a23_mem/p_mem[95][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20091 )
         );
  MUX \u_a23_mem/U20098  ( .IN0(\u_a23_mem/p_mem[63][3] ), .IN1(
        \u_a23_mem/p_mem[127][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20090 )
         );
  MUX \u_a23_mem/U20096  ( .IN0(\u_a23_mem/n20087 ), .IN1(\u_a23_mem/n20072 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20088 ) );
  MUX \u_a23_mem/U20095  ( .IN0(\u_a23_mem/n20086 ), .IN1(\u_a23_mem/n20079 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20087 ) );
  MUX \u_a23_mem/U20094  ( .IN0(\u_a23_mem/n20085 ), .IN1(\u_a23_mem/n20082 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20086 ) );
  MUX \u_a23_mem/U20093  ( .IN0(\u_a23_mem/n20084 ), .IN1(\u_a23_mem/n20083 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20085 ) );
  MUX \u_a23_mem/U20092  ( .IN0(\u_a23_mem/p_mem[2][3] ), .IN1(
        \u_a23_mem/p_mem[66][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20084 )
         );
  MUX \u_a23_mem/U20091  ( .IN0(\u_a23_mem/p_mem[34][3] ), .IN1(
        \u_a23_mem/p_mem[98][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20083 )
         );
  MUX \u_a23_mem/U20090  ( .IN0(\u_a23_mem/n20081 ), .IN1(\u_a23_mem/n20080 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20082 ) );
  MUX \u_a23_mem/U20089  ( .IN0(\u_a23_mem/p_mem[18][3] ), .IN1(
        \u_a23_mem/p_mem[82][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20081 )
         );
  MUX \u_a23_mem/U20088  ( .IN0(\u_a23_mem/p_mem[50][3] ), .IN1(
        \u_a23_mem/p_mem[114][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20080 )
         );
  MUX \u_a23_mem/U20087  ( .IN0(\u_a23_mem/n20078 ), .IN1(\u_a23_mem/n20075 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20079 ) );
  MUX \u_a23_mem/U20086  ( .IN0(\u_a23_mem/n20077 ), .IN1(\u_a23_mem/n20076 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20078 ) );
  MUX \u_a23_mem/U20085  ( .IN0(\u_a23_mem/p_mem[10][3] ), .IN1(
        \u_a23_mem/p_mem[74][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20077 )
         );
  MUX \u_a23_mem/U20084  ( .IN0(\u_a23_mem/p_mem[42][3] ), .IN1(
        \u_a23_mem/p_mem[106][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20076 )
         );
  MUX \u_a23_mem/U20083  ( .IN0(\u_a23_mem/n20074 ), .IN1(\u_a23_mem/n20073 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20075 ) );
  MUX \u_a23_mem/U20082  ( .IN0(\u_a23_mem/p_mem[26][3] ), .IN1(
        \u_a23_mem/p_mem[90][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20074 )
         );
  MUX \u_a23_mem/U20081  ( .IN0(\u_a23_mem/p_mem[58][3] ), .IN1(
        \u_a23_mem/p_mem[122][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20073 )
         );
  MUX \u_a23_mem/U20080  ( .IN0(\u_a23_mem/n20071 ), .IN1(\u_a23_mem/n20064 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20072 ) );
  MUX \u_a23_mem/U20079  ( .IN0(\u_a23_mem/n20070 ), .IN1(\u_a23_mem/n20067 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20071 ) );
  MUX \u_a23_mem/U20078  ( .IN0(\u_a23_mem/n20069 ), .IN1(\u_a23_mem/n20068 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20070 ) );
  MUX \u_a23_mem/U20077  ( .IN0(\u_a23_mem/p_mem[6][3] ), .IN1(
        \u_a23_mem/p_mem[70][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20069 )
         );
  MUX \u_a23_mem/U20076  ( .IN0(\u_a23_mem/p_mem[38][3] ), .IN1(
        \u_a23_mem/p_mem[102][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20068 )
         );
  MUX \u_a23_mem/U20075  ( .IN0(\u_a23_mem/n20066 ), .IN1(\u_a23_mem/n20065 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20067 ) );
  MUX \u_a23_mem/U20074  ( .IN0(\u_a23_mem/p_mem[22][3] ), .IN1(
        \u_a23_mem/p_mem[86][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20066 )
         );
  MUX \u_a23_mem/U20073  ( .IN0(\u_a23_mem/p_mem[54][3] ), .IN1(
        \u_a23_mem/p_mem[118][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20065 )
         );
  MUX \u_a23_mem/U20072  ( .IN0(\u_a23_mem/n20063 ), .IN1(\u_a23_mem/n20060 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20064 ) );
  MUX \u_a23_mem/U20071  ( .IN0(\u_a23_mem/n20062 ), .IN1(\u_a23_mem/n20061 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20063 ) );
  MUX \u_a23_mem/U20070  ( .IN0(\u_a23_mem/p_mem[14][3] ), .IN1(
        \u_a23_mem/p_mem[78][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20062 )
         );
  MUX \u_a23_mem/U20069  ( .IN0(\u_a23_mem/p_mem[46][3] ), .IN1(
        \u_a23_mem/p_mem[110][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20061 )
         );
  MUX \u_a23_mem/U20068  ( .IN0(\u_a23_mem/n20059 ), .IN1(\u_a23_mem/n20058 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20060 ) );
  MUX \u_a23_mem/U20067  ( .IN0(\u_a23_mem/p_mem[30][3] ), .IN1(
        \u_a23_mem/p_mem[94][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20059 )
         );
  MUX \u_a23_mem/U20066  ( .IN0(\u_a23_mem/p_mem[62][3] ), .IN1(
        \u_a23_mem/p_mem[126][3] ), .SEL(m_address[6]), .F(\u_a23_mem/n20058 )
         );
  MUX \u_a23_mem/U20033  ( .IN0(\u_a23_mem/n20025 ), .IN1(\u_a23_mem/n20010 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n20026 ) );
  MUX \u_a23_mem/U20032  ( .IN0(\u_a23_mem/n20024 ), .IN1(\u_a23_mem/n20017 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20025 ) );
  MUX \u_a23_mem/U20031  ( .IN0(\u_a23_mem/n20023 ), .IN1(\u_a23_mem/n20020 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20024 ) );
  MUX \u_a23_mem/U20030  ( .IN0(\u_a23_mem/n20022 ), .IN1(\u_a23_mem/n20021 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20023 ) );
  MUX \u_a23_mem/U20029  ( .IN0(\u_a23_mem/p_mem[1][2] ), .IN1(
        \u_a23_mem/p_mem[65][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n20022 )
         );
  MUX \u_a23_mem/U20028  ( .IN0(\u_a23_mem/p_mem[33][2] ), .IN1(
        \u_a23_mem/p_mem[97][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n20021 )
         );
  MUX \u_a23_mem/U20027  ( .IN0(\u_a23_mem/n20019 ), .IN1(\u_a23_mem/n20018 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20020 ) );
  MUX \u_a23_mem/U20026  ( .IN0(\u_a23_mem/p_mem[17][2] ), .IN1(
        \u_a23_mem/p_mem[81][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n20019 )
         );
  MUX \u_a23_mem/U20025  ( .IN0(\u_a23_mem/p_mem[49][2] ), .IN1(
        \u_a23_mem/p_mem[113][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n20018 )
         );
  MUX \u_a23_mem/U20024  ( .IN0(\u_a23_mem/n20016 ), .IN1(\u_a23_mem/n20013 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20017 ) );
  MUX \u_a23_mem/U20023  ( .IN0(\u_a23_mem/n20015 ), .IN1(\u_a23_mem/n20014 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20016 ) );
  MUX \u_a23_mem/U20022  ( .IN0(\u_a23_mem/p_mem[9][2] ), .IN1(
        \u_a23_mem/p_mem[73][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n20015 )
         );
  MUX \u_a23_mem/U20021  ( .IN0(\u_a23_mem/p_mem[41][2] ), .IN1(
        \u_a23_mem/p_mem[105][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n20014 )
         );
  MUX \u_a23_mem/U20020  ( .IN0(\u_a23_mem/n20012 ), .IN1(\u_a23_mem/n20011 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20013 ) );
  MUX \u_a23_mem/U20019  ( .IN0(\u_a23_mem/p_mem[25][2] ), .IN1(
        \u_a23_mem/p_mem[89][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n20012 )
         );
  MUX \u_a23_mem/U20018  ( .IN0(\u_a23_mem/p_mem[57][2] ), .IN1(
        \u_a23_mem/p_mem[121][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n20011 )
         );
  MUX \u_a23_mem/U20017  ( .IN0(\u_a23_mem/n20009 ), .IN1(\u_a23_mem/n20002 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n20010 ) );
  MUX \u_a23_mem/U20016  ( .IN0(\u_a23_mem/n20008 ), .IN1(\u_a23_mem/n20005 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20009 ) );
  MUX \u_a23_mem/U20015  ( .IN0(\u_a23_mem/n20007 ), .IN1(\u_a23_mem/n20006 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20008 ) );
  MUX \u_a23_mem/U20014  ( .IN0(\u_a23_mem/p_mem[5][2] ), .IN1(
        \u_a23_mem/p_mem[69][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n20007 )
         );
  MUX \u_a23_mem/U20013  ( .IN0(\u_a23_mem/p_mem[37][2] ), .IN1(
        \u_a23_mem/p_mem[101][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n20006 )
         );
  MUX \u_a23_mem/U20012  ( .IN0(\u_a23_mem/n20004 ), .IN1(\u_a23_mem/n20003 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20005 ) );
  MUX \u_a23_mem/U20011  ( .IN0(\u_a23_mem/p_mem[21][2] ), .IN1(
        \u_a23_mem/p_mem[85][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n20004 )
         );
  MUX \u_a23_mem/U20010  ( .IN0(\u_a23_mem/p_mem[53][2] ), .IN1(
        \u_a23_mem/p_mem[117][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n20003 )
         );
  MUX \u_a23_mem/U20009  ( .IN0(\u_a23_mem/n20001 ), .IN1(\u_a23_mem/n19998 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n20002 ) );
  MUX \u_a23_mem/U20008  ( .IN0(\u_a23_mem/n20000 ), .IN1(\u_a23_mem/n19999 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n20001 ) );
  MUX \u_a23_mem/U20007  ( .IN0(\u_a23_mem/p_mem[13][2] ), .IN1(
        \u_a23_mem/p_mem[77][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n20000 )
         );
  MUX \u_a23_mem/U20006  ( .IN0(\u_a23_mem/p_mem[45][2] ), .IN1(
        \u_a23_mem/p_mem[109][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19999 )
         );
  MUX \u_a23_mem/U20005  ( .IN0(\u_a23_mem/n19997 ), .IN1(\u_a23_mem/n19996 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19998 ) );
  MUX \u_a23_mem/U20004  ( .IN0(\u_a23_mem/p_mem[29][2] ), .IN1(
        \u_a23_mem/p_mem[93][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19997 )
         );
  MUX \u_a23_mem/U20003  ( .IN0(\u_a23_mem/p_mem[61][2] ), .IN1(
        \u_a23_mem/p_mem[125][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19996 )
         );
  MUX \u_a23_mem/U20002  ( .IN0(\u_a23_mem/n19994 ), .IN1(\u_a23_mem/n19979 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n19995 ) );
  MUX \u_a23_mem/U20001  ( .IN0(\u_a23_mem/n19993 ), .IN1(\u_a23_mem/n19986 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n19994 ) );
  MUX \u_a23_mem/U20000  ( .IN0(\u_a23_mem/n19992 ), .IN1(\u_a23_mem/n19989 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n19993 ) );
  MUX \u_a23_mem/U19999  ( .IN0(\u_a23_mem/n19991 ), .IN1(\u_a23_mem/n19990 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19992 ) );
  MUX \u_a23_mem/U19998  ( .IN0(\u_a23_mem/p_mem[3][2] ), .IN1(
        \u_a23_mem/p_mem[67][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19991 )
         );
  MUX \u_a23_mem/U19997  ( .IN0(\u_a23_mem/p_mem[35][2] ), .IN1(
        \u_a23_mem/p_mem[99][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19990 )
         );
  MUX \u_a23_mem/U19996  ( .IN0(\u_a23_mem/n19988 ), .IN1(\u_a23_mem/n19987 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19989 ) );
  MUX \u_a23_mem/U19995  ( .IN0(\u_a23_mem/p_mem[19][2] ), .IN1(
        \u_a23_mem/p_mem[83][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19988 )
         );
  MUX \u_a23_mem/U19994  ( .IN0(\u_a23_mem/p_mem[51][2] ), .IN1(
        \u_a23_mem/p_mem[115][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19987 )
         );
  MUX \u_a23_mem/U19993  ( .IN0(\u_a23_mem/n19985 ), .IN1(\u_a23_mem/n19982 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n19986 ) );
  MUX \u_a23_mem/U19992  ( .IN0(\u_a23_mem/n19984 ), .IN1(\u_a23_mem/n19983 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19985 ) );
  MUX \u_a23_mem/U19991  ( .IN0(\u_a23_mem/p_mem[11][2] ), .IN1(
        \u_a23_mem/p_mem[75][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19984 )
         );
  MUX \u_a23_mem/U19990  ( .IN0(\u_a23_mem/p_mem[43][2] ), .IN1(
        \u_a23_mem/p_mem[107][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19983 )
         );
  MUX \u_a23_mem/U19989  ( .IN0(\u_a23_mem/n19981 ), .IN1(\u_a23_mem/n19980 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19982 ) );
  MUX \u_a23_mem/U19988  ( .IN0(\u_a23_mem/p_mem[27][2] ), .IN1(
        \u_a23_mem/p_mem[91][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19981 )
         );
  MUX \u_a23_mem/U19987  ( .IN0(\u_a23_mem/p_mem[59][2] ), .IN1(
        \u_a23_mem/p_mem[123][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19980 )
         );
  MUX \u_a23_mem/U19986  ( .IN0(\u_a23_mem/n19978 ), .IN1(\u_a23_mem/n19971 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n19979 ) );
  MUX \u_a23_mem/U19985  ( .IN0(\u_a23_mem/n19977 ), .IN1(\u_a23_mem/n19974 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n19978 ) );
  MUX \u_a23_mem/U19984  ( .IN0(\u_a23_mem/n19976 ), .IN1(\u_a23_mem/n19975 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19977 ) );
  MUX \u_a23_mem/U19983  ( .IN0(\u_a23_mem/p_mem[7][2] ), .IN1(
        \u_a23_mem/p_mem[71][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19976 )
         );
  MUX \u_a23_mem/U19982  ( .IN0(\u_a23_mem/p_mem[39][2] ), .IN1(
        \u_a23_mem/p_mem[103][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19975 )
         );
  MUX \u_a23_mem/U19981  ( .IN0(\u_a23_mem/n19973 ), .IN1(\u_a23_mem/n19972 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19974 ) );
  MUX \u_a23_mem/U19980  ( .IN0(\u_a23_mem/p_mem[23][2] ), .IN1(
        \u_a23_mem/p_mem[87][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19973 )
         );
  MUX \u_a23_mem/U19979  ( .IN0(\u_a23_mem/p_mem[55][2] ), .IN1(
        \u_a23_mem/p_mem[119][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19972 )
         );
  MUX \u_a23_mem/U19978  ( .IN0(\u_a23_mem/n19970 ), .IN1(\u_a23_mem/n19967 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n19971 ) );
  MUX \u_a23_mem/U19977  ( .IN0(\u_a23_mem/n19969 ), .IN1(\u_a23_mem/n19968 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19970 ) );
  MUX \u_a23_mem/U19976  ( .IN0(\u_a23_mem/p_mem[15][2] ), .IN1(
        \u_a23_mem/p_mem[79][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19969 )
         );
  MUX \u_a23_mem/U19975  ( .IN0(\u_a23_mem/p_mem[47][2] ), .IN1(
        \u_a23_mem/p_mem[111][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19968 )
         );
  MUX \u_a23_mem/U19974  ( .IN0(\u_a23_mem/n19966 ), .IN1(\u_a23_mem/n19965 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19967 ) );
  MUX \u_a23_mem/U19973  ( .IN0(\u_a23_mem/p_mem[31][2] ), .IN1(
        \u_a23_mem/p_mem[95][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19966 )
         );
  MUX \u_a23_mem/U19972  ( .IN0(\u_a23_mem/p_mem[63][2] ), .IN1(
        \u_a23_mem/p_mem[127][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19965 )
         );
  MUX \u_a23_mem/U19970  ( .IN0(\u_a23_mem/n19962 ), .IN1(\u_a23_mem/n19947 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n19963 ) );
  MUX \u_a23_mem/U19969  ( .IN0(\u_a23_mem/n19961 ), .IN1(\u_a23_mem/n19954 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n19962 ) );
  MUX \u_a23_mem/U19968  ( .IN0(\u_a23_mem/n19960 ), .IN1(\u_a23_mem/n19957 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n19961 ) );
  MUX \u_a23_mem/U19967  ( .IN0(\u_a23_mem/n19959 ), .IN1(\u_a23_mem/n19958 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19960 ) );
  MUX \u_a23_mem/U19966  ( .IN0(\u_a23_mem/p_mem[2][2] ), .IN1(
        \u_a23_mem/p_mem[66][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19959 )
         );
  MUX \u_a23_mem/U19965  ( .IN0(\u_a23_mem/p_mem[34][2] ), .IN1(
        \u_a23_mem/p_mem[98][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19958 )
         );
  MUX \u_a23_mem/U19964  ( .IN0(\u_a23_mem/n19956 ), .IN1(\u_a23_mem/n19955 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19957 ) );
  MUX \u_a23_mem/U19963  ( .IN0(\u_a23_mem/p_mem[18][2] ), .IN1(
        \u_a23_mem/p_mem[82][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19956 )
         );
  MUX \u_a23_mem/U19962  ( .IN0(\u_a23_mem/p_mem[50][2] ), .IN1(
        \u_a23_mem/p_mem[114][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19955 )
         );
  MUX \u_a23_mem/U19961  ( .IN0(\u_a23_mem/n19953 ), .IN1(\u_a23_mem/n19950 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n19954 ) );
  MUX \u_a23_mem/U19960  ( .IN0(\u_a23_mem/n19952 ), .IN1(\u_a23_mem/n19951 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19953 ) );
  MUX \u_a23_mem/U19959  ( .IN0(\u_a23_mem/p_mem[10][2] ), .IN1(
        \u_a23_mem/p_mem[74][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19952 )
         );
  MUX \u_a23_mem/U19958  ( .IN0(\u_a23_mem/p_mem[42][2] ), .IN1(
        \u_a23_mem/p_mem[106][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19951 )
         );
  MUX \u_a23_mem/U19957  ( .IN0(\u_a23_mem/n19949 ), .IN1(\u_a23_mem/n19948 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19950 ) );
  MUX \u_a23_mem/U19956  ( .IN0(\u_a23_mem/p_mem[26][2] ), .IN1(
        \u_a23_mem/p_mem[90][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19949 )
         );
  MUX \u_a23_mem/U19955  ( .IN0(\u_a23_mem/p_mem[58][2] ), .IN1(
        \u_a23_mem/p_mem[122][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19948 )
         );
  MUX \u_a23_mem/U19954  ( .IN0(\u_a23_mem/n19946 ), .IN1(\u_a23_mem/n19939 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n19947 ) );
  MUX \u_a23_mem/U19953  ( .IN0(\u_a23_mem/n19945 ), .IN1(\u_a23_mem/n19942 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n19946 ) );
  MUX \u_a23_mem/U19952  ( .IN0(\u_a23_mem/n19944 ), .IN1(\u_a23_mem/n19943 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19945 ) );
  MUX \u_a23_mem/U19951  ( .IN0(\u_a23_mem/p_mem[6][2] ), .IN1(
        \u_a23_mem/p_mem[70][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19944 )
         );
  MUX \u_a23_mem/U19950  ( .IN0(\u_a23_mem/p_mem[38][2] ), .IN1(
        \u_a23_mem/p_mem[102][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19943 )
         );
  MUX \u_a23_mem/U19949  ( .IN0(\u_a23_mem/n19941 ), .IN1(\u_a23_mem/n19940 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19942 ) );
  MUX \u_a23_mem/U19948  ( .IN0(\u_a23_mem/p_mem[22][2] ), .IN1(
        \u_a23_mem/p_mem[86][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19941 )
         );
  MUX \u_a23_mem/U19947  ( .IN0(\u_a23_mem/p_mem[54][2] ), .IN1(
        \u_a23_mem/p_mem[118][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19940 )
         );
  MUX \u_a23_mem/U19946  ( .IN0(\u_a23_mem/n19938 ), .IN1(\u_a23_mem/n19935 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n19939 ) );
  MUX \u_a23_mem/U19945  ( .IN0(\u_a23_mem/n19937 ), .IN1(\u_a23_mem/n19936 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19938 ) );
  MUX \u_a23_mem/U19944  ( .IN0(\u_a23_mem/p_mem[14][2] ), .IN1(
        \u_a23_mem/p_mem[78][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19937 )
         );
  MUX \u_a23_mem/U19943  ( .IN0(\u_a23_mem/p_mem[46][2] ), .IN1(
        \u_a23_mem/p_mem[110][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19936 )
         );
  MUX \u_a23_mem/U19942  ( .IN0(\u_a23_mem/n19934 ), .IN1(\u_a23_mem/n19933 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19935 ) );
  MUX \u_a23_mem/U19941  ( .IN0(\u_a23_mem/p_mem[30][2] ), .IN1(
        \u_a23_mem/p_mem[94][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19934 )
         );
  MUX \u_a23_mem/U19940  ( .IN0(\u_a23_mem/p_mem[62][2] ), .IN1(
        \u_a23_mem/p_mem[126][2] ), .SEL(m_address[6]), .F(\u_a23_mem/n19933 )
         );
  MUX \u_a23_mem/U19907  ( .IN0(\u_a23_mem/n19900 ), .IN1(\u_a23_mem/n19885 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n19901 ) );
  MUX \u_a23_mem/U19906  ( .IN0(\u_a23_mem/n19899 ), .IN1(\u_a23_mem/n19892 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n19900 ) );
  MUX \u_a23_mem/U19905  ( .IN0(\u_a23_mem/n19898 ), .IN1(\u_a23_mem/n19895 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n19899 ) );
  MUX \u_a23_mem/U19904  ( .IN0(\u_a23_mem/n19897 ), .IN1(\u_a23_mem/n19896 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19898 ) );
  MUX \u_a23_mem/U19903  ( .IN0(\u_a23_mem/p_mem[1][1] ), .IN1(
        \u_a23_mem/p_mem[65][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19897 )
         );
  MUX \u_a23_mem/U19902  ( .IN0(\u_a23_mem/p_mem[33][1] ), .IN1(
        \u_a23_mem/p_mem[97][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19896 )
         );
  MUX \u_a23_mem/U19901  ( .IN0(\u_a23_mem/n19894 ), .IN1(\u_a23_mem/n19893 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19895 ) );
  MUX \u_a23_mem/U19900  ( .IN0(\u_a23_mem/p_mem[17][1] ), .IN1(
        \u_a23_mem/p_mem[81][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19894 )
         );
  MUX \u_a23_mem/U19899  ( .IN0(\u_a23_mem/p_mem[49][1] ), .IN1(
        \u_a23_mem/p_mem[113][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19893 )
         );
  MUX \u_a23_mem/U19898  ( .IN0(\u_a23_mem/n19891 ), .IN1(\u_a23_mem/n19888 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n19892 ) );
  MUX \u_a23_mem/U19897  ( .IN0(\u_a23_mem/n19890 ), .IN1(\u_a23_mem/n19889 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19891 ) );
  MUX \u_a23_mem/U19896  ( .IN0(\u_a23_mem/p_mem[9][1] ), .IN1(
        \u_a23_mem/p_mem[73][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19890 )
         );
  MUX \u_a23_mem/U19895  ( .IN0(\u_a23_mem/p_mem[41][1] ), .IN1(
        \u_a23_mem/p_mem[105][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19889 )
         );
  MUX \u_a23_mem/U19894  ( .IN0(\u_a23_mem/n19887 ), .IN1(\u_a23_mem/n19886 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19888 ) );
  MUX \u_a23_mem/U19893  ( .IN0(\u_a23_mem/p_mem[25][1] ), .IN1(
        \u_a23_mem/p_mem[89][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19887 )
         );
  MUX \u_a23_mem/U19892  ( .IN0(\u_a23_mem/p_mem[57][1] ), .IN1(
        \u_a23_mem/p_mem[121][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19886 )
         );
  MUX \u_a23_mem/U19891  ( .IN0(\u_a23_mem/n19884 ), .IN1(\u_a23_mem/n19877 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n19885 ) );
  MUX \u_a23_mem/U19890  ( .IN0(\u_a23_mem/n19883 ), .IN1(\u_a23_mem/n19880 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n19884 ) );
  MUX \u_a23_mem/U19889  ( .IN0(\u_a23_mem/n19882 ), .IN1(\u_a23_mem/n19881 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19883 ) );
  MUX \u_a23_mem/U19888  ( .IN0(\u_a23_mem/p_mem[5][1] ), .IN1(
        \u_a23_mem/p_mem[69][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19882 )
         );
  MUX \u_a23_mem/U19887  ( .IN0(\u_a23_mem/p_mem[37][1] ), .IN1(
        \u_a23_mem/p_mem[101][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19881 )
         );
  MUX \u_a23_mem/U19886  ( .IN0(\u_a23_mem/n19879 ), .IN1(\u_a23_mem/n19878 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19880 ) );
  MUX \u_a23_mem/U19885  ( .IN0(\u_a23_mem/p_mem[21][1] ), .IN1(
        \u_a23_mem/p_mem[85][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19879 )
         );
  MUX \u_a23_mem/U19884  ( .IN0(\u_a23_mem/p_mem[53][1] ), .IN1(
        \u_a23_mem/p_mem[117][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19878 )
         );
  MUX \u_a23_mem/U19883  ( .IN0(\u_a23_mem/n19876 ), .IN1(\u_a23_mem/n19873 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n19877 ) );
  MUX \u_a23_mem/U19882  ( .IN0(\u_a23_mem/n19875 ), .IN1(\u_a23_mem/n19874 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19876 ) );
  MUX \u_a23_mem/U19881  ( .IN0(\u_a23_mem/p_mem[13][1] ), .IN1(
        \u_a23_mem/p_mem[77][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19875 )
         );
  MUX \u_a23_mem/U19880  ( .IN0(\u_a23_mem/p_mem[45][1] ), .IN1(
        \u_a23_mem/p_mem[109][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19874 )
         );
  MUX \u_a23_mem/U19879  ( .IN0(\u_a23_mem/n19872 ), .IN1(\u_a23_mem/n19871 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19873 ) );
  MUX \u_a23_mem/U19878  ( .IN0(\u_a23_mem/p_mem[29][1] ), .IN1(
        \u_a23_mem/p_mem[93][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19872 )
         );
  MUX \u_a23_mem/U19877  ( .IN0(\u_a23_mem/p_mem[61][1] ), .IN1(
        \u_a23_mem/p_mem[125][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19871 )
         );
  MUX \u_a23_mem/U19876  ( .IN0(\u_a23_mem/n19869 ), .IN1(\u_a23_mem/n19854 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n19870 ) );
  MUX \u_a23_mem/U19875  ( .IN0(\u_a23_mem/n19868 ), .IN1(\u_a23_mem/n19861 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n19869 ) );
  MUX \u_a23_mem/U19874  ( .IN0(\u_a23_mem/n19867 ), .IN1(\u_a23_mem/n19864 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n19868 ) );
  MUX \u_a23_mem/U19873  ( .IN0(\u_a23_mem/n19866 ), .IN1(\u_a23_mem/n19865 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19867 ) );
  MUX \u_a23_mem/U19872  ( .IN0(\u_a23_mem/p_mem[3][1] ), .IN1(
        \u_a23_mem/p_mem[67][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19866 )
         );
  MUX \u_a23_mem/U19871  ( .IN0(\u_a23_mem/p_mem[35][1] ), .IN1(
        \u_a23_mem/p_mem[99][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19865 )
         );
  MUX \u_a23_mem/U19870  ( .IN0(\u_a23_mem/n19863 ), .IN1(\u_a23_mem/n19862 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19864 ) );
  MUX \u_a23_mem/U19869  ( .IN0(\u_a23_mem/p_mem[19][1] ), .IN1(
        \u_a23_mem/p_mem[83][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19863 )
         );
  MUX \u_a23_mem/U19868  ( .IN0(\u_a23_mem/p_mem[51][1] ), .IN1(
        \u_a23_mem/p_mem[115][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19862 )
         );
  MUX \u_a23_mem/U19867  ( .IN0(\u_a23_mem/n19860 ), .IN1(\u_a23_mem/n19857 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n19861 ) );
  MUX \u_a23_mem/U19866  ( .IN0(\u_a23_mem/n19859 ), .IN1(\u_a23_mem/n19858 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19860 ) );
  MUX \u_a23_mem/U19865  ( .IN0(\u_a23_mem/p_mem[11][1] ), .IN1(
        \u_a23_mem/p_mem[75][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19859 )
         );
  MUX \u_a23_mem/U19864  ( .IN0(\u_a23_mem/p_mem[43][1] ), .IN1(
        \u_a23_mem/p_mem[107][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19858 )
         );
  MUX \u_a23_mem/U19863  ( .IN0(\u_a23_mem/n19856 ), .IN1(\u_a23_mem/n19855 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19857 ) );
  MUX \u_a23_mem/U19862  ( .IN0(\u_a23_mem/p_mem[27][1] ), .IN1(
        \u_a23_mem/p_mem[91][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19856 )
         );
  MUX \u_a23_mem/U19861  ( .IN0(\u_a23_mem/p_mem[59][1] ), .IN1(
        \u_a23_mem/p_mem[123][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19855 )
         );
  MUX \u_a23_mem/U19860  ( .IN0(\u_a23_mem/n19853 ), .IN1(\u_a23_mem/n19846 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n19854 ) );
  MUX \u_a23_mem/U19859  ( .IN0(\u_a23_mem/n19852 ), .IN1(\u_a23_mem/n19849 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n19853 ) );
  MUX \u_a23_mem/U19858  ( .IN0(\u_a23_mem/n19851 ), .IN1(\u_a23_mem/n19850 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19852 ) );
  MUX \u_a23_mem/U19857  ( .IN0(\u_a23_mem/p_mem[7][1] ), .IN1(
        \u_a23_mem/p_mem[71][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19851 )
         );
  MUX \u_a23_mem/U19856  ( .IN0(\u_a23_mem/p_mem[39][1] ), .IN1(
        \u_a23_mem/p_mem[103][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19850 )
         );
  MUX \u_a23_mem/U19855  ( .IN0(\u_a23_mem/n19848 ), .IN1(\u_a23_mem/n19847 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19849 ) );
  MUX \u_a23_mem/U19854  ( .IN0(\u_a23_mem/p_mem[23][1] ), .IN1(
        \u_a23_mem/p_mem[87][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19848 )
         );
  MUX \u_a23_mem/U19853  ( .IN0(\u_a23_mem/p_mem[55][1] ), .IN1(
        \u_a23_mem/p_mem[119][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19847 )
         );
  MUX \u_a23_mem/U19852  ( .IN0(\u_a23_mem/n19845 ), .IN1(\u_a23_mem/n19842 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n19846 ) );
  MUX \u_a23_mem/U19851  ( .IN0(\u_a23_mem/n19844 ), .IN1(\u_a23_mem/n19843 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19845 ) );
  MUX \u_a23_mem/U19850  ( .IN0(\u_a23_mem/p_mem[15][1] ), .IN1(
        \u_a23_mem/p_mem[79][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19844 )
         );
  MUX \u_a23_mem/U19849  ( .IN0(\u_a23_mem/p_mem[47][1] ), .IN1(
        \u_a23_mem/p_mem[111][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19843 )
         );
  MUX \u_a23_mem/U19848  ( .IN0(\u_a23_mem/n19841 ), .IN1(\u_a23_mem/n19840 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19842 ) );
  MUX \u_a23_mem/U19847  ( .IN0(\u_a23_mem/p_mem[31][1] ), .IN1(
        \u_a23_mem/p_mem[95][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19841 )
         );
  MUX \u_a23_mem/U19846  ( .IN0(\u_a23_mem/p_mem[63][1] ), .IN1(
        \u_a23_mem/p_mem[127][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19840 )
         );
  MUX \u_a23_mem/U19844  ( .IN0(\u_a23_mem/n19837 ), .IN1(\u_a23_mem/n19822 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n19838 ) );
  MUX \u_a23_mem/U19843  ( .IN0(\u_a23_mem/n19836 ), .IN1(\u_a23_mem/n19829 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n19837 ) );
  MUX \u_a23_mem/U19842  ( .IN0(\u_a23_mem/n19835 ), .IN1(\u_a23_mem/n19832 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n19836 ) );
  MUX \u_a23_mem/U19841  ( .IN0(\u_a23_mem/n19834 ), .IN1(\u_a23_mem/n19833 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19835 ) );
  MUX \u_a23_mem/U19840  ( .IN0(\u_a23_mem/p_mem[2][1] ), .IN1(
        \u_a23_mem/p_mem[66][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19834 )
         );
  MUX \u_a23_mem/U19839  ( .IN0(\u_a23_mem/p_mem[34][1] ), .IN1(
        \u_a23_mem/p_mem[98][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19833 )
         );
  MUX \u_a23_mem/U19838  ( .IN0(\u_a23_mem/n19831 ), .IN1(\u_a23_mem/n19830 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19832 ) );
  MUX \u_a23_mem/U19837  ( .IN0(\u_a23_mem/p_mem[18][1] ), .IN1(
        \u_a23_mem/p_mem[82][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19831 )
         );
  MUX \u_a23_mem/U19836  ( .IN0(\u_a23_mem/p_mem[50][1] ), .IN1(
        \u_a23_mem/p_mem[114][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19830 )
         );
  MUX \u_a23_mem/U19835  ( .IN0(\u_a23_mem/n19828 ), .IN1(\u_a23_mem/n19825 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n19829 ) );
  MUX \u_a23_mem/U19834  ( .IN0(\u_a23_mem/n19827 ), .IN1(\u_a23_mem/n19826 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19828 ) );
  MUX \u_a23_mem/U19833  ( .IN0(\u_a23_mem/p_mem[10][1] ), .IN1(
        \u_a23_mem/p_mem[74][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19827 )
         );
  MUX \u_a23_mem/U19832  ( .IN0(\u_a23_mem/p_mem[42][1] ), .IN1(
        \u_a23_mem/p_mem[106][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19826 )
         );
  MUX \u_a23_mem/U19831  ( .IN0(\u_a23_mem/n19824 ), .IN1(\u_a23_mem/n19823 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19825 ) );
  MUX \u_a23_mem/U19830  ( .IN0(\u_a23_mem/p_mem[26][1] ), .IN1(
        \u_a23_mem/p_mem[90][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19824 )
         );
  MUX \u_a23_mem/U19829  ( .IN0(\u_a23_mem/p_mem[58][1] ), .IN1(
        \u_a23_mem/p_mem[122][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19823 )
         );
  MUX \u_a23_mem/U19828  ( .IN0(\u_a23_mem/n19821 ), .IN1(\u_a23_mem/n19814 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n19822 ) );
  MUX \u_a23_mem/U19827  ( .IN0(\u_a23_mem/n19820 ), .IN1(\u_a23_mem/n19817 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n19821 ) );
  MUX \u_a23_mem/U19826  ( .IN0(\u_a23_mem/n19819 ), .IN1(\u_a23_mem/n19818 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19820 ) );
  MUX \u_a23_mem/U19825  ( .IN0(\u_a23_mem/p_mem[6][1] ), .IN1(
        \u_a23_mem/p_mem[70][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19819 )
         );
  MUX \u_a23_mem/U19824  ( .IN0(\u_a23_mem/p_mem[38][1] ), .IN1(
        \u_a23_mem/p_mem[102][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19818 )
         );
  MUX \u_a23_mem/U19823  ( .IN0(\u_a23_mem/n19816 ), .IN1(\u_a23_mem/n19815 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19817 ) );
  MUX \u_a23_mem/U19822  ( .IN0(\u_a23_mem/p_mem[22][1] ), .IN1(
        \u_a23_mem/p_mem[86][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19816 )
         );
  MUX \u_a23_mem/U19821  ( .IN0(\u_a23_mem/p_mem[54][1] ), .IN1(
        \u_a23_mem/p_mem[118][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19815 )
         );
  MUX \u_a23_mem/U19820  ( .IN0(\u_a23_mem/n19813 ), .IN1(\u_a23_mem/n19810 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n19814 ) );
  MUX \u_a23_mem/U19819  ( .IN0(\u_a23_mem/n19812 ), .IN1(\u_a23_mem/n19811 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19813 ) );
  MUX \u_a23_mem/U19818  ( .IN0(\u_a23_mem/p_mem[14][1] ), .IN1(
        \u_a23_mem/p_mem[78][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19812 )
         );
  MUX \u_a23_mem/U19817  ( .IN0(\u_a23_mem/p_mem[46][1] ), .IN1(
        \u_a23_mem/p_mem[110][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19811 )
         );
  MUX \u_a23_mem/U19816  ( .IN0(\u_a23_mem/n19809 ), .IN1(\u_a23_mem/n19808 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19810 ) );
  MUX \u_a23_mem/U19815  ( .IN0(\u_a23_mem/p_mem[30][1] ), .IN1(
        \u_a23_mem/p_mem[94][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19809 )
         );
  MUX \u_a23_mem/U19814  ( .IN0(\u_a23_mem/p_mem[62][1] ), .IN1(
        \u_a23_mem/p_mem[126][1] ), .SEL(m_address[6]), .F(\u_a23_mem/n19808 )
         );
  MUX \u_a23_mem/U19781  ( .IN0(\u_a23_mem/n19775 ), .IN1(\u_a23_mem/n19760 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n19776 ) );
  MUX \u_a23_mem/U19780  ( .IN0(\u_a23_mem/n19774 ), .IN1(\u_a23_mem/n19767 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n19775 ) );
  MUX \u_a23_mem/U19779  ( .IN0(\u_a23_mem/n19773 ), .IN1(\u_a23_mem/n19770 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n19774 ) );
  MUX \u_a23_mem/U19778  ( .IN0(\u_a23_mem/n19772 ), .IN1(\u_a23_mem/n19771 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19773 ) );
  MUX \u_a23_mem/U19777  ( .IN0(\u_a23_mem/p_mem[1][0] ), .IN1(
        \u_a23_mem/p_mem[65][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19772 )
         );
  MUX \u_a23_mem/U19776  ( .IN0(\u_a23_mem/p_mem[33][0] ), .IN1(
        \u_a23_mem/p_mem[97][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19771 )
         );
  MUX \u_a23_mem/U19775  ( .IN0(\u_a23_mem/n19769 ), .IN1(\u_a23_mem/n19768 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19770 ) );
  MUX \u_a23_mem/U19774  ( .IN0(\u_a23_mem/p_mem[17][0] ), .IN1(
        \u_a23_mem/p_mem[81][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19769 )
         );
  MUX \u_a23_mem/U19773  ( .IN0(\u_a23_mem/p_mem[49][0] ), .IN1(
        \u_a23_mem/p_mem[113][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19768 )
         );
  MUX \u_a23_mem/U19772  ( .IN0(\u_a23_mem/n19766 ), .IN1(\u_a23_mem/n19763 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n19767 ) );
  MUX \u_a23_mem/U19771  ( .IN0(\u_a23_mem/n19765 ), .IN1(\u_a23_mem/n19764 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19766 ) );
  MUX \u_a23_mem/U19770  ( .IN0(\u_a23_mem/p_mem[9][0] ), .IN1(
        \u_a23_mem/p_mem[73][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19765 )
         );
  MUX \u_a23_mem/U19769  ( .IN0(\u_a23_mem/p_mem[41][0] ), .IN1(
        \u_a23_mem/p_mem[105][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19764 )
         );
  MUX \u_a23_mem/U19768  ( .IN0(\u_a23_mem/n19762 ), .IN1(\u_a23_mem/n19761 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19763 ) );
  MUX \u_a23_mem/U19767  ( .IN0(\u_a23_mem/p_mem[25][0] ), .IN1(
        \u_a23_mem/p_mem[89][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19762 )
         );
  MUX \u_a23_mem/U19766  ( .IN0(\u_a23_mem/p_mem[57][0] ), .IN1(
        \u_a23_mem/p_mem[121][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19761 )
         );
  MUX \u_a23_mem/U19765  ( .IN0(\u_a23_mem/n19759 ), .IN1(\u_a23_mem/n19752 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n19760 ) );
  MUX \u_a23_mem/U19764  ( .IN0(\u_a23_mem/n19758 ), .IN1(\u_a23_mem/n19755 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n19759 ) );
  MUX \u_a23_mem/U19763  ( .IN0(\u_a23_mem/n19757 ), .IN1(\u_a23_mem/n19756 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19758 ) );
  MUX \u_a23_mem/U19762  ( .IN0(\u_a23_mem/p_mem[5][0] ), .IN1(
        \u_a23_mem/p_mem[69][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19757 )
         );
  MUX \u_a23_mem/U19761  ( .IN0(\u_a23_mem/p_mem[37][0] ), .IN1(
        \u_a23_mem/p_mem[101][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19756 )
         );
  MUX \u_a23_mem/U19760  ( .IN0(\u_a23_mem/n19754 ), .IN1(\u_a23_mem/n19753 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19755 ) );
  MUX \u_a23_mem/U19759  ( .IN0(\u_a23_mem/p_mem[21][0] ), .IN1(
        \u_a23_mem/p_mem[85][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19754 )
         );
  MUX \u_a23_mem/U19758  ( .IN0(\u_a23_mem/p_mem[53][0] ), .IN1(
        \u_a23_mem/p_mem[117][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19753 )
         );
  MUX \u_a23_mem/U19757  ( .IN0(\u_a23_mem/n19751 ), .IN1(\u_a23_mem/n19748 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n19752 ) );
  MUX \u_a23_mem/U19756  ( .IN0(\u_a23_mem/n19750 ), .IN1(\u_a23_mem/n19749 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19751 ) );
  MUX \u_a23_mem/U19755  ( .IN0(\u_a23_mem/p_mem[13][0] ), .IN1(
        \u_a23_mem/p_mem[77][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19750 )
         );
  MUX \u_a23_mem/U19754  ( .IN0(\u_a23_mem/p_mem[45][0] ), .IN1(
        \u_a23_mem/p_mem[109][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19749 )
         );
  MUX \u_a23_mem/U19753  ( .IN0(\u_a23_mem/n19747 ), .IN1(\u_a23_mem/n19746 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19748 ) );
  MUX \u_a23_mem/U19752  ( .IN0(\u_a23_mem/p_mem[29][0] ), .IN1(
        \u_a23_mem/p_mem[93][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19747 )
         );
  MUX \u_a23_mem/U19751  ( .IN0(\u_a23_mem/p_mem[61][0] ), .IN1(
        \u_a23_mem/p_mem[125][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19746 )
         );
  MUX \u_a23_mem/U19750  ( .IN0(\u_a23_mem/n19744 ), .IN1(\u_a23_mem/n19729 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n19745 ) );
  MUX \u_a23_mem/U19749  ( .IN0(\u_a23_mem/n19743 ), .IN1(\u_a23_mem/n19736 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n19744 ) );
  MUX \u_a23_mem/U19748  ( .IN0(\u_a23_mem/n19742 ), .IN1(\u_a23_mem/n19739 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n19743 ) );
  MUX \u_a23_mem/U19747  ( .IN0(\u_a23_mem/n19741 ), .IN1(\u_a23_mem/n19740 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19742 ) );
  MUX \u_a23_mem/U19746  ( .IN0(\u_a23_mem/p_mem[3][0] ), .IN1(
        \u_a23_mem/p_mem[67][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19741 )
         );
  MUX \u_a23_mem/U19745  ( .IN0(\u_a23_mem/p_mem[35][0] ), .IN1(
        \u_a23_mem/p_mem[99][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19740 )
         );
  MUX \u_a23_mem/U19744  ( .IN0(\u_a23_mem/n19738 ), .IN1(\u_a23_mem/n19737 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19739 ) );
  MUX \u_a23_mem/U19743  ( .IN0(\u_a23_mem/p_mem[19][0] ), .IN1(
        \u_a23_mem/p_mem[83][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19738 )
         );
  MUX \u_a23_mem/U19742  ( .IN0(\u_a23_mem/p_mem[51][0] ), .IN1(
        \u_a23_mem/p_mem[115][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19737 )
         );
  MUX \u_a23_mem/U19741  ( .IN0(\u_a23_mem/n19735 ), .IN1(\u_a23_mem/n19732 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n19736 ) );
  MUX \u_a23_mem/U19740  ( .IN0(\u_a23_mem/n19734 ), .IN1(\u_a23_mem/n19733 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19735 ) );
  MUX \u_a23_mem/U19739  ( .IN0(\u_a23_mem/p_mem[11][0] ), .IN1(
        \u_a23_mem/p_mem[75][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19734 )
         );
  MUX \u_a23_mem/U19738  ( .IN0(\u_a23_mem/p_mem[43][0] ), .IN1(
        \u_a23_mem/p_mem[107][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19733 )
         );
  MUX \u_a23_mem/U19737  ( .IN0(\u_a23_mem/n19731 ), .IN1(\u_a23_mem/n19730 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19732 ) );
  MUX \u_a23_mem/U19736  ( .IN0(\u_a23_mem/p_mem[27][0] ), .IN1(
        \u_a23_mem/p_mem[91][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19731 )
         );
  MUX \u_a23_mem/U19735  ( .IN0(\u_a23_mem/p_mem[59][0] ), .IN1(
        \u_a23_mem/p_mem[123][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19730 )
         );
  MUX \u_a23_mem/U19734  ( .IN0(\u_a23_mem/n19728 ), .IN1(\u_a23_mem/n19721 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n19729 ) );
  MUX \u_a23_mem/U19733  ( .IN0(\u_a23_mem/n19727 ), .IN1(\u_a23_mem/n19724 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n19728 ) );
  MUX \u_a23_mem/U19732  ( .IN0(\u_a23_mem/n19726 ), .IN1(\u_a23_mem/n19725 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19727 ) );
  MUX \u_a23_mem/U19731  ( .IN0(\u_a23_mem/p_mem[7][0] ), .IN1(
        \u_a23_mem/p_mem[71][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19726 )
         );
  MUX \u_a23_mem/U19730  ( .IN0(\u_a23_mem/p_mem[39][0] ), .IN1(
        \u_a23_mem/p_mem[103][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19725 )
         );
  MUX \u_a23_mem/U19729  ( .IN0(\u_a23_mem/n19723 ), .IN1(\u_a23_mem/n19722 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19724 ) );
  MUX \u_a23_mem/U19728  ( .IN0(\u_a23_mem/p_mem[23][0] ), .IN1(
        \u_a23_mem/p_mem[87][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19723 )
         );
  MUX \u_a23_mem/U19727  ( .IN0(\u_a23_mem/p_mem[55][0] ), .IN1(
        \u_a23_mem/p_mem[119][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19722 )
         );
  MUX \u_a23_mem/U19726  ( .IN0(\u_a23_mem/n19720 ), .IN1(\u_a23_mem/n19717 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n19721 ) );
  MUX \u_a23_mem/U19725  ( .IN0(\u_a23_mem/n19719 ), .IN1(\u_a23_mem/n19718 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19720 ) );
  MUX \u_a23_mem/U19724  ( .IN0(\u_a23_mem/p_mem[15][0] ), .IN1(
        \u_a23_mem/p_mem[79][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19719 )
         );
  MUX \u_a23_mem/U19723  ( .IN0(\u_a23_mem/p_mem[47][0] ), .IN1(
        \u_a23_mem/p_mem[111][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19718 )
         );
  MUX \u_a23_mem/U19722  ( .IN0(\u_a23_mem/n19716 ), .IN1(\u_a23_mem/n19715 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19717 ) );
  MUX \u_a23_mem/U19721  ( .IN0(\u_a23_mem/p_mem[31][0] ), .IN1(
        \u_a23_mem/p_mem[95][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19716 )
         );
  MUX \u_a23_mem/U19720  ( .IN0(\u_a23_mem/p_mem[63][0] ), .IN1(
        \u_a23_mem/p_mem[127][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19715 )
         );
  MUX \u_a23_mem/U19718  ( .IN0(\u_a23_mem/n19712 ), .IN1(\u_a23_mem/n19697 ), 
        .SEL(m_address[2]), .F(\u_a23_mem/n19713 ) );
  MUX \u_a23_mem/U19717  ( .IN0(\u_a23_mem/n19711 ), .IN1(\u_a23_mem/n19704 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n19712 ) );
  MUX \u_a23_mem/U19716  ( .IN0(\u_a23_mem/n19710 ), .IN1(\u_a23_mem/n19707 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n19711 ) );
  MUX \u_a23_mem/U19715  ( .IN0(\u_a23_mem/n19709 ), .IN1(\u_a23_mem/n19708 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19710 ) );
  MUX \u_a23_mem/U19714  ( .IN0(\u_a23_mem/p_mem[2][0] ), .IN1(
        \u_a23_mem/p_mem[66][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19709 )
         );
  MUX \u_a23_mem/U19713  ( .IN0(\u_a23_mem/p_mem[34][0] ), .IN1(
        \u_a23_mem/p_mem[98][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19708 )
         );
  MUX \u_a23_mem/U19712  ( .IN0(\u_a23_mem/n19706 ), .IN1(\u_a23_mem/n19705 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19707 ) );
  MUX \u_a23_mem/U19711  ( .IN0(\u_a23_mem/p_mem[18][0] ), .IN1(
        \u_a23_mem/p_mem[82][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19706 )
         );
  MUX \u_a23_mem/U19710  ( .IN0(\u_a23_mem/p_mem[50][0] ), .IN1(
        \u_a23_mem/p_mem[114][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19705 )
         );
  MUX \u_a23_mem/U19709  ( .IN0(\u_a23_mem/n19703 ), .IN1(\u_a23_mem/n19700 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n19704 ) );
  MUX \u_a23_mem/U19708  ( .IN0(\u_a23_mem/n19702 ), .IN1(\u_a23_mem/n19701 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19703 ) );
  MUX \u_a23_mem/U19707  ( .IN0(\u_a23_mem/p_mem[10][0] ), .IN1(
        \u_a23_mem/p_mem[74][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19702 )
         );
  MUX \u_a23_mem/U19706  ( .IN0(\u_a23_mem/p_mem[42][0] ), .IN1(
        \u_a23_mem/p_mem[106][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19701 )
         );
  MUX \u_a23_mem/U19705  ( .IN0(\u_a23_mem/n19699 ), .IN1(\u_a23_mem/n19698 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19700 ) );
  MUX \u_a23_mem/U19704  ( .IN0(\u_a23_mem/p_mem[26][0] ), .IN1(
        \u_a23_mem/p_mem[90][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19699 )
         );
  MUX \u_a23_mem/U19703  ( .IN0(\u_a23_mem/p_mem[58][0] ), .IN1(
        \u_a23_mem/p_mem[122][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19698 )
         );
  MUX \u_a23_mem/U19702  ( .IN0(\u_a23_mem/n19696 ), .IN1(\u_a23_mem/n19689 ), 
        .SEL(m_address[3]), .F(\u_a23_mem/n19697 ) );
  MUX \u_a23_mem/U19701  ( .IN0(\u_a23_mem/n19695 ), .IN1(\u_a23_mem/n19692 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n19696 ) );
  MUX \u_a23_mem/U19700  ( .IN0(\u_a23_mem/n19694 ), .IN1(\u_a23_mem/n19693 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19695 ) );
  MUX \u_a23_mem/U19699  ( .IN0(\u_a23_mem/p_mem[6][0] ), .IN1(
        \u_a23_mem/p_mem[70][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19694 )
         );
  MUX \u_a23_mem/U19698  ( .IN0(\u_a23_mem/p_mem[38][0] ), .IN1(
        \u_a23_mem/p_mem[102][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19693 )
         );
  MUX \u_a23_mem/U19697  ( .IN0(\u_a23_mem/n19691 ), .IN1(\u_a23_mem/n19690 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19692 ) );
  MUX \u_a23_mem/U19696  ( .IN0(\u_a23_mem/p_mem[22][0] ), .IN1(
        \u_a23_mem/p_mem[86][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19691 )
         );
  MUX \u_a23_mem/U19695  ( .IN0(\u_a23_mem/p_mem[54][0] ), .IN1(
        \u_a23_mem/p_mem[118][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19690 )
         );
  MUX \u_a23_mem/U19694  ( .IN0(\u_a23_mem/n19688 ), .IN1(\u_a23_mem/n19685 ), 
        .SEL(m_address[4]), .F(\u_a23_mem/n19689 ) );
  MUX \u_a23_mem/U19693  ( .IN0(\u_a23_mem/n19687 ), .IN1(\u_a23_mem/n19686 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19688 ) );
  MUX \u_a23_mem/U19692  ( .IN0(\u_a23_mem/p_mem[14][0] ), .IN1(
        \u_a23_mem/p_mem[78][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19687 )
         );
  MUX \u_a23_mem/U19691  ( .IN0(\u_a23_mem/p_mem[46][0] ), .IN1(
        \u_a23_mem/p_mem[110][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19686 )
         );
  MUX \u_a23_mem/U19690  ( .IN0(\u_a23_mem/n19684 ), .IN1(\u_a23_mem/n19683 ), 
        .SEL(m_address[5]), .F(\u_a23_mem/n19685 ) );
  MUX \u_a23_mem/U19689  ( .IN0(\u_a23_mem/p_mem[30][0] ), .IN1(
        \u_a23_mem/p_mem[94][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19684 )
         );
  MUX \u_a23_mem/U19688  ( .IN0(\u_a23_mem/p_mem[62][0] ), .IN1(
        \u_a23_mem/p_mem[126][0] ), .SEL(m_address[6]), .F(\u_a23_mem/n19683 )
         );
  DFF \u_a23_mem/out_mem_reg[0][0]  ( .D(\u_a23_mem/n18372 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[0]) );
  DFF \u_a23_mem/out_mem_reg[0][1]  ( .D(\u_a23_mem/n18371 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[1]) );
  DFF \u_a23_mem/out_mem_reg[0][2]  ( .D(\u_a23_mem/n18370 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[2]) );
  DFF \u_a23_mem/out_mem_reg[0][3]  ( .D(\u_a23_mem/n18369 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[3]) );
  DFF \u_a23_mem/out_mem_reg[0][4]  ( .D(\u_a23_mem/n18368 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[4]) );
  DFF \u_a23_mem/out_mem_reg[0][5]  ( .D(\u_a23_mem/n18367 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[5]) );
  DFF \u_a23_mem/out_mem_reg[0][6]  ( .D(\u_a23_mem/n18366 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[6]) );
  DFF \u_a23_mem/out_mem_reg[0][7]  ( .D(\u_a23_mem/n18365 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[7]) );
  DFF \u_a23_mem/out_mem_reg[1][0]  ( .D(\u_a23_mem/n18364 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[8]) );
  DFF \u_a23_mem/out_mem_reg[1][1]  ( .D(\u_a23_mem/n18363 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[9]) );
  DFF \u_a23_mem/out_mem_reg[1][2]  ( .D(\u_a23_mem/n18362 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[10]) );
  DFF \u_a23_mem/out_mem_reg[1][3]  ( .D(\u_a23_mem/n18361 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[11]) );
  DFF \u_a23_mem/out_mem_reg[1][4]  ( .D(\u_a23_mem/n18360 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[12]) );
  DFF \u_a23_mem/out_mem_reg[1][5]  ( .D(\u_a23_mem/n18359 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[13]) );
  DFF \u_a23_mem/out_mem_reg[1][6]  ( .D(\u_a23_mem/n18358 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[14]) );
  DFF \u_a23_mem/out_mem_reg[1][7]  ( .D(\u_a23_mem/n18357 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[15]) );
  DFF \u_a23_mem/out_mem_reg[2][0]  ( .D(\u_a23_mem/n18356 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[16]) );
  DFF \u_a23_mem/out_mem_reg[2][1]  ( .D(\u_a23_mem/n18355 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[17]) );
  DFF \u_a23_mem/out_mem_reg[2][2]  ( .D(\u_a23_mem/n18354 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[18]) );
  DFF \u_a23_mem/out_mem_reg[2][3]  ( .D(\u_a23_mem/n18353 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[19]) );
  DFF \u_a23_mem/out_mem_reg[2][4]  ( .D(\u_a23_mem/n18352 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[20]) );
  DFF \u_a23_mem/out_mem_reg[2][5]  ( .D(\u_a23_mem/n18351 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[21]) );
  DFF \u_a23_mem/out_mem_reg[2][6]  ( .D(\u_a23_mem/n18350 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[22]) );
  DFF \u_a23_mem/out_mem_reg[2][7]  ( .D(\u_a23_mem/n18349 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[23]) );
  DFF \u_a23_mem/out_mem_reg[3][0]  ( .D(\u_a23_mem/n18348 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[24]) );
  DFF \u_a23_mem/out_mem_reg[3][1]  ( .D(\u_a23_mem/n18347 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[25]) );
  DFF \u_a23_mem/out_mem_reg[3][2]  ( .D(\u_a23_mem/n18346 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[26]) );
  DFF \u_a23_mem/out_mem_reg[3][3]  ( .D(\u_a23_mem/n18345 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[27]) );
  DFF \u_a23_mem/out_mem_reg[3][4]  ( .D(\u_a23_mem/n18344 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[28]) );
  DFF \u_a23_mem/out_mem_reg[3][5]  ( .D(\u_a23_mem/n18343 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[29]) );
  DFF \u_a23_mem/out_mem_reg[3][6]  ( .D(\u_a23_mem/n18342 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[30]) );
  DFF \u_a23_mem/out_mem_reg[3][7]  ( .D(\u_a23_mem/n18341 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[31]) );
  DFF \u_a23_mem/out_mem_reg[4][0]  ( .D(\u_a23_mem/n18340 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[32]) );
  DFF \u_a23_mem/out_mem_reg[4][1]  ( .D(\u_a23_mem/n18339 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[33]) );
  DFF \u_a23_mem/out_mem_reg[4][2]  ( .D(\u_a23_mem/n18338 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[34]) );
  DFF \u_a23_mem/out_mem_reg[4][3]  ( .D(\u_a23_mem/n18337 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[35]) );
  DFF \u_a23_mem/out_mem_reg[4][4]  ( .D(\u_a23_mem/n18336 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[36]) );
  DFF \u_a23_mem/out_mem_reg[4][5]  ( .D(\u_a23_mem/n18335 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[37]) );
  DFF \u_a23_mem/out_mem_reg[4][6]  ( .D(\u_a23_mem/n18334 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[38]) );
  DFF \u_a23_mem/out_mem_reg[4][7]  ( .D(\u_a23_mem/n18333 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[39]) );
  DFF \u_a23_mem/out_mem_reg[5][0]  ( .D(\u_a23_mem/n18332 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[40]) );
  DFF \u_a23_mem/out_mem_reg[5][1]  ( .D(\u_a23_mem/n18331 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[41]) );
  DFF \u_a23_mem/out_mem_reg[5][2]  ( .D(\u_a23_mem/n18330 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[42]) );
  DFF \u_a23_mem/out_mem_reg[5][3]  ( .D(\u_a23_mem/n18329 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[43]) );
  DFF \u_a23_mem/out_mem_reg[5][4]  ( .D(\u_a23_mem/n18328 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[44]) );
  DFF \u_a23_mem/out_mem_reg[5][5]  ( .D(\u_a23_mem/n18327 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[45]) );
  DFF \u_a23_mem/out_mem_reg[5][6]  ( .D(\u_a23_mem/n18326 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[46]) );
  DFF \u_a23_mem/out_mem_reg[5][7]  ( .D(\u_a23_mem/n18325 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[47]) );
  DFF \u_a23_mem/out_mem_reg[6][0]  ( .D(\u_a23_mem/n18324 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[48]) );
  DFF \u_a23_mem/out_mem_reg[6][1]  ( .D(\u_a23_mem/n18323 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[49]) );
  DFF \u_a23_mem/out_mem_reg[6][2]  ( .D(\u_a23_mem/n18322 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[50]) );
  DFF \u_a23_mem/out_mem_reg[6][3]  ( .D(\u_a23_mem/n18321 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[51]) );
  DFF \u_a23_mem/out_mem_reg[6][4]  ( .D(\u_a23_mem/n18320 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[52]) );
  DFF \u_a23_mem/out_mem_reg[6][5]  ( .D(\u_a23_mem/n18319 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[53]) );
  DFF \u_a23_mem/out_mem_reg[6][6]  ( .D(\u_a23_mem/n18318 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[54]) );
  DFF \u_a23_mem/out_mem_reg[6][7]  ( .D(\u_a23_mem/n18317 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[55]) );
  DFF \u_a23_mem/out_mem_reg[7][0]  ( .D(\u_a23_mem/n18316 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[56]) );
  DFF \u_a23_mem/out_mem_reg[7][1]  ( .D(\u_a23_mem/n18315 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[57]) );
  DFF \u_a23_mem/out_mem_reg[7][2]  ( .D(\u_a23_mem/n18314 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[58]) );
  DFF \u_a23_mem/out_mem_reg[7][3]  ( .D(\u_a23_mem/n18313 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[59]) );
  DFF \u_a23_mem/out_mem_reg[7][4]  ( .D(\u_a23_mem/n18312 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[60]) );
  DFF \u_a23_mem/out_mem_reg[7][5]  ( .D(\u_a23_mem/n18311 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[61]) );
  DFF \u_a23_mem/out_mem_reg[7][6]  ( .D(\u_a23_mem/n18310 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[62]) );
  DFF \u_a23_mem/out_mem_reg[7][7]  ( .D(\u_a23_mem/n18309 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[63]) );
  DFF \u_a23_mem/out_mem_reg[8][0]  ( .D(\u_a23_mem/n18308 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[64]) );
  DFF \u_a23_mem/out_mem_reg[8][1]  ( .D(\u_a23_mem/n18307 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[65]) );
  DFF \u_a23_mem/out_mem_reg[8][2]  ( .D(\u_a23_mem/n18306 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[66]) );
  DFF \u_a23_mem/out_mem_reg[8][3]  ( .D(\u_a23_mem/n18305 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[67]) );
  DFF \u_a23_mem/out_mem_reg[8][4]  ( .D(\u_a23_mem/n18304 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[68]) );
  DFF \u_a23_mem/out_mem_reg[8][5]  ( .D(\u_a23_mem/n18303 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[69]) );
  DFF \u_a23_mem/out_mem_reg[8][6]  ( .D(\u_a23_mem/n18302 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[70]) );
  DFF \u_a23_mem/out_mem_reg[8][7]  ( .D(\u_a23_mem/n18301 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[71]) );
  DFF \u_a23_mem/out_mem_reg[9][0]  ( .D(\u_a23_mem/n18300 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[72]) );
  DFF \u_a23_mem/out_mem_reg[9][1]  ( .D(\u_a23_mem/n18299 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[73]) );
  DFF \u_a23_mem/out_mem_reg[9][2]  ( .D(\u_a23_mem/n18298 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[74]) );
  DFF \u_a23_mem/out_mem_reg[9][3]  ( .D(\u_a23_mem/n18297 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[75]) );
  DFF \u_a23_mem/out_mem_reg[9][4]  ( .D(\u_a23_mem/n18296 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[76]) );
  DFF \u_a23_mem/out_mem_reg[9][5]  ( .D(\u_a23_mem/n18295 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[77]) );
  DFF \u_a23_mem/out_mem_reg[9][6]  ( .D(\u_a23_mem/n18294 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[78]) );
  DFF \u_a23_mem/out_mem_reg[9][7]  ( .D(\u_a23_mem/n18293 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(o[79]) );
  DFF \u_a23_mem/out_mem_reg[10][0]  ( .D(\u_a23_mem/n18292 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[80]) );
  DFF \u_a23_mem/out_mem_reg[10][1]  ( .D(\u_a23_mem/n18291 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[81]) );
  DFF \u_a23_mem/out_mem_reg[10][2]  ( .D(\u_a23_mem/n18290 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[82]) );
  DFF \u_a23_mem/out_mem_reg[10][3]  ( .D(\u_a23_mem/n18289 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[83]) );
  DFF \u_a23_mem/out_mem_reg[10][4]  ( .D(\u_a23_mem/n18288 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[84]) );
  DFF \u_a23_mem/out_mem_reg[10][5]  ( .D(\u_a23_mem/n18287 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[85]) );
  DFF \u_a23_mem/out_mem_reg[10][6]  ( .D(\u_a23_mem/n18286 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[86]) );
  DFF \u_a23_mem/out_mem_reg[10][7]  ( .D(\u_a23_mem/n18285 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[87]) );
  DFF \u_a23_mem/out_mem_reg[11][0]  ( .D(\u_a23_mem/n18284 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[88]) );
  DFF \u_a23_mem/out_mem_reg[11][1]  ( .D(\u_a23_mem/n18283 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[89]) );
  DFF \u_a23_mem/out_mem_reg[11][2]  ( .D(\u_a23_mem/n18282 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[90]) );
  DFF \u_a23_mem/out_mem_reg[11][3]  ( .D(\u_a23_mem/n18281 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[91]) );
  DFF \u_a23_mem/out_mem_reg[11][4]  ( .D(\u_a23_mem/n18280 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[92]) );
  DFF \u_a23_mem/out_mem_reg[11][5]  ( .D(\u_a23_mem/n18279 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[93]) );
  DFF \u_a23_mem/out_mem_reg[11][6]  ( .D(\u_a23_mem/n18278 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[94]) );
  DFF \u_a23_mem/out_mem_reg[11][7]  ( .D(\u_a23_mem/n18277 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[95]) );
  DFF \u_a23_mem/out_mem_reg[12][0]  ( .D(\u_a23_mem/n18276 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[96]) );
  DFF \u_a23_mem/out_mem_reg[12][1]  ( .D(\u_a23_mem/n18275 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[97]) );
  DFF \u_a23_mem/out_mem_reg[12][2]  ( .D(\u_a23_mem/n18274 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[98]) );
  DFF \u_a23_mem/out_mem_reg[12][3]  ( .D(\u_a23_mem/n18273 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[99]) );
  DFF \u_a23_mem/out_mem_reg[12][4]  ( .D(\u_a23_mem/n18272 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[100]) );
  DFF \u_a23_mem/out_mem_reg[12][5]  ( .D(\u_a23_mem/n18271 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[101]) );
  DFF \u_a23_mem/out_mem_reg[12][6]  ( .D(\u_a23_mem/n18270 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[102]) );
  DFF \u_a23_mem/out_mem_reg[12][7]  ( .D(\u_a23_mem/n18269 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[103]) );
  DFF \u_a23_mem/out_mem_reg[13][0]  ( .D(\u_a23_mem/n18268 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[104]) );
  DFF \u_a23_mem/out_mem_reg[13][1]  ( .D(\u_a23_mem/n18267 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[105]) );
  DFF \u_a23_mem/out_mem_reg[13][2]  ( .D(\u_a23_mem/n18266 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[106]) );
  DFF \u_a23_mem/out_mem_reg[13][3]  ( .D(\u_a23_mem/n18265 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[107]) );
  DFF \u_a23_mem/out_mem_reg[13][4]  ( .D(\u_a23_mem/n18264 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[108]) );
  DFF \u_a23_mem/out_mem_reg[13][5]  ( .D(\u_a23_mem/n18263 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[109]) );
  DFF \u_a23_mem/out_mem_reg[13][6]  ( .D(\u_a23_mem/n18262 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[110]) );
  DFF \u_a23_mem/out_mem_reg[13][7]  ( .D(\u_a23_mem/n18261 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[111]) );
  DFF \u_a23_mem/out_mem_reg[14][0]  ( .D(\u_a23_mem/n18260 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[112]) );
  DFF \u_a23_mem/out_mem_reg[14][1]  ( .D(\u_a23_mem/n18259 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[113]) );
  DFF \u_a23_mem/out_mem_reg[14][2]  ( .D(\u_a23_mem/n18258 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[114]) );
  DFF \u_a23_mem/out_mem_reg[14][3]  ( .D(\u_a23_mem/n18257 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[115]) );
  DFF \u_a23_mem/out_mem_reg[14][4]  ( .D(\u_a23_mem/n18256 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[116]) );
  DFF \u_a23_mem/out_mem_reg[14][5]  ( .D(\u_a23_mem/n18255 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[117]) );
  DFF \u_a23_mem/out_mem_reg[14][6]  ( .D(\u_a23_mem/n18254 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[118]) );
  DFF \u_a23_mem/out_mem_reg[14][7]  ( .D(\u_a23_mem/n18253 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[119]) );
  DFF \u_a23_mem/out_mem_reg[15][0]  ( .D(\u_a23_mem/n18252 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[120]) );
  DFF \u_a23_mem/out_mem_reg[15][1]  ( .D(\u_a23_mem/n18251 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[121]) );
  DFF \u_a23_mem/out_mem_reg[15][2]  ( .D(\u_a23_mem/n18250 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[122]) );
  DFF \u_a23_mem/out_mem_reg[15][3]  ( .D(\u_a23_mem/n18249 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[123]) );
  DFF \u_a23_mem/out_mem_reg[15][4]  ( .D(\u_a23_mem/n18248 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[124]) );
  DFF \u_a23_mem/out_mem_reg[15][5]  ( .D(\u_a23_mem/n18247 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[125]) );
  DFF \u_a23_mem/out_mem_reg[15][6]  ( .D(\u_a23_mem/n18246 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[126]) );
  DFF \u_a23_mem/out_mem_reg[15][7]  ( .D(\u_a23_mem/n18245 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[127]) );
  DFF \u_a23_mem/out_mem_reg[16][0]  ( .D(\u_a23_mem/n18244 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[128]) );
  DFF \u_a23_mem/out_mem_reg[16][1]  ( .D(\u_a23_mem/n18243 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[129]) );
  DFF \u_a23_mem/out_mem_reg[16][2]  ( .D(\u_a23_mem/n18242 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[130]) );
  DFF \u_a23_mem/out_mem_reg[16][3]  ( .D(\u_a23_mem/n18241 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[131]) );
  DFF \u_a23_mem/out_mem_reg[16][4]  ( .D(\u_a23_mem/n18240 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[132]) );
  DFF \u_a23_mem/out_mem_reg[16][5]  ( .D(\u_a23_mem/n18239 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[133]) );
  DFF \u_a23_mem/out_mem_reg[16][6]  ( .D(\u_a23_mem/n18238 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[134]) );
  DFF \u_a23_mem/out_mem_reg[16][7]  ( .D(\u_a23_mem/n18237 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[135]) );
  DFF \u_a23_mem/out_mem_reg[17][0]  ( .D(\u_a23_mem/n18236 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[136]) );
  DFF \u_a23_mem/out_mem_reg[17][1]  ( .D(\u_a23_mem/n18235 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[137]) );
  DFF \u_a23_mem/out_mem_reg[17][2]  ( .D(\u_a23_mem/n18234 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[138]) );
  DFF \u_a23_mem/out_mem_reg[17][3]  ( .D(\u_a23_mem/n18233 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[139]) );
  DFF \u_a23_mem/out_mem_reg[17][4]  ( .D(\u_a23_mem/n18232 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[140]) );
  DFF \u_a23_mem/out_mem_reg[17][5]  ( .D(\u_a23_mem/n18231 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[141]) );
  DFF \u_a23_mem/out_mem_reg[17][6]  ( .D(\u_a23_mem/n18230 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[142]) );
  DFF \u_a23_mem/out_mem_reg[17][7]  ( .D(\u_a23_mem/n18229 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[143]) );
  DFF \u_a23_mem/out_mem_reg[18][0]  ( .D(\u_a23_mem/n18228 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[144]) );
  DFF \u_a23_mem/out_mem_reg[18][1]  ( .D(\u_a23_mem/n18227 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[145]) );
  DFF \u_a23_mem/out_mem_reg[18][2]  ( .D(\u_a23_mem/n18226 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[146]) );
  DFF \u_a23_mem/out_mem_reg[18][3]  ( .D(\u_a23_mem/n18225 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[147]) );
  DFF \u_a23_mem/out_mem_reg[18][4]  ( .D(\u_a23_mem/n18224 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[148]) );
  DFF \u_a23_mem/out_mem_reg[18][5]  ( .D(\u_a23_mem/n18223 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[149]) );
  DFF \u_a23_mem/out_mem_reg[18][6]  ( .D(\u_a23_mem/n18222 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[150]) );
  DFF \u_a23_mem/out_mem_reg[18][7]  ( .D(\u_a23_mem/n18221 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[151]) );
  DFF \u_a23_mem/out_mem_reg[19][0]  ( .D(\u_a23_mem/n18220 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[152]) );
  DFF \u_a23_mem/out_mem_reg[19][1]  ( .D(\u_a23_mem/n18219 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[153]) );
  DFF \u_a23_mem/out_mem_reg[19][2]  ( .D(\u_a23_mem/n18218 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[154]) );
  DFF \u_a23_mem/out_mem_reg[19][3]  ( .D(\u_a23_mem/n18217 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[155]) );
  DFF \u_a23_mem/out_mem_reg[19][4]  ( .D(\u_a23_mem/n18216 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[156]) );
  DFF \u_a23_mem/out_mem_reg[19][5]  ( .D(\u_a23_mem/n18215 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[157]) );
  DFF \u_a23_mem/out_mem_reg[19][6]  ( .D(\u_a23_mem/n18214 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[158]) );
  DFF \u_a23_mem/out_mem_reg[19][7]  ( .D(\u_a23_mem/n18213 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[159]) );
  DFF \u_a23_mem/out_mem_reg[20][0]  ( .D(\u_a23_mem/n18212 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[160]) );
  DFF \u_a23_mem/out_mem_reg[20][1]  ( .D(\u_a23_mem/n18211 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[161]) );
  DFF \u_a23_mem/out_mem_reg[20][2]  ( .D(\u_a23_mem/n18210 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[162]) );
  DFF \u_a23_mem/out_mem_reg[20][3]  ( .D(\u_a23_mem/n18209 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[163]) );
  DFF \u_a23_mem/out_mem_reg[20][4]  ( .D(\u_a23_mem/n18208 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[164]) );
  DFF \u_a23_mem/out_mem_reg[20][5]  ( .D(\u_a23_mem/n18207 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[165]) );
  DFF \u_a23_mem/out_mem_reg[20][6]  ( .D(\u_a23_mem/n18206 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[166]) );
  DFF \u_a23_mem/out_mem_reg[20][7]  ( .D(\u_a23_mem/n18205 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[167]) );
  DFF \u_a23_mem/out_mem_reg[21][0]  ( .D(\u_a23_mem/n18204 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[168]) );
  DFF \u_a23_mem/out_mem_reg[21][1]  ( .D(\u_a23_mem/n18203 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[169]) );
  DFF \u_a23_mem/out_mem_reg[21][2]  ( .D(\u_a23_mem/n18202 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[170]) );
  DFF \u_a23_mem/out_mem_reg[21][3]  ( .D(\u_a23_mem/n18201 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[171]) );
  DFF \u_a23_mem/out_mem_reg[21][4]  ( .D(\u_a23_mem/n18200 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[172]) );
  DFF \u_a23_mem/out_mem_reg[21][5]  ( .D(\u_a23_mem/n18199 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[173]) );
  DFF \u_a23_mem/out_mem_reg[21][6]  ( .D(\u_a23_mem/n18198 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[174]) );
  DFF \u_a23_mem/out_mem_reg[21][7]  ( .D(\u_a23_mem/n18197 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[175]) );
  DFF \u_a23_mem/out_mem_reg[22][0]  ( .D(\u_a23_mem/n18196 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[176]) );
  DFF \u_a23_mem/out_mem_reg[22][1]  ( .D(\u_a23_mem/n18195 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[177]) );
  DFF \u_a23_mem/out_mem_reg[22][2]  ( .D(\u_a23_mem/n18194 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[178]) );
  DFF \u_a23_mem/out_mem_reg[22][3]  ( .D(\u_a23_mem/n18193 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[179]) );
  DFF \u_a23_mem/out_mem_reg[22][4]  ( .D(\u_a23_mem/n18192 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[180]) );
  DFF \u_a23_mem/out_mem_reg[22][5]  ( .D(\u_a23_mem/n18191 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[181]) );
  DFF \u_a23_mem/out_mem_reg[22][6]  ( .D(\u_a23_mem/n18190 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[182]) );
  DFF \u_a23_mem/out_mem_reg[22][7]  ( .D(\u_a23_mem/n18189 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[183]) );
  DFF \u_a23_mem/out_mem_reg[23][0]  ( .D(\u_a23_mem/n18188 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[184]) );
  DFF \u_a23_mem/out_mem_reg[23][1]  ( .D(\u_a23_mem/n18187 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[185]) );
  DFF \u_a23_mem/out_mem_reg[23][2]  ( .D(\u_a23_mem/n18186 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[186]) );
  DFF \u_a23_mem/out_mem_reg[23][3]  ( .D(\u_a23_mem/n18185 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[187]) );
  DFF \u_a23_mem/out_mem_reg[23][4]  ( .D(\u_a23_mem/n18184 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[188]) );
  DFF \u_a23_mem/out_mem_reg[23][5]  ( .D(\u_a23_mem/n18183 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[189]) );
  DFF \u_a23_mem/out_mem_reg[23][6]  ( .D(\u_a23_mem/n18182 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[190]) );
  DFF \u_a23_mem/out_mem_reg[23][7]  ( .D(\u_a23_mem/n18181 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[191]) );
  DFF \u_a23_mem/out_mem_reg[24][0]  ( .D(\u_a23_mem/n18180 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[192]) );
  DFF \u_a23_mem/out_mem_reg[24][1]  ( .D(\u_a23_mem/n18179 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[193]) );
  DFF \u_a23_mem/out_mem_reg[24][2]  ( .D(\u_a23_mem/n18178 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[194]) );
  DFF \u_a23_mem/out_mem_reg[24][3]  ( .D(\u_a23_mem/n18177 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[195]) );
  DFF \u_a23_mem/out_mem_reg[24][4]  ( .D(\u_a23_mem/n18176 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[196]) );
  DFF \u_a23_mem/out_mem_reg[24][5]  ( .D(\u_a23_mem/n18175 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[197]) );
  DFF \u_a23_mem/out_mem_reg[24][6]  ( .D(\u_a23_mem/n18174 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[198]) );
  DFF \u_a23_mem/out_mem_reg[24][7]  ( .D(\u_a23_mem/n18173 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[199]) );
  DFF \u_a23_mem/out_mem_reg[25][0]  ( .D(\u_a23_mem/n18172 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[200]) );
  DFF \u_a23_mem/out_mem_reg[25][1]  ( .D(\u_a23_mem/n18171 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[201]) );
  DFF \u_a23_mem/out_mem_reg[25][2]  ( .D(\u_a23_mem/n18170 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[202]) );
  DFF \u_a23_mem/out_mem_reg[25][3]  ( .D(\u_a23_mem/n18169 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[203]) );
  DFF \u_a23_mem/out_mem_reg[25][4]  ( .D(\u_a23_mem/n18168 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[204]) );
  DFF \u_a23_mem/out_mem_reg[25][5]  ( .D(\u_a23_mem/n18167 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[205]) );
  DFF \u_a23_mem/out_mem_reg[25][6]  ( .D(\u_a23_mem/n18166 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[206]) );
  DFF \u_a23_mem/out_mem_reg[25][7]  ( .D(\u_a23_mem/n18165 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[207]) );
  DFF \u_a23_mem/out_mem_reg[26][0]  ( .D(\u_a23_mem/n18164 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[208]) );
  DFF \u_a23_mem/out_mem_reg[26][1]  ( .D(\u_a23_mem/n18163 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[209]) );
  DFF \u_a23_mem/out_mem_reg[26][2]  ( .D(\u_a23_mem/n18162 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[210]) );
  DFF \u_a23_mem/out_mem_reg[26][3]  ( .D(\u_a23_mem/n18161 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[211]) );
  DFF \u_a23_mem/out_mem_reg[26][4]  ( .D(\u_a23_mem/n18160 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[212]) );
  DFF \u_a23_mem/out_mem_reg[26][5]  ( .D(\u_a23_mem/n18159 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[213]) );
  DFF \u_a23_mem/out_mem_reg[26][6]  ( .D(\u_a23_mem/n18158 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[214]) );
  DFF \u_a23_mem/out_mem_reg[26][7]  ( .D(\u_a23_mem/n18157 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[215]) );
  DFF \u_a23_mem/out_mem_reg[27][0]  ( .D(\u_a23_mem/n18156 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[216]) );
  DFF \u_a23_mem/out_mem_reg[27][1]  ( .D(\u_a23_mem/n18155 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[217]) );
  DFF \u_a23_mem/out_mem_reg[27][2]  ( .D(\u_a23_mem/n18154 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[218]) );
  DFF \u_a23_mem/out_mem_reg[27][3]  ( .D(\u_a23_mem/n18153 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[219]) );
  DFF \u_a23_mem/out_mem_reg[27][4]  ( .D(\u_a23_mem/n18152 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[220]) );
  DFF \u_a23_mem/out_mem_reg[27][5]  ( .D(\u_a23_mem/n18151 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[221]) );
  DFF \u_a23_mem/out_mem_reg[27][6]  ( .D(\u_a23_mem/n18150 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[222]) );
  DFF \u_a23_mem/out_mem_reg[27][7]  ( .D(\u_a23_mem/n18149 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[223]) );
  DFF \u_a23_mem/out_mem_reg[28][0]  ( .D(\u_a23_mem/n18148 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[224]) );
  DFF \u_a23_mem/out_mem_reg[28][1]  ( .D(\u_a23_mem/n18147 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[225]) );
  DFF \u_a23_mem/out_mem_reg[28][2]  ( .D(\u_a23_mem/n18146 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[226]) );
  DFF \u_a23_mem/out_mem_reg[28][3]  ( .D(\u_a23_mem/n18145 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[227]) );
  DFF \u_a23_mem/out_mem_reg[28][4]  ( .D(\u_a23_mem/n18144 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[228]) );
  DFF \u_a23_mem/out_mem_reg[28][5]  ( .D(\u_a23_mem/n18143 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[229]) );
  DFF \u_a23_mem/out_mem_reg[28][6]  ( .D(\u_a23_mem/n18142 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[230]) );
  DFF \u_a23_mem/out_mem_reg[28][7]  ( .D(\u_a23_mem/n18141 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[231]) );
  DFF \u_a23_mem/out_mem_reg[29][0]  ( .D(\u_a23_mem/n18140 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[232]) );
  DFF \u_a23_mem/out_mem_reg[29][1]  ( .D(\u_a23_mem/n18139 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[233]) );
  DFF \u_a23_mem/out_mem_reg[29][2]  ( .D(\u_a23_mem/n18138 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[234]) );
  DFF \u_a23_mem/out_mem_reg[29][3]  ( .D(\u_a23_mem/n18137 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[235]) );
  DFF \u_a23_mem/out_mem_reg[29][4]  ( .D(\u_a23_mem/n18136 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[236]) );
  DFF \u_a23_mem/out_mem_reg[29][5]  ( .D(\u_a23_mem/n18135 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[237]) );
  DFF \u_a23_mem/out_mem_reg[29][6]  ( .D(\u_a23_mem/n18134 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[238]) );
  DFF \u_a23_mem/out_mem_reg[29][7]  ( .D(\u_a23_mem/n18133 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[239]) );
  DFF \u_a23_mem/out_mem_reg[30][0]  ( .D(\u_a23_mem/n18132 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[240]) );
  DFF \u_a23_mem/out_mem_reg[30][1]  ( .D(\u_a23_mem/n18131 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[241]) );
  DFF \u_a23_mem/out_mem_reg[30][2]  ( .D(\u_a23_mem/n18130 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[242]) );
  DFF \u_a23_mem/out_mem_reg[30][3]  ( .D(\u_a23_mem/n18129 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[243]) );
  DFF \u_a23_mem/out_mem_reg[30][4]  ( .D(\u_a23_mem/n18128 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[244]) );
  DFF \u_a23_mem/out_mem_reg[30][5]  ( .D(\u_a23_mem/n18127 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[245]) );
  DFF \u_a23_mem/out_mem_reg[30][6]  ( .D(\u_a23_mem/n18126 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[246]) );
  DFF \u_a23_mem/out_mem_reg[30][7]  ( .D(\u_a23_mem/n18125 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[247]) );
  DFF \u_a23_mem/out_mem_reg[31][0]  ( .D(\u_a23_mem/n18124 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[248]) );
  DFF \u_a23_mem/out_mem_reg[31][1]  ( .D(\u_a23_mem/n18123 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[249]) );
  DFF \u_a23_mem/out_mem_reg[31][2]  ( .D(\u_a23_mem/n18122 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[250]) );
  DFF \u_a23_mem/out_mem_reg[31][3]  ( .D(\u_a23_mem/n18121 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[251]) );
  DFF \u_a23_mem/out_mem_reg[31][4]  ( .D(\u_a23_mem/n18120 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[252]) );
  DFF \u_a23_mem/out_mem_reg[31][5]  ( .D(\u_a23_mem/n18119 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[253]) );
  DFF \u_a23_mem/out_mem_reg[31][6]  ( .D(\u_a23_mem/n18118 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[254]) );
  DFF \u_a23_mem/out_mem_reg[31][7]  ( .D(\u_a23_mem/n18117 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(o[255]) );
  DFF \u_a23_mem/g_mem_reg[0][0]  ( .D(\u_a23_mem/g_mem[0][0] ), .CLK(clk), 
        .RST(rst), .I(g_init[0]), .Q(\u_a23_mem/g_mem[0][0] ) );
  DFF \u_a23_mem/g_mem_reg[0][1]  ( .D(\u_a23_mem/g_mem[0][1] ), .CLK(clk), 
        .RST(rst), .I(g_init[1]), .Q(\u_a23_mem/g_mem[0][1] ) );
  DFF \u_a23_mem/g_mem_reg[0][2]  ( .D(\u_a23_mem/g_mem[0][2] ), .CLK(clk), 
        .RST(rst), .I(g_init[2]), .Q(\u_a23_mem/g_mem[0][2] ) );
  DFF \u_a23_mem/g_mem_reg[0][3]  ( .D(\u_a23_mem/g_mem[0][3] ), .CLK(clk), 
        .RST(rst), .I(g_init[3]), .Q(\u_a23_mem/g_mem[0][3] ) );
  DFF \u_a23_mem/g_mem_reg[0][4]  ( .D(\u_a23_mem/g_mem[0][4] ), .CLK(clk), 
        .RST(rst), .I(g_init[4]), .Q(\u_a23_mem/g_mem[0][4] ) );
  DFF \u_a23_mem/g_mem_reg[0][5]  ( .D(\u_a23_mem/g_mem[0][5] ), .CLK(clk), 
        .RST(rst), .I(g_init[5]), .Q(\u_a23_mem/g_mem[0][5] ) );
  DFF \u_a23_mem/g_mem_reg[0][6]  ( .D(\u_a23_mem/g_mem[0][6] ), .CLK(clk), 
        .RST(rst), .I(g_init[6]), .Q(\u_a23_mem/g_mem[0][6] ) );
  DFF \u_a23_mem/g_mem_reg[0][7]  ( .D(\u_a23_mem/g_mem[0][7] ), .CLK(clk), 
        .RST(rst), .I(g_init[7]), .Q(\u_a23_mem/g_mem[0][7] ) );
  DFF \u_a23_mem/g_mem_reg[1][0]  ( .D(\u_a23_mem/g_mem[1][0] ), .CLK(clk), 
        .RST(rst), .I(g_init[8]), .Q(\u_a23_mem/g_mem[1][0] ) );
  DFF \u_a23_mem/g_mem_reg[1][1]  ( .D(\u_a23_mem/g_mem[1][1] ), .CLK(clk), 
        .RST(rst), .I(g_init[9]), .Q(\u_a23_mem/g_mem[1][1] ) );
  DFF \u_a23_mem/g_mem_reg[1][2]  ( .D(\u_a23_mem/g_mem[1][2] ), .CLK(clk), 
        .RST(rst), .I(g_init[10]), .Q(\u_a23_mem/g_mem[1][2] ) );
  DFF \u_a23_mem/g_mem_reg[1][3]  ( .D(\u_a23_mem/g_mem[1][3] ), .CLK(clk), 
        .RST(rst), .I(g_init[11]), .Q(\u_a23_mem/g_mem[1][3] ) );
  DFF \u_a23_mem/g_mem_reg[1][4]  ( .D(\u_a23_mem/g_mem[1][4] ), .CLK(clk), 
        .RST(rst), .I(g_init[12]), .Q(\u_a23_mem/g_mem[1][4] ) );
  DFF \u_a23_mem/g_mem_reg[1][5]  ( .D(\u_a23_mem/g_mem[1][5] ), .CLK(clk), 
        .RST(rst), .I(g_init[13]), .Q(\u_a23_mem/g_mem[1][5] ) );
  DFF \u_a23_mem/g_mem_reg[1][6]  ( .D(\u_a23_mem/g_mem[1][6] ), .CLK(clk), 
        .RST(rst), .I(g_init[14]), .Q(\u_a23_mem/g_mem[1][6] ) );
  DFF \u_a23_mem/g_mem_reg[1][7]  ( .D(\u_a23_mem/g_mem[1][7] ), .CLK(clk), 
        .RST(rst), .I(g_init[15]), .Q(\u_a23_mem/g_mem[1][7] ) );
  DFF \u_a23_mem/g_mem_reg[2][0]  ( .D(\u_a23_mem/g_mem[2][0] ), .CLK(clk), 
        .RST(rst), .I(g_init[16]), .Q(\u_a23_mem/g_mem[2][0] ) );
  DFF \u_a23_mem/g_mem_reg[2][1]  ( .D(\u_a23_mem/g_mem[2][1] ), .CLK(clk), 
        .RST(rst), .I(g_init[17]), .Q(\u_a23_mem/g_mem[2][1] ) );
  DFF \u_a23_mem/g_mem_reg[2][2]  ( .D(\u_a23_mem/g_mem[2][2] ), .CLK(clk), 
        .RST(rst), .I(g_init[18]), .Q(\u_a23_mem/g_mem[2][2] ) );
  DFF \u_a23_mem/g_mem_reg[2][3]  ( .D(\u_a23_mem/g_mem[2][3] ), .CLK(clk), 
        .RST(rst), .I(g_init[19]), .Q(\u_a23_mem/g_mem[2][3] ) );
  DFF \u_a23_mem/g_mem_reg[2][4]  ( .D(\u_a23_mem/g_mem[2][4] ), .CLK(clk), 
        .RST(rst), .I(g_init[20]), .Q(\u_a23_mem/g_mem[2][4] ) );
  DFF \u_a23_mem/g_mem_reg[2][5]  ( .D(\u_a23_mem/g_mem[2][5] ), .CLK(clk), 
        .RST(rst), .I(g_init[21]), .Q(\u_a23_mem/g_mem[2][5] ) );
  DFF \u_a23_mem/g_mem_reg[2][6]  ( .D(\u_a23_mem/g_mem[2][6] ), .CLK(clk), 
        .RST(rst), .I(g_init[22]), .Q(\u_a23_mem/g_mem[2][6] ) );
  DFF \u_a23_mem/g_mem_reg[2][7]  ( .D(\u_a23_mem/g_mem[2][7] ), .CLK(clk), 
        .RST(rst), .I(g_init[23]), .Q(\u_a23_mem/g_mem[2][7] ) );
  DFF \u_a23_mem/g_mem_reg[3][0]  ( .D(\u_a23_mem/g_mem[3][0] ), .CLK(clk), 
        .RST(rst), .I(g_init[24]), .Q(\u_a23_mem/g_mem[3][0] ) );
  DFF \u_a23_mem/g_mem_reg[3][1]  ( .D(\u_a23_mem/g_mem[3][1] ), .CLK(clk), 
        .RST(rst), .I(g_init[25]), .Q(\u_a23_mem/g_mem[3][1] ) );
  DFF \u_a23_mem/g_mem_reg[3][2]  ( .D(\u_a23_mem/g_mem[3][2] ), .CLK(clk), 
        .RST(rst), .I(g_init[26]), .Q(\u_a23_mem/g_mem[3][2] ) );
  DFF \u_a23_mem/g_mem_reg[3][3]  ( .D(\u_a23_mem/g_mem[3][3] ), .CLK(clk), 
        .RST(rst), .I(g_init[27]), .Q(\u_a23_mem/g_mem[3][3] ) );
  DFF \u_a23_mem/g_mem_reg[3][4]  ( .D(\u_a23_mem/g_mem[3][4] ), .CLK(clk), 
        .RST(rst), .I(g_init[28]), .Q(\u_a23_mem/g_mem[3][4] ) );
  DFF \u_a23_mem/g_mem_reg[3][5]  ( .D(\u_a23_mem/g_mem[3][5] ), .CLK(clk), 
        .RST(rst), .I(g_init[29]), .Q(\u_a23_mem/g_mem[3][5] ) );
  DFF \u_a23_mem/g_mem_reg[3][6]  ( .D(\u_a23_mem/g_mem[3][6] ), .CLK(clk), 
        .RST(rst), .I(g_init[30]), .Q(\u_a23_mem/g_mem[3][6] ) );
  DFF \u_a23_mem/g_mem_reg[3][7]  ( .D(\u_a23_mem/g_mem[3][7] ), .CLK(clk), 
        .RST(rst), .I(g_init[31]), .Q(\u_a23_mem/g_mem[3][7] ) );
  DFF \u_a23_mem/g_mem_reg[4][0]  ( .D(\u_a23_mem/g_mem[4][0] ), .CLK(clk), 
        .RST(rst), .I(g_init[32]), .Q(\u_a23_mem/g_mem[4][0] ) );
  DFF \u_a23_mem/g_mem_reg[4][1]  ( .D(\u_a23_mem/g_mem[4][1] ), .CLK(clk), 
        .RST(rst), .I(g_init[33]), .Q(\u_a23_mem/g_mem[4][1] ) );
  DFF \u_a23_mem/g_mem_reg[4][2]  ( .D(\u_a23_mem/g_mem[4][2] ), .CLK(clk), 
        .RST(rst), .I(g_init[34]), .Q(\u_a23_mem/g_mem[4][2] ) );
  DFF \u_a23_mem/g_mem_reg[4][3]  ( .D(\u_a23_mem/g_mem[4][3] ), .CLK(clk), 
        .RST(rst), .I(g_init[35]), .Q(\u_a23_mem/g_mem[4][3] ) );
  DFF \u_a23_mem/g_mem_reg[4][4]  ( .D(\u_a23_mem/g_mem[4][4] ), .CLK(clk), 
        .RST(rst), .I(g_init[36]), .Q(\u_a23_mem/g_mem[4][4] ) );
  DFF \u_a23_mem/g_mem_reg[4][5]  ( .D(\u_a23_mem/g_mem[4][5] ), .CLK(clk), 
        .RST(rst), .I(g_init[37]), .Q(\u_a23_mem/g_mem[4][5] ) );
  DFF \u_a23_mem/g_mem_reg[4][6]  ( .D(\u_a23_mem/g_mem[4][6] ), .CLK(clk), 
        .RST(rst), .I(g_init[38]), .Q(\u_a23_mem/g_mem[4][6] ) );
  DFF \u_a23_mem/g_mem_reg[4][7]  ( .D(\u_a23_mem/g_mem[4][7] ), .CLK(clk), 
        .RST(rst), .I(g_init[39]), .Q(\u_a23_mem/g_mem[4][7] ) );
  DFF \u_a23_mem/g_mem_reg[5][0]  ( .D(\u_a23_mem/g_mem[5][0] ), .CLK(clk), 
        .RST(rst), .I(g_init[40]), .Q(\u_a23_mem/g_mem[5][0] ) );
  DFF \u_a23_mem/g_mem_reg[5][1]  ( .D(\u_a23_mem/g_mem[5][1] ), .CLK(clk), 
        .RST(rst), .I(g_init[41]), .Q(\u_a23_mem/g_mem[5][1] ) );
  DFF \u_a23_mem/g_mem_reg[5][2]  ( .D(\u_a23_mem/g_mem[5][2] ), .CLK(clk), 
        .RST(rst), .I(g_init[42]), .Q(\u_a23_mem/g_mem[5][2] ) );
  DFF \u_a23_mem/g_mem_reg[5][3]  ( .D(\u_a23_mem/g_mem[5][3] ), .CLK(clk), 
        .RST(rst), .I(g_init[43]), .Q(\u_a23_mem/g_mem[5][3] ) );
  DFF \u_a23_mem/g_mem_reg[5][4]  ( .D(\u_a23_mem/g_mem[5][4] ), .CLK(clk), 
        .RST(rst), .I(g_init[44]), .Q(\u_a23_mem/g_mem[5][4] ) );
  DFF \u_a23_mem/g_mem_reg[5][5]  ( .D(\u_a23_mem/g_mem[5][5] ), .CLK(clk), 
        .RST(rst), .I(g_init[45]), .Q(\u_a23_mem/g_mem[5][5] ) );
  DFF \u_a23_mem/g_mem_reg[5][6]  ( .D(\u_a23_mem/g_mem[5][6] ), .CLK(clk), 
        .RST(rst), .I(g_init[46]), .Q(\u_a23_mem/g_mem[5][6] ) );
  DFF \u_a23_mem/g_mem_reg[5][7]  ( .D(\u_a23_mem/g_mem[5][7] ), .CLK(clk), 
        .RST(rst), .I(g_init[47]), .Q(\u_a23_mem/g_mem[5][7] ) );
  DFF \u_a23_mem/g_mem_reg[6][0]  ( .D(\u_a23_mem/g_mem[6][0] ), .CLK(clk), 
        .RST(rst), .I(g_init[48]), .Q(\u_a23_mem/g_mem[6][0] ) );
  DFF \u_a23_mem/g_mem_reg[6][1]  ( .D(\u_a23_mem/g_mem[6][1] ), .CLK(clk), 
        .RST(rst), .I(g_init[49]), .Q(\u_a23_mem/g_mem[6][1] ) );
  DFF \u_a23_mem/g_mem_reg[6][2]  ( .D(\u_a23_mem/g_mem[6][2] ), .CLK(clk), 
        .RST(rst), .I(g_init[50]), .Q(\u_a23_mem/g_mem[6][2] ) );
  DFF \u_a23_mem/g_mem_reg[6][3]  ( .D(\u_a23_mem/g_mem[6][3] ), .CLK(clk), 
        .RST(rst), .I(g_init[51]), .Q(\u_a23_mem/g_mem[6][3] ) );
  DFF \u_a23_mem/g_mem_reg[6][4]  ( .D(\u_a23_mem/g_mem[6][4] ), .CLK(clk), 
        .RST(rst), .I(g_init[52]), .Q(\u_a23_mem/g_mem[6][4] ) );
  DFF \u_a23_mem/g_mem_reg[6][5]  ( .D(\u_a23_mem/g_mem[6][5] ), .CLK(clk), 
        .RST(rst), .I(g_init[53]), .Q(\u_a23_mem/g_mem[6][5] ) );
  DFF \u_a23_mem/g_mem_reg[6][6]  ( .D(\u_a23_mem/g_mem[6][6] ), .CLK(clk), 
        .RST(rst), .I(g_init[54]), .Q(\u_a23_mem/g_mem[6][6] ) );
  DFF \u_a23_mem/g_mem_reg[6][7]  ( .D(\u_a23_mem/g_mem[6][7] ), .CLK(clk), 
        .RST(rst), .I(g_init[55]), .Q(\u_a23_mem/g_mem[6][7] ) );
  DFF \u_a23_mem/g_mem_reg[7][0]  ( .D(\u_a23_mem/g_mem[7][0] ), .CLK(clk), 
        .RST(rst), .I(g_init[56]), .Q(\u_a23_mem/g_mem[7][0] ) );
  DFF \u_a23_mem/g_mem_reg[7][1]  ( .D(\u_a23_mem/g_mem[7][1] ), .CLK(clk), 
        .RST(rst), .I(g_init[57]), .Q(\u_a23_mem/g_mem[7][1] ) );
  DFF \u_a23_mem/g_mem_reg[7][2]  ( .D(\u_a23_mem/g_mem[7][2] ), .CLK(clk), 
        .RST(rst), .I(g_init[58]), .Q(\u_a23_mem/g_mem[7][2] ) );
  DFF \u_a23_mem/g_mem_reg[7][3]  ( .D(\u_a23_mem/g_mem[7][3] ), .CLK(clk), 
        .RST(rst), .I(g_init[59]), .Q(\u_a23_mem/g_mem[7][3] ) );
  DFF \u_a23_mem/g_mem_reg[7][4]  ( .D(\u_a23_mem/g_mem[7][4] ), .CLK(clk), 
        .RST(rst), .I(g_init[60]), .Q(\u_a23_mem/g_mem[7][4] ) );
  DFF \u_a23_mem/g_mem_reg[7][5]  ( .D(\u_a23_mem/g_mem[7][5] ), .CLK(clk), 
        .RST(rst), .I(g_init[61]), .Q(\u_a23_mem/g_mem[7][5] ) );
  DFF \u_a23_mem/g_mem_reg[7][6]  ( .D(\u_a23_mem/g_mem[7][6] ), .CLK(clk), 
        .RST(rst), .I(g_init[62]), .Q(\u_a23_mem/g_mem[7][6] ) );
  DFF \u_a23_mem/g_mem_reg[7][7]  ( .D(\u_a23_mem/g_mem[7][7] ), .CLK(clk), 
        .RST(rst), .I(g_init[63]), .Q(\u_a23_mem/g_mem[7][7] ) );
  DFF \u_a23_mem/g_mem_reg[8][0]  ( .D(\u_a23_mem/g_mem[8][0] ), .CLK(clk), 
        .RST(rst), .I(g_init[64]), .Q(\u_a23_mem/g_mem[8][0] ) );
  DFF \u_a23_mem/g_mem_reg[8][1]  ( .D(\u_a23_mem/g_mem[8][1] ), .CLK(clk), 
        .RST(rst), .I(g_init[65]), .Q(\u_a23_mem/g_mem[8][1] ) );
  DFF \u_a23_mem/g_mem_reg[8][2]  ( .D(\u_a23_mem/g_mem[8][2] ), .CLK(clk), 
        .RST(rst), .I(g_init[66]), .Q(\u_a23_mem/g_mem[8][2] ) );
  DFF \u_a23_mem/g_mem_reg[8][3]  ( .D(\u_a23_mem/g_mem[8][3] ), .CLK(clk), 
        .RST(rst), .I(g_init[67]), .Q(\u_a23_mem/g_mem[8][3] ) );
  DFF \u_a23_mem/g_mem_reg[8][4]  ( .D(\u_a23_mem/g_mem[8][4] ), .CLK(clk), 
        .RST(rst), .I(g_init[68]), .Q(\u_a23_mem/g_mem[8][4] ) );
  DFF \u_a23_mem/g_mem_reg[8][5]  ( .D(\u_a23_mem/g_mem[8][5] ), .CLK(clk), 
        .RST(rst), .I(g_init[69]), .Q(\u_a23_mem/g_mem[8][5] ) );
  DFF \u_a23_mem/g_mem_reg[8][6]  ( .D(\u_a23_mem/g_mem[8][6] ), .CLK(clk), 
        .RST(rst), .I(g_init[70]), .Q(\u_a23_mem/g_mem[8][6] ) );
  DFF \u_a23_mem/g_mem_reg[8][7]  ( .D(\u_a23_mem/g_mem[8][7] ), .CLK(clk), 
        .RST(rst), .I(g_init[71]), .Q(\u_a23_mem/g_mem[8][7] ) );
  DFF \u_a23_mem/g_mem_reg[9][0]  ( .D(\u_a23_mem/g_mem[9][0] ), .CLK(clk), 
        .RST(rst), .I(g_init[72]), .Q(\u_a23_mem/g_mem[9][0] ) );
  DFF \u_a23_mem/g_mem_reg[9][1]  ( .D(\u_a23_mem/g_mem[9][1] ), .CLK(clk), 
        .RST(rst), .I(g_init[73]), .Q(\u_a23_mem/g_mem[9][1] ) );
  DFF \u_a23_mem/g_mem_reg[9][2]  ( .D(\u_a23_mem/g_mem[9][2] ), .CLK(clk), 
        .RST(rst), .I(g_init[74]), .Q(\u_a23_mem/g_mem[9][2] ) );
  DFF \u_a23_mem/g_mem_reg[9][3]  ( .D(\u_a23_mem/g_mem[9][3] ), .CLK(clk), 
        .RST(rst), .I(g_init[75]), .Q(\u_a23_mem/g_mem[9][3] ) );
  DFF \u_a23_mem/g_mem_reg[9][4]  ( .D(\u_a23_mem/g_mem[9][4] ), .CLK(clk), 
        .RST(rst), .I(g_init[76]), .Q(\u_a23_mem/g_mem[9][4] ) );
  DFF \u_a23_mem/g_mem_reg[9][5]  ( .D(\u_a23_mem/g_mem[9][5] ), .CLK(clk), 
        .RST(rst), .I(g_init[77]), .Q(\u_a23_mem/g_mem[9][5] ) );
  DFF \u_a23_mem/g_mem_reg[9][6]  ( .D(\u_a23_mem/g_mem[9][6] ), .CLK(clk), 
        .RST(rst), .I(g_init[78]), .Q(\u_a23_mem/g_mem[9][6] ) );
  DFF \u_a23_mem/g_mem_reg[9][7]  ( .D(\u_a23_mem/g_mem[9][7] ), .CLK(clk), 
        .RST(rst), .I(g_init[79]), .Q(\u_a23_mem/g_mem[9][7] ) );
  DFF \u_a23_mem/g_mem_reg[10][0]  ( .D(\u_a23_mem/g_mem[10][0] ), .CLK(clk), 
        .RST(rst), .I(g_init[80]), .Q(\u_a23_mem/g_mem[10][0] ) );
  DFF \u_a23_mem/g_mem_reg[10][1]  ( .D(\u_a23_mem/g_mem[10][1] ), .CLK(clk), 
        .RST(rst), .I(g_init[81]), .Q(\u_a23_mem/g_mem[10][1] ) );
  DFF \u_a23_mem/g_mem_reg[10][2]  ( .D(\u_a23_mem/g_mem[10][2] ), .CLK(clk), 
        .RST(rst), .I(g_init[82]), .Q(\u_a23_mem/g_mem[10][2] ) );
  DFF \u_a23_mem/g_mem_reg[10][3]  ( .D(\u_a23_mem/g_mem[10][3] ), .CLK(clk), 
        .RST(rst), .I(g_init[83]), .Q(\u_a23_mem/g_mem[10][3] ) );
  DFF \u_a23_mem/g_mem_reg[10][4]  ( .D(\u_a23_mem/g_mem[10][4] ), .CLK(clk), 
        .RST(rst), .I(g_init[84]), .Q(\u_a23_mem/g_mem[10][4] ) );
  DFF \u_a23_mem/g_mem_reg[10][5]  ( .D(\u_a23_mem/g_mem[10][5] ), .CLK(clk), 
        .RST(rst), .I(g_init[85]), .Q(\u_a23_mem/g_mem[10][5] ) );
  DFF \u_a23_mem/g_mem_reg[10][6]  ( .D(\u_a23_mem/g_mem[10][6] ), .CLK(clk), 
        .RST(rst), .I(g_init[86]), .Q(\u_a23_mem/g_mem[10][6] ) );
  DFF \u_a23_mem/g_mem_reg[10][7]  ( .D(\u_a23_mem/g_mem[10][7] ), .CLK(clk), 
        .RST(rst), .I(g_init[87]), .Q(\u_a23_mem/g_mem[10][7] ) );
  DFF \u_a23_mem/g_mem_reg[11][0]  ( .D(\u_a23_mem/g_mem[11][0] ), .CLK(clk), 
        .RST(rst), .I(g_init[88]), .Q(\u_a23_mem/g_mem[11][0] ) );
  DFF \u_a23_mem/g_mem_reg[11][1]  ( .D(\u_a23_mem/g_mem[11][1] ), .CLK(clk), 
        .RST(rst), .I(g_init[89]), .Q(\u_a23_mem/g_mem[11][1] ) );
  DFF \u_a23_mem/g_mem_reg[11][2]  ( .D(\u_a23_mem/g_mem[11][2] ), .CLK(clk), 
        .RST(rst), .I(g_init[90]), .Q(\u_a23_mem/g_mem[11][2] ) );
  DFF \u_a23_mem/g_mem_reg[11][3]  ( .D(\u_a23_mem/g_mem[11][3] ), .CLK(clk), 
        .RST(rst), .I(g_init[91]), .Q(\u_a23_mem/g_mem[11][3] ) );
  DFF \u_a23_mem/g_mem_reg[11][4]  ( .D(\u_a23_mem/g_mem[11][4] ), .CLK(clk), 
        .RST(rst), .I(g_init[92]), .Q(\u_a23_mem/g_mem[11][4] ) );
  DFF \u_a23_mem/g_mem_reg[11][5]  ( .D(\u_a23_mem/g_mem[11][5] ), .CLK(clk), 
        .RST(rst), .I(g_init[93]), .Q(\u_a23_mem/g_mem[11][5] ) );
  DFF \u_a23_mem/g_mem_reg[11][6]  ( .D(\u_a23_mem/g_mem[11][6] ), .CLK(clk), 
        .RST(rst), .I(g_init[94]), .Q(\u_a23_mem/g_mem[11][6] ) );
  DFF \u_a23_mem/g_mem_reg[11][7]  ( .D(\u_a23_mem/g_mem[11][7] ), .CLK(clk), 
        .RST(rst), .I(g_init[95]), .Q(\u_a23_mem/g_mem[11][7] ) );
  DFF \u_a23_mem/g_mem_reg[12][0]  ( .D(\u_a23_mem/g_mem[12][0] ), .CLK(clk), 
        .RST(rst), .I(g_init[96]), .Q(\u_a23_mem/g_mem[12][0] ) );
  DFF \u_a23_mem/g_mem_reg[12][1]  ( .D(\u_a23_mem/g_mem[12][1] ), .CLK(clk), 
        .RST(rst), .I(g_init[97]), .Q(\u_a23_mem/g_mem[12][1] ) );
  DFF \u_a23_mem/g_mem_reg[12][2]  ( .D(\u_a23_mem/g_mem[12][2] ), .CLK(clk), 
        .RST(rst), .I(g_init[98]), .Q(\u_a23_mem/g_mem[12][2] ) );
  DFF \u_a23_mem/g_mem_reg[12][3]  ( .D(\u_a23_mem/g_mem[12][3] ), .CLK(clk), 
        .RST(rst), .I(g_init[99]), .Q(\u_a23_mem/g_mem[12][3] ) );
  DFF \u_a23_mem/g_mem_reg[12][4]  ( .D(\u_a23_mem/g_mem[12][4] ), .CLK(clk), 
        .RST(rst), .I(g_init[100]), .Q(\u_a23_mem/g_mem[12][4] ) );
  DFF \u_a23_mem/g_mem_reg[12][5]  ( .D(\u_a23_mem/g_mem[12][5] ), .CLK(clk), 
        .RST(rst), .I(g_init[101]), .Q(\u_a23_mem/g_mem[12][5] ) );
  DFF \u_a23_mem/g_mem_reg[12][6]  ( .D(\u_a23_mem/g_mem[12][6] ), .CLK(clk), 
        .RST(rst), .I(g_init[102]), .Q(\u_a23_mem/g_mem[12][6] ) );
  DFF \u_a23_mem/g_mem_reg[12][7]  ( .D(\u_a23_mem/g_mem[12][7] ), .CLK(clk), 
        .RST(rst), .I(g_init[103]), .Q(\u_a23_mem/g_mem[12][7] ) );
  DFF \u_a23_mem/g_mem_reg[13][0]  ( .D(\u_a23_mem/g_mem[13][0] ), .CLK(clk), 
        .RST(rst), .I(g_init[104]), .Q(\u_a23_mem/g_mem[13][0] ) );
  DFF \u_a23_mem/g_mem_reg[13][1]  ( .D(\u_a23_mem/g_mem[13][1] ), .CLK(clk), 
        .RST(rst), .I(g_init[105]), .Q(\u_a23_mem/g_mem[13][1] ) );
  DFF \u_a23_mem/g_mem_reg[13][2]  ( .D(\u_a23_mem/g_mem[13][2] ), .CLK(clk), 
        .RST(rst), .I(g_init[106]), .Q(\u_a23_mem/g_mem[13][2] ) );
  DFF \u_a23_mem/g_mem_reg[13][3]  ( .D(\u_a23_mem/g_mem[13][3] ), .CLK(clk), 
        .RST(rst), .I(g_init[107]), .Q(\u_a23_mem/g_mem[13][3] ) );
  DFF \u_a23_mem/g_mem_reg[13][4]  ( .D(\u_a23_mem/g_mem[13][4] ), .CLK(clk), 
        .RST(rst), .I(g_init[108]), .Q(\u_a23_mem/g_mem[13][4] ) );
  DFF \u_a23_mem/g_mem_reg[13][5]  ( .D(\u_a23_mem/g_mem[13][5] ), .CLK(clk), 
        .RST(rst), .I(g_init[109]), .Q(\u_a23_mem/g_mem[13][5] ) );
  DFF \u_a23_mem/g_mem_reg[13][6]  ( .D(\u_a23_mem/g_mem[13][6] ), .CLK(clk), 
        .RST(rst), .I(g_init[110]), .Q(\u_a23_mem/g_mem[13][6] ) );
  DFF \u_a23_mem/g_mem_reg[13][7]  ( .D(\u_a23_mem/g_mem[13][7] ), .CLK(clk), 
        .RST(rst), .I(g_init[111]), .Q(\u_a23_mem/g_mem[13][7] ) );
  DFF \u_a23_mem/g_mem_reg[14][0]  ( .D(\u_a23_mem/g_mem[14][0] ), .CLK(clk), 
        .RST(rst), .I(g_init[112]), .Q(\u_a23_mem/g_mem[14][0] ) );
  DFF \u_a23_mem/g_mem_reg[14][1]  ( .D(\u_a23_mem/g_mem[14][1] ), .CLK(clk), 
        .RST(rst), .I(g_init[113]), .Q(\u_a23_mem/g_mem[14][1] ) );
  DFF \u_a23_mem/g_mem_reg[14][2]  ( .D(\u_a23_mem/g_mem[14][2] ), .CLK(clk), 
        .RST(rst), .I(g_init[114]), .Q(\u_a23_mem/g_mem[14][2] ) );
  DFF \u_a23_mem/g_mem_reg[14][3]  ( .D(\u_a23_mem/g_mem[14][3] ), .CLK(clk), 
        .RST(rst), .I(g_init[115]), .Q(\u_a23_mem/g_mem[14][3] ) );
  DFF \u_a23_mem/g_mem_reg[14][4]  ( .D(\u_a23_mem/g_mem[14][4] ), .CLK(clk), 
        .RST(rst), .I(g_init[116]), .Q(\u_a23_mem/g_mem[14][4] ) );
  DFF \u_a23_mem/g_mem_reg[14][5]  ( .D(\u_a23_mem/g_mem[14][5] ), .CLK(clk), 
        .RST(rst), .I(g_init[117]), .Q(\u_a23_mem/g_mem[14][5] ) );
  DFF \u_a23_mem/g_mem_reg[14][6]  ( .D(\u_a23_mem/g_mem[14][6] ), .CLK(clk), 
        .RST(rst), .I(g_init[118]), .Q(\u_a23_mem/g_mem[14][6] ) );
  DFF \u_a23_mem/g_mem_reg[14][7]  ( .D(\u_a23_mem/g_mem[14][7] ), .CLK(clk), 
        .RST(rst), .I(g_init[119]), .Q(\u_a23_mem/g_mem[14][7] ) );
  DFF \u_a23_mem/g_mem_reg[15][0]  ( .D(\u_a23_mem/g_mem[15][0] ), .CLK(clk), 
        .RST(rst), .I(g_init[120]), .Q(\u_a23_mem/g_mem[15][0] ) );
  DFF \u_a23_mem/g_mem_reg[15][1]  ( .D(\u_a23_mem/g_mem[15][1] ), .CLK(clk), 
        .RST(rst), .I(g_init[121]), .Q(\u_a23_mem/g_mem[15][1] ) );
  DFF \u_a23_mem/g_mem_reg[15][2]  ( .D(\u_a23_mem/g_mem[15][2] ), .CLK(clk), 
        .RST(rst), .I(g_init[122]), .Q(\u_a23_mem/g_mem[15][2] ) );
  DFF \u_a23_mem/g_mem_reg[15][3]  ( .D(\u_a23_mem/g_mem[15][3] ), .CLK(clk), 
        .RST(rst), .I(g_init[123]), .Q(\u_a23_mem/g_mem[15][3] ) );
  DFF \u_a23_mem/g_mem_reg[15][4]  ( .D(\u_a23_mem/g_mem[15][4] ), .CLK(clk), 
        .RST(rst), .I(g_init[124]), .Q(\u_a23_mem/g_mem[15][4] ) );
  DFF \u_a23_mem/g_mem_reg[15][5]  ( .D(\u_a23_mem/g_mem[15][5] ), .CLK(clk), 
        .RST(rst), .I(g_init[125]), .Q(\u_a23_mem/g_mem[15][5] ) );
  DFF \u_a23_mem/g_mem_reg[15][6]  ( .D(\u_a23_mem/g_mem[15][6] ), .CLK(clk), 
        .RST(rst), .I(g_init[126]), .Q(\u_a23_mem/g_mem[15][6] ) );
  DFF \u_a23_mem/g_mem_reg[15][7]  ( .D(\u_a23_mem/g_mem[15][7] ), .CLK(clk), 
        .RST(rst), .I(g_init[127]), .Q(\u_a23_mem/g_mem[15][7] ) );
  DFF \u_a23_mem/g_mem_reg[16][0]  ( .D(\u_a23_mem/g_mem[16][0] ), .CLK(clk), 
        .RST(rst), .I(g_init[128]), .Q(\u_a23_mem/g_mem[16][0] ) );
  DFF \u_a23_mem/g_mem_reg[16][1]  ( .D(\u_a23_mem/g_mem[16][1] ), .CLK(clk), 
        .RST(rst), .I(g_init[129]), .Q(\u_a23_mem/g_mem[16][1] ) );
  DFF \u_a23_mem/g_mem_reg[16][2]  ( .D(\u_a23_mem/g_mem[16][2] ), .CLK(clk), 
        .RST(rst), .I(g_init[130]), .Q(\u_a23_mem/g_mem[16][2] ) );
  DFF \u_a23_mem/g_mem_reg[16][3]  ( .D(\u_a23_mem/g_mem[16][3] ), .CLK(clk), 
        .RST(rst), .I(g_init[131]), .Q(\u_a23_mem/g_mem[16][3] ) );
  DFF \u_a23_mem/g_mem_reg[16][4]  ( .D(\u_a23_mem/g_mem[16][4] ), .CLK(clk), 
        .RST(rst), .I(g_init[132]), .Q(\u_a23_mem/g_mem[16][4] ) );
  DFF \u_a23_mem/g_mem_reg[16][5]  ( .D(\u_a23_mem/g_mem[16][5] ), .CLK(clk), 
        .RST(rst), .I(g_init[133]), .Q(\u_a23_mem/g_mem[16][5] ) );
  DFF \u_a23_mem/g_mem_reg[16][6]  ( .D(\u_a23_mem/g_mem[16][6] ), .CLK(clk), 
        .RST(rst), .I(g_init[134]), .Q(\u_a23_mem/g_mem[16][6] ) );
  DFF \u_a23_mem/g_mem_reg[16][7]  ( .D(\u_a23_mem/g_mem[16][7] ), .CLK(clk), 
        .RST(rst), .I(g_init[135]), .Q(\u_a23_mem/g_mem[16][7] ) );
  DFF \u_a23_mem/g_mem_reg[17][0]  ( .D(\u_a23_mem/g_mem[17][0] ), .CLK(clk), 
        .RST(rst), .I(g_init[136]), .Q(\u_a23_mem/g_mem[17][0] ) );
  DFF \u_a23_mem/g_mem_reg[17][1]  ( .D(\u_a23_mem/g_mem[17][1] ), .CLK(clk), 
        .RST(rst), .I(g_init[137]), .Q(\u_a23_mem/g_mem[17][1] ) );
  DFF \u_a23_mem/g_mem_reg[17][2]  ( .D(\u_a23_mem/g_mem[17][2] ), .CLK(clk), 
        .RST(rst), .I(g_init[138]), .Q(\u_a23_mem/g_mem[17][2] ) );
  DFF \u_a23_mem/g_mem_reg[17][3]  ( .D(\u_a23_mem/g_mem[17][3] ), .CLK(clk), 
        .RST(rst), .I(g_init[139]), .Q(\u_a23_mem/g_mem[17][3] ) );
  DFF \u_a23_mem/g_mem_reg[17][4]  ( .D(\u_a23_mem/g_mem[17][4] ), .CLK(clk), 
        .RST(rst), .I(g_init[140]), .Q(\u_a23_mem/g_mem[17][4] ) );
  DFF \u_a23_mem/g_mem_reg[17][5]  ( .D(\u_a23_mem/g_mem[17][5] ), .CLK(clk), 
        .RST(rst), .I(g_init[141]), .Q(\u_a23_mem/g_mem[17][5] ) );
  DFF \u_a23_mem/g_mem_reg[17][6]  ( .D(\u_a23_mem/g_mem[17][6] ), .CLK(clk), 
        .RST(rst), .I(g_init[142]), .Q(\u_a23_mem/g_mem[17][6] ) );
  DFF \u_a23_mem/g_mem_reg[17][7]  ( .D(\u_a23_mem/g_mem[17][7] ), .CLK(clk), 
        .RST(rst), .I(g_init[143]), .Q(\u_a23_mem/g_mem[17][7] ) );
  DFF \u_a23_mem/g_mem_reg[18][0]  ( .D(\u_a23_mem/g_mem[18][0] ), .CLK(clk), 
        .RST(rst), .I(g_init[144]), .Q(\u_a23_mem/g_mem[18][0] ) );
  DFF \u_a23_mem/g_mem_reg[18][1]  ( .D(\u_a23_mem/g_mem[18][1] ), .CLK(clk), 
        .RST(rst), .I(g_init[145]), .Q(\u_a23_mem/g_mem[18][1] ) );
  DFF \u_a23_mem/g_mem_reg[18][2]  ( .D(\u_a23_mem/g_mem[18][2] ), .CLK(clk), 
        .RST(rst), .I(g_init[146]), .Q(\u_a23_mem/g_mem[18][2] ) );
  DFF \u_a23_mem/g_mem_reg[18][3]  ( .D(\u_a23_mem/g_mem[18][3] ), .CLK(clk), 
        .RST(rst), .I(g_init[147]), .Q(\u_a23_mem/g_mem[18][3] ) );
  DFF \u_a23_mem/g_mem_reg[18][4]  ( .D(\u_a23_mem/g_mem[18][4] ), .CLK(clk), 
        .RST(rst), .I(g_init[148]), .Q(\u_a23_mem/g_mem[18][4] ) );
  DFF \u_a23_mem/g_mem_reg[18][5]  ( .D(\u_a23_mem/g_mem[18][5] ), .CLK(clk), 
        .RST(rst), .I(g_init[149]), .Q(\u_a23_mem/g_mem[18][5] ) );
  DFF \u_a23_mem/g_mem_reg[18][6]  ( .D(\u_a23_mem/g_mem[18][6] ), .CLK(clk), 
        .RST(rst), .I(g_init[150]), .Q(\u_a23_mem/g_mem[18][6] ) );
  DFF \u_a23_mem/g_mem_reg[18][7]  ( .D(\u_a23_mem/g_mem[18][7] ), .CLK(clk), 
        .RST(rst), .I(g_init[151]), .Q(\u_a23_mem/g_mem[18][7] ) );
  DFF \u_a23_mem/g_mem_reg[19][0]  ( .D(\u_a23_mem/g_mem[19][0] ), .CLK(clk), 
        .RST(rst), .I(g_init[152]), .Q(\u_a23_mem/g_mem[19][0] ) );
  DFF \u_a23_mem/g_mem_reg[19][1]  ( .D(\u_a23_mem/g_mem[19][1] ), .CLK(clk), 
        .RST(rst), .I(g_init[153]), .Q(\u_a23_mem/g_mem[19][1] ) );
  DFF \u_a23_mem/g_mem_reg[19][2]  ( .D(\u_a23_mem/g_mem[19][2] ), .CLK(clk), 
        .RST(rst), .I(g_init[154]), .Q(\u_a23_mem/g_mem[19][2] ) );
  DFF \u_a23_mem/g_mem_reg[19][3]  ( .D(\u_a23_mem/g_mem[19][3] ), .CLK(clk), 
        .RST(rst), .I(g_init[155]), .Q(\u_a23_mem/g_mem[19][3] ) );
  DFF \u_a23_mem/g_mem_reg[19][4]  ( .D(\u_a23_mem/g_mem[19][4] ), .CLK(clk), 
        .RST(rst), .I(g_init[156]), .Q(\u_a23_mem/g_mem[19][4] ) );
  DFF \u_a23_mem/g_mem_reg[19][5]  ( .D(\u_a23_mem/g_mem[19][5] ), .CLK(clk), 
        .RST(rst), .I(g_init[157]), .Q(\u_a23_mem/g_mem[19][5] ) );
  DFF \u_a23_mem/g_mem_reg[19][6]  ( .D(\u_a23_mem/g_mem[19][6] ), .CLK(clk), 
        .RST(rst), .I(g_init[158]), .Q(\u_a23_mem/g_mem[19][6] ) );
  DFF \u_a23_mem/g_mem_reg[19][7]  ( .D(\u_a23_mem/g_mem[19][7] ), .CLK(clk), 
        .RST(rst), .I(g_init[159]), .Q(\u_a23_mem/g_mem[19][7] ) );
  DFF \u_a23_mem/g_mem_reg[20][0]  ( .D(\u_a23_mem/g_mem[20][0] ), .CLK(clk), 
        .RST(rst), .I(g_init[160]), .Q(\u_a23_mem/g_mem[20][0] ) );
  DFF \u_a23_mem/g_mem_reg[20][1]  ( .D(\u_a23_mem/g_mem[20][1] ), .CLK(clk), 
        .RST(rst), .I(g_init[161]), .Q(\u_a23_mem/g_mem[20][1] ) );
  DFF \u_a23_mem/g_mem_reg[20][2]  ( .D(\u_a23_mem/g_mem[20][2] ), .CLK(clk), 
        .RST(rst), .I(g_init[162]), .Q(\u_a23_mem/g_mem[20][2] ) );
  DFF \u_a23_mem/g_mem_reg[20][3]  ( .D(\u_a23_mem/g_mem[20][3] ), .CLK(clk), 
        .RST(rst), .I(g_init[163]), .Q(\u_a23_mem/g_mem[20][3] ) );
  DFF \u_a23_mem/g_mem_reg[20][4]  ( .D(\u_a23_mem/g_mem[20][4] ), .CLK(clk), 
        .RST(rst), .I(g_init[164]), .Q(\u_a23_mem/g_mem[20][4] ) );
  DFF \u_a23_mem/g_mem_reg[20][5]  ( .D(\u_a23_mem/g_mem[20][5] ), .CLK(clk), 
        .RST(rst), .I(g_init[165]), .Q(\u_a23_mem/g_mem[20][5] ) );
  DFF \u_a23_mem/g_mem_reg[20][6]  ( .D(\u_a23_mem/g_mem[20][6] ), .CLK(clk), 
        .RST(rst), .I(g_init[166]), .Q(\u_a23_mem/g_mem[20][6] ) );
  DFF \u_a23_mem/g_mem_reg[20][7]  ( .D(\u_a23_mem/g_mem[20][7] ), .CLK(clk), 
        .RST(rst), .I(g_init[167]), .Q(\u_a23_mem/g_mem[20][7] ) );
  DFF \u_a23_mem/g_mem_reg[21][0]  ( .D(\u_a23_mem/g_mem[21][0] ), .CLK(clk), 
        .RST(rst), .I(g_init[168]), .Q(\u_a23_mem/g_mem[21][0] ) );
  DFF \u_a23_mem/g_mem_reg[21][1]  ( .D(\u_a23_mem/g_mem[21][1] ), .CLK(clk), 
        .RST(rst), .I(g_init[169]), .Q(\u_a23_mem/g_mem[21][1] ) );
  DFF \u_a23_mem/g_mem_reg[21][2]  ( .D(\u_a23_mem/g_mem[21][2] ), .CLK(clk), 
        .RST(rst), .I(g_init[170]), .Q(\u_a23_mem/g_mem[21][2] ) );
  DFF \u_a23_mem/g_mem_reg[21][3]  ( .D(\u_a23_mem/g_mem[21][3] ), .CLK(clk), 
        .RST(rst), .I(g_init[171]), .Q(\u_a23_mem/g_mem[21][3] ) );
  DFF \u_a23_mem/g_mem_reg[21][4]  ( .D(\u_a23_mem/g_mem[21][4] ), .CLK(clk), 
        .RST(rst), .I(g_init[172]), .Q(\u_a23_mem/g_mem[21][4] ) );
  DFF \u_a23_mem/g_mem_reg[21][5]  ( .D(\u_a23_mem/g_mem[21][5] ), .CLK(clk), 
        .RST(rst), .I(g_init[173]), .Q(\u_a23_mem/g_mem[21][5] ) );
  DFF \u_a23_mem/g_mem_reg[21][6]  ( .D(\u_a23_mem/g_mem[21][6] ), .CLK(clk), 
        .RST(rst), .I(g_init[174]), .Q(\u_a23_mem/g_mem[21][6] ) );
  DFF \u_a23_mem/g_mem_reg[21][7]  ( .D(\u_a23_mem/g_mem[21][7] ), .CLK(clk), 
        .RST(rst), .I(g_init[175]), .Q(\u_a23_mem/g_mem[21][7] ) );
  DFF \u_a23_mem/g_mem_reg[22][0]  ( .D(\u_a23_mem/g_mem[22][0] ), .CLK(clk), 
        .RST(rst), .I(g_init[176]), .Q(\u_a23_mem/g_mem[22][0] ) );
  DFF \u_a23_mem/g_mem_reg[22][1]  ( .D(\u_a23_mem/g_mem[22][1] ), .CLK(clk), 
        .RST(rst), .I(g_init[177]), .Q(\u_a23_mem/g_mem[22][1] ) );
  DFF \u_a23_mem/g_mem_reg[22][2]  ( .D(\u_a23_mem/g_mem[22][2] ), .CLK(clk), 
        .RST(rst), .I(g_init[178]), .Q(\u_a23_mem/g_mem[22][2] ) );
  DFF \u_a23_mem/g_mem_reg[22][3]  ( .D(\u_a23_mem/g_mem[22][3] ), .CLK(clk), 
        .RST(rst), .I(g_init[179]), .Q(\u_a23_mem/g_mem[22][3] ) );
  DFF \u_a23_mem/g_mem_reg[22][4]  ( .D(\u_a23_mem/g_mem[22][4] ), .CLK(clk), 
        .RST(rst), .I(g_init[180]), .Q(\u_a23_mem/g_mem[22][4] ) );
  DFF \u_a23_mem/g_mem_reg[22][5]  ( .D(\u_a23_mem/g_mem[22][5] ), .CLK(clk), 
        .RST(rst), .I(g_init[181]), .Q(\u_a23_mem/g_mem[22][5] ) );
  DFF \u_a23_mem/g_mem_reg[22][6]  ( .D(\u_a23_mem/g_mem[22][6] ), .CLK(clk), 
        .RST(rst), .I(g_init[182]), .Q(\u_a23_mem/g_mem[22][6] ) );
  DFF \u_a23_mem/g_mem_reg[22][7]  ( .D(\u_a23_mem/g_mem[22][7] ), .CLK(clk), 
        .RST(rst), .I(g_init[183]), .Q(\u_a23_mem/g_mem[22][7] ) );
  DFF \u_a23_mem/g_mem_reg[23][0]  ( .D(\u_a23_mem/g_mem[23][0] ), .CLK(clk), 
        .RST(rst), .I(g_init[184]), .Q(\u_a23_mem/g_mem[23][0] ) );
  DFF \u_a23_mem/g_mem_reg[23][1]  ( .D(\u_a23_mem/g_mem[23][1] ), .CLK(clk), 
        .RST(rst), .I(g_init[185]), .Q(\u_a23_mem/g_mem[23][1] ) );
  DFF \u_a23_mem/g_mem_reg[23][2]  ( .D(\u_a23_mem/g_mem[23][2] ), .CLK(clk), 
        .RST(rst), .I(g_init[186]), .Q(\u_a23_mem/g_mem[23][2] ) );
  DFF \u_a23_mem/g_mem_reg[23][3]  ( .D(\u_a23_mem/g_mem[23][3] ), .CLK(clk), 
        .RST(rst), .I(g_init[187]), .Q(\u_a23_mem/g_mem[23][3] ) );
  DFF \u_a23_mem/g_mem_reg[23][4]  ( .D(\u_a23_mem/g_mem[23][4] ), .CLK(clk), 
        .RST(rst), .I(g_init[188]), .Q(\u_a23_mem/g_mem[23][4] ) );
  DFF \u_a23_mem/g_mem_reg[23][5]  ( .D(\u_a23_mem/g_mem[23][5] ), .CLK(clk), 
        .RST(rst), .I(g_init[189]), .Q(\u_a23_mem/g_mem[23][5] ) );
  DFF \u_a23_mem/g_mem_reg[23][6]  ( .D(\u_a23_mem/g_mem[23][6] ), .CLK(clk), 
        .RST(rst), .I(g_init[190]), .Q(\u_a23_mem/g_mem[23][6] ) );
  DFF \u_a23_mem/g_mem_reg[23][7]  ( .D(\u_a23_mem/g_mem[23][7] ), .CLK(clk), 
        .RST(rst), .I(g_init[191]), .Q(\u_a23_mem/g_mem[23][7] ) );
  DFF \u_a23_mem/g_mem_reg[24][0]  ( .D(\u_a23_mem/g_mem[24][0] ), .CLK(clk), 
        .RST(rst), .I(g_init[192]), .Q(\u_a23_mem/g_mem[24][0] ) );
  DFF \u_a23_mem/g_mem_reg[24][1]  ( .D(\u_a23_mem/g_mem[24][1] ), .CLK(clk), 
        .RST(rst), .I(g_init[193]), .Q(\u_a23_mem/g_mem[24][1] ) );
  DFF \u_a23_mem/g_mem_reg[24][2]  ( .D(\u_a23_mem/g_mem[24][2] ), .CLK(clk), 
        .RST(rst), .I(g_init[194]), .Q(\u_a23_mem/g_mem[24][2] ) );
  DFF \u_a23_mem/g_mem_reg[24][3]  ( .D(\u_a23_mem/g_mem[24][3] ), .CLK(clk), 
        .RST(rst), .I(g_init[195]), .Q(\u_a23_mem/g_mem[24][3] ) );
  DFF \u_a23_mem/g_mem_reg[24][4]  ( .D(\u_a23_mem/g_mem[24][4] ), .CLK(clk), 
        .RST(rst), .I(g_init[196]), .Q(\u_a23_mem/g_mem[24][4] ) );
  DFF \u_a23_mem/g_mem_reg[24][5]  ( .D(\u_a23_mem/g_mem[24][5] ), .CLK(clk), 
        .RST(rst), .I(g_init[197]), .Q(\u_a23_mem/g_mem[24][5] ) );
  DFF \u_a23_mem/g_mem_reg[24][6]  ( .D(\u_a23_mem/g_mem[24][6] ), .CLK(clk), 
        .RST(rst), .I(g_init[198]), .Q(\u_a23_mem/g_mem[24][6] ) );
  DFF \u_a23_mem/g_mem_reg[24][7]  ( .D(\u_a23_mem/g_mem[24][7] ), .CLK(clk), 
        .RST(rst), .I(g_init[199]), .Q(\u_a23_mem/g_mem[24][7] ) );
  DFF \u_a23_mem/g_mem_reg[25][0]  ( .D(\u_a23_mem/g_mem[25][0] ), .CLK(clk), 
        .RST(rst), .I(g_init[200]), .Q(\u_a23_mem/g_mem[25][0] ) );
  DFF \u_a23_mem/g_mem_reg[25][1]  ( .D(\u_a23_mem/g_mem[25][1] ), .CLK(clk), 
        .RST(rst), .I(g_init[201]), .Q(\u_a23_mem/g_mem[25][1] ) );
  DFF \u_a23_mem/g_mem_reg[25][2]  ( .D(\u_a23_mem/g_mem[25][2] ), .CLK(clk), 
        .RST(rst), .I(g_init[202]), .Q(\u_a23_mem/g_mem[25][2] ) );
  DFF \u_a23_mem/g_mem_reg[25][3]  ( .D(\u_a23_mem/g_mem[25][3] ), .CLK(clk), 
        .RST(rst), .I(g_init[203]), .Q(\u_a23_mem/g_mem[25][3] ) );
  DFF \u_a23_mem/g_mem_reg[25][4]  ( .D(\u_a23_mem/g_mem[25][4] ), .CLK(clk), 
        .RST(rst), .I(g_init[204]), .Q(\u_a23_mem/g_mem[25][4] ) );
  DFF \u_a23_mem/g_mem_reg[25][5]  ( .D(\u_a23_mem/g_mem[25][5] ), .CLK(clk), 
        .RST(rst), .I(g_init[205]), .Q(\u_a23_mem/g_mem[25][5] ) );
  DFF \u_a23_mem/g_mem_reg[25][6]  ( .D(\u_a23_mem/g_mem[25][6] ), .CLK(clk), 
        .RST(rst), .I(g_init[206]), .Q(\u_a23_mem/g_mem[25][6] ) );
  DFF \u_a23_mem/g_mem_reg[25][7]  ( .D(\u_a23_mem/g_mem[25][7] ), .CLK(clk), 
        .RST(rst), .I(g_init[207]), .Q(\u_a23_mem/g_mem[25][7] ) );
  DFF \u_a23_mem/g_mem_reg[26][0]  ( .D(\u_a23_mem/g_mem[26][0] ), .CLK(clk), 
        .RST(rst), .I(g_init[208]), .Q(\u_a23_mem/g_mem[26][0] ) );
  DFF \u_a23_mem/g_mem_reg[26][1]  ( .D(\u_a23_mem/g_mem[26][1] ), .CLK(clk), 
        .RST(rst), .I(g_init[209]), .Q(\u_a23_mem/g_mem[26][1] ) );
  DFF \u_a23_mem/g_mem_reg[26][2]  ( .D(\u_a23_mem/g_mem[26][2] ), .CLK(clk), 
        .RST(rst), .I(g_init[210]), .Q(\u_a23_mem/g_mem[26][2] ) );
  DFF \u_a23_mem/g_mem_reg[26][3]  ( .D(\u_a23_mem/g_mem[26][3] ), .CLK(clk), 
        .RST(rst), .I(g_init[211]), .Q(\u_a23_mem/g_mem[26][3] ) );
  DFF \u_a23_mem/g_mem_reg[26][4]  ( .D(\u_a23_mem/g_mem[26][4] ), .CLK(clk), 
        .RST(rst), .I(g_init[212]), .Q(\u_a23_mem/g_mem[26][4] ) );
  DFF \u_a23_mem/g_mem_reg[26][5]  ( .D(\u_a23_mem/g_mem[26][5] ), .CLK(clk), 
        .RST(rst), .I(g_init[213]), .Q(\u_a23_mem/g_mem[26][5] ) );
  DFF \u_a23_mem/g_mem_reg[26][6]  ( .D(\u_a23_mem/g_mem[26][6] ), .CLK(clk), 
        .RST(rst), .I(g_init[214]), .Q(\u_a23_mem/g_mem[26][6] ) );
  DFF \u_a23_mem/g_mem_reg[26][7]  ( .D(\u_a23_mem/g_mem[26][7] ), .CLK(clk), 
        .RST(rst), .I(g_init[215]), .Q(\u_a23_mem/g_mem[26][7] ) );
  DFF \u_a23_mem/g_mem_reg[27][0]  ( .D(\u_a23_mem/g_mem[27][0] ), .CLK(clk), 
        .RST(rst), .I(g_init[216]), .Q(\u_a23_mem/g_mem[27][0] ) );
  DFF \u_a23_mem/g_mem_reg[27][1]  ( .D(\u_a23_mem/g_mem[27][1] ), .CLK(clk), 
        .RST(rst), .I(g_init[217]), .Q(\u_a23_mem/g_mem[27][1] ) );
  DFF \u_a23_mem/g_mem_reg[27][2]  ( .D(\u_a23_mem/g_mem[27][2] ), .CLK(clk), 
        .RST(rst), .I(g_init[218]), .Q(\u_a23_mem/g_mem[27][2] ) );
  DFF \u_a23_mem/g_mem_reg[27][3]  ( .D(\u_a23_mem/g_mem[27][3] ), .CLK(clk), 
        .RST(rst), .I(g_init[219]), .Q(\u_a23_mem/g_mem[27][3] ) );
  DFF \u_a23_mem/g_mem_reg[27][4]  ( .D(\u_a23_mem/g_mem[27][4] ), .CLK(clk), 
        .RST(rst), .I(g_init[220]), .Q(\u_a23_mem/g_mem[27][4] ) );
  DFF \u_a23_mem/g_mem_reg[27][5]  ( .D(\u_a23_mem/g_mem[27][5] ), .CLK(clk), 
        .RST(rst), .I(g_init[221]), .Q(\u_a23_mem/g_mem[27][5] ) );
  DFF \u_a23_mem/g_mem_reg[27][6]  ( .D(\u_a23_mem/g_mem[27][6] ), .CLK(clk), 
        .RST(rst), .I(g_init[222]), .Q(\u_a23_mem/g_mem[27][6] ) );
  DFF \u_a23_mem/g_mem_reg[27][7]  ( .D(\u_a23_mem/g_mem[27][7] ), .CLK(clk), 
        .RST(rst), .I(g_init[223]), .Q(\u_a23_mem/g_mem[27][7] ) );
  DFF \u_a23_mem/g_mem_reg[28][0]  ( .D(\u_a23_mem/g_mem[28][0] ), .CLK(clk), 
        .RST(rst), .I(g_init[224]), .Q(\u_a23_mem/g_mem[28][0] ) );
  DFF \u_a23_mem/g_mem_reg[28][1]  ( .D(\u_a23_mem/g_mem[28][1] ), .CLK(clk), 
        .RST(rst), .I(g_init[225]), .Q(\u_a23_mem/g_mem[28][1] ) );
  DFF \u_a23_mem/g_mem_reg[28][2]  ( .D(\u_a23_mem/g_mem[28][2] ), .CLK(clk), 
        .RST(rst), .I(g_init[226]), .Q(\u_a23_mem/g_mem[28][2] ) );
  DFF \u_a23_mem/g_mem_reg[28][3]  ( .D(\u_a23_mem/g_mem[28][3] ), .CLK(clk), 
        .RST(rst), .I(g_init[227]), .Q(\u_a23_mem/g_mem[28][3] ) );
  DFF \u_a23_mem/g_mem_reg[28][4]  ( .D(\u_a23_mem/g_mem[28][4] ), .CLK(clk), 
        .RST(rst), .I(g_init[228]), .Q(\u_a23_mem/g_mem[28][4] ) );
  DFF \u_a23_mem/g_mem_reg[28][5]  ( .D(\u_a23_mem/g_mem[28][5] ), .CLK(clk), 
        .RST(rst), .I(g_init[229]), .Q(\u_a23_mem/g_mem[28][5] ) );
  DFF \u_a23_mem/g_mem_reg[28][6]  ( .D(\u_a23_mem/g_mem[28][6] ), .CLK(clk), 
        .RST(rst), .I(g_init[230]), .Q(\u_a23_mem/g_mem[28][6] ) );
  DFF \u_a23_mem/g_mem_reg[28][7]  ( .D(\u_a23_mem/g_mem[28][7] ), .CLK(clk), 
        .RST(rst), .I(g_init[231]), .Q(\u_a23_mem/g_mem[28][7] ) );
  DFF \u_a23_mem/g_mem_reg[29][0]  ( .D(\u_a23_mem/g_mem[29][0] ), .CLK(clk), 
        .RST(rst), .I(g_init[232]), .Q(\u_a23_mem/g_mem[29][0] ) );
  DFF \u_a23_mem/g_mem_reg[29][1]  ( .D(\u_a23_mem/g_mem[29][1] ), .CLK(clk), 
        .RST(rst), .I(g_init[233]), .Q(\u_a23_mem/g_mem[29][1] ) );
  DFF \u_a23_mem/g_mem_reg[29][2]  ( .D(\u_a23_mem/g_mem[29][2] ), .CLK(clk), 
        .RST(rst), .I(g_init[234]), .Q(\u_a23_mem/g_mem[29][2] ) );
  DFF \u_a23_mem/g_mem_reg[29][3]  ( .D(\u_a23_mem/g_mem[29][3] ), .CLK(clk), 
        .RST(rst), .I(g_init[235]), .Q(\u_a23_mem/g_mem[29][3] ) );
  DFF \u_a23_mem/g_mem_reg[29][4]  ( .D(\u_a23_mem/g_mem[29][4] ), .CLK(clk), 
        .RST(rst), .I(g_init[236]), .Q(\u_a23_mem/g_mem[29][4] ) );
  DFF \u_a23_mem/g_mem_reg[29][5]  ( .D(\u_a23_mem/g_mem[29][5] ), .CLK(clk), 
        .RST(rst), .I(g_init[237]), .Q(\u_a23_mem/g_mem[29][5] ) );
  DFF \u_a23_mem/g_mem_reg[29][6]  ( .D(\u_a23_mem/g_mem[29][6] ), .CLK(clk), 
        .RST(rst), .I(g_init[238]), .Q(\u_a23_mem/g_mem[29][6] ) );
  DFF \u_a23_mem/g_mem_reg[29][7]  ( .D(\u_a23_mem/g_mem[29][7] ), .CLK(clk), 
        .RST(rst), .I(g_init[239]), .Q(\u_a23_mem/g_mem[29][7] ) );
  DFF \u_a23_mem/g_mem_reg[30][0]  ( .D(\u_a23_mem/g_mem[30][0] ), .CLK(clk), 
        .RST(rst), .I(g_init[240]), .Q(\u_a23_mem/g_mem[30][0] ) );
  DFF \u_a23_mem/g_mem_reg[30][1]  ( .D(\u_a23_mem/g_mem[30][1] ), .CLK(clk), 
        .RST(rst), .I(g_init[241]), .Q(\u_a23_mem/g_mem[30][1] ) );
  DFF \u_a23_mem/g_mem_reg[30][2]  ( .D(\u_a23_mem/g_mem[30][2] ), .CLK(clk), 
        .RST(rst), .I(g_init[242]), .Q(\u_a23_mem/g_mem[30][2] ) );
  DFF \u_a23_mem/g_mem_reg[30][3]  ( .D(\u_a23_mem/g_mem[30][3] ), .CLK(clk), 
        .RST(rst), .I(g_init[243]), .Q(\u_a23_mem/g_mem[30][3] ) );
  DFF \u_a23_mem/g_mem_reg[30][4]  ( .D(\u_a23_mem/g_mem[30][4] ), .CLK(clk), 
        .RST(rst), .I(g_init[244]), .Q(\u_a23_mem/g_mem[30][4] ) );
  DFF \u_a23_mem/g_mem_reg[30][5]  ( .D(\u_a23_mem/g_mem[30][5] ), .CLK(clk), 
        .RST(rst), .I(g_init[245]), .Q(\u_a23_mem/g_mem[30][5] ) );
  DFF \u_a23_mem/g_mem_reg[30][6]  ( .D(\u_a23_mem/g_mem[30][6] ), .CLK(clk), 
        .RST(rst), .I(g_init[246]), .Q(\u_a23_mem/g_mem[30][6] ) );
  DFF \u_a23_mem/g_mem_reg[30][7]  ( .D(\u_a23_mem/g_mem[30][7] ), .CLK(clk), 
        .RST(rst), .I(g_init[247]), .Q(\u_a23_mem/g_mem[30][7] ) );
  DFF \u_a23_mem/g_mem_reg[31][0]  ( .D(\u_a23_mem/g_mem[31][0] ), .CLK(clk), 
        .RST(rst), .I(g_init[248]), .Q(\u_a23_mem/g_mem[31][0] ) );
  DFF \u_a23_mem/g_mem_reg[31][1]  ( .D(\u_a23_mem/g_mem[31][1] ), .CLK(clk), 
        .RST(rst), .I(g_init[249]), .Q(\u_a23_mem/g_mem[31][1] ) );
  DFF \u_a23_mem/g_mem_reg[31][2]  ( .D(\u_a23_mem/g_mem[31][2] ), .CLK(clk), 
        .RST(rst), .I(g_init[250]), .Q(\u_a23_mem/g_mem[31][2] ) );
  DFF \u_a23_mem/g_mem_reg[31][3]  ( .D(\u_a23_mem/g_mem[31][3] ), .CLK(clk), 
        .RST(rst), .I(g_init[251]), .Q(\u_a23_mem/g_mem[31][3] ) );
  DFF \u_a23_mem/g_mem_reg[31][4]  ( .D(\u_a23_mem/g_mem[31][4] ), .CLK(clk), 
        .RST(rst), .I(g_init[252]), .Q(\u_a23_mem/g_mem[31][4] ) );
  DFF \u_a23_mem/g_mem_reg[31][5]  ( .D(\u_a23_mem/g_mem[31][5] ), .CLK(clk), 
        .RST(rst), .I(g_init[253]), .Q(\u_a23_mem/g_mem[31][5] ) );
  DFF \u_a23_mem/g_mem_reg[31][6]  ( .D(\u_a23_mem/g_mem[31][6] ), .CLK(clk), 
        .RST(rst), .I(g_init[254]), .Q(\u_a23_mem/g_mem[31][6] ) );
  DFF \u_a23_mem/g_mem_reg[31][7]  ( .D(\u_a23_mem/g_mem[31][7] ), .CLK(clk), 
        .RST(rst), .I(g_init[255]), .Q(\u_a23_mem/g_mem[31][7] ) );
  DFF \u_a23_mem/e_mem_reg[0][0]  ( .D(\u_a23_mem/e_mem[0][0] ), .CLK(clk), 
        .RST(rst), .I(e_init[0]), .Q(\u_a23_mem/e_mem[0][0] ) );
  DFF \u_a23_mem/e_mem_reg[0][1]  ( .D(\u_a23_mem/e_mem[0][1] ), .CLK(clk), 
        .RST(rst), .I(e_init[1]), .Q(\u_a23_mem/e_mem[0][1] ) );
  DFF \u_a23_mem/e_mem_reg[0][2]  ( .D(\u_a23_mem/e_mem[0][2] ), .CLK(clk), 
        .RST(rst), .I(e_init[2]), .Q(\u_a23_mem/e_mem[0][2] ) );
  DFF \u_a23_mem/e_mem_reg[0][3]  ( .D(\u_a23_mem/e_mem[0][3] ), .CLK(clk), 
        .RST(rst), .I(e_init[3]), .Q(\u_a23_mem/e_mem[0][3] ) );
  DFF \u_a23_mem/e_mem_reg[0][4]  ( .D(\u_a23_mem/e_mem[0][4] ), .CLK(clk), 
        .RST(rst), .I(e_init[4]), .Q(\u_a23_mem/e_mem[0][4] ) );
  DFF \u_a23_mem/e_mem_reg[0][5]  ( .D(\u_a23_mem/e_mem[0][5] ), .CLK(clk), 
        .RST(rst), .I(e_init[5]), .Q(\u_a23_mem/e_mem[0][5] ) );
  DFF \u_a23_mem/e_mem_reg[0][6]  ( .D(\u_a23_mem/e_mem[0][6] ), .CLK(clk), 
        .RST(rst), .I(e_init[6]), .Q(\u_a23_mem/e_mem[0][6] ) );
  DFF \u_a23_mem/e_mem_reg[0][7]  ( .D(\u_a23_mem/e_mem[0][7] ), .CLK(clk), 
        .RST(rst), .I(e_init[7]), .Q(\u_a23_mem/e_mem[0][7] ) );
  DFF \u_a23_mem/e_mem_reg[1][0]  ( .D(\u_a23_mem/e_mem[1][0] ), .CLK(clk), 
        .RST(rst), .I(e_init[8]), .Q(\u_a23_mem/e_mem[1][0] ) );
  DFF \u_a23_mem/e_mem_reg[1][1]  ( .D(\u_a23_mem/e_mem[1][1] ), .CLK(clk), 
        .RST(rst), .I(e_init[9]), .Q(\u_a23_mem/e_mem[1][1] ) );
  DFF \u_a23_mem/e_mem_reg[1][2]  ( .D(\u_a23_mem/e_mem[1][2] ), .CLK(clk), 
        .RST(rst), .I(e_init[10]), .Q(\u_a23_mem/e_mem[1][2] ) );
  DFF \u_a23_mem/e_mem_reg[1][3]  ( .D(\u_a23_mem/e_mem[1][3] ), .CLK(clk), 
        .RST(rst), .I(e_init[11]), .Q(\u_a23_mem/e_mem[1][3] ) );
  DFF \u_a23_mem/e_mem_reg[1][4]  ( .D(\u_a23_mem/e_mem[1][4] ), .CLK(clk), 
        .RST(rst), .I(e_init[12]), .Q(\u_a23_mem/e_mem[1][4] ) );
  DFF \u_a23_mem/e_mem_reg[1][5]  ( .D(\u_a23_mem/e_mem[1][5] ), .CLK(clk), 
        .RST(rst), .I(e_init[13]), .Q(\u_a23_mem/e_mem[1][5] ) );
  DFF \u_a23_mem/e_mem_reg[1][6]  ( .D(\u_a23_mem/e_mem[1][6] ), .CLK(clk), 
        .RST(rst), .I(e_init[14]), .Q(\u_a23_mem/e_mem[1][6] ) );
  DFF \u_a23_mem/e_mem_reg[1][7]  ( .D(\u_a23_mem/e_mem[1][7] ), .CLK(clk), 
        .RST(rst), .I(e_init[15]), .Q(\u_a23_mem/e_mem[1][7] ) );
  DFF \u_a23_mem/e_mem_reg[2][0]  ( .D(\u_a23_mem/e_mem[2][0] ), .CLK(clk), 
        .RST(rst), .I(e_init[16]), .Q(\u_a23_mem/e_mem[2][0] ) );
  DFF \u_a23_mem/e_mem_reg[2][1]  ( .D(\u_a23_mem/e_mem[2][1] ), .CLK(clk), 
        .RST(rst), .I(e_init[17]), .Q(\u_a23_mem/e_mem[2][1] ) );
  DFF \u_a23_mem/e_mem_reg[2][2]  ( .D(\u_a23_mem/e_mem[2][2] ), .CLK(clk), 
        .RST(rst), .I(e_init[18]), .Q(\u_a23_mem/e_mem[2][2] ) );
  DFF \u_a23_mem/e_mem_reg[2][3]  ( .D(\u_a23_mem/e_mem[2][3] ), .CLK(clk), 
        .RST(rst), .I(e_init[19]), .Q(\u_a23_mem/e_mem[2][3] ) );
  DFF \u_a23_mem/e_mem_reg[2][4]  ( .D(\u_a23_mem/e_mem[2][4] ), .CLK(clk), 
        .RST(rst), .I(e_init[20]), .Q(\u_a23_mem/e_mem[2][4] ) );
  DFF \u_a23_mem/e_mem_reg[2][5]  ( .D(\u_a23_mem/e_mem[2][5] ), .CLK(clk), 
        .RST(rst), .I(e_init[21]), .Q(\u_a23_mem/e_mem[2][5] ) );
  DFF \u_a23_mem/e_mem_reg[2][6]  ( .D(\u_a23_mem/e_mem[2][6] ), .CLK(clk), 
        .RST(rst), .I(e_init[22]), .Q(\u_a23_mem/e_mem[2][6] ) );
  DFF \u_a23_mem/e_mem_reg[2][7]  ( .D(\u_a23_mem/e_mem[2][7] ), .CLK(clk), 
        .RST(rst), .I(e_init[23]), .Q(\u_a23_mem/e_mem[2][7] ) );
  DFF \u_a23_mem/e_mem_reg[3][0]  ( .D(\u_a23_mem/e_mem[3][0] ), .CLK(clk), 
        .RST(rst), .I(e_init[24]), .Q(\u_a23_mem/e_mem[3][0] ) );
  DFF \u_a23_mem/e_mem_reg[3][1]  ( .D(\u_a23_mem/e_mem[3][1] ), .CLK(clk), 
        .RST(rst), .I(e_init[25]), .Q(\u_a23_mem/e_mem[3][1] ) );
  DFF \u_a23_mem/e_mem_reg[3][2]  ( .D(\u_a23_mem/e_mem[3][2] ), .CLK(clk), 
        .RST(rst), .I(e_init[26]), .Q(\u_a23_mem/e_mem[3][2] ) );
  DFF \u_a23_mem/e_mem_reg[3][3]  ( .D(\u_a23_mem/e_mem[3][3] ), .CLK(clk), 
        .RST(rst), .I(e_init[27]), .Q(\u_a23_mem/e_mem[3][3] ) );
  DFF \u_a23_mem/e_mem_reg[3][4]  ( .D(\u_a23_mem/e_mem[3][4] ), .CLK(clk), 
        .RST(rst), .I(e_init[28]), .Q(\u_a23_mem/e_mem[3][4] ) );
  DFF \u_a23_mem/e_mem_reg[3][5]  ( .D(\u_a23_mem/e_mem[3][5] ), .CLK(clk), 
        .RST(rst), .I(e_init[29]), .Q(\u_a23_mem/e_mem[3][5] ) );
  DFF \u_a23_mem/e_mem_reg[3][6]  ( .D(\u_a23_mem/e_mem[3][6] ), .CLK(clk), 
        .RST(rst), .I(e_init[30]), .Q(\u_a23_mem/e_mem[3][6] ) );
  DFF \u_a23_mem/e_mem_reg[3][7]  ( .D(\u_a23_mem/e_mem[3][7] ), .CLK(clk), 
        .RST(rst), .I(e_init[31]), .Q(\u_a23_mem/e_mem[3][7] ) );
  DFF \u_a23_mem/e_mem_reg[4][0]  ( .D(\u_a23_mem/e_mem[4][0] ), .CLK(clk), 
        .RST(rst), .I(e_init[32]), .Q(\u_a23_mem/e_mem[4][0] ) );
  DFF \u_a23_mem/e_mem_reg[4][1]  ( .D(\u_a23_mem/e_mem[4][1] ), .CLK(clk), 
        .RST(rst), .I(e_init[33]), .Q(\u_a23_mem/e_mem[4][1] ) );
  DFF \u_a23_mem/e_mem_reg[4][2]  ( .D(\u_a23_mem/e_mem[4][2] ), .CLK(clk), 
        .RST(rst), .I(e_init[34]), .Q(\u_a23_mem/e_mem[4][2] ) );
  DFF \u_a23_mem/e_mem_reg[4][3]  ( .D(\u_a23_mem/e_mem[4][3] ), .CLK(clk), 
        .RST(rst), .I(e_init[35]), .Q(\u_a23_mem/e_mem[4][3] ) );
  DFF \u_a23_mem/e_mem_reg[4][4]  ( .D(\u_a23_mem/e_mem[4][4] ), .CLK(clk), 
        .RST(rst), .I(e_init[36]), .Q(\u_a23_mem/e_mem[4][4] ) );
  DFF \u_a23_mem/e_mem_reg[4][5]  ( .D(\u_a23_mem/e_mem[4][5] ), .CLK(clk), 
        .RST(rst), .I(e_init[37]), .Q(\u_a23_mem/e_mem[4][5] ) );
  DFF \u_a23_mem/e_mem_reg[4][6]  ( .D(\u_a23_mem/e_mem[4][6] ), .CLK(clk), 
        .RST(rst), .I(e_init[38]), .Q(\u_a23_mem/e_mem[4][6] ) );
  DFF \u_a23_mem/e_mem_reg[4][7]  ( .D(\u_a23_mem/e_mem[4][7] ), .CLK(clk), 
        .RST(rst), .I(e_init[39]), .Q(\u_a23_mem/e_mem[4][7] ) );
  DFF \u_a23_mem/e_mem_reg[5][0]  ( .D(\u_a23_mem/e_mem[5][0] ), .CLK(clk), 
        .RST(rst), .I(e_init[40]), .Q(\u_a23_mem/e_mem[5][0] ) );
  DFF \u_a23_mem/e_mem_reg[5][1]  ( .D(\u_a23_mem/e_mem[5][1] ), .CLK(clk), 
        .RST(rst), .I(e_init[41]), .Q(\u_a23_mem/e_mem[5][1] ) );
  DFF \u_a23_mem/e_mem_reg[5][2]  ( .D(\u_a23_mem/e_mem[5][2] ), .CLK(clk), 
        .RST(rst), .I(e_init[42]), .Q(\u_a23_mem/e_mem[5][2] ) );
  DFF \u_a23_mem/e_mem_reg[5][3]  ( .D(\u_a23_mem/e_mem[5][3] ), .CLK(clk), 
        .RST(rst), .I(e_init[43]), .Q(\u_a23_mem/e_mem[5][3] ) );
  DFF \u_a23_mem/e_mem_reg[5][4]  ( .D(\u_a23_mem/e_mem[5][4] ), .CLK(clk), 
        .RST(rst), .I(e_init[44]), .Q(\u_a23_mem/e_mem[5][4] ) );
  DFF \u_a23_mem/e_mem_reg[5][5]  ( .D(\u_a23_mem/e_mem[5][5] ), .CLK(clk), 
        .RST(rst), .I(e_init[45]), .Q(\u_a23_mem/e_mem[5][5] ) );
  DFF \u_a23_mem/e_mem_reg[5][6]  ( .D(\u_a23_mem/e_mem[5][6] ), .CLK(clk), 
        .RST(rst), .I(e_init[46]), .Q(\u_a23_mem/e_mem[5][6] ) );
  DFF \u_a23_mem/e_mem_reg[5][7]  ( .D(\u_a23_mem/e_mem[5][7] ), .CLK(clk), 
        .RST(rst), .I(e_init[47]), .Q(\u_a23_mem/e_mem[5][7] ) );
  DFF \u_a23_mem/e_mem_reg[6][0]  ( .D(\u_a23_mem/e_mem[6][0] ), .CLK(clk), 
        .RST(rst), .I(e_init[48]), .Q(\u_a23_mem/e_mem[6][0] ) );
  DFF \u_a23_mem/e_mem_reg[6][1]  ( .D(\u_a23_mem/e_mem[6][1] ), .CLK(clk), 
        .RST(rst), .I(e_init[49]), .Q(\u_a23_mem/e_mem[6][1] ) );
  DFF \u_a23_mem/e_mem_reg[6][2]  ( .D(\u_a23_mem/e_mem[6][2] ), .CLK(clk), 
        .RST(rst), .I(e_init[50]), .Q(\u_a23_mem/e_mem[6][2] ) );
  DFF \u_a23_mem/e_mem_reg[6][3]  ( .D(\u_a23_mem/e_mem[6][3] ), .CLK(clk), 
        .RST(rst), .I(e_init[51]), .Q(\u_a23_mem/e_mem[6][3] ) );
  DFF \u_a23_mem/e_mem_reg[6][4]  ( .D(\u_a23_mem/e_mem[6][4] ), .CLK(clk), 
        .RST(rst), .I(e_init[52]), .Q(\u_a23_mem/e_mem[6][4] ) );
  DFF \u_a23_mem/e_mem_reg[6][5]  ( .D(\u_a23_mem/e_mem[6][5] ), .CLK(clk), 
        .RST(rst), .I(e_init[53]), .Q(\u_a23_mem/e_mem[6][5] ) );
  DFF \u_a23_mem/e_mem_reg[6][6]  ( .D(\u_a23_mem/e_mem[6][6] ), .CLK(clk), 
        .RST(rst), .I(e_init[54]), .Q(\u_a23_mem/e_mem[6][6] ) );
  DFF \u_a23_mem/e_mem_reg[6][7]  ( .D(\u_a23_mem/e_mem[6][7] ), .CLK(clk), 
        .RST(rst), .I(e_init[55]), .Q(\u_a23_mem/e_mem[6][7] ) );
  DFF \u_a23_mem/e_mem_reg[7][0]  ( .D(\u_a23_mem/e_mem[7][0] ), .CLK(clk), 
        .RST(rst), .I(e_init[56]), .Q(\u_a23_mem/e_mem[7][0] ) );
  DFF \u_a23_mem/e_mem_reg[7][1]  ( .D(\u_a23_mem/e_mem[7][1] ), .CLK(clk), 
        .RST(rst), .I(e_init[57]), .Q(\u_a23_mem/e_mem[7][1] ) );
  DFF \u_a23_mem/e_mem_reg[7][2]  ( .D(\u_a23_mem/e_mem[7][2] ), .CLK(clk), 
        .RST(rst), .I(e_init[58]), .Q(\u_a23_mem/e_mem[7][2] ) );
  DFF \u_a23_mem/e_mem_reg[7][3]  ( .D(\u_a23_mem/e_mem[7][3] ), .CLK(clk), 
        .RST(rst), .I(e_init[59]), .Q(\u_a23_mem/e_mem[7][3] ) );
  DFF \u_a23_mem/e_mem_reg[7][4]  ( .D(\u_a23_mem/e_mem[7][4] ), .CLK(clk), 
        .RST(rst), .I(e_init[60]), .Q(\u_a23_mem/e_mem[7][4] ) );
  DFF \u_a23_mem/e_mem_reg[7][5]  ( .D(\u_a23_mem/e_mem[7][5] ), .CLK(clk), 
        .RST(rst), .I(e_init[61]), .Q(\u_a23_mem/e_mem[7][5] ) );
  DFF \u_a23_mem/e_mem_reg[7][6]  ( .D(\u_a23_mem/e_mem[7][6] ), .CLK(clk), 
        .RST(rst), .I(e_init[62]), .Q(\u_a23_mem/e_mem[7][6] ) );
  DFF \u_a23_mem/e_mem_reg[7][7]  ( .D(\u_a23_mem/e_mem[7][7] ), .CLK(clk), 
        .RST(rst), .I(e_init[63]), .Q(\u_a23_mem/e_mem[7][7] ) );
  DFF \u_a23_mem/e_mem_reg[8][0]  ( .D(\u_a23_mem/e_mem[8][0] ), .CLK(clk), 
        .RST(rst), .I(e_init[64]), .Q(\u_a23_mem/e_mem[8][0] ) );
  DFF \u_a23_mem/e_mem_reg[8][1]  ( .D(\u_a23_mem/e_mem[8][1] ), .CLK(clk), 
        .RST(rst), .I(e_init[65]), .Q(\u_a23_mem/e_mem[8][1] ) );
  DFF \u_a23_mem/e_mem_reg[8][2]  ( .D(\u_a23_mem/e_mem[8][2] ), .CLK(clk), 
        .RST(rst), .I(e_init[66]), .Q(\u_a23_mem/e_mem[8][2] ) );
  DFF \u_a23_mem/e_mem_reg[8][3]  ( .D(\u_a23_mem/e_mem[8][3] ), .CLK(clk), 
        .RST(rst), .I(e_init[67]), .Q(\u_a23_mem/e_mem[8][3] ) );
  DFF \u_a23_mem/e_mem_reg[8][4]  ( .D(\u_a23_mem/e_mem[8][4] ), .CLK(clk), 
        .RST(rst), .I(e_init[68]), .Q(\u_a23_mem/e_mem[8][4] ) );
  DFF \u_a23_mem/e_mem_reg[8][5]  ( .D(\u_a23_mem/e_mem[8][5] ), .CLK(clk), 
        .RST(rst), .I(e_init[69]), .Q(\u_a23_mem/e_mem[8][5] ) );
  DFF \u_a23_mem/e_mem_reg[8][6]  ( .D(\u_a23_mem/e_mem[8][6] ), .CLK(clk), 
        .RST(rst), .I(e_init[70]), .Q(\u_a23_mem/e_mem[8][6] ) );
  DFF \u_a23_mem/e_mem_reg[8][7]  ( .D(\u_a23_mem/e_mem[8][7] ), .CLK(clk), 
        .RST(rst), .I(e_init[71]), .Q(\u_a23_mem/e_mem[8][7] ) );
  DFF \u_a23_mem/e_mem_reg[9][0]  ( .D(\u_a23_mem/e_mem[9][0] ), .CLK(clk), 
        .RST(rst), .I(e_init[72]), .Q(\u_a23_mem/e_mem[9][0] ) );
  DFF \u_a23_mem/e_mem_reg[9][1]  ( .D(\u_a23_mem/e_mem[9][1] ), .CLK(clk), 
        .RST(rst), .I(e_init[73]), .Q(\u_a23_mem/e_mem[9][1] ) );
  DFF \u_a23_mem/e_mem_reg[9][2]  ( .D(\u_a23_mem/e_mem[9][2] ), .CLK(clk), 
        .RST(rst), .I(e_init[74]), .Q(\u_a23_mem/e_mem[9][2] ) );
  DFF \u_a23_mem/e_mem_reg[9][3]  ( .D(\u_a23_mem/e_mem[9][3] ), .CLK(clk), 
        .RST(rst), .I(e_init[75]), .Q(\u_a23_mem/e_mem[9][3] ) );
  DFF \u_a23_mem/e_mem_reg[9][4]  ( .D(\u_a23_mem/e_mem[9][4] ), .CLK(clk), 
        .RST(rst), .I(e_init[76]), .Q(\u_a23_mem/e_mem[9][4] ) );
  DFF \u_a23_mem/e_mem_reg[9][5]  ( .D(\u_a23_mem/e_mem[9][5] ), .CLK(clk), 
        .RST(rst), .I(e_init[77]), .Q(\u_a23_mem/e_mem[9][5] ) );
  DFF \u_a23_mem/e_mem_reg[9][6]  ( .D(\u_a23_mem/e_mem[9][6] ), .CLK(clk), 
        .RST(rst), .I(e_init[78]), .Q(\u_a23_mem/e_mem[9][6] ) );
  DFF \u_a23_mem/e_mem_reg[9][7]  ( .D(\u_a23_mem/e_mem[9][7] ), .CLK(clk), 
        .RST(rst), .I(e_init[79]), .Q(\u_a23_mem/e_mem[9][7] ) );
  DFF \u_a23_mem/e_mem_reg[10][0]  ( .D(\u_a23_mem/e_mem[10][0] ), .CLK(clk), 
        .RST(rst), .I(e_init[80]), .Q(\u_a23_mem/e_mem[10][0] ) );
  DFF \u_a23_mem/e_mem_reg[10][1]  ( .D(\u_a23_mem/e_mem[10][1] ), .CLK(clk), 
        .RST(rst), .I(e_init[81]), .Q(\u_a23_mem/e_mem[10][1] ) );
  DFF \u_a23_mem/e_mem_reg[10][2]  ( .D(\u_a23_mem/e_mem[10][2] ), .CLK(clk), 
        .RST(rst), .I(e_init[82]), .Q(\u_a23_mem/e_mem[10][2] ) );
  DFF \u_a23_mem/e_mem_reg[10][3]  ( .D(\u_a23_mem/e_mem[10][3] ), .CLK(clk), 
        .RST(rst), .I(e_init[83]), .Q(\u_a23_mem/e_mem[10][3] ) );
  DFF \u_a23_mem/e_mem_reg[10][4]  ( .D(\u_a23_mem/e_mem[10][4] ), .CLK(clk), 
        .RST(rst), .I(e_init[84]), .Q(\u_a23_mem/e_mem[10][4] ) );
  DFF \u_a23_mem/e_mem_reg[10][5]  ( .D(\u_a23_mem/e_mem[10][5] ), .CLK(clk), 
        .RST(rst), .I(e_init[85]), .Q(\u_a23_mem/e_mem[10][5] ) );
  DFF \u_a23_mem/e_mem_reg[10][6]  ( .D(\u_a23_mem/e_mem[10][6] ), .CLK(clk), 
        .RST(rst), .I(e_init[86]), .Q(\u_a23_mem/e_mem[10][6] ) );
  DFF \u_a23_mem/e_mem_reg[10][7]  ( .D(\u_a23_mem/e_mem[10][7] ), .CLK(clk), 
        .RST(rst), .I(e_init[87]), .Q(\u_a23_mem/e_mem[10][7] ) );
  DFF \u_a23_mem/e_mem_reg[11][0]  ( .D(\u_a23_mem/e_mem[11][0] ), .CLK(clk), 
        .RST(rst), .I(e_init[88]), .Q(\u_a23_mem/e_mem[11][0] ) );
  DFF \u_a23_mem/e_mem_reg[11][1]  ( .D(\u_a23_mem/e_mem[11][1] ), .CLK(clk), 
        .RST(rst), .I(e_init[89]), .Q(\u_a23_mem/e_mem[11][1] ) );
  DFF \u_a23_mem/e_mem_reg[11][2]  ( .D(\u_a23_mem/e_mem[11][2] ), .CLK(clk), 
        .RST(rst), .I(e_init[90]), .Q(\u_a23_mem/e_mem[11][2] ) );
  DFF \u_a23_mem/e_mem_reg[11][3]  ( .D(\u_a23_mem/e_mem[11][3] ), .CLK(clk), 
        .RST(rst), .I(e_init[91]), .Q(\u_a23_mem/e_mem[11][3] ) );
  DFF \u_a23_mem/e_mem_reg[11][4]  ( .D(\u_a23_mem/e_mem[11][4] ), .CLK(clk), 
        .RST(rst), .I(e_init[92]), .Q(\u_a23_mem/e_mem[11][4] ) );
  DFF \u_a23_mem/e_mem_reg[11][5]  ( .D(\u_a23_mem/e_mem[11][5] ), .CLK(clk), 
        .RST(rst), .I(e_init[93]), .Q(\u_a23_mem/e_mem[11][5] ) );
  DFF \u_a23_mem/e_mem_reg[11][6]  ( .D(\u_a23_mem/e_mem[11][6] ), .CLK(clk), 
        .RST(rst), .I(e_init[94]), .Q(\u_a23_mem/e_mem[11][6] ) );
  DFF \u_a23_mem/e_mem_reg[11][7]  ( .D(\u_a23_mem/e_mem[11][7] ), .CLK(clk), 
        .RST(rst), .I(e_init[95]), .Q(\u_a23_mem/e_mem[11][7] ) );
  DFF \u_a23_mem/e_mem_reg[12][0]  ( .D(\u_a23_mem/e_mem[12][0] ), .CLK(clk), 
        .RST(rst), .I(e_init[96]), .Q(\u_a23_mem/e_mem[12][0] ) );
  DFF \u_a23_mem/e_mem_reg[12][1]  ( .D(\u_a23_mem/e_mem[12][1] ), .CLK(clk), 
        .RST(rst), .I(e_init[97]), .Q(\u_a23_mem/e_mem[12][1] ) );
  DFF \u_a23_mem/e_mem_reg[12][2]  ( .D(\u_a23_mem/e_mem[12][2] ), .CLK(clk), 
        .RST(rst), .I(e_init[98]), .Q(\u_a23_mem/e_mem[12][2] ) );
  DFF \u_a23_mem/e_mem_reg[12][3]  ( .D(\u_a23_mem/e_mem[12][3] ), .CLK(clk), 
        .RST(rst), .I(e_init[99]), .Q(\u_a23_mem/e_mem[12][3] ) );
  DFF \u_a23_mem/e_mem_reg[12][4]  ( .D(\u_a23_mem/e_mem[12][4] ), .CLK(clk), 
        .RST(rst), .I(e_init[100]), .Q(\u_a23_mem/e_mem[12][4] ) );
  DFF \u_a23_mem/e_mem_reg[12][5]  ( .D(\u_a23_mem/e_mem[12][5] ), .CLK(clk), 
        .RST(rst), .I(e_init[101]), .Q(\u_a23_mem/e_mem[12][5] ) );
  DFF \u_a23_mem/e_mem_reg[12][6]  ( .D(\u_a23_mem/e_mem[12][6] ), .CLK(clk), 
        .RST(rst), .I(e_init[102]), .Q(\u_a23_mem/e_mem[12][6] ) );
  DFF \u_a23_mem/e_mem_reg[12][7]  ( .D(\u_a23_mem/e_mem[12][7] ), .CLK(clk), 
        .RST(rst), .I(e_init[103]), .Q(\u_a23_mem/e_mem[12][7] ) );
  DFF \u_a23_mem/e_mem_reg[13][0]  ( .D(\u_a23_mem/e_mem[13][0] ), .CLK(clk), 
        .RST(rst), .I(e_init[104]), .Q(\u_a23_mem/e_mem[13][0] ) );
  DFF \u_a23_mem/e_mem_reg[13][1]  ( .D(\u_a23_mem/e_mem[13][1] ), .CLK(clk), 
        .RST(rst), .I(e_init[105]), .Q(\u_a23_mem/e_mem[13][1] ) );
  DFF \u_a23_mem/e_mem_reg[13][2]  ( .D(\u_a23_mem/e_mem[13][2] ), .CLK(clk), 
        .RST(rst), .I(e_init[106]), .Q(\u_a23_mem/e_mem[13][2] ) );
  DFF \u_a23_mem/e_mem_reg[13][3]  ( .D(\u_a23_mem/e_mem[13][3] ), .CLK(clk), 
        .RST(rst), .I(e_init[107]), .Q(\u_a23_mem/e_mem[13][3] ) );
  DFF \u_a23_mem/e_mem_reg[13][4]  ( .D(\u_a23_mem/e_mem[13][4] ), .CLK(clk), 
        .RST(rst), .I(e_init[108]), .Q(\u_a23_mem/e_mem[13][4] ) );
  DFF \u_a23_mem/e_mem_reg[13][5]  ( .D(\u_a23_mem/e_mem[13][5] ), .CLK(clk), 
        .RST(rst), .I(e_init[109]), .Q(\u_a23_mem/e_mem[13][5] ) );
  DFF \u_a23_mem/e_mem_reg[13][6]  ( .D(\u_a23_mem/e_mem[13][6] ), .CLK(clk), 
        .RST(rst), .I(e_init[110]), .Q(\u_a23_mem/e_mem[13][6] ) );
  DFF \u_a23_mem/e_mem_reg[13][7]  ( .D(\u_a23_mem/e_mem[13][7] ), .CLK(clk), 
        .RST(rst), .I(e_init[111]), .Q(\u_a23_mem/e_mem[13][7] ) );
  DFF \u_a23_mem/e_mem_reg[14][0]  ( .D(\u_a23_mem/e_mem[14][0] ), .CLK(clk), 
        .RST(rst), .I(e_init[112]), .Q(\u_a23_mem/e_mem[14][0] ) );
  DFF \u_a23_mem/e_mem_reg[14][1]  ( .D(\u_a23_mem/e_mem[14][1] ), .CLK(clk), 
        .RST(rst), .I(e_init[113]), .Q(\u_a23_mem/e_mem[14][1] ) );
  DFF \u_a23_mem/e_mem_reg[14][2]  ( .D(\u_a23_mem/e_mem[14][2] ), .CLK(clk), 
        .RST(rst), .I(e_init[114]), .Q(\u_a23_mem/e_mem[14][2] ) );
  DFF \u_a23_mem/e_mem_reg[14][3]  ( .D(\u_a23_mem/e_mem[14][3] ), .CLK(clk), 
        .RST(rst), .I(e_init[115]), .Q(\u_a23_mem/e_mem[14][3] ) );
  DFF \u_a23_mem/e_mem_reg[14][4]  ( .D(\u_a23_mem/e_mem[14][4] ), .CLK(clk), 
        .RST(rst), .I(e_init[116]), .Q(\u_a23_mem/e_mem[14][4] ) );
  DFF \u_a23_mem/e_mem_reg[14][5]  ( .D(\u_a23_mem/e_mem[14][5] ), .CLK(clk), 
        .RST(rst), .I(e_init[117]), .Q(\u_a23_mem/e_mem[14][5] ) );
  DFF \u_a23_mem/e_mem_reg[14][6]  ( .D(\u_a23_mem/e_mem[14][6] ), .CLK(clk), 
        .RST(rst), .I(e_init[118]), .Q(\u_a23_mem/e_mem[14][6] ) );
  DFF \u_a23_mem/e_mem_reg[14][7]  ( .D(\u_a23_mem/e_mem[14][7] ), .CLK(clk), 
        .RST(rst), .I(e_init[119]), .Q(\u_a23_mem/e_mem[14][7] ) );
  DFF \u_a23_mem/e_mem_reg[15][0]  ( .D(\u_a23_mem/e_mem[15][0] ), .CLK(clk), 
        .RST(rst), .I(e_init[120]), .Q(\u_a23_mem/e_mem[15][0] ) );
  DFF \u_a23_mem/e_mem_reg[15][1]  ( .D(\u_a23_mem/e_mem[15][1] ), .CLK(clk), 
        .RST(rst), .I(e_init[121]), .Q(\u_a23_mem/e_mem[15][1] ) );
  DFF \u_a23_mem/e_mem_reg[15][2]  ( .D(\u_a23_mem/e_mem[15][2] ), .CLK(clk), 
        .RST(rst), .I(e_init[122]), .Q(\u_a23_mem/e_mem[15][2] ) );
  DFF \u_a23_mem/e_mem_reg[15][3]  ( .D(\u_a23_mem/e_mem[15][3] ), .CLK(clk), 
        .RST(rst), .I(e_init[123]), .Q(\u_a23_mem/e_mem[15][3] ) );
  DFF \u_a23_mem/e_mem_reg[15][4]  ( .D(\u_a23_mem/e_mem[15][4] ), .CLK(clk), 
        .RST(rst), .I(e_init[124]), .Q(\u_a23_mem/e_mem[15][4] ) );
  DFF \u_a23_mem/e_mem_reg[15][5]  ( .D(\u_a23_mem/e_mem[15][5] ), .CLK(clk), 
        .RST(rst), .I(e_init[125]), .Q(\u_a23_mem/e_mem[15][5] ) );
  DFF \u_a23_mem/e_mem_reg[15][6]  ( .D(\u_a23_mem/e_mem[15][6] ), .CLK(clk), 
        .RST(rst), .I(e_init[126]), .Q(\u_a23_mem/e_mem[15][6] ) );
  DFF \u_a23_mem/e_mem_reg[15][7]  ( .D(\u_a23_mem/e_mem[15][7] ), .CLK(clk), 
        .RST(rst), .I(e_init[127]), .Q(\u_a23_mem/e_mem[15][7] ) );
  DFF \u_a23_mem/e_mem_reg[16][0]  ( .D(\u_a23_mem/e_mem[16][0] ), .CLK(clk), 
        .RST(rst), .I(e_init[128]), .Q(\u_a23_mem/e_mem[16][0] ) );
  DFF \u_a23_mem/e_mem_reg[16][1]  ( .D(\u_a23_mem/e_mem[16][1] ), .CLK(clk), 
        .RST(rst), .I(e_init[129]), .Q(\u_a23_mem/e_mem[16][1] ) );
  DFF \u_a23_mem/e_mem_reg[16][2]  ( .D(\u_a23_mem/e_mem[16][2] ), .CLK(clk), 
        .RST(rst), .I(e_init[130]), .Q(\u_a23_mem/e_mem[16][2] ) );
  DFF \u_a23_mem/e_mem_reg[16][3]  ( .D(\u_a23_mem/e_mem[16][3] ), .CLK(clk), 
        .RST(rst), .I(e_init[131]), .Q(\u_a23_mem/e_mem[16][3] ) );
  DFF \u_a23_mem/e_mem_reg[16][4]  ( .D(\u_a23_mem/e_mem[16][4] ), .CLK(clk), 
        .RST(rst), .I(e_init[132]), .Q(\u_a23_mem/e_mem[16][4] ) );
  DFF \u_a23_mem/e_mem_reg[16][5]  ( .D(\u_a23_mem/e_mem[16][5] ), .CLK(clk), 
        .RST(rst), .I(e_init[133]), .Q(\u_a23_mem/e_mem[16][5] ) );
  DFF \u_a23_mem/e_mem_reg[16][6]  ( .D(\u_a23_mem/e_mem[16][6] ), .CLK(clk), 
        .RST(rst), .I(e_init[134]), .Q(\u_a23_mem/e_mem[16][6] ) );
  DFF \u_a23_mem/e_mem_reg[16][7]  ( .D(\u_a23_mem/e_mem[16][7] ), .CLK(clk), 
        .RST(rst), .I(e_init[135]), .Q(\u_a23_mem/e_mem[16][7] ) );
  DFF \u_a23_mem/e_mem_reg[17][0]  ( .D(\u_a23_mem/e_mem[17][0] ), .CLK(clk), 
        .RST(rst), .I(e_init[136]), .Q(\u_a23_mem/e_mem[17][0] ) );
  DFF \u_a23_mem/e_mem_reg[17][1]  ( .D(\u_a23_mem/e_mem[17][1] ), .CLK(clk), 
        .RST(rst), .I(e_init[137]), .Q(\u_a23_mem/e_mem[17][1] ) );
  DFF \u_a23_mem/e_mem_reg[17][2]  ( .D(\u_a23_mem/e_mem[17][2] ), .CLK(clk), 
        .RST(rst), .I(e_init[138]), .Q(\u_a23_mem/e_mem[17][2] ) );
  DFF \u_a23_mem/e_mem_reg[17][3]  ( .D(\u_a23_mem/e_mem[17][3] ), .CLK(clk), 
        .RST(rst), .I(e_init[139]), .Q(\u_a23_mem/e_mem[17][3] ) );
  DFF \u_a23_mem/e_mem_reg[17][4]  ( .D(\u_a23_mem/e_mem[17][4] ), .CLK(clk), 
        .RST(rst), .I(e_init[140]), .Q(\u_a23_mem/e_mem[17][4] ) );
  DFF \u_a23_mem/e_mem_reg[17][5]  ( .D(\u_a23_mem/e_mem[17][5] ), .CLK(clk), 
        .RST(rst), .I(e_init[141]), .Q(\u_a23_mem/e_mem[17][5] ) );
  DFF \u_a23_mem/e_mem_reg[17][6]  ( .D(\u_a23_mem/e_mem[17][6] ), .CLK(clk), 
        .RST(rst), .I(e_init[142]), .Q(\u_a23_mem/e_mem[17][6] ) );
  DFF \u_a23_mem/e_mem_reg[17][7]  ( .D(\u_a23_mem/e_mem[17][7] ), .CLK(clk), 
        .RST(rst), .I(e_init[143]), .Q(\u_a23_mem/e_mem[17][7] ) );
  DFF \u_a23_mem/e_mem_reg[18][0]  ( .D(\u_a23_mem/e_mem[18][0] ), .CLK(clk), 
        .RST(rst), .I(e_init[144]), .Q(\u_a23_mem/e_mem[18][0] ) );
  DFF \u_a23_mem/e_mem_reg[18][1]  ( .D(\u_a23_mem/e_mem[18][1] ), .CLK(clk), 
        .RST(rst), .I(e_init[145]), .Q(\u_a23_mem/e_mem[18][1] ) );
  DFF \u_a23_mem/e_mem_reg[18][2]  ( .D(\u_a23_mem/e_mem[18][2] ), .CLK(clk), 
        .RST(rst), .I(e_init[146]), .Q(\u_a23_mem/e_mem[18][2] ) );
  DFF \u_a23_mem/e_mem_reg[18][3]  ( .D(\u_a23_mem/e_mem[18][3] ), .CLK(clk), 
        .RST(rst), .I(e_init[147]), .Q(\u_a23_mem/e_mem[18][3] ) );
  DFF \u_a23_mem/e_mem_reg[18][4]  ( .D(\u_a23_mem/e_mem[18][4] ), .CLK(clk), 
        .RST(rst), .I(e_init[148]), .Q(\u_a23_mem/e_mem[18][4] ) );
  DFF \u_a23_mem/e_mem_reg[18][5]  ( .D(\u_a23_mem/e_mem[18][5] ), .CLK(clk), 
        .RST(rst), .I(e_init[149]), .Q(\u_a23_mem/e_mem[18][5] ) );
  DFF \u_a23_mem/e_mem_reg[18][6]  ( .D(\u_a23_mem/e_mem[18][6] ), .CLK(clk), 
        .RST(rst), .I(e_init[150]), .Q(\u_a23_mem/e_mem[18][6] ) );
  DFF \u_a23_mem/e_mem_reg[18][7]  ( .D(\u_a23_mem/e_mem[18][7] ), .CLK(clk), 
        .RST(rst), .I(e_init[151]), .Q(\u_a23_mem/e_mem[18][7] ) );
  DFF \u_a23_mem/e_mem_reg[19][0]  ( .D(\u_a23_mem/e_mem[19][0] ), .CLK(clk), 
        .RST(rst), .I(e_init[152]), .Q(\u_a23_mem/e_mem[19][0] ) );
  DFF \u_a23_mem/e_mem_reg[19][1]  ( .D(\u_a23_mem/e_mem[19][1] ), .CLK(clk), 
        .RST(rst), .I(e_init[153]), .Q(\u_a23_mem/e_mem[19][1] ) );
  DFF \u_a23_mem/e_mem_reg[19][2]  ( .D(\u_a23_mem/e_mem[19][2] ), .CLK(clk), 
        .RST(rst), .I(e_init[154]), .Q(\u_a23_mem/e_mem[19][2] ) );
  DFF \u_a23_mem/e_mem_reg[19][3]  ( .D(\u_a23_mem/e_mem[19][3] ), .CLK(clk), 
        .RST(rst), .I(e_init[155]), .Q(\u_a23_mem/e_mem[19][3] ) );
  DFF \u_a23_mem/e_mem_reg[19][4]  ( .D(\u_a23_mem/e_mem[19][4] ), .CLK(clk), 
        .RST(rst), .I(e_init[156]), .Q(\u_a23_mem/e_mem[19][4] ) );
  DFF \u_a23_mem/e_mem_reg[19][5]  ( .D(\u_a23_mem/e_mem[19][5] ), .CLK(clk), 
        .RST(rst), .I(e_init[157]), .Q(\u_a23_mem/e_mem[19][5] ) );
  DFF \u_a23_mem/e_mem_reg[19][6]  ( .D(\u_a23_mem/e_mem[19][6] ), .CLK(clk), 
        .RST(rst), .I(e_init[158]), .Q(\u_a23_mem/e_mem[19][6] ) );
  DFF \u_a23_mem/e_mem_reg[19][7]  ( .D(\u_a23_mem/e_mem[19][7] ), .CLK(clk), 
        .RST(rst), .I(e_init[159]), .Q(\u_a23_mem/e_mem[19][7] ) );
  DFF \u_a23_mem/e_mem_reg[20][0]  ( .D(\u_a23_mem/e_mem[20][0] ), .CLK(clk), 
        .RST(rst), .I(e_init[160]), .Q(\u_a23_mem/e_mem[20][0] ) );
  DFF \u_a23_mem/e_mem_reg[20][1]  ( .D(\u_a23_mem/e_mem[20][1] ), .CLK(clk), 
        .RST(rst), .I(e_init[161]), .Q(\u_a23_mem/e_mem[20][1] ) );
  DFF \u_a23_mem/e_mem_reg[20][2]  ( .D(\u_a23_mem/e_mem[20][2] ), .CLK(clk), 
        .RST(rst), .I(e_init[162]), .Q(\u_a23_mem/e_mem[20][2] ) );
  DFF \u_a23_mem/e_mem_reg[20][3]  ( .D(\u_a23_mem/e_mem[20][3] ), .CLK(clk), 
        .RST(rst), .I(e_init[163]), .Q(\u_a23_mem/e_mem[20][3] ) );
  DFF \u_a23_mem/e_mem_reg[20][4]  ( .D(\u_a23_mem/e_mem[20][4] ), .CLK(clk), 
        .RST(rst), .I(e_init[164]), .Q(\u_a23_mem/e_mem[20][4] ) );
  DFF \u_a23_mem/e_mem_reg[20][5]  ( .D(\u_a23_mem/e_mem[20][5] ), .CLK(clk), 
        .RST(rst), .I(e_init[165]), .Q(\u_a23_mem/e_mem[20][5] ) );
  DFF \u_a23_mem/e_mem_reg[20][6]  ( .D(\u_a23_mem/e_mem[20][6] ), .CLK(clk), 
        .RST(rst), .I(e_init[166]), .Q(\u_a23_mem/e_mem[20][6] ) );
  DFF \u_a23_mem/e_mem_reg[20][7]  ( .D(\u_a23_mem/e_mem[20][7] ), .CLK(clk), 
        .RST(rst), .I(e_init[167]), .Q(\u_a23_mem/e_mem[20][7] ) );
  DFF \u_a23_mem/e_mem_reg[21][0]  ( .D(\u_a23_mem/e_mem[21][0] ), .CLK(clk), 
        .RST(rst), .I(e_init[168]), .Q(\u_a23_mem/e_mem[21][0] ) );
  DFF \u_a23_mem/e_mem_reg[21][1]  ( .D(\u_a23_mem/e_mem[21][1] ), .CLK(clk), 
        .RST(rst), .I(e_init[169]), .Q(\u_a23_mem/e_mem[21][1] ) );
  DFF \u_a23_mem/e_mem_reg[21][2]  ( .D(\u_a23_mem/e_mem[21][2] ), .CLK(clk), 
        .RST(rst), .I(e_init[170]), .Q(\u_a23_mem/e_mem[21][2] ) );
  DFF \u_a23_mem/e_mem_reg[21][3]  ( .D(\u_a23_mem/e_mem[21][3] ), .CLK(clk), 
        .RST(rst), .I(e_init[171]), .Q(\u_a23_mem/e_mem[21][3] ) );
  DFF \u_a23_mem/e_mem_reg[21][4]  ( .D(\u_a23_mem/e_mem[21][4] ), .CLK(clk), 
        .RST(rst), .I(e_init[172]), .Q(\u_a23_mem/e_mem[21][4] ) );
  DFF \u_a23_mem/e_mem_reg[21][5]  ( .D(\u_a23_mem/e_mem[21][5] ), .CLK(clk), 
        .RST(rst), .I(e_init[173]), .Q(\u_a23_mem/e_mem[21][5] ) );
  DFF \u_a23_mem/e_mem_reg[21][6]  ( .D(\u_a23_mem/e_mem[21][6] ), .CLK(clk), 
        .RST(rst), .I(e_init[174]), .Q(\u_a23_mem/e_mem[21][6] ) );
  DFF \u_a23_mem/e_mem_reg[21][7]  ( .D(\u_a23_mem/e_mem[21][7] ), .CLK(clk), 
        .RST(rst), .I(e_init[175]), .Q(\u_a23_mem/e_mem[21][7] ) );
  DFF \u_a23_mem/e_mem_reg[22][0]  ( .D(\u_a23_mem/e_mem[22][0] ), .CLK(clk), 
        .RST(rst), .I(e_init[176]), .Q(\u_a23_mem/e_mem[22][0] ) );
  DFF \u_a23_mem/e_mem_reg[22][1]  ( .D(\u_a23_mem/e_mem[22][1] ), .CLK(clk), 
        .RST(rst), .I(e_init[177]), .Q(\u_a23_mem/e_mem[22][1] ) );
  DFF \u_a23_mem/e_mem_reg[22][2]  ( .D(\u_a23_mem/e_mem[22][2] ), .CLK(clk), 
        .RST(rst), .I(e_init[178]), .Q(\u_a23_mem/e_mem[22][2] ) );
  DFF \u_a23_mem/e_mem_reg[22][3]  ( .D(\u_a23_mem/e_mem[22][3] ), .CLK(clk), 
        .RST(rst), .I(e_init[179]), .Q(\u_a23_mem/e_mem[22][3] ) );
  DFF \u_a23_mem/e_mem_reg[22][4]  ( .D(\u_a23_mem/e_mem[22][4] ), .CLK(clk), 
        .RST(rst), .I(e_init[180]), .Q(\u_a23_mem/e_mem[22][4] ) );
  DFF \u_a23_mem/e_mem_reg[22][5]  ( .D(\u_a23_mem/e_mem[22][5] ), .CLK(clk), 
        .RST(rst), .I(e_init[181]), .Q(\u_a23_mem/e_mem[22][5] ) );
  DFF \u_a23_mem/e_mem_reg[22][6]  ( .D(\u_a23_mem/e_mem[22][6] ), .CLK(clk), 
        .RST(rst), .I(e_init[182]), .Q(\u_a23_mem/e_mem[22][6] ) );
  DFF \u_a23_mem/e_mem_reg[22][7]  ( .D(\u_a23_mem/e_mem[22][7] ), .CLK(clk), 
        .RST(rst), .I(e_init[183]), .Q(\u_a23_mem/e_mem[22][7] ) );
  DFF \u_a23_mem/e_mem_reg[23][0]  ( .D(\u_a23_mem/e_mem[23][0] ), .CLK(clk), 
        .RST(rst), .I(e_init[184]), .Q(\u_a23_mem/e_mem[23][0] ) );
  DFF \u_a23_mem/e_mem_reg[23][1]  ( .D(\u_a23_mem/e_mem[23][1] ), .CLK(clk), 
        .RST(rst), .I(e_init[185]), .Q(\u_a23_mem/e_mem[23][1] ) );
  DFF \u_a23_mem/e_mem_reg[23][2]  ( .D(\u_a23_mem/e_mem[23][2] ), .CLK(clk), 
        .RST(rst), .I(e_init[186]), .Q(\u_a23_mem/e_mem[23][2] ) );
  DFF \u_a23_mem/e_mem_reg[23][3]  ( .D(\u_a23_mem/e_mem[23][3] ), .CLK(clk), 
        .RST(rst), .I(e_init[187]), .Q(\u_a23_mem/e_mem[23][3] ) );
  DFF \u_a23_mem/e_mem_reg[23][4]  ( .D(\u_a23_mem/e_mem[23][4] ), .CLK(clk), 
        .RST(rst), .I(e_init[188]), .Q(\u_a23_mem/e_mem[23][4] ) );
  DFF \u_a23_mem/e_mem_reg[23][5]  ( .D(\u_a23_mem/e_mem[23][5] ), .CLK(clk), 
        .RST(rst), .I(e_init[189]), .Q(\u_a23_mem/e_mem[23][5] ) );
  DFF \u_a23_mem/e_mem_reg[23][6]  ( .D(\u_a23_mem/e_mem[23][6] ), .CLK(clk), 
        .RST(rst), .I(e_init[190]), .Q(\u_a23_mem/e_mem[23][6] ) );
  DFF \u_a23_mem/e_mem_reg[23][7]  ( .D(\u_a23_mem/e_mem[23][7] ), .CLK(clk), 
        .RST(rst), .I(e_init[191]), .Q(\u_a23_mem/e_mem[23][7] ) );
  DFF \u_a23_mem/e_mem_reg[24][0]  ( .D(\u_a23_mem/e_mem[24][0] ), .CLK(clk), 
        .RST(rst), .I(e_init[192]), .Q(\u_a23_mem/e_mem[24][0] ) );
  DFF \u_a23_mem/e_mem_reg[24][1]  ( .D(\u_a23_mem/e_mem[24][1] ), .CLK(clk), 
        .RST(rst), .I(e_init[193]), .Q(\u_a23_mem/e_mem[24][1] ) );
  DFF \u_a23_mem/e_mem_reg[24][2]  ( .D(\u_a23_mem/e_mem[24][2] ), .CLK(clk), 
        .RST(rst), .I(e_init[194]), .Q(\u_a23_mem/e_mem[24][2] ) );
  DFF \u_a23_mem/e_mem_reg[24][3]  ( .D(\u_a23_mem/e_mem[24][3] ), .CLK(clk), 
        .RST(rst), .I(e_init[195]), .Q(\u_a23_mem/e_mem[24][3] ) );
  DFF \u_a23_mem/e_mem_reg[24][4]  ( .D(\u_a23_mem/e_mem[24][4] ), .CLK(clk), 
        .RST(rst), .I(e_init[196]), .Q(\u_a23_mem/e_mem[24][4] ) );
  DFF \u_a23_mem/e_mem_reg[24][5]  ( .D(\u_a23_mem/e_mem[24][5] ), .CLK(clk), 
        .RST(rst), .I(e_init[197]), .Q(\u_a23_mem/e_mem[24][5] ) );
  DFF \u_a23_mem/e_mem_reg[24][6]  ( .D(\u_a23_mem/e_mem[24][6] ), .CLK(clk), 
        .RST(rst), .I(e_init[198]), .Q(\u_a23_mem/e_mem[24][6] ) );
  DFF \u_a23_mem/e_mem_reg[24][7]  ( .D(\u_a23_mem/e_mem[24][7] ), .CLK(clk), 
        .RST(rst), .I(e_init[199]), .Q(\u_a23_mem/e_mem[24][7] ) );
  DFF \u_a23_mem/e_mem_reg[25][0]  ( .D(\u_a23_mem/e_mem[25][0] ), .CLK(clk), 
        .RST(rst), .I(e_init[200]), .Q(\u_a23_mem/e_mem[25][0] ) );
  DFF \u_a23_mem/e_mem_reg[25][1]  ( .D(\u_a23_mem/e_mem[25][1] ), .CLK(clk), 
        .RST(rst), .I(e_init[201]), .Q(\u_a23_mem/e_mem[25][1] ) );
  DFF \u_a23_mem/e_mem_reg[25][2]  ( .D(\u_a23_mem/e_mem[25][2] ), .CLK(clk), 
        .RST(rst), .I(e_init[202]), .Q(\u_a23_mem/e_mem[25][2] ) );
  DFF \u_a23_mem/e_mem_reg[25][3]  ( .D(\u_a23_mem/e_mem[25][3] ), .CLK(clk), 
        .RST(rst), .I(e_init[203]), .Q(\u_a23_mem/e_mem[25][3] ) );
  DFF \u_a23_mem/e_mem_reg[25][4]  ( .D(\u_a23_mem/e_mem[25][4] ), .CLK(clk), 
        .RST(rst), .I(e_init[204]), .Q(\u_a23_mem/e_mem[25][4] ) );
  DFF \u_a23_mem/e_mem_reg[25][5]  ( .D(\u_a23_mem/e_mem[25][5] ), .CLK(clk), 
        .RST(rst), .I(e_init[205]), .Q(\u_a23_mem/e_mem[25][5] ) );
  DFF \u_a23_mem/e_mem_reg[25][6]  ( .D(\u_a23_mem/e_mem[25][6] ), .CLK(clk), 
        .RST(rst), .I(e_init[206]), .Q(\u_a23_mem/e_mem[25][6] ) );
  DFF \u_a23_mem/e_mem_reg[25][7]  ( .D(\u_a23_mem/e_mem[25][7] ), .CLK(clk), 
        .RST(rst), .I(e_init[207]), .Q(\u_a23_mem/e_mem[25][7] ) );
  DFF \u_a23_mem/e_mem_reg[26][0]  ( .D(\u_a23_mem/e_mem[26][0] ), .CLK(clk), 
        .RST(rst), .I(e_init[208]), .Q(\u_a23_mem/e_mem[26][0] ) );
  DFF \u_a23_mem/e_mem_reg[26][1]  ( .D(\u_a23_mem/e_mem[26][1] ), .CLK(clk), 
        .RST(rst), .I(e_init[209]), .Q(\u_a23_mem/e_mem[26][1] ) );
  DFF \u_a23_mem/e_mem_reg[26][2]  ( .D(\u_a23_mem/e_mem[26][2] ), .CLK(clk), 
        .RST(rst), .I(e_init[210]), .Q(\u_a23_mem/e_mem[26][2] ) );
  DFF \u_a23_mem/e_mem_reg[26][3]  ( .D(\u_a23_mem/e_mem[26][3] ), .CLK(clk), 
        .RST(rst), .I(e_init[211]), .Q(\u_a23_mem/e_mem[26][3] ) );
  DFF \u_a23_mem/e_mem_reg[26][4]  ( .D(\u_a23_mem/e_mem[26][4] ), .CLK(clk), 
        .RST(rst), .I(e_init[212]), .Q(\u_a23_mem/e_mem[26][4] ) );
  DFF \u_a23_mem/e_mem_reg[26][5]  ( .D(\u_a23_mem/e_mem[26][5] ), .CLK(clk), 
        .RST(rst), .I(e_init[213]), .Q(\u_a23_mem/e_mem[26][5] ) );
  DFF \u_a23_mem/e_mem_reg[26][6]  ( .D(\u_a23_mem/e_mem[26][6] ), .CLK(clk), 
        .RST(rst), .I(e_init[214]), .Q(\u_a23_mem/e_mem[26][6] ) );
  DFF \u_a23_mem/e_mem_reg[26][7]  ( .D(\u_a23_mem/e_mem[26][7] ), .CLK(clk), 
        .RST(rst), .I(e_init[215]), .Q(\u_a23_mem/e_mem[26][7] ) );
  DFF \u_a23_mem/e_mem_reg[27][0]  ( .D(\u_a23_mem/e_mem[27][0] ), .CLK(clk), 
        .RST(rst), .I(e_init[216]), .Q(\u_a23_mem/e_mem[27][0] ) );
  DFF \u_a23_mem/e_mem_reg[27][1]  ( .D(\u_a23_mem/e_mem[27][1] ), .CLK(clk), 
        .RST(rst), .I(e_init[217]), .Q(\u_a23_mem/e_mem[27][1] ) );
  DFF \u_a23_mem/e_mem_reg[27][2]  ( .D(\u_a23_mem/e_mem[27][2] ), .CLK(clk), 
        .RST(rst), .I(e_init[218]), .Q(\u_a23_mem/e_mem[27][2] ) );
  DFF \u_a23_mem/e_mem_reg[27][3]  ( .D(\u_a23_mem/e_mem[27][3] ), .CLK(clk), 
        .RST(rst), .I(e_init[219]), .Q(\u_a23_mem/e_mem[27][3] ) );
  DFF \u_a23_mem/e_mem_reg[27][4]  ( .D(\u_a23_mem/e_mem[27][4] ), .CLK(clk), 
        .RST(rst), .I(e_init[220]), .Q(\u_a23_mem/e_mem[27][4] ) );
  DFF \u_a23_mem/e_mem_reg[27][5]  ( .D(\u_a23_mem/e_mem[27][5] ), .CLK(clk), 
        .RST(rst), .I(e_init[221]), .Q(\u_a23_mem/e_mem[27][5] ) );
  DFF \u_a23_mem/e_mem_reg[27][6]  ( .D(\u_a23_mem/e_mem[27][6] ), .CLK(clk), 
        .RST(rst), .I(e_init[222]), .Q(\u_a23_mem/e_mem[27][6] ) );
  DFF \u_a23_mem/e_mem_reg[27][7]  ( .D(\u_a23_mem/e_mem[27][7] ), .CLK(clk), 
        .RST(rst), .I(e_init[223]), .Q(\u_a23_mem/e_mem[27][7] ) );
  DFF \u_a23_mem/e_mem_reg[28][0]  ( .D(\u_a23_mem/e_mem[28][0] ), .CLK(clk), 
        .RST(rst), .I(e_init[224]), .Q(\u_a23_mem/e_mem[28][0] ) );
  DFF \u_a23_mem/e_mem_reg[28][1]  ( .D(\u_a23_mem/e_mem[28][1] ), .CLK(clk), 
        .RST(rst), .I(e_init[225]), .Q(\u_a23_mem/e_mem[28][1] ) );
  DFF \u_a23_mem/e_mem_reg[28][2]  ( .D(\u_a23_mem/e_mem[28][2] ), .CLK(clk), 
        .RST(rst), .I(e_init[226]), .Q(\u_a23_mem/e_mem[28][2] ) );
  DFF \u_a23_mem/e_mem_reg[28][3]  ( .D(\u_a23_mem/e_mem[28][3] ), .CLK(clk), 
        .RST(rst), .I(e_init[227]), .Q(\u_a23_mem/e_mem[28][3] ) );
  DFF \u_a23_mem/e_mem_reg[28][4]  ( .D(\u_a23_mem/e_mem[28][4] ), .CLK(clk), 
        .RST(rst), .I(e_init[228]), .Q(\u_a23_mem/e_mem[28][4] ) );
  DFF \u_a23_mem/e_mem_reg[28][5]  ( .D(\u_a23_mem/e_mem[28][5] ), .CLK(clk), 
        .RST(rst), .I(e_init[229]), .Q(\u_a23_mem/e_mem[28][5] ) );
  DFF \u_a23_mem/e_mem_reg[28][6]  ( .D(\u_a23_mem/e_mem[28][6] ), .CLK(clk), 
        .RST(rst), .I(e_init[230]), .Q(\u_a23_mem/e_mem[28][6] ) );
  DFF \u_a23_mem/e_mem_reg[28][7]  ( .D(\u_a23_mem/e_mem[28][7] ), .CLK(clk), 
        .RST(rst), .I(e_init[231]), .Q(\u_a23_mem/e_mem[28][7] ) );
  DFF \u_a23_mem/e_mem_reg[29][0]  ( .D(\u_a23_mem/e_mem[29][0] ), .CLK(clk), 
        .RST(rst), .I(e_init[232]), .Q(\u_a23_mem/e_mem[29][0] ) );
  DFF \u_a23_mem/e_mem_reg[29][1]  ( .D(\u_a23_mem/e_mem[29][1] ), .CLK(clk), 
        .RST(rst), .I(e_init[233]), .Q(\u_a23_mem/e_mem[29][1] ) );
  DFF \u_a23_mem/e_mem_reg[29][2]  ( .D(\u_a23_mem/e_mem[29][2] ), .CLK(clk), 
        .RST(rst), .I(e_init[234]), .Q(\u_a23_mem/e_mem[29][2] ) );
  DFF \u_a23_mem/e_mem_reg[29][3]  ( .D(\u_a23_mem/e_mem[29][3] ), .CLK(clk), 
        .RST(rst), .I(e_init[235]), .Q(\u_a23_mem/e_mem[29][3] ) );
  DFF \u_a23_mem/e_mem_reg[29][4]  ( .D(\u_a23_mem/e_mem[29][4] ), .CLK(clk), 
        .RST(rst), .I(e_init[236]), .Q(\u_a23_mem/e_mem[29][4] ) );
  DFF \u_a23_mem/e_mem_reg[29][5]  ( .D(\u_a23_mem/e_mem[29][5] ), .CLK(clk), 
        .RST(rst), .I(e_init[237]), .Q(\u_a23_mem/e_mem[29][5] ) );
  DFF \u_a23_mem/e_mem_reg[29][6]  ( .D(\u_a23_mem/e_mem[29][6] ), .CLK(clk), 
        .RST(rst), .I(e_init[238]), .Q(\u_a23_mem/e_mem[29][6] ) );
  DFF \u_a23_mem/e_mem_reg[29][7]  ( .D(\u_a23_mem/e_mem[29][7] ), .CLK(clk), 
        .RST(rst), .I(e_init[239]), .Q(\u_a23_mem/e_mem[29][7] ) );
  DFF \u_a23_mem/e_mem_reg[30][0]  ( .D(\u_a23_mem/e_mem[30][0] ), .CLK(clk), 
        .RST(rst), .I(e_init[240]), .Q(\u_a23_mem/e_mem[30][0] ) );
  DFF \u_a23_mem/e_mem_reg[30][1]  ( .D(\u_a23_mem/e_mem[30][1] ), .CLK(clk), 
        .RST(rst), .I(e_init[241]), .Q(\u_a23_mem/e_mem[30][1] ) );
  DFF \u_a23_mem/e_mem_reg[30][2]  ( .D(\u_a23_mem/e_mem[30][2] ), .CLK(clk), 
        .RST(rst), .I(e_init[242]), .Q(\u_a23_mem/e_mem[30][2] ) );
  DFF \u_a23_mem/e_mem_reg[30][3]  ( .D(\u_a23_mem/e_mem[30][3] ), .CLK(clk), 
        .RST(rst), .I(e_init[243]), .Q(\u_a23_mem/e_mem[30][3] ) );
  DFF \u_a23_mem/e_mem_reg[30][4]  ( .D(\u_a23_mem/e_mem[30][4] ), .CLK(clk), 
        .RST(rst), .I(e_init[244]), .Q(\u_a23_mem/e_mem[30][4] ) );
  DFF \u_a23_mem/e_mem_reg[30][5]  ( .D(\u_a23_mem/e_mem[30][5] ), .CLK(clk), 
        .RST(rst), .I(e_init[245]), .Q(\u_a23_mem/e_mem[30][5] ) );
  DFF \u_a23_mem/e_mem_reg[30][6]  ( .D(\u_a23_mem/e_mem[30][6] ), .CLK(clk), 
        .RST(rst), .I(e_init[246]), .Q(\u_a23_mem/e_mem[30][6] ) );
  DFF \u_a23_mem/e_mem_reg[30][7]  ( .D(\u_a23_mem/e_mem[30][7] ), .CLK(clk), 
        .RST(rst), .I(e_init[247]), .Q(\u_a23_mem/e_mem[30][7] ) );
  DFF \u_a23_mem/e_mem_reg[31][0]  ( .D(\u_a23_mem/e_mem[31][0] ), .CLK(clk), 
        .RST(rst), .I(e_init[248]), .Q(\u_a23_mem/e_mem[31][0] ) );
  DFF \u_a23_mem/e_mem_reg[31][1]  ( .D(\u_a23_mem/e_mem[31][1] ), .CLK(clk), 
        .RST(rst), .I(e_init[249]), .Q(\u_a23_mem/e_mem[31][1] ) );
  DFF \u_a23_mem/e_mem_reg[31][2]  ( .D(\u_a23_mem/e_mem[31][2] ), .CLK(clk), 
        .RST(rst), .I(e_init[250]), .Q(\u_a23_mem/e_mem[31][2] ) );
  DFF \u_a23_mem/e_mem_reg[31][3]  ( .D(\u_a23_mem/e_mem[31][3] ), .CLK(clk), 
        .RST(rst), .I(e_init[251]), .Q(\u_a23_mem/e_mem[31][3] ) );
  DFF \u_a23_mem/e_mem_reg[31][4]  ( .D(\u_a23_mem/e_mem[31][4] ), .CLK(clk), 
        .RST(rst), .I(e_init[252]), .Q(\u_a23_mem/e_mem[31][4] ) );
  DFF \u_a23_mem/e_mem_reg[31][5]  ( .D(\u_a23_mem/e_mem[31][5] ), .CLK(clk), 
        .RST(rst), .I(e_init[253]), .Q(\u_a23_mem/e_mem[31][5] ) );
  DFF \u_a23_mem/e_mem_reg[31][6]  ( .D(\u_a23_mem/e_mem[31][6] ), .CLK(clk), 
        .RST(rst), .I(e_init[254]), .Q(\u_a23_mem/e_mem[31][6] ) );
  DFF \u_a23_mem/e_mem_reg[31][7]  ( .D(\u_a23_mem/e_mem[31][7] ), .CLK(clk), 
        .RST(rst), .I(e_init[255]), .Q(\u_a23_mem/e_mem[31][7] ) );
  DFF \u_a23_mem/p_mem_reg[0][0]  ( .D(\u_a23_mem/n18380 ), .CLK(clk), .RST(
        rst), .I(p_init[0]), .Q(\u_a23_mem/p_mem[0][0] ) );
  DFF \u_a23_mem/p_mem_reg[0][1]  ( .D(\u_a23_mem/n18379 ), .CLK(clk), .RST(
        rst), .I(p_init[1]), .Q(\u_a23_mem/p_mem[0][1] ) );
  DFF \u_a23_mem/p_mem_reg[0][2]  ( .D(\u_a23_mem/n18378 ), .CLK(clk), .RST(
        rst), .I(p_init[2]), .Q(\u_a23_mem/p_mem[0][2] ) );
  DFF \u_a23_mem/p_mem_reg[0][3]  ( .D(\u_a23_mem/n18377 ), .CLK(clk), .RST(
        rst), .I(p_init[3]), .Q(\u_a23_mem/p_mem[0][3] ) );
  DFF \u_a23_mem/p_mem_reg[0][4]  ( .D(\u_a23_mem/n18376 ), .CLK(clk), .RST(
        rst), .I(p_init[4]), .Q(\u_a23_mem/p_mem[0][4] ) );
  DFF \u_a23_mem/p_mem_reg[0][5]  ( .D(\u_a23_mem/n18375 ), .CLK(clk), .RST(
        rst), .I(p_init[5]), .Q(\u_a23_mem/p_mem[0][5] ) );
  DFF \u_a23_mem/p_mem_reg[0][6]  ( .D(\u_a23_mem/n18374 ), .CLK(clk), .RST(
        rst), .I(p_init[6]), .Q(\u_a23_mem/p_mem[0][6] ) );
  DFF \u_a23_mem/p_mem_reg[0][7]  ( .D(\u_a23_mem/n18373 ), .CLK(clk), .RST(
        rst), .I(p_init[7]), .Q(\u_a23_mem/p_mem[0][7] ) );
  DFF \u_a23_mem/p_mem_reg[1][0]  ( .D(\u_a23_mem/n18388 ), .CLK(clk), .RST(
        rst), .I(p_init[8]), .Q(\u_a23_mem/p_mem[1][0] ) );
  DFF \u_a23_mem/p_mem_reg[1][1]  ( .D(\u_a23_mem/n18387 ), .CLK(clk), .RST(
        rst), .I(p_init[9]), .Q(\u_a23_mem/p_mem[1][1] ) );
  DFF \u_a23_mem/p_mem_reg[1][2]  ( .D(\u_a23_mem/n18386 ), .CLK(clk), .RST(
        rst), .I(p_init[10]), .Q(\u_a23_mem/p_mem[1][2] ) );
  DFF \u_a23_mem/p_mem_reg[1][3]  ( .D(\u_a23_mem/n18385 ), .CLK(clk), .RST(
        rst), .I(p_init[11]), .Q(\u_a23_mem/p_mem[1][3] ) );
  DFF \u_a23_mem/p_mem_reg[1][4]  ( .D(\u_a23_mem/n18384 ), .CLK(clk), .RST(
        rst), .I(p_init[12]), .Q(\u_a23_mem/p_mem[1][4] ) );
  DFF \u_a23_mem/p_mem_reg[1][5]  ( .D(\u_a23_mem/n18383 ), .CLK(clk), .RST(
        rst), .I(p_init[13]), .Q(\u_a23_mem/p_mem[1][5] ) );
  DFF \u_a23_mem/p_mem_reg[1][6]  ( .D(\u_a23_mem/n18382 ), .CLK(clk), .RST(
        rst), .I(p_init[14]), .Q(\u_a23_mem/p_mem[1][6] ) );
  DFF \u_a23_mem/p_mem_reg[1][7]  ( .D(\u_a23_mem/n18381 ), .CLK(clk), .RST(
        rst), .I(p_init[15]), .Q(\u_a23_mem/p_mem[1][7] ) );
  DFF \u_a23_mem/p_mem_reg[2][0]  ( .D(\u_a23_mem/n18396 ), .CLK(clk), .RST(
        rst), .I(p_init[16]), .Q(\u_a23_mem/p_mem[2][0] ) );
  DFF \u_a23_mem/p_mem_reg[2][1]  ( .D(\u_a23_mem/n18395 ), .CLK(clk), .RST(
        rst), .I(p_init[17]), .Q(\u_a23_mem/p_mem[2][1] ) );
  DFF \u_a23_mem/p_mem_reg[2][2]  ( .D(\u_a23_mem/n18394 ), .CLK(clk), .RST(
        rst), .I(p_init[18]), .Q(\u_a23_mem/p_mem[2][2] ) );
  DFF \u_a23_mem/p_mem_reg[2][3]  ( .D(\u_a23_mem/n18393 ), .CLK(clk), .RST(
        rst), .I(p_init[19]), .Q(\u_a23_mem/p_mem[2][3] ) );
  DFF \u_a23_mem/p_mem_reg[2][4]  ( .D(\u_a23_mem/n18392 ), .CLK(clk), .RST(
        rst), .I(p_init[20]), .Q(\u_a23_mem/p_mem[2][4] ) );
  DFF \u_a23_mem/p_mem_reg[2][5]  ( .D(\u_a23_mem/n18391 ), .CLK(clk), .RST(
        rst), .I(p_init[21]), .Q(\u_a23_mem/p_mem[2][5] ) );
  DFF \u_a23_mem/p_mem_reg[2][6]  ( .D(\u_a23_mem/n18390 ), .CLK(clk), .RST(
        rst), .I(p_init[22]), .Q(\u_a23_mem/p_mem[2][6] ) );
  DFF \u_a23_mem/p_mem_reg[2][7]  ( .D(\u_a23_mem/n18389 ), .CLK(clk), .RST(
        rst), .I(p_init[23]), .Q(\u_a23_mem/p_mem[2][7] ) );
  DFF \u_a23_mem/p_mem_reg[3][0]  ( .D(\u_a23_mem/n19396 ), .CLK(clk), .RST(
        rst), .I(p_init[24]), .Q(\u_a23_mem/p_mem[3][0] ) );
  DFF \u_a23_mem/p_mem_reg[3][1]  ( .D(\u_a23_mem/n19395 ), .CLK(clk), .RST(
        rst), .I(p_init[25]), .Q(\u_a23_mem/p_mem[3][1] ) );
  DFF \u_a23_mem/p_mem_reg[3][2]  ( .D(\u_a23_mem/n19394 ), .CLK(clk), .RST(
        rst), .I(p_init[26]), .Q(\u_a23_mem/p_mem[3][2] ) );
  DFF \u_a23_mem/p_mem_reg[3][3]  ( .D(\u_a23_mem/n19393 ), .CLK(clk), .RST(
        rst), .I(p_init[27]), .Q(\u_a23_mem/p_mem[3][3] ) );
  DFF \u_a23_mem/p_mem_reg[3][4]  ( .D(\u_a23_mem/n19392 ), .CLK(clk), .RST(
        rst), .I(p_init[28]), .Q(\u_a23_mem/p_mem[3][4] ) );
  DFF \u_a23_mem/p_mem_reg[3][5]  ( .D(\u_a23_mem/n19391 ), .CLK(clk), .RST(
        rst), .I(p_init[29]), .Q(\u_a23_mem/p_mem[3][5] ) );
  DFF \u_a23_mem/p_mem_reg[3][6]  ( .D(\u_a23_mem/n19390 ), .CLK(clk), .RST(
        rst), .I(p_init[30]), .Q(\u_a23_mem/p_mem[3][6] ) );
  DFF \u_a23_mem/p_mem_reg[3][7]  ( .D(\u_a23_mem/n19389 ), .CLK(clk), .RST(
        rst), .I(p_init[31]), .Q(\u_a23_mem/p_mem[3][7] ) );
  DFF \u_a23_mem/p_mem_reg[4][0]  ( .D(\u_a23_mem/n19388 ), .CLK(clk), .RST(
        rst), .I(p_init[32]), .Q(\u_a23_mem/p_mem[4][0] ) );
  DFF \u_a23_mem/p_mem_reg[4][1]  ( .D(\u_a23_mem/n19387 ), .CLK(clk), .RST(
        rst), .I(p_init[33]), .Q(\u_a23_mem/p_mem[4][1] ) );
  DFF \u_a23_mem/p_mem_reg[4][2]  ( .D(\u_a23_mem/n19386 ), .CLK(clk), .RST(
        rst), .I(p_init[34]), .Q(\u_a23_mem/p_mem[4][2] ) );
  DFF \u_a23_mem/p_mem_reg[4][3]  ( .D(\u_a23_mem/n19385 ), .CLK(clk), .RST(
        rst), .I(p_init[35]), .Q(\u_a23_mem/p_mem[4][3] ) );
  DFF \u_a23_mem/p_mem_reg[4][4]  ( .D(\u_a23_mem/n19384 ), .CLK(clk), .RST(
        rst), .I(p_init[36]), .Q(\u_a23_mem/p_mem[4][4] ) );
  DFF \u_a23_mem/p_mem_reg[4][5]  ( .D(\u_a23_mem/n19383 ), .CLK(clk), .RST(
        rst), .I(p_init[37]), .Q(\u_a23_mem/p_mem[4][5] ) );
  DFF \u_a23_mem/p_mem_reg[4][6]  ( .D(\u_a23_mem/n19382 ), .CLK(clk), .RST(
        rst), .I(p_init[38]), .Q(\u_a23_mem/p_mem[4][6] ) );
  DFF \u_a23_mem/p_mem_reg[4][7]  ( .D(\u_a23_mem/n19381 ), .CLK(clk), .RST(
        rst), .I(p_init[39]), .Q(\u_a23_mem/p_mem[4][7] ) );
  DFF \u_a23_mem/p_mem_reg[5][0]  ( .D(\u_a23_mem/n19380 ), .CLK(clk), .RST(
        rst), .I(p_init[40]), .Q(\u_a23_mem/p_mem[5][0] ) );
  DFF \u_a23_mem/p_mem_reg[5][1]  ( .D(\u_a23_mem/n19379 ), .CLK(clk), .RST(
        rst), .I(p_init[41]), .Q(\u_a23_mem/p_mem[5][1] ) );
  DFF \u_a23_mem/p_mem_reg[5][2]  ( .D(\u_a23_mem/n19378 ), .CLK(clk), .RST(
        rst), .I(p_init[42]), .Q(\u_a23_mem/p_mem[5][2] ) );
  DFF \u_a23_mem/p_mem_reg[5][3]  ( .D(\u_a23_mem/n19377 ), .CLK(clk), .RST(
        rst), .I(p_init[43]), .Q(\u_a23_mem/p_mem[5][3] ) );
  DFF \u_a23_mem/p_mem_reg[5][4]  ( .D(\u_a23_mem/n19376 ), .CLK(clk), .RST(
        rst), .I(p_init[44]), .Q(\u_a23_mem/p_mem[5][4] ) );
  DFF \u_a23_mem/p_mem_reg[5][5]  ( .D(\u_a23_mem/n19375 ), .CLK(clk), .RST(
        rst), .I(p_init[45]), .Q(\u_a23_mem/p_mem[5][5] ) );
  DFF \u_a23_mem/p_mem_reg[5][6]  ( .D(\u_a23_mem/n19374 ), .CLK(clk), .RST(
        rst), .I(p_init[46]), .Q(\u_a23_mem/p_mem[5][6] ) );
  DFF \u_a23_mem/p_mem_reg[5][7]  ( .D(\u_a23_mem/n19373 ), .CLK(clk), .RST(
        rst), .I(p_init[47]), .Q(\u_a23_mem/p_mem[5][7] ) );
  DFF \u_a23_mem/p_mem_reg[6][0]  ( .D(\u_a23_mem/n19372 ), .CLK(clk), .RST(
        rst), .I(p_init[48]), .Q(\u_a23_mem/p_mem[6][0] ) );
  DFF \u_a23_mem/p_mem_reg[6][1]  ( .D(\u_a23_mem/n19371 ), .CLK(clk), .RST(
        rst), .I(p_init[49]), .Q(\u_a23_mem/p_mem[6][1] ) );
  DFF \u_a23_mem/p_mem_reg[6][2]  ( .D(\u_a23_mem/n19370 ), .CLK(clk), .RST(
        rst), .I(p_init[50]), .Q(\u_a23_mem/p_mem[6][2] ) );
  DFF \u_a23_mem/p_mem_reg[6][3]  ( .D(\u_a23_mem/n19369 ), .CLK(clk), .RST(
        rst), .I(p_init[51]), .Q(\u_a23_mem/p_mem[6][3] ) );
  DFF \u_a23_mem/p_mem_reg[6][4]  ( .D(\u_a23_mem/n19368 ), .CLK(clk), .RST(
        rst), .I(p_init[52]), .Q(\u_a23_mem/p_mem[6][4] ) );
  DFF \u_a23_mem/p_mem_reg[6][5]  ( .D(\u_a23_mem/n19367 ), .CLK(clk), .RST(
        rst), .I(p_init[53]), .Q(\u_a23_mem/p_mem[6][5] ) );
  DFF \u_a23_mem/p_mem_reg[6][6]  ( .D(\u_a23_mem/n19366 ), .CLK(clk), .RST(
        rst), .I(p_init[54]), .Q(\u_a23_mem/p_mem[6][6] ) );
  DFF \u_a23_mem/p_mem_reg[6][7]  ( .D(\u_a23_mem/n19365 ), .CLK(clk), .RST(
        rst), .I(p_init[55]), .Q(\u_a23_mem/p_mem[6][7] ) );
  DFF \u_a23_mem/p_mem_reg[7][0]  ( .D(\u_a23_mem/n19364 ), .CLK(clk), .RST(
        rst), .I(p_init[56]), .Q(\u_a23_mem/p_mem[7][0] ) );
  DFF \u_a23_mem/p_mem_reg[7][1]  ( .D(\u_a23_mem/n19363 ), .CLK(clk), .RST(
        rst), .I(p_init[57]), .Q(\u_a23_mem/p_mem[7][1] ) );
  DFF \u_a23_mem/p_mem_reg[7][2]  ( .D(\u_a23_mem/n19362 ), .CLK(clk), .RST(
        rst), .I(p_init[58]), .Q(\u_a23_mem/p_mem[7][2] ) );
  DFF \u_a23_mem/p_mem_reg[7][3]  ( .D(\u_a23_mem/n19361 ), .CLK(clk), .RST(
        rst), .I(p_init[59]), .Q(\u_a23_mem/p_mem[7][3] ) );
  DFF \u_a23_mem/p_mem_reg[7][4]  ( .D(\u_a23_mem/n19360 ), .CLK(clk), .RST(
        rst), .I(p_init[60]), .Q(\u_a23_mem/p_mem[7][4] ) );
  DFF \u_a23_mem/p_mem_reg[7][5]  ( .D(\u_a23_mem/n19359 ), .CLK(clk), .RST(
        rst), .I(p_init[61]), .Q(\u_a23_mem/p_mem[7][5] ) );
  DFF \u_a23_mem/p_mem_reg[7][6]  ( .D(\u_a23_mem/n19358 ), .CLK(clk), .RST(
        rst), .I(p_init[62]), .Q(\u_a23_mem/p_mem[7][6] ) );
  DFF \u_a23_mem/p_mem_reg[7][7]  ( .D(\u_a23_mem/n19357 ), .CLK(clk), .RST(
        rst), .I(p_init[63]), .Q(\u_a23_mem/p_mem[7][7] ) );
  DFF \u_a23_mem/p_mem_reg[8][0]  ( .D(\u_a23_mem/n19356 ), .CLK(clk), .RST(
        rst), .I(p_init[64]), .Q(\u_a23_mem/p_mem[8][0] ) );
  DFF \u_a23_mem/p_mem_reg[8][1]  ( .D(\u_a23_mem/n19355 ), .CLK(clk), .RST(
        rst), .I(p_init[65]), .Q(\u_a23_mem/p_mem[8][1] ) );
  DFF \u_a23_mem/p_mem_reg[8][2]  ( .D(\u_a23_mem/n19354 ), .CLK(clk), .RST(
        rst), .I(p_init[66]), .Q(\u_a23_mem/p_mem[8][2] ) );
  DFF \u_a23_mem/p_mem_reg[8][3]  ( .D(\u_a23_mem/n19353 ), .CLK(clk), .RST(
        rst), .I(p_init[67]), .Q(\u_a23_mem/p_mem[8][3] ) );
  DFF \u_a23_mem/p_mem_reg[8][4]  ( .D(\u_a23_mem/n19352 ), .CLK(clk), .RST(
        rst), .I(p_init[68]), .Q(\u_a23_mem/p_mem[8][4] ) );
  DFF \u_a23_mem/p_mem_reg[8][5]  ( .D(\u_a23_mem/n19351 ), .CLK(clk), .RST(
        rst), .I(p_init[69]), .Q(\u_a23_mem/p_mem[8][5] ) );
  DFF \u_a23_mem/p_mem_reg[8][6]  ( .D(\u_a23_mem/n19350 ), .CLK(clk), .RST(
        rst), .I(p_init[70]), .Q(\u_a23_mem/p_mem[8][6] ) );
  DFF \u_a23_mem/p_mem_reg[8][7]  ( .D(\u_a23_mem/n19349 ), .CLK(clk), .RST(
        rst), .I(p_init[71]), .Q(\u_a23_mem/p_mem[8][7] ) );
  DFF \u_a23_mem/p_mem_reg[9][0]  ( .D(\u_a23_mem/n19348 ), .CLK(clk), .RST(
        rst), .I(p_init[72]), .Q(\u_a23_mem/p_mem[9][0] ) );
  DFF \u_a23_mem/p_mem_reg[9][1]  ( .D(\u_a23_mem/n19347 ), .CLK(clk), .RST(
        rst), .I(p_init[73]), .Q(\u_a23_mem/p_mem[9][1] ) );
  DFF \u_a23_mem/p_mem_reg[9][2]  ( .D(\u_a23_mem/n19346 ), .CLK(clk), .RST(
        rst), .I(p_init[74]), .Q(\u_a23_mem/p_mem[9][2] ) );
  DFF \u_a23_mem/p_mem_reg[9][3]  ( .D(\u_a23_mem/n19345 ), .CLK(clk), .RST(
        rst), .I(p_init[75]), .Q(\u_a23_mem/p_mem[9][3] ) );
  DFF \u_a23_mem/p_mem_reg[9][4]  ( .D(\u_a23_mem/n19344 ), .CLK(clk), .RST(
        rst), .I(p_init[76]), .Q(\u_a23_mem/p_mem[9][4] ) );
  DFF \u_a23_mem/p_mem_reg[9][5]  ( .D(\u_a23_mem/n19343 ), .CLK(clk), .RST(
        rst), .I(p_init[77]), .Q(\u_a23_mem/p_mem[9][5] ) );
  DFF \u_a23_mem/p_mem_reg[9][6]  ( .D(\u_a23_mem/n19342 ), .CLK(clk), .RST(
        rst), .I(p_init[78]), .Q(\u_a23_mem/p_mem[9][6] ) );
  DFF \u_a23_mem/p_mem_reg[9][7]  ( .D(\u_a23_mem/n19341 ), .CLK(clk), .RST(
        rst), .I(p_init[79]), .Q(\u_a23_mem/p_mem[9][7] ) );
  DFF \u_a23_mem/p_mem_reg[10][0]  ( .D(\u_a23_mem/n19340 ), .CLK(clk), .RST(
        rst), .I(p_init[80]), .Q(\u_a23_mem/p_mem[10][0] ) );
  DFF \u_a23_mem/p_mem_reg[10][1]  ( .D(\u_a23_mem/n19339 ), .CLK(clk), .RST(
        rst), .I(p_init[81]), .Q(\u_a23_mem/p_mem[10][1] ) );
  DFF \u_a23_mem/p_mem_reg[10][2]  ( .D(\u_a23_mem/n19338 ), .CLK(clk), .RST(
        rst), .I(p_init[82]), .Q(\u_a23_mem/p_mem[10][2] ) );
  DFF \u_a23_mem/p_mem_reg[10][3]  ( .D(\u_a23_mem/n19337 ), .CLK(clk), .RST(
        rst), .I(p_init[83]), .Q(\u_a23_mem/p_mem[10][3] ) );
  DFF \u_a23_mem/p_mem_reg[10][4]  ( .D(\u_a23_mem/n19336 ), .CLK(clk), .RST(
        rst), .I(p_init[84]), .Q(\u_a23_mem/p_mem[10][4] ) );
  DFF \u_a23_mem/p_mem_reg[10][5]  ( .D(\u_a23_mem/n19335 ), .CLK(clk), .RST(
        rst), .I(p_init[85]), .Q(\u_a23_mem/p_mem[10][5] ) );
  DFF \u_a23_mem/p_mem_reg[10][6]  ( .D(\u_a23_mem/n19334 ), .CLK(clk), .RST(
        rst), .I(p_init[86]), .Q(\u_a23_mem/p_mem[10][6] ) );
  DFF \u_a23_mem/p_mem_reg[10][7]  ( .D(\u_a23_mem/n19333 ), .CLK(clk), .RST(
        rst), .I(p_init[87]), .Q(\u_a23_mem/p_mem[10][7] ) );
  DFF \u_a23_mem/p_mem_reg[11][0]  ( .D(\u_a23_mem/n19332 ), .CLK(clk), .RST(
        rst), .I(p_init[88]), .Q(\u_a23_mem/p_mem[11][0] ) );
  DFF \u_a23_mem/p_mem_reg[11][1]  ( .D(\u_a23_mem/n19331 ), .CLK(clk), .RST(
        rst), .I(p_init[89]), .Q(\u_a23_mem/p_mem[11][1] ) );
  DFF \u_a23_mem/p_mem_reg[11][2]  ( .D(\u_a23_mem/n19330 ), .CLK(clk), .RST(
        rst), .I(p_init[90]), .Q(\u_a23_mem/p_mem[11][2] ) );
  DFF \u_a23_mem/p_mem_reg[11][3]  ( .D(\u_a23_mem/n19329 ), .CLK(clk), .RST(
        rst), .I(p_init[91]), .Q(\u_a23_mem/p_mem[11][3] ) );
  DFF \u_a23_mem/p_mem_reg[11][4]  ( .D(\u_a23_mem/n19328 ), .CLK(clk), .RST(
        rst), .I(p_init[92]), .Q(\u_a23_mem/p_mem[11][4] ) );
  DFF \u_a23_mem/p_mem_reg[11][5]  ( .D(\u_a23_mem/n19327 ), .CLK(clk), .RST(
        rst), .I(p_init[93]), .Q(\u_a23_mem/p_mem[11][5] ) );
  DFF \u_a23_mem/p_mem_reg[11][6]  ( .D(\u_a23_mem/n19326 ), .CLK(clk), .RST(
        rst), .I(p_init[94]), .Q(\u_a23_mem/p_mem[11][6] ) );
  DFF \u_a23_mem/p_mem_reg[11][7]  ( .D(\u_a23_mem/n19325 ), .CLK(clk), .RST(
        rst), .I(p_init[95]), .Q(\u_a23_mem/p_mem[11][7] ) );
  DFF \u_a23_mem/p_mem_reg[12][0]  ( .D(\u_a23_mem/n19324 ), .CLK(clk), .RST(
        rst), .I(p_init[96]), .Q(\u_a23_mem/p_mem[12][0] ) );
  DFF \u_a23_mem/p_mem_reg[12][1]  ( .D(\u_a23_mem/n19323 ), .CLK(clk), .RST(
        rst), .I(p_init[97]), .Q(\u_a23_mem/p_mem[12][1] ) );
  DFF \u_a23_mem/p_mem_reg[12][2]  ( .D(\u_a23_mem/n19322 ), .CLK(clk), .RST(
        rst), .I(p_init[98]), .Q(\u_a23_mem/p_mem[12][2] ) );
  DFF \u_a23_mem/p_mem_reg[12][3]  ( .D(\u_a23_mem/n19321 ), .CLK(clk), .RST(
        rst), .I(p_init[99]), .Q(\u_a23_mem/p_mem[12][3] ) );
  DFF \u_a23_mem/p_mem_reg[12][4]  ( .D(\u_a23_mem/n19320 ), .CLK(clk), .RST(
        rst), .I(p_init[100]), .Q(\u_a23_mem/p_mem[12][4] ) );
  DFF \u_a23_mem/p_mem_reg[12][5]  ( .D(\u_a23_mem/n19319 ), .CLK(clk), .RST(
        rst), .I(p_init[101]), .Q(\u_a23_mem/p_mem[12][5] ) );
  DFF \u_a23_mem/p_mem_reg[12][6]  ( .D(\u_a23_mem/n19318 ), .CLK(clk), .RST(
        rst), .I(p_init[102]), .Q(\u_a23_mem/p_mem[12][6] ) );
  DFF \u_a23_mem/p_mem_reg[12][7]  ( .D(\u_a23_mem/n19317 ), .CLK(clk), .RST(
        rst), .I(p_init[103]), .Q(\u_a23_mem/p_mem[12][7] ) );
  DFF \u_a23_mem/p_mem_reg[13][0]  ( .D(\u_a23_mem/n19316 ), .CLK(clk), .RST(
        rst), .I(p_init[104]), .Q(\u_a23_mem/p_mem[13][0] ) );
  DFF \u_a23_mem/p_mem_reg[13][1]  ( .D(\u_a23_mem/n19315 ), .CLK(clk), .RST(
        rst), .I(p_init[105]), .Q(\u_a23_mem/p_mem[13][1] ) );
  DFF \u_a23_mem/p_mem_reg[13][2]  ( .D(\u_a23_mem/n19314 ), .CLK(clk), .RST(
        rst), .I(p_init[106]), .Q(\u_a23_mem/p_mem[13][2] ) );
  DFF \u_a23_mem/p_mem_reg[13][3]  ( .D(\u_a23_mem/n19313 ), .CLK(clk), .RST(
        rst), .I(p_init[107]), .Q(\u_a23_mem/p_mem[13][3] ) );
  DFF \u_a23_mem/p_mem_reg[13][4]  ( .D(\u_a23_mem/n19312 ), .CLK(clk), .RST(
        rst), .I(p_init[108]), .Q(\u_a23_mem/p_mem[13][4] ) );
  DFF \u_a23_mem/p_mem_reg[13][5]  ( .D(\u_a23_mem/n19311 ), .CLK(clk), .RST(
        rst), .I(p_init[109]), .Q(\u_a23_mem/p_mem[13][5] ) );
  DFF \u_a23_mem/p_mem_reg[13][6]  ( .D(\u_a23_mem/n19310 ), .CLK(clk), .RST(
        rst), .I(p_init[110]), .Q(\u_a23_mem/p_mem[13][6] ) );
  DFF \u_a23_mem/p_mem_reg[13][7]  ( .D(\u_a23_mem/n19309 ), .CLK(clk), .RST(
        rst), .I(p_init[111]), .Q(\u_a23_mem/p_mem[13][7] ) );
  DFF \u_a23_mem/p_mem_reg[14][0]  ( .D(\u_a23_mem/n19308 ), .CLK(clk), .RST(
        rst), .I(p_init[112]), .Q(\u_a23_mem/p_mem[14][0] ) );
  DFF \u_a23_mem/p_mem_reg[14][1]  ( .D(\u_a23_mem/n19307 ), .CLK(clk), .RST(
        rst), .I(p_init[113]), .Q(\u_a23_mem/p_mem[14][1] ) );
  DFF \u_a23_mem/p_mem_reg[14][2]  ( .D(\u_a23_mem/n19306 ), .CLK(clk), .RST(
        rst), .I(p_init[114]), .Q(\u_a23_mem/p_mem[14][2] ) );
  DFF \u_a23_mem/p_mem_reg[14][3]  ( .D(\u_a23_mem/n19305 ), .CLK(clk), .RST(
        rst), .I(p_init[115]), .Q(\u_a23_mem/p_mem[14][3] ) );
  DFF \u_a23_mem/p_mem_reg[14][4]  ( .D(\u_a23_mem/n19304 ), .CLK(clk), .RST(
        rst), .I(p_init[116]), .Q(\u_a23_mem/p_mem[14][4] ) );
  DFF \u_a23_mem/p_mem_reg[14][5]  ( .D(\u_a23_mem/n19303 ), .CLK(clk), .RST(
        rst), .I(p_init[117]), .Q(\u_a23_mem/p_mem[14][5] ) );
  DFF \u_a23_mem/p_mem_reg[14][6]  ( .D(\u_a23_mem/n19302 ), .CLK(clk), .RST(
        rst), .I(p_init[118]), .Q(\u_a23_mem/p_mem[14][6] ) );
  DFF \u_a23_mem/p_mem_reg[14][7]  ( .D(\u_a23_mem/n19301 ), .CLK(clk), .RST(
        rst), .I(p_init[119]), .Q(\u_a23_mem/p_mem[14][7] ) );
  DFF \u_a23_mem/p_mem_reg[15][0]  ( .D(\u_a23_mem/n19300 ), .CLK(clk), .RST(
        rst), .I(p_init[120]), .Q(\u_a23_mem/p_mem[15][0] ) );
  DFF \u_a23_mem/p_mem_reg[15][1]  ( .D(\u_a23_mem/n19299 ), .CLK(clk), .RST(
        rst), .I(p_init[121]), .Q(\u_a23_mem/p_mem[15][1] ) );
  DFF \u_a23_mem/p_mem_reg[15][2]  ( .D(\u_a23_mem/n19298 ), .CLK(clk), .RST(
        rst), .I(p_init[122]), .Q(\u_a23_mem/p_mem[15][2] ) );
  DFF \u_a23_mem/p_mem_reg[15][3]  ( .D(\u_a23_mem/n19297 ), .CLK(clk), .RST(
        rst), .I(p_init[123]), .Q(\u_a23_mem/p_mem[15][3] ) );
  DFF \u_a23_mem/p_mem_reg[15][4]  ( .D(\u_a23_mem/n19296 ), .CLK(clk), .RST(
        rst), .I(p_init[124]), .Q(\u_a23_mem/p_mem[15][4] ) );
  DFF \u_a23_mem/p_mem_reg[15][5]  ( .D(\u_a23_mem/n19295 ), .CLK(clk), .RST(
        rst), .I(p_init[125]), .Q(\u_a23_mem/p_mem[15][5] ) );
  DFF \u_a23_mem/p_mem_reg[15][6]  ( .D(\u_a23_mem/n19294 ), .CLK(clk), .RST(
        rst), .I(p_init[126]), .Q(\u_a23_mem/p_mem[15][6] ) );
  DFF \u_a23_mem/p_mem_reg[15][7]  ( .D(\u_a23_mem/n19293 ), .CLK(clk), .RST(
        rst), .I(p_init[127]), .Q(\u_a23_mem/p_mem[15][7] ) );
  DFF \u_a23_mem/p_mem_reg[16][0]  ( .D(\u_a23_mem/n19292 ), .CLK(clk), .RST(
        rst), .I(p_init[128]), .Q(\u_a23_mem/p_mem[16][0] ) );
  DFF \u_a23_mem/p_mem_reg[16][1]  ( .D(\u_a23_mem/n19291 ), .CLK(clk), .RST(
        rst), .I(p_init[129]), .Q(\u_a23_mem/p_mem[16][1] ) );
  DFF \u_a23_mem/p_mem_reg[16][2]  ( .D(\u_a23_mem/n19290 ), .CLK(clk), .RST(
        rst), .I(p_init[130]), .Q(\u_a23_mem/p_mem[16][2] ) );
  DFF \u_a23_mem/p_mem_reg[16][3]  ( .D(\u_a23_mem/n19289 ), .CLK(clk), .RST(
        rst), .I(p_init[131]), .Q(\u_a23_mem/p_mem[16][3] ) );
  DFF \u_a23_mem/p_mem_reg[16][4]  ( .D(\u_a23_mem/n19288 ), .CLK(clk), .RST(
        rst), .I(p_init[132]), .Q(\u_a23_mem/p_mem[16][4] ) );
  DFF \u_a23_mem/p_mem_reg[16][5]  ( .D(\u_a23_mem/n19287 ), .CLK(clk), .RST(
        rst), .I(p_init[133]), .Q(\u_a23_mem/p_mem[16][5] ) );
  DFF \u_a23_mem/p_mem_reg[16][6]  ( .D(\u_a23_mem/n19286 ), .CLK(clk), .RST(
        rst), .I(p_init[134]), .Q(\u_a23_mem/p_mem[16][6] ) );
  DFF \u_a23_mem/p_mem_reg[16][7]  ( .D(\u_a23_mem/n19285 ), .CLK(clk), .RST(
        rst), .I(p_init[135]), .Q(\u_a23_mem/p_mem[16][7] ) );
  DFF \u_a23_mem/p_mem_reg[17][0]  ( .D(\u_a23_mem/n19284 ), .CLK(clk), .RST(
        rst), .I(p_init[136]), .Q(\u_a23_mem/p_mem[17][0] ) );
  DFF \u_a23_mem/p_mem_reg[17][1]  ( .D(\u_a23_mem/n19283 ), .CLK(clk), .RST(
        rst), .I(p_init[137]), .Q(\u_a23_mem/p_mem[17][1] ) );
  DFF \u_a23_mem/p_mem_reg[17][2]  ( .D(\u_a23_mem/n19282 ), .CLK(clk), .RST(
        rst), .I(p_init[138]), .Q(\u_a23_mem/p_mem[17][2] ) );
  DFF \u_a23_mem/p_mem_reg[17][3]  ( .D(\u_a23_mem/n19281 ), .CLK(clk), .RST(
        rst), .I(p_init[139]), .Q(\u_a23_mem/p_mem[17][3] ) );
  DFF \u_a23_mem/p_mem_reg[17][4]  ( .D(\u_a23_mem/n19280 ), .CLK(clk), .RST(
        rst), .I(p_init[140]), .Q(\u_a23_mem/p_mem[17][4] ) );
  DFF \u_a23_mem/p_mem_reg[17][5]  ( .D(\u_a23_mem/n19279 ), .CLK(clk), .RST(
        rst), .I(p_init[141]), .Q(\u_a23_mem/p_mem[17][5] ) );
  DFF \u_a23_mem/p_mem_reg[17][6]  ( .D(\u_a23_mem/n19278 ), .CLK(clk), .RST(
        rst), .I(p_init[142]), .Q(\u_a23_mem/p_mem[17][6] ) );
  DFF \u_a23_mem/p_mem_reg[17][7]  ( .D(\u_a23_mem/n19277 ), .CLK(clk), .RST(
        rst), .I(p_init[143]), .Q(\u_a23_mem/p_mem[17][7] ) );
  DFF \u_a23_mem/p_mem_reg[18][0]  ( .D(\u_a23_mem/n19276 ), .CLK(clk), .RST(
        rst), .I(p_init[144]), .Q(\u_a23_mem/p_mem[18][0] ) );
  DFF \u_a23_mem/p_mem_reg[18][1]  ( .D(\u_a23_mem/n19275 ), .CLK(clk), .RST(
        rst), .I(p_init[145]), .Q(\u_a23_mem/p_mem[18][1] ) );
  DFF \u_a23_mem/p_mem_reg[18][2]  ( .D(\u_a23_mem/n19274 ), .CLK(clk), .RST(
        rst), .I(p_init[146]), .Q(\u_a23_mem/p_mem[18][2] ) );
  DFF \u_a23_mem/p_mem_reg[18][3]  ( .D(\u_a23_mem/n19273 ), .CLK(clk), .RST(
        rst), .I(p_init[147]), .Q(\u_a23_mem/p_mem[18][3] ) );
  DFF \u_a23_mem/p_mem_reg[18][4]  ( .D(\u_a23_mem/n19272 ), .CLK(clk), .RST(
        rst), .I(p_init[148]), .Q(\u_a23_mem/p_mem[18][4] ) );
  DFF \u_a23_mem/p_mem_reg[18][5]  ( .D(\u_a23_mem/n19271 ), .CLK(clk), .RST(
        rst), .I(p_init[149]), .Q(\u_a23_mem/p_mem[18][5] ) );
  DFF \u_a23_mem/p_mem_reg[18][6]  ( .D(\u_a23_mem/n19270 ), .CLK(clk), .RST(
        rst), .I(p_init[150]), .Q(\u_a23_mem/p_mem[18][6] ) );
  DFF \u_a23_mem/p_mem_reg[18][7]  ( .D(\u_a23_mem/n19269 ), .CLK(clk), .RST(
        rst), .I(p_init[151]), .Q(\u_a23_mem/p_mem[18][7] ) );
  DFF \u_a23_mem/p_mem_reg[19][0]  ( .D(\u_a23_mem/n19268 ), .CLK(clk), .RST(
        rst), .I(p_init[152]), .Q(\u_a23_mem/p_mem[19][0] ) );
  DFF \u_a23_mem/p_mem_reg[19][1]  ( .D(\u_a23_mem/n19267 ), .CLK(clk), .RST(
        rst), .I(p_init[153]), .Q(\u_a23_mem/p_mem[19][1] ) );
  DFF \u_a23_mem/p_mem_reg[19][2]  ( .D(\u_a23_mem/n19266 ), .CLK(clk), .RST(
        rst), .I(p_init[154]), .Q(\u_a23_mem/p_mem[19][2] ) );
  DFF \u_a23_mem/p_mem_reg[19][3]  ( .D(\u_a23_mem/n19265 ), .CLK(clk), .RST(
        rst), .I(p_init[155]), .Q(\u_a23_mem/p_mem[19][3] ) );
  DFF \u_a23_mem/p_mem_reg[19][4]  ( .D(\u_a23_mem/n19264 ), .CLK(clk), .RST(
        rst), .I(p_init[156]), .Q(\u_a23_mem/p_mem[19][4] ) );
  DFF \u_a23_mem/p_mem_reg[19][5]  ( .D(\u_a23_mem/n19263 ), .CLK(clk), .RST(
        rst), .I(p_init[157]), .Q(\u_a23_mem/p_mem[19][5] ) );
  DFF \u_a23_mem/p_mem_reg[19][6]  ( .D(\u_a23_mem/n19262 ), .CLK(clk), .RST(
        rst), .I(p_init[158]), .Q(\u_a23_mem/p_mem[19][6] ) );
  DFF \u_a23_mem/p_mem_reg[19][7]  ( .D(\u_a23_mem/n19261 ), .CLK(clk), .RST(
        rst), .I(p_init[159]), .Q(\u_a23_mem/p_mem[19][7] ) );
  DFF \u_a23_mem/p_mem_reg[20][0]  ( .D(\u_a23_mem/n19260 ), .CLK(clk), .RST(
        rst), .I(p_init[160]), .Q(\u_a23_mem/p_mem[20][0] ) );
  DFF \u_a23_mem/p_mem_reg[20][1]  ( .D(\u_a23_mem/n19259 ), .CLK(clk), .RST(
        rst), .I(p_init[161]), .Q(\u_a23_mem/p_mem[20][1] ) );
  DFF \u_a23_mem/p_mem_reg[20][2]  ( .D(\u_a23_mem/n19258 ), .CLK(clk), .RST(
        rst), .I(p_init[162]), .Q(\u_a23_mem/p_mem[20][2] ) );
  DFF \u_a23_mem/p_mem_reg[20][3]  ( .D(\u_a23_mem/n19257 ), .CLK(clk), .RST(
        rst), .I(p_init[163]), .Q(\u_a23_mem/p_mem[20][3] ) );
  DFF \u_a23_mem/p_mem_reg[20][4]  ( .D(\u_a23_mem/n19256 ), .CLK(clk), .RST(
        rst), .I(p_init[164]), .Q(\u_a23_mem/p_mem[20][4] ) );
  DFF \u_a23_mem/p_mem_reg[20][5]  ( .D(\u_a23_mem/n19255 ), .CLK(clk), .RST(
        rst), .I(p_init[165]), .Q(\u_a23_mem/p_mem[20][5] ) );
  DFF \u_a23_mem/p_mem_reg[20][6]  ( .D(\u_a23_mem/n19254 ), .CLK(clk), .RST(
        rst), .I(p_init[166]), .Q(\u_a23_mem/p_mem[20][6] ) );
  DFF \u_a23_mem/p_mem_reg[20][7]  ( .D(\u_a23_mem/n19253 ), .CLK(clk), .RST(
        rst), .I(p_init[167]), .Q(\u_a23_mem/p_mem[20][7] ) );
  DFF \u_a23_mem/p_mem_reg[21][0]  ( .D(\u_a23_mem/n19252 ), .CLK(clk), .RST(
        rst), .I(p_init[168]), .Q(\u_a23_mem/p_mem[21][0] ) );
  DFF \u_a23_mem/p_mem_reg[21][1]  ( .D(\u_a23_mem/n19251 ), .CLK(clk), .RST(
        rst), .I(p_init[169]), .Q(\u_a23_mem/p_mem[21][1] ) );
  DFF \u_a23_mem/p_mem_reg[21][2]  ( .D(\u_a23_mem/n19250 ), .CLK(clk), .RST(
        rst), .I(p_init[170]), .Q(\u_a23_mem/p_mem[21][2] ) );
  DFF \u_a23_mem/p_mem_reg[21][3]  ( .D(\u_a23_mem/n19249 ), .CLK(clk), .RST(
        rst), .I(p_init[171]), .Q(\u_a23_mem/p_mem[21][3] ) );
  DFF \u_a23_mem/p_mem_reg[21][4]  ( .D(\u_a23_mem/n19248 ), .CLK(clk), .RST(
        rst), .I(p_init[172]), .Q(\u_a23_mem/p_mem[21][4] ) );
  DFF \u_a23_mem/p_mem_reg[21][5]  ( .D(\u_a23_mem/n19247 ), .CLK(clk), .RST(
        rst), .I(p_init[173]), .Q(\u_a23_mem/p_mem[21][5] ) );
  DFF \u_a23_mem/p_mem_reg[21][6]  ( .D(\u_a23_mem/n19246 ), .CLK(clk), .RST(
        rst), .I(p_init[174]), .Q(\u_a23_mem/p_mem[21][6] ) );
  DFF \u_a23_mem/p_mem_reg[21][7]  ( .D(\u_a23_mem/n19245 ), .CLK(clk), .RST(
        rst), .I(p_init[175]), .Q(\u_a23_mem/p_mem[21][7] ) );
  DFF \u_a23_mem/p_mem_reg[22][0]  ( .D(\u_a23_mem/n19244 ), .CLK(clk), .RST(
        rst), .I(p_init[176]), .Q(\u_a23_mem/p_mem[22][0] ) );
  DFF \u_a23_mem/p_mem_reg[22][1]  ( .D(\u_a23_mem/n19243 ), .CLK(clk), .RST(
        rst), .I(p_init[177]), .Q(\u_a23_mem/p_mem[22][1] ) );
  DFF \u_a23_mem/p_mem_reg[22][2]  ( .D(\u_a23_mem/n19242 ), .CLK(clk), .RST(
        rst), .I(p_init[178]), .Q(\u_a23_mem/p_mem[22][2] ) );
  DFF \u_a23_mem/p_mem_reg[22][3]  ( .D(\u_a23_mem/n19241 ), .CLK(clk), .RST(
        rst), .I(p_init[179]), .Q(\u_a23_mem/p_mem[22][3] ) );
  DFF \u_a23_mem/p_mem_reg[22][4]  ( .D(\u_a23_mem/n19240 ), .CLK(clk), .RST(
        rst), .I(p_init[180]), .Q(\u_a23_mem/p_mem[22][4] ) );
  DFF \u_a23_mem/p_mem_reg[22][5]  ( .D(\u_a23_mem/n19239 ), .CLK(clk), .RST(
        rst), .I(p_init[181]), .Q(\u_a23_mem/p_mem[22][5] ) );
  DFF \u_a23_mem/p_mem_reg[22][6]  ( .D(\u_a23_mem/n19238 ), .CLK(clk), .RST(
        rst), .I(p_init[182]), .Q(\u_a23_mem/p_mem[22][6] ) );
  DFF \u_a23_mem/p_mem_reg[22][7]  ( .D(\u_a23_mem/n19237 ), .CLK(clk), .RST(
        rst), .I(p_init[183]), .Q(\u_a23_mem/p_mem[22][7] ) );
  DFF \u_a23_mem/p_mem_reg[23][0]  ( .D(\u_a23_mem/n19236 ), .CLK(clk), .RST(
        rst), .I(p_init[184]), .Q(\u_a23_mem/p_mem[23][0] ) );
  DFF \u_a23_mem/p_mem_reg[23][1]  ( .D(\u_a23_mem/n19235 ), .CLK(clk), .RST(
        rst), .I(p_init[185]), .Q(\u_a23_mem/p_mem[23][1] ) );
  DFF \u_a23_mem/p_mem_reg[23][2]  ( .D(\u_a23_mem/n19234 ), .CLK(clk), .RST(
        rst), .I(p_init[186]), .Q(\u_a23_mem/p_mem[23][2] ) );
  DFF \u_a23_mem/p_mem_reg[23][3]  ( .D(\u_a23_mem/n19233 ), .CLK(clk), .RST(
        rst), .I(p_init[187]), .Q(\u_a23_mem/p_mem[23][3] ) );
  DFF \u_a23_mem/p_mem_reg[23][4]  ( .D(\u_a23_mem/n19232 ), .CLK(clk), .RST(
        rst), .I(p_init[188]), .Q(\u_a23_mem/p_mem[23][4] ) );
  DFF \u_a23_mem/p_mem_reg[23][5]  ( .D(\u_a23_mem/n19231 ), .CLK(clk), .RST(
        rst), .I(p_init[189]), .Q(\u_a23_mem/p_mem[23][5] ) );
  DFF \u_a23_mem/p_mem_reg[23][6]  ( .D(\u_a23_mem/n19230 ), .CLK(clk), .RST(
        rst), .I(p_init[190]), .Q(\u_a23_mem/p_mem[23][6] ) );
  DFF \u_a23_mem/p_mem_reg[23][7]  ( .D(\u_a23_mem/n19229 ), .CLK(clk), .RST(
        rst), .I(p_init[191]), .Q(\u_a23_mem/p_mem[23][7] ) );
  DFF \u_a23_mem/p_mem_reg[24][0]  ( .D(\u_a23_mem/n19228 ), .CLK(clk), .RST(
        rst), .I(p_init[192]), .Q(\u_a23_mem/p_mem[24][0] ) );
  DFF \u_a23_mem/p_mem_reg[24][1]  ( .D(\u_a23_mem/n19227 ), .CLK(clk), .RST(
        rst), .I(p_init[193]), .Q(\u_a23_mem/p_mem[24][1] ) );
  DFF \u_a23_mem/p_mem_reg[24][2]  ( .D(\u_a23_mem/n19226 ), .CLK(clk), .RST(
        rst), .I(p_init[194]), .Q(\u_a23_mem/p_mem[24][2] ) );
  DFF \u_a23_mem/p_mem_reg[24][3]  ( .D(\u_a23_mem/n19225 ), .CLK(clk), .RST(
        rst), .I(p_init[195]), .Q(\u_a23_mem/p_mem[24][3] ) );
  DFF \u_a23_mem/p_mem_reg[24][4]  ( .D(\u_a23_mem/n19224 ), .CLK(clk), .RST(
        rst), .I(p_init[196]), .Q(\u_a23_mem/p_mem[24][4] ) );
  DFF \u_a23_mem/p_mem_reg[24][5]  ( .D(\u_a23_mem/n19223 ), .CLK(clk), .RST(
        rst), .I(p_init[197]), .Q(\u_a23_mem/p_mem[24][5] ) );
  DFF \u_a23_mem/p_mem_reg[24][6]  ( .D(\u_a23_mem/n19222 ), .CLK(clk), .RST(
        rst), .I(p_init[198]), .Q(\u_a23_mem/p_mem[24][6] ) );
  DFF \u_a23_mem/p_mem_reg[24][7]  ( .D(\u_a23_mem/n19221 ), .CLK(clk), .RST(
        rst), .I(p_init[199]), .Q(\u_a23_mem/p_mem[24][7] ) );
  DFF \u_a23_mem/p_mem_reg[25][0]  ( .D(\u_a23_mem/n19220 ), .CLK(clk), .RST(
        rst), .I(p_init[200]), .Q(\u_a23_mem/p_mem[25][0] ) );
  DFF \u_a23_mem/p_mem_reg[25][1]  ( .D(\u_a23_mem/n19219 ), .CLK(clk), .RST(
        rst), .I(p_init[201]), .Q(\u_a23_mem/p_mem[25][1] ) );
  DFF \u_a23_mem/p_mem_reg[25][2]  ( .D(\u_a23_mem/n19218 ), .CLK(clk), .RST(
        rst), .I(p_init[202]), .Q(\u_a23_mem/p_mem[25][2] ) );
  DFF \u_a23_mem/p_mem_reg[25][3]  ( .D(\u_a23_mem/n19217 ), .CLK(clk), .RST(
        rst), .I(p_init[203]), .Q(\u_a23_mem/p_mem[25][3] ) );
  DFF \u_a23_mem/p_mem_reg[25][4]  ( .D(\u_a23_mem/n19216 ), .CLK(clk), .RST(
        rst), .I(p_init[204]), .Q(\u_a23_mem/p_mem[25][4] ) );
  DFF \u_a23_mem/p_mem_reg[25][5]  ( .D(\u_a23_mem/n19215 ), .CLK(clk), .RST(
        rst), .I(p_init[205]), .Q(\u_a23_mem/p_mem[25][5] ) );
  DFF \u_a23_mem/p_mem_reg[25][6]  ( .D(\u_a23_mem/n19214 ), .CLK(clk), .RST(
        rst), .I(p_init[206]), .Q(\u_a23_mem/p_mem[25][6] ) );
  DFF \u_a23_mem/p_mem_reg[25][7]  ( .D(\u_a23_mem/n19213 ), .CLK(clk), .RST(
        rst), .I(p_init[207]), .Q(\u_a23_mem/p_mem[25][7] ) );
  DFF \u_a23_mem/p_mem_reg[26][0]  ( .D(\u_a23_mem/n19212 ), .CLK(clk), .RST(
        rst), .I(p_init[208]), .Q(\u_a23_mem/p_mem[26][0] ) );
  DFF \u_a23_mem/p_mem_reg[26][1]  ( .D(\u_a23_mem/n19211 ), .CLK(clk), .RST(
        rst), .I(p_init[209]), .Q(\u_a23_mem/p_mem[26][1] ) );
  DFF \u_a23_mem/p_mem_reg[26][2]  ( .D(\u_a23_mem/n19210 ), .CLK(clk), .RST(
        rst), .I(p_init[210]), .Q(\u_a23_mem/p_mem[26][2] ) );
  DFF \u_a23_mem/p_mem_reg[26][3]  ( .D(\u_a23_mem/n19209 ), .CLK(clk), .RST(
        rst), .I(p_init[211]), .Q(\u_a23_mem/p_mem[26][3] ) );
  DFF \u_a23_mem/p_mem_reg[26][4]  ( .D(\u_a23_mem/n19208 ), .CLK(clk), .RST(
        rst), .I(p_init[212]), .Q(\u_a23_mem/p_mem[26][4] ) );
  DFF \u_a23_mem/p_mem_reg[26][5]  ( .D(\u_a23_mem/n19207 ), .CLK(clk), .RST(
        rst), .I(p_init[213]), .Q(\u_a23_mem/p_mem[26][5] ) );
  DFF \u_a23_mem/p_mem_reg[26][6]  ( .D(\u_a23_mem/n19206 ), .CLK(clk), .RST(
        rst), .I(p_init[214]), .Q(\u_a23_mem/p_mem[26][6] ) );
  DFF \u_a23_mem/p_mem_reg[26][7]  ( .D(\u_a23_mem/n19205 ), .CLK(clk), .RST(
        rst), .I(p_init[215]), .Q(\u_a23_mem/p_mem[26][7] ) );
  DFF \u_a23_mem/p_mem_reg[27][0]  ( .D(\u_a23_mem/n19204 ), .CLK(clk), .RST(
        rst), .I(p_init[216]), .Q(\u_a23_mem/p_mem[27][0] ) );
  DFF \u_a23_mem/p_mem_reg[27][1]  ( .D(\u_a23_mem/n19203 ), .CLK(clk), .RST(
        rst), .I(p_init[217]), .Q(\u_a23_mem/p_mem[27][1] ) );
  DFF \u_a23_mem/p_mem_reg[27][2]  ( .D(\u_a23_mem/n19202 ), .CLK(clk), .RST(
        rst), .I(p_init[218]), .Q(\u_a23_mem/p_mem[27][2] ) );
  DFF \u_a23_mem/p_mem_reg[27][3]  ( .D(\u_a23_mem/n19201 ), .CLK(clk), .RST(
        rst), .I(p_init[219]), .Q(\u_a23_mem/p_mem[27][3] ) );
  DFF \u_a23_mem/p_mem_reg[27][4]  ( .D(\u_a23_mem/n19200 ), .CLK(clk), .RST(
        rst), .I(p_init[220]), .Q(\u_a23_mem/p_mem[27][4] ) );
  DFF \u_a23_mem/p_mem_reg[27][5]  ( .D(\u_a23_mem/n19199 ), .CLK(clk), .RST(
        rst), .I(p_init[221]), .Q(\u_a23_mem/p_mem[27][5] ) );
  DFF \u_a23_mem/p_mem_reg[27][6]  ( .D(\u_a23_mem/n19198 ), .CLK(clk), .RST(
        rst), .I(p_init[222]), .Q(\u_a23_mem/p_mem[27][6] ) );
  DFF \u_a23_mem/p_mem_reg[27][7]  ( .D(\u_a23_mem/n19197 ), .CLK(clk), .RST(
        rst), .I(p_init[223]), .Q(\u_a23_mem/p_mem[27][7] ) );
  DFF \u_a23_mem/p_mem_reg[28][0]  ( .D(\u_a23_mem/n19196 ), .CLK(clk), .RST(
        rst), .I(p_init[224]), .Q(\u_a23_mem/p_mem[28][0] ) );
  DFF \u_a23_mem/p_mem_reg[28][1]  ( .D(\u_a23_mem/n19195 ), .CLK(clk), .RST(
        rst), .I(p_init[225]), .Q(\u_a23_mem/p_mem[28][1] ) );
  DFF \u_a23_mem/p_mem_reg[28][2]  ( .D(\u_a23_mem/n19194 ), .CLK(clk), .RST(
        rst), .I(p_init[226]), .Q(\u_a23_mem/p_mem[28][2] ) );
  DFF \u_a23_mem/p_mem_reg[28][3]  ( .D(\u_a23_mem/n19193 ), .CLK(clk), .RST(
        rst), .I(p_init[227]), .Q(\u_a23_mem/p_mem[28][3] ) );
  DFF \u_a23_mem/p_mem_reg[28][4]  ( .D(\u_a23_mem/n19192 ), .CLK(clk), .RST(
        rst), .I(p_init[228]), .Q(\u_a23_mem/p_mem[28][4] ) );
  DFF \u_a23_mem/p_mem_reg[28][5]  ( .D(\u_a23_mem/n19191 ), .CLK(clk), .RST(
        rst), .I(p_init[229]), .Q(\u_a23_mem/p_mem[28][5] ) );
  DFF \u_a23_mem/p_mem_reg[28][6]  ( .D(\u_a23_mem/n19190 ), .CLK(clk), .RST(
        rst), .I(p_init[230]), .Q(\u_a23_mem/p_mem[28][6] ) );
  DFF \u_a23_mem/p_mem_reg[28][7]  ( .D(\u_a23_mem/n19189 ), .CLK(clk), .RST(
        rst), .I(p_init[231]), .Q(\u_a23_mem/p_mem[28][7] ) );
  DFF \u_a23_mem/p_mem_reg[29][0]  ( .D(\u_a23_mem/n19188 ), .CLK(clk), .RST(
        rst), .I(p_init[232]), .Q(\u_a23_mem/p_mem[29][0] ) );
  DFF \u_a23_mem/p_mem_reg[29][1]  ( .D(\u_a23_mem/n19187 ), .CLK(clk), .RST(
        rst), .I(p_init[233]), .Q(\u_a23_mem/p_mem[29][1] ) );
  DFF \u_a23_mem/p_mem_reg[29][2]  ( .D(\u_a23_mem/n19186 ), .CLK(clk), .RST(
        rst), .I(p_init[234]), .Q(\u_a23_mem/p_mem[29][2] ) );
  DFF \u_a23_mem/p_mem_reg[29][3]  ( .D(\u_a23_mem/n19185 ), .CLK(clk), .RST(
        rst), .I(p_init[235]), .Q(\u_a23_mem/p_mem[29][3] ) );
  DFF \u_a23_mem/p_mem_reg[29][4]  ( .D(\u_a23_mem/n19184 ), .CLK(clk), .RST(
        rst), .I(p_init[236]), .Q(\u_a23_mem/p_mem[29][4] ) );
  DFF \u_a23_mem/p_mem_reg[29][5]  ( .D(\u_a23_mem/n19183 ), .CLK(clk), .RST(
        rst), .I(p_init[237]), .Q(\u_a23_mem/p_mem[29][5] ) );
  DFF \u_a23_mem/p_mem_reg[29][6]  ( .D(\u_a23_mem/n19182 ), .CLK(clk), .RST(
        rst), .I(p_init[238]), .Q(\u_a23_mem/p_mem[29][6] ) );
  DFF \u_a23_mem/p_mem_reg[29][7]  ( .D(\u_a23_mem/n19181 ), .CLK(clk), .RST(
        rst), .I(p_init[239]), .Q(\u_a23_mem/p_mem[29][7] ) );
  DFF \u_a23_mem/p_mem_reg[30][0]  ( .D(\u_a23_mem/n19180 ), .CLK(clk), .RST(
        rst), .I(p_init[240]), .Q(\u_a23_mem/p_mem[30][0] ) );
  DFF \u_a23_mem/p_mem_reg[30][1]  ( .D(\u_a23_mem/n19179 ), .CLK(clk), .RST(
        rst), .I(p_init[241]), .Q(\u_a23_mem/p_mem[30][1] ) );
  DFF \u_a23_mem/p_mem_reg[30][2]  ( .D(\u_a23_mem/n19178 ), .CLK(clk), .RST(
        rst), .I(p_init[242]), .Q(\u_a23_mem/p_mem[30][2] ) );
  DFF \u_a23_mem/p_mem_reg[30][3]  ( .D(\u_a23_mem/n19177 ), .CLK(clk), .RST(
        rst), .I(p_init[243]), .Q(\u_a23_mem/p_mem[30][3] ) );
  DFF \u_a23_mem/p_mem_reg[30][4]  ( .D(\u_a23_mem/n19176 ), .CLK(clk), .RST(
        rst), .I(p_init[244]), .Q(\u_a23_mem/p_mem[30][4] ) );
  DFF \u_a23_mem/p_mem_reg[30][5]  ( .D(\u_a23_mem/n19175 ), .CLK(clk), .RST(
        rst), .I(p_init[245]), .Q(\u_a23_mem/p_mem[30][5] ) );
  DFF \u_a23_mem/p_mem_reg[30][6]  ( .D(\u_a23_mem/n19174 ), .CLK(clk), .RST(
        rst), .I(p_init[246]), .Q(\u_a23_mem/p_mem[30][6] ) );
  DFF \u_a23_mem/p_mem_reg[30][7]  ( .D(\u_a23_mem/n19173 ), .CLK(clk), .RST(
        rst), .I(p_init[247]), .Q(\u_a23_mem/p_mem[30][7] ) );
  DFF \u_a23_mem/p_mem_reg[31][0]  ( .D(\u_a23_mem/n19172 ), .CLK(clk), .RST(
        rst), .I(p_init[248]), .Q(\u_a23_mem/p_mem[31][0] ) );
  DFF \u_a23_mem/p_mem_reg[31][1]  ( .D(\u_a23_mem/n19171 ), .CLK(clk), .RST(
        rst), .I(p_init[249]), .Q(\u_a23_mem/p_mem[31][1] ) );
  DFF \u_a23_mem/p_mem_reg[31][2]  ( .D(\u_a23_mem/n19170 ), .CLK(clk), .RST(
        rst), .I(p_init[250]), .Q(\u_a23_mem/p_mem[31][2] ) );
  DFF \u_a23_mem/p_mem_reg[31][3]  ( .D(\u_a23_mem/n19169 ), .CLK(clk), .RST(
        rst), .I(p_init[251]), .Q(\u_a23_mem/p_mem[31][3] ) );
  DFF \u_a23_mem/p_mem_reg[31][4]  ( .D(\u_a23_mem/n19168 ), .CLK(clk), .RST(
        rst), .I(p_init[252]), .Q(\u_a23_mem/p_mem[31][4] ) );
  DFF \u_a23_mem/p_mem_reg[31][5]  ( .D(\u_a23_mem/n19167 ), .CLK(clk), .RST(
        rst), .I(p_init[253]), .Q(\u_a23_mem/p_mem[31][5] ) );
  DFF \u_a23_mem/p_mem_reg[31][6]  ( .D(\u_a23_mem/n19166 ), .CLK(clk), .RST(
        rst), .I(p_init[254]), .Q(\u_a23_mem/p_mem[31][6] ) );
  DFF \u_a23_mem/p_mem_reg[31][7]  ( .D(\u_a23_mem/n19165 ), .CLK(clk), .RST(
        rst), .I(p_init[255]), .Q(\u_a23_mem/p_mem[31][7] ) );
  DFF \u_a23_mem/p_mem_reg[32][0]  ( .D(\u_a23_mem/n19164 ), .CLK(clk), .RST(
        rst), .I(p_init[256]), .Q(\u_a23_mem/p_mem[32][0] ) );
  DFF \u_a23_mem/p_mem_reg[32][1]  ( .D(\u_a23_mem/n19163 ), .CLK(clk), .RST(
        rst), .I(p_init[257]), .Q(\u_a23_mem/p_mem[32][1] ) );
  DFF \u_a23_mem/p_mem_reg[32][2]  ( .D(\u_a23_mem/n19162 ), .CLK(clk), .RST(
        rst), .I(p_init[258]), .Q(\u_a23_mem/p_mem[32][2] ) );
  DFF \u_a23_mem/p_mem_reg[32][3]  ( .D(\u_a23_mem/n19161 ), .CLK(clk), .RST(
        rst), .I(p_init[259]), .Q(\u_a23_mem/p_mem[32][3] ) );
  DFF \u_a23_mem/p_mem_reg[32][4]  ( .D(\u_a23_mem/n19160 ), .CLK(clk), .RST(
        rst), .I(p_init[260]), .Q(\u_a23_mem/p_mem[32][4] ) );
  DFF \u_a23_mem/p_mem_reg[32][5]  ( .D(\u_a23_mem/n19159 ), .CLK(clk), .RST(
        rst), .I(p_init[261]), .Q(\u_a23_mem/p_mem[32][5] ) );
  DFF \u_a23_mem/p_mem_reg[32][6]  ( .D(\u_a23_mem/n19158 ), .CLK(clk), .RST(
        rst), .I(p_init[262]), .Q(\u_a23_mem/p_mem[32][6] ) );
  DFF \u_a23_mem/p_mem_reg[32][7]  ( .D(\u_a23_mem/n19157 ), .CLK(clk), .RST(
        rst), .I(p_init[263]), .Q(\u_a23_mem/p_mem[32][7] ) );
  DFF \u_a23_mem/p_mem_reg[33][0]  ( .D(\u_a23_mem/n19156 ), .CLK(clk), .RST(
        rst), .I(p_init[264]), .Q(\u_a23_mem/p_mem[33][0] ) );
  DFF \u_a23_mem/p_mem_reg[33][1]  ( .D(\u_a23_mem/n19155 ), .CLK(clk), .RST(
        rst), .I(p_init[265]), .Q(\u_a23_mem/p_mem[33][1] ) );
  DFF \u_a23_mem/p_mem_reg[33][2]  ( .D(\u_a23_mem/n19154 ), .CLK(clk), .RST(
        rst), .I(p_init[266]), .Q(\u_a23_mem/p_mem[33][2] ) );
  DFF \u_a23_mem/p_mem_reg[33][3]  ( .D(\u_a23_mem/n19153 ), .CLK(clk), .RST(
        rst), .I(p_init[267]), .Q(\u_a23_mem/p_mem[33][3] ) );
  DFF \u_a23_mem/p_mem_reg[33][4]  ( .D(\u_a23_mem/n19152 ), .CLK(clk), .RST(
        rst), .I(p_init[268]), .Q(\u_a23_mem/p_mem[33][4] ) );
  DFF \u_a23_mem/p_mem_reg[33][5]  ( .D(\u_a23_mem/n19151 ), .CLK(clk), .RST(
        rst), .I(p_init[269]), .Q(\u_a23_mem/p_mem[33][5] ) );
  DFF \u_a23_mem/p_mem_reg[33][6]  ( .D(\u_a23_mem/n19150 ), .CLK(clk), .RST(
        rst), .I(p_init[270]), .Q(\u_a23_mem/p_mem[33][6] ) );
  DFF \u_a23_mem/p_mem_reg[33][7]  ( .D(\u_a23_mem/n19149 ), .CLK(clk), .RST(
        rst), .I(p_init[271]), .Q(\u_a23_mem/p_mem[33][7] ) );
  DFF \u_a23_mem/p_mem_reg[34][0]  ( .D(\u_a23_mem/n19148 ), .CLK(clk), .RST(
        rst), .I(p_init[272]), .Q(\u_a23_mem/p_mem[34][0] ) );
  DFF \u_a23_mem/p_mem_reg[34][1]  ( .D(\u_a23_mem/n19147 ), .CLK(clk), .RST(
        rst), .I(p_init[273]), .Q(\u_a23_mem/p_mem[34][1] ) );
  DFF \u_a23_mem/p_mem_reg[34][2]  ( .D(\u_a23_mem/n19146 ), .CLK(clk), .RST(
        rst), .I(p_init[274]), .Q(\u_a23_mem/p_mem[34][2] ) );
  DFF \u_a23_mem/p_mem_reg[34][3]  ( .D(\u_a23_mem/n19145 ), .CLK(clk), .RST(
        rst), .I(p_init[275]), .Q(\u_a23_mem/p_mem[34][3] ) );
  DFF \u_a23_mem/p_mem_reg[34][4]  ( .D(\u_a23_mem/n19144 ), .CLK(clk), .RST(
        rst), .I(p_init[276]), .Q(\u_a23_mem/p_mem[34][4] ) );
  DFF \u_a23_mem/p_mem_reg[34][5]  ( .D(\u_a23_mem/n19143 ), .CLK(clk), .RST(
        rst), .I(p_init[277]), .Q(\u_a23_mem/p_mem[34][5] ) );
  DFF \u_a23_mem/p_mem_reg[34][6]  ( .D(\u_a23_mem/n19142 ), .CLK(clk), .RST(
        rst), .I(p_init[278]), .Q(\u_a23_mem/p_mem[34][6] ) );
  DFF \u_a23_mem/p_mem_reg[34][7]  ( .D(\u_a23_mem/n19141 ), .CLK(clk), .RST(
        rst), .I(p_init[279]), .Q(\u_a23_mem/p_mem[34][7] ) );
  DFF \u_a23_mem/p_mem_reg[35][0]  ( .D(\u_a23_mem/n19140 ), .CLK(clk), .RST(
        rst), .I(p_init[280]), .Q(\u_a23_mem/p_mem[35][0] ) );
  DFF \u_a23_mem/p_mem_reg[35][1]  ( .D(\u_a23_mem/n19139 ), .CLK(clk), .RST(
        rst), .I(p_init[281]), .Q(\u_a23_mem/p_mem[35][1] ) );
  DFF \u_a23_mem/p_mem_reg[35][2]  ( .D(\u_a23_mem/n19138 ), .CLK(clk), .RST(
        rst), .I(p_init[282]), .Q(\u_a23_mem/p_mem[35][2] ) );
  DFF \u_a23_mem/p_mem_reg[35][3]  ( .D(\u_a23_mem/n19137 ), .CLK(clk), .RST(
        rst), .I(p_init[283]), .Q(\u_a23_mem/p_mem[35][3] ) );
  DFF \u_a23_mem/p_mem_reg[35][4]  ( .D(\u_a23_mem/n19136 ), .CLK(clk), .RST(
        rst), .I(p_init[284]), .Q(\u_a23_mem/p_mem[35][4] ) );
  DFF \u_a23_mem/p_mem_reg[35][5]  ( .D(\u_a23_mem/n19135 ), .CLK(clk), .RST(
        rst), .I(p_init[285]), .Q(\u_a23_mem/p_mem[35][5] ) );
  DFF \u_a23_mem/p_mem_reg[35][6]  ( .D(\u_a23_mem/n19134 ), .CLK(clk), .RST(
        rst), .I(p_init[286]), .Q(\u_a23_mem/p_mem[35][6] ) );
  DFF \u_a23_mem/p_mem_reg[35][7]  ( .D(\u_a23_mem/n19133 ), .CLK(clk), .RST(
        rst), .I(p_init[287]), .Q(\u_a23_mem/p_mem[35][7] ) );
  DFF \u_a23_mem/p_mem_reg[36][0]  ( .D(\u_a23_mem/n19132 ), .CLK(clk), .RST(
        rst), .I(p_init[288]), .Q(\u_a23_mem/p_mem[36][0] ) );
  DFF \u_a23_mem/p_mem_reg[36][1]  ( .D(\u_a23_mem/n19131 ), .CLK(clk), .RST(
        rst), .I(p_init[289]), .Q(\u_a23_mem/p_mem[36][1] ) );
  DFF \u_a23_mem/p_mem_reg[36][2]  ( .D(\u_a23_mem/n19130 ), .CLK(clk), .RST(
        rst), .I(p_init[290]), .Q(\u_a23_mem/p_mem[36][2] ) );
  DFF \u_a23_mem/p_mem_reg[36][3]  ( .D(\u_a23_mem/n19129 ), .CLK(clk), .RST(
        rst), .I(p_init[291]), .Q(\u_a23_mem/p_mem[36][3] ) );
  DFF \u_a23_mem/p_mem_reg[36][4]  ( .D(\u_a23_mem/n19128 ), .CLK(clk), .RST(
        rst), .I(p_init[292]), .Q(\u_a23_mem/p_mem[36][4] ) );
  DFF \u_a23_mem/p_mem_reg[36][5]  ( .D(\u_a23_mem/n19127 ), .CLK(clk), .RST(
        rst), .I(p_init[293]), .Q(\u_a23_mem/p_mem[36][5] ) );
  DFF \u_a23_mem/p_mem_reg[36][6]  ( .D(\u_a23_mem/n19126 ), .CLK(clk), .RST(
        rst), .I(p_init[294]), .Q(\u_a23_mem/p_mem[36][6] ) );
  DFF \u_a23_mem/p_mem_reg[36][7]  ( .D(\u_a23_mem/n19125 ), .CLK(clk), .RST(
        rst), .I(p_init[295]), .Q(\u_a23_mem/p_mem[36][7] ) );
  DFF \u_a23_mem/p_mem_reg[37][0]  ( .D(\u_a23_mem/n19124 ), .CLK(clk), .RST(
        rst), .I(p_init[296]), .Q(\u_a23_mem/p_mem[37][0] ) );
  DFF \u_a23_mem/p_mem_reg[37][1]  ( .D(\u_a23_mem/n19123 ), .CLK(clk), .RST(
        rst), .I(p_init[297]), .Q(\u_a23_mem/p_mem[37][1] ) );
  DFF \u_a23_mem/p_mem_reg[37][2]  ( .D(\u_a23_mem/n19122 ), .CLK(clk), .RST(
        rst), .I(p_init[298]), .Q(\u_a23_mem/p_mem[37][2] ) );
  DFF \u_a23_mem/p_mem_reg[37][3]  ( .D(\u_a23_mem/n19121 ), .CLK(clk), .RST(
        rst), .I(p_init[299]), .Q(\u_a23_mem/p_mem[37][3] ) );
  DFF \u_a23_mem/p_mem_reg[37][4]  ( .D(\u_a23_mem/n19120 ), .CLK(clk), .RST(
        rst), .I(p_init[300]), .Q(\u_a23_mem/p_mem[37][4] ) );
  DFF \u_a23_mem/p_mem_reg[37][5]  ( .D(\u_a23_mem/n19119 ), .CLK(clk), .RST(
        rst), .I(p_init[301]), .Q(\u_a23_mem/p_mem[37][5] ) );
  DFF \u_a23_mem/p_mem_reg[37][6]  ( .D(\u_a23_mem/n19118 ), .CLK(clk), .RST(
        rst), .I(p_init[302]), .Q(\u_a23_mem/p_mem[37][6] ) );
  DFF \u_a23_mem/p_mem_reg[37][7]  ( .D(\u_a23_mem/n19117 ), .CLK(clk), .RST(
        rst), .I(p_init[303]), .Q(\u_a23_mem/p_mem[37][7] ) );
  DFF \u_a23_mem/p_mem_reg[38][0]  ( .D(\u_a23_mem/n19116 ), .CLK(clk), .RST(
        rst), .I(p_init[304]), .Q(\u_a23_mem/p_mem[38][0] ) );
  DFF \u_a23_mem/p_mem_reg[38][1]  ( .D(\u_a23_mem/n19115 ), .CLK(clk), .RST(
        rst), .I(p_init[305]), .Q(\u_a23_mem/p_mem[38][1] ) );
  DFF \u_a23_mem/p_mem_reg[38][2]  ( .D(\u_a23_mem/n19114 ), .CLK(clk), .RST(
        rst), .I(p_init[306]), .Q(\u_a23_mem/p_mem[38][2] ) );
  DFF \u_a23_mem/p_mem_reg[38][3]  ( .D(\u_a23_mem/n19113 ), .CLK(clk), .RST(
        rst), .I(p_init[307]), .Q(\u_a23_mem/p_mem[38][3] ) );
  DFF \u_a23_mem/p_mem_reg[38][4]  ( .D(\u_a23_mem/n19112 ), .CLK(clk), .RST(
        rst), .I(p_init[308]), .Q(\u_a23_mem/p_mem[38][4] ) );
  DFF \u_a23_mem/p_mem_reg[38][5]  ( .D(\u_a23_mem/n19111 ), .CLK(clk), .RST(
        rst), .I(p_init[309]), .Q(\u_a23_mem/p_mem[38][5] ) );
  DFF \u_a23_mem/p_mem_reg[38][6]  ( .D(\u_a23_mem/n19110 ), .CLK(clk), .RST(
        rst), .I(p_init[310]), .Q(\u_a23_mem/p_mem[38][6] ) );
  DFF \u_a23_mem/p_mem_reg[38][7]  ( .D(\u_a23_mem/n19109 ), .CLK(clk), .RST(
        rst), .I(p_init[311]), .Q(\u_a23_mem/p_mem[38][7] ) );
  DFF \u_a23_mem/p_mem_reg[39][0]  ( .D(\u_a23_mem/n19108 ), .CLK(clk), .RST(
        rst), .I(p_init[312]), .Q(\u_a23_mem/p_mem[39][0] ) );
  DFF \u_a23_mem/p_mem_reg[39][1]  ( .D(\u_a23_mem/n19107 ), .CLK(clk), .RST(
        rst), .I(p_init[313]), .Q(\u_a23_mem/p_mem[39][1] ) );
  DFF \u_a23_mem/p_mem_reg[39][2]  ( .D(\u_a23_mem/n19106 ), .CLK(clk), .RST(
        rst), .I(p_init[314]), .Q(\u_a23_mem/p_mem[39][2] ) );
  DFF \u_a23_mem/p_mem_reg[39][3]  ( .D(\u_a23_mem/n19105 ), .CLK(clk), .RST(
        rst), .I(p_init[315]), .Q(\u_a23_mem/p_mem[39][3] ) );
  DFF \u_a23_mem/p_mem_reg[39][4]  ( .D(\u_a23_mem/n19104 ), .CLK(clk), .RST(
        rst), .I(p_init[316]), .Q(\u_a23_mem/p_mem[39][4] ) );
  DFF \u_a23_mem/p_mem_reg[39][5]  ( .D(\u_a23_mem/n19103 ), .CLK(clk), .RST(
        rst), .I(p_init[317]), .Q(\u_a23_mem/p_mem[39][5] ) );
  DFF \u_a23_mem/p_mem_reg[39][6]  ( .D(\u_a23_mem/n19102 ), .CLK(clk), .RST(
        rst), .I(p_init[318]), .Q(\u_a23_mem/p_mem[39][6] ) );
  DFF \u_a23_mem/p_mem_reg[39][7]  ( .D(\u_a23_mem/n19101 ), .CLK(clk), .RST(
        rst), .I(p_init[319]), .Q(\u_a23_mem/p_mem[39][7] ) );
  DFF \u_a23_mem/p_mem_reg[40][0]  ( .D(\u_a23_mem/n19100 ), .CLK(clk), .RST(
        rst), .I(p_init[320]), .Q(\u_a23_mem/p_mem[40][0] ) );
  DFF \u_a23_mem/p_mem_reg[40][1]  ( .D(\u_a23_mem/n19099 ), .CLK(clk), .RST(
        rst), .I(p_init[321]), .Q(\u_a23_mem/p_mem[40][1] ) );
  DFF \u_a23_mem/p_mem_reg[40][2]  ( .D(\u_a23_mem/n19098 ), .CLK(clk), .RST(
        rst), .I(p_init[322]), .Q(\u_a23_mem/p_mem[40][2] ) );
  DFF \u_a23_mem/p_mem_reg[40][3]  ( .D(\u_a23_mem/n19097 ), .CLK(clk), .RST(
        rst), .I(p_init[323]), .Q(\u_a23_mem/p_mem[40][3] ) );
  DFF \u_a23_mem/p_mem_reg[40][4]  ( .D(\u_a23_mem/n19096 ), .CLK(clk), .RST(
        rst), .I(p_init[324]), .Q(\u_a23_mem/p_mem[40][4] ) );
  DFF \u_a23_mem/p_mem_reg[40][5]  ( .D(\u_a23_mem/n19095 ), .CLK(clk), .RST(
        rst), .I(p_init[325]), .Q(\u_a23_mem/p_mem[40][5] ) );
  DFF \u_a23_mem/p_mem_reg[40][6]  ( .D(\u_a23_mem/n19094 ), .CLK(clk), .RST(
        rst), .I(p_init[326]), .Q(\u_a23_mem/p_mem[40][6] ) );
  DFF \u_a23_mem/p_mem_reg[40][7]  ( .D(\u_a23_mem/n19093 ), .CLK(clk), .RST(
        rst), .I(p_init[327]), .Q(\u_a23_mem/p_mem[40][7] ) );
  DFF \u_a23_mem/p_mem_reg[41][0]  ( .D(\u_a23_mem/n19092 ), .CLK(clk), .RST(
        rst), .I(p_init[328]), .Q(\u_a23_mem/p_mem[41][0] ) );
  DFF \u_a23_mem/p_mem_reg[41][1]  ( .D(\u_a23_mem/n19091 ), .CLK(clk), .RST(
        rst), .I(p_init[329]), .Q(\u_a23_mem/p_mem[41][1] ) );
  DFF \u_a23_mem/p_mem_reg[41][2]  ( .D(\u_a23_mem/n19090 ), .CLK(clk), .RST(
        rst), .I(p_init[330]), .Q(\u_a23_mem/p_mem[41][2] ) );
  DFF \u_a23_mem/p_mem_reg[41][3]  ( .D(\u_a23_mem/n19089 ), .CLK(clk), .RST(
        rst), .I(p_init[331]), .Q(\u_a23_mem/p_mem[41][3] ) );
  DFF \u_a23_mem/p_mem_reg[41][4]  ( .D(\u_a23_mem/n19088 ), .CLK(clk), .RST(
        rst), .I(p_init[332]), .Q(\u_a23_mem/p_mem[41][4] ) );
  DFF \u_a23_mem/p_mem_reg[41][5]  ( .D(\u_a23_mem/n19087 ), .CLK(clk), .RST(
        rst), .I(p_init[333]), .Q(\u_a23_mem/p_mem[41][5] ) );
  DFF \u_a23_mem/p_mem_reg[41][6]  ( .D(\u_a23_mem/n19086 ), .CLK(clk), .RST(
        rst), .I(p_init[334]), .Q(\u_a23_mem/p_mem[41][6] ) );
  DFF \u_a23_mem/p_mem_reg[41][7]  ( .D(\u_a23_mem/n19085 ), .CLK(clk), .RST(
        rst), .I(p_init[335]), .Q(\u_a23_mem/p_mem[41][7] ) );
  DFF \u_a23_mem/p_mem_reg[42][0]  ( .D(\u_a23_mem/n19084 ), .CLK(clk), .RST(
        rst), .I(p_init[336]), .Q(\u_a23_mem/p_mem[42][0] ) );
  DFF \u_a23_mem/p_mem_reg[42][1]  ( .D(\u_a23_mem/n19083 ), .CLK(clk), .RST(
        rst), .I(p_init[337]), .Q(\u_a23_mem/p_mem[42][1] ) );
  DFF \u_a23_mem/p_mem_reg[42][2]  ( .D(\u_a23_mem/n19082 ), .CLK(clk), .RST(
        rst), .I(p_init[338]), .Q(\u_a23_mem/p_mem[42][2] ) );
  DFF \u_a23_mem/p_mem_reg[42][3]  ( .D(\u_a23_mem/n19081 ), .CLK(clk), .RST(
        rst), .I(p_init[339]), .Q(\u_a23_mem/p_mem[42][3] ) );
  DFF \u_a23_mem/p_mem_reg[42][4]  ( .D(\u_a23_mem/n19080 ), .CLK(clk), .RST(
        rst), .I(p_init[340]), .Q(\u_a23_mem/p_mem[42][4] ) );
  DFF \u_a23_mem/p_mem_reg[42][5]  ( .D(\u_a23_mem/n19079 ), .CLK(clk), .RST(
        rst), .I(p_init[341]), .Q(\u_a23_mem/p_mem[42][5] ) );
  DFF \u_a23_mem/p_mem_reg[42][6]  ( .D(\u_a23_mem/n19078 ), .CLK(clk), .RST(
        rst), .I(p_init[342]), .Q(\u_a23_mem/p_mem[42][6] ) );
  DFF \u_a23_mem/p_mem_reg[42][7]  ( .D(\u_a23_mem/n19077 ), .CLK(clk), .RST(
        rst), .I(p_init[343]), .Q(\u_a23_mem/p_mem[42][7] ) );
  DFF \u_a23_mem/p_mem_reg[43][0]  ( .D(\u_a23_mem/n19076 ), .CLK(clk), .RST(
        rst), .I(p_init[344]), .Q(\u_a23_mem/p_mem[43][0] ) );
  DFF \u_a23_mem/p_mem_reg[43][1]  ( .D(\u_a23_mem/n19075 ), .CLK(clk), .RST(
        rst), .I(p_init[345]), .Q(\u_a23_mem/p_mem[43][1] ) );
  DFF \u_a23_mem/p_mem_reg[43][2]  ( .D(\u_a23_mem/n19074 ), .CLK(clk), .RST(
        rst), .I(p_init[346]), .Q(\u_a23_mem/p_mem[43][2] ) );
  DFF \u_a23_mem/p_mem_reg[43][3]  ( .D(\u_a23_mem/n19073 ), .CLK(clk), .RST(
        rst), .I(p_init[347]), .Q(\u_a23_mem/p_mem[43][3] ) );
  DFF \u_a23_mem/p_mem_reg[43][4]  ( .D(\u_a23_mem/n19072 ), .CLK(clk), .RST(
        rst), .I(p_init[348]), .Q(\u_a23_mem/p_mem[43][4] ) );
  DFF \u_a23_mem/p_mem_reg[43][5]  ( .D(\u_a23_mem/n19071 ), .CLK(clk), .RST(
        rst), .I(p_init[349]), .Q(\u_a23_mem/p_mem[43][5] ) );
  DFF \u_a23_mem/p_mem_reg[43][6]  ( .D(\u_a23_mem/n19070 ), .CLK(clk), .RST(
        rst), .I(p_init[350]), .Q(\u_a23_mem/p_mem[43][6] ) );
  DFF \u_a23_mem/p_mem_reg[43][7]  ( .D(\u_a23_mem/n19069 ), .CLK(clk), .RST(
        rst), .I(p_init[351]), .Q(\u_a23_mem/p_mem[43][7] ) );
  DFF \u_a23_mem/p_mem_reg[44][0]  ( .D(\u_a23_mem/n19068 ), .CLK(clk), .RST(
        rst), .I(p_init[352]), .Q(\u_a23_mem/p_mem[44][0] ) );
  DFF \u_a23_mem/p_mem_reg[44][1]  ( .D(\u_a23_mem/n19067 ), .CLK(clk), .RST(
        rst), .I(p_init[353]), .Q(\u_a23_mem/p_mem[44][1] ) );
  DFF \u_a23_mem/p_mem_reg[44][2]  ( .D(\u_a23_mem/n19066 ), .CLK(clk), .RST(
        rst), .I(p_init[354]), .Q(\u_a23_mem/p_mem[44][2] ) );
  DFF \u_a23_mem/p_mem_reg[44][3]  ( .D(\u_a23_mem/n19065 ), .CLK(clk), .RST(
        rst), .I(p_init[355]), .Q(\u_a23_mem/p_mem[44][3] ) );
  DFF \u_a23_mem/p_mem_reg[44][4]  ( .D(\u_a23_mem/n19064 ), .CLK(clk), .RST(
        rst), .I(p_init[356]), .Q(\u_a23_mem/p_mem[44][4] ) );
  DFF \u_a23_mem/p_mem_reg[44][5]  ( .D(\u_a23_mem/n19063 ), .CLK(clk), .RST(
        rst), .I(p_init[357]), .Q(\u_a23_mem/p_mem[44][5] ) );
  DFF \u_a23_mem/p_mem_reg[44][6]  ( .D(\u_a23_mem/n19062 ), .CLK(clk), .RST(
        rst), .I(p_init[358]), .Q(\u_a23_mem/p_mem[44][6] ) );
  DFF \u_a23_mem/p_mem_reg[44][7]  ( .D(\u_a23_mem/n19061 ), .CLK(clk), .RST(
        rst), .I(p_init[359]), .Q(\u_a23_mem/p_mem[44][7] ) );
  DFF \u_a23_mem/p_mem_reg[45][0]  ( .D(\u_a23_mem/n19060 ), .CLK(clk), .RST(
        rst), .I(p_init[360]), .Q(\u_a23_mem/p_mem[45][0] ) );
  DFF \u_a23_mem/p_mem_reg[45][1]  ( .D(\u_a23_mem/n19059 ), .CLK(clk), .RST(
        rst), .I(p_init[361]), .Q(\u_a23_mem/p_mem[45][1] ) );
  DFF \u_a23_mem/p_mem_reg[45][2]  ( .D(\u_a23_mem/n19058 ), .CLK(clk), .RST(
        rst), .I(p_init[362]), .Q(\u_a23_mem/p_mem[45][2] ) );
  DFF \u_a23_mem/p_mem_reg[45][3]  ( .D(\u_a23_mem/n19057 ), .CLK(clk), .RST(
        rst), .I(p_init[363]), .Q(\u_a23_mem/p_mem[45][3] ) );
  DFF \u_a23_mem/p_mem_reg[45][4]  ( .D(\u_a23_mem/n19056 ), .CLK(clk), .RST(
        rst), .I(p_init[364]), .Q(\u_a23_mem/p_mem[45][4] ) );
  DFF \u_a23_mem/p_mem_reg[45][5]  ( .D(\u_a23_mem/n19055 ), .CLK(clk), .RST(
        rst), .I(p_init[365]), .Q(\u_a23_mem/p_mem[45][5] ) );
  DFF \u_a23_mem/p_mem_reg[45][6]  ( .D(\u_a23_mem/n19054 ), .CLK(clk), .RST(
        rst), .I(p_init[366]), .Q(\u_a23_mem/p_mem[45][6] ) );
  DFF \u_a23_mem/p_mem_reg[45][7]  ( .D(\u_a23_mem/n19053 ), .CLK(clk), .RST(
        rst), .I(p_init[367]), .Q(\u_a23_mem/p_mem[45][7] ) );
  DFF \u_a23_mem/p_mem_reg[46][0]  ( .D(\u_a23_mem/n19052 ), .CLK(clk), .RST(
        rst), .I(p_init[368]), .Q(\u_a23_mem/p_mem[46][0] ) );
  DFF \u_a23_mem/p_mem_reg[46][1]  ( .D(\u_a23_mem/n19051 ), .CLK(clk), .RST(
        rst), .I(p_init[369]), .Q(\u_a23_mem/p_mem[46][1] ) );
  DFF \u_a23_mem/p_mem_reg[46][2]  ( .D(\u_a23_mem/n19050 ), .CLK(clk), .RST(
        rst), .I(p_init[370]), .Q(\u_a23_mem/p_mem[46][2] ) );
  DFF \u_a23_mem/p_mem_reg[46][3]  ( .D(\u_a23_mem/n19049 ), .CLK(clk), .RST(
        rst), .I(p_init[371]), .Q(\u_a23_mem/p_mem[46][3] ) );
  DFF \u_a23_mem/p_mem_reg[46][4]  ( .D(\u_a23_mem/n19048 ), .CLK(clk), .RST(
        rst), .I(p_init[372]), .Q(\u_a23_mem/p_mem[46][4] ) );
  DFF \u_a23_mem/p_mem_reg[46][5]  ( .D(\u_a23_mem/n19047 ), .CLK(clk), .RST(
        rst), .I(p_init[373]), .Q(\u_a23_mem/p_mem[46][5] ) );
  DFF \u_a23_mem/p_mem_reg[46][6]  ( .D(\u_a23_mem/n19046 ), .CLK(clk), .RST(
        rst), .I(p_init[374]), .Q(\u_a23_mem/p_mem[46][6] ) );
  DFF \u_a23_mem/p_mem_reg[46][7]  ( .D(\u_a23_mem/n19045 ), .CLK(clk), .RST(
        rst), .I(p_init[375]), .Q(\u_a23_mem/p_mem[46][7] ) );
  DFF \u_a23_mem/p_mem_reg[47][0]  ( .D(\u_a23_mem/n19044 ), .CLK(clk), .RST(
        rst), .I(p_init[376]), .Q(\u_a23_mem/p_mem[47][0] ) );
  DFF \u_a23_mem/p_mem_reg[47][1]  ( .D(\u_a23_mem/n19043 ), .CLK(clk), .RST(
        rst), .I(p_init[377]), .Q(\u_a23_mem/p_mem[47][1] ) );
  DFF \u_a23_mem/p_mem_reg[47][2]  ( .D(\u_a23_mem/n19042 ), .CLK(clk), .RST(
        rst), .I(p_init[378]), .Q(\u_a23_mem/p_mem[47][2] ) );
  DFF \u_a23_mem/p_mem_reg[47][3]  ( .D(\u_a23_mem/n19041 ), .CLK(clk), .RST(
        rst), .I(p_init[379]), .Q(\u_a23_mem/p_mem[47][3] ) );
  DFF \u_a23_mem/p_mem_reg[47][4]  ( .D(\u_a23_mem/n19040 ), .CLK(clk), .RST(
        rst), .I(p_init[380]), .Q(\u_a23_mem/p_mem[47][4] ) );
  DFF \u_a23_mem/p_mem_reg[47][5]  ( .D(\u_a23_mem/n19039 ), .CLK(clk), .RST(
        rst), .I(p_init[381]), .Q(\u_a23_mem/p_mem[47][5] ) );
  DFF \u_a23_mem/p_mem_reg[47][6]  ( .D(\u_a23_mem/n19038 ), .CLK(clk), .RST(
        rst), .I(p_init[382]), .Q(\u_a23_mem/p_mem[47][6] ) );
  DFF \u_a23_mem/p_mem_reg[47][7]  ( .D(\u_a23_mem/n19037 ), .CLK(clk), .RST(
        rst), .I(p_init[383]), .Q(\u_a23_mem/p_mem[47][7] ) );
  DFF \u_a23_mem/p_mem_reg[48][0]  ( .D(\u_a23_mem/n19036 ), .CLK(clk), .RST(
        rst), .I(p_init[384]), .Q(\u_a23_mem/p_mem[48][0] ) );
  DFF \u_a23_mem/p_mem_reg[48][1]  ( .D(\u_a23_mem/n19035 ), .CLK(clk), .RST(
        rst), .I(p_init[385]), .Q(\u_a23_mem/p_mem[48][1] ) );
  DFF \u_a23_mem/p_mem_reg[48][2]  ( .D(\u_a23_mem/n19034 ), .CLK(clk), .RST(
        rst), .I(p_init[386]), .Q(\u_a23_mem/p_mem[48][2] ) );
  DFF \u_a23_mem/p_mem_reg[48][3]  ( .D(\u_a23_mem/n19033 ), .CLK(clk), .RST(
        rst), .I(p_init[387]), .Q(\u_a23_mem/p_mem[48][3] ) );
  DFF \u_a23_mem/p_mem_reg[48][4]  ( .D(\u_a23_mem/n19032 ), .CLK(clk), .RST(
        rst), .I(p_init[388]), .Q(\u_a23_mem/p_mem[48][4] ) );
  DFF \u_a23_mem/p_mem_reg[48][5]  ( .D(\u_a23_mem/n19031 ), .CLK(clk), .RST(
        rst), .I(p_init[389]), .Q(\u_a23_mem/p_mem[48][5] ) );
  DFF \u_a23_mem/p_mem_reg[48][6]  ( .D(\u_a23_mem/n19030 ), .CLK(clk), .RST(
        rst), .I(p_init[390]), .Q(\u_a23_mem/p_mem[48][6] ) );
  DFF \u_a23_mem/p_mem_reg[48][7]  ( .D(\u_a23_mem/n19029 ), .CLK(clk), .RST(
        rst), .I(p_init[391]), .Q(\u_a23_mem/p_mem[48][7] ) );
  DFF \u_a23_mem/p_mem_reg[49][0]  ( .D(\u_a23_mem/n19028 ), .CLK(clk), .RST(
        rst), .I(p_init[392]), .Q(\u_a23_mem/p_mem[49][0] ) );
  DFF \u_a23_mem/p_mem_reg[49][1]  ( .D(\u_a23_mem/n19027 ), .CLK(clk), .RST(
        rst), .I(p_init[393]), .Q(\u_a23_mem/p_mem[49][1] ) );
  DFF \u_a23_mem/p_mem_reg[49][2]  ( .D(\u_a23_mem/n19026 ), .CLK(clk), .RST(
        rst), .I(p_init[394]), .Q(\u_a23_mem/p_mem[49][2] ) );
  DFF \u_a23_mem/p_mem_reg[49][3]  ( .D(\u_a23_mem/n19025 ), .CLK(clk), .RST(
        rst), .I(p_init[395]), .Q(\u_a23_mem/p_mem[49][3] ) );
  DFF \u_a23_mem/p_mem_reg[49][4]  ( .D(\u_a23_mem/n19024 ), .CLK(clk), .RST(
        rst), .I(p_init[396]), .Q(\u_a23_mem/p_mem[49][4] ) );
  DFF \u_a23_mem/p_mem_reg[49][5]  ( .D(\u_a23_mem/n19023 ), .CLK(clk), .RST(
        rst), .I(p_init[397]), .Q(\u_a23_mem/p_mem[49][5] ) );
  DFF \u_a23_mem/p_mem_reg[49][6]  ( .D(\u_a23_mem/n19022 ), .CLK(clk), .RST(
        rst), .I(p_init[398]), .Q(\u_a23_mem/p_mem[49][6] ) );
  DFF \u_a23_mem/p_mem_reg[49][7]  ( .D(\u_a23_mem/n19021 ), .CLK(clk), .RST(
        rst), .I(p_init[399]), .Q(\u_a23_mem/p_mem[49][7] ) );
  DFF \u_a23_mem/p_mem_reg[50][0]  ( .D(\u_a23_mem/n19020 ), .CLK(clk), .RST(
        rst), .I(p_init[400]), .Q(\u_a23_mem/p_mem[50][0] ) );
  DFF \u_a23_mem/p_mem_reg[50][1]  ( .D(\u_a23_mem/n19019 ), .CLK(clk), .RST(
        rst), .I(p_init[401]), .Q(\u_a23_mem/p_mem[50][1] ) );
  DFF \u_a23_mem/p_mem_reg[50][2]  ( .D(\u_a23_mem/n19018 ), .CLK(clk), .RST(
        rst), .I(p_init[402]), .Q(\u_a23_mem/p_mem[50][2] ) );
  DFF \u_a23_mem/p_mem_reg[50][3]  ( .D(\u_a23_mem/n19017 ), .CLK(clk), .RST(
        rst), .I(p_init[403]), .Q(\u_a23_mem/p_mem[50][3] ) );
  DFF \u_a23_mem/p_mem_reg[50][4]  ( .D(\u_a23_mem/n19016 ), .CLK(clk), .RST(
        rst), .I(p_init[404]), .Q(\u_a23_mem/p_mem[50][4] ) );
  DFF \u_a23_mem/p_mem_reg[50][5]  ( .D(\u_a23_mem/n19015 ), .CLK(clk), .RST(
        rst), .I(p_init[405]), .Q(\u_a23_mem/p_mem[50][5] ) );
  DFF \u_a23_mem/p_mem_reg[50][6]  ( .D(\u_a23_mem/n19014 ), .CLK(clk), .RST(
        rst), .I(p_init[406]), .Q(\u_a23_mem/p_mem[50][6] ) );
  DFF \u_a23_mem/p_mem_reg[50][7]  ( .D(\u_a23_mem/n19013 ), .CLK(clk), .RST(
        rst), .I(p_init[407]), .Q(\u_a23_mem/p_mem[50][7] ) );
  DFF \u_a23_mem/p_mem_reg[51][0]  ( .D(\u_a23_mem/n19012 ), .CLK(clk), .RST(
        rst), .I(p_init[408]), .Q(\u_a23_mem/p_mem[51][0] ) );
  DFF \u_a23_mem/p_mem_reg[51][1]  ( .D(\u_a23_mem/n19011 ), .CLK(clk), .RST(
        rst), .I(p_init[409]), .Q(\u_a23_mem/p_mem[51][1] ) );
  DFF \u_a23_mem/p_mem_reg[51][2]  ( .D(\u_a23_mem/n19010 ), .CLK(clk), .RST(
        rst), .I(p_init[410]), .Q(\u_a23_mem/p_mem[51][2] ) );
  DFF \u_a23_mem/p_mem_reg[51][3]  ( .D(\u_a23_mem/n19009 ), .CLK(clk), .RST(
        rst), .I(p_init[411]), .Q(\u_a23_mem/p_mem[51][3] ) );
  DFF \u_a23_mem/p_mem_reg[51][4]  ( .D(\u_a23_mem/n19008 ), .CLK(clk), .RST(
        rst), .I(p_init[412]), .Q(\u_a23_mem/p_mem[51][4] ) );
  DFF \u_a23_mem/p_mem_reg[51][5]  ( .D(\u_a23_mem/n19007 ), .CLK(clk), .RST(
        rst), .I(p_init[413]), .Q(\u_a23_mem/p_mem[51][5] ) );
  DFF \u_a23_mem/p_mem_reg[51][6]  ( .D(\u_a23_mem/n19006 ), .CLK(clk), .RST(
        rst), .I(p_init[414]), .Q(\u_a23_mem/p_mem[51][6] ) );
  DFF \u_a23_mem/p_mem_reg[51][7]  ( .D(\u_a23_mem/n19005 ), .CLK(clk), .RST(
        rst), .I(p_init[415]), .Q(\u_a23_mem/p_mem[51][7] ) );
  DFF \u_a23_mem/p_mem_reg[52][0]  ( .D(\u_a23_mem/n19004 ), .CLK(clk), .RST(
        rst), .I(p_init[416]), .Q(\u_a23_mem/p_mem[52][0] ) );
  DFF \u_a23_mem/p_mem_reg[52][1]  ( .D(\u_a23_mem/n19003 ), .CLK(clk), .RST(
        rst), .I(p_init[417]), .Q(\u_a23_mem/p_mem[52][1] ) );
  DFF \u_a23_mem/p_mem_reg[52][2]  ( .D(\u_a23_mem/n19002 ), .CLK(clk), .RST(
        rst), .I(p_init[418]), .Q(\u_a23_mem/p_mem[52][2] ) );
  DFF \u_a23_mem/p_mem_reg[52][3]  ( .D(\u_a23_mem/n19001 ), .CLK(clk), .RST(
        rst), .I(p_init[419]), .Q(\u_a23_mem/p_mem[52][3] ) );
  DFF \u_a23_mem/p_mem_reg[52][4]  ( .D(\u_a23_mem/n19000 ), .CLK(clk), .RST(
        rst), .I(p_init[420]), .Q(\u_a23_mem/p_mem[52][4] ) );
  DFF \u_a23_mem/p_mem_reg[52][5]  ( .D(\u_a23_mem/n18999 ), .CLK(clk), .RST(
        rst), .I(p_init[421]), .Q(\u_a23_mem/p_mem[52][5] ) );
  DFF \u_a23_mem/p_mem_reg[52][6]  ( .D(\u_a23_mem/n18998 ), .CLK(clk), .RST(
        rst), .I(p_init[422]), .Q(\u_a23_mem/p_mem[52][6] ) );
  DFF \u_a23_mem/p_mem_reg[52][7]  ( .D(\u_a23_mem/n18997 ), .CLK(clk), .RST(
        rst), .I(p_init[423]), .Q(\u_a23_mem/p_mem[52][7] ) );
  DFF \u_a23_mem/p_mem_reg[53][0]  ( .D(\u_a23_mem/n18996 ), .CLK(clk), .RST(
        rst), .I(p_init[424]), .Q(\u_a23_mem/p_mem[53][0] ) );
  DFF \u_a23_mem/p_mem_reg[53][1]  ( .D(\u_a23_mem/n18995 ), .CLK(clk), .RST(
        rst), .I(p_init[425]), .Q(\u_a23_mem/p_mem[53][1] ) );
  DFF \u_a23_mem/p_mem_reg[53][2]  ( .D(\u_a23_mem/n18994 ), .CLK(clk), .RST(
        rst), .I(p_init[426]), .Q(\u_a23_mem/p_mem[53][2] ) );
  DFF \u_a23_mem/p_mem_reg[53][3]  ( .D(\u_a23_mem/n18993 ), .CLK(clk), .RST(
        rst), .I(p_init[427]), .Q(\u_a23_mem/p_mem[53][3] ) );
  DFF \u_a23_mem/p_mem_reg[53][4]  ( .D(\u_a23_mem/n18992 ), .CLK(clk), .RST(
        rst), .I(p_init[428]), .Q(\u_a23_mem/p_mem[53][4] ) );
  DFF \u_a23_mem/p_mem_reg[53][5]  ( .D(\u_a23_mem/n18991 ), .CLK(clk), .RST(
        rst), .I(p_init[429]), .Q(\u_a23_mem/p_mem[53][5] ) );
  DFF \u_a23_mem/p_mem_reg[53][6]  ( .D(\u_a23_mem/n18990 ), .CLK(clk), .RST(
        rst), .I(p_init[430]), .Q(\u_a23_mem/p_mem[53][6] ) );
  DFF \u_a23_mem/p_mem_reg[53][7]  ( .D(\u_a23_mem/n18989 ), .CLK(clk), .RST(
        rst), .I(p_init[431]), .Q(\u_a23_mem/p_mem[53][7] ) );
  DFF \u_a23_mem/p_mem_reg[54][0]  ( .D(\u_a23_mem/n18988 ), .CLK(clk), .RST(
        rst), .I(p_init[432]), .Q(\u_a23_mem/p_mem[54][0] ) );
  DFF \u_a23_mem/p_mem_reg[54][1]  ( .D(\u_a23_mem/n18987 ), .CLK(clk), .RST(
        rst), .I(p_init[433]), .Q(\u_a23_mem/p_mem[54][1] ) );
  DFF \u_a23_mem/p_mem_reg[54][2]  ( .D(\u_a23_mem/n18986 ), .CLK(clk), .RST(
        rst), .I(p_init[434]), .Q(\u_a23_mem/p_mem[54][2] ) );
  DFF \u_a23_mem/p_mem_reg[54][3]  ( .D(\u_a23_mem/n18985 ), .CLK(clk), .RST(
        rst), .I(p_init[435]), .Q(\u_a23_mem/p_mem[54][3] ) );
  DFF \u_a23_mem/p_mem_reg[54][4]  ( .D(\u_a23_mem/n18984 ), .CLK(clk), .RST(
        rst), .I(p_init[436]), .Q(\u_a23_mem/p_mem[54][4] ) );
  DFF \u_a23_mem/p_mem_reg[54][5]  ( .D(\u_a23_mem/n18983 ), .CLK(clk), .RST(
        rst), .I(p_init[437]), .Q(\u_a23_mem/p_mem[54][5] ) );
  DFF \u_a23_mem/p_mem_reg[54][6]  ( .D(\u_a23_mem/n18982 ), .CLK(clk), .RST(
        rst), .I(p_init[438]), .Q(\u_a23_mem/p_mem[54][6] ) );
  DFF \u_a23_mem/p_mem_reg[54][7]  ( .D(\u_a23_mem/n18981 ), .CLK(clk), .RST(
        rst), .I(p_init[439]), .Q(\u_a23_mem/p_mem[54][7] ) );
  DFF \u_a23_mem/p_mem_reg[55][0]  ( .D(\u_a23_mem/n18980 ), .CLK(clk), .RST(
        rst), .I(p_init[440]), .Q(\u_a23_mem/p_mem[55][0] ) );
  DFF \u_a23_mem/p_mem_reg[55][1]  ( .D(\u_a23_mem/n18979 ), .CLK(clk), .RST(
        rst), .I(p_init[441]), .Q(\u_a23_mem/p_mem[55][1] ) );
  DFF \u_a23_mem/p_mem_reg[55][2]  ( .D(\u_a23_mem/n18978 ), .CLK(clk), .RST(
        rst), .I(p_init[442]), .Q(\u_a23_mem/p_mem[55][2] ) );
  DFF \u_a23_mem/p_mem_reg[55][3]  ( .D(\u_a23_mem/n18977 ), .CLK(clk), .RST(
        rst), .I(p_init[443]), .Q(\u_a23_mem/p_mem[55][3] ) );
  DFF \u_a23_mem/p_mem_reg[55][4]  ( .D(\u_a23_mem/n18976 ), .CLK(clk), .RST(
        rst), .I(p_init[444]), .Q(\u_a23_mem/p_mem[55][4] ) );
  DFF \u_a23_mem/p_mem_reg[55][5]  ( .D(\u_a23_mem/n18975 ), .CLK(clk), .RST(
        rst), .I(p_init[445]), .Q(\u_a23_mem/p_mem[55][5] ) );
  DFF \u_a23_mem/p_mem_reg[55][6]  ( .D(\u_a23_mem/n18974 ), .CLK(clk), .RST(
        rst), .I(p_init[446]), .Q(\u_a23_mem/p_mem[55][6] ) );
  DFF \u_a23_mem/p_mem_reg[55][7]  ( .D(\u_a23_mem/n18973 ), .CLK(clk), .RST(
        rst), .I(p_init[447]), .Q(\u_a23_mem/p_mem[55][7] ) );
  DFF \u_a23_mem/p_mem_reg[56][0]  ( .D(\u_a23_mem/n18972 ), .CLK(clk), .RST(
        rst), .I(p_init[448]), .Q(\u_a23_mem/p_mem[56][0] ) );
  DFF \u_a23_mem/p_mem_reg[56][1]  ( .D(\u_a23_mem/n18971 ), .CLK(clk), .RST(
        rst), .I(p_init[449]), .Q(\u_a23_mem/p_mem[56][1] ) );
  DFF \u_a23_mem/p_mem_reg[56][2]  ( .D(\u_a23_mem/n18970 ), .CLK(clk), .RST(
        rst), .I(p_init[450]), .Q(\u_a23_mem/p_mem[56][2] ) );
  DFF \u_a23_mem/p_mem_reg[56][3]  ( .D(\u_a23_mem/n18969 ), .CLK(clk), .RST(
        rst), .I(p_init[451]), .Q(\u_a23_mem/p_mem[56][3] ) );
  DFF \u_a23_mem/p_mem_reg[56][4]  ( .D(\u_a23_mem/n18968 ), .CLK(clk), .RST(
        rst), .I(p_init[452]), .Q(\u_a23_mem/p_mem[56][4] ) );
  DFF \u_a23_mem/p_mem_reg[56][5]  ( .D(\u_a23_mem/n18967 ), .CLK(clk), .RST(
        rst), .I(p_init[453]), .Q(\u_a23_mem/p_mem[56][5] ) );
  DFF \u_a23_mem/p_mem_reg[56][6]  ( .D(\u_a23_mem/n18966 ), .CLK(clk), .RST(
        rst), .I(p_init[454]), .Q(\u_a23_mem/p_mem[56][6] ) );
  DFF \u_a23_mem/p_mem_reg[56][7]  ( .D(\u_a23_mem/n18965 ), .CLK(clk), .RST(
        rst), .I(p_init[455]), .Q(\u_a23_mem/p_mem[56][7] ) );
  DFF \u_a23_mem/p_mem_reg[57][0]  ( .D(\u_a23_mem/n18964 ), .CLK(clk), .RST(
        rst), .I(p_init[456]), .Q(\u_a23_mem/p_mem[57][0] ) );
  DFF \u_a23_mem/p_mem_reg[57][1]  ( .D(\u_a23_mem/n18963 ), .CLK(clk), .RST(
        rst), .I(p_init[457]), .Q(\u_a23_mem/p_mem[57][1] ) );
  DFF \u_a23_mem/p_mem_reg[57][2]  ( .D(\u_a23_mem/n18962 ), .CLK(clk), .RST(
        rst), .I(p_init[458]), .Q(\u_a23_mem/p_mem[57][2] ) );
  DFF \u_a23_mem/p_mem_reg[57][3]  ( .D(\u_a23_mem/n18961 ), .CLK(clk), .RST(
        rst), .I(p_init[459]), .Q(\u_a23_mem/p_mem[57][3] ) );
  DFF \u_a23_mem/p_mem_reg[57][4]  ( .D(\u_a23_mem/n18960 ), .CLK(clk), .RST(
        rst), .I(p_init[460]), .Q(\u_a23_mem/p_mem[57][4] ) );
  DFF \u_a23_mem/p_mem_reg[57][5]  ( .D(\u_a23_mem/n18959 ), .CLK(clk), .RST(
        rst), .I(p_init[461]), .Q(\u_a23_mem/p_mem[57][5] ) );
  DFF \u_a23_mem/p_mem_reg[57][6]  ( .D(\u_a23_mem/n18958 ), .CLK(clk), .RST(
        rst), .I(p_init[462]), .Q(\u_a23_mem/p_mem[57][6] ) );
  DFF \u_a23_mem/p_mem_reg[57][7]  ( .D(\u_a23_mem/n18957 ), .CLK(clk), .RST(
        rst), .I(p_init[463]), .Q(\u_a23_mem/p_mem[57][7] ) );
  DFF \u_a23_mem/p_mem_reg[58][0]  ( .D(\u_a23_mem/n18956 ), .CLK(clk), .RST(
        rst), .I(p_init[464]), .Q(\u_a23_mem/p_mem[58][0] ) );
  DFF \u_a23_mem/p_mem_reg[58][1]  ( .D(\u_a23_mem/n18955 ), .CLK(clk), .RST(
        rst), .I(p_init[465]), .Q(\u_a23_mem/p_mem[58][1] ) );
  DFF \u_a23_mem/p_mem_reg[58][2]  ( .D(\u_a23_mem/n18954 ), .CLK(clk), .RST(
        rst), .I(p_init[466]), .Q(\u_a23_mem/p_mem[58][2] ) );
  DFF \u_a23_mem/p_mem_reg[58][3]  ( .D(\u_a23_mem/n18953 ), .CLK(clk), .RST(
        rst), .I(p_init[467]), .Q(\u_a23_mem/p_mem[58][3] ) );
  DFF \u_a23_mem/p_mem_reg[58][4]  ( .D(\u_a23_mem/n18952 ), .CLK(clk), .RST(
        rst), .I(p_init[468]), .Q(\u_a23_mem/p_mem[58][4] ) );
  DFF \u_a23_mem/p_mem_reg[58][5]  ( .D(\u_a23_mem/n18951 ), .CLK(clk), .RST(
        rst), .I(p_init[469]), .Q(\u_a23_mem/p_mem[58][5] ) );
  DFF \u_a23_mem/p_mem_reg[58][6]  ( .D(\u_a23_mem/n18950 ), .CLK(clk), .RST(
        rst), .I(p_init[470]), .Q(\u_a23_mem/p_mem[58][6] ) );
  DFF \u_a23_mem/p_mem_reg[58][7]  ( .D(\u_a23_mem/n18949 ), .CLK(clk), .RST(
        rst), .I(p_init[471]), .Q(\u_a23_mem/p_mem[58][7] ) );
  DFF \u_a23_mem/p_mem_reg[59][0]  ( .D(\u_a23_mem/n18948 ), .CLK(clk), .RST(
        rst), .I(p_init[472]), .Q(\u_a23_mem/p_mem[59][0] ) );
  DFF \u_a23_mem/p_mem_reg[59][1]  ( .D(\u_a23_mem/n18947 ), .CLK(clk), .RST(
        rst), .I(p_init[473]), .Q(\u_a23_mem/p_mem[59][1] ) );
  DFF \u_a23_mem/p_mem_reg[59][2]  ( .D(\u_a23_mem/n18946 ), .CLK(clk), .RST(
        rst), .I(p_init[474]), .Q(\u_a23_mem/p_mem[59][2] ) );
  DFF \u_a23_mem/p_mem_reg[59][3]  ( .D(\u_a23_mem/n18945 ), .CLK(clk), .RST(
        rst), .I(p_init[475]), .Q(\u_a23_mem/p_mem[59][3] ) );
  DFF \u_a23_mem/p_mem_reg[59][4]  ( .D(\u_a23_mem/n18944 ), .CLK(clk), .RST(
        rst), .I(p_init[476]), .Q(\u_a23_mem/p_mem[59][4] ) );
  DFF \u_a23_mem/p_mem_reg[59][5]  ( .D(\u_a23_mem/n18943 ), .CLK(clk), .RST(
        rst), .I(p_init[477]), .Q(\u_a23_mem/p_mem[59][5] ) );
  DFF \u_a23_mem/p_mem_reg[59][6]  ( .D(\u_a23_mem/n18942 ), .CLK(clk), .RST(
        rst), .I(p_init[478]), .Q(\u_a23_mem/p_mem[59][6] ) );
  DFF \u_a23_mem/p_mem_reg[59][7]  ( .D(\u_a23_mem/n18941 ), .CLK(clk), .RST(
        rst), .I(p_init[479]), .Q(\u_a23_mem/p_mem[59][7] ) );
  DFF \u_a23_mem/p_mem_reg[60][0]  ( .D(\u_a23_mem/n18940 ), .CLK(clk), .RST(
        rst), .I(p_init[480]), .Q(\u_a23_mem/p_mem[60][0] ) );
  DFF \u_a23_mem/p_mem_reg[60][1]  ( .D(\u_a23_mem/n18939 ), .CLK(clk), .RST(
        rst), .I(p_init[481]), .Q(\u_a23_mem/p_mem[60][1] ) );
  DFF \u_a23_mem/p_mem_reg[60][2]  ( .D(\u_a23_mem/n18938 ), .CLK(clk), .RST(
        rst), .I(p_init[482]), .Q(\u_a23_mem/p_mem[60][2] ) );
  DFF \u_a23_mem/p_mem_reg[60][3]  ( .D(\u_a23_mem/n18937 ), .CLK(clk), .RST(
        rst), .I(p_init[483]), .Q(\u_a23_mem/p_mem[60][3] ) );
  DFF \u_a23_mem/p_mem_reg[60][4]  ( .D(\u_a23_mem/n18936 ), .CLK(clk), .RST(
        rst), .I(p_init[484]), .Q(\u_a23_mem/p_mem[60][4] ) );
  DFF \u_a23_mem/p_mem_reg[60][5]  ( .D(\u_a23_mem/n18935 ), .CLK(clk), .RST(
        rst), .I(p_init[485]), .Q(\u_a23_mem/p_mem[60][5] ) );
  DFF \u_a23_mem/p_mem_reg[60][6]  ( .D(\u_a23_mem/n18934 ), .CLK(clk), .RST(
        rst), .I(p_init[486]), .Q(\u_a23_mem/p_mem[60][6] ) );
  DFF \u_a23_mem/p_mem_reg[60][7]  ( .D(\u_a23_mem/n18933 ), .CLK(clk), .RST(
        rst), .I(p_init[487]), .Q(\u_a23_mem/p_mem[60][7] ) );
  DFF \u_a23_mem/p_mem_reg[61][0]  ( .D(\u_a23_mem/n18932 ), .CLK(clk), .RST(
        rst), .I(p_init[488]), .Q(\u_a23_mem/p_mem[61][0] ) );
  DFF \u_a23_mem/p_mem_reg[61][1]  ( .D(\u_a23_mem/n18931 ), .CLK(clk), .RST(
        rst), .I(p_init[489]), .Q(\u_a23_mem/p_mem[61][1] ) );
  DFF \u_a23_mem/p_mem_reg[61][2]  ( .D(\u_a23_mem/n18930 ), .CLK(clk), .RST(
        rst), .I(p_init[490]), .Q(\u_a23_mem/p_mem[61][2] ) );
  DFF \u_a23_mem/p_mem_reg[61][3]  ( .D(\u_a23_mem/n18929 ), .CLK(clk), .RST(
        rst), .I(p_init[491]), .Q(\u_a23_mem/p_mem[61][3] ) );
  DFF \u_a23_mem/p_mem_reg[61][4]  ( .D(\u_a23_mem/n18928 ), .CLK(clk), .RST(
        rst), .I(p_init[492]), .Q(\u_a23_mem/p_mem[61][4] ) );
  DFF \u_a23_mem/p_mem_reg[61][5]  ( .D(\u_a23_mem/n18927 ), .CLK(clk), .RST(
        rst), .I(p_init[493]), .Q(\u_a23_mem/p_mem[61][5] ) );
  DFF \u_a23_mem/p_mem_reg[61][6]  ( .D(\u_a23_mem/n18926 ), .CLK(clk), .RST(
        rst), .I(p_init[494]), .Q(\u_a23_mem/p_mem[61][6] ) );
  DFF \u_a23_mem/p_mem_reg[61][7]  ( .D(\u_a23_mem/n18925 ), .CLK(clk), .RST(
        rst), .I(p_init[495]), .Q(\u_a23_mem/p_mem[61][7] ) );
  DFF \u_a23_mem/p_mem_reg[62][0]  ( .D(\u_a23_mem/n18924 ), .CLK(clk), .RST(
        rst), .I(p_init[496]), .Q(\u_a23_mem/p_mem[62][0] ) );
  DFF \u_a23_mem/p_mem_reg[62][1]  ( .D(\u_a23_mem/n18923 ), .CLK(clk), .RST(
        rst), .I(p_init[497]), .Q(\u_a23_mem/p_mem[62][1] ) );
  DFF \u_a23_mem/p_mem_reg[62][2]  ( .D(\u_a23_mem/n18922 ), .CLK(clk), .RST(
        rst), .I(p_init[498]), .Q(\u_a23_mem/p_mem[62][2] ) );
  DFF \u_a23_mem/p_mem_reg[62][3]  ( .D(\u_a23_mem/n18921 ), .CLK(clk), .RST(
        rst), .I(p_init[499]), .Q(\u_a23_mem/p_mem[62][3] ) );
  DFF \u_a23_mem/p_mem_reg[62][4]  ( .D(\u_a23_mem/n18920 ), .CLK(clk), .RST(
        rst), .I(p_init[500]), .Q(\u_a23_mem/p_mem[62][4] ) );
  DFF \u_a23_mem/p_mem_reg[62][5]  ( .D(\u_a23_mem/n18919 ), .CLK(clk), .RST(
        rst), .I(p_init[501]), .Q(\u_a23_mem/p_mem[62][5] ) );
  DFF \u_a23_mem/p_mem_reg[62][6]  ( .D(\u_a23_mem/n18918 ), .CLK(clk), .RST(
        rst), .I(p_init[502]), .Q(\u_a23_mem/p_mem[62][6] ) );
  DFF \u_a23_mem/p_mem_reg[62][7]  ( .D(\u_a23_mem/n18917 ), .CLK(clk), .RST(
        rst), .I(p_init[503]), .Q(\u_a23_mem/p_mem[62][7] ) );
  DFF \u_a23_mem/p_mem_reg[63][0]  ( .D(\u_a23_mem/n18916 ), .CLK(clk), .RST(
        rst), .I(p_init[504]), .Q(\u_a23_mem/p_mem[63][0] ) );
  DFF \u_a23_mem/p_mem_reg[63][1]  ( .D(\u_a23_mem/n18915 ), .CLK(clk), .RST(
        rst), .I(p_init[505]), .Q(\u_a23_mem/p_mem[63][1] ) );
  DFF \u_a23_mem/p_mem_reg[63][2]  ( .D(\u_a23_mem/n18914 ), .CLK(clk), .RST(
        rst), .I(p_init[506]), .Q(\u_a23_mem/p_mem[63][2] ) );
  DFF \u_a23_mem/p_mem_reg[63][3]  ( .D(\u_a23_mem/n18913 ), .CLK(clk), .RST(
        rst), .I(p_init[507]), .Q(\u_a23_mem/p_mem[63][3] ) );
  DFF \u_a23_mem/p_mem_reg[63][4]  ( .D(\u_a23_mem/n18912 ), .CLK(clk), .RST(
        rst), .I(p_init[508]), .Q(\u_a23_mem/p_mem[63][4] ) );
  DFF \u_a23_mem/p_mem_reg[63][5]  ( .D(\u_a23_mem/n18911 ), .CLK(clk), .RST(
        rst), .I(p_init[509]), .Q(\u_a23_mem/p_mem[63][5] ) );
  DFF \u_a23_mem/p_mem_reg[63][6]  ( .D(\u_a23_mem/n18910 ), .CLK(clk), .RST(
        rst), .I(p_init[510]), .Q(\u_a23_mem/p_mem[63][6] ) );
  DFF \u_a23_mem/p_mem_reg[63][7]  ( .D(\u_a23_mem/n18909 ), .CLK(clk), .RST(
        rst), .I(p_init[511]), .Q(\u_a23_mem/p_mem[63][7] ) );
  DFF \u_a23_mem/p_mem_reg[64][0]  ( .D(\u_a23_mem/n18908 ), .CLK(clk), .RST(
        rst), .I(p_init[512]), .Q(\u_a23_mem/p_mem[64][0] ) );
  DFF \u_a23_mem/p_mem_reg[64][1]  ( .D(\u_a23_mem/n18907 ), .CLK(clk), .RST(
        rst), .I(p_init[513]), .Q(\u_a23_mem/p_mem[64][1] ) );
  DFF \u_a23_mem/p_mem_reg[64][2]  ( .D(\u_a23_mem/n18906 ), .CLK(clk), .RST(
        rst), .I(p_init[514]), .Q(\u_a23_mem/p_mem[64][2] ) );
  DFF \u_a23_mem/p_mem_reg[64][3]  ( .D(\u_a23_mem/n18905 ), .CLK(clk), .RST(
        rst), .I(p_init[515]), .Q(\u_a23_mem/p_mem[64][3] ) );
  DFF \u_a23_mem/p_mem_reg[64][4]  ( .D(\u_a23_mem/n18904 ), .CLK(clk), .RST(
        rst), .I(p_init[516]), .Q(\u_a23_mem/p_mem[64][4] ) );
  DFF \u_a23_mem/p_mem_reg[64][5]  ( .D(\u_a23_mem/n18903 ), .CLK(clk), .RST(
        rst), .I(p_init[517]), .Q(\u_a23_mem/p_mem[64][5] ) );
  DFF \u_a23_mem/p_mem_reg[64][6]  ( .D(\u_a23_mem/n18902 ), .CLK(clk), .RST(
        rst), .I(p_init[518]), .Q(\u_a23_mem/p_mem[64][6] ) );
  DFF \u_a23_mem/p_mem_reg[64][7]  ( .D(\u_a23_mem/n18901 ), .CLK(clk), .RST(
        rst), .I(p_init[519]), .Q(\u_a23_mem/p_mem[64][7] ) );
  DFF \u_a23_mem/p_mem_reg[65][0]  ( .D(\u_a23_mem/n18900 ), .CLK(clk), .RST(
        rst), .I(p_init[520]), .Q(\u_a23_mem/p_mem[65][0] ) );
  DFF \u_a23_mem/p_mem_reg[65][1]  ( .D(\u_a23_mem/n18899 ), .CLK(clk), .RST(
        rst), .I(p_init[521]), .Q(\u_a23_mem/p_mem[65][1] ) );
  DFF \u_a23_mem/p_mem_reg[65][2]  ( .D(\u_a23_mem/n18898 ), .CLK(clk), .RST(
        rst), .I(p_init[522]), .Q(\u_a23_mem/p_mem[65][2] ) );
  DFF \u_a23_mem/p_mem_reg[65][3]  ( .D(\u_a23_mem/n18897 ), .CLK(clk), .RST(
        rst), .I(p_init[523]), .Q(\u_a23_mem/p_mem[65][3] ) );
  DFF \u_a23_mem/p_mem_reg[65][4]  ( .D(\u_a23_mem/n18896 ), .CLK(clk), .RST(
        rst), .I(p_init[524]), .Q(\u_a23_mem/p_mem[65][4] ) );
  DFF \u_a23_mem/p_mem_reg[65][5]  ( .D(\u_a23_mem/n18895 ), .CLK(clk), .RST(
        rst), .I(p_init[525]), .Q(\u_a23_mem/p_mem[65][5] ) );
  DFF \u_a23_mem/p_mem_reg[65][6]  ( .D(\u_a23_mem/n18894 ), .CLK(clk), .RST(
        rst), .I(p_init[526]), .Q(\u_a23_mem/p_mem[65][6] ) );
  DFF \u_a23_mem/p_mem_reg[65][7]  ( .D(\u_a23_mem/n18893 ), .CLK(clk), .RST(
        rst), .I(p_init[527]), .Q(\u_a23_mem/p_mem[65][7] ) );
  DFF \u_a23_mem/p_mem_reg[66][0]  ( .D(\u_a23_mem/n18892 ), .CLK(clk), .RST(
        rst), .I(p_init[528]), .Q(\u_a23_mem/p_mem[66][0] ) );
  DFF \u_a23_mem/p_mem_reg[66][1]  ( .D(\u_a23_mem/n18891 ), .CLK(clk), .RST(
        rst), .I(p_init[529]), .Q(\u_a23_mem/p_mem[66][1] ) );
  DFF \u_a23_mem/p_mem_reg[66][2]  ( .D(\u_a23_mem/n18890 ), .CLK(clk), .RST(
        rst), .I(p_init[530]), .Q(\u_a23_mem/p_mem[66][2] ) );
  DFF \u_a23_mem/p_mem_reg[66][3]  ( .D(\u_a23_mem/n18889 ), .CLK(clk), .RST(
        rst), .I(p_init[531]), .Q(\u_a23_mem/p_mem[66][3] ) );
  DFF \u_a23_mem/p_mem_reg[66][4]  ( .D(\u_a23_mem/n18888 ), .CLK(clk), .RST(
        rst), .I(p_init[532]), .Q(\u_a23_mem/p_mem[66][4] ) );
  DFF \u_a23_mem/p_mem_reg[66][5]  ( .D(\u_a23_mem/n18887 ), .CLK(clk), .RST(
        rst), .I(p_init[533]), .Q(\u_a23_mem/p_mem[66][5] ) );
  DFF \u_a23_mem/p_mem_reg[66][6]  ( .D(\u_a23_mem/n18886 ), .CLK(clk), .RST(
        rst), .I(p_init[534]), .Q(\u_a23_mem/p_mem[66][6] ) );
  DFF \u_a23_mem/p_mem_reg[66][7]  ( .D(\u_a23_mem/n18885 ), .CLK(clk), .RST(
        rst), .I(p_init[535]), .Q(\u_a23_mem/p_mem[66][7] ) );
  DFF \u_a23_mem/p_mem_reg[67][0]  ( .D(\u_a23_mem/n18884 ), .CLK(clk), .RST(
        rst), .I(p_init[536]), .Q(\u_a23_mem/p_mem[67][0] ) );
  DFF \u_a23_mem/p_mem_reg[67][1]  ( .D(\u_a23_mem/n18883 ), .CLK(clk), .RST(
        rst), .I(p_init[537]), .Q(\u_a23_mem/p_mem[67][1] ) );
  DFF \u_a23_mem/p_mem_reg[67][2]  ( .D(\u_a23_mem/n18882 ), .CLK(clk), .RST(
        rst), .I(p_init[538]), .Q(\u_a23_mem/p_mem[67][2] ) );
  DFF \u_a23_mem/p_mem_reg[67][3]  ( .D(\u_a23_mem/n18881 ), .CLK(clk), .RST(
        rst), .I(p_init[539]), .Q(\u_a23_mem/p_mem[67][3] ) );
  DFF \u_a23_mem/p_mem_reg[67][4]  ( .D(\u_a23_mem/n18880 ), .CLK(clk), .RST(
        rst), .I(p_init[540]), .Q(\u_a23_mem/p_mem[67][4] ) );
  DFF \u_a23_mem/p_mem_reg[67][5]  ( .D(\u_a23_mem/n18879 ), .CLK(clk), .RST(
        rst), .I(p_init[541]), .Q(\u_a23_mem/p_mem[67][5] ) );
  DFF \u_a23_mem/p_mem_reg[67][6]  ( .D(\u_a23_mem/n18878 ), .CLK(clk), .RST(
        rst), .I(p_init[542]), .Q(\u_a23_mem/p_mem[67][6] ) );
  DFF \u_a23_mem/p_mem_reg[67][7]  ( .D(\u_a23_mem/n18877 ), .CLK(clk), .RST(
        rst), .I(p_init[543]), .Q(\u_a23_mem/p_mem[67][7] ) );
  DFF \u_a23_mem/p_mem_reg[68][0]  ( .D(\u_a23_mem/n18876 ), .CLK(clk), .RST(
        rst), .I(p_init[544]), .Q(\u_a23_mem/p_mem[68][0] ) );
  DFF \u_a23_mem/p_mem_reg[68][1]  ( .D(\u_a23_mem/n18875 ), .CLK(clk), .RST(
        rst), .I(p_init[545]), .Q(\u_a23_mem/p_mem[68][1] ) );
  DFF \u_a23_mem/p_mem_reg[68][2]  ( .D(\u_a23_mem/n18874 ), .CLK(clk), .RST(
        rst), .I(p_init[546]), .Q(\u_a23_mem/p_mem[68][2] ) );
  DFF \u_a23_mem/p_mem_reg[68][3]  ( .D(\u_a23_mem/n18873 ), .CLK(clk), .RST(
        rst), .I(p_init[547]), .Q(\u_a23_mem/p_mem[68][3] ) );
  DFF \u_a23_mem/p_mem_reg[68][4]  ( .D(\u_a23_mem/n18872 ), .CLK(clk), .RST(
        rst), .I(p_init[548]), .Q(\u_a23_mem/p_mem[68][4] ) );
  DFF \u_a23_mem/p_mem_reg[68][5]  ( .D(\u_a23_mem/n18871 ), .CLK(clk), .RST(
        rst), .I(p_init[549]), .Q(\u_a23_mem/p_mem[68][5] ) );
  DFF \u_a23_mem/p_mem_reg[68][6]  ( .D(\u_a23_mem/n18870 ), .CLK(clk), .RST(
        rst), .I(p_init[550]), .Q(\u_a23_mem/p_mem[68][6] ) );
  DFF \u_a23_mem/p_mem_reg[68][7]  ( .D(\u_a23_mem/n18869 ), .CLK(clk), .RST(
        rst), .I(p_init[551]), .Q(\u_a23_mem/p_mem[68][7] ) );
  DFF \u_a23_mem/p_mem_reg[69][0]  ( .D(\u_a23_mem/n18868 ), .CLK(clk), .RST(
        rst), .I(p_init[552]), .Q(\u_a23_mem/p_mem[69][0] ) );
  DFF \u_a23_mem/p_mem_reg[69][1]  ( .D(\u_a23_mem/n18867 ), .CLK(clk), .RST(
        rst), .I(p_init[553]), .Q(\u_a23_mem/p_mem[69][1] ) );
  DFF \u_a23_mem/p_mem_reg[69][2]  ( .D(\u_a23_mem/n18866 ), .CLK(clk), .RST(
        rst), .I(p_init[554]), .Q(\u_a23_mem/p_mem[69][2] ) );
  DFF \u_a23_mem/p_mem_reg[69][3]  ( .D(\u_a23_mem/n18865 ), .CLK(clk), .RST(
        rst), .I(p_init[555]), .Q(\u_a23_mem/p_mem[69][3] ) );
  DFF \u_a23_mem/p_mem_reg[69][4]  ( .D(\u_a23_mem/n18864 ), .CLK(clk), .RST(
        rst), .I(p_init[556]), .Q(\u_a23_mem/p_mem[69][4] ) );
  DFF \u_a23_mem/p_mem_reg[69][5]  ( .D(\u_a23_mem/n18863 ), .CLK(clk), .RST(
        rst), .I(p_init[557]), .Q(\u_a23_mem/p_mem[69][5] ) );
  DFF \u_a23_mem/p_mem_reg[69][6]  ( .D(\u_a23_mem/n18862 ), .CLK(clk), .RST(
        rst), .I(p_init[558]), .Q(\u_a23_mem/p_mem[69][6] ) );
  DFF \u_a23_mem/p_mem_reg[69][7]  ( .D(\u_a23_mem/n18861 ), .CLK(clk), .RST(
        rst), .I(p_init[559]), .Q(\u_a23_mem/p_mem[69][7] ) );
  DFF \u_a23_mem/p_mem_reg[70][0]  ( .D(\u_a23_mem/n18860 ), .CLK(clk), .RST(
        rst), .I(p_init[560]), .Q(\u_a23_mem/p_mem[70][0] ) );
  DFF \u_a23_mem/p_mem_reg[70][1]  ( .D(\u_a23_mem/n18859 ), .CLK(clk), .RST(
        rst), .I(p_init[561]), .Q(\u_a23_mem/p_mem[70][1] ) );
  DFF \u_a23_mem/p_mem_reg[70][2]  ( .D(\u_a23_mem/n18858 ), .CLK(clk), .RST(
        rst), .I(p_init[562]), .Q(\u_a23_mem/p_mem[70][2] ) );
  DFF \u_a23_mem/p_mem_reg[70][3]  ( .D(\u_a23_mem/n18857 ), .CLK(clk), .RST(
        rst), .I(p_init[563]), .Q(\u_a23_mem/p_mem[70][3] ) );
  DFF \u_a23_mem/p_mem_reg[70][4]  ( .D(\u_a23_mem/n18856 ), .CLK(clk), .RST(
        rst), .I(p_init[564]), .Q(\u_a23_mem/p_mem[70][4] ) );
  DFF \u_a23_mem/p_mem_reg[70][5]  ( .D(\u_a23_mem/n18855 ), .CLK(clk), .RST(
        rst), .I(p_init[565]), .Q(\u_a23_mem/p_mem[70][5] ) );
  DFF \u_a23_mem/p_mem_reg[70][6]  ( .D(\u_a23_mem/n18854 ), .CLK(clk), .RST(
        rst), .I(p_init[566]), .Q(\u_a23_mem/p_mem[70][6] ) );
  DFF \u_a23_mem/p_mem_reg[70][7]  ( .D(\u_a23_mem/n18853 ), .CLK(clk), .RST(
        rst), .I(p_init[567]), .Q(\u_a23_mem/p_mem[70][7] ) );
  DFF \u_a23_mem/p_mem_reg[71][0]  ( .D(\u_a23_mem/n18852 ), .CLK(clk), .RST(
        rst), .I(p_init[568]), .Q(\u_a23_mem/p_mem[71][0] ) );
  DFF \u_a23_mem/p_mem_reg[71][1]  ( .D(\u_a23_mem/n18851 ), .CLK(clk), .RST(
        rst), .I(p_init[569]), .Q(\u_a23_mem/p_mem[71][1] ) );
  DFF \u_a23_mem/p_mem_reg[71][2]  ( .D(\u_a23_mem/n18850 ), .CLK(clk), .RST(
        rst), .I(p_init[570]), .Q(\u_a23_mem/p_mem[71][2] ) );
  DFF \u_a23_mem/p_mem_reg[71][3]  ( .D(\u_a23_mem/n18849 ), .CLK(clk), .RST(
        rst), .I(p_init[571]), .Q(\u_a23_mem/p_mem[71][3] ) );
  DFF \u_a23_mem/p_mem_reg[71][4]  ( .D(\u_a23_mem/n18848 ), .CLK(clk), .RST(
        rst), .I(p_init[572]), .Q(\u_a23_mem/p_mem[71][4] ) );
  DFF \u_a23_mem/p_mem_reg[71][5]  ( .D(\u_a23_mem/n18847 ), .CLK(clk), .RST(
        rst), .I(p_init[573]), .Q(\u_a23_mem/p_mem[71][5] ) );
  DFF \u_a23_mem/p_mem_reg[71][6]  ( .D(\u_a23_mem/n18846 ), .CLK(clk), .RST(
        rst), .I(p_init[574]), .Q(\u_a23_mem/p_mem[71][6] ) );
  DFF \u_a23_mem/p_mem_reg[71][7]  ( .D(\u_a23_mem/n18845 ), .CLK(clk), .RST(
        rst), .I(p_init[575]), .Q(\u_a23_mem/p_mem[71][7] ) );
  DFF \u_a23_mem/p_mem_reg[72][0]  ( .D(\u_a23_mem/n18844 ), .CLK(clk), .RST(
        rst), .I(p_init[576]), .Q(\u_a23_mem/p_mem[72][0] ) );
  DFF \u_a23_mem/p_mem_reg[72][1]  ( .D(\u_a23_mem/n18843 ), .CLK(clk), .RST(
        rst), .I(p_init[577]), .Q(\u_a23_mem/p_mem[72][1] ) );
  DFF \u_a23_mem/p_mem_reg[72][2]  ( .D(\u_a23_mem/n18842 ), .CLK(clk), .RST(
        rst), .I(p_init[578]), .Q(\u_a23_mem/p_mem[72][2] ) );
  DFF \u_a23_mem/p_mem_reg[72][3]  ( .D(\u_a23_mem/n18841 ), .CLK(clk), .RST(
        rst), .I(p_init[579]), .Q(\u_a23_mem/p_mem[72][3] ) );
  DFF \u_a23_mem/p_mem_reg[72][4]  ( .D(\u_a23_mem/n18840 ), .CLK(clk), .RST(
        rst), .I(p_init[580]), .Q(\u_a23_mem/p_mem[72][4] ) );
  DFF \u_a23_mem/p_mem_reg[72][5]  ( .D(\u_a23_mem/n18839 ), .CLK(clk), .RST(
        rst), .I(p_init[581]), .Q(\u_a23_mem/p_mem[72][5] ) );
  DFF \u_a23_mem/p_mem_reg[72][6]  ( .D(\u_a23_mem/n18838 ), .CLK(clk), .RST(
        rst), .I(p_init[582]), .Q(\u_a23_mem/p_mem[72][6] ) );
  DFF \u_a23_mem/p_mem_reg[72][7]  ( .D(\u_a23_mem/n18837 ), .CLK(clk), .RST(
        rst), .I(p_init[583]), .Q(\u_a23_mem/p_mem[72][7] ) );
  DFF \u_a23_mem/p_mem_reg[73][0]  ( .D(\u_a23_mem/n18836 ), .CLK(clk), .RST(
        rst), .I(p_init[584]), .Q(\u_a23_mem/p_mem[73][0] ) );
  DFF \u_a23_mem/p_mem_reg[73][1]  ( .D(\u_a23_mem/n18835 ), .CLK(clk), .RST(
        rst), .I(p_init[585]), .Q(\u_a23_mem/p_mem[73][1] ) );
  DFF \u_a23_mem/p_mem_reg[73][2]  ( .D(\u_a23_mem/n18834 ), .CLK(clk), .RST(
        rst), .I(p_init[586]), .Q(\u_a23_mem/p_mem[73][2] ) );
  DFF \u_a23_mem/p_mem_reg[73][3]  ( .D(\u_a23_mem/n18833 ), .CLK(clk), .RST(
        rst), .I(p_init[587]), .Q(\u_a23_mem/p_mem[73][3] ) );
  DFF \u_a23_mem/p_mem_reg[73][4]  ( .D(\u_a23_mem/n18832 ), .CLK(clk), .RST(
        rst), .I(p_init[588]), .Q(\u_a23_mem/p_mem[73][4] ) );
  DFF \u_a23_mem/p_mem_reg[73][5]  ( .D(\u_a23_mem/n18831 ), .CLK(clk), .RST(
        rst), .I(p_init[589]), .Q(\u_a23_mem/p_mem[73][5] ) );
  DFF \u_a23_mem/p_mem_reg[73][6]  ( .D(\u_a23_mem/n18830 ), .CLK(clk), .RST(
        rst), .I(p_init[590]), .Q(\u_a23_mem/p_mem[73][6] ) );
  DFF \u_a23_mem/p_mem_reg[73][7]  ( .D(\u_a23_mem/n18829 ), .CLK(clk), .RST(
        rst), .I(p_init[591]), .Q(\u_a23_mem/p_mem[73][7] ) );
  DFF \u_a23_mem/p_mem_reg[74][0]  ( .D(\u_a23_mem/n18828 ), .CLK(clk), .RST(
        rst), .I(p_init[592]), .Q(\u_a23_mem/p_mem[74][0] ) );
  DFF \u_a23_mem/p_mem_reg[74][1]  ( .D(\u_a23_mem/n18827 ), .CLK(clk), .RST(
        rst), .I(p_init[593]), .Q(\u_a23_mem/p_mem[74][1] ) );
  DFF \u_a23_mem/p_mem_reg[74][2]  ( .D(\u_a23_mem/n18826 ), .CLK(clk), .RST(
        rst), .I(p_init[594]), .Q(\u_a23_mem/p_mem[74][2] ) );
  DFF \u_a23_mem/p_mem_reg[74][3]  ( .D(\u_a23_mem/n18825 ), .CLK(clk), .RST(
        rst), .I(p_init[595]), .Q(\u_a23_mem/p_mem[74][3] ) );
  DFF \u_a23_mem/p_mem_reg[74][4]  ( .D(\u_a23_mem/n18824 ), .CLK(clk), .RST(
        rst), .I(p_init[596]), .Q(\u_a23_mem/p_mem[74][4] ) );
  DFF \u_a23_mem/p_mem_reg[74][5]  ( .D(\u_a23_mem/n18823 ), .CLK(clk), .RST(
        rst), .I(p_init[597]), .Q(\u_a23_mem/p_mem[74][5] ) );
  DFF \u_a23_mem/p_mem_reg[74][6]  ( .D(\u_a23_mem/n18822 ), .CLK(clk), .RST(
        rst), .I(p_init[598]), .Q(\u_a23_mem/p_mem[74][6] ) );
  DFF \u_a23_mem/p_mem_reg[74][7]  ( .D(\u_a23_mem/n18821 ), .CLK(clk), .RST(
        rst), .I(p_init[599]), .Q(\u_a23_mem/p_mem[74][7] ) );
  DFF \u_a23_mem/p_mem_reg[75][0]  ( .D(\u_a23_mem/n18820 ), .CLK(clk), .RST(
        rst), .I(p_init[600]), .Q(\u_a23_mem/p_mem[75][0] ) );
  DFF \u_a23_mem/p_mem_reg[75][1]  ( .D(\u_a23_mem/n18819 ), .CLK(clk), .RST(
        rst), .I(p_init[601]), .Q(\u_a23_mem/p_mem[75][1] ) );
  DFF \u_a23_mem/p_mem_reg[75][2]  ( .D(\u_a23_mem/n18818 ), .CLK(clk), .RST(
        rst), .I(p_init[602]), .Q(\u_a23_mem/p_mem[75][2] ) );
  DFF \u_a23_mem/p_mem_reg[75][3]  ( .D(\u_a23_mem/n18817 ), .CLK(clk), .RST(
        rst), .I(p_init[603]), .Q(\u_a23_mem/p_mem[75][3] ) );
  DFF \u_a23_mem/p_mem_reg[75][4]  ( .D(\u_a23_mem/n18816 ), .CLK(clk), .RST(
        rst), .I(p_init[604]), .Q(\u_a23_mem/p_mem[75][4] ) );
  DFF \u_a23_mem/p_mem_reg[75][5]  ( .D(\u_a23_mem/n18815 ), .CLK(clk), .RST(
        rst), .I(p_init[605]), .Q(\u_a23_mem/p_mem[75][5] ) );
  DFF \u_a23_mem/p_mem_reg[75][6]  ( .D(\u_a23_mem/n18814 ), .CLK(clk), .RST(
        rst), .I(p_init[606]), .Q(\u_a23_mem/p_mem[75][6] ) );
  DFF \u_a23_mem/p_mem_reg[75][7]  ( .D(\u_a23_mem/n18813 ), .CLK(clk), .RST(
        rst), .I(p_init[607]), .Q(\u_a23_mem/p_mem[75][7] ) );
  DFF \u_a23_mem/p_mem_reg[76][0]  ( .D(\u_a23_mem/n18812 ), .CLK(clk), .RST(
        rst), .I(p_init[608]), .Q(\u_a23_mem/p_mem[76][0] ) );
  DFF \u_a23_mem/p_mem_reg[76][1]  ( .D(\u_a23_mem/n18811 ), .CLK(clk), .RST(
        rst), .I(p_init[609]), .Q(\u_a23_mem/p_mem[76][1] ) );
  DFF \u_a23_mem/p_mem_reg[76][2]  ( .D(\u_a23_mem/n18810 ), .CLK(clk), .RST(
        rst), .I(p_init[610]), .Q(\u_a23_mem/p_mem[76][2] ) );
  DFF \u_a23_mem/p_mem_reg[76][3]  ( .D(\u_a23_mem/n18809 ), .CLK(clk), .RST(
        rst), .I(p_init[611]), .Q(\u_a23_mem/p_mem[76][3] ) );
  DFF \u_a23_mem/p_mem_reg[76][4]  ( .D(\u_a23_mem/n18808 ), .CLK(clk), .RST(
        rst), .I(p_init[612]), .Q(\u_a23_mem/p_mem[76][4] ) );
  DFF \u_a23_mem/p_mem_reg[76][5]  ( .D(\u_a23_mem/n18807 ), .CLK(clk), .RST(
        rst), .I(p_init[613]), .Q(\u_a23_mem/p_mem[76][5] ) );
  DFF \u_a23_mem/p_mem_reg[76][6]  ( .D(\u_a23_mem/n18806 ), .CLK(clk), .RST(
        rst), .I(p_init[614]), .Q(\u_a23_mem/p_mem[76][6] ) );
  DFF \u_a23_mem/p_mem_reg[76][7]  ( .D(\u_a23_mem/n18805 ), .CLK(clk), .RST(
        rst), .I(p_init[615]), .Q(\u_a23_mem/p_mem[76][7] ) );
  DFF \u_a23_mem/p_mem_reg[77][0]  ( .D(\u_a23_mem/n18804 ), .CLK(clk), .RST(
        rst), .I(p_init[616]), .Q(\u_a23_mem/p_mem[77][0] ) );
  DFF \u_a23_mem/p_mem_reg[77][1]  ( .D(\u_a23_mem/n18803 ), .CLK(clk), .RST(
        rst), .I(p_init[617]), .Q(\u_a23_mem/p_mem[77][1] ) );
  DFF \u_a23_mem/p_mem_reg[77][2]  ( .D(\u_a23_mem/n18802 ), .CLK(clk), .RST(
        rst), .I(p_init[618]), .Q(\u_a23_mem/p_mem[77][2] ) );
  DFF \u_a23_mem/p_mem_reg[77][3]  ( .D(\u_a23_mem/n18801 ), .CLK(clk), .RST(
        rst), .I(p_init[619]), .Q(\u_a23_mem/p_mem[77][3] ) );
  DFF \u_a23_mem/p_mem_reg[77][4]  ( .D(\u_a23_mem/n18800 ), .CLK(clk), .RST(
        rst), .I(p_init[620]), .Q(\u_a23_mem/p_mem[77][4] ) );
  DFF \u_a23_mem/p_mem_reg[77][5]  ( .D(\u_a23_mem/n18799 ), .CLK(clk), .RST(
        rst), .I(p_init[621]), .Q(\u_a23_mem/p_mem[77][5] ) );
  DFF \u_a23_mem/p_mem_reg[77][6]  ( .D(\u_a23_mem/n18798 ), .CLK(clk), .RST(
        rst), .I(p_init[622]), .Q(\u_a23_mem/p_mem[77][6] ) );
  DFF \u_a23_mem/p_mem_reg[77][7]  ( .D(\u_a23_mem/n18797 ), .CLK(clk), .RST(
        rst), .I(p_init[623]), .Q(\u_a23_mem/p_mem[77][7] ) );
  DFF \u_a23_mem/p_mem_reg[78][0]  ( .D(\u_a23_mem/n18796 ), .CLK(clk), .RST(
        rst), .I(p_init[624]), .Q(\u_a23_mem/p_mem[78][0] ) );
  DFF \u_a23_mem/p_mem_reg[78][1]  ( .D(\u_a23_mem/n18795 ), .CLK(clk), .RST(
        rst), .I(p_init[625]), .Q(\u_a23_mem/p_mem[78][1] ) );
  DFF \u_a23_mem/p_mem_reg[78][2]  ( .D(\u_a23_mem/n18794 ), .CLK(clk), .RST(
        rst), .I(p_init[626]), .Q(\u_a23_mem/p_mem[78][2] ) );
  DFF \u_a23_mem/p_mem_reg[78][3]  ( .D(\u_a23_mem/n18793 ), .CLK(clk), .RST(
        rst), .I(p_init[627]), .Q(\u_a23_mem/p_mem[78][3] ) );
  DFF \u_a23_mem/p_mem_reg[78][4]  ( .D(\u_a23_mem/n18792 ), .CLK(clk), .RST(
        rst), .I(p_init[628]), .Q(\u_a23_mem/p_mem[78][4] ) );
  DFF \u_a23_mem/p_mem_reg[78][5]  ( .D(\u_a23_mem/n18791 ), .CLK(clk), .RST(
        rst), .I(p_init[629]), .Q(\u_a23_mem/p_mem[78][5] ) );
  DFF \u_a23_mem/p_mem_reg[78][6]  ( .D(\u_a23_mem/n18790 ), .CLK(clk), .RST(
        rst), .I(p_init[630]), .Q(\u_a23_mem/p_mem[78][6] ) );
  DFF \u_a23_mem/p_mem_reg[78][7]  ( .D(\u_a23_mem/n18789 ), .CLK(clk), .RST(
        rst), .I(p_init[631]), .Q(\u_a23_mem/p_mem[78][7] ) );
  DFF \u_a23_mem/p_mem_reg[79][0]  ( .D(\u_a23_mem/n18788 ), .CLK(clk), .RST(
        rst), .I(p_init[632]), .Q(\u_a23_mem/p_mem[79][0] ) );
  DFF \u_a23_mem/p_mem_reg[79][1]  ( .D(\u_a23_mem/n18787 ), .CLK(clk), .RST(
        rst), .I(p_init[633]), .Q(\u_a23_mem/p_mem[79][1] ) );
  DFF \u_a23_mem/p_mem_reg[79][2]  ( .D(\u_a23_mem/n18786 ), .CLK(clk), .RST(
        rst), .I(p_init[634]), .Q(\u_a23_mem/p_mem[79][2] ) );
  DFF \u_a23_mem/p_mem_reg[79][3]  ( .D(\u_a23_mem/n18785 ), .CLK(clk), .RST(
        rst), .I(p_init[635]), .Q(\u_a23_mem/p_mem[79][3] ) );
  DFF \u_a23_mem/p_mem_reg[79][4]  ( .D(\u_a23_mem/n18784 ), .CLK(clk), .RST(
        rst), .I(p_init[636]), .Q(\u_a23_mem/p_mem[79][4] ) );
  DFF \u_a23_mem/p_mem_reg[79][5]  ( .D(\u_a23_mem/n18783 ), .CLK(clk), .RST(
        rst), .I(p_init[637]), .Q(\u_a23_mem/p_mem[79][5] ) );
  DFF \u_a23_mem/p_mem_reg[79][6]  ( .D(\u_a23_mem/n18782 ), .CLK(clk), .RST(
        rst), .I(p_init[638]), .Q(\u_a23_mem/p_mem[79][6] ) );
  DFF \u_a23_mem/p_mem_reg[79][7]  ( .D(\u_a23_mem/n18781 ), .CLK(clk), .RST(
        rst), .I(p_init[639]), .Q(\u_a23_mem/p_mem[79][7] ) );
  DFF \u_a23_mem/p_mem_reg[80][0]  ( .D(\u_a23_mem/n18780 ), .CLK(clk), .RST(
        rst), .I(p_init[640]), .Q(\u_a23_mem/p_mem[80][0] ) );
  DFF \u_a23_mem/p_mem_reg[80][1]  ( .D(\u_a23_mem/n18779 ), .CLK(clk), .RST(
        rst), .I(p_init[641]), .Q(\u_a23_mem/p_mem[80][1] ) );
  DFF \u_a23_mem/p_mem_reg[80][2]  ( .D(\u_a23_mem/n18778 ), .CLK(clk), .RST(
        rst), .I(p_init[642]), .Q(\u_a23_mem/p_mem[80][2] ) );
  DFF \u_a23_mem/p_mem_reg[80][3]  ( .D(\u_a23_mem/n18777 ), .CLK(clk), .RST(
        rst), .I(p_init[643]), .Q(\u_a23_mem/p_mem[80][3] ) );
  DFF \u_a23_mem/p_mem_reg[80][4]  ( .D(\u_a23_mem/n18776 ), .CLK(clk), .RST(
        rst), .I(p_init[644]), .Q(\u_a23_mem/p_mem[80][4] ) );
  DFF \u_a23_mem/p_mem_reg[80][5]  ( .D(\u_a23_mem/n18775 ), .CLK(clk), .RST(
        rst), .I(p_init[645]), .Q(\u_a23_mem/p_mem[80][5] ) );
  DFF \u_a23_mem/p_mem_reg[80][6]  ( .D(\u_a23_mem/n18774 ), .CLK(clk), .RST(
        rst), .I(p_init[646]), .Q(\u_a23_mem/p_mem[80][6] ) );
  DFF \u_a23_mem/p_mem_reg[80][7]  ( .D(\u_a23_mem/n18773 ), .CLK(clk), .RST(
        rst), .I(p_init[647]), .Q(\u_a23_mem/p_mem[80][7] ) );
  DFF \u_a23_mem/p_mem_reg[81][0]  ( .D(\u_a23_mem/n18772 ), .CLK(clk), .RST(
        rst), .I(p_init[648]), .Q(\u_a23_mem/p_mem[81][0] ) );
  DFF \u_a23_mem/p_mem_reg[81][1]  ( .D(\u_a23_mem/n18771 ), .CLK(clk), .RST(
        rst), .I(p_init[649]), .Q(\u_a23_mem/p_mem[81][1] ) );
  DFF \u_a23_mem/p_mem_reg[81][2]  ( .D(\u_a23_mem/n18770 ), .CLK(clk), .RST(
        rst), .I(p_init[650]), .Q(\u_a23_mem/p_mem[81][2] ) );
  DFF \u_a23_mem/p_mem_reg[81][3]  ( .D(\u_a23_mem/n18769 ), .CLK(clk), .RST(
        rst), .I(p_init[651]), .Q(\u_a23_mem/p_mem[81][3] ) );
  DFF \u_a23_mem/p_mem_reg[81][4]  ( .D(\u_a23_mem/n18768 ), .CLK(clk), .RST(
        rst), .I(p_init[652]), .Q(\u_a23_mem/p_mem[81][4] ) );
  DFF \u_a23_mem/p_mem_reg[81][5]  ( .D(\u_a23_mem/n18767 ), .CLK(clk), .RST(
        rst), .I(p_init[653]), .Q(\u_a23_mem/p_mem[81][5] ) );
  DFF \u_a23_mem/p_mem_reg[81][6]  ( .D(\u_a23_mem/n18766 ), .CLK(clk), .RST(
        rst), .I(p_init[654]), .Q(\u_a23_mem/p_mem[81][6] ) );
  DFF \u_a23_mem/p_mem_reg[81][7]  ( .D(\u_a23_mem/n18765 ), .CLK(clk), .RST(
        rst), .I(p_init[655]), .Q(\u_a23_mem/p_mem[81][7] ) );
  DFF \u_a23_mem/p_mem_reg[82][0]  ( .D(\u_a23_mem/n18764 ), .CLK(clk), .RST(
        rst), .I(p_init[656]), .Q(\u_a23_mem/p_mem[82][0] ) );
  DFF \u_a23_mem/p_mem_reg[82][1]  ( .D(\u_a23_mem/n18763 ), .CLK(clk), .RST(
        rst), .I(p_init[657]), .Q(\u_a23_mem/p_mem[82][1] ) );
  DFF \u_a23_mem/p_mem_reg[82][2]  ( .D(\u_a23_mem/n18762 ), .CLK(clk), .RST(
        rst), .I(p_init[658]), .Q(\u_a23_mem/p_mem[82][2] ) );
  DFF \u_a23_mem/p_mem_reg[82][3]  ( .D(\u_a23_mem/n18761 ), .CLK(clk), .RST(
        rst), .I(p_init[659]), .Q(\u_a23_mem/p_mem[82][3] ) );
  DFF \u_a23_mem/p_mem_reg[82][4]  ( .D(\u_a23_mem/n18760 ), .CLK(clk), .RST(
        rst), .I(p_init[660]), .Q(\u_a23_mem/p_mem[82][4] ) );
  DFF \u_a23_mem/p_mem_reg[82][5]  ( .D(\u_a23_mem/n18759 ), .CLK(clk), .RST(
        rst), .I(p_init[661]), .Q(\u_a23_mem/p_mem[82][5] ) );
  DFF \u_a23_mem/p_mem_reg[82][6]  ( .D(\u_a23_mem/n18758 ), .CLK(clk), .RST(
        rst), .I(p_init[662]), .Q(\u_a23_mem/p_mem[82][6] ) );
  DFF \u_a23_mem/p_mem_reg[82][7]  ( .D(\u_a23_mem/n18757 ), .CLK(clk), .RST(
        rst), .I(p_init[663]), .Q(\u_a23_mem/p_mem[82][7] ) );
  DFF \u_a23_mem/p_mem_reg[83][0]  ( .D(\u_a23_mem/n18756 ), .CLK(clk), .RST(
        rst), .I(p_init[664]), .Q(\u_a23_mem/p_mem[83][0] ) );
  DFF \u_a23_mem/p_mem_reg[83][1]  ( .D(\u_a23_mem/n18755 ), .CLK(clk), .RST(
        rst), .I(p_init[665]), .Q(\u_a23_mem/p_mem[83][1] ) );
  DFF \u_a23_mem/p_mem_reg[83][2]  ( .D(\u_a23_mem/n18754 ), .CLK(clk), .RST(
        rst), .I(p_init[666]), .Q(\u_a23_mem/p_mem[83][2] ) );
  DFF \u_a23_mem/p_mem_reg[83][3]  ( .D(\u_a23_mem/n18753 ), .CLK(clk), .RST(
        rst), .I(p_init[667]), .Q(\u_a23_mem/p_mem[83][3] ) );
  DFF \u_a23_mem/p_mem_reg[83][4]  ( .D(\u_a23_mem/n18752 ), .CLK(clk), .RST(
        rst), .I(p_init[668]), .Q(\u_a23_mem/p_mem[83][4] ) );
  DFF \u_a23_mem/p_mem_reg[83][5]  ( .D(\u_a23_mem/n18751 ), .CLK(clk), .RST(
        rst), .I(p_init[669]), .Q(\u_a23_mem/p_mem[83][5] ) );
  DFF \u_a23_mem/p_mem_reg[83][6]  ( .D(\u_a23_mem/n18750 ), .CLK(clk), .RST(
        rst), .I(p_init[670]), .Q(\u_a23_mem/p_mem[83][6] ) );
  DFF \u_a23_mem/p_mem_reg[83][7]  ( .D(\u_a23_mem/n18749 ), .CLK(clk), .RST(
        rst), .I(p_init[671]), .Q(\u_a23_mem/p_mem[83][7] ) );
  DFF \u_a23_mem/p_mem_reg[84][0]  ( .D(\u_a23_mem/n18748 ), .CLK(clk), .RST(
        rst), .I(p_init[672]), .Q(\u_a23_mem/p_mem[84][0] ) );
  DFF \u_a23_mem/p_mem_reg[84][1]  ( .D(\u_a23_mem/n18747 ), .CLK(clk), .RST(
        rst), .I(p_init[673]), .Q(\u_a23_mem/p_mem[84][1] ) );
  DFF \u_a23_mem/p_mem_reg[84][2]  ( .D(\u_a23_mem/n18746 ), .CLK(clk), .RST(
        rst), .I(p_init[674]), .Q(\u_a23_mem/p_mem[84][2] ) );
  DFF \u_a23_mem/p_mem_reg[84][3]  ( .D(\u_a23_mem/n18745 ), .CLK(clk), .RST(
        rst), .I(p_init[675]), .Q(\u_a23_mem/p_mem[84][3] ) );
  DFF \u_a23_mem/p_mem_reg[84][4]  ( .D(\u_a23_mem/n18744 ), .CLK(clk), .RST(
        rst), .I(p_init[676]), .Q(\u_a23_mem/p_mem[84][4] ) );
  DFF \u_a23_mem/p_mem_reg[84][5]  ( .D(\u_a23_mem/n18743 ), .CLK(clk), .RST(
        rst), .I(p_init[677]), .Q(\u_a23_mem/p_mem[84][5] ) );
  DFF \u_a23_mem/p_mem_reg[84][6]  ( .D(\u_a23_mem/n18742 ), .CLK(clk), .RST(
        rst), .I(p_init[678]), .Q(\u_a23_mem/p_mem[84][6] ) );
  DFF \u_a23_mem/p_mem_reg[84][7]  ( .D(\u_a23_mem/n18741 ), .CLK(clk), .RST(
        rst), .I(p_init[679]), .Q(\u_a23_mem/p_mem[84][7] ) );
  DFF \u_a23_mem/p_mem_reg[85][0]  ( .D(\u_a23_mem/n18740 ), .CLK(clk), .RST(
        rst), .I(p_init[680]), .Q(\u_a23_mem/p_mem[85][0] ) );
  DFF \u_a23_mem/p_mem_reg[85][1]  ( .D(\u_a23_mem/n18739 ), .CLK(clk), .RST(
        rst), .I(p_init[681]), .Q(\u_a23_mem/p_mem[85][1] ) );
  DFF \u_a23_mem/p_mem_reg[85][2]  ( .D(\u_a23_mem/n18738 ), .CLK(clk), .RST(
        rst), .I(p_init[682]), .Q(\u_a23_mem/p_mem[85][2] ) );
  DFF \u_a23_mem/p_mem_reg[85][3]  ( .D(\u_a23_mem/n18737 ), .CLK(clk), .RST(
        rst), .I(p_init[683]), .Q(\u_a23_mem/p_mem[85][3] ) );
  DFF \u_a23_mem/p_mem_reg[85][4]  ( .D(\u_a23_mem/n18736 ), .CLK(clk), .RST(
        rst), .I(p_init[684]), .Q(\u_a23_mem/p_mem[85][4] ) );
  DFF \u_a23_mem/p_mem_reg[85][5]  ( .D(\u_a23_mem/n18735 ), .CLK(clk), .RST(
        rst), .I(p_init[685]), .Q(\u_a23_mem/p_mem[85][5] ) );
  DFF \u_a23_mem/p_mem_reg[85][6]  ( .D(\u_a23_mem/n18734 ), .CLK(clk), .RST(
        rst), .I(p_init[686]), .Q(\u_a23_mem/p_mem[85][6] ) );
  DFF \u_a23_mem/p_mem_reg[85][7]  ( .D(\u_a23_mem/n18733 ), .CLK(clk), .RST(
        rst), .I(p_init[687]), .Q(\u_a23_mem/p_mem[85][7] ) );
  DFF \u_a23_mem/p_mem_reg[86][0]  ( .D(\u_a23_mem/n18732 ), .CLK(clk), .RST(
        rst), .I(p_init[688]), .Q(\u_a23_mem/p_mem[86][0] ) );
  DFF \u_a23_mem/p_mem_reg[86][1]  ( .D(\u_a23_mem/n18731 ), .CLK(clk), .RST(
        rst), .I(p_init[689]), .Q(\u_a23_mem/p_mem[86][1] ) );
  DFF \u_a23_mem/p_mem_reg[86][2]  ( .D(\u_a23_mem/n18730 ), .CLK(clk), .RST(
        rst), .I(p_init[690]), .Q(\u_a23_mem/p_mem[86][2] ) );
  DFF \u_a23_mem/p_mem_reg[86][3]  ( .D(\u_a23_mem/n18729 ), .CLK(clk), .RST(
        rst), .I(p_init[691]), .Q(\u_a23_mem/p_mem[86][3] ) );
  DFF \u_a23_mem/p_mem_reg[86][4]  ( .D(\u_a23_mem/n18728 ), .CLK(clk), .RST(
        rst), .I(p_init[692]), .Q(\u_a23_mem/p_mem[86][4] ) );
  DFF \u_a23_mem/p_mem_reg[86][5]  ( .D(\u_a23_mem/n18727 ), .CLK(clk), .RST(
        rst), .I(p_init[693]), .Q(\u_a23_mem/p_mem[86][5] ) );
  DFF \u_a23_mem/p_mem_reg[86][6]  ( .D(\u_a23_mem/n18726 ), .CLK(clk), .RST(
        rst), .I(p_init[694]), .Q(\u_a23_mem/p_mem[86][6] ) );
  DFF \u_a23_mem/p_mem_reg[86][7]  ( .D(\u_a23_mem/n18725 ), .CLK(clk), .RST(
        rst), .I(p_init[695]), .Q(\u_a23_mem/p_mem[86][7] ) );
  DFF \u_a23_mem/p_mem_reg[87][0]  ( .D(\u_a23_mem/n18724 ), .CLK(clk), .RST(
        rst), .I(p_init[696]), .Q(\u_a23_mem/p_mem[87][0] ) );
  DFF \u_a23_mem/p_mem_reg[87][1]  ( .D(\u_a23_mem/n18723 ), .CLK(clk), .RST(
        rst), .I(p_init[697]), .Q(\u_a23_mem/p_mem[87][1] ) );
  DFF \u_a23_mem/p_mem_reg[87][2]  ( .D(\u_a23_mem/n18722 ), .CLK(clk), .RST(
        rst), .I(p_init[698]), .Q(\u_a23_mem/p_mem[87][2] ) );
  DFF \u_a23_mem/p_mem_reg[87][3]  ( .D(\u_a23_mem/n18721 ), .CLK(clk), .RST(
        rst), .I(p_init[699]), .Q(\u_a23_mem/p_mem[87][3] ) );
  DFF \u_a23_mem/p_mem_reg[87][4]  ( .D(\u_a23_mem/n18720 ), .CLK(clk), .RST(
        rst), .I(p_init[700]), .Q(\u_a23_mem/p_mem[87][4] ) );
  DFF \u_a23_mem/p_mem_reg[87][5]  ( .D(\u_a23_mem/n18719 ), .CLK(clk), .RST(
        rst), .I(p_init[701]), .Q(\u_a23_mem/p_mem[87][5] ) );
  DFF \u_a23_mem/p_mem_reg[87][6]  ( .D(\u_a23_mem/n18718 ), .CLK(clk), .RST(
        rst), .I(p_init[702]), .Q(\u_a23_mem/p_mem[87][6] ) );
  DFF \u_a23_mem/p_mem_reg[87][7]  ( .D(\u_a23_mem/n18717 ), .CLK(clk), .RST(
        rst), .I(p_init[703]), .Q(\u_a23_mem/p_mem[87][7] ) );
  DFF \u_a23_mem/p_mem_reg[88][0]  ( .D(\u_a23_mem/n18716 ), .CLK(clk), .RST(
        rst), .I(p_init[704]), .Q(\u_a23_mem/p_mem[88][0] ) );
  DFF \u_a23_mem/p_mem_reg[88][1]  ( .D(\u_a23_mem/n18715 ), .CLK(clk), .RST(
        rst), .I(p_init[705]), .Q(\u_a23_mem/p_mem[88][1] ) );
  DFF \u_a23_mem/p_mem_reg[88][2]  ( .D(\u_a23_mem/n18714 ), .CLK(clk), .RST(
        rst), .I(p_init[706]), .Q(\u_a23_mem/p_mem[88][2] ) );
  DFF \u_a23_mem/p_mem_reg[88][3]  ( .D(\u_a23_mem/n18713 ), .CLK(clk), .RST(
        rst), .I(p_init[707]), .Q(\u_a23_mem/p_mem[88][3] ) );
  DFF \u_a23_mem/p_mem_reg[88][4]  ( .D(\u_a23_mem/n18712 ), .CLK(clk), .RST(
        rst), .I(p_init[708]), .Q(\u_a23_mem/p_mem[88][4] ) );
  DFF \u_a23_mem/p_mem_reg[88][5]  ( .D(\u_a23_mem/n18711 ), .CLK(clk), .RST(
        rst), .I(p_init[709]), .Q(\u_a23_mem/p_mem[88][5] ) );
  DFF \u_a23_mem/p_mem_reg[88][6]  ( .D(\u_a23_mem/n18710 ), .CLK(clk), .RST(
        rst), .I(p_init[710]), .Q(\u_a23_mem/p_mem[88][6] ) );
  DFF \u_a23_mem/p_mem_reg[88][7]  ( .D(\u_a23_mem/n18709 ), .CLK(clk), .RST(
        rst), .I(p_init[711]), .Q(\u_a23_mem/p_mem[88][7] ) );
  DFF \u_a23_mem/p_mem_reg[89][0]  ( .D(\u_a23_mem/n18708 ), .CLK(clk), .RST(
        rst), .I(p_init[712]), .Q(\u_a23_mem/p_mem[89][0] ) );
  DFF \u_a23_mem/p_mem_reg[89][1]  ( .D(\u_a23_mem/n18707 ), .CLK(clk), .RST(
        rst), .I(p_init[713]), .Q(\u_a23_mem/p_mem[89][1] ) );
  DFF \u_a23_mem/p_mem_reg[89][2]  ( .D(\u_a23_mem/n18706 ), .CLK(clk), .RST(
        rst), .I(p_init[714]), .Q(\u_a23_mem/p_mem[89][2] ) );
  DFF \u_a23_mem/p_mem_reg[89][3]  ( .D(\u_a23_mem/n18705 ), .CLK(clk), .RST(
        rst), .I(p_init[715]), .Q(\u_a23_mem/p_mem[89][3] ) );
  DFF \u_a23_mem/p_mem_reg[89][4]  ( .D(\u_a23_mem/n18704 ), .CLK(clk), .RST(
        rst), .I(p_init[716]), .Q(\u_a23_mem/p_mem[89][4] ) );
  DFF \u_a23_mem/p_mem_reg[89][5]  ( .D(\u_a23_mem/n18703 ), .CLK(clk), .RST(
        rst), .I(p_init[717]), .Q(\u_a23_mem/p_mem[89][5] ) );
  DFF \u_a23_mem/p_mem_reg[89][6]  ( .D(\u_a23_mem/n18702 ), .CLK(clk), .RST(
        rst), .I(p_init[718]), .Q(\u_a23_mem/p_mem[89][6] ) );
  DFF \u_a23_mem/p_mem_reg[89][7]  ( .D(\u_a23_mem/n18701 ), .CLK(clk), .RST(
        rst), .I(p_init[719]), .Q(\u_a23_mem/p_mem[89][7] ) );
  DFF \u_a23_mem/p_mem_reg[90][0]  ( .D(\u_a23_mem/n18700 ), .CLK(clk), .RST(
        rst), .I(p_init[720]), .Q(\u_a23_mem/p_mem[90][0] ) );
  DFF \u_a23_mem/p_mem_reg[90][1]  ( .D(\u_a23_mem/n18699 ), .CLK(clk), .RST(
        rst), .I(p_init[721]), .Q(\u_a23_mem/p_mem[90][1] ) );
  DFF \u_a23_mem/p_mem_reg[90][2]  ( .D(\u_a23_mem/n18698 ), .CLK(clk), .RST(
        rst), .I(p_init[722]), .Q(\u_a23_mem/p_mem[90][2] ) );
  DFF \u_a23_mem/p_mem_reg[90][3]  ( .D(\u_a23_mem/n18697 ), .CLK(clk), .RST(
        rst), .I(p_init[723]), .Q(\u_a23_mem/p_mem[90][3] ) );
  DFF \u_a23_mem/p_mem_reg[90][4]  ( .D(\u_a23_mem/n18696 ), .CLK(clk), .RST(
        rst), .I(p_init[724]), .Q(\u_a23_mem/p_mem[90][4] ) );
  DFF \u_a23_mem/p_mem_reg[90][5]  ( .D(\u_a23_mem/n18695 ), .CLK(clk), .RST(
        rst), .I(p_init[725]), .Q(\u_a23_mem/p_mem[90][5] ) );
  DFF \u_a23_mem/p_mem_reg[90][6]  ( .D(\u_a23_mem/n18694 ), .CLK(clk), .RST(
        rst), .I(p_init[726]), .Q(\u_a23_mem/p_mem[90][6] ) );
  DFF \u_a23_mem/p_mem_reg[90][7]  ( .D(\u_a23_mem/n18693 ), .CLK(clk), .RST(
        rst), .I(p_init[727]), .Q(\u_a23_mem/p_mem[90][7] ) );
  DFF \u_a23_mem/p_mem_reg[91][0]  ( .D(\u_a23_mem/n18692 ), .CLK(clk), .RST(
        rst), .I(p_init[728]), .Q(\u_a23_mem/p_mem[91][0] ) );
  DFF \u_a23_mem/p_mem_reg[91][1]  ( .D(\u_a23_mem/n18691 ), .CLK(clk), .RST(
        rst), .I(p_init[729]), .Q(\u_a23_mem/p_mem[91][1] ) );
  DFF \u_a23_mem/p_mem_reg[91][2]  ( .D(\u_a23_mem/n18690 ), .CLK(clk), .RST(
        rst), .I(p_init[730]), .Q(\u_a23_mem/p_mem[91][2] ) );
  DFF \u_a23_mem/p_mem_reg[91][3]  ( .D(\u_a23_mem/n18689 ), .CLK(clk), .RST(
        rst), .I(p_init[731]), .Q(\u_a23_mem/p_mem[91][3] ) );
  DFF \u_a23_mem/p_mem_reg[91][4]  ( .D(\u_a23_mem/n18688 ), .CLK(clk), .RST(
        rst), .I(p_init[732]), .Q(\u_a23_mem/p_mem[91][4] ) );
  DFF \u_a23_mem/p_mem_reg[91][5]  ( .D(\u_a23_mem/n18687 ), .CLK(clk), .RST(
        rst), .I(p_init[733]), .Q(\u_a23_mem/p_mem[91][5] ) );
  DFF \u_a23_mem/p_mem_reg[91][6]  ( .D(\u_a23_mem/n18686 ), .CLK(clk), .RST(
        rst), .I(p_init[734]), .Q(\u_a23_mem/p_mem[91][6] ) );
  DFF \u_a23_mem/p_mem_reg[91][7]  ( .D(\u_a23_mem/n18685 ), .CLK(clk), .RST(
        rst), .I(p_init[735]), .Q(\u_a23_mem/p_mem[91][7] ) );
  DFF \u_a23_mem/p_mem_reg[92][0]  ( .D(\u_a23_mem/n18684 ), .CLK(clk), .RST(
        rst), .I(p_init[736]), .Q(\u_a23_mem/p_mem[92][0] ) );
  DFF \u_a23_mem/p_mem_reg[92][1]  ( .D(\u_a23_mem/n18683 ), .CLK(clk), .RST(
        rst), .I(p_init[737]), .Q(\u_a23_mem/p_mem[92][1] ) );
  DFF \u_a23_mem/p_mem_reg[92][2]  ( .D(\u_a23_mem/n18682 ), .CLK(clk), .RST(
        rst), .I(p_init[738]), .Q(\u_a23_mem/p_mem[92][2] ) );
  DFF \u_a23_mem/p_mem_reg[92][3]  ( .D(\u_a23_mem/n18681 ), .CLK(clk), .RST(
        rst), .I(p_init[739]), .Q(\u_a23_mem/p_mem[92][3] ) );
  DFF \u_a23_mem/p_mem_reg[92][4]  ( .D(\u_a23_mem/n18680 ), .CLK(clk), .RST(
        rst), .I(p_init[740]), .Q(\u_a23_mem/p_mem[92][4] ) );
  DFF \u_a23_mem/p_mem_reg[92][5]  ( .D(\u_a23_mem/n18679 ), .CLK(clk), .RST(
        rst), .I(p_init[741]), .Q(\u_a23_mem/p_mem[92][5] ) );
  DFF \u_a23_mem/p_mem_reg[92][6]  ( .D(\u_a23_mem/n18678 ), .CLK(clk), .RST(
        rst), .I(p_init[742]), .Q(\u_a23_mem/p_mem[92][6] ) );
  DFF \u_a23_mem/p_mem_reg[92][7]  ( .D(\u_a23_mem/n18677 ), .CLK(clk), .RST(
        rst), .I(p_init[743]), .Q(\u_a23_mem/p_mem[92][7] ) );
  DFF \u_a23_mem/p_mem_reg[93][0]  ( .D(\u_a23_mem/n18676 ), .CLK(clk), .RST(
        rst), .I(p_init[744]), .Q(\u_a23_mem/p_mem[93][0] ) );
  DFF \u_a23_mem/p_mem_reg[93][1]  ( .D(\u_a23_mem/n18675 ), .CLK(clk), .RST(
        rst), .I(p_init[745]), .Q(\u_a23_mem/p_mem[93][1] ) );
  DFF \u_a23_mem/p_mem_reg[93][2]  ( .D(\u_a23_mem/n18674 ), .CLK(clk), .RST(
        rst), .I(p_init[746]), .Q(\u_a23_mem/p_mem[93][2] ) );
  DFF \u_a23_mem/p_mem_reg[93][3]  ( .D(\u_a23_mem/n18673 ), .CLK(clk), .RST(
        rst), .I(p_init[747]), .Q(\u_a23_mem/p_mem[93][3] ) );
  DFF \u_a23_mem/p_mem_reg[93][4]  ( .D(\u_a23_mem/n18672 ), .CLK(clk), .RST(
        rst), .I(p_init[748]), .Q(\u_a23_mem/p_mem[93][4] ) );
  DFF \u_a23_mem/p_mem_reg[93][5]  ( .D(\u_a23_mem/n18671 ), .CLK(clk), .RST(
        rst), .I(p_init[749]), .Q(\u_a23_mem/p_mem[93][5] ) );
  DFF \u_a23_mem/p_mem_reg[93][6]  ( .D(\u_a23_mem/n18670 ), .CLK(clk), .RST(
        rst), .I(p_init[750]), .Q(\u_a23_mem/p_mem[93][6] ) );
  DFF \u_a23_mem/p_mem_reg[93][7]  ( .D(\u_a23_mem/n18669 ), .CLK(clk), .RST(
        rst), .I(p_init[751]), .Q(\u_a23_mem/p_mem[93][7] ) );
  DFF \u_a23_mem/p_mem_reg[94][0]  ( .D(\u_a23_mem/n18668 ), .CLK(clk), .RST(
        rst), .I(p_init[752]), .Q(\u_a23_mem/p_mem[94][0] ) );
  DFF \u_a23_mem/p_mem_reg[94][1]  ( .D(\u_a23_mem/n18667 ), .CLK(clk), .RST(
        rst), .I(p_init[753]), .Q(\u_a23_mem/p_mem[94][1] ) );
  DFF \u_a23_mem/p_mem_reg[94][2]  ( .D(\u_a23_mem/n18666 ), .CLK(clk), .RST(
        rst), .I(p_init[754]), .Q(\u_a23_mem/p_mem[94][2] ) );
  DFF \u_a23_mem/p_mem_reg[94][3]  ( .D(\u_a23_mem/n18665 ), .CLK(clk), .RST(
        rst), .I(p_init[755]), .Q(\u_a23_mem/p_mem[94][3] ) );
  DFF \u_a23_mem/p_mem_reg[94][4]  ( .D(\u_a23_mem/n18664 ), .CLK(clk), .RST(
        rst), .I(p_init[756]), .Q(\u_a23_mem/p_mem[94][4] ) );
  DFF \u_a23_mem/p_mem_reg[94][5]  ( .D(\u_a23_mem/n18663 ), .CLK(clk), .RST(
        rst), .I(p_init[757]), .Q(\u_a23_mem/p_mem[94][5] ) );
  DFF \u_a23_mem/p_mem_reg[94][6]  ( .D(\u_a23_mem/n18662 ), .CLK(clk), .RST(
        rst), .I(p_init[758]), .Q(\u_a23_mem/p_mem[94][6] ) );
  DFF \u_a23_mem/p_mem_reg[94][7]  ( .D(\u_a23_mem/n18661 ), .CLK(clk), .RST(
        rst), .I(p_init[759]), .Q(\u_a23_mem/p_mem[94][7] ) );
  DFF \u_a23_mem/p_mem_reg[95][0]  ( .D(\u_a23_mem/n18660 ), .CLK(clk), .RST(
        rst), .I(p_init[760]), .Q(\u_a23_mem/p_mem[95][0] ) );
  DFF \u_a23_mem/p_mem_reg[95][1]  ( .D(\u_a23_mem/n18659 ), .CLK(clk), .RST(
        rst), .I(p_init[761]), .Q(\u_a23_mem/p_mem[95][1] ) );
  DFF \u_a23_mem/p_mem_reg[95][2]  ( .D(\u_a23_mem/n18658 ), .CLK(clk), .RST(
        rst), .I(p_init[762]), .Q(\u_a23_mem/p_mem[95][2] ) );
  DFF \u_a23_mem/p_mem_reg[95][3]  ( .D(\u_a23_mem/n18657 ), .CLK(clk), .RST(
        rst), .I(p_init[763]), .Q(\u_a23_mem/p_mem[95][3] ) );
  DFF \u_a23_mem/p_mem_reg[95][4]  ( .D(\u_a23_mem/n18656 ), .CLK(clk), .RST(
        rst), .I(p_init[764]), .Q(\u_a23_mem/p_mem[95][4] ) );
  DFF \u_a23_mem/p_mem_reg[95][5]  ( .D(\u_a23_mem/n18655 ), .CLK(clk), .RST(
        rst), .I(p_init[765]), .Q(\u_a23_mem/p_mem[95][5] ) );
  DFF \u_a23_mem/p_mem_reg[95][6]  ( .D(\u_a23_mem/n18654 ), .CLK(clk), .RST(
        rst), .I(p_init[766]), .Q(\u_a23_mem/p_mem[95][6] ) );
  DFF \u_a23_mem/p_mem_reg[95][7]  ( .D(\u_a23_mem/n18653 ), .CLK(clk), .RST(
        rst), .I(p_init[767]), .Q(\u_a23_mem/p_mem[95][7] ) );
  DFF \u_a23_mem/p_mem_reg[96][0]  ( .D(\u_a23_mem/n18652 ), .CLK(clk), .RST(
        rst), .I(p_init[768]), .Q(\u_a23_mem/p_mem[96][0] ) );
  DFF \u_a23_mem/p_mem_reg[96][1]  ( .D(\u_a23_mem/n18651 ), .CLK(clk), .RST(
        rst), .I(p_init[769]), .Q(\u_a23_mem/p_mem[96][1] ) );
  DFF \u_a23_mem/p_mem_reg[96][2]  ( .D(\u_a23_mem/n18650 ), .CLK(clk), .RST(
        rst), .I(p_init[770]), .Q(\u_a23_mem/p_mem[96][2] ) );
  DFF \u_a23_mem/p_mem_reg[96][3]  ( .D(\u_a23_mem/n18649 ), .CLK(clk), .RST(
        rst), .I(p_init[771]), .Q(\u_a23_mem/p_mem[96][3] ) );
  DFF \u_a23_mem/p_mem_reg[96][4]  ( .D(\u_a23_mem/n18648 ), .CLK(clk), .RST(
        rst), .I(p_init[772]), .Q(\u_a23_mem/p_mem[96][4] ) );
  DFF \u_a23_mem/p_mem_reg[96][5]  ( .D(\u_a23_mem/n18647 ), .CLK(clk), .RST(
        rst), .I(p_init[773]), .Q(\u_a23_mem/p_mem[96][5] ) );
  DFF \u_a23_mem/p_mem_reg[96][6]  ( .D(\u_a23_mem/n18646 ), .CLK(clk), .RST(
        rst), .I(p_init[774]), .Q(\u_a23_mem/p_mem[96][6] ) );
  DFF \u_a23_mem/p_mem_reg[96][7]  ( .D(\u_a23_mem/n18645 ), .CLK(clk), .RST(
        rst), .I(p_init[775]), .Q(\u_a23_mem/p_mem[96][7] ) );
  DFF \u_a23_mem/p_mem_reg[97][0]  ( .D(\u_a23_mem/n18644 ), .CLK(clk), .RST(
        rst), .I(p_init[776]), .Q(\u_a23_mem/p_mem[97][0] ) );
  DFF \u_a23_mem/p_mem_reg[97][1]  ( .D(\u_a23_mem/n18643 ), .CLK(clk), .RST(
        rst), .I(p_init[777]), .Q(\u_a23_mem/p_mem[97][1] ) );
  DFF \u_a23_mem/p_mem_reg[97][2]  ( .D(\u_a23_mem/n18642 ), .CLK(clk), .RST(
        rst), .I(p_init[778]), .Q(\u_a23_mem/p_mem[97][2] ) );
  DFF \u_a23_mem/p_mem_reg[97][3]  ( .D(\u_a23_mem/n18641 ), .CLK(clk), .RST(
        rst), .I(p_init[779]), .Q(\u_a23_mem/p_mem[97][3] ) );
  DFF \u_a23_mem/p_mem_reg[97][4]  ( .D(\u_a23_mem/n18640 ), .CLK(clk), .RST(
        rst), .I(p_init[780]), .Q(\u_a23_mem/p_mem[97][4] ) );
  DFF \u_a23_mem/p_mem_reg[97][5]  ( .D(\u_a23_mem/n18639 ), .CLK(clk), .RST(
        rst), .I(p_init[781]), .Q(\u_a23_mem/p_mem[97][5] ) );
  DFF \u_a23_mem/p_mem_reg[97][6]  ( .D(\u_a23_mem/n18638 ), .CLK(clk), .RST(
        rst), .I(p_init[782]), .Q(\u_a23_mem/p_mem[97][6] ) );
  DFF \u_a23_mem/p_mem_reg[97][7]  ( .D(\u_a23_mem/n18637 ), .CLK(clk), .RST(
        rst), .I(p_init[783]), .Q(\u_a23_mem/p_mem[97][7] ) );
  DFF \u_a23_mem/p_mem_reg[98][0]  ( .D(\u_a23_mem/n18636 ), .CLK(clk), .RST(
        rst), .I(p_init[784]), .Q(\u_a23_mem/p_mem[98][0] ) );
  DFF \u_a23_mem/p_mem_reg[98][1]  ( .D(\u_a23_mem/n18635 ), .CLK(clk), .RST(
        rst), .I(p_init[785]), .Q(\u_a23_mem/p_mem[98][1] ) );
  DFF \u_a23_mem/p_mem_reg[98][2]  ( .D(\u_a23_mem/n18634 ), .CLK(clk), .RST(
        rst), .I(p_init[786]), .Q(\u_a23_mem/p_mem[98][2] ) );
  DFF \u_a23_mem/p_mem_reg[98][3]  ( .D(\u_a23_mem/n18633 ), .CLK(clk), .RST(
        rst), .I(p_init[787]), .Q(\u_a23_mem/p_mem[98][3] ) );
  DFF \u_a23_mem/p_mem_reg[98][4]  ( .D(\u_a23_mem/n18632 ), .CLK(clk), .RST(
        rst), .I(p_init[788]), .Q(\u_a23_mem/p_mem[98][4] ) );
  DFF \u_a23_mem/p_mem_reg[98][5]  ( .D(\u_a23_mem/n18631 ), .CLK(clk), .RST(
        rst), .I(p_init[789]), .Q(\u_a23_mem/p_mem[98][5] ) );
  DFF \u_a23_mem/p_mem_reg[98][6]  ( .D(\u_a23_mem/n18630 ), .CLK(clk), .RST(
        rst), .I(p_init[790]), .Q(\u_a23_mem/p_mem[98][6] ) );
  DFF \u_a23_mem/p_mem_reg[98][7]  ( .D(\u_a23_mem/n18629 ), .CLK(clk), .RST(
        rst), .I(p_init[791]), .Q(\u_a23_mem/p_mem[98][7] ) );
  DFF \u_a23_mem/p_mem_reg[99][0]  ( .D(\u_a23_mem/n18628 ), .CLK(clk), .RST(
        rst), .I(p_init[792]), .Q(\u_a23_mem/p_mem[99][0] ) );
  DFF \u_a23_mem/p_mem_reg[99][1]  ( .D(\u_a23_mem/n18627 ), .CLK(clk), .RST(
        rst), .I(p_init[793]), .Q(\u_a23_mem/p_mem[99][1] ) );
  DFF \u_a23_mem/p_mem_reg[99][2]  ( .D(\u_a23_mem/n18626 ), .CLK(clk), .RST(
        rst), .I(p_init[794]), .Q(\u_a23_mem/p_mem[99][2] ) );
  DFF \u_a23_mem/p_mem_reg[99][3]  ( .D(\u_a23_mem/n18625 ), .CLK(clk), .RST(
        rst), .I(p_init[795]), .Q(\u_a23_mem/p_mem[99][3] ) );
  DFF \u_a23_mem/p_mem_reg[99][4]  ( .D(\u_a23_mem/n18624 ), .CLK(clk), .RST(
        rst), .I(p_init[796]), .Q(\u_a23_mem/p_mem[99][4] ) );
  DFF \u_a23_mem/p_mem_reg[99][5]  ( .D(\u_a23_mem/n18623 ), .CLK(clk), .RST(
        rst), .I(p_init[797]), .Q(\u_a23_mem/p_mem[99][5] ) );
  DFF \u_a23_mem/p_mem_reg[99][6]  ( .D(\u_a23_mem/n18622 ), .CLK(clk), .RST(
        rst), .I(p_init[798]), .Q(\u_a23_mem/p_mem[99][6] ) );
  DFF \u_a23_mem/p_mem_reg[99][7]  ( .D(\u_a23_mem/n18621 ), .CLK(clk), .RST(
        rst), .I(p_init[799]), .Q(\u_a23_mem/p_mem[99][7] ) );
  DFF \u_a23_mem/p_mem_reg[100][0]  ( .D(\u_a23_mem/n18620 ), .CLK(clk), .RST(
        rst), .I(p_init[800]), .Q(\u_a23_mem/p_mem[100][0] ) );
  DFF \u_a23_mem/p_mem_reg[100][1]  ( .D(\u_a23_mem/n18619 ), .CLK(clk), .RST(
        rst), .I(p_init[801]), .Q(\u_a23_mem/p_mem[100][1] ) );
  DFF \u_a23_mem/p_mem_reg[100][2]  ( .D(\u_a23_mem/n18618 ), .CLK(clk), .RST(
        rst), .I(p_init[802]), .Q(\u_a23_mem/p_mem[100][2] ) );
  DFF \u_a23_mem/p_mem_reg[100][3]  ( .D(\u_a23_mem/n18617 ), .CLK(clk), .RST(
        rst), .I(p_init[803]), .Q(\u_a23_mem/p_mem[100][3] ) );
  DFF \u_a23_mem/p_mem_reg[100][4]  ( .D(\u_a23_mem/n18616 ), .CLK(clk), .RST(
        rst), .I(p_init[804]), .Q(\u_a23_mem/p_mem[100][4] ) );
  DFF \u_a23_mem/p_mem_reg[100][5]  ( .D(\u_a23_mem/n18615 ), .CLK(clk), .RST(
        rst), .I(p_init[805]), .Q(\u_a23_mem/p_mem[100][5] ) );
  DFF \u_a23_mem/p_mem_reg[100][6]  ( .D(\u_a23_mem/n18614 ), .CLK(clk), .RST(
        rst), .I(p_init[806]), .Q(\u_a23_mem/p_mem[100][6] ) );
  DFF \u_a23_mem/p_mem_reg[100][7]  ( .D(\u_a23_mem/n18613 ), .CLK(clk), .RST(
        rst), .I(p_init[807]), .Q(\u_a23_mem/p_mem[100][7] ) );
  DFF \u_a23_mem/p_mem_reg[101][0]  ( .D(\u_a23_mem/n18612 ), .CLK(clk), .RST(
        rst), .I(p_init[808]), .Q(\u_a23_mem/p_mem[101][0] ) );
  DFF \u_a23_mem/p_mem_reg[101][1]  ( .D(\u_a23_mem/n18611 ), .CLK(clk), .RST(
        rst), .I(p_init[809]), .Q(\u_a23_mem/p_mem[101][1] ) );
  DFF \u_a23_mem/p_mem_reg[101][2]  ( .D(\u_a23_mem/n18610 ), .CLK(clk), .RST(
        rst), .I(p_init[810]), .Q(\u_a23_mem/p_mem[101][2] ) );
  DFF \u_a23_mem/p_mem_reg[101][3]  ( .D(\u_a23_mem/n18609 ), .CLK(clk), .RST(
        rst), .I(p_init[811]), .Q(\u_a23_mem/p_mem[101][3] ) );
  DFF \u_a23_mem/p_mem_reg[101][4]  ( .D(\u_a23_mem/n18608 ), .CLK(clk), .RST(
        rst), .I(p_init[812]), .Q(\u_a23_mem/p_mem[101][4] ) );
  DFF \u_a23_mem/p_mem_reg[101][5]  ( .D(\u_a23_mem/n18607 ), .CLK(clk), .RST(
        rst), .I(p_init[813]), .Q(\u_a23_mem/p_mem[101][5] ) );
  DFF \u_a23_mem/p_mem_reg[101][6]  ( .D(\u_a23_mem/n18606 ), .CLK(clk), .RST(
        rst), .I(p_init[814]), .Q(\u_a23_mem/p_mem[101][6] ) );
  DFF \u_a23_mem/p_mem_reg[101][7]  ( .D(\u_a23_mem/n18605 ), .CLK(clk), .RST(
        rst), .I(p_init[815]), .Q(\u_a23_mem/p_mem[101][7] ) );
  DFF \u_a23_mem/p_mem_reg[102][0]  ( .D(\u_a23_mem/n18604 ), .CLK(clk), .RST(
        rst), .I(p_init[816]), .Q(\u_a23_mem/p_mem[102][0] ) );
  DFF \u_a23_mem/p_mem_reg[102][1]  ( .D(\u_a23_mem/n18603 ), .CLK(clk), .RST(
        rst), .I(p_init[817]), .Q(\u_a23_mem/p_mem[102][1] ) );
  DFF \u_a23_mem/p_mem_reg[102][2]  ( .D(\u_a23_mem/n18602 ), .CLK(clk), .RST(
        rst), .I(p_init[818]), .Q(\u_a23_mem/p_mem[102][2] ) );
  DFF \u_a23_mem/p_mem_reg[102][3]  ( .D(\u_a23_mem/n18601 ), .CLK(clk), .RST(
        rst), .I(p_init[819]), .Q(\u_a23_mem/p_mem[102][3] ) );
  DFF \u_a23_mem/p_mem_reg[102][4]  ( .D(\u_a23_mem/n18600 ), .CLK(clk), .RST(
        rst), .I(p_init[820]), .Q(\u_a23_mem/p_mem[102][4] ) );
  DFF \u_a23_mem/p_mem_reg[102][5]  ( .D(\u_a23_mem/n18599 ), .CLK(clk), .RST(
        rst), .I(p_init[821]), .Q(\u_a23_mem/p_mem[102][5] ) );
  DFF \u_a23_mem/p_mem_reg[102][6]  ( .D(\u_a23_mem/n18598 ), .CLK(clk), .RST(
        rst), .I(p_init[822]), .Q(\u_a23_mem/p_mem[102][6] ) );
  DFF \u_a23_mem/p_mem_reg[102][7]  ( .D(\u_a23_mem/n18597 ), .CLK(clk), .RST(
        rst), .I(p_init[823]), .Q(\u_a23_mem/p_mem[102][7] ) );
  DFF \u_a23_mem/p_mem_reg[103][0]  ( .D(\u_a23_mem/n18596 ), .CLK(clk), .RST(
        rst), .I(p_init[824]), .Q(\u_a23_mem/p_mem[103][0] ) );
  DFF \u_a23_mem/p_mem_reg[103][1]  ( .D(\u_a23_mem/n18595 ), .CLK(clk), .RST(
        rst), .I(p_init[825]), .Q(\u_a23_mem/p_mem[103][1] ) );
  DFF \u_a23_mem/p_mem_reg[103][2]  ( .D(\u_a23_mem/n18594 ), .CLK(clk), .RST(
        rst), .I(p_init[826]), .Q(\u_a23_mem/p_mem[103][2] ) );
  DFF \u_a23_mem/p_mem_reg[103][3]  ( .D(\u_a23_mem/n18593 ), .CLK(clk), .RST(
        rst), .I(p_init[827]), .Q(\u_a23_mem/p_mem[103][3] ) );
  DFF \u_a23_mem/p_mem_reg[103][4]  ( .D(\u_a23_mem/n18592 ), .CLK(clk), .RST(
        rst), .I(p_init[828]), .Q(\u_a23_mem/p_mem[103][4] ) );
  DFF \u_a23_mem/p_mem_reg[103][5]  ( .D(\u_a23_mem/n18591 ), .CLK(clk), .RST(
        rst), .I(p_init[829]), .Q(\u_a23_mem/p_mem[103][5] ) );
  DFF \u_a23_mem/p_mem_reg[103][6]  ( .D(\u_a23_mem/n18590 ), .CLK(clk), .RST(
        rst), .I(p_init[830]), .Q(\u_a23_mem/p_mem[103][6] ) );
  DFF \u_a23_mem/p_mem_reg[103][7]  ( .D(\u_a23_mem/n18589 ), .CLK(clk), .RST(
        rst), .I(p_init[831]), .Q(\u_a23_mem/p_mem[103][7] ) );
  DFF \u_a23_mem/p_mem_reg[104][0]  ( .D(\u_a23_mem/n18588 ), .CLK(clk), .RST(
        rst), .I(p_init[832]), .Q(\u_a23_mem/p_mem[104][0] ) );
  DFF \u_a23_mem/p_mem_reg[104][1]  ( .D(\u_a23_mem/n18587 ), .CLK(clk), .RST(
        rst), .I(p_init[833]), .Q(\u_a23_mem/p_mem[104][1] ) );
  DFF \u_a23_mem/p_mem_reg[104][2]  ( .D(\u_a23_mem/n18586 ), .CLK(clk), .RST(
        rst), .I(p_init[834]), .Q(\u_a23_mem/p_mem[104][2] ) );
  DFF \u_a23_mem/p_mem_reg[104][3]  ( .D(\u_a23_mem/n18585 ), .CLK(clk), .RST(
        rst), .I(p_init[835]), .Q(\u_a23_mem/p_mem[104][3] ) );
  DFF \u_a23_mem/p_mem_reg[104][4]  ( .D(\u_a23_mem/n18584 ), .CLK(clk), .RST(
        rst), .I(p_init[836]), .Q(\u_a23_mem/p_mem[104][4] ) );
  DFF \u_a23_mem/p_mem_reg[104][5]  ( .D(\u_a23_mem/n18583 ), .CLK(clk), .RST(
        rst), .I(p_init[837]), .Q(\u_a23_mem/p_mem[104][5] ) );
  DFF \u_a23_mem/p_mem_reg[104][6]  ( .D(\u_a23_mem/n18582 ), .CLK(clk), .RST(
        rst), .I(p_init[838]), .Q(\u_a23_mem/p_mem[104][6] ) );
  DFF \u_a23_mem/p_mem_reg[104][7]  ( .D(\u_a23_mem/n18581 ), .CLK(clk), .RST(
        rst), .I(p_init[839]), .Q(\u_a23_mem/p_mem[104][7] ) );
  DFF \u_a23_mem/p_mem_reg[105][0]  ( .D(\u_a23_mem/n18580 ), .CLK(clk), .RST(
        rst), .I(p_init[840]), .Q(\u_a23_mem/p_mem[105][0] ) );
  DFF \u_a23_mem/p_mem_reg[105][1]  ( .D(\u_a23_mem/n18579 ), .CLK(clk), .RST(
        rst), .I(p_init[841]), .Q(\u_a23_mem/p_mem[105][1] ) );
  DFF \u_a23_mem/p_mem_reg[105][2]  ( .D(\u_a23_mem/n18578 ), .CLK(clk), .RST(
        rst), .I(p_init[842]), .Q(\u_a23_mem/p_mem[105][2] ) );
  DFF \u_a23_mem/p_mem_reg[105][3]  ( .D(\u_a23_mem/n18577 ), .CLK(clk), .RST(
        rst), .I(p_init[843]), .Q(\u_a23_mem/p_mem[105][3] ) );
  DFF \u_a23_mem/p_mem_reg[105][4]  ( .D(\u_a23_mem/n18576 ), .CLK(clk), .RST(
        rst), .I(p_init[844]), .Q(\u_a23_mem/p_mem[105][4] ) );
  DFF \u_a23_mem/p_mem_reg[105][5]  ( .D(\u_a23_mem/n18575 ), .CLK(clk), .RST(
        rst), .I(p_init[845]), .Q(\u_a23_mem/p_mem[105][5] ) );
  DFF \u_a23_mem/p_mem_reg[105][6]  ( .D(\u_a23_mem/n18574 ), .CLK(clk), .RST(
        rst), .I(p_init[846]), .Q(\u_a23_mem/p_mem[105][6] ) );
  DFF \u_a23_mem/p_mem_reg[105][7]  ( .D(\u_a23_mem/n18573 ), .CLK(clk), .RST(
        rst), .I(p_init[847]), .Q(\u_a23_mem/p_mem[105][7] ) );
  DFF \u_a23_mem/p_mem_reg[106][0]  ( .D(\u_a23_mem/n18572 ), .CLK(clk), .RST(
        rst), .I(p_init[848]), .Q(\u_a23_mem/p_mem[106][0] ) );
  DFF \u_a23_mem/p_mem_reg[106][1]  ( .D(\u_a23_mem/n18571 ), .CLK(clk), .RST(
        rst), .I(p_init[849]), .Q(\u_a23_mem/p_mem[106][1] ) );
  DFF \u_a23_mem/p_mem_reg[106][2]  ( .D(\u_a23_mem/n18570 ), .CLK(clk), .RST(
        rst), .I(p_init[850]), .Q(\u_a23_mem/p_mem[106][2] ) );
  DFF \u_a23_mem/p_mem_reg[106][3]  ( .D(\u_a23_mem/n18569 ), .CLK(clk), .RST(
        rst), .I(p_init[851]), .Q(\u_a23_mem/p_mem[106][3] ) );
  DFF \u_a23_mem/p_mem_reg[106][4]  ( .D(\u_a23_mem/n18568 ), .CLK(clk), .RST(
        rst), .I(p_init[852]), .Q(\u_a23_mem/p_mem[106][4] ) );
  DFF \u_a23_mem/p_mem_reg[106][5]  ( .D(\u_a23_mem/n18567 ), .CLK(clk), .RST(
        rst), .I(p_init[853]), .Q(\u_a23_mem/p_mem[106][5] ) );
  DFF \u_a23_mem/p_mem_reg[106][6]  ( .D(\u_a23_mem/n18566 ), .CLK(clk), .RST(
        rst), .I(p_init[854]), .Q(\u_a23_mem/p_mem[106][6] ) );
  DFF \u_a23_mem/p_mem_reg[106][7]  ( .D(\u_a23_mem/n18565 ), .CLK(clk), .RST(
        rst), .I(p_init[855]), .Q(\u_a23_mem/p_mem[106][7] ) );
  DFF \u_a23_mem/p_mem_reg[107][0]  ( .D(\u_a23_mem/n18564 ), .CLK(clk), .RST(
        rst), .I(p_init[856]), .Q(\u_a23_mem/p_mem[107][0] ) );
  DFF \u_a23_mem/p_mem_reg[107][1]  ( .D(\u_a23_mem/n18563 ), .CLK(clk), .RST(
        rst), .I(p_init[857]), .Q(\u_a23_mem/p_mem[107][1] ) );
  DFF \u_a23_mem/p_mem_reg[107][2]  ( .D(\u_a23_mem/n18562 ), .CLK(clk), .RST(
        rst), .I(p_init[858]), .Q(\u_a23_mem/p_mem[107][2] ) );
  DFF \u_a23_mem/p_mem_reg[107][3]  ( .D(\u_a23_mem/n18561 ), .CLK(clk), .RST(
        rst), .I(p_init[859]), .Q(\u_a23_mem/p_mem[107][3] ) );
  DFF \u_a23_mem/p_mem_reg[107][4]  ( .D(\u_a23_mem/n18560 ), .CLK(clk), .RST(
        rst), .I(p_init[860]), .Q(\u_a23_mem/p_mem[107][4] ) );
  DFF \u_a23_mem/p_mem_reg[107][5]  ( .D(\u_a23_mem/n18559 ), .CLK(clk), .RST(
        rst), .I(p_init[861]), .Q(\u_a23_mem/p_mem[107][5] ) );
  DFF \u_a23_mem/p_mem_reg[107][6]  ( .D(\u_a23_mem/n18558 ), .CLK(clk), .RST(
        rst), .I(p_init[862]), .Q(\u_a23_mem/p_mem[107][6] ) );
  DFF \u_a23_mem/p_mem_reg[107][7]  ( .D(\u_a23_mem/n18557 ), .CLK(clk), .RST(
        rst), .I(p_init[863]), .Q(\u_a23_mem/p_mem[107][7] ) );
  DFF \u_a23_mem/p_mem_reg[108][0]  ( .D(\u_a23_mem/n18556 ), .CLK(clk), .RST(
        rst), .I(p_init[864]), .Q(\u_a23_mem/p_mem[108][0] ) );
  DFF \u_a23_mem/p_mem_reg[108][1]  ( .D(\u_a23_mem/n18555 ), .CLK(clk), .RST(
        rst), .I(p_init[865]), .Q(\u_a23_mem/p_mem[108][1] ) );
  DFF \u_a23_mem/p_mem_reg[108][2]  ( .D(\u_a23_mem/n18554 ), .CLK(clk), .RST(
        rst), .I(p_init[866]), .Q(\u_a23_mem/p_mem[108][2] ) );
  DFF \u_a23_mem/p_mem_reg[108][3]  ( .D(\u_a23_mem/n18553 ), .CLK(clk), .RST(
        rst), .I(p_init[867]), .Q(\u_a23_mem/p_mem[108][3] ) );
  DFF \u_a23_mem/p_mem_reg[108][4]  ( .D(\u_a23_mem/n18552 ), .CLK(clk), .RST(
        rst), .I(p_init[868]), .Q(\u_a23_mem/p_mem[108][4] ) );
  DFF \u_a23_mem/p_mem_reg[108][5]  ( .D(\u_a23_mem/n18551 ), .CLK(clk), .RST(
        rst), .I(p_init[869]), .Q(\u_a23_mem/p_mem[108][5] ) );
  DFF \u_a23_mem/p_mem_reg[108][6]  ( .D(\u_a23_mem/n18550 ), .CLK(clk), .RST(
        rst), .I(p_init[870]), .Q(\u_a23_mem/p_mem[108][6] ) );
  DFF \u_a23_mem/p_mem_reg[108][7]  ( .D(\u_a23_mem/n18549 ), .CLK(clk), .RST(
        rst), .I(p_init[871]), .Q(\u_a23_mem/p_mem[108][7] ) );
  DFF \u_a23_mem/p_mem_reg[109][0]  ( .D(\u_a23_mem/n18548 ), .CLK(clk), .RST(
        rst), .I(p_init[872]), .Q(\u_a23_mem/p_mem[109][0] ) );
  DFF \u_a23_mem/p_mem_reg[109][1]  ( .D(\u_a23_mem/n18547 ), .CLK(clk), .RST(
        rst), .I(p_init[873]), .Q(\u_a23_mem/p_mem[109][1] ) );
  DFF \u_a23_mem/p_mem_reg[109][2]  ( .D(\u_a23_mem/n18546 ), .CLK(clk), .RST(
        rst), .I(p_init[874]), .Q(\u_a23_mem/p_mem[109][2] ) );
  DFF \u_a23_mem/p_mem_reg[109][3]  ( .D(\u_a23_mem/n18545 ), .CLK(clk), .RST(
        rst), .I(p_init[875]), .Q(\u_a23_mem/p_mem[109][3] ) );
  DFF \u_a23_mem/p_mem_reg[109][4]  ( .D(\u_a23_mem/n18544 ), .CLK(clk), .RST(
        rst), .I(p_init[876]), .Q(\u_a23_mem/p_mem[109][4] ) );
  DFF \u_a23_mem/p_mem_reg[109][5]  ( .D(\u_a23_mem/n18543 ), .CLK(clk), .RST(
        rst), .I(p_init[877]), .Q(\u_a23_mem/p_mem[109][5] ) );
  DFF \u_a23_mem/p_mem_reg[109][6]  ( .D(\u_a23_mem/n18542 ), .CLK(clk), .RST(
        rst), .I(p_init[878]), .Q(\u_a23_mem/p_mem[109][6] ) );
  DFF \u_a23_mem/p_mem_reg[109][7]  ( .D(\u_a23_mem/n18541 ), .CLK(clk), .RST(
        rst), .I(p_init[879]), .Q(\u_a23_mem/p_mem[109][7] ) );
  DFF \u_a23_mem/p_mem_reg[110][0]  ( .D(\u_a23_mem/n18540 ), .CLK(clk), .RST(
        rst), .I(p_init[880]), .Q(\u_a23_mem/p_mem[110][0] ) );
  DFF \u_a23_mem/p_mem_reg[110][1]  ( .D(\u_a23_mem/n18539 ), .CLK(clk), .RST(
        rst), .I(p_init[881]), .Q(\u_a23_mem/p_mem[110][1] ) );
  DFF \u_a23_mem/p_mem_reg[110][2]  ( .D(\u_a23_mem/n18538 ), .CLK(clk), .RST(
        rst), .I(p_init[882]), .Q(\u_a23_mem/p_mem[110][2] ) );
  DFF \u_a23_mem/p_mem_reg[110][3]  ( .D(\u_a23_mem/n18537 ), .CLK(clk), .RST(
        rst), .I(p_init[883]), .Q(\u_a23_mem/p_mem[110][3] ) );
  DFF \u_a23_mem/p_mem_reg[110][4]  ( .D(\u_a23_mem/n18536 ), .CLK(clk), .RST(
        rst), .I(p_init[884]), .Q(\u_a23_mem/p_mem[110][4] ) );
  DFF \u_a23_mem/p_mem_reg[110][5]  ( .D(\u_a23_mem/n18535 ), .CLK(clk), .RST(
        rst), .I(p_init[885]), .Q(\u_a23_mem/p_mem[110][5] ) );
  DFF \u_a23_mem/p_mem_reg[110][6]  ( .D(\u_a23_mem/n18534 ), .CLK(clk), .RST(
        rst), .I(p_init[886]), .Q(\u_a23_mem/p_mem[110][6] ) );
  DFF \u_a23_mem/p_mem_reg[110][7]  ( .D(\u_a23_mem/n18533 ), .CLK(clk), .RST(
        rst), .I(p_init[887]), .Q(\u_a23_mem/p_mem[110][7] ) );
  DFF \u_a23_mem/p_mem_reg[111][0]  ( .D(\u_a23_mem/n18532 ), .CLK(clk), .RST(
        rst), .I(p_init[888]), .Q(\u_a23_mem/p_mem[111][0] ) );
  DFF \u_a23_mem/p_mem_reg[111][1]  ( .D(\u_a23_mem/n18531 ), .CLK(clk), .RST(
        rst), .I(p_init[889]), .Q(\u_a23_mem/p_mem[111][1] ) );
  DFF \u_a23_mem/p_mem_reg[111][2]  ( .D(\u_a23_mem/n18530 ), .CLK(clk), .RST(
        rst), .I(p_init[890]), .Q(\u_a23_mem/p_mem[111][2] ) );
  DFF \u_a23_mem/p_mem_reg[111][3]  ( .D(\u_a23_mem/n18529 ), .CLK(clk), .RST(
        rst), .I(p_init[891]), .Q(\u_a23_mem/p_mem[111][3] ) );
  DFF \u_a23_mem/p_mem_reg[111][4]  ( .D(\u_a23_mem/n18528 ), .CLK(clk), .RST(
        rst), .I(p_init[892]), .Q(\u_a23_mem/p_mem[111][4] ) );
  DFF \u_a23_mem/p_mem_reg[111][5]  ( .D(\u_a23_mem/n18527 ), .CLK(clk), .RST(
        rst), .I(p_init[893]), .Q(\u_a23_mem/p_mem[111][5] ) );
  DFF \u_a23_mem/p_mem_reg[111][6]  ( .D(\u_a23_mem/n18526 ), .CLK(clk), .RST(
        rst), .I(p_init[894]), .Q(\u_a23_mem/p_mem[111][6] ) );
  DFF \u_a23_mem/p_mem_reg[111][7]  ( .D(\u_a23_mem/n18525 ), .CLK(clk), .RST(
        rst), .I(p_init[895]), .Q(\u_a23_mem/p_mem[111][7] ) );
  DFF \u_a23_mem/p_mem_reg[112][0]  ( .D(\u_a23_mem/n18524 ), .CLK(clk), .RST(
        rst), .I(p_init[896]), .Q(\u_a23_mem/p_mem[112][0] ) );
  DFF \u_a23_mem/p_mem_reg[112][1]  ( .D(\u_a23_mem/n18523 ), .CLK(clk), .RST(
        rst), .I(p_init[897]), .Q(\u_a23_mem/p_mem[112][1] ) );
  DFF \u_a23_mem/p_mem_reg[112][2]  ( .D(\u_a23_mem/n18522 ), .CLK(clk), .RST(
        rst), .I(p_init[898]), .Q(\u_a23_mem/p_mem[112][2] ) );
  DFF \u_a23_mem/p_mem_reg[112][3]  ( .D(\u_a23_mem/n18521 ), .CLK(clk), .RST(
        rst), .I(p_init[899]), .Q(\u_a23_mem/p_mem[112][3] ) );
  DFF \u_a23_mem/p_mem_reg[112][4]  ( .D(\u_a23_mem/n18520 ), .CLK(clk), .RST(
        rst), .I(p_init[900]), .Q(\u_a23_mem/p_mem[112][4] ) );
  DFF \u_a23_mem/p_mem_reg[112][5]  ( .D(\u_a23_mem/n18519 ), .CLK(clk), .RST(
        rst), .I(p_init[901]), .Q(\u_a23_mem/p_mem[112][5] ) );
  DFF \u_a23_mem/p_mem_reg[112][6]  ( .D(\u_a23_mem/n18518 ), .CLK(clk), .RST(
        rst), .I(p_init[902]), .Q(\u_a23_mem/p_mem[112][6] ) );
  DFF \u_a23_mem/p_mem_reg[112][7]  ( .D(\u_a23_mem/n18517 ), .CLK(clk), .RST(
        rst), .I(p_init[903]), .Q(\u_a23_mem/p_mem[112][7] ) );
  DFF \u_a23_mem/p_mem_reg[113][0]  ( .D(\u_a23_mem/n18516 ), .CLK(clk), .RST(
        rst), .I(p_init[904]), .Q(\u_a23_mem/p_mem[113][0] ) );
  DFF \u_a23_mem/p_mem_reg[113][1]  ( .D(\u_a23_mem/n18515 ), .CLK(clk), .RST(
        rst), .I(p_init[905]), .Q(\u_a23_mem/p_mem[113][1] ) );
  DFF \u_a23_mem/p_mem_reg[113][2]  ( .D(\u_a23_mem/n18514 ), .CLK(clk), .RST(
        rst), .I(p_init[906]), .Q(\u_a23_mem/p_mem[113][2] ) );
  DFF \u_a23_mem/p_mem_reg[113][3]  ( .D(\u_a23_mem/n18513 ), .CLK(clk), .RST(
        rst), .I(p_init[907]), .Q(\u_a23_mem/p_mem[113][3] ) );
  DFF \u_a23_mem/p_mem_reg[113][4]  ( .D(\u_a23_mem/n18512 ), .CLK(clk), .RST(
        rst), .I(p_init[908]), .Q(\u_a23_mem/p_mem[113][4] ) );
  DFF \u_a23_mem/p_mem_reg[113][5]  ( .D(\u_a23_mem/n18511 ), .CLK(clk), .RST(
        rst), .I(p_init[909]), .Q(\u_a23_mem/p_mem[113][5] ) );
  DFF \u_a23_mem/p_mem_reg[113][6]  ( .D(\u_a23_mem/n18510 ), .CLK(clk), .RST(
        rst), .I(p_init[910]), .Q(\u_a23_mem/p_mem[113][6] ) );
  DFF \u_a23_mem/p_mem_reg[113][7]  ( .D(\u_a23_mem/n18509 ), .CLK(clk), .RST(
        rst), .I(p_init[911]), .Q(\u_a23_mem/p_mem[113][7] ) );
  DFF \u_a23_mem/p_mem_reg[114][0]  ( .D(\u_a23_mem/n18508 ), .CLK(clk), .RST(
        rst), .I(p_init[912]), .Q(\u_a23_mem/p_mem[114][0] ) );
  DFF \u_a23_mem/p_mem_reg[114][1]  ( .D(\u_a23_mem/n18507 ), .CLK(clk), .RST(
        rst), .I(p_init[913]), .Q(\u_a23_mem/p_mem[114][1] ) );
  DFF \u_a23_mem/p_mem_reg[114][2]  ( .D(\u_a23_mem/n18506 ), .CLK(clk), .RST(
        rst), .I(p_init[914]), .Q(\u_a23_mem/p_mem[114][2] ) );
  DFF \u_a23_mem/p_mem_reg[114][3]  ( .D(\u_a23_mem/n18505 ), .CLK(clk), .RST(
        rst), .I(p_init[915]), .Q(\u_a23_mem/p_mem[114][3] ) );
  DFF \u_a23_mem/p_mem_reg[114][4]  ( .D(\u_a23_mem/n18504 ), .CLK(clk), .RST(
        rst), .I(p_init[916]), .Q(\u_a23_mem/p_mem[114][4] ) );
  DFF \u_a23_mem/p_mem_reg[114][5]  ( .D(\u_a23_mem/n18503 ), .CLK(clk), .RST(
        rst), .I(p_init[917]), .Q(\u_a23_mem/p_mem[114][5] ) );
  DFF \u_a23_mem/p_mem_reg[114][6]  ( .D(\u_a23_mem/n18502 ), .CLK(clk), .RST(
        rst), .I(p_init[918]), .Q(\u_a23_mem/p_mem[114][6] ) );
  DFF \u_a23_mem/p_mem_reg[114][7]  ( .D(\u_a23_mem/n18501 ), .CLK(clk), .RST(
        rst), .I(p_init[919]), .Q(\u_a23_mem/p_mem[114][7] ) );
  DFF \u_a23_mem/p_mem_reg[115][0]  ( .D(\u_a23_mem/n18500 ), .CLK(clk), .RST(
        rst), .I(p_init[920]), .Q(\u_a23_mem/p_mem[115][0] ) );
  DFF \u_a23_mem/p_mem_reg[115][1]  ( .D(\u_a23_mem/n18499 ), .CLK(clk), .RST(
        rst), .I(p_init[921]), .Q(\u_a23_mem/p_mem[115][1] ) );
  DFF \u_a23_mem/p_mem_reg[115][2]  ( .D(\u_a23_mem/n18498 ), .CLK(clk), .RST(
        rst), .I(p_init[922]), .Q(\u_a23_mem/p_mem[115][2] ) );
  DFF \u_a23_mem/p_mem_reg[115][3]  ( .D(\u_a23_mem/n18497 ), .CLK(clk), .RST(
        rst), .I(p_init[923]), .Q(\u_a23_mem/p_mem[115][3] ) );
  DFF \u_a23_mem/p_mem_reg[115][4]  ( .D(\u_a23_mem/n18496 ), .CLK(clk), .RST(
        rst), .I(p_init[924]), .Q(\u_a23_mem/p_mem[115][4] ) );
  DFF \u_a23_mem/p_mem_reg[115][5]  ( .D(\u_a23_mem/n18495 ), .CLK(clk), .RST(
        rst), .I(p_init[925]), .Q(\u_a23_mem/p_mem[115][5] ) );
  DFF \u_a23_mem/p_mem_reg[115][6]  ( .D(\u_a23_mem/n18494 ), .CLK(clk), .RST(
        rst), .I(p_init[926]), .Q(\u_a23_mem/p_mem[115][6] ) );
  DFF \u_a23_mem/p_mem_reg[115][7]  ( .D(\u_a23_mem/n18493 ), .CLK(clk), .RST(
        rst), .I(p_init[927]), .Q(\u_a23_mem/p_mem[115][7] ) );
  DFF \u_a23_mem/p_mem_reg[116][0]  ( .D(\u_a23_mem/n18492 ), .CLK(clk), .RST(
        rst), .I(p_init[928]), .Q(\u_a23_mem/p_mem[116][0] ) );
  DFF \u_a23_mem/p_mem_reg[116][1]  ( .D(\u_a23_mem/n18491 ), .CLK(clk), .RST(
        rst), .I(p_init[929]), .Q(\u_a23_mem/p_mem[116][1] ) );
  DFF \u_a23_mem/p_mem_reg[116][2]  ( .D(\u_a23_mem/n18490 ), .CLK(clk), .RST(
        rst), .I(p_init[930]), .Q(\u_a23_mem/p_mem[116][2] ) );
  DFF \u_a23_mem/p_mem_reg[116][3]  ( .D(\u_a23_mem/n18489 ), .CLK(clk), .RST(
        rst), .I(p_init[931]), .Q(\u_a23_mem/p_mem[116][3] ) );
  DFF \u_a23_mem/p_mem_reg[116][4]  ( .D(\u_a23_mem/n18488 ), .CLK(clk), .RST(
        rst), .I(p_init[932]), .Q(\u_a23_mem/p_mem[116][4] ) );
  DFF \u_a23_mem/p_mem_reg[116][5]  ( .D(\u_a23_mem/n18487 ), .CLK(clk), .RST(
        rst), .I(p_init[933]), .Q(\u_a23_mem/p_mem[116][5] ) );
  DFF \u_a23_mem/p_mem_reg[116][6]  ( .D(\u_a23_mem/n18486 ), .CLK(clk), .RST(
        rst), .I(p_init[934]), .Q(\u_a23_mem/p_mem[116][6] ) );
  DFF \u_a23_mem/p_mem_reg[116][7]  ( .D(\u_a23_mem/n18485 ), .CLK(clk), .RST(
        rst), .I(p_init[935]), .Q(\u_a23_mem/p_mem[116][7] ) );
  DFF \u_a23_mem/p_mem_reg[117][0]  ( .D(\u_a23_mem/n18484 ), .CLK(clk), .RST(
        rst), .I(p_init[936]), .Q(\u_a23_mem/p_mem[117][0] ) );
  DFF \u_a23_mem/p_mem_reg[117][1]  ( .D(\u_a23_mem/n18483 ), .CLK(clk), .RST(
        rst), .I(p_init[937]), .Q(\u_a23_mem/p_mem[117][1] ) );
  DFF \u_a23_mem/p_mem_reg[117][2]  ( .D(\u_a23_mem/n18482 ), .CLK(clk), .RST(
        rst), .I(p_init[938]), .Q(\u_a23_mem/p_mem[117][2] ) );
  DFF \u_a23_mem/p_mem_reg[117][3]  ( .D(\u_a23_mem/n18481 ), .CLK(clk), .RST(
        rst), .I(p_init[939]), .Q(\u_a23_mem/p_mem[117][3] ) );
  DFF \u_a23_mem/p_mem_reg[117][4]  ( .D(\u_a23_mem/n18480 ), .CLK(clk), .RST(
        rst), .I(p_init[940]), .Q(\u_a23_mem/p_mem[117][4] ) );
  DFF \u_a23_mem/p_mem_reg[117][5]  ( .D(\u_a23_mem/n18479 ), .CLK(clk), .RST(
        rst), .I(p_init[941]), .Q(\u_a23_mem/p_mem[117][5] ) );
  DFF \u_a23_mem/p_mem_reg[117][6]  ( .D(\u_a23_mem/n18478 ), .CLK(clk), .RST(
        rst), .I(p_init[942]), .Q(\u_a23_mem/p_mem[117][6] ) );
  DFF \u_a23_mem/p_mem_reg[117][7]  ( .D(\u_a23_mem/n18477 ), .CLK(clk), .RST(
        rst), .I(p_init[943]), .Q(\u_a23_mem/p_mem[117][7] ) );
  DFF \u_a23_mem/p_mem_reg[118][0]  ( .D(\u_a23_mem/n18476 ), .CLK(clk), .RST(
        rst), .I(p_init[944]), .Q(\u_a23_mem/p_mem[118][0] ) );
  DFF \u_a23_mem/p_mem_reg[118][1]  ( .D(\u_a23_mem/n18475 ), .CLK(clk), .RST(
        rst), .I(p_init[945]), .Q(\u_a23_mem/p_mem[118][1] ) );
  DFF \u_a23_mem/p_mem_reg[118][2]  ( .D(\u_a23_mem/n18474 ), .CLK(clk), .RST(
        rst), .I(p_init[946]), .Q(\u_a23_mem/p_mem[118][2] ) );
  DFF \u_a23_mem/p_mem_reg[118][3]  ( .D(\u_a23_mem/n18473 ), .CLK(clk), .RST(
        rst), .I(p_init[947]), .Q(\u_a23_mem/p_mem[118][3] ) );
  DFF \u_a23_mem/p_mem_reg[118][4]  ( .D(\u_a23_mem/n18472 ), .CLK(clk), .RST(
        rst), .I(p_init[948]), .Q(\u_a23_mem/p_mem[118][4] ) );
  DFF \u_a23_mem/p_mem_reg[118][5]  ( .D(\u_a23_mem/n18471 ), .CLK(clk), .RST(
        rst), .I(p_init[949]), .Q(\u_a23_mem/p_mem[118][5] ) );
  DFF \u_a23_mem/p_mem_reg[118][6]  ( .D(\u_a23_mem/n18470 ), .CLK(clk), .RST(
        rst), .I(p_init[950]), .Q(\u_a23_mem/p_mem[118][6] ) );
  DFF \u_a23_mem/p_mem_reg[118][7]  ( .D(\u_a23_mem/n18469 ), .CLK(clk), .RST(
        rst), .I(p_init[951]), .Q(\u_a23_mem/p_mem[118][7] ) );
  DFF \u_a23_mem/p_mem_reg[119][0]  ( .D(\u_a23_mem/n18468 ), .CLK(clk), .RST(
        rst), .I(p_init[952]), .Q(\u_a23_mem/p_mem[119][0] ) );
  DFF \u_a23_mem/p_mem_reg[119][1]  ( .D(\u_a23_mem/n18467 ), .CLK(clk), .RST(
        rst), .I(p_init[953]), .Q(\u_a23_mem/p_mem[119][1] ) );
  DFF \u_a23_mem/p_mem_reg[119][2]  ( .D(\u_a23_mem/n18466 ), .CLK(clk), .RST(
        rst), .I(p_init[954]), .Q(\u_a23_mem/p_mem[119][2] ) );
  DFF \u_a23_mem/p_mem_reg[119][3]  ( .D(\u_a23_mem/n18465 ), .CLK(clk), .RST(
        rst), .I(p_init[955]), .Q(\u_a23_mem/p_mem[119][3] ) );
  DFF \u_a23_mem/p_mem_reg[119][4]  ( .D(\u_a23_mem/n18464 ), .CLK(clk), .RST(
        rst), .I(p_init[956]), .Q(\u_a23_mem/p_mem[119][4] ) );
  DFF \u_a23_mem/p_mem_reg[119][5]  ( .D(\u_a23_mem/n18463 ), .CLK(clk), .RST(
        rst), .I(p_init[957]), .Q(\u_a23_mem/p_mem[119][5] ) );
  DFF \u_a23_mem/p_mem_reg[119][6]  ( .D(\u_a23_mem/n18462 ), .CLK(clk), .RST(
        rst), .I(p_init[958]), .Q(\u_a23_mem/p_mem[119][6] ) );
  DFF \u_a23_mem/p_mem_reg[119][7]  ( .D(\u_a23_mem/n18461 ), .CLK(clk), .RST(
        rst), .I(p_init[959]), .Q(\u_a23_mem/p_mem[119][7] ) );
  DFF \u_a23_mem/p_mem_reg[120][0]  ( .D(\u_a23_mem/n18460 ), .CLK(clk), .RST(
        rst), .I(p_init[960]), .Q(\u_a23_mem/p_mem[120][0] ) );
  DFF \u_a23_mem/p_mem_reg[120][1]  ( .D(\u_a23_mem/n18459 ), .CLK(clk), .RST(
        rst), .I(p_init[961]), .Q(\u_a23_mem/p_mem[120][1] ) );
  DFF \u_a23_mem/p_mem_reg[120][2]  ( .D(\u_a23_mem/n18458 ), .CLK(clk), .RST(
        rst), .I(p_init[962]), .Q(\u_a23_mem/p_mem[120][2] ) );
  DFF \u_a23_mem/p_mem_reg[120][3]  ( .D(\u_a23_mem/n18457 ), .CLK(clk), .RST(
        rst), .I(p_init[963]), .Q(\u_a23_mem/p_mem[120][3] ) );
  DFF \u_a23_mem/p_mem_reg[120][4]  ( .D(\u_a23_mem/n18456 ), .CLK(clk), .RST(
        rst), .I(p_init[964]), .Q(\u_a23_mem/p_mem[120][4] ) );
  DFF \u_a23_mem/p_mem_reg[120][5]  ( .D(\u_a23_mem/n18455 ), .CLK(clk), .RST(
        rst), .I(p_init[965]), .Q(\u_a23_mem/p_mem[120][5] ) );
  DFF \u_a23_mem/p_mem_reg[120][6]  ( .D(\u_a23_mem/n18454 ), .CLK(clk), .RST(
        rst), .I(p_init[966]), .Q(\u_a23_mem/p_mem[120][6] ) );
  DFF \u_a23_mem/p_mem_reg[120][7]  ( .D(\u_a23_mem/n18453 ), .CLK(clk), .RST(
        rst), .I(p_init[967]), .Q(\u_a23_mem/p_mem[120][7] ) );
  DFF \u_a23_mem/p_mem_reg[121][0]  ( .D(\u_a23_mem/n18452 ), .CLK(clk), .RST(
        rst), .I(p_init[968]), .Q(\u_a23_mem/p_mem[121][0] ) );
  DFF \u_a23_mem/p_mem_reg[121][1]  ( .D(\u_a23_mem/n18451 ), .CLK(clk), .RST(
        rst), .I(p_init[969]), .Q(\u_a23_mem/p_mem[121][1] ) );
  DFF \u_a23_mem/p_mem_reg[121][2]  ( .D(\u_a23_mem/n18450 ), .CLK(clk), .RST(
        rst), .I(p_init[970]), .Q(\u_a23_mem/p_mem[121][2] ) );
  DFF \u_a23_mem/p_mem_reg[121][3]  ( .D(\u_a23_mem/n18449 ), .CLK(clk), .RST(
        rst), .I(p_init[971]), .Q(\u_a23_mem/p_mem[121][3] ) );
  DFF \u_a23_mem/p_mem_reg[121][4]  ( .D(\u_a23_mem/n18448 ), .CLK(clk), .RST(
        rst), .I(p_init[972]), .Q(\u_a23_mem/p_mem[121][4] ) );
  DFF \u_a23_mem/p_mem_reg[121][5]  ( .D(\u_a23_mem/n18447 ), .CLK(clk), .RST(
        rst), .I(p_init[973]), .Q(\u_a23_mem/p_mem[121][5] ) );
  DFF \u_a23_mem/p_mem_reg[121][6]  ( .D(\u_a23_mem/n18446 ), .CLK(clk), .RST(
        rst), .I(p_init[974]), .Q(\u_a23_mem/p_mem[121][6] ) );
  DFF \u_a23_mem/p_mem_reg[121][7]  ( .D(\u_a23_mem/n18445 ), .CLK(clk), .RST(
        rst), .I(p_init[975]), .Q(\u_a23_mem/p_mem[121][7] ) );
  DFF \u_a23_mem/p_mem_reg[122][0]  ( .D(\u_a23_mem/n18444 ), .CLK(clk), .RST(
        rst), .I(p_init[976]), .Q(\u_a23_mem/p_mem[122][0] ) );
  DFF \u_a23_mem/p_mem_reg[122][1]  ( .D(\u_a23_mem/n18443 ), .CLK(clk), .RST(
        rst), .I(p_init[977]), .Q(\u_a23_mem/p_mem[122][1] ) );
  DFF \u_a23_mem/p_mem_reg[122][2]  ( .D(\u_a23_mem/n18442 ), .CLK(clk), .RST(
        rst), .I(p_init[978]), .Q(\u_a23_mem/p_mem[122][2] ) );
  DFF \u_a23_mem/p_mem_reg[122][3]  ( .D(\u_a23_mem/n18441 ), .CLK(clk), .RST(
        rst), .I(p_init[979]), .Q(\u_a23_mem/p_mem[122][3] ) );
  DFF \u_a23_mem/p_mem_reg[122][4]  ( .D(\u_a23_mem/n18440 ), .CLK(clk), .RST(
        rst), .I(p_init[980]), .Q(\u_a23_mem/p_mem[122][4] ) );
  DFF \u_a23_mem/p_mem_reg[122][5]  ( .D(\u_a23_mem/n18439 ), .CLK(clk), .RST(
        rst), .I(p_init[981]), .Q(\u_a23_mem/p_mem[122][5] ) );
  DFF \u_a23_mem/p_mem_reg[122][6]  ( .D(\u_a23_mem/n18438 ), .CLK(clk), .RST(
        rst), .I(p_init[982]), .Q(\u_a23_mem/p_mem[122][6] ) );
  DFF \u_a23_mem/p_mem_reg[122][7]  ( .D(\u_a23_mem/n18437 ), .CLK(clk), .RST(
        rst), .I(p_init[983]), .Q(\u_a23_mem/p_mem[122][7] ) );
  DFF \u_a23_mem/p_mem_reg[123][0]  ( .D(\u_a23_mem/n18436 ), .CLK(clk), .RST(
        rst), .I(p_init[984]), .Q(\u_a23_mem/p_mem[123][0] ) );
  DFF \u_a23_mem/p_mem_reg[123][1]  ( .D(\u_a23_mem/n18435 ), .CLK(clk), .RST(
        rst), .I(p_init[985]), .Q(\u_a23_mem/p_mem[123][1] ) );
  DFF \u_a23_mem/p_mem_reg[123][2]  ( .D(\u_a23_mem/n18434 ), .CLK(clk), .RST(
        rst), .I(p_init[986]), .Q(\u_a23_mem/p_mem[123][2] ) );
  DFF \u_a23_mem/p_mem_reg[123][3]  ( .D(\u_a23_mem/n18433 ), .CLK(clk), .RST(
        rst), .I(p_init[987]), .Q(\u_a23_mem/p_mem[123][3] ) );
  DFF \u_a23_mem/p_mem_reg[123][4]  ( .D(\u_a23_mem/n18432 ), .CLK(clk), .RST(
        rst), .I(p_init[988]), .Q(\u_a23_mem/p_mem[123][4] ) );
  DFF \u_a23_mem/p_mem_reg[123][5]  ( .D(\u_a23_mem/n18431 ), .CLK(clk), .RST(
        rst), .I(p_init[989]), .Q(\u_a23_mem/p_mem[123][5] ) );
  DFF \u_a23_mem/p_mem_reg[123][6]  ( .D(\u_a23_mem/n18430 ), .CLK(clk), .RST(
        rst), .I(p_init[990]), .Q(\u_a23_mem/p_mem[123][6] ) );
  DFF \u_a23_mem/p_mem_reg[123][7]  ( .D(\u_a23_mem/n18429 ), .CLK(clk), .RST(
        rst), .I(p_init[991]), .Q(\u_a23_mem/p_mem[123][7] ) );
  DFF \u_a23_mem/p_mem_reg[124][0]  ( .D(\u_a23_mem/n18428 ), .CLK(clk), .RST(
        rst), .I(p_init[992]), .Q(\u_a23_mem/p_mem[124][0] ) );
  DFF \u_a23_mem/p_mem_reg[124][1]  ( .D(\u_a23_mem/n18427 ), .CLK(clk), .RST(
        rst), .I(p_init[993]), .Q(\u_a23_mem/p_mem[124][1] ) );
  DFF \u_a23_mem/p_mem_reg[124][2]  ( .D(\u_a23_mem/n18426 ), .CLK(clk), .RST(
        rst), .I(p_init[994]), .Q(\u_a23_mem/p_mem[124][2] ) );
  DFF \u_a23_mem/p_mem_reg[124][3]  ( .D(\u_a23_mem/n18425 ), .CLK(clk), .RST(
        rst), .I(p_init[995]), .Q(\u_a23_mem/p_mem[124][3] ) );
  DFF \u_a23_mem/p_mem_reg[124][4]  ( .D(\u_a23_mem/n18424 ), .CLK(clk), .RST(
        rst), .I(p_init[996]), .Q(\u_a23_mem/p_mem[124][4] ) );
  DFF \u_a23_mem/p_mem_reg[124][5]  ( .D(\u_a23_mem/n18423 ), .CLK(clk), .RST(
        rst), .I(p_init[997]), .Q(\u_a23_mem/p_mem[124][5] ) );
  DFF \u_a23_mem/p_mem_reg[124][6]  ( .D(\u_a23_mem/n18422 ), .CLK(clk), .RST(
        rst), .I(p_init[998]), .Q(\u_a23_mem/p_mem[124][6] ) );
  DFF \u_a23_mem/p_mem_reg[124][7]  ( .D(\u_a23_mem/n18421 ), .CLK(clk), .RST(
        rst), .I(p_init[999]), .Q(\u_a23_mem/p_mem[124][7] ) );
  DFF \u_a23_mem/p_mem_reg[125][0]  ( .D(\u_a23_mem/n18420 ), .CLK(clk), .RST(
        rst), .I(p_init[1000]), .Q(\u_a23_mem/p_mem[125][0] ) );
  DFF \u_a23_mem/p_mem_reg[125][1]  ( .D(\u_a23_mem/n18419 ), .CLK(clk), .RST(
        rst), .I(p_init[1001]), .Q(\u_a23_mem/p_mem[125][1] ) );
  DFF \u_a23_mem/p_mem_reg[125][2]  ( .D(\u_a23_mem/n18418 ), .CLK(clk), .RST(
        rst), .I(p_init[1002]), .Q(\u_a23_mem/p_mem[125][2] ) );
  DFF \u_a23_mem/p_mem_reg[125][3]  ( .D(\u_a23_mem/n18417 ), .CLK(clk), .RST(
        rst), .I(p_init[1003]), .Q(\u_a23_mem/p_mem[125][3] ) );
  DFF \u_a23_mem/p_mem_reg[125][4]  ( .D(\u_a23_mem/n18416 ), .CLK(clk), .RST(
        rst), .I(p_init[1004]), .Q(\u_a23_mem/p_mem[125][4] ) );
  DFF \u_a23_mem/p_mem_reg[125][5]  ( .D(\u_a23_mem/n18415 ), .CLK(clk), .RST(
        rst), .I(p_init[1005]), .Q(\u_a23_mem/p_mem[125][5] ) );
  DFF \u_a23_mem/p_mem_reg[125][6]  ( .D(\u_a23_mem/n18414 ), .CLK(clk), .RST(
        rst), .I(p_init[1006]), .Q(\u_a23_mem/p_mem[125][6] ) );
  DFF \u_a23_mem/p_mem_reg[125][7]  ( .D(\u_a23_mem/n18413 ), .CLK(clk), .RST(
        rst), .I(p_init[1007]), .Q(\u_a23_mem/p_mem[125][7] ) );
  DFF \u_a23_mem/p_mem_reg[126][0]  ( .D(\u_a23_mem/n18412 ), .CLK(clk), .RST(
        rst), .I(p_init[1008]), .Q(\u_a23_mem/p_mem[126][0] ) );
  DFF \u_a23_mem/p_mem_reg[126][1]  ( .D(\u_a23_mem/n18411 ), .CLK(clk), .RST(
        rst), .I(p_init[1009]), .Q(\u_a23_mem/p_mem[126][1] ) );
  DFF \u_a23_mem/p_mem_reg[126][2]  ( .D(\u_a23_mem/n18410 ), .CLK(clk), .RST(
        rst), .I(p_init[1010]), .Q(\u_a23_mem/p_mem[126][2] ) );
  DFF \u_a23_mem/p_mem_reg[126][3]  ( .D(\u_a23_mem/n18409 ), .CLK(clk), .RST(
        rst), .I(p_init[1011]), .Q(\u_a23_mem/p_mem[126][3] ) );
  DFF \u_a23_mem/p_mem_reg[126][4]  ( .D(\u_a23_mem/n18408 ), .CLK(clk), .RST(
        rst), .I(p_init[1012]), .Q(\u_a23_mem/p_mem[126][4] ) );
  DFF \u_a23_mem/p_mem_reg[126][5]  ( .D(\u_a23_mem/n18407 ), .CLK(clk), .RST(
        rst), .I(p_init[1013]), .Q(\u_a23_mem/p_mem[126][5] ) );
  DFF \u_a23_mem/p_mem_reg[126][6]  ( .D(\u_a23_mem/n18406 ), .CLK(clk), .RST(
        rst), .I(p_init[1014]), .Q(\u_a23_mem/p_mem[126][6] ) );
  DFF \u_a23_mem/p_mem_reg[126][7]  ( .D(\u_a23_mem/n18405 ), .CLK(clk), .RST(
        rst), .I(p_init[1015]), .Q(\u_a23_mem/p_mem[126][7] ) );
  DFF \u_a23_mem/p_mem_reg[127][0]  ( .D(\u_a23_mem/n18404 ), .CLK(clk), .RST(
        rst), .I(p_init[1016]), .Q(\u_a23_mem/p_mem[127][0] ) );
  DFF \u_a23_mem/p_mem_reg[127][1]  ( .D(\u_a23_mem/n18403 ), .CLK(clk), .RST(
        rst), .I(p_init[1017]), .Q(\u_a23_mem/p_mem[127][1] ) );
  DFF \u_a23_mem/p_mem_reg[127][2]  ( .D(\u_a23_mem/n18402 ), .CLK(clk), .RST(
        rst), .I(p_init[1018]), .Q(\u_a23_mem/p_mem[127][2] ) );
  DFF \u_a23_mem/p_mem_reg[127][3]  ( .D(\u_a23_mem/n18401 ), .CLK(clk), .RST(
        rst), .I(p_init[1019]), .Q(\u_a23_mem/p_mem[127][3] ) );
  DFF \u_a23_mem/p_mem_reg[127][4]  ( .D(\u_a23_mem/n18400 ), .CLK(clk), .RST(
        rst), .I(p_init[1020]), .Q(\u_a23_mem/p_mem[127][4] ) );
  DFF \u_a23_mem/p_mem_reg[127][5]  ( .D(\u_a23_mem/n18399 ), .CLK(clk), .RST(
        rst), .I(p_init[1021]), .Q(\u_a23_mem/p_mem[127][5] ) );
  DFF \u_a23_mem/p_mem_reg[127][6]  ( .D(\u_a23_mem/n18398 ), .CLK(clk), .RST(
        rst), .I(p_init[1022]), .Q(\u_a23_mem/p_mem[127][6] ) );
  DFF \u_a23_mem/p_mem_reg[127][7]  ( .D(\u_a23_mem/n18397 ), .CLK(clk), .RST(
        rst), .I(p_init[1023]), .Q(\u_a23_mem/p_mem[127][7] ) );
  DFF \u_a23_mem/stack_mem_reg[0][0]  ( .D(\u_a23_mem/n19652 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[0][0] ) );
  DFF \u_a23_mem/stack_mem_reg[0][1]  ( .D(\u_a23_mem/n19651 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[0][1] ) );
  DFF \u_a23_mem/stack_mem_reg[0][2]  ( .D(\u_a23_mem/n19650 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[0][2] ) );
  DFF \u_a23_mem/stack_mem_reg[0][3]  ( .D(\u_a23_mem/n19649 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[0][3] ) );
  DFF \u_a23_mem/stack_mem_reg[0][4]  ( .D(\u_a23_mem/n19648 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[0][4] ) );
  DFF \u_a23_mem/stack_mem_reg[0][5]  ( .D(\u_a23_mem/n19647 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[0][5] ) );
  DFF \u_a23_mem/stack_mem_reg[0][6]  ( .D(\u_a23_mem/n19646 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[0][6] ) );
  DFF \u_a23_mem/stack_mem_reg[0][7]  ( .D(\u_a23_mem/n19645 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[0][7] ) );
  DFF \u_a23_mem/stack_mem_reg[1][0]  ( .D(\u_a23_mem/n19644 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[1][0] ) );
  DFF \u_a23_mem/stack_mem_reg[1][1]  ( .D(\u_a23_mem/n19643 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[1][1] ) );
  DFF \u_a23_mem/stack_mem_reg[1][2]  ( .D(\u_a23_mem/n19642 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[1][2] ) );
  DFF \u_a23_mem/stack_mem_reg[1][3]  ( .D(\u_a23_mem/n19641 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[1][3] ) );
  DFF \u_a23_mem/stack_mem_reg[1][4]  ( .D(\u_a23_mem/n19640 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[1][4] ) );
  DFF \u_a23_mem/stack_mem_reg[1][5]  ( .D(\u_a23_mem/n19639 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[1][5] ) );
  DFF \u_a23_mem/stack_mem_reg[1][6]  ( .D(\u_a23_mem/n19638 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[1][6] ) );
  DFF \u_a23_mem/stack_mem_reg[1][7]  ( .D(\u_a23_mem/n19637 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[1][7] ) );
  DFF \u_a23_mem/stack_mem_reg[2][0]  ( .D(\u_a23_mem/n19636 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[2][0] ) );
  DFF \u_a23_mem/stack_mem_reg[2][1]  ( .D(\u_a23_mem/n19635 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[2][1] ) );
  DFF \u_a23_mem/stack_mem_reg[2][2]  ( .D(\u_a23_mem/n19634 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[2][2] ) );
  DFF \u_a23_mem/stack_mem_reg[2][3]  ( .D(\u_a23_mem/n19633 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[2][3] ) );
  DFF \u_a23_mem/stack_mem_reg[2][4]  ( .D(\u_a23_mem/n19632 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[2][4] ) );
  DFF \u_a23_mem/stack_mem_reg[2][5]  ( .D(\u_a23_mem/n19631 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[2][5] ) );
  DFF \u_a23_mem/stack_mem_reg[2][6]  ( .D(\u_a23_mem/n19630 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[2][6] ) );
  DFF \u_a23_mem/stack_mem_reg[2][7]  ( .D(\u_a23_mem/n19629 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[2][7] ) );
  DFF \u_a23_mem/stack_mem_reg[3][0]  ( .D(\u_a23_mem/n19628 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[3][0] ) );
  DFF \u_a23_mem/stack_mem_reg[3][1]  ( .D(\u_a23_mem/n19627 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[3][1] ) );
  DFF \u_a23_mem/stack_mem_reg[3][2]  ( .D(\u_a23_mem/n19626 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[3][2] ) );
  DFF \u_a23_mem/stack_mem_reg[3][3]  ( .D(\u_a23_mem/n19625 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[3][3] ) );
  DFF \u_a23_mem/stack_mem_reg[3][4]  ( .D(\u_a23_mem/n19624 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[3][4] ) );
  DFF \u_a23_mem/stack_mem_reg[3][5]  ( .D(\u_a23_mem/n19623 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[3][5] ) );
  DFF \u_a23_mem/stack_mem_reg[3][6]  ( .D(\u_a23_mem/n19622 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[3][6] ) );
  DFF \u_a23_mem/stack_mem_reg[3][7]  ( .D(\u_a23_mem/n19621 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[3][7] ) );
  DFF \u_a23_mem/stack_mem_reg[4][0]  ( .D(\u_a23_mem/n19620 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[4][0] ) );
  DFF \u_a23_mem/stack_mem_reg[4][1]  ( .D(\u_a23_mem/n19619 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[4][1] ) );
  DFF \u_a23_mem/stack_mem_reg[4][2]  ( .D(\u_a23_mem/n19618 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[4][2] ) );
  DFF \u_a23_mem/stack_mem_reg[4][3]  ( .D(\u_a23_mem/n19617 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[4][3] ) );
  DFF \u_a23_mem/stack_mem_reg[4][4]  ( .D(\u_a23_mem/n19616 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[4][4] ) );
  DFF \u_a23_mem/stack_mem_reg[4][5]  ( .D(\u_a23_mem/n19615 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[4][5] ) );
  DFF \u_a23_mem/stack_mem_reg[4][6]  ( .D(\u_a23_mem/n19614 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[4][6] ) );
  DFF \u_a23_mem/stack_mem_reg[4][7]  ( .D(\u_a23_mem/n19613 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[4][7] ) );
  DFF \u_a23_mem/stack_mem_reg[5][0]  ( .D(\u_a23_mem/n19612 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[5][0] ) );
  DFF \u_a23_mem/stack_mem_reg[5][1]  ( .D(\u_a23_mem/n19611 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[5][1] ) );
  DFF \u_a23_mem/stack_mem_reg[5][2]  ( .D(\u_a23_mem/n19610 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[5][2] ) );
  DFF \u_a23_mem/stack_mem_reg[5][3]  ( .D(\u_a23_mem/n19609 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[5][3] ) );
  DFF \u_a23_mem/stack_mem_reg[5][4]  ( .D(\u_a23_mem/n19608 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[5][4] ) );
  DFF \u_a23_mem/stack_mem_reg[5][5]  ( .D(\u_a23_mem/n19607 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[5][5] ) );
  DFF \u_a23_mem/stack_mem_reg[5][6]  ( .D(\u_a23_mem/n19606 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[5][6] ) );
  DFF \u_a23_mem/stack_mem_reg[5][7]  ( .D(\u_a23_mem/n19605 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[5][7] ) );
  DFF \u_a23_mem/stack_mem_reg[6][0]  ( .D(\u_a23_mem/n19604 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[6][0] ) );
  DFF \u_a23_mem/stack_mem_reg[6][1]  ( .D(\u_a23_mem/n19603 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[6][1] ) );
  DFF \u_a23_mem/stack_mem_reg[6][2]  ( .D(\u_a23_mem/n19602 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[6][2] ) );
  DFF \u_a23_mem/stack_mem_reg[6][3]  ( .D(\u_a23_mem/n19601 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[6][3] ) );
  DFF \u_a23_mem/stack_mem_reg[6][4]  ( .D(\u_a23_mem/n19600 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[6][4] ) );
  DFF \u_a23_mem/stack_mem_reg[6][5]  ( .D(\u_a23_mem/n19599 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[6][5] ) );
  DFF \u_a23_mem/stack_mem_reg[6][6]  ( .D(\u_a23_mem/n19598 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[6][6] ) );
  DFF \u_a23_mem/stack_mem_reg[6][7]  ( .D(\u_a23_mem/n19597 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[6][7] ) );
  DFF \u_a23_mem/stack_mem_reg[7][0]  ( .D(\u_a23_mem/n19596 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[7][0] ) );
  DFF \u_a23_mem/stack_mem_reg[7][1]  ( .D(\u_a23_mem/n19595 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[7][1] ) );
  DFF \u_a23_mem/stack_mem_reg[7][2]  ( .D(\u_a23_mem/n19594 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[7][2] ) );
  DFF \u_a23_mem/stack_mem_reg[7][3]  ( .D(\u_a23_mem/n19593 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[7][3] ) );
  DFF \u_a23_mem/stack_mem_reg[7][4]  ( .D(\u_a23_mem/n19592 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[7][4] ) );
  DFF \u_a23_mem/stack_mem_reg[7][5]  ( .D(\u_a23_mem/n19591 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[7][5] ) );
  DFF \u_a23_mem/stack_mem_reg[7][6]  ( .D(\u_a23_mem/n19590 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[7][6] ) );
  DFF \u_a23_mem/stack_mem_reg[7][7]  ( .D(\u_a23_mem/n19589 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[7][7] ) );
  DFF \u_a23_mem/stack_mem_reg[8][0]  ( .D(\u_a23_mem/n19588 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[8][0] ) );
  DFF \u_a23_mem/stack_mem_reg[8][1]  ( .D(\u_a23_mem/n19587 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[8][1] ) );
  DFF \u_a23_mem/stack_mem_reg[8][2]  ( .D(\u_a23_mem/n19586 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[8][2] ) );
  DFF \u_a23_mem/stack_mem_reg[8][3]  ( .D(\u_a23_mem/n19585 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[8][3] ) );
  DFF \u_a23_mem/stack_mem_reg[8][4]  ( .D(\u_a23_mem/n19584 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[8][4] ) );
  DFF \u_a23_mem/stack_mem_reg[8][5]  ( .D(\u_a23_mem/n19583 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[8][5] ) );
  DFF \u_a23_mem/stack_mem_reg[8][6]  ( .D(\u_a23_mem/n19582 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[8][6] ) );
  DFF \u_a23_mem/stack_mem_reg[8][7]  ( .D(\u_a23_mem/n19581 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[8][7] ) );
  DFF \u_a23_mem/stack_mem_reg[9][0]  ( .D(\u_a23_mem/n19580 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[9][0] ) );
  DFF \u_a23_mem/stack_mem_reg[9][1]  ( .D(\u_a23_mem/n19579 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[9][1] ) );
  DFF \u_a23_mem/stack_mem_reg[9][2]  ( .D(\u_a23_mem/n19578 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[9][2] ) );
  DFF \u_a23_mem/stack_mem_reg[9][3]  ( .D(\u_a23_mem/n19577 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[9][3] ) );
  DFF \u_a23_mem/stack_mem_reg[9][4]  ( .D(\u_a23_mem/n19576 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[9][4] ) );
  DFF \u_a23_mem/stack_mem_reg[9][5]  ( .D(\u_a23_mem/n19575 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[9][5] ) );
  DFF \u_a23_mem/stack_mem_reg[9][6]  ( .D(\u_a23_mem/n19574 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[9][6] ) );
  DFF \u_a23_mem/stack_mem_reg[9][7]  ( .D(\u_a23_mem/n19573 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[9][7] ) );
  DFF \u_a23_mem/stack_mem_reg[10][0]  ( .D(\u_a23_mem/n19572 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[10][0] ) );
  DFF \u_a23_mem/stack_mem_reg[10][1]  ( .D(\u_a23_mem/n19571 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[10][1] ) );
  DFF \u_a23_mem/stack_mem_reg[10][2]  ( .D(\u_a23_mem/n19570 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[10][2] ) );
  DFF \u_a23_mem/stack_mem_reg[10][3]  ( .D(\u_a23_mem/n19569 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[10][3] ) );
  DFF \u_a23_mem/stack_mem_reg[10][4]  ( .D(\u_a23_mem/n19568 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[10][4] ) );
  DFF \u_a23_mem/stack_mem_reg[10][5]  ( .D(\u_a23_mem/n19567 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[10][5] ) );
  DFF \u_a23_mem/stack_mem_reg[10][6]  ( .D(\u_a23_mem/n19566 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[10][6] ) );
  DFF \u_a23_mem/stack_mem_reg[10][7]  ( .D(\u_a23_mem/n19565 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[10][7] ) );
  DFF \u_a23_mem/stack_mem_reg[11][0]  ( .D(\u_a23_mem/n19564 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[11][0] ) );
  DFF \u_a23_mem/stack_mem_reg[11][1]  ( .D(\u_a23_mem/n19563 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[11][1] ) );
  DFF \u_a23_mem/stack_mem_reg[11][2]  ( .D(\u_a23_mem/n19562 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[11][2] ) );
  DFF \u_a23_mem/stack_mem_reg[11][3]  ( .D(\u_a23_mem/n19561 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[11][3] ) );
  DFF \u_a23_mem/stack_mem_reg[11][4]  ( .D(\u_a23_mem/n19560 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[11][4] ) );
  DFF \u_a23_mem/stack_mem_reg[11][5]  ( .D(\u_a23_mem/n19559 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[11][5] ) );
  DFF \u_a23_mem/stack_mem_reg[11][6]  ( .D(\u_a23_mem/n19558 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[11][6] ) );
  DFF \u_a23_mem/stack_mem_reg[11][7]  ( .D(\u_a23_mem/n19557 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[11][7] ) );
  DFF \u_a23_mem/stack_mem_reg[12][0]  ( .D(\u_a23_mem/n19556 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[12][0] ) );
  DFF \u_a23_mem/stack_mem_reg[12][1]  ( .D(\u_a23_mem/n19555 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[12][1] ) );
  DFF \u_a23_mem/stack_mem_reg[12][2]  ( .D(\u_a23_mem/n19554 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[12][2] ) );
  DFF \u_a23_mem/stack_mem_reg[12][3]  ( .D(\u_a23_mem/n19553 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[12][3] ) );
  DFF \u_a23_mem/stack_mem_reg[12][4]  ( .D(\u_a23_mem/n19552 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[12][4] ) );
  DFF \u_a23_mem/stack_mem_reg[12][5]  ( .D(\u_a23_mem/n19551 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[12][5] ) );
  DFF \u_a23_mem/stack_mem_reg[12][6]  ( .D(\u_a23_mem/n19550 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[12][6] ) );
  DFF \u_a23_mem/stack_mem_reg[12][7]  ( .D(\u_a23_mem/n19549 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[12][7] ) );
  DFF \u_a23_mem/stack_mem_reg[13][0]  ( .D(\u_a23_mem/n19548 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[13][0] ) );
  DFF \u_a23_mem/stack_mem_reg[13][1]  ( .D(\u_a23_mem/n19547 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[13][1] ) );
  DFF \u_a23_mem/stack_mem_reg[13][2]  ( .D(\u_a23_mem/n19546 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[13][2] ) );
  DFF \u_a23_mem/stack_mem_reg[13][3]  ( .D(\u_a23_mem/n19545 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[13][3] ) );
  DFF \u_a23_mem/stack_mem_reg[13][4]  ( .D(\u_a23_mem/n19544 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[13][4] ) );
  DFF \u_a23_mem/stack_mem_reg[13][5]  ( .D(\u_a23_mem/n19543 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[13][5] ) );
  DFF \u_a23_mem/stack_mem_reg[13][6]  ( .D(\u_a23_mem/n19542 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[13][6] ) );
  DFF \u_a23_mem/stack_mem_reg[13][7]  ( .D(\u_a23_mem/n19541 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[13][7] ) );
  DFF \u_a23_mem/stack_mem_reg[14][0]  ( .D(\u_a23_mem/n19540 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[14][0] ) );
  DFF \u_a23_mem/stack_mem_reg[14][1]  ( .D(\u_a23_mem/n19539 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[14][1] ) );
  DFF \u_a23_mem/stack_mem_reg[14][2]  ( .D(\u_a23_mem/n19538 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[14][2] ) );
  DFF \u_a23_mem/stack_mem_reg[14][3]  ( .D(\u_a23_mem/n19537 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[14][3] ) );
  DFF \u_a23_mem/stack_mem_reg[14][4]  ( .D(\u_a23_mem/n19536 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[14][4] ) );
  DFF \u_a23_mem/stack_mem_reg[14][5]  ( .D(\u_a23_mem/n19535 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[14][5] ) );
  DFF \u_a23_mem/stack_mem_reg[14][6]  ( .D(\u_a23_mem/n19534 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[14][6] ) );
  DFF \u_a23_mem/stack_mem_reg[14][7]  ( .D(\u_a23_mem/n19533 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[14][7] ) );
  DFF \u_a23_mem/stack_mem_reg[15][0]  ( .D(\u_a23_mem/n19532 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[15][0] ) );
  DFF \u_a23_mem/stack_mem_reg[15][1]  ( .D(\u_a23_mem/n19531 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[15][1] ) );
  DFF \u_a23_mem/stack_mem_reg[15][2]  ( .D(\u_a23_mem/n19530 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[15][2] ) );
  DFF \u_a23_mem/stack_mem_reg[15][3]  ( .D(\u_a23_mem/n19529 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[15][3] ) );
  DFF \u_a23_mem/stack_mem_reg[15][4]  ( .D(\u_a23_mem/n19528 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[15][4] ) );
  DFF \u_a23_mem/stack_mem_reg[15][5]  ( .D(\u_a23_mem/n19527 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[15][5] ) );
  DFF \u_a23_mem/stack_mem_reg[15][6]  ( .D(\u_a23_mem/n19526 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[15][6] ) );
  DFF \u_a23_mem/stack_mem_reg[15][7]  ( .D(\u_a23_mem/n19525 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[15][7] ) );
  DFF \u_a23_mem/stack_mem_reg[16][0]  ( .D(\u_a23_mem/n19524 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[16][0] ) );
  DFF \u_a23_mem/stack_mem_reg[16][1]  ( .D(\u_a23_mem/n19523 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[16][1] ) );
  DFF \u_a23_mem/stack_mem_reg[16][2]  ( .D(\u_a23_mem/n19522 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[16][2] ) );
  DFF \u_a23_mem/stack_mem_reg[16][3]  ( .D(\u_a23_mem/n19521 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[16][3] ) );
  DFF \u_a23_mem/stack_mem_reg[16][4]  ( .D(\u_a23_mem/n19520 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[16][4] ) );
  DFF \u_a23_mem/stack_mem_reg[16][5]  ( .D(\u_a23_mem/n19519 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[16][5] ) );
  DFF \u_a23_mem/stack_mem_reg[16][6]  ( .D(\u_a23_mem/n19518 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[16][6] ) );
  DFF \u_a23_mem/stack_mem_reg[16][7]  ( .D(\u_a23_mem/n19517 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[16][7] ) );
  DFF \u_a23_mem/stack_mem_reg[17][0]  ( .D(\u_a23_mem/n19516 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[17][0] ) );
  DFF \u_a23_mem/stack_mem_reg[17][1]  ( .D(\u_a23_mem/n19515 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[17][1] ) );
  DFF \u_a23_mem/stack_mem_reg[17][2]  ( .D(\u_a23_mem/n19514 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[17][2] ) );
  DFF \u_a23_mem/stack_mem_reg[17][3]  ( .D(\u_a23_mem/n19513 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[17][3] ) );
  DFF \u_a23_mem/stack_mem_reg[17][4]  ( .D(\u_a23_mem/n19512 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[17][4] ) );
  DFF \u_a23_mem/stack_mem_reg[17][5]  ( .D(\u_a23_mem/n19511 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[17][5] ) );
  DFF \u_a23_mem/stack_mem_reg[17][6]  ( .D(\u_a23_mem/n19510 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[17][6] ) );
  DFF \u_a23_mem/stack_mem_reg[17][7]  ( .D(\u_a23_mem/n19509 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[17][7] ) );
  DFF \u_a23_mem/stack_mem_reg[18][0]  ( .D(\u_a23_mem/n19508 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[18][0] ) );
  DFF \u_a23_mem/stack_mem_reg[18][1]  ( .D(\u_a23_mem/n19507 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[18][1] ) );
  DFF \u_a23_mem/stack_mem_reg[18][2]  ( .D(\u_a23_mem/n19506 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[18][2] ) );
  DFF \u_a23_mem/stack_mem_reg[18][3]  ( .D(\u_a23_mem/n19505 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[18][3] ) );
  DFF \u_a23_mem/stack_mem_reg[18][4]  ( .D(\u_a23_mem/n19504 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[18][4] ) );
  DFF \u_a23_mem/stack_mem_reg[18][5]  ( .D(\u_a23_mem/n19503 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[18][5] ) );
  DFF \u_a23_mem/stack_mem_reg[18][6]  ( .D(\u_a23_mem/n19502 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[18][6] ) );
  DFF \u_a23_mem/stack_mem_reg[18][7]  ( .D(\u_a23_mem/n19501 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[18][7] ) );
  DFF \u_a23_mem/stack_mem_reg[19][0]  ( .D(\u_a23_mem/n19500 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[19][0] ) );
  DFF \u_a23_mem/stack_mem_reg[19][1]  ( .D(\u_a23_mem/n19499 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[19][1] ) );
  DFF \u_a23_mem/stack_mem_reg[19][2]  ( .D(\u_a23_mem/n19498 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[19][2] ) );
  DFF \u_a23_mem/stack_mem_reg[19][3]  ( .D(\u_a23_mem/n19497 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[19][3] ) );
  DFF \u_a23_mem/stack_mem_reg[19][4]  ( .D(\u_a23_mem/n19496 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[19][4] ) );
  DFF \u_a23_mem/stack_mem_reg[19][5]  ( .D(\u_a23_mem/n19495 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[19][5] ) );
  DFF \u_a23_mem/stack_mem_reg[19][6]  ( .D(\u_a23_mem/n19494 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[19][6] ) );
  DFF \u_a23_mem/stack_mem_reg[19][7]  ( .D(\u_a23_mem/n19493 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[19][7] ) );
  DFF \u_a23_mem/stack_mem_reg[20][0]  ( .D(\u_a23_mem/n19492 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[20][0] ) );
  DFF \u_a23_mem/stack_mem_reg[20][1]  ( .D(\u_a23_mem/n19491 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[20][1] ) );
  DFF \u_a23_mem/stack_mem_reg[20][2]  ( .D(\u_a23_mem/n19490 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[20][2] ) );
  DFF \u_a23_mem/stack_mem_reg[20][3]  ( .D(\u_a23_mem/n19489 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[20][3] ) );
  DFF \u_a23_mem/stack_mem_reg[20][4]  ( .D(\u_a23_mem/n19488 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[20][4] ) );
  DFF \u_a23_mem/stack_mem_reg[20][5]  ( .D(\u_a23_mem/n19487 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[20][5] ) );
  DFF \u_a23_mem/stack_mem_reg[20][6]  ( .D(\u_a23_mem/n19486 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[20][6] ) );
  DFF \u_a23_mem/stack_mem_reg[20][7]  ( .D(\u_a23_mem/n19485 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[20][7] ) );
  DFF \u_a23_mem/stack_mem_reg[21][0]  ( .D(\u_a23_mem/n19484 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[21][0] ) );
  DFF \u_a23_mem/stack_mem_reg[21][1]  ( .D(\u_a23_mem/n19483 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[21][1] ) );
  DFF \u_a23_mem/stack_mem_reg[21][2]  ( .D(\u_a23_mem/n19482 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[21][2] ) );
  DFF \u_a23_mem/stack_mem_reg[21][3]  ( .D(\u_a23_mem/n19481 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[21][3] ) );
  DFF \u_a23_mem/stack_mem_reg[21][4]  ( .D(\u_a23_mem/n19480 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[21][4] ) );
  DFF \u_a23_mem/stack_mem_reg[21][5]  ( .D(\u_a23_mem/n19479 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[21][5] ) );
  DFF \u_a23_mem/stack_mem_reg[21][6]  ( .D(\u_a23_mem/n19478 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[21][6] ) );
  DFF \u_a23_mem/stack_mem_reg[21][7]  ( .D(\u_a23_mem/n19477 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[21][7] ) );
  DFF \u_a23_mem/stack_mem_reg[22][0]  ( .D(\u_a23_mem/n19476 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[22][0] ) );
  DFF \u_a23_mem/stack_mem_reg[22][1]  ( .D(\u_a23_mem/n19475 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[22][1] ) );
  DFF \u_a23_mem/stack_mem_reg[22][2]  ( .D(\u_a23_mem/n19474 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[22][2] ) );
  DFF \u_a23_mem/stack_mem_reg[22][3]  ( .D(\u_a23_mem/n19473 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[22][3] ) );
  DFF \u_a23_mem/stack_mem_reg[22][4]  ( .D(\u_a23_mem/n19472 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[22][4] ) );
  DFF \u_a23_mem/stack_mem_reg[22][5]  ( .D(\u_a23_mem/n19471 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[22][5] ) );
  DFF \u_a23_mem/stack_mem_reg[22][6]  ( .D(\u_a23_mem/n19470 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[22][6] ) );
  DFF \u_a23_mem/stack_mem_reg[22][7]  ( .D(\u_a23_mem/n19469 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[22][7] ) );
  DFF \u_a23_mem/stack_mem_reg[23][0]  ( .D(\u_a23_mem/n19468 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[23][0] ) );
  DFF \u_a23_mem/stack_mem_reg[23][1]  ( .D(\u_a23_mem/n19467 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[23][1] ) );
  DFF \u_a23_mem/stack_mem_reg[23][2]  ( .D(\u_a23_mem/n19466 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[23][2] ) );
  DFF \u_a23_mem/stack_mem_reg[23][3]  ( .D(\u_a23_mem/n19465 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[23][3] ) );
  DFF \u_a23_mem/stack_mem_reg[23][4]  ( .D(\u_a23_mem/n19464 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[23][4] ) );
  DFF \u_a23_mem/stack_mem_reg[23][5]  ( .D(\u_a23_mem/n19463 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[23][5] ) );
  DFF \u_a23_mem/stack_mem_reg[23][6]  ( .D(\u_a23_mem/n19462 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[23][6] ) );
  DFF \u_a23_mem/stack_mem_reg[23][7]  ( .D(\u_a23_mem/n19461 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[23][7] ) );
  DFF \u_a23_mem/stack_mem_reg[24][0]  ( .D(\u_a23_mem/n19460 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[24][0] ) );
  DFF \u_a23_mem/stack_mem_reg[24][1]  ( .D(\u_a23_mem/n19459 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[24][1] ) );
  DFF \u_a23_mem/stack_mem_reg[24][2]  ( .D(\u_a23_mem/n19458 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[24][2] ) );
  DFF \u_a23_mem/stack_mem_reg[24][3]  ( .D(\u_a23_mem/n19457 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[24][3] ) );
  DFF \u_a23_mem/stack_mem_reg[24][4]  ( .D(\u_a23_mem/n19456 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[24][4] ) );
  DFF \u_a23_mem/stack_mem_reg[24][5]  ( .D(\u_a23_mem/n19455 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[24][5] ) );
  DFF \u_a23_mem/stack_mem_reg[24][6]  ( .D(\u_a23_mem/n19454 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[24][6] ) );
  DFF \u_a23_mem/stack_mem_reg[24][7]  ( .D(\u_a23_mem/n19453 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[24][7] ) );
  DFF \u_a23_mem/stack_mem_reg[25][0]  ( .D(\u_a23_mem/n19452 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[25][0] ) );
  DFF \u_a23_mem/stack_mem_reg[25][1]  ( .D(\u_a23_mem/n19451 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[25][1] ) );
  DFF \u_a23_mem/stack_mem_reg[25][2]  ( .D(\u_a23_mem/n19450 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[25][2] ) );
  DFF \u_a23_mem/stack_mem_reg[25][3]  ( .D(\u_a23_mem/n19449 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[25][3] ) );
  DFF \u_a23_mem/stack_mem_reg[25][4]  ( .D(\u_a23_mem/n19448 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[25][4] ) );
  DFF \u_a23_mem/stack_mem_reg[25][5]  ( .D(\u_a23_mem/n19447 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[25][5] ) );
  DFF \u_a23_mem/stack_mem_reg[25][6]  ( .D(\u_a23_mem/n19446 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[25][6] ) );
  DFF \u_a23_mem/stack_mem_reg[25][7]  ( .D(\u_a23_mem/n19445 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[25][7] ) );
  DFF \u_a23_mem/stack_mem_reg[26][0]  ( .D(\u_a23_mem/n19444 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[26][0] ) );
  DFF \u_a23_mem/stack_mem_reg[26][1]  ( .D(\u_a23_mem/n19443 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[26][1] ) );
  DFF \u_a23_mem/stack_mem_reg[26][2]  ( .D(\u_a23_mem/n19442 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[26][2] ) );
  DFF \u_a23_mem/stack_mem_reg[26][3]  ( .D(\u_a23_mem/n19441 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[26][3] ) );
  DFF \u_a23_mem/stack_mem_reg[26][4]  ( .D(\u_a23_mem/n19440 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[26][4] ) );
  DFF \u_a23_mem/stack_mem_reg[26][5]  ( .D(\u_a23_mem/n19439 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[26][5] ) );
  DFF \u_a23_mem/stack_mem_reg[26][6]  ( .D(\u_a23_mem/n19438 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[26][6] ) );
  DFF \u_a23_mem/stack_mem_reg[26][7]  ( .D(\u_a23_mem/n19437 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[26][7] ) );
  DFF \u_a23_mem/stack_mem_reg[27][0]  ( .D(\u_a23_mem/n19436 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[27][0] ) );
  DFF \u_a23_mem/stack_mem_reg[27][1]  ( .D(\u_a23_mem/n19435 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[27][1] ) );
  DFF \u_a23_mem/stack_mem_reg[27][2]  ( .D(\u_a23_mem/n19434 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[27][2] ) );
  DFF \u_a23_mem/stack_mem_reg[27][3]  ( .D(\u_a23_mem/n19433 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[27][3] ) );
  DFF \u_a23_mem/stack_mem_reg[27][4]  ( .D(\u_a23_mem/n19432 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[27][4] ) );
  DFF \u_a23_mem/stack_mem_reg[27][5]  ( .D(\u_a23_mem/n19431 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[27][5] ) );
  DFF \u_a23_mem/stack_mem_reg[27][6]  ( .D(\u_a23_mem/n19430 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[27][6] ) );
  DFF \u_a23_mem/stack_mem_reg[27][7]  ( .D(\u_a23_mem/n19429 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[27][7] ) );
  DFF \u_a23_mem/stack_mem_reg[28][0]  ( .D(\u_a23_mem/n19428 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[28][0] ) );
  DFF \u_a23_mem/stack_mem_reg[28][1]  ( .D(\u_a23_mem/n19427 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[28][1] ) );
  DFF \u_a23_mem/stack_mem_reg[28][2]  ( .D(\u_a23_mem/n19426 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[28][2] ) );
  DFF \u_a23_mem/stack_mem_reg[28][3]  ( .D(\u_a23_mem/n19425 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[28][3] ) );
  DFF \u_a23_mem/stack_mem_reg[28][4]  ( .D(\u_a23_mem/n19424 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[28][4] ) );
  DFF \u_a23_mem/stack_mem_reg[28][5]  ( .D(\u_a23_mem/n19423 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[28][5] ) );
  DFF \u_a23_mem/stack_mem_reg[28][6]  ( .D(\u_a23_mem/n19422 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[28][6] ) );
  DFF \u_a23_mem/stack_mem_reg[28][7]  ( .D(\u_a23_mem/n19421 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[28][7] ) );
  DFF \u_a23_mem/stack_mem_reg[29][0]  ( .D(\u_a23_mem/n19420 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[29][0] ) );
  DFF \u_a23_mem/stack_mem_reg[29][1]  ( .D(\u_a23_mem/n19419 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[29][1] ) );
  DFF \u_a23_mem/stack_mem_reg[29][2]  ( .D(\u_a23_mem/n19418 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[29][2] ) );
  DFF \u_a23_mem/stack_mem_reg[29][3]  ( .D(\u_a23_mem/n19417 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[29][3] ) );
  DFF \u_a23_mem/stack_mem_reg[29][4]  ( .D(\u_a23_mem/n19416 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[29][4] ) );
  DFF \u_a23_mem/stack_mem_reg[29][5]  ( .D(\u_a23_mem/n19415 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[29][5] ) );
  DFF \u_a23_mem/stack_mem_reg[29][6]  ( .D(\u_a23_mem/n19414 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[29][6] ) );
  DFF \u_a23_mem/stack_mem_reg[29][7]  ( .D(\u_a23_mem/n19413 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[29][7] ) );
  DFF \u_a23_mem/stack_mem_reg[30][0]  ( .D(\u_a23_mem/n19412 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[30][0] ) );
  DFF \u_a23_mem/stack_mem_reg[30][1]  ( .D(\u_a23_mem/n19411 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[30][1] ) );
  DFF \u_a23_mem/stack_mem_reg[30][2]  ( .D(\u_a23_mem/n19410 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[30][2] ) );
  DFF \u_a23_mem/stack_mem_reg[30][3]  ( .D(\u_a23_mem/n19409 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[30][3] ) );
  DFF \u_a23_mem/stack_mem_reg[30][4]  ( .D(\u_a23_mem/n19408 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[30][4] ) );
  DFF \u_a23_mem/stack_mem_reg[30][5]  ( .D(\u_a23_mem/n19407 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[30][5] ) );
  DFF \u_a23_mem/stack_mem_reg[30][6]  ( .D(\u_a23_mem/n19406 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[30][6] ) );
  DFF \u_a23_mem/stack_mem_reg[30][7]  ( .D(\u_a23_mem/n19405 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[30][7] ) );
  DFF \u_a23_mem/stack_mem_reg[31][0]  ( .D(\u_a23_mem/n19404 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[31][0] ) );
  DFF \u_a23_mem/stack_mem_reg[31][1]  ( .D(\u_a23_mem/n19403 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[31][1] ) );
  DFF \u_a23_mem/stack_mem_reg[31][2]  ( .D(\u_a23_mem/n19402 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[31][2] ) );
  DFF \u_a23_mem/stack_mem_reg[31][3]  ( .D(\u_a23_mem/n19401 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[31][3] ) );
  DFF \u_a23_mem/stack_mem_reg[31][4]  ( .D(\u_a23_mem/n19400 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[31][4] ) );
  DFF \u_a23_mem/stack_mem_reg[31][5]  ( .D(\u_a23_mem/n19399 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[31][5] ) );
  DFF \u_a23_mem/stack_mem_reg[31][6]  ( .D(\u_a23_mem/n19398 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[31][6] ) );
  DFF \u_a23_mem/stack_mem_reg[31][7]  ( .D(\u_a23_mem/n19397 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_mem/stack_mem[31][7] ) );
  DFF \u_a23_core/u_decode/o_imm32_reg[9]  ( .D(
        \u_a23_core/u_decode/imm32_nxt[9] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm32[9] ) );
  DFF \u_a23_core/u_decode/o_imm32_reg[7]  ( .D(
        \u_a23_core/u_decode/imm32_nxt[7] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm32[7] ) );
  DFF \u_a23_core/u_decode/o_imm32_reg[5]  ( .D(
        \u_a23_core/u_decode/imm32_nxt[5] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm32[5] ) );
  DFF \u_a23_core/u_decode/o_imm32_reg[3]  ( .D(
        \u_a23_core/u_decode/imm32_nxt[3] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm32[3] ) );
  DFF \u_a23_core/u_decode/o_imm32_reg[31]  ( .D(
        \u_a23_core/u_decode/imm32_nxt[31] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm32[31] ) );
  DFF \u_a23_core/u_decode/o_imm32_reg[29]  ( .D(
        \u_a23_core/u_decode/imm32_nxt[29] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm32[29] ) );
  DFF \u_a23_core/u_decode/o_imm32_reg[27]  ( .D(
        \u_a23_core/u_decode/imm32_nxt[27] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm32[27] ) );
  DFF \u_a23_core/u_decode/o_imm32_reg[25]  ( .D(
        \u_a23_core/u_decode/imm32_nxt[25] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm32[25] ) );
  DFF \u_a23_core/u_decode/o_imm32_reg[23]  ( .D(
        \u_a23_core/u_decode/imm32_nxt[23] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm32[23] ) );
  DFF \u_a23_core/u_decode/o_imm32_reg[21]  ( .D(
        \u_a23_core/u_decode/imm32_nxt[21] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm32[21] ) );
  DFF \u_a23_core/u_decode/o_imm32_reg[1]  ( .D(
        \u_a23_core/u_decode/imm32_nxt[1] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm32[1] ) );
  DFF \u_a23_core/u_decode/o_imm32_reg[19]  ( .D(
        \u_a23_core/u_decode/imm32_nxt[19] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm32[19] ) );
  DFF \u_a23_core/u_decode/o_imm32_reg[17]  ( .D(
        \u_a23_core/u_decode/imm32_nxt[17] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm32[17] ) );
  DFF \u_a23_core/u_decode/o_imm32_reg[15]  ( .D(
        \u_a23_core/u_decode/imm32_nxt[15] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm32[15] ) );
  DFF \u_a23_core/u_decode/o_imm32_reg[13]  ( .D(
        \u_a23_core/u_decode/imm32_nxt[13] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm32[13] ) );
  DFF \u_a23_core/u_decode/o_imm32_reg[11]  ( .D(
        \u_a23_core/u_decode/imm32_nxt[11] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm32[11] ) );
  DFF \u_a23_core/u_decode/address_sel_r_reg[0]  ( .D(
        \u_a23_core/u_decode/address_sel_nxt[0] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\u_a23_core/address_sel[0] ) );
  DFF \u_a23_core/u_decode/address_sel_r_reg[2]  ( .D(
        \u_a23_core/u_decode/address_sel_nxt[2] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\u_a23_core/address_sel[2] ) );
  DFF \u_a23_core/u_decode/o_write_data_wen_reg  ( .D(
        \u_a23_core/u_decode/write_data_wen_nxt ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\u_a23_core/write_data_wen ) );
  DFF \u_a23_core/u_decode/o_reg_bank_wen_reg[0]  ( .D(
        \u_a23_core/u_decode/N1089 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/reg_bank_wen[0] ) );
  DFF \u_a23_core/u_decode/o_reg_bank_wen_reg[4]  ( .D(
        \u_a23_core/u_decode/n1508 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/reg_bank_wen[4] ) );
  DFF \u_a23_core/u_decode/o_reg_bank_wen_reg[12]  ( .D(
        \u_a23_core/u_decode/n1502 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/reg_bank_wen[12] ) );
  DFF \u_a23_core/u_decode/o_reg_bank_wen_reg[8]  ( .D(
        \u_a23_core/u_decode/n1498 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/reg_bank_wen[8] ) );
  DFF \u_a23_core/u_decode/o_reg_bank_wen_reg[7]  ( .D(
        \u_a23_core/u_decode/n1511 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/reg_bank_wen[7] ) );
  DFF \u_a23_core/u_decode/o_reg_bank_wen_reg[3]  ( .D(
        \u_a23_core/u_decode/n1507 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/reg_bank_wen[3] ) );
  DFF \u_a23_core/u_decode/o_reg_bank_wen_reg[11]  ( .D(
        \u_a23_core/u_decode/n1501 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/reg_bank_wen[11] ) );
  DFF \u_a23_core/u_decode/o_reg_bank_wen_reg[6]  ( .D(
        \u_a23_core/u_decode/n1510 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/reg_bank_wen[6] ) );
  DFF \u_a23_core/u_decode/o_reg_bank_wen_reg[2]  ( .D(
        \u_a23_core/u_decode/n1506 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/reg_bank_wen[2] ) );
  DFF \u_a23_core/u_decode/o_reg_bank_wen_reg[14]  ( .D(
        \u_a23_core/u_decode/n1504 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/reg_bank_wen[14] ) );
  DFF \u_a23_core/u_decode/o_reg_bank_wen_reg[10]  ( .D(
        \u_a23_core/u_decode/n1500 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/reg_bank_wen[10] ) );
  DFF \u_a23_core/u_decode/o_reg_bank_wen_reg[5]  ( .D(
        \u_a23_core/u_decode/n1509 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/reg_bank_wen[5] ) );
  DFF \u_a23_core/u_decode/o_reg_bank_wen_reg[1]  ( .D(
        \u_a23_core/u_decode/n1505 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/reg_bank_wen[1] ) );
  DFF \u_a23_core/u_decode/o_reg_bank_wen_reg[13]  ( .D(
        \u_a23_core/u_decode/n1503 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/reg_bank_wen[13] ) );
  DFF \u_a23_core/u_decode/o_reg_bank_wen_reg[9]  ( .D(
        \u_a23_core/u_decode/n1499 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/reg_bank_wen[9] ) );
  DFF \u_a23_core/u_decode/o_barrel_shift_data_sel_reg[0]  ( .D(
        \u_a23_core/u_decode/barrel_shift_data_sel_nxt[0] ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\u_a23_core/barrel_shift_data_sel[0] ) );
  DFF \u_a23_core/u_decode/saved_current_instruction_reg[27]  ( .D(
        \u_a23_core/u_decode/n1481 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/saved_current_instruction[27] ) );
  DFF \u_a23_core/u_decode/o_status_bits_sel_reg[2]  ( .D(
        \u_a23_core/u_decode/status_bits_sel_nxt[2] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/status_bits_sel[2] ) );
  DFF \u_a23_core/u_decode/o_status_bits_sel_reg[0]  ( .D(
        \u_a23_core/u_decode/status_bits_sel_nxt_0 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/status_bits_sel[0] ) );
  DFF \u_a23_core/u_decode/o_rds_sel_reg[0]  ( .D(\u_a23_core/rds_sel_nxt[0] ), 
        .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/rds_sel[0] ) );
  DFF \u_a23_core/u_decode/o_rds_sel_reg[1]  ( .D(\u_a23_core/rds_sel_nxt[1] ), 
        .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/rds_sel[1] ) );
  DFF \u_a23_core/u_decode/o_rds_sel_reg[2]  ( .D(\u_a23_core/rds_sel_nxt[2] ), 
        .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/rds_sel[2] ) );
  DFF \u_a23_core/u_decode/o_rds_sel_reg[3]  ( .D(\u_a23_core/rds_sel_nxt[3] ), 
        .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/rds_sel[3] ) );
  DFF \u_a23_core/u_decode/o_alu_function_reg[7]  ( .D(
        \u_a23_core/u_decode/alu_function_nxt[7] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\u_a23_core/alu_function[7] ) );
  DFF \u_a23_core/u_decode/o_alu_function_reg[6]  ( .D(
        \u_a23_core/u_decode/alu_function_nxt[6] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\u_a23_core/alu_function[6] ) );
  DFF \u_a23_core/u_decode/o_alu_function_reg[5]  ( .D(
        \u_a23_core/u_decode/alu_function_nxt[5] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\u_a23_core/alu_function[5] ) );
  DFF \u_a23_core/u_decode/o_alu_function_reg[0]  ( .D(
        \u_a23_core/u_decode/alu_function_nxt[0] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\u_a23_core/alu_function[0] ) );
  DFF \u_a23_core/u_decode/pc_sel_r_reg[0]  ( .D(
        \u_a23_core/u_decode/pc_sel_nxt[0] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/pc_sel[0] ) );
  DFF \u_a23_core/u_decode/o_alu_function_reg[1]  ( .D(
        \u_a23_core/u_decode/alu_function_nxt[1] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\u_a23_core/alu_function[1] ) );
  DFF \u_a23_core/u_decode/o_alu_function_reg[2]  ( .D(
        \u_a23_core/u_decode/alu_function_nxt[2] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\u_a23_core/alu_function[2] ) );
  DFF \u_a23_core/u_decode/o_alu_function_reg[3]  ( .D(
        \u_a23_core/u_decode/alu_function_nxt[3] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\u_a23_core/alu_function[3] ) );
  DFF \u_a23_core/u_decode/o_alu_function_reg[4]  ( .D(
        \u_a23_core/u_decode/alu_function_nxt[4] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\u_a23_core/alu_function[4] ) );
  DFF \u_a23_core/u_decode/o_alu_function_reg[8]  ( .D(
        \u_a23_core/u_decode/alu_function_nxt[8] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\u_a23_core/alu_function[8] ) );
  DFF \u_a23_core/u_decode/o_shift_imm_zero_reg  ( .D(
        \u_a23_core/u_decode/shift_imm_zero_nxt ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\u_a23_core/shift_imm_zero ) );
  DFF \u_a23_core/u_decode/o_barrel_shift_amount_sel_reg[0]  ( .D(
        \u_a23_core/u_decode/barrel_shift_amount_sel_nxt[0] ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_core/barrel_shift_amount_sel[0] ) );
  DFF \u_a23_core/u_decode/o_barrel_shift_amount_sel_reg[1]  ( .D(
        \u_a23_core/u_decode/barrel_shift_amount_sel_nxt[1] ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_core/barrel_shift_amount_sel[1] ) );
  DFF \u_a23_core/u_decode/o_barrel_shift_data_sel_reg[1]  ( .D(
        \u_a23_core/u_decode/barrel_shift_data_sel_nxt[1] ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\u_a23_core/barrel_shift_data_sel[1] ) );
  DFF \u_a23_core/u_decode/o_barrel_shift_function_reg[0]  ( .D(
        \u_a23_core/u_decode/barrel_shift_function_nxt[0] ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\u_a23_core/barrel_shift_function[0] ) );
  DFF \u_a23_core/u_decode/o_barrel_shift_function_reg[1]  ( .D(
        \u_a23_core/u_decode/barrel_shift_function_nxt[1] ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\u_a23_core/barrel_shift_function[1] ) );
  DFF \u_a23_core/u_decode/o_use_carry_in_reg  ( .D(
        \u_a23_core/u_decode/use_carry_in_nxt ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/use_carry_in ) );
  DFF \u_a23_core/u_decode/o_status_bits_flags_wen_reg  ( .D(
        \u_a23_core/u_decode/status_bits_flags_wen_nxt ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/status_bits_flags_wen ) );
  DFF \u_a23_core/u_decode/o_imm32_reg[2]  ( .D(
        \u_a23_core/u_decode/imm32_nxt[2] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm32[2] ) );
  DFF \u_a23_core/u_decode/o_imm32_reg[4]  ( .D(
        \u_a23_core/u_decode/imm32_nxt[4] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm32[4] ) );
  DFF \u_a23_core/u_decode/o_imm32_reg[6]  ( .D(
        \u_a23_core/u_decode/imm32_nxt[6] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm32[6] ) );
  DFF \u_a23_core/u_decode/o_imm32_reg[8]  ( .D(
        \u_a23_core/u_decode/imm32_nxt[8] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm32[8] ) );
  DFF \u_a23_core/u_decode/o_imm32_reg[20]  ( .D(
        \u_a23_core/u_decode/imm32_nxt[20] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm32[20] ) );
  DFF \u_a23_core/u_decode/o_imm32_reg[18]  ( .D(
        \u_a23_core/u_decode/imm32_nxt[18] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm32[18] ) );
  DFF \u_a23_core/u_decode/o_imm32_reg[0]  ( .D(
        \u_a23_core/u_decode/imm32_nxt[0] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm32[0] ) );
  DFF \u_a23_core/u_decode/o_imm32_reg[30]  ( .D(
        \u_a23_core/u_decode/imm32_nxt[30] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm32[30] ) );
  DFF \u_a23_core/u_decode/o_imm32_reg[28]  ( .D(
        \u_a23_core/u_decode/imm32_nxt[28] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm32[28] ) );
  DFF \u_a23_core/u_decode/o_imm32_reg[26]  ( .D(
        \u_a23_core/u_decode/imm32_nxt[26] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm32[26] ) );
  DFF \u_a23_core/u_decode/o_imm32_reg[10]  ( .D(
        \u_a23_core/u_decode/imm32_nxt[10] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm32[10] ) );
  DFF \u_a23_core/u_decode/o_imm32_reg[12]  ( .D(
        \u_a23_core/u_decode/imm32_nxt[12] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm32[12] ) );
  DFF \u_a23_core/u_decode/o_imm32_reg[14]  ( .D(
        \u_a23_core/u_decode/imm32_nxt[14] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm32[14] ) );
  DFF \u_a23_core/u_decode/o_imm32_reg[16]  ( .D(
        \u_a23_core/u_decode/imm32_nxt[16] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm32[16] ) );
  DFF \u_a23_core/u_decode/o_imm32_reg[22]  ( .D(
        \u_a23_core/u_decode/imm32_nxt[22] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm32[22] ) );
  DFF \u_a23_core/u_decode/o_imm32_reg[24]  ( .D(
        \u_a23_core/u_decode/imm32_nxt[24] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm32[24] ) );
  DFF \u_a23_core/u_decode/address_sel_r_reg[3]  ( .D(
        \u_a23_core/u_decode/pc_sel_nxt[1] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/address_sel[3] ) );
  DFF \u_a23_core/u_decode/pc_sel_r_reg[1]  ( .D(
        \u_a23_core/u_decode/pc_sel_nxt[1] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/pc_sel[1] ) );
  DFF \u_a23_core/u_decode/o_rn_sel_reg[0]  ( .D(\u_a23_core/rn_sel_nxt[0] ), 
        .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/rn_sel[0] ) );
  DFF \u_a23_core/u_decode/o_rn_sel_reg[1]  ( .D(\u_a23_core/rn_sel_nxt[1] ), 
        .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/rn_sel[1] ) );
  DFF \u_a23_core/u_decode/o_rn_sel_reg[3]  ( .D(\u_a23_core/rn_sel_nxt[3] ), 
        .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/rn_sel[3] ) );
  DFF \u_a23_core/u_decode/o_rn_sel_reg[2]  ( .D(\u_a23_core/rn_sel_nxt[2] ), 
        .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/rn_sel[2] ) );
  DFF \u_a23_core/u_decode/o_reg_write_sel_reg[0]  ( .D(
        \u_a23_core/u_decode/reg_write_sel_nxt[0] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\u_a23_core/reg_write_sel[0] ) );
  DFF \u_a23_core/u_decode/condition_r_reg[3]  ( .D(
        \u_a23_core/u_decode/n1427 ), .CLK(clk), .RST(rst), .I(1'b1), .Q(
        \u_a23_core/condition[3] ) );
  DFF \u_a23_core/u_decode/condition_r_reg[2]  ( .D(
        \u_a23_core/u_decode/n1429 ), .CLK(clk), .RST(rst), .I(1'b1), .Q(
        \u_a23_core/condition[2] ) );
  DFF \u_a23_core/u_decode/condition_r_reg[1]  ( .D(
        \u_a23_core/u_decode/n1431 ), .CLK(clk), .RST(rst), .I(1'b1), .Q(
        \u_a23_core/condition[1] ) );
  DFF \u_a23_core/u_decode/condition_r_reg[0]  ( .D(
        \u_a23_core/u_decode/n1433 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/condition[0] ) );
  DFF \u_a23_core/u_decode/saved_current_instruction_reg[15]  ( .D(
        \u_a23_core/u_decode/n1465 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/saved_current_instruction[15] ) );
  DFF \u_a23_core/u_decode/mtrans_reg_d2_reg[0]  ( .D(
        \u_a23_core/u_decode/mtrans_reg_d1[0] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_decode/mtrans_reg_d2[0] ) );
  DFF \u_a23_core/u_decode/mtrans_reg_d1_reg[0]  ( .D(
        \u_a23_core/u_decode/N384 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/mtrans_reg_d1[0] ) );
  DFF \u_a23_core/u_decode/saved_current_instruction_reg[14]  ( .D(
        \u_a23_core/u_decode/n1466 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/saved_current_instruction[14] ) );
  DFF \u_a23_core/u_decode/mtrans_reg_d2_reg[1]  ( .D(
        \u_a23_core/u_decode/mtrans_reg_d1[1] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_decode/mtrans_reg_d2[1] ) );
  DFF \u_a23_core/u_decode/mtrans_reg_d1_reg[1]  ( .D(
        \u_a23_core/u_decode/N348 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/mtrans_reg_d1[1] ) );
  DFF \u_a23_core/u_decode/saved_current_instruction_reg[13]  ( .D(
        \u_a23_core/u_decode/n1467 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/saved_current_instruction[13] ) );
  DFF \u_a23_core/u_decode/saved_current_instruction_reg[12]  ( .D(
        \u_a23_core/u_decode/n1468 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/saved_current_instruction[12] ) );
  DFF \u_a23_core/u_decode/mtrans_reg_d2_reg[2]  ( .D(
        \u_a23_core/u_decode/mtrans_reg_d1[2] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_decode/mtrans_reg_d2[2] ) );
  DFF \u_a23_core/u_decode/mtrans_reg_d1_reg[2]  ( .D(
        \u_a23_core/u_decode/N319 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/mtrans_reg_d1[2] ) );
  DFF \u_a23_core/u_decode/o_imm_shift_amount_reg[4]  ( .D(
        \u_a23_core/u_decode/instruction[11] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm_shift_amount[4] ) );
  DFF \u_a23_core/u_decode/saved_current_instruction_reg[11]  ( .D(
        \u_a23_core/u_decode/n1469 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/saved_current_instruction[11] ) );
  DFF \u_a23_core/u_decode/o_imm_shift_amount_reg[3]  ( .D(
        \u_a23_core/u_decode/instruction[10] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm_shift_amount[3] ) );
  DFF \u_a23_core/u_decode/saved_current_instruction_reg[10]  ( .D(
        \u_a23_core/u_decode/n1470 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/saved_current_instruction[10] ) );
  DFF \u_a23_core/u_decode/o_imm_shift_amount_reg[2]  ( .D(
        \u_a23_core/u_decode/instruction[9] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm_shift_amount[2] ) );
  DFF \u_a23_core/u_decode/saved_current_instruction_reg[9]  ( .D(
        \u_a23_core/u_decode/n1471 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/saved_current_instruction[9] ) );
  DFF \u_a23_core/u_decode/o_imm_shift_amount_reg[1]  ( .D(
        \u_a23_core/u_decode/instruction[8] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm_shift_amount[1] ) );
  DFF \u_a23_core/u_decode/saved_current_instruction_reg[8]  ( .D(
        \u_a23_core/u_decode/n1472 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/saved_current_instruction[8] ) );
  DFF \u_a23_core/u_decode/mtrans_reg_d2_reg[3]  ( .D(
        \u_a23_core/u_decode/mtrans_reg_d1[3] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_decode/mtrans_reg_d2[3] ) );
  DFF \u_a23_core/u_decode/mtrans_reg_d1_reg[3]  ( .D(
        \u_a23_core/u_decode/N298 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/mtrans_reg_d1[3] ) );
  DFF \u_a23_core/u_decode/o_multiply_function_reg[1]  ( .D(
        \u_a23_core/u_decode/n1493 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/multiply_function[1] ) );
  DFF \u_a23_core/u_decode/address_sel_r_reg[1]  ( .D(
        \u_a23_core/u_decode/address_sel_nxt[1] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\u_a23_core/address_sel[1] ) );
  DFF \u_a23_core/u_decode/o_multiply_function_reg[0]  ( .D(
        \u_a23_core/u_decode/n1494 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/multiply_function[0] ) );
  DFF \u_a23_core/u_decode/pre_fetch_instruction_reg[31]  ( .D(
        \u_a23_core/u_decode/n1434 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/pre_fetch_instruction[31] ) );
  DFF \u_a23_core/u_decode/pre_fetch_instruction_reg[30]  ( .D(
        \u_a23_core/u_decode/n1435 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/pre_fetch_instruction[30] ) );
  DFF \u_a23_core/u_decode/pre_fetch_instruction_reg[29]  ( .D(
        \u_a23_core/u_decode/n1436 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/pre_fetch_instruction[29] ) );
  DFF \u_a23_core/u_decode/pre_fetch_instruction_reg[28]  ( .D(
        \u_a23_core/u_decode/n1437 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/pre_fetch_instruction[28] ) );
  DFF \u_a23_core/u_decode/pre_fetch_instruction_reg[27]  ( .D(
        \u_a23_core/u_decode/n1438 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/pre_fetch_instruction[27] ) );
  DFF \u_a23_core/u_decode/saved_current_instruction_reg[26]  ( .D(
        \u_a23_core/u_decode/n1482 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/saved_current_instruction[26] ) );
  DFF \u_a23_core/u_decode/pre_fetch_instruction_reg[26]  ( .D(
        \u_a23_core/u_decode/n1439 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/pre_fetch_instruction[26] ) );
  DFF \u_a23_core/u_decode/saved_current_instruction_reg[25]  ( .D(
        \u_a23_core/u_decode/n1483 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/saved_current_instruction[25] ) );
  DFF \u_a23_core/u_decode/pre_fetch_instruction_reg[25]  ( .D(
        \u_a23_core/u_decode/n1440 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/pre_fetch_instruction[25] ) );
  DFF \u_a23_core/u_decode/saved_current_instruction_reg[24]  ( .D(
        \u_a23_core/u_decode/n1484 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/saved_current_instruction[24] ) );
  DFF \u_a23_core/u_decode/pre_fetch_instruction_reg[24]  ( .D(
        \u_a23_core/u_decode/n1441 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/pre_fetch_instruction[24] ) );
  DFF \u_a23_core/u_decode/saved_current_instruction_reg[23]  ( .D(
        \u_a23_core/u_decode/n1485 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/saved_current_instruction[23] ) );
  DFF \u_a23_core/u_decode/pre_fetch_instruction_reg[23]  ( .D(
        \u_a23_core/u_decode/n1442 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/pre_fetch_instruction[23] ) );
  DFF \u_a23_core/u_decode/saved_current_instruction_reg[22]  ( .D(
        \u_a23_core/u_decode/n1486 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/saved_current_instruction[22] ) );
  DFF \u_a23_core/u_decode/o_byte_enable_sel_reg[0]  ( .D(
        \u_a23_core/u_decode/byte_enable_sel_nxt[0] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/byte_enable_sel[0] ) );
  DFF \u_a23_core/u_decode/pre_fetch_instruction_reg[22]  ( .D(
        \u_a23_core/u_decode/n1443 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/pre_fetch_instruction[22] ) );
  DFF \u_a23_core/u_decode/saved_current_instruction_reg[21]  ( .D(
        \u_a23_core/u_decode/n1487 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/saved_current_instruction[21] ) );
  DFF \u_a23_core/u_decode/pre_fetch_instruction_reg[21]  ( .D(
        \u_a23_core/u_decode/n1444 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/pre_fetch_instruction[21] ) );
  DFF \u_a23_core/u_decode/saved_current_instruction_reg[20]  ( .D(
        \u_a23_core/u_decode/n1488 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/saved_current_instruction[20] ) );
  DFF \u_a23_core/u_decode/pre_fetch_instruction_reg[20]  ( .D(
        \u_a23_core/u_decode/n1445 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/pre_fetch_instruction[20] ) );
  DFF \u_a23_core/u_decode/saved_current_instruction_reg[19]  ( .D(
        \u_a23_core/u_decode/n1489 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/saved_current_instruction[19] ) );
  DFF \u_a23_core/u_decode/pre_fetch_instruction_reg[19]  ( .D(
        \u_a23_core/u_decode/n1446 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/pre_fetch_instruction[19] ) );
  DFF \u_a23_core/u_decode/saved_current_instruction_reg[18]  ( .D(
        \u_a23_core/u_decode/n1490 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/saved_current_instruction[18] ) );
  DFF \u_a23_core/u_decode/pre_fetch_instruction_reg[18]  ( .D(
        \u_a23_core/u_decode/n1447 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/pre_fetch_instruction[18] ) );
  DFF \u_a23_core/u_decode/saved_current_instruction_reg[17]  ( .D(
        \u_a23_core/u_decode/n1491 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/saved_current_instruction[17] ) );
  DFF \u_a23_core/u_decode/pre_fetch_instruction_reg[17]  ( .D(
        \u_a23_core/u_decode/n1448 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/pre_fetch_instruction[17] ) );
  DFF \u_a23_core/u_decode/saved_current_instruction_reg[16]  ( .D(
        \u_a23_core/u_decode/n1492 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/saved_current_instruction[16] ) );
  DFF \u_a23_core/u_decode/pre_fetch_instruction_reg[16]  ( .D(
        \u_a23_core/u_decode/n1449 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/pre_fetch_instruction[16] ) );
  DFF \u_a23_core/u_decode/pre_fetch_instruction_reg[15]  ( .D(
        \u_a23_core/u_decode/n1450 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/pre_fetch_instruction[15] ) );
  DFF \u_a23_core/u_decode/pre_fetch_instruction_reg[14]  ( .D(
        \u_a23_core/u_decode/n1451 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/pre_fetch_instruction[14] ) );
  DFF \u_a23_core/u_decode/pre_fetch_instruction_reg[13]  ( .D(
        \u_a23_core/u_decode/n1452 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/pre_fetch_instruction[13] ) );
  DFF \u_a23_core/u_decode/pre_fetch_instruction_reg[12]  ( .D(
        \u_a23_core/u_decode/n1453 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/pre_fetch_instruction[12] ) );
  DFF \u_a23_core/u_decode/pre_fetch_instruction_reg[11]  ( .D(
        \u_a23_core/u_decode/n1454 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/pre_fetch_instruction[11] ) );
  DFF \u_a23_core/u_decode/pre_fetch_instruction_reg[10]  ( .D(
        \u_a23_core/u_decode/n1455 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/pre_fetch_instruction[10] ) );
  DFF \u_a23_core/u_decode/pre_fetch_instruction_reg[9]  ( .D(
        \u_a23_core/u_decode/n1456 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/pre_fetch_instruction[9] ) );
  DFF \u_a23_core/u_decode/pre_fetch_instruction_reg[8]  ( .D(
        \u_a23_core/u_decode/n1457 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/pre_fetch_instruction[8] ) );
  DFF \u_a23_core/u_decode/pre_fetch_instruction_reg[7]  ( .D(
        \u_a23_core/u_decode/n1458 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/pre_fetch_instruction[7] ) );
  DFF \u_a23_core/u_decode/saved_current_instruction_reg[6]  ( .D(
        \u_a23_core/u_decode/n1474 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/saved_current_instruction[6] ) );
  DFF \u_a23_core/u_decode/pre_fetch_instruction_reg[6]  ( .D(
        \u_a23_core/u_decode/n1459 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/pre_fetch_instruction[6] ) );
  DFF \u_a23_core/u_decode/saved_current_instruction_reg[5]  ( .D(
        \u_a23_core/u_decode/n1475 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/saved_current_instruction[5] ) );
  DFF \u_a23_core/u_decode/pre_fetch_instruction_reg[5]  ( .D(
        \u_a23_core/u_decode/n1460 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/pre_fetch_instruction[5] ) );
  DFF \u_a23_core/u_decode/saved_current_instruction_reg[4]  ( .D(
        \u_a23_core/u_decode/n1476 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/saved_current_instruction[4] ) );
  DFF \u_a23_core/u_decode/pre_fetch_instruction_reg[4]  ( .D(
        \u_a23_core/u_decode/n1461 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/pre_fetch_instruction[4] ) );
  DFF \u_a23_core/u_decode/saved_current_instruction_reg[3]  ( .D(
        \u_a23_core/u_decode/n1477 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/saved_current_instruction[3] ) );
  DFF \u_a23_core/u_decode/o_rm_sel_reg[3]  ( .D(\u_a23_core/rm_sel_nxt[3] ), 
        .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/rm_sel[3] ) );
  DFF \u_a23_core/u_decode/pre_fetch_instruction_reg[3]  ( .D(
        \u_a23_core/u_decode/n1462 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/pre_fetch_instruction[3] ) );
  DFF \u_a23_core/u_decode/saved_current_instruction_reg[2]  ( .D(
        \u_a23_core/u_decode/n1478 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/saved_current_instruction[2] ) );
  DFF \u_a23_core/u_decode/o_rm_sel_reg[2]  ( .D(\u_a23_core/rm_sel_nxt[2] ), 
        .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/rm_sel[2] ) );
  DFF \u_a23_core/u_decode/pre_fetch_instruction_reg[2]  ( .D(
        \u_a23_core/u_decode/n1463 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/pre_fetch_instruction[2] ) );
  DFF \u_a23_core/u_decode/pre_fetch_instruction_reg[1]  ( .D(
        \u_a23_core/u_decode/n1464 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/pre_fetch_instruction[1] ) );
  DFF \u_a23_core/u_decode/o_reg_write_sel_reg[1]  ( .D(n16637), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\u_a23_core/reg_write_sel[1] ) );
  DFF \u_a23_core/u_decode/control_state_reg[3]  ( .D(
        \u_a23_core/u_decode/control_state_nxt[3] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\u_a23_core/u_decode/control_state[3] ) );
  DFF \u_a23_core/u_decode/control_state_reg[4]  ( .D(
        \u_a23_core/u_decode/control_state_nxt[4] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\u_a23_core/u_decode/control_state[4] ) );
  DFF \u_a23_core/u_decode/o_imm_shift_amount_reg[0]  ( .D(
        \u_a23_core/u_decode/instruction[7] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/imm_shift_amount[0] ) );
  DFF \u_a23_core/u_decode/saved_current_instruction_reg[7]  ( .D(
        \u_a23_core/u_decode/n1473 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/saved_current_instruction[7] ) );
  DFF \u_a23_core/u_decode/saved_current_instruction_reg[0]  ( .D(
        \u_a23_core/u_decode/n1480 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/saved_current_instruction[0] ) );
  DFF \u_a23_core/u_decode/control_state_reg[1]  ( .D(
        \u_a23_core/u_decode/control_state_nxt[1] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\u_a23_core/u_decode/control_state[1] ) );
  DFF \u_a23_core/u_decode/control_state_reg[2]  ( .D(
        \u_a23_core/u_decode/control_state_nxt[2] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\u_a23_core/u_decode/control_state[2] ) );
  DFF \u_a23_core/u_decode/pc_wen_r_reg  ( .D(\u_a23_core/u_decode/pc_wen_nxt ), .CLK(clk), .RST(rst), .I(1'b1), .Q(\u_a23_core/pc_wen ) );
  DFF \u_a23_core/u_decode/control_state_reg[0]  ( .D(
        \u_a23_core/u_decode/control_state_nxt[0] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\u_a23_core/u_decode/control_state[0] ) );
  DFF \u_a23_core/u_decode/o_rm_sel_reg[1]  ( .D(\u_a23_core/rm_sel_nxt[1] ), 
        .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/rm_sel[1] ) );
  DFF \u_a23_core/u_decode/saved_current_instruction_reg[1]  ( .D(
        \u_a23_core/u_decode/n1479 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/saved_current_instruction[1] ) );
  DFF \u_a23_core/u_decode/o_rm_sel_reg[0]  ( .D(\u_a23_core/rm_sel_nxt[0] ), 
        .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/rm_sel[0] ) );
  DFF \u_a23_core/u_decode/pre_fetch_instruction_reg[0]  ( .D(
        \u_a23_core/u_decode/n1495 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_decode/pre_fetch_instruction[0] ) );
  DFF \u_a23_core/u_decode/o_read_data_alignment_reg[3]  ( .D(
        \u_a23_core/u_execute/address_plus4[0] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\u_a23_core/read_data_alignment[3] ) );
  DFF \u_a23_core/u_decode/o_read_data_alignment_reg[4]  ( .D(
        \u_a23_core/execute_address[1] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/read_data_alignment[4] ) );
  DFF \u_a23_core/u_decode/o_read_data_reg[0]  ( .D(\u_a23_core/read_data[0] ), 
        .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/read_data_s2[0] ) );
  DFF \u_a23_core/u_decode/o_read_data_reg[1]  ( .D(\u_a23_core/read_data[1] ), 
        .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/read_data_s2[1] ) );
  DFF \u_a23_core/u_decode/o_read_data_reg[2]  ( .D(\u_a23_core/read_data[2] ), 
        .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/read_data_s2[2] ) );
  DFF \u_a23_core/u_decode/o_read_data_reg[3]  ( .D(\u_a23_core/read_data[3] ), 
        .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/read_data_s2[3] ) );
  DFF \u_a23_core/u_decode/o_read_data_reg[4]  ( .D(\u_a23_core/read_data[4] ), 
        .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/read_data_s2[4] ) );
  DFF \u_a23_core/u_decode/o_read_data_reg[5]  ( .D(\u_a23_core/read_data[5] ), 
        .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/read_data_s2[5] ) );
  DFF \u_a23_core/u_decode/o_read_data_reg[6]  ( .D(\u_a23_core/read_data[6] ), 
        .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/read_data_s2[6] ) );
  DFF \u_a23_core/u_decode/o_read_data_reg[7]  ( .D(\u_a23_core/read_data[7] ), 
        .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/read_data_s2[7] ) );
  DFF \u_a23_core/u_decode/o_read_data_reg[8]  ( .D(\u_a23_core/read_data[8] ), 
        .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/read_data_s2[8] ) );
  DFF \u_a23_core/u_decode/o_read_data_reg[9]  ( .D(\u_a23_core/read_data[9] ), 
        .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/read_data_s2[9] ) );
  DFF \u_a23_core/u_decode/o_read_data_reg[10]  ( .D(
        \u_a23_core/read_data[10] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/read_data_s2[10] ) );
  DFF \u_a23_core/u_decode/o_read_data_reg[11]  ( .D(
        \u_a23_core/read_data[11] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/read_data_s2[11] ) );
  DFF \u_a23_core/u_decode/o_read_data_reg[12]  ( .D(
        \u_a23_core/read_data[12] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/read_data_s2[12] ) );
  DFF \u_a23_core/u_decode/o_read_data_reg[13]  ( .D(
        \u_a23_core/read_data[13] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/read_data_s2[13] ) );
  DFF \u_a23_core/u_decode/o_read_data_reg[14]  ( .D(
        \u_a23_core/read_data[14] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/read_data_s2[14] ) );
  DFF \u_a23_core/u_decode/o_read_data_reg[15]  ( .D(
        \u_a23_core/read_data[15] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/read_data_s2[15] ) );
  DFF \u_a23_core/u_decode/o_read_data_reg[16]  ( .D(
        \u_a23_core/read_data[16] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/read_data_s2[16] ) );
  DFF \u_a23_core/u_decode/o_read_data_reg[17]  ( .D(
        \u_a23_core/read_data[17] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/read_data_s2[17] ) );
  DFF \u_a23_core/u_decode/o_read_data_reg[18]  ( .D(
        \u_a23_core/read_data[18] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/read_data_s2[18] ) );
  DFF \u_a23_core/u_decode/o_read_data_reg[19]  ( .D(
        \u_a23_core/read_data[19] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/read_data_s2[19] ) );
  DFF \u_a23_core/u_decode/o_read_data_reg[20]  ( .D(
        \u_a23_core/read_data[20] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/read_data_s2[20] ) );
  DFF \u_a23_core/u_decode/o_read_data_reg[21]  ( .D(
        \u_a23_core/read_data[21] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/read_data_s2[21] ) );
  DFF \u_a23_core/u_decode/o_read_data_reg[22]  ( .D(
        \u_a23_core/read_data[22] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/read_data_s2[22] ) );
  DFF \u_a23_core/u_decode/o_read_data_reg[23]  ( .D(
        \u_a23_core/read_data[23] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/read_data_s2[23] ) );
  DFF \u_a23_core/u_decode/o_read_data_reg[24]  ( .D(
        \u_a23_core/read_data[24] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/read_data_s2[24] ) );
  DFF \u_a23_core/u_decode/o_read_data_reg[25]  ( .D(
        \u_a23_core/read_data[25] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/read_data_s2[25] ) );
  DFF \u_a23_core/u_decode/o_read_data_reg[26]  ( .D(
        \u_a23_core/read_data[26] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/read_data_s2[26] ) );
  DFF \u_a23_core/u_decode/o_read_data_reg[27]  ( .D(
        \u_a23_core/read_data[27] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/read_data_s2[27] ) );
  DFF \u_a23_core/u_decode/o_read_data_reg[28]  ( .D(
        \u_a23_core/read_data[28] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/read_data_s2[28] ) );
  DFF \u_a23_core/u_decode/o_read_data_reg[29]  ( .D(
        \u_a23_core/read_data[29] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/read_data_s2[29] ) );
  DFF \u_a23_core/u_decode/o_read_data_reg[30]  ( .D(
        \u_a23_core/read_data[30] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/read_data_s2[30] ) );
  DFF \u_a23_core/u_decode/o_read_data_reg[31]  ( .D(
        \u_a23_core/read_data[31] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/read_data_s2[31] ) );
  DFF \u_a23_core/u_execute/o_write_data_reg[0]  ( .D(
        \u_a23_core/u_execute/rs[0] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        m_write[0]) );
  DFF \u_a23_core/u_execute/o_write_data_reg[1]  ( .D(
        \u_a23_core/u_execute/rs[1] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        m_write[1]) );
  DFF \u_a23_core/u_execute/o_write_data_reg[2]  ( .D(
        \u_a23_core/u_execute/write_data_nxt[2] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_write[2]) );
  DFF \u_a23_core/u_execute/o_write_data_reg[3]  ( .D(
        \u_a23_core/u_execute/write_data_nxt[3] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_write[3]) );
  DFF \u_a23_core/u_execute/o_write_data_reg[4]  ( .D(
        \u_a23_core/u_execute/write_data_nxt[4] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_write[4]) );
  DFF \u_a23_core/u_execute/o_write_data_reg[5]  ( .D(
        \u_a23_core/u_execute/write_data_nxt[5] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_write[5]) );
  DFF \u_a23_core/u_execute/o_write_data_reg[6]  ( .D(
        \u_a23_core/u_execute/write_data_nxt[6] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_write[6]) );
  DFF \u_a23_core/u_execute/o_write_data_reg[7]  ( .D(
        \u_a23_core/u_execute/write_data_nxt[7] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_write[7]) );
  DFF \u_a23_core/u_execute/o_write_data_reg[8]  ( .D(
        \u_a23_core/u_execute/write_data_nxt[8] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_write[8]) );
  DFF \u_a23_core/u_execute/o_write_data_reg[9]  ( .D(
        \u_a23_core/u_execute/write_data_nxt[9] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_write[9]) );
  DFF \u_a23_core/u_execute/o_write_data_reg[10]  ( .D(
        \u_a23_core/u_execute/write_data_nxt[10] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_write[10]) );
  DFF \u_a23_core/u_execute/o_write_data_reg[11]  ( .D(
        \u_a23_core/u_execute/write_data_nxt[11] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_write[11]) );
  DFF \u_a23_core/u_execute/o_write_data_reg[12]  ( .D(
        \u_a23_core/u_execute/write_data_nxt[12] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_write[12]) );
  DFF \u_a23_core/u_execute/o_write_data_reg[13]  ( .D(
        \u_a23_core/u_execute/write_data_nxt[13] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_write[13]) );
  DFF \u_a23_core/u_execute/o_write_data_reg[14]  ( .D(
        \u_a23_core/u_execute/write_data_nxt[14] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_write[14]) );
  DFF \u_a23_core/u_execute/o_write_data_reg[15]  ( .D(
        \u_a23_core/u_execute/write_data_nxt[15] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_write[15]) );
  DFF \u_a23_core/u_execute/o_write_data_reg[16]  ( .D(
        \u_a23_core/u_execute/write_data_nxt[16] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_write[16]) );
  DFF \u_a23_core/u_execute/o_write_data_reg[17]  ( .D(
        \u_a23_core/u_execute/write_data_nxt[17] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_write[17]) );
  DFF \u_a23_core/u_execute/o_write_data_reg[18]  ( .D(
        \u_a23_core/u_execute/write_data_nxt[18] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_write[18]) );
  DFF \u_a23_core/u_execute/o_write_data_reg[19]  ( .D(
        \u_a23_core/u_execute/write_data_nxt[19] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_write[19]) );
  DFF \u_a23_core/u_execute/o_write_data_reg[20]  ( .D(
        \u_a23_core/u_execute/write_data_nxt[20] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_write[20]) );
  DFF \u_a23_core/u_execute/o_write_data_reg[21]  ( .D(
        \u_a23_core/u_execute/write_data_nxt[21] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_write[21]) );
  DFF \u_a23_core/u_execute/o_write_data_reg[22]  ( .D(
        \u_a23_core/u_execute/write_data_nxt[22] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_write[22]) );
  DFF \u_a23_core/u_execute/o_write_data_reg[23]  ( .D(
        \u_a23_core/u_execute/write_data_nxt[23] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_write[23]) );
  DFF \u_a23_core/u_execute/o_write_data_reg[24]  ( .D(
        \u_a23_core/u_execute/write_data_nxt[24] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_write[24]) );
  DFF \u_a23_core/u_execute/o_write_data_reg[25]  ( .D(
        \u_a23_core/u_execute/write_data_nxt[25] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_write[25]) );
  DFF \u_a23_core/u_execute/o_write_data_reg[26]  ( .D(
        \u_a23_core/u_execute/write_data_nxt[26] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_write[26]) );
  DFF \u_a23_core/u_execute/o_write_data_reg[27]  ( .D(
        \u_a23_core/u_execute/write_data_nxt[27] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_write[27]) );
  DFF \u_a23_core/u_execute/o_write_data_reg[28]  ( .D(
        \u_a23_core/u_execute/write_data_nxt[28] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_write[28]) );
  DFF \u_a23_core/u_execute/o_write_data_reg[29]  ( .D(
        \u_a23_core/u_execute/write_data_nxt[29] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_write[29]) );
  DFF \u_a23_core/u_execute/o_write_data_reg[30]  ( .D(
        \u_a23_core/u_execute/write_data_nxt[30] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_write[30]) );
  DFF \u_a23_core/u_execute/o_write_data_reg[31]  ( .D(
        \u_a23_core/u_execute/write_data_nxt[31] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_write[31]) );
  DFF \u_a23_core/u_execute/o_write_enable_reg  ( .D(
        \u_a23_core/u_execute/write_enable_nxt ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_write_en) );
  DFF \u_a23_core/u_execute/address_r_reg[30]  ( .D(
        \u_a23_core/execute_address_nxt[30] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(m_address[30]) );
  DFF \u_a23_core/u_execute/address_r_reg[29]  ( .D(
        \u_a23_core/execute_address_nxt[29] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(m_address[29]) );
  DFF \u_a23_core/u_execute/address_r_reg[28]  ( .D(
        \u_a23_core/execute_address_nxt[28] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(m_address[28]) );
  DFF \u_a23_core/u_execute/address_r_reg[27]  ( .D(
        \u_a23_core/execute_address_nxt[27] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(m_address[27]) );
  DFF \u_a23_core/u_execute/address_r_reg[26]  ( .D(
        \u_a23_core/execute_address_nxt[26] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(m_address[26]) );
  DFF \u_a23_core/u_execute/address_r_reg[25]  ( .D(
        \u_a23_core/execute_address_nxt[25] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(m_address[25]) );
  DFF \u_a23_core/u_execute/address_r_reg[24]  ( .D(
        \u_a23_core/execute_address_nxt[24] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(m_address[24]) );
  DFF \u_a23_core/u_execute/address_r_reg[23]  ( .D(
        \u_a23_core/execute_address_nxt[23] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(m_address[23]) );
  DFF \u_a23_core/u_execute/address_r_reg[22]  ( .D(
        \u_a23_core/execute_address_nxt[22] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(m_address[22]) );
  DFF \u_a23_core/u_execute/address_r_reg[21]  ( .D(
        \u_a23_core/execute_address_nxt[21] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(m_address[21]) );
  DFF \u_a23_core/u_execute/address_r_reg[20]  ( .D(
        \u_a23_core/execute_address_nxt[20] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(m_address[20]) );
  DFF \u_a23_core/u_execute/address_r_reg[19]  ( .D(
        \u_a23_core/execute_address_nxt[19] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(m_address[19]) );
  DFF \u_a23_core/u_execute/address_r_reg[18]  ( .D(
        \u_a23_core/execute_address_nxt[18] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(m_address[18]) );
  DFF \u_a23_core/u_execute/address_r_reg[17]  ( .D(
        \u_a23_core/execute_address_nxt[17] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(m_address[17]) );
  DFF \u_a23_core/u_execute/address_r_reg[16]  ( .D(
        \u_a23_core/execute_address_nxt[16] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(m_address[16]) );
  DFF \u_a23_core/u_execute/address_r_reg[15]  ( .D(
        \u_a23_core/execute_address_nxt[15] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(m_address[15]) );
  DFF \u_a23_core/u_execute/address_r_reg[14]  ( .D(
        \u_a23_core/execute_address_nxt[14] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(m_address[14]) );
  DFF \u_a23_core/u_execute/address_r_reg[13]  ( .D(
        \u_a23_core/execute_address_nxt[13] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(m_address[13]) );
  DFF \u_a23_core/u_execute/address_r_reg[12]  ( .D(
        \u_a23_core/execute_address_nxt[12] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(m_address[12]) );
  DFF \u_a23_core/u_execute/address_r_reg[11]  ( .D(
        \u_a23_core/execute_address_nxt[11] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(m_address[11]) );
  DFF \u_a23_core/u_execute/address_r_reg[10]  ( .D(
        \u_a23_core/execute_address_nxt[10] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(m_address[10]) );
  DFF \u_a23_core/u_execute/address_r_reg[9]  ( .D(
        \u_a23_core/execute_address_nxt[9] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(m_address[9]) );
  DFF \u_a23_core/u_execute/address_r_reg[8]  ( .D(
        \u_a23_core/execute_address_nxt[8] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(m_address[8]) );
  DFF \u_a23_core/u_execute/address_r_reg[7]  ( .D(
        \u_a23_core/execute_address_nxt[7] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(m_address[7]) );
  DFF \u_a23_core/u_execute/address_r_reg[6]  ( .D(
        \u_a23_core/execute_address_nxt[6] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(m_address[6]) );
  DFF \u_a23_core/u_execute/address_r_reg[5]  ( .D(
        \u_a23_core/execute_address_nxt[5] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(m_address[5]) );
  DFF \u_a23_core/u_execute/address_r_reg[4]  ( .D(
        \u_a23_core/execute_address_nxt[4] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(m_address[4]) );
  DFF \u_a23_core/u_execute/address_r_reg[3]  ( .D(
        \u_a23_core/execute_address_nxt[3] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(m_address[3]) );
  DFF \u_a23_core/u_execute/address_r_reg[2]  ( .D(
        \u_a23_core/execute_address_nxt[2] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(m_address[2]) );
  DFF \u_a23_core/u_execute/o_byte_enable_reg[2]  ( .D(
        \u_a23_core/u_execute/byte_enable_nxt[2] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_byte_enable[2]) );
  DFF \u_a23_core/u_execute/o_byte_enable_reg[3]  ( .D(
        \u_a23_core/u_execute/byte_enable_nxt[3] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_byte_enable[3]) );
  DFF \u_a23_core/u_execute/o_byte_enable_reg[1]  ( .D(
        \u_a23_core/u_execute/byte_enable_nxt[1] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_byte_enable[1]) );
  DFF \u_a23_core/u_execute/o_byte_enable_reg[0]  ( .D(
        \u_a23_core/u_execute/byte_enable_nxt[0] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(m_byte_enable[0]) );
  DFF \u_a23_core/u_execute/address_r_reg[1]  ( .D(
        \u_a23_core/execute_address_nxt[1] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/execute_address[1] ) );
  DFF \u_a23_core/u_execute/address_r_reg[0]  ( .D(
        \u_a23_core/execute_address_nxt[0] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\u_a23_core/u_execute/address_plus4[0] ) );
  DFF \u_a23_core/u_execute/address_r_reg[31]  ( .D(
        \u_a23_core/execute_address_nxt[31] ), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(m_address[31]) );
  DFF \u_a23_core/u_execute/status_bits_flags_reg[2]  ( .D(
        \u_a23_core/u_execute/n1074 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_execute/save_int_pc_m4[30] ) );
  DFF \u_a23_core/u_execute/status_bits_flags_reg[1]  ( .D(
        \u_a23_core/u_execute/n1075 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_execute/save_int_pc_m4[29] ) );
  DFF \u_a23_core/u_execute/status_bits_flags_reg[3]  ( .D(
        \u_a23_core/u_execute/n1073 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_execute/save_int_pc_m4[31] ) );
  DFF \u_a23_core/u_execute/status_bits_flags_reg[0]  ( .D(
        \u_a23_core/u_execute/n1076 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \u_a23_core/u_execute/save_int_pc_m4[28] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[66]  ( .D(
        \u_a23_core/u_execute/u_multiply/n544 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[66] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[67]  ( .D(
        \u_a23_core/u_execute/u_multiply/n543 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[67] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[65]  ( .D(
        \u_a23_core/u_execute/u_multiply/n545 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[65] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[64]  ( .D(
        \u_a23_core/u_execute/u_multiply/n546 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[64] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[63]  ( .D(
        \u_a23_core/u_execute/u_multiply/n547 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[63] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[62]  ( .D(
        \u_a23_core/u_execute/u_multiply/n548 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[62] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[61]  ( .D(
        \u_a23_core/u_execute/u_multiply/n549 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[61] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[60]  ( .D(
        \u_a23_core/u_execute/u_multiply/n550 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[60] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[59]  ( .D(
        \u_a23_core/u_execute/u_multiply/n551 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[59] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[58]  ( .D(
        \u_a23_core/u_execute/u_multiply/n552 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[58] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[57]  ( .D(
        \u_a23_core/u_execute/u_multiply/n553 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[57] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[56]  ( .D(
        \u_a23_core/u_execute/u_multiply/n554 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[56] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[55]  ( .D(
        \u_a23_core/u_execute/u_multiply/n555 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[55] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[54]  ( .D(
        \u_a23_core/u_execute/u_multiply/n556 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[54] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[53]  ( .D(
        \u_a23_core/u_execute/u_multiply/n557 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[53] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[52]  ( .D(
        \u_a23_core/u_execute/u_multiply/n558 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[52] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[51]  ( .D(
        \u_a23_core/u_execute/u_multiply/n559 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[51] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[50]  ( .D(
        \u_a23_core/u_execute/u_multiply/n560 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[50] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[49]  ( .D(
        \u_a23_core/u_execute/u_multiply/n561 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[49] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[48]  ( .D(
        \u_a23_core/u_execute/u_multiply/n562 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[48] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[47]  ( .D(
        \u_a23_core/u_execute/u_multiply/n563 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[47] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[46]  ( .D(
        \u_a23_core/u_execute/u_multiply/n564 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[46] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[45]  ( .D(
        \u_a23_core/u_execute/u_multiply/n565 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[45] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[44]  ( .D(
        \u_a23_core/u_execute/u_multiply/n566 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[44] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[43]  ( .D(
        \u_a23_core/u_execute/u_multiply/n567 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[43] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[42]  ( .D(
        \u_a23_core/u_execute/u_multiply/n568 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[42] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[41]  ( .D(
        \u_a23_core/u_execute/u_multiply/n569 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[41] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[40]  ( .D(
        \u_a23_core/u_execute/u_multiply/n570 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[40] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[39]  ( .D(
        \u_a23_core/u_execute/u_multiply/n571 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[39] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[38]  ( .D(
        \u_a23_core/u_execute/u_multiply/n572 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[38] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[37]  ( .D(
        \u_a23_core/u_execute/u_multiply/n573 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[37] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[36]  ( .D(
        \u_a23_core/u_execute/u_multiply/n574 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[36] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[35]  ( .D(
        \u_a23_core/u_execute/u_multiply/n575 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[35] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[34]  ( .D(
        \u_a23_core/u_execute/u_multiply/n576 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[34] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[1]  ( .D(
        \u_a23_core/u_execute/u_multiply/n608 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/multiply_out[0] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[2]  ( .D(
        \u_a23_core/u_execute/u_multiply/n607 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/multiply_out[1] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[3]  ( .D(
        \u_a23_core/u_execute/u_multiply/n606 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/multiply_out[2] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[4]  ( .D(
        \u_a23_core/u_execute/u_multiply/n605 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/multiply_out[3] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[5]  ( .D(
        \u_a23_core/u_execute/u_multiply/n604 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/multiply_out[4] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[6]  ( .D(
        \u_a23_core/u_execute/u_multiply/n603 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/multiply_out[5] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[7]  ( .D(
        \u_a23_core/u_execute/u_multiply/n602 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/multiply_out[6] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[8]  ( .D(
        \u_a23_core/u_execute/u_multiply/n601 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/multiply_out[7] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[9]  ( .D(
        \u_a23_core/u_execute/u_multiply/n600 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/multiply_out[8] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[10]  ( .D(
        \u_a23_core/u_execute/u_multiply/n599 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/multiply_out[9] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[11]  ( .D(
        \u_a23_core/u_execute/u_multiply/n598 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/multiply_out[10] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[12]  ( .D(
        \u_a23_core/u_execute/u_multiply/n597 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/multiply_out[11] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[13]  ( .D(
        \u_a23_core/u_execute/u_multiply/n596 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/multiply_out[12] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[14]  ( .D(
        \u_a23_core/u_execute/u_multiply/n595 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/multiply_out[13] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[15]  ( .D(
        \u_a23_core/u_execute/u_multiply/n594 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/multiply_out[14] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[16]  ( .D(
        \u_a23_core/u_execute/u_multiply/n593 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/multiply_out[15] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[17]  ( .D(
        \u_a23_core/u_execute/u_multiply/n592 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/multiply_out[16] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[18]  ( .D(
        \u_a23_core/u_execute/u_multiply/n591 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/multiply_out[17] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[19]  ( .D(
        \u_a23_core/u_execute/u_multiply/n590 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/multiply_out[18] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[20]  ( .D(
        \u_a23_core/u_execute/u_multiply/n589 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/multiply_out[19] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[21]  ( .D(
        \u_a23_core/u_execute/u_multiply/n588 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/multiply_out[20] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[22]  ( .D(
        \u_a23_core/u_execute/u_multiply/n587 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/multiply_out[21] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[23]  ( .D(
        \u_a23_core/u_execute/u_multiply/n586 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/multiply_out[22] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[24]  ( .D(
        \u_a23_core/u_execute/u_multiply/n585 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/multiply_out[23] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[25]  ( .D(
        \u_a23_core/u_execute/u_multiply/n584 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/multiply_out[24] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[26]  ( .D(
        \u_a23_core/u_execute/u_multiply/n583 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/multiply_out[25] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[27]  ( .D(
        \u_a23_core/u_execute/u_multiply/n582 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/multiply_out[26] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[28]  ( .D(
        \u_a23_core/u_execute/u_multiply/n581 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/multiply_out[27] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[29]  ( .D(
        \u_a23_core/u_execute/u_multiply/n580 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/multiply_out[28] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[30]  ( .D(
        \u_a23_core/u_execute/u_multiply/n579 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/multiply_out[29] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[31]  ( .D(
        \u_a23_core/u_execute/u_multiply/n578 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/multiply_out[30] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[32]  ( .D(
        \u_a23_core/u_execute/u_multiply/n577 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/multiply_out[31] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[33]  ( .D(
        \u_a23_core/u_execute/u_multiply/n609 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product[33] ) );
  DFF \u_a23_core/u_execute/u_multiply/product_reg[0]  ( .D(
        \u_a23_core/u_execute/u_multiply/n610 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/product_0 ) );
  DFF \u_a23_core/u_execute/u_multiply/o_done_reg  ( .D(
        \u_a23_core/u_execute/u_multiply/n499 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/multiply_done ) );
  DFF \u_a23_core/u_execute/u_multiply/count_reg[5]  ( .D(
        \u_a23_core/u_execute/u_multiply/n501 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/count[5] ) );
  DFF \u_a23_core/u_execute/u_multiply/count_reg[4]  ( .D(
        \u_a23_core/u_execute/u_multiply/n503 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/count[4] ) );
  DFF \u_a23_core/u_execute/u_multiply/count_reg[3]  ( .D(
        \u_a23_core/u_execute/u_multiply/n505 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/count[3] ) );
  DFF \u_a23_core/u_execute/u_multiply/count_reg[2]  ( .D(
        \u_a23_core/u_execute/u_multiply/n507 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/count[2] ) );
  DFF \u_a23_core/u_execute/u_multiply/count_reg[1]  ( .D(
        \u_a23_core/u_execute/u_multiply/n509 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/count[1] ) );
  DFF \u_a23_core/u_execute/u_multiply/count_reg[0]  ( .D(
        \u_a23_core/u_execute/u_multiply/n611 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(\u_a23_core/u_execute/u_multiply/count[0] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r10_reg[0]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n3975 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r10[0] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r10_reg[1]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n3977 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r10[1] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r10_reg[2]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n3979 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r10[2] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r10_reg[3]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n3981 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r10[3] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r10_reg[4]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n3983 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r10[4] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r10_reg[5]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n3985 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r10[5] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r10_reg[6]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n3987 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r10[6] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r10_reg[7]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n3989 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r10[7] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r10_reg[8]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n3991 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r10[8] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r10_reg[9]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n3993 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r10[9] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r10_reg[10]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n3995 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r10[10] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r10_reg[11]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n3997 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r10[11] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r10_reg[12]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n3999 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r10[12] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r10_reg[13]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4001 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r10[13] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r10_reg[14]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4003 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r10[14] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r10_reg[15]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4005 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r10[15] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r10_reg[16]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4007 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r10[16] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r10_reg[17]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4009 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r10[17] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r10_reg[18]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4011 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r10[18] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r10_reg[19]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4013 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r10[19] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r10_reg[20]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4015 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r10[20] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r10_reg[21]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4017 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r10[21] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r10_reg[22]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4019 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r10[22] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r10_reg[23]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4021 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r10[23] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r10_reg[24]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4023 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r10[24] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r10_reg[25]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4025 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r10[25] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r10_reg[26]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4027 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r10[26] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r10_reg[27]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4029 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r10[27] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r10_reg[28]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4031 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r10[28] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r10_reg[29]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4033 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r10[29] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r10_reg[30]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4035 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r10[30] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r10_reg[31]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4037 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r10[31] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r9_reg[0]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4039 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r9[0] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r9_reg[1]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4041 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r9[1] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r9_reg[2]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4043 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r9[2] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r9_reg[3]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4045 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r9[3] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r9_reg[4]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4047 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r9[4] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r9_reg[5]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4049 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r9[5] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r9_reg[6]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4051 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r9[6] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r9_reg[7]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4053 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r9[7] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r9_reg[8]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4055 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r9[8] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r9_reg[9]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4057 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r9[9] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r9_reg[10]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4059 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r9[10] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r9_reg[11]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4061 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r9[11] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r9_reg[12]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4063 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r9[12] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r9_reg[13]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4065 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r9[13] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r9_reg[14]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4067 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r9[14] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r9_reg[15]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4069 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r9[15] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r9_reg[16]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4071 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r9[16] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r9_reg[17]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4073 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r9[17] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r9_reg[18]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4075 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r9[18] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r9_reg[19]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4077 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r9[19] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r9_reg[20]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4079 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r9[20] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r9_reg[21]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4081 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r9[21] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r9_reg[22]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4083 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r9[22] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r9_reg[23]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4085 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r9[23] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r9_reg[24]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4087 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r9[24] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r9_reg[25]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4089 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r9[25] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r9_reg[26]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4091 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r9[26] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r9_reg[27]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4093 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r9[27] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r9_reg[28]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4095 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r9[28] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r9_reg[29]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4097 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r9[29] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r9_reg[30]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4099 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r9[30] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r9_reg[31]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4101 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r9[31] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r8_reg[0]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4103 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r8[0] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r8_reg[1]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4105 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r8[1] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r8_reg[2]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4107 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r8[2] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r8_reg[3]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4109 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r8[3] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r8_reg[4]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4111 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r8[4] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r8_reg[5]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4113 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r8[5] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r8_reg[6]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4115 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r8[6] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r8_reg[7]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4117 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r8[7] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r8_reg[8]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4119 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r8[8] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r8_reg[9]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4121 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r8[9] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r8_reg[10]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4123 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r8[10] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r8_reg[11]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4125 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r8[11] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r8_reg[12]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4127 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r8[12] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r8_reg[13]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4129 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r8[13] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r8_reg[14]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4131 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r8[14] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r8_reg[15]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4133 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r8[15] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r8_reg[16]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4135 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r8[16] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r8_reg[17]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4137 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r8[17] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r8_reg[18]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4139 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r8[18] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r8_reg[19]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4141 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r8[19] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r8_reg[20]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4143 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r8[20] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r8_reg[21]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4145 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r8[21] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r8_reg[22]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4147 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r8[22] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r8_reg[23]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4149 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r8[23] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r8_reg[24]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4151 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r8[24] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r8_reg[25]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4153 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r8[25] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r8_reg[26]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4155 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r8[26] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r8_reg[27]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4157 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r8[27] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r8_reg[28]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4159 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r8[28] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r8_reg[29]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4161 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r8[29] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r8_reg[30]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4163 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r8[30] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r8_reg[31]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4165 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r8[31] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r7_reg[0]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4167 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r7[0] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r7_reg[1]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4169 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r7[1] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r7_reg[2]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4171 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r7[2] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r7_reg[3]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4173 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r7[3] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r7_reg[4]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4175 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r7[4] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r7_reg[5]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4177 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r7[5] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r7_reg[6]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4179 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r7[6] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r7_reg[7]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4181 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r7[7] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r7_reg[8]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4183 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r7[8] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r7_reg[9]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4185 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r7[9] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r7_reg[10]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4187 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r7[10] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r7_reg[11]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4189 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r7[11] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r7_reg[12]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4191 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r7[12] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r7_reg[13]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4193 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r7[13] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r7_reg[14]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4195 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r7[14] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r7_reg[15]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4197 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r7[15] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r7_reg[16]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4199 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r7[16] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r7_reg[17]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4201 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r7[17] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r7_reg[18]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4203 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r7[18] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r7_reg[19]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4205 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r7[19] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r7_reg[20]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4207 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r7[20] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r7_reg[21]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4209 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r7[21] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r7_reg[22]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4211 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r7[22] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r7_reg[23]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4213 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r7[23] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r7_reg[24]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4215 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r7[24] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r7_reg[25]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4217 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r7[25] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r7_reg[26]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4219 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r7[26] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r7_reg[27]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4221 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r7[27] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r7_reg[28]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4223 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r7[28] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r7_reg[29]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4225 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r7[29] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r7_reg[30]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4227 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r7[30] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r7_reg[31]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4229 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r7[31] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r6_reg[0]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4231 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r6[0] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r6_reg[1]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4233 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r6[1] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r6_reg[2]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4235 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r6[2] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r6_reg[3]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4237 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r6[3] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r6_reg[4]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4239 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r6[4] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r6_reg[5]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4241 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r6[5] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r6_reg[6]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4243 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r6[6] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r6_reg[7]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4245 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r6[7] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r6_reg[8]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4247 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r6[8] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r6_reg[9]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4249 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r6[9] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r6_reg[10]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4251 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r6[10] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r6_reg[11]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4253 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r6[11] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r6_reg[12]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4255 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r6[12] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r6_reg[13]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4257 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r6[13] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r6_reg[14]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4259 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r6[14] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r6_reg[15]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4261 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r6[15] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r6_reg[16]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4263 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r6[16] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r6_reg[17]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4265 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r6[17] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r6_reg[18]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4267 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r6[18] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r6_reg[19]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4269 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r6[19] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r6_reg[20]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4271 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r6[20] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r6_reg[21]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4273 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r6[21] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r6_reg[22]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4275 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r6[22] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r6_reg[23]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4277 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r6[23] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r6_reg[24]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4279 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r6[24] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r6_reg[25]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4281 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r6[25] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r6_reg[26]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4283 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r6[26] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r6_reg[27]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4285 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r6[27] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r6_reg[28]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4287 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r6[28] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r6_reg[29]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4289 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r6[29] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r6_reg[30]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4291 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r6[30] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r6_reg[31]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4293 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r6[31] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r5_reg[0]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4295 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r5[0] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r5_reg[1]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4297 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r5[1] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r5_reg[2]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4299 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r5[2] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r5_reg[3]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4301 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r5[3] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r5_reg[4]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4303 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r5[4] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r5_reg[5]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4305 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r5[5] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r5_reg[6]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4307 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r5[6] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r5_reg[7]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4309 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r5[7] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r5_reg[8]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4311 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r5[8] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r5_reg[9]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4313 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r5[9] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r5_reg[10]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4315 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r5[10] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r5_reg[11]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4317 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r5[11] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r5_reg[12]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4319 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r5[12] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r5_reg[13]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4321 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r5[13] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r5_reg[14]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4323 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r5[14] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r5_reg[15]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4325 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r5[15] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r5_reg[16]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4327 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r5[16] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r5_reg[17]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4329 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r5[17] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r5_reg[18]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4331 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r5[18] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r5_reg[19]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4333 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r5[19] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r5_reg[20]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4335 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r5[20] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r5_reg[21]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4337 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r5[21] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r5_reg[22]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4339 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r5[22] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r5_reg[23]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4341 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r5[23] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r5_reg[24]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4343 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r5[24] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r5_reg[25]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4345 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r5[25] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r5_reg[26]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4347 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r5[26] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r5_reg[27]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4349 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r5[27] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r5_reg[28]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4351 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r5[28] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r5_reg[29]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4353 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r5[29] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r5_reg[30]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4355 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r5[30] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r5_reg[31]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4357 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r5[31] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r4_reg[0]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4359 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r4[0] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r4_reg[1]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4361 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r4[1] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r4_reg[2]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4363 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r4[2] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r4_reg[3]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4365 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r4[3] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r4_reg[4]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4367 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r4[4] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r4_reg[5]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4369 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r4[5] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r4_reg[6]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4371 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r4[6] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r4_reg[7]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4373 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r4[7] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r4_reg[8]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4375 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r4[8] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r4_reg[9]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4377 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r4[9] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r4_reg[10]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4379 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r4[10] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r4_reg[11]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4381 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r4[11] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r4_reg[12]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4383 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r4[12] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r4_reg[13]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4385 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r4[13] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r4_reg[14]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4387 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r4[14] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r4_reg[15]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4389 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r4[15] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r4_reg[16]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4391 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r4[16] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r4_reg[17]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4393 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r4[17] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r4_reg[18]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4395 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r4[18] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r4_reg[19]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4397 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r4[19] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r4_reg[20]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4399 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r4[20] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r4_reg[21]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4401 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r4[21] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r4_reg[22]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4403 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r4[22] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r4_reg[23]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4405 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r4[23] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r4_reg[24]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4407 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r4[24] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r4_reg[25]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4409 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r4[25] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r4_reg[26]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4411 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r4[26] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r4_reg[27]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4413 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r4[27] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r4_reg[28]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4415 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r4[28] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r4_reg[29]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4417 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r4[29] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r4_reg[30]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4419 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r4[30] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r4_reg[31]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4421 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r4[31] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r3_reg[0]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4423 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r3[0] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r3_reg[1]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4425 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r3[1] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r3_reg[2]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4427 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r3[2] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r3_reg[3]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4429 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r3[3] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r3_reg[4]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4431 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r3[4] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r3_reg[5]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4433 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r3[5] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r3_reg[6]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4435 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r3[6] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r3_reg[7]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4437 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r3[7] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r3_reg[8]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4439 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r3[8] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r3_reg[9]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4441 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r3[9] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r3_reg[10]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4443 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r3[10] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r3_reg[11]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4445 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r3[11] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r3_reg[12]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4447 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r3[12] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r3_reg[13]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4449 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r3[13] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r3_reg[14]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4451 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r3[14] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r3_reg[15]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4453 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r3[15] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r3_reg[16]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4455 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r3[16] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r3_reg[17]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4457 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r3[17] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r3_reg[18]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4459 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r3[18] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r3_reg[19]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4461 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r3[19] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r3_reg[20]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4463 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r3[20] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r3_reg[21]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4465 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r3[21] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r3_reg[22]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4467 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r3[22] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r3_reg[23]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4469 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r3[23] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r3_reg[24]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4471 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r3[24] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r3_reg[25]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4473 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r3[25] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r3_reg[26]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4475 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r3[26] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r3_reg[27]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4477 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r3[27] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r3_reg[28]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4479 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r3[28] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r3_reg[29]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4481 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r3[29] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r3_reg[30]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4483 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r3[30] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r3_reg[31]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4485 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r3[31] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r2_reg[0]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4487 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r2[0] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r2_reg[1]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4489 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r2[1] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r2_reg[2]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4491 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r2[2] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r2_reg[3]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4493 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r2[3] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r2_reg[4]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4495 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r2[4] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r2_reg[5]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4497 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r2[5] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r2_reg[6]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4499 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r2[6] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r2_reg[7]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4501 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r2[7] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r2_reg[8]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4503 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r2[8] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r2_reg[9]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4505 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r2[9] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r2_reg[10]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4507 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r2[10] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r2_reg[11]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4509 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r2[11] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r2_reg[12]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4511 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r2[12] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r2_reg[13]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4513 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r2[13] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r2_reg[14]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4515 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r2[14] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r2_reg[15]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4517 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r2[15] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r2_reg[16]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4519 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r2[16] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r2_reg[17]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4521 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r2[17] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r2_reg[18]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4523 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r2[18] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r2_reg[19]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4525 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r2[19] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r2_reg[20]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4527 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r2[20] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r2_reg[21]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4529 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r2[21] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r2_reg[22]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4531 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r2[22] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r2_reg[23]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4533 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r2[23] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r2_reg[24]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4535 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r2[24] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r2_reg[25]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4537 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r2[25] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r2_reg[26]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4539 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r2[26] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r2_reg[27]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4541 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r2[27] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r2_reg[28]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4543 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r2[28] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r2_reg[29]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4545 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r2[29] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r2_reg[30]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4547 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r2[30] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r2_reg[31]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4549 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r2[31] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r1_reg[0]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4551 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r1[0] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r1_reg[1]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4553 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r1[1] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r1_reg[2]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4555 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r1[2] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r1_reg[3]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4557 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r1[3] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r1_reg[4]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4559 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r1[4] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r1_reg[5]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4561 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r1[5] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r1_reg[6]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4563 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r1[6] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r1_reg[7]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4565 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r1[7] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r1_reg[8]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4567 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r1[8] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r1_reg[9]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4569 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r1[9] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r1_reg[10]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4571 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r1[10] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r1_reg[11]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4573 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r1[11] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r1_reg[12]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4575 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r1[12] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r1_reg[13]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4577 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r1[13] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r1_reg[14]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4579 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r1[14] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r1_reg[15]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4581 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r1[15] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r1_reg[16]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4583 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r1[16] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r1_reg[17]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4585 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r1[17] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r1_reg[18]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4587 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r1[18] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r1_reg[19]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4589 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r1[19] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r1_reg[20]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4591 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r1[20] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r1_reg[21]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4593 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r1[21] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r1_reg[22]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4595 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r1[22] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r1_reg[23]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4597 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r1[23] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r1_reg[24]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4599 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r1[24] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r1_reg[25]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4601 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r1[25] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r1_reg[26]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4603 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r1[26] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r1_reg[27]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4605 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r1[27] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r1_reg[28]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4607 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r1[28] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r1_reg[29]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4609 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r1[29] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r1_reg[30]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4611 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r1[30] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r1_reg[31]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4613 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r1[31] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r0_reg[0]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4615 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r0[0] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r0_reg[1]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4617 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r0[1] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r0_reg[2]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4619 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r0[2] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r0_reg[3]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4621 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r0[3] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r0_reg[4]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4623 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r0[4] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r0_reg[5]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4625 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r0[5] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r0_reg[6]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4627 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r0[6] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r0_reg[7]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4629 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r0[7] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r0_reg[8]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4631 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r0[8] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r0_reg[9]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4633 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r0[9] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r0_reg[10]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4635 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r0[10] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r0_reg[11]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4637 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r0[11] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r0_reg[12]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4639 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r0[12] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r0_reg[13]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4641 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r0[13] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r0_reg[14]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4643 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r0[14] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r0_reg[15]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4645 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r0[15] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r0_reg[16]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4647 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r0[16] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r0_reg[17]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4649 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r0[17] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r0_reg[18]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4651 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r0[18] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r0_reg[19]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4653 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r0[19] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r0_reg[20]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4655 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r0[20] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r0_reg[21]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4657 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r0[21] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r0_reg[22]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4659 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r0[22] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r0_reg[23]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4661 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r0[23] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r0_reg[24]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4663 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r0[24] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r0_reg[25]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4665 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r0[25] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r0_reg[26]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4667 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r0[26] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r0_reg[27]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4669 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r0[27] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r0_reg[28]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4671 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r0[28] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r0_reg[29]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4673 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r0[29] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r0_reg[30]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4675 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r0[30] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r0_reg[31]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4677 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r0[31] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r15_reg[0]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4679 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/pc[2] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r15_reg[1]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4681 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/pc[3] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r15_reg[2]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4683 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/pc[4] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r15_reg[3]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4685 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/pc[5] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r15_reg[4]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4687 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/pc[6] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r15_reg[5]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4689 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/pc[7] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r15_reg[6]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4691 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/pc[8] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r15_reg[7]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4693 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/pc[9] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r15_reg[8]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4695 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/pc[10] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r15_reg[9]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4697 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/pc[11] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r15_reg[10]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4699 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/pc[12] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r15_reg[11]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4701 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/pc[13] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r15_reg[12]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4703 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/pc[14] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r15_reg[13]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4705 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/pc[15] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r15_reg[14]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4707 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/pc[16] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r15_reg[15]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4709 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/pc[17] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r15_reg[16]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4711 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/pc[18] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r15_reg[17]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4713 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/pc[19] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r15_reg[18]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4715 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/pc[20] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r15_reg[19]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4717 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/pc[21] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r15_reg[20]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4719 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/pc[22] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r15_reg[21]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4721 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/pc[23] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r15_reg[22]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4723 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/pc[24] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r15_reg[23]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4725 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/pc[25] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r12_reg[0]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4727 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r12[0] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r12_reg[1]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4729 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r12[1] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r12_reg[2]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4731 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r12[2] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r12_reg[3]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4733 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r12[3] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r12_reg[4]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4735 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r12[4] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r12_reg[5]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4737 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r12[5] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r12_reg[6]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4739 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r12[6] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r12_reg[7]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4741 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r12[7] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r12_reg[8]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4743 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r12[8] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r12_reg[9]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4745 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r12[9] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r12_reg[10]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4747 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r12[10] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r12_reg[11]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4749 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r12[11] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r12_reg[12]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4751 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r12[12] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r12_reg[13]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4753 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r12[13] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r12_reg[14]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4755 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r12[14] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r12_reg[15]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4757 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r12[15] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r12_reg[16]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4759 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r12[16] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r12_reg[17]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4761 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r12[17] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r12_reg[18]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4763 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r12[18] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r12_reg[19]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4765 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r12[19] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r12_reg[20]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4767 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r12[20] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r12_reg[21]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4769 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r12[21] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r12_reg[22]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4771 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r12[22] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r12_reg[23]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4773 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r12[23] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r12_reg[24]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4775 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r12[24] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r12_reg[25]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4777 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r12[25] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r12_reg[26]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4779 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r12[26] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r12_reg[27]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4781 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r12[27] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r12_reg[28]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4783 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r12[28] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r12_reg[29]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4785 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r12[29] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r12_reg[30]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4787 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r12[30] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r12_reg[31]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4789 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r12[31] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r13_reg[0]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4791 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r13[0] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r13_reg[1]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4793 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r13[1] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r13_reg[2]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4795 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r13[2] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r13_reg[3]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4797 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r13[3] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r13_reg[4]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4799 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r13[4] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r13_reg[5]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4801 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r13[5] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r13_reg[6]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4803 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r13[6] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r13_reg[7]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4805 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r13[7] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r13_reg[8]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4807 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r13[8] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r13_reg[9]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4809 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r13[9] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r13_reg[10]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4811 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r13[10] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r13_reg[11]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4813 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r13[11] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r13_reg[12]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4815 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r13[12] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r13_reg[13]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4817 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r13[13] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r13_reg[14]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4819 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r13[14] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r13_reg[15]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4821 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r13[15] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r13_reg[16]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4823 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r13[16] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r13_reg[17]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4825 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r13[17] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r13_reg[18]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4827 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r13[18] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r13_reg[19]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4829 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r13[19] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r13_reg[20]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4831 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r13[20] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r13_reg[21]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4833 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r13[21] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r13_reg[22]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4835 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r13[22] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r13_reg[23]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4837 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r13[23] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r13_reg[24]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4839 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r13[24] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r13_reg[25]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4841 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r13[25] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r13_reg[26]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4843 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r13[26] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r13_reg[27]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4845 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r13[27] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r13_reg[28]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4847 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r13[28] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r13_reg[29]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4849 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r13[29] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r13_reg[30]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4851 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r13[30] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r13_reg[31]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4853 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r13[31] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r14_reg[0]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4855 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r14[0] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r14_reg[1]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4857 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r14[1] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r14_reg[2]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4859 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r14[2] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r14_reg[3]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4861 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r14[3] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r14_reg[4]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4863 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r14[4] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r14_reg[5]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4865 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r14[5] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r14_reg[6]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4867 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r14[6] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r14_reg[7]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4869 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r14[7] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r14_reg[8]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4871 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r14[8] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r14_reg[9]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4873 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r14[9] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r14_reg[10]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4875 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r14[10] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r14_reg[11]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4877 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r14[11] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r14_reg[12]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4879 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r14[12] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r14_reg[13]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4881 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r14[13] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r14_reg[14]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4883 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r14[14] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r14_reg[15]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4885 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r14[15] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r14_reg[16]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4887 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r14[16] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r14_reg[17]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4889 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r14[17] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r14_reg[18]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4891 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r14[18] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r14_reg[19]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4893 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r14[19] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r14_reg[20]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4895 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r14[20] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r14_reg[21]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4897 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r14[21] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r14_reg[22]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4899 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r14[22] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r14_reg[23]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4901 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r14[23] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r14_reg[24]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4903 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r14[24] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r14_reg[25]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4905 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r14[25] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r14_reg[26]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4907 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r14[26] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r14_reg[27]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4909 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r14[27] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r14_reg[28]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4911 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r14[28] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r14_reg[29]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4913 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r14[29] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r14_reg[30]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4915 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r14[30] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r14_reg[31]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4917 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r14[31] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r11_reg[0]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4919 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r11[0] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r11_reg[1]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4921 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r11[1] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r11_reg[2]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4923 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r11[2] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r11_reg[3]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4925 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r11[3] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r11_reg[4]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4927 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r11[4] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r11_reg[5]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4929 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r11[5] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r11_reg[6]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4931 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r11[6] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r11_reg[7]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4933 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r11[7] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r11_reg[8]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4935 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r11[8] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r11_reg[9]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4937 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r11[9] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r11_reg[10]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4939 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r11[10] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r11_reg[11]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4941 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r11[11] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r11_reg[12]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4943 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r11[12] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r11_reg[13]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4945 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r11[13] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r11_reg[14]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4947 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r11[14] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r11_reg[15]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4949 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r11[15] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r11_reg[16]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4951 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r11[16] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r11_reg[17]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4953 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r11[17] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r11_reg[18]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4955 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r11[18] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r11_reg[19]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4957 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r11[19] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r11_reg[20]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4959 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r11[20] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r11_reg[21]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4961 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r11[21] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r11_reg[22]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4963 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r11[22] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r11_reg[23]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4965 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r11[23] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r11_reg[24]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4967 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r11[24] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r11_reg[25]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4969 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r11[25] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r11_reg[26]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4971 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r11[26] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r11_reg[27]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4973 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r11[27] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r11_reg[28]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4975 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r11[28] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r11_reg[29]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4977 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r11[29] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r11_reg[30]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4979 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r11[30] ) );
  DFF \u_a23_core/u_execute/u_register_bank/r11_reg[31]  ( .D(
        \u_a23_core/u_execute/u_register_bank/n4981 ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\u_a23_core/u_execute/u_register_bank/r11[31] ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_90/U1_1_1  ( .IN0(n16636), .IN1(
        n16635), .COUT(\u_a23_core/u_execute/u_multiply/add_90/carry[2] ), 
        .SUM(\u_a23_core/u_execute/u_multiply/multiplier_bar[1] ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_90/U1_1_2  ( .IN0(n16625), .IN1(
        \u_a23_core/u_execute/u_multiply/add_90/carry[2] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_90/carry[3] ), .SUM(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[2] ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_90/U1_1_3  ( .IN0(n16628), .IN1(
        \u_a23_core/u_execute/u_multiply/add_90/carry[3] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_90/carry[4] ), .SUM(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[3] ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_90/U1_1_4  ( .IN0(n16629), .IN1(
        \u_a23_core/u_execute/u_multiply/add_90/carry[4] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_90/carry[5] ), .SUM(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[4] ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_90/U1_1_5  ( .IN0(n16630), .IN1(
        \u_a23_core/u_execute/u_multiply/add_90/carry[5] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_90/carry[6] ), .SUM(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[5] ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_90/U1_1_6  ( .IN0(n16631), .IN1(
        \u_a23_core/u_execute/u_multiply/add_90/carry[6] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_90/carry[7] ), .SUM(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[6] ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_90/U1_1_7  ( .IN0(n16632), .IN1(
        \u_a23_core/u_execute/u_multiply/add_90/carry[7] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_90/carry[8] ), .SUM(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[7] ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_90/U1_1_8  ( .IN0(n16633), .IN1(
        \u_a23_core/u_execute/u_multiply/add_90/carry[8] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_90/carry[9] ), .SUM(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[8] ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_90/U1_1_9  ( .IN0(n16634), .IN1(
        \u_a23_core/u_execute/u_multiply/add_90/carry[9] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_90/carry[10] ), .SUM(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[9] ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_90/U1_1_10  ( .IN0(n16605), 
        .IN1(\u_a23_core/u_execute/u_multiply/add_90/carry[10] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_90/carry[11] ), .SUM(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[10] ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_90/U1_1_11  ( .IN0(n16606), 
        .IN1(\u_a23_core/u_execute/u_multiply/add_90/carry[11] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_90/carry[12] ), .SUM(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[11] ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_90/U1_1_12  ( .IN0(n16607), 
        .IN1(\u_a23_core/u_execute/u_multiply/add_90/carry[12] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_90/carry[13] ), .SUM(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[12] ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_90/U1_1_13  ( .IN0(n16608), 
        .IN1(\u_a23_core/u_execute/u_multiply/add_90/carry[13] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_90/carry[14] ), .SUM(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[13] ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_90/U1_1_14  ( .IN0(n16609), 
        .IN1(\u_a23_core/u_execute/u_multiply/add_90/carry[14] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_90/carry[15] ), .SUM(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[14] ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_90/U1_1_15  ( .IN0(n16610), 
        .IN1(\u_a23_core/u_execute/u_multiply/add_90/carry[15] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_90/carry[16] ), .SUM(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[15] ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_90/U1_1_16  ( .IN0(n16611), 
        .IN1(\u_a23_core/u_execute/u_multiply/add_90/carry[16] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_90/carry[17] ), .SUM(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[16] ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_90/U1_1_17  ( .IN0(n16612), 
        .IN1(\u_a23_core/u_execute/u_multiply/add_90/carry[17] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_90/carry[18] ), .SUM(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[17] ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_90/U1_1_18  ( .IN0(n16613), 
        .IN1(\u_a23_core/u_execute/u_multiply/add_90/carry[18] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_90/carry[19] ), .SUM(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[18] ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_90/U1_1_19  ( .IN0(n16614), 
        .IN1(\u_a23_core/u_execute/u_multiply/add_90/carry[19] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_90/carry[20] ), .SUM(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[19] ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_90/U1_1_20  ( .IN0(n16615), 
        .IN1(\u_a23_core/u_execute/u_multiply/add_90/carry[20] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_90/carry[21] ), .SUM(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[20] ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_90/U1_1_21  ( .IN0(n16616), 
        .IN1(\u_a23_core/u_execute/u_multiply/add_90/carry[21] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_90/carry[22] ), .SUM(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[21] ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_90/U1_1_22  ( .IN0(n16617), 
        .IN1(\u_a23_core/u_execute/u_multiply/add_90/carry[22] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_90/carry[23] ), .SUM(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[22] ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_90/U1_1_23  ( .IN0(n16618), 
        .IN1(\u_a23_core/u_execute/u_multiply/add_90/carry[23] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_90/carry[24] ), .SUM(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[23] ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_90/U1_1_24  ( .IN0(n16619), 
        .IN1(\u_a23_core/u_execute/u_multiply/add_90/carry[24] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_90/carry[25] ), .SUM(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[24] ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_90/U1_1_25  ( .IN0(n16620), 
        .IN1(\u_a23_core/u_execute/u_multiply/add_90/carry[25] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_90/carry[26] ), .SUM(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[25] ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_90/U1_1_26  ( .IN0(n16621), 
        .IN1(\u_a23_core/u_execute/u_multiply/add_90/carry[26] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_90/carry[27] ), .SUM(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[26] ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_90/U1_1_27  ( .IN0(n16622), 
        .IN1(\u_a23_core/u_execute/u_multiply/add_90/carry[27] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_90/carry[28] ), .SUM(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[27] ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_90/U1_1_28  ( .IN0(n16623), 
        .IN1(\u_a23_core/u_execute/u_multiply/add_90/carry[28] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_90/carry[29] ), .SUM(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[28] ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_90/U1_1_29  ( .IN0(n16624), 
        .IN1(\u_a23_core/u_execute/u_multiply/add_90/carry[29] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_90/carry[30] ), .SUM(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[29] ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_90/U1_1_30  ( .IN0(n16626), 
        .IN1(\u_a23_core/u_execute/u_multiply/add_90/carry[30] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_90/carry[31] ), .SUM(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[30] ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_90/U1_1_31  ( .IN0(n16627), 
        .IN1(\u_a23_core/u_execute/u_multiply/add_90/carry[31] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_90/carry[32] ), .SUM(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[31] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_100/U1_1  ( .CIN(
        \u_a23_core/u_execute/u_multiply/product[35] ), .IN0(
        \u_a23_core/u_execute/u_multiply/sum34_b[1] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_100/carry[1] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_100/carry[2] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum[1] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_100/U1_2  ( .CIN(
        \u_a23_core/u_execute/u_multiply/product[36] ), .IN0(
        \u_a23_core/u_execute/u_multiply/sum34_b[2] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_100/carry[2] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_100/carry[3] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum[2] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_100/U1_3  ( .CIN(
        \u_a23_core/u_execute/u_multiply/product[37] ), .IN0(
        \u_a23_core/u_execute/u_multiply/sum34_b[3] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_100/carry[3] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_100/carry[4] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum[3] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_100/U1_4  ( .CIN(
        \u_a23_core/u_execute/u_multiply/product[38] ), .IN0(
        \u_a23_core/u_execute/u_multiply/sum34_b[4] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_100/carry[4] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_100/carry[5] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum[4] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_100/U1_5  ( .CIN(
        \u_a23_core/u_execute/u_multiply/product[39] ), .IN0(
        \u_a23_core/u_execute/u_multiply/sum34_b[5] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_100/carry[5] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_100/carry[6] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum[5] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_100/U1_6  ( .CIN(
        \u_a23_core/u_execute/u_multiply/product[40] ), .IN0(
        \u_a23_core/u_execute/u_multiply/sum34_b[6] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_100/carry[6] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_100/carry[7] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum[6] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_100/U1_7  ( .CIN(
        \u_a23_core/u_execute/u_multiply/product[41] ), .IN0(
        \u_a23_core/u_execute/u_multiply/sum34_b[7] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_100/carry[7] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_100/carry[8] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum[7] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_100/U1_8  ( .CIN(
        \u_a23_core/u_execute/u_multiply/product[42] ), .IN0(
        \u_a23_core/u_execute/u_multiply/sum34_b[8] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_100/carry[8] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_100/carry[9] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum[8] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_100/U1_9  ( .CIN(
        \u_a23_core/u_execute/u_multiply/product[43] ), .IN0(
        \u_a23_core/u_execute/u_multiply/sum34_b[9] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_100/carry[9] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_100/carry[10] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum[9] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_100/U1_10  ( .CIN(
        \u_a23_core/u_execute/u_multiply/product[44] ), .IN0(
        \u_a23_core/u_execute/u_multiply/sum34_b[10] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_100/carry[10] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_100/carry[11] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum[10] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_100/U1_11  ( .CIN(
        \u_a23_core/u_execute/u_multiply/product[45] ), .IN0(
        \u_a23_core/u_execute/u_multiply/sum34_b[11] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_100/carry[11] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_100/carry[12] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum[11] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_100/U1_12  ( .CIN(
        \u_a23_core/u_execute/u_multiply/product[46] ), .IN0(
        \u_a23_core/u_execute/u_multiply/sum34_b[12] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_100/carry[12] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_100/carry[13] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum[12] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_100/U1_13  ( .CIN(
        \u_a23_core/u_execute/u_multiply/product[47] ), .IN0(
        \u_a23_core/u_execute/u_multiply/sum34_b[13] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_100/carry[13] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_100/carry[14] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum[13] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_100/U1_14  ( .CIN(
        \u_a23_core/u_execute/u_multiply/product[48] ), .IN0(
        \u_a23_core/u_execute/u_multiply/sum34_b[14] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_100/carry[14] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_100/carry[15] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum[14] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_100/U1_15  ( .CIN(
        \u_a23_core/u_execute/u_multiply/product[49] ), .IN0(
        \u_a23_core/u_execute/u_multiply/sum34_b[15] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_100/carry[15] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_100/carry[16] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum[15] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_100/U1_16  ( .CIN(
        \u_a23_core/u_execute/u_multiply/product[50] ), .IN0(
        \u_a23_core/u_execute/u_multiply/sum34_b[16] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_100/carry[16] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_100/carry[17] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum[16] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_100/U1_17  ( .CIN(
        \u_a23_core/u_execute/u_multiply/product[51] ), .IN0(
        \u_a23_core/u_execute/u_multiply/sum34_b[17] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_100/carry[17] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_100/carry[18] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum[17] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_100/U1_18  ( .CIN(
        \u_a23_core/u_execute/u_multiply/product[52] ), .IN0(
        \u_a23_core/u_execute/u_multiply/sum34_b[18] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_100/carry[18] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_100/carry[19] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum[18] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_100/U1_19  ( .CIN(
        \u_a23_core/u_execute/u_multiply/product[53] ), .IN0(
        \u_a23_core/u_execute/u_multiply/sum34_b[19] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_100/carry[19] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_100/carry[20] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum[19] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_100/U1_20  ( .CIN(
        \u_a23_core/u_execute/u_multiply/product[54] ), .IN0(
        \u_a23_core/u_execute/u_multiply/sum34_b[20] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_100/carry[20] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_100/carry[21] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum[20] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_100/U1_21  ( .CIN(
        \u_a23_core/u_execute/u_multiply/product[55] ), .IN0(
        \u_a23_core/u_execute/u_multiply/sum34_b[21] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_100/carry[21] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_100/carry[22] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum[21] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_100/U1_22  ( .CIN(
        \u_a23_core/u_execute/u_multiply/product[56] ), .IN0(
        \u_a23_core/u_execute/u_multiply/sum34_b[22] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_100/carry[22] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_100/carry[23] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum[22] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_100/U1_23  ( .CIN(
        \u_a23_core/u_execute/u_multiply/product[57] ), .IN0(
        \u_a23_core/u_execute/u_multiply/sum34_b[23] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_100/carry[23] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_100/carry[24] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum[23] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_100/U1_24  ( .CIN(
        \u_a23_core/u_execute/u_multiply/product[58] ), .IN0(
        \u_a23_core/u_execute/u_multiply/sum34_b[24] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_100/carry[24] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_100/carry[25] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum[24] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_100/U1_25  ( .CIN(
        \u_a23_core/u_execute/u_multiply/product[59] ), .IN0(
        \u_a23_core/u_execute/u_multiply/sum34_b[25] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_100/carry[25] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_100/carry[26] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum[25] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_100/U1_26  ( .CIN(
        \u_a23_core/u_execute/u_multiply/product[60] ), .IN0(
        \u_a23_core/u_execute/u_multiply/sum34_b[26] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_100/carry[26] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_100/carry[27] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum[26] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_100/U1_27  ( .CIN(
        \u_a23_core/u_execute/u_multiply/product[61] ), .IN0(
        \u_a23_core/u_execute/u_multiply/sum34_b[27] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_100/carry[27] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_100/carry[28] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum[27] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_100/U1_28  ( .CIN(
        \u_a23_core/u_execute/u_multiply/product[62] ), .IN0(
        \u_a23_core/u_execute/u_multiply/sum34_b[28] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_100/carry[28] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_100/carry[29] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum[28] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_100/U1_29  ( .CIN(
        \u_a23_core/u_execute/u_multiply/product[63] ), .IN0(
        \u_a23_core/u_execute/u_multiply/sum34_b[29] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_100/carry[29] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_100/carry[30] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum[29] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_100/U1_30  ( .CIN(
        \u_a23_core/u_execute/u_multiply/product[64] ), .IN0(
        \u_a23_core/u_execute/u_multiply/sum34_b[30] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_100/carry[30] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_100/carry[31] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum[30] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_100/U1_31  ( .CIN(
        \u_a23_core/u_execute/u_multiply/product[65] ), .IN0(
        \u_a23_core/u_execute/u_multiply/sum34_b[31] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_100/carry[31] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_100/carry[32] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum[31] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_100/U1_32  ( .CIN(
        \u_a23_core/u_execute/u_multiply/product[66] ), .IN0(
        \u_a23_core/u_execute/u_multiply/sum34_b[33] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_100/carry[32] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_100/carry[33] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum[32] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_100/U1_33  ( .CIN(
        \u_a23_core/u_execute/u_multiply/product[67] ), .IN0(
        \u_a23_core/u_execute/u_multiply/sum34_b[33] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_100/carry[33] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum[33] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_105/U1_1  ( .CIN(
        \u_a23_core/u_execute/multiply_out[1] ), .IN0(
        \u_a23_core/u_execute/rs[1] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_105/carry[1] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_105/carry[2] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum_acc1[1] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_105/U1_2  ( .CIN(
        \u_a23_core/u_execute/multiply_out[2] ), .IN0(
        \u_a23_core/u_execute/rs[2] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_105/carry[2] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_105/carry[3] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum_acc1[2] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_105/U1_3  ( .CIN(
        \u_a23_core/u_execute/multiply_out[3] ), .IN0(
        \u_a23_core/u_execute/rs[3] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_105/carry[3] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_105/carry[4] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum_acc1[3] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_105/U1_4  ( .CIN(
        \u_a23_core/u_execute/multiply_out[4] ), .IN0(
        \u_a23_core/u_execute/rs[4] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_105/carry[4] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_105/carry[5] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum_acc1[4] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_105/U1_5  ( .CIN(
        \u_a23_core/u_execute/multiply_out[5] ), .IN0(
        \u_a23_core/u_execute/rs[5] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_105/carry[5] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_105/carry[6] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum_acc1[5] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_105/U1_6  ( .CIN(
        \u_a23_core/u_execute/multiply_out[6] ), .IN0(
        \u_a23_core/u_execute/rs[6] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_105/carry[6] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_105/carry[7] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum_acc1[6] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_105/U1_7  ( .CIN(
        \u_a23_core/u_execute/multiply_out[7] ), .IN0(
        \u_a23_core/u_execute/rs[7] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_105/carry[7] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_105/carry[8] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum_acc1[7] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_105/U1_8  ( .CIN(
        \u_a23_core/u_execute/multiply_out[8] ), .IN0(
        \u_a23_core/u_execute/rs[8] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_105/carry[8] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_105/carry[9] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum_acc1[8] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_105/U1_9  ( .CIN(
        \u_a23_core/u_execute/multiply_out[9] ), .IN0(
        \u_a23_core/u_execute/rs[9] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_105/carry[9] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_105/carry[10] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum_acc1[9] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_105/U1_10  ( .CIN(
        \u_a23_core/u_execute/multiply_out[10] ), .IN0(
        \u_a23_core/u_execute/rs[10] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_105/carry[10] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_105/carry[11] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum_acc1[10] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_105/U1_11  ( .CIN(
        \u_a23_core/u_execute/multiply_out[11] ), .IN0(
        \u_a23_core/u_execute/rs[11] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_105/carry[11] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_105/carry[12] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum_acc1[11] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_105/U1_12  ( .CIN(
        \u_a23_core/u_execute/multiply_out[12] ), .IN0(
        \u_a23_core/u_execute/rs[12] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_105/carry[12] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_105/carry[13] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum_acc1[12] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_105/U1_13  ( .CIN(
        \u_a23_core/u_execute/multiply_out[13] ), .IN0(
        \u_a23_core/u_execute/rs[13] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_105/carry[13] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_105/carry[14] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum_acc1[13] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_105/U1_14  ( .CIN(
        \u_a23_core/u_execute/multiply_out[14] ), .IN0(
        \u_a23_core/u_execute/rs[14] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_105/carry[14] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_105/carry[15] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum_acc1[14] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_105/U1_15  ( .CIN(
        \u_a23_core/u_execute/multiply_out[15] ), .IN0(
        \u_a23_core/u_execute/rs[15] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_105/carry[15] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_105/carry[16] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum_acc1[15] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_105/U1_16  ( .CIN(
        \u_a23_core/u_execute/multiply_out[16] ), .IN0(
        \u_a23_core/u_execute/rs[16] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_105/carry[16] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_105/carry[17] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum_acc1[16] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_105/U1_17  ( .CIN(
        \u_a23_core/u_execute/multiply_out[17] ), .IN0(
        \u_a23_core/u_execute/rs[17] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_105/carry[17] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_105/carry[18] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum_acc1[17] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_105/U1_18  ( .CIN(
        \u_a23_core/u_execute/multiply_out[18] ), .IN0(
        \u_a23_core/u_execute/rs[18] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_105/carry[18] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_105/carry[19] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum_acc1[18] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_105/U1_19  ( .CIN(
        \u_a23_core/u_execute/multiply_out[19] ), .IN0(
        \u_a23_core/u_execute/rs[19] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_105/carry[19] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_105/carry[20] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum_acc1[19] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_105/U1_20  ( .CIN(
        \u_a23_core/u_execute/multiply_out[20] ), .IN0(
        \u_a23_core/u_execute/rs[20] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_105/carry[20] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_105/carry[21] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum_acc1[20] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_105/U1_21  ( .CIN(
        \u_a23_core/u_execute/multiply_out[21] ), .IN0(
        \u_a23_core/u_execute/rs[21] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_105/carry[21] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_105/carry[22] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum_acc1[21] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_105/U1_22  ( .CIN(
        \u_a23_core/u_execute/multiply_out[22] ), .IN0(
        \u_a23_core/u_execute/rs[22] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_105/carry[22] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_105/carry[23] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum_acc1[22] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_105/U1_23  ( .CIN(
        \u_a23_core/u_execute/multiply_out[23] ), .IN0(
        \u_a23_core/u_execute/rs[23] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_105/carry[23] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_105/carry[24] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum_acc1[23] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_105/U1_24  ( .CIN(
        \u_a23_core/u_execute/multiply_out[24] ), .IN0(
        \u_a23_core/u_execute/rs[24] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_105/carry[24] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_105/carry[25] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum_acc1[24] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_105/U1_25  ( .CIN(
        \u_a23_core/u_execute/multiply_out[25] ), .IN0(
        \u_a23_core/u_execute/rs[25] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_105/carry[25] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_105/carry[26] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum_acc1[25] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_105/U1_26  ( .CIN(
        \u_a23_core/u_execute/multiply_out[26] ), .IN0(
        \u_a23_core/u_execute/rs[26] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_105/carry[26] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_105/carry[27] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum_acc1[26] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_105/U1_27  ( .CIN(
        \u_a23_core/u_execute/multiply_out[27] ), .IN0(
        \u_a23_core/u_execute/rs[27] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_105/carry[27] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_105/carry[28] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum_acc1[27] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_105/U1_28  ( .CIN(
        \u_a23_core/u_execute/multiply_out[28] ), .IN0(
        \u_a23_core/u_execute/rs[28] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_105/carry[28] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_105/carry[29] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum_acc1[28] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_105/U1_29  ( .CIN(
        \u_a23_core/u_execute/multiply_out[29] ), .IN0(
        \u_a23_core/u_execute/rs[29] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_105/carry[29] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_105/carry[30] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum_acc1[29] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_105/U1_30  ( .CIN(
        \u_a23_core/u_execute/multiply_out[30] ), .IN0(
        \u_a23_core/u_execute/rs[30] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_105/carry[30] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_105/carry[31] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum_acc1[30] ) );
  FADDER \u_a23_core/u_execute/u_multiply/add_105/U1_31  ( .CIN(
        \u_a23_core/u_execute/multiply_out[31] ), .IN0(
        \u_a23_core/u_execute/rs[31] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_105/carry[31] ), .SUM(
        \u_a23_core/u_execute/u_multiply/sum_acc1[31] ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_139/U1_1_1  ( .IN0(
        \u_a23_core/u_execute/u_multiply/count[1] ), .IN1(
        \u_a23_core/u_execute/u_multiply/count[0] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_139/carry[2] ), .SUM(
        \u_a23_core/u_execute/u_multiply/N55 ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_139/U1_1_2  ( .IN0(
        \u_a23_core/u_execute/u_multiply/count[2] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_139/carry[2] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_139/carry[3] ), .SUM(
        \u_a23_core/u_execute/u_multiply/N56 ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_139/U1_1_3  ( .IN0(
        \u_a23_core/u_execute/u_multiply/count[3] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_139/carry[3] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_139/carry[4] ), .SUM(
        \u_a23_core/u_execute/u_multiply/N57 ) );
  HADDER \u_a23_core/u_execute/u_multiply/add_139/U1_1_4  ( .IN0(
        \u_a23_core/u_execute/u_multiply/count[4] ), .IN1(
        \u_a23_core/u_execute/u_multiply/add_139/carry[4] ), .COUT(
        \u_a23_core/u_execute/u_multiply/add_139/carry[5] ), .SUM(
        \u_a23_core/u_execute/u_multiply/N58 ) );
  FADDER \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/U1_0  ( .CIN(
        \u_a23_core/u_execute/u_alu/a[0] ), .IN0(
        \u_a23_core/u_execute/u_alu/b_not[0] ), .IN1(
        \u_a23_core/u_execute/u_alu/carry_in ), .COUT(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[1] ), .SUM(
        \u_a23_core/u_execute/u_alu/fadder_out[0] ) );
  FADDER \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/U1_1  ( .CIN(
        \u_a23_core/u_execute/u_alu/a[1] ), .IN0(
        \u_a23_core/u_execute/u_alu/b_not[1] ), .IN1(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[1] ), .COUT(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[2] ), .SUM(
        \u_a23_core/u_execute/u_alu/fadder_out[1] ) );
  FADDER \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/U1_2  ( .CIN(
        \u_a23_core/u_execute/u_alu/a[2] ), .IN0(
        \u_a23_core/u_execute/u_alu/b_not[2] ), .IN1(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[2] ), .COUT(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[3] ), .SUM(
        \u_a23_core/u_execute/u_alu/fadder_out[2] ) );
  FADDER \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/U1_3  ( .CIN(
        \u_a23_core/u_execute/u_alu/a[3] ), .IN0(
        \u_a23_core/u_execute/u_alu/b_not[3] ), .IN1(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[3] ), .COUT(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[4] ), .SUM(
        \u_a23_core/u_execute/u_alu/fadder_out[3] ) );
  FADDER \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/U1_4  ( .CIN(
        \u_a23_core/u_execute/u_alu/a[4] ), .IN0(
        \u_a23_core/u_execute/u_alu/b_not[4] ), .IN1(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[4] ), .COUT(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[5] ), .SUM(
        \u_a23_core/u_execute/u_alu/fadder_out[4] ) );
  FADDER \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/U1_5  ( .CIN(
        \u_a23_core/u_execute/u_alu/a[5] ), .IN0(
        \u_a23_core/u_execute/u_alu/b_not[5] ), .IN1(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[5] ), .COUT(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[6] ), .SUM(
        \u_a23_core/u_execute/u_alu/fadder_out[5] ) );
  FADDER \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/U1_6  ( .CIN(
        \u_a23_core/u_execute/u_alu/a[6] ), .IN0(
        \u_a23_core/u_execute/u_alu/b_not[6] ), .IN1(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[6] ), .COUT(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[7] ), .SUM(
        \u_a23_core/u_execute/u_alu/fadder_out[6] ) );
  FADDER \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/U1_7  ( .CIN(
        \u_a23_core/u_execute/u_alu/a[7] ), .IN0(
        \u_a23_core/u_execute/u_alu/b_not[7] ), .IN1(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[7] ), .COUT(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[8] ), .SUM(
        \u_a23_core/u_execute/u_alu/fadder_out[7] ) );
  FADDER \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/U1_8  ( .CIN(
        \u_a23_core/u_execute/u_alu/a[8] ), .IN0(
        \u_a23_core/u_execute/u_alu/b_not[8] ), .IN1(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[8] ), .COUT(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[9] ), .SUM(
        \u_a23_core/u_execute/u_alu/fadder_out[8] ) );
  FADDER \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/U1_9  ( .CIN(
        \u_a23_core/u_execute/u_alu/a[9] ), .IN0(
        \u_a23_core/u_execute/u_alu/b_not[9] ), .IN1(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[9] ), .COUT(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[10] ), .SUM(
        \u_a23_core/u_execute/u_alu/fadder_out[9] ) );
  FADDER \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/U1_10  ( .CIN(
        \u_a23_core/u_execute/u_alu/a[10] ), .IN0(
        \u_a23_core/u_execute/u_alu/b_not[10] ), .IN1(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[10] ), .COUT(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[11] ), .SUM(
        \u_a23_core/u_execute/u_alu/fadder_out[10] ) );
  FADDER \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/U1_11  ( .CIN(
        \u_a23_core/u_execute/u_alu/a[11] ), .IN0(
        \u_a23_core/u_execute/u_alu/b_not[11] ), .IN1(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[11] ), .COUT(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[12] ), .SUM(
        \u_a23_core/u_execute/u_alu/fadder_out[11] ) );
  FADDER \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/U1_12  ( .CIN(
        \u_a23_core/u_execute/u_alu/a[12] ), .IN0(
        \u_a23_core/u_execute/u_alu/b_not[12] ), .IN1(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[12] ), .COUT(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[13] ), .SUM(
        \u_a23_core/u_execute/u_alu/fadder_out[12] ) );
  FADDER \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/U1_13  ( .CIN(
        \u_a23_core/u_execute/u_alu/a[13] ), .IN0(
        \u_a23_core/u_execute/u_alu/b_not[13] ), .IN1(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[13] ), .COUT(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[14] ), .SUM(
        \u_a23_core/u_execute/u_alu/fadder_out[13] ) );
  FADDER \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/U1_14  ( .CIN(
        \u_a23_core/u_execute/u_alu/a[14] ), .IN0(
        \u_a23_core/u_execute/u_alu/b_not[14] ), .IN1(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[14] ), .COUT(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[15] ), .SUM(
        \u_a23_core/u_execute/u_alu/fadder_out[14] ) );
  FADDER \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/U1_15  ( .CIN(
        \u_a23_core/u_execute/u_alu/a[15] ), .IN0(
        \u_a23_core/u_execute/u_alu/b_not[15] ), .IN1(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[15] ), .COUT(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[16] ), .SUM(
        \u_a23_core/u_execute/u_alu/fadder_out[15] ) );
  FADDER \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/U1_16  ( .CIN(
        \u_a23_core/u_execute/u_alu/a[16] ), .IN0(
        \u_a23_core/u_execute/u_alu/b_not[16] ), .IN1(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[16] ), .COUT(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[17] ), .SUM(
        \u_a23_core/u_execute/u_alu/fadder_out[16] ) );
  FADDER \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/U1_17  ( .CIN(
        \u_a23_core/u_execute/u_alu/a[17] ), .IN0(
        \u_a23_core/u_execute/u_alu/b_not[17] ), .IN1(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[17] ), .COUT(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[18] ), .SUM(
        \u_a23_core/u_execute/u_alu/fadder_out[17] ) );
  FADDER \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/U1_18  ( .CIN(
        \u_a23_core/u_execute/u_alu/a[18] ), .IN0(
        \u_a23_core/u_execute/u_alu/b_not[18] ), .IN1(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[18] ), .COUT(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[19] ), .SUM(
        \u_a23_core/u_execute/u_alu/fadder_out[18] ) );
  FADDER \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/U1_19  ( .CIN(
        \u_a23_core/u_execute/u_alu/a[19] ), .IN0(
        \u_a23_core/u_execute/u_alu/b_not[19] ), .IN1(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[19] ), .COUT(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[20] ), .SUM(
        \u_a23_core/u_execute/u_alu/fadder_out[19] ) );
  FADDER \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/U1_20  ( .CIN(
        \u_a23_core/u_execute/u_alu/a[20] ), .IN0(
        \u_a23_core/u_execute/u_alu/b_not[20] ), .IN1(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[20] ), .COUT(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[21] ), .SUM(
        \u_a23_core/u_execute/u_alu/fadder_out[20] ) );
  FADDER \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/U1_21  ( .CIN(
        \u_a23_core/u_execute/u_alu/a[21] ), .IN0(
        \u_a23_core/u_execute/u_alu/b_not[21] ), .IN1(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[21] ), .COUT(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[22] ), .SUM(
        \u_a23_core/u_execute/u_alu/fadder_out[21] ) );
  FADDER \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/U1_22  ( .CIN(
        \u_a23_core/u_execute/u_alu/a[22] ), .IN0(
        \u_a23_core/u_execute/u_alu/b_not[22] ), .IN1(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[22] ), .COUT(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[23] ), .SUM(
        \u_a23_core/u_execute/u_alu/fadder_out[22] ) );
  FADDER \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/U1_23  ( .CIN(
        \u_a23_core/u_execute/u_alu/a[23] ), .IN0(
        \u_a23_core/u_execute/u_alu/b_not[23] ), .IN1(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[23] ), .COUT(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[24] ), .SUM(
        \u_a23_core/u_execute/u_alu/fadder_out[23] ) );
  FADDER \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/U1_24  ( .CIN(
        \u_a23_core/u_execute/u_alu/a[24] ), .IN0(
        \u_a23_core/u_execute/u_alu/b_not[24] ), .IN1(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[24] ), .COUT(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[25] ), .SUM(
        \u_a23_core/u_execute/u_alu/fadder_out[24] ) );
  FADDER \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/U1_25  ( .CIN(
        \u_a23_core/u_execute/u_alu/a[25] ), .IN0(
        \u_a23_core/u_execute/u_alu/b_not[25] ), .IN1(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[25] ), .COUT(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[26] ), .SUM(
        \u_a23_core/u_execute/u_alu/fadder_out[25] ) );
  FADDER \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/U1_26  ( .CIN(
        \u_a23_core/u_execute/u_alu/a[26] ), .IN0(
        \u_a23_core/u_execute/u_alu/b_not[26] ), .IN1(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[26] ), .COUT(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[27] ), .SUM(
        \u_a23_core/u_execute/u_alu/fadder_out[26] ) );
  FADDER \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/U1_27  ( .CIN(
        \u_a23_core/u_execute/u_alu/a[27] ), .IN0(
        \u_a23_core/u_execute/u_alu/b_not[27] ), .IN1(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[27] ), .COUT(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[28] ), .SUM(
        \u_a23_core/u_execute/u_alu/fadder_out[27] ) );
  FADDER \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/U1_28  ( .CIN(
        \u_a23_core/u_execute/u_alu/a[28] ), .IN0(
        \u_a23_core/u_execute/u_alu/b_not[28] ), .IN1(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[28] ), .COUT(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[29] ), .SUM(
        \u_a23_core/u_execute/u_alu/fadder_out[28] ) );
  FADDER \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/U1_29  ( .CIN(
        \u_a23_core/u_execute/u_alu/a[29] ), .IN0(
        \u_a23_core/u_execute/u_alu/b_not[29] ), .IN1(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[29] ), .COUT(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[30] ), .SUM(
        \u_a23_core/u_execute/u_alu/fadder_out[29] ) );
  FADDER \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/U1_30  ( .CIN(
        \u_a23_core/u_execute/u_alu/a[30] ), .IN0(
        \u_a23_core/u_execute/u_alu/b_not[30] ), .IN1(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[30] ), .COUT(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[31] ), .SUM(
        \u_a23_core/u_execute/u_alu/fadder_out[30] ) );
  FADDER \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/U1_31  ( .CIN(
        \u_a23_core/u_execute/u_alu/a[31] ), .IN0(
        \u_a23_core/u_execute/u_alu/b_not[31] ), .IN1(
        \u_a23_core/u_execute/u_alu/add_1_root_add_121_2/carry[31] ), .COUT(
        \u_a23_core/u_execute/u_alu/fadder_out[32] ), .SUM(
        \u_a23_core/u_execute/u_alu/fadder_out[31] ) );
  FADDER \u_a23_core/u_decode/add_11_root_add_415_15/U1_0  ( .CIN(
        \u_a23_core/u_decode/instruction[5] ), .IN0(
        \u_a23_core/u_decode/instruction[4] ), .IN1(
        \u_a23_core/u_decode/instruction[6] ), .COUT(
        \u_a23_core/u_decode/N528 ), .SUM(\u_a23_core/u_decode/N527 ) );
  FADDER \u_a23_core/u_decode/add_10_root_add_415_15/U1_0  ( .CIN(
        \u_a23_core/rm_sel_nxt[2] ), .IN0(\u_a23_core/rm_sel_nxt[1] ), .IN1(
        \u_a23_core/rm_sel_nxt[3] ), .COUT(\u_a23_core/u_decode/N533 ), .SUM(
        \u_a23_core/u_decode/N532 ) );
  FADDER \u_a23_core/u_decode/add_9_root_add_415_15/U1_0  ( .CIN(
        \u_a23_core/u_decode/N518 ), .IN0(\u_a23_core/u_decode/N520 ), .IN1(
        \u_a23_core/rm_sel_nxt[0] ), .COUT(
        \u_a23_core/u_decode/add_9_root_add_415_15/carry[1] ), .SUM(
        \u_a23_core/u_decode/N537 ) );
  FADDER \u_a23_core/u_decode/add_9_root_add_415_15/U1_1  ( .CIN(
        \u_a23_core/u_decode/N519 ), .IN0(\u_a23_core/u_decode/N521 ), .IN1(
        \u_a23_core/u_decode/add_9_root_add_415_15/carry[1] ), .COUT(
        \u_a23_core/u_decode/N539 ), .SUM(\u_a23_core/u_decode/N538 ) );
  FADDER \u_a23_core/u_decode/add_8_root_add_415_15/U1_1  ( .CIN(
        \u_a23_core/u_decode/N524 ), .IN0(\u_a23_core/u_decode/N528 ), .IN1(
        \u_a23_core/u_decode/add_8_root_add_415_15/carry[1] ), .COUT(
        \u_a23_core/u_decode/N544 ), .SUM(\u_a23_core/u_decode/N543 ) );
  FADDER \u_a23_core/u_decode/add_7_root_add_415_15/U1_1  ( .CIN(
        \u_a23_core/u_decode/N533 ), .IN0(\u_a23_core/u_decode/N538 ), .IN1(
        \u_a23_core/u_decode/add_7_root_add_415_15/carry[1] ), .COUT(
        \u_a23_core/u_decode/add_7_root_add_415_15/carry[2] ), .SUM(
        \u_a23_core/u_decode/N548 ) );
  FADDER \u_a23_core/u_decode/add_6_root_add_415_15/U1_1  ( .CIN(
        \u_a23_core/u_decode/N543 ), .IN0(\u_a23_core/u_decode/N548 ), .IN1(
        \u_a23_core/u_decode/add_6_root_add_415_15/carry[1] ), .COUT(
        \u_a23_core/u_decode/add_6_root_add_415_15/carry[2] ), .SUM(
        \u_a23_core/u_decode/mtrans_num_registers[1] ) );
  FADDER \u_a23_core/u_decode/add_6_root_add_415_15/U1_2  ( .CIN(
        \u_a23_core/u_decode/N544 ), .IN0(\u_a23_core/u_decode/N549 ), .IN1(
        \u_a23_core/u_decode/add_6_root_add_415_15/carry[2] ), .COUT(
        \u_a23_core/u_decode/add_6_root_add_415_15/carry[3] ), .SUM(
        \u_a23_core/u_decode/mtrans_num_registers[2] ) );
  OR U1 ( .A(\u_a23_core/u_execute/sub_166/carry[10] ), .B(
        \u_a23_core/u_execute/pc[10] ), .Z(
        \u_a23_core/u_execute/sub_166/carry[11] ) );
  XNOR U2 ( .A(\u_a23_core/u_execute/pc[10] ), .B(
        \u_a23_core/u_execute/sub_166/carry[10] ), .Z(
        \u_a23_core/u_execute/pc_minus4[10] ) );
  OR U3 ( .A(\u_a23_core/u_execute/sub_166/carry[11] ), .B(
        \u_a23_core/u_execute/pc[11] ), .Z(
        \u_a23_core/u_execute/sub_166/carry[12] ) );
  XNOR U4 ( .A(\u_a23_core/u_execute/pc[11] ), .B(
        \u_a23_core/u_execute/sub_166/carry[11] ), .Z(
        \u_a23_core/u_execute/pc_minus4[11] ) );
  OR U5 ( .A(\u_a23_core/u_execute/sub_166/carry[12] ), .B(
        \u_a23_core/u_execute/pc[12] ), .Z(
        \u_a23_core/u_execute/sub_166/carry[13] ) );
  XNOR U6 ( .A(\u_a23_core/u_execute/pc[12] ), .B(
        \u_a23_core/u_execute/sub_166/carry[12] ), .Z(
        \u_a23_core/u_execute/pc_minus4[12] ) );
  OR U7 ( .A(\u_a23_core/u_execute/sub_166/carry[13] ), .B(
        \u_a23_core/u_execute/pc[13] ), .Z(
        \u_a23_core/u_execute/sub_166/carry[14] ) );
  XNOR U8 ( .A(\u_a23_core/u_execute/pc[13] ), .B(
        \u_a23_core/u_execute/sub_166/carry[13] ), .Z(
        \u_a23_core/u_execute/pc_minus4[13] ) );
  OR U9 ( .A(\u_a23_core/u_execute/sub_166/carry[14] ), .B(
        \u_a23_core/u_execute/pc[14] ), .Z(
        \u_a23_core/u_execute/sub_166/carry[15] ) );
  XNOR U10 ( .A(\u_a23_core/u_execute/pc[14] ), .B(
        \u_a23_core/u_execute/sub_166/carry[14] ), .Z(
        \u_a23_core/u_execute/pc_minus4[14] ) );
  OR U11 ( .A(\u_a23_core/u_execute/sub_166/carry[15] ), .B(
        \u_a23_core/u_execute/pc[15] ), .Z(
        \u_a23_core/u_execute/sub_166/carry[16] ) );
  XNOR U12 ( .A(\u_a23_core/u_execute/pc[15] ), .B(
        \u_a23_core/u_execute/sub_166/carry[15] ), .Z(
        \u_a23_core/u_execute/pc_minus4[15] ) );
  OR U13 ( .A(\u_a23_core/u_execute/sub_166/carry[16] ), .B(
        \u_a23_core/u_execute/pc[16] ), .Z(
        \u_a23_core/u_execute/sub_166/carry[17] ) );
  XNOR U14 ( .A(\u_a23_core/u_execute/pc[16] ), .B(
        \u_a23_core/u_execute/sub_166/carry[16] ), .Z(
        \u_a23_core/u_execute/pc_minus4[16] ) );
  OR U15 ( .A(\u_a23_core/u_execute/sub_166/carry[17] ), .B(
        \u_a23_core/u_execute/pc[17] ), .Z(
        \u_a23_core/u_execute/sub_166/carry[18] ) );
  XNOR U16 ( .A(\u_a23_core/u_execute/pc[17] ), .B(
        \u_a23_core/u_execute/sub_166/carry[17] ), .Z(
        \u_a23_core/u_execute/pc_minus4[17] ) );
  OR U17 ( .A(\u_a23_core/u_execute/sub_166/carry[18] ), .B(
        \u_a23_core/u_execute/pc[18] ), .Z(
        \u_a23_core/u_execute/sub_166/carry[19] ) );
  XNOR U18 ( .A(\u_a23_core/u_execute/pc[18] ), .B(
        \u_a23_core/u_execute/sub_166/carry[18] ), .Z(
        \u_a23_core/u_execute/pc_minus4[18] ) );
  OR U19 ( .A(\u_a23_core/u_execute/sub_166/carry[19] ), .B(
        \u_a23_core/u_execute/pc[19] ), .Z(
        \u_a23_core/u_execute/sub_166/carry[20] ) );
  XNOR U20 ( .A(\u_a23_core/u_execute/pc[19] ), .B(
        \u_a23_core/u_execute/sub_166/carry[19] ), .Z(
        \u_a23_core/u_execute/pc_minus4[19] ) );
  OR U21 ( .A(\u_a23_core/u_execute/sub_166/carry[20] ), .B(
        \u_a23_core/u_execute/pc[20] ), .Z(
        \u_a23_core/u_execute/sub_166/carry[21] ) );
  XNOR U22 ( .A(\u_a23_core/u_execute/pc[20] ), .B(
        \u_a23_core/u_execute/sub_166/carry[20] ), .Z(
        \u_a23_core/u_execute/pc_minus4[20] ) );
  OR U23 ( .A(\u_a23_core/u_execute/sub_166/carry[21] ), .B(
        \u_a23_core/u_execute/pc[21] ), .Z(
        \u_a23_core/u_execute/sub_166/carry[22] ) );
  XNOR U24 ( .A(\u_a23_core/u_execute/pc[21] ), .B(
        \u_a23_core/u_execute/sub_166/carry[21] ), .Z(
        \u_a23_core/u_execute/pc_minus4[21] ) );
  OR U25 ( .A(\u_a23_core/u_execute/sub_166/carry[22] ), .B(
        \u_a23_core/u_execute/pc[22] ), .Z(
        \u_a23_core/u_execute/sub_166/carry[23] ) );
  XNOR U26 ( .A(\u_a23_core/u_execute/pc[22] ), .B(
        \u_a23_core/u_execute/sub_166/carry[22] ), .Z(
        \u_a23_core/u_execute/pc_minus4[22] ) );
  OR U27 ( .A(\u_a23_core/u_execute/sub_166/carry[23] ), .B(
        \u_a23_core/u_execute/pc[23] ), .Z(
        \u_a23_core/u_execute/sub_166/carry[24] ) );
  XNOR U28 ( .A(\u_a23_core/u_execute/pc[23] ), .B(
        \u_a23_core/u_execute/sub_166/carry[23] ), .Z(
        \u_a23_core/u_execute/pc_minus4[23] ) );
  OR U29 ( .A(\u_a23_core/u_execute/sub_166/carry[24] ), .B(
        \u_a23_core/u_execute/pc[24] ), .Z(
        \u_a23_core/u_execute/sub_166/carry[25] ) );
  XNOR U30 ( .A(\u_a23_core/u_execute/pc[24] ), .B(
        \u_a23_core/u_execute/sub_166/carry[24] ), .Z(
        \u_a23_core/u_execute/pc_minus4[24] ) );
  OR U31 ( .A(\u_a23_core/u_execute/sub_166/carry[25] ), .B(
        \u_a23_core/u_execute/pc[25] ), .Z(
        \u_a23_core/u_execute/sub_166/carry[26] ) );
  XNOR U32 ( .A(\u_a23_core/u_execute/pc[25] ), .B(
        \u_a23_core/u_execute/sub_166/carry[25] ), .Z(
        \u_a23_core/u_execute/pc_minus4[25] ) );
  OR U33 ( .A(\u_a23_core/u_execute/pc[2] ), .B(\u_a23_core/u_execute/pc[3] ), 
        .Z(\u_a23_core/u_execute/sub_166/carry[4] ) );
  XNOR U34 ( .A(\u_a23_core/u_execute/pc[3] ), .B(\u_a23_core/u_execute/pc[2] ), .Z(\u_a23_core/u_execute/pc_minus4[3] ) );
  OR U35 ( .A(\u_a23_core/u_execute/sub_166/carry[4] ), .B(
        \u_a23_core/u_execute/pc[4] ), .Z(
        \u_a23_core/u_execute/sub_166/carry[5] ) );
  XNOR U36 ( .A(\u_a23_core/u_execute/pc[4] ), .B(
        \u_a23_core/u_execute/sub_166/carry[4] ), .Z(
        \u_a23_core/u_execute/pc_minus4[4] ) );
  OR U37 ( .A(\u_a23_core/u_execute/sub_166/carry[5] ), .B(
        \u_a23_core/u_execute/pc[5] ), .Z(
        \u_a23_core/u_execute/sub_166/carry[6] ) );
  XNOR U38 ( .A(\u_a23_core/u_execute/pc[5] ), .B(
        \u_a23_core/u_execute/sub_166/carry[5] ), .Z(
        \u_a23_core/u_execute/pc_minus4[5] ) );
  OR U39 ( .A(\u_a23_core/u_execute/sub_166/carry[6] ), .B(
        \u_a23_core/u_execute/pc[6] ), .Z(
        \u_a23_core/u_execute/sub_166/carry[7] ) );
  XNOR U40 ( .A(\u_a23_core/u_execute/pc[6] ), .B(
        \u_a23_core/u_execute/sub_166/carry[6] ), .Z(
        \u_a23_core/u_execute/pc_minus4[6] ) );
  OR U41 ( .A(\u_a23_core/u_execute/sub_166/carry[7] ), .B(
        \u_a23_core/u_execute/pc[7] ), .Z(
        \u_a23_core/u_execute/sub_166/carry[8] ) );
  XNOR U42 ( .A(\u_a23_core/u_execute/pc[7] ), .B(
        \u_a23_core/u_execute/sub_166/carry[7] ), .Z(
        \u_a23_core/u_execute/pc_minus4[7] ) );
  OR U43 ( .A(\u_a23_core/u_execute/sub_166/carry[8] ), .B(
        \u_a23_core/u_execute/pc[8] ), .Z(
        \u_a23_core/u_execute/sub_166/carry[9] ) );
  XNOR U44 ( .A(\u_a23_core/u_execute/pc[8] ), .B(
        \u_a23_core/u_execute/sub_166/carry[8] ), .Z(
        \u_a23_core/u_execute/pc_minus4[8] ) );
  OR U45 ( .A(\u_a23_core/u_execute/sub_166/carry[9] ), .B(
        \u_a23_core/u_execute/pc[9] ), .Z(
        \u_a23_core/u_execute/sub_166/carry[10] ) );
  XNOR U46 ( .A(\u_a23_core/u_execute/pc[9] ), .B(
        \u_a23_core/u_execute/sub_166/carry[9] ), .Z(
        \u_a23_core/u_execute/pc_minus4[9] ) );
  AND U47 ( .A(\u_a23_core/u_execute/u_multiply/product[34] ), .B(
        \u_a23_core/u_execute/u_multiply/sum34_b[0] ), .Z(
        \u_a23_core/u_execute/u_multiply/add_100/carry[1] ) );
  XOR U48 ( .A(\u_a23_core/u_execute/u_multiply/sum34_b[0] ), .B(
        \u_a23_core/u_execute/u_multiply/product[34] ), .Z(
        \u_a23_core/u_execute/u_multiply/sum[0] ) );
  AND U49 ( .A(\u_a23_core/u_execute/multiply_out[0] ), .B(
        \u_a23_core/u_execute/rs[0] ), .Z(
        \u_a23_core/u_execute/u_multiply/add_105/carry[1] ) );
  XOR U50 ( .A(\u_a23_core/u_execute/rs[0] ), .B(
        \u_a23_core/u_execute/multiply_out[0] ), .Z(
        \u_a23_core/u_execute/u_multiply/sum_acc1[0] ) );
  AND U51 ( .A(\u_a23_core/u_execute/pc[2] ), .B(\u_a23_core/u_execute/pc[3] ), 
        .Z(\u_a23_core/u_execute/add_165/carry[4] ) );
  XOR U52 ( .A(\u_a23_core/u_execute/pc[3] ), .B(\u_a23_core/u_execute/pc[2] ), 
        .Z(\u_a23_core/u_execute/pc_plus4[3] ) );
  AND U53 ( .A(\u_a23_core/u_execute/add_165/carry[4] ), .B(
        \u_a23_core/u_execute/pc[4] ), .Z(
        \u_a23_core/u_execute/add_165/carry[5] ) );
  XOR U54 ( .A(\u_a23_core/u_execute/pc[4] ), .B(
        \u_a23_core/u_execute/add_165/carry[4] ), .Z(
        \u_a23_core/u_execute/pc_plus4[4] ) );
  AND U55 ( .A(\u_a23_core/u_execute/add_165/carry[5] ), .B(
        \u_a23_core/u_execute/pc[5] ), .Z(
        \u_a23_core/u_execute/add_165/carry[6] ) );
  XOR U56 ( .A(\u_a23_core/u_execute/pc[5] ), .B(
        \u_a23_core/u_execute/add_165/carry[5] ), .Z(
        \u_a23_core/u_execute/pc_plus4[5] ) );
  AND U57 ( .A(\u_a23_core/u_execute/add_165/carry[6] ), .B(
        \u_a23_core/u_execute/pc[6] ), .Z(
        \u_a23_core/u_execute/add_165/carry[7] ) );
  XOR U58 ( .A(\u_a23_core/u_execute/pc[6] ), .B(
        \u_a23_core/u_execute/add_165/carry[6] ), .Z(
        \u_a23_core/u_execute/pc_plus4[6] ) );
  AND U59 ( .A(\u_a23_core/u_execute/add_165/carry[7] ), .B(
        \u_a23_core/u_execute/pc[7] ), .Z(
        \u_a23_core/u_execute/add_165/carry[8] ) );
  XOR U60 ( .A(\u_a23_core/u_execute/pc[7] ), .B(
        \u_a23_core/u_execute/add_165/carry[7] ), .Z(
        \u_a23_core/u_execute/pc_plus4[7] ) );
  AND U61 ( .A(\u_a23_core/u_execute/add_165/carry[8] ), .B(
        \u_a23_core/u_execute/pc[8] ), .Z(
        \u_a23_core/u_execute/add_165/carry[9] ) );
  XOR U62 ( .A(\u_a23_core/u_execute/pc[8] ), .B(
        \u_a23_core/u_execute/add_165/carry[8] ), .Z(
        \u_a23_core/u_execute/pc_plus4[8] ) );
  AND U63 ( .A(\u_a23_core/u_execute/add_165/carry[9] ), .B(
        \u_a23_core/u_execute/pc[9] ), .Z(
        \u_a23_core/u_execute/add_165/carry[10] ) );
  XOR U64 ( .A(\u_a23_core/u_execute/pc[9] ), .B(
        \u_a23_core/u_execute/add_165/carry[9] ), .Z(
        \u_a23_core/u_execute/pc_plus4[9] ) );
  AND U65 ( .A(\u_a23_core/u_execute/add_165/carry[10] ), .B(
        \u_a23_core/u_execute/pc[10] ), .Z(
        \u_a23_core/u_execute/add_165/carry[11] ) );
  XOR U66 ( .A(\u_a23_core/u_execute/pc[10] ), .B(
        \u_a23_core/u_execute/add_165/carry[10] ), .Z(
        \u_a23_core/u_execute/pc_plus4[10] ) );
  AND U67 ( .A(\u_a23_core/u_execute/add_165/carry[11] ), .B(
        \u_a23_core/u_execute/pc[11] ), .Z(
        \u_a23_core/u_execute/add_165/carry[12] ) );
  XOR U68 ( .A(\u_a23_core/u_execute/pc[11] ), .B(
        \u_a23_core/u_execute/add_165/carry[11] ), .Z(
        \u_a23_core/u_execute/pc_plus4[11] ) );
  AND U69 ( .A(\u_a23_core/u_execute/add_165/carry[12] ), .B(
        \u_a23_core/u_execute/pc[12] ), .Z(
        \u_a23_core/u_execute/add_165/carry[13] ) );
  XOR U70 ( .A(\u_a23_core/u_execute/pc[12] ), .B(
        \u_a23_core/u_execute/add_165/carry[12] ), .Z(
        \u_a23_core/u_execute/pc_plus4[12] ) );
  AND U71 ( .A(\u_a23_core/u_execute/add_165/carry[13] ), .B(
        \u_a23_core/u_execute/pc[13] ), .Z(
        \u_a23_core/u_execute/add_165/carry[14] ) );
  XOR U72 ( .A(\u_a23_core/u_execute/pc[13] ), .B(
        \u_a23_core/u_execute/add_165/carry[13] ), .Z(
        \u_a23_core/u_execute/pc_plus4[13] ) );
  AND U73 ( .A(\u_a23_core/u_execute/add_165/carry[14] ), .B(
        \u_a23_core/u_execute/pc[14] ), .Z(
        \u_a23_core/u_execute/add_165/carry[15] ) );
  XOR U74 ( .A(\u_a23_core/u_execute/pc[14] ), .B(
        \u_a23_core/u_execute/add_165/carry[14] ), .Z(
        \u_a23_core/u_execute/pc_plus4[14] ) );
  AND U75 ( .A(\u_a23_core/u_execute/add_165/carry[15] ), .B(
        \u_a23_core/u_execute/pc[15] ), .Z(
        \u_a23_core/u_execute/add_165/carry[16] ) );
  XOR U76 ( .A(\u_a23_core/u_execute/pc[15] ), .B(
        \u_a23_core/u_execute/add_165/carry[15] ), .Z(
        \u_a23_core/u_execute/pc_plus4[15] ) );
  AND U77 ( .A(\u_a23_core/u_execute/add_165/carry[16] ), .B(
        \u_a23_core/u_execute/pc[16] ), .Z(
        \u_a23_core/u_execute/add_165/carry[17] ) );
  XOR U78 ( .A(\u_a23_core/u_execute/pc[16] ), .B(
        \u_a23_core/u_execute/add_165/carry[16] ), .Z(
        \u_a23_core/u_execute/pc_plus4[16] ) );
  AND U79 ( .A(\u_a23_core/u_execute/add_165/carry[17] ), .B(
        \u_a23_core/u_execute/pc[17] ), .Z(
        \u_a23_core/u_execute/add_165/carry[18] ) );
  XOR U80 ( .A(\u_a23_core/u_execute/pc[17] ), .B(
        \u_a23_core/u_execute/add_165/carry[17] ), .Z(
        \u_a23_core/u_execute/pc_plus4[17] ) );
  AND U81 ( .A(\u_a23_core/u_execute/add_165/carry[18] ), .B(
        \u_a23_core/u_execute/pc[18] ), .Z(
        \u_a23_core/u_execute/add_165/carry[19] ) );
  XOR U82 ( .A(\u_a23_core/u_execute/pc[18] ), .B(
        \u_a23_core/u_execute/add_165/carry[18] ), .Z(
        \u_a23_core/u_execute/pc_plus4[18] ) );
  AND U83 ( .A(\u_a23_core/u_execute/add_165/carry[19] ), .B(
        \u_a23_core/u_execute/pc[19] ), .Z(
        \u_a23_core/u_execute/add_165/carry[20] ) );
  XOR U84 ( .A(\u_a23_core/u_execute/pc[19] ), .B(
        \u_a23_core/u_execute/add_165/carry[19] ), .Z(
        \u_a23_core/u_execute/pc_plus4[19] ) );
  AND U85 ( .A(\u_a23_core/u_execute/add_165/carry[20] ), .B(
        \u_a23_core/u_execute/pc[20] ), .Z(
        \u_a23_core/u_execute/add_165/carry[21] ) );
  XOR U86 ( .A(\u_a23_core/u_execute/pc[20] ), .B(
        \u_a23_core/u_execute/add_165/carry[20] ), .Z(
        \u_a23_core/u_execute/pc_plus4[20] ) );
  AND U87 ( .A(\u_a23_core/u_execute/add_165/carry[21] ), .B(
        \u_a23_core/u_execute/pc[21] ), .Z(
        \u_a23_core/u_execute/add_165/carry[22] ) );
  XOR U88 ( .A(\u_a23_core/u_execute/pc[21] ), .B(
        \u_a23_core/u_execute/add_165/carry[21] ), .Z(
        \u_a23_core/u_execute/pc_plus4[21] ) );
  AND U89 ( .A(\u_a23_core/u_execute/add_165/carry[22] ), .B(
        \u_a23_core/u_execute/pc[22] ), .Z(
        \u_a23_core/u_execute/add_165/carry[23] ) );
  XOR U90 ( .A(\u_a23_core/u_execute/pc[22] ), .B(
        \u_a23_core/u_execute/add_165/carry[22] ), .Z(
        \u_a23_core/u_execute/pc_plus4[22] ) );
  AND U91 ( .A(\u_a23_core/u_execute/add_165/carry[23] ), .B(
        \u_a23_core/u_execute/pc[23] ), .Z(
        \u_a23_core/u_execute/add_165/carry[24] ) );
  XOR U92 ( .A(\u_a23_core/u_execute/pc[23] ), .B(
        \u_a23_core/u_execute/add_165/carry[23] ), .Z(
        \u_a23_core/u_execute/pc_plus4[23] ) );
  AND U93 ( .A(\u_a23_core/u_execute/add_165/carry[24] ), .B(
        \u_a23_core/u_execute/pc[24] ), .Z(
        \u_a23_core/u_execute/add_165/carry[25] ) );
  XOR U94 ( .A(\u_a23_core/u_execute/pc[24] ), .B(
        \u_a23_core/u_execute/add_165/carry[24] ), .Z(
        \u_a23_core/u_execute/pc_plus4[24] ) );
  AND U95 ( .A(\u_a23_core/u_execute/pc[25] ), .B(
        \u_a23_core/u_execute/add_165/carry[25] ), .Z(
        \u_a23_core/u_execute/pc_plus4[26] ) );
  XOR U96 ( .A(\u_a23_core/u_execute/pc[25] ), .B(
        \u_a23_core/u_execute/add_165/carry[25] ), .Z(
        \u_a23_core/u_execute/pc_plus4[25] ) );
  AND U97 ( .A(m_address[2]), .B(m_address[3]), .Z(
        \u_a23_core/u_execute/add_167/carry[4] ) );
  XOR U98 ( .A(m_address[3]), .B(m_address[2]), .Z(
        \u_a23_core/u_execute/address_plus4[3] ) );
  AND U99 ( .A(\u_a23_core/u_execute/add_167/carry[4] ), .B(m_address[4]), .Z(
        \u_a23_core/u_execute/add_167/carry[5] ) );
  XOR U100 ( .A(m_address[4]), .B(\u_a23_core/u_execute/add_167/carry[4] ), 
        .Z(\u_a23_core/u_execute/address_plus4[4] ) );
  AND U101 ( .A(\u_a23_core/u_execute/add_167/carry[5] ), .B(m_address[5]), 
        .Z(\u_a23_core/u_execute/add_167/carry[6] ) );
  XOR U102 ( .A(m_address[5]), .B(\u_a23_core/u_execute/add_167/carry[5] ), 
        .Z(\u_a23_core/u_execute/address_plus4[5] ) );
  AND U103 ( .A(\u_a23_core/u_execute/add_167/carry[6] ), .B(m_address[6]), 
        .Z(\u_a23_core/u_execute/add_167/carry[7] ) );
  XOR U104 ( .A(m_address[6]), .B(\u_a23_core/u_execute/add_167/carry[6] ), 
        .Z(\u_a23_core/u_execute/address_plus4[6] ) );
  AND U105 ( .A(\u_a23_core/u_execute/add_167/carry[7] ), .B(m_address[7]), 
        .Z(\u_a23_core/u_execute/add_167/carry[8] ) );
  XOR U106 ( .A(m_address[7]), .B(\u_a23_core/u_execute/add_167/carry[7] ), 
        .Z(\u_a23_core/u_execute/address_plus4[7] ) );
  AND U107 ( .A(\u_a23_core/u_execute/add_167/carry[8] ), .B(m_address[8]), 
        .Z(\u_a23_core/u_execute/add_167/carry[9] ) );
  XOR U108 ( .A(m_address[8]), .B(\u_a23_core/u_execute/add_167/carry[8] ), 
        .Z(\u_a23_core/u_execute/address_plus4[8] ) );
  AND U109 ( .A(\u_a23_core/u_execute/add_167/carry[9] ), .B(m_address[9]), 
        .Z(\u_a23_core/u_execute/add_167/carry[10] ) );
  XOR U110 ( .A(m_address[9]), .B(\u_a23_core/u_execute/add_167/carry[9] ), 
        .Z(\u_a23_core/u_execute/address_plus4[9] ) );
  AND U111 ( .A(\u_a23_core/u_execute/add_167/carry[10] ), .B(m_address[10]), 
        .Z(\u_a23_core/u_execute/add_167/carry[11] ) );
  XOR U112 ( .A(m_address[10]), .B(\u_a23_core/u_execute/add_167/carry[10] ), 
        .Z(\u_a23_core/u_execute/address_plus4[10] ) );
  AND U113 ( .A(\u_a23_core/u_execute/add_167/carry[11] ), .B(m_address[11]), 
        .Z(\u_a23_core/u_execute/add_167/carry[12] ) );
  XOR U114 ( .A(m_address[11]), .B(\u_a23_core/u_execute/add_167/carry[11] ), 
        .Z(\u_a23_core/u_execute/address_plus4[11] ) );
  AND U115 ( .A(\u_a23_core/u_execute/add_167/carry[12] ), .B(m_address[12]), 
        .Z(\u_a23_core/u_execute/add_167/carry[13] ) );
  XOR U116 ( .A(m_address[12]), .B(\u_a23_core/u_execute/add_167/carry[12] ), 
        .Z(\u_a23_core/u_execute/address_plus4[12] ) );
  AND U117 ( .A(\u_a23_core/u_execute/add_167/carry[13] ), .B(m_address[13]), 
        .Z(\u_a23_core/u_execute/add_167/carry[14] ) );
  XOR U118 ( .A(m_address[13]), .B(\u_a23_core/u_execute/add_167/carry[13] ), 
        .Z(\u_a23_core/u_execute/address_plus4[13] ) );
  AND U119 ( .A(\u_a23_core/u_execute/add_167/carry[14] ), .B(m_address[14]), 
        .Z(\u_a23_core/u_execute/add_167/carry[15] ) );
  XOR U120 ( .A(m_address[14]), .B(\u_a23_core/u_execute/add_167/carry[14] ), 
        .Z(\u_a23_core/u_execute/address_plus4[14] ) );
  AND U121 ( .A(\u_a23_core/u_execute/add_167/carry[15] ), .B(m_address[15]), 
        .Z(\u_a23_core/u_execute/add_167/carry[16] ) );
  XOR U122 ( .A(m_address[15]), .B(\u_a23_core/u_execute/add_167/carry[15] ), 
        .Z(\u_a23_core/u_execute/address_plus4[15] ) );
  AND U123 ( .A(\u_a23_core/u_execute/add_167/carry[16] ), .B(m_address[16]), 
        .Z(\u_a23_core/u_execute/add_167/carry[17] ) );
  XOR U124 ( .A(m_address[16]), .B(\u_a23_core/u_execute/add_167/carry[16] ), 
        .Z(\u_a23_core/u_execute/address_plus4[16] ) );
  AND U125 ( .A(\u_a23_core/u_execute/add_167/carry[17] ), .B(m_address[17]), 
        .Z(\u_a23_core/u_execute/add_167/carry[18] ) );
  XOR U126 ( .A(m_address[17]), .B(\u_a23_core/u_execute/add_167/carry[17] ), 
        .Z(\u_a23_core/u_execute/address_plus4[17] ) );
  AND U127 ( .A(\u_a23_core/u_execute/add_167/carry[18] ), .B(m_address[18]), 
        .Z(\u_a23_core/u_execute/add_167/carry[19] ) );
  XOR U128 ( .A(m_address[18]), .B(\u_a23_core/u_execute/add_167/carry[18] ), 
        .Z(\u_a23_core/u_execute/address_plus4[18] ) );
  AND U129 ( .A(\u_a23_core/u_execute/add_167/carry[19] ), .B(m_address[19]), 
        .Z(\u_a23_core/u_execute/add_167/carry[20] ) );
  XOR U130 ( .A(m_address[19]), .B(\u_a23_core/u_execute/add_167/carry[19] ), 
        .Z(\u_a23_core/u_execute/address_plus4[19] ) );
  AND U131 ( .A(\u_a23_core/u_execute/add_167/carry[20] ), .B(m_address[20]), 
        .Z(\u_a23_core/u_execute/add_167/carry[21] ) );
  XOR U132 ( .A(m_address[20]), .B(\u_a23_core/u_execute/add_167/carry[20] ), 
        .Z(\u_a23_core/u_execute/address_plus4[20] ) );
  AND U133 ( .A(\u_a23_core/u_execute/add_167/carry[21] ), .B(m_address[21]), 
        .Z(\u_a23_core/u_execute/add_167/carry[22] ) );
  XOR U134 ( .A(m_address[21]), .B(\u_a23_core/u_execute/add_167/carry[21] ), 
        .Z(\u_a23_core/u_execute/address_plus4[21] ) );
  AND U135 ( .A(\u_a23_core/u_execute/add_167/carry[22] ), .B(m_address[22]), 
        .Z(\u_a23_core/u_execute/add_167/carry[23] ) );
  XOR U136 ( .A(m_address[22]), .B(\u_a23_core/u_execute/add_167/carry[22] ), 
        .Z(\u_a23_core/u_execute/address_plus4[22] ) );
  AND U137 ( .A(\u_a23_core/u_execute/add_167/carry[23] ), .B(m_address[23]), 
        .Z(\u_a23_core/u_execute/add_167/carry[24] ) );
  XOR U138 ( .A(m_address[23]), .B(\u_a23_core/u_execute/add_167/carry[23] ), 
        .Z(\u_a23_core/u_execute/address_plus4[23] ) );
  AND U139 ( .A(\u_a23_core/u_execute/add_167/carry[24] ), .B(m_address[24]), 
        .Z(\u_a23_core/u_execute/add_167/carry[25] ) );
  XOR U140 ( .A(m_address[24]), .B(\u_a23_core/u_execute/add_167/carry[24] ), 
        .Z(\u_a23_core/u_execute/address_plus4[24] ) );
  AND U141 ( .A(\u_a23_core/u_execute/add_167/carry[25] ), .B(m_address[25]), 
        .Z(\u_a23_core/u_execute/add_167/carry[26] ) );
  XOR U142 ( .A(m_address[25]), .B(\u_a23_core/u_execute/add_167/carry[25] ), 
        .Z(\u_a23_core/u_execute/address_plus4[25] ) );
  AND U143 ( .A(\u_a23_core/u_execute/add_167/carry[26] ), .B(m_address[26]), 
        .Z(\u_a23_core/u_execute/add_167/carry[27] ) );
  XOR U144 ( .A(m_address[26]), .B(\u_a23_core/u_execute/add_167/carry[26] ), 
        .Z(\u_a23_core/u_execute/address_plus4[26] ) );
  AND U145 ( .A(\u_a23_core/u_execute/add_167/carry[27] ), .B(m_address[27]), 
        .Z(\u_a23_core/u_execute/add_167/carry[28] ) );
  XOR U146 ( .A(m_address[27]), .B(\u_a23_core/u_execute/add_167/carry[27] ), 
        .Z(\u_a23_core/u_execute/address_plus4[27] ) );
  AND U147 ( .A(\u_a23_core/u_execute/add_167/carry[28] ), .B(m_address[28]), 
        .Z(\u_a23_core/u_execute/add_167/carry[29] ) );
  XOR U148 ( .A(m_address[28]), .B(\u_a23_core/u_execute/add_167/carry[28] ), 
        .Z(\u_a23_core/u_execute/address_plus4[28] ) );
  AND U149 ( .A(\u_a23_core/u_execute/add_167/carry[29] ), .B(m_address[29]), 
        .Z(\u_a23_core/u_execute/add_167/carry[30] ) );
  XOR U150 ( .A(m_address[29]), .B(\u_a23_core/u_execute/add_167/carry[29] ), 
        .Z(\u_a23_core/u_execute/address_plus4[29] ) );
  AND U151 ( .A(\u_a23_core/u_execute/add_167/carry[30] ), .B(m_address[30]), 
        .Z(\u_a23_core/u_execute/add_167/carry[31] ) );
  XOR U152 ( .A(m_address[30]), .B(\u_a23_core/u_execute/add_167/carry[30] ), 
        .Z(\u_a23_core/u_execute/address_plus4[30] ) );
  XOR U153 ( .A(m_address[31]), .B(\u_a23_core/u_execute/add_167/carry[31] ), 
        .Z(\u_a23_core/u_execute/address_plus4[31] ) );
  AND U154 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[2] ), .B(
        \u_a23_core/u_execute/alu_out_pc_filtered[3] ), .Z(
        \u_a23_core/u_execute/add_168/carry[4] ) );
  XOR U155 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[3] ), .B(
        \u_a23_core/u_execute/alu_out_pc_filtered[2] ), .Z(
        \u_a23_core/u_execute/alu_plus4[3] ) );
  AND U156 ( .A(\u_a23_core/u_execute/add_168/carry[4] ), .B(
        \u_a23_core/u_execute/alu_out_pc_filtered[4] ), .Z(
        \u_a23_core/u_execute/add_168/carry[5] ) );
  XOR U157 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[4] ), .B(
        \u_a23_core/u_execute/add_168/carry[4] ), .Z(
        \u_a23_core/u_execute/alu_plus4[4] ) );
  AND U158 ( .A(\u_a23_core/u_execute/add_168/carry[5] ), .B(
        \u_a23_core/u_execute/alu_out_pc_filtered[5] ), .Z(
        \u_a23_core/u_execute/add_168/carry[6] ) );
  XOR U159 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[5] ), .B(
        \u_a23_core/u_execute/add_168/carry[5] ), .Z(
        \u_a23_core/u_execute/alu_plus4[5] ) );
  AND U160 ( .A(\u_a23_core/u_execute/add_168/carry[6] ), .B(
        \u_a23_core/u_execute/alu_out_pc_filtered[6] ), .Z(
        \u_a23_core/u_execute/add_168/carry[7] ) );
  XOR U161 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[6] ), .B(
        \u_a23_core/u_execute/add_168/carry[6] ), .Z(
        \u_a23_core/u_execute/alu_plus4[6] ) );
  AND U162 ( .A(\u_a23_core/u_execute/add_168/carry[7] ), .B(
        \u_a23_core/u_execute/alu_out_pc_filtered[7] ), .Z(
        \u_a23_core/u_execute/add_168/carry[8] ) );
  XOR U163 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[7] ), .B(
        \u_a23_core/u_execute/add_168/carry[7] ), .Z(
        \u_a23_core/u_execute/alu_plus4[7] ) );
  AND U164 ( .A(\u_a23_core/u_execute/add_168/carry[8] ), .B(
        \u_a23_core/u_execute/alu_out_pc_filtered[8] ), .Z(
        \u_a23_core/u_execute/add_168/carry[9] ) );
  XOR U165 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[8] ), .B(
        \u_a23_core/u_execute/add_168/carry[8] ), .Z(
        \u_a23_core/u_execute/alu_plus4[8] ) );
  AND U166 ( .A(\u_a23_core/u_execute/add_168/carry[9] ), .B(
        \u_a23_core/u_execute/alu_out_pc_filtered[9] ), .Z(
        \u_a23_core/u_execute/add_168/carry[10] ) );
  XOR U167 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[9] ), .B(
        \u_a23_core/u_execute/add_168/carry[9] ), .Z(
        \u_a23_core/u_execute/alu_plus4[9] ) );
  AND U168 ( .A(\u_a23_core/u_execute/add_168/carry[10] ), .B(
        \u_a23_core/u_execute/alu_out_pc_filtered[10] ), .Z(
        \u_a23_core/u_execute/add_168/carry[11] ) );
  XOR U169 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[10] ), .B(
        \u_a23_core/u_execute/add_168/carry[10] ), .Z(
        \u_a23_core/u_execute/alu_plus4[10] ) );
  AND U170 ( .A(\u_a23_core/u_execute/add_168/carry[11] ), .B(
        \u_a23_core/u_execute/alu_out_pc_filtered[11] ), .Z(
        \u_a23_core/u_execute/add_168/carry[12] ) );
  XOR U171 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[11] ), .B(
        \u_a23_core/u_execute/add_168/carry[11] ), .Z(
        \u_a23_core/u_execute/alu_plus4[11] ) );
  AND U172 ( .A(\u_a23_core/u_execute/add_168/carry[12] ), .B(
        \u_a23_core/u_execute/alu_out_pc_filtered[12] ), .Z(
        \u_a23_core/u_execute/add_168/carry[13] ) );
  XOR U173 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[12] ), .B(
        \u_a23_core/u_execute/add_168/carry[12] ), .Z(
        \u_a23_core/u_execute/alu_plus4[12] ) );
  AND U174 ( .A(\u_a23_core/u_execute/add_168/carry[13] ), .B(
        \u_a23_core/u_execute/alu_out_pc_filtered[13] ), .Z(
        \u_a23_core/u_execute/add_168/carry[14] ) );
  XOR U175 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[13] ), .B(
        \u_a23_core/u_execute/add_168/carry[13] ), .Z(
        \u_a23_core/u_execute/alu_plus4[13] ) );
  AND U176 ( .A(\u_a23_core/u_execute/add_168/carry[14] ), .B(
        \u_a23_core/u_execute/alu_out_pc_filtered[14] ), .Z(
        \u_a23_core/u_execute/add_168/carry[15] ) );
  XOR U177 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[14] ), .B(
        \u_a23_core/u_execute/add_168/carry[14] ), .Z(
        \u_a23_core/u_execute/alu_plus4[14] ) );
  AND U178 ( .A(\u_a23_core/u_execute/add_168/carry[15] ), .B(
        \u_a23_core/u_execute/alu_out_pc_filtered[15] ), .Z(
        \u_a23_core/u_execute/add_168/carry[16] ) );
  XOR U179 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[15] ), .B(
        \u_a23_core/u_execute/add_168/carry[15] ), .Z(
        \u_a23_core/u_execute/alu_plus4[15] ) );
  AND U180 ( .A(\u_a23_core/u_execute/add_168/carry[16] ), .B(
        \u_a23_core/u_execute/alu_out_pc_filtered[16] ), .Z(
        \u_a23_core/u_execute/add_168/carry[17] ) );
  XOR U181 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[16] ), .B(
        \u_a23_core/u_execute/add_168/carry[16] ), .Z(
        \u_a23_core/u_execute/alu_plus4[16] ) );
  AND U182 ( .A(\u_a23_core/u_execute/add_168/carry[17] ), .B(
        \u_a23_core/u_execute/alu_out_pc_filtered[17] ), .Z(
        \u_a23_core/u_execute/add_168/carry[18] ) );
  XOR U183 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[17] ), .B(
        \u_a23_core/u_execute/add_168/carry[17] ), .Z(
        \u_a23_core/u_execute/alu_plus4[17] ) );
  AND U184 ( .A(\u_a23_core/u_execute/add_168/carry[18] ), .B(
        \u_a23_core/u_execute/alu_out_pc_filtered[18] ), .Z(
        \u_a23_core/u_execute/add_168/carry[19] ) );
  XOR U185 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[18] ), .B(
        \u_a23_core/u_execute/add_168/carry[18] ), .Z(
        \u_a23_core/u_execute/alu_plus4[18] ) );
  AND U186 ( .A(\u_a23_core/u_execute/add_168/carry[19] ), .B(
        \u_a23_core/u_execute/alu_out_pc_filtered[19] ), .Z(
        \u_a23_core/u_execute/add_168/carry[20] ) );
  XOR U187 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[19] ), .B(
        \u_a23_core/u_execute/add_168/carry[19] ), .Z(
        \u_a23_core/u_execute/alu_plus4[19] ) );
  AND U188 ( .A(\u_a23_core/u_execute/add_168/carry[20] ), .B(
        \u_a23_core/u_execute/alu_out_pc_filtered[20] ), .Z(
        \u_a23_core/u_execute/add_168/carry[21] ) );
  XOR U189 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[20] ), .B(
        \u_a23_core/u_execute/add_168/carry[20] ), .Z(
        \u_a23_core/u_execute/alu_plus4[20] ) );
  AND U190 ( .A(\u_a23_core/u_execute/add_168/carry[21] ), .B(
        \u_a23_core/u_execute/alu_out_pc_filtered[21] ), .Z(
        \u_a23_core/u_execute/add_168/carry[22] ) );
  XOR U191 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[21] ), .B(
        \u_a23_core/u_execute/add_168/carry[21] ), .Z(
        \u_a23_core/u_execute/alu_plus4[21] ) );
  AND U192 ( .A(\u_a23_core/u_execute/add_168/carry[22] ), .B(
        \u_a23_core/u_execute/alu_out_pc_filtered[22] ), .Z(
        \u_a23_core/u_execute/add_168/carry[23] ) );
  XOR U193 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[22] ), .B(
        \u_a23_core/u_execute/add_168/carry[22] ), .Z(
        \u_a23_core/u_execute/alu_plus4[22] ) );
  AND U194 ( .A(\u_a23_core/u_execute/add_168/carry[23] ), .B(
        \u_a23_core/u_execute/alu_out_pc_filtered[23] ), .Z(
        \u_a23_core/u_execute/add_168/carry[24] ) );
  XOR U195 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[23] ), .B(
        \u_a23_core/u_execute/add_168/carry[23] ), .Z(
        \u_a23_core/u_execute/alu_plus4[23] ) );
  AND U196 ( .A(\u_a23_core/u_execute/add_168/carry[24] ), .B(
        \u_a23_core/u_execute/alu_out_pc_filtered[24] ), .Z(
        \u_a23_core/u_execute/add_168/carry[25] ) );
  XOR U197 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[24] ), .B(
        \u_a23_core/u_execute/add_168/carry[24] ), .Z(
        \u_a23_core/u_execute/alu_plus4[24] ) );
  AND U198 ( .A(\u_a23_core/u_execute/add_168/carry[25] ), .B(
        \u_a23_core/u_execute/alu_out_pc_filtered[25] ), .Z(
        \u_a23_core/u_execute/add_168/carry[26] ) );
  XOR U199 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[25] ), .B(
        \u_a23_core/u_execute/add_168/carry[25] ), .Z(
        \u_a23_core/u_execute/alu_plus4[25] ) );
  AND U200 ( .A(\u_a23_core/u_execute/add_168/carry[26] ), .B(
        \u_a23_core/u_execute/alu_out[26] ), .Z(
        \u_a23_core/u_execute/add_168/carry[27] ) );
  XOR U201 ( .A(\u_a23_core/u_execute/alu_out[26] ), .B(
        \u_a23_core/u_execute/add_168/carry[26] ), .Z(
        \u_a23_core/u_execute/alu_plus4[26] ) );
  AND U202 ( .A(\u_a23_core/u_execute/add_168/carry[27] ), .B(
        \u_a23_core/u_execute/alu_out[27] ), .Z(
        \u_a23_core/u_execute/add_168/carry[28] ) );
  XOR U203 ( .A(\u_a23_core/u_execute/alu_out[27] ), .B(
        \u_a23_core/u_execute/add_168/carry[27] ), .Z(
        \u_a23_core/u_execute/alu_plus4[27] ) );
  AND U204 ( .A(\u_a23_core/u_execute/add_168/carry[28] ), .B(
        \u_a23_core/u_execute/alu_out[28] ), .Z(
        \u_a23_core/u_execute/add_168/carry[29] ) );
  XOR U205 ( .A(\u_a23_core/u_execute/alu_out[28] ), .B(
        \u_a23_core/u_execute/add_168/carry[28] ), .Z(
        \u_a23_core/u_execute/alu_plus4[28] ) );
  AND U206 ( .A(\u_a23_core/u_execute/add_168/carry[29] ), .B(
        \u_a23_core/u_execute/alu_out[29] ), .Z(
        \u_a23_core/u_execute/add_168/carry[30] ) );
  XOR U207 ( .A(\u_a23_core/u_execute/alu_out[29] ), .B(
        \u_a23_core/u_execute/add_168/carry[29] ), .Z(
        \u_a23_core/u_execute/alu_plus4[29] ) );
  AND U208 ( .A(\u_a23_core/u_execute/add_168/carry[30] ), .B(
        \u_a23_core/u_execute/alu_out[30] ), .Z(
        \u_a23_core/u_execute/add_168/carry[31] ) );
  XOR U209 ( .A(\u_a23_core/u_execute/alu_out[30] ), .B(
        \u_a23_core/u_execute/add_168/carry[30] ), .Z(
        \u_a23_core/u_execute/alu_plus4[30] ) );
  XOR U210 ( .A(\u_a23_core/u_execute/alu_out[31] ), .B(
        \u_a23_core/u_execute/add_168/carry[31] ), .Z(
        \u_a23_core/u_execute/alu_plus4[31] ) );
  AND U211 ( .A(\u_a23_core/u_execute/rn[2] ), .B(\u_a23_core/u_execute/rn[3] ), .Z(\u_a23_core/u_execute/add_169/carry[4] ) );
  XOR U212 ( .A(\u_a23_core/u_execute/rn[3] ), .B(\u_a23_core/u_execute/rn[2] ), .Z(\u_a23_core/u_execute/rn_plus4[3] ) );
  AND U213 ( .A(\u_a23_core/u_execute/add_169/carry[4] ), .B(
        \u_a23_core/u_execute/rn[4] ), .Z(
        \u_a23_core/u_execute/add_169/carry[5] ) );
  XOR U214 ( .A(\u_a23_core/u_execute/rn[4] ), .B(
        \u_a23_core/u_execute/add_169/carry[4] ), .Z(
        \u_a23_core/u_execute/rn_plus4[4] ) );
  AND U215 ( .A(\u_a23_core/u_execute/add_169/carry[5] ), .B(
        \u_a23_core/u_execute/rn[5] ), .Z(
        \u_a23_core/u_execute/add_169/carry[6] ) );
  XOR U216 ( .A(\u_a23_core/u_execute/rn[5] ), .B(
        \u_a23_core/u_execute/add_169/carry[5] ), .Z(
        \u_a23_core/u_execute/rn_plus4[5] ) );
  AND U217 ( .A(\u_a23_core/u_execute/add_169/carry[6] ), .B(
        \u_a23_core/u_execute/rn[6] ), .Z(
        \u_a23_core/u_execute/add_169/carry[7] ) );
  XOR U218 ( .A(\u_a23_core/u_execute/rn[6] ), .B(
        \u_a23_core/u_execute/add_169/carry[6] ), .Z(
        \u_a23_core/u_execute/rn_plus4[6] ) );
  AND U219 ( .A(\u_a23_core/u_execute/add_169/carry[7] ), .B(
        \u_a23_core/u_execute/rn[7] ), .Z(
        \u_a23_core/u_execute/add_169/carry[8] ) );
  XOR U220 ( .A(\u_a23_core/u_execute/rn[7] ), .B(
        \u_a23_core/u_execute/add_169/carry[7] ), .Z(
        \u_a23_core/u_execute/rn_plus4[7] ) );
  AND U221 ( .A(\u_a23_core/u_execute/add_169/carry[8] ), .B(
        \u_a23_core/u_execute/rn[8] ), .Z(
        \u_a23_core/u_execute/add_169/carry[9] ) );
  XOR U222 ( .A(\u_a23_core/u_execute/rn[8] ), .B(
        \u_a23_core/u_execute/add_169/carry[8] ), .Z(
        \u_a23_core/u_execute/rn_plus4[8] ) );
  AND U223 ( .A(\u_a23_core/u_execute/add_169/carry[9] ), .B(
        \u_a23_core/u_execute/rn[9] ), .Z(
        \u_a23_core/u_execute/add_169/carry[10] ) );
  XOR U224 ( .A(\u_a23_core/u_execute/rn[9] ), .B(
        \u_a23_core/u_execute/add_169/carry[9] ), .Z(
        \u_a23_core/u_execute/rn_plus4[9] ) );
  AND U225 ( .A(\u_a23_core/u_execute/add_169/carry[10] ), .B(
        \u_a23_core/u_execute/rn[10] ), .Z(
        \u_a23_core/u_execute/add_169/carry[11] ) );
  XOR U226 ( .A(\u_a23_core/u_execute/rn[10] ), .B(
        \u_a23_core/u_execute/add_169/carry[10] ), .Z(
        \u_a23_core/u_execute/rn_plus4[10] ) );
  AND U227 ( .A(\u_a23_core/u_execute/add_169/carry[11] ), .B(
        \u_a23_core/u_execute/rn[11] ), .Z(
        \u_a23_core/u_execute/add_169/carry[12] ) );
  XOR U228 ( .A(\u_a23_core/u_execute/rn[11] ), .B(
        \u_a23_core/u_execute/add_169/carry[11] ), .Z(
        \u_a23_core/u_execute/rn_plus4[11] ) );
  AND U229 ( .A(\u_a23_core/u_execute/add_169/carry[12] ), .B(
        \u_a23_core/u_execute/rn[12] ), .Z(
        \u_a23_core/u_execute/add_169/carry[13] ) );
  XOR U230 ( .A(\u_a23_core/u_execute/rn[12] ), .B(
        \u_a23_core/u_execute/add_169/carry[12] ), .Z(
        \u_a23_core/u_execute/rn_plus4[12] ) );
  AND U231 ( .A(\u_a23_core/u_execute/add_169/carry[13] ), .B(
        \u_a23_core/u_execute/rn[13] ), .Z(
        \u_a23_core/u_execute/add_169/carry[14] ) );
  XOR U232 ( .A(\u_a23_core/u_execute/rn[13] ), .B(
        \u_a23_core/u_execute/add_169/carry[13] ), .Z(
        \u_a23_core/u_execute/rn_plus4[13] ) );
  AND U233 ( .A(\u_a23_core/u_execute/add_169/carry[14] ), .B(
        \u_a23_core/u_execute/rn[14] ), .Z(
        \u_a23_core/u_execute/add_169/carry[15] ) );
  XOR U234 ( .A(\u_a23_core/u_execute/rn[14] ), .B(
        \u_a23_core/u_execute/add_169/carry[14] ), .Z(
        \u_a23_core/u_execute/rn_plus4[14] ) );
  AND U235 ( .A(\u_a23_core/u_execute/add_169/carry[15] ), .B(
        \u_a23_core/u_execute/rn[15] ), .Z(
        \u_a23_core/u_execute/add_169/carry[16] ) );
  XOR U236 ( .A(\u_a23_core/u_execute/rn[15] ), .B(
        \u_a23_core/u_execute/add_169/carry[15] ), .Z(
        \u_a23_core/u_execute/rn_plus4[15] ) );
  AND U237 ( .A(\u_a23_core/u_execute/add_169/carry[16] ), .B(
        \u_a23_core/u_execute/rn[16] ), .Z(
        \u_a23_core/u_execute/add_169/carry[17] ) );
  XOR U238 ( .A(\u_a23_core/u_execute/rn[16] ), .B(
        \u_a23_core/u_execute/add_169/carry[16] ), .Z(
        \u_a23_core/u_execute/rn_plus4[16] ) );
  AND U239 ( .A(\u_a23_core/u_execute/add_169/carry[17] ), .B(
        \u_a23_core/u_execute/rn[17] ), .Z(
        \u_a23_core/u_execute/add_169/carry[18] ) );
  XOR U240 ( .A(\u_a23_core/u_execute/rn[17] ), .B(
        \u_a23_core/u_execute/add_169/carry[17] ), .Z(
        \u_a23_core/u_execute/rn_plus4[17] ) );
  AND U241 ( .A(\u_a23_core/u_execute/add_169/carry[18] ), .B(
        \u_a23_core/u_execute/rn[18] ), .Z(
        \u_a23_core/u_execute/add_169/carry[19] ) );
  XOR U242 ( .A(\u_a23_core/u_execute/rn[18] ), .B(
        \u_a23_core/u_execute/add_169/carry[18] ), .Z(
        \u_a23_core/u_execute/rn_plus4[18] ) );
  AND U243 ( .A(\u_a23_core/u_execute/add_169/carry[19] ), .B(
        \u_a23_core/u_execute/rn[19] ), .Z(
        \u_a23_core/u_execute/add_169/carry[20] ) );
  XOR U244 ( .A(\u_a23_core/u_execute/rn[19] ), .B(
        \u_a23_core/u_execute/add_169/carry[19] ), .Z(
        \u_a23_core/u_execute/rn_plus4[19] ) );
  AND U245 ( .A(\u_a23_core/u_execute/add_169/carry[20] ), .B(
        \u_a23_core/u_execute/rn[20] ), .Z(
        \u_a23_core/u_execute/add_169/carry[21] ) );
  XOR U246 ( .A(\u_a23_core/u_execute/rn[20] ), .B(
        \u_a23_core/u_execute/add_169/carry[20] ), .Z(
        \u_a23_core/u_execute/rn_plus4[20] ) );
  AND U247 ( .A(\u_a23_core/u_execute/add_169/carry[21] ), .B(
        \u_a23_core/u_execute/rn[21] ), .Z(
        \u_a23_core/u_execute/add_169/carry[22] ) );
  XOR U248 ( .A(\u_a23_core/u_execute/rn[21] ), .B(
        \u_a23_core/u_execute/add_169/carry[21] ), .Z(
        \u_a23_core/u_execute/rn_plus4[21] ) );
  AND U249 ( .A(\u_a23_core/u_execute/add_169/carry[22] ), .B(
        \u_a23_core/u_execute/rn[22] ), .Z(
        \u_a23_core/u_execute/add_169/carry[23] ) );
  XOR U250 ( .A(\u_a23_core/u_execute/rn[22] ), .B(
        \u_a23_core/u_execute/add_169/carry[22] ), .Z(
        \u_a23_core/u_execute/rn_plus4[22] ) );
  AND U251 ( .A(\u_a23_core/u_execute/add_169/carry[23] ), .B(
        \u_a23_core/u_execute/rn[23] ), .Z(
        \u_a23_core/u_execute/add_169/carry[24] ) );
  XOR U252 ( .A(\u_a23_core/u_execute/rn[23] ), .B(
        \u_a23_core/u_execute/add_169/carry[23] ), .Z(
        \u_a23_core/u_execute/rn_plus4[23] ) );
  AND U253 ( .A(\u_a23_core/u_execute/add_169/carry[24] ), .B(
        \u_a23_core/u_execute/rn[24] ), .Z(
        \u_a23_core/u_execute/add_169/carry[25] ) );
  XOR U254 ( .A(\u_a23_core/u_execute/rn[24] ), .B(
        \u_a23_core/u_execute/add_169/carry[24] ), .Z(
        \u_a23_core/u_execute/rn_plus4[24] ) );
  AND U255 ( .A(\u_a23_core/u_execute/add_169/carry[25] ), .B(
        \u_a23_core/u_execute/rn[25] ), .Z(
        \u_a23_core/u_execute/add_169/carry[26] ) );
  XOR U256 ( .A(\u_a23_core/u_execute/rn[25] ), .B(
        \u_a23_core/u_execute/add_169/carry[25] ), .Z(
        \u_a23_core/u_execute/rn_plus4[25] ) );
  AND U257 ( .A(\u_a23_core/u_execute/add_169/carry[26] ), .B(
        \u_a23_core/u_execute/rn[26] ), .Z(
        \u_a23_core/u_execute/add_169/carry[27] ) );
  XOR U258 ( .A(\u_a23_core/u_execute/rn[26] ), .B(
        \u_a23_core/u_execute/add_169/carry[26] ), .Z(
        \u_a23_core/u_execute/rn_plus4[26] ) );
  AND U259 ( .A(\u_a23_core/u_execute/add_169/carry[27] ), .B(
        \u_a23_core/u_execute/rn[27] ), .Z(
        \u_a23_core/u_execute/add_169/carry[28] ) );
  XOR U260 ( .A(\u_a23_core/u_execute/rn[27] ), .B(
        \u_a23_core/u_execute/add_169/carry[27] ), .Z(
        \u_a23_core/u_execute/rn_plus4[27] ) );
  AND U261 ( .A(\u_a23_core/u_execute/add_169/carry[28] ), .B(
        \u_a23_core/u_execute/rn[28] ), .Z(
        \u_a23_core/u_execute/add_169/carry[29] ) );
  XOR U262 ( .A(\u_a23_core/u_execute/rn[28] ), .B(
        \u_a23_core/u_execute/add_169/carry[28] ), .Z(
        \u_a23_core/u_execute/rn_plus4[28] ) );
  AND U263 ( .A(\u_a23_core/u_execute/add_169/carry[29] ), .B(
        \u_a23_core/u_execute/rn[29] ), .Z(
        \u_a23_core/u_execute/add_169/carry[30] ) );
  XOR U264 ( .A(\u_a23_core/u_execute/rn[29] ), .B(
        \u_a23_core/u_execute/add_169/carry[29] ), .Z(
        \u_a23_core/u_execute/rn_plus4[29] ) );
  AND U265 ( .A(\u_a23_core/u_execute/add_169/carry[30] ), .B(
        \u_a23_core/u_execute/rn[30] ), .Z(
        \u_a23_core/u_execute/add_169/carry[31] ) );
  XOR U266 ( .A(\u_a23_core/u_execute/rn[30] ), .B(
        \u_a23_core/u_execute/add_169/carry[30] ), .Z(
        \u_a23_core/u_execute/rn_plus4[30] ) );
  XOR U267 ( .A(\u_a23_core/u_execute/rn[31] ), .B(
        \u_a23_core/u_execute/add_169/carry[31] ), .Z(
        \u_a23_core/u_execute/rn_plus4[31] ) );
  AND U268 ( .A(\u_a23_core/u_decode/N527 ), .B(\u_a23_core/u_decode/N523 ), 
        .Z(\u_a23_core/u_decode/add_8_root_add_415_15/carry[1] ) );
  XOR U269 ( .A(\u_a23_core/u_decode/N527 ), .B(\u_a23_core/u_decode/N523 ), 
        .Z(\u_a23_core/u_decode/N542 ) );
  AND U270 ( .A(\u_a23_core/u_decode/N537 ), .B(\u_a23_core/u_decode/N532 ), 
        .Z(\u_a23_core/u_decode/add_7_root_add_415_15/carry[1] ) );
  XOR U271 ( .A(\u_a23_core/u_decode/N537 ), .B(\u_a23_core/u_decode/N532 ), 
        .Z(\u_a23_core/u_decode/N547 ) );
  AND U272 ( .A(\u_a23_core/u_decode/N539 ), .B(
        \u_a23_core/u_decode/add_7_root_add_415_15/carry[2] ), .Z(
        \u_a23_core/u_decode/N550 ) );
  XOR U273 ( .A(\u_a23_core/u_decode/N539 ), .B(
        \u_a23_core/u_decode/add_7_root_add_415_15/carry[2] ), .Z(
        \u_a23_core/u_decode/N549 ) );
  AND U274 ( .A(\u_a23_core/u_decode/N542 ), .B(\u_a23_core/u_decode/N547 ), 
        .Z(\u_a23_core/u_decode/add_6_root_add_415_15/carry[1] ) );
  XOR U275 ( .A(\u_a23_core/u_decode/N547 ), .B(\u_a23_core/u_decode/N542 ), 
        .Z(\u_a23_core/u_decode/mtrans_num_registers[0] ) );
  AND U276 ( .A(\u_a23_core/u_decode/N550 ), .B(
        \u_a23_core/u_decode/add_6_root_add_415_15/carry[3] ), .Z(
        \u_a23_core/u_decode/mtrans_num_registers[4] ) );
  XOR U277 ( .A(\u_a23_core/u_decode/N550 ), .B(
        \u_a23_core/u_decode/add_6_root_add_415_15/carry[3] ), .Z(
        \u_a23_core/u_decode/mtrans_num_registers[3] ) );
  MUX U278 ( .IN0(\u_a23_mem/stack_mem[0][0] ), .IN1(m_write[0]), .SEL(n1), 
        .F(\u_a23_mem/n19652 ) );
  MUX U279 ( .IN0(\u_a23_mem/stack_mem[0][1] ), .IN1(m_write[1]), .SEL(n1), 
        .F(\u_a23_mem/n19651 ) );
  MUX U280 ( .IN0(\u_a23_mem/stack_mem[0][2] ), .IN1(m_write[2]), .SEL(n1), 
        .F(\u_a23_mem/n19650 ) );
  MUX U281 ( .IN0(\u_a23_mem/stack_mem[0][3] ), .IN1(m_write[3]), .SEL(n1), 
        .F(\u_a23_mem/n19649 ) );
  MUX U282 ( .IN0(\u_a23_mem/stack_mem[0][4] ), .IN1(m_write[4]), .SEL(n1), 
        .F(\u_a23_mem/n19648 ) );
  MUX U283 ( .IN0(\u_a23_mem/stack_mem[0][5] ), .IN1(m_write[5]), .SEL(n1), 
        .F(\u_a23_mem/n19647 ) );
  MUX U284 ( .IN0(\u_a23_mem/stack_mem[0][6] ), .IN1(m_write[6]), .SEL(n1), 
        .F(\u_a23_mem/n19646 ) );
  MUX U285 ( .IN0(\u_a23_mem/stack_mem[0][7] ), .IN1(m_write[7]), .SEL(n1), 
        .F(\u_a23_mem/n19645 ) );
  NOR U286 ( .A(n2), .B(n3), .Z(n1) );
  NAND U287 ( .A(n4), .B(n5), .Z(\u_a23_mem/n19644 ) );
  NAND U288 ( .A(n6), .B(\u_a23_mem/stack_mem[1][0] ), .Z(n5) );
  AND U289 ( .A(n7), .B(n8), .Z(n4) );
  NANDN U290 ( .B(n3), .A(n9), .Z(n8) );
  OR U291 ( .A(n10), .B(n11), .Z(n7) );
  NAND U292 ( .A(n12), .B(n13), .Z(\u_a23_mem/n19643 ) );
  NAND U293 ( .A(n6), .B(\u_a23_mem/stack_mem[1][1] ), .Z(n13) );
  AND U294 ( .A(n14), .B(n15), .Z(n12) );
  NANDN U295 ( .B(n3), .A(n16), .Z(n15) );
  OR U296 ( .A(n10), .B(n17), .Z(n14) );
  NAND U297 ( .A(n18), .B(n19), .Z(\u_a23_mem/n19642 ) );
  NAND U298 ( .A(n6), .B(\u_a23_mem/stack_mem[1][2] ), .Z(n19) );
  AND U299 ( .A(n20), .B(n21), .Z(n18) );
  NANDN U300 ( .B(n3), .A(n22), .Z(n21) );
  OR U301 ( .A(n10), .B(n23), .Z(n20) );
  NAND U302 ( .A(n24), .B(n25), .Z(\u_a23_mem/n19641 ) );
  NAND U303 ( .A(n6), .B(\u_a23_mem/stack_mem[1][3] ), .Z(n25) );
  AND U304 ( .A(n26), .B(n27), .Z(n24) );
  NANDN U305 ( .B(n3), .A(n28), .Z(n27) );
  OR U306 ( .A(n10), .B(n29), .Z(n26) );
  NAND U307 ( .A(n30), .B(n31), .Z(\u_a23_mem/n19640 ) );
  NAND U308 ( .A(n6), .B(\u_a23_mem/stack_mem[1][4] ), .Z(n31) );
  AND U309 ( .A(n32), .B(n33), .Z(n30) );
  NANDN U310 ( .B(n3), .A(n34), .Z(n33) );
  OR U311 ( .A(n10), .B(n35), .Z(n32) );
  NAND U312 ( .A(n36), .B(n37), .Z(\u_a23_mem/n19639 ) );
  NAND U313 ( .A(n6), .B(\u_a23_mem/stack_mem[1][5] ), .Z(n37) );
  AND U314 ( .A(n38), .B(n39), .Z(n36) );
  NANDN U315 ( .B(n3), .A(n40), .Z(n39) );
  OR U316 ( .A(n10), .B(n41), .Z(n38) );
  NAND U317 ( .A(n42), .B(n43), .Z(\u_a23_mem/n19638 ) );
  NAND U318 ( .A(n6), .B(\u_a23_mem/stack_mem[1][6] ), .Z(n43) );
  AND U319 ( .A(n44), .B(n45), .Z(n42) );
  NANDN U320 ( .B(n3), .A(n46), .Z(n45) );
  OR U321 ( .A(n10), .B(n47), .Z(n44) );
  NAND U322 ( .A(n48), .B(n49), .Z(\u_a23_mem/n19637 ) );
  NAND U323 ( .A(n6), .B(\u_a23_mem/stack_mem[1][7] ), .Z(n49) );
  NANDN U324 ( .B(n3), .A(n50), .Z(n6) );
  AND U325 ( .A(n51), .B(n52), .Z(n48) );
  NANDN U326 ( .B(n3), .A(n53), .Z(n52) );
  OR U327 ( .A(n10), .B(n54), .Z(n51) );
  NAND U328 ( .A(n55), .B(n56), .Z(\u_a23_mem/n19636 ) );
  NAND U329 ( .A(n57), .B(\u_a23_mem/stack_mem[2][0] ), .Z(n56) );
  AND U330 ( .A(n58), .B(n59), .Z(n55) );
  NANDN U331 ( .B(n3), .A(n60), .Z(n59) );
  OR U332 ( .A(n11), .B(n61), .Z(n58) );
  NAND U333 ( .A(n62), .B(n63), .Z(\u_a23_mem/n19635 ) );
  NAND U334 ( .A(n57), .B(\u_a23_mem/stack_mem[2][1] ), .Z(n63) );
  AND U335 ( .A(n64), .B(n65), .Z(n62) );
  NANDN U336 ( .B(n3), .A(n66), .Z(n65) );
  OR U337 ( .A(n17), .B(n61), .Z(n64) );
  NAND U338 ( .A(n67), .B(n68), .Z(\u_a23_mem/n19634 ) );
  NAND U339 ( .A(n57), .B(\u_a23_mem/stack_mem[2][2] ), .Z(n68) );
  AND U340 ( .A(n69), .B(n70), .Z(n67) );
  NANDN U341 ( .B(n3), .A(n71), .Z(n70) );
  OR U342 ( .A(n23), .B(n61), .Z(n69) );
  NAND U343 ( .A(n72), .B(n73), .Z(\u_a23_mem/n19633 ) );
  NAND U344 ( .A(n57), .B(\u_a23_mem/stack_mem[2][3] ), .Z(n73) );
  AND U345 ( .A(n74), .B(n75), .Z(n72) );
  NANDN U346 ( .B(n3), .A(n76), .Z(n75) );
  OR U347 ( .A(n29), .B(n61), .Z(n74) );
  NAND U348 ( .A(n77), .B(n78), .Z(\u_a23_mem/n19632 ) );
  NAND U349 ( .A(n57), .B(\u_a23_mem/stack_mem[2][4] ), .Z(n78) );
  AND U350 ( .A(n79), .B(n80), .Z(n77) );
  NANDN U351 ( .B(n3), .A(n81), .Z(n80) );
  OR U352 ( .A(n35), .B(n61), .Z(n79) );
  NAND U353 ( .A(n82), .B(n83), .Z(\u_a23_mem/n19631 ) );
  NAND U354 ( .A(n57), .B(\u_a23_mem/stack_mem[2][5] ), .Z(n83) );
  AND U355 ( .A(n84), .B(n85), .Z(n82) );
  NANDN U356 ( .B(n3), .A(n86), .Z(n85) );
  OR U357 ( .A(n41), .B(n61), .Z(n84) );
  NAND U358 ( .A(n87), .B(n88), .Z(\u_a23_mem/n19630 ) );
  NAND U359 ( .A(n57), .B(\u_a23_mem/stack_mem[2][6] ), .Z(n88) );
  AND U360 ( .A(n89), .B(n90), .Z(n87) );
  NANDN U361 ( .B(n3), .A(n91), .Z(n90) );
  OR U362 ( .A(n47), .B(n61), .Z(n89) );
  NAND U363 ( .A(n92), .B(n93), .Z(\u_a23_mem/n19629 ) );
  NAND U364 ( .A(n57), .B(\u_a23_mem/stack_mem[2][7] ), .Z(n93) );
  NANDN U365 ( .B(n94), .A(n95), .Z(n57) );
  AND U366 ( .A(n96), .B(n97), .Z(n92) );
  NANDN U367 ( .B(n3), .A(n98), .Z(n97) );
  OR U368 ( .A(n54), .B(n61), .Z(n96) );
  NAND U369 ( .A(n99), .B(n100), .Z(\u_a23_mem/n19628 ) );
  NAND U370 ( .A(n101), .B(\u_a23_mem/stack_mem[3][0] ), .Z(n100) );
  AND U371 ( .A(n102), .B(n103), .Z(n99) );
  NANDN U372 ( .B(n3), .A(n104), .Z(n103) );
  OR U373 ( .A(n11), .B(n105), .Z(n102) );
  NAND U374 ( .A(n106), .B(n107), .Z(\u_a23_mem/n19627 ) );
  NAND U375 ( .A(n101), .B(\u_a23_mem/stack_mem[3][1] ), .Z(n107) );
  AND U376 ( .A(n108), .B(n109), .Z(n106) );
  NANDN U377 ( .B(n3), .A(n110), .Z(n109) );
  OR U378 ( .A(n17), .B(n105), .Z(n108) );
  NAND U379 ( .A(n111), .B(n112), .Z(\u_a23_mem/n19626 ) );
  NAND U380 ( .A(n101), .B(\u_a23_mem/stack_mem[3][2] ), .Z(n112) );
  AND U381 ( .A(n113), .B(n114), .Z(n111) );
  NANDN U382 ( .B(n3), .A(n115), .Z(n114) );
  OR U383 ( .A(n23), .B(n105), .Z(n113) );
  NAND U384 ( .A(n116), .B(n117), .Z(\u_a23_mem/n19625 ) );
  NAND U385 ( .A(n101), .B(\u_a23_mem/stack_mem[3][3] ), .Z(n117) );
  AND U386 ( .A(n118), .B(n119), .Z(n116) );
  NANDN U387 ( .B(n3), .A(n120), .Z(n119) );
  OR U388 ( .A(n29), .B(n105), .Z(n118) );
  NAND U389 ( .A(n121), .B(n122), .Z(\u_a23_mem/n19624 ) );
  NAND U390 ( .A(n101), .B(\u_a23_mem/stack_mem[3][4] ), .Z(n122) );
  AND U391 ( .A(n123), .B(n124), .Z(n121) );
  NANDN U392 ( .B(n3), .A(n125), .Z(n124) );
  OR U393 ( .A(n35), .B(n105), .Z(n123) );
  NAND U394 ( .A(n126), .B(n127), .Z(\u_a23_mem/n19623 ) );
  NAND U395 ( .A(n101), .B(\u_a23_mem/stack_mem[3][5] ), .Z(n127) );
  AND U396 ( .A(n128), .B(n129), .Z(n126) );
  NANDN U397 ( .B(n3), .A(n130), .Z(n129) );
  OR U398 ( .A(n41), .B(n105), .Z(n128) );
  NAND U399 ( .A(n131), .B(n132), .Z(\u_a23_mem/n19622 ) );
  NAND U400 ( .A(n101), .B(\u_a23_mem/stack_mem[3][6] ), .Z(n132) );
  AND U401 ( .A(n133), .B(n134), .Z(n131) );
  NANDN U402 ( .B(n3), .A(n135), .Z(n134) );
  OR U403 ( .A(n47), .B(n105), .Z(n133) );
  NAND U404 ( .A(n136), .B(n137), .Z(\u_a23_mem/n19621 ) );
  NAND U405 ( .A(n101), .B(\u_a23_mem/stack_mem[3][7] ), .Z(n137) );
  OR U406 ( .A(n138), .B(n139), .Z(n101) );
  AND U407 ( .A(n140), .B(n141), .Z(n136) );
  NANDN U408 ( .B(n3), .A(n142), .Z(n141) );
  NAND U409 ( .A(n143), .B(n95), .Z(n3) );
  OR U410 ( .A(n54), .B(n105), .Z(n140) );
  NAND U411 ( .A(n144), .B(n145), .Z(\u_a23_mem/n19620 ) );
  OR U412 ( .A(n11), .B(n146), .Z(n145) );
  NAND U413 ( .A(n147), .B(\u_a23_mem/stack_mem[4][0] ), .Z(n144) );
  NAND U414 ( .A(n148), .B(n149), .Z(\u_a23_mem/n19619 ) );
  OR U415 ( .A(n17), .B(n146), .Z(n149) );
  NAND U416 ( .A(n147), .B(\u_a23_mem/stack_mem[4][1] ), .Z(n148) );
  NAND U417 ( .A(n150), .B(n151), .Z(\u_a23_mem/n19618 ) );
  OR U418 ( .A(n23), .B(n146), .Z(n151) );
  NAND U419 ( .A(n147), .B(\u_a23_mem/stack_mem[4][2] ), .Z(n150) );
  NAND U420 ( .A(n152), .B(n153), .Z(\u_a23_mem/n19617 ) );
  OR U421 ( .A(n29), .B(n146), .Z(n153) );
  NAND U422 ( .A(n147), .B(\u_a23_mem/stack_mem[4][3] ), .Z(n152) );
  NAND U423 ( .A(n154), .B(n155), .Z(\u_a23_mem/n19616 ) );
  OR U424 ( .A(n35), .B(n146), .Z(n155) );
  NAND U425 ( .A(n147), .B(\u_a23_mem/stack_mem[4][4] ), .Z(n154) );
  NAND U426 ( .A(n156), .B(n157), .Z(\u_a23_mem/n19615 ) );
  OR U427 ( .A(n41), .B(n146), .Z(n157) );
  NAND U428 ( .A(n147), .B(\u_a23_mem/stack_mem[4][5] ), .Z(n156) );
  NAND U429 ( .A(n158), .B(n159), .Z(\u_a23_mem/n19614 ) );
  OR U430 ( .A(n47), .B(n146), .Z(n159) );
  NAND U431 ( .A(n147), .B(\u_a23_mem/stack_mem[4][6] ), .Z(n158) );
  NAND U432 ( .A(n160), .B(n161), .Z(\u_a23_mem/n19613 ) );
  OR U433 ( .A(n54), .B(n146), .Z(n161) );
  NAND U434 ( .A(n147), .B(\u_a23_mem/stack_mem[4][7] ), .Z(n160) );
  NANDN U435 ( .B(n162), .A(n163), .Z(n147) );
  NAND U436 ( .A(n164), .B(n165), .Z(\u_a23_mem/n19612 ) );
  NAND U437 ( .A(n166), .B(\u_a23_mem/stack_mem[5][0] ), .Z(n165) );
  AND U438 ( .A(n167), .B(n168), .Z(n164) );
  NANDN U439 ( .B(n169), .A(n9), .Z(n168) );
  OR U440 ( .A(n11), .B(n170), .Z(n167) );
  NAND U441 ( .A(n171), .B(n172), .Z(\u_a23_mem/n19611 ) );
  NAND U442 ( .A(n166), .B(\u_a23_mem/stack_mem[5][1] ), .Z(n172) );
  AND U443 ( .A(n173), .B(n174), .Z(n171) );
  NANDN U444 ( .B(n169), .A(n16), .Z(n174) );
  OR U445 ( .A(n17), .B(n170), .Z(n173) );
  NAND U446 ( .A(n175), .B(n176), .Z(\u_a23_mem/n19610 ) );
  NAND U447 ( .A(n166), .B(\u_a23_mem/stack_mem[5][2] ), .Z(n176) );
  AND U448 ( .A(n177), .B(n178), .Z(n175) );
  NANDN U449 ( .B(n169), .A(n22), .Z(n178) );
  OR U450 ( .A(n23), .B(n170), .Z(n177) );
  NAND U451 ( .A(n179), .B(n180), .Z(\u_a23_mem/n19609 ) );
  NAND U452 ( .A(n166), .B(\u_a23_mem/stack_mem[5][3] ), .Z(n180) );
  AND U453 ( .A(n181), .B(n182), .Z(n179) );
  NANDN U454 ( .B(n169), .A(n28), .Z(n182) );
  OR U455 ( .A(n29), .B(n170), .Z(n181) );
  NAND U456 ( .A(n183), .B(n184), .Z(\u_a23_mem/n19608 ) );
  NAND U457 ( .A(n166), .B(\u_a23_mem/stack_mem[5][4] ), .Z(n184) );
  AND U458 ( .A(n185), .B(n186), .Z(n183) );
  NANDN U459 ( .B(n169), .A(n34), .Z(n186) );
  OR U460 ( .A(n35), .B(n170), .Z(n185) );
  NAND U461 ( .A(n187), .B(n188), .Z(\u_a23_mem/n19607 ) );
  NAND U462 ( .A(n166), .B(\u_a23_mem/stack_mem[5][5] ), .Z(n188) );
  AND U463 ( .A(n189), .B(n190), .Z(n187) );
  NANDN U464 ( .B(n169), .A(n40), .Z(n190) );
  OR U465 ( .A(n41), .B(n170), .Z(n189) );
  NAND U466 ( .A(n191), .B(n192), .Z(\u_a23_mem/n19606 ) );
  NAND U467 ( .A(n166), .B(\u_a23_mem/stack_mem[5][6] ), .Z(n192) );
  AND U468 ( .A(n193), .B(n194), .Z(n191) );
  NANDN U469 ( .B(n169), .A(n46), .Z(n194) );
  OR U470 ( .A(n47), .B(n170), .Z(n193) );
  NAND U471 ( .A(n195), .B(n196), .Z(\u_a23_mem/n19605 ) );
  NAND U472 ( .A(n166), .B(\u_a23_mem/stack_mem[5][7] ), .Z(n196) );
  NANDN U473 ( .B(n197), .A(n163), .Z(n166) );
  AND U474 ( .A(n198), .B(n199), .Z(n195) );
  NANDN U475 ( .B(n169), .A(n53), .Z(n199) );
  OR U476 ( .A(n54), .B(n170), .Z(n198) );
  NAND U477 ( .A(n200), .B(n201), .Z(\u_a23_mem/n19604 ) );
  NAND U478 ( .A(n202), .B(\u_a23_mem/stack_mem[6][0] ), .Z(n201) );
  AND U479 ( .A(n203), .B(n204), .Z(n200) );
  NANDN U480 ( .B(n169), .A(n60), .Z(n204) );
  OR U481 ( .A(n11), .B(n205), .Z(n203) );
  NAND U482 ( .A(n206), .B(n207), .Z(\u_a23_mem/n19603 ) );
  NAND U483 ( .A(n202), .B(\u_a23_mem/stack_mem[6][1] ), .Z(n207) );
  AND U484 ( .A(n208), .B(n209), .Z(n206) );
  NANDN U485 ( .B(n169), .A(n66), .Z(n209) );
  OR U486 ( .A(n17), .B(n205), .Z(n208) );
  NAND U487 ( .A(n210), .B(n211), .Z(\u_a23_mem/n19602 ) );
  NAND U488 ( .A(n202), .B(\u_a23_mem/stack_mem[6][2] ), .Z(n211) );
  AND U489 ( .A(n212), .B(n213), .Z(n210) );
  NANDN U490 ( .B(n169), .A(n71), .Z(n213) );
  OR U491 ( .A(n23), .B(n205), .Z(n212) );
  NAND U492 ( .A(n214), .B(n215), .Z(\u_a23_mem/n19601 ) );
  NAND U493 ( .A(n202), .B(\u_a23_mem/stack_mem[6][3] ), .Z(n215) );
  AND U494 ( .A(n216), .B(n217), .Z(n214) );
  NANDN U495 ( .B(n169), .A(n76), .Z(n217) );
  OR U496 ( .A(n29), .B(n205), .Z(n216) );
  NAND U497 ( .A(n218), .B(n219), .Z(\u_a23_mem/n19600 ) );
  NAND U498 ( .A(n202), .B(\u_a23_mem/stack_mem[6][4] ), .Z(n219) );
  AND U499 ( .A(n220), .B(n221), .Z(n218) );
  NANDN U500 ( .B(n169), .A(n81), .Z(n221) );
  OR U501 ( .A(n35), .B(n205), .Z(n220) );
  NAND U502 ( .A(n222), .B(n223), .Z(\u_a23_mem/n19599 ) );
  NAND U503 ( .A(n202), .B(\u_a23_mem/stack_mem[6][5] ), .Z(n223) );
  AND U504 ( .A(n224), .B(n225), .Z(n222) );
  NANDN U505 ( .B(n169), .A(n86), .Z(n225) );
  OR U506 ( .A(n41), .B(n205), .Z(n224) );
  NAND U507 ( .A(n226), .B(n227), .Z(\u_a23_mem/n19598 ) );
  NAND U508 ( .A(n202), .B(\u_a23_mem/stack_mem[6][6] ), .Z(n227) );
  AND U509 ( .A(n228), .B(n229), .Z(n226) );
  NANDN U510 ( .B(n169), .A(n91), .Z(n229) );
  OR U511 ( .A(n47), .B(n205), .Z(n228) );
  NAND U512 ( .A(n230), .B(n231), .Z(\u_a23_mem/n19597 ) );
  NAND U513 ( .A(n202), .B(\u_a23_mem/stack_mem[6][7] ), .Z(n231) );
  NANDN U514 ( .B(n232), .A(n163), .Z(n202) );
  AND U515 ( .A(n233), .B(n234), .Z(n230) );
  NANDN U516 ( .B(n169), .A(n98), .Z(n234) );
  OR U517 ( .A(n54), .B(n205), .Z(n233) );
  NAND U518 ( .A(n235), .B(n236), .Z(\u_a23_mem/n19596 ) );
  NAND U519 ( .A(n237), .B(\u_a23_mem/stack_mem[7][0] ), .Z(n236) );
  AND U520 ( .A(n238), .B(n239), .Z(n235) );
  NANDN U521 ( .B(n169), .A(n104), .Z(n239) );
  OR U522 ( .A(n11), .B(n240), .Z(n238) );
  NAND U523 ( .A(n241), .B(n242), .Z(\u_a23_mem/n19595 ) );
  NAND U524 ( .A(n237), .B(\u_a23_mem/stack_mem[7][1] ), .Z(n242) );
  AND U525 ( .A(n243), .B(n244), .Z(n241) );
  NANDN U526 ( .B(n169), .A(n110), .Z(n244) );
  OR U527 ( .A(n17), .B(n240), .Z(n243) );
  NAND U528 ( .A(n245), .B(n246), .Z(\u_a23_mem/n19594 ) );
  NAND U529 ( .A(n237), .B(\u_a23_mem/stack_mem[7][2] ), .Z(n246) );
  AND U530 ( .A(n247), .B(n248), .Z(n245) );
  NANDN U531 ( .B(n169), .A(n115), .Z(n248) );
  OR U532 ( .A(n23), .B(n240), .Z(n247) );
  NAND U533 ( .A(n249), .B(n250), .Z(\u_a23_mem/n19593 ) );
  NAND U534 ( .A(n237), .B(\u_a23_mem/stack_mem[7][3] ), .Z(n250) );
  AND U535 ( .A(n251), .B(n252), .Z(n249) );
  NANDN U536 ( .B(n169), .A(n120), .Z(n252) );
  OR U537 ( .A(n29), .B(n240), .Z(n251) );
  NAND U538 ( .A(n253), .B(n254), .Z(\u_a23_mem/n19592 ) );
  NAND U539 ( .A(n237), .B(\u_a23_mem/stack_mem[7][4] ), .Z(n254) );
  AND U540 ( .A(n255), .B(n256), .Z(n253) );
  NANDN U541 ( .B(n169), .A(n125), .Z(n256) );
  OR U542 ( .A(n35), .B(n240), .Z(n255) );
  NAND U543 ( .A(n257), .B(n258), .Z(\u_a23_mem/n19591 ) );
  NAND U544 ( .A(n237), .B(\u_a23_mem/stack_mem[7][5] ), .Z(n258) );
  AND U545 ( .A(n259), .B(n260), .Z(n257) );
  NANDN U546 ( .B(n169), .A(n130), .Z(n260) );
  OR U547 ( .A(n41), .B(n240), .Z(n259) );
  NAND U548 ( .A(n261), .B(n262), .Z(\u_a23_mem/n19590 ) );
  NAND U549 ( .A(n237), .B(\u_a23_mem/stack_mem[7][6] ), .Z(n262) );
  AND U550 ( .A(n263), .B(n264), .Z(n261) );
  NANDN U551 ( .B(n169), .A(n135), .Z(n264) );
  OR U552 ( .A(n47), .B(n240), .Z(n263) );
  NAND U553 ( .A(n265), .B(n266), .Z(\u_a23_mem/n19589 ) );
  NAND U554 ( .A(n237), .B(\u_a23_mem/stack_mem[7][7] ), .Z(n266) );
  NANDN U555 ( .B(n138), .A(n163), .Z(n237) );
  AND U556 ( .A(n267), .B(n268), .Z(n265) );
  NANDN U557 ( .B(n169), .A(n142), .Z(n268) );
  NAND U558 ( .A(n163), .B(n95), .Z(n169) );
  OR U559 ( .A(n54), .B(n240), .Z(n267) );
  NAND U560 ( .A(n269), .B(n270), .Z(\u_a23_mem/n19588 ) );
  OR U561 ( .A(n11), .B(n271), .Z(n270) );
  NAND U562 ( .A(n272), .B(\u_a23_mem/stack_mem[8][0] ), .Z(n269) );
  NAND U563 ( .A(n273), .B(n274), .Z(\u_a23_mem/n19587 ) );
  OR U564 ( .A(n17), .B(n271), .Z(n274) );
  NAND U565 ( .A(n272), .B(\u_a23_mem/stack_mem[8][1] ), .Z(n273) );
  NAND U566 ( .A(n275), .B(n276), .Z(\u_a23_mem/n19586 ) );
  OR U567 ( .A(n23), .B(n271), .Z(n276) );
  NAND U568 ( .A(n272), .B(\u_a23_mem/stack_mem[8][2] ), .Z(n275) );
  NAND U569 ( .A(n277), .B(n278), .Z(\u_a23_mem/n19585 ) );
  OR U570 ( .A(n29), .B(n271), .Z(n278) );
  NAND U571 ( .A(n272), .B(\u_a23_mem/stack_mem[8][3] ), .Z(n277) );
  NAND U572 ( .A(n279), .B(n280), .Z(\u_a23_mem/n19584 ) );
  OR U573 ( .A(n35), .B(n271), .Z(n280) );
  NAND U574 ( .A(n272), .B(\u_a23_mem/stack_mem[8][4] ), .Z(n279) );
  NAND U575 ( .A(n281), .B(n282), .Z(\u_a23_mem/n19583 ) );
  OR U576 ( .A(n41), .B(n271), .Z(n282) );
  NAND U577 ( .A(n272), .B(\u_a23_mem/stack_mem[8][5] ), .Z(n281) );
  NAND U578 ( .A(n283), .B(n284), .Z(\u_a23_mem/n19582 ) );
  OR U579 ( .A(n47), .B(n271), .Z(n284) );
  NAND U580 ( .A(n272), .B(\u_a23_mem/stack_mem[8][6] ), .Z(n283) );
  NAND U581 ( .A(n285), .B(n286), .Z(\u_a23_mem/n19581 ) );
  OR U582 ( .A(n54), .B(n271), .Z(n286) );
  NAND U583 ( .A(n272), .B(\u_a23_mem/stack_mem[8][7] ), .Z(n285) );
  NANDN U584 ( .B(n162), .A(n287), .Z(n272) );
  NAND U585 ( .A(n288), .B(n289), .Z(\u_a23_mem/n19580 ) );
  NAND U586 ( .A(n290), .B(\u_a23_mem/stack_mem[9][0] ), .Z(n289) );
  AND U587 ( .A(n291), .B(n292), .Z(n288) );
  NANDN U588 ( .B(n293), .A(n9), .Z(n292) );
  OR U589 ( .A(n11), .B(n294), .Z(n291) );
  NAND U590 ( .A(n295), .B(n296), .Z(\u_a23_mem/n19579 ) );
  NAND U591 ( .A(n290), .B(\u_a23_mem/stack_mem[9][1] ), .Z(n296) );
  AND U592 ( .A(n297), .B(n298), .Z(n295) );
  NANDN U593 ( .B(n293), .A(n16), .Z(n298) );
  OR U594 ( .A(n17), .B(n294), .Z(n297) );
  NAND U595 ( .A(n299), .B(n300), .Z(\u_a23_mem/n19578 ) );
  NAND U596 ( .A(n290), .B(\u_a23_mem/stack_mem[9][2] ), .Z(n300) );
  AND U597 ( .A(n301), .B(n302), .Z(n299) );
  NANDN U598 ( .B(n293), .A(n22), .Z(n302) );
  OR U599 ( .A(n23), .B(n294), .Z(n301) );
  NAND U600 ( .A(n303), .B(n304), .Z(\u_a23_mem/n19577 ) );
  NAND U601 ( .A(n290), .B(\u_a23_mem/stack_mem[9][3] ), .Z(n304) );
  AND U602 ( .A(n305), .B(n306), .Z(n303) );
  NANDN U603 ( .B(n293), .A(n28), .Z(n306) );
  OR U604 ( .A(n29), .B(n294), .Z(n305) );
  NAND U605 ( .A(n307), .B(n308), .Z(\u_a23_mem/n19576 ) );
  NAND U606 ( .A(n290), .B(\u_a23_mem/stack_mem[9][4] ), .Z(n308) );
  AND U607 ( .A(n309), .B(n310), .Z(n307) );
  NANDN U608 ( .B(n293), .A(n34), .Z(n310) );
  OR U609 ( .A(n35), .B(n294), .Z(n309) );
  NAND U610 ( .A(n311), .B(n312), .Z(\u_a23_mem/n19575 ) );
  NAND U611 ( .A(n290), .B(\u_a23_mem/stack_mem[9][5] ), .Z(n312) );
  AND U612 ( .A(n313), .B(n314), .Z(n311) );
  NANDN U613 ( .B(n293), .A(n40), .Z(n314) );
  OR U614 ( .A(n41), .B(n294), .Z(n313) );
  NAND U615 ( .A(n315), .B(n316), .Z(\u_a23_mem/n19574 ) );
  NAND U616 ( .A(n290), .B(\u_a23_mem/stack_mem[9][6] ), .Z(n316) );
  AND U617 ( .A(n317), .B(n318), .Z(n315) );
  NANDN U618 ( .B(n293), .A(n46), .Z(n318) );
  OR U619 ( .A(n47), .B(n294), .Z(n317) );
  NAND U620 ( .A(n319), .B(n320), .Z(\u_a23_mem/n19573 ) );
  NAND U621 ( .A(n290), .B(\u_a23_mem/stack_mem[9][7] ), .Z(n320) );
  NANDN U622 ( .B(n197), .A(n287), .Z(n290) );
  AND U623 ( .A(n321), .B(n322), .Z(n319) );
  NANDN U624 ( .B(n293), .A(n53), .Z(n322) );
  OR U625 ( .A(n54), .B(n294), .Z(n321) );
  NAND U626 ( .A(n323), .B(n324), .Z(\u_a23_mem/n19572 ) );
  NAND U627 ( .A(n325), .B(\u_a23_mem/stack_mem[10][0] ), .Z(n324) );
  AND U628 ( .A(n326), .B(n327), .Z(n323) );
  NANDN U629 ( .B(n293), .A(n60), .Z(n327) );
  OR U630 ( .A(n11), .B(n328), .Z(n326) );
  NAND U631 ( .A(n329), .B(n330), .Z(\u_a23_mem/n19571 ) );
  NAND U632 ( .A(n325), .B(\u_a23_mem/stack_mem[10][1] ), .Z(n330) );
  AND U633 ( .A(n331), .B(n332), .Z(n329) );
  NANDN U634 ( .B(n293), .A(n66), .Z(n332) );
  OR U635 ( .A(n17), .B(n328), .Z(n331) );
  NAND U636 ( .A(n333), .B(n334), .Z(\u_a23_mem/n19570 ) );
  NAND U637 ( .A(n325), .B(\u_a23_mem/stack_mem[10][2] ), .Z(n334) );
  AND U638 ( .A(n335), .B(n336), .Z(n333) );
  NANDN U639 ( .B(n293), .A(n71), .Z(n336) );
  OR U640 ( .A(n23), .B(n328), .Z(n335) );
  NAND U641 ( .A(n337), .B(n338), .Z(\u_a23_mem/n19569 ) );
  NAND U642 ( .A(n325), .B(\u_a23_mem/stack_mem[10][3] ), .Z(n338) );
  AND U643 ( .A(n339), .B(n340), .Z(n337) );
  NANDN U644 ( .B(n293), .A(n76), .Z(n340) );
  OR U645 ( .A(n29), .B(n328), .Z(n339) );
  NAND U646 ( .A(n341), .B(n342), .Z(\u_a23_mem/n19568 ) );
  NAND U647 ( .A(n325), .B(\u_a23_mem/stack_mem[10][4] ), .Z(n342) );
  AND U648 ( .A(n343), .B(n344), .Z(n341) );
  NANDN U649 ( .B(n293), .A(n81), .Z(n344) );
  OR U650 ( .A(n35), .B(n328), .Z(n343) );
  NAND U651 ( .A(n345), .B(n346), .Z(\u_a23_mem/n19567 ) );
  NAND U652 ( .A(n325), .B(\u_a23_mem/stack_mem[10][5] ), .Z(n346) );
  AND U653 ( .A(n347), .B(n348), .Z(n345) );
  NANDN U654 ( .B(n293), .A(n86), .Z(n348) );
  OR U655 ( .A(n41), .B(n328), .Z(n347) );
  NAND U656 ( .A(n349), .B(n350), .Z(\u_a23_mem/n19566 ) );
  NAND U657 ( .A(n325), .B(\u_a23_mem/stack_mem[10][6] ), .Z(n350) );
  AND U658 ( .A(n351), .B(n352), .Z(n349) );
  NANDN U659 ( .B(n293), .A(n91), .Z(n352) );
  OR U660 ( .A(n47), .B(n328), .Z(n351) );
  NAND U661 ( .A(n353), .B(n354), .Z(\u_a23_mem/n19565 ) );
  NAND U662 ( .A(n325), .B(\u_a23_mem/stack_mem[10][7] ), .Z(n354) );
  NANDN U663 ( .B(n232), .A(n287), .Z(n325) );
  AND U664 ( .A(n355), .B(n356), .Z(n353) );
  NANDN U665 ( .B(n293), .A(n98), .Z(n356) );
  OR U666 ( .A(n54), .B(n328), .Z(n355) );
  NAND U667 ( .A(n357), .B(n358), .Z(\u_a23_mem/n19564 ) );
  NAND U668 ( .A(n359), .B(\u_a23_mem/stack_mem[11][0] ), .Z(n358) );
  AND U669 ( .A(n360), .B(n361), .Z(n357) );
  NANDN U670 ( .B(n293), .A(n104), .Z(n361) );
  OR U671 ( .A(n11), .B(n362), .Z(n360) );
  NAND U672 ( .A(n363), .B(n364), .Z(\u_a23_mem/n19563 ) );
  NAND U673 ( .A(n359), .B(\u_a23_mem/stack_mem[11][1] ), .Z(n364) );
  AND U674 ( .A(n365), .B(n366), .Z(n363) );
  NANDN U675 ( .B(n293), .A(n110), .Z(n366) );
  OR U676 ( .A(n17), .B(n362), .Z(n365) );
  NAND U677 ( .A(n367), .B(n368), .Z(\u_a23_mem/n19562 ) );
  NAND U678 ( .A(n359), .B(\u_a23_mem/stack_mem[11][2] ), .Z(n368) );
  AND U679 ( .A(n369), .B(n370), .Z(n367) );
  NANDN U680 ( .B(n293), .A(n115), .Z(n370) );
  OR U681 ( .A(n23), .B(n362), .Z(n369) );
  NAND U682 ( .A(n371), .B(n372), .Z(\u_a23_mem/n19561 ) );
  NAND U683 ( .A(n359), .B(\u_a23_mem/stack_mem[11][3] ), .Z(n372) );
  AND U684 ( .A(n373), .B(n374), .Z(n371) );
  NANDN U685 ( .B(n293), .A(n120), .Z(n374) );
  OR U686 ( .A(n29), .B(n362), .Z(n373) );
  NAND U687 ( .A(n375), .B(n376), .Z(\u_a23_mem/n19560 ) );
  NAND U688 ( .A(n359), .B(\u_a23_mem/stack_mem[11][4] ), .Z(n376) );
  AND U689 ( .A(n377), .B(n378), .Z(n375) );
  NANDN U690 ( .B(n293), .A(n125), .Z(n378) );
  OR U691 ( .A(n35), .B(n362), .Z(n377) );
  NAND U692 ( .A(n379), .B(n380), .Z(\u_a23_mem/n19559 ) );
  NAND U693 ( .A(n359), .B(\u_a23_mem/stack_mem[11][5] ), .Z(n380) );
  AND U694 ( .A(n381), .B(n382), .Z(n379) );
  NANDN U695 ( .B(n293), .A(n130), .Z(n382) );
  OR U696 ( .A(n41), .B(n362), .Z(n381) );
  NAND U697 ( .A(n383), .B(n384), .Z(\u_a23_mem/n19558 ) );
  NAND U698 ( .A(n359), .B(\u_a23_mem/stack_mem[11][6] ), .Z(n384) );
  AND U699 ( .A(n385), .B(n386), .Z(n383) );
  NANDN U700 ( .B(n293), .A(n135), .Z(n386) );
  OR U701 ( .A(n47), .B(n362), .Z(n385) );
  NAND U702 ( .A(n387), .B(n388), .Z(\u_a23_mem/n19557 ) );
  NAND U703 ( .A(n359), .B(\u_a23_mem/stack_mem[11][7] ), .Z(n388) );
  NANDN U704 ( .B(n138), .A(n287), .Z(n359) );
  AND U705 ( .A(n389), .B(n390), .Z(n387) );
  NANDN U706 ( .B(n293), .A(n142), .Z(n390) );
  NAND U707 ( .A(n287), .B(n95), .Z(n293) );
  OR U708 ( .A(n54), .B(n362), .Z(n389) );
  NAND U709 ( .A(n391), .B(n392), .Z(\u_a23_mem/n19556 ) );
  OR U710 ( .A(n11), .B(n393), .Z(n392) );
  NAND U711 ( .A(n394), .B(\u_a23_mem/stack_mem[12][0] ), .Z(n391) );
  NAND U712 ( .A(n395), .B(n396), .Z(\u_a23_mem/n19555 ) );
  OR U713 ( .A(n17), .B(n393), .Z(n396) );
  NAND U714 ( .A(n394), .B(\u_a23_mem/stack_mem[12][1] ), .Z(n395) );
  NAND U715 ( .A(n397), .B(n398), .Z(\u_a23_mem/n19554 ) );
  OR U716 ( .A(n23), .B(n393), .Z(n398) );
  NAND U717 ( .A(n394), .B(\u_a23_mem/stack_mem[12][2] ), .Z(n397) );
  NAND U718 ( .A(n399), .B(n400), .Z(\u_a23_mem/n19553 ) );
  OR U719 ( .A(n29), .B(n393), .Z(n400) );
  NAND U720 ( .A(n394), .B(\u_a23_mem/stack_mem[12][3] ), .Z(n399) );
  NAND U721 ( .A(n401), .B(n402), .Z(\u_a23_mem/n19552 ) );
  OR U722 ( .A(n35), .B(n393), .Z(n402) );
  NAND U723 ( .A(n394), .B(\u_a23_mem/stack_mem[12][4] ), .Z(n401) );
  NAND U724 ( .A(n403), .B(n404), .Z(\u_a23_mem/n19551 ) );
  OR U725 ( .A(n41), .B(n393), .Z(n404) );
  NAND U726 ( .A(n394), .B(\u_a23_mem/stack_mem[12][5] ), .Z(n403) );
  NAND U727 ( .A(n405), .B(n406), .Z(\u_a23_mem/n19550 ) );
  OR U728 ( .A(n47), .B(n393), .Z(n406) );
  NAND U729 ( .A(n394), .B(\u_a23_mem/stack_mem[12][6] ), .Z(n405) );
  NAND U730 ( .A(n407), .B(n408), .Z(\u_a23_mem/n19549 ) );
  OR U731 ( .A(n54), .B(n393), .Z(n408) );
  NAND U732 ( .A(n394), .B(\u_a23_mem/stack_mem[12][7] ), .Z(n407) );
  NANDN U733 ( .B(n162), .A(n409), .Z(n394) );
  NAND U734 ( .A(n410), .B(n411), .Z(\u_a23_mem/n19548 ) );
  NAND U735 ( .A(n412), .B(\u_a23_mem/stack_mem[13][0] ), .Z(n411) );
  AND U736 ( .A(n413), .B(n414), .Z(n410) );
  NANDN U737 ( .B(n415), .A(n9), .Z(n414) );
  OR U738 ( .A(n11), .B(n416), .Z(n413) );
  NAND U739 ( .A(n417), .B(n418), .Z(\u_a23_mem/n19547 ) );
  NAND U740 ( .A(n412), .B(\u_a23_mem/stack_mem[13][1] ), .Z(n418) );
  AND U741 ( .A(n419), .B(n420), .Z(n417) );
  NANDN U742 ( .B(n415), .A(n16), .Z(n420) );
  OR U743 ( .A(n17), .B(n416), .Z(n419) );
  NAND U744 ( .A(n421), .B(n422), .Z(\u_a23_mem/n19546 ) );
  NAND U745 ( .A(n412), .B(\u_a23_mem/stack_mem[13][2] ), .Z(n422) );
  AND U746 ( .A(n423), .B(n424), .Z(n421) );
  NANDN U747 ( .B(n415), .A(n22), .Z(n424) );
  OR U748 ( .A(n23), .B(n416), .Z(n423) );
  NAND U749 ( .A(n425), .B(n426), .Z(\u_a23_mem/n19545 ) );
  NAND U750 ( .A(n412), .B(\u_a23_mem/stack_mem[13][3] ), .Z(n426) );
  AND U751 ( .A(n427), .B(n428), .Z(n425) );
  NANDN U752 ( .B(n415), .A(n28), .Z(n428) );
  OR U753 ( .A(n29), .B(n416), .Z(n427) );
  NAND U754 ( .A(n429), .B(n430), .Z(\u_a23_mem/n19544 ) );
  NAND U755 ( .A(n412), .B(\u_a23_mem/stack_mem[13][4] ), .Z(n430) );
  AND U756 ( .A(n431), .B(n432), .Z(n429) );
  NANDN U757 ( .B(n415), .A(n34), .Z(n432) );
  OR U758 ( .A(n35), .B(n416), .Z(n431) );
  NAND U759 ( .A(n433), .B(n434), .Z(\u_a23_mem/n19543 ) );
  NAND U760 ( .A(n412), .B(\u_a23_mem/stack_mem[13][5] ), .Z(n434) );
  AND U761 ( .A(n435), .B(n436), .Z(n433) );
  NANDN U762 ( .B(n415), .A(n40), .Z(n436) );
  OR U763 ( .A(n41), .B(n416), .Z(n435) );
  NAND U764 ( .A(n437), .B(n438), .Z(\u_a23_mem/n19542 ) );
  NAND U765 ( .A(n412), .B(\u_a23_mem/stack_mem[13][6] ), .Z(n438) );
  AND U766 ( .A(n439), .B(n440), .Z(n437) );
  NANDN U767 ( .B(n415), .A(n46), .Z(n440) );
  OR U768 ( .A(n47), .B(n416), .Z(n439) );
  NAND U769 ( .A(n441), .B(n442), .Z(\u_a23_mem/n19541 ) );
  NAND U770 ( .A(n412), .B(\u_a23_mem/stack_mem[13][7] ), .Z(n442) );
  NANDN U771 ( .B(n197), .A(n409), .Z(n412) );
  AND U772 ( .A(n443), .B(n444), .Z(n441) );
  NANDN U773 ( .B(n415), .A(n53), .Z(n444) );
  OR U774 ( .A(n54), .B(n416), .Z(n443) );
  NAND U775 ( .A(n445), .B(n446), .Z(\u_a23_mem/n19540 ) );
  NAND U776 ( .A(n447), .B(\u_a23_mem/stack_mem[14][0] ), .Z(n446) );
  AND U777 ( .A(n448), .B(n449), .Z(n445) );
  NANDN U778 ( .B(n415), .A(n60), .Z(n449) );
  OR U779 ( .A(n11), .B(n450), .Z(n448) );
  NAND U780 ( .A(n451), .B(n452), .Z(\u_a23_mem/n19539 ) );
  NAND U781 ( .A(n447), .B(\u_a23_mem/stack_mem[14][1] ), .Z(n452) );
  AND U782 ( .A(n453), .B(n454), .Z(n451) );
  NANDN U783 ( .B(n415), .A(n66), .Z(n454) );
  OR U784 ( .A(n17), .B(n450), .Z(n453) );
  NAND U785 ( .A(n455), .B(n456), .Z(\u_a23_mem/n19538 ) );
  NAND U786 ( .A(n447), .B(\u_a23_mem/stack_mem[14][2] ), .Z(n456) );
  AND U787 ( .A(n457), .B(n458), .Z(n455) );
  NANDN U788 ( .B(n415), .A(n71), .Z(n458) );
  OR U789 ( .A(n23), .B(n450), .Z(n457) );
  NAND U790 ( .A(n459), .B(n460), .Z(\u_a23_mem/n19537 ) );
  NAND U791 ( .A(n447), .B(\u_a23_mem/stack_mem[14][3] ), .Z(n460) );
  AND U792 ( .A(n461), .B(n462), .Z(n459) );
  NANDN U793 ( .B(n415), .A(n76), .Z(n462) );
  OR U794 ( .A(n29), .B(n450), .Z(n461) );
  NAND U795 ( .A(n463), .B(n464), .Z(\u_a23_mem/n19536 ) );
  NAND U796 ( .A(n447), .B(\u_a23_mem/stack_mem[14][4] ), .Z(n464) );
  AND U797 ( .A(n465), .B(n466), .Z(n463) );
  NANDN U798 ( .B(n415), .A(n81), .Z(n466) );
  OR U799 ( .A(n35), .B(n450), .Z(n465) );
  NAND U800 ( .A(n467), .B(n468), .Z(\u_a23_mem/n19535 ) );
  NAND U801 ( .A(n447), .B(\u_a23_mem/stack_mem[14][5] ), .Z(n468) );
  AND U802 ( .A(n469), .B(n470), .Z(n467) );
  NANDN U803 ( .B(n415), .A(n86), .Z(n470) );
  OR U804 ( .A(n41), .B(n450), .Z(n469) );
  NAND U805 ( .A(n471), .B(n472), .Z(\u_a23_mem/n19534 ) );
  NAND U806 ( .A(n447), .B(\u_a23_mem/stack_mem[14][6] ), .Z(n472) );
  AND U807 ( .A(n473), .B(n474), .Z(n471) );
  NANDN U808 ( .B(n415), .A(n91), .Z(n474) );
  OR U809 ( .A(n47), .B(n450), .Z(n473) );
  NAND U810 ( .A(n475), .B(n476), .Z(\u_a23_mem/n19533 ) );
  NAND U811 ( .A(n447), .B(\u_a23_mem/stack_mem[14][7] ), .Z(n476) );
  NANDN U812 ( .B(n232), .A(n409), .Z(n447) );
  AND U813 ( .A(n477), .B(n478), .Z(n475) );
  NANDN U814 ( .B(n415), .A(n98), .Z(n478) );
  OR U815 ( .A(n54), .B(n450), .Z(n477) );
  NAND U816 ( .A(n479), .B(n480), .Z(\u_a23_mem/n19532 ) );
  NAND U817 ( .A(n481), .B(\u_a23_mem/stack_mem[15][0] ), .Z(n480) );
  AND U818 ( .A(n482), .B(n483), .Z(n479) );
  NANDN U819 ( .B(n415), .A(n104), .Z(n483) );
  OR U820 ( .A(n11), .B(n484), .Z(n482) );
  NAND U821 ( .A(n485), .B(n486), .Z(\u_a23_mem/n19531 ) );
  NAND U822 ( .A(n481), .B(\u_a23_mem/stack_mem[15][1] ), .Z(n486) );
  AND U823 ( .A(n487), .B(n488), .Z(n485) );
  NANDN U824 ( .B(n415), .A(n110), .Z(n488) );
  OR U825 ( .A(n17), .B(n484), .Z(n487) );
  NAND U826 ( .A(n489), .B(n490), .Z(\u_a23_mem/n19530 ) );
  NAND U827 ( .A(n481), .B(\u_a23_mem/stack_mem[15][2] ), .Z(n490) );
  AND U828 ( .A(n491), .B(n492), .Z(n489) );
  NANDN U829 ( .B(n415), .A(n115), .Z(n492) );
  OR U830 ( .A(n23), .B(n484), .Z(n491) );
  NAND U831 ( .A(n493), .B(n494), .Z(\u_a23_mem/n19529 ) );
  NAND U832 ( .A(n481), .B(\u_a23_mem/stack_mem[15][3] ), .Z(n494) );
  AND U833 ( .A(n495), .B(n496), .Z(n493) );
  NANDN U834 ( .B(n415), .A(n120), .Z(n496) );
  OR U835 ( .A(n29), .B(n484), .Z(n495) );
  NAND U836 ( .A(n497), .B(n498), .Z(\u_a23_mem/n19528 ) );
  NAND U837 ( .A(n481), .B(\u_a23_mem/stack_mem[15][4] ), .Z(n498) );
  AND U838 ( .A(n499), .B(n500), .Z(n497) );
  NANDN U839 ( .B(n415), .A(n125), .Z(n500) );
  OR U840 ( .A(n35), .B(n484), .Z(n499) );
  NAND U841 ( .A(n501), .B(n502), .Z(\u_a23_mem/n19527 ) );
  NAND U842 ( .A(n481), .B(\u_a23_mem/stack_mem[15][5] ), .Z(n502) );
  AND U843 ( .A(n503), .B(n504), .Z(n501) );
  NANDN U844 ( .B(n415), .A(n130), .Z(n504) );
  OR U845 ( .A(n41), .B(n484), .Z(n503) );
  NAND U846 ( .A(n505), .B(n506), .Z(\u_a23_mem/n19526 ) );
  NAND U847 ( .A(n481), .B(\u_a23_mem/stack_mem[15][6] ), .Z(n506) );
  AND U848 ( .A(n507), .B(n508), .Z(n505) );
  NANDN U849 ( .B(n415), .A(n135), .Z(n508) );
  OR U850 ( .A(n47), .B(n484), .Z(n507) );
  NAND U851 ( .A(n509), .B(n510), .Z(\u_a23_mem/n19525 ) );
  NAND U852 ( .A(n481), .B(\u_a23_mem/stack_mem[15][7] ), .Z(n510) );
  NANDN U853 ( .B(n138), .A(n409), .Z(n481) );
  AND U854 ( .A(n511), .B(n512), .Z(n509) );
  NANDN U855 ( .B(n415), .A(n142), .Z(n512) );
  NAND U856 ( .A(n409), .B(n95), .Z(n415) );
  OR U857 ( .A(n54), .B(n484), .Z(n511) );
  NAND U858 ( .A(n513), .B(n514), .Z(\u_a23_mem/n19524 ) );
  OR U859 ( .A(n11), .B(n515), .Z(n514) );
  NAND U860 ( .A(n516), .B(\u_a23_mem/stack_mem[16][0] ), .Z(n513) );
  NAND U861 ( .A(n517), .B(n518), .Z(\u_a23_mem/n19523 ) );
  OR U862 ( .A(n17), .B(n515), .Z(n518) );
  NAND U863 ( .A(n516), .B(\u_a23_mem/stack_mem[16][1] ), .Z(n517) );
  NAND U864 ( .A(n519), .B(n520), .Z(\u_a23_mem/n19522 ) );
  OR U865 ( .A(n23), .B(n515), .Z(n520) );
  NAND U866 ( .A(n516), .B(\u_a23_mem/stack_mem[16][2] ), .Z(n519) );
  NAND U867 ( .A(n521), .B(n522), .Z(\u_a23_mem/n19521 ) );
  OR U868 ( .A(n29), .B(n515), .Z(n522) );
  NAND U869 ( .A(n516), .B(\u_a23_mem/stack_mem[16][3] ), .Z(n521) );
  NAND U870 ( .A(n523), .B(n524), .Z(\u_a23_mem/n19520 ) );
  OR U871 ( .A(n35), .B(n515), .Z(n524) );
  NAND U872 ( .A(n516), .B(\u_a23_mem/stack_mem[16][4] ), .Z(n523) );
  NAND U873 ( .A(n525), .B(n526), .Z(\u_a23_mem/n19519 ) );
  OR U874 ( .A(n41), .B(n515), .Z(n526) );
  NAND U875 ( .A(n516), .B(\u_a23_mem/stack_mem[16][5] ), .Z(n525) );
  NAND U876 ( .A(n527), .B(n528), .Z(\u_a23_mem/n19518 ) );
  OR U877 ( .A(n47), .B(n515), .Z(n528) );
  NAND U878 ( .A(n516), .B(\u_a23_mem/stack_mem[16][6] ), .Z(n527) );
  NAND U879 ( .A(n529), .B(n530), .Z(\u_a23_mem/n19517 ) );
  OR U880 ( .A(n54), .B(n515), .Z(n530) );
  NAND U881 ( .A(n516), .B(\u_a23_mem/stack_mem[16][7] ), .Z(n529) );
  NANDN U882 ( .B(n162), .A(n531), .Z(n516) );
  NAND U883 ( .A(n532), .B(n533), .Z(\u_a23_mem/n19516 ) );
  NAND U884 ( .A(n534), .B(\u_a23_mem/stack_mem[17][0] ), .Z(n533) );
  AND U885 ( .A(n535), .B(n536), .Z(n532) );
  NANDN U886 ( .B(n537), .A(n9), .Z(n536) );
  OR U887 ( .A(n11), .B(n538), .Z(n535) );
  NAND U888 ( .A(n539), .B(n540), .Z(\u_a23_mem/n19515 ) );
  NAND U889 ( .A(n534), .B(\u_a23_mem/stack_mem[17][1] ), .Z(n540) );
  AND U890 ( .A(n541), .B(n542), .Z(n539) );
  NANDN U891 ( .B(n537), .A(n16), .Z(n542) );
  OR U892 ( .A(n17), .B(n538), .Z(n541) );
  NAND U893 ( .A(n543), .B(n544), .Z(\u_a23_mem/n19514 ) );
  NAND U894 ( .A(n534), .B(\u_a23_mem/stack_mem[17][2] ), .Z(n544) );
  AND U895 ( .A(n545), .B(n546), .Z(n543) );
  NANDN U896 ( .B(n537), .A(n22), .Z(n546) );
  OR U897 ( .A(n23), .B(n538), .Z(n545) );
  NAND U898 ( .A(n547), .B(n548), .Z(\u_a23_mem/n19513 ) );
  NAND U899 ( .A(n534), .B(\u_a23_mem/stack_mem[17][3] ), .Z(n548) );
  AND U900 ( .A(n549), .B(n550), .Z(n547) );
  NANDN U901 ( .B(n537), .A(n28), .Z(n550) );
  OR U902 ( .A(n29), .B(n538), .Z(n549) );
  NAND U903 ( .A(n551), .B(n552), .Z(\u_a23_mem/n19512 ) );
  NAND U904 ( .A(n534), .B(\u_a23_mem/stack_mem[17][4] ), .Z(n552) );
  AND U905 ( .A(n553), .B(n554), .Z(n551) );
  NANDN U906 ( .B(n537), .A(n34), .Z(n554) );
  OR U907 ( .A(n35), .B(n538), .Z(n553) );
  NAND U908 ( .A(n555), .B(n556), .Z(\u_a23_mem/n19511 ) );
  NAND U909 ( .A(n534), .B(\u_a23_mem/stack_mem[17][5] ), .Z(n556) );
  AND U910 ( .A(n557), .B(n558), .Z(n555) );
  NANDN U911 ( .B(n537), .A(n40), .Z(n558) );
  OR U912 ( .A(n41), .B(n538), .Z(n557) );
  NAND U913 ( .A(n559), .B(n560), .Z(\u_a23_mem/n19510 ) );
  NAND U914 ( .A(n534), .B(\u_a23_mem/stack_mem[17][6] ), .Z(n560) );
  AND U915 ( .A(n561), .B(n562), .Z(n559) );
  NANDN U916 ( .B(n537), .A(n46), .Z(n562) );
  OR U917 ( .A(n47), .B(n538), .Z(n561) );
  NAND U918 ( .A(n563), .B(n564), .Z(\u_a23_mem/n19509 ) );
  NAND U919 ( .A(n534), .B(\u_a23_mem/stack_mem[17][7] ), .Z(n564) );
  NANDN U920 ( .B(n197), .A(n531), .Z(n534) );
  AND U921 ( .A(n565), .B(n566), .Z(n563) );
  NANDN U922 ( .B(n537), .A(n53), .Z(n566) );
  OR U923 ( .A(n54), .B(n538), .Z(n565) );
  NAND U924 ( .A(n567), .B(n568), .Z(\u_a23_mem/n19508 ) );
  NAND U925 ( .A(n569), .B(\u_a23_mem/stack_mem[18][0] ), .Z(n568) );
  AND U926 ( .A(n570), .B(n571), .Z(n567) );
  NANDN U927 ( .B(n537), .A(n60), .Z(n571) );
  OR U928 ( .A(n11), .B(n572), .Z(n570) );
  NAND U929 ( .A(n573), .B(n574), .Z(\u_a23_mem/n19507 ) );
  NAND U930 ( .A(n569), .B(\u_a23_mem/stack_mem[18][1] ), .Z(n574) );
  AND U931 ( .A(n575), .B(n576), .Z(n573) );
  NANDN U932 ( .B(n537), .A(n66), .Z(n576) );
  OR U933 ( .A(n17), .B(n572), .Z(n575) );
  NAND U934 ( .A(n577), .B(n578), .Z(\u_a23_mem/n19506 ) );
  NAND U935 ( .A(n569), .B(\u_a23_mem/stack_mem[18][2] ), .Z(n578) );
  AND U936 ( .A(n579), .B(n580), .Z(n577) );
  NANDN U937 ( .B(n537), .A(n71), .Z(n580) );
  OR U938 ( .A(n23), .B(n572), .Z(n579) );
  NAND U939 ( .A(n581), .B(n582), .Z(\u_a23_mem/n19505 ) );
  NAND U940 ( .A(n569), .B(\u_a23_mem/stack_mem[18][3] ), .Z(n582) );
  AND U941 ( .A(n583), .B(n584), .Z(n581) );
  NANDN U942 ( .B(n537), .A(n76), .Z(n584) );
  OR U943 ( .A(n29), .B(n572), .Z(n583) );
  NAND U944 ( .A(n585), .B(n586), .Z(\u_a23_mem/n19504 ) );
  NAND U945 ( .A(n569), .B(\u_a23_mem/stack_mem[18][4] ), .Z(n586) );
  AND U946 ( .A(n587), .B(n588), .Z(n585) );
  NANDN U947 ( .B(n537), .A(n81), .Z(n588) );
  OR U948 ( .A(n35), .B(n572), .Z(n587) );
  NAND U949 ( .A(n589), .B(n590), .Z(\u_a23_mem/n19503 ) );
  NAND U950 ( .A(n569), .B(\u_a23_mem/stack_mem[18][5] ), .Z(n590) );
  AND U951 ( .A(n591), .B(n592), .Z(n589) );
  NANDN U952 ( .B(n537), .A(n86), .Z(n592) );
  OR U953 ( .A(n41), .B(n572), .Z(n591) );
  NAND U954 ( .A(n593), .B(n594), .Z(\u_a23_mem/n19502 ) );
  NAND U955 ( .A(n569), .B(\u_a23_mem/stack_mem[18][6] ), .Z(n594) );
  AND U956 ( .A(n595), .B(n596), .Z(n593) );
  NANDN U957 ( .B(n537), .A(n91), .Z(n596) );
  OR U958 ( .A(n47), .B(n572), .Z(n595) );
  NAND U959 ( .A(n597), .B(n598), .Z(\u_a23_mem/n19501 ) );
  NAND U960 ( .A(n569), .B(\u_a23_mem/stack_mem[18][7] ), .Z(n598) );
  NANDN U961 ( .B(n232), .A(n531), .Z(n569) );
  AND U962 ( .A(n599), .B(n600), .Z(n597) );
  NANDN U963 ( .B(n537), .A(n98), .Z(n600) );
  OR U964 ( .A(n54), .B(n572), .Z(n599) );
  NAND U965 ( .A(n601), .B(n602), .Z(\u_a23_mem/n19500 ) );
  NAND U966 ( .A(n603), .B(\u_a23_mem/stack_mem[19][0] ), .Z(n602) );
  AND U967 ( .A(n604), .B(n605), .Z(n601) );
  NANDN U968 ( .B(n537), .A(n104), .Z(n605) );
  OR U969 ( .A(n11), .B(n606), .Z(n604) );
  NAND U970 ( .A(n607), .B(n608), .Z(\u_a23_mem/n19499 ) );
  NAND U971 ( .A(n603), .B(\u_a23_mem/stack_mem[19][1] ), .Z(n608) );
  AND U972 ( .A(n609), .B(n610), .Z(n607) );
  NANDN U973 ( .B(n537), .A(n110), .Z(n610) );
  OR U974 ( .A(n17), .B(n606), .Z(n609) );
  NAND U975 ( .A(n611), .B(n612), .Z(\u_a23_mem/n19498 ) );
  NAND U976 ( .A(n603), .B(\u_a23_mem/stack_mem[19][2] ), .Z(n612) );
  AND U977 ( .A(n613), .B(n614), .Z(n611) );
  NANDN U978 ( .B(n537), .A(n115), .Z(n614) );
  OR U979 ( .A(n23), .B(n606), .Z(n613) );
  NAND U980 ( .A(n615), .B(n616), .Z(\u_a23_mem/n19497 ) );
  NAND U981 ( .A(n603), .B(\u_a23_mem/stack_mem[19][3] ), .Z(n616) );
  AND U982 ( .A(n617), .B(n618), .Z(n615) );
  NANDN U983 ( .B(n537), .A(n120), .Z(n618) );
  OR U984 ( .A(n29), .B(n606), .Z(n617) );
  NAND U985 ( .A(n619), .B(n620), .Z(\u_a23_mem/n19496 ) );
  NAND U986 ( .A(n603), .B(\u_a23_mem/stack_mem[19][4] ), .Z(n620) );
  AND U987 ( .A(n621), .B(n622), .Z(n619) );
  NANDN U988 ( .B(n537), .A(n125), .Z(n622) );
  OR U989 ( .A(n35), .B(n606), .Z(n621) );
  NAND U990 ( .A(n623), .B(n624), .Z(\u_a23_mem/n19495 ) );
  NAND U991 ( .A(n603), .B(\u_a23_mem/stack_mem[19][5] ), .Z(n624) );
  AND U992 ( .A(n625), .B(n626), .Z(n623) );
  NANDN U993 ( .B(n537), .A(n130), .Z(n626) );
  OR U994 ( .A(n41), .B(n606), .Z(n625) );
  NAND U995 ( .A(n627), .B(n628), .Z(\u_a23_mem/n19494 ) );
  NAND U996 ( .A(n603), .B(\u_a23_mem/stack_mem[19][6] ), .Z(n628) );
  AND U997 ( .A(n629), .B(n630), .Z(n627) );
  NANDN U998 ( .B(n537), .A(n135), .Z(n630) );
  OR U999 ( .A(n47), .B(n606), .Z(n629) );
  NAND U1000 ( .A(n631), .B(n632), .Z(\u_a23_mem/n19493 ) );
  NAND U1001 ( .A(n603), .B(\u_a23_mem/stack_mem[19][7] ), .Z(n632) );
  NANDN U1002 ( .B(n138), .A(n531), .Z(n603) );
  AND U1003 ( .A(n633), .B(n634), .Z(n631) );
  NANDN U1004 ( .B(n537), .A(n142), .Z(n634) );
  NAND U1005 ( .A(n531), .B(n95), .Z(n537) );
  OR U1006 ( .A(n54), .B(n606), .Z(n633) );
  NAND U1007 ( .A(n635), .B(n636), .Z(\u_a23_mem/n19492 ) );
  OR U1008 ( .A(n11), .B(n637), .Z(n636) );
  NAND U1009 ( .A(n638), .B(\u_a23_mem/stack_mem[20][0] ), .Z(n635) );
  NAND U1010 ( .A(n639), .B(n640), .Z(\u_a23_mem/n19491 ) );
  OR U1011 ( .A(n17), .B(n637), .Z(n640) );
  NAND U1012 ( .A(n638), .B(\u_a23_mem/stack_mem[20][1] ), .Z(n639) );
  NAND U1013 ( .A(n641), .B(n642), .Z(\u_a23_mem/n19490 ) );
  OR U1014 ( .A(n23), .B(n637), .Z(n642) );
  NAND U1015 ( .A(n638), .B(\u_a23_mem/stack_mem[20][2] ), .Z(n641) );
  NAND U1016 ( .A(n643), .B(n644), .Z(\u_a23_mem/n19489 ) );
  OR U1017 ( .A(n29), .B(n637), .Z(n644) );
  NAND U1018 ( .A(n638), .B(\u_a23_mem/stack_mem[20][3] ), .Z(n643) );
  NAND U1019 ( .A(n645), .B(n646), .Z(\u_a23_mem/n19488 ) );
  OR U1020 ( .A(n35), .B(n637), .Z(n646) );
  NAND U1021 ( .A(n638), .B(\u_a23_mem/stack_mem[20][4] ), .Z(n645) );
  NAND U1022 ( .A(n647), .B(n648), .Z(\u_a23_mem/n19487 ) );
  OR U1023 ( .A(n41), .B(n637), .Z(n648) );
  NAND U1024 ( .A(n638), .B(\u_a23_mem/stack_mem[20][5] ), .Z(n647) );
  NAND U1025 ( .A(n649), .B(n650), .Z(\u_a23_mem/n19486 ) );
  OR U1026 ( .A(n47), .B(n637), .Z(n650) );
  NAND U1027 ( .A(n638), .B(\u_a23_mem/stack_mem[20][6] ), .Z(n649) );
  NAND U1028 ( .A(n651), .B(n652), .Z(\u_a23_mem/n19485 ) );
  OR U1029 ( .A(n54), .B(n637), .Z(n652) );
  NAND U1030 ( .A(n638), .B(\u_a23_mem/stack_mem[20][7] ), .Z(n651) );
  NANDN U1031 ( .B(n162), .A(n653), .Z(n638) );
  NAND U1032 ( .A(n654), .B(n655), .Z(\u_a23_mem/n19484 ) );
  NAND U1033 ( .A(n656), .B(\u_a23_mem/stack_mem[21][0] ), .Z(n655) );
  AND U1034 ( .A(n657), .B(n658), .Z(n654) );
  NANDN U1035 ( .B(n659), .A(n9), .Z(n658) );
  OR U1036 ( .A(n11), .B(n660), .Z(n657) );
  NAND U1037 ( .A(n661), .B(n662), .Z(\u_a23_mem/n19483 ) );
  NAND U1038 ( .A(n656), .B(\u_a23_mem/stack_mem[21][1] ), .Z(n662) );
  AND U1039 ( .A(n663), .B(n664), .Z(n661) );
  NANDN U1040 ( .B(n659), .A(n16), .Z(n664) );
  OR U1041 ( .A(n17), .B(n660), .Z(n663) );
  NAND U1042 ( .A(n665), .B(n666), .Z(\u_a23_mem/n19482 ) );
  NAND U1043 ( .A(n656), .B(\u_a23_mem/stack_mem[21][2] ), .Z(n666) );
  AND U1044 ( .A(n667), .B(n668), .Z(n665) );
  NANDN U1045 ( .B(n659), .A(n22), .Z(n668) );
  OR U1046 ( .A(n23), .B(n660), .Z(n667) );
  NAND U1047 ( .A(n669), .B(n670), .Z(\u_a23_mem/n19481 ) );
  NAND U1048 ( .A(n656), .B(\u_a23_mem/stack_mem[21][3] ), .Z(n670) );
  AND U1049 ( .A(n671), .B(n672), .Z(n669) );
  NANDN U1050 ( .B(n659), .A(n28), .Z(n672) );
  OR U1051 ( .A(n29), .B(n660), .Z(n671) );
  NAND U1052 ( .A(n673), .B(n674), .Z(\u_a23_mem/n19480 ) );
  NAND U1053 ( .A(n656), .B(\u_a23_mem/stack_mem[21][4] ), .Z(n674) );
  AND U1054 ( .A(n675), .B(n676), .Z(n673) );
  NANDN U1055 ( .B(n659), .A(n34), .Z(n676) );
  OR U1056 ( .A(n35), .B(n660), .Z(n675) );
  NAND U1057 ( .A(n677), .B(n678), .Z(\u_a23_mem/n19479 ) );
  NAND U1058 ( .A(n656), .B(\u_a23_mem/stack_mem[21][5] ), .Z(n678) );
  AND U1059 ( .A(n679), .B(n680), .Z(n677) );
  NANDN U1060 ( .B(n659), .A(n40), .Z(n680) );
  OR U1061 ( .A(n41), .B(n660), .Z(n679) );
  NAND U1062 ( .A(n681), .B(n682), .Z(\u_a23_mem/n19478 ) );
  NAND U1063 ( .A(n656), .B(\u_a23_mem/stack_mem[21][6] ), .Z(n682) );
  AND U1064 ( .A(n683), .B(n684), .Z(n681) );
  NANDN U1065 ( .B(n659), .A(n46), .Z(n684) );
  OR U1066 ( .A(n47), .B(n660), .Z(n683) );
  NAND U1067 ( .A(n685), .B(n686), .Z(\u_a23_mem/n19477 ) );
  NAND U1068 ( .A(n656), .B(\u_a23_mem/stack_mem[21][7] ), .Z(n686) );
  NANDN U1069 ( .B(n197), .A(n653), .Z(n656) );
  AND U1070 ( .A(n687), .B(n688), .Z(n685) );
  NANDN U1071 ( .B(n659), .A(n53), .Z(n688) );
  OR U1072 ( .A(n54), .B(n660), .Z(n687) );
  NAND U1073 ( .A(n689), .B(n690), .Z(\u_a23_mem/n19476 ) );
  NAND U1074 ( .A(n691), .B(\u_a23_mem/stack_mem[22][0] ), .Z(n690) );
  AND U1075 ( .A(n692), .B(n693), .Z(n689) );
  NANDN U1076 ( .B(n659), .A(n60), .Z(n693) );
  OR U1077 ( .A(n11), .B(n694), .Z(n692) );
  NAND U1078 ( .A(n695), .B(n696), .Z(\u_a23_mem/n19475 ) );
  NAND U1079 ( .A(n691), .B(\u_a23_mem/stack_mem[22][1] ), .Z(n696) );
  AND U1080 ( .A(n697), .B(n698), .Z(n695) );
  NANDN U1081 ( .B(n659), .A(n66), .Z(n698) );
  OR U1082 ( .A(n17), .B(n694), .Z(n697) );
  NAND U1083 ( .A(n699), .B(n700), .Z(\u_a23_mem/n19474 ) );
  NAND U1084 ( .A(n691), .B(\u_a23_mem/stack_mem[22][2] ), .Z(n700) );
  AND U1085 ( .A(n701), .B(n702), .Z(n699) );
  NANDN U1086 ( .B(n659), .A(n71), .Z(n702) );
  OR U1087 ( .A(n23), .B(n694), .Z(n701) );
  NAND U1088 ( .A(n703), .B(n704), .Z(\u_a23_mem/n19473 ) );
  NAND U1089 ( .A(n691), .B(\u_a23_mem/stack_mem[22][3] ), .Z(n704) );
  AND U1090 ( .A(n705), .B(n706), .Z(n703) );
  NANDN U1091 ( .B(n659), .A(n76), .Z(n706) );
  OR U1092 ( .A(n29), .B(n694), .Z(n705) );
  NAND U1093 ( .A(n707), .B(n708), .Z(\u_a23_mem/n19472 ) );
  NAND U1094 ( .A(n691), .B(\u_a23_mem/stack_mem[22][4] ), .Z(n708) );
  AND U1095 ( .A(n709), .B(n710), .Z(n707) );
  NANDN U1096 ( .B(n659), .A(n81), .Z(n710) );
  OR U1097 ( .A(n35), .B(n694), .Z(n709) );
  NAND U1098 ( .A(n711), .B(n712), .Z(\u_a23_mem/n19471 ) );
  NAND U1099 ( .A(n691), .B(\u_a23_mem/stack_mem[22][5] ), .Z(n712) );
  AND U1100 ( .A(n713), .B(n714), .Z(n711) );
  NANDN U1101 ( .B(n659), .A(n86), .Z(n714) );
  OR U1102 ( .A(n41), .B(n694), .Z(n713) );
  NAND U1103 ( .A(n715), .B(n716), .Z(\u_a23_mem/n19470 ) );
  NAND U1104 ( .A(n691), .B(\u_a23_mem/stack_mem[22][6] ), .Z(n716) );
  AND U1105 ( .A(n717), .B(n718), .Z(n715) );
  NANDN U1106 ( .B(n659), .A(n91), .Z(n718) );
  OR U1107 ( .A(n47), .B(n694), .Z(n717) );
  NAND U1108 ( .A(n719), .B(n720), .Z(\u_a23_mem/n19469 ) );
  NAND U1109 ( .A(n691), .B(\u_a23_mem/stack_mem[22][7] ), .Z(n720) );
  NANDN U1110 ( .B(n232), .A(n653), .Z(n691) );
  AND U1111 ( .A(n721), .B(n722), .Z(n719) );
  NANDN U1112 ( .B(n659), .A(n98), .Z(n722) );
  OR U1113 ( .A(n54), .B(n694), .Z(n721) );
  NAND U1114 ( .A(n723), .B(n724), .Z(\u_a23_mem/n19468 ) );
  NAND U1115 ( .A(n725), .B(\u_a23_mem/stack_mem[23][0] ), .Z(n724) );
  AND U1116 ( .A(n726), .B(n727), .Z(n723) );
  NANDN U1117 ( .B(n659), .A(n104), .Z(n727) );
  OR U1118 ( .A(n11), .B(n728), .Z(n726) );
  NAND U1119 ( .A(n729), .B(n730), .Z(\u_a23_mem/n19467 ) );
  NAND U1120 ( .A(n725), .B(\u_a23_mem/stack_mem[23][1] ), .Z(n730) );
  AND U1121 ( .A(n731), .B(n732), .Z(n729) );
  NANDN U1122 ( .B(n659), .A(n110), .Z(n732) );
  OR U1123 ( .A(n17), .B(n728), .Z(n731) );
  NAND U1124 ( .A(n733), .B(n734), .Z(\u_a23_mem/n19466 ) );
  NAND U1125 ( .A(n725), .B(\u_a23_mem/stack_mem[23][2] ), .Z(n734) );
  AND U1126 ( .A(n735), .B(n736), .Z(n733) );
  NANDN U1127 ( .B(n659), .A(n115), .Z(n736) );
  OR U1128 ( .A(n23), .B(n728), .Z(n735) );
  NAND U1129 ( .A(n737), .B(n738), .Z(\u_a23_mem/n19465 ) );
  NAND U1130 ( .A(n725), .B(\u_a23_mem/stack_mem[23][3] ), .Z(n738) );
  AND U1131 ( .A(n739), .B(n740), .Z(n737) );
  NANDN U1132 ( .B(n659), .A(n120), .Z(n740) );
  OR U1133 ( .A(n29), .B(n728), .Z(n739) );
  NAND U1134 ( .A(n741), .B(n742), .Z(\u_a23_mem/n19464 ) );
  NAND U1135 ( .A(n725), .B(\u_a23_mem/stack_mem[23][4] ), .Z(n742) );
  AND U1136 ( .A(n743), .B(n744), .Z(n741) );
  NANDN U1137 ( .B(n659), .A(n125), .Z(n744) );
  OR U1138 ( .A(n35), .B(n728), .Z(n743) );
  NAND U1139 ( .A(n745), .B(n746), .Z(\u_a23_mem/n19463 ) );
  NAND U1140 ( .A(n725), .B(\u_a23_mem/stack_mem[23][5] ), .Z(n746) );
  AND U1141 ( .A(n747), .B(n748), .Z(n745) );
  NANDN U1142 ( .B(n659), .A(n130), .Z(n748) );
  OR U1143 ( .A(n41), .B(n728), .Z(n747) );
  NAND U1144 ( .A(n749), .B(n750), .Z(\u_a23_mem/n19462 ) );
  NAND U1145 ( .A(n725), .B(\u_a23_mem/stack_mem[23][6] ), .Z(n750) );
  AND U1146 ( .A(n751), .B(n752), .Z(n749) );
  NANDN U1147 ( .B(n659), .A(n135), .Z(n752) );
  OR U1148 ( .A(n47), .B(n728), .Z(n751) );
  NAND U1149 ( .A(n753), .B(n754), .Z(\u_a23_mem/n19461 ) );
  NAND U1150 ( .A(n725), .B(\u_a23_mem/stack_mem[23][7] ), .Z(n754) );
  NANDN U1151 ( .B(n138), .A(n653), .Z(n725) );
  AND U1152 ( .A(n755), .B(n756), .Z(n753) );
  NANDN U1153 ( .B(n659), .A(n142), .Z(n756) );
  NAND U1154 ( .A(n653), .B(n95), .Z(n659) );
  OR U1155 ( .A(n54), .B(n728), .Z(n755) );
  NAND U1156 ( .A(n757), .B(n758), .Z(\u_a23_mem/n19460 ) );
  OR U1157 ( .A(n11), .B(n759), .Z(n758) );
  NAND U1158 ( .A(n760), .B(\u_a23_mem/stack_mem[24][0] ), .Z(n757) );
  NAND U1159 ( .A(n761), .B(n762), .Z(\u_a23_mem/n19459 ) );
  OR U1160 ( .A(n17), .B(n759), .Z(n762) );
  NAND U1161 ( .A(n760), .B(\u_a23_mem/stack_mem[24][1] ), .Z(n761) );
  NAND U1162 ( .A(n763), .B(n764), .Z(\u_a23_mem/n19458 ) );
  OR U1163 ( .A(n23), .B(n759), .Z(n764) );
  NAND U1164 ( .A(n760), .B(\u_a23_mem/stack_mem[24][2] ), .Z(n763) );
  NAND U1165 ( .A(n765), .B(n766), .Z(\u_a23_mem/n19457 ) );
  OR U1166 ( .A(n29), .B(n759), .Z(n766) );
  NAND U1167 ( .A(n760), .B(\u_a23_mem/stack_mem[24][3] ), .Z(n765) );
  NAND U1168 ( .A(n767), .B(n768), .Z(\u_a23_mem/n19456 ) );
  OR U1169 ( .A(n35), .B(n759), .Z(n768) );
  NAND U1170 ( .A(n760), .B(\u_a23_mem/stack_mem[24][4] ), .Z(n767) );
  NAND U1171 ( .A(n769), .B(n770), .Z(\u_a23_mem/n19455 ) );
  OR U1172 ( .A(n41), .B(n759), .Z(n770) );
  NAND U1173 ( .A(n760), .B(\u_a23_mem/stack_mem[24][5] ), .Z(n769) );
  NAND U1174 ( .A(n771), .B(n772), .Z(\u_a23_mem/n19454 ) );
  OR U1175 ( .A(n47), .B(n759), .Z(n772) );
  NAND U1176 ( .A(n760), .B(\u_a23_mem/stack_mem[24][6] ), .Z(n771) );
  NAND U1177 ( .A(n773), .B(n774), .Z(\u_a23_mem/n19453 ) );
  OR U1178 ( .A(n54), .B(n759), .Z(n774) );
  NAND U1179 ( .A(n760), .B(\u_a23_mem/stack_mem[24][7] ), .Z(n773) );
  OR U1180 ( .A(n162), .B(n775), .Z(n760) );
  NAND U1181 ( .A(n776), .B(n777), .Z(\u_a23_mem/n19452 ) );
  NAND U1182 ( .A(n778), .B(\u_a23_mem/stack_mem[25][0] ), .Z(n777) );
  AND U1183 ( .A(n779), .B(n780), .Z(n776) );
  NANDN U1184 ( .B(n781), .A(n9), .Z(n780) );
  OR U1185 ( .A(n11), .B(n782), .Z(n779) );
  NAND U1186 ( .A(n783), .B(n784), .Z(\u_a23_mem/n19451 ) );
  NAND U1187 ( .A(n778), .B(\u_a23_mem/stack_mem[25][1] ), .Z(n784) );
  AND U1188 ( .A(n785), .B(n786), .Z(n783) );
  NANDN U1189 ( .B(n781), .A(n16), .Z(n786) );
  OR U1190 ( .A(n17), .B(n782), .Z(n785) );
  NAND U1191 ( .A(n787), .B(n788), .Z(\u_a23_mem/n19450 ) );
  NAND U1192 ( .A(n778), .B(\u_a23_mem/stack_mem[25][2] ), .Z(n788) );
  AND U1193 ( .A(n789), .B(n790), .Z(n787) );
  NANDN U1194 ( .B(n781), .A(n22), .Z(n790) );
  OR U1195 ( .A(n23), .B(n782), .Z(n789) );
  NAND U1196 ( .A(n791), .B(n792), .Z(\u_a23_mem/n19449 ) );
  NAND U1197 ( .A(n778), .B(\u_a23_mem/stack_mem[25][3] ), .Z(n792) );
  AND U1198 ( .A(n793), .B(n794), .Z(n791) );
  NANDN U1199 ( .B(n781), .A(n28), .Z(n794) );
  OR U1200 ( .A(n29), .B(n782), .Z(n793) );
  NAND U1201 ( .A(n795), .B(n796), .Z(\u_a23_mem/n19448 ) );
  NAND U1202 ( .A(n778), .B(\u_a23_mem/stack_mem[25][4] ), .Z(n796) );
  AND U1203 ( .A(n797), .B(n798), .Z(n795) );
  NANDN U1204 ( .B(n781), .A(n34), .Z(n798) );
  OR U1205 ( .A(n35), .B(n782), .Z(n797) );
  NAND U1206 ( .A(n799), .B(n800), .Z(\u_a23_mem/n19447 ) );
  NAND U1207 ( .A(n778), .B(\u_a23_mem/stack_mem[25][5] ), .Z(n800) );
  AND U1208 ( .A(n801), .B(n802), .Z(n799) );
  NANDN U1209 ( .B(n781), .A(n40), .Z(n802) );
  OR U1210 ( .A(n41), .B(n782), .Z(n801) );
  NAND U1211 ( .A(n803), .B(n804), .Z(\u_a23_mem/n19446 ) );
  NAND U1212 ( .A(n778), .B(\u_a23_mem/stack_mem[25][6] ), .Z(n804) );
  AND U1213 ( .A(n805), .B(n806), .Z(n803) );
  NANDN U1214 ( .B(n781), .A(n46), .Z(n806) );
  OR U1215 ( .A(n47), .B(n782), .Z(n805) );
  NAND U1216 ( .A(n807), .B(n808), .Z(\u_a23_mem/n19445 ) );
  NAND U1217 ( .A(n778), .B(\u_a23_mem/stack_mem[25][7] ), .Z(n808) );
  OR U1218 ( .A(n197), .B(n775), .Z(n778) );
  AND U1219 ( .A(n809), .B(n810), .Z(n807) );
  NANDN U1220 ( .B(n781), .A(n53), .Z(n810) );
  OR U1221 ( .A(n54), .B(n782), .Z(n809) );
  NAND U1222 ( .A(n811), .B(n812), .Z(\u_a23_mem/n19444 ) );
  NAND U1223 ( .A(n813), .B(\u_a23_mem/stack_mem[26][0] ), .Z(n812) );
  AND U1224 ( .A(n814), .B(n815), .Z(n811) );
  NANDN U1225 ( .B(n781), .A(n60), .Z(n815) );
  OR U1226 ( .A(n11), .B(n816), .Z(n814) );
  NAND U1227 ( .A(n817), .B(n818), .Z(\u_a23_mem/n19443 ) );
  NAND U1228 ( .A(n813), .B(\u_a23_mem/stack_mem[26][1] ), .Z(n818) );
  AND U1229 ( .A(n819), .B(n820), .Z(n817) );
  NANDN U1230 ( .B(n781), .A(n66), .Z(n820) );
  OR U1231 ( .A(n17), .B(n816), .Z(n819) );
  NAND U1232 ( .A(n821), .B(n822), .Z(\u_a23_mem/n19442 ) );
  NAND U1233 ( .A(n813), .B(\u_a23_mem/stack_mem[26][2] ), .Z(n822) );
  AND U1234 ( .A(n823), .B(n824), .Z(n821) );
  NANDN U1235 ( .B(n781), .A(n71), .Z(n824) );
  OR U1236 ( .A(n23), .B(n816), .Z(n823) );
  NAND U1237 ( .A(n825), .B(n826), .Z(\u_a23_mem/n19441 ) );
  NAND U1238 ( .A(n813), .B(\u_a23_mem/stack_mem[26][3] ), .Z(n826) );
  AND U1239 ( .A(n827), .B(n828), .Z(n825) );
  NANDN U1240 ( .B(n781), .A(n76), .Z(n828) );
  OR U1241 ( .A(n29), .B(n816), .Z(n827) );
  NAND U1242 ( .A(n829), .B(n830), .Z(\u_a23_mem/n19440 ) );
  NAND U1243 ( .A(n813), .B(\u_a23_mem/stack_mem[26][4] ), .Z(n830) );
  AND U1244 ( .A(n831), .B(n832), .Z(n829) );
  NANDN U1245 ( .B(n781), .A(n81), .Z(n832) );
  OR U1246 ( .A(n35), .B(n816), .Z(n831) );
  NAND U1247 ( .A(n833), .B(n834), .Z(\u_a23_mem/n19439 ) );
  NAND U1248 ( .A(n813), .B(\u_a23_mem/stack_mem[26][5] ), .Z(n834) );
  AND U1249 ( .A(n835), .B(n836), .Z(n833) );
  NANDN U1250 ( .B(n781), .A(n86), .Z(n836) );
  OR U1251 ( .A(n41), .B(n816), .Z(n835) );
  NAND U1252 ( .A(n837), .B(n838), .Z(\u_a23_mem/n19438 ) );
  NAND U1253 ( .A(n813), .B(\u_a23_mem/stack_mem[26][6] ), .Z(n838) );
  AND U1254 ( .A(n839), .B(n840), .Z(n837) );
  NANDN U1255 ( .B(n781), .A(n91), .Z(n840) );
  OR U1256 ( .A(n47), .B(n816), .Z(n839) );
  NAND U1257 ( .A(n841), .B(n842), .Z(\u_a23_mem/n19437 ) );
  NAND U1258 ( .A(n813), .B(\u_a23_mem/stack_mem[26][7] ), .Z(n842) );
  OR U1259 ( .A(n232), .B(n775), .Z(n813) );
  AND U1260 ( .A(n843), .B(n844), .Z(n841) );
  NANDN U1261 ( .B(n781), .A(n98), .Z(n844) );
  OR U1262 ( .A(n54), .B(n816), .Z(n843) );
  NAND U1263 ( .A(n845), .B(n846), .Z(\u_a23_mem/n19436 ) );
  NAND U1264 ( .A(n847), .B(\u_a23_mem/stack_mem[27][0] ), .Z(n846) );
  AND U1265 ( .A(n848), .B(n849), .Z(n845) );
  NANDN U1266 ( .B(n781), .A(n104), .Z(n849) );
  OR U1267 ( .A(n11), .B(n850), .Z(n848) );
  NAND U1268 ( .A(n851), .B(n852), .Z(\u_a23_mem/n19435 ) );
  NAND U1269 ( .A(n847), .B(\u_a23_mem/stack_mem[27][1] ), .Z(n852) );
  AND U1270 ( .A(n853), .B(n854), .Z(n851) );
  NANDN U1271 ( .B(n781), .A(n110), .Z(n854) );
  OR U1272 ( .A(n17), .B(n850), .Z(n853) );
  NAND U1273 ( .A(n855), .B(n856), .Z(\u_a23_mem/n19434 ) );
  NAND U1274 ( .A(n847), .B(\u_a23_mem/stack_mem[27][2] ), .Z(n856) );
  AND U1275 ( .A(n857), .B(n858), .Z(n855) );
  NANDN U1276 ( .B(n781), .A(n115), .Z(n858) );
  OR U1277 ( .A(n23), .B(n850), .Z(n857) );
  NAND U1278 ( .A(n859), .B(n860), .Z(\u_a23_mem/n19433 ) );
  NAND U1279 ( .A(n847), .B(\u_a23_mem/stack_mem[27][3] ), .Z(n860) );
  AND U1280 ( .A(n861), .B(n862), .Z(n859) );
  NANDN U1281 ( .B(n781), .A(n120), .Z(n862) );
  OR U1282 ( .A(n29), .B(n850), .Z(n861) );
  NAND U1283 ( .A(n863), .B(n864), .Z(\u_a23_mem/n19432 ) );
  NAND U1284 ( .A(n847), .B(\u_a23_mem/stack_mem[27][4] ), .Z(n864) );
  AND U1285 ( .A(n865), .B(n866), .Z(n863) );
  NANDN U1286 ( .B(n781), .A(n125), .Z(n866) );
  OR U1287 ( .A(n35), .B(n850), .Z(n865) );
  NAND U1288 ( .A(n867), .B(n868), .Z(\u_a23_mem/n19431 ) );
  NAND U1289 ( .A(n847), .B(\u_a23_mem/stack_mem[27][5] ), .Z(n868) );
  AND U1290 ( .A(n869), .B(n870), .Z(n867) );
  NANDN U1291 ( .B(n781), .A(n130), .Z(n870) );
  OR U1292 ( .A(n41), .B(n850), .Z(n869) );
  NAND U1293 ( .A(n871), .B(n872), .Z(\u_a23_mem/n19430 ) );
  NAND U1294 ( .A(n847), .B(\u_a23_mem/stack_mem[27][6] ), .Z(n872) );
  AND U1295 ( .A(n873), .B(n874), .Z(n871) );
  NANDN U1296 ( .B(n781), .A(n135), .Z(n874) );
  OR U1297 ( .A(n47), .B(n850), .Z(n873) );
  NAND U1298 ( .A(n875), .B(n876), .Z(\u_a23_mem/n19429 ) );
  NAND U1299 ( .A(n847), .B(\u_a23_mem/stack_mem[27][7] ), .Z(n876) );
  OR U1300 ( .A(n138), .B(n775), .Z(n847) );
  AND U1301 ( .A(n877), .B(n878), .Z(n875) );
  NANDN U1302 ( .B(n781), .A(n142), .Z(n878) );
  NAND U1303 ( .A(n879), .B(n95), .Z(n781) );
  OR U1304 ( .A(n54), .B(n850), .Z(n877) );
  NAND U1305 ( .A(n880), .B(n881), .Z(\u_a23_mem/n19428 ) );
  OR U1306 ( .A(n11), .B(n882), .Z(n881) );
  NAND U1307 ( .A(n883), .B(\u_a23_mem/stack_mem[28][0] ), .Z(n880) );
  NAND U1308 ( .A(n884), .B(n885), .Z(\u_a23_mem/n19427 ) );
  OR U1309 ( .A(n17), .B(n882), .Z(n885) );
  NAND U1310 ( .A(n883), .B(\u_a23_mem/stack_mem[28][1] ), .Z(n884) );
  NAND U1311 ( .A(n886), .B(n887), .Z(\u_a23_mem/n19426 ) );
  OR U1312 ( .A(n23), .B(n882), .Z(n887) );
  NAND U1313 ( .A(n883), .B(\u_a23_mem/stack_mem[28][2] ), .Z(n886) );
  NAND U1314 ( .A(n888), .B(n889), .Z(\u_a23_mem/n19425 ) );
  OR U1315 ( .A(n29), .B(n882), .Z(n889) );
  NAND U1316 ( .A(n883), .B(\u_a23_mem/stack_mem[28][3] ), .Z(n888) );
  NAND U1317 ( .A(n890), .B(n891), .Z(\u_a23_mem/n19424 ) );
  OR U1318 ( .A(n35), .B(n882), .Z(n891) );
  NAND U1319 ( .A(n883), .B(\u_a23_mem/stack_mem[28][4] ), .Z(n890) );
  NAND U1320 ( .A(n892), .B(n893), .Z(\u_a23_mem/n19423 ) );
  OR U1321 ( .A(n41), .B(n882), .Z(n893) );
  NAND U1322 ( .A(n883), .B(\u_a23_mem/stack_mem[28][5] ), .Z(n892) );
  NAND U1323 ( .A(n894), .B(n895), .Z(\u_a23_mem/n19422 ) );
  OR U1324 ( .A(n47), .B(n882), .Z(n895) );
  NAND U1325 ( .A(n883), .B(\u_a23_mem/stack_mem[28][6] ), .Z(n894) );
  NAND U1326 ( .A(n896), .B(n897), .Z(\u_a23_mem/n19421 ) );
  OR U1327 ( .A(n54), .B(n882), .Z(n897) );
  NAND U1328 ( .A(n883), .B(\u_a23_mem/stack_mem[28][7] ), .Z(n896) );
  OR U1329 ( .A(n162), .B(n898), .Z(n883) );
  NAND U1330 ( .A(n95), .B(n899), .Z(n162) );
  NAND U1331 ( .A(n900), .B(n901), .Z(\u_a23_mem/n19420 ) );
  NAND U1332 ( .A(n902), .B(\u_a23_mem/stack_mem[29][0] ), .Z(n901) );
  AND U1333 ( .A(n903), .B(n904), .Z(n900) );
  NANDN U1334 ( .B(n905), .A(n9), .Z(n904) );
  OR U1335 ( .A(n11), .B(n906), .Z(n903) );
  NAND U1336 ( .A(n907), .B(n908), .Z(\u_a23_mem/n19419 ) );
  NAND U1337 ( .A(n902), .B(\u_a23_mem/stack_mem[29][1] ), .Z(n908) );
  AND U1338 ( .A(n909), .B(n910), .Z(n907) );
  NANDN U1339 ( .B(n905), .A(n16), .Z(n910) );
  OR U1340 ( .A(n17), .B(n906), .Z(n909) );
  NAND U1341 ( .A(n911), .B(n912), .Z(\u_a23_mem/n19418 ) );
  NAND U1342 ( .A(n902), .B(\u_a23_mem/stack_mem[29][2] ), .Z(n912) );
  AND U1343 ( .A(n913), .B(n914), .Z(n911) );
  NANDN U1344 ( .B(n905), .A(n22), .Z(n914) );
  OR U1345 ( .A(n23), .B(n906), .Z(n913) );
  NAND U1346 ( .A(n915), .B(n916), .Z(\u_a23_mem/n19417 ) );
  NAND U1347 ( .A(n902), .B(\u_a23_mem/stack_mem[29][3] ), .Z(n916) );
  AND U1348 ( .A(n917), .B(n918), .Z(n915) );
  NANDN U1349 ( .B(n905), .A(n28), .Z(n918) );
  OR U1350 ( .A(n29), .B(n906), .Z(n917) );
  NAND U1351 ( .A(n919), .B(n920), .Z(\u_a23_mem/n19416 ) );
  NAND U1352 ( .A(n902), .B(\u_a23_mem/stack_mem[29][4] ), .Z(n920) );
  AND U1353 ( .A(n921), .B(n922), .Z(n919) );
  NANDN U1354 ( .B(n905), .A(n34), .Z(n922) );
  OR U1355 ( .A(n35), .B(n906), .Z(n921) );
  NAND U1356 ( .A(n923), .B(n924), .Z(\u_a23_mem/n19415 ) );
  NAND U1357 ( .A(n902), .B(\u_a23_mem/stack_mem[29][5] ), .Z(n924) );
  AND U1358 ( .A(n925), .B(n926), .Z(n923) );
  NANDN U1359 ( .B(n905), .A(n40), .Z(n926) );
  OR U1360 ( .A(n41), .B(n906), .Z(n925) );
  NAND U1361 ( .A(n927), .B(n928), .Z(\u_a23_mem/n19414 ) );
  NAND U1362 ( .A(n902), .B(\u_a23_mem/stack_mem[29][6] ), .Z(n928) );
  AND U1363 ( .A(n929), .B(n930), .Z(n927) );
  NANDN U1364 ( .B(n905), .A(n46), .Z(n930) );
  OR U1365 ( .A(n47), .B(n906), .Z(n929) );
  NAND U1366 ( .A(n931), .B(n932), .Z(\u_a23_mem/n19413 ) );
  NAND U1367 ( .A(n902), .B(\u_a23_mem/stack_mem[29][7] ), .Z(n932) );
  OR U1368 ( .A(n197), .B(n898), .Z(n902) );
  NAND U1369 ( .A(n95), .B(n933), .Z(n197) );
  AND U1370 ( .A(n934), .B(n935), .Z(n931) );
  NANDN U1371 ( .B(n905), .A(n53), .Z(n935) );
  OR U1372 ( .A(n54), .B(n906), .Z(n934) );
  NAND U1373 ( .A(n936), .B(n937), .Z(\u_a23_mem/n19412 ) );
  NAND U1374 ( .A(n938), .B(\u_a23_mem/stack_mem[30][0] ), .Z(n937) );
  AND U1375 ( .A(n939), .B(n940), .Z(n936) );
  NANDN U1376 ( .B(n905), .A(n60), .Z(n940) );
  OR U1377 ( .A(n11), .B(n941), .Z(n939) );
  NAND U1378 ( .A(n942), .B(n943), .Z(\u_a23_mem/n19411 ) );
  NAND U1379 ( .A(n938), .B(\u_a23_mem/stack_mem[30][1] ), .Z(n943) );
  AND U1380 ( .A(n944), .B(n945), .Z(n942) );
  NANDN U1381 ( .B(n905), .A(n66), .Z(n945) );
  OR U1382 ( .A(n17), .B(n941), .Z(n944) );
  NAND U1383 ( .A(n946), .B(n947), .Z(\u_a23_mem/n19410 ) );
  NAND U1384 ( .A(n938), .B(\u_a23_mem/stack_mem[30][2] ), .Z(n947) );
  AND U1385 ( .A(n948), .B(n949), .Z(n946) );
  NANDN U1386 ( .B(n905), .A(n71), .Z(n949) );
  OR U1387 ( .A(n23), .B(n941), .Z(n948) );
  NAND U1388 ( .A(n950), .B(n951), .Z(\u_a23_mem/n19409 ) );
  NAND U1389 ( .A(n938), .B(\u_a23_mem/stack_mem[30][3] ), .Z(n951) );
  AND U1390 ( .A(n952), .B(n953), .Z(n950) );
  NANDN U1391 ( .B(n905), .A(n76), .Z(n953) );
  OR U1392 ( .A(n29), .B(n941), .Z(n952) );
  NAND U1393 ( .A(n954), .B(n955), .Z(\u_a23_mem/n19408 ) );
  NAND U1394 ( .A(n938), .B(\u_a23_mem/stack_mem[30][4] ), .Z(n955) );
  AND U1395 ( .A(n956), .B(n957), .Z(n954) );
  NANDN U1396 ( .B(n905), .A(n81), .Z(n957) );
  OR U1397 ( .A(n35), .B(n941), .Z(n956) );
  NAND U1398 ( .A(n958), .B(n959), .Z(\u_a23_mem/n19407 ) );
  NAND U1399 ( .A(n938), .B(\u_a23_mem/stack_mem[30][5] ), .Z(n959) );
  AND U1400 ( .A(n960), .B(n961), .Z(n958) );
  NANDN U1401 ( .B(n905), .A(n86), .Z(n961) );
  OR U1402 ( .A(n41), .B(n941), .Z(n960) );
  NAND U1403 ( .A(n962), .B(n963), .Z(\u_a23_mem/n19406 ) );
  NAND U1404 ( .A(n938), .B(\u_a23_mem/stack_mem[30][6] ), .Z(n963) );
  AND U1405 ( .A(n964), .B(n965), .Z(n962) );
  NANDN U1406 ( .B(n905), .A(n91), .Z(n965) );
  OR U1407 ( .A(n47), .B(n941), .Z(n964) );
  NAND U1408 ( .A(n966), .B(n967), .Z(\u_a23_mem/n19405 ) );
  NAND U1409 ( .A(n938), .B(\u_a23_mem/stack_mem[30][7] ), .Z(n967) );
  OR U1410 ( .A(n232), .B(n898), .Z(n938) );
  NAND U1411 ( .A(n95), .B(n968), .Z(n232) );
  AND U1412 ( .A(n969), .B(n970), .Z(n966) );
  NANDN U1413 ( .B(n905), .A(n98), .Z(n970) );
  OR U1414 ( .A(n54), .B(n941), .Z(n969) );
  NAND U1415 ( .A(n971), .B(n972), .Z(\u_a23_mem/n19404 ) );
  NAND U1416 ( .A(n973), .B(\u_a23_mem/stack_mem[31][0] ), .Z(n972) );
  AND U1417 ( .A(n974), .B(n975), .Z(n971) );
  NANDN U1418 ( .B(n905), .A(n104), .Z(n975) );
  NANDN U1419 ( .B(n11), .A(n976), .Z(n974) );
  NAND U1420 ( .A(n95), .B(m_write[0]), .Z(n11) );
  NAND U1421 ( .A(n977), .B(n978), .Z(\u_a23_mem/n19403 ) );
  NAND U1422 ( .A(n973), .B(\u_a23_mem/stack_mem[31][1] ), .Z(n978) );
  AND U1423 ( .A(n979), .B(n980), .Z(n977) );
  NANDN U1424 ( .B(n905), .A(n110), .Z(n980) );
  NANDN U1425 ( .B(n17), .A(n976), .Z(n979) );
  NAND U1426 ( .A(n95), .B(m_write[1]), .Z(n17) );
  NAND U1427 ( .A(n981), .B(n982), .Z(\u_a23_mem/n19402 ) );
  NAND U1428 ( .A(n973), .B(\u_a23_mem/stack_mem[31][2] ), .Z(n982) );
  AND U1429 ( .A(n983), .B(n984), .Z(n981) );
  NANDN U1430 ( .B(n905), .A(n115), .Z(n984) );
  NANDN U1431 ( .B(n23), .A(n976), .Z(n983) );
  NAND U1432 ( .A(n95), .B(m_write[2]), .Z(n23) );
  NAND U1433 ( .A(n985), .B(n986), .Z(\u_a23_mem/n19401 ) );
  NAND U1434 ( .A(n973), .B(\u_a23_mem/stack_mem[31][3] ), .Z(n986) );
  AND U1435 ( .A(n987), .B(n988), .Z(n985) );
  NANDN U1436 ( .B(n905), .A(n120), .Z(n988) );
  NANDN U1437 ( .B(n29), .A(n976), .Z(n987) );
  NAND U1438 ( .A(n95), .B(m_write[3]), .Z(n29) );
  NAND U1439 ( .A(n989), .B(n990), .Z(\u_a23_mem/n19400 ) );
  NAND U1440 ( .A(n973), .B(\u_a23_mem/stack_mem[31][4] ), .Z(n990) );
  AND U1441 ( .A(n991), .B(n992), .Z(n989) );
  NANDN U1442 ( .B(n905), .A(n125), .Z(n992) );
  NANDN U1443 ( .B(n35), .A(n976), .Z(n991) );
  NAND U1444 ( .A(n95), .B(m_write[4]), .Z(n35) );
  NAND U1445 ( .A(n993), .B(n994), .Z(\u_a23_mem/n19399 ) );
  NAND U1446 ( .A(n973), .B(\u_a23_mem/stack_mem[31][5] ), .Z(n994) );
  AND U1447 ( .A(n995), .B(n996), .Z(n993) );
  NANDN U1448 ( .B(n905), .A(n130), .Z(n996) );
  NANDN U1449 ( .B(n41), .A(n976), .Z(n995) );
  NAND U1450 ( .A(n95), .B(m_write[5]), .Z(n41) );
  NAND U1451 ( .A(n997), .B(n998), .Z(\u_a23_mem/n19398 ) );
  NAND U1452 ( .A(n973), .B(\u_a23_mem/stack_mem[31][6] ), .Z(n998) );
  AND U1453 ( .A(n999), .B(n1000), .Z(n997) );
  NANDN U1454 ( .B(n905), .A(n135), .Z(n1000) );
  NANDN U1455 ( .B(n47), .A(n976), .Z(n999) );
  NAND U1456 ( .A(n95), .B(m_write[6]), .Z(n47) );
  NAND U1457 ( .A(n1001), .B(n1002), .Z(\u_a23_mem/n19397 ) );
  NAND U1458 ( .A(n973), .B(\u_a23_mem/stack_mem[31][7] ), .Z(n1002) );
  OR U1459 ( .A(n138), .B(n898), .Z(n973) );
  NAND U1460 ( .A(n95), .B(n1003), .Z(n138) );
  AND U1461 ( .A(n1004), .B(n1005), .Z(n1001) );
  NANDN U1462 ( .B(n905), .A(n142), .Z(n1005) );
  NAND U1463 ( .A(n1006), .B(n95), .Z(n905) );
  NANDN U1464 ( .B(n54), .A(n976), .Z(n1004) );
  NAND U1465 ( .A(m_write[7]), .B(n95), .Z(n54) );
  AND U1466 ( .A(m_write_en), .B(n1007), .Z(n95) );
  NAND U1467 ( .A(n1008), .B(n1009), .Z(\u_a23_mem/n19396 ) );
  OR U1468 ( .A(n1010), .B(n1011), .Z(n1009) );
  AND U1469 ( .A(n1012), .B(n1013), .Z(n1008) );
  NAND U1470 ( .A(n1014), .B(\u_a23_mem/p_mem[3][0] ), .Z(n1013) );
  NANDN U1471 ( .B(n1015), .A(n1016), .Z(n1012) );
  NAND U1472 ( .A(n1017), .B(n1018), .Z(\u_a23_mem/n19395 ) );
  OR U1473 ( .A(n1010), .B(n1019), .Z(n1018) );
  AND U1474 ( .A(n1020), .B(n1021), .Z(n1017) );
  NAND U1475 ( .A(n1014), .B(\u_a23_mem/p_mem[3][1] ), .Z(n1021) );
  NANDN U1476 ( .B(n1022), .A(n1016), .Z(n1020) );
  NAND U1477 ( .A(n1023), .B(n1024), .Z(\u_a23_mem/n19394 ) );
  OR U1478 ( .A(n1010), .B(n1025), .Z(n1024) );
  AND U1479 ( .A(n1026), .B(n1027), .Z(n1023) );
  NAND U1480 ( .A(n1014), .B(\u_a23_mem/p_mem[3][2] ), .Z(n1027) );
  NANDN U1481 ( .B(n1028), .A(n1016), .Z(n1026) );
  NAND U1482 ( .A(n1029), .B(n1030), .Z(\u_a23_mem/n19393 ) );
  OR U1483 ( .A(n1010), .B(n1031), .Z(n1030) );
  AND U1484 ( .A(n1032), .B(n1033), .Z(n1029) );
  NAND U1485 ( .A(n1014), .B(\u_a23_mem/p_mem[3][3] ), .Z(n1033) );
  NANDN U1486 ( .B(n1034), .A(n1016), .Z(n1032) );
  NAND U1487 ( .A(n1035), .B(n1036), .Z(\u_a23_mem/n19392 ) );
  OR U1488 ( .A(n1010), .B(n1037), .Z(n1036) );
  AND U1489 ( .A(n1038), .B(n1039), .Z(n1035) );
  NAND U1490 ( .A(n1014), .B(\u_a23_mem/p_mem[3][4] ), .Z(n1039) );
  NANDN U1491 ( .B(n1040), .A(n1016), .Z(n1038) );
  NAND U1492 ( .A(n1041), .B(n1042), .Z(\u_a23_mem/n19391 ) );
  OR U1493 ( .A(n1010), .B(n1043), .Z(n1042) );
  AND U1494 ( .A(n1044), .B(n1045), .Z(n1041) );
  NAND U1495 ( .A(n1014), .B(\u_a23_mem/p_mem[3][5] ), .Z(n1045) );
  NANDN U1496 ( .B(n1046), .A(n1016), .Z(n1044) );
  NAND U1497 ( .A(n1047), .B(n1048), .Z(\u_a23_mem/n19390 ) );
  OR U1498 ( .A(n1049), .B(n1010), .Z(n1048) );
  AND U1499 ( .A(n1050), .B(n1051), .Z(n1047) );
  NAND U1500 ( .A(n1014), .B(\u_a23_mem/p_mem[3][6] ), .Z(n1051) );
  NANDN U1501 ( .B(n1052), .A(n1016), .Z(n1050) );
  NAND U1502 ( .A(n1053), .B(n1054), .Z(\u_a23_mem/n19389 ) );
  NANDN U1503 ( .B(n1010), .A(n1055), .Z(n1054) );
  NAND U1504 ( .A(n1016), .B(n1056), .Z(n1010) );
  AND U1505 ( .A(n1057), .B(n1058), .Z(n1053) );
  NAND U1506 ( .A(n1014), .B(\u_a23_mem/p_mem[3][7] ), .Z(n1058) );
  OR U1507 ( .A(n1059), .B(n1060), .Z(n1014) );
  IV U1508 ( .A(n1016), .Z(n1060) );
  NAND U1509 ( .A(n1016), .B(n1061), .Z(n1057) );
  NAND U1510 ( .A(n1062), .B(n1063), .Z(\u_a23_mem/n19388 ) );
  NAND U1511 ( .A(n1064), .B(\u_a23_mem/p_mem[4][0] ), .Z(n1063) );
  OR U1512 ( .A(n1011), .B(n1065), .Z(n1062) );
  NAND U1513 ( .A(n1066), .B(n1067), .Z(\u_a23_mem/n19387 ) );
  NAND U1514 ( .A(n1064), .B(\u_a23_mem/p_mem[4][1] ), .Z(n1067) );
  OR U1515 ( .A(n1019), .B(n1065), .Z(n1066) );
  NAND U1516 ( .A(n1068), .B(n1069), .Z(\u_a23_mem/n19386 ) );
  NAND U1517 ( .A(n1064), .B(\u_a23_mem/p_mem[4][2] ), .Z(n1069) );
  OR U1518 ( .A(n1025), .B(n1065), .Z(n1068) );
  NAND U1519 ( .A(n1070), .B(n1071), .Z(\u_a23_mem/n19385 ) );
  NAND U1520 ( .A(n1064), .B(\u_a23_mem/p_mem[4][3] ), .Z(n1071) );
  OR U1521 ( .A(n1031), .B(n1065), .Z(n1070) );
  NAND U1522 ( .A(n1072), .B(n1073), .Z(\u_a23_mem/n19384 ) );
  NAND U1523 ( .A(n1064), .B(\u_a23_mem/p_mem[4][4] ), .Z(n1073) );
  OR U1524 ( .A(n1037), .B(n1065), .Z(n1072) );
  NAND U1525 ( .A(n1074), .B(n1075), .Z(\u_a23_mem/n19383 ) );
  NAND U1526 ( .A(n1064), .B(\u_a23_mem/p_mem[4][5] ), .Z(n1075) );
  OR U1527 ( .A(n1043), .B(n1065), .Z(n1074) );
  NAND U1528 ( .A(n1076), .B(n1077), .Z(\u_a23_mem/n19382 ) );
  NAND U1529 ( .A(n1064), .B(\u_a23_mem/p_mem[4][6] ), .Z(n1077) );
  OR U1530 ( .A(n1049), .B(n1065), .Z(n1076) );
  NAND U1531 ( .A(n1078), .B(n1079), .Z(\u_a23_mem/n19381 ) );
  NAND U1532 ( .A(n1064), .B(\u_a23_mem/p_mem[4][7] ), .Z(n1079) );
  NANDN U1533 ( .B(n1080), .A(n1081), .Z(n1064) );
  NANDN U1534 ( .B(n1065), .A(n1055), .Z(n1078) );
  NANDN U1535 ( .B(n2), .A(n1081), .Z(n1065) );
  NAND U1536 ( .A(n1082), .B(n1083), .Z(\u_a23_mem/n19380 ) );
  OR U1537 ( .A(n1011), .B(n1084), .Z(n1083) );
  AND U1538 ( .A(n1085), .B(n1086), .Z(n1082) );
  NANDN U1539 ( .B(n1087), .A(n1081), .Z(n1086) );
  NAND U1540 ( .A(n1088), .B(\u_a23_mem/p_mem[5][0] ), .Z(n1085) );
  NAND U1541 ( .A(n1089), .B(n1090), .Z(\u_a23_mem/n19379 ) );
  OR U1542 ( .A(n1019), .B(n1084), .Z(n1090) );
  AND U1543 ( .A(n1091), .B(n1092), .Z(n1089) );
  NANDN U1544 ( .B(n1093), .A(n1081), .Z(n1092) );
  NAND U1545 ( .A(n1088), .B(\u_a23_mem/p_mem[5][1] ), .Z(n1091) );
  NAND U1546 ( .A(n1094), .B(n1095), .Z(\u_a23_mem/n19378 ) );
  OR U1547 ( .A(n1025), .B(n1084), .Z(n1095) );
  AND U1548 ( .A(n1096), .B(n1097), .Z(n1094) );
  NANDN U1549 ( .B(n1098), .A(n1081), .Z(n1097) );
  NAND U1550 ( .A(n1088), .B(\u_a23_mem/p_mem[5][2] ), .Z(n1096) );
  NAND U1551 ( .A(n1099), .B(n1100), .Z(\u_a23_mem/n19377 ) );
  OR U1552 ( .A(n1031), .B(n1084), .Z(n1100) );
  AND U1553 ( .A(n1101), .B(n1102), .Z(n1099) );
  NANDN U1554 ( .B(n1103), .A(n1081), .Z(n1102) );
  NAND U1555 ( .A(n1088), .B(\u_a23_mem/p_mem[5][3] ), .Z(n1101) );
  NAND U1556 ( .A(n1104), .B(n1105), .Z(\u_a23_mem/n19376 ) );
  OR U1557 ( .A(n1037), .B(n1084), .Z(n1105) );
  AND U1558 ( .A(n1106), .B(n1107), .Z(n1104) );
  NANDN U1559 ( .B(n1108), .A(n1081), .Z(n1107) );
  NAND U1560 ( .A(n1088), .B(\u_a23_mem/p_mem[5][4] ), .Z(n1106) );
  NAND U1561 ( .A(n1109), .B(n1110), .Z(\u_a23_mem/n19375 ) );
  OR U1562 ( .A(n1043), .B(n1084), .Z(n1110) );
  AND U1563 ( .A(n1111), .B(n1112), .Z(n1109) );
  NANDN U1564 ( .B(n1113), .A(n1081), .Z(n1112) );
  NAND U1565 ( .A(n1088), .B(\u_a23_mem/p_mem[5][5] ), .Z(n1111) );
  NAND U1566 ( .A(n1114), .B(n1115), .Z(\u_a23_mem/n19374 ) );
  OR U1567 ( .A(n1049), .B(n1084), .Z(n1115) );
  AND U1568 ( .A(n1116), .B(n1117), .Z(n1114) );
  NANDN U1569 ( .B(n1118), .A(n1081), .Z(n1117) );
  NAND U1570 ( .A(n1088), .B(\u_a23_mem/p_mem[5][6] ), .Z(n1116) );
  NAND U1571 ( .A(n1119), .B(n1120), .Z(\u_a23_mem/n19373 ) );
  NANDN U1572 ( .B(n1084), .A(n1055), .Z(n1120) );
  NAND U1573 ( .A(n1121), .B(n1081), .Z(n1084) );
  AND U1574 ( .A(n1122), .B(n1123), .Z(n1119) );
  NANDN U1575 ( .B(n1124), .A(n1081), .Z(n1123) );
  NAND U1576 ( .A(n1088), .B(\u_a23_mem/p_mem[5][7] ), .Z(n1122) );
  NANDN U1577 ( .B(n1125), .A(n1081), .Z(n1088) );
  NAND U1578 ( .A(n1126), .B(n1127), .Z(\u_a23_mem/n19372 ) );
  OR U1579 ( .A(n1011), .B(n1128), .Z(n1127) );
  AND U1580 ( .A(n1129), .B(n1130), .Z(n1126) );
  NANDN U1581 ( .B(n1131), .A(n1081), .Z(n1130) );
  NAND U1582 ( .A(n1132), .B(\u_a23_mem/p_mem[6][0] ), .Z(n1129) );
  NAND U1583 ( .A(n1133), .B(n1134), .Z(\u_a23_mem/n19371 ) );
  OR U1584 ( .A(n1019), .B(n1128), .Z(n1134) );
  AND U1585 ( .A(n1135), .B(n1136), .Z(n1133) );
  NANDN U1586 ( .B(n1137), .A(n1081), .Z(n1136) );
  NAND U1587 ( .A(n1132), .B(\u_a23_mem/p_mem[6][1] ), .Z(n1135) );
  NAND U1588 ( .A(n1138), .B(n1139), .Z(\u_a23_mem/n19370 ) );
  OR U1589 ( .A(n1025), .B(n1128), .Z(n1139) );
  AND U1590 ( .A(n1140), .B(n1141), .Z(n1138) );
  NANDN U1591 ( .B(n1142), .A(n1081), .Z(n1141) );
  NAND U1592 ( .A(n1132), .B(\u_a23_mem/p_mem[6][2] ), .Z(n1140) );
  NAND U1593 ( .A(n1143), .B(n1144), .Z(\u_a23_mem/n19369 ) );
  OR U1594 ( .A(n1031), .B(n1128), .Z(n1144) );
  AND U1595 ( .A(n1145), .B(n1146), .Z(n1143) );
  NANDN U1596 ( .B(n1147), .A(n1081), .Z(n1146) );
  NAND U1597 ( .A(n1132), .B(\u_a23_mem/p_mem[6][3] ), .Z(n1145) );
  NAND U1598 ( .A(n1148), .B(n1149), .Z(\u_a23_mem/n19368 ) );
  OR U1599 ( .A(n1037), .B(n1128), .Z(n1149) );
  AND U1600 ( .A(n1150), .B(n1151), .Z(n1148) );
  NANDN U1601 ( .B(n1152), .A(n1081), .Z(n1151) );
  NAND U1602 ( .A(n1132), .B(\u_a23_mem/p_mem[6][4] ), .Z(n1150) );
  NAND U1603 ( .A(n1153), .B(n1154), .Z(\u_a23_mem/n19367 ) );
  OR U1604 ( .A(n1043), .B(n1128), .Z(n1154) );
  AND U1605 ( .A(n1155), .B(n1156), .Z(n1153) );
  NANDN U1606 ( .B(n1157), .A(n1081), .Z(n1156) );
  NAND U1607 ( .A(n1132), .B(\u_a23_mem/p_mem[6][5] ), .Z(n1155) );
  NAND U1608 ( .A(n1158), .B(n1159), .Z(\u_a23_mem/n19366 ) );
  OR U1609 ( .A(n1049), .B(n1128), .Z(n1159) );
  AND U1610 ( .A(n1160), .B(n1161), .Z(n1158) );
  NANDN U1611 ( .B(n1162), .A(n1081), .Z(n1161) );
  NAND U1612 ( .A(n1132), .B(\u_a23_mem/p_mem[6][6] ), .Z(n1160) );
  NAND U1613 ( .A(n1163), .B(n1164), .Z(\u_a23_mem/n19365 ) );
  NANDN U1614 ( .B(n1128), .A(n1055), .Z(n1164) );
  NAND U1615 ( .A(n1165), .B(n1081), .Z(n1128) );
  AND U1616 ( .A(n1166), .B(n1167), .Z(n1163) );
  NANDN U1617 ( .B(n1168), .A(n1081), .Z(n1167) );
  NAND U1618 ( .A(n1132), .B(\u_a23_mem/p_mem[6][7] ), .Z(n1166) );
  NANDN U1619 ( .B(n1169), .A(n1081), .Z(n1132) );
  NAND U1620 ( .A(n1170), .B(n1171), .Z(\u_a23_mem/n19364 ) );
  OR U1621 ( .A(n1011), .B(n1172), .Z(n1171) );
  AND U1622 ( .A(n1173), .B(n1174), .Z(n1170) );
  NAND U1623 ( .A(n1175), .B(\u_a23_mem/p_mem[7][0] ), .Z(n1174) );
  NANDN U1624 ( .B(n1015), .A(n1081), .Z(n1173) );
  NAND U1625 ( .A(n1176), .B(n1177), .Z(\u_a23_mem/n19363 ) );
  OR U1626 ( .A(n1019), .B(n1172), .Z(n1177) );
  AND U1627 ( .A(n1178), .B(n1179), .Z(n1176) );
  NAND U1628 ( .A(n1175), .B(\u_a23_mem/p_mem[7][1] ), .Z(n1179) );
  NANDN U1629 ( .B(n1022), .A(n1081), .Z(n1178) );
  NAND U1630 ( .A(n1180), .B(n1181), .Z(\u_a23_mem/n19362 ) );
  OR U1631 ( .A(n1025), .B(n1172), .Z(n1181) );
  AND U1632 ( .A(n1182), .B(n1183), .Z(n1180) );
  NAND U1633 ( .A(n1175), .B(\u_a23_mem/p_mem[7][2] ), .Z(n1183) );
  NANDN U1634 ( .B(n1028), .A(n1081), .Z(n1182) );
  NAND U1635 ( .A(n1184), .B(n1185), .Z(\u_a23_mem/n19361 ) );
  OR U1636 ( .A(n1031), .B(n1172), .Z(n1185) );
  AND U1637 ( .A(n1186), .B(n1187), .Z(n1184) );
  NAND U1638 ( .A(n1175), .B(\u_a23_mem/p_mem[7][3] ), .Z(n1187) );
  NANDN U1639 ( .B(n1034), .A(n1081), .Z(n1186) );
  NAND U1640 ( .A(n1188), .B(n1189), .Z(\u_a23_mem/n19360 ) );
  OR U1641 ( .A(n1037), .B(n1172), .Z(n1189) );
  AND U1642 ( .A(n1190), .B(n1191), .Z(n1188) );
  NAND U1643 ( .A(n1175), .B(\u_a23_mem/p_mem[7][4] ), .Z(n1191) );
  NANDN U1644 ( .B(n1040), .A(n1081), .Z(n1190) );
  NAND U1645 ( .A(n1192), .B(n1193), .Z(\u_a23_mem/n19359 ) );
  OR U1646 ( .A(n1043), .B(n1172), .Z(n1193) );
  AND U1647 ( .A(n1194), .B(n1195), .Z(n1192) );
  NAND U1648 ( .A(n1175), .B(\u_a23_mem/p_mem[7][5] ), .Z(n1195) );
  NANDN U1649 ( .B(n1046), .A(n1081), .Z(n1194) );
  NAND U1650 ( .A(n1196), .B(n1197), .Z(\u_a23_mem/n19358 ) );
  OR U1651 ( .A(n1049), .B(n1172), .Z(n1197) );
  AND U1652 ( .A(n1198), .B(n1199), .Z(n1196) );
  NAND U1653 ( .A(n1175), .B(\u_a23_mem/p_mem[7][6] ), .Z(n1199) );
  NANDN U1654 ( .B(n1052), .A(n1081), .Z(n1198) );
  NAND U1655 ( .A(n1200), .B(n1201), .Z(\u_a23_mem/n19357 ) );
  NANDN U1656 ( .B(n1172), .A(n1055), .Z(n1201) );
  NAND U1657 ( .A(n1056), .B(n1081), .Z(n1172) );
  AND U1658 ( .A(n1202), .B(n1203), .Z(n1200) );
  NAND U1659 ( .A(n1175), .B(\u_a23_mem/p_mem[7][7] ), .Z(n1203) );
  NANDN U1660 ( .B(n1059), .A(n1081), .Z(n1175) );
  NAND U1661 ( .A(n1061), .B(n1081), .Z(n1202) );
  ANDN U1662 ( .A(n1204), .B(n1205), .Z(n1081) );
  NAND U1663 ( .A(n1206), .B(n1207), .Z(\u_a23_mem/n19356 ) );
  NAND U1664 ( .A(n1208), .B(\u_a23_mem/p_mem[8][0] ), .Z(n1207) );
  OR U1665 ( .A(n1011), .B(n1209), .Z(n1206) );
  NAND U1666 ( .A(n1210), .B(n1211), .Z(\u_a23_mem/n19355 ) );
  NAND U1667 ( .A(n1208), .B(\u_a23_mem/p_mem[8][1] ), .Z(n1211) );
  OR U1668 ( .A(n1019), .B(n1209), .Z(n1210) );
  NAND U1669 ( .A(n1212), .B(n1213), .Z(\u_a23_mem/n19354 ) );
  NAND U1670 ( .A(n1208), .B(\u_a23_mem/p_mem[8][2] ), .Z(n1213) );
  OR U1671 ( .A(n1025), .B(n1209), .Z(n1212) );
  NAND U1672 ( .A(n1214), .B(n1215), .Z(\u_a23_mem/n19353 ) );
  NAND U1673 ( .A(n1208), .B(\u_a23_mem/p_mem[8][3] ), .Z(n1215) );
  OR U1674 ( .A(n1031), .B(n1209), .Z(n1214) );
  NAND U1675 ( .A(n1216), .B(n1217), .Z(\u_a23_mem/n19352 ) );
  NAND U1676 ( .A(n1208), .B(\u_a23_mem/p_mem[8][4] ), .Z(n1217) );
  OR U1677 ( .A(n1037), .B(n1209), .Z(n1216) );
  NAND U1678 ( .A(n1218), .B(n1219), .Z(\u_a23_mem/n19351 ) );
  NAND U1679 ( .A(n1208), .B(\u_a23_mem/p_mem[8][5] ), .Z(n1219) );
  OR U1680 ( .A(n1043), .B(n1209), .Z(n1218) );
  NAND U1681 ( .A(n1220), .B(n1221), .Z(\u_a23_mem/n19350 ) );
  NAND U1682 ( .A(n1208), .B(\u_a23_mem/p_mem[8][6] ), .Z(n1221) );
  OR U1683 ( .A(n1049), .B(n1209), .Z(n1220) );
  NAND U1684 ( .A(n1222), .B(n1223), .Z(\u_a23_mem/n19349 ) );
  NAND U1685 ( .A(n1208), .B(\u_a23_mem/p_mem[8][7] ), .Z(n1223) );
  NANDN U1686 ( .B(n1080), .A(n1224), .Z(n1208) );
  NANDN U1687 ( .B(n1209), .A(n1055), .Z(n1222) );
  NANDN U1688 ( .B(n2), .A(n1224), .Z(n1209) );
  NAND U1689 ( .A(n1225), .B(n1226), .Z(\u_a23_mem/n19348 ) );
  OR U1690 ( .A(n1011), .B(n1227), .Z(n1226) );
  AND U1691 ( .A(n1228), .B(n1229), .Z(n1225) );
  NANDN U1692 ( .B(n1087), .A(n1224), .Z(n1229) );
  NAND U1693 ( .A(n1230), .B(\u_a23_mem/p_mem[9][0] ), .Z(n1228) );
  NAND U1694 ( .A(n1231), .B(n1232), .Z(\u_a23_mem/n19347 ) );
  OR U1695 ( .A(n1019), .B(n1227), .Z(n1232) );
  AND U1696 ( .A(n1233), .B(n1234), .Z(n1231) );
  NANDN U1697 ( .B(n1093), .A(n1224), .Z(n1234) );
  NAND U1698 ( .A(n1230), .B(\u_a23_mem/p_mem[9][1] ), .Z(n1233) );
  NAND U1699 ( .A(n1235), .B(n1236), .Z(\u_a23_mem/n19346 ) );
  OR U1700 ( .A(n1025), .B(n1227), .Z(n1236) );
  AND U1701 ( .A(n1237), .B(n1238), .Z(n1235) );
  NANDN U1702 ( .B(n1098), .A(n1224), .Z(n1238) );
  NAND U1703 ( .A(n1230), .B(\u_a23_mem/p_mem[9][2] ), .Z(n1237) );
  NAND U1704 ( .A(n1239), .B(n1240), .Z(\u_a23_mem/n19345 ) );
  OR U1705 ( .A(n1031), .B(n1227), .Z(n1240) );
  AND U1706 ( .A(n1241), .B(n1242), .Z(n1239) );
  NANDN U1707 ( .B(n1103), .A(n1224), .Z(n1242) );
  NAND U1708 ( .A(n1230), .B(\u_a23_mem/p_mem[9][3] ), .Z(n1241) );
  NAND U1709 ( .A(n1243), .B(n1244), .Z(\u_a23_mem/n19344 ) );
  OR U1710 ( .A(n1037), .B(n1227), .Z(n1244) );
  AND U1711 ( .A(n1245), .B(n1246), .Z(n1243) );
  NANDN U1712 ( .B(n1108), .A(n1224), .Z(n1246) );
  NAND U1713 ( .A(n1230), .B(\u_a23_mem/p_mem[9][4] ), .Z(n1245) );
  NAND U1714 ( .A(n1247), .B(n1248), .Z(\u_a23_mem/n19343 ) );
  OR U1715 ( .A(n1043), .B(n1227), .Z(n1248) );
  AND U1716 ( .A(n1249), .B(n1250), .Z(n1247) );
  NANDN U1717 ( .B(n1113), .A(n1224), .Z(n1250) );
  NAND U1718 ( .A(n1230), .B(\u_a23_mem/p_mem[9][5] ), .Z(n1249) );
  NAND U1719 ( .A(n1251), .B(n1252), .Z(\u_a23_mem/n19342 ) );
  OR U1720 ( .A(n1049), .B(n1227), .Z(n1252) );
  AND U1721 ( .A(n1253), .B(n1254), .Z(n1251) );
  NANDN U1722 ( .B(n1118), .A(n1224), .Z(n1254) );
  NAND U1723 ( .A(n1230), .B(\u_a23_mem/p_mem[9][6] ), .Z(n1253) );
  NAND U1724 ( .A(n1255), .B(n1256), .Z(\u_a23_mem/n19341 ) );
  NANDN U1725 ( .B(n1227), .A(n1055), .Z(n1256) );
  NAND U1726 ( .A(n1121), .B(n1224), .Z(n1227) );
  AND U1727 ( .A(n1257), .B(n1258), .Z(n1255) );
  NANDN U1728 ( .B(n1124), .A(n1224), .Z(n1258) );
  NAND U1729 ( .A(n1230), .B(\u_a23_mem/p_mem[9][7] ), .Z(n1257) );
  NANDN U1730 ( .B(n1125), .A(n1224), .Z(n1230) );
  NAND U1731 ( .A(n1259), .B(n1260), .Z(\u_a23_mem/n19340 ) );
  OR U1732 ( .A(n1011), .B(n1261), .Z(n1260) );
  AND U1733 ( .A(n1262), .B(n1263), .Z(n1259) );
  NANDN U1734 ( .B(n1131), .A(n1224), .Z(n1263) );
  NAND U1735 ( .A(n1264), .B(\u_a23_mem/p_mem[10][0] ), .Z(n1262) );
  NAND U1736 ( .A(n1265), .B(n1266), .Z(\u_a23_mem/n19339 ) );
  OR U1737 ( .A(n1019), .B(n1261), .Z(n1266) );
  AND U1738 ( .A(n1267), .B(n1268), .Z(n1265) );
  NANDN U1739 ( .B(n1137), .A(n1224), .Z(n1268) );
  NAND U1740 ( .A(n1264), .B(\u_a23_mem/p_mem[10][1] ), .Z(n1267) );
  NAND U1741 ( .A(n1269), .B(n1270), .Z(\u_a23_mem/n19338 ) );
  OR U1742 ( .A(n1025), .B(n1261), .Z(n1270) );
  AND U1743 ( .A(n1271), .B(n1272), .Z(n1269) );
  NANDN U1744 ( .B(n1142), .A(n1224), .Z(n1272) );
  NAND U1745 ( .A(n1264), .B(\u_a23_mem/p_mem[10][2] ), .Z(n1271) );
  NAND U1746 ( .A(n1273), .B(n1274), .Z(\u_a23_mem/n19337 ) );
  OR U1747 ( .A(n1031), .B(n1261), .Z(n1274) );
  AND U1748 ( .A(n1275), .B(n1276), .Z(n1273) );
  NANDN U1749 ( .B(n1147), .A(n1224), .Z(n1276) );
  NAND U1750 ( .A(n1264), .B(\u_a23_mem/p_mem[10][3] ), .Z(n1275) );
  NAND U1751 ( .A(n1277), .B(n1278), .Z(\u_a23_mem/n19336 ) );
  OR U1752 ( .A(n1037), .B(n1261), .Z(n1278) );
  AND U1753 ( .A(n1279), .B(n1280), .Z(n1277) );
  NANDN U1754 ( .B(n1152), .A(n1224), .Z(n1280) );
  NAND U1755 ( .A(n1264), .B(\u_a23_mem/p_mem[10][4] ), .Z(n1279) );
  NAND U1756 ( .A(n1281), .B(n1282), .Z(\u_a23_mem/n19335 ) );
  OR U1757 ( .A(n1043), .B(n1261), .Z(n1282) );
  AND U1758 ( .A(n1283), .B(n1284), .Z(n1281) );
  NANDN U1759 ( .B(n1157), .A(n1224), .Z(n1284) );
  NAND U1760 ( .A(n1264), .B(\u_a23_mem/p_mem[10][5] ), .Z(n1283) );
  NAND U1761 ( .A(n1285), .B(n1286), .Z(\u_a23_mem/n19334 ) );
  OR U1762 ( .A(n1049), .B(n1261), .Z(n1286) );
  AND U1763 ( .A(n1287), .B(n1288), .Z(n1285) );
  NANDN U1764 ( .B(n1162), .A(n1224), .Z(n1288) );
  NAND U1765 ( .A(n1264), .B(\u_a23_mem/p_mem[10][6] ), .Z(n1287) );
  NAND U1766 ( .A(n1289), .B(n1290), .Z(\u_a23_mem/n19333 ) );
  NANDN U1767 ( .B(n1261), .A(n1055), .Z(n1290) );
  NAND U1768 ( .A(n1165), .B(n1224), .Z(n1261) );
  AND U1769 ( .A(n1291), .B(n1292), .Z(n1289) );
  NANDN U1770 ( .B(n1168), .A(n1224), .Z(n1292) );
  NAND U1771 ( .A(n1264), .B(\u_a23_mem/p_mem[10][7] ), .Z(n1291) );
  NANDN U1772 ( .B(n1169), .A(n1224), .Z(n1264) );
  NAND U1773 ( .A(n1293), .B(n1294), .Z(\u_a23_mem/n19332 ) );
  OR U1774 ( .A(n1011), .B(n1295), .Z(n1294) );
  AND U1775 ( .A(n1296), .B(n1297), .Z(n1293) );
  NAND U1776 ( .A(n1298), .B(\u_a23_mem/p_mem[11][0] ), .Z(n1297) );
  NANDN U1777 ( .B(n1015), .A(n1224), .Z(n1296) );
  NAND U1778 ( .A(n1299), .B(n1300), .Z(\u_a23_mem/n19331 ) );
  OR U1779 ( .A(n1019), .B(n1295), .Z(n1300) );
  AND U1780 ( .A(n1301), .B(n1302), .Z(n1299) );
  NAND U1781 ( .A(n1298), .B(\u_a23_mem/p_mem[11][1] ), .Z(n1302) );
  NANDN U1782 ( .B(n1022), .A(n1224), .Z(n1301) );
  NAND U1783 ( .A(n1303), .B(n1304), .Z(\u_a23_mem/n19330 ) );
  OR U1784 ( .A(n1025), .B(n1295), .Z(n1304) );
  AND U1785 ( .A(n1305), .B(n1306), .Z(n1303) );
  NAND U1786 ( .A(n1298), .B(\u_a23_mem/p_mem[11][2] ), .Z(n1306) );
  NANDN U1787 ( .B(n1028), .A(n1224), .Z(n1305) );
  NAND U1788 ( .A(n1307), .B(n1308), .Z(\u_a23_mem/n19329 ) );
  OR U1789 ( .A(n1031), .B(n1295), .Z(n1308) );
  AND U1790 ( .A(n1309), .B(n1310), .Z(n1307) );
  NAND U1791 ( .A(n1298), .B(\u_a23_mem/p_mem[11][3] ), .Z(n1310) );
  NANDN U1792 ( .B(n1034), .A(n1224), .Z(n1309) );
  NAND U1793 ( .A(n1311), .B(n1312), .Z(\u_a23_mem/n19328 ) );
  OR U1794 ( .A(n1037), .B(n1295), .Z(n1312) );
  AND U1795 ( .A(n1313), .B(n1314), .Z(n1311) );
  NAND U1796 ( .A(n1298), .B(\u_a23_mem/p_mem[11][4] ), .Z(n1314) );
  NANDN U1797 ( .B(n1040), .A(n1224), .Z(n1313) );
  NAND U1798 ( .A(n1315), .B(n1316), .Z(\u_a23_mem/n19327 ) );
  OR U1799 ( .A(n1043), .B(n1295), .Z(n1316) );
  AND U1800 ( .A(n1317), .B(n1318), .Z(n1315) );
  NAND U1801 ( .A(n1298), .B(\u_a23_mem/p_mem[11][5] ), .Z(n1318) );
  NANDN U1802 ( .B(n1046), .A(n1224), .Z(n1317) );
  NAND U1803 ( .A(n1319), .B(n1320), .Z(\u_a23_mem/n19326 ) );
  OR U1804 ( .A(n1049), .B(n1295), .Z(n1320) );
  AND U1805 ( .A(n1321), .B(n1322), .Z(n1319) );
  NAND U1806 ( .A(n1298), .B(\u_a23_mem/p_mem[11][6] ), .Z(n1322) );
  NANDN U1807 ( .B(n1052), .A(n1224), .Z(n1321) );
  NAND U1808 ( .A(n1323), .B(n1324), .Z(\u_a23_mem/n19325 ) );
  NANDN U1809 ( .B(n1295), .A(n1055), .Z(n1324) );
  NAND U1810 ( .A(n1056), .B(n1224), .Z(n1295) );
  AND U1811 ( .A(n1325), .B(n1326), .Z(n1323) );
  NAND U1812 ( .A(n1298), .B(\u_a23_mem/p_mem[11][7] ), .Z(n1326) );
  NANDN U1813 ( .B(n1059), .A(n1224), .Z(n1298) );
  NAND U1814 ( .A(n1061), .B(n1224), .Z(n1325) );
  ANDN U1815 ( .A(n1327), .B(n1205), .Z(n1224) );
  NAND U1816 ( .A(n1328), .B(n1329), .Z(\u_a23_mem/n19324 ) );
  NAND U1817 ( .A(n1330), .B(\u_a23_mem/p_mem[12][0] ), .Z(n1329) );
  OR U1818 ( .A(n1011), .B(n1331), .Z(n1328) );
  NAND U1819 ( .A(n1332), .B(n1333), .Z(\u_a23_mem/n19323 ) );
  NAND U1820 ( .A(n1330), .B(\u_a23_mem/p_mem[12][1] ), .Z(n1333) );
  OR U1821 ( .A(n1019), .B(n1331), .Z(n1332) );
  NAND U1822 ( .A(n1334), .B(n1335), .Z(\u_a23_mem/n19322 ) );
  NAND U1823 ( .A(n1330), .B(\u_a23_mem/p_mem[12][2] ), .Z(n1335) );
  OR U1824 ( .A(n1025), .B(n1331), .Z(n1334) );
  NAND U1825 ( .A(n1336), .B(n1337), .Z(\u_a23_mem/n19321 ) );
  NAND U1826 ( .A(n1330), .B(\u_a23_mem/p_mem[12][3] ), .Z(n1337) );
  OR U1827 ( .A(n1031), .B(n1331), .Z(n1336) );
  NAND U1828 ( .A(n1338), .B(n1339), .Z(\u_a23_mem/n19320 ) );
  NAND U1829 ( .A(n1330), .B(\u_a23_mem/p_mem[12][4] ), .Z(n1339) );
  OR U1830 ( .A(n1037), .B(n1331), .Z(n1338) );
  NAND U1831 ( .A(n1340), .B(n1341), .Z(\u_a23_mem/n19319 ) );
  NAND U1832 ( .A(n1330), .B(\u_a23_mem/p_mem[12][5] ), .Z(n1341) );
  OR U1833 ( .A(n1043), .B(n1331), .Z(n1340) );
  NAND U1834 ( .A(n1342), .B(n1343), .Z(\u_a23_mem/n19318 ) );
  NAND U1835 ( .A(n1330), .B(\u_a23_mem/p_mem[12][6] ), .Z(n1343) );
  OR U1836 ( .A(n1049), .B(n1331), .Z(n1342) );
  NAND U1837 ( .A(n1344), .B(n1345), .Z(\u_a23_mem/n19317 ) );
  NAND U1838 ( .A(n1330), .B(\u_a23_mem/p_mem[12][7] ), .Z(n1345) );
  NANDN U1839 ( .B(n1080), .A(n1346), .Z(n1330) );
  NANDN U1840 ( .B(n1331), .A(n1055), .Z(n1344) );
  NANDN U1841 ( .B(n2), .A(n1346), .Z(n1331) );
  NAND U1842 ( .A(n1347), .B(n1348), .Z(\u_a23_mem/n19316 ) );
  OR U1843 ( .A(n1011), .B(n1349), .Z(n1348) );
  AND U1844 ( .A(n1350), .B(n1351), .Z(n1347) );
  NANDN U1845 ( .B(n1087), .A(n1346), .Z(n1351) );
  NAND U1846 ( .A(n1352), .B(\u_a23_mem/p_mem[13][0] ), .Z(n1350) );
  NAND U1847 ( .A(n1353), .B(n1354), .Z(\u_a23_mem/n19315 ) );
  OR U1848 ( .A(n1019), .B(n1349), .Z(n1354) );
  AND U1849 ( .A(n1355), .B(n1356), .Z(n1353) );
  NANDN U1850 ( .B(n1093), .A(n1346), .Z(n1356) );
  NAND U1851 ( .A(n1352), .B(\u_a23_mem/p_mem[13][1] ), .Z(n1355) );
  NAND U1852 ( .A(n1357), .B(n1358), .Z(\u_a23_mem/n19314 ) );
  OR U1853 ( .A(n1025), .B(n1349), .Z(n1358) );
  AND U1854 ( .A(n1359), .B(n1360), .Z(n1357) );
  NANDN U1855 ( .B(n1098), .A(n1346), .Z(n1360) );
  NAND U1856 ( .A(n1352), .B(\u_a23_mem/p_mem[13][2] ), .Z(n1359) );
  NAND U1857 ( .A(n1361), .B(n1362), .Z(\u_a23_mem/n19313 ) );
  OR U1858 ( .A(n1031), .B(n1349), .Z(n1362) );
  AND U1859 ( .A(n1363), .B(n1364), .Z(n1361) );
  NANDN U1860 ( .B(n1103), .A(n1346), .Z(n1364) );
  NAND U1861 ( .A(n1352), .B(\u_a23_mem/p_mem[13][3] ), .Z(n1363) );
  NAND U1862 ( .A(n1365), .B(n1366), .Z(\u_a23_mem/n19312 ) );
  OR U1863 ( .A(n1037), .B(n1349), .Z(n1366) );
  AND U1864 ( .A(n1367), .B(n1368), .Z(n1365) );
  NANDN U1865 ( .B(n1108), .A(n1346), .Z(n1368) );
  NAND U1866 ( .A(n1352), .B(\u_a23_mem/p_mem[13][4] ), .Z(n1367) );
  NAND U1867 ( .A(n1369), .B(n1370), .Z(\u_a23_mem/n19311 ) );
  OR U1868 ( .A(n1043), .B(n1349), .Z(n1370) );
  AND U1869 ( .A(n1371), .B(n1372), .Z(n1369) );
  NANDN U1870 ( .B(n1113), .A(n1346), .Z(n1372) );
  NAND U1871 ( .A(n1352), .B(\u_a23_mem/p_mem[13][5] ), .Z(n1371) );
  NAND U1872 ( .A(n1373), .B(n1374), .Z(\u_a23_mem/n19310 ) );
  OR U1873 ( .A(n1049), .B(n1349), .Z(n1374) );
  AND U1874 ( .A(n1375), .B(n1376), .Z(n1373) );
  NANDN U1875 ( .B(n1118), .A(n1346), .Z(n1376) );
  NAND U1876 ( .A(n1352), .B(\u_a23_mem/p_mem[13][6] ), .Z(n1375) );
  NAND U1877 ( .A(n1377), .B(n1378), .Z(\u_a23_mem/n19309 ) );
  NANDN U1878 ( .B(n1349), .A(n1055), .Z(n1378) );
  NAND U1879 ( .A(n1121), .B(n1346), .Z(n1349) );
  AND U1880 ( .A(n1379), .B(n1380), .Z(n1377) );
  NANDN U1881 ( .B(n1124), .A(n1346), .Z(n1380) );
  NAND U1882 ( .A(n1352), .B(\u_a23_mem/p_mem[13][7] ), .Z(n1379) );
  NANDN U1883 ( .B(n1125), .A(n1346), .Z(n1352) );
  NAND U1884 ( .A(n1381), .B(n1382), .Z(\u_a23_mem/n19308 ) );
  OR U1885 ( .A(n1011), .B(n1383), .Z(n1382) );
  AND U1886 ( .A(n1384), .B(n1385), .Z(n1381) );
  NANDN U1887 ( .B(n1131), .A(n1346), .Z(n1385) );
  NAND U1888 ( .A(n1386), .B(\u_a23_mem/p_mem[14][0] ), .Z(n1384) );
  NAND U1889 ( .A(n1387), .B(n1388), .Z(\u_a23_mem/n19307 ) );
  OR U1890 ( .A(n1019), .B(n1383), .Z(n1388) );
  AND U1891 ( .A(n1389), .B(n1390), .Z(n1387) );
  NANDN U1892 ( .B(n1137), .A(n1346), .Z(n1390) );
  NAND U1893 ( .A(n1386), .B(\u_a23_mem/p_mem[14][1] ), .Z(n1389) );
  NAND U1894 ( .A(n1391), .B(n1392), .Z(\u_a23_mem/n19306 ) );
  OR U1895 ( .A(n1025), .B(n1383), .Z(n1392) );
  AND U1896 ( .A(n1393), .B(n1394), .Z(n1391) );
  NANDN U1897 ( .B(n1142), .A(n1346), .Z(n1394) );
  NAND U1898 ( .A(n1386), .B(\u_a23_mem/p_mem[14][2] ), .Z(n1393) );
  NAND U1899 ( .A(n1395), .B(n1396), .Z(\u_a23_mem/n19305 ) );
  OR U1900 ( .A(n1031), .B(n1383), .Z(n1396) );
  AND U1901 ( .A(n1397), .B(n1398), .Z(n1395) );
  NANDN U1902 ( .B(n1147), .A(n1346), .Z(n1398) );
  NAND U1903 ( .A(n1386), .B(\u_a23_mem/p_mem[14][3] ), .Z(n1397) );
  NAND U1904 ( .A(n1399), .B(n1400), .Z(\u_a23_mem/n19304 ) );
  OR U1905 ( .A(n1037), .B(n1383), .Z(n1400) );
  AND U1906 ( .A(n1401), .B(n1402), .Z(n1399) );
  NANDN U1907 ( .B(n1152), .A(n1346), .Z(n1402) );
  NAND U1908 ( .A(n1386), .B(\u_a23_mem/p_mem[14][4] ), .Z(n1401) );
  NAND U1909 ( .A(n1403), .B(n1404), .Z(\u_a23_mem/n19303 ) );
  OR U1910 ( .A(n1043), .B(n1383), .Z(n1404) );
  AND U1911 ( .A(n1405), .B(n1406), .Z(n1403) );
  NANDN U1912 ( .B(n1157), .A(n1346), .Z(n1406) );
  NAND U1913 ( .A(n1386), .B(\u_a23_mem/p_mem[14][5] ), .Z(n1405) );
  NAND U1914 ( .A(n1407), .B(n1408), .Z(\u_a23_mem/n19302 ) );
  OR U1915 ( .A(n1049), .B(n1383), .Z(n1408) );
  AND U1916 ( .A(n1409), .B(n1410), .Z(n1407) );
  NANDN U1917 ( .B(n1162), .A(n1346), .Z(n1410) );
  NAND U1918 ( .A(n1386), .B(\u_a23_mem/p_mem[14][6] ), .Z(n1409) );
  NAND U1919 ( .A(n1411), .B(n1412), .Z(\u_a23_mem/n19301 ) );
  NANDN U1920 ( .B(n1383), .A(n1055), .Z(n1412) );
  NAND U1921 ( .A(n1165), .B(n1346), .Z(n1383) );
  AND U1922 ( .A(n1413), .B(n1414), .Z(n1411) );
  NANDN U1923 ( .B(n1168), .A(n1346), .Z(n1414) );
  NAND U1924 ( .A(n1386), .B(\u_a23_mem/p_mem[14][7] ), .Z(n1413) );
  NANDN U1925 ( .B(n1169), .A(n1346), .Z(n1386) );
  NAND U1926 ( .A(n1415), .B(n1416), .Z(\u_a23_mem/n19300 ) );
  OR U1927 ( .A(n1011), .B(n1417), .Z(n1416) );
  AND U1928 ( .A(n1418), .B(n1419), .Z(n1415) );
  NAND U1929 ( .A(n1420), .B(\u_a23_mem/p_mem[15][0] ), .Z(n1419) );
  NANDN U1930 ( .B(n1015), .A(n1346), .Z(n1418) );
  NAND U1931 ( .A(n1421), .B(n1422), .Z(\u_a23_mem/n19299 ) );
  OR U1932 ( .A(n1019), .B(n1417), .Z(n1422) );
  AND U1933 ( .A(n1423), .B(n1424), .Z(n1421) );
  NAND U1934 ( .A(n1420), .B(\u_a23_mem/p_mem[15][1] ), .Z(n1424) );
  NANDN U1935 ( .B(n1022), .A(n1346), .Z(n1423) );
  NAND U1936 ( .A(n1425), .B(n1426), .Z(\u_a23_mem/n19298 ) );
  OR U1937 ( .A(n1025), .B(n1417), .Z(n1426) );
  AND U1938 ( .A(n1427), .B(n1428), .Z(n1425) );
  NAND U1939 ( .A(n1420), .B(\u_a23_mem/p_mem[15][2] ), .Z(n1428) );
  NANDN U1940 ( .B(n1028), .A(n1346), .Z(n1427) );
  NAND U1941 ( .A(n1429), .B(n1430), .Z(\u_a23_mem/n19297 ) );
  OR U1942 ( .A(n1031), .B(n1417), .Z(n1430) );
  AND U1943 ( .A(n1431), .B(n1432), .Z(n1429) );
  NAND U1944 ( .A(n1420), .B(\u_a23_mem/p_mem[15][3] ), .Z(n1432) );
  NANDN U1945 ( .B(n1034), .A(n1346), .Z(n1431) );
  NAND U1946 ( .A(n1433), .B(n1434), .Z(\u_a23_mem/n19296 ) );
  OR U1947 ( .A(n1037), .B(n1417), .Z(n1434) );
  AND U1948 ( .A(n1435), .B(n1436), .Z(n1433) );
  NAND U1949 ( .A(n1420), .B(\u_a23_mem/p_mem[15][4] ), .Z(n1436) );
  NANDN U1950 ( .B(n1040), .A(n1346), .Z(n1435) );
  NAND U1951 ( .A(n1437), .B(n1438), .Z(\u_a23_mem/n19295 ) );
  OR U1952 ( .A(n1043), .B(n1417), .Z(n1438) );
  AND U1953 ( .A(n1439), .B(n1440), .Z(n1437) );
  NAND U1954 ( .A(n1420), .B(\u_a23_mem/p_mem[15][5] ), .Z(n1440) );
  NANDN U1955 ( .B(n1046), .A(n1346), .Z(n1439) );
  NAND U1956 ( .A(n1441), .B(n1442), .Z(\u_a23_mem/n19294 ) );
  OR U1957 ( .A(n1049), .B(n1417), .Z(n1442) );
  AND U1958 ( .A(n1443), .B(n1444), .Z(n1441) );
  NAND U1959 ( .A(n1420), .B(\u_a23_mem/p_mem[15][6] ), .Z(n1444) );
  NANDN U1960 ( .B(n1052), .A(n1346), .Z(n1443) );
  NAND U1961 ( .A(n1445), .B(n1446), .Z(\u_a23_mem/n19293 ) );
  NANDN U1962 ( .B(n1417), .A(n1055), .Z(n1446) );
  NAND U1963 ( .A(n1056), .B(n1346), .Z(n1417) );
  AND U1964 ( .A(n1447), .B(n1448), .Z(n1445) );
  NAND U1965 ( .A(n1420), .B(\u_a23_mem/p_mem[15][7] ), .Z(n1448) );
  NANDN U1966 ( .B(n1059), .A(n1346), .Z(n1420) );
  NAND U1967 ( .A(n1061), .B(n1346), .Z(n1447) );
  ANDN U1968 ( .A(n1449), .B(n1205), .Z(n1346) );
  NAND U1969 ( .A(n1450), .B(n1451), .Z(\u_a23_mem/n19292 ) );
  NAND U1970 ( .A(n1452), .B(\u_a23_mem/p_mem[16][0] ), .Z(n1451) );
  OR U1971 ( .A(n1011), .B(n1453), .Z(n1450) );
  NAND U1972 ( .A(n1454), .B(n1455), .Z(\u_a23_mem/n19291 ) );
  NAND U1973 ( .A(n1452), .B(\u_a23_mem/p_mem[16][1] ), .Z(n1455) );
  OR U1974 ( .A(n1019), .B(n1453), .Z(n1454) );
  NAND U1975 ( .A(n1456), .B(n1457), .Z(\u_a23_mem/n19290 ) );
  NAND U1976 ( .A(n1452), .B(\u_a23_mem/p_mem[16][2] ), .Z(n1457) );
  OR U1977 ( .A(n1025), .B(n1453), .Z(n1456) );
  NAND U1978 ( .A(n1458), .B(n1459), .Z(\u_a23_mem/n19289 ) );
  NAND U1979 ( .A(n1452), .B(\u_a23_mem/p_mem[16][3] ), .Z(n1459) );
  OR U1980 ( .A(n1031), .B(n1453), .Z(n1458) );
  NAND U1981 ( .A(n1460), .B(n1461), .Z(\u_a23_mem/n19288 ) );
  NAND U1982 ( .A(n1452), .B(\u_a23_mem/p_mem[16][4] ), .Z(n1461) );
  OR U1983 ( .A(n1037), .B(n1453), .Z(n1460) );
  NAND U1984 ( .A(n1462), .B(n1463), .Z(\u_a23_mem/n19287 ) );
  NAND U1985 ( .A(n1452), .B(\u_a23_mem/p_mem[16][5] ), .Z(n1463) );
  OR U1986 ( .A(n1043), .B(n1453), .Z(n1462) );
  NAND U1987 ( .A(n1464), .B(n1465), .Z(\u_a23_mem/n19286 ) );
  NAND U1988 ( .A(n1452), .B(\u_a23_mem/p_mem[16][6] ), .Z(n1465) );
  OR U1989 ( .A(n1049), .B(n1453), .Z(n1464) );
  NAND U1990 ( .A(n1466), .B(n1467), .Z(\u_a23_mem/n19285 ) );
  NAND U1991 ( .A(n1452), .B(\u_a23_mem/p_mem[16][7] ), .Z(n1467) );
  NANDN U1992 ( .B(n1080), .A(n1468), .Z(n1452) );
  NANDN U1993 ( .B(n1453), .A(n1055), .Z(n1466) );
  NANDN U1994 ( .B(n2), .A(n1468), .Z(n1453) );
  NAND U1995 ( .A(n1469), .B(n1470), .Z(\u_a23_mem/n19284 ) );
  OR U1996 ( .A(n1011), .B(n1471), .Z(n1470) );
  AND U1997 ( .A(n1472), .B(n1473), .Z(n1469) );
  NANDN U1998 ( .B(n1087), .A(n1468), .Z(n1473) );
  NAND U1999 ( .A(n1474), .B(\u_a23_mem/p_mem[17][0] ), .Z(n1472) );
  NAND U2000 ( .A(n1475), .B(n1476), .Z(\u_a23_mem/n19283 ) );
  OR U2001 ( .A(n1019), .B(n1471), .Z(n1476) );
  AND U2002 ( .A(n1477), .B(n1478), .Z(n1475) );
  NANDN U2003 ( .B(n1093), .A(n1468), .Z(n1478) );
  NAND U2004 ( .A(n1474), .B(\u_a23_mem/p_mem[17][1] ), .Z(n1477) );
  NAND U2005 ( .A(n1479), .B(n1480), .Z(\u_a23_mem/n19282 ) );
  OR U2006 ( .A(n1025), .B(n1471), .Z(n1480) );
  AND U2007 ( .A(n1481), .B(n1482), .Z(n1479) );
  NANDN U2008 ( .B(n1098), .A(n1468), .Z(n1482) );
  NAND U2009 ( .A(n1474), .B(\u_a23_mem/p_mem[17][2] ), .Z(n1481) );
  NAND U2010 ( .A(n1483), .B(n1484), .Z(\u_a23_mem/n19281 ) );
  OR U2011 ( .A(n1031), .B(n1471), .Z(n1484) );
  AND U2012 ( .A(n1485), .B(n1486), .Z(n1483) );
  NANDN U2013 ( .B(n1103), .A(n1468), .Z(n1486) );
  NAND U2014 ( .A(n1474), .B(\u_a23_mem/p_mem[17][3] ), .Z(n1485) );
  NAND U2015 ( .A(n1487), .B(n1488), .Z(\u_a23_mem/n19280 ) );
  OR U2016 ( .A(n1037), .B(n1471), .Z(n1488) );
  AND U2017 ( .A(n1489), .B(n1490), .Z(n1487) );
  NANDN U2018 ( .B(n1108), .A(n1468), .Z(n1490) );
  NAND U2019 ( .A(n1474), .B(\u_a23_mem/p_mem[17][4] ), .Z(n1489) );
  NAND U2020 ( .A(n1491), .B(n1492), .Z(\u_a23_mem/n19279 ) );
  OR U2021 ( .A(n1043), .B(n1471), .Z(n1492) );
  AND U2022 ( .A(n1493), .B(n1494), .Z(n1491) );
  NANDN U2023 ( .B(n1113), .A(n1468), .Z(n1494) );
  NAND U2024 ( .A(n1474), .B(\u_a23_mem/p_mem[17][5] ), .Z(n1493) );
  NAND U2025 ( .A(n1495), .B(n1496), .Z(\u_a23_mem/n19278 ) );
  OR U2026 ( .A(n1049), .B(n1471), .Z(n1496) );
  AND U2027 ( .A(n1497), .B(n1498), .Z(n1495) );
  NANDN U2028 ( .B(n1118), .A(n1468), .Z(n1498) );
  NAND U2029 ( .A(n1474), .B(\u_a23_mem/p_mem[17][6] ), .Z(n1497) );
  NAND U2030 ( .A(n1499), .B(n1500), .Z(\u_a23_mem/n19277 ) );
  NANDN U2031 ( .B(n1471), .A(n1055), .Z(n1500) );
  NAND U2032 ( .A(n1121), .B(n1468), .Z(n1471) );
  AND U2033 ( .A(n1501), .B(n1502), .Z(n1499) );
  NANDN U2034 ( .B(n1124), .A(n1468), .Z(n1502) );
  NAND U2035 ( .A(n1474), .B(\u_a23_mem/p_mem[17][7] ), .Z(n1501) );
  NANDN U2036 ( .B(n1125), .A(n1468), .Z(n1474) );
  NAND U2037 ( .A(n1503), .B(n1504), .Z(\u_a23_mem/n19276 ) );
  OR U2038 ( .A(n1011), .B(n1505), .Z(n1504) );
  AND U2039 ( .A(n1506), .B(n1507), .Z(n1503) );
  NANDN U2040 ( .B(n1131), .A(n1468), .Z(n1507) );
  NAND U2041 ( .A(n1508), .B(\u_a23_mem/p_mem[18][0] ), .Z(n1506) );
  NAND U2042 ( .A(n1509), .B(n1510), .Z(\u_a23_mem/n19275 ) );
  OR U2043 ( .A(n1019), .B(n1505), .Z(n1510) );
  AND U2044 ( .A(n1511), .B(n1512), .Z(n1509) );
  NANDN U2045 ( .B(n1137), .A(n1468), .Z(n1512) );
  NAND U2046 ( .A(n1508), .B(\u_a23_mem/p_mem[18][1] ), .Z(n1511) );
  NAND U2047 ( .A(n1513), .B(n1514), .Z(\u_a23_mem/n19274 ) );
  OR U2048 ( .A(n1025), .B(n1505), .Z(n1514) );
  AND U2049 ( .A(n1515), .B(n1516), .Z(n1513) );
  NANDN U2050 ( .B(n1142), .A(n1468), .Z(n1516) );
  NAND U2051 ( .A(n1508), .B(\u_a23_mem/p_mem[18][2] ), .Z(n1515) );
  NAND U2052 ( .A(n1517), .B(n1518), .Z(\u_a23_mem/n19273 ) );
  OR U2053 ( .A(n1031), .B(n1505), .Z(n1518) );
  AND U2054 ( .A(n1519), .B(n1520), .Z(n1517) );
  NANDN U2055 ( .B(n1147), .A(n1468), .Z(n1520) );
  NAND U2056 ( .A(n1508), .B(\u_a23_mem/p_mem[18][3] ), .Z(n1519) );
  NAND U2057 ( .A(n1521), .B(n1522), .Z(\u_a23_mem/n19272 ) );
  OR U2058 ( .A(n1037), .B(n1505), .Z(n1522) );
  AND U2059 ( .A(n1523), .B(n1524), .Z(n1521) );
  NANDN U2060 ( .B(n1152), .A(n1468), .Z(n1524) );
  NAND U2061 ( .A(n1508), .B(\u_a23_mem/p_mem[18][4] ), .Z(n1523) );
  NAND U2062 ( .A(n1525), .B(n1526), .Z(\u_a23_mem/n19271 ) );
  OR U2063 ( .A(n1043), .B(n1505), .Z(n1526) );
  AND U2064 ( .A(n1527), .B(n1528), .Z(n1525) );
  NANDN U2065 ( .B(n1157), .A(n1468), .Z(n1528) );
  NAND U2066 ( .A(n1508), .B(\u_a23_mem/p_mem[18][5] ), .Z(n1527) );
  NAND U2067 ( .A(n1529), .B(n1530), .Z(\u_a23_mem/n19270 ) );
  OR U2068 ( .A(n1049), .B(n1505), .Z(n1530) );
  AND U2069 ( .A(n1531), .B(n1532), .Z(n1529) );
  NANDN U2070 ( .B(n1162), .A(n1468), .Z(n1532) );
  NAND U2071 ( .A(n1508), .B(\u_a23_mem/p_mem[18][6] ), .Z(n1531) );
  NAND U2072 ( .A(n1533), .B(n1534), .Z(\u_a23_mem/n19269 ) );
  NANDN U2073 ( .B(n1505), .A(n1055), .Z(n1534) );
  NAND U2074 ( .A(n1165), .B(n1468), .Z(n1505) );
  AND U2075 ( .A(n1535), .B(n1536), .Z(n1533) );
  NANDN U2076 ( .B(n1168), .A(n1468), .Z(n1536) );
  NAND U2077 ( .A(n1508), .B(\u_a23_mem/p_mem[18][7] ), .Z(n1535) );
  NANDN U2078 ( .B(n1169), .A(n1468), .Z(n1508) );
  NAND U2079 ( .A(n1537), .B(n1538), .Z(\u_a23_mem/n19268 ) );
  OR U2080 ( .A(n1011), .B(n1539), .Z(n1538) );
  AND U2081 ( .A(n1540), .B(n1541), .Z(n1537) );
  NAND U2082 ( .A(n1542), .B(\u_a23_mem/p_mem[19][0] ), .Z(n1541) );
  NANDN U2083 ( .B(n1015), .A(n1468), .Z(n1540) );
  NAND U2084 ( .A(n1543), .B(n1544), .Z(\u_a23_mem/n19267 ) );
  OR U2085 ( .A(n1019), .B(n1539), .Z(n1544) );
  AND U2086 ( .A(n1545), .B(n1546), .Z(n1543) );
  NAND U2087 ( .A(n1542), .B(\u_a23_mem/p_mem[19][1] ), .Z(n1546) );
  NANDN U2088 ( .B(n1022), .A(n1468), .Z(n1545) );
  NAND U2089 ( .A(n1547), .B(n1548), .Z(\u_a23_mem/n19266 ) );
  OR U2090 ( .A(n1025), .B(n1539), .Z(n1548) );
  AND U2091 ( .A(n1549), .B(n1550), .Z(n1547) );
  NAND U2092 ( .A(n1542), .B(\u_a23_mem/p_mem[19][2] ), .Z(n1550) );
  NANDN U2093 ( .B(n1028), .A(n1468), .Z(n1549) );
  NAND U2094 ( .A(n1551), .B(n1552), .Z(\u_a23_mem/n19265 ) );
  OR U2095 ( .A(n1031), .B(n1539), .Z(n1552) );
  AND U2096 ( .A(n1553), .B(n1554), .Z(n1551) );
  NAND U2097 ( .A(n1542), .B(\u_a23_mem/p_mem[19][3] ), .Z(n1554) );
  NANDN U2098 ( .B(n1034), .A(n1468), .Z(n1553) );
  NAND U2099 ( .A(n1555), .B(n1556), .Z(\u_a23_mem/n19264 ) );
  OR U2100 ( .A(n1037), .B(n1539), .Z(n1556) );
  AND U2101 ( .A(n1557), .B(n1558), .Z(n1555) );
  NAND U2102 ( .A(n1542), .B(\u_a23_mem/p_mem[19][4] ), .Z(n1558) );
  NANDN U2103 ( .B(n1040), .A(n1468), .Z(n1557) );
  NAND U2104 ( .A(n1559), .B(n1560), .Z(\u_a23_mem/n19263 ) );
  OR U2105 ( .A(n1043), .B(n1539), .Z(n1560) );
  AND U2106 ( .A(n1561), .B(n1562), .Z(n1559) );
  NAND U2107 ( .A(n1542), .B(\u_a23_mem/p_mem[19][5] ), .Z(n1562) );
  NANDN U2108 ( .B(n1046), .A(n1468), .Z(n1561) );
  NAND U2109 ( .A(n1563), .B(n1564), .Z(\u_a23_mem/n19262 ) );
  OR U2110 ( .A(n1049), .B(n1539), .Z(n1564) );
  AND U2111 ( .A(n1565), .B(n1566), .Z(n1563) );
  NAND U2112 ( .A(n1542), .B(\u_a23_mem/p_mem[19][6] ), .Z(n1566) );
  NANDN U2113 ( .B(n1052), .A(n1468), .Z(n1565) );
  NAND U2114 ( .A(n1567), .B(n1568), .Z(\u_a23_mem/n19261 ) );
  NANDN U2115 ( .B(n1539), .A(n1055), .Z(n1568) );
  NAND U2116 ( .A(n1056), .B(n1468), .Z(n1539) );
  AND U2117 ( .A(n1569), .B(n1570), .Z(n1567) );
  NAND U2118 ( .A(n1542), .B(\u_a23_mem/p_mem[19][7] ), .Z(n1570) );
  NANDN U2119 ( .B(n1059), .A(n1468), .Z(n1542) );
  NAND U2120 ( .A(n1061), .B(n1468), .Z(n1569) );
  ANDN U2121 ( .A(n1571), .B(n1572), .Z(n1468) );
  NAND U2122 ( .A(n1573), .B(n1574), .Z(\u_a23_mem/n19260 ) );
  NAND U2123 ( .A(n1575), .B(\u_a23_mem/p_mem[20][0] ), .Z(n1574) );
  OR U2124 ( .A(n1011), .B(n1576), .Z(n1573) );
  NAND U2125 ( .A(n1577), .B(n1578), .Z(\u_a23_mem/n19259 ) );
  NAND U2126 ( .A(n1575), .B(\u_a23_mem/p_mem[20][1] ), .Z(n1578) );
  OR U2127 ( .A(n1019), .B(n1576), .Z(n1577) );
  NAND U2128 ( .A(n1579), .B(n1580), .Z(\u_a23_mem/n19258 ) );
  NAND U2129 ( .A(n1575), .B(\u_a23_mem/p_mem[20][2] ), .Z(n1580) );
  OR U2130 ( .A(n1025), .B(n1576), .Z(n1579) );
  NAND U2131 ( .A(n1581), .B(n1582), .Z(\u_a23_mem/n19257 ) );
  NAND U2132 ( .A(n1575), .B(\u_a23_mem/p_mem[20][3] ), .Z(n1582) );
  OR U2133 ( .A(n1031), .B(n1576), .Z(n1581) );
  NAND U2134 ( .A(n1583), .B(n1584), .Z(\u_a23_mem/n19256 ) );
  NAND U2135 ( .A(n1575), .B(\u_a23_mem/p_mem[20][4] ), .Z(n1584) );
  OR U2136 ( .A(n1037), .B(n1576), .Z(n1583) );
  NAND U2137 ( .A(n1585), .B(n1586), .Z(\u_a23_mem/n19255 ) );
  NAND U2138 ( .A(n1575), .B(\u_a23_mem/p_mem[20][5] ), .Z(n1586) );
  OR U2139 ( .A(n1043), .B(n1576), .Z(n1585) );
  NAND U2140 ( .A(n1587), .B(n1588), .Z(\u_a23_mem/n19254 ) );
  NAND U2141 ( .A(n1575), .B(\u_a23_mem/p_mem[20][6] ), .Z(n1588) );
  OR U2142 ( .A(n1049), .B(n1576), .Z(n1587) );
  NAND U2143 ( .A(n1589), .B(n1590), .Z(\u_a23_mem/n19253 ) );
  NAND U2144 ( .A(n1575), .B(\u_a23_mem/p_mem[20][7] ), .Z(n1590) );
  NANDN U2145 ( .B(n1080), .A(n1591), .Z(n1575) );
  NANDN U2146 ( .B(n1576), .A(n1055), .Z(n1589) );
  NANDN U2147 ( .B(n2), .A(n1591), .Z(n1576) );
  NAND U2148 ( .A(n1592), .B(n1593), .Z(\u_a23_mem/n19252 ) );
  OR U2149 ( .A(n1011), .B(n1594), .Z(n1593) );
  AND U2150 ( .A(n1595), .B(n1596), .Z(n1592) );
  NANDN U2151 ( .B(n1087), .A(n1591), .Z(n1596) );
  NAND U2152 ( .A(n1597), .B(\u_a23_mem/p_mem[21][0] ), .Z(n1595) );
  NAND U2153 ( .A(n1598), .B(n1599), .Z(\u_a23_mem/n19251 ) );
  OR U2154 ( .A(n1019), .B(n1594), .Z(n1599) );
  AND U2155 ( .A(n1600), .B(n1601), .Z(n1598) );
  NANDN U2156 ( .B(n1093), .A(n1591), .Z(n1601) );
  NAND U2157 ( .A(n1597), .B(\u_a23_mem/p_mem[21][1] ), .Z(n1600) );
  NAND U2158 ( .A(n1602), .B(n1603), .Z(\u_a23_mem/n19250 ) );
  OR U2159 ( .A(n1025), .B(n1594), .Z(n1603) );
  AND U2160 ( .A(n1604), .B(n1605), .Z(n1602) );
  NANDN U2161 ( .B(n1098), .A(n1591), .Z(n1605) );
  NAND U2162 ( .A(n1597), .B(\u_a23_mem/p_mem[21][2] ), .Z(n1604) );
  NAND U2163 ( .A(n1606), .B(n1607), .Z(\u_a23_mem/n19249 ) );
  OR U2164 ( .A(n1031), .B(n1594), .Z(n1607) );
  AND U2165 ( .A(n1608), .B(n1609), .Z(n1606) );
  NANDN U2166 ( .B(n1103), .A(n1591), .Z(n1609) );
  NAND U2167 ( .A(n1597), .B(\u_a23_mem/p_mem[21][3] ), .Z(n1608) );
  NAND U2168 ( .A(n1610), .B(n1611), .Z(\u_a23_mem/n19248 ) );
  OR U2169 ( .A(n1037), .B(n1594), .Z(n1611) );
  AND U2170 ( .A(n1612), .B(n1613), .Z(n1610) );
  NANDN U2171 ( .B(n1108), .A(n1591), .Z(n1613) );
  NAND U2172 ( .A(n1597), .B(\u_a23_mem/p_mem[21][4] ), .Z(n1612) );
  NAND U2173 ( .A(n1614), .B(n1615), .Z(\u_a23_mem/n19247 ) );
  OR U2174 ( .A(n1043), .B(n1594), .Z(n1615) );
  AND U2175 ( .A(n1616), .B(n1617), .Z(n1614) );
  NANDN U2176 ( .B(n1113), .A(n1591), .Z(n1617) );
  NAND U2177 ( .A(n1597), .B(\u_a23_mem/p_mem[21][5] ), .Z(n1616) );
  NAND U2178 ( .A(n1618), .B(n1619), .Z(\u_a23_mem/n19246 ) );
  OR U2179 ( .A(n1049), .B(n1594), .Z(n1619) );
  AND U2180 ( .A(n1620), .B(n1621), .Z(n1618) );
  NANDN U2181 ( .B(n1118), .A(n1591), .Z(n1621) );
  NAND U2182 ( .A(n1597), .B(\u_a23_mem/p_mem[21][6] ), .Z(n1620) );
  NAND U2183 ( .A(n1622), .B(n1623), .Z(\u_a23_mem/n19245 ) );
  NANDN U2184 ( .B(n1594), .A(n1055), .Z(n1623) );
  NAND U2185 ( .A(n1121), .B(n1591), .Z(n1594) );
  AND U2186 ( .A(n1624), .B(n1625), .Z(n1622) );
  NANDN U2187 ( .B(n1124), .A(n1591), .Z(n1625) );
  NAND U2188 ( .A(n1597), .B(\u_a23_mem/p_mem[21][7] ), .Z(n1624) );
  NANDN U2189 ( .B(n1125), .A(n1591), .Z(n1597) );
  NAND U2190 ( .A(n1626), .B(n1627), .Z(\u_a23_mem/n19244 ) );
  OR U2191 ( .A(n1011), .B(n1628), .Z(n1627) );
  AND U2192 ( .A(n1629), .B(n1630), .Z(n1626) );
  NANDN U2193 ( .B(n1131), .A(n1591), .Z(n1630) );
  NAND U2194 ( .A(n1631), .B(\u_a23_mem/p_mem[22][0] ), .Z(n1629) );
  NAND U2195 ( .A(n1632), .B(n1633), .Z(\u_a23_mem/n19243 ) );
  OR U2196 ( .A(n1019), .B(n1628), .Z(n1633) );
  AND U2197 ( .A(n1634), .B(n1635), .Z(n1632) );
  NANDN U2198 ( .B(n1137), .A(n1591), .Z(n1635) );
  NAND U2199 ( .A(n1631), .B(\u_a23_mem/p_mem[22][1] ), .Z(n1634) );
  NAND U2200 ( .A(n1636), .B(n1637), .Z(\u_a23_mem/n19242 ) );
  OR U2201 ( .A(n1025), .B(n1628), .Z(n1637) );
  AND U2202 ( .A(n1638), .B(n1639), .Z(n1636) );
  NANDN U2203 ( .B(n1142), .A(n1591), .Z(n1639) );
  NAND U2204 ( .A(n1631), .B(\u_a23_mem/p_mem[22][2] ), .Z(n1638) );
  NAND U2205 ( .A(n1640), .B(n1641), .Z(\u_a23_mem/n19241 ) );
  OR U2206 ( .A(n1031), .B(n1628), .Z(n1641) );
  AND U2207 ( .A(n1642), .B(n1643), .Z(n1640) );
  NANDN U2208 ( .B(n1147), .A(n1591), .Z(n1643) );
  NAND U2209 ( .A(n1631), .B(\u_a23_mem/p_mem[22][3] ), .Z(n1642) );
  NAND U2210 ( .A(n1644), .B(n1645), .Z(\u_a23_mem/n19240 ) );
  OR U2211 ( .A(n1037), .B(n1628), .Z(n1645) );
  AND U2212 ( .A(n1646), .B(n1647), .Z(n1644) );
  NANDN U2213 ( .B(n1152), .A(n1591), .Z(n1647) );
  NAND U2214 ( .A(n1631), .B(\u_a23_mem/p_mem[22][4] ), .Z(n1646) );
  NAND U2215 ( .A(n1648), .B(n1649), .Z(\u_a23_mem/n19239 ) );
  OR U2216 ( .A(n1043), .B(n1628), .Z(n1649) );
  AND U2217 ( .A(n1650), .B(n1651), .Z(n1648) );
  NANDN U2218 ( .B(n1157), .A(n1591), .Z(n1651) );
  NAND U2219 ( .A(n1631), .B(\u_a23_mem/p_mem[22][5] ), .Z(n1650) );
  NAND U2220 ( .A(n1652), .B(n1653), .Z(\u_a23_mem/n19238 ) );
  OR U2221 ( .A(n1049), .B(n1628), .Z(n1653) );
  AND U2222 ( .A(n1654), .B(n1655), .Z(n1652) );
  NANDN U2223 ( .B(n1162), .A(n1591), .Z(n1655) );
  NAND U2224 ( .A(n1631), .B(\u_a23_mem/p_mem[22][6] ), .Z(n1654) );
  NAND U2225 ( .A(n1656), .B(n1657), .Z(\u_a23_mem/n19237 ) );
  NANDN U2226 ( .B(n1628), .A(n1055), .Z(n1657) );
  NAND U2227 ( .A(n1165), .B(n1591), .Z(n1628) );
  AND U2228 ( .A(n1658), .B(n1659), .Z(n1656) );
  NANDN U2229 ( .B(n1168), .A(n1591), .Z(n1659) );
  NAND U2230 ( .A(n1631), .B(\u_a23_mem/p_mem[22][7] ), .Z(n1658) );
  NANDN U2231 ( .B(n1169), .A(n1591), .Z(n1631) );
  NAND U2232 ( .A(n1660), .B(n1661), .Z(\u_a23_mem/n19236 ) );
  OR U2233 ( .A(n1011), .B(n1662), .Z(n1661) );
  AND U2234 ( .A(n1663), .B(n1664), .Z(n1660) );
  NAND U2235 ( .A(n1665), .B(\u_a23_mem/p_mem[23][0] ), .Z(n1664) );
  NANDN U2236 ( .B(n1015), .A(n1591), .Z(n1663) );
  NAND U2237 ( .A(n1666), .B(n1667), .Z(\u_a23_mem/n19235 ) );
  OR U2238 ( .A(n1019), .B(n1662), .Z(n1667) );
  AND U2239 ( .A(n1668), .B(n1669), .Z(n1666) );
  NAND U2240 ( .A(n1665), .B(\u_a23_mem/p_mem[23][1] ), .Z(n1669) );
  NANDN U2241 ( .B(n1022), .A(n1591), .Z(n1668) );
  NAND U2242 ( .A(n1670), .B(n1671), .Z(\u_a23_mem/n19234 ) );
  OR U2243 ( .A(n1025), .B(n1662), .Z(n1671) );
  AND U2244 ( .A(n1672), .B(n1673), .Z(n1670) );
  NAND U2245 ( .A(n1665), .B(\u_a23_mem/p_mem[23][2] ), .Z(n1673) );
  NANDN U2246 ( .B(n1028), .A(n1591), .Z(n1672) );
  NAND U2247 ( .A(n1674), .B(n1675), .Z(\u_a23_mem/n19233 ) );
  OR U2248 ( .A(n1031), .B(n1662), .Z(n1675) );
  AND U2249 ( .A(n1676), .B(n1677), .Z(n1674) );
  NAND U2250 ( .A(n1665), .B(\u_a23_mem/p_mem[23][3] ), .Z(n1677) );
  NANDN U2251 ( .B(n1034), .A(n1591), .Z(n1676) );
  NAND U2252 ( .A(n1678), .B(n1679), .Z(\u_a23_mem/n19232 ) );
  OR U2253 ( .A(n1037), .B(n1662), .Z(n1679) );
  AND U2254 ( .A(n1680), .B(n1681), .Z(n1678) );
  NAND U2255 ( .A(n1665), .B(\u_a23_mem/p_mem[23][4] ), .Z(n1681) );
  NANDN U2256 ( .B(n1040), .A(n1591), .Z(n1680) );
  NAND U2257 ( .A(n1682), .B(n1683), .Z(\u_a23_mem/n19231 ) );
  OR U2258 ( .A(n1043), .B(n1662), .Z(n1683) );
  AND U2259 ( .A(n1684), .B(n1685), .Z(n1682) );
  NAND U2260 ( .A(n1665), .B(\u_a23_mem/p_mem[23][5] ), .Z(n1685) );
  NANDN U2261 ( .B(n1046), .A(n1591), .Z(n1684) );
  NAND U2262 ( .A(n1686), .B(n1687), .Z(\u_a23_mem/n19230 ) );
  OR U2263 ( .A(n1049), .B(n1662), .Z(n1687) );
  AND U2264 ( .A(n1688), .B(n1689), .Z(n1686) );
  NAND U2265 ( .A(n1665), .B(\u_a23_mem/p_mem[23][6] ), .Z(n1689) );
  NANDN U2266 ( .B(n1052), .A(n1591), .Z(n1688) );
  NAND U2267 ( .A(n1690), .B(n1691), .Z(\u_a23_mem/n19229 ) );
  NANDN U2268 ( .B(n1662), .A(n1055), .Z(n1691) );
  NAND U2269 ( .A(n1056), .B(n1591), .Z(n1662) );
  AND U2270 ( .A(n1692), .B(n1693), .Z(n1690) );
  NAND U2271 ( .A(n1665), .B(\u_a23_mem/p_mem[23][7] ), .Z(n1693) );
  NANDN U2272 ( .B(n1059), .A(n1591), .Z(n1665) );
  NAND U2273 ( .A(n1061), .B(n1591), .Z(n1692) );
  ANDN U2274 ( .A(n1694), .B(n1572), .Z(n1591) );
  NAND U2275 ( .A(n1695), .B(n1696), .Z(\u_a23_mem/n19228 ) );
  NAND U2276 ( .A(n1697), .B(\u_a23_mem/p_mem[24][0] ), .Z(n1696) );
  OR U2277 ( .A(n1011), .B(n1698), .Z(n1695) );
  NAND U2278 ( .A(n1699), .B(n1700), .Z(\u_a23_mem/n19227 ) );
  NAND U2279 ( .A(n1697), .B(\u_a23_mem/p_mem[24][1] ), .Z(n1700) );
  OR U2280 ( .A(n1019), .B(n1698), .Z(n1699) );
  NAND U2281 ( .A(n1701), .B(n1702), .Z(\u_a23_mem/n19226 ) );
  NAND U2282 ( .A(n1697), .B(\u_a23_mem/p_mem[24][2] ), .Z(n1702) );
  OR U2283 ( .A(n1025), .B(n1698), .Z(n1701) );
  NAND U2284 ( .A(n1703), .B(n1704), .Z(\u_a23_mem/n19225 ) );
  NAND U2285 ( .A(n1697), .B(\u_a23_mem/p_mem[24][3] ), .Z(n1704) );
  OR U2286 ( .A(n1031), .B(n1698), .Z(n1703) );
  NAND U2287 ( .A(n1705), .B(n1706), .Z(\u_a23_mem/n19224 ) );
  NAND U2288 ( .A(n1697), .B(\u_a23_mem/p_mem[24][4] ), .Z(n1706) );
  OR U2289 ( .A(n1037), .B(n1698), .Z(n1705) );
  NAND U2290 ( .A(n1707), .B(n1708), .Z(\u_a23_mem/n19223 ) );
  NAND U2291 ( .A(n1697), .B(\u_a23_mem/p_mem[24][5] ), .Z(n1708) );
  OR U2292 ( .A(n1043), .B(n1698), .Z(n1707) );
  NAND U2293 ( .A(n1709), .B(n1710), .Z(\u_a23_mem/n19222 ) );
  NAND U2294 ( .A(n1697), .B(\u_a23_mem/p_mem[24][6] ), .Z(n1710) );
  OR U2295 ( .A(n1049), .B(n1698), .Z(n1709) );
  NAND U2296 ( .A(n1711), .B(n1712), .Z(\u_a23_mem/n19221 ) );
  NAND U2297 ( .A(n1697), .B(\u_a23_mem/p_mem[24][7] ), .Z(n1712) );
  NANDN U2298 ( .B(n1080), .A(n1713), .Z(n1697) );
  NANDN U2299 ( .B(n1698), .A(n1055), .Z(n1711) );
  NANDN U2300 ( .B(n2), .A(n1713), .Z(n1698) );
  NAND U2301 ( .A(n1714), .B(n1715), .Z(\u_a23_mem/n19220 ) );
  OR U2302 ( .A(n1011), .B(n1716), .Z(n1715) );
  AND U2303 ( .A(n1717), .B(n1718), .Z(n1714) );
  NANDN U2304 ( .B(n1087), .A(n1713), .Z(n1718) );
  NAND U2305 ( .A(n1719), .B(\u_a23_mem/p_mem[25][0] ), .Z(n1717) );
  NAND U2306 ( .A(n1720), .B(n1721), .Z(\u_a23_mem/n19219 ) );
  OR U2307 ( .A(n1019), .B(n1716), .Z(n1721) );
  AND U2308 ( .A(n1722), .B(n1723), .Z(n1720) );
  NANDN U2309 ( .B(n1093), .A(n1713), .Z(n1723) );
  NAND U2310 ( .A(n1719), .B(\u_a23_mem/p_mem[25][1] ), .Z(n1722) );
  NAND U2311 ( .A(n1724), .B(n1725), .Z(\u_a23_mem/n19218 ) );
  OR U2312 ( .A(n1025), .B(n1716), .Z(n1725) );
  AND U2313 ( .A(n1726), .B(n1727), .Z(n1724) );
  NANDN U2314 ( .B(n1098), .A(n1713), .Z(n1727) );
  NAND U2315 ( .A(n1719), .B(\u_a23_mem/p_mem[25][2] ), .Z(n1726) );
  NAND U2316 ( .A(n1728), .B(n1729), .Z(\u_a23_mem/n19217 ) );
  OR U2317 ( .A(n1031), .B(n1716), .Z(n1729) );
  AND U2318 ( .A(n1730), .B(n1731), .Z(n1728) );
  NANDN U2319 ( .B(n1103), .A(n1713), .Z(n1731) );
  NAND U2320 ( .A(n1719), .B(\u_a23_mem/p_mem[25][3] ), .Z(n1730) );
  NAND U2321 ( .A(n1732), .B(n1733), .Z(\u_a23_mem/n19216 ) );
  OR U2322 ( .A(n1037), .B(n1716), .Z(n1733) );
  AND U2323 ( .A(n1734), .B(n1735), .Z(n1732) );
  NANDN U2324 ( .B(n1108), .A(n1713), .Z(n1735) );
  NAND U2325 ( .A(n1719), .B(\u_a23_mem/p_mem[25][4] ), .Z(n1734) );
  NAND U2326 ( .A(n1736), .B(n1737), .Z(\u_a23_mem/n19215 ) );
  OR U2327 ( .A(n1043), .B(n1716), .Z(n1737) );
  AND U2328 ( .A(n1738), .B(n1739), .Z(n1736) );
  NANDN U2329 ( .B(n1113), .A(n1713), .Z(n1739) );
  NAND U2330 ( .A(n1719), .B(\u_a23_mem/p_mem[25][5] ), .Z(n1738) );
  NAND U2331 ( .A(n1740), .B(n1741), .Z(\u_a23_mem/n19214 ) );
  OR U2332 ( .A(n1049), .B(n1716), .Z(n1741) );
  AND U2333 ( .A(n1742), .B(n1743), .Z(n1740) );
  NANDN U2334 ( .B(n1118), .A(n1713), .Z(n1743) );
  NAND U2335 ( .A(n1719), .B(\u_a23_mem/p_mem[25][6] ), .Z(n1742) );
  NAND U2336 ( .A(n1744), .B(n1745), .Z(\u_a23_mem/n19213 ) );
  NANDN U2337 ( .B(n1716), .A(n1055), .Z(n1745) );
  NAND U2338 ( .A(n1121), .B(n1713), .Z(n1716) );
  AND U2339 ( .A(n1746), .B(n1747), .Z(n1744) );
  NANDN U2340 ( .B(n1124), .A(n1713), .Z(n1747) );
  NAND U2341 ( .A(n1719), .B(\u_a23_mem/p_mem[25][7] ), .Z(n1746) );
  NANDN U2342 ( .B(n1125), .A(n1713), .Z(n1719) );
  NAND U2343 ( .A(n1748), .B(n1749), .Z(\u_a23_mem/n19212 ) );
  OR U2344 ( .A(n1011), .B(n1750), .Z(n1749) );
  AND U2345 ( .A(n1751), .B(n1752), .Z(n1748) );
  NANDN U2346 ( .B(n1131), .A(n1713), .Z(n1752) );
  NAND U2347 ( .A(n1753), .B(\u_a23_mem/p_mem[26][0] ), .Z(n1751) );
  NAND U2348 ( .A(n1754), .B(n1755), .Z(\u_a23_mem/n19211 ) );
  OR U2349 ( .A(n1019), .B(n1750), .Z(n1755) );
  AND U2350 ( .A(n1756), .B(n1757), .Z(n1754) );
  NANDN U2351 ( .B(n1137), .A(n1713), .Z(n1757) );
  NAND U2352 ( .A(n1753), .B(\u_a23_mem/p_mem[26][1] ), .Z(n1756) );
  NAND U2353 ( .A(n1758), .B(n1759), .Z(\u_a23_mem/n19210 ) );
  OR U2354 ( .A(n1025), .B(n1750), .Z(n1759) );
  AND U2355 ( .A(n1760), .B(n1761), .Z(n1758) );
  NANDN U2356 ( .B(n1142), .A(n1713), .Z(n1761) );
  NAND U2357 ( .A(n1753), .B(\u_a23_mem/p_mem[26][2] ), .Z(n1760) );
  NAND U2358 ( .A(n1762), .B(n1763), .Z(\u_a23_mem/n19209 ) );
  OR U2359 ( .A(n1031), .B(n1750), .Z(n1763) );
  AND U2360 ( .A(n1764), .B(n1765), .Z(n1762) );
  NANDN U2361 ( .B(n1147), .A(n1713), .Z(n1765) );
  NAND U2362 ( .A(n1753), .B(\u_a23_mem/p_mem[26][3] ), .Z(n1764) );
  NAND U2363 ( .A(n1766), .B(n1767), .Z(\u_a23_mem/n19208 ) );
  OR U2364 ( .A(n1037), .B(n1750), .Z(n1767) );
  AND U2365 ( .A(n1768), .B(n1769), .Z(n1766) );
  NANDN U2366 ( .B(n1152), .A(n1713), .Z(n1769) );
  NAND U2367 ( .A(n1753), .B(\u_a23_mem/p_mem[26][4] ), .Z(n1768) );
  NAND U2368 ( .A(n1770), .B(n1771), .Z(\u_a23_mem/n19207 ) );
  OR U2369 ( .A(n1043), .B(n1750), .Z(n1771) );
  AND U2370 ( .A(n1772), .B(n1773), .Z(n1770) );
  NANDN U2371 ( .B(n1157), .A(n1713), .Z(n1773) );
  NAND U2372 ( .A(n1753), .B(\u_a23_mem/p_mem[26][5] ), .Z(n1772) );
  NAND U2373 ( .A(n1774), .B(n1775), .Z(\u_a23_mem/n19206 ) );
  OR U2374 ( .A(n1049), .B(n1750), .Z(n1775) );
  AND U2375 ( .A(n1776), .B(n1777), .Z(n1774) );
  NANDN U2376 ( .B(n1162), .A(n1713), .Z(n1777) );
  NAND U2377 ( .A(n1753), .B(\u_a23_mem/p_mem[26][6] ), .Z(n1776) );
  NAND U2378 ( .A(n1778), .B(n1779), .Z(\u_a23_mem/n19205 ) );
  NANDN U2379 ( .B(n1750), .A(n1055), .Z(n1779) );
  NAND U2380 ( .A(n1165), .B(n1713), .Z(n1750) );
  AND U2381 ( .A(n1780), .B(n1781), .Z(n1778) );
  NANDN U2382 ( .B(n1168), .A(n1713), .Z(n1781) );
  NAND U2383 ( .A(n1753), .B(\u_a23_mem/p_mem[26][7] ), .Z(n1780) );
  NANDN U2384 ( .B(n1169), .A(n1713), .Z(n1753) );
  NAND U2385 ( .A(n1782), .B(n1783), .Z(\u_a23_mem/n19204 ) );
  OR U2386 ( .A(n1011), .B(n1784), .Z(n1783) );
  AND U2387 ( .A(n1785), .B(n1786), .Z(n1782) );
  NAND U2388 ( .A(n1787), .B(\u_a23_mem/p_mem[27][0] ), .Z(n1786) );
  NANDN U2389 ( .B(n1015), .A(n1713), .Z(n1785) );
  NAND U2390 ( .A(n1788), .B(n1789), .Z(\u_a23_mem/n19203 ) );
  OR U2391 ( .A(n1019), .B(n1784), .Z(n1789) );
  AND U2392 ( .A(n1790), .B(n1791), .Z(n1788) );
  NAND U2393 ( .A(n1787), .B(\u_a23_mem/p_mem[27][1] ), .Z(n1791) );
  NANDN U2394 ( .B(n1022), .A(n1713), .Z(n1790) );
  NAND U2395 ( .A(n1792), .B(n1793), .Z(\u_a23_mem/n19202 ) );
  OR U2396 ( .A(n1025), .B(n1784), .Z(n1793) );
  AND U2397 ( .A(n1794), .B(n1795), .Z(n1792) );
  NAND U2398 ( .A(n1787), .B(\u_a23_mem/p_mem[27][2] ), .Z(n1795) );
  NANDN U2399 ( .B(n1028), .A(n1713), .Z(n1794) );
  NAND U2400 ( .A(n1796), .B(n1797), .Z(\u_a23_mem/n19201 ) );
  OR U2401 ( .A(n1031), .B(n1784), .Z(n1797) );
  AND U2402 ( .A(n1798), .B(n1799), .Z(n1796) );
  NAND U2403 ( .A(n1787), .B(\u_a23_mem/p_mem[27][3] ), .Z(n1799) );
  NANDN U2404 ( .B(n1034), .A(n1713), .Z(n1798) );
  NAND U2405 ( .A(n1800), .B(n1801), .Z(\u_a23_mem/n19200 ) );
  OR U2406 ( .A(n1037), .B(n1784), .Z(n1801) );
  AND U2407 ( .A(n1802), .B(n1803), .Z(n1800) );
  NAND U2408 ( .A(n1787), .B(\u_a23_mem/p_mem[27][4] ), .Z(n1803) );
  NANDN U2409 ( .B(n1040), .A(n1713), .Z(n1802) );
  NAND U2410 ( .A(n1804), .B(n1805), .Z(\u_a23_mem/n19199 ) );
  OR U2411 ( .A(n1043), .B(n1784), .Z(n1805) );
  AND U2412 ( .A(n1806), .B(n1807), .Z(n1804) );
  NAND U2413 ( .A(n1787), .B(\u_a23_mem/p_mem[27][5] ), .Z(n1807) );
  NANDN U2414 ( .B(n1046), .A(n1713), .Z(n1806) );
  NAND U2415 ( .A(n1808), .B(n1809), .Z(\u_a23_mem/n19198 ) );
  OR U2416 ( .A(n1049), .B(n1784), .Z(n1809) );
  AND U2417 ( .A(n1810), .B(n1811), .Z(n1808) );
  NAND U2418 ( .A(n1787), .B(\u_a23_mem/p_mem[27][6] ), .Z(n1811) );
  NANDN U2419 ( .B(n1052), .A(n1713), .Z(n1810) );
  NAND U2420 ( .A(n1812), .B(n1813), .Z(\u_a23_mem/n19197 ) );
  NANDN U2421 ( .B(n1784), .A(n1055), .Z(n1813) );
  NAND U2422 ( .A(n1056), .B(n1713), .Z(n1784) );
  AND U2423 ( .A(n1814), .B(n1815), .Z(n1812) );
  NAND U2424 ( .A(n1787), .B(\u_a23_mem/p_mem[27][7] ), .Z(n1815) );
  NANDN U2425 ( .B(n1059), .A(n1713), .Z(n1787) );
  NAND U2426 ( .A(n1061), .B(n1713), .Z(n1814) );
  ANDN U2427 ( .A(n1816), .B(n1572), .Z(n1713) );
  NAND U2428 ( .A(n1817), .B(n1818), .Z(\u_a23_mem/n19196 ) );
  NAND U2429 ( .A(n1819), .B(\u_a23_mem/p_mem[28][0] ), .Z(n1818) );
  OR U2430 ( .A(n1011), .B(n1820), .Z(n1817) );
  NAND U2431 ( .A(n1821), .B(n1822), .Z(\u_a23_mem/n19195 ) );
  NAND U2432 ( .A(n1819), .B(\u_a23_mem/p_mem[28][1] ), .Z(n1822) );
  OR U2433 ( .A(n1019), .B(n1820), .Z(n1821) );
  NAND U2434 ( .A(n1823), .B(n1824), .Z(\u_a23_mem/n19194 ) );
  NAND U2435 ( .A(n1819), .B(\u_a23_mem/p_mem[28][2] ), .Z(n1824) );
  OR U2436 ( .A(n1025), .B(n1820), .Z(n1823) );
  NAND U2437 ( .A(n1825), .B(n1826), .Z(\u_a23_mem/n19193 ) );
  NAND U2438 ( .A(n1819), .B(\u_a23_mem/p_mem[28][3] ), .Z(n1826) );
  OR U2439 ( .A(n1031), .B(n1820), .Z(n1825) );
  NAND U2440 ( .A(n1827), .B(n1828), .Z(\u_a23_mem/n19192 ) );
  NAND U2441 ( .A(n1819), .B(\u_a23_mem/p_mem[28][4] ), .Z(n1828) );
  OR U2442 ( .A(n1037), .B(n1820), .Z(n1827) );
  NAND U2443 ( .A(n1829), .B(n1830), .Z(\u_a23_mem/n19191 ) );
  NAND U2444 ( .A(n1819), .B(\u_a23_mem/p_mem[28][5] ), .Z(n1830) );
  OR U2445 ( .A(n1043), .B(n1820), .Z(n1829) );
  NAND U2446 ( .A(n1831), .B(n1832), .Z(\u_a23_mem/n19190 ) );
  NAND U2447 ( .A(n1819), .B(\u_a23_mem/p_mem[28][6] ), .Z(n1832) );
  OR U2448 ( .A(n1049), .B(n1820), .Z(n1831) );
  NAND U2449 ( .A(n1833), .B(n1834), .Z(\u_a23_mem/n19189 ) );
  NAND U2450 ( .A(n1819), .B(\u_a23_mem/p_mem[28][7] ), .Z(n1834) );
  NANDN U2451 ( .B(n1080), .A(n1835), .Z(n1819) );
  NANDN U2452 ( .B(n1820), .A(n1055), .Z(n1833) );
  NANDN U2453 ( .B(n2), .A(n1835), .Z(n1820) );
  NAND U2454 ( .A(n1836), .B(n1837), .Z(\u_a23_mem/n19188 ) );
  OR U2455 ( .A(n1011), .B(n1838), .Z(n1837) );
  AND U2456 ( .A(n1839), .B(n1840), .Z(n1836) );
  NANDN U2457 ( .B(n1087), .A(n1835), .Z(n1840) );
  NAND U2458 ( .A(n1841), .B(\u_a23_mem/p_mem[29][0] ), .Z(n1839) );
  NAND U2459 ( .A(n1842), .B(n1843), .Z(\u_a23_mem/n19187 ) );
  OR U2460 ( .A(n1019), .B(n1838), .Z(n1843) );
  AND U2461 ( .A(n1844), .B(n1845), .Z(n1842) );
  NANDN U2462 ( .B(n1093), .A(n1835), .Z(n1845) );
  NAND U2463 ( .A(n1841), .B(\u_a23_mem/p_mem[29][1] ), .Z(n1844) );
  NAND U2464 ( .A(n1846), .B(n1847), .Z(\u_a23_mem/n19186 ) );
  OR U2465 ( .A(n1025), .B(n1838), .Z(n1847) );
  AND U2466 ( .A(n1848), .B(n1849), .Z(n1846) );
  NANDN U2467 ( .B(n1098), .A(n1835), .Z(n1849) );
  NAND U2468 ( .A(n1841), .B(\u_a23_mem/p_mem[29][2] ), .Z(n1848) );
  NAND U2469 ( .A(n1850), .B(n1851), .Z(\u_a23_mem/n19185 ) );
  OR U2470 ( .A(n1031), .B(n1838), .Z(n1851) );
  AND U2471 ( .A(n1852), .B(n1853), .Z(n1850) );
  NANDN U2472 ( .B(n1103), .A(n1835), .Z(n1853) );
  NAND U2473 ( .A(n1841), .B(\u_a23_mem/p_mem[29][3] ), .Z(n1852) );
  NAND U2474 ( .A(n1854), .B(n1855), .Z(\u_a23_mem/n19184 ) );
  OR U2475 ( .A(n1037), .B(n1838), .Z(n1855) );
  AND U2476 ( .A(n1856), .B(n1857), .Z(n1854) );
  NANDN U2477 ( .B(n1108), .A(n1835), .Z(n1857) );
  NAND U2478 ( .A(n1841), .B(\u_a23_mem/p_mem[29][4] ), .Z(n1856) );
  NAND U2479 ( .A(n1858), .B(n1859), .Z(\u_a23_mem/n19183 ) );
  OR U2480 ( .A(n1043), .B(n1838), .Z(n1859) );
  AND U2481 ( .A(n1860), .B(n1861), .Z(n1858) );
  NANDN U2482 ( .B(n1113), .A(n1835), .Z(n1861) );
  NAND U2483 ( .A(n1841), .B(\u_a23_mem/p_mem[29][5] ), .Z(n1860) );
  NAND U2484 ( .A(n1862), .B(n1863), .Z(\u_a23_mem/n19182 ) );
  OR U2485 ( .A(n1049), .B(n1838), .Z(n1863) );
  AND U2486 ( .A(n1864), .B(n1865), .Z(n1862) );
  NANDN U2487 ( .B(n1118), .A(n1835), .Z(n1865) );
  NAND U2488 ( .A(n1841), .B(\u_a23_mem/p_mem[29][6] ), .Z(n1864) );
  NAND U2489 ( .A(n1866), .B(n1867), .Z(\u_a23_mem/n19181 ) );
  NANDN U2490 ( .B(n1838), .A(n1055), .Z(n1867) );
  NAND U2491 ( .A(n1121), .B(n1835), .Z(n1838) );
  AND U2492 ( .A(n1868), .B(n1869), .Z(n1866) );
  NANDN U2493 ( .B(n1124), .A(n1835), .Z(n1869) );
  NAND U2494 ( .A(n1841), .B(\u_a23_mem/p_mem[29][7] ), .Z(n1868) );
  NANDN U2495 ( .B(n1125), .A(n1835), .Z(n1841) );
  NAND U2496 ( .A(n1870), .B(n1871), .Z(\u_a23_mem/n19180 ) );
  OR U2497 ( .A(n1011), .B(n1872), .Z(n1871) );
  AND U2498 ( .A(n1873), .B(n1874), .Z(n1870) );
  NANDN U2499 ( .B(n1131), .A(n1835), .Z(n1874) );
  NAND U2500 ( .A(n1875), .B(\u_a23_mem/p_mem[30][0] ), .Z(n1873) );
  NAND U2501 ( .A(n1876), .B(n1877), .Z(\u_a23_mem/n19179 ) );
  OR U2502 ( .A(n1019), .B(n1872), .Z(n1877) );
  AND U2503 ( .A(n1878), .B(n1879), .Z(n1876) );
  NANDN U2504 ( .B(n1137), .A(n1835), .Z(n1879) );
  NAND U2505 ( .A(n1875), .B(\u_a23_mem/p_mem[30][1] ), .Z(n1878) );
  NAND U2506 ( .A(n1880), .B(n1881), .Z(\u_a23_mem/n19178 ) );
  OR U2507 ( .A(n1025), .B(n1872), .Z(n1881) );
  AND U2508 ( .A(n1882), .B(n1883), .Z(n1880) );
  NANDN U2509 ( .B(n1142), .A(n1835), .Z(n1883) );
  NAND U2510 ( .A(n1875), .B(\u_a23_mem/p_mem[30][2] ), .Z(n1882) );
  NAND U2511 ( .A(n1884), .B(n1885), .Z(\u_a23_mem/n19177 ) );
  OR U2512 ( .A(n1031), .B(n1872), .Z(n1885) );
  AND U2513 ( .A(n1886), .B(n1887), .Z(n1884) );
  NANDN U2514 ( .B(n1147), .A(n1835), .Z(n1887) );
  NAND U2515 ( .A(n1875), .B(\u_a23_mem/p_mem[30][3] ), .Z(n1886) );
  NAND U2516 ( .A(n1888), .B(n1889), .Z(\u_a23_mem/n19176 ) );
  OR U2517 ( .A(n1037), .B(n1872), .Z(n1889) );
  AND U2518 ( .A(n1890), .B(n1891), .Z(n1888) );
  NANDN U2519 ( .B(n1152), .A(n1835), .Z(n1891) );
  NAND U2520 ( .A(n1875), .B(\u_a23_mem/p_mem[30][4] ), .Z(n1890) );
  NAND U2521 ( .A(n1892), .B(n1893), .Z(\u_a23_mem/n19175 ) );
  OR U2522 ( .A(n1043), .B(n1872), .Z(n1893) );
  AND U2523 ( .A(n1894), .B(n1895), .Z(n1892) );
  NANDN U2524 ( .B(n1157), .A(n1835), .Z(n1895) );
  NAND U2525 ( .A(n1875), .B(\u_a23_mem/p_mem[30][5] ), .Z(n1894) );
  NAND U2526 ( .A(n1896), .B(n1897), .Z(\u_a23_mem/n19174 ) );
  OR U2527 ( .A(n1049), .B(n1872), .Z(n1897) );
  AND U2528 ( .A(n1898), .B(n1899), .Z(n1896) );
  NANDN U2529 ( .B(n1162), .A(n1835), .Z(n1899) );
  NAND U2530 ( .A(n1875), .B(\u_a23_mem/p_mem[30][6] ), .Z(n1898) );
  NAND U2531 ( .A(n1900), .B(n1901), .Z(\u_a23_mem/n19173 ) );
  NANDN U2532 ( .B(n1872), .A(n1055), .Z(n1901) );
  NAND U2533 ( .A(n1165), .B(n1835), .Z(n1872) );
  AND U2534 ( .A(n1902), .B(n1903), .Z(n1900) );
  NANDN U2535 ( .B(n1168), .A(n1835), .Z(n1903) );
  NAND U2536 ( .A(n1875), .B(\u_a23_mem/p_mem[30][7] ), .Z(n1902) );
  NANDN U2537 ( .B(n1169), .A(n1835), .Z(n1875) );
  NAND U2538 ( .A(n1904), .B(n1905), .Z(\u_a23_mem/n19172 ) );
  OR U2539 ( .A(n1011), .B(n1906), .Z(n1905) );
  AND U2540 ( .A(n1907), .B(n1908), .Z(n1904) );
  NAND U2541 ( .A(n1909), .B(\u_a23_mem/p_mem[31][0] ), .Z(n1908) );
  NANDN U2542 ( .B(n1015), .A(n1835), .Z(n1907) );
  NAND U2543 ( .A(n1910), .B(n1911), .Z(\u_a23_mem/n19171 ) );
  OR U2544 ( .A(n1019), .B(n1906), .Z(n1911) );
  AND U2545 ( .A(n1912), .B(n1913), .Z(n1910) );
  NAND U2546 ( .A(n1909), .B(\u_a23_mem/p_mem[31][1] ), .Z(n1913) );
  NANDN U2547 ( .B(n1022), .A(n1835), .Z(n1912) );
  NAND U2548 ( .A(n1914), .B(n1915), .Z(\u_a23_mem/n19170 ) );
  OR U2549 ( .A(n1025), .B(n1906), .Z(n1915) );
  AND U2550 ( .A(n1916), .B(n1917), .Z(n1914) );
  NAND U2551 ( .A(n1909), .B(\u_a23_mem/p_mem[31][2] ), .Z(n1917) );
  NANDN U2552 ( .B(n1028), .A(n1835), .Z(n1916) );
  NAND U2553 ( .A(n1918), .B(n1919), .Z(\u_a23_mem/n19169 ) );
  OR U2554 ( .A(n1031), .B(n1906), .Z(n1919) );
  AND U2555 ( .A(n1920), .B(n1921), .Z(n1918) );
  NAND U2556 ( .A(n1909), .B(\u_a23_mem/p_mem[31][3] ), .Z(n1921) );
  NANDN U2557 ( .B(n1034), .A(n1835), .Z(n1920) );
  NAND U2558 ( .A(n1922), .B(n1923), .Z(\u_a23_mem/n19168 ) );
  OR U2559 ( .A(n1037), .B(n1906), .Z(n1923) );
  AND U2560 ( .A(n1924), .B(n1925), .Z(n1922) );
  NAND U2561 ( .A(n1909), .B(\u_a23_mem/p_mem[31][4] ), .Z(n1925) );
  NANDN U2562 ( .B(n1040), .A(n1835), .Z(n1924) );
  NAND U2563 ( .A(n1926), .B(n1927), .Z(\u_a23_mem/n19167 ) );
  OR U2564 ( .A(n1043), .B(n1906), .Z(n1927) );
  AND U2565 ( .A(n1928), .B(n1929), .Z(n1926) );
  NAND U2566 ( .A(n1909), .B(\u_a23_mem/p_mem[31][5] ), .Z(n1929) );
  NANDN U2567 ( .B(n1046), .A(n1835), .Z(n1928) );
  NAND U2568 ( .A(n1930), .B(n1931), .Z(\u_a23_mem/n19166 ) );
  OR U2569 ( .A(n1049), .B(n1906), .Z(n1931) );
  AND U2570 ( .A(n1932), .B(n1933), .Z(n1930) );
  NAND U2571 ( .A(n1909), .B(\u_a23_mem/p_mem[31][6] ), .Z(n1933) );
  NANDN U2572 ( .B(n1052), .A(n1835), .Z(n1932) );
  NAND U2573 ( .A(n1934), .B(n1935), .Z(\u_a23_mem/n19165 ) );
  NANDN U2574 ( .B(n1906), .A(n1055), .Z(n1935) );
  NAND U2575 ( .A(n1056), .B(n1835), .Z(n1906) );
  AND U2576 ( .A(n1936), .B(n1937), .Z(n1934) );
  NAND U2577 ( .A(n1909), .B(\u_a23_mem/p_mem[31][7] ), .Z(n1937) );
  NANDN U2578 ( .B(n1059), .A(n1835), .Z(n1909) );
  NAND U2579 ( .A(n1061), .B(n1835), .Z(n1936) );
  NOR U2580 ( .A(n1938), .B(n1572), .Z(n1835) );
  NANDN U2581 ( .B(n1939), .A(n1940), .Z(n1572) );
  NAND U2582 ( .A(n1941), .B(n1942), .Z(\u_a23_mem/n19164 ) );
  NAND U2583 ( .A(n1943), .B(\u_a23_mem/p_mem[32][0] ), .Z(n1942) );
  OR U2584 ( .A(n1011), .B(n1944), .Z(n1941) );
  NAND U2585 ( .A(n1945), .B(n1946), .Z(\u_a23_mem/n19163 ) );
  NAND U2586 ( .A(n1943), .B(\u_a23_mem/p_mem[32][1] ), .Z(n1946) );
  OR U2587 ( .A(n1019), .B(n1944), .Z(n1945) );
  NAND U2588 ( .A(n1947), .B(n1948), .Z(\u_a23_mem/n19162 ) );
  NAND U2589 ( .A(n1943), .B(\u_a23_mem/p_mem[32][2] ), .Z(n1948) );
  OR U2590 ( .A(n1025), .B(n1944), .Z(n1947) );
  NAND U2591 ( .A(n1949), .B(n1950), .Z(\u_a23_mem/n19161 ) );
  NAND U2592 ( .A(n1943), .B(\u_a23_mem/p_mem[32][3] ), .Z(n1950) );
  OR U2593 ( .A(n1031), .B(n1944), .Z(n1949) );
  NAND U2594 ( .A(n1951), .B(n1952), .Z(\u_a23_mem/n19160 ) );
  NAND U2595 ( .A(n1943), .B(\u_a23_mem/p_mem[32][4] ), .Z(n1952) );
  OR U2596 ( .A(n1037), .B(n1944), .Z(n1951) );
  NAND U2597 ( .A(n1953), .B(n1954), .Z(\u_a23_mem/n19159 ) );
  NAND U2598 ( .A(n1943), .B(\u_a23_mem/p_mem[32][5] ), .Z(n1954) );
  OR U2599 ( .A(n1043), .B(n1944), .Z(n1953) );
  NAND U2600 ( .A(n1955), .B(n1956), .Z(\u_a23_mem/n19158 ) );
  NAND U2601 ( .A(n1943), .B(\u_a23_mem/p_mem[32][6] ), .Z(n1956) );
  OR U2602 ( .A(n1049), .B(n1944), .Z(n1955) );
  NAND U2603 ( .A(n1957), .B(n1958), .Z(\u_a23_mem/n19157 ) );
  NAND U2604 ( .A(n1943), .B(\u_a23_mem/p_mem[32][7] ), .Z(n1958) );
  NANDN U2605 ( .B(n1080), .A(n1959), .Z(n1943) );
  NANDN U2606 ( .B(n1944), .A(n1055), .Z(n1957) );
  NANDN U2607 ( .B(n2), .A(n1959), .Z(n1944) );
  NAND U2608 ( .A(n1960), .B(n1961), .Z(\u_a23_mem/n19156 ) );
  OR U2609 ( .A(n1011), .B(n1962), .Z(n1961) );
  AND U2610 ( .A(n1963), .B(n1964), .Z(n1960) );
  NANDN U2611 ( .B(n1087), .A(n1959), .Z(n1964) );
  NAND U2612 ( .A(n1965), .B(\u_a23_mem/p_mem[33][0] ), .Z(n1963) );
  NAND U2613 ( .A(n1966), .B(n1967), .Z(\u_a23_mem/n19155 ) );
  OR U2614 ( .A(n1019), .B(n1962), .Z(n1967) );
  AND U2615 ( .A(n1968), .B(n1969), .Z(n1966) );
  NANDN U2616 ( .B(n1093), .A(n1959), .Z(n1969) );
  NAND U2617 ( .A(n1965), .B(\u_a23_mem/p_mem[33][1] ), .Z(n1968) );
  NAND U2618 ( .A(n1970), .B(n1971), .Z(\u_a23_mem/n19154 ) );
  OR U2619 ( .A(n1025), .B(n1962), .Z(n1971) );
  AND U2620 ( .A(n1972), .B(n1973), .Z(n1970) );
  NANDN U2621 ( .B(n1098), .A(n1959), .Z(n1973) );
  NAND U2622 ( .A(n1965), .B(\u_a23_mem/p_mem[33][2] ), .Z(n1972) );
  NAND U2623 ( .A(n1974), .B(n1975), .Z(\u_a23_mem/n19153 ) );
  OR U2624 ( .A(n1031), .B(n1962), .Z(n1975) );
  AND U2625 ( .A(n1976), .B(n1977), .Z(n1974) );
  NANDN U2626 ( .B(n1103), .A(n1959), .Z(n1977) );
  NAND U2627 ( .A(n1965), .B(\u_a23_mem/p_mem[33][3] ), .Z(n1976) );
  NAND U2628 ( .A(n1978), .B(n1979), .Z(\u_a23_mem/n19152 ) );
  OR U2629 ( .A(n1037), .B(n1962), .Z(n1979) );
  AND U2630 ( .A(n1980), .B(n1981), .Z(n1978) );
  NANDN U2631 ( .B(n1108), .A(n1959), .Z(n1981) );
  NAND U2632 ( .A(n1965), .B(\u_a23_mem/p_mem[33][4] ), .Z(n1980) );
  NAND U2633 ( .A(n1982), .B(n1983), .Z(\u_a23_mem/n19151 ) );
  OR U2634 ( .A(n1043), .B(n1962), .Z(n1983) );
  AND U2635 ( .A(n1984), .B(n1985), .Z(n1982) );
  NANDN U2636 ( .B(n1113), .A(n1959), .Z(n1985) );
  NAND U2637 ( .A(n1965), .B(\u_a23_mem/p_mem[33][5] ), .Z(n1984) );
  NAND U2638 ( .A(n1986), .B(n1987), .Z(\u_a23_mem/n19150 ) );
  OR U2639 ( .A(n1049), .B(n1962), .Z(n1987) );
  AND U2640 ( .A(n1988), .B(n1989), .Z(n1986) );
  NANDN U2641 ( .B(n1118), .A(n1959), .Z(n1989) );
  NAND U2642 ( .A(n1965), .B(\u_a23_mem/p_mem[33][6] ), .Z(n1988) );
  NAND U2643 ( .A(n1990), .B(n1991), .Z(\u_a23_mem/n19149 ) );
  NANDN U2644 ( .B(n1962), .A(n1055), .Z(n1991) );
  NAND U2645 ( .A(n1121), .B(n1959), .Z(n1962) );
  AND U2646 ( .A(n1992), .B(n1993), .Z(n1990) );
  NANDN U2647 ( .B(n1124), .A(n1959), .Z(n1993) );
  NAND U2648 ( .A(n1965), .B(\u_a23_mem/p_mem[33][7] ), .Z(n1992) );
  NANDN U2649 ( .B(n1125), .A(n1959), .Z(n1965) );
  NAND U2650 ( .A(n1994), .B(n1995), .Z(\u_a23_mem/n19148 ) );
  OR U2651 ( .A(n1011), .B(n1996), .Z(n1995) );
  AND U2652 ( .A(n1997), .B(n1998), .Z(n1994) );
  NANDN U2653 ( .B(n1131), .A(n1959), .Z(n1998) );
  NAND U2654 ( .A(n1999), .B(\u_a23_mem/p_mem[34][0] ), .Z(n1997) );
  NAND U2655 ( .A(n2000), .B(n2001), .Z(\u_a23_mem/n19147 ) );
  OR U2656 ( .A(n1019), .B(n1996), .Z(n2001) );
  AND U2657 ( .A(n2002), .B(n2003), .Z(n2000) );
  NANDN U2658 ( .B(n1137), .A(n1959), .Z(n2003) );
  NAND U2659 ( .A(n1999), .B(\u_a23_mem/p_mem[34][1] ), .Z(n2002) );
  NAND U2660 ( .A(n2004), .B(n2005), .Z(\u_a23_mem/n19146 ) );
  OR U2661 ( .A(n1025), .B(n1996), .Z(n2005) );
  AND U2662 ( .A(n2006), .B(n2007), .Z(n2004) );
  NANDN U2663 ( .B(n1142), .A(n1959), .Z(n2007) );
  NAND U2664 ( .A(n1999), .B(\u_a23_mem/p_mem[34][2] ), .Z(n2006) );
  NAND U2665 ( .A(n2008), .B(n2009), .Z(\u_a23_mem/n19145 ) );
  OR U2666 ( .A(n1031), .B(n1996), .Z(n2009) );
  AND U2667 ( .A(n2010), .B(n2011), .Z(n2008) );
  NANDN U2668 ( .B(n1147), .A(n1959), .Z(n2011) );
  NAND U2669 ( .A(n1999), .B(\u_a23_mem/p_mem[34][3] ), .Z(n2010) );
  NAND U2670 ( .A(n2012), .B(n2013), .Z(\u_a23_mem/n19144 ) );
  OR U2671 ( .A(n1037), .B(n1996), .Z(n2013) );
  AND U2672 ( .A(n2014), .B(n2015), .Z(n2012) );
  NANDN U2673 ( .B(n1152), .A(n1959), .Z(n2015) );
  NAND U2674 ( .A(n1999), .B(\u_a23_mem/p_mem[34][4] ), .Z(n2014) );
  NAND U2675 ( .A(n2016), .B(n2017), .Z(\u_a23_mem/n19143 ) );
  OR U2676 ( .A(n1043), .B(n1996), .Z(n2017) );
  AND U2677 ( .A(n2018), .B(n2019), .Z(n2016) );
  NANDN U2678 ( .B(n1157), .A(n1959), .Z(n2019) );
  NAND U2679 ( .A(n1999), .B(\u_a23_mem/p_mem[34][5] ), .Z(n2018) );
  NAND U2680 ( .A(n2020), .B(n2021), .Z(\u_a23_mem/n19142 ) );
  OR U2681 ( .A(n1049), .B(n1996), .Z(n2021) );
  AND U2682 ( .A(n2022), .B(n2023), .Z(n2020) );
  NANDN U2683 ( .B(n1162), .A(n1959), .Z(n2023) );
  NAND U2684 ( .A(n1999), .B(\u_a23_mem/p_mem[34][6] ), .Z(n2022) );
  NAND U2685 ( .A(n2024), .B(n2025), .Z(\u_a23_mem/n19141 ) );
  NANDN U2686 ( .B(n1996), .A(n1055), .Z(n2025) );
  NAND U2687 ( .A(n1165), .B(n1959), .Z(n1996) );
  AND U2688 ( .A(n2026), .B(n2027), .Z(n2024) );
  NANDN U2689 ( .B(n1168), .A(n1959), .Z(n2027) );
  NAND U2690 ( .A(n1999), .B(\u_a23_mem/p_mem[34][7] ), .Z(n2026) );
  NANDN U2691 ( .B(n1169), .A(n1959), .Z(n1999) );
  NAND U2692 ( .A(n2028), .B(n2029), .Z(\u_a23_mem/n19140 ) );
  OR U2693 ( .A(n1011), .B(n2030), .Z(n2029) );
  AND U2694 ( .A(n2031), .B(n2032), .Z(n2028) );
  NAND U2695 ( .A(n2033), .B(\u_a23_mem/p_mem[35][0] ), .Z(n2032) );
  NANDN U2696 ( .B(n1015), .A(n1959), .Z(n2031) );
  NAND U2697 ( .A(n2034), .B(n2035), .Z(\u_a23_mem/n19139 ) );
  OR U2698 ( .A(n1019), .B(n2030), .Z(n2035) );
  AND U2699 ( .A(n2036), .B(n2037), .Z(n2034) );
  NAND U2700 ( .A(n2033), .B(\u_a23_mem/p_mem[35][1] ), .Z(n2037) );
  NANDN U2701 ( .B(n1022), .A(n1959), .Z(n2036) );
  NAND U2702 ( .A(n2038), .B(n2039), .Z(\u_a23_mem/n19138 ) );
  OR U2703 ( .A(n1025), .B(n2030), .Z(n2039) );
  AND U2704 ( .A(n2040), .B(n2041), .Z(n2038) );
  NAND U2705 ( .A(n2033), .B(\u_a23_mem/p_mem[35][2] ), .Z(n2041) );
  NANDN U2706 ( .B(n1028), .A(n1959), .Z(n2040) );
  NAND U2707 ( .A(n2042), .B(n2043), .Z(\u_a23_mem/n19137 ) );
  OR U2708 ( .A(n1031), .B(n2030), .Z(n2043) );
  AND U2709 ( .A(n2044), .B(n2045), .Z(n2042) );
  NAND U2710 ( .A(n2033), .B(\u_a23_mem/p_mem[35][3] ), .Z(n2045) );
  NANDN U2711 ( .B(n1034), .A(n1959), .Z(n2044) );
  NAND U2712 ( .A(n2046), .B(n2047), .Z(\u_a23_mem/n19136 ) );
  OR U2713 ( .A(n1037), .B(n2030), .Z(n2047) );
  AND U2714 ( .A(n2048), .B(n2049), .Z(n2046) );
  NAND U2715 ( .A(n2033), .B(\u_a23_mem/p_mem[35][4] ), .Z(n2049) );
  NANDN U2716 ( .B(n1040), .A(n1959), .Z(n2048) );
  NAND U2717 ( .A(n2050), .B(n2051), .Z(\u_a23_mem/n19135 ) );
  OR U2718 ( .A(n1043), .B(n2030), .Z(n2051) );
  AND U2719 ( .A(n2052), .B(n2053), .Z(n2050) );
  NAND U2720 ( .A(n2033), .B(\u_a23_mem/p_mem[35][5] ), .Z(n2053) );
  NANDN U2721 ( .B(n1046), .A(n1959), .Z(n2052) );
  NAND U2722 ( .A(n2054), .B(n2055), .Z(\u_a23_mem/n19134 ) );
  OR U2723 ( .A(n1049), .B(n2030), .Z(n2055) );
  AND U2724 ( .A(n2056), .B(n2057), .Z(n2054) );
  NAND U2725 ( .A(n2033), .B(\u_a23_mem/p_mem[35][6] ), .Z(n2057) );
  NANDN U2726 ( .B(n1052), .A(n1959), .Z(n2056) );
  NAND U2727 ( .A(n2058), .B(n2059), .Z(\u_a23_mem/n19133 ) );
  NANDN U2728 ( .B(n2030), .A(n1055), .Z(n2059) );
  NAND U2729 ( .A(n1056), .B(n1959), .Z(n2030) );
  AND U2730 ( .A(n2060), .B(n2061), .Z(n2058) );
  NAND U2731 ( .A(n2033), .B(\u_a23_mem/p_mem[35][7] ), .Z(n2061) );
  NANDN U2732 ( .B(n1059), .A(n1959), .Z(n2033) );
  NAND U2733 ( .A(n1061), .B(n1959), .Z(n2060) );
  ANDN U2734 ( .A(n1571), .B(n2062), .Z(n1959) );
  NAND U2735 ( .A(n2063), .B(n2064), .Z(\u_a23_mem/n19132 ) );
  NAND U2736 ( .A(n2065), .B(\u_a23_mem/p_mem[36][0] ), .Z(n2064) );
  OR U2737 ( .A(n1011), .B(n2066), .Z(n2063) );
  NAND U2738 ( .A(n2067), .B(n2068), .Z(\u_a23_mem/n19131 ) );
  NAND U2739 ( .A(n2065), .B(\u_a23_mem/p_mem[36][1] ), .Z(n2068) );
  OR U2740 ( .A(n1019), .B(n2066), .Z(n2067) );
  NAND U2741 ( .A(n2069), .B(n2070), .Z(\u_a23_mem/n19130 ) );
  NAND U2742 ( .A(n2065), .B(\u_a23_mem/p_mem[36][2] ), .Z(n2070) );
  OR U2743 ( .A(n1025), .B(n2066), .Z(n2069) );
  NAND U2744 ( .A(n2071), .B(n2072), .Z(\u_a23_mem/n19129 ) );
  NAND U2745 ( .A(n2065), .B(\u_a23_mem/p_mem[36][3] ), .Z(n2072) );
  OR U2746 ( .A(n1031), .B(n2066), .Z(n2071) );
  NAND U2747 ( .A(n2073), .B(n2074), .Z(\u_a23_mem/n19128 ) );
  NAND U2748 ( .A(n2065), .B(\u_a23_mem/p_mem[36][4] ), .Z(n2074) );
  OR U2749 ( .A(n1037), .B(n2066), .Z(n2073) );
  NAND U2750 ( .A(n2075), .B(n2076), .Z(\u_a23_mem/n19127 ) );
  NAND U2751 ( .A(n2065), .B(\u_a23_mem/p_mem[36][5] ), .Z(n2076) );
  OR U2752 ( .A(n1043), .B(n2066), .Z(n2075) );
  NAND U2753 ( .A(n2077), .B(n2078), .Z(\u_a23_mem/n19126 ) );
  NAND U2754 ( .A(n2065), .B(\u_a23_mem/p_mem[36][6] ), .Z(n2078) );
  OR U2755 ( .A(n1049), .B(n2066), .Z(n2077) );
  NAND U2756 ( .A(n2079), .B(n2080), .Z(\u_a23_mem/n19125 ) );
  NAND U2757 ( .A(n2065), .B(\u_a23_mem/p_mem[36][7] ), .Z(n2080) );
  NANDN U2758 ( .B(n1080), .A(n2081), .Z(n2065) );
  NANDN U2759 ( .B(n2066), .A(n1055), .Z(n2079) );
  NANDN U2760 ( .B(n2), .A(n2081), .Z(n2066) );
  NAND U2761 ( .A(n2082), .B(n2083), .Z(\u_a23_mem/n19124 ) );
  OR U2762 ( .A(n1011), .B(n2084), .Z(n2083) );
  AND U2763 ( .A(n2085), .B(n2086), .Z(n2082) );
  NANDN U2764 ( .B(n1087), .A(n2081), .Z(n2086) );
  NAND U2765 ( .A(n2087), .B(\u_a23_mem/p_mem[37][0] ), .Z(n2085) );
  NAND U2766 ( .A(n2088), .B(n2089), .Z(\u_a23_mem/n19123 ) );
  OR U2767 ( .A(n1019), .B(n2084), .Z(n2089) );
  AND U2768 ( .A(n2090), .B(n2091), .Z(n2088) );
  NANDN U2769 ( .B(n1093), .A(n2081), .Z(n2091) );
  NAND U2770 ( .A(n2087), .B(\u_a23_mem/p_mem[37][1] ), .Z(n2090) );
  NAND U2771 ( .A(n2092), .B(n2093), .Z(\u_a23_mem/n19122 ) );
  OR U2772 ( .A(n1025), .B(n2084), .Z(n2093) );
  AND U2773 ( .A(n2094), .B(n2095), .Z(n2092) );
  NANDN U2774 ( .B(n1098), .A(n2081), .Z(n2095) );
  NAND U2775 ( .A(n2087), .B(\u_a23_mem/p_mem[37][2] ), .Z(n2094) );
  NAND U2776 ( .A(n2096), .B(n2097), .Z(\u_a23_mem/n19121 ) );
  OR U2777 ( .A(n1031), .B(n2084), .Z(n2097) );
  AND U2778 ( .A(n2098), .B(n2099), .Z(n2096) );
  NANDN U2779 ( .B(n1103), .A(n2081), .Z(n2099) );
  NAND U2780 ( .A(n2087), .B(\u_a23_mem/p_mem[37][3] ), .Z(n2098) );
  NAND U2781 ( .A(n2100), .B(n2101), .Z(\u_a23_mem/n19120 ) );
  OR U2782 ( .A(n1037), .B(n2084), .Z(n2101) );
  AND U2783 ( .A(n2102), .B(n2103), .Z(n2100) );
  NANDN U2784 ( .B(n1108), .A(n2081), .Z(n2103) );
  NAND U2785 ( .A(n2087), .B(\u_a23_mem/p_mem[37][4] ), .Z(n2102) );
  NAND U2786 ( .A(n2104), .B(n2105), .Z(\u_a23_mem/n19119 ) );
  OR U2787 ( .A(n1043), .B(n2084), .Z(n2105) );
  AND U2788 ( .A(n2106), .B(n2107), .Z(n2104) );
  NANDN U2789 ( .B(n1113), .A(n2081), .Z(n2107) );
  NAND U2790 ( .A(n2087), .B(\u_a23_mem/p_mem[37][5] ), .Z(n2106) );
  NAND U2791 ( .A(n2108), .B(n2109), .Z(\u_a23_mem/n19118 ) );
  OR U2792 ( .A(n1049), .B(n2084), .Z(n2109) );
  AND U2793 ( .A(n2110), .B(n2111), .Z(n2108) );
  NANDN U2794 ( .B(n1118), .A(n2081), .Z(n2111) );
  NAND U2795 ( .A(n2087), .B(\u_a23_mem/p_mem[37][6] ), .Z(n2110) );
  NAND U2796 ( .A(n2112), .B(n2113), .Z(\u_a23_mem/n19117 ) );
  NANDN U2797 ( .B(n2084), .A(n1055), .Z(n2113) );
  NAND U2798 ( .A(n1121), .B(n2081), .Z(n2084) );
  AND U2799 ( .A(n2114), .B(n2115), .Z(n2112) );
  NANDN U2800 ( .B(n1124), .A(n2081), .Z(n2115) );
  NAND U2801 ( .A(n2087), .B(\u_a23_mem/p_mem[37][7] ), .Z(n2114) );
  NANDN U2802 ( .B(n1125), .A(n2081), .Z(n2087) );
  NAND U2803 ( .A(n2116), .B(n2117), .Z(\u_a23_mem/n19116 ) );
  OR U2804 ( .A(n1011), .B(n2118), .Z(n2117) );
  AND U2805 ( .A(n2119), .B(n2120), .Z(n2116) );
  NANDN U2806 ( .B(n1131), .A(n2081), .Z(n2120) );
  NAND U2807 ( .A(n2121), .B(\u_a23_mem/p_mem[38][0] ), .Z(n2119) );
  NAND U2808 ( .A(n2122), .B(n2123), .Z(\u_a23_mem/n19115 ) );
  OR U2809 ( .A(n1019), .B(n2118), .Z(n2123) );
  AND U2810 ( .A(n2124), .B(n2125), .Z(n2122) );
  NANDN U2811 ( .B(n1137), .A(n2081), .Z(n2125) );
  NAND U2812 ( .A(n2121), .B(\u_a23_mem/p_mem[38][1] ), .Z(n2124) );
  NAND U2813 ( .A(n2126), .B(n2127), .Z(\u_a23_mem/n19114 ) );
  OR U2814 ( .A(n1025), .B(n2118), .Z(n2127) );
  AND U2815 ( .A(n2128), .B(n2129), .Z(n2126) );
  NANDN U2816 ( .B(n1142), .A(n2081), .Z(n2129) );
  NAND U2817 ( .A(n2121), .B(\u_a23_mem/p_mem[38][2] ), .Z(n2128) );
  NAND U2818 ( .A(n2130), .B(n2131), .Z(\u_a23_mem/n19113 ) );
  OR U2819 ( .A(n1031), .B(n2118), .Z(n2131) );
  AND U2820 ( .A(n2132), .B(n2133), .Z(n2130) );
  NANDN U2821 ( .B(n1147), .A(n2081), .Z(n2133) );
  NAND U2822 ( .A(n2121), .B(\u_a23_mem/p_mem[38][3] ), .Z(n2132) );
  NAND U2823 ( .A(n2134), .B(n2135), .Z(\u_a23_mem/n19112 ) );
  OR U2824 ( .A(n1037), .B(n2118), .Z(n2135) );
  AND U2825 ( .A(n2136), .B(n2137), .Z(n2134) );
  NANDN U2826 ( .B(n1152), .A(n2081), .Z(n2137) );
  NAND U2827 ( .A(n2121), .B(\u_a23_mem/p_mem[38][4] ), .Z(n2136) );
  NAND U2828 ( .A(n2138), .B(n2139), .Z(\u_a23_mem/n19111 ) );
  OR U2829 ( .A(n1043), .B(n2118), .Z(n2139) );
  AND U2830 ( .A(n2140), .B(n2141), .Z(n2138) );
  NANDN U2831 ( .B(n1157), .A(n2081), .Z(n2141) );
  NAND U2832 ( .A(n2121), .B(\u_a23_mem/p_mem[38][5] ), .Z(n2140) );
  NAND U2833 ( .A(n2142), .B(n2143), .Z(\u_a23_mem/n19110 ) );
  OR U2834 ( .A(n1049), .B(n2118), .Z(n2143) );
  AND U2835 ( .A(n2144), .B(n2145), .Z(n2142) );
  NANDN U2836 ( .B(n1162), .A(n2081), .Z(n2145) );
  NAND U2837 ( .A(n2121), .B(\u_a23_mem/p_mem[38][6] ), .Z(n2144) );
  NAND U2838 ( .A(n2146), .B(n2147), .Z(\u_a23_mem/n19109 ) );
  NANDN U2839 ( .B(n2118), .A(n1055), .Z(n2147) );
  NAND U2840 ( .A(n1165), .B(n2081), .Z(n2118) );
  AND U2841 ( .A(n2148), .B(n2149), .Z(n2146) );
  NANDN U2842 ( .B(n1168), .A(n2081), .Z(n2149) );
  NAND U2843 ( .A(n2121), .B(\u_a23_mem/p_mem[38][7] ), .Z(n2148) );
  NANDN U2844 ( .B(n1169), .A(n2081), .Z(n2121) );
  NAND U2845 ( .A(n2150), .B(n2151), .Z(\u_a23_mem/n19108 ) );
  OR U2846 ( .A(n1011), .B(n2152), .Z(n2151) );
  AND U2847 ( .A(n2153), .B(n2154), .Z(n2150) );
  NAND U2848 ( .A(n2155), .B(\u_a23_mem/p_mem[39][0] ), .Z(n2154) );
  NANDN U2849 ( .B(n1015), .A(n2081), .Z(n2153) );
  NAND U2850 ( .A(n2156), .B(n2157), .Z(\u_a23_mem/n19107 ) );
  OR U2851 ( .A(n1019), .B(n2152), .Z(n2157) );
  AND U2852 ( .A(n2158), .B(n2159), .Z(n2156) );
  NAND U2853 ( .A(n2155), .B(\u_a23_mem/p_mem[39][1] ), .Z(n2159) );
  NANDN U2854 ( .B(n1022), .A(n2081), .Z(n2158) );
  NAND U2855 ( .A(n2160), .B(n2161), .Z(\u_a23_mem/n19106 ) );
  OR U2856 ( .A(n1025), .B(n2152), .Z(n2161) );
  AND U2857 ( .A(n2162), .B(n2163), .Z(n2160) );
  NAND U2858 ( .A(n2155), .B(\u_a23_mem/p_mem[39][2] ), .Z(n2163) );
  NANDN U2859 ( .B(n1028), .A(n2081), .Z(n2162) );
  NAND U2860 ( .A(n2164), .B(n2165), .Z(\u_a23_mem/n19105 ) );
  OR U2861 ( .A(n1031), .B(n2152), .Z(n2165) );
  AND U2862 ( .A(n2166), .B(n2167), .Z(n2164) );
  NAND U2863 ( .A(n2155), .B(\u_a23_mem/p_mem[39][3] ), .Z(n2167) );
  NANDN U2864 ( .B(n1034), .A(n2081), .Z(n2166) );
  NAND U2865 ( .A(n2168), .B(n2169), .Z(\u_a23_mem/n19104 ) );
  OR U2866 ( .A(n1037), .B(n2152), .Z(n2169) );
  AND U2867 ( .A(n2170), .B(n2171), .Z(n2168) );
  NAND U2868 ( .A(n2155), .B(\u_a23_mem/p_mem[39][4] ), .Z(n2171) );
  NANDN U2869 ( .B(n1040), .A(n2081), .Z(n2170) );
  NAND U2870 ( .A(n2172), .B(n2173), .Z(\u_a23_mem/n19103 ) );
  OR U2871 ( .A(n1043), .B(n2152), .Z(n2173) );
  AND U2872 ( .A(n2174), .B(n2175), .Z(n2172) );
  NAND U2873 ( .A(n2155), .B(\u_a23_mem/p_mem[39][5] ), .Z(n2175) );
  NANDN U2874 ( .B(n1046), .A(n2081), .Z(n2174) );
  NAND U2875 ( .A(n2176), .B(n2177), .Z(\u_a23_mem/n19102 ) );
  OR U2876 ( .A(n1049), .B(n2152), .Z(n2177) );
  AND U2877 ( .A(n2178), .B(n2179), .Z(n2176) );
  NAND U2878 ( .A(n2155), .B(\u_a23_mem/p_mem[39][6] ), .Z(n2179) );
  NANDN U2879 ( .B(n1052), .A(n2081), .Z(n2178) );
  NAND U2880 ( .A(n2180), .B(n2181), .Z(\u_a23_mem/n19101 ) );
  NANDN U2881 ( .B(n2152), .A(n1055), .Z(n2181) );
  NAND U2882 ( .A(n1056), .B(n2081), .Z(n2152) );
  AND U2883 ( .A(n2182), .B(n2183), .Z(n2180) );
  NAND U2884 ( .A(n2155), .B(\u_a23_mem/p_mem[39][7] ), .Z(n2183) );
  NANDN U2885 ( .B(n1059), .A(n2081), .Z(n2155) );
  NAND U2886 ( .A(n1061), .B(n2081), .Z(n2182) );
  AND U2887 ( .A(n1694), .B(n2184), .Z(n2081) );
  NAND U2888 ( .A(n2185), .B(n2186), .Z(\u_a23_mem/n19100 ) );
  NAND U2889 ( .A(n2187), .B(\u_a23_mem/p_mem[40][0] ), .Z(n2186) );
  OR U2890 ( .A(n1011), .B(n2188), .Z(n2185) );
  NAND U2891 ( .A(n2189), .B(n2190), .Z(\u_a23_mem/n19099 ) );
  NAND U2892 ( .A(n2187), .B(\u_a23_mem/p_mem[40][1] ), .Z(n2190) );
  OR U2893 ( .A(n1019), .B(n2188), .Z(n2189) );
  NAND U2894 ( .A(n2191), .B(n2192), .Z(\u_a23_mem/n19098 ) );
  NAND U2895 ( .A(n2187), .B(\u_a23_mem/p_mem[40][2] ), .Z(n2192) );
  OR U2896 ( .A(n1025), .B(n2188), .Z(n2191) );
  NAND U2897 ( .A(n2193), .B(n2194), .Z(\u_a23_mem/n19097 ) );
  NAND U2898 ( .A(n2187), .B(\u_a23_mem/p_mem[40][3] ), .Z(n2194) );
  OR U2899 ( .A(n1031), .B(n2188), .Z(n2193) );
  NAND U2900 ( .A(n2195), .B(n2196), .Z(\u_a23_mem/n19096 ) );
  NAND U2901 ( .A(n2187), .B(\u_a23_mem/p_mem[40][4] ), .Z(n2196) );
  OR U2902 ( .A(n1037), .B(n2188), .Z(n2195) );
  NAND U2903 ( .A(n2197), .B(n2198), .Z(\u_a23_mem/n19095 ) );
  NAND U2904 ( .A(n2187), .B(\u_a23_mem/p_mem[40][5] ), .Z(n2198) );
  OR U2905 ( .A(n1043), .B(n2188), .Z(n2197) );
  NAND U2906 ( .A(n2199), .B(n2200), .Z(\u_a23_mem/n19094 ) );
  NAND U2907 ( .A(n2187), .B(\u_a23_mem/p_mem[40][6] ), .Z(n2200) );
  OR U2908 ( .A(n1049), .B(n2188), .Z(n2199) );
  NAND U2909 ( .A(n2201), .B(n2202), .Z(\u_a23_mem/n19093 ) );
  NAND U2910 ( .A(n2187), .B(\u_a23_mem/p_mem[40][7] ), .Z(n2202) );
  NANDN U2911 ( .B(n1080), .A(n2203), .Z(n2187) );
  NANDN U2912 ( .B(n2188), .A(n1055), .Z(n2201) );
  NANDN U2913 ( .B(n2), .A(n2203), .Z(n2188) );
  NAND U2914 ( .A(n2204), .B(n2205), .Z(\u_a23_mem/n19092 ) );
  OR U2915 ( .A(n1011), .B(n2206), .Z(n2205) );
  AND U2916 ( .A(n2207), .B(n2208), .Z(n2204) );
  NANDN U2917 ( .B(n1087), .A(n2203), .Z(n2208) );
  NAND U2918 ( .A(n2209), .B(\u_a23_mem/p_mem[41][0] ), .Z(n2207) );
  NAND U2919 ( .A(n2210), .B(n2211), .Z(\u_a23_mem/n19091 ) );
  OR U2920 ( .A(n1019), .B(n2206), .Z(n2211) );
  AND U2921 ( .A(n2212), .B(n2213), .Z(n2210) );
  NANDN U2922 ( .B(n1093), .A(n2203), .Z(n2213) );
  NAND U2923 ( .A(n2209), .B(\u_a23_mem/p_mem[41][1] ), .Z(n2212) );
  NAND U2924 ( .A(n2214), .B(n2215), .Z(\u_a23_mem/n19090 ) );
  OR U2925 ( .A(n1025), .B(n2206), .Z(n2215) );
  AND U2926 ( .A(n2216), .B(n2217), .Z(n2214) );
  NANDN U2927 ( .B(n1098), .A(n2203), .Z(n2217) );
  NAND U2928 ( .A(n2209), .B(\u_a23_mem/p_mem[41][2] ), .Z(n2216) );
  NAND U2929 ( .A(n2218), .B(n2219), .Z(\u_a23_mem/n19089 ) );
  OR U2930 ( .A(n1031), .B(n2206), .Z(n2219) );
  AND U2931 ( .A(n2220), .B(n2221), .Z(n2218) );
  NANDN U2932 ( .B(n1103), .A(n2203), .Z(n2221) );
  NAND U2933 ( .A(n2209), .B(\u_a23_mem/p_mem[41][3] ), .Z(n2220) );
  NAND U2934 ( .A(n2222), .B(n2223), .Z(\u_a23_mem/n19088 ) );
  OR U2935 ( .A(n1037), .B(n2206), .Z(n2223) );
  AND U2936 ( .A(n2224), .B(n2225), .Z(n2222) );
  NANDN U2937 ( .B(n1108), .A(n2203), .Z(n2225) );
  NAND U2938 ( .A(n2209), .B(\u_a23_mem/p_mem[41][4] ), .Z(n2224) );
  NAND U2939 ( .A(n2226), .B(n2227), .Z(\u_a23_mem/n19087 ) );
  OR U2940 ( .A(n1043), .B(n2206), .Z(n2227) );
  AND U2941 ( .A(n2228), .B(n2229), .Z(n2226) );
  NANDN U2942 ( .B(n1113), .A(n2203), .Z(n2229) );
  NAND U2943 ( .A(n2209), .B(\u_a23_mem/p_mem[41][5] ), .Z(n2228) );
  NAND U2944 ( .A(n2230), .B(n2231), .Z(\u_a23_mem/n19086 ) );
  OR U2945 ( .A(n1049), .B(n2206), .Z(n2231) );
  AND U2946 ( .A(n2232), .B(n2233), .Z(n2230) );
  NANDN U2947 ( .B(n1118), .A(n2203), .Z(n2233) );
  NAND U2948 ( .A(n2209), .B(\u_a23_mem/p_mem[41][6] ), .Z(n2232) );
  NAND U2949 ( .A(n2234), .B(n2235), .Z(\u_a23_mem/n19085 ) );
  NANDN U2950 ( .B(n2206), .A(n1055), .Z(n2235) );
  NAND U2951 ( .A(n1121), .B(n2203), .Z(n2206) );
  AND U2952 ( .A(n2236), .B(n2237), .Z(n2234) );
  NANDN U2953 ( .B(n1124), .A(n2203), .Z(n2237) );
  NAND U2954 ( .A(n2209), .B(\u_a23_mem/p_mem[41][7] ), .Z(n2236) );
  NANDN U2955 ( .B(n1125), .A(n2203), .Z(n2209) );
  NAND U2956 ( .A(n2238), .B(n2239), .Z(\u_a23_mem/n19084 ) );
  OR U2957 ( .A(n1011), .B(n2240), .Z(n2239) );
  AND U2958 ( .A(n2241), .B(n2242), .Z(n2238) );
  NANDN U2959 ( .B(n1131), .A(n2203), .Z(n2242) );
  NAND U2960 ( .A(n2243), .B(\u_a23_mem/p_mem[42][0] ), .Z(n2241) );
  NAND U2961 ( .A(n2244), .B(n2245), .Z(\u_a23_mem/n19083 ) );
  OR U2962 ( .A(n1019), .B(n2240), .Z(n2245) );
  AND U2963 ( .A(n2246), .B(n2247), .Z(n2244) );
  NANDN U2964 ( .B(n1137), .A(n2203), .Z(n2247) );
  NAND U2965 ( .A(n2243), .B(\u_a23_mem/p_mem[42][1] ), .Z(n2246) );
  NAND U2966 ( .A(n2248), .B(n2249), .Z(\u_a23_mem/n19082 ) );
  OR U2967 ( .A(n1025), .B(n2240), .Z(n2249) );
  AND U2968 ( .A(n2250), .B(n2251), .Z(n2248) );
  NANDN U2969 ( .B(n1142), .A(n2203), .Z(n2251) );
  NAND U2970 ( .A(n2243), .B(\u_a23_mem/p_mem[42][2] ), .Z(n2250) );
  NAND U2971 ( .A(n2252), .B(n2253), .Z(\u_a23_mem/n19081 ) );
  OR U2972 ( .A(n1031), .B(n2240), .Z(n2253) );
  AND U2973 ( .A(n2254), .B(n2255), .Z(n2252) );
  NANDN U2974 ( .B(n1147), .A(n2203), .Z(n2255) );
  NAND U2975 ( .A(n2243), .B(\u_a23_mem/p_mem[42][3] ), .Z(n2254) );
  NAND U2976 ( .A(n2256), .B(n2257), .Z(\u_a23_mem/n19080 ) );
  OR U2977 ( .A(n1037), .B(n2240), .Z(n2257) );
  AND U2978 ( .A(n2258), .B(n2259), .Z(n2256) );
  NANDN U2979 ( .B(n1152), .A(n2203), .Z(n2259) );
  NAND U2980 ( .A(n2243), .B(\u_a23_mem/p_mem[42][4] ), .Z(n2258) );
  NAND U2981 ( .A(n2260), .B(n2261), .Z(\u_a23_mem/n19079 ) );
  OR U2982 ( .A(n1043), .B(n2240), .Z(n2261) );
  AND U2983 ( .A(n2262), .B(n2263), .Z(n2260) );
  NANDN U2984 ( .B(n1157), .A(n2203), .Z(n2263) );
  NAND U2985 ( .A(n2243), .B(\u_a23_mem/p_mem[42][5] ), .Z(n2262) );
  NAND U2986 ( .A(n2264), .B(n2265), .Z(\u_a23_mem/n19078 ) );
  OR U2987 ( .A(n1049), .B(n2240), .Z(n2265) );
  AND U2988 ( .A(n2266), .B(n2267), .Z(n2264) );
  NANDN U2989 ( .B(n1162), .A(n2203), .Z(n2267) );
  NAND U2990 ( .A(n2243), .B(\u_a23_mem/p_mem[42][6] ), .Z(n2266) );
  NAND U2991 ( .A(n2268), .B(n2269), .Z(\u_a23_mem/n19077 ) );
  NANDN U2992 ( .B(n2240), .A(n1055), .Z(n2269) );
  NAND U2993 ( .A(n1165), .B(n2203), .Z(n2240) );
  AND U2994 ( .A(n2270), .B(n2271), .Z(n2268) );
  NANDN U2995 ( .B(n1168), .A(n2203), .Z(n2271) );
  NAND U2996 ( .A(n2243), .B(\u_a23_mem/p_mem[42][7] ), .Z(n2270) );
  NANDN U2997 ( .B(n1169), .A(n2203), .Z(n2243) );
  NAND U2998 ( .A(n2272), .B(n2273), .Z(\u_a23_mem/n19076 ) );
  OR U2999 ( .A(n1011), .B(n2274), .Z(n2273) );
  AND U3000 ( .A(n2275), .B(n2276), .Z(n2272) );
  NAND U3001 ( .A(n2277), .B(\u_a23_mem/p_mem[43][0] ), .Z(n2276) );
  NANDN U3002 ( .B(n1015), .A(n2203), .Z(n2275) );
  NAND U3003 ( .A(n2278), .B(n2279), .Z(\u_a23_mem/n19075 ) );
  OR U3004 ( .A(n1019), .B(n2274), .Z(n2279) );
  AND U3005 ( .A(n2280), .B(n2281), .Z(n2278) );
  NAND U3006 ( .A(n2277), .B(\u_a23_mem/p_mem[43][1] ), .Z(n2281) );
  NANDN U3007 ( .B(n1022), .A(n2203), .Z(n2280) );
  NAND U3008 ( .A(n2282), .B(n2283), .Z(\u_a23_mem/n19074 ) );
  OR U3009 ( .A(n1025), .B(n2274), .Z(n2283) );
  AND U3010 ( .A(n2284), .B(n2285), .Z(n2282) );
  NAND U3011 ( .A(n2277), .B(\u_a23_mem/p_mem[43][2] ), .Z(n2285) );
  NANDN U3012 ( .B(n1028), .A(n2203), .Z(n2284) );
  NAND U3013 ( .A(n2286), .B(n2287), .Z(\u_a23_mem/n19073 ) );
  OR U3014 ( .A(n1031), .B(n2274), .Z(n2287) );
  AND U3015 ( .A(n2288), .B(n2289), .Z(n2286) );
  NAND U3016 ( .A(n2277), .B(\u_a23_mem/p_mem[43][3] ), .Z(n2289) );
  NANDN U3017 ( .B(n1034), .A(n2203), .Z(n2288) );
  NAND U3018 ( .A(n2290), .B(n2291), .Z(\u_a23_mem/n19072 ) );
  OR U3019 ( .A(n1037), .B(n2274), .Z(n2291) );
  AND U3020 ( .A(n2292), .B(n2293), .Z(n2290) );
  NAND U3021 ( .A(n2277), .B(\u_a23_mem/p_mem[43][4] ), .Z(n2293) );
  NANDN U3022 ( .B(n1040), .A(n2203), .Z(n2292) );
  NAND U3023 ( .A(n2294), .B(n2295), .Z(\u_a23_mem/n19071 ) );
  OR U3024 ( .A(n1043), .B(n2274), .Z(n2295) );
  AND U3025 ( .A(n2296), .B(n2297), .Z(n2294) );
  NAND U3026 ( .A(n2277), .B(\u_a23_mem/p_mem[43][5] ), .Z(n2297) );
  NANDN U3027 ( .B(n1046), .A(n2203), .Z(n2296) );
  NAND U3028 ( .A(n2298), .B(n2299), .Z(\u_a23_mem/n19070 ) );
  OR U3029 ( .A(n1049), .B(n2274), .Z(n2299) );
  AND U3030 ( .A(n2300), .B(n2301), .Z(n2298) );
  NAND U3031 ( .A(n2277), .B(\u_a23_mem/p_mem[43][6] ), .Z(n2301) );
  NANDN U3032 ( .B(n1052), .A(n2203), .Z(n2300) );
  NAND U3033 ( .A(n2302), .B(n2303), .Z(\u_a23_mem/n19069 ) );
  NANDN U3034 ( .B(n2274), .A(n1055), .Z(n2303) );
  NAND U3035 ( .A(n1056), .B(n2203), .Z(n2274) );
  AND U3036 ( .A(n2304), .B(n2305), .Z(n2302) );
  NAND U3037 ( .A(n2277), .B(\u_a23_mem/p_mem[43][7] ), .Z(n2305) );
  NANDN U3038 ( .B(n1059), .A(n2203), .Z(n2277) );
  NAND U3039 ( .A(n1061), .B(n2203), .Z(n2304) );
  AND U3040 ( .A(n1816), .B(n2184), .Z(n2203) );
  NAND U3041 ( .A(n2306), .B(n2307), .Z(\u_a23_mem/n19068 ) );
  NAND U3042 ( .A(n2308), .B(\u_a23_mem/p_mem[44][0] ), .Z(n2307) );
  OR U3043 ( .A(n1011), .B(n2309), .Z(n2306) );
  NAND U3044 ( .A(n2310), .B(n2311), .Z(\u_a23_mem/n19067 ) );
  NAND U3045 ( .A(n2308), .B(\u_a23_mem/p_mem[44][1] ), .Z(n2311) );
  OR U3046 ( .A(n1019), .B(n2309), .Z(n2310) );
  NAND U3047 ( .A(n2312), .B(n2313), .Z(\u_a23_mem/n19066 ) );
  NAND U3048 ( .A(n2308), .B(\u_a23_mem/p_mem[44][2] ), .Z(n2313) );
  OR U3049 ( .A(n1025), .B(n2309), .Z(n2312) );
  NAND U3050 ( .A(n2314), .B(n2315), .Z(\u_a23_mem/n19065 ) );
  NAND U3051 ( .A(n2308), .B(\u_a23_mem/p_mem[44][3] ), .Z(n2315) );
  OR U3052 ( .A(n1031), .B(n2309), .Z(n2314) );
  NAND U3053 ( .A(n2316), .B(n2317), .Z(\u_a23_mem/n19064 ) );
  NAND U3054 ( .A(n2308), .B(\u_a23_mem/p_mem[44][4] ), .Z(n2317) );
  OR U3055 ( .A(n1037), .B(n2309), .Z(n2316) );
  NAND U3056 ( .A(n2318), .B(n2319), .Z(\u_a23_mem/n19063 ) );
  NAND U3057 ( .A(n2308), .B(\u_a23_mem/p_mem[44][5] ), .Z(n2319) );
  OR U3058 ( .A(n1043), .B(n2309), .Z(n2318) );
  NAND U3059 ( .A(n2320), .B(n2321), .Z(\u_a23_mem/n19062 ) );
  NAND U3060 ( .A(n2308), .B(\u_a23_mem/p_mem[44][6] ), .Z(n2321) );
  OR U3061 ( .A(n1049), .B(n2309), .Z(n2320) );
  NAND U3062 ( .A(n2322), .B(n2323), .Z(\u_a23_mem/n19061 ) );
  NAND U3063 ( .A(n2308), .B(\u_a23_mem/p_mem[44][7] ), .Z(n2323) );
  NANDN U3064 ( .B(n1080), .A(n2324), .Z(n2308) );
  NANDN U3065 ( .B(n2309), .A(n1055), .Z(n2322) );
  NANDN U3066 ( .B(n2), .A(n2324), .Z(n2309) );
  NAND U3067 ( .A(n2325), .B(n2326), .Z(\u_a23_mem/n19060 ) );
  OR U3068 ( .A(n1011), .B(n2327), .Z(n2326) );
  AND U3069 ( .A(n2328), .B(n2329), .Z(n2325) );
  NANDN U3070 ( .B(n1087), .A(n2324), .Z(n2329) );
  NAND U3071 ( .A(n2330), .B(\u_a23_mem/p_mem[45][0] ), .Z(n2328) );
  NAND U3072 ( .A(n2331), .B(n2332), .Z(\u_a23_mem/n19059 ) );
  OR U3073 ( .A(n1019), .B(n2327), .Z(n2332) );
  AND U3074 ( .A(n2333), .B(n2334), .Z(n2331) );
  NANDN U3075 ( .B(n1093), .A(n2324), .Z(n2334) );
  NAND U3076 ( .A(n2330), .B(\u_a23_mem/p_mem[45][1] ), .Z(n2333) );
  NAND U3077 ( .A(n2335), .B(n2336), .Z(\u_a23_mem/n19058 ) );
  OR U3078 ( .A(n1025), .B(n2327), .Z(n2336) );
  AND U3079 ( .A(n2337), .B(n2338), .Z(n2335) );
  NANDN U3080 ( .B(n1098), .A(n2324), .Z(n2338) );
  NAND U3081 ( .A(n2330), .B(\u_a23_mem/p_mem[45][2] ), .Z(n2337) );
  NAND U3082 ( .A(n2339), .B(n2340), .Z(\u_a23_mem/n19057 ) );
  OR U3083 ( .A(n1031), .B(n2327), .Z(n2340) );
  AND U3084 ( .A(n2341), .B(n2342), .Z(n2339) );
  NANDN U3085 ( .B(n1103), .A(n2324), .Z(n2342) );
  NAND U3086 ( .A(n2330), .B(\u_a23_mem/p_mem[45][3] ), .Z(n2341) );
  NAND U3087 ( .A(n2343), .B(n2344), .Z(\u_a23_mem/n19056 ) );
  OR U3088 ( .A(n1037), .B(n2327), .Z(n2344) );
  AND U3089 ( .A(n2345), .B(n2346), .Z(n2343) );
  NANDN U3090 ( .B(n1108), .A(n2324), .Z(n2346) );
  NAND U3091 ( .A(n2330), .B(\u_a23_mem/p_mem[45][4] ), .Z(n2345) );
  NAND U3092 ( .A(n2347), .B(n2348), .Z(\u_a23_mem/n19055 ) );
  OR U3093 ( .A(n1043), .B(n2327), .Z(n2348) );
  AND U3094 ( .A(n2349), .B(n2350), .Z(n2347) );
  NANDN U3095 ( .B(n1113), .A(n2324), .Z(n2350) );
  NAND U3096 ( .A(n2330), .B(\u_a23_mem/p_mem[45][5] ), .Z(n2349) );
  NAND U3097 ( .A(n2351), .B(n2352), .Z(\u_a23_mem/n19054 ) );
  OR U3098 ( .A(n1049), .B(n2327), .Z(n2352) );
  AND U3099 ( .A(n2353), .B(n2354), .Z(n2351) );
  NANDN U3100 ( .B(n1118), .A(n2324), .Z(n2354) );
  NAND U3101 ( .A(n2330), .B(\u_a23_mem/p_mem[45][6] ), .Z(n2353) );
  NAND U3102 ( .A(n2355), .B(n2356), .Z(\u_a23_mem/n19053 ) );
  NANDN U3103 ( .B(n2327), .A(n1055), .Z(n2356) );
  NAND U3104 ( .A(n1121), .B(n2324), .Z(n2327) );
  AND U3105 ( .A(n2357), .B(n2358), .Z(n2355) );
  NANDN U3106 ( .B(n1124), .A(n2324), .Z(n2358) );
  NAND U3107 ( .A(n2330), .B(\u_a23_mem/p_mem[45][7] ), .Z(n2357) );
  NANDN U3108 ( .B(n1125), .A(n2324), .Z(n2330) );
  NAND U3109 ( .A(n2359), .B(n2360), .Z(\u_a23_mem/n19052 ) );
  OR U3110 ( .A(n1011), .B(n2361), .Z(n2360) );
  AND U3111 ( .A(n2362), .B(n2363), .Z(n2359) );
  NANDN U3112 ( .B(n1131), .A(n2324), .Z(n2363) );
  NAND U3113 ( .A(n2364), .B(\u_a23_mem/p_mem[46][0] ), .Z(n2362) );
  NAND U3114 ( .A(n2365), .B(n2366), .Z(\u_a23_mem/n19051 ) );
  OR U3115 ( .A(n1019), .B(n2361), .Z(n2366) );
  AND U3116 ( .A(n2367), .B(n2368), .Z(n2365) );
  NANDN U3117 ( .B(n1137), .A(n2324), .Z(n2368) );
  NAND U3118 ( .A(n2364), .B(\u_a23_mem/p_mem[46][1] ), .Z(n2367) );
  NAND U3119 ( .A(n2369), .B(n2370), .Z(\u_a23_mem/n19050 ) );
  OR U3120 ( .A(n1025), .B(n2361), .Z(n2370) );
  AND U3121 ( .A(n2371), .B(n2372), .Z(n2369) );
  NANDN U3122 ( .B(n1142), .A(n2324), .Z(n2372) );
  NAND U3123 ( .A(n2364), .B(\u_a23_mem/p_mem[46][2] ), .Z(n2371) );
  NAND U3124 ( .A(n2373), .B(n2374), .Z(\u_a23_mem/n19049 ) );
  OR U3125 ( .A(n1031), .B(n2361), .Z(n2374) );
  AND U3126 ( .A(n2375), .B(n2376), .Z(n2373) );
  NANDN U3127 ( .B(n1147), .A(n2324), .Z(n2376) );
  NAND U3128 ( .A(n2364), .B(\u_a23_mem/p_mem[46][3] ), .Z(n2375) );
  NAND U3129 ( .A(n2377), .B(n2378), .Z(\u_a23_mem/n19048 ) );
  OR U3130 ( .A(n1037), .B(n2361), .Z(n2378) );
  AND U3131 ( .A(n2379), .B(n2380), .Z(n2377) );
  NANDN U3132 ( .B(n1152), .A(n2324), .Z(n2380) );
  NAND U3133 ( .A(n2364), .B(\u_a23_mem/p_mem[46][4] ), .Z(n2379) );
  NAND U3134 ( .A(n2381), .B(n2382), .Z(\u_a23_mem/n19047 ) );
  OR U3135 ( .A(n1043), .B(n2361), .Z(n2382) );
  AND U3136 ( .A(n2383), .B(n2384), .Z(n2381) );
  NANDN U3137 ( .B(n1157), .A(n2324), .Z(n2384) );
  NAND U3138 ( .A(n2364), .B(\u_a23_mem/p_mem[46][5] ), .Z(n2383) );
  NAND U3139 ( .A(n2385), .B(n2386), .Z(\u_a23_mem/n19046 ) );
  OR U3140 ( .A(n1049), .B(n2361), .Z(n2386) );
  AND U3141 ( .A(n2387), .B(n2388), .Z(n2385) );
  NANDN U3142 ( .B(n1162), .A(n2324), .Z(n2388) );
  NAND U3143 ( .A(n2364), .B(\u_a23_mem/p_mem[46][6] ), .Z(n2387) );
  NAND U3144 ( .A(n2389), .B(n2390), .Z(\u_a23_mem/n19045 ) );
  NANDN U3145 ( .B(n2361), .A(n1055), .Z(n2390) );
  NAND U3146 ( .A(n1165), .B(n2324), .Z(n2361) );
  AND U3147 ( .A(n2391), .B(n2392), .Z(n2389) );
  NANDN U3148 ( .B(n1168), .A(n2324), .Z(n2392) );
  NAND U3149 ( .A(n2364), .B(\u_a23_mem/p_mem[46][7] ), .Z(n2391) );
  NANDN U3150 ( .B(n1169), .A(n2324), .Z(n2364) );
  NAND U3151 ( .A(n2393), .B(n2394), .Z(\u_a23_mem/n19044 ) );
  OR U3152 ( .A(n1011), .B(n2395), .Z(n2394) );
  AND U3153 ( .A(n2396), .B(n2397), .Z(n2393) );
  NAND U3154 ( .A(n2398), .B(\u_a23_mem/p_mem[47][0] ), .Z(n2397) );
  NANDN U3155 ( .B(n1015), .A(n2324), .Z(n2396) );
  NAND U3156 ( .A(n2399), .B(n2400), .Z(\u_a23_mem/n19043 ) );
  OR U3157 ( .A(n1019), .B(n2395), .Z(n2400) );
  AND U3158 ( .A(n2401), .B(n2402), .Z(n2399) );
  NAND U3159 ( .A(n2398), .B(\u_a23_mem/p_mem[47][1] ), .Z(n2402) );
  NANDN U3160 ( .B(n1022), .A(n2324), .Z(n2401) );
  NAND U3161 ( .A(n2403), .B(n2404), .Z(\u_a23_mem/n19042 ) );
  OR U3162 ( .A(n1025), .B(n2395), .Z(n2404) );
  AND U3163 ( .A(n2405), .B(n2406), .Z(n2403) );
  NAND U3164 ( .A(n2398), .B(\u_a23_mem/p_mem[47][2] ), .Z(n2406) );
  NANDN U3165 ( .B(n1028), .A(n2324), .Z(n2405) );
  NAND U3166 ( .A(n2407), .B(n2408), .Z(\u_a23_mem/n19041 ) );
  OR U3167 ( .A(n1031), .B(n2395), .Z(n2408) );
  AND U3168 ( .A(n2409), .B(n2410), .Z(n2407) );
  NAND U3169 ( .A(n2398), .B(\u_a23_mem/p_mem[47][3] ), .Z(n2410) );
  NANDN U3170 ( .B(n1034), .A(n2324), .Z(n2409) );
  NAND U3171 ( .A(n2411), .B(n2412), .Z(\u_a23_mem/n19040 ) );
  OR U3172 ( .A(n1037), .B(n2395), .Z(n2412) );
  AND U3173 ( .A(n2413), .B(n2414), .Z(n2411) );
  NAND U3174 ( .A(n2398), .B(\u_a23_mem/p_mem[47][4] ), .Z(n2414) );
  NANDN U3175 ( .B(n1040), .A(n2324), .Z(n2413) );
  NAND U3176 ( .A(n2415), .B(n2416), .Z(\u_a23_mem/n19039 ) );
  OR U3177 ( .A(n1043), .B(n2395), .Z(n2416) );
  AND U3178 ( .A(n2417), .B(n2418), .Z(n2415) );
  NAND U3179 ( .A(n2398), .B(\u_a23_mem/p_mem[47][5] ), .Z(n2418) );
  NANDN U3180 ( .B(n1046), .A(n2324), .Z(n2417) );
  NAND U3181 ( .A(n2419), .B(n2420), .Z(\u_a23_mem/n19038 ) );
  OR U3182 ( .A(n1049), .B(n2395), .Z(n2420) );
  AND U3183 ( .A(n2421), .B(n2422), .Z(n2419) );
  NAND U3184 ( .A(n2398), .B(\u_a23_mem/p_mem[47][6] ), .Z(n2422) );
  NANDN U3185 ( .B(n1052), .A(n2324), .Z(n2421) );
  NAND U3186 ( .A(n2423), .B(n2424), .Z(\u_a23_mem/n19037 ) );
  NANDN U3187 ( .B(n2395), .A(n1055), .Z(n2424) );
  NAND U3188 ( .A(n1056), .B(n2324), .Z(n2395) );
  AND U3189 ( .A(n2425), .B(n2426), .Z(n2423) );
  NAND U3190 ( .A(n2398), .B(\u_a23_mem/p_mem[47][7] ), .Z(n2426) );
  NANDN U3191 ( .B(n1059), .A(n2324), .Z(n2398) );
  NAND U3192 ( .A(n1061), .B(n2324), .Z(n2425) );
  NOR U3193 ( .A(n2062), .B(n1938), .Z(n2324) );
  IV U3194 ( .A(n2184), .Z(n2062) );
  ANDN U3195 ( .A(n2427), .B(n2428), .Z(n2184) );
  AND U3196 ( .A(n1939), .B(n2429), .Z(n2427) );
  NAND U3197 ( .A(n2430), .B(n2431), .Z(\u_a23_mem/n19036 ) );
  NAND U3198 ( .A(n2432), .B(\u_a23_mem/p_mem[48][0] ), .Z(n2431) );
  OR U3199 ( .A(n1011), .B(n2433), .Z(n2430) );
  NAND U3200 ( .A(n2434), .B(n2435), .Z(\u_a23_mem/n19035 ) );
  NAND U3201 ( .A(n2432), .B(\u_a23_mem/p_mem[48][1] ), .Z(n2435) );
  OR U3202 ( .A(n1019), .B(n2433), .Z(n2434) );
  NAND U3203 ( .A(n2436), .B(n2437), .Z(\u_a23_mem/n19034 ) );
  NAND U3204 ( .A(n2432), .B(\u_a23_mem/p_mem[48][2] ), .Z(n2437) );
  OR U3205 ( .A(n1025), .B(n2433), .Z(n2436) );
  NAND U3206 ( .A(n2438), .B(n2439), .Z(\u_a23_mem/n19033 ) );
  NAND U3207 ( .A(n2432), .B(\u_a23_mem/p_mem[48][3] ), .Z(n2439) );
  OR U3208 ( .A(n1031), .B(n2433), .Z(n2438) );
  NAND U3209 ( .A(n2440), .B(n2441), .Z(\u_a23_mem/n19032 ) );
  NAND U3210 ( .A(n2432), .B(\u_a23_mem/p_mem[48][4] ), .Z(n2441) );
  OR U3211 ( .A(n1037), .B(n2433), .Z(n2440) );
  NAND U3212 ( .A(n2442), .B(n2443), .Z(\u_a23_mem/n19031 ) );
  NAND U3213 ( .A(n2432), .B(\u_a23_mem/p_mem[48][5] ), .Z(n2443) );
  OR U3214 ( .A(n1043), .B(n2433), .Z(n2442) );
  NAND U3215 ( .A(n2444), .B(n2445), .Z(\u_a23_mem/n19030 ) );
  NAND U3216 ( .A(n2432), .B(\u_a23_mem/p_mem[48][6] ), .Z(n2445) );
  OR U3217 ( .A(n1049), .B(n2433), .Z(n2444) );
  NAND U3218 ( .A(n2446), .B(n2447), .Z(\u_a23_mem/n19029 ) );
  NAND U3219 ( .A(n2432), .B(\u_a23_mem/p_mem[48][7] ), .Z(n2447) );
  NANDN U3220 ( .B(n1080), .A(n2448), .Z(n2432) );
  NANDN U3221 ( .B(n2433), .A(n1055), .Z(n2446) );
  NANDN U3222 ( .B(n2), .A(n2448), .Z(n2433) );
  NAND U3223 ( .A(n2449), .B(n2450), .Z(\u_a23_mem/n19028 ) );
  OR U3224 ( .A(n1011), .B(n2451), .Z(n2450) );
  AND U3225 ( .A(n2452), .B(n2453), .Z(n2449) );
  NANDN U3226 ( .B(n1087), .A(n2448), .Z(n2453) );
  NAND U3227 ( .A(n2454), .B(\u_a23_mem/p_mem[49][0] ), .Z(n2452) );
  NAND U3228 ( .A(n2455), .B(n2456), .Z(\u_a23_mem/n19027 ) );
  OR U3229 ( .A(n1019), .B(n2451), .Z(n2456) );
  AND U3230 ( .A(n2457), .B(n2458), .Z(n2455) );
  NANDN U3231 ( .B(n1093), .A(n2448), .Z(n2458) );
  NAND U3232 ( .A(n2454), .B(\u_a23_mem/p_mem[49][1] ), .Z(n2457) );
  NAND U3233 ( .A(n2459), .B(n2460), .Z(\u_a23_mem/n19026 ) );
  OR U3234 ( .A(n1025), .B(n2451), .Z(n2460) );
  AND U3235 ( .A(n2461), .B(n2462), .Z(n2459) );
  NANDN U3236 ( .B(n1098), .A(n2448), .Z(n2462) );
  NAND U3237 ( .A(n2454), .B(\u_a23_mem/p_mem[49][2] ), .Z(n2461) );
  NAND U3238 ( .A(n2463), .B(n2464), .Z(\u_a23_mem/n19025 ) );
  OR U3239 ( .A(n1031), .B(n2451), .Z(n2464) );
  AND U3240 ( .A(n2465), .B(n2466), .Z(n2463) );
  NANDN U3241 ( .B(n1103), .A(n2448), .Z(n2466) );
  NAND U3242 ( .A(n2454), .B(\u_a23_mem/p_mem[49][3] ), .Z(n2465) );
  NAND U3243 ( .A(n2467), .B(n2468), .Z(\u_a23_mem/n19024 ) );
  OR U3244 ( .A(n1037), .B(n2451), .Z(n2468) );
  AND U3245 ( .A(n2469), .B(n2470), .Z(n2467) );
  NANDN U3246 ( .B(n1108), .A(n2448), .Z(n2470) );
  NAND U3247 ( .A(n2454), .B(\u_a23_mem/p_mem[49][4] ), .Z(n2469) );
  NAND U3248 ( .A(n2471), .B(n2472), .Z(\u_a23_mem/n19023 ) );
  OR U3249 ( .A(n1043), .B(n2451), .Z(n2472) );
  AND U3250 ( .A(n2473), .B(n2474), .Z(n2471) );
  NANDN U3251 ( .B(n1113), .A(n2448), .Z(n2474) );
  NAND U3252 ( .A(n2454), .B(\u_a23_mem/p_mem[49][5] ), .Z(n2473) );
  NAND U3253 ( .A(n2475), .B(n2476), .Z(\u_a23_mem/n19022 ) );
  OR U3254 ( .A(n1049), .B(n2451), .Z(n2476) );
  AND U3255 ( .A(n2477), .B(n2478), .Z(n2475) );
  NANDN U3256 ( .B(n1118), .A(n2448), .Z(n2478) );
  NAND U3257 ( .A(n2454), .B(\u_a23_mem/p_mem[49][6] ), .Z(n2477) );
  NAND U3258 ( .A(n2479), .B(n2480), .Z(\u_a23_mem/n19021 ) );
  NANDN U3259 ( .B(n2451), .A(n1055), .Z(n2480) );
  NAND U3260 ( .A(n1121), .B(n2448), .Z(n2451) );
  AND U3261 ( .A(n2481), .B(n2482), .Z(n2479) );
  NANDN U3262 ( .B(n1124), .A(n2448), .Z(n2482) );
  NAND U3263 ( .A(n2454), .B(\u_a23_mem/p_mem[49][7] ), .Z(n2481) );
  NANDN U3264 ( .B(n1125), .A(n2448), .Z(n2454) );
  NAND U3265 ( .A(n2483), .B(n2484), .Z(\u_a23_mem/n19020 ) );
  OR U3266 ( .A(n1011), .B(n2485), .Z(n2484) );
  AND U3267 ( .A(n2486), .B(n2487), .Z(n2483) );
  NANDN U3268 ( .B(n1131), .A(n2448), .Z(n2487) );
  NAND U3269 ( .A(n2488), .B(\u_a23_mem/p_mem[50][0] ), .Z(n2486) );
  NAND U3270 ( .A(n2489), .B(n2490), .Z(\u_a23_mem/n19019 ) );
  OR U3271 ( .A(n1019), .B(n2485), .Z(n2490) );
  AND U3272 ( .A(n2491), .B(n2492), .Z(n2489) );
  NANDN U3273 ( .B(n1137), .A(n2448), .Z(n2492) );
  NAND U3274 ( .A(n2488), .B(\u_a23_mem/p_mem[50][1] ), .Z(n2491) );
  NAND U3275 ( .A(n2493), .B(n2494), .Z(\u_a23_mem/n19018 ) );
  OR U3276 ( .A(n1025), .B(n2485), .Z(n2494) );
  AND U3277 ( .A(n2495), .B(n2496), .Z(n2493) );
  NANDN U3278 ( .B(n1142), .A(n2448), .Z(n2496) );
  NAND U3279 ( .A(n2488), .B(\u_a23_mem/p_mem[50][2] ), .Z(n2495) );
  NAND U3280 ( .A(n2497), .B(n2498), .Z(\u_a23_mem/n19017 ) );
  OR U3281 ( .A(n1031), .B(n2485), .Z(n2498) );
  AND U3282 ( .A(n2499), .B(n2500), .Z(n2497) );
  NANDN U3283 ( .B(n1147), .A(n2448), .Z(n2500) );
  NAND U3284 ( .A(n2488), .B(\u_a23_mem/p_mem[50][3] ), .Z(n2499) );
  NAND U3285 ( .A(n2501), .B(n2502), .Z(\u_a23_mem/n19016 ) );
  OR U3286 ( .A(n1037), .B(n2485), .Z(n2502) );
  AND U3287 ( .A(n2503), .B(n2504), .Z(n2501) );
  NANDN U3288 ( .B(n1152), .A(n2448), .Z(n2504) );
  NAND U3289 ( .A(n2488), .B(\u_a23_mem/p_mem[50][4] ), .Z(n2503) );
  NAND U3290 ( .A(n2505), .B(n2506), .Z(\u_a23_mem/n19015 ) );
  OR U3291 ( .A(n1043), .B(n2485), .Z(n2506) );
  AND U3292 ( .A(n2507), .B(n2508), .Z(n2505) );
  NANDN U3293 ( .B(n1157), .A(n2448), .Z(n2508) );
  NAND U3294 ( .A(n2488), .B(\u_a23_mem/p_mem[50][5] ), .Z(n2507) );
  NAND U3295 ( .A(n2509), .B(n2510), .Z(\u_a23_mem/n19014 ) );
  OR U3296 ( .A(n1049), .B(n2485), .Z(n2510) );
  AND U3297 ( .A(n2511), .B(n2512), .Z(n2509) );
  NANDN U3298 ( .B(n1162), .A(n2448), .Z(n2512) );
  NAND U3299 ( .A(n2488), .B(\u_a23_mem/p_mem[50][6] ), .Z(n2511) );
  NAND U3300 ( .A(n2513), .B(n2514), .Z(\u_a23_mem/n19013 ) );
  NANDN U3301 ( .B(n2485), .A(n1055), .Z(n2514) );
  NAND U3302 ( .A(n1165), .B(n2448), .Z(n2485) );
  AND U3303 ( .A(n2515), .B(n2516), .Z(n2513) );
  NANDN U3304 ( .B(n1168), .A(n2448), .Z(n2516) );
  NAND U3305 ( .A(n2488), .B(\u_a23_mem/p_mem[50][7] ), .Z(n2515) );
  NANDN U3306 ( .B(n1169), .A(n2448), .Z(n2488) );
  NAND U3307 ( .A(n2517), .B(n2518), .Z(\u_a23_mem/n19012 ) );
  OR U3308 ( .A(n1011), .B(n2519), .Z(n2518) );
  AND U3309 ( .A(n2520), .B(n2521), .Z(n2517) );
  NAND U3310 ( .A(n2522), .B(\u_a23_mem/p_mem[51][0] ), .Z(n2521) );
  NANDN U3311 ( .B(n1015), .A(n2448), .Z(n2520) );
  NAND U3312 ( .A(n2523), .B(n2524), .Z(\u_a23_mem/n19011 ) );
  OR U3313 ( .A(n1019), .B(n2519), .Z(n2524) );
  AND U3314 ( .A(n2525), .B(n2526), .Z(n2523) );
  NAND U3315 ( .A(n2522), .B(\u_a23_mem/p_mem[51][1] ), .Z(n2526) );
  NANDN U3316 ( .B(n1022), .A(n2448), .Z(n2525) );
  NAND U3317 ( .A(n2527), .B(n2528), .Z(\u_a23_mem/n19010 ) );
  OR U3318 ( .A(n1025), .B(n2519), .Z(n2528) );
  AND U3319 ( .A(n2529), .B(n2530), .Z(n2527) );
  NAND U3320 ( .A(n2522), .B(\u_a23_mem/p_mem[51][2] ), .Z(n2530) );
  NANDN U3321 ( .B(n1028), .A(n2448), .Z(n2529) );
  NAND U3322 ( .A(n2531), .B(n2532), .Z(\u_a23_mem/n19009 ) );
  OR U3323 ( .A(n1031), .B(n2519), .Z(n2532) );
  AND U3324 ( .A(n2533), .B(n2534), .Z(n2531) );
  NAND U3325 ( .A(n2522), .B(\u_a23_mem/p_mem[51][3] ), .Z(n2534) );
  NANDN U3326 ( .B(n1034), .A(n2448), .Z(n2533) );
  NAND U3327 ( .A(n2535), .B(n2536), .Z(\u_a23_mem/n19008 ) );
  OR U3328 ( .A(n1037), .B(n2519), .Z(n2536) );
  AND U3329 ( .A(n2537), .B(n2538), .Z(n2535) );
  NAND U3330 ( .A(n2522), .B(\u_a23_mem/p_mem[51][4] ), .Z(n2538) );
  NANDN U3331 ( .B(n1040), .A(n2448), .Z(n2537) );
  NAND U3332 ( .A(n2539), .B(n2540), .Z(\u_a23_mem/n19007 ) );
  OR U3333 ( .A(n1043), .B(n2519), .Z(n2540) );
  AND U3334 ( .A(n2541), .B(n2542), .Z(n2539) );
  NAND U3335 ( .A(n2522), .B(\u_a23_mem/p_mem[51][5] ), .Z(n2542) );
  NANDN U3336 ( .B(n1046), .A(n2448), .Z(n2541) );
  NAND U3337 ( .A(n2543), .B(n2544), .Z(\u_a23_mem/n19006 ) );
  OR U3338 ( .A(n1049), .B(n2519), .Z(n2544) );
  AND U3339 ( .A(n2545), .B(n2546), .Z(n2543) );
  NAND U3340 ( .A(n2522), .B(\u_a23_mem/p_mem[51][6] ), .Z(n2546) );
  NANDN U3341 ( .B(n1052), .A(n2448), .Z(n2545) );
  NAND U3342 ( .A(n2547), .B(n2548), .Z(\u_a23_mem/n19005 ) );
  NANDN U3343 ( .B(n2519), .A(n1055), .Z(n2548) );
  NAND U3344 ( .A(n1056), .B(n2448), .Z(n2519) );
  AND U3345 ( .A(n2549), .B(n2550), .Z(n2547) );
  NAND U3346 ( .A(n2522), .B(\u_a23_mem/p_mem[51][7] ), .Z(n2550) );
  NANDN U3347 ( .B(n1059), .A(n2448), .Z(n2522) );
  NAND U3348 ( .A(n1061), .B(n2448), .Z(n2549) );
  ANDN U3349 ( .A(n1571), .B(n2551), .Z(n2448) );
  NAND U3350 ( .A(n2552), .B(n2553), .Z(\u_a23_mem/n19004 ) );
  NAND U3351 ( .A(n2554), .B(\u_a23_mem/p_mem[52][0] ), .Z(n2553) );
  OR U3352 ( .A(n1011), .B(n2555), .Z(n2552) );
  NAND U3353 ( .A(n2556), .B(n2557), .Z(\u_a23_mem/n19003 ) );
  NAND U3354 ( .A(n2554), .B(\u_a23_mem/p_mem[52][1] ), .Z(n2557) );
  OR U3355 ( .A(n1019), .B(n2555), .Z(n2556) );
  NAND U3356 ( .A(n2558), .B(n2559), .Z(\u_a23_mem/n19002 ) );
  NAND U3357 ( .A(n2554), .B(\u_a23_mem/p_mem[52][2] ), .Z(n2559) );
  OR U3358 ( .A(n1025), .B(n2555), .Z(n2558) );
  NAND U3359 ( .A(n2560), .B(n2561), .Z(\u_a23_mem/n19001 ) );
  NAND U3360 ( .A(n2554), .B(\u_a23_mem/p_mem[52][3] ), .Z(n2561) );
  OR U3361 ( .A(n1031), .B(n2555), .Z(n2560) );
  NAND U3362 ( .A(n2562), .B(n2563), .Z(\u_a23_mem/n19000 ) );
  NAND U3363 ( .A(n2554), .B(\u_a23_mem/p_mem[52][4] ), .Z(n2563) );
  OR U3364 ( .A(n1037), .B(n2555), .Z(n2562) );
  NAND U3365 ( .A(n2564), .B(n2565), .Z(\u_a23_mem/n18999 ) );
  NAND U3366 ( .A(n2554), .B(\u_a23_mem/p_mem[52][5] ), .Z(n2565) );
  OR U3367 ( .A(n1043), .B(n2555), .Z(n2564) );
  NAND U3368 ( .A(n2566), .B(n2567), .Z(\u_a23_mem/n18998 ) );
  NAND U3369 ( .A(n2554), .B(\u_a23_mem/p_mem[52][6] ), .Z(n2567) );
  OR U3370 ( .A(n1049), .B(n2555), .Z(n2566) );
  NAND U3371 ( .A(n2568), .B(n2569), .Z(\u_a23_mem/n18997 ) );
  NAND U3372 ( .A(n2554), .B(\u_a23_mem/p_mem[52][7] ), .Z(n2569) );
  NANDN U3373 ( .B(n1080), .A(n2570), .Z(n2554) );
  NANDN U3374 ( .B(n2555), .A(n1055), .Z(n2568) );
  NANDN U3375 ( .B(n2), .A(n2570), .Z(n2555) );
  NAND U3376 ( .A(n2571), .B(n2572), .Z(\u_a23_mem/n18996 ) );
  OR U3377 ( .A(n1011), .B(n2573), .Z(n2572) );
  AND U3378 ( .A(n2574), .B(n2575), .Z(n2571) );
  NANDN U3379 ( .B(n1087), .A(n2570), .Z(n2575) );
  NAND U3380 ( .A(n2576), .B(\u_a23_mem/p_mem[53][0] ), .Z(n2574) );
  NAND U3381 ( .A(n2577), .B(n2578), .Z(\u_a23_mem/n18995 ) );
  OR U3382 ( .A(n1019), .B(n2573), .Z(n2578) );
  AND U3383 ( .A(n2579), .B(n2580), .Z(n2577) );
  NANDN U3384 ( .B(n1093), .A(n2570), .Z(n2580) );
  NAND U3385 ( .A(n2576), .B(\u_a23_mem/p_mem[53][1] ), .Z(n2579) );
  NAND U3386 ( .A(n2581), .B(n2582), .Z(\u_a23_mem/n18994 ) );
  OR U3387 ( .A(n1025), .B(n2573), .Z(n2582) );
  AND U3388 ( .A(n2583), .B(n2584), .Z(n2581) );
  NANDN U3389 ( .B(n1098), .A(n2570), .Z(n2584) );
  NAND U3390 ( .A(n2576), .B(\u_a23_mem/p_mem[53][2] ), .Z(n2583) );
  NAND U3391 ( .A(n2585), .B(n2586), .Z(\u_a23_mem/n18993 ) );
  OR U3392 ( .A(n1031), .B(n2573), .Z(n2586) );
  AND U3393 ( .A(n2587), .B(n2588), .Z(n2585) );
  NANDN U3394 ( .B(n1103), .A(n2570), .Z(n2588) );
  NAND U3395 ( .A(n2576), .B(\u_a23_mem/p_mem[53][3] ), .Z(n2587) );
  NAND U3396 ( .A(n2589), .B(n2590), .Z(\u_a23_mem/n18992 ) );
  OR U3397 ( .A(n1037), .B(n2573), .Z(n2590) );
  AND U3398 ( .A(n2591), .B(n2592), .Z(n2589) );
  NANDN U3399 ( .B(n1108), .A(n2570), .Z(n2592) );
  NAND U3400 ( .A(n2576), .B(\u_a23_mem/p_mem[53][4] ), .Z(n2591) );
  NAND U3401 ( .A(n2593), .B(n2594), .Z(\u_a23_mem/n18991 ) );
  OR U3402 ( .A(n1043), .B(n2573), .Z(n2594) );
  AND U3403 ( .A(n2595), .B(n2596), .Z(n2593) );
  NANDN U3404 ( .B(n1113), .A(n2570), .Z(n2596) );
  NAND U3405 ( .A(n2576), .B(\u_a23_mem/p_mem[53][5] ), .Z(n2595) );
  NAND U3406 ( .A(n2597), .B(n2598), .Z(\u_a23_mem/n18990 ) );
  OR U3407 ( .A(n1049), .B(n2573), .Z(n2598) );
  AND U3408 ( .A(n2599), .B(n2600), .Z(n2597) );
  NANDN U3409 ( .B(n1118), .A(n2570), .Z(n2600) );
  NAND U3410 ( .A(n2576), .B(\u_a23_mem/p_mem[53][6] ), .Z(n2599) );
  NAND U3411 ( .A(n2601), .B(n2602), .Z(\u_a23_mem/n18989 ) );
  NANDN U3412 ( .B(n2573), .A(n1055), .Z(n2602) );
  NAND U3413 ( .A(n1121), .B(n2570), .Z(n2573) );
  AND U3414 ( .A(n2603), .B(n2604), .Z(n2601) );
  NANDN U3415 ( .B(n1124), .A(n2570), .Z(n2604) );
  NAND U3416 ( .A(n2576), .B(\u_a23_mem/p_mem[53][7] ), .Z(n2603) );
  NANDN U3417 ( .B(n1125), .A(n2570), .Z(n2576) );
  NAND U3418 ( .A(n2605), .B(n2606), .Z(\u_a23_mem/n18988 ) );
  OR U3419 ( .A(n1011), .B(n2607), .Z(n2606) );
  AND U3420 ( .A(n2608), .B(n2609), .Z(n2605) );
  NANDN U3421 ( .B(n1131), .A(n2570), .Z(n2609) );
  NAND U3422 ( .A(n2610), .B(\u_a23_mem/p_mem[54][0] ), .Z(n2608) );
  NAND U3423 ( .A(n2611), .B(n2612), .Z(\u_a23_mem/n18987 ) );
  OR U3424 ( .A(n1019), .B(n2607), .Z(n2612) );
  AND U3425 ( .A(n2613), .B(n2614), .Z(n2611) );
  NANDN U3426 ( .B(n1137), .A(n2570), .Z(n2614) );
  NAND U3427 ( .A(n2610), .B(\u_a23_mem/p_mem[54][1] ), .Z(n2613) );
  NAND U3428 ( .A(n2615), .B(n2616), .Z(\u_a23_mem/n18986 ) );
  OR U3429 ( .A(n1025), .B(n2607), .Z(n2616) );
  AND U3430 ( .A(n2617), .B(n2618), .Z(n2615) );
  NANDN U3431 ( .B(n1142), .A(n2570), .Z(n2618) );
  NAND U3432 ( .A(n2610), .B(\u_a23_mem/p_mem[54][2] ), .Z(n2617) );
  NAND U3433 ( .A(n2619), .B(n2620), .Z(\u_a23_mem/n18985 ) );
  OR U3434 ( .A(n1031), .B(n2607), .Z(n2620) );
  AND U3435 ( .A(n2621), .B(n2622), .Z(n2619) );
  NANDN U3436 ( .B(n1147), .A(n2570), .Z(n2622) );
  NAND U3437 ( .A(n2610), .B(\u_a23_mem/p_mem[54][3] ), .Z(n2621) );
  NAND U3438 ( .A(n2623), .B(n2624), .Z(\u_a23_mem/n18984 ) );
  OR U3439 ( .A(n1037), .B(n2607), .Z(n2624) );
  AND U3440 ( .A(n2625), .B(n2626), .Z(n2623) );
  NANDN U3441 ( .B(n1152), .A(n2570), .Z(n2626) );
  NAND U3442 ( .A(n2610), .B(\u_a23_mem/p_mem[54][4] ), .Z(n2625) );
  NAND U3443 ( .A(n2627), .B(n2628), .Z(\u_a23_mem/n18983 ) );
  OR U3444 ( .A(n1043), .B(n2607), .Z(n2628) );
  AND U3445 ( .A(n2629), .B(n2630), .Z(n2627) );
  NANDN U3446 ( .B(n1157), .A(n2570), .Z(n2630) );
  NAND U3447 ( .A(n2610), .B(\u_a23_mem/p_mem[54][5] ), .Z(n2629) );
  NAND U3448 ( .A(n2631), .B(n2632), .Z(\u_a23_mem/n18982 ) );
  OR U3449 ( .A(n1049), .B(n2607), .Z(n2632) );
  AND U3450 ( .A(n2633), .B(n2634), .Z(n2631) );
  NANDN U3451 ( .B(n1162), .A(n2570), .Z(n2634) );
  NAND U3452 ( .A(n2610), .B(\u_a23_mem/p_mem[54][6] ), .Z(n2633) );
  NAND U3453 ( .A(n2635), .B(n2636), .Z(\u_a23_mem/n18981 ) );
  NANDN U3454 ( .B(n2607), .A(n1055), .Z(n2636) );
  NAND U3455 ( .A(n1165), .B(n2570), .Z(n2607) );
  AND U3456 ( .A(n2637), .B(n2638), .Z(n2635) );
  NANDN U3457 ( .B(n1168), .A(n2570), .Z(n2638) );
  NAND U3458 ( .A(n2610), .B(\u_a23_mem/p_mem[54][7] ), .Z(n2637) );
  NANDN U3459 ( .B(n1169), .A(n2570), .Z(n2610) );
  NAND U3460 ( .A(n2639), .B(n2640), .Z(\u_a23_mem/n18980 ) );
  OR U3461 ( .A(n1011), .B(n2641), .Z(n2640) );
  AND U3462 ( .A(n2642), .B(n2643), .Z(n2639) );
  NAND U3463 ( .A(n2644), .B(\u_a23_mem/p_mem[55][0] ), .Z(n2643) );
  NANDN U3464 ( .B(n1015), .A(n2570), .Z(n2642) );
  NAND U3465 ( .A(n2645), .B(n2646), .Z(\u_a23_mem/n18979 ) );
  OR U3466 ( .A(n1019), .B(n2641), .Z(n2646) );
  AND U3467 ( .A(n2647), .B(n2648), .Z(n2645) );
  NAND U3468 ( .A(n2644), .B(\u_a23_mem/p_mem[55][1] ), .Z(n2648) );
  NANDN U3469 ( .B(n1022), .A(n2570), .Z(n2647) );
  NAND U3470 ( .A(n2649), .B(n2650), .Z(\u_a23_mem/n18978 ) );
  OR U3471 ( .A(n1025), .B(n2641), .Z(n2650) );
  AND U3472 ( .A(n2651), .B(n2652), .Z(n2649) );
  NAND U3473 ( .A(n2644), .B(\u_a23_mem/p_mem[55][2] ), .Z(n2652) );
  NANDN U3474 ( .B(n1028), .A(n2570), .Z(n2651) );
  NAND U3475 ( .A(n2653), .B(n2654), .Z(\u_a23_mem/n18977 ) );
  OR U3476 ( .A(n1031), .B(n2641), .Z(n2654) );
  AND U3477 ( .A(n2655), .B(n2656), .Z(n2653) );
  NAND U3478 ( .A(n2644), .B(\u_a23_mem/p_mem[55][3] ), .Z(n2656) );
  NANDN U3479 ( .B(n1034), .A(n2570), .Z(n2655) );
  NAND U3480 ( .A(n2657), .B(n2658), .Z(\u_a23_mem/n18976 ) );
  OR U3481 ( .A(n1037), .B(n2641), .Z(n2658) );
  AND U3482 ( .A(n2659), .B(n2660), .Z(n2657) );
  NAND U3483 ( .A(n2644), .B(\u_a23_mem/p_mem[55][4] ), .Z(n2660) );
  NANDN U3484 ( .B(n1040), .A(n2570), .Z(n2659) );
  NAND U3485 ( .A(n2661), .B(n2662), .Z(\u_a23_mem/n18975 ) );
  OR U3486 ( .A(n1043), .B(n2641), .Z(n2662) );
  AND U3487 ( .A(n2663), .B(n2664), .Z(n2661) );
  NAND U3488 ( .A(n2644), .B(\u_a23_mem/p_mem[55][5] ), .Z(n2664) );
  NANDN U3489 ( .B(n1046), .A(n2570), .Z(n2663) );
  NAND U3490 ( .A(n2665), .B(n2666), .Z(\u_a23_mem/n18974 ) );
  OR U3491 ( .A(n1049), .B(n2641), .Z(n2666) );
  AND U3492 ( .A(n2667), .B(n2668), .Z(n2665) );
  NAND U3493 ( .A(n2644), .B(\u_a23_mem/p_mem[55][6] ), .Z(n2668) );
  NANDN U3494 ( .B(n1052), .A(n2570), .Z(n2667) );
  NAND U3495 ( .A(n2669), .B(n2670), .Z(\u_a23_mem/n18973 ) );
  NANDN U3496 ( .B(n2641), .A(n1055), .Z(n2670) );
  NAND U3497 ( .A(n1056), .B(n2570), .Z(n2641) );
  AND U3498 ( .A(n2671), .B(n2672), .Z(n2669) );
  NAND U3499 ( .A(n2644), .B(\u_a23_mem/p_mem[55][7] ), .Z(n2672) );
  NANDN U3500 ( .B(n1059), .A(n2570), .Z(n2644) );
  NAND U3501 ( .A(n1061), .B(n2570), .Z(n2671) );
  AND U3502 ( .A(n1694), .B(n2673), .Z(n2570) );
  NAND U3503 ( .A(n2674), .B(n2675), .Z(\u_a23_mem/n18972 ) );
  NAND U3504 ( .A(n2676), .B(\u_a23_mem/p_mem[56][0] ), .Z(n2675) );
  OR U3505 ( .A(n1011), .B(n2677), .Z(n2674) );
  NAND U3506 ( .A(n2678), .B(n2679), .Z(\u_a23_mem/n18971 ) );
  NAND U3507 ( .A(n2676), .B(\u_a23_mem/p_mem[56][1] ), .Z(n2679) );
  OR U3508 ( .A(n1019), .B(n2677), .Z(n2678) );
  NAND U3509 ( .A(n2680), .B(n2681), .Z(\u_a23_mem/n18970 ) );
  NAND U3510 ( .A(n2676), .B(\u_a23_mem/p_mem[56][2] ), .Z(n2681) );
  OR U3511 ( .A(n1025), .B(n2677), .Z(n2680) );
  NAND U3512 ( .A(n2682), .B(n2683), .Z(\u_a23_mem/n18969 ) );
  NAND U3513 ( .A(n2676), .B(\u_a23_mem/p_mem[56][3] ), .Z(n2683) );
  OR U3514 ( .A(n1031), .B(n2677), .Z(n2682) );
  NAND U3515 ( .A(n2684), .B(n2685), .Z(\u_a23_mem/n18968 ) );
  NAND U3516 ( .A(n2676), .B(\u_a23_mem/p_mem[56][4] ), .Z(n2685) );
  OR U3517 ( .A(n1037), .B(n2677), .Z(n2684) );
  NAND U3518 ( .A(n2686), .B(n2687), .Z(\u_a23_mem/n18967 ) );
  NAND U3519 ( .A(n2676), .B(\u_a23_mem/p_mem[56][5] ), .Z(n2687) );
  OR U3520 ( .A(n1043), .B(n2677), .Z(n2686) );
  NAND U3521 ( .A(n2688), .B(n2689), .Z(\u_a23_mem/n18966 ) );
  NAND U3522 ( .A(n2676), .B(\u_a23_mem/p_mem[56][6] ), .Z(n2689) );
  OR U3523 ( .A(n1049), .B(n2677), .Z(n2688) );
  NAND U3524 ( .A(n2690), .B(n2691), .Z(\u_a23_mem/n18965 ) );
  NAND U3525 ( .A(n2676), .B(\u_a23_mem/p_mem[56][7] ), .Z(n2691) );
  NANDN U3526 ( .B(n1080), .A(n2692), .Z(n2676) );
  NANDN U3527 ( .B(n2677), .A(n1055), .Z(n2690) );
  NANDN U3528 ( .B(n2), .A(n2692), .Z(n2677) );
  NAND U3529 ( .A(n2693), .B(n2694), .Z(\u_a23_mem/n18964 ) );
  OR U3530 ( .A(n1011), .B(n2695), .Z(n2694) );
  AND U3531 ( .A(n2696), .B(n2697), .Z(n2693) );
  NANDN U3532 ( .B(n1087), .A(n2692), .Z(n2697) );
  NAND U3533 ( .A(n2698), .B(\u_a23_mem/p_mem[57][0] ), .Z(n2696) );
  NAND U3534 ( .A(n2699), .B(n2700), .Z(\u_a23_mem/n18963 ) );
  OR U3535 ( .A(n1019), .B(n2695), .Z(n2700) );
  AND U3536 ( .A(n2701), .B(n2702), .Z(n2699) );
  NANDN U3537 ( .B(n1093), .A(n2692), .Z(n2702) );
  NAND U3538 ( .A(n2698), .B(\u_a23_mem/p_mem[57][1] ), .Z(n2701) );
  NAND U3539 ( .A(n2703), .B(n2704), .Z(\u_a23_mem/n18962 ) );
  OR U3540 ( .A(n1025), .B(n2695), .Z(n2704) );
  AND U3541 ( .A(n2705), .B(n2706), .Z(n2703) );
  NANDN U3542 ( .B(n1098), .A(n2692), .Z(n2706) );
  NAND U3543 ( .A(n2698), .B(\u_a23_mem/p_mem[57][2] ), .Z(n2705) );
  NAND U3544 ( .A(n2707), .B(n2708), .Z(\u_a23_mem/n18961 ) );
  OR U3545 ( .A(n1031), .B(n2695), .Z(n2708) );
  AND U3546 ( .A(n2709), .B(n2710), .Z(n2707) );
  NANDN U3547 ( .B(n1103), .A(n2692), .Z(n2710) );
  NAND U3548 ( .A(n2698), .B(\u_a23_mem/p_mem[57][3] ), .Z(n2709) );
  NAND U3549 ( .A(n2711), .B(n2712), .Z(\u_a23_mem/n18960 ) );
  OR U3550 ( .A(n1037), .B(n2695), .Z(n2712) );
  AND U3551 ( .A(n2713), .B(n2714), .Z(n2711) );
  NANDN U3552 ( .B(n1108), .A(n2692), .Z(n2714) );
  NAND U3553 ( .A(n2698), .B(\u_a23_mem/p_mem[57][4] ), .Z(n2713) );
  NAND U3554 ( .A(n2715), .B(n2716), .Z(\u_a23_mem/n18959 ) );
  OR U3555 ( .A(n1043), .B(n2695), .Z(n2716) );
  AND U3556 ( .A(n2717), .B(n2718), .Z(n2715) );
  NANDN U3557 ( .B(n1113), .A(n2692), .Z(n2718) );
  NAND U3558 ( .A(n2698), .B(\u_a23_mem/p_mem[57][5] ), .Z(n2717) );
  NAND U3559 ( .A(n2719), .B(n2720), .Z(\u_a23_mem/n18958 ) );
  OR U3560 ( .A(n1049), .B(n2695), .Z(n2720) );
  AND U3561 ( .A(n2721), .B(n2722), .Z(n2719) );
  NANDN U3562 ( .B(n1118), .A(n2692), .Z(n2722) );
  NAND U3563 ( .A(n2698), .B(\u_a23_mem/p_mem[57][6] ), .Z(n2721) );
  NAND U3564 ( .A(n2723), .B(n2724), .Z(\u_a23_mem/n18957 ) );
  NANDN U3565 ( .B(n2695), .A(n1055), .Z(n2724) );
  NAND U3566 ( .A(n1121), .B(n2692), .Z(n2695) );
  AND U3567 ( .A(n2725), .B(n2726), .Z(n2723) );
  NANDN U3568 ( .B(n1124), .A(n2692), .Z(n2726) );
  NAND U3569 ( .A(n2698), .B(\u_a23_mem/p_mem[57][7] ), .Z(n2725) );
  NANDN U3570 ( .B(n1125), .A(n2692), .Z(n2698) );
  NAND U3571 ( .A(n2727), .B(n2728), .Z(\u_a23_mem/n18956 ) );
  OR U3572 ( .A(n1011), .B(n2729), .Z(n2728) );
  AND U3573 ( .A(n2730), .B(n2731), .Z(n2727) );
  NANDN U3574 ( .B(n1131), .A(n2692), .Z(n2731) );
  NAND U3575 ( .A(n2732), .B(\u_a23_mem/p_mem[58][0] ), .Z(n2730) );
  NAND U3576 ( .A(n2733), .B(n2734), .Z(\u_a23_mem/n18955 ) );
  OR U3577 ( .A(n1019), .B(n2729), .Z(n2734) );
  AND U3578 ( .A(n2735), .B(n2736), .Z(n2733) );
  NANDN U3579 ( .B(n1137), .A(n2692), .Z(n2736) );
  NAND U3580 ( .A(n2732), .B(\u_a23_mem/p_mem[58][1] ), .Z(n2735) );
  NAND U3581 ( .A(n2737), .B(n2738), .Z(\u_a23_mem/n18954 ) );
  OR U3582 ( .A(n1025), .B(n2729), .Z(n2738) );
  AND U3583 ( .A(n2739), .B(n2740), .Z(n2737) );
  NANDN U3584 ( .B(n1142), .A(n2692), .Z(n2740) );
  NAND U3585 ( .A(n2732), .B(\u_a23_mem/p_mem[58][2] ), .Z(n2739) );
  NAND U3586 ( .A(n2741), .B(n2742), .Z(\u_a23_mem/n18953 ) );
  OR U3587 ( .A(n1031), .B(n2729), .Z(n2742) );
  AND U3588 ( .A(n2743), .B(n2744), .Z(n2741) );
  NANDN U3589 ( .B(n1147), .A(n2692), .Z(n2744) );
  NAND U3590 ( .A(n2732), .B(\u_a23_mem/p_mem[58][3] ), .Z(n2743) );
  NAND U3591 ( .A(n2745), .B(n2746), .Z(\u_a23_mem/n18952 ) );
  OR U3592 ( .A(n1037), .B(n2729), .Z(n2746) );
  AND U3593 ( .A(n2747), .B(n2748), .Z(n2745) );
  NANDN U3594 ( .B(n1152), .A(n2692), .Z(n2748) );
  NAND U3595 ( .A(n2732), .B(\u_a23_mem/p_mem[58][4] ), .Z(n2747) );
  NAND U3596 ( .A(n2749), .B(n2750), .Z(\u_a23_mem/n18951 ) );
  OR U3597 ( .A(n1043), .B(n2729), .Z(n2750) );
  AND U3598 ( .A(n2751), .B(n2752), .Z(n2749) );
  NANDN U3599 ( .B(n1157), .A(n2692), .Z(n2752) );
  NAND U3600 ( .A(n2732), .B(\u_a23_mem/p_mem[58][5] ), .Z(n2751) );
  NAND U3601 ( .A(n2753), .B(n2754), .Z(\u_a23_mem/n18950 ) );
  OR U3602 ( .A(n1049), .B(n2729), .Z(n2754) );
  AND U3603 ( .A(n2755), .B(n2756), .Z(n2753) );
  NANDN U3604 ( .B(n1162), .A(n2692), .Z(n2756) );
  NAND U3605 ( .A(n2732), .B(\u_a23_mem/p_mem[58][6] ), .Z(n2755) );
  NAND U3606 ( .A(n2757), .B(n2758), .Z(\u_a23_mem/n18949 ) );
  NANDN U3607 ( .B(n2729), .A(n1055), .Z(n2758) );
  NAND U3608 ( .A(n1165), .B(n2692), .Z(n2729) );
  AND U3609 ( .A(n2759), .B(n2760), .Z(n2757) );
  NANDN U3610 ( .B(n1168), .A(n2692), .Z(n2760) );
  NAND U3611 ( .A(n2732), .B(\u_a23_mem/p_mem[58][7] ), .Z(n2759) );
  NANDN U3612 ( .B(n1169), .A(n2692), .Z(n2732) );
  NAND U3613 ( .A(n2761), .B(n2762), .Z(\u_a23_mem/n18948 ) );
  OR U3614 ( .A(n1011), .B(n2763), .Z(n2762) );
  AND U3615 ( .A(n2764), .B(n2765), .Z(n2761) );
  NAND U3616 ( .A(n2766), .B(\u_a23_mem/p_mem[59][0] ), .Z(n2765) );
  NANDN U3617 ( .B(n1015), .A(n2692), .Z(n2764) );
  NAND U3618 ( .A(n2767), .B(n2768), .Z(\u_a23_mem/n18947 ) );
  OR U3619 ( .A(n1019), .B(n2763), .Z(n2768) );
  AND U3620 ( .A(n2769), .B(n2770), .Z(n2767) );
  NAND U3621 ( .A(n2766), .B(\u_a23_mem/p_mem[59][1] ), .Z(n2770) );
  NANDN U3622 ( .B(n1022), .A(n2692), .Z(n2769) );
  NAND U3623 ( .A(n2771), .B(n2772), .Z(\u_a23_mem/n18946 ) );
  OR U3624 ( .A(n1025), .B(n2763), .Z(n2772) );
  AND U3625 ( .A(n2773), .B(n2774), .Z(n2771) );
  NAND U3626 ( .A(n2766), .B(\u_a23_mem/p_mem[59][2] ), .Z(n2774) );
  NANDN U3627 ( .B(n1028), .A(n2692), .Z(n2773) );
  NAND U3628 ( .A(n2775), .B(n2776), .Z(\u_a23_mem/n18945 ) );
  OR U3629 ( .A(n1031), .B(n2763), .Z(n2776) );
  AND U3630 ( .A(n2777), .B(n2778), .Z(n2775) );
  NAND U3631 ( .A(n2766), .B(\u_a23_mem/p_mem[59][3] ), .Z(n2778) );
  NANDN U3632 ( .B(n1034), .A(n2692), .Z(n2777) );
  NAND U3633 ( .A(n2779), .B(n2780), .Z(\u_a23_mem/n18944 ) );
  OR U3634 ( .A(n1037), .B(n2763), .Z(n2780) );
  AND U3635 ( .A(n2781), .B(n2782), .Z(n2779) );
  NAND U3636 ( .A(n2766), .B(\u_a23_mem/p_mem[59][4] ), .Z(n2782) );
  NANDN U3637 ( .B(n1040), .A(n2692), .Z(n2781) );
  NAND U3638 ( .A(n2783), .B(n2784), .Z(\u_a23_mem/n18943 ) );
  OR U3639 ( .A(n1043), .B(n2763), .Z(n2784) );
  AND U3640 ( .A(n2785), .B(n2786), .Z(n2783) );
  NAND U3641 ( .A(n2766), .B(\u_a23_mem/p_mem[59][5] ), .Z(n2786) );
  NANDN U3642 ( .B(n1046), .A(n2692), .Z(n2785) );
  NAND U3643 ( .A(n2787), .B(n2788), .Z(\u_a23_mem/n18942 ) );
  OR U3644 ( .A(n1049), .B(n2763), .Z(n2788) );
  AND U3645 ( .A(n2789), .B(n2790), .Z(n2787) );
  NAND U3646 ( .A(n2766), .B(\u_a23_mem/p_mem[59][6] ), .Z(n2790) );
  NANDN U3647 ( .B(n1052), .A(n2692), .Z(n2789) );
  NAND U3648 ( .A(n2791), .B(n2792), .Z(\u_a23_mem/n18941 ) );
  NANDN U3649 ( .B(n2763), .A(n1055), .Z(n2792) );
  NAND U3650 ( .A(n1056), .B(n2692), .Z(n2763) );
  AND U3651 ( .A(n2793), .B(n2794), .Z(n2791) );
  NAND U3652 ( .A(n2766), .B(\u_a23_mem/p_mem[59][7] ), .Z(n2794) );
  NANDN U3653 ( .B(n1059), .A(n2692), .Z(n2766) );
  NAND U3654 ( .A(n1061), .B(n2692), .Z(n2793) );
  AND U3655 ( .A(n1816), .B(n2673), .Z(n2692) );
  NAND U3656 ( .A(n2795), .B(n2796), .Z(\u_a23_mem/n18940 ) );
  NAND U3657 ( .A(n2797), .B(\u_a23_mem/p_mem[60][0] ), .Z(n2796) );
  OR U3658 ( .A(n1011), .B(n2798), .Z(n2795) );
  NAND U3659 ( .A(n2799), .B(n2800), .Z(\u_a23_mem/n18939 ) );
  NAND U3660 ( .A(n2797), .B(\u_a23_mem/p_mem[60][1] ), .Z(n2800) );
  OR U3661 ( .A(n1019), .B(n2798), .Z(n2799) );
  NAND U3662 ( .A(n2801), .B(n2802), .Z(\u_a23_mem/n18938 ) );
  NAND U3663 ( .A(n2797), .B(\u_a23_mem/p_mem[60][2] ), .Z(n2802) );
  OR U3664 ( .A(n1025), .B(n2798), .Z(n2801) );
  NAND U3665 ( .A(n2803), .B(n2804), .Z(\u_a23_mem/n18937 ) );
  NAND U3666 ( .A(n2797), .B(\u_a23_mem/p_mem[60][3] ), .Z(n2804) );
  OR U3667 ( .A(n1031), .B(n2798), .Z(n2803) );
  NAND U3668 ( .A(n2805), .B(n2806), .Z(\u_a23_mem/n18936 ) );
  NAND U3669 ( .A(n2797), .B(\u_a23_mem/p_mem[60][4] ), .Z(n2806) );
  OR U3670 ( .A(n1037), .B(n2798), .Z(n2805) );
  NAND U3671 ( .A(n2807), .B(n2808), .Z(\u_a23_mem/n18935 ) );
  NAND U3672 ( .A(n2797), .B(\u_a23_mem/p_mem[60][5] ), .Z(n2808) );
  OR U3673 ( .A(n1043), .B(n2798), .Z(n2807) );
  NAND U3674 ( .A(n2809), .B(n2810), .Z(\u_a23_mem/n18934 ) );
  NAND U3675 ( .A(n2797), .B(\u_a23_mem/p_mem[60][6] ), .Z(n2810) );
  OR U3676 ( .A(n1049), .B(n2798), .Z(n2809) );
  NAND U3677 ( .A(n2811), .B(n2812), .Z(\u_a23_mem/n18933 ) );
  NAND U3678 ( .A(n2797), .B(\u_a23_mem/p_mem[60][7] ), .Z(n2812) );
  NANDN U3679 ( .B(n1080), .A(n2813), .Z(n2797) );
  NANDN U3680 ( .B(n2798), .A(n1055), .Z(n2811) );
  NANDN U3681 ( .B(n2), .A(n2813), .Z(n2798) );
  NAND U3682 ( .A(n2814), .B(n2815), .Z(\u_a23_mem/n18932 ) );
  OR U3683 ( .A(n1011), .B(n2816), .Z(n2815) );
  AND U3684 ( .A(n2817), .B(n2818), .Z(n2814) );
  NANDN U3685 ( .B(n1087), .A(n2813), .Z(n2818) );
  NAND U3686 ( .A(n2819), .B(\u_a23_mem/p_mem[61][0] ), .Z(n2817) );
  NAND U3687 ( .A(n2820), .B(n2821), .Z(\u_a23_mem/n18931 ) );
  OR U3688 ( .A(n1019), .B(n2816), .Z(n2821) );
  AND U3689 ( .A(n2822), .B(n2823), .Z(n2820) );
  NANDN U3690 ( .B(n1093), .A(n2813), .Z(n2823) );
  NAND U3691 ( .A(n2819), .B(\u_a23_mem/p_mem[61][1] ), .Z(n2822) );
  NAND U3692 ( .A(n2824), .B(n2825), .Z(\u_a23_mem/n18930 ) );
  OR U3693 ( .A(n1025), .B(n2816), .Z(n2825) );
  AND U3694 ( .A(n2826), .B(n2827), .Z(n2824) );
  NANDN U3695 ( .B(n1098), .A(n2813), .Z(n2827) );
  NAND U3696 ( .A(n2819), .B(\u_a23_mem/p_mem[61][2] ), .Z(n2826) );
  NAND U3697 ( .A(n2828), .B(n2829), .Z(\u_a23_mem/n18929 ) );
  OR U3698 ( .A(n1031), .B(n2816), .Z(n2829) );
  AND U3699 ( .A(n2830), .B(n2831), .Z(n2828) );
  NANDN U3700 ( .B(n1103), .A(n2813), .Z(n2831) );
  NAND U3701 ( .A(n2819), .B(\u_a23_mem/p_mem[61][3] ), .Z(n2830) );
  NAND U3702 ( .A(n2832), .B(n2833), .Z(\u_a23_mem/n18928 ) );
  OR U3703 ( .A(n1037), .B(n2816), .Z(n2833) );
  AND U3704 ( .A(n2834), .B(n2835), .Z(n2832) );
  NANDN U3705 ( .B(n1108), .A(n2813), .Z(n2835) );
  NAND U3706 ( .A(n2819), .B(\u_a23_mem/p_mem[61][4] ), .Z(n2834) );
  NAND U3707 ( .A(n2836), .B(n2837), .Z(\u_a23_mem/n18927 ) );
  OR U3708 ( .A(n1043), .B(n2816), .Z(n2837) );
  AND U3709 ( .A(n2838), .B(n2839), .Z(n2836) );
  NANDN U3710 ( .B(n1113), .A(n2813), .Z(n2839) );
  NAND U3711 ( .A(n2819), .B(\u_a23_mem/p_mem[61][5] ), .Z(n2838) );
  NAND U3712 ( .A(n2840), .B(n2841), .Z(\u_a23_mem/n18926 ) );
  OR U3713 ( .A(n1049), .B(n2816), .Z(n2841) );
  AND U3714 ( .A(n2842), .B(n2843), .Z(n2840) );
  NANDN U3715 ( .B(n1118), .A(n2813), .Z(n2843) );
  NAND U3716 ( .A(n2819), .B(\u_a23_mem/p_mem[61][6] ), .Z(n2842) );
  NAND U3717 ( .A(n2844), .B(n2845), .Z(\u_a23_mem/n18925 ) );
  NANDN U3718 ( .B(n2816), .A(n1055), .Z(n2845) );
  NAND U3719 ( .A(n1121), .B(n2813), .Z(n2816) );
  AND U3720 ( .A(n2846), .B(n2847), .Z(n2844) );
  NANDN U3721 ( .B(n1124), .A(n2813), .Z(n2847) );
  NAND U3722 ( .A(n2819), .B(\u_a23_mem/p_mem[61][7] ), .Z(n2846) );
  NANDN U3723 ( .B(n1125), .A(n2813), .Z(n2819) );
  NAND U3724 ( .A(n2848), .B(n2849), .Z(\u_a23_mem/n18924 ) );
  OR U3725 ( .A(n1011), .B(n2850), .Z(n2849) );
  AND U3726 ( .A(n2851), .B(n2852), .Z(n2848) );
  NANDN U3727 ( .B(n1131), .A(n2813), .Z(n2852) );
  NAND U3728 ( .A(n2853), .B(\u_a23_mem/p_mem[62][0] ), .Z(n2851) );
  NAND U3729 ( .A(n2854), .B(n2855), .Z(\u_a23_mem/n18923 ) );
  OR U3730 ( .A(n1019), .B(n2850), .Z(n2855) );
  AND U3731 ( .A(n2856), .B(n2857), .Z(n2854) );
  NANDN U3732 ( .B(n1137), .A(n2813), .Z(n2857) );
  NAND U3733 ( .A(n2853), .B(\u_a23_mem/p_mem[62][1] ), .Z(n2856) );
  NAND U3734 ( .A(n2858), .B(n2859), .Z(\u_a23_mem/n18922 ) );
  OR U3735 ( .A(n1025), .B(n2850), .Z(n2859) );
  AND U3736 ( .A(n2860), .B(n2861), .Z(n2858) );
  NANDN U3737 ( .B(n1142), .A(n2813), .Z(n2861) );
  NAND U3738 ( .A(n2853), .B(\u_a23_mem/p_mem[62][2] ), .Z(n2860) );
  NAND U3739 ( .A(n2862), .B(n2863), .Z(\u_a23_mem/n18921 ) );
  OR U3740 ( .A(n1031), .B(n2850), .Z(n2863) );
  AND U3741 ( .A(n2864), .B(n2865), .Z(n2862) );
  NANDN U3742 ( .B(n1147), .A(n2813), .Z(n2865) );
  NAND U3743 ( .A(n2853), .B(\u_a23_mem/p_mem[62][3] ), .Z(n2864) );
  NAND U3744 ( .A(n2866), .B(n2867), .Z(\u_a23_mem/n18920 ) );
  OR U3745 ( .A(n1037), .B(n2850), .Z(n2867) );
  AND U3746 ( .A(n2868), .B(n2869), .Z(n2866) );
  NANDN U3747 ( .B(n1152), .A(n2813), .Z(n2869) );
  NAND U3748 ( .A(n2853), .B(\u_a23_mem/p_mem[62][4] ), .Z(n2868) );
  NAND U3749 ( .A(n2870), .B(n2871), .Z(\u_a23_mem/n18919 ) );
  OR U3750 ( .A(n1043), .B(n2850), .Z(n2871) );
  AND U3751 ( .A(n2872), .B(n2873), .Z(n2870) );
  NANDN U3752 ( .B(n1157), .A(n2813), .Z(n2873) );
  NAND U3753 ( .A(n2853), .B(\u_a23_mem/p_mem[62][5] ), .Z(n2872) );
  NAND U3754 ( .A(n2874), .B(n2875), .Z(\u_a23_mem/n18918 ) );
  OR U3755 ( .A(n1049), .B(n2850), .Z(n2875) );
  AND U3756 ( .A(n2876), .B(n2877), .Z(n2874) );
  NANDN U3757 ( .B(n1162), .A(n2813), .Z(n2877) );
  NAND U3758 ( .A(n2853), .B(\u_a23_mem/p_mem[62][6] ), .Z(n2876) );
  NAND U3759 ( .A(n2878), .B(n2879), .Z(\u_a23_mem/n18917 ) );
  NANDN U3760 ( .B(n2850), .A(n1055), .Z(n2879) );
  NAND U3761 ( .A(n1165), .B(n2813), .Z(n2850) );
  AND U3762 ( .A(n2880), .B(n2881), .Z(n2878) );
  NANDN U3763 ( .B(n1168), .A(n2813), .Z(n2881) );
  NAND U3764 ( .A(n2853), .B(\u_a23_mem/p_mem[62][7] ), .Z(n2880) );
  NANDN U3765 ( .B(n1169), .A(n2813), .Z(n2853) );
  NAND U3766 ( .A(n2882), .B(n2883), .Z(\u_a23_mem/n18916 ) );
  OR U3767 ( .A(n1011), .B(n2884), .Z(n2883) );
  AND U3768 ( .A(n2885), .B(n2886), .Z(n2882) );
  NAND U3769 ( .A(n2887), .B(\u_a23_mem/p_mem[63][0] ), .Z(n2886) );
  NANDN U3770 ( .B(n1015), .A(n2813), .Z(n2885) );
  NAND U3771 ( .A(n2888), .B(n2889), .Z(\u_a23_mem/n18915 ) );
  OR U3772 ( .A(n1019), .B(n2884), .Z(n2889) );
  AND U3773 ( .A(n2890), .B(n2891), .Z(n2888) );
  NAND U3774 ( .A(n2887), .B(\u_a23_mem/p_mem[63][1] ), .Z(n2891) );
  NANDN U3775 ( .B(n1022), .A(n2813), .Z(n2890) );
  NAND U3776 ( .A(n2892), .B(n2893), .Z(\u_a23_mem/n18914 ) );
  OR U3777 ( .A(n1025), .B(n2884), .Z(n2893) );
  AND U3778 ( .A(n2894), .B(n2895), .Z(n2892) );
  NAND U3779 ( .A(n2887), .B(\u_a23_mem/p_mem[63][2] ), .Z(n2895) );
  NANDN U3780 ( .B(n1028), .A(n2813), .Z(n2894) );
  NAND U3781 ( .A(n2896), .B(n2897), .Z(\u_a23_mem/n18913 ) );
  OR U3782 ( .A(n1031), .B(n2884), .Z(n2897) );
  AND U3783 ( .A(n2898), .B(n2899), .Z(n2896) );
  NAND U3784 ( .A(n2887), .B(\u_a23_mem/p_mem[63][3] ), .Z(n2899) );
  NANDN U3785 ( .B(n1034), .A(n2813), .Z(n2898) );
  NAND U3786 ( .A(n2900), .B(n2901), .Z(\u_a23_mem/n18912 ) );
  OR U3787 ( .A(n1037), .B(n2884), .Z(n2901) );
  AND U3788 ( .A(n2902), .B(n2903), .Z(n2900) );
  NAND U3789 ( .A(n2887), .B(\u_a23_mem/p_mem[63][4] ), .Z(n2903) );
  NANDN U3790 ( .B(n1040), .A(n2813), .Z(n2902) );
  NAND U3791 ( .A(n2904), .B(n2905), .Z(\u_a23_mem/n18911 ) );
  OR U3792 ( .A(n1043), .B(n2884), .Z(n2905) );
  AND U3793 ( .A(n2906), .B(n2907), .Z(n2904) );
  NAND U3794 ( .A(n2887), .B(\u_a23_mem/p_mem[63][5] ), .Z(n2907) );
  NANDN U3795 ( .B(n1046), .A(n2813), .Z(n2906) );
  NAND U3796 ( .A(n2908), .B(n2909), .Z(\u_a23_mem/n18910 ) );
  OR U3797 ( .A(n1049), .B(n2884), .Z(n2909) );
  AND U3798 ( .A(n2910), .B(n2911), .Z(n2908) );
  NAND U3799 ( .A(n2887), .B(\u_a23_mem/p_mem[63][6] ), .Z(n2911) );
  NANDN U3800 ( .B(n1052), .A(n2813), .Z(n2910) );
  NAND U3801 ( .A(n2912), .B(n2913), .Z(\u_a23_mem/n18909 ) );
  NANDN U3802 ( .B(n2884), .A(n1055), .Z(n2913) );
  NAND U3803 ( .A(n1056), .B(n2813), .Z(n2884) );
  AND U3804 ( .A(n2914), .B(n2915), .Z(n2912) );
  NAND U3805 ( .A(n2887), .B(\u_a23_mem/p_mem[63][7] ), .Z(n2915) );
  NANDN U3806 ( .B(n1059), .A(n2813), .Z(n2887) );
  NAND U3807 ( .A(n1061), .B(n2813), .Z(n2914) );
  NOR U3808 ( .A(n2551), .B(n1938), .Z(n2813) );
  IV U3809 ( .A(n2673), .Z(n2551) );
  ANDN U3810 ( .A(n2916), .B(n2428), .Z(n2673) );
  AND U3811 ( .A(n2429), .B(m_address[4]), .Z(n2916) );
  NAND U3812 ( .A(n2917), .B(n2918), .Z(\u_a23_mem/n18908 ) );
  NAND U3813 ( .A(n2919), .B(\u_a23_mem/p_mem[64][0] ), .Z(n2918) );
  OR U3814 ( .A(n1011), .B(n2920), .Z(n2917) );
  NAND U3815 ( .A(n2921), .B(n2922), .Z(\u_a23_mem/n18907 ) );
  NAND U3816 ( .A(n2919), .B(\u_a23_mem/p_mem[64][1] ), .Z(n2922) );
  OR U3817 ( .A(n1019), .B(n2920), .Z(n2921) );
  NAND U3818 ( .A(n2923), .B(n2924), .Z(\u_a23_mem/n18906 ) );
  NAND U3819 ( .A(n2919), .B(\u_a23_mem/p_mem[64][2] ), .Z(n2924) );
  OR U3820 ( .A(n1025), .B(n2920), .Z(n2923) );
  NAND U3821 ( .A(n2925), .B(n2926), .Z(\u_a23_mem/n18905 ) );
  NAND U3822 ( .A(n2919), .B(\u_a23_mem/p_mem[64][3] ), .Z(n2926) );
  OR U3823 ( .A(n1031), .B(n2920), .Z(n2925) );
  NAND U3824 ( .A(n2927), .B(n2928), .Z(\u_a23_mem/n18904 ) );
  NAND U3825 ( .A(n2919), .B(\u_a23_mem/p_mem[64][4] ), .Z(n2928) );
  OR U3826 ( .A(n1037), .B(n2920), .Z(n2927) );
  NAND U3827 ( .A(n2929), .B(n2930), .Z(\u_a23_mem/n18903 ) );
  NAND U3828 ( .A(n2919), .B(\u_a23_mem/p_mem[64][5] ), .Z(n2930) );
  OR U3829 ( .A(n1043), .B(n2920), .Z(n2929) );
  NAND U3830 ( .A(n2931), .B(n2932), .Z(\u_a23_mem/n18902 ) );
  NAND U3831 ( .A(n2919), .B(\u_a23_mem/p_mem[64][6] ), .Z(n2932) );
  OR U3832 ( .A(n1049), .B(n2920), .Z(n2931) );
  NAND U3833 ( .A(n2933), .B(n2934), .Z(\u_a23_mem/n18901 ) );
  NAND U3834 ( .A(n2919), .B(\u_a23_mem/p_mem[64][7] ), .Z(n2934) );
  NAND U3835 ( .A(n2935), .B(n2936), .Z(n2919) );
  AND U3836 ( .A(n2937), .B(n2938), .Z(n2935) );
  NANDN U3837 ( .B(n2920), .A(n1055), .Z(n2933) );
  NANDN U3838 ( .B(n2), .A(n2939), .Z(n2920) );
  NAND U3839 ( .A(n2940), .B(n2941), .Z(\u_a23_mem/n18900 ) );
  OR U3840 ( .A(n1011), .B(n2942), .Z(n2941) );
  AND U3841 ( .A(n2943), .B(n2944), .Z(n2940) );
  NANDN U3842 ( .B(n1087), .A(n2939), .Z(n2944) );
  NAND U3843 ( .A(n2945), .B(\u_a23_mem/p_mem[65][0] ), .Z(n2943) );
  NAND U3844 ( .A(n2946), .B(n2947), .Z(\u_a23_mem/n18899 ) );
  OR U3845 ( .A(n1019), .B(n2942), .Z(n2947) );
  AND U3846 ( .A(n2948), .B(n2949), .Z(n2946) );
  NANDN U3847 ( .B(n1093), .A(n2939), .Z(n2949) );
  NAND U3848 ( .A(n2945), .B(\u_a23_mem/p_mem[65][1] ), .Z(n2948) );
  NAND U3849 ( .A(n2950), .B(n2951), .Z(\u_a23_mem/n18898 ) );
  OR U3850 ( .A(n1025), .B(n2942), .Z(n2951) );
  AND U3851 ( .A(n2952), .B(n2953), .Z(n2950) );
  NANDN U3852 ( .B(n1098), .A(n2939), .Z(n2953) );
  NAND U3853 ( .A(n2945), .B(\u_a23_mem/p_mem[65][2] ), .Z(n2952) );
  NAND U3854 ( .A(n2954), .B(n2955), .Z(\u_a23_mem/n18897 ) );
  OR U3855 ( .A(n1031), .B(n2942), .Z(n2955) );
  AND U3856 ( .A(n2956), .B(n2957), .Z(n2954) );
  NANDN U3857 ( .B(n1103), .A(n2939), .Z(n2957) );
  NAND U3858 ( .A(n2945), .B(\u_a23_mem/p_mem[65][3] ), .Z(n2956) );
  NAND U3859 ( .A(n2958), .B(n2959), .Z(\u_a23_mem/n18896 ) );
  OR U3860 ( .A(n1037), .B(n2942), .Z(n2959) );
  AND U3861 ( .A(n2960), .B(n2961), .Z(n2958) );
  NANDN U3862 ( .B(n1108), .A(n2939), .Z(n2961) );
  NAND U3863 ( .A(n2945), .B(\u_a23_mem/p_mem[65][4] ), .Z(n2960) );
  NAND U3864 ( .A(n2962), .B(n2963), .Z(\u_a23_mem/n18895 ) );
  OR U3865 ( .A(n1043), .B(n2942), .Z(n2963) );
  AND U3866 ( .A(n2964), .B(n2965), .Z(n2962) );
  NANDN U3867 ( .B(n1113), .A(n2939), .Z(n2965) );
  NAND U3868 ( .A(n2945), .B(\u_a23_mem/p_mem[65][5] ), .Z(n2964) );
  NAND U3869 ( .A(n2966), .B(n2967), .Z(\u_a23_mem/n18894 ) );
  OR U3870 ( .A(n1049), .B(n2942), .Z(n2967) );
  AND U3871 ( .A(n2968), .B(n2969), .Z(n2966) );
  NANDN U3872 ( .B(n1118), .A(n2939), .Z(n2969) );
  NAND U3873 ( .A(n2945), .B(\u_a23_mem/p_mem[65][6] ), .Z(n2968) );
  NAND U3874 ( .A(n2970), .B(n2971), .Z(\u_a23_mem/n18893 ) );
  NANDN U3875 ( .B(n2942), .A(n1055), .Z(n2971) );
  NAND U3876 ( .A(n1121), .B(n2939), .Z(n2942) );
  AND U3877 ( .A(n2972), .B(n2973), .Z(n2970) );
  NANDN U3878 ( .B(n1124), .A(n2939), .Z(n2973) );
  NAND U3879 ( .A(n2945), .B(\u_a23_mem/p_mem[65][7] ), .Z(n2972) );
  NAND U3880 ( .A(n2974), .B(n2936), .Z(n2945) );
  AND U3881 ( .A(n2975), .B(n2976), .Z(n2936) );
  AND U3882 ( .A(n2977), .B(n2978), .Z(n2976) );
  ANDN U3883 ( .A(n2939), .B(n2979), .Z(n2975) );
  AND U3884 ( .A(n2980), .B(n2938), .Z(n2974) );
  NAND U3885 ( .A(n2981), .B(n2982), .Z(\u_a23_mem/n18892 ) );
  OR U3886 ( .A(n1011), .B(n2983), .Z(n2982) );
  AND U3887 ( .A(n2984), .B(n2985), .Z(n2981) );
  NANDN U3888 ( .B(n1131), .A(n2939), .Z(n2985) );
  NAND U3889 ( .A(n2986), .B(\u_a23_mem/p_mem[66][0] ), .Z(n2984) );
  NAND U3890 ( .A(n2987), .B(n2988), .Z(\u_a23_mem/n18891 ) );
  OR U3891 ( .A(n1019), .B(n2983), .Z(n2988) );
  AND U3892 ( .A(n2989), .B(n2990), .Z(n2987) );
  NANDN U3893 ( .B(n1137), .A(n2939), .Z(n2990) );
  NAND U3894 ( .A(n2986), .B(\u_a23_mem/p_mem[66][1] ), .Z(n2989) );
  NAND U3895 ( .A(n2991), .B(n2992), .Z(\u_a23_mem/n18890 ) );
  OR U3896 ( .A(n1025), .B(n2983), .Z(n2992) );
  AND U3897 ( .A(n2993), .B(n2994), .Z(n2991) );
  NANDN U3898 ( .B(n1142), .A(n2939), .Z(n2994) );
  NAND U3899 ( .A(n2986), .B(\u_a23_mem/p_mem[66][2] ), .Z(n2993) );
  NAND U3900 ( .A(n2995), .B(n2996), .Z(\u_a23_mem/n18889 ) );
  OR U3901 ( .A(n1031), .B(n2983), .Z(n2996) );
  AND U3902 ( .A(n2997), .B(n2998), .Z(n2995) );
  NANDN U3903 ( .B(n1147), .A(n2939), .Z(n2998) );
  NAND U3904 ( .A(n2986), .B(\u_a23_mem/p_mem[66][3] ), .Z(n2997) );
  NAND U3905 ( .A(n2999), .B(n3000), .Z(\u_a23_mem/n18888 ) );
  OR U3906 ( .A(n1037), .B(n2983), .Z(n3000) );
  AND U3907 ( .A(n3001), .B(n3002), .Z(n2999) );
  NANDN U3908 ( .B(n1152), .A(n2939), .Z(n3002) );
  NAND U3909 ( .A(n2986), .B(\u_a23_mem/p_mem[66][4] ), .Z(n3001) );
  NAND U3910 ( .A(n3003), .B(n3004), .Z(\u_a23_mem/n18887 ) );
  OR U3911 ( .A(n1043), .B(n2983), .Z(n3004) );
  AND U3912 ( .A(n3005), .B(n3006), .Z(n3003) );
  NANDN U3913 ( .B(n1157), .A(n2939), .Z(n3006) );
  NAND U3914 ( .A(n2986), .B(\u_a23_mem/p_mem[66][5] ), .Z(n3005) );
  NAND U3915 ( .A(n3007), .B(n3008), .Z(\u_a23_mem/n18886 ) );
  OR U3916 ( .A(n1049), .B(n2983), .Z(n3008) );
  AND U3917 ( .A(n3009), .B(n3010), .Z(n3007) );
  NANDN U3918 ( .B(n1162), .A(n2939), .Z(n3010) );
  NAND U3919 ( .A(n2986), .B(\u_a23_mem/p_mem[66][6] ), .Z(n3009) );
  NAND U3920 ( .A(n3011), .B(n3012), .Z(\u_a23_mem/n18885 ) );
  NANDN U3921 ( .B(n2983), .A(n1055), .Z(n3012) );
  NAND U3922 ( .A(n1165), .B(n2939), .Z(n2983) );
  AND U3923 ( .A(n3013), .B(n3014), .Z(n3011) );
  NANDN U3924 ( .B(n1168), .A(n2939), .Z(n3014) );
  NAND U3925 ( .A(n2986), .B(\u_a23_mem/p_mem[66][7] ), .Z(n3013) );
  NANDN U3926 ( .B(n1169), .A(n2939), .Z(n2986) );
  NAND U3927 ( .A(n3015), .B(n3016), .Z(\u_a23_mem/n18884 ) );
  OR U3928 ( .A(n1011), .B(n3017), .Z(n3016) );
  AND U3929 ( .A(n3018), .B(n3019), .Z(n3015) );
  NAND U3930 ( .A(n3020), .B(\u_a23_mem/p_mem[67][0] ), .Z(n3019) );
  NANDN U3931 ( .B(n1015), .A(n2939), .Z(n3018) );
  NAND U3932 ( .A(n3021), .B(n3022), .Z(\u_a23_mem/n18883 ) );
  OR U3933 ( .A(n1019), .B(n3017), .Z(n3022) );
  AND U3934 ( .A(n3023), .B(n3024), .Z(n3021) );
  NAND U3935 ( .A(n3020), .B(\u_a23_mem/p_mem[67][1] ), .Z(n3024) );
  NANDN U3936 ( .B(n1022), .A(n2939), .Z(n3023) );
  NAND U3937 ( .A(n3025), .B(n3026), .Z(\u_a23_mem/n18882 ) );
  OR U3938 ( .A(n1025), .B(n3017), .Z(n3026) );
  AND U3939 ( .A(n3027), .B(n3028), .Z(n3025) );
  NAND U3940 ( .A(n3020), .B(\u_a23_mem/p_mem[67][2] ), .Z(n3028) );
  NANDN U3941 ( .B(n1028), .A(n2939), .Z(n3027) );
  NAND U3942 ( .A(n3029), .B(n3030), .Z(\u_a23_mem/n18881 ) );
  OR U3943 ( .A(n1031), .B(n3017), .Z(n3030) );
  AND U3944 ( .A(n3031), .B(n3032), .Z(n3029) );
  NAND U3945 ( .A(n3020), .B(\u_a23_mem/p_mem[67][3] ), .Z(n3032) );
  NANDN U3946 ( .B(n1034), .A(n2939), .Z(n3031) );
  NAND U3947 ( .A(n3033), .B(n3034), .Z(\u_a23_mem/n18880 ) );
  OR U3948 ( .A(n1037), .B(n3017), .Z(n3034) );
  AND U3949 ( .A(n3035), .B(n3036), .Z(n3033) );
  NAND U3950 ( .A(n3020), .B(\u_a23_mem/p_mem[67][4] ), .Z(n3036) );
  NANDN U3951 ( .B(n1040), .A(n2939), .Z(n3035) );
  NAND U3952 ( .A(n3037), .B(n3038), .Z(\u_a23_mem/n18879 ) );
  OR U3953 ( .A(n1043), .B(n3017), .Z(n3038) );
  AND U3954 ( .A(n3039), .B(n3040), .Z(n3037) );
  NAND U3955 ( .A(n3020), .B(\u_a23_mem/p_mem[67][5] ), .Z(n3040) );
  NANDN U3956 ( .B(n1046), .A(n2939), .Z(n3039) );
  NAND U3957 ( .A(n3041), .B(n3042), .Z(\u_a23_mem/n18878 ) );
  OR U3958 ( .A(n1049), .B(n3017), .Z(n3042) );
  AND U3959 ( .A(n3043), .B(n3044), .Z(n3041) );
  NAND U3960 ( .A(n3020), .B(\u_a23_mem/p_mem[67][6] ), .Z(n3044) );
  NANDN U3961 ( .B(n1052), .A(n2939), .Z(n3043) );
  NAND U3962 ( .A(n3045), .B(n3046), .Z(\u_a23_mem/n18877 ) );
  NANDN U3963 ( .B(n3017), .A(n1055), .Z(n3046) );
  NAND U3964 ( .A(n1056), .B(n2939), .Z(n3017) );
  AND U3965 ( .A(n3047), .B(n3048), .Z(n3045) );
  NAND U3966 ( .A(n3020), .B(\u_a23_mem/p_mem[67][7] ), .Z(n3048) );
  NANDN U3967 ( .B(n1059), .A(n2939), .Z(n3020) );
  NAND U3968 ( .A(n1061), .B(n2939), .Z(n3047) );
  ANDN U3969 ( .A(n1571), .B(n3049), .Z(n2939) );
  NAND U3970 ( .A(n3050), .B(n3051), .Z(\u_a23_mem/n18876 ) );
  NAND U3971 ( .A(n3052), .B(\u_a23_mem/p_mem[68][0] ), .Z(n3051) );
  OR U3972 ( .A(n1011), .B(n3053), .Z(n3050) );
  NAND U3973 ( .A(n3054), .B(n3055), .Z(\u_a23_mem/n18875 ) );
  NAND U3974 ( .A(n3052), .B(\u_a23_mem/p_mem[68][1] ), .Z(n3055) );
  OR U3975 ( .A(n1019), .B(n3053), .Z(n3054) );
  NAND U3976 ( .A(n3056), .B(n3057), .Z(\u_a23_mem/n18874 ) );
  NAND U3977 ( .A(n3052), .B(\u_a23_mem/p_mem[68][2] ), .Z(n3057) );
  OR U3978 ( .A(n1025), .B(n3053), .Z(n3056) );
  NAND U3979 ( .A(n3058), .B(n3059), .Z(\u_a23_mem/n18873 ) );
  NAND U3980 ( .A(n3052), .B(\u_a23_mem/p_mem[68][3] ), .Z(n3059) );
  OR U3981 ( .A(n1031), .B(n3053), .Z(n3058) );
  NAND U3982 ( .A(n3060), .B(n3061), .Z(\u_a23_mem/n18872 ) );
  NAND U3983 ( .A(n3052), .B(\u_a23_mem/p_mem[68][4] ), .Z(n3061) );
  OR U3984 ( .A(n1037), .B(n3053), .Z(n3060) );
  NAND U3985 ( .A(n3062), .B(n3063), .Z(\u_a23_mem/n18871 ) );
  NAND U3986 ( .A(n3052), .B(\u_a23_mem/p_mem[68][5] ), .Z(n3063) );
  OR U3987 ( .A(n1043), .B(n3053), .Z(n3062) );
  NAND U3988 ( .A(n3064), .B(n3065), .Z(\u_a23_mem/n18870 ) );
  NAND U3989 ( .A(n3052), .B(\u_a23_mem/p_mem[68][6] ), .Z(n3065) );
  OR U3990 ( .A(n1049), .B(n3053), .Z(n3064) );
  NAND U3991 ( .A(n3066), .B(n3067), .Z(\u_a23_mem/n18869 ) );
  NAND U3992 ( .A(n3052), .B(\u_a23_mem/p_mem[68][7] ), .Z(n3067) );
  NANDN U3993 ( .B(n1080), .A(n3068), .Z(n3052) );
  NANDN U3994 ( .B(n3053), .A(n1055), .Z(n3066) );
  NANDN U3995 ( .B(n2), .A(n3068), .Z(n3053) );
  NAND U3996 ( .A(n3069), .B(n3070), .Z(\u_a23_mem/n18868 ) );
  OR U3997 ( .A(n1011), .B(n3071), .Z(n3070) );
  AND U3998 ( .A(n3072), .B(n3073), .Z(n3069) );
  NANDN U3999 ( .B(n1087), .A(n3068), .Z(n3073) );
  NAND U4000 ( .A(n3074), .B(\u_a23_mem/p_mem[69][0] ), .Z(n3072) );
  NAND U4001 ( .A(n3075), .B(n3076), .Z(\u_a23_mem/n18867 ) );
  OR U4002 ( .A(n1019), .B(n3071), .Z(n3076) );
  AND U4003 ( .A(n3077), .B(n3078), .Z(n3075) );
  NANDN U4004 ( .B(n1093), .A(n3068), .Z(n3078) );
  NAND U4005 ( .A(n3074), .B(\u_a23_mem/p_mem[69][1] ), .Z(n3077) );
  NAND U4006 ( .A(n3079), .B(n3080), .Z(\u_a23_mem/n18866 ) );
  OR U4007 ( .A(n1025), .B(n3071), .Z(n3080) );
  AND U4008 ( .A(n3081), .B(n3082), .Z(n3079) );
  NANDN U4009 ( .B(n1098), .A(n3068), .Z(n3082) );
  NAND U4010 ( .A(n3074), .B(\u_a23_mem/p_mem[69][2] ), .Z(n3081) );
  NAND U4011 ( .A(n3083), .B(n3084), .Z(\u_a23_mem/n18865 ) );
  OR U4012 ( .A(n1031), .B(n3071), .Z(n3084) );
  AND U4013 ( .A(n3085), .B(n3086), .Z(n3083) );
  NANDN U4014 ( .B(n1103), .A(n3068), .Z(n3086) );
  NAND U4015 ( .A(n3074), .B(\u_a23_mem/p_mem[69][3] ), .Z(n3085) );
  NAND U4016 ( .A(n3087), .B(n3088), .Z(\u_a23_mem/n18864 ) );
  OR U4017 ( .A(n1037), .B(n3071), .Z(n3088) );
  AND U4018 ( .A(n3089), .B(n3090), .Z(n3087) );
  NANDN U4019 ( .B(n1108), .A(n3068), .Z(n3090) );
  NAND U4020 ( .A(n3074), .B(\u_a23_mem/p_mem[69][4] ), .Z(n3089) );
  NAND U4021 ( .A(n3091), .B(n3092), .Z(\u_a23_mem/n18863 ) );
  OR U4022 ( .A(n1043), .B(n3071), .Z(n3092) );
  AND U4023 ( .A(n3093), .B(n3094), .Z(n3091) );
  NANDN U4024 ( .B(n1113), .A(n3068), .Z(n3094) );
  NAND U4025 ( .A(n3074), .B(\u_a23_mem/p_mem[69][5] ), .Z(n3093) );
  NAND U4026 ( .A(n3095), .B(n3096), .Z(\u_a23_mem/n18862 ) );
  OR U4027 ( .A(n1049), .B(n3071), .Z(n3096) );
  AND U4028 ( .A(n3097), .B(n3098), .Z(n3095) );
  NANDN U4029 ( .B(n1118), .A(n3068), .Z(n3098) );
  NAND U4030 ( .A(n3074), .B(\u_a23_mem/p_mem[69][6] ), .Z(n3097) );
  NAND U4031 ( .A(n3099), .B(n3100), .Z(\u_a23_mem/n18861 ) );
  NANDN U4032 ( .B(n3071), .A(n1055), .Z(n3100) );
  NAND U4033 ( .A(n1121), .B(n3068), .Z(n3071) );
  AND U4034 ( .A(n3101), .B(n3102), .Z(n3099) );
  NANDN U4035 ( .B(n1124), .A(n3068), .Z(n3102) );
  NAND U4036 ( .A(n3074), .B(\u_a23_mem/p_mem[69][7] ), .Z(n3101) );
  NANDN U4037 ( .B(n1125), .A(n3068), .Z(n3074) );
  NAND U4038 ( .A(n3103), .B(n3104), .Z(\u_a23_mem/n18860 ) );
  OR U4039 ( .A(n1011), .B(n3105), .Z(n3104) );
  AND U4040 ( .A(n3106), .B(n3107), .Z(n3103) );
  NANDN U4041 ( .B(n1131), .A(n3068), .Z(n3107) );
  NAND U4042 ( .A(n3108), .B(\u_a23_mem/p_mem[70][0] ), .Z(n3106) );
  NAND U4043 ( .A(n3109), .B(n3110), .Z(\u_a23_mem/n18859 ) );
  OR U4044 ( .A(n1019), .B(n3105), .Z(n3110) );
  AND U4045 ( .A(n3111), .B(n3112), .Z(n3109) );
  NANDN U4046 ( .B(n1137), .A(n3068), .Z(n3112) );
  NAND U4047 ( .A(n3108), .B(\u_a23_mem/p_mem[70][1] ), .Z(n3111) );
  NAND U4048 ( .A(n3113), .B(n3114), .Z(\u_a23_mem/n18858 ) );
  OR U4049 ( .A(n1025), .B(n3105), .Z(n3114) );
  AND U4050 ( .A(n3115), .B(n3116), .Z(n3113) );
  NANDN U4051 ( .B(n1142), .A(n3068), .Z(n3116) );
  NAND U4052 ( .A(n3108), .B(\u_a23_mem/p_mem[70][2] ), .Z(n3115) );
  NAND U4053 ( .A(n3117), .B(n3118), .Z(\u_a23_mem/n18857 ) );
  OR U4054 ( .A(n1031), .B(n3105), .Z(n3118) );
  AND U4055 ( .A(n3119), .B(n3120), .Z(n3117) );
  NANDN U4056 ( .B(n1147), .A(n3068), .Z(n3120) );
  NAND U4057 ( .A(n3108), .B(\u_a23_mem/p_mem[70][3] ), .Z(n3119) );
  NAND U4058 ( .A(n3121), .B(n3122), .Z(\u_a23_mem/n18856 ) );
  OR U4059 ( .A(n1037), .B(n3105), .Z(n3122) );
  AND U4060 ( .A(n3123), .B(n3124), .Z(n3121) );
  NANDN U4061 ( .B(n1152), .A(n3068), .Z(n3124) );
  NAND U4062 ( .A(n3108), .B(\u_a23_mem/p_mem[70][4] ), .Z(n3123) );
  NAND U4063 ( .A(n3125), .B(n3126), .Z(\u_a23_mem/n18855 ) );
  OR U4064 ( .A(n1043), .B(n3105), .Z(n3126) );
  AND U4065 ( .A(n3127), .B(n3128), .Z(n3125) );
  NANDN U4066 ( .B(n1157), .A(n3068), .Z(n3128) );
  NAND U4067 ( .A(n3108), .B(\u_a23_mem/p_mem[70][5] ), .Z(n3127) );
  NAND U4068 ( .A(n3129), .B(n3130), .Z(\u_a23_mem/n18854 ) );
  OR U4069 ( .A(n1049), .B(n3105), .Z(n3130) );
  AND U4070 ( .A(n3131), .B(n3132), .Z(n3129) );
  NANDN U4071 ( .B(n1162), .A(n3068), .Z(n3132) );
  NAND U4072 ( .A(n3108), .B(\u_a23_mem/p_mem[70][6] ), .Z(n3131) );
  NAND U4073 ( .A(n3133), .B(n3134), .Z(\u_a23_mem/n18853 ) );
  NANDN U4074 ( .B(n3105), .A(n1055), .Z(n3134) );
  NAND U4075 ( .A(n1165), .B(n3068), .Z(n3105) );
  AND U4076 ( .A(n3135), .B(n3136), .Z(n3133) );
  NANDN U4077 ( .B(n1168), .A(n3068), .Z(n3136) );
  NAND U4078 ( .A(n3108), .B(\u_a23_mem/p_mem[70][7] ), .Z(n3135) );
  NANDN U4079 ( .B(n1169), .A(n3068), .Z(n3108) );
  NAND U4080 ( .A(n3137), .B(n3138), .Z(\u_a23_mem/n18852 ) );
  OR U4081 ( .A(n1011), .B(n3139), .Z(n3138) );
  AND U4082 ( .A(n3140), .B(n3141), .Z(n3137) );
  NAND U4083 ( .A(n3142), .B(\u_a23_mem/p_mem[71][0] ), .Z(n3141) );
  NANDN U4084 ( .B(n1015), .A(n3068), .Z(n3140) );
  NAND U4085 ( .A(n3143), .B(n3144), .Z(\u_a23_mem/n18851 ) );
  OR U4086 ( .A(n1019), .B(n3139), .Z(n3144) );
  AND U4087 ( .A(n3145), .B(n3146), .Z(n3143) );
  NAND U4088 ( .A(n3142), .B(\u_a23_mem/p_mem[71][1] ), .Z(n3146) );
  NANDN U4089 ( .B(n1022), .A(n3068), .Z(n3145) );
  NAND U4090 ( .A(n3147), .B(n3148), .Z(\u_a23_mem/n18850 ) );
  OR U4091 ( .A(n1025), .B(n3139), .Z(n3148) );
  AND U4092 ( .A(n3149), .B(n3150), .Z(n3147) );
  NAND U4093 ( .A(n3142), .B(\u_a23_mem/p_mem[71][2] ), .Z(n3150) );
  NANDN U4094 ( .B(n1028), .A(n3068), .Z(n3149) );
  NAND U4095 ( .A(n3151), .B(n3152), .Z(\u_a23_mem/n18849 ) );
  OR U4096 ( .A(n1031), .B(n3139), .Z(n3152) );
  AND U4097 ( .A(n3153), .B(n3154), .Z(n3151) );
  NAND U4098 ( .A(n3142), .B(\u_a23_mem/p_mem[71][3] ), .Z(n3154) );
  NANDN U4099 ( .B(n1034), .A(n3068), .Z(n3153) );
  NAND U4100 ( .A(n3155), .B(n3156), .Z(\u_a23_mem/n18848 ) );
  OR U4101 ( .A(n1037), .B(n3139), .Z(n3156) );
  AND U4102 ( .A(n3157), .B(n3158), .Z(n3155) );
  NAND U4103 ( .A(n3142), .B(\u_a23_mem/p_mem[71][4] ), .Z(n3158) );
  NANDN U4104 ( .B(n1040), .A(n3068), .Z(n3157) );
  NAND U4105 ( .A(n3159), .B(n3160), .Z(\u_a23_mem/n18847 ) );
  OR U4106 ( .A(n1043), .B(n3139), .Z(n3160) );
  AND U4107 ( .A(n3161), .B(n3162), .Z(n3159) );
  NAND U4108 ( .A(n3142), .B(\u_a23_mem/p_mem[71][5] ), .Z(n3162) );
  NANDN U4109 ( .B(n1046), .A(n3068), .Z(n3161) );
  NAND U4110 ( .A(n3163), .B(n3164), .Z(\u_a23_mem/n18846 ) );
  OR U4111 ( .A(n1049), .B(n3139), .Z(n3164) );
  AND U4112 ( .A(n3165), .B(n3166), .Z(n3163) );
  NAND U4113 ( .A(n3142), .B(\u_a23_mem/p_mem[71][6] ), .Z(n3166) );
  NANDN U4114 ( .B(n1052), .A(n3068), .Z(n3165) );
  NAND U4115 ( .A(n3167), .B(n3168), .Z(\u_a23_mem/n18845 ) );
  NANDN U4116 ( .B(n3139), .A(n1055), .Z(n3168) );
  NAND U4117 ( .A(n1056), .B(n3068), .Z(n3139) );
  AND U4118 ( .A(n3169), .B(n3170), .Z(n3167) );
  NAND U4119 ( .A(n3142), .B(\u_a23_mem/p_mem[71][7] ), .Z(n3170) );
  NANDN U4120 ( .B(n1059), .A(n3068), .Z(n3142) );
  NAND U4121 ( .A(n1061), .B(n3068), .Z(n3169) );
  AND U4122 ( .A(n1694), .B(n3171), .Z(n3068) );
  NAND U4123 ( .A(n3172), .B(n3173), .Z(\u_a23_mem/n18844 ) );
  NAND U4124 ( .A(n3174), .B(\u_a23_mem/p_mem[72][0] ), .Z(n3173) );
  OR U4125 ( .A(n1011), .B(n3175), .Z(n3172) );
  NAND U4126 ( .A(n3176), .B(n3177), .Z(\u_a23_mem/n18843 ) );
  NAND U4127 ( .A(n3174), .B(\u_a23_mem/p_mem[72][1] ), .Z(n3177) );
  OR U4128 ( .A(n1019), .B(n3175), .Z(n3176) );
  NAND U4129 ( .A(n3178), .B(n3179), .Z(\u_a23_mem/n18842 ) );
  NAND U4130 ( .A(n3174), .B(\u_a23_mem/p_mem[72][2] ), .Z(n3179) );
  OR U4131 ( .A(n1025), .B(n3175), .Z(n3178) );
  NAND U4132 ( .A(n3180), .B(n3181), .Z(\u_a23_mem/n18841 ) );
  NAND U4133 ( .A(n3174), .B(\u_a23_mem/p_mem[72][3] ), .Z(n3181) );
  OR U4134 ( .A(n1031), .B(n3175), .Z(n3180) );
  NAND U4135 ( .A(n3182), .B(n3183), .Z(\u_a23_mem/n18840 ) );
  NAND U4136 ( .A(n3174), .B(\u_a23_mem/p_mem[72][4] ), .Z(n3183) );
  OR U4137 ( .A(n1037), .B(n3175), .Z(n3182) );
  NAND U4138 ( .A(n3184), .B(n3185), .Z(\u_a23_mem/n18839 ) );
  NAND U4139 ( .A(n3174), .B(\u_a23_mem/p_mem[72][5] ), .Z(n3185) );
  OR U4140 ( .A(n1043), .B(n3175), .Z(n3184) );
  NAND U4141 ( .A(n3186), .B(n3187), .Z(\u_a23_mem/n18838 ) );
  NAND U4142 ( .A(n3174), .B(\u_a23_mem/p_mem[72][6] ), .Z(n3187) );
  OR U4143 ( .A(n1049), .B(n3175), .Z(n3186) );
  NAND U4144 ( .A(n3188), .B(n3189), .Z(\u_a23_mem/n18837 ) );
  NAND U4145 ( .A(n3174), .B(\u_a23_mem/p_mem[72][7] ), .Z(n3189) );
  NANDN U4146 ( .B(n1080), .A(n3190), .Z(n3174) );
  NANDN U4147 ( .B(n3175), .A(n1055), .Z(n3188) );
  NANDN U4148 ( .B(n2), .A(n3190), .Z(n3175) );
  NAND U4149 ( .A(n3191), .B(n3192), .Z(\u_a23_mem/n18836 ) );
  OR U4150 ( .A(n1011), .B(n3193), .Z(n3192) );
  AND U4151 ( .A(n3194), .B(n3195), .Z(n3191) );
  NANDN U4152 ( .B(n1087), .A(n3190), .Z(n3195) );
  NAND U4153 ( .A(n3196), .B(\u_a23_mem/p_mem[73][0] ), .Z(n3194) );
  NAND U4154 ( .A(n3197), .B(n3198), .Z(\u_a23_mem/n18835 ) );
  OR U4155 ( .A(n1019), .B(n3193), .Z(n3198) );
  AND U4156 ( .A(n3199), .B(n3200), .Z(n3197) );
  NANDN U4157 ( .B(n1093), .A(n3190), .Z(n3200) );
  NAND U4158 ( .A(n3196), .B(\u_a23_mem/p_mem[73][1] ), .Z(n3199) );
  NAND U4159 ( .A(n3201), .B(n3202), .Z(\u_a23_mem/n18834 ) );
  OR U4160 ( .A(n1025), .B(n3193), .Z(n3202) );
  AND U4161 ( .A(n3203), .B(n3204), .Z(n3201) );
  NANDN U4162 ( .B(n1098), .A(n3190), .Z(n3204) );
  NAND U4163 ( .A(n3196), .B(\u_a23_mem/p_mem[73][2] ), .Z(n3203) );
  NAND U4164 ( .A(n3205), .B(n3206), .Z(\u_a23_mem/n18833 ) );
  OR U4165 ( .A(n1031), .B(n3193), .Z(n3206) );
  AND U4166 ( .A(n3207), .B(n3208), .Z(n3205) );
  NANDN U4167 ( .B(n1103), .A(n3190), .Z(n3208) );
  NAND U4168 ( .A(n3196), .B(\u_a23_mem/p_mem[73][3] ), .Z(n3207) );
  NAND U4169 ( .A(n3209), .B(n3210), .Z(\u_a23_mem/n18832 ) );
  OR U4170 ( .A(n1037), .B(n3193), .Z(n3210) );
  AND U4171 ( .A(n3211), .B(n3212), .Z(n3209) );
  NANDN U4172 ( .B(n1108), .A(n3190), .Z(n3212) );
  NAND U4173 ( .A(n3196), .B(\u_a23_mem/p_mem[73][4] ), .Z(n3211) );
  NAND U4174 ( .A(n3213), .B(n3214), .Z(\u_a23_mem/n18831 ) );
  OR U4175 ( .A(n1043), .B(n3193), .Z(n3214) );
  AND U4176 ( .A(n3215), .B(n3216), .Z(n3213) );
  NANDN U4177 ( .B(n1113), .A(n3190), .Z(n3216) );
  NAND U4178 ( .A(n3196), .B(\u_a23_mem/p_mem[73][5] ), .Z(n3215) );
  NAND U4179 ( .A(n3217), .B(n3218), .Z(\u_a23_mem/n18830 ) );
  OR U4180 ( .A(n1049), .B(n3193), .Z(n3218) );
  AND U4181 ( .A(n3219), .B(n3220), .Z(n3217) );
  NANDN U4182 ( .B(n1118), .A(n3190), .Z(n3220) );
  NAND U4183 ( .A(n3196), .B(\u_a23_mem/p_mem[73][6] ), .Z(n3219) );
  NAND U4184 ( .A(n3221), .B(n3222), .Z(\u_a23_mem/n18829 ) );
  NANDN U4185 ( .B(n3193), .A(n1055), .Z(n3222) );
  NAND U4186 ( .A(n1121), .B(n3190), .Z(n3193) );
  AND U4187 ( .A(n3223), .B(n3224), .Z(n3221) );
  NANDN U4188 ( .B(n1124), .A(n3190), .Z(n3224) );
  NAND U4189 ( .A(n3196), .B(\u_a23_mem/p_mem[73][7] ), .Z(n3223) );
  NANDN U4190 ( .B(n1125), .A(n3190), .Z(n3196) );
  NAND U4191 ( .A(n3225), .B(n3226), .Z(\u_a23_mem/n18828 ) );
  OR U4192 ( .A(n1011), .B(n3227), .Z(n3226) );
  AND U4193 ( .A(n3228), .B(n3229), .Z(n3225) );
  NANDN U4194 ( .B(n1131), .A(n3190), .Z(n3229) );
  NAND U4195 ( .A(n3230), .B(\u_a23_mem/p_mem[74][0] ), .Z(n3228) );
  NAND U4196 ( .A(n3231), .B(n3232), .Z(\u_a23_mem/n18827 ) );
  OR U4197 ( .A(n1019), .B(n3227), .Z(n3232) );
  AND U4198 ( .A(n3233), .B(n3234), .Z(n3231) );
  NANDN U4199 ( .B(n1137), .A(n3190), .Z(n3234) );
  NAND U4200 ( .A(n3230), .B(\u_a23_mem/p_mem[74][1] ), .Z(n3233) );
  NAND U4201 ( .A(n3235), .B(n3236), .Z(\u_a23_mem/n18826 ) );
  OR U4202 ( .A(n1025), .B(n3227), .Z(n3236) );
  AND U4203 ( .A(n3237), .B(n3238), .Z(n3235) );
  NANDN U4204 ( .B(n1142), .A(n3190), .Z(n3238) );
  NAND U4205 ( .A(n3230), .B(\u_a23_mem/p_mem[74][2] ), .Z(n3237) );
  NAND U4206 ( .A(n3239), .B(n3240), .Z(\u_a23_mem/n18825 ) );
  OR U4207 ( .A(n1031), .B(n3227), .Z(n3240) );
  AND U4208 ( .A(n3241), .B(n3242), .Z(n3239) );
  NANDN U4209 ( .B(n1147), .A(n3190), .Z(n3242) );
  NAND U4210 ( .A(n3230), .B(\u_a23_mem/p_mem[74][3] ), .Z(n3241) );
  NAND U4211 ( .A(n3243), .B(n3244), .Z(\u_a23_mem/n18824 ) );
  OR U4212 ( .A(n1037), .B(n3227), .Z(n3244) );
  AND U4213 ( .A(n3245), .B(n3246), .Z(n3243) );
  NANDN U4214 ( .B(n1152), .A(n3190), .Z(n3246) );
  NAND U4215 ( .A(n3230), .B(\u_a23_mem/p_mem[74][4] ), .Z(n3245) );
  NAND U4216 ( .A(n3247), .B(n3248), .Z(\u_a23_mem/n18823 ) );
  OR U4217 ( .A(n1043), .B(n3227), .Z(n3248) );
  AND U4218 ( .A(n3249), .B(n3250), .Z(n3247) );
  NANDN U4219 ( .B(n1157), .A(n3190), .Z(n3250) );
  NAND U4220 ( .A(n3230), .B(\u_a23_mem/p_mem[74][5] ), .Z(n3249) );
  NAND U4221 ( .A(n3251), .B(n3252), .Z(\u_a23_mem/n18822 ) );
  OR U4222 ( .A(n1049), .B(n3227), .Z(n3252) );
  AND U4223 ( .A(n3253), .B(n3254), .Z(n3251) );
  NANDN U4224 ( .B(n1162), .A(n3190), .Z(n3254) );
  NAND U4225 ( .A(n3230), .B(\u_a23_mem/p_mem[74][6] ), .Z(n3253) );
  NAND U4226 ( .A(n3255), .B(n3256), .Z(\u_a23_mem/n18821 ) );
  NANDN U4227 ( .B(n3227), .A(n1055), .Z(n3256) );
  NAND U4228 ( .A(n1165), .B(n3190), .Z(n3227) );
  AND U4229 ( .A(n3257), .B(n3258), .Z(n3255) );
  NANDN U4230 ( .B(n1168), .A(n3190), .Z(n3258) );
  NAND U4231 ( .A(n3230), .B(\u_a23_mem/p_mem[74][7] ), .Z(n3257) );
  NANDN U4232 ( .B(n1169), .A(n3190), .Z(n3230) );
  NAND U4233 ( .A(n3259), .B(n3260), .Z(\u_a23_mem/n18820 ) );
  OR U4234 ( .A(n1011), .B(n3261), .Z(n3260) );
  AND U4235 ( .A(n3262), .B(n3263), .Z(n3259) );
  NAND U4236 ( .A(n3264), .B(\u_a23_mem/p_mem[75][0] ), .Z(n3263) );
  NANDN U4237 ( .B(n1015), .A(n3190), .Z(n3262) );
  NAND U4238 ( .A(n3265), .B(n3266), .Z(\u_a23_mem/n18819 ) );
  OR U4239 ( .A(n1019), .B(n3261), .Z(n3266) );
  AND U4240 ( .A(n3267), .B(n3268), .Z(n3265) );
  NAND U4241 ( .A(n3264), .B(\u_a23_mem/p_mem[75][1] ), .Z(n3268) );
  NANDN U4242 ( .B(n1022), .A(n3190), .Z(n3267) );
  NAND U4243 ( .A(n3269), .B(n3270), .Z(\u_a23_mem/n18818 ) );
  OR U4244 ( .A(n1025), .B(n3261), .Z(n3270) );
  AND U4245 ( .A(n3271), .B(n3272), .Z(n3269) );
  NAND U4246 ( .A(n3264), .B(\u_a23_mem/p_mem[75][2] ), .Z(n3272) );
  NANDN U4247 ( .B(n1028), .A(n3190), .Z(n3271) );
  NAND U4248 ( .A(n3273), .B(n3274), .Z(\u_a23_mem/n18817 ) );
  OR U4249 ( .A(n1031), .B(n3261), .Z(n3274) );
  AND U4250 ( .A(n3275), .B(n3276), .Z(n3273) );
  NAND U4251 ( .A(n3264), .B(\u_a23_mem/p_mem[75][3] ), .Z(n3276) );
  NANDN U4252 ( .B(n1034), .A(n3190), .Z(n3275) );
  NAND U4253 ( .A(n3277), .B(n3278), .Z(\u_a23_mem/n18816 ) );
  OR U4254 ( .A(n1037), .B(n3261), .Z(n3278) );
  AND U4255 ( .A(n3279), .B(n3280), .Z(n3277) );
  NAND U4256 ( .A(n3264), .B(\u_a23_mem/p_mem[75][4] ), .Z(n3280) );
  NANDN U4257 ( .B(n1040), .A(n3190), .Z(n3279) );
  NAND U4258 ( .A(n3281), .B(n3282), .Z(\u_a23_mem/n18815 ) );
  OR U4259 ( .A(n1043), .B(n3261), .Z(n3282) );
  AND U4260 ( .A(n3283), .B(n3284), .Z(n3281) );
  NAND U4261 ( .A(n3264), .B(\u_a23_mem/p_mem[75][5] ), .Z(n3284) );
  NANDN U4262 ( .B(n1046), .A(n3190), .Z(n3283) );
  NAND U4263 ( .A(n3285), .B(n3286), .Z(\u_a23_mem/n18814 ) );
  OR U4264 ( .A(n1049), .B(n3261), .Z(n3286) );
  AND U4265 ( .A(n3287), .B(n3288), .Z(n3285) );
  NAND U4266 ( .A(n3264), .B(\u_a23_mem/p_mem[75][6] ), .Z(n3288) );
  NANDN U4267 ( .B(n1052), .A(n3190), .Z(n3287) );
  NAND U4268 ( .A(n3289), .B(n3290), .Z(\u_a23_mem/n18813 ) );
  NANDN U4269 ( .B(n3261), .A(n1055), .Z(n3290) );
  NAND U4270 ( .A(n1056), .B(n3190), .Z(n3261) );
  AND U4271 ( .A(n3291), .B(n3292), .Z(n3289) );
  NAND U4272 ( .A(n3264), .B(\u_a23_mem/p_mem[75][7] ), .Z(n3292) );
  NANDN U4273 ( .B(n1059), .A(n3190), .Z(n3264) );
  NAND U4274 ( .A(n1061), .B(n3190), .Z(n3291) );
  AND U4275 ( .A(n1816), .B(n3171), .Z(n3190) );
  NAND U4276 ( .A(n3293), .B(n3294), .Z(\u_a23_mem/n18812 ) );
  NAND U4277 ( .A(n3295), .B(\u_a23_mem/p_mem[76][0] ), .Z(n3294) );
  OR U4278 ( .A(n1011), .B(n3296), .Z(n3293) );
  NAND U4279 ( .A(n3297), .B(n3298), .Z(\u_a23_mem/n18811 ) );
  NAND U4280 ( .A(n3295), .B(\u_a23_mem/p_mem[76][1] ), .Z(n3298) );
  OR U4281 ( .A(n1019), .B(n3296), .Z(n3297) );
  NAND U4282 ( .A(n3299), .B(n3300), .Z(\u_a23_mem/n18810 ) );
  NAND U4283 ( .A(n3295), .B(\u_a23_mem/p_mem[76][2] ), .Z(n3300) );
  OR U4284 ( .A(n1025), .B(n3296), .Z(n3299) );
  NAND U4285 ( .A(n3301), .B(n3302), .Z(\u_a23_mem/n18809 ) );
  NAND U4286 ( .A(n3295), .B(\u_a23_mem/p_mem[76][3] ), .Z(n3302) );
  OR U4287 ( .A(n1031), .B(n3296), .Z(n3301) );
  NAND U4288 ( .A(n3303), .B(n3304), .Z(\u_a23_mem/n18808 ) );
  NAND U4289 ( .A(n3295), .B(\u_a23_mem/p_mem[76][4] ), .Z(n3304) );
  OR U4290 ( .A(n1037), .B(n3296), .Z(n3303) );
  NAND U4291 ( .A(n3305), .B(n3306), .Z(\u_a23_mem/n18807 ) );
  NAND U4292 ( .A(n3295), .B(\u_a23_mem/p_mem[76][5] ), .Z(n3306) );
  OR U4293 ( .A(n1043), .B(n3296), .Z(n3305) );
  NAND U4294 ( .A(n3307), .B(n3308), .Z(\u_a23_mem/n18806 ) );
  NAND U4295 ( .A(n3295), .B(\u_a23_mem/p_mem[76][6] ), .Z(n3308) );
  OR U4296 ( .A(n1049), .B(n3296), .Z(n3307) );
  NAND U4297 ( .A(n3309), .B(n3310), .Z(\u_a23_mem/n18805 ) );
  NAND U4298 ( .A(n3295), .B(\u_a23_mem/p_mem[76][7] ), .Z(n3310) );
  NANDN U4299 ( .B(n1080), .A(n3311), .Z(n3295) );
  NANDN U4300 ( .B(n3296), .A(n1055), .Z(n3309) );
  NANDN U4301 ( .B(n2), .A(n3311), .Z(n3296) );
  NAND U4302 ( .A(n3312), .B(n3313), .Z(\u_a23_mem/n18804 ) );
  OR U4303 ( .A(n1011), .B(n3314), .Z(n3313) );
  AND U4304 ( .A(n3315), .B(n3316), .Z(n3312) );
  NANDN U4305 ( .B(n1087), .A(n3311), .Z(n3316) );
  NAND U4306 ( .A(n3317), .B(\u_a23_mem/p_mem[77][0] ), .Z(n3315) );
  NAND U4307 ( .A(n3318), .B(n3319), .Z(\u_a23_mem/n18803 ) );
  OR U4308 ( .A(n1019), .B(n3314), .Z(n3319) );
  AND U4309 ( .A(n3320), .B(n3321), .Z(n3318) );
  NANDN U4310 ( .B(n1093), .A(n3311), .Z(n3321) );
  NAND U4311 ( .A(n3317), .B(\u_a23_mem/p_mem[77][1] ), .Z(n3320) );
  NAND U4312 ( .A(n3322), .B(n3323), .Z(\u_a23_mem/n18802 ) );
  OR U4313 ( .A(n1025), .B(n3314), .Z(n3323) );
  AND U4314 ( .A(n3324), .B(n3325), .Z(n3322) );
  NANDN U4315 ( .B(n1098), .A(n3311), .Z(n3325) );
  NAND U4316 ( .A(n3317), .B(\u_a23_mem/p_mem[77][2] ), .Z(n3324) );
  NAND U4317 ( .A(n3326), .B(n3327), .Z(\u_a23_mem/n18801 ) );
  OR U4318 ( .A(n1031), .B(n3314), .Z(n3327) );
  AND U4319 ( .A(n3328), .B(n3329), .Z(n3326) );
  NANDN U4320 ( .B(n1103), .A(n3311), .Z(n3329) );
  NAND U4321 ( .A(n3317), .B(\u_a23_mem/p_mem[77][3] ), .Z(n3328) );
  NAND U4322 ( .A(n3330), .B(n3331), .Z(\u_a23_mem/n18800 ) );
  OR U4323 ( .A(n1037), .B(n3314), .Z(n3331) );
  AND U4324 ( .A(n3332), .B(n3333), .Z(n3330) );
  NANDN U4325 ( .B(n1108), .A(n3311), .Z(n3333) );
  NAND U4326 ( .A(n3317), .B(\u_a23_mem/p_mem[77][4] ), .Z(n3332) );
  NAND U4327 ( .A(n3334), .B(n3335), .Z(\u_a23_mem/n18799 ) );
  OR U4328 ( .A(n1043), .B(n3314), .Z(n3335) );
  AND U4329 ( .A(n3336), .B(n3337), .Z(n3334) );
  NANDN U4330 ( .B(n1113), .A(n3311), .Z(n3337) );
  NAND U4331 ( .A(n3317), .B(\u_a23_mem/p_mem[77][5] ), .Z(n3336) );
  NAND U4332 ( .A(n3338), .B(n3339), .Z(\u_a23_mem/n18798 ) );
  OR U4333 ( .A(n1049), .B(n3314), .Z(n3339) );
  AND U4334 ( .A(n3340), .B(n3341), .Z(n3338) );
  NANDN U4335 ( .B(n1118), .A(n3311), .Z(n3341) );
  NAND U4336 ( .A(n3317), .B(\u_a23_mem/p_mem[77][6] ), .Z(n3340) );
  NAND U4337 ( .A(n3342), .B(n3343), .Z(\u_a23_mem/n18797 ) );
  NANDN U4338 ( .B(n3314), .A(n1055), .Z(n3343) );
  NAND U4339 ( .A(n1121), .B(n3311), .Z(n3314) );
  AND U4340 ( .A(n3344), .B(n3345), .Z(n3342) );
  NANDN U4341 ( .B(n1124), .A(n3311), .Z(n3345) );
  NAND U4342 ( .A(n3317), .B(\u_a23_mem/p_mem[77][7] ), .Z(n3344) );
  NANDN U4343 ( .B(n1125), .A(n3311), .Z(n3317) );
  NAND U4344 ( .A(n3346), .B(n3347), .Z(\u_a23_mem/n18796 ) );
  OR U4345 ( .A(n1011), .B(n3348), .Z(n3347) );
  AND U4346 ( .A(n3349), .B(n3350), .Z(n3346) );
  NANDN U4347 ( .B(n1131), .A(n3311), .Z(n3350) );
  NAND U4348 ( .A(n3351), .B(\u_a23_mem/p_mem[78][0] ), .Z(n3349) );
  NAND U4349 ( .A(n3352), .B(n3353), .Z(\u_a23_mem/n18795 ) );
  OR U4350 ( .A(n1019), .B(n3348), .Z(n3353) );
  AND U4351 ( .A(n3354), .B(n3355), .Z(n3352) );
  NANDN U4352 ( .B(n1137), .A(n3311), .Z(n3355) );
  NAND U4353 ( .A(n3351), .B(\u_a23_mem/p_mem[78][1] ), .Z(n3354) );
  NAND U4354 ( .A(n3356), .B(n3357), .Z(\u_a23_mem/n18794 ) );
  OR U4355 ( .A(n1025), .B(n3348), .Z(n3357) );
  AND U4356 ( .A(n3358), .B(n3359), .Z(n3356) );
  NANDN U4357 ( .B(n1142), .A(n3311), .Z(n3359) );
  NAND U4358 ( .A(n3351), .B(\u_a23_mem/p_mem[78][2] ), .Z(n3358) );
  NAND U4359 ( .A(n3360), .B(n3361), .Z(\u_a23_mem/n18793 ) );
  OR U4360 ( .A(n1031), .B(n3348), .Z(n3361) );
  AND U4361 ( .A(n3362), .B(n3363), .Z(n3360) );
  NANDN U4362 ( .B(n1147), .A(n3311), .Z(n3363) );
  NAND U4363 ( .A(n3351), .B(\u_a23_mem/p_mem[78][3] ), .Z(n3362) );
  NAND U4364 ( .A(n3364), .B(n3365), .Z(\u_a23_mem/n18792 ) );
  OR U4365 ( .A(n1037), .B(n3348), .Z(n3365) );
  AND U4366 ( .A(n3366), .B(n3367), .Z(n3364) );
  NANDN U4367 ( .B(n1152), .A(n3311), .Z(n3367) );
  NAND U4368 ( .A(n3351), .B(\u_a23_mem/p_mem[78][4] ), .Z(n3366) );
  NAND U4369 ( .A(n3368), .B(n3369), .Z(\u_a23_mem/n18791 ) );
  OR U4370 ( .A(n1043), .B(n3348), .Z(n3369) );
  AND U4371 ( .A(n3370), .B(n3371), .Z(n3368) );
  NANDN U4372 ( .B(n1157), .A(n3311), .Z(n3371) );
  NAND U4373 ( .A(n3351), .B(\u_a23_mem/p_mem[78][5] ), .Z(n3370) );
  NAND U4374 ( .A(n3372), .B(n3373), .Z(\u_a23_mem/n18790 ) );
  OR U4375 ( .A(n1049), .B(n3348), .Z(n3373) );
  AND U4376 ( .A(n3374), .B(n3375), .Z(n3372) );
  NANDN U4377 ( .B(n1162), .A(n3311), .Z(n3375) );
  NAND U4378 ( .A(n3351), .B(\u_a23_mem/p_mem[78][6] ), .Z(n3374) );
  NAND U4379 ( .A(n3376), .B(n3377), .Z(\u_a23_mem/n18789 ) );
  NANDN U4380 ( .B(n3348), .A(n1055), .Z(n3377) );
  NAND U4381 ( .A(n1165), .B(n3311), .Z(n3348) );
  AND U4382 ( .A(n3378), .B(n3379), .Z(n3376) );
  NANDN U4383 ( .B(n1168), .A(n3311), .Z(n3379) );
  NAND U4384 ( .A(n3351), .B(\u_a23_mem/p_mem[78][7] ), .Z(n3378) );
  NANDN U4385 ( .B(n1169), .A(n3311), .Z(n3351) );
  NAND U4386 ( .A(n3380), .B(n3381), .Z(\u_a23_mem/n18788 ) );
  OR U4387 ( .A(n1011), .B(n3382), .Z(n3381) );
  AND U4388 ( .A(n3383), .B(n3384), .Z(n3380) );
  NAND U4389 ( .A(n3385), .B(\u_a23_mem/p_mem[79][0] ), .Z(n3384) );
  NANDN U4390 ( .B(n1015), .A(n3311), .Z(n3383) );
  NAND U4391 ( .A(n3386), .B(n3387), .Z(\u_a23_mem/n18787 ) );
  OR U4392 ( .A(n1019), .B(n3382), .Z(n3387) );
  AND U4393 ( .A(n3388), .B(n3389), .Z(n3386) );
  NAND U4394 ( .A(n3385), .B(\u_a23_mem/p_mem[79][1] ), .Z(n3389) );
  NANDN U4395 ( .B(n1022), .A(n3311), .Z(n3388) );
  NAND U4396 ( .A(n3390), .B(n3391), .Z(\u_a23_mem/n18786 ) );
  OR U4397 ( .A(n1025), .B(n3382), .Z(n3391) );
  AND U4398 ( .A(n3392), .B(n3393), .Z(n3390) );
  NAND U4399 ( .A(n3385), .B(\u_a23_mem/p_mem[79][2] ), .Z(n3393) );
  NANDN U4400 ( .B(n1028), .A(n3311), .Z(n3392) );
  NAND U4401 ( .A(n3394), .B(n3395), .Z(\u_a23_mem/n18785 ) );
  OR U4402 ( .A(n1031), .B(n3382), .Z(n3395) );
  AND U4403 ( .A(n3396), .B(n3397), .Z(n3394) );
  NAND U4404 ( .A(n3385), .B(\u_a23_mem/p_mem[79][3] ), .Z(n3397) );
  NANDN U4405 ( .B(n1034), .A(n3311), .Z(n3396) );
  NAND U4406 ( .A(n3398), .B(n3399), .Z(\u_a23_mem/n18784 ) );
  OR U4407 ( .A(n1037), .B(n3382), .Z(n3399) );
  AND U4408 ( .A(n3400), .B(n3401), .Z(n3398) );
  NAND U4409 ( .A(n3385), .B(\u_a23_mem/p_mem[79][4] ), .Z(n3401) );
  NANDN U4410 ( .B(n1040), .A(n3311), .Z(n3400) );
  NAND U4411 ( .A(n3402), .B(n3403), .Z(\u_a23_mem/n18783 ) );
  OR U4412 ( .A(n1043), .B(n3382), .Z(n3403) );
  AND U4413 ( .A(n3404), .B(n3405), .Z(n3402) );
  NAND U4414 ( .A(n3385), .B(\u_a23_mem/p_mem[79][5] ), .Z(n3405) );
  NANDN U4415 ( .B(n1046), .A(n3311), .Z(n3404) );
  NAND U4416 ( .A(n3406), .B(n3407), .Z(\u_a23_mem/n18782 ) );
  OR U4417 ( .A(n1049), .B(n3382), .Z(n3407) );
  AND U4418 ( .A(n3408), .B(n3409), .Z(n3406) );
  NAND U4419 ( .A(n3385), .B(\u_a23_mem/p_mem[79][6] ), .Z(n3409) );
  NANDN U4420 ( .B(n1052), .A(n3311), .Z(n3408) );
  NAND U4421 ( .A(n3410), .B(n3411), .Z(\u_a23_mem/n18781 ) );
  NANDN U4422 ( .B(n3382), .A(n1055), .Z(n3411) );
  NAND U4423 ( .A(n1056), .B(n3311), .Z(n3382) );
  AND U4424 ( .A(n3412), .B(n3413), .Z(n3410) );
  NAND U4425 ( .A(n3385), .B(\u_a23_mem/p_mem[79][7] ), .Z(n3413) );
  NANDN U4426 ( .B(n1059), .A(n3311), .Z(n3385) );
  NAND U4427 ( .A(n1061), .B(n3311), .Z(n3412) );
  NOR U4428 ( .A(n3049), .B(n1938), .Z(n3311) );
  IV U4429 ( .A(n3171), .Z(n3049) );
  ANDN U4430 ( .A(n3414), .B(n2429), .Z(n3171) );
  AND U4431 ( .A(n1939), .B(n2428), .Z(n3414) );
  NAND U4432 ( .A(n3415), .B(n3416), .Z(\u_a23_mem/n18780 ) );
  NAND U4433 ( .A(n3417), .B(\u_a23_mem/p_mem[80][0] ), .Z(n3416) );
  OR U4434 ( .A(n1011), .B(n3418), .Z(n3415) );
  NAND U4435 ( .A(n3419), .B(n3420), .Z(\u_a23_mem/n18779 ) );
  NAND U4436 ( .A(n3417), .B(\u_a23_mem/p_mem[80][1] ), .Z(n3420) );
  OR U4437 ( .A(n1019), .B(n3418), .Z(n3419) );
  NAND U4438 ( .A(n3421), .B(n3422), .Z(\u_a23_mem/n18778 ) );
  NAND U4439 ( .A(n3417), .B(\u_a23_mem/p_mem[80][2] ), .Z(n3422) );
  OR U4440 ( .A(n1025), .B(n3418), .Z(n3421) );
  NAND U4441 ( .A(n3423), .B(n3424), .Z(\u_a23_mem/n18777 ) );
  NAND U4442 ( .A(n3417), .B(\u_a23_mem/p_mem[80][3] ), .Z(n3424) );
  OR U4443 ( .A(n1031), .B(n3418), .Z(n3423) );
  NAND U4444 ( .A(n3425), .B(n3426), .Z(\u_a23_mem/n18776 ) );
  NAND U4445 ( .A(n3417), .B(\u_a23_mem/p_mem[80][4] ), .Z(n3426) );
  OR U4446 ( .A(n1037), .B(n3418), .Z(n3425) );
  NAND U4447 ( .A(n3427), .B(n3428), .Z(\u_a23_mem/n18775 ) );
  NAND U4448 ( .A(n3417), .B(\u_a23_mem/p_mem[80][5] ), .Z(n3428) );
  OR U4449 ( .A(n1043), .B(n3418), .Z(n3427) );
  NAND U4450 ( .A(n3429), .B(n3430), .Z(\u_a23_mem/n18774 ) );
  NAND U4451 ( .A(n3417), .B(\u_a23_mem/p_mem[80][6] ), .Z(n3430) );
  OR U4452 ( .A(n1049), .B(n3418), .Z(n3429) );
  NAND U4453 ( .A(n3431), .B(n3432), .Z(\u_a23_mem/n18773 ) );
  NAND U4454 ( .A(n3417), .B(\u_a23_mem/p_mem[80][7] ), .Z(n3432) );
  NANDN U4455 ( .B(n1080), .A(n3433), .Z(n3417) );
  NANDN U4456 ( .B(n3418), .A(n1055), .Z(n3431) );
  NANDN U4457 ( .B(n2), .A(n3433), .Z(n3418) );
  NAND U4458 ( .A(n3434), .B(n3435), .Z(\u_a23_mem/n18772 ) );
  OR U4459 ( .A(n1011), .B(n3436), .Z(n3435) );
  AND U4460 ( .A(n3437), .B(n3438), .Z(n3434) );
  NANDN U4461 ( .B(n1087), .A(n3433), .Z(n3438) );
  NAND U4462 ( .A(n3439), .B(\u_a23_mem/p_mem[81][0] ), .Z(n3437) );
  NAND U4463 ( .A(n3440), .B(n3441), .Z(\u_a23_mem/n18771 ) );
  OR U4464 ( .A(n1019), .B(n3436), .Z(n3441) );
  AND U4465 ( .A(n3442), .B(n3443), .Z(n3440) );
  NANDN U4466 ( .B(n1093), .A(n3433), .Z(n3443) );
  NAND U4467 ( .A(n3439), .B(\u_a23_mem/p_mem[81][1] ), .Z(n3442) );
  NAND U4468 ( .A(n3444), .B(n3445), .Z(\u_a23_mem/n18770 ) );
  OR U4469 ( .A(n1025), .B(n3436), .Z(n3445) );
  AND U4470 ( .A(n3446), .B(n3447), .Z(n3444) );
  NANDN U4471 ( .B(n1098), .A(n3433), .Z(n3447) );
  NAND U4472 ( .A(n3439), .B(\u_a23_mem/p_mem[81][2] ), .Z(n3446) );
  NAND U4473 ( .A(n3448), .B(n3449), .Z(\u_a23_mem/n18769 ) );
  OR U4474 ( .A(n1031), .B(n3436), .Z(n3449) );
  AND U4475 ( .A(n3450), .B(n3451), .Z(n3448) );
  NANDN U4476 ( .B(n1103), .A(n3433), .Z(n3451) );
  NAND U4477 ( .A(n3439), .B(\u_a23_mem/p_mem[81][3] ), .Z(n3450) );
  NAND U4478 ( .A(n3452), .B(n3453), .Z(\u_a23_mem/n18768 ) );
  OR U4479 ( .A(n1037), .B(n3436), .Z(n3453) );
  AND U4480 ( .A(n3454), .B(n3455), .Z(n3452) );
  NANDN U4481 ( .B(n1108), .A(n3433), .Z(n3455) );
  NAND U4482 ( .A(n3439), .B(\u_a23_mem/p_mem[81][4] ), .Z(n3454) );
  NAND U4483 ( .A(n3456), .B(n3457), .Z(\u_a23_mem/n18767 ) );
  OR U4484 ( .A(n1043), .B(n3436), .Z(n3457) );
  AND U4485 ( .A(n3458), .B(n3459), .Z(n3456) );
  NANDN U4486 ( .B(n1113), .A(n3433), .Z(n3459) );
  NAND U4487 ( .A(n3439), .B(\u_a23_mem/p_mem[81][5] ), .Z(n3458) );
  NAND U4488 ( .A(n3460), .B(n3461), .Z(\u_a23_mem/n18766 ) );
  OR U4489 ( .A(n1049), .B(n3436), .Z(n3461) );
  AND U4490 ( .A(n3462), .B(n3463), .Z(n3460) );
  NANDN U4491 ( .B(n1118), .A(n3433), .Z(n3463) );
  NAND U4492 ( .A(n3439), .B(\u_a23_mem/p_mem[81][6] ), .Z(n3462) );
  NAND U4493 ( .A(n3464), .B(n3465), .Z(\u_a23_mem/n18765 ) );
  NANDN U4494 ( .B(n3436), .A(n1055), .Z(n3465) );
  NAND U4495 ( .A(n1121), .B(n3433), .Z(n3436) );
  AND U4496 ( .A(n3466), .B(n3467), .Z(n3464) );
  NANDN U4497 ( .B(n1124), .A(n3433), .Z(n3467) );
  NAND U4498 ( .A(n3439), .B(\u_a23_mem/p_mem[81][7] ), .Z(n3466) );
  NANDN U4499 ( .B(n1125), .A(n3433), .Z(n3439) );
  NAND U4500 ( .A(n3468), .B(n3469), .Z(\u_a23_mem/n18764 ) );
  OR U4501 ( .A(n1011), .B(n3470), .Z(n3469) );
  AND U4502 ( .A(n3471), .B(n3472), .Z(n3468) );
  NANDN U4503 ( .B(n1131), .A(n3433), .Z(n3472) );
  NAND U4504 ( .A(n3473), .B(\u_a23_mem/p_mem[82][0] ), .Z(n3471) );
  NAND U4505 ( .A(n3474), .B(n3475), .Z(\u_a23_mem/n18763 ) );
  OR U4506 ( .A(n1019), .B(n3470), .Z(n3475) );
  AND U4507 ( .A(n3476), .B(n3477), .Z(n3474) );
  NANDN U4508 ( .B(n1137), .A(n3433), .Z(n3477) );
  NAND U4509 ( .A(n3473), .B(\u_a23_mem/p_mem[82][1] ), .Z(n3476) );
  NAND U4510 ( .A(n3478), .B(n3479), .Z(\u_a23_mem/n18762 ) );
  OR U4511 ( .A(n1025), .B(n3470), .Z(n3479) );
  AND U4512 ( .A(n3480), .B(n3481), .Z(n3478) );
  NANDN U4513 ( .B(n1142), .A(n3433), .Z(n3481) );
  NAND U4514 ( .A(n3473), .B(\u_a23_mem/p_mem[82][2] ), .Z(n3480) );
  NAND U4515 ( .A(n3482), .B(n3483), .Z(\u_a23_mem/n18761 ) );
  OR U4516 ( .A(n1031), .B(n3470), .Z(n3483) );
  AND U4517 ( .A(n3484), .B(n3485), .Z(n3482) );
  NANDN U4518 ( .B(n1147), .A(n3433), .Z(n3485) );
  NAND U4519 ( .A(n3473), .B(\u_a23_mem/p_mem[82][3] ), .Z(n3484) );
  NAND U4520 ( .A(n3486), .B(n3487), .Z(\u_a23_mem/n18760 ) );
  OR U4521 ( .A(n1037), .B(n3470), .Z(n3487) );
  AND U4522 ( .A(n3488), .B(n3489), .Z(n3486) );
  NANDN U4523 ( .B(n1152), .A(n3433), .Z(n3489) );
  NAND U4524 ( .A(n3473), .B(\u_a23_mem/p_mem[82][4] ), .Z(n3488) );
  NAND U4525 ( .A(n3490), .B(n3491), .Z(\u_a23_mem/n18759 ) );
  OR U4526 ( .A(n1043), .B(n3470), .Z(n3491) );
  AND U4527 ( .A(n3492), .B(n3493), .Z(n3490) );
  NANDN U4528 ( .B(n1157), .A(n3433), .Z(n3493) );
  NAND U4529 ( .A(n3473), .B(\u_a23_mem/p_mem[82][5] ), .Z(n3492) );
  NAND U4530 ( .A(n3494), .B(n3495), .Z(\u_a23_mem/n18758 ) );
  OR U4531 ( .A(n1049), .B(n3470), .Z(n3495) );
  AND U4532 ( .A(n3496), .B(n3497), .Z(n3494) );
  NANDN U4533 ( .B(n1162), .A(n3433), .Z(n3497) );
  NAND U4534 ( .A(n3473), .B(\u_a23_mem/p_mem[82][6] ), .Z(n3496) );
  NAND U4535 ( .A(n3498), .B(n3499), .Z(\u_a23_mem/n18757 ) );
  NANDN U4536 ( .B(n3470), .A(n1055), .Z(n3499) );
  NAND U4537 ( .A(n1165), .B(n3433), .Z(n3470) );
  AND U4538 ( .A(n3500), .B(n3501), .Z(n3498) );
  NANDN U4539 ( .B(n1168), .A(n3433), .Z(n3501) );
  NAND U4540 ( .A(n3473), .B(\u_a23_mem/p_mem[82][7] ), .Z(n3500) );
  NANDN U4541 ( .B(n1169), .A(n3433), .Z(n3473) );
  NAND U4542 ( .A(n3502), .B(n3503), .Z(\u_a23_mem/n18756 ) );
  OR U4543 ( .A(n1011), .B(n3504), .Z(n3503) );
  AND U4544 ( .A(n3505), .B(n3506), .Z(n3502) );
  NAND U4545 ( .A(n3507), .B(\u_a23_mem/p_mem[83][0] ), .Z(n3506) );
  NANDN U4546 ( .B(n1015), .A(n3433), .Z(n3505) );
  NAND U4547 ( .A(n3508), .B(n3509), .Z(\u_a23_mem/n18755 ) );
  OR U4548 ( .A(n1019), .B(n3504), .Z(n3509) );
  AND U4549 ( .A(n3510), .B(n3511), .Z(n3508) );
  NAND U4550 ( .A(n3507), .B(\u_a23_mem/p_mem[83][1] ), .Z(n3511) );
  NANDN U4551 ( .B(n1022), .A(n3433), .Z(n3510) );
  NAND U4552 ( .A(n3512), .B(n3513), .Z(\u_a23_mem/n18754 ) );
  OR U4553 ( .A(n1025), .B(n3504), .Z(n3513) );
  AND U4554 ( .A(n3514), .B(n3515), .Z(n3512) );
  NAND U4555 ( .A(n3507), .B(\u_a23_mem/p_mem[83][2] ), .Z(n3515) );
  NANDN U4556 ( .B(n1028), .A(n3433), .Z(n3514) );
  NAND U4557 ( .A(n3516), .B(n3517), .Z(\u_a23_mem/n18753 ) );
  OR U4558 ( .A(n1031), .B(n3504), .Z(n3517) );
  AND U4559 ( .A(n3518), .B(n3519), .Z(n3516) );
  NAND U4560 ( .A(n3507), .B(\u_a23_mem/p_mem[83][3] ), .Z(n3519) );
  NANDN U4561 ( .B(n1034), .A(n3433), .Z(n3518) );
  NAND U4562 ( .A(n3520), .B(n3521), .Z(\u_a23_mem/n18752 ) );
  OR U4563 ( .A(n1037), .B(n3504), .Z(n3521) );
  AND U4564 ( .A(n3522), .B(n3523), .Z(n3520) );
  NAND U4565 ( .A(n3507), .B(\u_a23_mem/p_mem[83][4] ), .Z(n3523) );
  NANDN U4566 ( .B(n1040), .A(n3433), .Z(n3522) );
  NAND U4567 ( .A(n3524), .B(n3525), .Z(\u_a23_mem/n18751 ) );
  OR U4568 ( .A(n1043), .B(n3504), .Z(n3525) );
  AND U4569 ( .A(n3526), .B(n3527), .Z(n3524) );
  NAND U4570 ( .A(n3507), .B(\u_a23_mem/p_mem[83][5] ), .Z(n3527) );
  NANDN U4571 ( .B(n1046), .A(n3433), .Z(n3526) );
  NAND U4572 ( .A(n3528), .B(n3529), .Z(\u_a23_mem/n18750 ) );
  OR U4573 ( .A(n1049), .B(n3504), .Z(n3529) );
  AND U4574 ( .A(n3530), .B(n3531), .Z(n3528) );
  NAND U4575 ( .A(n3507), .B(\u_a23_mem/p_mem[83][6] ), .Z(n3531) );
  NANDN U4576 ( .B(n1052), .A(n3433), .Z(n3530) );
  NAND U4577 ( .A(n3532), .B(n3533), .Z(\u_a23_mem/n18749 ) );
  NANDN U4578 ( .B(n3504), .A(n1055), .Z(n3533) );
  NAND U4579 ( .A(n1056), .B(n3433), .Z(n3504) );
  AND U4580 ( .A(n3534), .B(n3535), .Z(n3532) );
  NAND U4581 ( .A(n3507), .B(\u_a23_mem/p_mem[83][7] ), .Z(n3535) );
  NANDN U4582 ( .B(n1059), .A(n3433), .Z(n3507) );
  NAND U4583 ( .A(n1061), .B(n3433), .Z(n3534) );
  ANDN U4584 ( .A(n1571), .B(n3536), .Z(n3433) );
  NAND U4585 ( .A(n3537), .B(n3538), .Z(\u_a23_mem/n18748 ) );
  NAND U4586 ( .A(n3539), .B(\u_a23_mem/p_mem[84][0] ), .Z(n3538) );
  OR U4587 ( .A(n1011), .B(n3540), .Z(n3537) );
  NAND U4588 ( .A(n3541), .B(n3542), .Z(\u_a23_mem/n18747 ) );
  NAND U4589 ( .A(n3539), .B(\u_a23_mem/p_mem[84][1] ), .Z(n3542) );
  OR U4590 ( .A(n1019), .B(n3540), .Z(n3541) );
  NAND U4591 ( .A(n3543), .B(n3544), .Z(\u_a23_mem/n18746 ) );
  NAND U4592 ( .A(n3539), .B(\u_a23_mem/p_mem[84][2] ), .Z(n3544) );
  OR U4593 ( .A(n1025), .B(n3540), .Z(n3543) );
  NAND U4594 ( .A(n3545), .B(n3546), .Z(\u_a23_mem/n18745 ) );
  NAND U4595 ( .A(n3539), .B(\u_a23_mem/p_mem[84][3] ), .Z(n3546) );
  OR U4596 ( .A(n1031), .B(n3540), .Z(n3545) );
  NAND U4597 ( .A(n3547), .B(n3548), .Z(\u_a23_mem/n18744 ) );
  NAND U4598 ( .A(n3539), .B(\u_a23_mem/p_mem[84][4] ), .Z(n3548) );
  OR U4599 ( .A(n1037), .B(n3540), .Z(n3547) );
  NAND U4600 ( .A(n3549), .B(n3550), .Z(\u_a23_mem/n18743 ) );
  NAND U4601 ( .A(n3539), .B(\u_a23_mem/p_mem[84][5] ), .Z(n3550) );
  OR U4602 ( .A(n1043), .B(n3540), .Z(n3549) );
  NAND U4603 ( .A(n3551), .B(n3552), .Z(\u_a23_mem/n18742 ) );
  NAND U4604 ( .A(n3539), .B(\u_a23_mem/p_mem[84][6] ), .Z(n3552) );
  OR U4605 ( .A(n1049), .B(n3540), .Z(n3551) );
  NAND U4606 ( .A(n3553), .B(n3554), .Z(\u_a23_mem/n18741 ) );
  NAND U4607 ( .A(n3539), .B(\u_a23_mem/p_mem[84][7] ), .Z(n3554) );
  NANDN U4608 ( .B(n1080), .A(n3555), .Z(n3539) );
  NANDN U4609 ( .B(n3540), .A(n1055), .Z(n3553) );
  NANDN U4610 ( .B(n2), .A(n3555), .Z(n3540) );
  NAND U4611 ( .A(n3556), .B(n3557), .Z(\u_a23_mem/n18740 ) );
  OR U4612 ( .A(n1011), .B(n3558), .Z(n3557) );
  AND U4613 ( .A(n3559), .B(n3560), .Z(n3556) );
  NANDN U4614 ( .B(n1087), .A(n3555), .Z(n3560) );
  NAND U4615 ( .A(n3561), .B(\u_a23_mem/p_mem[85][0] ), .Z(n3559) );
  NAND U4616 ( .A(n3562), .B(n3563), .Z(\u_a23_mem/n18739 ) );
  OR U4617 ( .A(n1019), .B(n3558), .Z(n3563) );
  AND U4618 ( .A(n3564), .B(n3565), .Z(n3562) );
  NANDN U4619 ( .B(n1093), .A(n3555), .Z(n3565) );
  NAND U4620 ( .A(n3561), .B(\u_a23_mem/p_mem[85][1] ), .Z(n3564) );
  NAND U4621 ( .A(n3566), .B(n3567), .Z(\u_a23_mem/n18738 ) );
  OR U4622 ( .A(n1025), .B(n3558), .Z(n3567) );
  AND U4623 ( .A(n3568), .B(n3569), .Z(n3566) );
  NANDN U4624 ( .B(n1098), .A(n3555), .Z(n3569) );
  NAND U4625 ( .A(n3561), .B(\u_a23_mem/p_mem[85][2] ), .Z(n3568) );
  NAND U4626 ( .A(n3570), .B(n3571), .Z(\u_a23_mem/n18737 ) );
  OR U4627 ( .A(n1031), .B(n3558), .Z(n3571) );
  AND U4628 ( .A(n3572), .B(n3573), .Z(n3570) );
  NANDN U4629 ( .B(n1103), .A(n3555), .Z(n3573) );
  NAND U4630 ( .A(n3561), .B(\u_a23_mem/p_mem[85][3] ), .Z(n3572) );
  NAND U4631 ( .A(n3574), .B(n3575), .Z(\u_a23_mem/n18736 ) );
  OR U4632 ( .A(n1037), .B(n3558), .Z(n3575) );
  AND U4633 ( .A(n3576), .B(n3577), .Z(n3574) );
  NANDN U4634 ( .B(n1108), .A(n3555), .Z(n3577) );
  NAND U4635 ( .A(n3561), .B(\u_a23_mem/p_mem[85][4] ), .Z(n3576) );
  NAND U4636 ( .A(n3578), .B(n3579), .Z(\u_a23_mem/n18735 ) );
  OR U4637 ( .A(n1043), .B(n3558), .Z(n3579) );
  AND U4638 ( .A(n3580), .B(n3581), .Z(n3578) );
  NANDN U4639 ( .B(n1113), .A(n3555), .Z(n3581) );
  NAND U4640 ( .A(n3561), .B(\u_a23_mem/p_mem[85][5] ), .Z(n3580) );
  NAND U4641 ( .A(n3582), .B(n3583), .Z(\u_a23_mem/n18734 ) );
  OR U4642 ( .A(n1049), .B(n3558), .Z(n3583) );
  AND U4643 ( .A(n3584), .B(n3585), .Z(n3582) );
  NANDN U4644 ( .B(n1118), .A(n3555), .Z(n3585) );
  NAND U4645 ( .A(n3561), .B(\u_a23_mem/p_mem[85][6] ), .Z(n3584) );
  NAND U4646 ( .A(n3586), .B(n3587), .Z(\u_a23_mem/n18733 ) );
  NANDN U4647 ( .B(n3558), .A(n1055), .Z(n3587) );
  NAND U4648 ( .A(n1121), .B(n3555), .Z(n3558) );
  AND U4649 ( .A(n3588), .B(n3589), .Z(n3586) );
  NANDN U4650 ( .B(n1124), .A(n3555), .Z(n3589) );
  NAND U4651 ( .A(n3561), .B(\u_a23_mem/p_mem[85][7] ), .Z(n3588) );
  NANDN U4652 ( .B(n1125), .A(n3555), .Z(n3561) );
  NAND U4653 ( .A(n3590), .B(n3591), .Z(\u_a23_mem/n18732 ) );
  OR U4654 ( .A(n1011), .B(n3592), .Z(n3591) );
  AND U4655 ( .A(n3593), .B(n3594), .Z(n3590) );
  NANDN U4656 ( .B(n1131), .A(n3555), .Z(n3594) );
  NAND U4657 ( .A(n3595), .B(\u_a23_mem/p_mem[86][0] ), .Z(n3593) );
  NAND U4658 ( .A(n3596), .B(n3597), .Z(\u_a23_mem/n18731 ) );
  OR U4659 ( .A(n1019), .B(n3592), .Z(n3597) );
  AND U4660 ( .A(n3598), .B(n3599), .Z(n3596) );
  NANDN U4661 ( .B(n1137), .A(n3555), .Z(n3599) );
  NAND U4662 ( .A(n3595), .B(\u_a23_mem/p_mem[86][1] ), .Z(n3598) );
  NAND U4663 ( .A(n3600), .B(n3601), .Z(\u_a23_mem/n18730 ) );
  OR U4664 ( .A(n1025), .B(n3592), .Z(n3601) );
  AND U4665 ( .A(n3602), .B(n3603), .Z(n3600) );
  NANDN U4666 ( .B(n1142), .A(n3555), .Z(n3603) );
  NAND U4667 ( .A(n3595), .B(\u_a23_mem/p_mem[86][2] ), .Z(n3602) );
  NAND U4668 ( .A(n3604), .B(n3605), .Z(\u_a23_mem/n18729 ) );
  OR U4669 ( .A(n1031), .B(n3592), .Z(n3605) );
  AND U4670 ( .A(n3606), .B(n3607), .Z(n3604) );
  NANDN U4671 ( .B(n1147), .A(n3555), .Z(n3607) );
  NAND U4672 ( .A(n3595), .B(\u_a23_mem/p_mem[86][3] ), .Z(n3606) );
  NAND U4673 ( .A(n3608), .B(n3609), .Z(\u_a23_mem/n18728 ) );
  OR U4674 ( .A(n1037), .B(n3592), .Z(n3609) );
  AND U4675 ( .A(n3610), .B(n3611), .Z(n3608) );
  NANDN U4676 ( .B(n1152), .A(n3555), .Z(n3611) );
  NAND U4677 ( .A(n3595), .B(\u_a23_mem/p_mem[86][4] ), .Z(n3610) );
  NAND U4678 ( .A(n3612), .B(n3613), .Z(\u_a23_mem/n18727 ) );
  OR U4679 ( .A(n1043), .B(n3592), .Z(n3613) );
  AND U4680 ( .A(n3614), .B(n3615), .Z(n3612) );
  NANDN U4681 ( .B(n1157), .A(n3555), .Z(n3615) );
  NAND U4682 ( .A(n3595), .B(\u_a23_mem/p_mem[86][5] ), .Z(n3614) );
  NAND U4683 ( .A(n3616), .B(n3617), .Z(\u_a23_mem/n18726 ) );
  OR U4684 ( .A(n1049), .B(n3592), .Z(n3617) );
  AND U4685 ( .A(n3618), .B(n3619), .Z(n3616) );
  NANDN U4686 ( .B(n1162), .A(n3555), .Z(n3619) );
  NAND U4687 ( .A(n3595), .B(\u_a23_mem/p_mem[86][6] ), .Z(n3618) );
  NAND U4688 ( .A(n3620), .B(n3621), .Z(\u_a23_mem/n18725 ) );
  NANDN U4689 ( .B(n3592), .A(n1055), .Z(n3621) );
  NAND U4690 ( .A(n1165), .B(n3555), .Z(n3592) );
  AND U4691 ( .A(n3622), .B(n3623), .Z(n3620) );
  NANDN U4692 ( .B(n1168), .A(n3555), .Z(n3623) );
  NAND U4693 ( .A(n3595), .B(\u_a23_mem/p_mem[86][7] ), .Z(n3622) );
  NANDN U4694 ( .B(n1169), .A(n3555), .Z(n3595) );
  NAND U4695 ( .A(n3624), .B(n3625), .Z(\u_a23_mem/n18724 ) );
  OR U4696 ( .A(n1011), .B(n3626), .Z(n3625) );
  AND U4697 ( .A(n3627), .B(n3628), .Z(n3624) );
  NAND U4698 ( .A(n3629), .B(\u_a23_mem/p_mem[87][0] ), .Z(n3628) );
  NANDN U4699 ( .B(n1015), .A(n3555), .Z(n3627) );
  NAND U4700 ( .A(n3630), .B(n3631), .Z(\u_a23_mem/n18723 ) );
  OR U4701 ( .A(n1019), .B(n3626), .Z(n3631) );
  AND U4702 ( .A(n3632), .B(n3633), .Z(n3630) );
  NAND U4703 ( .A(n3629), .B(\u_a23_mem/p_mem[87][1] ), .Z(n3633) );
  NANDN U4704 ( .B(n1022), .A(n3555), .Z(n3632) );
  NAND U4705 ( .A(n3634), .B(n3635), .Z(\u_a23_mem/n18722 ) );
  OR U4706 ( .A(n1025), .B(n3626), .Z(n3635) );
  AND U4707 ( .A(n3636), .B(n3637), .Z(n3634) );
  NAND U4708 ( .A(n3629), .B(\u_a23_mem/p_mem[87][2] ), .Z(n3637) );
  NANDN U4709 ( .B(n1028), .A(n3555), .Z(n3636) );
  NAND U4710 ( .A(n3638), .B(n3639), .Z(\u_a23_mem/n18721 ) );
  OR U4711 ( .A(n1031), .B(n3626), .Z(n3639) );
  AND U4712 ( .A(n3640), .B(n3641), .Z(n3638) );
  NAND U4713 ( .A(n3629), .B(\u_a23_mem/p_mem[87][3] ), .Z(n3641) );
  NANDN U4714 ( .B(n1034), .A(n3555), .Z(n3640) );
  NAND U4715 ( .A(n3642), .B(n3643), .Z(\u_a23_mem/n18720 ) );
  OR U4716 ( .A(n1037), .B(n3626), .Z(n3643) );
  AND U4717 ( .A(n3644), .B(n3645), .Z(n3642) );
  NAND U4718 ( .A(n3629), .B(\u_a23_mem/p_mem[87][4] ), .Z(n3645) );
  NANDN U4719 ( .B(n1040), .A(n3555), .Z(n3644) );
  NAND U4720 ( .A(n3646), .B(n3647), .Z(\u_a23_mem/n18719 ) );
  OR U4721 ( .A(n1043), .B(n3626), .Z(n3647) );
  AND U4722 ( .A(n3648), .B(n3649), .Z(n3646) );
  NAND U4723 ( .A(n3629), .B(\u_a23_mem/p_mem[87][5] ), .Z(n3649) );
  NANDN U4724 ( .B(n1046), .A(n3555), .Z(n3648) );
  NAND U4725 ( .A(n3650), .B(n3651), .Z(\u_a23_mem/n18718 ) );
  OR U4726 ( .A(n1049), .B(n3626), .Z(n3651) );
  AND U4727 ( .A(n3652), .B(n3653), .Z(n3650) );
  NAND U4728 ( .A(n3629), .B(\u_a23_mem/p_mem[87][6] ), .Z(n3653) );
  NANDN U4729 ( .B(n1052), .A(n3555), .Z(n3652) );
  NAND U4730 ( .A(n3654), .B(n3655), .Z(\u_a23_mem/n18717 ) );
  NANDN U4731 ( .B(n3626), .A(n1055), .Z(n3655) );
  NAND U4732 ( .A(n1056), .B(n3555), .Z(n3626) );
  AND U4733 ( .A(n3656), .B(n3657), .Z(n3654) );
  NAND U4734 ( .A(n3629), .B(\u_a23_mem/p_mem[87][7] ), .Z(n3657) );
  NANDN U4735 ( .B(n1059), .A(n3555), .Z(n3629) );
  NAND U4736 ( .A(n1061), .B(n3555), .Z(n3656) );
  AND U4737 ( .A(n1694), .B(n3658), .Z(n3555) );
  NAND U4738 ( .A(n3659), .B(n3660), .Z(\u_a23_mem/n18716 ) );
  NAND U4739 ( .A(n3661), .B(\u_a23_mem/p_mem[88][0] ), .Z(n3660) );
  OR U4740 ( .A(n1011), .B(n3662), .Z(n3659) );
  NAND U4741 ( .A(n3663), .B(n3664), .Z(\u_a23_mem/n18715 ) );
  NAND U4742 ( .A(n3661), .B(\u_a23_mem/p_mem[88][1] ), .Z(n3664) );
  OR U4743 ( .A(n1019), .B(n3662), .Z(n3663) );
  NAND U4744 ( .A(n3665), .B(n3666), .Z(\u_a23_mem/n18714 ) );
  NAND U4745 ( .A(n3661), .B(\u_a23_mem/p_mem[88][2] ), .Z(n3666) );
  OR U4746 ( .A(n1025), .B(n3662), .Z(n3665) );
  NAND U4747 ( .A(n3667), .B(n3668), .Z(\u_a23_mem/n18713 ) );
  NAND U4748 ( .A(n3661), .B(\u_a23_mem/p_mem[88][3] ), .Z(n3668) );
  OR U4749 ( .A(n1031), .B(n3662), .Z(n3667) );
  NAND U4750 ( .A(n3669), .B(n3670), .Z(\u_a23_mem/n18712 ) );
  NAND U4751 ( .A(n3661), .B(\u_a23_mem/p_mem[88][4] ), .Z(n3670) );
  OR U4752 ( .A(n1037), .B(n3662), .Z(n3669) );
  NAND U4753 ( .A(n3671), .B(n3672), .Z(\u_a23_mem/n18711 ) );
  NAND U4754 ( .A(n3661), .B(\u_a23_mem/p_mem[88][5] ), .Z(n3672) );
  OR U4755 ( .A(n1043), .B(n3662), .Z(n3671) );
  NAND U4756 ( .A(n3673), .B(n3674), .Z(\u_a23_mem/n18710 ) );
  NAND U4757 ( .A(n3661), .B(\u_a23_mem/p_mem[88][6] ), .Z(n3674) );
  OR U4758 ( .A(n1049), .B(n3662), .Z(n3673) );
  NAND U4759 ( .A(n3675), .B(n3676), .Z(\u_a23_mem/n18709 ) );
  NAND U4760 ( .A(n3661), .B(\u_a23_mem/p_mem[88][7] ), .Z(n3676) );
  NANDN U4761 ( .B(n1080), .A(n3677), .Z(n3661) );
  NANDN U4762 ( .B(n3662), .A(n1055), .Z(n3675) );
  NANDN U4763 ( .B(n2), .A(n3677), .Z(n3662) );
  NAND U4764 ( .A(n3678), .B(n3679), .Z(\u_a23_mem/n18708 ) );
  OR U4765 ( .A(n1011), .B(n3680), .Z(n3679) );
  AND U4766 ( .A(n3681), .B(n3682), .Z(n3678) );
  NANDN U4767 ( .B(n1087), .A(n3677), .Z(n3682) );
  NAND U4768 ( .A(n3683), .B(\u_a23_mem/p_mem[89][0] ), .Z(n3681) );
  NAND U4769 ( .A(n3684), .B(n3685), .Z(\u_a23_mem/n18707 ) );
  OR U4770 ( .A(n1019), .B(n3680), .Z(n3685) );
  AND U4771 ( .A(n3686), .B(n3687), .Z(n3684) );
  NANDN U4772 ( .B(n1093), .A(n3677), .Z(n3687) );
  NAND U4773 ( .A(n3683), .B(\u_a23_mem/p_mem[89][1] ), .Z(n3686) );
  NAND U4774 ( .A(n3688), .B(n3689), .Z(\u_a23_mem/n18706 ) );
  OR U4775 ( .A(n1025), .B(n3680), .Z(n3689) );
  AND U4776 ( .A(n3690), .B(n3691), .Z(n3688) );
  NANDN U4777 ( .B(n1098), .A(n3677), .Z(n3691) );
  NAND U4778 ( .A(n3683), .B(\u_a23_mem/p_mem[89][2] ), .Z(n3690) );
  NAND U4779 ( .A(n3692), .B(n3693), .Z(\u_a23_mem/n18705 ) );
  OR U4780 ( .A(n1031), .B(n3680), .Z(n3693) );
  AND U4781 ( .A(n3694), .B(n3695), .Z(n3692) );
  NANDN U4782 ( .B(n1103), .A(n3677), .Z(n3695) );
  NAND U4783 ( .A(n3683), .B(\u_a23_mem/p_mem[89][3] ), .Z(n3694) );
  NAND U4784 ( .A(n3696), .B(n3697), .Z(\u_a23_mem/n18704 ) );
  OR U4785 ( .A(n1037), .B(n3680), .Z(n3697) );
  AND U4786 ( .A(n3698), .B(n3699), .Z(n3696) );
  NANDN U4787 ( .B(n1108), .A(n3677), .Z(n3699) );
  NAND U4788 ( .A(n3683), .B(\u_a23_mem/p_mem[89][4] ), .Z(n3698) );
  NAND U4789 ( .A(n3700), .B(n3701), .Z(\u_a23_mem/n18703 ) );
  OR U4790 ( .A(n1043), .B(n3680), .Z(n3701) );
  AND U4791 ( .A(n3702), .B(n3703), .Z(n3700) );
  NANDN U4792 ( .B(n1113), .A(n3677), .Z(n3703) );
  NAND U4793 ( .A(n3683), .B(\u_a23_mem/p_mem[89][5] ), .Z(n3702) );
  NAND U4794 ( .A(n3704), .B(n3705), .Z(\u_a23_mem/n18702 ) );
  OR U4795 ( .A(n1049), .B(n3680), .Z(n3705) );
  AND U4796 ( .A(n3706), .B(n3707), .Z(n3704) );
  NANDN U4797 ( .B(n1118), .A(n3677), .Z(n3707) );
  NAND U4798 ( .A(n3683), .B(\u_a23_mem/p_mem[89][6] ), .Z(n3706) );
  NAND U4799 ( .A(n3708), .B(n3709), .Z(\u_a23_mem/n18701 ) );
  NANDN U4800 ( .B(n3680), .A(n1055), .Z(n3709) );
  NAND U4801 ( .A(n1121), .B(n3677), .Z(n3680) );
  AND U4802 ( .A(n3710), .B(n3711), .Z(n3708) );
  NANDN U4803 ( .B(n1124), .A(n3677), .Z(n3711) );
  NAND U4804 ( .A(n3683), .B(\u_a23_mem/p_mem[89][7] ), .Z(n3710) );
  NANDN U4805 ( .B(n1125), .A(n3677), .Z(n3683) );
  NAND U4806 ( .A(n3712), .B(n3713), .Z(\u_a23_mem/n18700 ) );
  OR U4807 ( .A(n1011), .B(n3714), .Z(n3713) );
  AND U4808 ( .A(n3715), .B(n3716), .Z(n3712) );
  NANDN U4809 ( .B(n1131), .A(n3677), .Z(n3716) );
  NAND U4810 ( .A(n3717), .B(\u_a23_mem/p_mem[90][0] ), .Z(n3715) );
  NAND U4811 ( .A(n3718), .B(n3719), .Z(\u_a23_mem/n18699 ) );
  OR U4812 ( .A(n1019), .B(n3714), .Z(n3719) );
  AND U4813 ( .A(n3720), .B(n3721), .Z(n3718) );
  NANDN U4814 ( .B(n1137), .A(n3677), .Z(n3721) );
  NAND U4815 ( .A(n3717), .B(\u_a23_mem/p_mem[90][1] ), .Z(n3720) );
  NAND U4816 ( .A(n3722), .B(n3723), .Z(\u_a23_mem/n18698 ) );
  OR U4817 ( .A(n1025), .B(n3714), .Z(n3723) );
  AND U4818 ( .A(n3724), .B(n3725), .Z(n3722) );
  NANDN U4819 ( .B(n1142), .A(n3677), .Z(n3725) );
  NAND U4820 ( .A(n3717), .B(\u_a23_mem/p_mem[90][2] ), .Z(n3724) );
  NAND U4821 ( .A(n3726), .B(n3727), .Z(\u_a23_mem/n18697 ) );
  OR U4822 ( .A(n1031), .B(n3714), .Z(n3727) );
  AND U4823 ( .A(n3728), .B(n3729), .Z(n3726) );
  NANDN U4824 ( .B(n1147), .A(n3677), .Z(n3729) );
  NAND U4825 ( .A(n3717), .B(\u_a23_mem/p_mem[90][3] ), .Z(n3728) );
  NAND U4826 ( .A(n3730), .B(n3731), .Z(\u_a23_mem/n18696 ) );
  OR U4827 ( .A(n1037), .B(n3714), .Z(n3731) );
  AND U4828 ( .A(n3732), .B(n3733), .Z(n3730) );
  NANDN U4829 ( .B(n1152), .A(n3677), .Z(n3733) );
  NAND U4830 ( .A(n3717), .B(\u_a23_mem/p_mem[90][4] ), .Z(n3732) );
  NAND U4831 ( .A(n3734), .B(n3735), .Z(\u_a23_mem/n18695 ) );
  OR U4832 ( .A(n1043), .B(n3714), .Z(n3735) );
  AND U4833 ( .A(n3736), .B(n3737), .Z(n3734) );
  NANDN U4834 ( .B(n1157), .A(n3677), .Z(n3737) );
  NAND U4835 ( .A(n3717), .B(\u_a23_mem/p_mem[90][5] ), .Z(n3736) );
  NAND U4836 ( .A(n3738), .B(n3739), .Z(\u_a23_mem/n18694 ) );
  OR U4837 ( .A(n1049), .B(n3714), .Z(n3739) );
  AND U4838 ( .A(n3740), .B(n3741), .Z(n3738) );
  NANDN U4839 ( .B(n1162), .A(n3677), .Z(n3741) );
  NAND U4840 ( .A(n3717), .B(\u_a23_mem/p_mem[90][6] ), .Z(n3740) );
  NAND U4841 ( .A(n3742), .B(n3743), .Z(\u_a23_mem/n18693 ) );
  NANDN U4842 ( .B(n3714), .A(n1055), .Z(n3743) );
  NAND U4843 ( .A(n1165), .B(n3677), .Z(n3714) );
  AND U4844 ( .A(n3744), .B(n3745), .Z(n3742) );
  NANDN U4845 ( .B(n1168), .A(n3677), .Z(n3745) );
  NAND U4846 ( .A(n3717), .B(\u_a23_mem/p_mem[90][7] ), .Z(n3744) );
  NANDN U4847 ( .B(n1169), .A(n3677), .Z(n3717) );
  NAND U4848 ( .A(n3746), .B(n3747), .Z(\u_a23_mem/n18692 ) );
  OR U4849 ( .A(n1011), .B(n3748), .Z(n3747) );
  AND U4850 ( .A(n3749), .B(n3750), .Z(n3746) );
  NAND U4851 ( .A(n3751), .B(\u_a23_mem/p_mem[91][0] ), .Z(n3750) );
  NANDN U4852 ( .B(n1015), .A(n3677), .Z(n3749) );
  NAND U4853 ( .A(n3752), .B(n3753), .Z(\u_a23_mem/n18691 ) );
  OR U4854 ( .A(n1019), .B(n3748), .Z(n3753) );
  AND U4855 ( .A(n3754), .B(n3755), .Z(n3752) );
  NAND U4856 ( .A(n3751), .B(\u_a23_mem/p_mem[91][1] ), .Z(n3755) );
  NANDN U4857 ( .B(n1022), .A(n3677), .Z(n3754) );
  NAND U4858 ( .A(n3756), .B(n3757), .Z(\u_a23_mem/n18690 ) );
  OR U4859 ( .A(n1025), .B(n3748), .Z(n3757) );
  AND U4860 ( .A(n3758), .B(n3759), .Z(n3756) );
  NAND U4861 ( .A(n3751), .B(\u_a23_mem/p_mem[91][2] ), .Z(n3759) );
  NANDN U4862 ( .B(n1028), .A(n3677), .Z(n3758) );
  NAND U4863 ( .A(n3760), .B(n3761), .Z(\u_a23_mem/n18689 ) );
  OR U4864 ( .A(n1031), .B(n3748), .Z(n3761) );
  AND U4865 ( .A(n3762), .B(n3763), .Z(n3760) );
  NAND U4866 ( .A(n3751), .B(\u_a23_mem/p_mem[91][3] ), .Z(n3763) );
  NANDN U4867 ( .B(n1034), .A(n3677), .Z(n3762) );
  NAND U4868 ( .A(n3764), .B(n3765), .Z(\u_a23_mem/n18688 ) );
  OR U4869 ( .A(n1037), .B(n3748), .Z(n3765) );
  AND U4870 ( .A(n3766), .B(n3767), .Z(n3764) );
  NAND U4871 ( .A(n3751), .B(\u_a23_mem/p_mem[91][4] ), .Z(n3767) );
  NANDN U4872 ( .B(n1040), .A(n3677), .Z(n3766) );
  NAND U4873 ( .A(n3768), .B(n3769), .Z(\u_a23_mem/n18687 ) );
  OR U4874 ( .A(n1043), .B(n3748), .Z(n3769) );
  AND U4875 ( .A(n3770), .B(n3771), .Z(n3768) );
  NAND U4876 ( .A(n3751), .B(\u_a23_mem/p_mem[91][5] ), .Z(n3771) );
  NANDN U4877 ( .B(n1046), .A(n3677), .Z(n3770) );
  NAND U4878 ( .A(n3772), .B(n3773), .Z(\u_a23_mem/n18686 ) );
  OR U4879 ( .A(n1049), .B(n3748), .Z(n3773) );
  AND U4880 ( .A(n3774), .B(n3775), .Z(n3772) );
  NAND U4881 ( .A(n3751), .B(\u_a23_mem/p_mem[91][6] ), .Z(n3775) );
  NANDN U4882 ( .B(n1052), .A(n3677), .Z(n3774) );
  NAND U4883 ( .A(n3776), .B(n3777), .Z(\u_a23_mem/n18685 ) );
  NANDN U4884 ( .B(n3748), .A(n1055), .Z(n3777) );
  NAND U4885 ( .A(n1056), .B(n3677), .Z(n3748) );
  AND U4886 ( .A(n3778), .B(n3779), .Z(n3776) );
  NAND U4887 ( .A(n3751), .B(\u_a23_mem/p_mem[91][7] ), .Z(n3779) );
  NANDN U4888 ( .B(n1059), .A(n3677), .Z(n3751) );
  NAND U4889 ( .A(n1061), .B(n3677), .Z(n3778) );
  AND U4890 ( .A(n1816), .B(n3658), .Z(n3677) );
  NAND U4891 ( .A(n3780), .B(n3781), .Z(\u_a23_mem/n18684 ) );
  NAND U4892 ( .A(n3782), .B(\u_a23_mem/p_mem[92][0] ), .Z(n3781) );
  OR U4893 ( .A(n1011), .B(n3783), .Z(n3780) );
  NAND U4894 ( .A(n3784), .B(n3785), .Z(\u_a23_mem/n18683 ) );
  NAND U4895 ( .A(n3782), .B(\u_a23_mem/p_mem[92][1] ), .Z(n3785) );
  OR U4896 ( .A(n1019), .B(n3783), .Z(n3784) );
  NAND U4897 ( .A(n3786), .B(n3787), .Z(\u_a23_mem/n18682 ) );
  NAND U4898 ( .A(n3782), .B(\u_a23_mem/p_mem[92][2] ), .Z(n3787) );
  OR U4899 ( .A(n1025), .B(n3783), .Z(n3786) );
  NAND U4900 ( .A(n3788), .B(n3789), .Z(\u_a23_mem/n18681 ) );
  NAND U4901 ( .A(n3782), .B(\u_a23_mem/p_mem[92][3] ), .Z(n3789) );
  OR U4902 ( .A(n1031), .B(n3783), .Z(n3788) );
  NAND U4903 ( .A(n3790), .B(n3791), .Z(\u_a23_mem/n18680 ) );
  NAND U4904 ( .A(n3782), .B(\u_a23_mem/p_mem[92][4] ), .Z(n3791) );
  OR U4905 ( .A(n1037), .B(n3783), .Z(n3790) );
  NAND U4906 ( .A(n3792), .B(n3793), .Z(\u_a23_mem/n18679 ) );
  NAND U4907 ( .A(n3782), .B(\u_a23_mem/p_mem[92][5] ), .Z(n3793) );
  OR U4908 ( .A(n1043), .B(n3783), .Z(n3792) );
  NAND U4909 ( .A(n3794), .B(n3795), .Z(\u_a23_mem/n18678 ) );
  NAND U4910 ( .A(n3782), .B(\u_a23_mem/p_mem[92][6] ), .Z(n3795) );
  OR U4911 ( .A(n1049), .B(n3783), .Z(n3794) );
  NAND U4912 ( .A(n3796), .B(n3797), .Z(\u_a23_mem/n18677 ) );
  NAND U4913 ( .A(n3782), .B(\u_a23_mem/p_mem[92][7] ), .Z(n3797) );
  NANDN U4914 ( .B(n1080), .A(n3798), .Z(n3782) );
  NANDN U4915 ( .B(n3783), .A(n1055), .Z(n3796) );
  NANDN U4916 ( .B(n2), .A(n3798), .Z(n3783) );
  NAND U4917 ( .A(n3799), .B(n3800), .Z(\u_a23_mem/n18676 ) );
  OR U4918 ( .A(n1011), .B(n3801), .Z(n3800) );
  AND U4919 ( .A(n3802), .B(n3803), .Z(n3799) );
  NANDN U4920 ( .B(n1087), .A(n3798), .Z(n3803) );
  NAND U4921 ( .A(n3804), .B(\u_a23_mem/p_mem[93][0] ), .Z(n3802) );
  NAND U4922 ( .A(n3805), .B(n3806), .Z(\u_a23_mem/n18675 ) );
  OR U4923 ( .A(n1019), .B(n3801), .Z(n3806) );
  AND U4924 ( .A(n3807), .B(n3808), .Z(n3805) );
  NANDN U4925 ( .B(n1093), .A(n3798), .Z(n3808) );
  NAND U4926 ( .A(n3804), .B(\u_a23_mem/p_mem[93][1] ), .Z(n3807) );
  NAND U4927 ( .A(n3809), .B(n3810), .Z(\u_a23_mem/n18674 ) );
  OR U4928 ( .A(n1025), .B(n3801), .Z(n3810) );
  AND U4929 ( .A(n3811), .B(n3812), .Z(n3809) );
  NANDN U4930 ( .B(n1098), .A(n3798), .Z(n3812) );
  NAND U4931 ( .A(n3804), .B(\u_a23_mem/p_mem[93][2] ), .Z(n3811) );
  NAND U4932 ( .A(n3813), .B(n3814), .Z(\u_a23_mem/n18673 ) );
  OR U4933 ( .A(n1031), .B(n3801), .Z(n3814) );
  AND U4934 ( .A(n3815), .B(n3816), .Z(n3813) );
  NANDN U4935 ( .B(n1103), .A(n3798), .Z(n3816) );
  NAND U4936 ( .A(n3804), .B(\u_a23_mem/p_mem[93][3] ), .Z(n3815) );
  NAND U4937 ( .A(n3817), .B(n3818), .Z(\u_a23_mem/n18672 ) );
  OR U4938 ( .A(n1037), .B(n3801), .Z(n3818) );
  AND U4939 ( .A(n3819), .B(n3820), .Z(n3817) );
  NANDN U4940 ( .B(n1108), .A(n3798), .Z(n3820) );
  NAND U4941 ( .A(n3804), .B(\u_a23_mem/p_mem[93][4] ), .Z(n3819) );
  NAND U4942 ( .A(n3821), .B(n3822), .Z(\u_a23_mem/n18671 ) );
  OR U4943 ( .A(n1043), .B(n3801), .Z(n3822) );
  AND U4944 ( .A(n3823), .B(n3824), .Z(n3821) );
  NANDN U4945 ( .B(n1113), .A(n3798), .Z(n3824) );
  NAND U4946 ( .A(n3804), .B(\u_a23_mem/p_mem[93][5] ), .Z(n3823) );
  NAND U4947 ( .A(n3825), .B(n3826), .Z(\u_a23_mem/n18670 ) );
  OR U4948 ( .A(n1049), .B(n3801), .Z(n3826) );
  AND U4949 ( .A(n3827), .B(n3828), .Z(n3825) );
  NANDN U4950 ( .B(n1118), .A(n3798), .Z(n3828) );
  NAND U4951 ( .A(n3804), .B(\u_a23_mem/p_mem[93][6] ), .Z(n3827) );
  NAND U4952 ( .A(n3829), .B(n3830), .Z(\u_a23_mem/n18669 ) );
  NANDN U4953 ( .B(n3801), .A(n1055), .Z(n3830) );
  NAND U4954 ( .A(n1121), .B(n3798), .Z(n3801) );
  AND U4955 ( .A(n3831), .B(n3832), .Z(n3829) );
  NANDN U4956 ( .B(n1124), .A(n3798), .Z(n3832) );
  NAND U4957 ( .A(n3804), .B(\u_a23_mem/p_mem[93][7] ), .Z(n3831) );
  NANDN U4958 ( .B(n1125), .A(n3798), .Z(n3804) );
  NAND U4959 ( .A(n3833), .B(n3834), .Z(\u_a23_mem/n18668 ) );
  OR U4960 ( .A(n1011), .B(n3835), .Z(n3834) );
  AND U4961 ( .A(n3836), .B(n3837), .Z(n3833) );
  NANDN U4962 ( .B(n1131), .A(n3798), .Z(n3837) );
  NAND U4963 ( .A(n3838), .B(\u_a23_mem/p_mem[94][0] ), .Z(n3836) );
  NAND U4964 ( .A(n3839), .B(n3840), .Z(\u_a23_mem/n18667 ) );
  OR U4965 ( .A(n1019), .B(n3835), .Z(n3840) );
  AND U4966 ( .A(n3841), .B(n3842), .Z(n3839) );
  NANDN U4967 ( .B(n1137), .A(n3798), .Z(n3842) );
  NAND U4968 ( .A(n3838), .B(\u_a23_mem/p_mem[94][1] ), .Z(n3841) );
  NAND U4969 ( .A(n3843), .B(n3844), .Z(\u_a23_mem/n18666 ) );
  OR U4970 ( .A(n1025), .B(n3835), .Z(n3844) );
  AND U4971 ( .A(n3845), .B(n3846), .Z(n3843) );
  NANDN U4972 ( .B(n1142), .A(n3798), .Z(n3846) );
  NAND U4973 ( .A(n3838), .B(\u_a23_mem/p_mem[94][2] ), .Z(n3845) );
  NAND U4974 ( .A(n3847), .B(n3848), .Z(\u_a23_mem/n18665 ) );
  OR U4975 ( .A(n1031), .B(n3835), .Z(n3848) );
  AND U4976 ( .A(n3849), .B(n3850), .Z(n3847) );
  NANDN U4977 ( .B(n1147), .A(n3798), .Z(n3850) );
  NAND U4978 ( .A(n3838), .B(\u_a23_mem/p_mem[94][3] ), .Z(n3849) );
  NAND U4979 ( .A(n3851), .B(n3852), .Z(\u_a23_mem/n18664 ) );
  OR U4980 ( .A(n1037), .B(n3835), .Z(n3852) );
  AND U4981 ( .A(n3853), .B(n3854), .Z(n3851) );
  NANDN U4982 ( .B(n1152), .A(n3798), .Z(n3854) );
  NAND U4983 ( .A(n3838), .B(\u_a23_mem/p_mem[94][4] ), .Z(n3853) );
  NAND U4984 ( .A(n3855), .B(n3856), .Z(\u_a23_mem/n18663 ) );
  OR U4985 ( .A(n1043), .B(n3835), .Z(n3856) );
  AND U4986 ( .A(n3857), .B(n3858), .Z(n3855) );
  NANDN U4987 ( .B(n1157), .A(n3798), .Z(n3858) );
  NAND U4988 ( .A(n3838), .B(\u_a23_mem/p_mem[94][5] ), .Z(n3857) );
  NAND U4989 ( .A(n3859), .B(n3860), .Z(\u_a23_mem/n18662 ) );
  OR U4990 ( .A(n1049), .B(n3835), .Z(n3860) );
  AND U4991 ( .A(n3861), .B(n3862), .Z(n3859) );
  NANDN U4992 ( .B(n1162), .A(n3798), .Z(n3862) );
  NAND U4993 ( .A(n3838), .B(\u_a23_mem/p_mem[94][6] ), .Z(n3861) );
  NAND U4994 ( .A(n3863), .B(n3864), .Z(\u_a23_mem/n18661 ) );
  NANDN U4995 ( .B(n3835), .A(n1055), .Z(n3864) );
  NAND U4996 ( .A(n1165), .B(n3798), .Z(n3835) );
  AND U4997 ( .A(n3865), .B(n3866), .Z(n3863) );
  NANDN U4998 ( .B(n1168), .A(n3798), .Z(n3866) );
  NAND U4999 ( .A(n3838), .B(\u_a23_mem/p_mem[94][7] ), .Z(n3865) );
  NANDN U5000 ( .B(n1169), .A(n3798), .Z(n3838) );
  NAND U5001 ( .A(n3867), .B(n3868), .Z(\u_a23_mem/n18660 ) );
  OR U5002 ( .A(n1011), .B(n3869), .Z(n3868) );
  AND U5003 ( .A(n3870), .B(n3871), .Z(n3867) );
  NAND U5004 ( .A(n3872), .B(\u_a23_mem/p_mem[95][0] ), .Z(n3871) );
  NANDN U5005 ( .B(n1015), .A(n3798), .Z(n3870) );
  NAND U5006 ( .A(n3873), .B(n3874), .Z(\u_a23_mem/n18659 ) );
  OR U5007 ( .A(n1019), .B(n3869), .Z(n3874) );
  AND U5008 ( .A(n3875), .B(n3876), .Z(n3873) );
  NAND U5009 ( .A(n3872), .B(\u_a23_mem/p_mem[95][1] ), .Z(n3876) );
  NANDN U5010 ( .B(n1022), .A(n3798), .Z(n3875) );
  NAND U5011 ( .A(n3877), .B(n3878), .Z(\u_a23_mem/n18658 ) );
  OR U5012 ( .A(n1025), .B(n3869), .Z(n3878) );
  AND U5013 ( .A(n3879), .B(n3880), .Z(n3877) );
  NAND U5014 ( .A(n3872), .B(\u_a23_mem/p_mem[95][2] ), .Z(n3880) );
  NANDN U5015 ( .B(n1028), .A(n3798), .Z(n3879) );
  NAND U5016 ( .A(n3881), .B(n3882), .Z(\u_a23_mem/n18657 ) );
  OR U5017 ( .A(n1031), .B(n3869), .Z(n3882) );
  AND U5018 ( .A(n3883), .B(n3884), .Z(n3881) );
  NAND U5019 ( .A(n3872), .B(\u_a23_mem/p_mem[95][3] ), .Z(n3884) );
  NANDN U5020 ( .B(n1034), .A(n3798), .Z(n3883) );
  NAND U5021 ( .A(n3885), .B(n3886), .Z(\u_a23_mem/n18656 ) );
  OR U5022 ( .A(n1037), .B(n3869), .Z(n3886) );
  AND U5023 ( .A(n3887), .B(n3888), .Z(n3885) );
  NAND U5024 ( .A(n3872), .B(\u_a23_mem/p_mem[95][4] ), .Z(n3888) );
  NANDN U5025 ( .B(n1040), .A(n3798), .Z(n3887) );
  NAND U5026 ( .A(n3889), .B(n3890), .Z(\u_a23_mem/n18655 ) );
  OR U5027 ( .A(n1043), .B(n3869), .Z(n3890) );
  AND U5028 ( .A(n3891), .B(n3892), .Z(n3889) );
  NAND U5029 ( .A(n3872), .B(\u_a23_mem/p_mem[95][5] ), .Z(n3892) );
  NANDN U5030 ( .B(n1046), .A(n3798), .Z(n3891) );
  NAND U5031 ( .A(n3893), .B(n3894), .Z(\u_a23_mem/n18654 ) );
  OR U5032 ( .A(n1049), .B(n3869), .Z(n3894) );
  AND U5033 ( .A(n3895), .B(n3896), .Z(n3893) );
  NAND U5034 ( .A(n3872), .B(\u_a23_mem/p_mem[95][6] ), .Z(n3896) );
  NANDN U5035 ( .B(n1052), .A(n3798), .Z(n3895) );
  NAND U5036 ( .A(n3897), .B(n3898), .Z(\u_a23_mem/n18653 ) );
  NANDN U5037 ( .B(n3869), .A(n1055), .Z(n3898) );
  NAND U5038 ( .A(n1056), .B(n3798), .Z(n3869) );
  AND U5039 ( .A(n3899), .B(n3900), .Z(n3897) );
  NAND U5040 ( .A(n3872), .B(\u_a23_mem/p_mem[95][7] ), .Z(n3900) );
  NANDN U5041 ( .B(n1059), .A(n3798), .Z(n3872) );
  NAND U5042 ( .A(n1061), .B(n3798), .Z(n3899) );
  NOR U5043 ( .A(n3536), .B(n1938), .Z(n3798) );
  IV U5044 ( .A(n3658), .Z(n3536) );
  ANDN U5045 ( .A(n3901), .B(n2429), .Z(n3658) );
  AND U5046 ( .A(n2428), .B(m_address[4]), .Z(n3901) );
  NAND U5047 ( .A(n3902), .B(n3903), .Z(\u_a23_mem/n18652 ) );
  NAND U5048 ( .A(n3904), .B(\u_a23_mem/p_mem[96][0] ), .Z(n3903) );
  OR U5049 ( .A(n1011), .B(n3905), .Z(n3902) );
  NAND U5050 ( .A(n3906), .B(n3907), .Z(\u_a23_mem/n18651 ) );
  NAND U5051 ( .A(n3904), .B(\u_a23_mem/p_mem[96][1] ), .Z(n3907) );
  OR U5052 ( .A(n1019), .B(n3905), .Z(n3906) );
  NAND U5053 ( .A(n3908), .B(n3909), .Z(\u_a23_mem/n18650 ) );
  NAND U5054 ( .A(n3904), .B(\u_a23_mem/p_mem[96][2] ), .Z(n3909) );
  OR U5055 ( .A(n1025), .B(n3905), .Z(n3908) );
  NAND U5056 ( .A(n3910), .B(n3911), .Z(\u_a23_mem/n18649 ) );
  NAND U5057 ( .A(n3904), .B(\u_a23_mem/p_mem[96][3] ), .Z(n3911) );
  OR U5058 ( .A(n1031), .B(n3905), .Z(n3910) );
  NAND U5059 ( .A(n3912), .B(n3913), .Z(\u_a23_mem/n18648 ) );
  NAND U5060 ( .A(n3904), .B(\u_a23_mem/p_mem[96][4] ), .Z(n3913) );
  OR U5061 ( .A(n1037), .B(n3905), .Z(n3912) );
  NAND U5062 ( .A(n3914), .B(n3915), .Z(\u_a23_mem/n18647 ) );
  NAND U5063 ( .A(n3904), .B(\u_a23_mem/p_mem[96][5] ), .Z(n3915) );
  OR U5064 ( .A(n1043), .B(n3905), .Z(n3914) );
  NAND U5065 ( .A(n3916), .B(n3917), .Z(\u_a23_mem/n18646 ) );
  NAND U5066 ( .A(n3904), .B(\u_a23_mem/p_mem[96][6] ), .Z(n3917) );
  OR U5067 ( .A(n1049), .B(n3905), .Z(n3916) );
  NAND U5068 ( .A(n3918), .B(n3919), .Z(\u_a23_mem/n18645 ) );
  NAND U5069 ( .A(n3904), .B(\u_a23_mem/p_mem[96][7] ), .Z(n3919) );
  NANDN U5070 ( .B(n1080), .A(n3920), .Z(n3904) );
  NANDN U5071 ( .B(n3905), .A(n1055), .Z(n3918) );
  NANDN U5072 ( .B(n2), .A(n3920), .Z(n3905) );
  NAND U5073 ( .A(n3921), .B(n3922), .Z(\u_a23_mem/n18644 ) );
  OR U5074 ( .A(n1011), .B(n3923), .Z(n3922) );
  AND U5075 ( .A(n3924), .B(n3925), .Z(n3921) );
  NANDN U5076 ( .B(n1087), .A(n3920), .Z(n3925) );
  NAND U5077 ( .A(n3926), .B(\u_a23_mem/p_mem[97][0] ), .Z(n3924) );
  NAND U5078 ( .A(n3927), .B(n3928), .Z(\u_a23_mem/n18643 ) );
  OR U5079 ( .A(n1019), .B(n3923), .Z(n3928) );
  AND U5080 ( .A(n3929), .B(n3930), .Z(n3927) );
  NANDN U5081 ( .B(n1093), .A(n3920), .Z(n3930) );
  NAND U5082 ( .A(n3926), .B(\u_a23_mem/p_mem[97][1] ), .Z(n3929) );
  NAND U5083 ( .A(n3931), .B(n3932), .Z(\u_a23_mem/n18642 ) );
  OR U5084 ( .A(n1025), .B(n3923), .Z(n3932) );
  AND U5085 ( .A(n3933), .B(n3934), .Z(n3931) );
  NANDN U5086 ( .B(n1098), .A(n3920), .Z(n3934) );
  NAND U5087 ( .A(n3926), .B(\u_a23_mem/p_mem[97][2] ), .Z(n3933) );
  NAND U5088 ( .A(n3935), .B(n3936), .Z(\u_a23_mem/n18641 ) );
  OR U5089 ( .A(n1031), .B(n3923), .Z(n3936) );
  AND U5090 ( .A(n3937), .B(n3938), .Z(n3935) );
  NANDN U5091 ( .B(n1103), .A(n3920), .Z(n3938) );
  NAND U5092 ( .A(n3926), .B(\u_a23_mem/p_mem[97][3] ), .Z(n3937) );
  NAND U5093 ( .A(n3939), .B(n3940), .Z(\u_a23_mem/n18640 ) );
  OR U5094 ( .A(n1037), .B(n3923), .Z(n3940) );
  AND U5095 ( .A(n3941), .B(n3942), .Z(n3939) );
  NANDN U5096 ( .B(n1108), .A(n3920), .Z(n3942) );
  NAND U5097 ( .A(n3926), .B(\u_a23_mem/p_mem[97][4] ), .Z(n3941) );
  NAND U5098 ( .A(n3943), .B(n3944), .Z(\u_a23_mem/n18639 ) );
  OR U5099 ( .A(n1043), .B(n3923), .Z(n3944) );
  AND U5100 ( .A(n3945), .B(n3946), .Z(n3943) );
  NANDN U5101 ( .B(n1113), .A(n3920), .Z(n3946) );
  NAND U5102 ( .A(n3926), .B(\u_a23_mem/p_mem[97][5] ), .Z(n3945) );
  NAND U5103 ( .A(n3947), .B(n3948), .Z(\u_a23_mem/n18638 ) );
  OR U5104 ( .A(n1049), .B(n3923), .Z(n3948) );
  AND U5105 ( .A(n3949), .B(n3950), .Z(n3947) );
  NANDN U5106 ( .B(n1118), .A(n3920), .Z(n3950) );
  NAND U5107 ( .A(n3926), .B(\u_a23_mem/p_mem[97][6] ), .Z(n3949) );
  NAND U5108 ( .A(n3951), .B(n3952), .Z(\u_a23_mem/n18637 ) );
  NANDN U5109 ( .B(n3923), .A(n1055), .Z(n3952) );
  NAND U5110 ( .A(n1121), .B(n3920), .Z(n3923) );
  AND U5111 ( .A(n3953), .B(n3954), .Z(n3951) );
  NANDN U5112 ( .B(n1124), .A(n3920), .Z(n3954) );
  NAND U5113 ( .A(n3926), .B(\u_a23_mem/p_mem[97][7] ), .Z(n3953) );
  NANDN U5114 ( .B(n1125), .A(n3920), .Z(n3926) );
  NAND U5115 ( .A(n3955), .B(n3956), .Z(\u_a23_mem/n18636 ) );
  OR U5116 ( .A(n1011), .B(n3957), .Z(n3956) );
  AND U5117 ( .A(n3958), .B(n3959), .Z(n3955) );
  NANDN U5118 ( .B(n1131), .A(n3920), .Z(n3959) );
  NAND U5119 ( .A(n3960), .B(\u_a23_mem/p_mem[98][0] ), .Z(n3958) );
  NAND U5120 ( .A(n3961), .B(n3962), .Z(\u_a23_mem/n18635 ) );
  OR U5121 ( .A(n1019), .B(n3957), .Z(n3962) );
  AND U5122 ( .A(n3963), .B(n3964), .Z(n3961) );
  NANDN U5123 ( .B(n1137), .A(n3920), .Z(n3964) );
  NAND U5124 ( .A(n3960), .B(\u_a23_mem/p_mem[98][1] ), .Z(n3963) );
  NAND U5125 ( .A(n3965), .B(n3966), .Z(\u_a23_mem/n18634 ) );
  OR U5126 ( .A(n1025), .B(n3957), .Z(n3966) );
  AND U5127 ( .A(n3967), .B(n3968), .Z(n3965) );
  NANDN U5128 ( .B(n1142), .A(n3920), .Z(n3968) );
  NAND U5129 ( .A(n3960), .B(\u_a23_mem/p_mem[98][2] ), .Z(n3967) );
  NAND U5130 ( .A(n3969), .B(n3970), .Z(\u_a23_mem/n18633 ) );
  OR U5131 ( .A(n1031), .B(n3957), .Z(n3970) );
  AND U5132 ( .A(n3971), .B(n3972), .Z(n3969) );
  NANDN U5133 ( .B(n1147), .A(n3920), .Z(n3972) );
  NAND U5134 ( .A(n3960), .B(\u_a23_mem/p_mem[98][3] ), .Z(n3971) );
  NAND U5135 ( .A(n3973), .B(n3974), .Z(\u_a23_mem/n18632 ) );
  OR U5136 ( .A(n1037), .B(n3957), .Z(n3974) );
  AND U5137 ( .A(n3975), .B(n3976), .Z(n3973) );
  NANDN U5138 ( .B(n1152), .A(n3920), .Z(n3976) );
  NAND U5139 ( .A(n3960), .B(\u_a23_mem/p_mem[98][4] ), .Z(n3975) );
  NAND U5140 ( .A(n3977), .B(n3978), .Z(\u_a23_mem/n18631 ) );
  OR U5141 ( .A(n1043), .B(n3957), .Z(n3978) );
  AND U5142 ( .A(n3979), .B(n3980), .Z(n3977) );
  NANDN U5143 ( .B(n1157), .A(n3920), .Z(n3980) );
  NAND U5144 ( .A(n3960), .B(\u_a23_mem/p_mem[98][5] ), .Z(n3979) );
  NAND U5145 ( .A(n3981), .B(n3982), .Z(\u_a23_mem/n18630 ) );
  OR U5146 ( .A(n1049), .B(n3957), .Z(n3982) );
  AND U5147 ( .A(n3983), .B(n3984), .Z(n3981) );
  NANDN U5148 ( .B(n1162), .A(n3920), .Z(n3984) );
  NAND U5149 ( .A(n3960), .B(\u_a23_mem/p_mem[98][6] ), .Z(n3983) );
  NAND U5150 ( .A(n3985), .B(n3986), .Z(\u_a23_mem/n18629 ) );
  NANDN U5151 ( .B(n3957), .A(n1055), .Z(n3986) );
  NAND U5152 ( .A(n1165), .B(n3920), .Z(n3957) );
  AND U5153 ( .A(n3987), .B(n3988), .Z(n3985) );
  NANDN U5154 ( .B(n1168), .A(n3920), .Z(n3988) );
  NAND U5155 ( .A(n3960), .B(\u_a23_mem/p_mem[98][7] ), .Z(n3987) );
  NANDN U5156 ( .B(n1169), .A(n3920), .Z(n3960) );
  NAND U5157 ( .A(n3989), .B(n3990), .Z(\u_a23_mem/n18628 ) );
  OR U5158 ( .A(n1011), .B(n3991), .Z(n3990) );
  AND U5159 ( .A(n3992), .B(n3993), .Z(n3989) );
  NAND U5160 ( .A(n3994), .B(\u_a23_mem/p_mem[99][0] ), .Z(n3993) );
  NANDN U5161 ( .B(n1015), .A(n3920), .Z(n3992) );
  NAND U5162 ( .A(n3995), .B(n3996), .Z(\u_a23_mem/n18627 ) );
  OR U5163 ( .A(n1019), .B(n3991), .Z(n3996) );
  AND U5164 ( .A(n3997), .B(n3998), .Z(n3995) );
  NAND U5165 ( .A(n3994), .B(\u_a23_mem/p_mem[99][1] ), .Z(n3998) );
  NANDN U5166 ( .B(n1022), .A(n3920), .Z(n3997) );
  NAND U5167 ( .A(n3999), .B(n4000), .Z(\u_a23_mem/n18626 ) );
  OR U5168 ( .A(n1025), .B(n3991), .Z(n4000) );
  AND U5169 ( .A(n4001), .B(n4002), .Z(n3999) );
  NAND U5170 ( .A(n3994), .B(\u_a23_mem/p_mem[99][2] ), .Z(n4002) );
  NANDN U5171 ( .B(n1028), .A(n3920), .Z(n4001) );
  NAND U5172 ( .A(n4003), .B(n4004), .Z(\u_a23_mem/n18625 ) );
  OR U5173 ( .A(n1031), .B(n3991), .Z(n4004) );
  AND U5174 ( .A(n4005), .B(n4006), .Z(n4003) );
  NAND U5175 ( .A(n3994), .B(\u_a23_mem/p_mem[99][3] ), .Z(n4006) );
  NANDN U5176 ( .B(n1034), .A(n3920), .Z(n4005) );
  NAND U5177 ( .A(n4007), .B(n4008), .Z(\u_a23_mem/n18624 ) );
  OR U5178 ( .A(n1037), .B(n3991), .Z(n4008) );
  AND U5179 ( .A(n4009), .B(n4010), .Z(n4007) );
  NAND U5180 ( .A(n3994), .B(\u_a23_mem/p_mem[99][4] ), .Z(n4010) );
  NANDN U5181 ( .B(n1040), .A(n3920), .Z(n4009) );
  NAND U5182 ( .A(n4011), .B(n4012), .Z(\u_a23_mem/n18623 ) );
  OR U5183 ( .A(n1043), .B(n3991), .Z(n4012) );
  AND U5184 ( .A(n4013), .B(n4014), .Z(n4011) );
  NAND U5185 ( .A(n3994), .B(\u_a23_mem/p_mem[99][5] ), .Z(n4014) );
  NANDN U5186 ( .B(n1046), .A(n3920), .Z(n4013) );
  NAND U5187 ( .A(n4015), .B(n4016), .Z(\u_a23_mem/n18622 ) );
  OR U5188 ( .A(n1049), .B(n3991), .Z(n4016) );
  AND U5189 ( .A(n4017), .B(n4018), .Z(n4015) );
  NAND U5190 ( .A(n3994), .B(\u_a23_mem/p_mem[99][6] ), .Z(n4018) );
  NANDN U5191 ( .B(n1052), .A(n3920), .Z(n4017) );
  NAND U5192 ( .A(n4019), .B(n4020), .Z(\u_a23_mem/n18621 ) );
  NANDN U5193 ( .B(n3991), .A(n1055), .Z(n4020) );
  NAND U5194 ( .A(n1056), .B(n3920), .Z(n3991) );
  AND U5195 ( .A(n4021), .B(n4022), .Z(n4019) );
  NAND U5196 ( .A(n3994), .B(\u_a23_mem/p_mem[99][7] ), .Z(n4022) );
  NANDN U5197 ( .B(n1059), .A(n3920), .Z(n3994) );
  NAND U5198 ( .A(n1061), .B(n3920), .Z(n4021) );
  ANDN U5199 ( .A(n1571), .B(n4023), .Z(n3920) );
  NAND U5200 ( .A(n4024), .B(n4025), .Z(\u_a23_mem/n18620 ) );
  NAND U5201 ( .A(n4026), .B(\u_a23_mem/p_mem[100][0] ), .Z(n4025) );
  OR U5202 ( .A(n1011), .B(n4027), .Z(n4024) );
  NAND U5203 ( .A(n4028), .B(n4029), .Z(\u_a23_mem/n18619 ) );
  NAND U5204 ( .A(n4026), .B(\u_a23_mem/p_mem[100][1] ), .Z(n4029) );
  OR U5205 ( .A(n1019), .B(n4027), .Z(n4028) );
  NAND U5206 ( .A(n4030), .B(n4031), .Z(\u_a23_mem/n18618 ) );
  NAND U5207 ( .A(n4026), .B(\u_a23_mem/p_mem[100][2] ), .Z(n4031) );
  OR U5208 ( .A(n1025), .B(n4027), .Z(n4030) );
  NAND U5209 ( .A(n4032), .B(n4033), .Z(\u_a23_mem/n18617 ) );
  NAND U5210 ( .A(n4026), .B(\u_a23_mem/p_mem[100][3] ), .Z(n4033) );
  OR U5211 ( .A(n1031), .B(n4027), .Z(n4032) );
  NAND U5212 ( .A(n4034), .B(n4035), .Z(\u_a23_mem/n18616 ) );
  NAND U5213 ( .A(n4026), .B(\u_a23_mem/p_mem[100][4] ), .Z(n4035) );
  OR U5214 ( .A(n1037), .B(n4027), .Z(n4034) );
  NAND U5215 ( .A(n4036), .B(n4037), .Z(\u_a23_mem/n18615 ) );
  NAND U5216 ( .A(n4026), .B(\u_a23_mem/p_mem[100][5] ), .Z(n4037) );
  OR U5217 ( .A(n1043), .B(n4027), .Z(n4036) );
  NAND U5218 ( .A(n4038), .B(n4039), .Z(\u_a23_mem/n18614 ) );
  NAND U5219 ( .A(n4026), .B(\u_a23_mem/p_mem[100][6] ), .Z(n4039) );
  OR U5220 ( .A(n1049), .B(n4027), .Z(n4038) );
  NAND U5221 ( .A(n4040), .B(n4041), .Z(\u_a23_mem/n18613 ) );
  NAND U5222 ( .A(n4026), .B(\u_a23_mem/p_mem[100][7] ), .Z(n4041) );
  NANDN U5223 ( .B(n1080), .A(n4042), .Z(n4026) );
  NANDN U5224 ( .B(n4027), .A(n1055), .Z(n4040) );
  NANDN U5225 ( .B(n2), .A(n4042), .Z(n4027) );
  NAND U5226 ( .A(n4043), .B(n4044), .Z(\u_a23_mem/n18612 ) );
  OR U5227 ( .A(n1011), .B(n4045), .Z(n4044) );
  AND U5228 ( .A(n4046), .B(n4047), .Z(n4043) );
  NANDN U5229 ( .B(n1087), .A(n4042), .Z(n4047) );
  NAND U5230 ( .A(n4048), .B(\u_a23_mem/p_mem[101][0] ), .Z(n4046) );
  NAND U5231 ( .A(n4049), .B(n4050), .Z(\u_a23_mem/n18611 ) );
  OR U5232 ( .A(n1019), .B(n4045), .Z(n4050) );
  AND U5233 ( .A(n4051), .B(n4052), .Z(n4049) );
  NANDN U5234 ( .B(n1093), .A(n4042), .Z(n4052) );
  NAND U5235 ( .A(n4048), .B(\u_a23_mem/p_mem[101][1] ), .Z(n4051) );
  NAND U5236 ( .A(n4053), .B(n4054), .Z(\u_a23_mem/n18610 ) );
  OR U5237 ( .A(n1025), .B(n4045), .Z(n4054) );
  AND U5238 ( .A(n4055), .B(n4056), .Z(n4053) );
  NANDN U5239 ( .B(n1098), .A(n4042), .Z(n4056) );
  NAND U5240 ( .A(n4048), .B(\u_a23_mem/p_mem[101][2] ), .Z(n4055) );
  NAND U5241 ( .A(n4057), .B(n4058), .Z(\u_a23_mem/n18609 ) );
  OR U5242 ( .A(n1031), .B(n4045), .Z(n4058) );
  AND U5243 ( .A(n4059), .B(n4060), .Z(n4057) );
  NANDN U5244 ( .B(n1103), .A(n4042), .Z(n4060) );
  NAND U5245 ( .A(n4048), .B(\u_a23_mem/p_mem[101][3] ), .Z(n4059) );
  NAND U5246 ( .A(n4061), .B(n4062), .Z(\u_a23_mem/n18608 ) );
  OR U5247 ( .A(n1037), .B(n4045), .Z(n4062) );
  AND U5248 ( .A(n4063), .B(n4064), .Z(n4061) );
  NANDN U5249 ( .B(n1108), .A(n4042), .Z(n4064) );
  NAND U5250 ( .A(n4048), .B(\u_a23_mem/p_mem[101][4] ), .Z(n4063) );
  NAND U5251 ( .A(n4065), .B(n4066), .Z(\u_a23_mem/n18607 ) );
  OR U5252 ( .A(n1043), .B(n4045), .Z(n4066) );
  AND U5253 ( .A(n4067), .B(n4068), .Z(n4065) );
  NANDN U5254 ( .B(n1113), .A(n4042), .Z(n4068) );
  NAND U5255 ( .A(n4048), .B(\u_a23_mem/p_mem[101][5] ), .Z(n4067) );
  NAND U5256 ( .A(n4069), .B(n4070), .Z(\u_a23_mem/n18606 ) );
  OR U5257 ( .A(n1049), .B(n4045), .Z(n4070) );
  AND U5258 ( .A(n4071), .B(n4072), .Z(n4069) );
  NANDN U5259 ( .B(n1118), .A(n4042), .Z(n4072) );
  NAND U5260 ( .A(n4048), .B(\u_a23_mem/p_mem[101][6] ), .Z(n4071) );
  NAND U5261 ( .A(n4073), .B(n4074), .Z(\u_a23_mem/n18605 ) );
  NANDN U5262 ( .B(n4045), .A(n1055), .Z(n4074) );
  NAND U5263 ( .A(n1121), .B(n4042), .Z(n4045) );
  AND U5264 ( .A(n4075), .B(n4076), .Z(n4073) );
  NANDN U5265 ( .B(n1124), .A(n4042), .Z(n4076) );
  NAND U5266 ( .A(n4048), .B(\u_a23_mem/p_mem[101][7] ), .Z(n4075) );
  NANDN U5267 ( .B(n1125), .A(n4042), .Z(n4048) );
  NAND U5268 ( .A(n4077), .B(n4078), .Z(\u_a23_mem/n18604 ) );
  OR U5269 ( .A(n1011), .B(n4079), .Z(n4078) );
  AND U5270 ( .A(n4080), .B(n4081), .Z(n4077) );
  NANDN U5271 ( .B(n1131), .A(n4042), .Z(n4081) );
  NAND U5272 ( .A(n4082), .B(\u_a23_mem/p_mem[102][0] ), .Z(n4080) );
  NAND U5273 ( .A(n4083), .B(n4084), .Z(\u_a23_mem/n18603 ) );
  OR U5274 ( .A(n1019), .B(n4079), .Z(n4084) );
  AND U5275 ( .A(n4085), .B(n4086), .Z(n4083) );
  NANDN U5276 ( .B(n1137), .A(n4042), .Z(n4086) );
  NAND U5277 ( .A(n4082), .B(\u_a23_mem/p_mem[102][1] ), .Z(n4085) );
  NAND U5278 ( .A(n4087), .B(n4088), .Z(\u_a23_mem/n18602 ) );
  OR U5279 ( .A(n1025), .B(n4079), .Z(n4088) );
  AND U5280 ( .A(n4089), .B(n4090), .Z(n4087) );
  NANDN U5281 ( .B(n1142), .A(n4042), .Z(n4090) );
  NAND U5282 ( .A(n4082), .B(\u_a23_mem/p_mem[102][2] ), .Z(n4089) );
  NAND U5283 ( .A(n4091), .B(n4092), .Z(\u_a23_mem/n18601 ) );
  OR U5284 ( .A(n1031), .B(n4079), .Z(n4092) );
  AND U5285 ( .A(n4093), .B(n4094), .Z(n4091) );
  NANDN U5286 ( .B(n1147), .A(n4042), .Z(n4094) );
  NAND U5287 ( .A(n4082), .B(\u_a23_mem/p_mem[102][3] ), .Z(n4093) );
  NAND U5288 ( .A(n4095), .B(n4096), .Z(\u_a23_mem/n18600 ) );
  OR U5289 ( .A(n1037), .B(n4079), .Z(n4096) );
  AND U5290 ( .A(n4097), .B(n4098), .Z(n4095) );
  NANDN U5291 ( .B(n1152), .A(n4042), .Z(n4098) );
  NAND U5292 ( .A(n4082), .B(\u_a23_mem/p_mem[102][4] ), .Z(n4097) );
  NAND U5293 ( .A(n4099), .B(n4100), .Z(\u_a23_mem/n18599 ) );
  OR U5294 ( .A(n1043), .B(n4079), .Z(n4100) );
  AND U5295 ( .A(n4101), .B(n4102), .Z(n4099) );
  NANDN U5296 ( .B(n1157), .A(n4042), .Z(n4102) );
  NAND U5297 ( .A(n4082), .B(\u_a23_mem/p_mem[102][5] ), .Z(n4101) );
  NAND U5298 ( .A(n4103), .B(n4104), .Z(\u_a23_mem/n18598 ) );
  OR U5299 ( .A(n1049), .B(n4079), .Z(n4104) );
  AND U5300 ( .A(n4105), .B(n4106), .Z(n4103) );
  NANDN U5301 ( .B(n1162), .A(n4042), .Z(n4106) );
  NAND U5302 ( .A(n4082), .B(\u_a23_mem/p_mem[102][6] ), .Z(n4105) );
  NAND U5303 ( .A(n4107), .B(n4108), .Z(\u_a23_mem/n18597 ) );
  NANDN U5304 ( .B(n4079), .A(n1055), .Z(n4108) );
  NAND U5305 ( .A(n1165), .B(n4042), .Z(n4079) );
  AND U5306 ( .A(n4109), .B(n4110), .Z(n4107) );
  NANDN U5307 ( .B(n1168), .A(n4042), .Z(n4110) );
  NAND U5308 ( .A(n4082), .B(\u_a23_mem/p_mem[102][7] ), .Z(n4109) );
  NANDN U5309 ( .B(n1169), .A(n4042), .Z(n4082) );
  NAND U5310 ( .A(n4111), .B(n4112), .Z(\u_a23_mem/n18596 ) );
  OR U5311 ( .A(n1011), .B(n4113), .Z(n4112) );
  AND U5312 ( .A(n4114), .B(n4115), .Z(n4111) );
  NAND U5313 ( .A(n4116), .B(\u_a23_mem/p_mem[103][0] ), .Z(n4115) );
  NANDN U5314 ( .B(n1015), .A(n4042), .Z(n4114) );
  NAND U5315 ( .A(n4117), .B(n4118), .Z(\u_a23_mem/n18595 ) );
  OR U5316 ( .A(n1019), .B(n4113), .Z(n4118) );
  AND U5317 ( .A(n4119), .B(n4120), .Z(n4117) );
  NAND U5318 ( .A(n4116), .B(\u_a23_mem/p_mem[103][1] ), .Z(n4120) );
  NANDN U5319 ( .B(n1022), .A(n4042), .Z(n4119) );
  NAND U5320 ( .A(n4121), .B(n4122), .Z(\u_a23_mem/n18594 ) );
  OR U5321 ( .A(n1025), .B(n4113), .Z(n4122) );
  AND U5322 ( .A(n4123), .B(n4124), .Z(n4121) );
  NAND U5323 ( .A(n4116), .B(\u_a23_mem/p_mem[103][2] ), .Z(n4124) );
  NANDN U5324 ( .B(n1028), .A(n4042), .Z(n4123) );
  NAND U5325 ( .A(n4125), .B(n4126), .Z(\u_a23_mem/n18593 ) );
  OR U5326 ( .A(n1031), .B(n4113), .Z(n4126) );
  AND U5327 ( .A(n4127), .B(n4128), .Z(n4125) );
  NAND U5328 ( .A(n4116), .B(\u_a23_mem/p_mem[103][3] ), .Z(n4128) );
  NANDN U5329 ( .B(n1034), .A(n4042), .Z(n4127) );
  NAND U5330 ( .A(n4129), .B(n4130), .Z(\u_a23_mem/n18592 ) );
  OR U5331 ( .A(n1037), .B(n4113), .Z(n4130) );
  AND U5332 ( .A(n4131), .B(n4132), .Z(n4129) );
  NAND U5333 ( .A(n4116), .B(\u_a23_mem/p_mem[103][4] ), .Z(n4132) );
  NANDN U5334 ( .B(n1040), .A(n4042), .Z(n4131) );
  NAND U5335 ( .A(n4133), .B(n4134), .Z(\u_a23_mem/n18591 ) );
  OR U5336 ( .A(n1043), .B(n4113), .Z(n4134) );
  AND U5337 ( .A(n4135), .B(n4136), .Z(n4133) );
  NAND U5338 ( .A(n4116), .B(\u_a23_mem/p_mem[103][5] ), .Z(n4136) );
  NANDN U5339 ( .B(n1046), .A(n4042), .Z(n4135) );
  NAND U5340 ( .A(n4137), .B(n4138), .Z(\u_a23_mem/n18590 ) );
  OR U5341 ( .A(n1049), .B(n4113), .Z(n4138) );
  AND U5342 ( .A(n4139), .B(n4140), .Z(n4137) );
  NAND U5343 ( .A(n4116), .B(\u_a23_mem/p_mem[103][6] ), .Z(n4140) );
  NANDN U5344 ( .B(n1052), .A(n4042), .Z(n4139) );
  NAND U5345 ( .A(n4141), .B(n4142), .Z(\u_a23_mem/n18589 ) );
  NANDN U5346 ( .B(n4113), .A(n1055), .Z(n4142) );
  NAND U5347 ( .A(n1056), .B(n4042), .Z(n4113) );
  AND U5348 ( .A(n4143), .B(n4144), .Z(n4141) );
  NAND U5349 ( .A(n4116), .B(\u_a23_mem/p_mem[103][7] ), .Z(n4144) );
  NANDN U5350 ( .B(n1059), .A(n4042), .Z(n4116) );
  NAND U5351 ( .A(n1061), .B(n4042), .Z(n4143) );
  ANDN U5352 ( .A(n1694), .B(n4023), .Z(n4042) );
  ANDN U5353 ( .A(n4145), .B(n4146), .Z(n1694) );
  AND U5354 ( .A(n4147), .B(n4148), .Z(n4145) );
  NAND U5355 ( .A(n4149), .B(n4150), .Z(\u_a23_mem/n18588 ) );
  NAND U5356 ( .A(n4151), .B(\u_a23_mem/p_mem[104][0] ), .Z(n4150) );
  OR U5357 ( .A(n1011), .B(n4152), .Z(n4149) );
  NAND U5358 ( .A(n4153), .B(n4154), .Z(\u_a23_mem/n18587 ) );
  NAND U5359 ( .A(n4151), .B(\u_a23_mem/p_mem[104][1] ), .Z(n4154) );
  OR U5360 ( .A(n1019), .B(n4152), .Z(n4153) );
  NAND U5361 ( .A(n4155), .B(n4156), .Z(\u_a23_mem/n18586 ) );
  NAND U5362 ( .A(n4151), .B(\u_a23_mem/p_mem[104][2] ), .Z(n4156) );
  OR U5363 ( .A(n1025), .B(n4152), .Z(n4155) );
  NAND U5364 ( .A(n4157), .B(n4158), .Z(\u_a23_mem/n18585 ) );
  NAND U5365 ( .A(n4151), .B(\u_a23_mem/p_mem[104][3] ), .Z(n4158) );
  OR U5366 ( .A(n1031), .B(n4152), .Z(n4157) );
  NAND U5367 ( .A(n4159), .B(n4160), .Z(\u_a23_mem/n18584 ) );
  NAND U5368 ( .A(n4151), .B(\u_a23_mem/p_mem[104][4] ), .Z(n4160) );
  OR U5369 ( .A(n1037), .B(n4152), .Z(n4159) );
  NAND U5370 ( .A(n4161), .B(n4162), .Z(\u_a23_mem/n18583 ) );
  NAND U5371 ( .A(n4151), .B(\u_a23_mem/p_mem[104][5] ), .Z(n4162) );
  OR U5372 ( .A(n1043), .B(n4152), .Z(n4161) );
  NAND U5373 ( .A(n4163), .B(n4164), .Z(\u_a23_mem/n18582 ) );
  NAND U5374 ( .A(n4151), .B(\u_a23_mem/p_mem[104][6] ), .Z(n4164) );
  OR U5375 ( .A(n1049), .B(n4152), .Z(n4163) );
  NAND U5376 ( .A(n4165), .B(n4166), .Z(\u_a23_mem/n18581 ) );
  NAND U5377 ( .A(n4151), .B(\u_a23_mem/p_mem[104][7] ), .Z(n4166) );
  NANDN U5378 ( .B(n1080), .A(n4167), .Z(n4151) );
  NANDN U5379 ( .B(n4152), .A(n1055), .Z(n4165) );
  NANDN U5380 ( .B(n2), .A(n4167), .Z(n4152) );
  NAND U5381 ( .A(n4168), .B(n4169), .Z(\u_a23_mem/n18580 ) );
  OR U5382 ( .A(n1011), .B(n4170), .Z(n4169) );
  AND U5383 ( .A(n4171), .B(n4172), .Z(n4168) );
  NANDN U5384 ( .B(n1087), .A(n4167), .Z(n4172) );
  NAND U5385 ( .A(n4173), .B(\u_a23_mem/p_mem[105][0] ), .Z(n4171) );
  NAND U5386 ( .A(n4174), .B(n4175), .Z(\u_a23_mem/n18579 ) );
  OR U5387 ( .A(n1019), .B(n4170), .Z(n4175) );
  AND U5388 ( .A(n4176), .B(n4177), .Z(n4174) );
  NANDN U5389 ( .B(n1093), .A(n4167), .Z(n4177) );
  NAND U5390 ( .A(n4173), .B(\u_a23_mem/p_mem[105][1] ), .Z(n4176) );
  NAND U5391 ( .A(n4178), .B(n4179), .Z(\u_a23_mem/n18578 ) );
  OR U5392 ( .A(n1025), .B(n4170), .Z(n4179) );
  AND U5393 ( .A(n4180), .B(n4181), .Z(n4178) );
  NANDN U5394 ( .B(n1098), .A(n4167), .Z(n4181) );
  NAND U5395 ( .A(n4173), .B(\u_a23_mem/p_mem[105][2] ), .Z(n4180) );
  NAND U5396 ( .A(n4182), .B(n4183), .Z(\u_a23_mem/n18577 ) );
  OR U5397 ( .A(n1031), .B(n4170), .Z(n4183) );
  AND U5398 ( .A(n4184), .B(n4185), .Z(n4182) );
  NANDN U5399 ( .B(n1103), .A(n4167), .Z(n4185) );
  NAND U5400 ( .A(n4173), .B(\u_a23_mem/p_mem[105][3] ), .Z(n4184) );
  NAND U5401 ( .A(n4186), .B(n4187), .Z(\u_a23_mem/n18576 ) );
  OR U5402 ( .A(n1037), .B(n4170), .Z(n4187) );
  AND U5403 ( .A(n4188), .B(n4189), .Z(n4186) );
  NANDN U5404 ( .B(n1108), .A(n4167), .Z(n4189) );
  NAND U5405 ( .A(n4173), .B(\u_a23_mem/p_mem[105][4] ), .Z(n4188) );
  NAND U5406 ( .A(n4190), .B(n4191), .Z(\u_a23_mem/n18575 ) );
  OR U5407 ( .A(n1043), .B(n4170), .Z(n4191) );
  AND U5408 ( .A(n4192), .B(n4193), .Z(n4190) );
  NANDN U5409 ( .B(n1113), .A(n4167), .Z(n4193) );
  NAND U5410 ( .A(n4173), .B(\u_a23_mem/p_mem[105][5] ), .Z(n4192) );
  NAND U5411 ( .A(n4194), .B(n4195), .Z(\u_a23_mem/n18574 ) );
  OR U5412 ( .A(n1049), .B(n4170), .Z(n4195) );
  AND U5413 ( .A(n4196), .B(n4197), .Z(n4194) );
  NANDN U5414 ( .B(n1118), .A(n4167), .Z(n4197) );
  NAND U5415 ( .A(n4173), .B(\u_a23_mem/p_mem[105][6] ), .Z(n4196) );
  NAND U5416 ( .A(n4198), .B(n4199), .Z(\u_a23_mem/n18573 ) );
  NANDN U5417 ( .B(n4170), .A(n1055), .Z(n4199) );
  NAND U5418 ( .A(n1121), .B(n4167), .Z(n4170) );
  AND U5419 ( .A(n4200), .B(n4201), .Z(n4198) );
  NANDN U5420 ( .B(n1124), .A(n4167), .Z(n4201) );
  NAND U5421 ( .A(n4173), .B(\u_a23_mem/p_mem[105][7] ), .Z(n4200) );
  NANDN U5422 ( .B(n1125), .A(n4167), .Z(n4173) );
  NAND U5423 ( .A(n4202), .B(n4203), .Z(\u_a23_mem/n18572 ) );
  OR U5424 ( .A(n1011), .B(n4204), .Z(n4203) );
  AND U5425 ( .A(n4205), .B(n4206), .Z(n4202) );
  NANDN U5426 ( .B(n1131), .A(n4167), .Z(n4206) );
  NAND U5427 ( .A(n4207), .B(\u_a23_mem/p_mem[106][0] ), .Z(n4205) );
  NAND U5428 ( .A(n4208), .B(n4209), .Z(\u_a23_mem/n18571 ) );
  OR U5429 ( .A(n1019), .B(n4204), .Z(n4209) );
  AND U5430 ( .A(n4210), .B(n4211), .Z(n4208) );
  NANDN U5431 ( .B(n1137), .A(n4167), .Z(n4211) );
  NAND U5432 ( .A(n4207), .B(\u_a23_mem/p_mem[106][1] ), .Z(n4210) );
  NAND U5433 ( .A(n4212), .B(n4213), .Z(\u_a23_mem/n18570 ) );
  OR U5434 ( .A(n1025), .B(n4204), .Z(n4213) );
  AND U5435 ( .A(n4214), .B(n4215), .Z(n4212) );
  NANDN U5436 ( .B(n1142), .A(n4167), .Z(n4215) );
  NAND U5437 ( .A(n4207), .B(\u_a23_mem/p_mem[106][2] ), .Z(n4214) );
  NAND U5438 ( .A(n4216), .B(n4217), .Z(\u_a23_mem/n18569 ) );
  OR U5439 ( .A(n1031), .B(n4204), .Z(n4217) );
  AND U5440 ( .A(n4218), .B(n4219), .Z(n4216) );
  NANDN U5441 ( .B(n1147), .A(n4167), .Z(n4219) );
  NAND U5442 ( .A(n4207), .B(\u_a23_mem/p_mem[106][3] ), .Z(n4218) );
  NAND U5443 ( .A(n4220), .B(n4221), .Z(\u_a23_mem/n18568 ) );
  OR U5444 ( .A(n1037), .B(n4204), .Z(n4221) );
  AND U5445 ( .A(n4222), .B(n4223), .Z(n4220) );
  NANDN U5446 ( .B(n1152), .A(n4167), .Z(n4223) );
  NAND U5447 ( .A(n4207), .B(\u_a23_mem/p_mem[106][4] ), .Z(n4222) );
  NAND U5448 ( .A(n4224), .B(n4225), .Z(\u_a23_mem/n18567 ) );
  OR U5449 ( .A(n1043), .B(n4204), .Z(n4225) );
  AND U5450 ( .A(n4226), .B(n4227), .Z(n4224) );
  NANDN U5451 ( .B(n1157), .A(n4167), .Z(n4227) );
  NAND U5452 ( .A(n4207), .B(\u_a23_mem/p_mem[106][5] ), .Z(n4226) );
  NAND U5453 ( .A(n4228), .B(n4229), .Z(\u_a23_mem/n18566 ) );
  OR U5454 ( .A(n1049), .B(n4204), .Z(n4229) );
  AND U5455 ( .A(n4230), .B(n4231), .Z(n4228) );
  NANDN U5456 ( .B(n1162), .A(n4167), .Z(n4231) );
  NAND U5457 ( .A(n4207), .B(\u_a23_mem/p_mem[106][6] ), .Z(n4230) );
  NAND U5458 ( .A(n4232), .B(n4233), .Z(\u_a23_mem/n18565 ) );
  NANDN U5459 ( .B(n4204), .A(n1055), .Z(n4233) );
  NAND U5460 ( .A(n1165), .B(n4167), .Z(n4204) );
  AND U5461 ( .A(n4234), .B(n4235), .Z(n4232) );
  NANDN U5462 ( .B(n1168), .A(n4167), .Z(n4235) );
  NAND U5463 ( .A(n4207), .B(\u_a23_mem/p_mem[106][7] ), .Z(n4234) );
  NANDN U5464 ( .B(n1169), .A(n4167), .Z(n4207) );
  NAND U5465 ( .A(n4236), .B(n4237), .Z(\u_a23_mem/n18564 ) );
  OR U5466 ( .A(n1011), .B(n4238), .Z(n4237) );
  AND U5467 ( .A(n4239), .B(n4240), .Z(n4236) );
  NAND U5468 ( .A(n4241), .B(\u_a23_mem/p_mem[107][0] ), .Z(n4240) );
  NANDN U5469 ( .B(n1015), .A(n4167), .Z(n4239) );
  NAND U5470 ( .A(n4242), .B(n4243), .Z(\u_a23_mem/n18563 ) );
  OR U5471 ( .A(n1019), .B(n4238), .Z(n4243) );
  AND U5472 ( .A(n4244), .B(n4245), .Z(n4242) );
  NAND U5473 ( .A(n4241), .B(\u_a23_mem/p_mem[107][1] ), .Z(n4245) );
  NANDN U5474 ( .B(n1022), .A(n4167), .Z(n4244) );
  NAND U5475 ( .A(n4246), .B(n4247), .Z(\u_a23_mem/n18562 ) );
  OR U5476 ( .A(n1025), .B(n4238), .Z(n4247) );
  AND U5477 ( .A(n4248), .B(n4249), .Z(n4246) );
  NAND U5478 ( .A(n4241), .B(\u_a23_mem/p_mem[107][2] ), .Z(n4249) );
  NANDN U5479 ( .B(n1028), .A(n4167), .Z(n4248) );
  NAND U5480 ( .A(n4250), .B(n4251), .Z(\u_a23_mem/n18561 ) );
  OR U5481 ( .A(n1031), .B(n4238), .Z(n4251) );
  AND U5482 ( .A(n4252), .B(n4253), .Z(n4250) );
  NAND U5483 ( .A(n4241), .B(\u_a23_mem/p_mem[107][3] ), .Z(n4253) );
  NANDN U5484 ( .B(n1034), .A(n4167), .Z(n4252) );
  NAND U5485 ( .A(n4254), .B(n4255), .Z(\u_a23_mem/n18560 ) );
  OR U5486 ( .A(n1037), .B(n4238), .Z(n4255) );
  AND U5487 ( .A(n4256), .B(n4257), .Z(n4254) );
  NAND U5488 ( .A(n4241), .B(\u_a23_mem/p_mem[107][4] ), .Z(n4257) );
  NANDN U5489 ( .B(n1040), .A(n4167), .Z(n4256) );
  NAND U5490 ( .A(n4258), .B(n4259), .Z(\u_a23_mem/n18559 ) );
  OR U5491 ( .A(n1043), .B(n4238), .Z(n4259) );
  AND U5492 ( .A(n4260), .B(n4261), .Z(n4258) );
  NAND U5493 ( .A(n4241), .B(\u_a23_mem/p_mem[107][5] ), .Z(n4261) );
  NANDN U5494 ( .B(n1046), .A(n4167), .Z(n4260) );
  NAND U5495 ( .A(n4262), .B(n4263), .Z(\u_a23_mem/n18558 ) );
  OR U5496 ( .A(n1049), .B(n4238), .Z(n4263) );
  AND U5497 ( .A(n4264), .B(n4265), .Z(n4262) );
  NAND U5498 ( .A(n4241), .B(\u_a23_mem/p_mem[107][6] ), .Z(n4265) );
  NANDN U5499 ( .B(n1052), .A(n4167), .Z(n4264) );
  NAND U5500 ( .A(n4266), .B(n4267), .Z(\u_a23_mem/n18557 ) );
  NANDN U5501 ( .B(n4238), .A(n1055), .Z(n4267) );
  NAND U5502 ( .A(n1056), .B(n4167), .Z(n4238) );
  AND U5503 ( .A(n4268), .B(n4269), .Z(n4266) );
  NAND U5504 ( .A(n4241), .B(\u_a23_mem/p_mem[107][7] ), .Z(n4269) );
  NANDN U5505 ( .B(n1059), .A(n4167), .Z(n4241) );
  NAND U5506 ( .A(n1061), .B(n4167), .Z(n4268) );
  ANDN U5507 ( .A(n1816), .B(n4023), .Z(n4167) );
  ANDN U5508 ( .A(n4270), .B(n4147), .Z(n1816) );
  AND U5509 ( .A(n4146), .B(n4148), .Z(n4270) );
  NAND U5510 ( .A(n4271), .B(n4272), .Z(\u_a23_mem/n18556 ) );
  NAND U5511 ( .A(n4273), .B(\u_a23_mem/p_mem[108][0] ), .Z(n4272) );
  OR U5512 ( .A(n1011), .B(n4274), .Z(n4271) );
  NAND U5513 ( .A(n4275), .B(n4276), .Z(\u_a23_mem/n18555 ) );
  NAND U5514 ( .A(n4273), .B(\u_a23_mem/p_mem[108][1] ), .Z(n4276) );
  OR U5515 ( .A(n1019), .B(n4274), .Z(n4275) );
  NAND U5516 ( .A(n4277), .B(n4278), .Z(\u_a23_mem/n18554 ) );
  NAND U5517 ( .A(n4273), .B(\u_a23_mem/p_mem[108][2] ), .Z(n4278) );
  OR U5518 ( .A(n1025), .B(n4274), .Z(n4277) );
  NAND U5519 ( .A(n4279), .B(n4280), .Z(\u_a23_mem/n18553 ) );
  NAND U5520 ( .A(n4273), .B(\u_a23_mem/p_mem[108][3] ), .Z(n4280) );
  OR U5521 ( .A(n1031), .B(n4274), .Z(n4279) );
  NAND U5522 ( .A(n4281), .B(n4282), .Z(\u_a23_mem/n18552 ) );
  NAND U5523 ( .A(n4273), .B(\u_a23_mem/p_mem[108][4] ), .Z(n4282) );
  OR U5524 ( .A(n1037), .B(n4274), .Z(n4281) );
  NAND U5525 ( .A(n4283), .B(n4284), .Z(\u_a23_mem/n18551 ) );
  NAND U5526 ( .A(n4273), .B(\u_a23_mem/p_mem[108][5] ), .Z(n4284) );
  OR U5527 ( .A(n1043), .B(n4274), .Z(n4283) );
  NAND U5528 ( .A(n4285), .B(n4286), .Z(\u_a23_mem/n18550 ) );
  NAND U5529 ( .A(n4273), .B(\u_a23_mem/p_mem[108][6] ), .Z(n4286) );
  OR U5530 ( .A(n1049), .B(n4274), .Z(n4285) );
  NAND U5531 ( .A(n4287), .B(n4288), .Z(\u_a23_mem/n18549 ) );
  NAND U5532 ( .A(n4273), .B(\u_a23_mem/p_mem[108][7] ), .Z(n4288) );
  NANDN U5533 ( .B(n1080), .A(n4289), .Z(n4273) );
  NANDN U5534 ( .B(n4274), .A(n1055), .Z(n4287) );
  NANDN U5535 ( .B(n2), .A(n4289), .Z(n4274) );
  NAND U5536 ( .A(n4290), .B(n4291), .Z(\u_a23_mem/n18548 ) );
  OR U5537 ( .A(n1011), .B(n4292), .Z(n4291) );
  AND U5538 ( .A(n4293), .B(n4294), .Z(n4290) );
  NANDN U5539 ( .B(n1087), .A(n4289), .Z(n4294) );
  NAND U5540 ( .A(n4295), .B(\u_a23_mem/p_mem[109][0] ), .Z(n4293) );
  NAND U5541 ( .A(n4296), .B(n4297), .Z(\u_a23_mem/n18547 ) );
  OR U5542 ( .A(n1019), .B(n4292), .Z(n4297) );
  AND U5543 ( .A(n4298), .B(n4299), .Z(n4296) );
  NANDN U5544 ( .B(n1093), .A(n4289), .Z(n4299) );
  NAND U5545 ( .A(n4295), .B(\u_a23_mem/p_mem[109][1] ), .Z(n4298) );
  NAND U5546 ( .A(n4300), .B(n4301), .Z(\u_a23_mem/n18546 ) );
  OR U5547 ( .A(n1025), .B(n4292), .Z(n4301) );
  AND U5548 ( .A(n4302), .B(n4303), .Z(n4300) );
  NANDN U5549 ( .B(n1098), .A(n4289), .Z(n4303) );
  NAND U5550 ( .A(n4295), .B(\u_a23_mem/p_mem[109][2] ), .Z(n4302) );
  NAND U5551 ( .A(n4304), .B(n4305), .Z(\u_a23_mem/n18545 ) );
  OR U5552 ( .A(n1031), .B(n4292), .Z(n4305) );
  AND U5553 ( .A(n4306), .B(n4307), .Z(n4304) );
  NANDN U5554 ( .B(n1103), .A(n4289), .Z(n4307) );
  NAND U5555 ( .A(n4295), .B(\u_a23_mem/p_mem[109][3] ), .Z(n4306) );
  NAND U5556 ( .A(n4308), .B(n4309), .Z(\u_a23_mem/n18544 ) );
  OR U5557 ( .A(n1037), .B(n4292), .Z(n4309) );
  AND U5558 ( .A(n4310), .B(n4311), .Z(n4308) );
  NANDN U5559 ( .B(n1108), .A(n4289), .Z(n4311) );
  NAND U5560 ( .A(n4295), .B(\u_a23_mem/p_mem[109][4] ), .Z(n4310) );
  NAND U5561 ( .A(n4312), .B(n4313), .Z(\u_a23_mem/n18543 ) );
  OR U5562 ( .A(n1043), .B(n4292), .Z(n4313) );
  AND U5563 ( .A(n4314), .B(n4315), .Z(n4312) );
  NANDN U5564 ( .B(n1113), .A(n4289), .Z(n4315) );
  NAND U5565 ( .A(n4295), .B(\u_a23_mem/p_mem[109][5] ), .Z(n4314) );
  NAND U5566 ( .A(n4316), .B(n4317), .Z(\u_a23_mem/n18542 ) );
  OR U5567 ( .A(n1049), .B(n4292), .Z(n4317) );
  AND U5568 ( .A(n4318), .B(n4319), .Z(n4316) );
  NANDN U5569 ( .B(n1118), .A(n4289), .Z(n4319) );
  NAND U5570 ( .A(n4295), .B(\u_a23_mem/p_mem[109][6] ), .Z(n4318) );
  NAND U5571 ( .A(n4320), .B(n4321), .Z(\u_a23_mem/n18541 ) );
  NANDN U5572 ( .B(n4292), .A(n1055), .Z(n4321) );
  NAND U5573 ( .A(n1121), .B(n4289), .Z(n4292) );
  AND U5574 ( .A(n4322), .B(n4323), .Z(n4320) );
  NANDN U5575 ( .B(n1124), .A(n4289), .Z(n4323) );
  NAND U5576 ( .A(n4295), .B(\u_a23_mem/p_mem[109][7] ), .Z(n4322) );
  NANDN U5577 ( .B(n1125), .A(n4289), .Z(n4295) );
  NAND U5578 ( .A(n4324), .B(n4325), .Z(\u_a23_mem/n18540 ) );
  OR U5579 ( .A(n1011), .B(n4326), .Z(n4325) );
  AND U5580 ( .A(n4327), .B(n4328), .Z(n4324) );
  NANDN U5581 ( .B(n1131), .A(n4289), .Z(n4328) );
  NAND U5582 ( .A(n4329), .B(\u_a23_mem/p_mem[110][0] ), .Z(n4327) );
  NAND U5583 ( .A(n4330), .B(n4331), .Z(\u_a23_mem/n18539 ) );
  OR U5584 ( .A(n1019), .B(n4326), .Z(n4331) );
  AND U5585 ( .A(n4332), .B(n4333), .Z(n4330) );
  NANDN U5586 ( .B(n1137), .A(n4289), .Z(n4333) );
  NAND U5587 ( .A(n4329), .B(\u_a23_mem/p_mem[110][1] ), .Z(n4332) );
  NAND U5588 ( .A(n4334), .B(n4335), .Z(\u_a23_mem/n18538 ) );
  OR U5589 ( .A(n1025), .B(n4326), .Z(n4335) );
  AND U5590 ( .A(n4336), .B(n4337), .Z(n4334) );
  NANDN U5591 ( .B(n1142), .A(n4289), .Z(n4337) );
  NAND U5592 ( .A(n4329), .B(\u_a23_mem/p_mem[110][2] ), .Z(n4336) );
  NAND U5593 ( .A(n4338), .B(n4339), .Z(\u_a23_mem/n18537 ) );
  OR U5594 ( .A(n1031), .B(n4326), .Z(n4339) );
  AND U5595 ( .A(n4340), .B(n4341), .Z(n4338) );
  NANDN U5596 ( .B(n1147), .A(n4289), .Z(n4341) );
  NAND U5597 ( .A(n4329), .B(\u_a23_mem/p_mem[110][3] ), .Z(n4340) );
  NAND U5598 ( .A(n4342), .B(n4343), .Z(\u_a23_mem/n18536 ) );
  OR U5599 ( .A(n1037), .B(n4326), .Z(n4343) );
  AND U5600 ( .A(n4344), .B(n4345), .Z(n4342) );
  NANDN U5601 ( .B(n1152), .A(n4289), .Z(n4345) );
  NAND U5602 ( .A(n4329), .B(\u_a23_mem/p_mem[110][4] ), .Z(n4344) );
  NAND U5603 ( .A(n4346), .B(n4347), .Z(\u_a23_mem/n18535 ) );
  OR U5604 ( .A(n1043), .B(n4326), .Z(n4347) );
  AND U5605 ( .A(n4348), .B(n4349), .Z(n4346) );
  NANDN U5606 ( .B(n1157), .A(n4289), .Z(n4349) );
  NAND U5607 ( .A(n4329), .B(\u_a23_mem/p_mem[110][5] ), .Z(n4348) );
  NAND U5608 ( .A(n4350), .B(n4351), .Z(\u_a23_mem/n18534 ) );
  OR U5609 ( .A(n1049), .B(n4326), .Z(n4351) );
  AND U5610 ( .A(n4352), .B(n4353), .Z(n4350) );
  NANDN U5611 ( .B(n1162), .A(n4289), .Z(n4353) );
  NAND U5612 ( .A(n4329), .B(\u_a23_mem/p_mem[110][6] ), .Z(n4352) );
  NAND U5613 ( .A(n4354), .B(n4355), .Z(\u_a23_mem/n18533 ) );
  NANDN U5614 ( .B(n4326), .A(n1055), .Z(n4355) );
  NAND U5615 ( .A(n1165), .B(n4289), .Z(n4326) );
  AND U5616 ( .A(n4356), .B(n4357), .Z(n4354) );
  NANDN U5617 ( .B(n1168), .A(n4289), .Z(n4357) );
  NAND U5618 ( .A(n4329), .B(\u_a23_mem/p_mem[110][7] ), .Z(n4356) );
  NANDN U5619 ( .B(n1169), .A(n4289), .Z(n4329) );
  NAND U5620 ( .A(n4358), .B(n4359), .Z(\u_a23_mem/n18532 ) );
  OR U5621 ( .A(n1011), .B(n4360), .Z(n4359) );
  AND U5622 ( .A(n4361), .B(n4362), .Z(n4358) );
  NAND U5623 ( .A(n4363), .B(\u_a23_mem/p_mem[111][0] ), .Z(n4362) );
  NANDN U5624 ( .B(n1015), .A(n4289), .Z(n4361) );
  NAND U5625 ( .A(n4364), .B(n4365), .Z(\u_a23_mem/n18531 ) );
  OR U5626 ( .A(n1019), .B(n4360), .Z(n4365) );
  AND U5627 ( .A(n4366), .B(n4367), .Z(n4364) );
  NAND U5628 ( .A(n4363), .B(\u_a23_mem/p_mem[111][1] ), .Z(n4367) );
  NANDN U5629 ( .B(n1022), .A(n4289), .Z(n4366) );
  NAND U5630 ( .A(n4368), .B(n4369), .Z(\u_a23_mem/n18530 ) );
  OR U5631 ( .A(n1025), .B(n4360), .Z(n4369) );
  AND U5632 ( .A(n4370), .B(n4371), .Z(n4368) );
  NAND U5633 ( .A(n4363), .B(\u_a23_mem/p_mem[111][2] ), .Z(n4371) );
  NANDN U5634 ( .B(n1028), .A(n4289), .Z(n4370) );
  NAND U5635 ( .A(n4372), .B(n4373), .Z(\u_a23_mem/n18529 ) );
  OR U5636 ( .A(n1031), .B(n4360), .Z(n4373) );
  AND U5637 ( .A(n4374), .B(n4375), .Z(n4372) );
  NAND U5638 ( .A(n4363), .B(\u_a23_mem/p_mem[111][3] ), .Z(n4375) );
  NANDN U5639 ( .B(n1034), .A(n4289), .Z(n4374) );
  NAND U5640 ( .A(n4376), .B(n4377), .Z(\u_a23_mem/n18528 ) );
  OR U5641 ( .A(n1037), .B(n4360), .Z(n4377) );
  AND U5642 ( .A(n4378), .B(n4379), .Z(n4376) );
  NAND U5643 ( .A(n4363), .B(\u_a23_mem/p_mem[111][4] ), .Z(n4379) );
  NANDN U5644 ( .B(n1040), .A(n4289), .Z(n4378) );
  NAND U5645 ( .A(n4380), .B(n4381), .Z(\u_a23_mem/n18527 ) );
  OR U5646 ( .A(n1043), .B(n4360), .Z(n4381) );
  AND U5647 ( .A(n4382), .B(n4383), .Z(n4380) );
  NAND U5648 ( .A(n4363), .B(\u_a23_mem/p_mem[111][5] ), .Z(n4383) );
  NANDN U5649 ( .B(n1046), .A(n4289), .Z(n4382) );
  NAND U5650 ( .A(n4384), .B(n4385), .Z(\u_a23_mem/n18526 ) );
  OR U5651 ( .A(n1049), .B(n4360), .Z(n4385) );
  AND U5652 ( .A(n4386), .B(n4387), .Z(n4384) );
  NAND U5653 ( .A(n4363), .B(\u_a23_mem/p_mem[111][6] ), .Z(n4387) );
  NANDN U5654 ( .B(n1052), .A(n4289), .Z(n4386) );
  NAND U5655 ( .A(n4388), .B(n4389), .Z(\u_a23_mem/n18525 ) );
  NANDN U5656 ( .B(n4360), .A(n1055), .Z(n4389) );
  NAND U5657 ( .A(n1056), .B(n4289), .Z(n4360) );
  AND U5658 ( .A(n4390), .B(n4391), .Z(n4388) );
  NAND U5659 ( .A(n4363), .B(\u_a23_mem/p_mem[111][7] ), .Z(n4391) );
  NANDN U5660 ( .B(n1059), .A(n4289), .Z(n4363) );
  NAND U5661 ( .A(n1061), .B(n4289), .Z(n4390) );
  NOR U5662 ( .A(n1938), .B(n4023), .Z(n4289) );
  NAND U5663 ( .A(m_address[6]), .B(n4392), .Z(n4023) );
  AND U5664 ( .A(n1939), .B(m_address[5]), .Z(n4392) );
  NANDN U5665 ( .B(n4147), .A(n4393), .Z(n1938) );
  AND U5666 ( .A(n4148), .B(m_address[2]), .Z(n4393) );
  NAND U5667 ( .A(n4394), .B(n4395), .Z(\u_a23_mem/n18524 ) );
  NAND U5668 ( .A(n4396), .B(\u_a23_mem/p_mem[112][0] ), .Z(n4395) );
  OR U5669 ( .A(n1011), .B(n4397), .Z(n4394) );
  NAND U5670 ( .A(n4398), .B(n4399), .Z(\u_a23_mem/n18523 ) );
  NAND U5671 ( .A(n4396), .B(\u_a23_mem/p_mem[112][1] ), .Z(n4399) );
  OR U5672 ( .A(n1019), .B(n4397), .Z(n4398) );
  NAND U5673 ( .A(n4400), .B(n4401), .Z(\u_a23_mem/n18522 ) );
  NAND U5674 ( .A(n4396), .B(\u_a23_mem/p_mem[112][2] ), .Z(n4401) );
  OR U5675 ( .A(n1025), .B(n4397), .Z(n4400) );
  NAND U5676 ( .A(n4402), .B(n4403), .Z(\u_a23_mem/n18521 ) );
  NAND U5677 ( .A(n4396), .B(\u_a23_mem/p_mem[112][3] ), .Z(n4403) );
  OR U5678 ( .A(n1031), .B(n4397), .Z(n4402) );
  NAND U5679 ( .A(n4404), .B(n4405), .Z(\u_a23_mem/n18520 ) );
  NAND U5680 ( .A(n4396), .B(\u_a23_mem/p_mem[112][4] ), .Z(n4405) );
  OR U5681 ( .A(n1037), .B(n4397), .Z(n4404) );
  NAND U5682 ( .A(n4406), .B(n4407), .Z(\u_a23_mem/n18519 ) );
  NAND U5683 ( .A(n4396), .B(\u_a23_mem/p_mem[112][5] ), .Z(n4407) );
  OR U5684 ( .A(n1043), .B(n4397), .Z(n4406) );
  NAND U5685 ( .A(n4408), .B(n4409), .Z(\u_a23_mem/n18518 ) );
  NAND U5686 ( .A(n4396), .B(\u_a23_mem/p_mem[112][6] ), .Z(n4409) );
  OR U5687 ( .A(n1049), .B(n4397), .Z(n4408) );
  NAND U5688 ( .A(n4410), .B(n4411), .Z(\u_a23_mem/n18517 ) );
  NAND U5689 ( .A(n4396), .B(\u_a23_mem/p_mem[112][7] ), .Z(n4411) );
  NANDN U5690 ( .B(n1080), .A(n4412), .Z(n4396) );
  NANDN U5691 ( .B(n4397), .A(n1055), .Z(n4410) );
  NANDN U5692 ( .B(n2), .A(n4412), .Z(n4397) );
  NAND U5693 ( .A(n4413), .B(n4414), .Z(\u_a23_mem/n18516 ) );
  OR U5694 ( .A(n1011), .B(n4415), .Z(n4414) );
  AND U5695 ( .A(n4416), .B(n4417), .Z(n4413) );
  NANDN U5696 ( .B(n1087), .A(n4412), .Z(n4417) );
  NAND U5697 ( .A(n4418), .B(\u_a23_mem/p_mem[113][0] ), .Z(n4416) );
  NAND U5698 ( .A(n4419), .B(n4420), .Z(\u_a23_mem/n18515 ) );
  OR U5699 ( .A(n1019), .B(n4415), .Z(n4420) );
  AND U5700 ( .A(n4421), .B(n4422), .Z(n4419) );
  NANDN U5701 ( .B(n1093), .A(n4412), .Z(n4422) );
  NAND U5702 ( .A(n4418), .B(\u_a23_mem/p_mem[113][1] ), .Z(n4421) );
  NAND U5703 ( .A(n4423), .B(n4424), .Z(\u_a23_mem/n18514 ) );
  OR U5704 ( .A(n1025), .B(n4415), .Z(n4424) );
  AND U5705 ( .A(n4425), .B(n4426), .Z(n4423) );
  NANDN U5706 ( .B(n1098), .A(n4412), .Z(n4426) );
  NAND U5707 ( .A(n4418), .B(\u_a23_mem/p_mem[113][2] ), .Z(n4425) );
  NAND U5708 ( .A(n4427), .B(n4428), .Z(\u_a23_mem/n18513 ) );
  OR U5709 ( .A(n1031), .B(n4415), .Z(n4428) );
  AND U5710 ( .A(n4429), .B(n4430), .Z(n4427) );
  NANDN U5711 ( .B(n1103), .A(n4412), .Z(n4430) );
  NAND U5712 ( .A(n4418), .B(\u_a23_mem/p_mem[113][3] ), .Z(n4429) );
  NAND U5713 ( .A(n4431), .B(n4432), .Z(\u_a23_mem/n18512 ) );
  OR U5714 ( .A(n1037), .B(n4415), .Z(n4432) );
  AND U5715 ( .A(n4433), .B(n4434), .Z(n4431) );
  NANDN U5716 ( .B(n1108), .A(n4412), .Z(n4434) );
  NAND U5717 ( .A(n4418), .B(\u_a23_mem/p_mem[113][4] ), .Z(n4433) );
  NAND U5718 ( .A(n4435), .B(n4436), .Z(\u_a23_mem/n18511 ) );
  OR U5719 ( .A(n1043), .B(n4415), .Z(n4436) );
  AND U5720 ( .A(n4437), .B(n4438), .Z(n4435) );
  NANDN U5721 ( .B(n1113), .A(n4412), .Z(n4438) );
  NAND U5722 ( .A(n4418), .B(\u_a23_mem/p_mem[113][5] ), .Z(n4437) );
  NAND U5723 ( .A(n4439), .B(n4440), .Z(\u_a23_mem/n18510 ) );
  OR U5724 ( .A(n1049), .B(n4415), .Z(n4440) );
  AND U5725 ( .A(n4441), .B(n4442), .Z(n4439) );
  NANDN U5726 ( .B(n1118), .A(n4412), .Z(n4442) );
  NAND U5727 ( .A(n4418), .B(\u_a23_mem/p_mem[113][6] ), .Z(n4441) );
  NAND U5728 ( .A(n4443), .B(n4444), .Z(\u_a23_mem/n18509 ) );
  NANDN U5729 ( .B(n4415), .A(n1055), .Z(n4444) );
  NAND U5730 ( .A(n1121), .B(n4412), .Z(n4415) );
  AND U5731 ( .A(n4445), .B(n4446), .Z(n4443) );
  NANDN U5732 ( .B(n1124), .A(n4412), .Z(n4446) );
  NAND U5733 ( .A(n4418), .B(\u_a23_mem/p_mem[113][7] ), .Z(n4445) );
  NANDN U5734 ( .B(n1125), .A(n4412), .Z(n4418) );
  NAND U5735 ( .A(n4447), .B(n4448), .Z(\u_a23_mem/n18508 ) );
  OR U5736 ( .A(n1011), .B(n4449), .Z(n4448) );
  AND U5737 ( .A(n4450), .B(n4451), .Z(n4447) );
  NANDN U5738 ( .B(n1131), .A(n4412), .Z(n4451) );
  NAND U5739 ( .A(n4452), .B(\u_a23_mem/p_mem[114][0] ), .Z(n4450) );
  NAND U5740 ( .A(n4453), .B(n4454), .Z(\u_a23_mem/n18507 ) );
  OR U5741 ( .A(n1019), .B(n4449), .Z(n4454) );
  AND U5742 ( .A(n4455), .B(n4456), .Z(n4453) );
  NANDN U5743 ( .B(n1137), .A(n4412), .Z(n4456) );
  NAND U5744 ( .A(n4452), .B(\u_a23_mem/p_mem[114][1] ), .Z(n4455) );
  NAND U5745 ( .A(n4457), .B(n4458), .Z(\u_a23_mem/n18506 ) );
  OR U5746 ( .A(n1025), .B(n4449), .Z(n4458) );
  AND U5747 ( .A(n4459), .B(n4460), .Z(n4457) );
  NANDN U5748 ( .B(n1142), .A(n4412), .Z(n4460) );
  NAND U5749 ( .A(n4452), .B(\u_a23_mem/p_mem[114][2] ), .Z(n4459) );
  NAND U5750 ( .A(n4461), .B(n4462), .Z(\u_a23_mem/n18505 ) );
  OR U5751 ( .A(n1031), .B(n4449), .Z(n4462) );
  AND U5752 ( .A(n4463), .B(n4464), .Z(n4461) );
  NANDN U5753 ( .B(n1147), .A(n4412), .Z(n4464) );
  NAND U5754 ( .A(n4452), .B(\u_a23_mem/p_mem[114][3] ), .Z(n4463) );
  NAND U5755 ( .A(n4465), .B(n4466), .Z(\u_a23_mem/n18504 ) );
  OR U5756 ( .A(n1037), .B(n4449), .Z(n4466) );
  AND U5757 ( .A(n4467), .B(n4468), .Z(n4465) );
  NANDN U5758 ( .B(n1152), .A(n4412), .Z(n4468) );
  NAND U5759 ( .A(n4452), .B(\u_a23_mem/p_mem[114][4] ), .Z(n4467) );
  NAND U5760 ( .A(n4469), .B(n4470), .Z(\u_a23_mem/n18503 ) );
  OR U5761 ( .A(n1043), .B(n4449), .Z(n4470) );
  AND U5762 ( .A(n4471), .B(n4472), .Z(n4469) );
  NANDN U5763 ( .B(n1157), .A(n4412), .Z(n4472) );
  NAND U5764 ( .A(n4452), .B(\u_a23_mem/p_mem[114][5] ), .Z(n4471) );
  NAND U5765 ( .A(n4473), .B(n4474), .Z(\u_a23_mem/n18502 ) );
  OR U5766 ( .A(n1049), .B(n4449), .Z(n4474) );
  AND U5767 ( .A(n4475), .B(n4476), .Z(n4473) );
  NANDN U5768 ( .B(n1162), .A(n4412), .Z(n4476) );
  NAND U5769 ( .A(n4452), .B(\u_a23_mem/p_mem[114][6] ), .Z(n4475) );
  NAND U5770 ( .A(n4477), .B(n4478), .Z(\u_a23_mem/n18501 ) );
  NANDN U5771 ( .B(n4449), .A(n1055), .Z(n4478) );
  NAND U5772 ( .A(n1165), .B(n4412), .Z(n4449) );
  AND U5773 ( .A(n4479), .B(n4480), .Z(n4477) );
  NANDN U5774 ( .B(n1168), .A(n4412), .Z(n4480) );
  NAND U5775 ( .A(n4452), .B(\u_a23_mem/p_mem[114][7] ), .Z(n4479) );
  NANDN U5776 ( .B(n1169), .A(n4412), .Z(n4452) );
  NAND U5777 ( .A(n4481), .B(n4482), .Z(\u_a23_mem/n18500 ) );
  OR U5778 ( .A(n1011), .B(n4483), .Z(n4482) );
  AND U5779 ( .A(n4484), .B(n4485), .Z(n4481) );
  NAND U5780 ( .A(n4486), .B(\u_a23_mem/p_mem[115][0] ), .Z(n4485) );
  NANDN U5781 ( .B(n1015), .A(n4412), .Z(n4484) );
  NAND U5782 ( .A(n4487), .B(n4488), .Z(\u_a23_mem/n18499 ) );
  OR U5783 ( .A(n1019), .B(n4483), .Z(n4488) );
  AND U5784 ( .A(n4489), .B(n4490), .Z(n4487) );
  NAND U5785 ( .A(n4486), .B(\u_a23_mem/p_mem[115][1] ), .Z(n4490) );
  NANDN U5786 ( .B(n1022), .A(n4412), .Z(n4489) );
  NAND U5787 ( .A(n4491), .B(n4492), .Z(\u_a23_mem/n18498 ) );
  OR U5788 ( .A(n1025), .B(n4483), .Z(n4492) );
  AND U5789 ( .A(n4493), .B(n4494), .Z(n4491) );
  NAND U5790 ( .A(n4486), .B(\u_a23_mem/p_mem[115][2] ), .Z(n4494) );
  NANDN U5791 ( .B(n1028), .A(n4412), .Z(n4493) );
  NAND U5792 ( .A(n4495), .B(n4496), .Z(\u_a23_mem/n18497 ) );
  OR U5793 ( .A(n1031), .B(n4483), .Z(n4496) );
  AND U5794 ( .A(n4497), .B(n4498), .Z(n4495) );
  NAND U5795 ( .A(n4486), .B(\u_a23_mem/p_mem[115][3] ), .Z(n4498) );
  NANDN U5796 ( .B(n1034), .A(n4412), .Z(n4497) );
  NAND U5797 ( .A(n4499), .B(n4500), .Z(\u_a23_mem/n18496 ) );
  OR U5798 ( .A(n1037), .B(n4483), .Z(n4500) );
  AND U5799 ( .A(n4501), .B(n4502), .Z(n4499) );
  NAND U5800 ( .A(n4486), .B(\u_a23_mem/p_mem[115][4] ), .Z(n4502) );
  NANDN U5801 ( .B(n1040), .A(n4412), .Z(n4501) );
  NAND U5802 ( .A(n4503), .B(n4504), .Z(\u_a23_mem/n18495 ) );
  OR U5803 ( .A(n1043), .B(n4483), .Z(n4504) );
  AND U5804 ( .A(n4505), .B(n4506), .Z(n4503) );
  NAND U5805 ( .A(n4486), .B(\u_a23_mem/p_mem[115][5] ), .Z(n4506) );
  NANDN U5806 ( .B(n1046), .A(n4412), .Z(n4505) );
  NAND U5807 ( .A(n4507), .B(n4508), .Z(\u_a23_mem/n18494 ) );
  OR U5808 ( .A(n1049), .B(n4483), .Z(n4508) );
  AND U5809 ( .A(n4509), .B(n4510), .Z(n4507) );
  NAND U5810 ( .A(n4486), .B(\u_a23_mem/p_mem[115][6] ), .Z(n4510) );
  NANDN U5811 ( .B(n1052), .A(n4412), .Z(n4509) );
  NAND U5812 ( .A(n4511), .B(n4512), .Z(\u_a23_mem/n18493 ) );
  NANDN U5813 ( .B(n4483), .A(n1055), .Z(n4512) );
  NAND U5814 ( .A(n1056), .B(n4412), .Z(n4483) );
  AND U5815 ( .A(n4513), .B(n4514), .Z(n4511) );
  NAND U5816 ( .A(n4486), .B(\u_a23_mem/p_mem[115][7] ), .Z(n4514) );
  NANDN U5817 ( .B(n1059), .A(n4412), .Z(n4486) );
  NAND U5818 ( .A(n1061), .B(n4412), .Z(n4513) );
  AND U5819 ( .A(n4515), .B(n4516), .Z(n4412) );
  AND U5820 ( .A(n1571), .B(m_address[4]), .Z(n4516) );
  ANDN U5821 ( .A(n4517), .B(n4518), .Z(n1571) );
  NAND U5822 ( .A(n4519), .B(n4520), .Z(\u_a23_mem/n18492 ) );
  NAND U5823 ( .A(n4521), .B(\u_a23_mem/p_mem[116][0] ), .Z(n4520) );
  OR U5824 ( .A(n1011), .B(n4522), .Z(n4519) );
  NAND U5825 ( .A(n4523), .B(n4524), .Z(\u_a23_mem/n18491 ) );
  NAND U5826 ( .A(n4521), .B(\u_a23_mem/p_mem[116][1] ), .Z(n4524) );
  OR U5827 ( .A(n1019), .B(n4522), .Z(n4523) );
  NAND U5828 ( .A(n4525), .B(n4526), .Z(\u_a23_mem/n18490 ) );
  NAND U5829 ( .A(n4521), .B(\u_a23_mem/p_mem[116][2] ), .Z(n4526) );
  OR U5830 ( .A(n1025), .B(n4522), .Z(n4525) );
  NAND U5831 ( .A(n4527), .B(n4528), .Z(\u_a23_mem/n18489 ) );
  NAND U5832 ( .A(n4521), .B(\u_a23_mem/p_mem[116][3] ), .Z(n4528) );
  OR U5833 ( .A(n1031), .B(n4522), .Z(n4527) );
  NAND U5834 ( .A(n4529), .B(n4530), .Z(\u_a23_mem/n18488 ) );
  NAND U5835 ( .A(n4521), .B(\u_a23_mem/p_mem[116][4] ), .Z(n4530) );
  OR U5836 ( .A(n1037), .B(n4522), .Z(n4529) );
  NAND U5837 ( .A(n4531), .B(n4532), .Z(\u_a23_mem/n18487 ) );
  NAND U5838 ( .A(n4521), .B(\u_a23_mem/p_mem[116][5] ), .Z(n4532) );
  OR U5839 ( .A(n1043), .B(n4522), .Z(n4531) );
  NAND U5840 ( .A(n4533), .B(n4534), .Z(\u_a23_mem/n18486 ) );
  NAND U5841 ( .A(n4521), .B(\u_a23_mem/p_mem[116][6] ), .Z(n4534) );
  OR U5842 ( .A(n1049), .B(n4522), .Z(n4533) );
  NAND U5843 ( .A(n4535), .B(n4536), .Z(\u_a23_mem/n18485 ) );
  NAND U5844 ( .A(n4521), .B(\u_a23_mem/p_mem[116][7] ), .Z(n4536) );
  NANDN U5845 ( .B(n1080), .A(n4537), .Z(n4521) );
  NANDN U5846 ( .B(n4522), .A(n1055), .Z(n4535) );
  NANDN U5847 ( .B(n2), .A(n4537), .Z(n4522) );
  NAND U5848 ( .A(n4538), .B(n4539), .Z(\u_a23_mem/n18484 ) );
  OR U5849 ( .A(n1011), .B(n4540), .Z(n4539) );
  AND U5850 ( .A(n4541), .B(n4542), .Z(n4538) );
  NANDN U5851 ( .B(n1087), .A(n4537), .Z(n4542) );
  NAND U5852 ( .A(n4543), .B(\u_a23_mem/p_mem[117][0] ), .Z(n4541) );
  NAND U5853 ( .A(n4544), .B(n4545), .Z(\u_a23_mem/n18483 ) );
  OR U5854 ( .A(n1019), .B(n4540), .Z(n4545) );
  AND U5855 ( .A(n4546), .B(n4547), .Z(n4544) );
  NANDN U5856 ( .B(n1093), .A(n4537), .Z(n4547) );
  NAND U5857 ( .A(n4543), .B(\u_a23_mem/p_mem[117][1] ), .Z(n4546) );
  NAND U5858 ( .A(n4548), .B(n4549), .Z(\u_a23_mem/n18482 ) );
  OR U5859 ( .A(n1025), .B(n4540), .Z(n4549) );
  AND U5860 ( .A(n4550), .B(n4551), .Z(n4548) );
  NANDN U5861 ( .B(n1098), .A(n4537), .Z(n4551) );
  NAND U5862 ( .A(n4543), .B(\u_a23_mem/p_mem[117][2] ), .Z(n4550) );
  NAND U5863 ( .A(n4552), .B(n4553), .Z(\u_a23_mem/n18481 ) );
  OR U5864 ( .A(n1031), .B(n4540), .Z(n4553) );
  AND U5865 ( .A(n4554), .B(n4555), .Z(n4552) );
  NANDN U5866 ( .B(n1103), .A(n4537), .Z(n4555) );
  NAND U5867 ( .A(n4543), .B(\u_a23_mem/p_mem[117][3] ), .Z(n4554) );
  NAND U5868 ( .A(n4556), .B(n4557), .Z(\u_a23_mem/n18480 ) );
  OR U5869 ( .A(n1037), .B(n4540), .Z(n4557) );
  AND U5870 ( .A(n4558), .B(n4559), .Z(n4556) );
  NANDN U5871 ( .B(n1108), .A(n4537), .Z(n4559) );
  NAND U5872 ( .A(n4543), .B(\u_a23_mem/p_mem[117][4] ), .Z(n4558) );
  NAND U5873 ( .A(n4560), .B(n4561), .Z(\u_a23_mem/n18479 ) );
  OR U5874 ( .A(n1043), .B(n4540), .Z(n4561) );
  AND U5875 ( .A(n4562), .B(n4563), .Z(n4560) );
  NANDN U5876 ( .B(n1113), .A(n4537), .Z(n4563) );
  NAND U5877 ( .A(n4543), .B(\u_a23_mem/p_mem[117][5] ), .Z(n4562) );
  NAND U5878 ( .A(n4564), .B(n4565), .Z(\u_a23_mem/n18478 ) );
  OR U5879 ( .A(n1049), .B(n4540), .Z(n4565) );
  AND U5880 ( .A(n4566), .B(n4567), .Z(n4564) );
  NANDN U5881 ( .B(n1118), .A(n4537), .Z(n4567) );
  NAND U5882 ( .A(n4543), .B(\u_a23_mem/p_mem[117][6] ), .Z(n4566) );
  NAND U5883 ( .A(n4568), .B(n4569), .Z(\u_a23_mem/n18477 ) );
  NANDN U5884 ( .B(n4540), .A(n1055), .Z(n4569) );
  NAND U5885 ( .A(n1121), .B(n4537), .Z(n4540) );
  AND U5886 ( .A(n4570), .B(n4571), .Z(n4568) );
  NANDN U5887 ( .B(n1124), .A(n4537), .Z(n4571) );
  NAND U5888 ( .A(n4543), .B(\u_a23_mem/p_mem[117][7] ), .Z(n4570) );
  NANDN U5889 ( .B(n1125), .A(n4537), .Z(n4543) );
  NAND U5890 ( .A(n4572), .B(n4573), .Z(\u_a23_mem/n18476 ) );
  OR U5891 ( .A(n1011), .B(n4574), .Z(n4573) );
  AND U5892 ( .A(n4575), .B(n4576), .Z(n4572) );
  NANDN U5893 ( .B(n1131), .A(n4537), .Z(n4576) );
  NAND U5894 ( .A(n4577), .B(\u_a23_mem/p_mem[118][0] ), .Z(n4575) );
  NAND U5895 ( .A(n4578), .B(n4579), .Z(\u_a23_mem/n18475 ) );
  OR U5896 ( .A(n1019), .B(n4574), .Z(n4579) );
  AND U5897 ( .A(n4580), .B(n4581), .Z(n4578) );
  NANDN U5898 ( .B(n1137), .A(n4537), .Z(n4581) );
  NAND U5899 ( .A(n4577), .B(\u_a23_mem/p_mem[118][1] ), .Z(n4580) );
  NAND U5900 ( .A(n4582), .B(n4583), .Z(\u_a23_mem/n18474 ) );
  OR U5901 ( .A(n1025), .B(n4574), .Z(n4583) );
  AND U5902 ( .A(n4584), .B(n4585), .Z(n4582) );
  NANDN U5903 ( .B(n1142), .A(n4537), .Z(n4585) );
  NAND U5904 ( .A(n4577), .B(\u_a23_mem/p_mem[118][2] ), .Z(n4584) );
  NAND U5905 ( .A(n4586), .B(n4587), .Z(\u_a23_mem/n18473 ) );
  OR U5906 ( .A(n1031), .B(n4574), .Z(n4587) );
  AND U5907 ( .A(n4588), .B(n4589), .Z(n4586) );
  NANDN U5908 ( .B(n1147), .A(n4537), .Z(n4589) );
  NAND U5909 ( .A(n4577), .B(\u_a23_mem/p_mem[118][3] ), .Z(n4588) );
  NAND U5910 ( .A(n4590), .B(n4591), .Z(\u_a23_mem/n18472 ) );
  OR U5911 ( .A(n1037), .B(n4574), .Z(n4591) );
  AND U5912 ( .A(n4592), .B(n4593), .Z(n4590) );
  NANDN U5913 ( .B(n1152), .A(n4537), .Z(n4593) );
  NAND U5914 ( .A(n4577), .B(\u_a23_mem/p_mem[118][4] ), .Z(n4592) );
  NAND U5915 ( .A(n4594), .B(n4595), .Z(\u_a23_mem/n18471 ) );
  OR U5916 ( .A(n1043), .B(n4574), .Z(n4595) );
  AND U5917 ( .A(n4596), .B(n4597), .Z(n4594) );
  NANDN U5918 ( .B(n1157), .A(n4537), .Z(n4597) );
  NAND U5919 ( .A(n4577), .B(\u_a23_mem/p_mem[118][5] ), .Z(n4596) );
  NAND U5920 ( .A(n4598), .B(n4599), .Z(\u_a23_mem/n18470 ) );
  OR U5921 ( .A(n1049), .B(n4574), .Z(n4599) );
  AND U5922 ( .A(n4600), .B(n4601), .Z(n4598) );
  NANDN U5923 ( .B(n1162), .A(n4537), .Z(n4601) );
  NAND U5924 ( .A(n4577), .B(\u_a23_mem/p_mem[118][6] ), .Z(n4600) );
  NAND U5925 ( .A(n4602), .B(n4603), .Z(\u_a23_mem/n18469 ) );
  NANDN U5926 ( .B(n4574), .A(n1055), .Z(n4603) );
  NAND U5927 ( .A(n1165), .B(n4537), .Z(n4574) );
  AND U5928 ( .A(n4604), .B(n4605), .Z(n4602) );
  NANDN U5929 ( .B(n1168), .A(n4537), .Z(n4605) );
  NAND U5930 ( .A(n4577), .B(\u_a23_mem/p_mem[118][7] ), .Z(n4604) );
  NANDN U5931 ( .B(n1169), .A(n4537), .Z(n4577) );
  NAND U5932 ( .A(n4606), .B(n4607), .Z(\u_a23_mem/n18468 ) );
  OR U5933 ( .A(n1011), .B(n4608), .Z(n4607) );
  AND U5934 ( .A(n4609), .B(n4610), .Z(n4606) );
  NAND U5935 ( .A(n4611), .B(\u_a23_mem/p_mem[119][0] ), .Z(n4610) );
  NANDN U5936 ( .B(n1015), .A(n4537), .Z(n4609) );
  NAND U5937 ( .A(n4612), .B(n4613), .Z(\u_a23_mem/n18467 ) );
  OR U5938 ( .A(n1019), .B(n4608), .Z(n4613) );
  AND U5939 ( .A(n4614), .B(n4615), .Z(n4612) );
  NAND U5940 ( .A(n4611), .B(\u_a23_mem/p_mem[119][1] ), .Z(n4615) );
  NANDN U5941 ( .B(n1022), .A(n4537), .Z(n4614) );
  NAND U5942 ( .A(n4616), .B(n4617), .Z(\u_a23_mem/n18466 ) );
  OR U5943 ( .A(n1025), .B(n4608), .Z(n4617) );
  AND U5944 ( .A(n4618), .B(n4619), .Z(n4616) );
  NAND U5945 ( .A(n4611), .B(\u_a23_mem/p_mem[119][2] ), .Z(n4619) );
  NANDN U5946 ( .B(n1028), .A(n4537), .Z(n4618) );
  NAND U5947 ( .A(n4620), .B(n4621), .Z(\u_a23_mem/n18465 ) );
  OR U5948 ( .A(n1031), .B(n4608), .Z(n4621) );
  AND U5949 ( .A(n4622), .B(n4623), .Z(n4620) );
  NAND U5950 ( .A(n4611), .B(\u_a23_mem/p_mem[119][3] ), .Z(n4623) );
  NANDN U5951 ( .B(n1034), .A(n4537), .Z(n4622) );
  NAND U5952 ( .A(n4624), .B(n4625), .Z(\u_a23_mem/n18464 ) );
  OR U5953 ( .A(n1037), .B(n4608), .Z(n4625) );
  AND U5954 ( .A(n4626), .B(n4627), .Z(n4624) );
  NAND U5955 ( .A(n4611), .B(\u_a23_mem/p_mem[119][4] ), .Z(n4627) );
  NANDN U5956 ( .B(n1040), .A(n4537), .Z(n4626) );
  NAND U5957 ( .A(n4628), .B(n4629), .Z(\u_a23_mem/n18463 ) );
  OR U5958 ( .A(n1043), .B(n4608), .Z(n4629) );
  AND U5959 ( .A(n4630), .B(n4631), .Z(n4628) );
  NAND U5960 ( .A(n4611), .B(\u_a23_mem/p_mem[119][5] ), .Z(n4631) );
  NANDN U5961 ( .B(n1046), .A(n4537), .Z(n4630) );
  NAND U5962 ( .A(n4632), .B(n4633), .Z(\u_a23_mem/n18462 ) );
  OR U5963 ( .A(n1049), .B(n4608), .Z(n4633) );
  AND U5964 ( .A(n4634), .B(n4635), .Z(n4632) );
  NAND U5965 ( .A(n4611), .B(\u_a23_mem/p_mem[119][6] ), .Z(n4635) );
  NANDN U5966 ( .B(n1052), .A(n4537), .Z(n4634) );
  NAND U5967 ( .A(n4636), .B(n4637), .Z(\u_a23_mem/n18461 ) );
  NANDN U5968 ( .B(n4608), .A(n1055), .Z(n4637) );
  NAND U5969 ( .A(n1056), .B(n4537), .Z(n4608) );
  AND U5970 ( .A(n4638), .B(n4639), .Z(n4636) );
  NAND U5971 ( .A(n4611), .B(\u_a23_mem/p_mem[119][7] ), .Z(n4639) );
  NANDN U5972 ( .B(n1059), .A(n4537), .Z(n4611) );
  NAND U5973 ( .A(n1061), .B(n4537), .Z(n4638) );
  ANDN U5974 ( .A(n1204), .B(n4640), .Z(n4537) );
  AND U5975 ( .A(n4147), .B(m_address[2]), .Z(n1204) );
  NAND U5976 ( .A(n4641), .B(n4642), .Z(\u_a23_mem/n18460 ) );
  NAND U5977 ( .A(n4643), .B(\u_a23_mem/p_mem[120][0] ), .Z(n4642) );
  OR U5978 ( .A(n1011), .B(n4644), .Z(n4641) );
  NAND U5979 ( .A(n4645), .B(n4646), .Z(\u_a23_mem/n18459 ) );
  NAND U5980 ( .A(n4643), .B(\u_a23_mem/p_mem[120][1] ), .Z(n4646) );
  OR U5981 ( .A(n1019), .B(n4644), .Z(n4645) );
  NAND U5982 ( .A(n4647), .B(n4648), .Z(\u_a23_mem/n18458 ) );
  NAND U5983 ( .A(n4643), .B(\u_a23_mem/p_mem[120][2] ), .Z(n4648) );
  OR U5984 ( .A(n1025), .B(n4644), .Z(n4647) );
  NAND U5985 ( .A(n4649), .B(n4650), .Z(\u_a23_mem/n18457 ) );
  NAND U5986 ( .A(n4643), .B(\u_a23_mem/p_mem[120][3] ), .Z(n4650) );
  OR U5987 ( .A(n1031), .B(n4644), .Z(n4649) );
  NAND U5988 ( .A(n4651), .B(n4652), .Z(\u_a23_mem/n18456 ) );
  NAND U5989 ( .A(n4643), .B(\u_a23_mem/p_mem[120][4] ), .Z(n4652) );
  OR U5990 ( .A(n1037), .B(n4644), .Z(n4651) );
  NAND U5991 ( .A(n4653), .B(n4654), .Z(\u_a23_mem/n18455 ) );
  NAND U5992 ( .A(n4643), .B(\u_a23_mem/p_mem[120][5] ), .Z(n4654) );
  OR U5993 ( .A(n1043), .B(n4644), .Z(n4653) );
  NAND U5994 ( .A(n4655), .B(n4656), .Z(\u_a23_mem/n18454 ) );
  NAND U5995 ( .A(n4643), .B(\u_a23_mem/p_mem[120][6] ), .Z(n4656) );
  OR U5996 ( .A(n1049), .B(n4644), .Z(n4655) );
  NAND U5997 ( .A(n4657), .B(n4658), .Z(\u_a23_mem/n18453 ) );
  NAND U5998 ( .A(n4643), .B(\u_a23_mem/p_mem[120][7] ), .Z(n4658) );
  NANDN U5999 ( .B(n1080), .A(n4659), .Z(n4643) );
  NANDN U6000 ( .B(n4644), .A(n1055), .Z(n4657) );
  NANDN U6001 ( .B(n2), .A(n4659), .Z(n4644) );
  NAND U6002 ( .A(n4660), .B(n4661), .Z(\u_a23_mem/n18452 ) );
  OR U6003 ( .A(n1011), .B(n4662), .Z(n4661) );
  AND U6004 ( .A(n4663), .B(n4664), .Z(n4660) );
  NANDN U6005 ( .B(n1087), .A(n4659), .Z(n4664) );
  NAND U6006 ( .A(n4665), .B(\u_a23_mem/p_mem[121][0] ), .Z(n4663) );
  NAND U6007 ( .A(n4666), .B(n4667), .Z(\u_a23_mem/n18451 ) );
  OR U6008 ( .A(n1019), .B(n4662), .Z(n4667) );
  AND U6009 ( .A(n4668), .B(n4669), .Z(n4666) );
  NANDN U6010 ( .B(n1093), .A(n4659), .Z(n4669) );
  NAND U6011 ( .A(n4665), .B(\u_a23_mem/p_mem[121][1] ), .Z(n4668) );
  NAND U6012 ( .A(n4670), .B(n4671), .Z(\u_a23_mem/n18450 ) );
  OR U6013 ( .A(n1025), .B(n4662), .Z(n4671) );
  AND U6014 ( .A(n4672), .B(n4673), .Z(n4670) );
  NANDN U6015 ( .B(n1098), .A(n4659), .Z(n4673) );
  NAND U6016 ( .A(n4665), .B(\u_a23_mem/p_mem[121][2] ), .Z(n4672) );
  NAND U6017 ( .A(n4674), .B(n4675), .Z(\u_a23_mem/n18449 ) );
  OR U6018 ( .A(n1031), .B(n4662), .Z(n4675) );
  AND U6019 ( .A(n4676), .B(n4677), .Z(n4674) );
  NANDN U6020 ( .B(n1103), .A(n4659), .Z(n4677) );
  NAND U6021 ( .A(n4665), .B(\u_a23_mem/p_mem[121][3] ), .Z(n4676) );
  NAND U6022 ( .A(n4678), .B(n4679), .Z(\u_a23_mem/n18448 ) );
  OR U6023 ( .A(n1037), .B(n4662), .Z(n4679) );
  AND U6024 ( .A(n4680), .B(n4681), .Z(n4678) );
  NANDN U6025 ( .B(n1108), .A(n4659), .Z(n4681) );
  NAND U6026 ( .A(n4665), .B(\u_a23_mem/p_mem[121][4] ), .Z(n4680) );
  NAND U6027 ( .A(n4682), .B(n4683), .Z(\u_a23_mem/n18447 ) );
  OR U6028 ( .A(n1043), .B(n4662), .Z(n4683) );
  AND U6029 ( .A(n4684), .B(n4685), .Z(n4682) );
  NANDN U6030 ( .B(n1113), .A(n4659), .Z(n4685) );
  NAND U6031 ( .A(n4665), .B(\u_a23_mem/p_mem[121][5] ), .Z(n4684) );
  NAND U6032 ( .A(n4686), .B(n4687), .Z(\u_a23_mem/n18446 ) );
  OR U6033 ( .A(n1049), .B(n4662), .Z(n4687) );
  AND U6034 ( .A(n4688), .B(n4689), .Z(n4686) );
  NANDN U6035 ( .B(n1118), .A(n4659), .Z(n4689) );
  NAND U6036 ( .A(n4665), .B(\u_a23_mem/p_mem[121][6] ), .Z(n4688) );
  NAND U6037 ( .A(n4690), .B(n4691), .Z(\u_a23_mem/n18445 ) );
  NANDN U6038 ( .B(n4662), .A(n1055), .Z(n4691) );
  NAND U6039 ( .A(n1121), .B(n4659), .Z(n4662) );
  AND U6040 ( .A(n4692), .B(n4693), .Z(n4690) );
  NANDN U6041 ( .B(n1124), .A(n4659), .Z(n4693) );
  NAND U6042 ( .A(n4665), .B(\u_a23_mem/p_mem[121][7] ), .Z(n4692) );
  NANDN U6043 ( .B(n1125), .A(n4659), .Z(n4665) );
  NAND U6044 ( .A(n4694), .B(n4695), .Z(\u_a23_mem/n18444 ) );
  OR U6045 ( .A(n1011), .B(n4696), .Z(n4695) );
  AND U6046 ( .A(n4697), .B(n4698), .Z(n4694) );
  NANDN U6047 ( .B(n1131), .A(n4659), .Z(n4698) );
  NAND U6048 ( .A(n4699), .B(\u_a23_mem/p_mem[122][0] ), .Z(n4697) );
  NAND U6049 ( .A(n4700), .B(n4701), .Z(\u_a23_mem/n18443 ) );
  OR U6050 ( .A(n1019), .B(n4696), .Z(n4701) );
  AND U6051 ( .A(n4702), .B(n4703), .Z(n4700) );
  NANDN U6052 ( .B(n1137), .A(n4659), .Z(n4703) );
  NAND U6053 ( .A(n4699), .B(\u_a23_mem/p_mem[122][1] ), .Z(n4702) );
  NAND U6054 ( .A(n4704), .B(n4705), .Z(\u_a23_mem/n18442 ) );
  OR U6055 ( .A(n1025), .B(n4696), .Z(n4705) );
  AND U6056 ( .A(n4706), .B(n4707), .Z(n4704) );
  NANDN U6057 ( .B(n1142), .A(n4659), .Z(n4707) );
  NAND U6058 ( .A(n4699), .B(\u_a23_mem/p_mem[122][2] ), .Z(n4706) );
  NAND U6059 ( .A(n4708), .B(n4709), .Z(\u_a23_mem/n18441 ) );
  OR U6060 ( .A(n1031), .B(n4696), .Z(n4709) );
  AND U6061 ( .A(n4710), .B(n4711), .Z(n4708) );
  NANDN U6062 ( .B(n1147), .A(n4659), .Z(n4711) );
  NAND U6063 ( .A(n4699), .B(\u_a23_mem/p_mem[122][3] ), .Z(n4710) );
  NAND U6064 ( .A(n4712), .B(n4713), .Z(\u_a23_mem/n18440 ) );
  OR U6065 ( .A(n1037), .B(n4696), .Z(n4713) );
  AND U6066 ( .A(n4714), .B(n4715), .Z(n4712) );
  NANDN U6067 ( .B(n1152), .A(n4659), .Z(n4715) );
  NAND U6068 ( .A(n4699), .B(\u_a23_mem/p_mem[122][4] ), .Z(n4714) );
  NAND U6069 ( .A(n4716), .B(n4717), .Z(\u_a23_mem/n18439 ) );
  OR U6070 ( .A(n1043), .B(n4696), .Z(n4717) );
  AND U6071 ( .A(n4718), .B(n4719), .Z(n4716) );
  NANDN U6072 ( .B(n1157), .A(n4659), .Z(n4719) );
  NAND U6073 ( .A(n4699), .B(\u_a23_mem/p_mem[122][5] ), .Z(n4718) );
  NAND U6074 ( .A(n4720), .B(n4721), .Z(\u_a23_mem/n18438 ) );
  OR U6075 ( .A(n1049), .B(n4696), .Z(n4721) );
  AND U6076 ( .A(n4722), .B(n4723), .Z(n4720) );
  NANDN U6077 ( .B(n1162), .A(n4659), .Z(n4723) );
  NAND U6078 ( .A(n4699), .B(\u_a23_mem/p_mem[122][6] ), .Z(n4722) );
  NAND U6079 ( .A(n4724), .B(n4725), .Z(\u_a23_mem/n18437 ) );
  NANDN U6080 ( .B(n4696), .A(n1055), .Z(n4725) );
  NAND U6081 ( .A(n1165), .B(n4659), .Z(n4696) );
  AND U6082 ( .A(n4726), .B(n4727), .Z(n4724) );
  NANDN U6083 ( .B(n1168), .A(n4659), .Z(n4727) );
  NAND U6084 ( .A(n4699), .B(\u_a23_mem/p_mem[122][7] ), .Z(n4726) );
  NANDN U6085 ( .B(n1169), .A(n4659), .Z(n4699) );
  NAND U6086 ( .A(n4728), .B(n4729), .Z(\u_a23_mem/n18436 ) );
  OR U6087 ( .A(n1011), .B(n4730), .Z(n4729) );
  AND U6088 ( .A(n4731), .B(n4732), .Z(n4728) );
  NAND U6089 ( .A(n4733), .B(\u_a23_mem/p_mem[123][0] ), .Z(n4732) );
  NANDN U6090 ( .B(n1015), .A(n4659), .Z(n4731) );
  NAND U6091 ( .A(n4734), .B(n4735), .Z(\u_a23_mem/n18435 ) );
  OR U6092 ( .A(n1019), .B(n4730), .Z(n4735) );
  AND U6093 ( .A(n4736), .B(n4737), .Z(n4734) );
  NAND U6094 ( .A(n4733), .B(\u_a23_mem/p_mem[123][1] ), .Z(n4737) );
  NANDN U6095 ( .B(n1022), .A(n4659), .Z(n4736) );
  NAND U6096 ( .A(n4738), .B(n4739), .Z(\u_a23_mem/n18434 ) );
  OR U6097 ( .A(n1025), .B(n4730), .Z(n4739) );
  AND U6098 ( .A(n4740), .B(n4741), .Z(n4738) );
  NAND U6099 ( .A(n4733), .B(\u_a23_mem/p_mem[123][2] ), .Z(n4741) );
  NANDN U6100 ( .B(n1028), .A(n4659), .Z(n4740) );
  NAND U6101 ( .A(n4742), .B(n4743), .Z(\u_a23_mem/n18433 ) );
  OR U6102 ( .A(n1031), .B(n4730), .Z(n4743) );
  AND U6103 ( .A(n4744), .B(n4745), .Z(n4742) );
  NAND U6104 ( .A(n4733), .B(\u_a23_mem/p_mem[123][3] ), .Z(n4745) );
  NANDN U6105 ( .B(n1034), .A(n4659), .Z(n4744) );
  NAND U6106 ( .A(n4746), .B(n4747), .Z(\u_a23_mem/n18432 ) );
  OR U6107 ( .A(n1037), .B(n4730), .Z(n4747) );
  AND U6108 ( .A(n4748), .B(n4749), .Z(n4746) );
  NAND U6109 ( .A(n4733), .B(\u_a23_mem/p_mem[123][4] ), .Z(n4749) );
  NANDN U6110 ( .B(n1040), .A(n4659), .Z(n4748) );
  NAND U6111 ( .A(n4750), .B(n4751), .Z(\u_a23_mem/n18431 ) );
  OR U6112 ( .A(n1043), .B(n4730), .Z(n4751) );
  AND U6113 ( .A(n4752), .B(n4753), .Z(n4750) );
  NAND U6114 ( .A(n4733), .B(\u_a23_mem/p_mem[123][5] ), .Z(n4753) );
  NANDN U6115 ( .B(n1046), .A(n4659), .Z(n4752) );
  NAND U6116 ( .A(n4754), .B(n4755), .Z(\u_a23_mem/n18430 ) );
  OR U6117 ( .A(n1049), .B(n4730), .Z(n4755) );
  AND U6118 ( .A(n4756), .B(n4757), .Z(n4754) );
  NAND U6119 ( .A(n4733), .B(\u_a23_mem/p_mem[123][6] ), .Z(n4757) );
  NANDN U6120 ( .B(n1052), .A(n4659), .Z(n4756) );
  NAND U6121 ( .A(n4758), .B(n4759), .Z(\u_a23_mem/n18429 ) );
  NANDN U6122 ( .B(n4730), .A(n1055), .Z(n4759) );
  NAND U6123 ( .A(n1056), .B(n4659), .Z(n4730) );
  AND U6124 ( .A(n4760), .B(n4761), .Z(n4758) );
  NAND U6125 ( .A(n4733), .B(\u_a23_mem/p_mem[123][7] ), .Z(n4761) );
  NANDN U6126 ( .B(n1059), .A(n4659), .Z(n4733) );
  NAND U6127 ( .A(n1061), .B(n4659), .Z(n4760) );
  ANDN U6128 ( .A(n1327), .B(n4640), .Z(n4659) );
  AND U6129 ( .A(n4146), .B(m_address[3]), .Z(n1327) );
  NAND U6130 ( .A(n4762), .B(n4763), .Z(\u_a23_mem/n18428 ) );
  NAND U6131 ( .A(n4764), .B(\u_a23_mem/p_mem[124][0] ), .Z(n4763) );
  OR U6132 ( .A(n1011), .B(n4765), .Z(n4762) );
  NAND U6133 ( .A(n4766), .B(n4767), .Z(\u_a23_mem/n18427 ) );
  NAND U6134 ( .A(n4764), .B(\u_a23_mem/p_mem[124][1] ), .Z(n4767) );
  OR U6135 ( .A(n1019), .B(n4765), .Z(n4766) );
  NAND U6136 ( .A(n4768), .B(n4769), .Z(\u_a23_mem/n18426 ) );
  NAND U6137 ( .A(n4764), .B(\u_a23_mem/p_mem[124][2] ), .Z(n4769) );
  OR U6138 ( .A(n1025), .B(n4765), .Z(n4768) );
  NAND U6139 ( .A(n4770), .B(n4771), .Z(\u_a23_mem/n18425 ) );
  NAND U6140 ( .A(n4764), .B(\u_a23_mem/p_mem[124][3] ), .Z(n4771) );
  OR U6141 ( .A(n1031), .B(n4765), .Z(n4770) );
  NAND U6142 ( .A(n4772), .B(n4773), .Z(\u_a23_mem/n18424 ) );
  NAND U6143 ( .A(n4764), .B(\u_a23_mem/p_mem[124][4] ), .Z(n4773) );
  OR U6144 ( .A(n1037), .B(n4765), .Z(n4772) );
  NAND U6145 ( .A(n4774), .B(n4775), .Z(\u_a23_mem/n18423 ) );
  NAND U6146 ( .A(n4764), .B(\u_a23_mem/p_mem[124][5] ), .Z(n4775) );
  OR U6147 ( .A(n1043), .B(n4765), .Z(n4774) );
  NAND U6148 ( .A(n4776), .B(n4777), .Z(\u_a23_mem/n18422 ) );
  NAND U6149 ( .A(n4764), .B(\u_a23_mem/p_mem[124][6] ), .Z(n4777) );
  OR U6150 ( .A(n1049), .B(n4765), .Z(n4776) );
  NAND U6151 ( .A(n4778), .B(n4779), .Z(\u_a23_mem/n18421 ) );
  NAND U6152 ( .A(n4764), .B(\u_a23_mem/p_mem[124][7] ), .Z(n4779) );
  OR U6153 ( .A(n1080), .B(n4780), .Z(n4764) );
  NAND U6154 ( .A(n2938), .B(n899), .Z(n1080) );
  NANDN U6155 ( .B(n4765), .A(n1055), .Z(n4778) );
  OR U6156 ( .A(n2), .B(n4780), .Z(n4765) );
  NAND U6157 ( .A(n4781), .B(n4782), .Z(\u_a23_mem/n18420 ) );
  OR U6158 ( .A(n1011), .B(n4783), .Z(n4782) );
  AND U6159 ( .A(n4784), .B(n4785), .Z(n4781) );
  NANDN U6160 ( .B(n1087), .A(n4786), .Z(n4785) );
  NAND U6161 ( .A(n2938), .B(n9), .Z(n1087) );
  NAND U6162 ( .A(n4787), .B(\u_a23_mem/p_mem[125][0] ), .Z(n4784) );
  NAND U6163 ( .A(n4788), .B(n4789), .Z(\u_a23_mem/n18419 ) );
  OR U6164 ( .A(n1019), .B(n4783), .Z(n4789) );
  AND U6165 ( .A(n4790), .B(n4791), .Z(n4788) );
  NANDN U6166 ( .B(n1093), .A(n4786), .Z(n4791) );
  NAND U6167 ( .A(n2938), .B(n16), .Z(n1093) );
  NAND U6168 ( .A(n4787), .B(\u_a23_mem/p_mem[125][1] ), .Z(n4790) );
  NAND U6169 ( .A(n4792), .B(n4793), .Z(\u_a23_mem/n18418 ) );
  OR U6170 ( .A(n1025), .B(n4783), .Z(n4793) );
  AND U6171 ( .A(n4794), .B(n4795), .Z(n4792) );
  NANDN U6172 ( .B(n1098), .A(n4786), .Z(n4795) );
  NAND U6173 ( .A(n2938), .B(n22), .Z(n1098) );
  NAND U6174 ( .A(n4787), .B(\u_a23_mem/p_mem[125][2] ), .Z(n4794) );
  NAND U6175 ( .A(n4796), .B(n4797), .Z(\u_a23_mem/n18417 ) );
  OR U6176 ( .A(n1031), .B(n4783), .Z(n4797) );
  AND U6177 ( .A(n4798), .B(n4799), .Z(n4796) );
  NANDN U6178 ( .B(n1103), .A(n4786), .Z(n4799) );
  NAND U6179 ( .A(n2938), .B(n28), .Z(n1103) );
  NAND U6180 ( .A(n4787), .B(\u_a23_mem/p_mem[125][3] ), .Z(n4798) );
  NAND U6181 ( .A(n4800), .B(n4801), .Z(\u_a23_mem/n18416 ) );
  OR U6182 ( .A(n1037), .B(n4783), .Z(n4801) );
  AND U6183 ( .A(n4802), .B(n4803), .Z(n4800) );
  NANDN U6184 ( .B(n1108), .A(n4786), .Z(n4803) );
  NAND U6185 ( .A(n2938), .B(n34), .Z(n1108) );
  NAND U6186 ( .A(n4787), .B(\u_a23_mem/p_mem[125][4] ), .Z(n4802) );
  NAND U6187 ( .A(n4804), .B(n4805), .Z(\u_a23_mem/n18415 ) );
  OR U6188 ( .A(n1043), .B(n4783), .Z(n4805) );
  AND U6189 ( .A(n4806), .B(n4807), .Z(n4804) );
  NANDN U6190 ( .B(n1113), .A(n4786), .Z(n4807) );
  NAND U6191 ( .A(n2938), .B(n40), .Z(n1113) );
  NAND U6192 ( .A(n4787), .B(\u_a23_mem/p_mem[125][5] ), .Z(n4806) );
  NAND U6193 ( .A(n4808), .B(n4809), .Z(\u_a23_mem/n18414 ) );
  OR U6194 ( .A(n1049), .B(n4783), .Z(n4809) );
  AND U6195 ( .A(n4810), .B(n4811), .Z(n4808) );
  NANDN U6196 ( .B(n1118), .A(n4786), .Z(n4811) );
  NAND U6197 ( .A(n2938), .B(n46), .Z(n1118) );
  NAND U6198 ( .A(n4787), .B(\u_a23_mem/p_mem[125][6] ), .Z(n4810) );
  NAND U6199 ( .A(n4812), .B(n4813), .Z(\u_a23_mem/n18413 ) );
  NANDN U6200 ( .B(n4783), .A(n1055), .Z(n4813) );
  NAND U6201 ( .A(n4786), .B(n1121), .Z(n4783) );
  AND U6202 ( .A(n4814), .B(n4815), .Z(n4812) );
  NANDN U6203 ( .B(n1124), .A(n4786), .Z(n4815) );
  NAND U6204 ( .A(n2938), .B(n53), .Z(n1124) );
  NAND U6205 ( .A(n4787), .B(\u_a23_mem/p_mem[125][7] ), .Z(n4814) );
  OR U6206 ( .A(n1125), .B(n4780), .Z(n4787) );
  NAND U6207 ( .A(n2938), .B(n933), .Z(n1125) );
  NAND U6208 ( .A(n4816), .B(n4817), .Z(\u_a23_mem/n18412 ) );
  OR U6209 ( .A(n1011), .B(n4818), .Z(n4817) );
  AND U6210 ( .A(n4819), .B(n4820), .Z(n4816) );
  NANDN U6211 ( .B(n1131), .A(n4786), .Z(n4820) );
  NAND U6212 ( .A(n2938), .B(n60), .Z(n1131) );
  NAND U6213 ( .A(n4821), .B(\u_a23_mem/p_mem[126][0] ), .Z(n4819) );
  NAND U6214 ( .A(n4822), .B(n4823), .Z(\u_a23_mem/n18411 ) );
  OR U6215 ( .A(n1019), .B(n4818), .Z(n4823) );
  AND U6216 ( .A(n4824), .B(n4825), .Z(n4822) );
  NANDN U6217 ( .B(n1137), .A(n4786), .Z(n4825) );
  NAND U6218 ( .A(n2938), .B(n66), .Z(n1137) );
  NAND U6219 ( .A(n4821), .B(\u_a23_mem/p_mem[126][1] ), .Z(n4824) );
  NAND U6220 ( .A(n4826), .B(n4827), .Z(\u_a23_mem/n18410 ) );
  OR U6221 ( .A(n1025), .B(n4818), .Z(n4827) );
  AND U6222 ( .A(n4828), .B(n4829), .Z(n4826) );
  NANDN U6223 ( .B(n1142), .A(n4786), .Z(n4829) );
  NAND U6224 ( .A(n2938), .B(n71), .Z(n1142) );
  NAND U6225 ( .A(n4821), .B(\u_a23_mem/p_mem[126][2] ), .Z(n4828) );
  NAND U6226 ( .A(n4830), .B(n4831), .Z(\u_a23_mem/n18409 ) );
  OR U6227 ( .A(n1031), .B(n4818), .Z(n4831) );
  AND U6228 ( .A(n4832), .B(n4833), .Z(n4830) );
  NANDN U6229 ( .B(n1147), .A(n4786), .Z(n4833) );
  NAND U6230 ( .A(n2938), .B(n76), .Z(n1147) );
  NAND U6231 ( .A(n4821), .B(\u_a23_mem/p_mem[126][3] ), .Z(n4832) );
  NAND U6232 ( .A(n4834), .B(n4835), .Z(\u_a23_mem/n18408 ) );
  OR U6233 ( .A(n1037), .B(n4818), .Z(n4835) );
  AND U6234 ( .A(n4836), .B(n4837), .Z(n4834) );
  NANDN U6235 ( .B(n1152), .A(n4786), .Z(n4837) );
  NAND U6236 ( .A(n2938), .B(n81), .Z(n1152) );
  NAND U6237 ( .A(n4821), .B(\u_a23_mem/p_mem[126][4] ), .Z(n4836) );
  NAND U6238 ( .A(n4838), .B(n4839), .Z(\u_a23_mem/n18407 ) );
  OR U6239 ( .A(n1043), .B(n4818), .Z(n4839) );
  AND U6240 ( .A(n4840), .B(n4841), .Z(n4838) );
  NANDN U6241 ( .B(n1157), .A(n4786), .Z(n4841) );
  NAND U6242 ( .A(n2938), .B(n86), .Z(n1157) );
  NAND U6243 ( .A(n4821), .B(\u_a23_mem/p_mem[126][5] ), .Z(n4840) );
  NAND U6244 ( .A(n4842), .B(n4843), .Z(\u_a23_mem/n18406 ) );
  OR U6245 ( .A(n4818), .B(n1049), .Z(n4843) );
  AND U6246 ( .A(n4844), .B(n4845), .Z(n4842) );
  NANDN U6247 ( .B(n1162), .A(n4786), .Z(n4845) );
  NAND U6248 ( .A(n2938), .B(n91), .Z(n1162) );
  NAND U6249 ( .A(n4821), .B(\u_a23_mem/p_mem[126][6] ), .Z(n4844) );
  NAND U6250 ( .A(n4846), .B(n4847), .Z(\u_a23_mem/n18405 ) );
  NANDN U6251 ( .B(n4818), .A(n1055), .Z(n4847) );
  NAND U6252 ( .A(n4786), .B(n1165), .Z(n4818) );
  AND U6253 ( .A(n4848), .B(n4849), .Z(n4846) );
  NANDN U6254 ( .B(n1168), .A(n4786), .Z(n4849) );
  NAND U6255 ( .A(n2938), .B(n98), .Z(n1168) );
  NAND U6256 ( .A(n4821), .B(\u_a23_mem/p_mem[126][7] ), .Z(n4848) );
  OR U6257 ( .A(n1169), .B(n4780), .Z(n4821) );
  NAND U6258 ( .A(n2938), .B(n968), .Z(n1169) );
  NAND U6259 ( .A(n4850), .B(n4851), .Z(\u_a23_mem/n18404 ) );
  NANDN U6260 ( .B(n1011), .A(n4852), .Z(n4851) );
  NAND U6261 ( .A(n2938), .B(m_write[0]), .Z(n1011) );
  AND U6262 ( .A(n4853), .B(n4854), .Z(n4850) );
  NAND U6263 ( .A(n4855), .B(\u_a23_mem/p_mem[127][0] ), .Z(n4854) );
  NANDN U6264 ( .B(n1015), .A(n4786), .Z(n4853) );
  NAND U6265 ( .A(n2938), .B(n104), .Z(n1015) );
  NAND U6266 ( .A(n4856), .B(n4857), .Z(\u_a23_mem/n18403 ) );
  NANDN U6267 ( .B(n1019), .A(n4852), .Z(n4857) );
  NAND U6268 ( .A(n2938), .B(m_write[1]), .Z(n1019) );
  AND U6269 ( .A(n4858), .B(n4859), .Z(n4856) );
  NAND U6270 ( .A(n4855), .B(\u_a23_mem/p_mem[127][1] ), .Z(n4859) );
  NANDN U6271 ( .B(n1022), .A(n4786), .Z(n4858) );
  NAND U6272 ( .A(n2938), .B(n110), .Z(n1022) );
  NAND U6273 ( .A(n4860), .B(n4861), .Z(\u_a23_mem/n18402 ) );
  NANDN U6274 ( .B(n1025), .A(n4852), .Z(n4861) );
  NAND U6275 ( .A(n2938), .B(m_write[2]), .Z(n1025) );
  AND U6276 ( .A(n4862), .B(n4863), .Z(n4860) );
  NAND U6277 ( .A(n4855), .B(\u_a23_mem/p_mem[127][2] ), .Z(n4863) );
  NANDN U6278 ( .B(n1028), .A(n4786), .Z(n4862) );
  NAND U6279 ( .A(n2938), .B(n115), .Z(n1028) );
  NAND U6280 ( .A(n4864), .B(n4865), .Z(\u_a23_mem/n18401 ) );
  NANDN U6281 ( .B(n1031), .A(n4852), .Z(n4865) );
  NAND U6282 ( .A(n2938), .B(m_write[3]), .Z(n1031) );
  AND U6283 ( .A(n4866), .B(n4867), .Z(n4864) );
  NAND U6284 ( .A(n4855), .B(\u_a23_mem/p_mem[127][3] ), .Z(n4867) );
  NANDN U6285 ( .B(n1034), .A(n4786), .Z(n4866) );
  NAND U6286 ( .A(n2938), .B(n120), .Z(n1034) );
  NAND U6287 ( .A(n4868), .B(n4869), .Z(\u_a23_mem/n18400 ) );
  NANDN U6288 ( .B(n1037), .A(n4852), .Z(n4869) );
  NAND U6289 ( .A(n2938), .B(m_write[4]), .Z(n1037) );
  AND U6290 ( .A(n4870), .B(n4871), .Z(n4868) );
  NAND U6291 ( .A(n4855), .B(\u_a23_mem/p_mem[127][4] ), .Z(n4871) );
  NANDN U6292 ( .B(n1040), .A(n4786), .Z(n4870) );
  NAND U6293 ( .A(n2938), .B(n125), .Z(n1040) );
  NAND U6294 ( .A(n4872), .B(n4873), .Z(\u_a23_mem/n18399 ) );
  NANDN U6295 ( .B(n1043), .A(n4852), .Z(n4873) );
  NAND U6296 ( .A(n2938), .B(m_write[5]), .Z(n1043) );
  AND U6297 ( .A(n4874), .B(n4875), .Z(n4872) );
  NAND U6298 ( .A(n4855), .B(\u_a23_mem/p_mem[127][5] ), .Z(n4875) );
  NANDN U6299 ( .B(n1046), .A(n4786), .Z(n4874) );
  NAND U6300 ( .A(n2938), .B(n130), .Z(n1046) );
  NAND U6301 ( .A(n4876), .B(n4877), .Z(\u_a23_mem/n18398 ) );
  NANDN U6302 ( .B(n1049), .A(n4852), .Z(n4877) );
  NAND U6303 ( .A(n2938), .B(m_write[6]), .Z(n1049) );
  AND U6304 ( .A(n4878), .B(n4879), .Z(n4876) );
  NAND U6305 ( .A(n4855), .B(\u_a23_mem/p_mem[127][6] ), .Z(n4879) );
  NANDN U6306 ( .B(n1052), .A(n4786), .Z(n4878) );
  NAND U6307 ( .A(n2938), .B(n135), .Z(n1052) );
  NAND U6308 ( .A(n4880), .B(n4881), .Z(\u_a23_mem/n18397 ) );
  NAND U6309 ( .A(n4852), .B(n1055), .Z(n4881) );
  ANDN U6310 ( .A(m_write[7]), .B(n4882), .Z(n1055) );
  ANDN U6311 ( .A(n4786), .B(n2977), .Z(n4852) );
  AND U6312 ( .A(n4883), .B(n4884), .Z(n4880) );
  NAND U6313 ( .A(n4855), .B(\u_a23_mem/p_mem[127][7] ), .Z(n4884) );
  OR U6314 ( .A(n1059), .B(n4780), .Z(n4855) );
  NAND U6315 ( .A(n2938), .B(n1003), .Z(n1059) );
  NAND U6316 ( .A(n4786), .B(n1061), .Z(n4883) );
  ANDN U6317 ( .A(n142), .B(n4882), .Z(n1061) );
  IV U6318 ( .A(n4780), .Z(n4786) );
  NANDN U6319 ( .B(n4640), .A(n1449), .Z(n4780) );
  AND U6320 ( .A(m_address[2]), .B(m_address[3]), .Z(n1449) );
  NAND U6321 ( .A(n4515), .B(n4885), .Z(n4640) );
  AND U6322 ( .A(n4148), .B(m_address[4]), .Z(n4885) );
  AND U6323 ( .A(m_address[5]), .B(m_address[6]), .Z(n4515) );
  NAND U6324 ( .A(n4886), .B(n4887), .Z(\u_a23_mem/n18396 ) );
  NAND U6325 ( .A(n4888), .B(\u_a23_mem/p_mem[2][0] ), .Z(n4887) );
  AND U6326 ( .A(n4889), .B(n4890), .Z(n4886) );
  NANDN U6327 ( .B(n4891), .A(n60), .Z(n4890) );
  NANDN U6328 ( .B(n4892), .A(m_write[0]), .Z(n4889) );
  NAND U6329 ( .A(n4893), .B(n4894), .Z(\u_a23_mem/n18395 ) );
  NAND U6330 ( .A(n4888), .B(\u_a23_mem/p_mem[2][1] ), .Z(n4894) );
  AND U6331 ( .A(n4895), .B(n4896), .Z(n4893) );
  NANDN U6332 ( .B(n4891), .A(n66), .Z(n4896) );
  NANDN U6333 ( .B(n4892), .A(m_write[1]), .Z(n4895) );
  NAND U6334 ( .A(n4897), .B(n4898), .Z(\u_a23_mem/n18394 ) );
  NAND U6335 ( .A(n4888), .B(\u_a23_mem/p_mem[2][2] ), .Z(n4898) );
  AND U6336 ( .A(n4899), .B(n4900), .Z(n4897) );
  NANDN U6337 ( .B(n4891), .A(n71), .Z(n4900) );
  NANDN U6338 ( .B(n4892), .A(m_write[2]), .Z(n4899) );
  NAND U6339 ( .A(n4901), .B(n4902), .Z(\u_a23_mem/n18393 ) );
  NAND U6340 ( .A(n4888), .B(\u_a23_mem/p_mem[2][3] ), .Z(n4902) );
  AND U6341 ( .A(n4903), .B(n4904), .Z(n4901) );
  NANDN U6342 ( .B(n4891), .A(n76), .Z(n4904) );
  NANDN U6343 ( .B(n4892), .A(m_write[3]), .Z(n4903) );
  NAND U6344 ( .A(n4905), .B(n4906), .Z(\u_a23_mem/n18392 ) );
  NAND U6345 ( .A(n4888), .B(\u_a23_mem/p_mem[2][4] ), .Z(n4906) );
  AND U6346 ( .A(n4907), .B(n4908), .Z(n4905) );
  NANDN U6347 ( .B(n4891), .A(n81), .Z(n4908) );
  NANDN U6348 ( .B(n4892), .A(m_write[4]), .Z(n4907) );
  NAND U6349 ( .A(n4909), .B(n4910), .Z(\u_a23_mem/n18391 ) );
  NAND U6350 ( .A(n4888), .B(\u_a23_mem/p_mem[2][5] ), .Z(n4910) );
  AND U6351 ( .A(n4911), .B(n4912), .Z(n4909) );
  NANDN U6352 ( .B(n4891), .A(n86), .Z(n4912) );
  NANDN U6353 ( .B(n4892), .A(m_write[5]), .Z(n4911) );
  NAND U6354 ( .A(n4913), .B(n4914), .Z(\u_a23_mem/n18390 ) );
  NAND U6355 ( .A(n4888), .B(\u_a23_mem/p_mem[2][6] ), .Z(n4914) );
  AND U6356 ( .A(n4915), .B(n4916), .Z(n4913) );
  NANDN U6357 ( .B(n4891), .A(n91), .Z(n4916) );
  NANDN U6358 ( .B(n4892), .A(m_write[6]), .Z(n4915) );
  NAND U6359 ( .A(n4917), .B(n4918), .Z(\u_a23_mem/n18389 ) );
  NAND U6360 ( .A(n4888), .B(\u_a23_mem/p_mem[2][7] ), .Z(n4918) );
  NANDN U6361 ( .B(n4882), .A(n4919), .Z(n4888) );
  ANDN U6362 ( .A(n1016), .B(n4920), .Z(n4919) );
  AND U6363 ( .A(n4921), .B(n4922), .Z(n4917) );
  NANDN U6364 ( .B(n4891), .A(n98), .Z(n4922) );
  NAND U6365 ( .A(n1016), .B(n2938), .Z(n4891) );
  NANDN U6366 ( .B(n4892), .A(m_write[7]), .Z(n4921) );
  NAND U6367 ( .A(n2938), .B(n4923), .Z(n4892) );
  AND U6368 ( .A(n1016), .B(n1165), .Z(n4923) );
  NAND U6369 ( .A(n4924), .B(n4925), .Z(\u_a23_mem/n18388 ) );
  NAND U6370 ( .A(n4926), .B(\u_a23_mem/p_mem[1][0] ), .Z(n4925) );
  AND U6371 ( .A(n4927), .B(n4928), .Z(n4924) );
  NAND U6372 ( .A(n9), .B(n4929), .Z(n4928) );
  NANDN U6373 ( .B(n4930), .A(m_write[0]), .Z(n4927) );
  NAND U6374 ( .A(n4931), .B(n4932), .Z(\u_a23_mem/n18387 ) );
  NAND U6375 ( .A(n4926), .B(\u_a23_mem/p_mem[1][1] ), .Z(n4932) );
  AND U6376 ( .A(n4933), .B(n4934), .Z(n4931) );
  NAND U6377 ( .A(n16), .B(n4929), .Z(n4934) );
  NANDN U6378 ( .B(n4930), .A(m_write[1]), .Z(n4933) );
  NAND U6379 ( .A(n4935), .B(n4936), .Z(\u_a23_mem/n18386 ) );
  NAND U6380 ( .A(n4926), .B(\u_a23_mem/p_mem[1][2] ), .Z(n4936) );
  AND U6381 ( .A(n4937), .B(n4938), .Z(n4935) );
  NAND U6382 ( .A(n22), .B(n4929), .Z(n4938) );
  NANDN U6383 ( .B(n4930), .A(m_write[2]), .Z(n4937) );
  NAND U6384 ( .A(n4939), .B(n4940), .Z(\u_a23_mem/n18385 ) );
  NAND U6385 ( .A(n4926), .B(\u_a23_mem/p_mem[1][3] ), .Z(n4940) );
  AND U6386 ( .A(n4941), .B(n4942), .Z(n4939) );
  NAND U6387 ( .A(n28), .B(n4929), .Z(n4942) );
  NANDN U6388 ( .B(n4930), .A(m_write[3]), .Z(n4941) );
  NAND U6389 ( .A(n4943), .B(n4944), .Z(\u_a23_mem/n18384 ) );
  NAND U6390 ( .A(n4926), .B(\u_a23_mem/p_mem[1][4] ), .Z(n4944) );
  AND U6391 ( .A(n4945), .B(n4946), .Z(n4943) );
  NAND U6392 ( .A(n34), .B(n4929), .Z(n4946) );
  NANDN U6393 ( .B(n4930), .A(m_write[4]), .Z(n4945) );
  NAND U6394 ( .A(n4947), .B(n4948), .Z(\u_a23_mem/n18383 ) );
  NAND U6395 ( .A(n4926), .B(\u_a23_mem/p_mem[1][5] ), .Z(n4948) );
  AND U6396 ( .A(n4949), .B(n4950), .Z(n4947) );
  NAND U6397 ( .A(n40), .B(n4929), .Z(n4950) );
  NANDN U6398 ( .B(n4930), .A(m_write[5]), .Z(n4949) );
  NAND U6399 ( .A(n4951), .B(n4952), .Z(\u_a23_mem/n18382 ) );
  NAND U6400 ( .A(n4926), .B(\u_a23_mem/p_mem[1][6] ), .Z(n4952) );
  AND U6401 ( .A(n4953), .B(n4954), .Z(n4951) );
  NAND U6402 ( .A(n46), .B(n4929), .Z(n4954) );
  NANDN U6403 ( .B(n4930), .A(m_write[6]), .Z(n4953) );
  NAND U6404 ( .A(n4955), .B(n4956), .Z(\u_a23_mem/n18381 ) );
  NAND U6405 ( .A(n4926), .B(\u_a23_mem/p_mem[1][7] ), .Z(n4956) );
  NANDN U6406 ( .B(n4882), .A(n4957), .Z(n4926) );
  AND U6407 ( .A(n50), .B(n1016), .Z(n4957) );
  AND U6408 ( .A(n4958), .B(n4959), .Z(n4955) );
  NAND U6409 ( .A(n53), .B(n4929), .Z(n4959) );
  NANDN U6410 ( .B(n4930), .A(m_write[7]), .Z(n4958) );
  NAND U6411 ( .A(n2938), .B(n4960), .Z(n4930) );
  AND U6412 ( .A(n1016), .B(n1121), .Z(n4960) );
  IV U6413 ( .A(n4882), .Z(n2938) );
  MUX U6414 ( .IN0(\u_a23_mem/p_mem[0][0] ), .IN1(m_write[0]), .SEL(n4961), 
        .F(\u_a23_mem/n18380 ) );
  MUX U6415 ( .IN0(\u_a23_mem/p_mem[0][1] ), .IN1(m_write[1]), .SEL(n4961), 
        .F(\u_a23_mem/n18379 ) );
  MUX U6416 ( .IN0(\u_a23_mem/p_mem[0][2] ), .IN1(m_write[2]), .SEL(n4961), 
        .F(\u_a23_mem/n18378 ) );
  MUX U6417 ( .IN0(\u_a23_mem/p_mem[0][3] ), .IN1(m_write[3]), .SEL(n4961), 
        .F(\u_a23_mem/n18377 ) );
  MUX U6418 ( .IN0(\u_a23_mem/p_mem[0][4] ), .IN1(m_write[4]), .SEL(n4961), 
        .F(\u_a23_mem/n18376 ) );
  MUX U6419 ( .IN0(\u_a23_mem/p_mem[0][5] ), .IN1(m_write[5]), .SEL(n4961), 
        .F(\u_a23_mem/n18375 ) );
  MUX U6420 ( .IN0(\u_a23_mem/p_mem[0][6] ), .IN1(m_write[6]), .SEL(n4961), 
        .F(\u_a23_mem/n18374 ) );
  MUX U6421 ( .IN0(\u_a23_mem/p_mem[0][7] ), .IN1(m_write[7]), .SEL(n4961), 
        .F(\u_a23_mem/n18373 ) );
  ANDN U6422 ( .A(n4929), .B(n2), .Z(n4961) );
  ANDN U6423 ( .A(n1016), .B(n4882), .Z(n4929) );
  NANDN U6424 ( .B(n4962), .A(m_write_en), .Z(n4882) );
  ANDN U6425 ( .A(n4517), .B(n1205), .Z(n1016) );
  NANDN U6426 ( .B(m_address[4]), .A(n4963), .Z(n1205) );
  AND U6427 ( .A(n4146), .B(n4147), .Z(n4517) );
  MUX U6428 ( .IN0(o[0]), .IN1(m_write[0]), .SEL(n4964), .F(\u_a23_mem/n18372 ) );
  MUX U6429 ( .IN0(o[1]), .IN1(m_write[1]), .SEL(n4964), .F(\u_a23_mem/n18371 ) );
  MUX U6430 ( .IN0(o[2]), .IN1(m_write[2]), .SEL(n4964), .F(\u_a23_mem/n18370 ) );
  MUX U6431 ( .IN0(o[3]), .IN1(m_write[3]), .SEL(n4964), .F(\u_a23_mem/n18369 ) );
  MUX U6432 ( .IN0(o[4]), .IN1(m_write[4]), .SEL(n4964), .F(\u_a23_mem/n18368 ) );
  MUX U6433 ( .IN0(o[5]), .IN1(m_write[5]), .SEL(n4964), .F(\u_a23_mem/n18367 ) );
  MUX U6434 ( .IN0(o[6]), .IN1(m_write[6]), .SEL(n4964), .F(\u_a23_mem/n18366 ) );
  MUX U6435 ( .IN0(o[7]), .IN1(m_write[7]), .SEL(n4964), .F(\u_a23_mem/n18365 ) );
  NOR U6436 ( .A(n4965), .B(n2), .Z(n4964) );
  NAND U6437 ( .A(n4966), .B(n4967), .Z(\u_a23_mem/n18364 ) );
  NAND U6438 ( .A(n4968), .B(o[8]), .Z(n4967) );
  AND U6439 ( .A(n4969), .B(n4970), .Z(n4966) );
  NAND U6440 ( .A(n4971), .B(n9), .Z(n4970) );
  OR U6441 ( .A(n10), .B(n4972), .Z(n4969) );
  NAND U6442 ( .A(n4973), .B(n4974), .Z(\u_a23_mem/n18363 ) );
  NAND U6443 ( .A(n4968), .B(o[9]), .Z(n4974) );
  AND U6444 ( .A(n4975), .B(n4976), .Z(n4973) );
  NAND U6445 ( .A(n4971), .B(n16), .Z(n4976) );
  OR U6446 ( .A(n10), .B(n4977), .Z(n4975) );
  NAND U6447 ( .A(n4978), .B(n4979), .Z(\u_a23_mem/n18362 ) );
  NAND U6448 ( .A(n4968), .B(o[10]), .Z(n4979) );
  AND U6449 ( .A(n4980), .B(n4981), .Z(n4978) );
  NAND U6450 ( .A(n4971), .B(n22), .Z(n4981) );
  OR U6451 ( .A(n10), .B(n4982), .Z(n4980) );
  NAND U6452 ( .A(n4983), .B(n4984), .Z(\u_a23_mem/n18361 ) );
  NAND U6453 ( .A(n4968), .B(o[11]), .Z(n4984) );
  AND U6454 ( .A(n4985), .B(n4986), .Z(n4983) );
  NAND U6455 ( .A(n4971), .B(n28), .Z(n4986) );
  OR U6456 ( .A(n10), .B(n4987), .Z(n4985) );
  NAND U6457 ( .A(n4988), .B(n4989), .Z(\u_a23_mem/n18360 ) );
  NAND U6458 ( .A(n4968), .B(o[12]), .Z(n4989) );
  AND U6459 ( .A(n4990), .B(n4991), .Z(n4988) );
  NAND U6460 ( .A(n4971), .B(n34), .Z(n4991) );
  OR U6461 ( .A(n10), .B(n4992), .Z(n4990) );
  NAND U6462 ( .A(n4993), .B(n4994), .Z(\u_a23_mem/n18359 ) );
  NAND U6463 ( .A(n4968), .B(o[13]), .Z(n4994) );
  AND U6464 ( .A(n4995), .B(n4996), .Z(n4993) );
  NAND U6465 ( .A(n4971), .B(n40), .Z(n4996) );
  OR U6466 ( .A(n10), .B(n4997), .Z(n4995) );
  NAND U6467 ( .A(n4998), .B(n4999), .Z(\u_a23_mem/n18358 ) );
  NAND U6468 ( .A(n4968), .B(o[14]), .Z(n4999) );
  AND U6469 ( .A(n5000), .B(n5001), .Z(n4998) );
  NAND U6470 ( .A(n4971), .B(n46), .Z(n5001) );
  OR U6471 ( .A(n5002), .B(n10), .Z(n5000) );
  NAND U6472 ( .A(n5003), .B(n5004), .Z(\u_a23_mem/n18357 ) );
  NAND U6473 ( .A(n4968), .B(o[15]), .Z(n5004) );
  NANDN U6474 ( .B(n4965), .A(n50), .Z(n4968) );
  ANDN U6475 ( .A(n5005), .B(n5006), .Z(n50) );
  NAND U6476 ( .A(n2937), .B(n2), .Z(n5005) );
  IV U6477 ( .A(n4971), .Z(n4965) );
  AND U6478 ( .A(n5007), .B(n5008), .Z(n5003) );
  NAND U6479 ( .A(n4971), .B(n53), .Z(n5008) );
  NANDN U6480 ( .B(n10), .A(n5009), .Z(n5007) );
  NAND U6481 ( .A(n143), .B(n1121), .Z(n10) );
  NAND U6482 ( .A(n5010), .B(n5011), .Z(\u_a23_mem/n18356 ) );
  NAND U6483 ( .A(n5012), .B(o[16]), .Z(n5011) );
  AND U6484 ( .A(n5013), .B(n5014), .Z(n5010) );
  NAND U6485 ( .A(n4971), .B(n60), .Z(n5014) );
  OR U6486 ( .A(n61), .B(n4972), .Z(n5013) );
  NAND U6487 ( .A(n5015), .B(n5016), .Z(\u_a23_mem/n18355 ) );
  NAND U6488 ( .A(n5012), .B(o[17]), .Z(n5016) );
  AND U6489 ( .A(n5017), .B(n5018), .Z(n5015) );
  NAND U6490 ( .A(n4971), .B(n66), .Z(n5018) );
  OR U6491 ( .A(n61), .B(n4977), .Z(n5017) );
  NAND U6492 ( .A(n5019), .B(n5020), .Z(\u_a23_mem/n18354 ) );
  NAND U6493 ( .A(n5012), .B(o[18]), .Z(n5020) );
  AND U6494 ( .A(n5021), .B(n5022), .Z(n5019) );
  NAND U6495 ( .A(n4971), .B(n71), .Z(n5022) );
  OR U6496 ( .A(n61), .B(n4982), .Z(n5021) );
  NAND U6497 ( .A(n5023), .B(n5024), .Z(\u_a23_mem/n18353 ) );
  NAND U6498 ( .A(n5012), .B(o[19]), .Z(n5024) );
  AND U6499 ( .A(n5025), .B(n5026), .Z(n5023) );
  NAND U6500 ( .A(n4971), .B(n76), .Z(n5026) );
  OR U6501 ( .A(n61), .B(n4987), .Z(n5025) );
  NAND U6502 ( .A(n5027), .B(n5028), .Z(\u_a23_mem/n18352 ) );
  NAND U6503 ( .A(n5012), .B(o[20]), .Z(n5028) );
  AND U6504 ( .A(n5029), .B(n5030), .Z(n5027) );
  NAND U6505 ( .A(n4971), .B(n81), .Z(n5030) );
  OR U6506 ( .A(n61), .B(n4992), .Z(n5029) );
  NAND U6507 ( .A(n5031), .B(n5032), .Z(\u_a23_mem/n18351 ) );
  NAND U6508 ( .A(n5012), .B(o[21]), .Z(n5032) );
  AND U6509 ( .A(n5033), .B(n5034), .Z(n5031) );
  NAND U6510 ( .A(n4971), .B(n86), .Z(n5034) );
  OR U6511 ( .A(n61), .B(n4997), .Z(n5033) );
  NAND U6512 ( .A(n5035), .B(n5036), .Z(\u_a23_mem/n18350 ) );
  NAND U6513 ( .A(n5012), .B(o[22]), .Z(n5036) );
  AND U6514 ( .A(n5037), .B(n5038), .Z(n5035) );
  NAND U6515 ( .A(n4971), .B(n91), .Z(n5038) );
  OR U6516 ( .A(n61), .B(n5002), .Z(n5037) );
  NAND U6517 ( .A(n5039), .B(n5040), .Z(\u_a23_mem/n18349 ) );
  NAND U6518 ( .A(n5012), .B(o[23]), .Z(n5040) );
  OR U6519 ( .A(n94), .B(n5041), .Z(n5012) );
  NANDN U6520 ( .B(n4920), .A(n143), .Z(n94) );
  NAND U6521 ( .A(n5042), .B(n5043), .Z(n4920) );
  AND U6522 ( .A(n2980), .B(n2937), .Z(n5042) );
  AND U6523 ( .A(n5044), .B(n5045), .Z(n5039) );
  NAND U6524 ( .A(n4971), .B(n98), .Z(n5045) );
  NANDN U6525 ( .B(n61), .A(n5009), .Z(n5044) );
  NAND U6526 ( .A(n143), .B(n1165), .Z(n61) );
  NAND U6527 ( .A(n5046), .B(n5047), .Z(\u_a23_mem/n18348 ) );
  NAND U6528 ( .A(n5048), .B(o[24]), .Z(n5047) );
  AND U6529 ( .A(n5049), .B(n5050), .Z(n5046) );
  NAND U6530 ( .A(n4971), .B(n104), .Z(n5050) );
  OR U6531 ( .A(n105), .B(n4972), .Z(n5049) );
  NAND U6532 ( .A(n5051), .B(n5052), .Z(\u_a23_mem/n18347 ) );
  NAND U6533 ( .A(n5048), .B(o[25]), .Z(n5052) );
  AND U6534 ( .A(n5053), .B(n5054), .Z(n5051) );
  NAND U6535 ( .A(n4971), .B(n110), .Z(n5054) );
  OR U6536 ( .A(n105), .B(n4977), .Z(n5053) );
  NAND U6537 ( .A(n5055), .B(n5056), .Z(\u_a23_mem/n18346 ) );
  NAND U6538 ( .A(n5048), .B(o[26]), .Z(n5056) );
  AND U6539 ( .A(n5057), .B(n5058), .Z(n5055) );
  NAND U6540 ( .A(n4971), .B(n115), .Z(n5058) );
  OR U6541 ( .A(n105), .B(n4982), .Z(n5057) );
  NAND U6542 ( .A(n5059), .B(n5060), .Z(\u_a23_mem/n18345 ) );
  NAND U6543 ( .A(n5048), .B(o[27]), .Z(n5060) );
  AND U6544 ( .A(n5061), .B(n5062), .Z(n5059) );
  NAND U6545 ( .A(n4971), .B(n120), .Z(n5062) );
  OR U6546 ( .A(n105), .B(n4987), .Z(n5061) );
  NAND U6547 ( .A(n5063), .B(n5064), .Z(\u_a23_mem/n18344 ) );
  NAND U6548 ( .A(n5048), .B(o[28]), .Z(n5064) );
  AND U6549 ( .A(n5065), .B(n5066), .Z(n5063) );
  NAND U6550 ( .A(n4971), .B(n125), .Z(n5066) );
  OR U6551 ( .A(n105), .B(n4992), .Z(n5065) );
  NAND U6552 ( .A(n5067), .B(n5068), .Z(\u_a23_mem/n18343 ) );
  NAND U6553 ( .A(n5048), .B(o[29]), .Z(n5068) );
  AND U6554 ( .A(n5069), .B(n5070), .Z(n5067) );
  NAND U6555 ( .A(n4971), .B(n130), .Z(n5070) );
  OR U6556 ( .A(n105), .B(n4997), .Z(n5069) );
  NAND U6557 ( .A(n5071), .B(n5072), .Z(\u_a23_mem/n18342 ) );
  NAND U6558 ( .A(n5048), .B(o[30]), .Z(n5072) );
  AND U6559 ( .A(n5073), .B(n5074), .Z(n5071) );
  NAND U6560 ( .A(n4971), .B(n135), .Z(n5074) );
  OR U6561 ( .A(n105), .B(n5002), .Z(n5073) );
  NAND U6562 ( .A(n5075), .B(n5076), .Z(\u_a23_mem/n18341 ) );
  NAND U6563 ( .A(n5048), .B(o[31]), .Z(n5076) );
  NANDN U6564 ( .B(n139), .A(n5077), .Z(n5048) );
  AND U6565 ( .A(n5078), .B(n5079), .Z(n5075) );
  NAND U6566 ( .A(n4971), .B(n142), .Z(n5079) );
  NOR U6567 ( .A(n139), .B(n5041), .Z(n4971) );
  NANDN U6568 ( .B(n105), .A(n5009), .Z(n5078) );
  NAND U6569 ( .A(n143), .B(n1056), .Z(n105) );
  IV U6570 ( .A(n139), .Z(n143) );
  NAND U6571 ( .A(n5080), .B(n5081), .Z(n139) );
  NAND U6572 ( .A(n5082), .B(n5083), .Z(\u_a23_mem/n18340 ) );
  OR U6573 ( .A(n146), .B(n4972), .Z(n5083) );
  NAND U6574 ( .A(n5084), .B(o[32]), .Z(n5082) );
  NAND U6575 ( .A(n5085), .B(n5086), .Z(\u_a23_mem/n18339 ) );
  OR U6576 ( .A(n146), .B(n4977), .Z(n5086) );
  NAND U6577 ( .A(n5084), .B(o[33]), .Z(n5085) );
  NAND U6578 ( .A(n5087), .B(n5088), .Z(\u_a23_mem/n18338 ) );
  OR U6579 ( .A(n146), .B(n4982), .Z(n5088) );
  NAND U6580 ( .A(n5084), .B(o[34]), .Z(n5087) );
  NAND U6581 ( .A(n5089), .B(n5090), .Z(\u_a23_mem/n18337 ) );
  OR U6582 ( .A(n146), .B(n4987), .Z(n5090) );
  NAND U6583 ( .A(n5084), .B(o[35]), .Z(n5089) );
  NAND U6584 ( .A(n5091), .B(n5092), .Z(\u_a23_mem/n18336 ) );
  OR U6585 ( .A(n146), .B(n4992), .Z(n5092) );
  NAND U6586 ( .A(n5084), .B(o[36]), .Z(n5091) );
  NAND U6587 ( .A(n5093), .B(n5094), .Z(\u_a23_mem/n18335 ) );
  OR U6588 ( .A(n146), .B(n4997), .Z(n5094) );
  NAND U6589 ( .A(n5084), .B(o[37]), .Z(n5093) );
  NAND U6590 ( .A(n5095), .B(n5096), .Z(\u_a23_mem/n18334 ) );
  OR U6591 ( .A(n146), .B(n5002), .Z(n5096) );
  NAND U6592 ( .A(n5084), .B(o[38]), .Z(n5095) );
  NAND U6593 ( .A(n5097), .B(n5098), .Z(\u_a23_mem/n18333 ) );
  NANDN U6594 ( .B(n146), .A(n5009), .Z(n5098) );
  NANDN U6595 ( .B(n2), .A(n163), .Z(n146) );
  NAND U6596 ( .A(n5084), .B(o[39]), .Z(n5097) );
  NANDN U6597 ( .B(n5099), .A(n163), .Z(n5084) );
  NAND U6598 ( .A(n5100), .B(n5101), .Z(\u_a23_mem/n18332 ) );
  NAND U6599 ( .A(n5102), .B(o[40]), .Z(n5101) );
  AND U6600 ( .A(n5103), .B(n5104), .Z(n5100) );
  NANDN U6601 ( .B(n5105), .A(n9), .Z(n5104) );
  OR U6602 ( .A(n170), .B(n4972), .Z(n5103) );
  NAND U6603 ( .A(n5106), .B(n5107), .Z(\u_a23_mem/n18331 ) );
  NAND U6604 ( .A(n5102), .B(o[41]), .Z(n5107) );
  AND U6605 ( .A(n5108), .B(n5109), .Z(n5106) );
  NANDN U6606 ( .B(n5105), .A(n16), .Z(n5109) );
  OR U6607 ( .A(n170), .B(n4977), .Z(n5108) );
  NAND U6608 ( .A(n5110), .B(n5111), .Z(\u_a23_mem/n18330 ) );
  NAND U6609 ( .A(n5102), .B(o[42]), .Z(n5111) );
  AND U6610 ( .A(n5112), .B(n5113), .Z(n5110) );
  NANDN U6611 ( .B(n5105), .A(n22), .Z(n5113) );
  OR U6612 ( .A(n170), .B(n4982), .Z(n5112) );
  NAND U6613 ( .A(n5114), .B(n5115), .Z(\u_a23_mem/n18329 ) );
  NAND U6614 ( .A(n5102), .B(o[43]), .Z(n5115) );
  AND U6615 ( .A(n5116), .B(n5117), .Z(n5114) );
  NANDN U6616 ( .B(n5105), .A(n28), .Z(n5117) );
  OR U6617 ( .A(n170), .B(n4987), .Z(n5116) );
  NAND U6618 ( .A(n5118), .B(n5119), .Z(\u_a23_mem/n18328 ) );
  NAND U6619 ( .A(n5102), .B(o[44]), .Z(n5119) );
  AND U6620 ( .A(n5120), .B(n5121), .Z(n5118) );
  NANDN U6621 ( .B(n5105), .A(n34), .Z(n5121) );
  OR U6622 ( .A(n170), .B(n4992), .Z(n5120) );
  NAND U6623 ( .A(n5122), .B(n5123), .Z(\u_a23_mem/n18327 ) );
  NAND U6624 ( .A(n5102), .B(o[45]), .Z(n5123) );
  AND U6625 ( .A(n5124), .B(n5125), .Z(n5122) );
  NANDN U6626 ( .B(n5105), .A(n40), .Z(n5125) );
  OR U6627 ( .A(n170), .B(n4997), .Z(n5124) );
  NAND U6628 ( .A(n5126), .B(n5127), .Z(\u_a23_mem/n18326 ) );
  NAND U6629 ( .A(n5102), .B(o[46]), .Z(n5127) );
  AND U6630 ( .A(n5128), .B(n5129), .Z(n5126) );
  NANDN U6631 ( .B(n5105), .A(n46), .Z(n5129) );
  OR U6632 ( .A(n170), .B(n5002), .Z(n5128) );
  NAND U6633 ( .A(n5130), .B(n5131), .Z(\u_a23_mem/n18325 ) );
  NAND U6634 ( .A(n5102), .B(o[47]), .Z(n5131) );
  NANDN U6635 ( .B(n5132), .A(n163), .Z(n5102) );
  AND U6636 ( .A(n5133), .B(n5134), .Z(n5130) );
  NANDN U6637 ( .B(n5105), .A(n53), .Z(n5134) );
  NANDN U6638 ( .B(n170), .A(n5009), .Z(n5133) );
  NAND U6639 ( .A(n1121), .B(n163), .Z(n170) );
  NAND U6640 ( .A(n5135), .B(n5136), .Z(\u_a23_mem/n18324 ) );
  NAND U6641 ( .A(n5137), .B(o[48]), .Z(n5136) );
  AND U6642 ( .A(n5138), .B(n5139), .Z(n5135) );
  NANDN U6643 ( .B(n5105), .A(n60), .Z(n5139) );
  OR U6644 ( .A(n205), .B(n4972), .Z(n5138) );
  NAND U6645 ( .A(n5140), .B(n5141), .Z(\u_a23_mem/n18323 ) );
  NAND U6646 ( .A(n5137), .B(o[49]), .Z(n5141) );
  AND U6647 ( .A(n5142), .B(n5143), .Z(n5140) );
  NANDN U6648 ( .B(n5105), .A(n66), .Z(n5143) );
  OR U6649 ( .A(n205), .B(n4977), .Z(n5142) );
  NAND U6650 ( .A(n5144), .B(n5145), .Z(\u_a23_mem/n18322 ) );
  NAND U6651 ( .A(n5137), .B(o[50]), .Z(n5145) );
  AND U6652 ( .A(n5146), .B(n5147), .Z(n5144) );
  NANDN U6653 ( .B(n5105), .A(n71), .Z(n5147) );
  OR U6654 ( .A(n205), .B(n4982), .Z(n5146) );
  NAND U6655 ( .A(n5148), .B(n5149), .Z(\u_a23_mem/n18321 ) );
  NAND U6656 ( .A(n5137), .B(o[51]), .Z(n5149) );
  AND U6657 ( .A(n5150), .B(n5151), .Z(n5148) );
  NANDN U6658 ( .B(n5105), .A(n76), .Z(n5151) );
  OR U6659 ( .A(n205), .B(n4987), .Z(n5150) );
  NAND U6660 ( .A(n5152), .B(n5153), .Z(\u_a23_mem/n18320 ) );
  NAND U6661 ( .A(n5137), .B(o[52]), .Z(n5153) );
  AND U6662 ( .A(n5154), .B(n5155), .Z(n5152) );
  NANDN U6663 ( .B(n5105), .A(n81), .Z(n5155) );
  OR U6664 ( .A(n205), .B(n4992), .Z(n5154) );
  NAND U6665 ( .A(n5156), .B(n5157), .Z(\u_a23_mem/n18319 ) );
  NAND U6666 ( .A(n5137), .B(o[53]), .Z(n5157) );
  AND U6667 ( .A(n5158), .B(n5159), .Z(n5156) );
  NANDN U6668 ( .B(n5105), .A(n86), .Z(n5159) );
  OR U6669 ( .A(n205), .B(n4997), .Z(n5158) );
  NAND U6670 ( .A(n5160), .B(n5161), .Z(\u_a23_mem/n18318 ) );
  NAND U6671 ( .A(n5137), .B(o[54]), .Z(n5161) );
  AND U6672 ( .A(n5162), .B(n5163), .Z(n5160) );
  NANDN U6673 ( .B(n5105), .A(n91), .Z(n5163) );
  OR U6674 ( .A(n205), .B(n5002), .Z(n5162) );
  NAND U6675 ( .A(n5164), .B(n5165), .Z(\u_a23_mem/n18317 ) );
  NAND U6676 ( .A(n5137), .B(o[55]), .Z(n5165) );
  NANDN U6677 ( .B(n5166), .A(n163), .Z(n5137) );
  AND U6678 ( .A(n5167), .B(n5168), .Z(n5164) );
  NANDN U6679 ( .B(n5105), .A(n98), .Z(n5168) );
  NANDN U6680 ( .B(n205), .A(n5009), .Z(n5167) );
  NAND U6681 ( .A(n1165), .B(n163), .Z(n205) );
  NAND U6682 ( .A(n5169), .B(n5170), .Z(\u_a23_mem/n18316 ) );
  NAND U6683 ( .A(n5171), .B(o[56]), .Z(n5170) );
  AND U6684 ( .A(n5172), .B(n5173), .Z(n5169) );
  NANDN U6685 ( .B(n5105), .A(n104), .Z(n5173) );
  OR U6686 ( .A(n240), .B(n4972), .Z(n5172) );
  NAND U6687 ( .A(n5174), .B(n5175), .Z(\u_a23_mem/n18315 ) );
  NAND U6688 ( .A(n5171), .B(o[57]), .Z(n5175) );
  AND U6689 ( .A(n5176), .B(n5177), .Z(n5174) );
  NANDN U6690 ( .B(n5105), .A(n110), .Z(n5177) );
  OR U6691 ( .A(n240), .B(n4977), .Z(n5176) );
  NAND U6692 ( .A(n5178), .B(n5179), .Z(\u_a23_mem/n18314 ) );
  NAND U6693 ( .A(n5171), .B(o[58]), .Z(n5179) );
  AND U6694 ( .A(n5180), .B(n5181), .Z(n5178) );
  NANDN U6695 ( .B(n5105), .A(n115), .Z(n5181) );
  OR U6696 ( .A(n240), .B(n4982), .Z(n5180) );
  NAND U6697 ( .A(n5182), .B(n5183), .Z(\u_a23_mem/n18313 ) );
  NAND U6698 ( .A(n5171), .B(o[59]), .Z(n5183) );
  AND U6699 ( .A(n5184), .B(n5185), .Z(n5182) );
  NANDN U6700 ( .B(n5105), .A(n120), .Z(n5185) );
  OR U6701 ( .A(n240), .B(n4987), .Z(n5184) );
  NAND U6702 ( .A(n5186), .B(n5187), .Z(\u_a23_mem/n18312 ) );
  NAND U6703 ( .A(n5171), .B(o[60]), .Z(n5187) );
  AND U6704 ( .A(n5188), .B(n5189), .Z(n5186) );
  NANDN U6705 ( .B(n5105), .A(n125), .Z(n5189) );
  OR U6706 ( .A(n240), .B(n4992), .Z(n5188) );
  NAND U6707 ( .A(n5190), .B(n5191), .Z(\u_a23_mem/n18311 ) );
  NAND U6708 ( .A(n5171), .B(o[61]), .Z(n5191) );
  AND U6709 ( .A(n5192), .B(n5193), .Z(n5190) );
  NANDN U6710 ( .B(n5105), .A(n130), .Z(n5193) );
  OR U6711 ( .A(n240), .B(n4997), .Z(n5192) );
  NAND U6712 ( .A(n5194), .B(n5195), .Z(\u_a23_mem/n18310 ) );
  NAND U6713 ( .A(n5171), .B(o[62]), .Z(n5195) );
  AND U6714 ( .A(n5196), .B(n5197), .Z(n5194) );
  NANDN U6715 ( .B(n5105), .A(n135), .Z(n5197) );
  OR U6716 ( .A(n240), .B(n5002), .Z(n5196) );
  NAND U6717 ( .A(n5198), .B(n5199), .Z(\u_a23_mem/n18309 ) );
  NAND U6718 ( .A(n5171), .B(o[63]), .Z(n5199) );
  NAND U6719 ( .A(n163), .B(n5077), .Z(n5171) );
  AND U6720 ( .A(n5200), .B(n5201), .Z(n5198) );
  NANDN U6721 ( .B(n5105), .A(n142), .Z(n5201) );
  NAND U6722 ( .A(n5202), .B(n163), .Z(n5105) );
  NANDN U6723 ( .B(n240), .A(n5009), .Z(n5200) );
  NAND U6724 ( .A(n1056), .B(n163), .Z(n240) );
  AND U6725 ( .A(n5080), .B(n5203), .Z(n163) );
  AND U6726 ( .A(n4147), .B(n1939), .Z(n5080) );
  NAND U6727 ( .A(n5204), .B(n5205), .Z(\u_a23_mem/n18308 ) );
  OR U6728 ( .A(n271), .B(n4972), .Z(n5205) );
  NAND U6729 ( .A(n5206), .B(o[64]), .Z(n5204) );
  NAND U6730 ( .A(n5207), .B(n5208), .Z(\u_a23_mem/n18307 ) );
  OR U6731 ( .A(n271), .B(n4977), .Z(n5208) );
  NAND U6732 ( .A(n5206), .B(o[65]), .Z(n5207) );
  NAND U6733 ( .A(n5209), .B(n5210), .Z(\u_a23_mem/n18306 ) );
  OR U6734 ( .A(n271), .B(n4982), .Z(n5210) );
  NAND U6735 ( .A(n5206), .B(o[66]), .Z(n5209) );
  NAND U6736 ( .A(n5211), .B(n5212), .Z(\u_a23_mem/n18305 ) );
  OR U6737 ( .A(n271), .B(n4987), .Z(n5212) );
  NAND U6738 ( .A(n5206), .B(o[67]), .Z(n5211) );
  NAND U6739 ( .A(n5213), .B(n5214), .Z(\u_a23_mem/n18304 ) );
  OR U6740 ( .A(n271), .B(n4992), .Z(n5214) );
  NAND U6741 ( .A(n5206), .B(o[68]), .Z(n5213) );
  NAND U6742 ( .A(n5215), .B(n5216), .Z(\u_a23_mem/n18303 ) );
  OR U6743 ( .A(n271), .B(n4997), .Z(n5216) );
  NAND U6744 ( .A(n5206), .B(o[69]), .Z(n5215) );
  NAND U6745 ( .A(n5217), .B(n5218), .Z(\u_a23_mem/n18302 ) );
  OR U6746 ( .A(n271), .B(n5002), .Z(n5218) );
  NAND U6747 ( .A(n5206), .B(o[70]), .Z(n5217) );
  NAND U6748 ( .A(n5219), .B(n5220), .Z(\u_a23_mem/n18301 ) );
  NANDN U6749 ( .B(n271), .A(n5009), .Z(n5220) );
  NANDN U6750 ( .B(n2), .A(n287), .Z(n271) );
  NAND U6751 ( .A(n5206), .B(o[71]), .Z(n5219) );
  NANDN U6752 ( .B(n5099), .A(n287), .Z(n5206) );
  NAND U6753 ( .A(n5221), .B(n5222), .Z(\u_a23_mem/n18300 ) );
  NAND U6754 ( .A(n5223), .B(o[72]), .Z(n5222) );
  AND U6755 ( .A(n5224), .B(n5225), .Z(n5221) );
  NANDN U6756 ( .B(n5226), .A(n9), .Z(n5225) );
  OR U6757 ( .A(n294), .B(n4972), .Z(n5224) );
  NAND U6758 ( .A(n5227), .B(n5228), .Z(\u_a23_mem/n18299 ) );
  NAND U6759 ( .A(n5223), .B(o[73]), .Z(n5228) );
  AND U6760 ( .A(n5229), .B(n5230), .Z(n5227) );
  NANDN U6761 ( .B(n5226), .A(n16), .Z(n5230) );
  OR U6762 ( .A(n294), .B(n4977), .Z(n5229) );
  NAND U6763 ( .A(n5231), .B(n5232), .Z(\u_a23_mem/n18298 ) );
  NAND U6764 ( .A(n5223), .B(o[74]), .Z(n5232) );
  AND U6765 ( .A(n5233), .B(n5234), .Z(n5231) );
  NANDN U6766 ( .B(n5226), .A(n22), .Z(n5234) );
  OR U6767 ( .A(n294), .B(n4982), .Z(n5233) );
  NAND U6768 ( .A(n5235), .B(n5236), .Z(\u_a23_mem/n18297 ) );
  NAND U6769 ( .A(n5223), .B(o[75]), .Z(n5236) );
  AND U6770 ( .A(n5237), .B(n5238), .Z(n5235) );
  NANDN U6771 ( .B(n5226), .A(n28), .Z(n5238) );
  OR U6772 ( .A(n294), .B(n4987), .Z(n5237) );
  NAND U6773 ( .A(n5239), .B(n5240), .Z(\u_a23_mem/n18296 ) );
  NAND U6774 ( .A(n5223), .B(o[76]), .Z(n5240) );
  AND U6775 ( .A(n5241), .B(n5242), .Z(n5239) );
  NANDN U6776 ( .B(n5226), .A(n34), .Z(n5242) );
  OR U6777 ( .A(n294), .B(n4992), .Z(n5241) );
  NAND U6778 ( .A(n5243), .B(n5244), .Z(\u_a23_mem/n18295 ) );
  NAND U6779 ( .A(n5223), .B(o[77]), .Z(n5244) );
  AND U6780 ( .A(n5245), .B(n5246), .Z(n5243) );
  NANDN U6781 ( .B(n5226), .A(n40), .Z(n5246) );
  OR U6782 ( .A(n294), .B(n4997), .Z(n5245) );
  NAND U6783 ( .A(n5247), .B(n5248), .Z(\u_a23_mem/n18294 ) );
  NAND U6784 ( .A(n5223), .B(o[78]), .Z(n5248) );
  AND U6785 ( .A(n5249), .B(n5250), .Z(n5247) );
  NANDN U6786 ( .B(n5226), .A(n46), .Z(n5250) );
  OR U6787 ( .A(n294), .B(n5002), .Z(n5249) );
  NAND U6788 ( .A(n5251), .B(n5252), .Z(\u_a23_mem/n18293 ) );
  NAND U6789 ( .A(n5223), .B(o[79]), .Z(n5252) );
  NANDN U6790 ( .B(n5132), .A(n287), .Z(n5223) );
  AND U6791 ( .A(n5253), .B(n5254), .Z(n5251) );
  NANDN U6792 ( .B(n5226), .A(n53), .Z(n5254) );
  NANDN U6793 ( .B(n294), .A(n5009), .Z(n5253) );
  NAND U6794 ( .A(n1121), .B(n287), .Z(n294) );
  NAND U6795 ( .A(n5255), .B(n5256), .Z(\u_a23_mem/n18292 ) );
  NAND U6796 ( .A(n5257), .B(o[80]), .Z(n5256) );
  AND U6797 ( .A(n5258), .B(n5259), .Z(n5255) );
  NANDN U6798 ( .B(n5226), .A(n60), .Z(n5259) );
  OR U6799 ( .A(n328), .B(n4972), .Z(n5258) );
  NAND U6800 ( .A(n5260), .B(n5261), .Z(\u_a23_mem/n18291 ) );
  NAND U6801 ( .A(n5257), .B(o[81]), .Z(n5261) );
  AND U6802 ( .A(n5262), .B(n5263), .Z(n5260) );
  NANDN U6803 ( .B(n5226), .A(n66), .Z(n5263) );
  OR U6804 ( .A(n328), .B(n4977), .Z(n5262) );
  NAND U6805 ( .A(n5264), .B(n5265), .Z(\u_a23_mem/n18290 ) );
  NAND U6806 ( .A(n5257), .B(o[82]), .Z(n5265) );
  AND U6807 ( .A(n5266), .B(n5267), .Z(n5264) );
  NANDN U6808 ( .B(n5226), .A(n71), .Z(n5267) );
  OR U6809 ( .A(n328), .B(n4982), .Z(n5266) );
  NAND U6810 ( .A(n5268), .B(n5269), .Z(\u_a23_mem/n18289 ) );
  NAND U6811 ( .A(n5257), .B(o[83]), .Z(n5269) );
  AND U6812 ( .A(n5270), .B(n5271), .Z(n5268) );
  NANDN U6813 ( .B(n5226), .A(n76), .Z(n5271) );
  OR U6814 ( .A(n328), .B(n4987), .Z(n5270) );
  NAND U6815 ( .A(n5272), .B(n5273), .Z(\u_a23_mem/n18288 ) );
  NAND U6816 ( .A(n5257), .B(o[84]), .Z(n5273) );
  AND U6817 ( .A(n5274), .B(n5275), .Z(n5272) );
  NANDN U6818 ( .B(n5226), .A(n81), .Z(n5275) );
  OR U6819 ( .A(n328), .B(n4992), .Z(n5274) );
  NAND U6820 ( .A(n5276), .B(n5277), .Z(\u_a23_mem/n18287 ) );
  NAND U6821 ( .A(n5257), .B(o[85]), .Z(n5277) );
  AND U6822 ( .A(n5278), .B(n5279), .Z(n5276) );
  NANDN U6823 ( .B(n5226), .A(n86), .Z(n5279) );
  OR U6824 ( .A(n328), .B(n4997), .Z(n5278) );
  NAND U6825 ( .A(n5280), .B(n5281), .Z(\u_a23_mem/n18286 ) );
  NAND U6826 ( .A(n5257), .B(o[86]), .Z(n5281) );
  AND U6827 ( .A(n5282), .B(n5283), .Z(n5280) );
  NANDN U6828 ( .B(n5226), .A(n91), .Z(n5283) );
  OR U6829 ( .A(n328), .B(n5002), .Z(n5282) );
  NAND U6830 ( .A(n5284), .B(n5285), .Z(\u_a23_mem/n18285 ) );
  NAND U6831 ( .A(n5257), .B(o[87]), .Z(n5285) );
  NANDN U6832 ( .B(n5166), .A(n287), .Z(n5257) );
  AND U6833 ( .A(n5286), .B(n5287), .Z(n5284) );
  NANDN U6834 ( .B(n5226), .A(n98), .Z(n5287) );
  NANDN U6835 ( .B(n328), .A(n5009), .Z(n5286) );
  NAND U6836 ( .A(n1165), .B(n287), .Z(n328) );
  NAND U6837 ( .A(n5288), .B(n5289), .Z(\u_a23_mem/n18284 ) );
  NAND U6838 ( .A(n5290), .B(o[88]), .Z(n5289) );
  AND U6839 ( .A(n5291), .B(n5292), .Z(n5288) );
  NANDN U6840 ( .B(n5226), .A(n104), .Z(n5292) );
  OR U6841 ( .A(n362), .B(n4972), .Z(n5291) );
  NAND U6842 ( .A(n5293), .B(n5294), .Z(\u_a23_mem/n18283 ) );
  NAND U6843 ( .A(n5290), .B(o[89]), .Z(n5294) );
  AND U6844 ( .A(n5295), .B(n5296), .Z(n5293) );
  NANDN U6845 ( .B(n5226), .A(n110), .Z(n5296) );
  OR U6846 ( .A(n362), .B(n4977), .Z(n5295) );
  NAND U6847 ( .A(n5297), .B(n5298), .Z(\u_a23_mem/n18282 ) );
  NAND U6848 ( .A(n5290), .B(o[90]), .Z(n5298) );
  AND U6849 ( .A(n5299), .B(n5300), .Z(n5297) );
  NANDN U6850 ( .B(n5226), .A(n115), .Z(n5300) );
  OR U6851 ( .A(n362), .B(n4982), .Z(n5299) );
  NAND U6852 ( .A(n5301), .B(n5302), .Z(\u_a23_mem/n18281 ) );
  NAND U6853 ( .A(n5290), .B(o[91]), .Z(n5302) );
  AND U6854 ( .A(n5303), .B(n5304), .Z(n5301) );
  NANDN U6855 ( .B(n5226), .A(n120), .Z(n5304) );
  OR U6856 ( .A(n362), .B(n4987), .Z(n5303) );
  NAND U6857 ( .A(n5305), .B(n5306), .Z(\u_a23_mem/n18280 ) );
  NAND U6858 ( .A(n5290), .B(o[92]), .Z(n5306) );
  AND U6859 ( .A(n5307), .B(n5308), .Z(n5305) );
  NANDN U6860 ( .B(n5226), .A(n125), .Z(n5308) );
  OR U6861 ( .A(n362), .B(n4992), .Z(n5307) );
  NAND U6862 ( .A(n5309), .B(n5310), .Z(\u_a23_mem/n18279 ) );
  NAND U6863 ( .A(n5290), .B(o[93]), .Z(n5310) );
  AND U6864 ( .A(n5311), .B(n5312), .Z(n5309) );
  NANDN U6865 ( .B(n5226), .A(n130), .Z(n5312) );
  OR U6866 ( .A(n362), .B(n4997), .Z(n5311) );
  NAND U6867 ( .A(n5313), .B(n5314), .Z(\u_a23_mem/n18278 ) );
  NAND U6868 ( .A(n5290), .B(o[94]), .Z(n5314) );
  AND U6869 ( .A(n5315), .B(n5316), .Z(n5313) );
  NANDN U6870 ( .B(n5226), .A(n135), .Z(n5316) );
  OR U6871 ( .A(n362), .B(n5002), .Z(n5315) );
  NAND U6872 ( .A(n5317), .B(n5318), .Z(\u_a23_mem/n18277 ) );
  NAND U6873 ( .A(n5290), .B(o[95]), .Z(n5318) );
  NAND U6874 ( .A(n287), .B(n5077), .Z(n5290) );
  AND U6875 ( .A(n5319), .B(n5320), .Z(n5317) );
  NANDN U6876 ( .B(n5226), .A(n142), .Z(n5320) );
  NAND U6877 ( .A(n5202), .B(n287), .Z(n5226) );
  NANDN U6878 ( .B(n362), .A(n5009), .Z(n5319) );
  NAND U6879 ( .A(n1056), .B(n287), .Z(n362) );
  ANDN U6880 ( .A(n5321), .B(n4147), .Z(n287) );
  AND U6881 ( .A(n5081), .B(n1939), .Z(n5321) );
  NAND U6882 ( .A(n5322), .B(n5323), .Z(\u_a23_mem/n18276 ) );
  OR U6883 ( .A(n393), .B(n4972), .Z(n5323) );
  NAND U6884 ( .A(n5324), .B(o[96]), .Z(n5322) );
  NAND U6885 ( .A(n5325), .B(n5326), .Z(\u_a23_mem/n18275 ) );
  OR U6886 ( .A(n393), .B(n4977), .Z(n5326) );
  NAND U6887 ( .A(n5324), .B(o[97]), .Z(n5325) );
  NAND U6888 ( .A(n5327), .B(n5328), .Z(\u_a23_mem/n18274 ) );
  OR U6889 ( .A(n393), .B(n4982), .Z(n5328) );
  NAND U6890 ( .A(n5324), .B(o[98]), .Z(n5327) );
  NAND U6891 ( .A(n5329), .B(n5330), .Z(\u_a23_mem/n18273 ) );
  OR U6892 ( .A(n393), .B(n4987), .Z(n5330) );
  NAND U6893 ( .A(n5324), .B(o[99]), .Z(n5329) );
  NAND U6894 ( .A(n5331), .B(n5332), .Z(\u_a23_mem/n18272 ) );
  OR U6895 ( .A(n393), .B(n4992), .Z(n5332) );
  NAND U6896 ( .A(n5324), .B(o[100]), .Z(n5331) );
  NAND U6897 ( .A(n5333), .B(n5334), .Z(\u_a23_mem/n18271 ) );
  OR U6898 ( .A(n393), .B(n4997), .Z(n5334) );
  NAND U6899 ( .A(n5324), .B(o[101]), .Z(n5333) );
  NAND U6900 ( .A(n5335), .B(n5336), .Z(\u_a23_mem/n18270 ) );
  OR U6901 ( .A(n393), .B(n5002), .Z(n5336) );
  NAND U6902 ( .A(n5324), .B(o[102]), .Z(n5335) );
  NAND U6903 ( .A(n5337), .B(n5338), .Z(\u_a23_mem/n18269 ) );
  NANDN U6904 ( .B(n393), .A(n5009), .Z(n5338) );
  NANDN U6905 ( .B(n2), .A(n409), .Z(n393) );
  NAND U6906 ( .A(n5324), .B(o[103]), .Z(n5337) );
  NANDN U6907 ( .B(n5099), .A(n409), .Z(n5324) );
  NAND U6908 ( .A(n5339), .B(n5340), .Z(\u_a23_mem/n18268 ) );
  NAND U6909 ( .A(n5341), .B(o[104]), .Z(n5340) );
  AND U6910 ( .A(n5342), .B(n5343), .Z(n5339) );
  NANDN U6911 ( .B(n5344), .A(n9), .Z(n5343) );
  OR U6912 ( .A(n416), .B(n4972), .Z(n5342) );
  NAND U6913 ( .A(n5345), .B(n5346), .Z(\u_a23_mem/n18267 ) );
  NAND U6914 ( .A(n5341), .B(o[105]), .Z(n5346) );
  AND U6915 ( .A(n5347), .B(n5348), .Z(n5345) );
  NANDN U6916 ( .B(n5344), .A(n16), .Z(n5348) );
  OR U6917 ( .A(n416), .B(n4977), .Z(n5347) );
  NAND U6918 ( .A(n5349), .B(n5350), .Z(\u_a23_mem/n18266 ) );
  NAND U6919 ( .A(n5341), .B(o[106]), .Z(n5350) );
  AND U6920 ( .A(n5351), .B(n5352), .Z(n5349) );
  NANDN U6921 ( .B(n5344), .A(n22), .Z(n5352) );
  OR U6922 ( .A(n416), .B(n4982), .Z(n5351) );
  NAND U6923 ( .A(n5353), .B(n5354), .Z(\u_a23_mem/n18265 ) );
  NAND U6924 ( .A(n5341), .B(o[107]), .Z(n5354) );
  AND U6925 ( .A(n5355), .B(n5356), .Z(n5353) );
  NANDN U6926 ( .B(n5344), .A(n28), .Z(n5356) );
  OR U6927 ( .A(n416), .B(n4987), .Z(n5355) );
  NAND U6928 ( .A(n5357), .B(n5358), .Z(\u_a23_mem/n18264 ) );
  NAND U6929 ( .A(n5341), .B(o[108]), .Z(n5358) );
  AND U6930 ( .A(n5359), .B(n5360), .Z(n5357) );
  NANDN U6931 ( .B(n5344), .A(n34), .Z(n5360) );
  OR U6932 ( .A(n416), .B(n4992), .Z(n5359) );
  NAND U6933 ( .A(n5361), .B(n5362), .Z(\u_a23_mem/n18263 ) );
  NAND U6934 ( .A(n5341), .B(o[109]), .Z(n5362) );
  AND U6935 ( .A(n5363), .B(n5364), .Z(n5361) );
  NANDN U6936 ( .B(n5344), .A(n40), .Z(n5364) );
  OR U6937 ( .A(n416), .B(n4997), .Z(n5363) );
  NAND U6938 ( .A(n5365), .B(n5366), .Z(\u_a23_mem/n18262 ) );
  NAND U6939 ( .A(n5341), .B(o[110]), .Z(n5366) );
  AND U6940 ( .A(n5367), .B(n5368), .Z(n5365) );
  NANDN U6941 ( .B(n5344), .A(n46), .Z(n5368) );
  OR U6942 ( .A(n416), .B(n5002), .Z(n5367) );
  NAND U6943 ( .A(n5369), .B(n5370), .Z(\u_a23_mem/n18261 ) );
  NAND U6944 ( .A(n5341), .B(o[111]), .Z(n5370) );
  NANDN U6945 ( .B(n5132), .A(n409), .Z(n5341) );
  AND U6946 ( .A(n5371), .B(n5372), .Z(n5369) );
  NANDN U6947 ( .B(n5344), .A(n53), .Z(n5372) );
  NANDN U6948 ( .B(n416), .A(n5009), .Z(n5371) );
  NAND U6949 ( .A(n1121), .B(n409), .Z(n416) );
  NAND U6950 ( .A(n5373), .B(n5374), .Z(\u_a23_mem/n18260 ) );
  NAND U6951 ( .A(n5375), .B(o[112]), .Z(n5374) );
  AND U6952 ( .A(n5376), .B(n5377), .Z(n5373) );
  NANDN U6953 ( .B(n5344), .A(n60), .Z(n5377) );
  OR U6954 ( .A(n450), .B(n4972), .Z(n5376) );
  NAND U6955 ( .A(n5378), .B(n5379), .Z(\u_a23_mem/n18259 ) );
  NAND U6956 ( .A(n5375), .B(o[113]), .Z(n5379) );
  AND U6957 ( .A(n5380), .B(n5381), .Z(n5378) );
  NANDN U6958 ( .B(n5344), .A(n66), .Z(n5381) );
  OR U6959 ( .A(n450), .B(n4977), .Z(n5380) );
  NAND U6960 ( .A(n5382), .B(n5383), .Z(\u_a23_mem/n18258 ) );
  NAND U6961 ( .A(n5375), .B(o[114]), .Z(n5383) );
  AND U6962 ( .A(n5384), .B(n5385), .Z(n5382) );
  NANDN U6963 ( .B(n5344), .A(n71), .Z(n5385) );
  OR U6964 ( .A(n450), .B(n4982), .Z(n5384) );
  NAND U6965 ( .A(n5386), .B(n5387), .Z(\u_a23_mem/n18257 ) );
  NAND U6966 ( .A(n5375), .B(o[115]), .Z(n5387) );
  AND U6967 ( .A(n5388), .B(n5389), .Z(n5386) );
  NANDN U6968 ( .B(n5344), .A(n76), .Z(n5389) );
  OR U6969 ( .A(n450), .B(n4987), .Z(n5388) );
  NAND U6970 ( .A(n5390), .B(n5391), .Z(\u_a23_mem/n18256 ) );
  NAND U6971 ( .A(n5375), .B(o[116]), .Z(n5391) );
  AND U6972 ( .A(n5392), .B(n5393), .Z(n5390) );
  NANDN U6973 ( .B(n5344), .A(n81), .Z(n5393) );
  OR U6974 ( .A(n450), .B(n4992), .Z(n5392) );
  NAND U6975 ( .A(n5394), .B(n5395), .Z(\u_a23_mem/n18255 ) );
  NAND U6976 ( .A(n5375), .B(o[117]), .Z(n5395) );
  AND U6977 ( .A(n5396), .B(n5397), .Z(n5394) );
  NANDN U6978 ( .B(n5344), .A(n86), .Z(n5397) );
  OR U6979 ( .A(n450), .B(n4997), .Z(n5396) );
  NAND U6980 ( .A(n5398), .B(n5399), .Z(\u_a23_mem/n18254 ) );
  NAND U6981 ( .A(n5375), .B(o[118]), .Z(n5399) );
  AND U6982 ( .A(n5400), .B(n5401), .Z(n5398) );
  NANDN U6983 ( .B(n5344), .A(n91), .Z(n5401) );
  OR U6984 ( .A(n450), .B(n5002), .Z(n5400) );
  NAND U6985 ( .A(n5402), .B(n5403), .Z(\u_a23_mem/n18253 ) );
  NAND U6986 ( .A(n5375), .B(o[119]), .Z(n5403) );
  NANDN U6987 ( .B(n5166), .A(n409), .Z(n5375) );
  AND U6988 ( .A(n5404), .B(n5405), .Z(n5402) );
  NANDN U6989 ( .B(n5344), .A(n98), .Z(n5405) );
  NANDN U6990 ( .B(n450), .A(n5009), .Z(n5404) );
  NAND U6991 ( .A(n1165), .B(n409), .Z(n450) );
  NAND U6992 ( .A(n5406), .B(n5407), .Z(\u_a23_mem/n18252 ) );
  NAND U6993 ( .A(n5408), .B(o[120]), .Z(n5407) );
  AND U6994 ( .A(n5409), .B(n5410), .Z(n5406) );
  NANDN U6995 ( .B(n5344), .A(n104), .Z(n5410) );
  OR U6996 ( .A(n484), .B(n4972), .Z(n5409) );
  NAND U6997 ( .A(n5411), .B(n5412), .Z(\u_a23_mem/n18251 ) );
  NAND U6998 ( .A(n5408), .B(o[121]), .Z(n5412) );
  AND U6999 ( .A(n5413), .B(n5414), .Z(n5411) );
  NANDN U7000 ( .B(n5344), .A(n110), .Z(n5414) );
  OR U7001 ( .A(n484), .B(n4977), .Z(n5413) );
  NAND U7002 ( .A(n5415), .B(n5416), .Z(\u_a23_mem/n18250 ) );
  NAND U7003 ( .A(n5408), .B(o[122]), .Z(n5416) );
  AND U7004 ( .A(n5417), .B(n5418), .Z(n5415) );
  NANDN U7005 ( .B(n5344), .A(n115), .Z(n5418) );
  OR U7006 ( .A(n484), .B(n4982), .Z(n5417) );
  NAND U7007 ( .A(n5419), .B(n5420), .Z(\u_a23_mem/n18249 ) );
  NAND U7008 ( .A(n5408), .B(o[123]), .Z(n5420) );
  AND U7009 ( .A(n5421), .B(n5422), .Z(n5419) );
  NANDN U7010 ( .B(n5344), .A(n120), .Z(n5422) );
  OR U7011 ( .A(n484), .B(n4987), .Z(n5421) );
  NAND U7012 ( .A(n5423), .B(n5424), .Z(\u_a23_mem/n18248 ) );
  NAND U7013 ( .A(n5408), .B(o[124]), .Z(n5424) );
  AND U7014 ( .A(n5425), .B(n5426), .Z(n5423) );
  NANDN U7015 ( .B(n5344), .A(n125), .Z(n5426) );
  OR U7016 ( .A(n484), .B(n4992), .Z(n5425) );
  NAND U7017 ( .A(n5427), .B(n5428), .Z(\u_a23_mem/n18247 ) );
  NAND U7018 ( .A(n5408), .B(o[125]), .Z(n5428) );
  AND U7019 ( .A(n5429), .B(n5430), .Z(n5427) );
  NANDN U7020 ( .B(n5344), .A(n130), .Z(n5430) );
  OR U7021 ( .A(n484), .B(n4997), .Z(n5429) );
  NAND U7022 ( .A(n5431), .B(n5432), .Z(\u_a23_mem/n18246 ) );
  NAND U7023 ( .A(n5408), .B(o[126]), .Z(n5432) );
  AND U7024 ( .A(n5433), .B(n5434), .Z(n5431) );
  NANDN U7025 ( .B(n5344), .A(n135), .Z(n5434) );
  OR U7026 ( .A(n484), .B(n5002), .Z(n5433) );
  NAND U7027 ( .A(n5435), .B(n5436), .Z(\u_a23_mem/n18245 ) );
  NAND U7028 ( .A(n5408), .B(o[127]), .Z(n5436) );
  NAND U7029 ( .A(n409), .B(n5077), .Z(n5408) );
  AND U7030 ( .A(n5437), .B(n5438), .Z(n5435) );
  NANDN U7031 ( .B(n5344), .A(n142), .Z(n5438) );
  NAND U7032 ( .A(n5202), .B(n409), .Z(n5344) );
  NANDN U7033 ( .B(n484), .A(n5009), .Z(n5437) );
  NAND U7034 ( .A(n1056), .B(n409), .Z(n484) );
  ANDN U7035 ( .A(n5439), .B(n4147), .Z(n409) );
  AND U7036 ( .A(n5203), .B(n1939), .Z(n5439) );
  NAND U7037 ( .A(n5440), .B(n5441), .Z(\u_a23_mem/n18244 ) );
  OR U7038 ( .A(n515), .B(n4972), .Z(n5441) );
  NAND U7039 ( .A(n5442), .B(o[128]), .Z(n5440) );
  NAND U7040 ( .A(n5443), .B(n5444), .Z(\u_a23_mem/n18243 ) );
  OR U7041 ( .A(n515), .B(n4977), .Z(n5444) );
  NAND U7042 ( .A(n5442), .B(o[129]), .Z(n5443) );
  NAND U7043 ( .A(n5445), .B(n5446), .Z(\u_a23_mem/n18242 ) );
  OR U7044 ( .A(n515), .B(n4982), .Z(n5446) );
  NAND U7045 ( .A(n5442), .B(o[130]), .Z(n5445) );
  NAND U7046 ( .A(n5447), .B(n5448), .Z(\u_a23_mem/n18241 ) );
  OR U7047 ( .A(n515), .B(n4987), .Z(n5448) );
  NAND U7048 ( .A(n5442), .B(o[131]), .Z(n5447) );
  NAND U7049 ( .A(n5449), .B(n5450), .Z(\u_a23_mem/n18240 ) );
  OR U7050 ( .A(n515), .B(n4992), .Z(n5450) );
  NAND U7051 ( .A(n5442), .B(o[132]), .Z(n5449) );
  NAND U7052 ( .A(n5451), .B(n5452), .Z(\u_a23_mem/n18239 ) );
  OR U7053 ( .A(n515), .B(n4997), .Z(n5452) );
  NAND U7054 ( .A(n5442), .B(o[133]), .Z(n5451) );
  NAND U7055 ( .A(n5453), .B(n5454), .Z(\u_a23_mem/n18238 ) );
  OR U7056 ( .A(n515), .B(n5002), .Z(n5454) );
  NAND U7057 ( .A(n5442), .B(o[134]), .Z(n5453) );
  NAND U7058 ( .A(n5455), .B(n5456), .Z(\u_a23_mem/n18237 ) );
  NANDN U7059 ( .B(n515), .A(n5009), .Z(n5456) );
  NANDN U7060 ( .B(n2), .A(n531), .Z(n515) );
  NAND U7061 ( .A(n5442), .B(o[135]), .Z(n5455) );
  NANDN U7062 ( .B(n5099), .A(n531), .Z(n5442) );
  NAND U7063 ( .A(n5457), .B(n5458), .Z(\u_a23_mem/n18236 ) );
  NAND U7064 ( .A(n5459), .B(o[136]), .Z(n5458) );
  AND U7065 ( .A(n5460), .B(n5461), .Z(n5457) );
  NANDN U7066 ( .B(n5462), .A(n9), .Z(n5461) );
  OR U7067 ( .A(n538), .B(n4972), .Z(n5460) );
  NAND U7068 ( .A(n5463), .B(n5464), .Z(\u_a23_mem/n18235 ) );
  NAND U7069 ( .A(n5459), .B(o[137]), .Z(n5464) );
  AND U7070 ( .A(n5465), .B(n5466), .Z(n5463) );
  NANDN U7071 ( .B(n5462), .A(n16), .Z(n5466) );
  OR U7072 ( .A(n538), .B(n4977), .Z(n5465) );
  NAND U7073 ( .A(n5467), .B(n5468), .Z(\u_a23_mem/n18234 ) );
  NAND U7074 ( .A(n5459), .B(o[138]), .Z(n5468) );
  AND U7075 ( .A(n5469), .B(n5470), .Z(n5467) );
  NANDN U7076 ( .B(n5462), .A(n22), .Z(n5470) );
  OR U7077 ( .A(n538), .B(n4982), .Z(n5469) );
  NAND U7078 ( .A(n5471), .B(n5472), .Z(\u_a23_mem/n18233 ) );
  NAND U7079 ( .A(n5459), .B(o[139]), .Z(n5472) );
  AND U7080 ( .A(n5473), .B(n5474), .Z(n5471) );
  NANDN U7081 ( .B(n5462), .A(n28), .Z(n5474) );
  OR U7082 ( .A(n538), .B(n4987), .Z(n5473) );
  NAND U7083 ( .A(n5475), .B(n5476), .Z(\u_a23_mem/n18232 ) );
  NAND U7084 ( .A(n5459), .B(o[140]), .Z(n5476) );
  AND U7085 ( .A(n5477), .B(n5478), .Z(n5475) );
  NANDN U7086 ( .B(n5462), .A(n34), .Z(n5478) );
  OR U7087 ( .A(n538), .B(n4992), .Z(n5477) );
  NAND U7088 ( .A(n5479), .B(n5480), .Z(\u_a23_mem/n18231 ) );
  NAND U7089 ( .A(n5459), .B(o[141]), .Z(n5480) );
  AND U7090 ( .A(n5481), .B(n5482), .Z(n5479) );
  NANDN U7091 ( .B(n5462), .A(n40), .Z(n5482) );
  OR U7092 ( .A(n538), .B(n4997), .Z(n5481) );
  NAND U7093 ( .A(n5483), .B(n5484), .Z(\u_a23_mem/n18230 ) );
  NAND U7094 ( .A(n5459), .B(o[142]), .Z(n5484) );
  AND U7095 ( .A(n5485), .B(n5486), .Z(n5483) );
  NANDN U7096 ( .B(n5462), .A(n46), .Z(n5486) );
  OR U7097 ( .A(n538), .B(n5002), .Z(n5485) );
  NAND U7098 ( .A(n5487), .B(n5488), .Z(\u_a23_mem/n18229 ) );
  NAND U7099 ( .A(n5459), .B(o[143]), .Z(n5488) );
  NANDN U7100 ( .B(n5132), .A(n531), .Z(n5459) );
  AND U7101 ( .A(n5489), .B(n5490), .Z(n5487) );
  NANDN U7102 ( .B(n5462), .A(n53), .Z(n5490) );
  NANDN U7103 ( .B(n538), .A(n5009), .Z(n5489) );
  NAND U7104 ( .A(n1121), .B(n531), .Z(n538) );
  NAND U7105 ( .A(n5491), .B(n5492), .Z(\u_a23_mem/n18228 ) );
  NAND U7106 ( .A(n5493), .B(o[144]), .Z(n5492) );
  AND U7107 ( .A(n5494), .B(n5495), .Z(n5491) );
  NANDN U7108 ( .B(n5462), .A(n60), .Z(n5495) );
  OR U7109 ( .A(n572), .B(n4972), .Z(n5494) );
  NAND U7110 ( .A(n5496), .B(n5497), .Z(\u_a23_mem/n18227 ) );
  NAND U7111 ( .A(n5493), .B(o[145]), .Z(n5497) );
  AND U7112 ( .A(n5498), .B(n5499), .Z(n5496) );
  NANDN U7113 ( .B(n5462), .A(n66), .Z(n5499) );
  OR U7114 ( .A(n572), .B(n4977), .Z(n5498) );
  NAND U7115 ( .A(n5500), .B(n5501), .Z(\u_a23_mem/n18226 ) );
  NAND U7116 ( .A(n5493), .B(o[146]), .Z(n5501) );
  AND U7117 ( .A(n5502), .B(n5503), .Z(n5500) );
  NANDN U7118 ( .B(n5462), .A(n71), .Z(n5503) );
  OR U7119 ( .A(n572), .B(n4982), .Z(n5502) );
  NAND U7120 ( .A(n5504), .B(n5505), .Z(\u_a23_mem/n18225 ) );
  NAND U7121 ( .A(n5493), .B(o[147]), .Z(n5505) );
  AND U7122 ( .A(n5506), .B(n5507), .Z(n5504) );
  NANDN U7123 ( .B(n5462), .A(n76), .Z(n5507) );
  OR U7124 ( .A(n572), .B(n4987), .Z(n5506) );
  NAND U7125 ( .A(n5508), .B(n5509), .Z(\u_a23_mem/n18224 ) );
  NAND U7126 ( .A(n5493), .B(o[148]), .Z(n5509) );
  AND U7127 ( .A(n5510), .B(n5511), .Z(n5508) );
  NANDN U7128 ( .B(n5462), .A(n81), .Z(n5511) );
  OR U7129 ( .A(n572), .B(n4992), .Z(n5510) );
  NAND U7130 ( .A(n5512), .B(n5513), .Z(\u_a23_mem/n18223 ) );
  NAND U7131 ( .A(n5493), .B(o[149]), .Z(n5513) );
  AND U7132 ( .A(n5514), .B(n5515), .Z(n5512) );
  NANDN U7133 ( .B(n5462), .A(n86), .Z(n5515) );
  OR U7134 ( .A(n572), .B(n4997), .Z(n5514) );
  NAND U7135 ( .A(n5516), .B(n5517), .Z(\u_a23_mem/n18222 ) );
  NAND U7136 ( .A(n5493), .B(o[150]), .Z(n5517) );
  AND U7137 ( .A(n5518), .B(n5519), .Z(n5516) );
  NANDN U7138 ( .B(n5462), .A(n91), .Z(n5519) );
  OR U7139 ( .A(n572), .B(n5002), .Z(n5518) );
  NAND U7140 ( .A(n5520), .B(n5521), .Z(\u_a23_mem/n18221 ) );
  NAND U7141 ( .A(n5493), .B(o[151]), .Z(n5521) );
  NANDN U7142 ( .B(n5166), .A(n531), .Z(n5493) );
  AND U7143 ( .A(n5522), .B(n5523), .Z(n5520) );
  NANDN U7144 ( .B(n5462), .A(n98), .Z(n5523) );
  NANDN U7145 ( .B(n572), .A(n5009), .Z(n5522) );
  NAND U7146 ( .A(n1165), .B(n531), .Z(n572) );
  NAND U7147 ( .A(n5524), .B(n5525), .Z(\u_a23_mem/n18220 ) );
  NAND U7148 ( .A(n5526), .B(o[152]), .Z(n5525) );
  AND U7149 ( .A(n5527), .B(n5528), .Z(n5524) );
  NANDN U7150 ( .B(n5462), .A(n104), .Z(n5528) );
  OR U7151 ( .A(n606), .B(n4972), .Z(n5527) );
  NAND U7152 ( .A(n5529), .B(n5530), .Z(\u_a23_mem/n18219 ) );
  NAND U7153 ( .A(n5526), .B(o[153]), .Z(n5530) );
  AND U7154 ( .A(n5531), .B(n5532), .Z(n5529) );
  NANDN U7155 ( .B(n5462), .A(n110), .Z(n5532) );
  OR U7156 ( .A(n606), .B(n4977), .Z(n5531) );
  NAND U7157 ( .A(n5533), .B(n5534), .Z(\u_a23_mem/n18218 ) );
  NAND U7158 ( .A(n5526), .B(o[154]), .Z(n5534) );
  AND U7159 ( .A(n5535), .B(n5536), .Z(n5533) );
  NANDN U7160 ( .B(n5462), .A(n115), .Z(n5536) );
  OR U7161 ( .A(n606), .B(n4982), .Z(n5535) );
  NAND U7162 ( .A(n5537), .B(n5538), .Z(\u_a23_mem/n18217 ) );
  NAND U7163 ( .A(n5526), .B(o[155]), .Z(n5538) );
  AND U7164 ( .A(n5539), .B(n5540), .Z(n5537) );
  NANDN U7165 ( .B(n5462), .A(n120), .Z(n5540) );
  OR U7166 ( .A(n606), .B(n4987), .Z(n5539) );
  NAND U7167 ( .A(n5541), .B(n5542), .Z(\u_a23_mem/n18216 ) );
  NAND U7168 ( .A(n5526), .B(o[156]), .Z(n5542) );
  AND U7169 ( .A(n5543), .B(n5544), .Z(n5541) );
  NANDN U7170 ( .B(n5462), .A(n125), .Z(n5544) );
  OR U7171 ( .A(n606), .B(n4992), .Z(n5543) );
  NAND U7172 ( .A(n5545), .B(n5546), .Z(\u_a23_mem/n18215 ) );
  NAND U7173 ( .A(n5526), .B(o[157]), .Z(n5546) );
  AND U7174 ( .A(n5547), .B(n5548), .Z(n5545) );
  NANDN U7175 ( .B(n5462), .A(n130), .Z(n5548) );
  OR U7176 ( .A(n606), .B(n4997), .Z(n5547) );
  NAND U7177 ( .A(n5549), .B(n5550), .Z(\u_a23_mem/n18214 ) );
  NAND U7178 ( .A(n5526), .B(o[158]), .Z(n5550) );
  AND U7179 ( .A(n5551), .B(n5552), .Z(n5549) );
  NANDN U7180 ( .B(n5462), .A(n135), .Z(n5552) );
  OR U7181 ( .A(n606), .B(n5002), .Z(n5551) );
  NAND U7182 ( .A(n5553), .B(n5554), .Z(\u_a23_mem/n18213 ) );
  NAND U7183 ( .A(n5526), .B(o[159]), .Z(n5554) );
  NAND U7184 ( .A(n531), .B(n5077), .Z(n5526) );
  AND U7185 ( .A(n5555), .B(n5556), .Z(n5553) );
  NANDN U7186 ( .B(n5462), .A(n142), .Z(n5556) );
  NAND U7187 ( .A(n5202), .B(n531), .Z(n5462) );
  NANDN U7188 ( .B(n606), .A(n5009), .Z(n5555) );
  NAND U7189 ( .A(n1056), .B(n531), .Z(n606) );
  ANDN U7190 ( .A(n5557), .B(n1939), .Z(n531) );
  AND U7191 ( .A(n5081), .B(n4147), .Z(n5557) );
  NAND U7192 ( .A(n5558), .B(n5559), .Z(\u_a23_mem/n18212 ) );
  OR U7193 ( .A(n637), .B(n4972), .Z(n5559) );
  NAND U7194 ( .A(n5560), .B(o[160]), .Z(n5558) );
  NAND U7195 ( .A(n5561), .B(n5562), .Z(\u_a23_mem/n18211 ) );
  OR U7196 ( .A(n637), .B(n4977), .Z(n5562) );
  NAND U7197 ( .A(n5560), .B(o[161]), .Z(n5561) );
  NAND U7198 ( .A(n5563), .B(n5564), .Z(\u_a23_mem/n18210 ) );
  OR U7199 ( .A(n637), .B(n4982), .Z(n5564) );
  NAND U7200 ( .A(n5560), .B(o[162]), .Z(n5563) );
  NAND U7201 ( .A(n5565), .B(n5566), .Z(\u_a23_mem/n18209 ) );
  OR U7202 ( .A(n637), .B(n4987), .Z(n5566) );
  NAND U7203 ( .A(n5560), .B(o[163]), .Z(n5565) );
  NAND U7204 ( .A(n5567), .B(n5568), .Z(\u_a23_mem/n18208 ) );
  OR U7205 ( .A(n637), .B(n4992), .Z(n5568) );
  NAND U7206 ( .A(n5560), .B(o[164]), .Z(n5567) );
  NAND U7207 ( .A(n5569), .B(n5570), .Z(\u_a23_mem/n18207 ) );
  OR U7208 ( .A(n637), .B(n4997), .Z(n5570) );
  NAND U7209 ( .A(n5560), .B(o[165]), .Z(n5569) );
  NAND U7210 ( .A(n5571), .B(n5572), .Z(\u_a23_mem/n18206 ) );
  OR U7211 ( .A(n637), .B(n5002), .Z(n5572) );
  NAND U7212 ( .A(n5560), .B(o[166]), .Z(n5571) );
  NAND U7213 ( .A(n5573), .B(n5574), .Z(\u_a23_mem/n18205 ) );
  NANDN U7214 ( .B(n637), .A(n5009), .Z(n5574) );
  NANDN U7215 ( .B(n2), .A(n653), .Z(n637) );
  NAND U7216 ( .A(n5560), .B(o[167]), .Z(n5573) );
  NANDN U7217 ( .B(n5099), .A(n653), .Z(n5560) );
  NAND U7218 ( .A(n5575), .B(n5576), .Z(\u_a23_mem/n18204 ) );
  NAND U7219 ( .A(n5577), .B(o[168]), .Z(n5576) );
  AND U7220 ( .A(n5578), .B(n5579), .Z(n5575) );
  NANDN U7221 ( .B(n5580), .A(n9), .Z(n5579) );
  OR U7222 ( .A(n660), .B(n4972), .Z(n5578) );
  NAND U7223 ( .A(n5581), .B(n5582), .Z(\u_a23_mem/n18203 ) );
  NAND U7224 ( .A(n5577), .B(o[169]), .Z(n5582) );
  AND U7225 ( .A(n5583), .B(n5584), .Z(n5581) );
  NANDN U7226 ( .B(n5580), .A(n16), .Z(n5584) );
  OR U7227 ( .A(n660), .B(n4977), .Z(n5583) );
  NAND U7228 ( .A(n5585), .B(n5586), .Z(\u_a23_mem/n18202 ) );
  NAND U7229 ( .A(n5577), .B(o[170]), .Z(n5586) );
  AND U7230 ( .A(n5587), .B(n5588), .Z(n5585) );
  NANDN U7231 ( .B(n5580), .A(n22), .Z(n5588) );
  OR U7232 ( .A(n660), .B(n4982), .Z(n5587) );
  NAND U7233 ( .A(n5589), .B(n5590), .Z(\u_a23_mem/n18201 ) );
  NAND U7234 ( .A(n5577), .B(o[171]), .Z(n5590) );
  AND U7235 ( .A(n5591), .B(n5592), .Z(n5589) );
  NANDN U7236 ( .B(n5580), .A(n28), .Z(n5592) );
  OR U7237 ( .A(n660), .B(n4987), .Z(n5591) );
  NAND U7238 ( .A(n5593), .B(n5594), .Z(\u_a23_mem/n18200 ) );
  NAND U7239 ( .A(n5577), .B(o[172]), .Z(n5594) );
  AND U7240 ( .A(n5595), .B(n5596), .Z(n5593) );
  NANDN U7241 ( .B(n5580), .A(n34), .Z(n5596) );
  OR U7242 ( .A(n660), .B(n4992), .Z(n5595) );
  NAND U7243 ( .A(n5597), .B(n5598), .Z(\u_a23_mem/n18199 ) );
  NAND U7244 ( .A(n5577), .B(o[173]), .Z(n5598) );
  AND U7245 ( .A(n5599), .B(n5600), .Z(n5597) );
  NANDN U7246 ( .B(n5580), .A(n40), .Z(n5600) );
  OR U7247 ( .A(n660), .B(n4997), .Z(n5599) );
  NAND U7248 ( .A(n5601), .B(n5602), .Z(\u_a23_mem/n18198 ) );
  NAND U7249 ( .A(n5577), .B(o[174]), .Z(n5602) );
  AND U7250 ( .A(n5603), .B(n5604), .Z(n5601) );
  NANDN U7251 ( .B(n5580), .A(n46), .Z(n5604) );
  OR U7252 ( .A(n660), .B(n5002), .Z(n5603) );
  NAND U7253 ( .A(n5605), .B(n5606), .Z(\u_a23_mem/n18197 ) );
  NAND U7254 ( .A(n5577), .B(o[175]), .Z(n5606) );
  NANDN U7255 ( .B(n5132), .A(n653), .Z(n5577) );
  AND U7256 ( .A(n5607), .B(n5608), .Z(n5605) );
  NANDN U7257 ( .B(n5580), .A(n53), .Z(n5608) );
  NANDN U7258 ( .B(n660), .A(n5009), .Z(n5607) );
  NAND U7259 ( .A(n1121), .B(n653), .Z(n660) );
  NAND U7260 ( .A(n5609), .B(n5610), .Z(\u_a23_mem/n18196 ) );
  NAND U7261 ( .A(n5611), .B(o[176]), .Z(n5610) );
  AND U7262 ( .A(n5612), .B(n5613), .Z(n5609) );
  NANDN U7263 ( .B(n5580), .A(n60), .Z(n5613) );
  OR U7264 ( .A(n694), .B(n4972), .Z(n5612) );
  NAND U7265 ( .A(n5614), .B(n5615), .Z(\u_a23_mem/n18195 ) );
  NAND U7266 ( .A(n5611), .B(o[177]), .Z(n5615) );
  AND U7267 ( .A(n5616), .B(n5617), .Z(n5614) );
  NANDN U7268 ( .B(n5580), .A(n66), .Z(n5617) );
  OR U7269 ( .A(n694), .B(n4977), .Z(n5616) );
  NAND U7270 ( .A(n5618), .B(n5619), .Z(\u_a23_mem/n18194 ) );
  NAND U7271 ( .A(n5611), .B(o[178]), .Z(n5619) );
  AND U7272 ( .A(n5620), .B(n5621), .Z(n5618) );
  NANDN U7273 ( .B(n5580), .A(n71), .Z(n5621) );
  OR U7274 ( .A(n694), .B(n4982), .Z(n5620) );
  NAND U7275 ( .A(n5622), .B(n5623), .Z(\u_a23_mem/n18193 ) );
  NAND U7276 ( .A(n5611), .B(o[179]), .Z(n5623) );
  AND U7277 ( .A(n5624), .B(n5625), .Z(n5622) );
  NANDN U7278 ( .B(n5580), .A(n76), .Z(n5625) );
  OR U7279 ( .A(n694), .B(n4987), .Z(n5624) );
  NAND U7280 ( .A(n5626), .B(n5627), .Z(\u_a23_mem/n18192 ) );
  NAND U7281 ( .A(n5611), .B(o[180]), .Z(n5627) );
  AND U7282 ( .A(n5628), .B(n5629), .Z(n5626) );
  NANDN U7283 ( .B(n5580), .A(n81), .Z(n5629) );
  OR U7284 ( .A(n694), .B(n4992), .Z(n5628) );
  NAND U7285 ( .A(n5630), .B(n5631), .Z(\u_a23_mem/n18191 ) );
  NAND U7286 ( .A(n5611), .B(o[181]), .Z(n5631) );
  AND U7287 ( .A(n5632), .B(n5633), .Z(n5630) );
  NANDN U7288 ( .B(n5580), .A(n86), .Z(n5633) );
  OR U7289 ( .A(n694), .B(n4997), .Z(n5632) );
  NAND U7290 ( .A(n5634), .B(n5635), .Z(\u_a23_mem/n18190 ) );
  NAND U7291 ( .A(n5611), .B(o[182]), .Z(n5635) );
  AND U7292 ( .A(n5636), .B(n5637), .Z(n5634) );
  NANDN U7293 ( .B(n5580), .A(n91), .Z(n5637) );
  OR U7294 ( .A(n694), .B(n5002), .Z(n5636) );
  NAND U7295 ( .A(n5638), .B(n5639), .Z(\u_a23_mem/n18189 ) );
  NAND U7296 ( .A(n5611), .B(o[183]), .Z(n5639) );
  NANDN U7297 ( .B(n5166), .A(n653), .Z(n5611) );
  AND U7298 ( .A(n5640), .B(n5641), .Z(n5638) );
  NANDN U7299 ( .B(n5580), .A(n98), .Z(n5641) );
  NANDN U7300 ( .B(n694), .A(n5009), .Z(n5640) );
  NAND U7301 ( .A(n1165), .B(n653), .Z(n694) );
  NAND U7302 ( .A(n5642), .B(n5643), .Z(\u_a23_mem/n18188 ) );
  NAND U7303 ( .A(n5644), .B(o[184]), .Z(n5643) );
  AND U7304 ( .A(n5645), .B(n5646), .Z(n5642) );
  NANDN U7305 ( .B(n5580), .A(n104), .Z(n5646) );
  OR U7306 ( .A(n728), .B(n4972), .Z(n5645) );
  NAND U7307 ( .A(n5647), .B(n5648), .Z(\u_a23_mem/n18187 ) );
  NAND U7308 ( .A(n5644), .B(o[185]), .Z(n5648) );
  AND U7309 ( .A(n5649), .B(n5650), .Z(n5647) );
  NANDN U7310 ( .B(n5580), .A(n110), .Z(n5650) );
  OR U7311 ( .A(n728), .B(n4977), .Z(n5649) );
  NAND U7312 ( .A(n5651), .B(n5652), .Z(\u_a23_mem/n18186 ) );
  NAND U7313 ( .A(n5644), .B(o[186]), .Z(n5652) );
  AND U7314 ( .A(n5653), .B(n5654), .Z(n5651) );
  NANDN U7315 ( .B(n5580), .A(n115), .Z(n5654) );
  OR U7316 ( .A(n728), .B(n4982), .Z(n5653) );
  NAND U7317 ( .A(n5655), .B(n5656), .Z(\u_a23_mem/n18185 ) );
  NAND U7318 ( .A(n5644), .B(o[187]), .Z(n5656) );
  AND U7319 ( .A(n5657), .B(n5658), .Z(n5655) );
  NANDN U7320 ( .B(n5580), .A(n120), .Z(n5658) );
  OR U7321 ( .A(n728), .B(n4987), .Z(n5657) );
  NAND U7322 ( .A(n5659), .B(n5660), .Z(\u_a23_mem/n18184 ) );
  NAND U7323 ( .A(n5644), .B(o[188]), .Z(n5660) );
  AND U7324 ( .A(n5661), .B(n5662), .Z(n5659) );
  NANDN U7325 ( .B(n5580), .A(n125), .Z(n5662) );
  OR U7326 ( .A(n728), .B(n4992), .Z(n5661) );
  NAND U7327 ( .A(n5663), .B(n5664), .Z(\u_a23_mem/n18183 ) );
  NAND U7328 ( .A(n5644), .B(o[189]), .Z(n5664) );
  AND U7329 ( .A(n5665), .B(n5666), .Z(n5663) );
  NANDN U7330 ( .B(n5580), .A(n130), .Z(n5666) );
  OR U7331 ( .A(n728), .B(n4997), .Z(n5665) );
  NAND U7332 ( .A(n5667), .B(n5668), .Z(\u_a23_mem/n18182 ) );
  NAND U7333 ( .A(n5644), .B(o[190]), .Z(n5668) );
  AND U7334 ( .A(n5669), .B(n5670), .Z(n5667) );
  NANDN U7335 ( .B(n5580), .A(n135), .Z(n5670) );
  OR U7336 ( .A(n728), .B(n5002), .Z(n5669) );
  NAND U7337 ( .A(n5671), .B(n5672), .Z(\u_a23_mem/n18181 ) );
  NAND U7338 ( .A(n5644), .B(o[191]), .Z(n5672) );
  NAND U7339 ( .A(n653), .B(n5077), .Z(n5644) );
  AND U7340 ( .A(n5673), .B(n5674), .Z(n5671) );
  NANDN U7341 ( .B(n5580), .A(n142), .Z(n5674) );
  NAND U7342 ( .A(n5202), .B(n653), .Z(n5580) );
  NANDN U7343 ( .B(n728), .A(n5009), .Z(n5673) );
  NAND U7344 ( .A(n1056), .B(n653), .Z(n728) );
  ANDN U7345 ( .A(n5675), .B(n1939), .Z(n653) );
  AND U7346 ( .A(n5203), .B(n4147), .Z(n5675) );
  IV U7347 ( .A(m_address[3]), .Z(n4147) );
  NAND U7348 ( .A(n5676), .B(n5677), .Z(\u_a23_mem/n18180 ) );
  OR U7349 ( .A(n759), .B(n4972), .Z(n5677) );
  NAND U7350 ( .A(n5678), .B(o[192]), .Z(n5676) );
  NAND U7351 ( .A(n5679), .B(n5680), .Z(\u_a23_mem/n18179 ) );
  OR U7352 ( .A(n759), .B(n4977), .Z(n5680) );
  NAND U7353 ( .A(n5678), .B(o[193]), .Z(n5679) );
  NAND U7354 ( .A(n5681), .B(n5682), .Z(\u_a23_mem/n18178 ) );
  OR U7355 ( .A(n759), .B(n4982), .Z(n5682) );
  NAND U7356 ( .A(n5678), .B(o[194]), .Z(n5681) );
  NAND U7357 ( .A(n5683), .B(n5684), .Z(\u_a23_mem/n18177 ) );
  OR U7358 ( .A(n759), .B(n4987), .Z(n5684) );
  NAND U7359 ( .A(n5678), .B(o[195]), .Z(n5683) );
  NAND U7360 ( .A(n5685), .B(n5686), .Z(\u_a23_mem/n18176 ) );
  OR U7361 ( .A(n759), .B(n4992), .Z(n5686) );
  NAND U7362 ( .A(n5678), .B(o[196]), .Z(n5685) );
  NAND U7363 ( .A(n5687), .B(n5688), .Z(\u_a23_mem/n18175 ) );
  OR U7364 ( .A(n759), .B(n4997), .Z(n5688) );
  NAND U7365 ( .A(n5678), .B(o[197]), .Z(n5687) );
  NAND U7366 ( .A(n5689), .B(n5690), .Z(\u_a23_mem/n18174 ) );
  OR U7367 ( .A(n759), .B(n5002), .Z(n5690) );
  NAND U7368 ( .A(n5678), .B(o[198]), .Z(n5689) );
  NAND U7369 ( .A(n5691), .B(n5692), .Z(\u_a23_mem/n18173 ) );
  NANDN U7370 ( .B(n759), .A(n5009), .Z(n5692) );
  OR U7371 ( .A(n2), .B(n775), .Z(n759) );
  NAND U7372 ( .A(n5678), .B(o[199]), .Z(n5691) );
  OR U7373 ( .A(n5099), .B(n775), .Z(n5678) );
  NAND U7374 ( .A(n5693), .B(n5694), .Z(\u_a23_mem/n18172 ) );
  NAND U7375 ( .A(n5695), .B(o[200]), .Z(n5694) );
  AND U7376 ( .A(n5696), .B(n5697), .Z(n5693) );
  NANDN U7377 ( .B(n5698), .A(n9), .Z(n5697) );
  OR U7378 ( .A(n782), .B(n4972), .Z(n5696) );
  NAND U7379 ( .A(n5699), .B(n5700), .Z(\u_a23_mem/n18171 ) );
  NAND U7380 ( .A(n5695), .B(o[201]), .Z(n5700) );
  AND U7381 ( .A(n5701), .B(n5702), .Z(n5699) );
  NANDN U7382 ( .B(n5698), .A(n16), .Z(n5702) );
  OR U7383 ( .A(n782), .B(n4977), .Z(n5701) );
  NAND U7384 ( .A(n5703), .B(n5704), .Z(\u_a23_mem/n18170 ) );
  NAND U7385 ( .A(n5695), .B(o[202]), .Z(n5704) );
  AND U7386 ( .A(n5705), .B(n5706), .Z(n5703) );
  NANDN U7387 ( .B(n5698), .A(n22), .Z(n5706) );
  OR U7388 ( .A(n782), .B(n4982), .Z(n5705) );
  NAND U7389 ( .A(n5707), .B(n5708), .Z(\u_a23_mem/n18169 ) );
  NAND U7390 ( .A(n5695), .B(o[203]), .Z(n5708) );
  AND U7391 ( .A(n5709), .B(n5710), .Z(n5707) );
  NANDN U7392 ( .B(n5698), .A(n28), .Z(n5710) );
  OR U7393 ( .A(n782), .B(n4987), .Z(n5709) );
  NAND U7394 ( .A(n5711), .B(n5712), .Z(\u_a23_mem/n18168 ) );
  NAND U7395 ( .A(n5695), .B(o[204]), .Z(n5712) );
  AND U7396 ( .A(n5713), .B(n5714), .Z(n5711) );
  NANDN U7397 ( .B(n5698), .A(n34), .Z(n5714) );
  OR U7398 ( .A(n782), .B(n4992), .Z(n5713) );
  NAND U7399 ( .A(n5715), .B(n5716), .Z(\u_a23_mem/n18167 ) );
  NAND U7400 ( .A(n5695), .B(o[205]), .Z(n5716) );
  AND U7401 ( .A(n5717), .B(n5718), .Z(n5715) );
  NANDN U7402 ( .B(n5698), .A(n40), .Z(n5718) );
  OR U7403 ( .A(n782), .B(n4997), .Z(n5717) );
  NAND U7404 ( .A(n5719), .B(n5720), .Z(\u_a23_mem/n18166 ) );
  NAND U7405 ( .A(n5695), .B(o[206]), .Z(n5720) );
  AND U7406 ( .A(n5721), .B(n5722), .Z(n5719) );
  NANDN U7407 ( .B(n5698), .A(n46), .Z(n5722) );
  OR U7408 ( .A(n782), .B(n5002), .Z(n5721) );
  NAND U7409 ( .A(n5723), .B(n5724), .Z(\u_a23_mem/n18165 ) );
  NAND U7410 ( .A(n5695), .B(o[207]), .Z(n5724) );
  OR U7411 ( .A(n5132), .B(n775), .Z(n5695) );
  AND U7412 ( .A(n5725), .B(n5726), .Z(n5723) );
  NANDN U7413 ( .B(n5698), .A(n53), .Z(n5726) );
  NANDN U7414 ( .B(n782), .A(n5009), .Z(n5725) );
  NAND U7415 ( .A(n879), .B(n1121), .Z(n782) );
  NAND U7416 ( .A(n5727), .B(n5728), .Z(\u_a23_mem/n18164 ) );
  NAND U7417 ( .A(n5729), .B(o[208]), .Z(n5728) );
  AND U7418 ( .A(n5730), .B(n5731), .Z(n5727) );
  NANDN U7419 ( .B(n5698), .A(n60), .Z(n5731) );
  OR U7420 ( .A(n816), .B(n4972), .Z(n5730) );
  NAND U7421 ( .A(n5732), .B(n5733), .Z(\u_a23_mem/n18163 ) );
  NAND U7422 ( .A(n5729), .B(o[209]), .Z(n5733) );
  AND U7423 ( .A(n5734), .B(n5735), .Z(n5732) );
  NANDN U7424 ( .B(n5698), .A(n66), .Z(n5735) );
  OR U7425 ( .A(n816), .B(n4977), .Z(n5734) );
  NAND U7426 ( .A(n5736), .B(n5737), .Z(\u_a23_mem/n18162 ) );
  NAND U7427 ( .A(n5729), .B(o[210]), .Z(n5737) );
  AND U7428 ( .A(n5738), .B(n5739), .Z(n5736) );
  NANDN U7429 ( .B(n5698), .A(n71), .Z(n5739) );
  OR U7430 ( .A(n816), .B(n4982), .Z(n5738) );
  NAND U7431 ( .A(n5740), .B(n5741), .Z(\u_a23_mem/n18161 ) );
  NAND U7432 ( .A(n5729), .B(o[211]), .Z(n5741) );
  AND U7433 ( .A(n5742), .B(n5743), .Z(n5740) );
  NANDN U7434 ( .B(n5698), .A(n76), .Z(n5743) );
  OR U7435 ( .A(n816), .B(n4987), .Z(n5742) );
  NAND U7436 ( .A(n5744), .B(n5745), .Z(\u_a23_mem/n18160 ) );
  NAND U7437 ( .A(n5729), .B(o[212]), .Z(n5745) );
  AND U7438 ( .A(n5746), .B(n5747), .Z(n5744) );
  NANDN U7439 ( .B(n5698), .A(n81), .Z(n5747) );
  OR U7440 ( .A(n816), .B(n4992), .Z(n5746) );
  NAND U7441 ( .A(n5748), .B(n5749), .Z(\u_a23_mem/n18159 ) );
  NAND U7442 ( .A(n5729), .B(o[213]), .Z(n5749) );
  AND U7443 ( .A(n5750), .B(n5751), .Z(n5748) );
  NANDN U7444 ( .B(n5698), .A(n86), .Z(n5751) );
  OR U7445 ( .A(n816), .B(n4997), .Z(n5750) );
  NAND U7446 ( .A(n5752), .B(n5753), .Z(\u_a23_mem/n18158 ) );
  NAND U7447 ( .A(n5729), .B(o[214]), .Z(n5753) );
  AND U7448 ( .A(n5754), .B(n5755), .Z(n5752) );
  NANDN U7449 ( .B(n5698), .A(n91), .Z(n5755) );
  OR U7450 ( .A(n816), .B(n5002), .Z(n5754) );
  NAND U7451 ( .A(n5756), .B(n5757), .Z(\u_a23_mem/n18157 ) );
  NAND U7452 ( .A(n5729), .B(o[215]), .Z(n5757) );
  OR U7453 ( .A(n5166), .B(n775), .Z(n5729) );
  AND U7454 ( .A(n5758), .B(n5759), .Z(n5756) );
  NANDN U7455 ( .B(n5698), .A(n98), .Z(n5759) );
  NANDN U7456 ( .B(n816), .A(n5009), .Z(n5758) );
  NAND U7457 ( .A(n879), .B(n1165), .Z(n816) );
  NAND U7458 ( .A(n5760), .B(n5761), .Z(\u_a23_mem/n18156 ) );
  NAND U7459 ( .A(n5762), .B(o[216]), .Z(n5761) );
  AND U7460 ( .A(n5763), .B(n5764), .Z(n5760) );
  NANDN U7461 ( .B(n5698), .A(n104), .Z(n5764) );
  OR U7462 ( .A(n850), .B(n4972), .Z(n5763) );
  NAND U7463 ( .A(n5765), .B(n5766), .Z(\u_a23_mem/n18155 ) );
  NAND U7464 ( .A(n5762), .B(o[217]), .Z(n5766) );
  AND U7465 ( .A(n5767), .B(n5768), .Z(n5765) );
  NANDN U7466 ( .B(n5698), .A(n110), .Z(n5768) );
  OR U7467 ( .A(n850), .B(n4977), .Z(n5767) );
  NAND U7468 ( .A(n5769), .B(n5770), .Z(\u_a23_mem/n18154 ) );
  NAND U7469 ( .A(n5762), .B(o[218]), .Z(n5770) );
  AND U7470 ( .A(n5771), .B(n5772), .Z(n5769) );
  NANDN U7471 ( .B(n5698), .A(n115), .Z(n5772) );
  OR U7472 ( .A(n850), .B(n4982), .Z(n5771) );
  NAND U7473 ( .A(n5773), .B(n5774), .Z(\u_a23_mem/n18153 ) );
  NAND U7474 ( .A(n5762), .B(o[219]), .Z(n5774) );
  AND U7475 ( .A(n5775), .B(n5776), .Z(n5773) );
  NANDN U7476 ( .B(n5698), .A(n120), .Z(n5776) );
  OR U7477 ( .A(n850), .B(n4987), .Z(n5775) );
  NAND U7478 ( .A(n5777), .B(n5778), .Z(\u_a23_mem/n18152 ) );
  NAND U7479 ( .A(n5762), .B(o[220]), .Z(n5778) );
  AND U7480 ( .A(n5779), .B(n5780), .Z(n5777) );
  NANDN U7481 ( .B(n5698), .A(n125), .Z(n5780) );
  OR U7482 ( .A(n850), .B(n4992), .Z(n5779) );
  NAND U7483 ( .A(n5781), .B(n5782), .Z(\u_a23_mem/n18151 ) );
  NAND U7484 ( .A(n5762), .B(o[221]), .Z(n5782) );
  AND U7485 ( .A(n5783), .B(n5784), .Z(n5781) );
  NANDN U7486 ( .B(n5698), .A(n130), .Z(n5784) );
  OR U7487 ( .A(n850), .B(n4997), .Z(n5783) );
  NAND U7488 ( .A(n5785), .B(n5786), .Z(\u_a23_mem/n18150 ) );
  NAND U7489 ( .A(n5762), .B(o[222]), .Z(n5786) );
  AND U7490 ( .A(n5787), .B(n5788), .Z(n5785) );
  NANDN U7491 ( .B(n5698), .A(n135), .Z(n5788) );
  OR U7492 ( .A(n850), .B(n5002), .Z(n5787) );
  NAND U7493 ( .A(n5789), .B(n5790), .Z(\u_a23_mem/n18149 ) );
  NAND U7494 ( .A(n5762), .B(o[223]), .Z(n5790) );
  NANDN U7495 ( .B(n775), .A(n5077), .Z(n5762) );
  IV U7496 ( .A(n879), .Z(n775) );
  AND U7497 ( .A(n5791), .B(n5792), .Z(n5789) );
  NANDN U7498 ( .B(n5698), .A(n142), .Z(n5792) );
  NAND U7499 ( .A(n879), .B(n5202), .Z(n5698) );
  NANDN U7500 ( .B(n850), .A(n5009), .Z(n5791) );
  NAND U7501 ( .A(n879), .B(n1056), .Z(n850) );
  IV U7502 ( .A(n2977), .Z(n1056) );
  NAND U7503 ( .A(n5793), .B(n5794), .Z(\u_a23_mem/n18148 ) );
  OR U7504 ( .A(n882), .B(n4972), .Z(n5794) );
  NAND U7505 ( .A(n5795), .B(o[224]), .Z(n5793) );
  NAND U7506 ( .A(n5796), .B(n5797), .Z(\u_a23_mem/n18147 ) );
  OR U7507 ( .A(n882), .B(n4977), .Z(n5797) );
  NAND U7508 ( .A(n5795), .B(o[225]), .Z(n5796) );
  NAND U7509 ( .A(n5798), .B(n5799), .Z(\u_a23_mem/n18146 ) );
  OR U7510 ( .A(n882), .B(n4982), .Z(n5799) );
  NAND U7511 ( .A(n5795), .B(o[226]), .Z(n5798) );
  NAND U7512 ( .A(n5800), .B(n5801), .Z(\u_a23_mem/n18145 ) );
  OR U7513 ( .A(n882), .B(n4987), .Z(n5801) );
  NAND U7514 ( .A(n5795), .B(o[227]), .Z(n5800) );
  NAND U7515 ( .A(n5802), .B(n5803), .Z(\u_a23_mem/n18144 ) );
  OR U7516 ( .A(n882), .B(n4992), .Z(n5803) );
  NAND U7517 ( .A(n5795), .B(o[228]), .Z(n5802) );
  NAND U7518 ( .A(n5804), .B(n5805), .Z(\u_a23_mem/n18143 ) );
  OR U7519 ( .A(n882), .B(n4997), .Z(n5805) );
  NAND U7520 ( .A(n5795), .B(o[229]), .Z(n5804) );
  NAND U7521 ( .A(n5806), .B(n5807), .Z(\u_a23_mem/n18142 ) );
  OR U7522 ( .A(n882), .B(n5002), .Z(n5807) );
  NAND U7523 ( .A(n5795), .B(o[230]), .Z(n5806) );
  NAND U7524 ( .A(n5808), .B(n5809), .Z(\u_a23_mem/n18141 ) );
  NANDN U7525 ( .B(n882), .A(n5009), .Z(n5809) );
  OR U7526 ( .A(n2), .B(n898), .Z(n882) );
  NAND U7527 ( .A(n5795), .B(o[231]), .Z(n5808) );
  OR U7528 ( .A(n5099), .B(n898), .Z(n5795) );
  NAND U7529 ( .A(n5202), .B(n899), .Z(n5099) );
  AND U7530 ( .A(n5810), .B(n2977), .Z(n899) );
  NAND U7531 ( .A(n5811), .B(n5812), .Z(\u_a23_mem/n18140 ) );
  NAND U7532 ( .A(n5813), .B(o[232]), .Z(n5812) );
  AND U7533 ( .A(n5814), .B(n5815), .Z(n5811) );
  NAND U7534 ( .A(n5816), .B(n9), .Z(n5815) );
  AND U7535 ( .A(n5817), .B(m_write[8]), .Z(n9) );
  OR U7536 ( .A(n906), .B(n4972), .Z(n5814) );
  NAND U7537 ( .A(n5818), .B(n5819), .Z(\u_a23_mem/n18139 ) );
  NAND U7538 ( .A(n5813), .B(o[233]), .Z(n5819) );
  AND U7539 ( .A(n5820), .B(n5821), .Z(n5818) );
  NAND U7540 ( .A(n5816), .B(n16), .Z(n5821) );
  AND U7541 ( .A(n5817), .B(m_write[9]), .Z(n16) );
  OR U7542 ( .A(n906), .B(n4977), .Z(n5820) );
  NAND U7543 ( .A(n5822), .B(n5823), .Z(\u_a23_mem/n18138 ) );
  NAND U7544 ( .A(n5813), .B(o[234]), .Z(n5823) );
  AND U7545 ( .A(n5824), .B(n5825), .Z(n5822) );
  NAND U7546 ( .A(n5816), .B(n22), .Z(n5825) );
  AND U7547 ( .A(n5817), .B(m_write[10]), .Z(n22) );
  OR U7548 ( .A(n906), .B(n4982), .Z(n5824) );
  NAND U7549 ( .A(n5826), .B(n5827), .Z(\u_a23_mem/n18137 ) );
  NAND U7550 ( .A(n5813), .B(o[235]), .Z(n5827) );
  AND U7551 ( .A(n5828), .B(n5829), .Z(n5826) );
  NAND U7552 ( .A(n5816), .B(n28), .Z(n5829) );
  AND U7553 ( .A(n5817), .B(m_write[11]), .Z(n28) );
  OR U7554 ( .A(n906), .B(n4987), .Z(n5828) );
  NAND U7555 ( .A(n5830), .B(n5831), .Z(\u_a23_mem/n18136 ) );
  NAND U7556 ( .A(n5813), .B(o[236]), .Z(n5831) );
  AND U7557 ( .A(n5832), .B(n5833), .Z(n5830) );
  NAND U7558 ( .A(n5816), .B(n34), .Z(n5833) );
  AND U7559 ( .A(n5817), .B(m_write[12]), .Z(n34) );
  OR U7560 ( .A(n906), .B(n4992), .Z(n5832) );
  NAND U7561 ( .A(n5834), .B(n5835), .Z(\u_a23_mem/n18135 ) );
  NAND U7562 ( .A(n5813), .B(o[237]), .Z(n5835) );
  AND U7563 ( .A(n5836), .B(n5837), .Z(n5834) );
  NAND U7564 ( .A(n5816), .B(n40), .Z(n5837) );
  AND U7565 ( .A(n5817), .B(m_write[13]), .Z(n40) );
  OR U7566 ( .A(n906), .B(n4997), .Z(n5836) );
  NAND U7567 ( .A(n5838), .B(n5839), .Z(\u_a23_mem/n18134 ) );
  NAND U7568 ( .A(n5813), .B(o[238]), .Z(n5839) );
  AND U7569 ( .A(n5840), .B(n5841), .Z(n5838) );
  NAND U7570 ( .A(n5816), .B(n46), .Z(n5841) );
  AND U7571 ( .A(n5817), .B(m_write[14]), .Z(n46) );
  OR U7572 ( .A(n906), .B(n5002), .Z(n5840) );
  NAND U7573 ( .A(n5842), .B(n5843), .Z(\u_a23_mem/n18133 ) );
  NAND U7574 ( .A(n5813), .B(o[239]), .Z(n5843) );
  OR U7575 ( .A(n5132), .B(n898), .Z(n5813) );
  NAND U7576 ( .A(n5202), .B(n933), .Z(n5132) );
  ANDN U7577 ( .A(n5844), .B(n1165), .Z(n933) );
  AND U7578 ( .A(n5845), .B(n5846), .Z(n5842) );
  NAND U7579 ( .A(n5816), .B(n53), .Z(n5846) );
  AND U7580 ( .A(n5817), .B(m_write[15]), .Z(n53) );
  NANDN U7581 ( .B(n906), .A(n5009), .Z(n5845) );
  NAND U7582 ( .A(n1006), .B(n1121), .Z(n906) );
  IV U7583 ( .A(n2937), .Z(n1121) );
  NAND U7584 ( .A(n5847), .B(n5848), .Z(\u_a23_mem/n18132 ) );
  NAND U7585 ( .A(n5849), .B(o[240]), .Z(n5848) );
  AND U7586 ( .A(n5850), .B(n5851), .Z(n5847) );
  NAND U7587 ( .A(n5816), .B(n60), .Z(n5851) );
  AND U7588 ( .A(n5817), .B(m_write[16]), .Z(n60) );
  OR U7589 ( .A(n941), .B(n4972), .Z(n5850) );
  NAND U7590 ( .A(n5852), .B(n5853), .Z(\u_a23_mem/n18131 ) );
  NAND U7591 ( .A(n5849), .B(o[241]), .Z(n5853) );
  AND U7592 ( .A(n5854), .B(n5855), .Z(n5852) );
  NAND U7593 ( .A(n5816), .B(n66), .Z(n5855) );
  AND U7594 ( .A(n5817), .B(m_write[17]), .Z(n66) );
  OR U7595 ( .A(n941), .B(n4977), .Z(n5854) );
  NAND U7596 ( .A(n5856), .B(n5857), .Z(\u_a23_mem/n18130 ) );
  NAND U7597 ( .A(n5849), .B(o[242]), .Z(n5857) );
  AND U7598 ( .A(n5858), .B(n5859), .Z(n5856) );
  NAND U7599 ( .A(n5816), .B(n71), .Z(n5859) );
  AND U7600 ( .A(n5817), .B(m_write[18]), .Z(n71) );
  OR U7601 ( .A(n941), .B(n4982), .Z(n5858) );
  NAND U7602 ( .A(n5860), .B(n5861), .Z(\u_a23_mem/n18129 ) );
  NAND U7603 ( .A(n5849), .B(o[243]), .Z(n5861) );
  AND U7604 ( .A(n5862), .B(n5863), .Z(n5860) );
  NAND U7605 ( .A(n5816), .B(n76), .Z(n5863) );
  AND U7606 ( .A(n5817), .B(m_write[19]), .Z(n76) );
  OR U7607 ( .A(n941), .B(n4987), .Z(n5862) );
  NAND U7608 ( .A(n5864), .B(n5865), .Z(\u_a23_mem/n18128 ) );
  NAND U7609 ( .A(n5849), .B(o[244]), .Z(n5865) );
  AND U7610 ( .A(n5866), .B(n5867), .Z(n5864) );
  NAND U7611 ( .A(n5816), .B(n81), .Z(n5867) );
  AND U7612 ( .A(n5817), .B(m_write[20]), .Z(n81) );
  OR U7613 ( .A(n941), .B(n4992), .Z(n5866) );
  NAND U7614 ( .A(n5868), .B(n5869), .Z(\u_a23_mem/n18127 ) );
  NAND U7615 ( .A(n5849), .B(o[245]), .Z(n5869) );
  AND U7616 ( .A(n5870), .B(n5871), .Z(n5868) );
  NAND U7617 ( .A(n5816), .B(n86), .Z(n5871) );
  AND U7618 ( .A(n5817), .B(m_write[21]), .Z(n86) );
  OR U7619 ( .A(n941), .B(n4997), .Z(n5870) );
  NAND U7620 ( .A(n5872), .B(n5873), .Z(\u_a23_mem/n18126 ) );
  NAND U7621 ( .A(n5849), .B(o[246]), .Z(n5873) );
  AND U7622 ( .A(n5874), .B(n5875), .Z(n5872) );
  NAND U7623 ( .A(n5816), .B(n91), .Z(n5875) );
  AND U7624 ( .A(n5817), .B(m_write[22]), .Z(n91) );
  OR U7625 ( .A(n941), .B(n5002), .Z(n5874) );
  NAND U7626 ( .A(n5876), .B(n5877), .Z(\u_a23_mem/n18125 ) );
  NAND U7627 ( .A(n5849), .B(o[247]), .Z(n5877) );
  OR U7628 ( .A(n5166), .B(n898), .Z(n5849) );
  NAND U7629 ( .A(n5202), .B(n968), .Z(n5166) );
  AND U7630 ( .A(n5844), .B(n2937), .Z(n968) );
  ANDN U7631 ( .A(n5878), .B(n2979), .Z(n5844) );
  AND U7632 ( .A(n2977), .B(n2980), .Z(n5878) );
  AND U7633 ( .A(n5879), .B(n5880), .Z(n5876) );
  NAND U7634 ( .A(n5816), .B(n98), .Z(n5880) );
  AND U7635 ( .A(n5817), .B(m_write[23]), .Z(n98) );
  NANDN U7636 ( .B(n941), .A(n5009), .Z(n5879) );
  NAND U7637 ( .A(n1006), .B(n1165), .Z(n941) );
  IV U7638 ( .A(n2978), .Z(n1165) );
  NAND U7639 ( .A(n5881), .B(n5882), .Z(\u_a23_mem/n18124 ) );
  NAND U7640 ( .A(n5883), .B(o[248]), .Z(n5882) );
  AND U7641 ( .A(n5884), .B(n5885), .Z(n5881) );
  NAND U7642 ( .A(n5816), .B(n104), .Z(n5885) );
  AND U7643 ( .A(n5817), .B(m_write[24]), .Z(n104) );
  NANDN U7644 ( .B(n4972), .A(n976), .Z(n5884) );
  NAND U7645 ( .A(n5202), .B(m_write[0]), .Z(n4972) );
  NAND U7646 ( .A(n5886), .B(n5887), .Z(\u_a23_mem/n18123 ) );
  NAND U7647 ( .A(n5883), .B(o[249]), .Z(n5887) );
  AND U7648 ( .A(n5888), .B(n5889), .Z(n5886) );
  NAND U7649 ( .A(n5816), .B(n110), .Z(n5889) );
  AND U7650 ( .A(n5817), .B(m_write[25]), .Z(n110) );
  NANDN U7651 ( .B(n4977), .A(n976), .Z(n5888) );
  NAND U7652 ( .A(n5202), .B(m_write[1]), .Z(n4977) );
  NAND U7653 ( .A(n5890), .B(n5891), .Z(\u_a23_mem/n18122 ) );
  NAND U7654 ( .A(n5883), .B(o[250]), .Z(n5891) );
  AND U7655 ( .A(n5892), .B(n5893), .Z(n5890) );
  NAND U7656 ( .A(n5816), .B(n115), .Z(n5893) );
  AND U7657 ( .A(n5817), .B(m_write[26]), .Z(n115) );
  NANDN U7658 ( .B(n4982), .A(n976), .Z(n5892) );
  NAND U7659 ( .A(n5202), .B(m_write[2]), .Z(n4982) );
  NAND U7660 ( .A(n5894), .B(n5895), .Z(\u_a23_mem/n18121 ) );
  NAND U7661 ( .A(n5883), .B(o[251]), .Z(n5895) );
  AND U7662 ( .A(n5896), .B(n5897), .Z(n5894) );
  NAND U7663 ( .A(n5816), .B(n120), .Z(n5897) );
  AND U7664 ( .A(n5817), .B(m_write[27]), .Z(n120) );
  NANDN U7665 ( .B(n4987), .A(n976), .Z(n5896) );
  NAND U7666 ( .A(n5202), .B(m_write[3]), .Z(n4987) );
  NAND U7667 ( .A(n5898), .B(n5899), .Z(\u_a23_mem/n18120 ) );
  NAND U7668 ( .A(n5883), .B(o[252]), .Z(n5899) );
  AND U7669 ( .A(n5900), .B(n5901), .Z(n5898) );
  NAND U7670 ( .A(n5816), .B(n125), .Z(n5901) );
  AND U7671 ( .A(n5817), .B(m_write[28]), .Z(n125) );
  NANDN U7672 ( .B(n4992), .A(n976), .Z(n5900) );
  NAND U7673 ( .A(n5202), .B(m_write[4]), .Z(n4992) );
  NAND U7674 ( .A(n5902), .B(n5903), .Z(\u_a23_mem/n18119 ) );
  NAND U7675 ( .A(n5883), .B(o[253]), .Z(n5903) );
  AND U7676 ( .A(n5904), .B(n5905), .Z(n5902) );
  NAND U7677 ( .A(n5816), .B(n130), .Z(n5905) );
  AND U7678 ( .A(n5817), .B(m_write[29]), .Z(n130) );
  NANDN U7679 ( .B(n4997), .A(n976), .Z(n5904) );
  NAND U7680 ( .A(n5202), .B(m_write[5]), .Z(n4997) );
  NAND U7681 ( .A(n5906), .B(n5907), .Z(\u_a23_mem/n18118 ) );
  NAND U7682 ( .A(n5883), .B(o[254]), .Z(n5907) );
  AND U7683 ( .A(n5908), .B(n5909), .Z(n5906) );
  NAND U7684 ( .A(n5816), .B(n135), .Z(n5909) );
  AND U7685 ( .A(n5817), .B(m_write[30]), .Z(n135) );
  NANDN U7686 ( .B(n5002), .A(n976), .Z(n5908) );
  NAND U7687 ( .A(n5202), .B(m_write[6]), .Z(n5002) );
  NAND U7688 ( .A(n5910), .B(n5911), .Z(\u_a23_mem/n18117 ) );
  NAND U7689 ( .A(n5883), .B(o[255]), .Z(n5911) );
  NANDN U7690 ( .B(n898), .A(n5077), .Z(n5883) );
  AND U7691 ( .A(n1003), .B(n5202), .Z(n5077) );
  ANDN U7692 ( .A(n5810), .B(n5006), .Z(n1003) );
  ANDN U7693 ( .A(n5912), .B(n2979), .Z(n5810) );
  ANDN U7694 ( .A(n2977), .B(n5043), .Z(n2979) );
  NAND U7695 ( .A(n2937), .B(n5913), .Z(n5043) );
  AND U7696 ( .A(n2), .B(n2978), .Z(n5913) );
  NOR U7697 ( .A(n5006), .B(n5817), .Z(n2) );
  IV U7698 ( .A(n2980), .Z(n5006) );
  NAND U7699 ( .A(n5914), .B(n5915), .Z(n2980) );
  AND U7700 ( .A(m_byte_enable[0]), .B(n5916), .Z(n5914) );
  AND U7701 ( .A(n2978), .B(n2937), .Z(n5912) );
  NAND U7702 ( .A(n5917), .B(n5915), .Z(n2937) );
  AND U7703 ( .A(n5918), .B(n5919), .Z(n5915) );
  ANDN U7704 ( .A(m_byte_enable[1]), .B(m_byte_enable[0]), .Z(n5917) );
  NAND U7705 ( .A(n5920), .B(n5921), .Z(n2978) );
  AND U7706 ( .A(n5916), .B(n5919), .Z(n5921) );
  IV U7707 ( .A(m_byte_enable[3]), .Z(n5919) );
  ANDN U7708 ( .A(m_byte_enable[2]), .B(m_byte_enable[0]), .Z(n5920) );
  AND U7709 ( .A(n5922), .B(n5923), .Z(n5910) );
  NAND U7710 ( .A(n142), .B(n5816), .Z(n5923) );
  ANDN U7711 ( .A(n5202), .B(n898), .Z(n5816) );
  IV U7712 ( .A(n1006), .Z(n898) );
  AND U7713 ( .A(n5817), .B(m_write[31]), .Z(n142) );
  AND U7714 ( .A(n5924), .B(n5925), .Z(n5817) );
  AND U7715 ( .A(m_byte_enable[0]), .B(m_byte_enable[1]), .Z(n5925) );
  AND U7716 ( .A(m_byte_enable[2]), .B(m_byte_enable[3]), .Z(n5924) );
  NAND U7717 ( .A(n5009), .B(n976), .Z(n5922) );
  ANDN U7718 ( .A(n1006), .B(n2977), .Z(n976) );
  NAND U7719 ( .A(n5926), .B(n5927), .Z(n2977) );
  AND U7720 ( .A(n5916), .B(n5918), .Z(n5927) );
  IV U7721 ( .A(m_byte_enable[2]), .Z(n5918) );
  IV U7722 ( .A(m_byte_enable[1]), .Z(n5916) );
  ANDN U7723 ( .A(m_byte_enable[3]), .B(m_byte_enable[0]), .Z(n5926) );
  ANDN U7724 ( .A(n5928), .B(n1939), .Z(n1006) );
  AND U7725 ( .A(n5203), .B(m_address[3]), .Z(n5928) );
  AND U7726 ( .A(n4963), .B(m_address[2]), .Z(n5203) );
  ANDN U7727 ( .A(m_write[7]), .B(n5041), .Z(n5009) );
  IV U7728 ( .A(n5202), .Z(n5041) );
  AND U7729 ( .A(m_write_en), .B(n5929), .Z(n5202) );
  AND U7730 ( .A(\u_a23_core/write_data_wen ), .B(n5930), .Z(
        \u_a23_core/u_execute/write_enable_nxt ) );
  NAND U7731 ( .A(n5931), .B(n5932), .Z(
        \u_a23_core/u_execute/write_data_nxt[9] ) );
  NAND U7732 ( .A(n5933), .B(n5934), .Z(n5932) );
  AND U7733 ( .A(n5935), .B(n5936), .Z(n5931) );
  NAND U7734 ( .A(n5937), .B(n5938), .Z(n5936) );
  NAND U7735 ( .A(n5939), .B(n5940), .Z(
        \u_a23_core/u_execute/write_data_nxt[8] ) );
  NAND U7736 ( .A(n5933), .B(n5941), .Z(n5940) );
  AND U7737 ( .A(n5942), .B(n5943), .Z(n5939) );
  NAND U7738 ( .A(n5944), .B(n5938), .Z(n5943) );
  NAND U7739 ( .A(n5945), .B(n5946), .Z(
        \u_a23_core/u_execute/write_data_nxt[31] ) );
  NAND U7740 ( .A(n5933), .B(\u_a23_core/u_execute/rs[31] ), .Z(n5946) );
  AND U7741 ( .A(n5947), .B(n5948), .Z(n5945) );
  NAND U7742 ( .A(\u_a23_core/u_execute/save_int_pc_m4[31] ), .B(n5938), .Z(
        n5948) );
  NAND U7743 ( .A(n5949), .B(n5950), .Z(
        \u_a23_core/u_execute/write_data_nxt[30] ) );
  NAND U7744 ( .A(n5933), .B(\u_a23_core/u_execute/rs[30] ), .Z(n5950) );
  AND U7745 ( .A(n5951), .B(n5952), .Z(n5949) );
  NAND U7746 ( .A(\u_a23_core/u_execute/save_int_pc_m4[30] ), .B(n5938), .Z(
        n5952) );
  NAND U7747 ( .A(n5953), .B(n5954), .Z(
        \u_a23_core/u_execute/write_data_nxt[29] ) );
  NAND U7748 ( .A(n5933), .B(\u_a23_core/u_execute/rs[29] ), .Z(n5954) );
  AND U7749 ( .A(n5955), .B(n5956), .Z(n5953) );
  NAND U7750 ( .A(\u_a23_core/u_execute/save_int_pc_m4[29] ), .B(n5938), .Z(
        n5956) );
  NAND U7751 ( .A(n5957), .B(n5958), .Z(
        \u_a23_core/u_execute/write_data_nxt[28] ) );
  NAND U7752 ( .A(n5933), .B(\u_a23_core/u_execute/rs[28] ), .Z(n5958) );
  AND U7753 ( .A(n5959), .B(n5960), .Z(n5957) );
  NAND U7754 ( .A(\u_a23_core/u_execute/save_int_pc_m4[28] ), .B(n5938), .Z(
        n5960) );
  NAND U7755 ( .A(n5961), .B(n5962), .Z(
        \u_a23_core/u_execute/write_data_nxt[27] ) );
  NAND U7756 ( .A(n5933), .B(\u_a23_core/u_execute/rs[27] ), .Z(n5962) );
  ANDN U7757 ( .A(n5963), .B(n5938), .Z(n5961) );
  NAND U7758 ( .A(n5964), .B(n5965), .Z(
        \u_a23_core/u_execute/write_data_nxt[26] ) );
  NAND U7759 ( .A(n5933), .B(\u_a23_core/u_execute/rs[26] ), .Z(n5965) );
  ANDN U7760 ( .A(n5966), .B(n5938), .Z(n5964) );
  NAND U7761 ( .A(n5967), .B(n5968), .Z(
        \u_a23_core/u_execute/write_data_nxt[25] ) );
  NAND U7762 ( .A(n5933), .B(n5969), .Z(n5968) );
  AND U7763 ( .A(n5935), .B(n5970), .Z(n5967) );
  NAND U7764 ( .A(n5971), .B(n5938), .Z(n5970) );
  NAND U7765 ( .A(n5972), .B(n5973), .Z(
        \u_a23_core/u_execute/write_data_nxt[24] ) );
  NAND U7766 ( .A(n5933), .B(n5974), .Z(n5973) );
  AND U7767 ( .A(n5942), .B(n5975), .Z(n5972) );
  NAND U7768 ( .A(n5976), .B(n5938), .Z(n5975) );
  NAND U7769 ( .A(n5977), .B(n5978), .Z(
        \u_a23_core/u_execute/write_data_nxt[23] ) );
  NAND U7770 ( .A(n5933), .B(n5979), .Z(n5978) );
  AND U7771 ( .A(n5947), .B(n5980), .Z(n5977) );
  NAND U7772 ( .A(n5981), .B(n5938), .Z(n5980) );
  NAND U7773 ( .A(n5982), .B(n5983), .Z(
        \u_a23_core/u_execute/write_data_nxt[22] ) );
  NAND U7774 ( .A(n5933), .B(n5984), .Z(n5983) );
  AND U7775 ( .A(n5951), .B(n5985), .Z(n5982) );
  NAND U7776 ( .A(n5986), .B(n5938), .Z(n5985) );
  NAND U7777 ( .A(n5987), .B(n5988), .Z(
        \u_a23_core/u_execute/write_data_nxt[21] ) );
  NAND U7778 ( .A(n5933), .B(n5989), .Z(n5988) );
  AND U7779 ( .A(n5955), .B(n5990), .Z(n5987) );
  NAND U7780 ( .A(n5991), .B(n5938), .Z(n5990) );
  NAND U7781 ( .A(n5992), .B(n5993), .Z(
        \u_a23_core/u_execute/write_data_nxt[20] ) );
  NAND U7782 ( .A(n5933), .B(n5994), .Z(n5993) );
  AND U7783 ( .A(n5959), .B(n5995), .Z(n5992) );
  NAND U7784 ( .A(n5996), .B(n5938), .Z(n5995) );
  NAND U7785 ( .A(n5997), .B(n5998), .Z(
        \u_a23_core/u_execute/write_data_nxt[19] ) );
  NAND U7786 ( .A(n5933), .B(n5999), .Z(n5998) );
  AND U7787 ( .A(n5963), .B(n6000), .Z(n5997) );
  NAND U7788 ( .A(n6001), .B(n5938), .Z(n6000) );
  NAND U7789 ( .A(n6002), .B(n6003), .Z(
        \u_a23_core/u_execute/write_data_nxt[18] ) );
  NAND U7790 ( .A(n5933), .B(n6004), .Z(n6003) );
  AND U7791 ( .A(n5966), .B(n6005), .Z(n6002) );
  NAND U7792 ( .A(n6006), .B(n5938), .Z(n6005) );
  NAND U7793 ( .A(n6007), .B(n6008), .Z(
        \u_a23_core/u_execute/write_data_nxt[17] ) );
  NAND U7794 ( .A(n5933), .B(n6009), .Z(n6008) );
  AND U7795 ( .A(n5935), .B(n6010), .Z(n6007) );
  NAND U7796 ( .A(n6011), .B(n5938), .Z(n6010) );
  NANDN U7797 ( .B(n5933), .A(\u_a23_core/u_execute/rs[1] ), .Z(n5935) );
  NAND U7798 ( .A(n6012), .B(n6013), .Z(
        \u_a23_core/u_execute/write_data_nxt[16] ) );
  NAND U7799 ( .A(n5933), .B(n6014), .Z(n6013) );
  AND U7800 ( .A(n5942), .B(n6015), .Z(n6012) );
  NAND U7801 ( .A(n6016), .B(n5938), .Z(n6015) );
  NANDN U7802 ( .B(n5933), .A(\u_a23_core/u_execute/rs[0] ), .Z(n5942) );
  NAND U7803 ( .A(n6017), .B(n6018), .Z(
        \u_a23_core/u_execute/write_data_nxt[15] ) );
  NAND U7804 ( .A(n5933), .B(n6019), .Z(n6018) );
  AND U7805 ( .A(n5947), .B(n6020), .Z(n6017) );
  NAND U7806 ( .A(n6021), .B(n5938), .Z(n6020) );
  NANDN U7807 ( .B(n5933), .A(\u_a23_core/u_execute/write_data_nxt[7] ), .Z(
        n5947) );
  NAND U7808 ( .A(n6022), .B(n6023), .Z(
        \u_a23_core/u_execute/write_data_nxt[7] ) );
  NAND U7809 ( .A(n6024), .B(n6025), .Z(n6022) );
  NAND U7810 ( .A(n6026), .B(n6027), .Z(
        \u_a23_core/u_execute/write_data_nxt[14] ) );
  NAND U7811 ( .A(n5933), .B(n6028), .Z(n6027) );
  AND U7812 ( .A(n5951), .B(n6029), .Z(n6026) );
  NAND U7813 ( .A(n6030), .B(n5938), .Z(n6029) );
  NANDN U7814 ( .B(n5933), .A(\u_a23_core/u_execute/write_data_nxt[6] ), .Z(
        n5951) );
  NAND U7815 ( .A(n6031), .B(n6032), .Z(
        \u_a23_core/u_execute/write_data_nxt[6] ) );
  NAND U7816 ( .A(n6033), .B(n6025), .Z(n6031) );
  NAND U7817 ( .A(n6034), .B(n6035), .Z(
        \u_a23_core/u_execute/write_data_nxt[13] ) );
  NAND U7818 ( .A(n5933), .B(n6036), .Z(n6035) );
  AND U7819 ( .A(n5955), .B(n6037), .Z(n6034) );
  NAND U7820 ( .A(n6038), .B(n5938), .Z(n6037) );
  NANDN U7821 ( .B(n5933), .A(\u_a23_core/u_execute/write_data_nxt[5] ), .Z(
        n5955) );
  NAND U7822 ( .A(n6039), .B(n6040), .Z(
        \u_a23_core/u_execute/write_data_nxt[5] ) );
  NAND U7823 ( .A(n6041), .B(n6025), .Z(n6039) );
  NAND U7824 ( .A(n6042), .B(n6043), .Z(
        \u_a23_core/u_execute/write_data_nxt[12] ) );
  NAND U7825 ( .A(n5933), .B(n6044), .Z(n6043) );
  AND U7826 ( .A(n5959), .B(n6045), .Z(n6042) );
  NAND U7827 ( .A(n6046), .B(n5938), .Z(n6045) );
  NANDN U7828 ( .B(n5933), .A(\u_a23_core/u_execute/write_data_nxt[4] ), .Z(
        n5959) );
  NAND U7829 ( .A(n6047), .B(n6048), .Z(
        \u_a23_core/u_execute/write_data_nxt[4] ) );
  NAND U7830 ( .A(n6049), .B(n6025), .Z(n6047) );
  NAND U7831 ( .A(n6050), .B(n6051), .Z(
        \u_a23_core/u_execute/write_data_nxt[11] ) );
  NAND U7832 ( .A(n5933), .B(n6052), .Z(n6051) );
  AND U7833 ( .A(n5963), .B(n6053), .Z(n6050) );
  NAND U7834 ( .A(n6054), .B(n5938), .Z(n6053) );
  NANDN U7835 ( .B(n5933), .A(\u_a23_core/u_execute/write_data_nxt[3] ), .Z(
        n5963) );
  NAND U7836 ( .A(n6055), .B(n6056), .Z(
        \u_a23_core/u_execute/write_data_nxt[3] ) );
  NAND U7837 ( .A(n6057), .B(n6025), .Z(n6055) );
  NAND U7838 ( .A(n6058), .B(n6059), .Z(
        \u_a23_core/u_execute/write_data_nxt[10] ) );
  NAND U7839 ( .A(n5933), .B(n6060), .Z(n6059) );
  AND U7840 ( .A(n5966), .B(n6061), .Z(n6058) );
  NAND U7841 ( .A(n6062), .B(n5938), .Z(n6061) );
  ANDN U7842 ( .A(n6025), .B(\u_a23_core/byte_enable_sel[0] ), .Z(n5938) );
  NANDN U7843 ( .B(n5933), .A(\u_a23_core/u_execute/write_data_nxt[2] ), .Z(
        n5966) );
  NAND U7844 ( .A(n6063), .B(n6064), .Z(
        \u_a23_core/u_execute/write_data_nxt[2] ) );
  NAND U7845 ( .A(n6065), .B(n6025), .Z(n6063) );
  IV U7846 ( .A(\u_a23_core/byte_enable_sel[0] ), .Z(n5933) );
  MUX U7847 ( .IN0(\u_a23_core/u_execute/u_register_bank/r11[31] ), .IN1(n6066), .SEL(n6067), .F(\u_a23_core/u_execute/u_register_bank/n4981 ) );
  MUX U7848 ( .IN0(\u_a23_core/u_execute/u_register_bank/r11[30] ), .IN1(n6068), .SEL(n6067), .F(\u_a23_core/u_execute/u_register_bank/n4979 ) );
  MUX U7849 ( .IN0(\u_a23_core/u_execute/u_register_bank/r11[29] ), .IN1(n6069), .SEL(n6067), .F(\u_a23_core/u_execute/u_register_bank/n4977 ) );
  MUX U7850 ( .IN0(\u_a23_core/u_execute/u_register_bank/r11[28] ), .IN1(n6070), .SEL(n6067), .F(\u_a23_core/u_execute/u_register_bank/n4975 ) );
  MUX U7851 ( .IN0(\u_a23_core/u_execute/u_register_bank/r11[27] ), .IN1(n6071), .SEL(n6067), .F(\u_a23_core/u_execute/u_register_bank/n4973 ) );
  MUX U7852 ( .IN0(\u_a23_core/u_execute/u_register_bank/r11[26] ), .IN1(n6072), .SEL(n6067), .F(\u_a23_core/u_execute/u_register_bank/n4971 ) );
  MUX U7853 ( .IN0(\u_a23_core/u_execute/u_register_bank/r11[25] ), .IN1(n6073), .SEL(n6067), .F(\u_a23_core/u_execute/u_register_bank/n4969 ) );
  MUX U7854 ( .IN0(\u_a23_core/u_execute/u_register_bank/r11[24] ), .IN1(n6074), .SEL(n6067), .F(\u_a23_core/u_execute/u_register_bank/n4967 ) );
  MUX U7855 ( .IN0(\u_a23_core/u_execute/u_register_bank/r11[23] ), .IN1(n6075), .SEL(n6067), .F(\u_a23_core/u_execute/u_register_bank/n4965 ) );
  MUX U7856 ( .IN0(\u_a23_core/u_execute/u_register_bank/r11[22] ), .IN1(n6076), .SEL(n6067), .F(\u_a23_core/u_execute/u_register_bank/n4963 ) );
  MUX U7857 ( .IN0(\u_a23_core/u_execute/u_register_bank/r11[21] ), .IN1(n6077), .SEL(n6067), .F(\u_a23_core/u_execute/u_register_bank/n4961 ) );
  MUX U7858 ( .IN0(\u_a23_core/u_execute/u_register_bank/r11[20] ), .IN1(n6078), .SEL(n6067), .F(\u_a23_core/u_execute/u_register_bank/n4959 ) );
  MUX U7859 ( .IN0(\u_a23_core/u_execute/u_register_bank/r11[19] ), .IN1(n6079), .SEL(n6067), .F(\u_a23_core/u_execute/u_register_bank/n4957 ) );
  MUX U7860 ( .IN0(\u_a23_core/u_execute/u_register_bank/r11[18] ), .IN1(n6080), .SEL(n6067), .F(\u_a23_core/u_execute/u_register_bank/n4955 ) );
  MUX U7861 ( .IN0(\u_a23_core/u_execute/u_register_bank/r11[17] ), .IN1(n6081), .SEL(n6067), .F(\u_a23_core/u_execute/u_register_bank/n4953 ) );
  MUX U7862 ( .IN0(\u_a23_core/u_execute/u_register_bank/r11[16] ), .IN1(n6082), .SEL(n6067), .F(\u_a23_core/u_execute/u_register_bank/n4951 ) );
  MUX U7863 ( .IN0(\u_a23_core/u_execute/u_register_bank/r11[15] ), .IN1(n6083), .SEL(n6067), .F(\u_a23_core/u_execute/u_register_bank/n4949 ) );
  MUX U7864 ( .IN0(\u_a23_core/u_execute/u_register_bank/r11[14] ), .IN1(n6084), .SEL(n6067), .F(\u_a23_core/u_execute/u_register_bank/n4947 ) );
  MUX U7865 ( .IN0(\u_a23_core/u_execute/u_register_bank/r11[13] ), .IN1(n6085), .SEL(n6067), .F(\u_a23_core/u_execute/u_register_bank/n4945 ) );
  MUX U7866 ( .IN0(\u_a23_core/u_execute/u_register_bank/r11[12] ), .IN1(n6086), .SEL(n6067), .F(\u_a23_core/u_execute/u_register_bank/n4943 ) );
  MUX U7867 ( .IN0(\u_a23_core/u_execute/u_register_bank/r11[11] ), .IN1(n6087), .SEL(n6067), .F(\u_a23_core/u_execute/u_register_bank/n4941 ) );
  MUX U7868 ( .IN0(\u_a23_core/u_execute/u_register_bank/r11[10] ), .IN1(n6088), .SEL(n6067), .F(\u_a23_core/u_execute/u_register_bank/n4939 ) );
  MUX U7869 ( .IN0(\u_a23_core/u_execute/u_register_bank/r11[9] ), .IN1(n6089), 
        .SEL(n6067), .F(\u_a23_core/u_execute/u_register_bank/n4937 ) );
  MUX U7870 ( .IN0(\u_a23_core/u_execute/u_register_bank/r11[8] ), .IN1(n6090), 
        .SEL(n6067), .F(\u_a23_core/u_execute/u_register_bank/n4935 ) );
  MUX U7871 ( .IN0(\u_a23_core/u_execute/u_register_bank/r11[7] ), .IN1(n6091), 
        .SEL(n6067), .F(\u_a23_core/u_execute/u_register_bank/n4933 ) );
  MUX U7872 ( .IN0(\u_a23_core/u_execute/u_register_bank/r11[6] ), .IN1(n6092), 
        .SEL(n6067), .F(\u_a23_core/u_execute/u_register_bank/n4931 ) );
  MUX U7873 ( .IN0(\u_a23_core/u_execute/u_register_bank/r11[5] ), .IN1(n6093), 
        .SEL(n6067), .F(\u_a23_core/u_execute/u_register_bank/n4929 ) );
  MUX U7874 ( .IN0(\u_a23_core/u_execute/u_register_bank/r11[4] ), .IN1(n6094), 
        .SEL(n6067), .F(\u_a23_core/u_execute/u_register_bank/n4927 ) );
  MUX U7875 ( .IN0(\u_a23_core/u_execute/u_register_bank/r11[3] ), .IN1(n6095), 
        .SEL(n6067), .F(\u_a23_core/u_execute/u_register_bank/n4925 ) );
  MUX U7876 ( .IN0(\u_a23_core/u_execute/u_register_bank/r11[2] ), .IN1(n6096), 
        .SEL(n6067), .F(\u_a23_core/u_execute/u_register_bank/n4923 ) );
  MUX U7877 ( .IN0(\u_a23_core/u_execute/u_register_bank/r11[1] ), .IN1(n6097), 
        .SEL(n6067), .F(\u_a23_core/u_execute/u_register_bank/n4921 ) );
  MUX U7878 ( .IN0(\u_a23_core/u_execute/u_register_bank/r11[0] ), .IN1(n6098), 
        .SEL(n6067), .F(\u_a23_core/u_execute/u_register_bank/n4919 ) );
  ANDN U7879 ( .A(\u_a23_core/reg_bank_wen[11] ), .B(n6099), .Z(n6067) );
  MUX U7880 ( .IN0(\u_a23_core/u_execute/u_register_bank/r14[31] ), .IN1(n6066), .SEL(n6100), .F(\u_a23_core/u_execute/u_register_bank/n4917 ) );
  MUX U7881 ( .IN0(\u_a23_core/u_execute/u_register_bank/r14[30] ), .IN1(n6068), .SEL(n6100), .F(\u_a23_core/u_execute/u_register_bank/n4915 ) );
  MUX U7882 ( .IN0(\u_a23_core/u_execute/u_register_bank/r14[29] ), .IN1(n6069), .SEL(n6100), .F(\u_a23_core/u_execute/u_register_bank/n4913 ) );
  MUX U7883 ( .IN0(\u_a23_core/u_execute/u_register_bank/r14[28] ), .IN1(n6070), .SEL(n6100), .F(\u_a23_core/u_execute/u_register_bank/n4911 ) );
  MUX U7884 ( .IN0(\u_a23_core/u_execute/u_register_bank/r14[27] ), .IN1(n6071), .SEL(n6100), .F(\u_a23_core/u_execute/u_register_bank/n4909 ) );
  MUX U7885 ( .IN0(\u_a23_core/u_execute/u_register_bank/r14[26] ), .IN1(n6072), .SEL(n6100), .F(\u_a23_core/u_execute/u_register_bank/n4907 ) );
  MUX U7886 ( .IN0(\u_a23_core/u_execute/u_register_bank/r14[25] ), .IN1(n6073), .SEL(n6100), .F(\u_a23_core/u_execute/u_register_bank/n4905 ) );
  MUX U7887 ( .IN0(\u_a23_core/u_execute/u_register_bank/r14[24] ), .IN1(n6074), .SEL(n6100), .F(\u_a23_core/u_execute/u_register_bank/n4903 ) );
  MUX U7888 ( .IN0(\u_a23_core/u_execute/u_register_bank/r14[23] ), .IN1(n6075), .SEL(n6100), .F(\u_a23_core/u_execute/u_register_bank/n4901 ) );
  MUX U7889 ( .IN0(\u_a23_core/u_execute/u_register_bank/r14[22] ), .IN1(n6076), .SEL(n6100), .F(\u_a23_core/u_execute/u_register_bank/n4899 ) );
  MUX U7890 ( .IN0(\u_a23_core/u_execute/u_register_bank/r14[21] ), .IN1(n6077), .SEL(n6100), .F(\u_a23_core/u_execute/u_register_bank/n4897 ) );
  MUX U7891 ( .IN0(\u_a23_core/u_execute/u_register_bank/r14[20] ), .IN1(n6078), .SEL(n6100), .F(\u_a23_core/u_execute/u_register_bank/n4895 ) );
  MUX U7892 ( .IN0(\u_a23_core/u_execute/u_register_bank/r14[19] ), .IN1(n6079), .SEL(n6100), .F(\u_a23_core/u_execute/u_register_bank/n4893 ) );
  MUX U7893 ( .IN0(\u_a23_core/u_execute/u_register_bank/r14[18] ), .IN1(n6080), .SEL(n6100), .F(\u_a23_core/u_execute/u_register_bank/n4891 ) );
  MUX U7894 ( .IN0(\u_a23_core/u_execute/u_register_bank/r14[17] ), .IN1(n6081), .SEL(n6100), .F(\u_a23_core/u_execute/u_register_bank/n4889 ) );
  MUX U7895 ( .IN0(\u_a23_core/u_execute/u_register_bank/r14[16] ), .IN1(n6082), .SEL(n6100), .F(\u_a23_core/u_execute/u_register_bank/n4887 ) );
  MUX U7896 ( .IN0(\u_a23_core/u_execute/u_register_bank/r14[15] ), .IN1(n6083), .SEL(n6100), .F(\u_a23_core/u_execute/u_register_bank/n4885 ) );
  MUX U7897 ( .IN0(\u_a23_core/u_execute/u_register_bank/r14[14] ), .IN1(n6084), .SEL(n6100), .F(\u_a23_core/u_execute/u_register_bank/n4883 ) );
  MUX U7898 ( .IN0(\u_a23_core/u_execute/u_register_bank/r14[13] ), .IN1(n6085), .SEL(n6100), .F(\u_a23_core/u_execute/u_register_bank/n4881 ) );
  MUX U7899 ( .IN0(\u_a23_core/u_execute/u_register_bank/r14[12] ), .IN1(n6086), .SEL(n6100), .F(\u_a23_core/u_execute/u_register_bank/n4879 ) );
  MUX U7900 ( .IN0(\u_a23_core/u_execute/u_register_bank/r14[11] ), .IN1(n6087), .SEL(n6100), .F(\u_a23_core/u_execute/u_register_bank/n4877 ) );
  MUX U7901 ( .IN0(\u_a23_core/u_execute/u_register_bank/r14[10] ), .IN1(n6088), .SEL(n6100), .F(\u_a23_core/u_execute/u_register_bank/n4875 ) );
  MUX U7902 ( .IN0(\u_a23_core/u_execute/u_register_bank/r14[9] ), .IN1(n6089), 
        .SEL(n6100), .F(\u_a23_core/u_execute/u_register_bank/n4873 ) );
  MUX U7903 ( .IN0(\u_a23_core/u_execute/u_register_bank/r14[8] ), .IN1(n6090), 
        .SEL(n6100), .F(\u_a23_core/u_execute/u_register_bank/n4871 ) );
  MUX U7904 ( .IN0(\u_a23_core/u_execute/u_register_bank/r14[7] ), .IN1(n6091), 
        .SEL(n6100), .F(\u_a23_core/u_execute/u_register_bank/n4869 ) );
  MUX U7905 ( .IN0(\u_a23_core/u_execute/u_register_bank/r14[6] ), .IN1(n6092), 
        .SEL(n6100), .F(\u_a23_core/u_execute/u_register_bank/n4867 ) );
  MUX U7906 ( .IN0(\u_a23_core/u_execute/u_register_bank/r14[5] ), .IN1(n6093), 
        .SEL(n6100), .F(\u_a23_core/u_execute/u_register_bank/n4865 ) );
  MUX U7907 ( .IN0(\u_a23_core/u_execute/u_register_bank/r14[4] ), .IN1(n6094), 
        .SEL(n6100), .F(\u_a23_core/u_execute/u_register_bank/n4863 ) );
  MUX U7908 ( .IN0(\u_a23_core/u_execute/u_register_bank/r14[3] ), .IN1(n6095), 
        .SEL(n6100), .F(\u_a23_core/u_execute/u_register_bank/n4861 ) );
  MUX U7909 ( .IN0(\u_a23_core/u_execute/u_register_bank/r14[2] ), .IN1(n6096), 
        .SEL(n6100), .F(\u_a23_core/u_execute/u_register_bank/n4859 ) );
  MUX U7910 ( .IN0(\u_a23_core/u_execute/u_register_bank/r14[1] ), .IN1(n6097), 
        .SEL(n6100), .F(\u_a23_core/u_execute/u_register_bank/n4857 ) );
  MUX U7911 ( .IN0(\u_a23_core/u_execute/u_register_bank/r14[0] ), .IN1(n6098), 
        .SEL(n6100), .F(\u_a23_core/u_execute/u_register_bank/n4855 ) );
  ANDN U7912 ( .A(\u_a23_core/reg_bank_wen[14] ), .B(n6099), .Z(n6100) );
  MUX U7913 ( .IN0(\u_a23_core/u_execute/u_register_bank/r13[31] ), .IN1(n6066), .SEL(n6101), .F(\u_a23_core/u_execute/u_register_bank/n4853 ) );
  MUX U7914 ( .IN0(\u_a23_core/u_execute/u_register_bank/r13[30] ), .IN1(n6068), .SEL(n6101), .F(\u_a23_core/u_execute/u_register_bank/n4851 ) );
  MUX U7915 ( .IN0(\u_a23_core/u_execute/u_register_bank/r13[29] ), .IN1(n6069), .SEL(n6101), .F(\u_a23_core/u_execute/u_register_bank/n4849 ) );
  MUX U7916 ( .IN0(\u_a23_core/u_execute/u_register_bank/r13[28] ), .IN1(n6070), .SEL(n6101), .F(\u_a23_core/u_execute/u_register_bank/n4847 ) );
  MUX U7917 ( .IN0(\u_a23_core/u_execute/u_register_bank/r13[27] ), .IN1(n6071), .SEL(n6101), .F(\u_a23_core/u_execute/u_register_bank/n4845 ) );
  MUX U7918 ( .IN0(\u_a23_core/u_execute/u_register_bank/r13[26] ), .IN1(n6072), .SEL(n6101), .F(\u_a23_core/u_execute/u_register_bank/n4843 ) );
  MUX U7919 ( .IN0(\u_a23_core/u_execute/u_register_bank/r13[25] ), .IN1(n6073), .SEL(n6101), .F(\u_a23_core/u_execute/u_register_bank/n4841 ) );
  MUX U7920 ( .IN0(\u_a23_core/u_execute/u_register_bank/r13[24] ), .IN1(n6074), .SEL(n6101), .F(\u_a23_core/u_execute/u_register_bank/n4839 ) );
  MUX U7921 ( .IN0(\u_a23_core/u_execute/u_register_bank/r13[23] ), .IN1(n6075), .SEL(n6101), .F(\u_a23_core/u_execute/u_register_bank/n4837 ) );
  MUX U7922 ( .IN0(\u_a23_core/u_execute/u_register_bank/r13[22] ), .IN1(n6076), .SEL(n6101), .F(\u_a23_core/u_execute/u_register_bank/n4835 ) );
  MUX U7923 ( .IN0(\u_a23_core/u_execute/u_register_bank/r13[21] ), .IN1(n6077), .SEL(n6101), .F(\u_a23_core/u_execute/u_register_bank/n4833 ) );
  MUX U7924 ( .IN0(\u_a23_core/u_execute/u_register_bank/r13[20] ), .IN1(n6078), .SEL(n6101), .F(\u_a23_core/u_execute/u_register_bank/n4831 ) );
  MUX U7925 ( .IN0(\u_a23_core/u_execute/u_register_bank/r13[19] ), .IN1(n6079), .SEL(n6101), .F(\u_a23_core/u_execute/u_register_bank/n4829 ) );
  MUX U7926 ( .IN0(\u_a23_core/u_execute/u_register_bank/r13[18] ), .IN1(n6080), .SEL(n6101), .F(\u_a23_core/u_execute/u_register_bank/n4827 ) );
  MUX U7927 ( .IN0(\u_a23_core/u_execute/u_register_bank/r13[17] ), .IN1(n6081), .SEL(n6101), .F(\u_a23_core/u_execute/u_register_bank/n4825 ) );
  MUX U7928 ( .IN0(\u_a23_core/u_execute/u_register_bank/r13[16] ), .IN1(n6082), .SEL(n6101), .F(\u_a23_core/u_execute/u_register_bank/n4823 ) );
  MUX U7929 ( .IN0(\u_a23_core/u_execute/u_register_bank/r13[15] ), .IN1(n6083), .SEL(n6101), .F(\u_a23_core/u_execute/u_register_bank/n4821 ) );
  MUX U7930 ( .IN0(\u_a23_core/u_execute/u_register_bank/r13[14] ), .IN1(n6084), .SEL(n6101), .F(\u_a23_core/u_execute/u_register_bank/n4819 ) );
  MUX U7931 ( .IN0(\u_a23_core/u_execute/u_register_bank/r13[13] ), .IN1(n6085), .SEL(n6101), .F(\u_a23_core/u_execute/u_register_bank/n4817 ) );
  MUX U7932 ( .IN0(\u_a23_core/u_execute/u_register_bank/r13[12] ), .IN1(n6086), .SEL(n6101), .F(\u_a23_core/u_execute/u_register_bank/n4815 ) );
  MUX U7933 ( .IN0(\u_a23_core/u_execute/u_register_bank/r13[11] ), .IN1(n6087), .SEL(n6101), .F(\u_a23_core/u_execute/u_register_bank/n4813 ) );
  MUX U7934 ( .IN0(\u_a23_core/u_execute/u_register_bank/r13[10] ), .IN1(n6088), .SEL(n6101), .F(\u_a23_core/u_execute/u_register_bank/n4811 ) );
  MUX U7935 ( .IN0(\u_a23_core/u_execute/u_register_bank/r13[9] ), .IN1(n6089), 
        .SEL(n6101), .F(\u_a23_core/u_execute/u_register_bank/n4809 ) );
  MUX U7936 ( .IN0(\u_a23_core/u_execute/u_register_bank/r13[8] ), .IN1(n6090), 
        .SEL(n6101), .F(\u_a23_core/u_execute/u_register_bank/n4807 ) );
  MUX U7937 ( .IN0(\u_a23_core/u_execute/u_register_bank/r13[7] ), .IN1(n6091), 
        .SEL(n6101), .F(\u_a23_core/u_execute/u_register_bank/n4805 ) );
  MUX U7938 ( .IN0(\u_a23_core/u_execute/u_register_bank/r13[6] ), .IN1(n6092), 
        .SEL(n6101), .F(\u_a23_core/u_execute/u_register_bank/n4803 ) );
  MUX U7939 ( .IN0(\u_a23_core/u_execute/u_register_bank/r13[5] ), .IN1(n6093), 
        .SEL(n6101), .F(\u_a23_core/u_execute/u_register_bank/n4801 ) );
  MUX U7940 ( .IN0(\u_a23_core/u_execute/u_register_bank/r13[4] ), .IN1(n6094), 
        .SEL(n6101), .F(\u_a23_core/u_execute/u_register_bank/n4799 ) );
  MUX U7941 ( .IN0(\u_a23_core/u_execute/u_register_bank/r13[3] ), .IN1(n6095), 
        .SEL(n6101), .F(\u_a23_core/u_execute/u_register_bank/n4797 ) );
  MUX U7942 ( .IN0(\u_a23_core/u_execute/u_register_bank/r13[2] ), .IN1(n6096), 
        .SEL(n6101), .F(\u_a23_core/u_execute/u_register_bank/n4795 ) );
  MUX U7943 ( .IN0(\u_a23_core/u_execute/u_register_bank/r13[1] ), .IN1(n6097), 
        .SEL(n6101), .F(\u_a23_core/u_execute/u_register_bank/n4793 ) );
  MUX U7944 ( .IN0(\u_a23_core/u_execute/u_register_bank/r13[0] ), .IN1(n6098), 
        .SEL(n6101), .F(\u_a23_core/u_execute/u_register_bank/n4791 ) );
  ANDN U7945 ( .A(\u_a23_core/reg_bank_wen[13] ), .B(n6099), .Z(n6101) );
  MUX U7946 ( .IN0(\u_a23_core/u_execute/u_register_bank/r12[31] ), .IN1(n6066), .SEL(n6102), .F(\u_a23_core/u_execute/u_register_bank/n4789 ) );
  MUX U7947 ( .IN0(\u_a23_core/u_execute/u_register_bank/r12[30] ), .IN1(n6068), .SEL(n6102), .F(\u_a23_core/u_execute/u_register_bank/n4787 ) );
  MUX U7948 ( .IN0(\u_a23_core/u_execute/u_register_bank/r12[29] ), .IN1(n6069), .SEL(n6102), .F(\u_a23_core/u_execute/u_register_bank/n4785 ) );
  MUX U7949 ( .IN0(\u_a23_core/u_execute/u_register_bank/r12[28] ), .IN1(n6070), .SEL(n6102), .F(\u_a23_core/u_execute/u_register_bank/n4783 ) );
  MUX U7950 ( .IN0(\u_a23_core/u_execute/u_register_bank/r12[27] ), .IN1(n6071), .SEL(n6102), .F(\u_a23_core/u_execute/u_register_bank/n4781 ) );
  MUX U7951 ( .IN0(\u_a23_core/u_execute/u_register_bank/r12[26] ), .IN1(n6072), .SEL(n6102), .F(\u_a23_core/u_execute/u_register_bank/n4779 ) );
  MUX U7952 ( .IN0(\u_a23_core/u_execute/u_register_bank/r12[25] ), .IN1(n6073), .SEL(n6102), .F(\u_a23_core/u_execute/u_register_bank/n4777 ) );
  MUX U7953 ( .IN0(\u_a23_core/u_execute/u_register_bank/r12[24] ), .IN1(n6074), .SEL(n6102), .F(\u_a23_core/u_execute/u_register_bank/n4775 ) );
  MUX U7954 ( .IN0(\u_a23_core/u_execute/u_register_bank/r12[23] ), .IN1(n6075), .SEL(n6102), .F(\u_a23_core/u_execute/u_register_bank/n4773 ) );
  MUX U7955 ( .IN0(\u_a23_core/u_execute/u_register_bank/r12[22] ), .IN1(n6076), .SEL(n6102), .F(\u_a23_core/u_execute/u_register_bank/n4771 ) );
  MUX U7956 ( .IN0(\u_a23_core/u_execute/u_register_bank/r12[21] ), .IN1(n6077), .SEL(n6102), .F(\u_a23_core/u_execute/u_register_bank/n4769 ) );
  MUX U7957 ( .IN0(\u_a23_core/u_execute/u_register_bank/r12[20] ), .IN1(n6078), .SEL(n6102), .F(\u_a23_core/u_execute/u_register_bank/n4767 ) );
  MUX U7958 ( .IN0(\u_a23_core/u_execute/u_register_bank/r12[19] ), .IN1(n6079), .SEL(n6102), .F(\u_a23_core/u_execute/u_register_bank/n4765 ) );
  MUX U7959 ( .IN0(\u_a23_core/u_execute/u_register_bank/r12[18] ), .IN1(n6080), .SEL(n6102), .F(\u_a23_core/u_execute/u_register_bank/n4763 ) );
  MUX U7960 ( .IN0(\u_a23_core/u_execute/u_register_bank/r12[17] ), .IN1(n6081), .SEL(n6102), .F(\u_a23_core/u_execute/u_register_bank/n4761 ) );
  MUX U7961 ( .IN0(\u_a23_core/u_execute/u_register_bank/r12[16] ), .IN1(n6082), .SEL(n6102), .F(\u_a23_core/u_execute/u_register_bank/n4759 ) );
  MUX U7962 ( .IN0(\u_a23_core/u_execute/u_register_bank/r12[15] ), .IN1(n6083), .SEL(n6102), .F(\u_a23_core/u_execute/u_register_bank/n4757 ) );
  MUX U7963 ( .IN0(\u_a23_core/u_execute/u_register_bank/r12[14] ), .IN1(n6084), .SEL(n6102), .F(\u_a23_core/u_execute/u_register_bank/n4755 ) );
  MUX U7964 ( .IN0(\u_a23_core/u_execute/u_register_bank/r12[13] ), .IN1(n6085), .SEL(n6102), .F(\u_a23_core/u_execute/u_register_bank/n4753 ) );
  MUX U7965 ( .IN0(\u_a23_core/u_execute/u_register_bank/r12[12] ), .IN1(n6086), .SEL(n6102), .F(\u_a23_core/u_execute/u_register_bank/n4751 ) );
  MUX U7966 ( .IN0(\u_a23_core/u_execute/u_register_bank/r12[11] ), .IN1(n6087), .SEL(n6102), .F(\u_a23_core/u_execute/u_register_bank/n4749 ) );
  MUX U7967 ( .IN0(\u_a23_core/u_execute/u_register_bank/r12[10] ), .IN1(n6088), .SEL(n6102), .F(\u_a23_core/u_execute/u_register_bank/n4747 ) );
  MUX U7968 ( .IN0(\u_a23_core/u_execute/u_register_bank/r12[9] ), .IN1(n6089), 
        .SEL(n6102), .F(\u_a23_core/u_execute/u_register_bank/n4745 ) );
  MUX U7969 ( .IN0(\u_a23_core/u_execute/u_register_bank/r12[8] ), .IN1(n6090), 
        .SEL(n6102), .F(\u_a23_core/u_execute/u_register_bank/n4743 ) );
  MUX U7970 ( .IN0(\u_a23_core/u_execute/u_register_bank/r12[7] ), .IN1(n6091), 
        .SEL(n6102), .F(\u_a23_core/u_execute/u_register_bank/n4741 ) );
  MUX U7971 ( .IN0(\u_a23_core/u_execute/u_register_bank/r12[6] ), .IN1(n6092), 
        .SEL(n6102), .F(\u_a23_core/u_execute/u_register_bank/n4739 ) );
  MUX U7972 ( .IN0(\u_a23_core/u_execute/u_register_bank/r12[5] ), .IN1(n6093), 
        .SEL(n6102), .F(\u_a23_core/u_execute/u_register_bank/n4737 ) );
  MUX U7973 ( .IN0(\u_a23_core/u_execute/u_register_bank/r12[4] ), .IN1(n6094), 
        .SEL(n6102), .F(\u_a23_core/u_execute/u_register_bank/n4735 ) );
  MUX U7974 ( .IN0(\u_a23_core/u_execute/u_register_bank/r12[3] ), .IN1(n6095), 
        .SEL(n6102), .F(\u_a23_core/u_execute/u_register_bank/n4733 ) );
  MUX U7975 ( .IN0(\u_a23_core/u_execute/u_register_bank/r12[2] ), .IN1(n6096), 
        .SEL(n6102), .F(\u_a23_core/u_execute/u_register_bank/n4731 ) );
  MUX U7976 ( .IN0(\u_a23_core/u_execute/u_register_bank/r12[1] ), .IN1(n6097), 
        .SEL(n6102), .F(\u_a23_core/u_execute/u_register_bank/n4729 ) );
  MUX U7977 ( .IN0(\u_a23_core/u_execute/u_register_bank/r12[0] ), .IN1(n6098), 
        .SEL(n6102), .F(\u_a23_core/u_execute/u_register_bank/n4727 ) );
  ANDN U7978 ( .A(\u_a23_core/reg_bank_wen[12] ), .B(n6099), .Z(n6102) );
  MUX U7979 ( .IN0(\u_a23_core/u_execute/pc[25] ), .IN1(n5971), .SEL(
        \u_a23_core/pc_wen ), .F(\u_a23_core/u_execute/u_register_bank/n4725 )
         );
  NAND U7980 ( .A(n6103), .B(n6104), .Z(n5971) );
  NAND U7981 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[25] ), .B(n6105), 
        .Z(n6104) );
  AND U7982 ( .A(n6106), .B(n6107), .Z(n6103) );
  NAND U7983 ( .A(n6108), .B(\u_a23_core/u_execute/pc_plus4[25] ), .Z(n6107)
         );
  NANDN U7984 ( .B(n6109), .A(\u_a23_core/u_execute/pc_minus4[25] ), .Z(n6106)
         );
  MUX U7985 ( .IN0(\u_a23_core/u_execute/pc[24] ), .IN1(n5976), .SEL(
        \u_a23_core/pc_wen ), .F(\u_a23_core/u_execute/u_register_bank/n4723 )
         );
  NAND U7986 ( .A(n6110), .B(n6111), .Z(n5976) );
  NAND U7987 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[24] ), .B(n6105), 
        .Z(n6111) );
  AND U7988 ( .A(n6112), .B(n6113), .Z(n6110) );
  NAND U7989 ( .A(n6108), .B(\u_a23_core/u_execute/pc_plus4[24] ), .Z(n6113)
         );
  NANDN U7990 ( .B(n6109), .A(\u_a23_core/u_execute/pc_minus4[24] ), .Z(n6112)
         );
  MUX U7991 ( .IN0(\u_a23_core/u_execute/pc[23] ), .IN1(n5981), .SEL(
        \u_a23_core/pc_wen ), .F(\u_a23_core/u_execute/u_register_bank/n4721 )
         );
  NAND U7992 ( .A(n6114), .B(n6115), .Z(n5981) );
  NAND U7993 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[23] ), .B(n6105), 
        .Z(n6115) );
  AND U7994 ( .A(n6116), .B(n6117), .Z(n6114) );
  NAND U7995 ( .A(n6108), .B(\u_a23_core/u_execute/pc_plus4[23] ), .Z(n6117)
         );
  NANDN U7996 ( .B(n6109), .A(\u_a23_core/u_execute/pc_minus4[23] ), .Z(n6116)
         );
  MUX U7997 ( .IN0(\u_a23_core/u_execute/pc[22] ), .IN1(n5986), .SEL(
        \u_a23_core/pc_wen ), .F(\u_a23_core/u_execute/u_register_bank/n4719 )
         );
  NAND U7998 ( .A(n6118), .B(n6119), .Z(n5986) );
  NAND U7999 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[22] ), .B(n6105), 
        .Z(n6119) );
  AND U8000 ( .A(n6120), .B(n6121), .Z(n6118) );
  NAND U8001 ( .A(n6108), .B(\u_a23_core/u_execute/pc_plus4[22] ), .Z(n6121)
         );
  NANDN U8002 ( .B(n6109), .A(\u_a23_core/u_execute/pc_minus4[22] ), .Z(n6120)
         );
  MUX U8003 ( .IN0(\u_a23_core/u_execute/pc[21] ), .IN1(n5991), .SEL(
        \u_a23_core/pc_wen ), .F(\u_a23_core/u_execute/u_register_bank/n4717 )
         );
  NAND U8004 ( .A(n6122), .B(n6123), .Z(n5991) );
  NAND U8005 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[21] ), .B(n6105), 
        .Z(n6123) );
  AND U8006 ( .A(n6124), .B(n6125), .Z(n6122) );
  NAND U8007 ( .A(n6108), .B(\u_a23_core/u_execute/pc_plus4[21] ), .Z(n6125)
         );
  NANDN U8008 ( .B(n6109), .A(\u_a23_core/u_execute/pc_minus4[21] ), .Z(n6124)
         );
  MUX U8009 ( .IN0(\u_a23_core/u_execute/pc[20] ), .IN1(n5996), .SEL(
        \u_a23_core/pc_wen ), .F(\u_a23_core/u_execute/u_register_bank/n4715 )
         );
  NAND U8010 ( .A(n6126), .B(n6127), .Z(n5996) );
  NAND U8011 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[20] ), .B(n6105), 
        .Z(n6127) );
  AND U8012 ( .A(n6128), .B(n6129), .Z(n6126) );
  NAND U8013 ( .A(n6108), .B(\u_a23_core/u_execute/pc_plus4[20] ), .Z(n6129)
         );
  NANDN U8014 ( .B(n6109), .A(\u_a23_core/u_execute/pc_minus4[20] ), .Z(n6128)
         );
  MUX U8015 ( .IN0(\u_a23_core/u_execute/pc[19] ), .IN1(n6001), .SEL(
        \u_a23_core/pc_wen ), .F(\u_a23_core/u_execute/u_register_bank/n4713 )
         );
  NAND U8016 ( .A(n6130), .B(n6131), .Z(n6001) );
  NAND U8017 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[19] ), .B(n6105), 
        .Z(n6131) );
  AND U8018 ( .A(n6132), .B(n6133), .Z(n6130) );
  NAND U8019 ( .A(n6108), .B(\u_a23_core/u_execute/pc_plus4[19] ), .Z(n6133)
         );
  NANDN U8020 ( .B(n6109), .A(\u_a23_core/u_execute/pc_minus4[19] ), .Z(n6132)
         );
  MUX U8021 ( .IN0(\u_a23_core/u_execute/pc[18] ), .IN1(n6006), .SEL(
        \u_a23_core/pc_wen ), .F(\u_a23_core/u_execute/u_register_bank/n4711 )
         );
  NAND U8022 ( .A(n6134), .B(n6135), .Z(n6006) );
  NAND U8023 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[18] ), .B(n6105), 
        .Z(n6135) );
  AND U8024 ( .A(n6136), .B(n6137), .Z(n6134) );
  NAND U8025 ( .A(n6108), .B(\u_a23_core/u_execute/pc_plus4[18] ), .Z(n6137)
         );
  NANDN U8026 ( .B(n6109), .A(\u_a23_core/u_execute/pc_minus4[18] ), .Z(n6136)
         );
  MUX U8027 ( .IN0(\u_a23_core/u_execute/pc[17] ), .IN1(n6011), .SEL(
        \u_a23_core/pc_wen ), .F(\u_a23_core/u_execute/u_register_bank/n4709 )
         );
  NAND U8028 ( .A(n6138), .B(n6139), .Z(n6011) );
  NAND U8029 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[17] ), .B(n6105), 
        .Z(n6139) );
  AND U8030 ( .A(n6140), .B(n6141), .Z(n6138) );
  NAND U8031 ( .A(n6108), .B(\u_a23_core/u_execute/pc_plus4[17] ), .Z(n6141)
         );
  NANDN U8032 ( .B(n6109), .A(\u_a23_core/u_execute/pc_minus4[17] ), .Z(n6140)
         );
  MUX U8033 ( .IN0(\u_a23_core/u_execute/pc[16] ), .IN1(n6016), .SEL(
        \u_a23_core/pc_wen ), .F(\u_a23_core/u_execute/u_register_bank/n4707 )
         );
  NAND U8034 ( .A(n6142), .B(n6143), .Z(n6016) );
  NAND U8035 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[16] ), .B(n6105), 
        .Z(n6143) );
  AND U8036 ( .A(n6144), .B(n6145), .Z(n6142) );
  NAND U8037 ( .A(n6108), .B(\u_a23_core/u_execute/pc_plus4[16] ), .Z(n6145)
         );
  NANDN U8038 ( .B(n6109), .A(\u_a23_core/u_execute/pc_minus4[16] ), .Z(n6144)
         );
  MUX U8039 ( .IN0(\u_a23_core/u_execute/pc[15] ), .IN1(n6021), .SEL(
        \u_a23_core/pc_wen ), .F(\u_a23_core/u_execute/u_register_bank/n4705 )
         );
  NAND U8040 ( .A(n6146), .B(n6147), .Z(n6021) );
  NAND U8041 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[15] ), .B(n6105), 
        .Z(n6147) );
  AND U8042 ( .A(n6148), .B(n6149), .Z(n6146) );
  NAND U8043 ( .A(n6108), .B(\u_a23_core/u_execute/pc_plus4[15] ), .Z(n6149)
         );
  NANDN U8044 ( .B(n6109), .A(\u_a23_core/u_execute/pc_minus4[15] ), .Z(n6148)
         );
  MUX U8045 ( .IN0(\u_a23_core/u_execute/pc[14] ), .IN1(n6030), .SEL(
        \u_a23_core/pc_wen ), .F(\u_a23_core/u_execute/u_register_bank/n4703 )
         );
  NAND U8046 ( .A(n6150), .B(n6151), .Z(n6030) );
  NAND U8047 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[14] ), .B(n6105), 
        .Z(n6151) );
  AND U8048 ( .A(n6152), .B(n6153), .Z(n6150) );
  NAND U8049 ( .A(n6108), .B(\u_a23_core/u_execute/pc_plus4[14] ), .Z(n6153)
         );
  NANDN U8050 ( .B(n6109), .A(\u_a23_core/u_execute/pc_minus4[14] ), .Z(n6152)
         );
  MUX U8051 ( .IN0(\u_a23_core/u_execute/pc[13] ), .IN1(n6038), .SEL(
        \u_a23_core/pc_wen ), .F(\u_a23_core/u_execute/u_register_bank/n4701 )
         );
  NAND U8052 ( .A(n6154), .B(n6155), .Z(n6038) );
  NAND U8053 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[13] ), .B(n6105), 
        .Z(n6155) );
  AND U8054 ( .A(n6156), .B(n6157), .Z(n6154) );
  NAND U8055 ( .A(n6108), .B(\u_a23_core/u_execute/pc_plus4[13] ), .Z(n6157)
         );
  NANDN U8056 ( .B(n6109), .A(\u_a23_core/u_execute/pc_minus4[13] ), .Z(n6156)
         );
  MUX U8057 ( .IN0(\u_a23_core/u_execute/pc[12] ), .IN1(n6046), .SEL(
        \u_a23_core/pc_wen ), .F(\u_a23_core/u_execute/u_register_bank/n4699 )
         );
  NAND U8058 ( .A(n6158), .B(n6159), .Z(n6046) );
  NAND U8059 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[12] ), .B(n6105), 
        .Z(n6159) );
  AND U8060 ( .A(n6160), .B(n6161), .Z(n6158) );
  NAND U8061 ( .A(n6108), .B(\u_a23_core/u_execute/pc_plus4[12] ), .Z(n6161)
         );
  NANDN U8062 ( .B(n6109), .A(\u_a23_core/u_execute/pc_minus4[12] ), .Z(n6160)
         );
  MUX U8063 ( .IN0(\u_a23_core/u_execute/pc[11] ), .IN1(n6054), .SEL(
        \u_a23_core/pc_wen ), .F(\u_a23_core/u_execute/u_register_bank/n4697 )
         );
  NAND U8064 ( .A(n6162), .B(n6163), .Z(n6054) );
  NAND U8065 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[11] ), .B(n6105), 
        .Z(n6163) );
  AND U8066 ( .A(n6164), .B(n6165), .Z(n6162) );
  NAND U8067 ( .A(n6108), .B(\u_a23_core/u_execute/pc_plus4[11] ), .Z(n6165)
         );
  NANDN U8068 ( .B(n6109), .A(\u_a23_core/u_execute/pc_minus4[11] ), .Z(n6164)
         );
  MUX U8069 ( .IN0(\u_a23_core/u_execute/pc[10] ), .IN1(n6062), .SEL(
        \u_a23_core/pc_wen ), .F(\u_a23_core/u_execute/u_register_bank/n4695 )
         );
  NAND U8070 ( .A(n6166), .B(n6167), .Z(n6062) );
  NAND U8071 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[10] ), .B(n6105), 
        .Z(n6167) );
  AND U8072 ( .A(n6168), .B(n6169), .Z(n6166) );
  NAND U8073 ( .A(n6108), .B(\u_a23_core/u_execute/pc_plus4[10] ), .Z(n6169)
         );
  NANDN U8074 ( .B(n6109), .A(\u_a23_core/u_execute/pc_minus4[10] ), .Z(n6168)
         );
  MUX U8075 ( .IN0(\u_a23_core/u_execute/pc[9] ), .IN1(n5937), .SEL(
        \u_a23_core/pc_wen ), .F(\u_a23_core/u_execute/u_register_bank/n4693 )
         );
  NAND U8076 ( .A(n6170), .B(n6171), .Z(n5937) );
  NAND U8077 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[9] ), .B(n6105), 
        .Z(n6171) );
  AND U8078 ( .A(n6172), .B(n6173), .Z(n6170) );
  NAND U8079 ( .A(n6108), .B(\u_a23_core/u_execute/pc_plus4[9] ), .Z(n6173) );
  NANDN U8080 ( .B(n6109), .A(\u_a23_core/u_execute/pc_minus4[9] ), .Z(n6172)
         );
  MUX U8081 ( .IN0(\u_a23_core/u_execute/pc[8] ), .IN1(n5944), .SEL(
        \u_a23_core/pc_wen ), .F(\u_a23_core/u_execute/u_register_bank/n4691 )
         );
  NAND U8082 ( .A(n6174), .B(n6175), .Z(n5944) );
  NAND U8083 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[8] ), .B(n6105), 
        .Z(n6175) );
  AND U8084 ( .A(n6176), .B(n6177), .Z(n6174) );
  NAND U8085 ( .A(n6108), .B(\u_a23_core/u_execute/pc_plus4[8] ), .Z(n6177) );
  NANDN U8086 ( .B(n6109), .A(\u_a23_core/u_execute/pc_minus4[8] ), .Z(n6176)
         );
  MUX U8087 ( .IN0(\u_a23_core/u_execute/pc[7] ), .IN1(n6024), .SEL(
        \u_a23_core/pc_wen ), .F(\u_a23_core/u_execute/u_register_bank/n4689 )
         );
  NAND U8088 ( .A(n6178), .B(n6179), .Z(n6024) );
  NAND U8089 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[7] ), .B(n6105), 
        .Z(n6179) );
  AND U8090 ( .A(n6180), .B(n6181), .Z(n6178) );
  NAND U8091 ( .A(n6108), .B(\u_a23_core/u_execute/pc_plus4[7] ), .Z(n6181) );
  NANDN U8092 ( .B(n6109), .A(\u_a23_core/u_execute/pc_minus4[7] ), .Z(n6180)
         );
  MUX U8093 ( .IN0(\u_a23_core/u_execute/pc[6] ), .IN1(n6033), .SEL(
        \u_a23_core/pc_wen ), .F(\u_a23_core/u_execute/u_register_bank/n4687 )
         );
  NAND U8094 ( .A(n6182), .B(n6183), .Z(n6033) );
  NAND U8095 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[6] ), .B(n6105), 
        .Z(n6183) );
  AND U8096 ( .A(n6184), .B(n6185), .Z(n6182) );
  NAND U8097 ( .A(n6108), .B(\u_a23_core/u_execute/pc_plus4[6] ), .Z(n6185) );
  NANDN U8098 ( .B(n6109), .A(\u_a23_core/u_execute/pc_minus4[6] ), .Z(n6184)
         );
  MUX U8099 ( .IN0(\u_a23_core/u_execute/pc[5] ), .IN1(n6041), .SEL(
        \u_a23_core/pc_wen ), .F(\u_a23_core/u_execute/u_register_bank/n4685 )
         );
  NAND U8100 ( .A(n6186), .B(n6187), .Z(n6041) );
  NAND U8101 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[5] ), .B(n6105), 
        .Z(n6187) );
  AND U8102 ( .A(n6188), .B(n6189), .Z(n6186) );
  NAND U8103 ( .A(n6108), .B(\u_a23_core/u_execute/pc_plus4[5] ), .Z(n6189) );
  NANDN U8104 ( .B(n6109), .A(\u_a23_core/u_execute/pc_minus4[5] ), .Z(n6188)
         );
  MUX U8105 ( .IN0(\u_a23_core/u_execute/pc[4] ), .IN1(n6049), .SEL(
        \u_a23_core/pc_wen ), .F(\u_a23_core/u_execute/u_register_bank/n4683 )
         );
  NAND U8106 ( .A(n6190), .B(n6191), .Z(n6049) );
  NAND U8107 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[4] ), .B(n6105), 
        .Z(n6191) );
  AND U8108 ( .A(n6192), .B(n6193), .Z(n6190) );
  NAND U8109 ( .A(n6108), .B(\u_a23_core/u_execute/pc_plus4[4] ), .Z(n6193) );
  NANDN U8110 ( .B(n6109), .A(\u_a23_core/u_execute/pc_minus4[4] ), .Z(n6192)
         );
  MUX U8111 ( .IN0(\u_a23_core/u_execute/pc[3] ), .IN1(n6057), .SEL(
        \u_a23_core/pc_wen ), .F(\u_a23_core/u_execute/u_register_bank/n4681 )
         );
  NAND U8112 ( .A(n6194), .B(n6195), .Z(n6057) );
  NAND U8113 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[3] ), .B(n6105), 
        .Z(n6195) );
  AND U8114 ( .A(n6196), .B(n6197), .Z(n6194) );
  NAND U8115 ( .A(n6108), .B(\u_a23_core/u_execute/pc_plus4[3] ), .Z(n6197) );
  IV U8116 ( .A(n6198), .Z(n6108) );
  NANDN U8117 ( .B(n6109), .A(\u_a23_core/u_execute/pc_minus4[3] ), .Z(n6196)
         );
  MUX U8118 ( .IN0(\u_a23_core/u_execute/pc[2] ), .IN1(n6065), .SEL(
        \u_a23_core/pc_wen ), .F(\u_a23_core/u_execute/u_register_bank/n4679 )
         );
  NAND U8119 ( .A(n6199), .B(n6200), .Z(n6065) );
  NAND U8120 ( .A(n6201), .B(n6202), .Z(n6200) );
  NAND U8121 ( .A(n6198), .B(n6109), .Z(n6202) );
  NAND U8122 ( .A(n6099), .B(\u_a23_core/pc_sel[1] ), .Z(n6109) );
  OR U8123 ( .A(\u_a23_core/pc_sel[1] ), .B(\u_a23_core/pc_sel[0] ), .Z(n6198)
         );
  NAND U8124 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[2] ), .B(n6105), 
        .Z(n6199) );
  MUX U8125 ( .IN0(\u_a23_core/pc_sel[0] ), .IN1(n5930), .SEL(
        \u_a23_core/pc_sel[1] ), .F(n6105) );
  MUX U8126 ( .IN0(\u_a23_core/u_execute/u_register_bank/r0[31] ), .IN1(n6066), 
        .SEL(n6203), .F(\u_a23_core/u_execute/u_register_bank/n4677 ) );
  MUX U8127 ( .IN0(\u_a23_core/u_execute/u_register_bank/r0[30] ), .IN1(n6068), 
        .SEL(n6203), .F(\u_a23_core/u_execute/u_register_bank/n4675 ) );
  MUX U8128 ( .IN0(\u_a23_core/u_execute/u_register_bank/r0[29] ), .IN1(n6069), 
        .SEL(n6203), .F(\u_a23_core/u_execute/u_register_bank/n4673 ) );
  MUX U8129 ( .IN0(\u_a23_core/u_execute/u_register_bank/r0[28] ), .IN1(n6070), 
        .SEL(n6203), .F(\u_a23_core/u_execute/u_register_bank/n4671 ) );
  MUX U8130 ( .IN0(\u_a23_core/u_execute/u_register_bank/r0[27] ), .IN1(n6071), 
        .SEL(n6203), .F(\u_a23_core/u_execute/u_register_bank/n4669 ) );
  MUX U8131 ( .IN0(\u_a23_core/u_execute/u_register_bank/r0[26] ), .IN1(n6072), 
        .SEL(n6203), .F(\u_a23_core/u_execute/u_register_bank/n4667 ) );
  MUX U8132 ( .IN0(\u_a23_core/u_execute/u_register_bank/r0[25] ), .IN1(n6073), 
        .SEL(n6203), .F(\u_a23_core/u_execute/u_register_bank/n4665 ) );
  MUX U8133 ( .IN0(\u_a23_core/u_execute/u_register_bank/r0[24] ), .IN1(n6074), 
        .SEL(n6203), .F(\u_a23_core/u_execute/u_register_bank/n4663 ) );
  MUX U8134 ( .IN0(\u_a23_core/u_execute/u_register_bank/r0[23] ), .IN1(n6075), 
        .SEL(n6203), .F(\u_a23_core/u_execute/u_register_bank/n4661 ) );
  MUX U8135 ( .IN0(\u_a23_core/u_execute/u_register_bank/r0[22] ), .IN1(n6076), 
        .SEL(n6203), .F(\u_a23_core/u_execute/u_register_bank/n4659 ) );
  MUX U8136 ( .IN0(\u_a23_core/u_execute/u_register_bank/r0[21] ), .IN1(n6077), 
        .SEL(n6203), .F(\u_a23_core/u_execute/u_register_bank/n4657 ) );
  MUX U8137 ( .IN0(\u_a23_core/u_execute/u_register_bank/r0[20] ), .IN1(n6078), 
        .SEL(n6203), .F(\u_a23_core/u_execute/u_register_bank/n4655 ) );
  MUX U8138 ( .IN0(\u_a23_core/u_execute/u_register_bank/r0[19] ), .IN1(n6079), 
        .SEL(n6203), .F(\u_a23_core/u_execute/u_register_bank/n4653 ) );
  MUX U8139 ( .IN0(\u_a23_core/u_execute/u_register_bank/r0[18] ), .IN1(n6080), 
        .SEL(n6203), .F(\u_a23_core/u_execute/u_register_bank/n4651 ) );
  MUX U8140 ( .IN0(\u_a23_core/u_execute/u_register_bank/r0[17] ), .IN1(n6081), 
        .SEL(n6203), .F(\u_a23_core/u_execute/u_register_bank/n4649 ) );
  MUX U8141 ( .IN0(\u_a23_core/u_execute/u_register_bank/r0[16] ), .IN1(n6082), 
        .SEL(n6203), .F(\u_a23_core/u_execute/u_register_bank/n4647 ) );
  MUX U8142 ( .IN0(\u_a23_core/u_execute/u_register_bank/r0[15] ), .IN1(n6083), 
        .SEL(n6203), .F(\u_a23_core/u_execute/u_register_bank/n4645 ) );
  MUX U8143 ( .IN0(\u_a23_core/u_execute/u_register_bank/r0[14] ), .IN1(n6084), 
        .SEL(n6203), .F(\u_a23_core/u_execute/u_register_bank/n4643 ) );
  MUX U8144 ( .IN0(\u_a23_core/u_execute/u_register_bank/r0[13] ), .IN1(n6085), 
        .SEL(n6203), .F(\u_a23_core/u_execute/u_register_bank/n4641 ) );
  MUX U8145 ( .IN0(\u_a23_core/u_execute/u_register_bank/r0[12] ), .IN1(n6086), 
        .SEL(n6203), .F(\u_a23_core/u_execute/u_register_bank/n4639 ) );
  MUX U8146 ( .IN0(\u_a23_core/u_execute/u_register_bank/r0[11] ), .IN1(n6087), 
        .SEL(n6203), .F(\u_a23_core/u_execute/u_register_bank/n4637 ) );
  MUX U8147 ( .IN0(\u_a23_core/u_execute/u_register_bank/r0[10] ), .IN1(n6088), 
        .SEL(n6203), .F(\u_a23_core/u_execute/u_register_bank/n4635 ) );
  MUX U8148 ( .IN0(\u_a23_core/u_execute/u_register_bank/r0[9] ), .IN1(n6089), 
        .SEL(n6203), .F(\u_a23_core/u_execute/u_register_bank/n4633 ) );
  MUX U8149 ( .IN0(\u_a23_core/u_execute/u_register_bank/r0[8] ), .IN1(n6090), 
        .SEL(n6203), .F(\u_a23_core/u_execute/u_register_bank/n4631 ) );
  MUX U8150 ( .IN0(\u_a23_core/u_execute/u_register_bank/r0[7] ), .IN1(n6091), 
        .SEL(n6203), .F(\u_a23_core/u_execute/u_register_bank/n4629 ) );
  MUX U8151 ( .IN0(\u_a23_core/u_execute/u_register_bank/r0[6] ), .IN1(n6092), 
        .SEL(n6203), .F(\u_a23_core/u_execute/u_register_bank/n4627 ) );
  MUX U8152 ( .IN0(\u_a23_core/u_execute/u_register_bank/r0[5] ), .IN1(n6093), 
        .SEL(n6203), .F(\u_a23_core/u_execute/u_register_bank/n4625 ) );
  MUX U8153 ( .IN0(\u_a23_core/u_execute/u_register_bank/r0[4] ), .IN1(n6094), 
        .SEL(n6203), .F(\u_a23_core/u_execute/u_register_bank/n4623 ) );
  MUX U8154 ( .IN0(\u_a23_core/u_execute/u_register_bank/r0[3] ), .IN1(n6095), 
        .SEL(n6203), .F(\u_a23_core/u_execute/u_register_bank/n4621 ) );
  MUX U8155 ( .IN0(\u_a23_core/u_execute/u_register_bank/r0[2] ), .IN1(n6096), 
        .SEL(n6203), .F(\u_a23_core/u_execute/u_register_bank/n4619 ) );
  MUX U8156 ( .IN0(\u_a23_core/u_execute/u_register_bank/r0[1] ), .IN1(n6097), 
        .SEL(n6203), .F(\u_a23_core/u_execute/u_register_bank/n4617 ) );
  MUX U8157 ( .IN0(\u_a23_core/u_execute/u_register_bank/r0[0] ), .IN1(n6098), 
        .SEL(n6203), .F(\u_a23_core/u_execute/u_register_bank/n4615 ) );
  ANDN U8158 ( .A(\u_a23_core/reg_bank_wen[0] ), .B(n6099), .Z(n6203) );
  MUX U8159 ( .IN0(\u_a23_core/u_execute/u_register_bank/r1[31] ), .IN1(n6066), 
        .SEL(n6204), .F(\u_a23_core/u_execute/u_register_bank/n4613 ) );
  MUX U8160 ( .IN0(\u_a23_core/u_execute/u_register_bank/r1[30] ), .IN1(n6068), 
        .SEL(n6204), .F(\u_a23_core/u_execute/u_register_bank/n4611 ) );
  MUX U8161 ( .IN0(\u_a23_core/u_execute/u_register_bank/r1[29] ), .IN1(n6069), 
        .SEL(n6204), .F(\u_a23_core/u_execute/u_register_bank/n4609 ) );
  MUX U8162 ( .IN0(\u_a23_core/u_execute/u_register_bank/r1[28] ), .IN1(n6070), 
        .SEL(n6204), .F(\u_a23_core/u_execute/u_register_bank/n4607 ) );
  MUX U8163 ( .IN0(\u_a23_core/u_execute/u_register_bank/r1[27] ), .IN1(n6071), 
        .SEL(n6204), .F(\u_a23_core/u_execute/u_register_bank/n4605 ) );
  MUX U8164 ( .IN0(\u_a23_core/u_execute/u_register_bank/r1[26] ), .IN1(n6072), 
        .SEL(n6204), .F(\u_a23_core/u_execute/u_register_bank/n4603 ) );
  MUX U8165 ( .IN0(\u_a23_core/u_execute/u_register_bank/r1[25] ), .IN1(n6073), 
        .SEL(n6204), .F(\u_a23_core/u_execute/u_register_bank/n4601 ) );
  MUX U8166 ( .IN0(\u_a23_core/u_execute/u_register_bank/r1[24] ), .IN1(n6074), 
        .SEL(n6204), .F(\u_a23_core/u_execute/u_register_bank/n4599 ) );
  MUX U8167 ( .IN0(\u_a23_core/u_execute/u_register_bank/r1[23] ), .IN1(n6075), 
        .SEL(n6204), .F(\u_a23_core/u_execute/u_register_bank/n4597 ) );
  MUX U8168 ( .IN0(\u_a23_core/u_execute/u_register_bank/r1[22] ), .IN1(n6076), 
        .SEL(n6204), .F(\u_a23_core/u_execute/u_register_bank/n4595 ) );
  MUX U8169 ( .IN0(\u_a23_core/u_execute/u_register_bank/r1[21] ), .IN1(n6077), 
        .SEL(n6204), .F(\u_a23_core/u_execute/u_register_bank/n4593 ) );
  MUX U8170 ( .IN0(\u_a23_core/u_execute/u_register_bank/r1[20] ), .IN1(n6078), 
        .SEL(n6204), .F(\u_a23_core/u_execute/u_register_bank/n4591 ) );
  MUX U8171 ( .IN0(\u_a23_core/u_execute/u_register_bank/r1[19] ), .IN1(n6079), 
        .SEL(n6204), .F(\u_a23_core/u_execute/u_register_bank/n4589 ) );
  MUX U8172 ( .IN0(\u_a23_core/u_execute/u_register_bank/r1[18] ), .IN1(n6080), 
        .SEL(n6204), .F(\u_a23_core/u_execute/u_register_bank/n4587 ) );
  MUX U8173 ( .IN0(\u_a23_core/u_execute/u_register_bank/r1[17] ), .IN1(n6081), 
        .SEL(n6204), .F(\u_a23_core/u_execute/u_register_bank/n4585 ) );
  MUX U8174 ( .IN0(\u_a23_core/u_execute/u_register_bank/r1[16] ), .IN1(n6082), 
        .SEL(n6204), .F(\u_a23_core/u_execute/u_register_bank/n4583 ) );
  MUX U8175 ( .IN0(\u_a23_core/u_execute/u_register_bank/r1[15] ), .IN1(n6083), 
        .SEL(n6204), .F(\u_a23_core/u_execute/u_register_bank/n4581 ) );
  MUX U8176 ( .IN0(\u_a23_core/u_execute/u_register_bank/r1[14] ), .IN1(n6084), 
        .SEL(n6204), .F(\u_a23_core/u_execute/u_register_bank/n4579 ) );
  MUX U8177 ( .IN0(\u_a23_core/u_execute/u_register_bank/r1[13] ), .IN1(n6085), 
        .SEL(n6204), .F(\u_a23_core/u_execute/u_register_bank/n4577 ) );
  MUX U8178 ( .IN0(\u_a23_core/u_execute/u_register_bank/r1[12] ), .IN1(n6086), 
        .SEL(n6204), .F(\u_a23_core/u_execute/u_register_bank/n4575 ) );
  MUX U8179 ( .IN0(\u_a23_core/u_execute/u_register_bank/r1[11] ), .IN1(n6087), 
        .SEL(n6204), .F(\u_a23_core/u_execute/u_register_bank/n4573 ) );
  MUX U8180 ( .IN0(\u_a23_core/u_execute/u_register_bank/r1[10] ), .IN1(n6088), 
        .SEL(n6204), .F(\u_a23_core/u_execute/u_register_bank/n4571 ) );
  MUX U8181 ( .IN0(\u_a23_core/u_execute/u_register_bank/r1[9] ), .IN1(n6089), 
        .SEL(n6204), .F(\u_a23_core/u_execute/u_register_bank/n4569 ) );
  MUX U8182 ( .IN0(\u_a23_core/u_execute/u_register_bank/r1[8] ), .IN1(n6090), 
        .SEL(n6204), .F(\u_a23_core/u_execute/u_register_bank/n4567 ) );
  MUX U8183 ( .IN0(\u_a23_core/u_execute/u_register_bank/r1[7] ), .IN1(n6091), 
        .SEL(n6204), .F(\u_a23_core/u_execute/u_register_bank/n4565 ) );
  MUX U8184 ( .IN0(\u_a23_core/u_execute/u_register_bank/r1[6] ), .IN1(n6092), 
        .SEL(n6204), .F(\u_a23_core/u_execute/u_register_bank/n4563 ) );
  MUX U8185 ( .IN0(\u_a23_core/u_execute/u_register_bank/r1[5] ), .IN1(n6093), 
        .SEL(n6204), .F(\u_a23_core/u_execute/u_register_bank/n4561 ) );
  MUX U8186 ( .IN0(\u_a23_core/u_execute/u_register_bank/r1[4] ), .IN1(n6094), 
        .SEL(n6204), .F(\u_a23_core/u_execute/u_register_bank/n4559 ) );
  MUX U8187 ( .IN0(\u_a23_core/u_execute/u_register_bank/r1[3] ), .IN1(n6095), 
        .SEL(n6204), .F(\u_a23_core/u_execute/u_register_bank/n4557 ) );
  MUX U8188 ( .IN0(\u_a23_core/u_execute/u_register_bank/r1[2] ), .IN1(n6096), 
        .SEL(n6204), .F(\u_a23_core/u_execute/u_register_bank/n4555 ) );
  MUX U8189 ( .IN0(\u_a23_core/u_execute/u_register_bank/r1[1] ), .IN1(n6097), 
        .SEL(n6204), .F(\u_a23_core/u_execute/u_register_bank/n4553 ) );
  MUX U8190 ( .IN0(\u_a23_core/u_execute/u_register_bank/r1[0] ), .IN1(n6098), 
        .SEL(n6204), .F(\u_a23_core/u_execute/u_register_bank/n4551 ) );
  ANDN U8191 ( .A(\u_a23_core/reg_bank_wen[1] ), .B(n6099), .Z(n6204) );
  MUX U8192 ( .IN0(\u_a23_core/u_execute/u_register_bank/r2[31] ), .IN1(n6066), 
        .SEL(n6205), .F(\u_a23_core/u_execute/u_register_bank/n4549 ) );
  MUX U8193 ( .IN0(\u_a23_core/u_execute/u_register_bank/r2[30] ), .IN1(n6068), 
        .SEL(n6205), .F(\u_a23_core/u_execute/u_register_bank/n4547 ) );
  MUX U8194 ( .IN0(\u_a23_core/u_execute/u_register_bank/r2[29] ), .IN1(n6069), 
        .SEL(n6205), .F(\u_a23_core/u_execute/u_register_bank/n4545 ) );
  MUX U8195 ( .IN0(\u_a23_core/u_execute/u_register_bank/r2[28] ), .IN1(n6070), 
        .SEL(n6205), .F(\u_a23_core/u_execute/u_register_bank/n4543 ) );
  MUX U8196 ( .IN0(\u_a23_core/u_execute/u_register_bank/r2[27] ), .IN1(n6071), 
        .SEL(n6205), .F(\u_a23_core/u_execute/u_register_bank/n4541 ) );
  MUX U8197 ( .IN0(\u_a23_core/u_execute/u_register_bank/r2[26] ), .IN1(n6072), 
        .SEL(n6205), .F(\u_a23_core/u_execute/u_register_bank/n4539 ) );
  MUX U8198 ( .IN0(\u_a23_core/u_execute/u_register_bank/r2[25] ), .IN1(n6073), 
        .SEL(n6205), .F(\u_a23_core/u_execute/u_register_bank/n4537 ) );
  MUX U8199 ( .IN0(\u_a23_core/u_execute/u_register_bank/r2[24] ), .IN1(n6074), 
        .SEL(n6205), .F(\u_a23_core/u_execute/u_register_bank/n4535 ) );
  MUX U8200 ( .IN0(\u_a23_core/u_execute/u_register_bank/r2[23] ), .IN1(n6075), 
        .SEL(n6205), .F(\u_a23_core/u_execute/u_register_bank/n4533 ) );
  MUX U8201 ( .IN0(\u_a23_core/u_execute/u_register_bank/r2[22] ), .IN1(n6076), 
        .SEL(n6205), .F(\u_a23_core/u_execute/u_register_bank/n4531 ) );
  MUX U8202 ( .IN0(\u_a23_core/u_execute/u_register_bank/r2[21] ), .IN1(n6077), 
        .SEL(n6205), .F(\u_a23_core/u_execute/u_register_bank/n4529 ) );
  MUX U8203 ( .IN0(\u_a23_core/u_execute/u_register_bank/r2[20] ), .IN1(n6078), 
        .SEL(n6205), .F(\u_a23_core/u_execute/u_register_bank/n4527 ) );
  MUX U8204 ( .IN0(\u_a23_core/u_execute/u_register_bank/r2[19] ), .IN1(n6079), 
        .SEL(n6205), .F(\u_a23_core/u_execute/u_register_bank/n4525 ) );
  MUX U8205 ( .IN0(\u_a23_core/u_execute/u_register_bank/r2[18] ), .IN1(n6080), 
        .SEL(n6205), .F(\u_a23_core/u_execute/u_register_bank/n4523 ) );
  MUX U8206 ( .IN0(\u_a23_core/u_execute/u_register_bank/r2[17] ), .IN1(n6081), 
        .SEL(n6205), .F(\u_a23_core/u_execute/u_register_bank/n4521 ) );
  MUX U8207 ( .IN0(\u_a23_core/u_execute/u_register_bank/r2[16] ), .IN1(n6082), 
        .SEL(n6205), .F(\u_a23_core/u_execute/u_register_bank/n4519 ) );
  MUX U8208 ( .IN0(\u_a23_core/u_execute/u_register_bank/r2[15] ), .IN1(n6083), 
        .SEL(n6205), .F(\u_a23_core/u_execute/u_register_bank/n4517 ) );
  MUX U8209 ( .IN0(\u_a23_core/u_execute/u_register_bank/r2[14] ), .IN1(n6084), 
        .SEL(n6205), .F(\u_a23_core/u_execute/u_register_bank/n4515 ) );
  MUX U8210 ( .IN0(\u_a23_core/u_execute/u_register_bank/r2[13] ), .IN1(n6085), 
        .SEL(n6205), .F(\u_a23_core/u_execute/u_register_bank/n4513 ) );
  MUX U8211 ( .IN0(\u_a23_core/u_execute/u_register_bank/r2[12] ), .IN1(n6086), 
        .SEL(n6205), .F(\u_a23_core/u_execute/u_register_bank/n4511 ) );
  MUX U8212 ( .IN0(\u_a23_core/u_execute/u_register_bank/r2[11] ), .IN1(n6087), 
        .SEL(n6205), .F(\u_a23_core/u_execute/u_register_bank/n4509 ) );
  MUX U8213 ( .IN0(\u_a23_core/u_execute/u_register_bank/r2[10] ), .IN1(n6088), 
        .SEL(n6205), .F(\u_a23_core/u_execute/u_register_bank/n4507 ) );
  MUX U8214 ( .IN0(\u_a23_core/u_execute/u_register_bank/r2[9] ), .IN1(n6089), 
        .SEL(n6205), .F(\u_a23_core/u_execute/u_register_bank/n4505 ) );
  MUX U8215 ( .IN0(\u_a23_core/u_execute/u_register_bank/r2[8] ), .IN1(n6090), 
        .SEL(n6205), .F(\u_a23_core/u_execute/u_register_bank/n4503 ) );
  MUX U8216 ( .IN0(\u_a23_core/u_execute/u_register_bank/r2[7] ), .IN1(n6091), 
        .SEL(n6205), .F(\u_a23_core/u_execute/u_register_bank/n4501 ) );
  MUX U8217 ( .IN0(\u_a23_core/u_execute/u_register_bank/r2[6] ), .IN1(n6092), 
        .SEL(n6205), .F(\u_a23_core/u_execute/u_register_bank/n4499 ) );
  MUX U8218 ( .IN0(\u_a23_core/u_execute/u_register_bank/r2[5] ), .IN1(n6093), 
        .SEL(n6205), .F(\u_a23_core/u_execute/u_register_bank/n4497 ) );
  MUX U8219 ( .IN0(\u_a23_core/u_execute/u_register_bank/r2[4] ), .IN1(n6094), 
        .SEL(n6205), .F(\u_a23_core/u_execute/u_register_bank/n4495 ) );
  MUX U8220 ( .IN0(\u_a23_core/u_execute/u_register_bank/r2[3] ), .IN1(n6095), 
        .SEL(n6205), .F(\u_a23_core/u_execute/u_register_bank/n4493 ) );
  MUX U8221 ( .IN0(\u_a23_core/u_execute/u_register_bank/r2[2] ), .IN1(n6096), 
        .SEL(n6205), .F(\u_a23_core/u_execute/u_register_bank/n4491 ) );
  MUX U8222 ( .IN0(\u_a23_core/u_execute/u_register_bank/r2[1] ), .IN1(n6097), 
        .SEL(n6205), .F(\u_a23_core/u_execute/u_register_bank/n4489 ) );
  MUX U8223 ( .IN0(\u_a23_core/u_execute/u_register_bank/r2[0] ), .IN1(n6098), 
        .SEL(n6205), .F(\u_a23_core/u_execute/u_register_bank/n4487 ) );
  ANDN U8224 ( .A(\u_a23_core/reg_bank_wen[2] ), .B(n6099), .Z(n6205) );
  MUX U8225 ( .IN0(\u_a23_core/u_execute/u_register_bank/r3[31] ), .IN1(n6066), 
        .SEL(n6206), .F(\u_a23_core/u_execute/u_register_bank/n4485 ) );
  MUX U8226 ( .IN0(\u_a23_core/u_execute/u_register_bank/r3[30] ), .IN1(n6068), 
        .SEL(n6206), .F(\u_a23_core/u_execute/u_register_bank/n4483 ) );
  MUX U8227 ( .IN0(\u_a23_core/u_execute/u_register_bank/r3[29] ), .IN1(n6069), 
        .SEL(n6206), .F(\u_a23_core/u_execute/u_register_bank/n4481 ) );
  MUX U8228 ( .IN0(\u_a23_core/u_execute/u_register_bank/r3[28] ), .IN1(n6070), 
        .SEL(n6206), .F(\u_a23_core/u_execute/u_register_bank/n4479 ) );
  MUX U8229 ( .IN0(\u_a23_core/u_execute/u_register_bank/r3[27] ), .IN1(n6071), 
        .SEL(n6206), .F(\u_a23_core/u_execute/u_register_bank/n4477 ) );
  MUX U8230 ( .IN0(\u_a23_core/u_execute/u_register_bank/r3[26] ), .IN1(n6072), 
        .SEL(n6206), .F(\u_a23_core/u_execute/u_register_bank/n4475 ) );
  MUX U8231 ( .IN0(\u_a23_core/u_execute/u_register_bank/r3[25] ), .IN1(n6073), 
        .SEL(n6206), .F(\u_a23_core/u_execute/u_register_bank/n4473 ) );
  MUX U8232 ( .IN0(\u_a23_core/u_execute/u_register_bank/r3[24] ), .IN1(n6074), 
        .SEL(n6206), .F(\u_a23_core/u_execute/u_register_bank/n4471 ) );
  MUX U8233 ( .IN0(\u_a23_core/u_execute/u_register_bank/r3[23] ), .IN1(n6075), 
        .SEL(n6206), .F(\u_a23_core/u_execute/u_register_bank/n4469 ) );
  MUX U8234 ( .IN0(\u_a23_core/u_execute/u_register_bank/r3[22] ), .IN1(n6076), 
        .SEL(n6206), .F(\u_a23_core/u_execute/u_register_bank/n4467 ) );
  MUX U8235 ( .IN0(\u_a23_core/u_execute/u_register_bank/r3[21] ), .IN1(n6077), 
        .SEL(n6206), .F(\u_a23_core/u_execute/u_register_bank/n4465 ) );
  MUX U8236 ( .IN0(\u_a23_core/u_execute/u_register_bank/r3[20] ), .IN1(n6078), 
        .SEL(n6206), .F(\u_a23_core/u_execute/u_register_bank/n4463 ) );
  MUX U8237 ( .IN0(\u_a23_core/u_execute/u_register_bank/r3[19] ), .IN1(n6079), 
        .SEL(n6206), .F(\u_a23_core/u_execute/u_register_bank/n4461 ) );
  MUX U8238 ( .IN0(\u_a23_core/u_execute/u_register_bank/r3[18] ), .IN1(n6080), 
        .SEL(n6206), .F(\u_a23_core/u_execute/u_register_bank/n4459 ) );
  MUX U8239 ( .IN0(\u_a23_core/u_execute/u_register_bank/r3[17] ), .IN1(n6081), 
        .SEL(n6206), .F(\u_a23_core/u_execute/u_register_bank/n4457 ) );
  MUX U8240 ( .IN0(\u_a23_core/u_execute/u_register_bank/r3[16] ), .IN1(n6082), 
        .SEL(n6206), .F(\u_a23_core/u_execute/u_register_bank/n4455 ) );
  MUX U8241 ( .IN0(\u_a23_core/u_execute/u_register_bank/r3[15] ), .IN1(n6083), 
        .SEL(n6206), .F(\u_a23_core/u_execute/u_register_bank/n4453 ) );
  MUX U8242 ( .IN0(\u_a23_core/u_execute/u_register_bank/r3[14] ), .IN1(n6084), 
        .SEL(n6206), .F(\u_a23_core/u_execute/u_register_bank/n4451 ) );
  MUX U8243 ( .IN0(\u_a23_core/u_execute/u_register_bank/r3[13] ), .IN1(n6085), 
        .SEL(n6206), .F(\u_a23_core/u_execute/u_register_bank/n4449 ) );
  MUX U8244 ( .IN0(\u_a23_core/u_execute/u_register_bank/r3[12] ), .IN1(n6086), 
        .SEL(n6206), .F(\u_a23_core/u_execute/u_register_bank/n4447 ) );
  MUX U8245 ( .IN0(\u_a23_core/u_execute/u_register_bank/r3[11] ), .IN1(n6087), 
        .SEL(n6206), .F(\u_a23_core/u_execute/u_register_bank/n4445 ) );
  MUX U8246 ( .IN0(\u_a23_core/u_execute/u_register_bank/r3[10] ), .IN1(n6088), 
        .SEL(n6206), .F(\u_a23_core/u_execute/u_register_bank/n4443 ) );
  MUX U8247 ( .IN0(\u_a23_core/u_execute/u_register_bank/r3[9] ), .IN1(n6089), 
        .SEL(n6206), .F(\u_a23_core/u_execute/u_register_bank/n4441 ) );
  MUX U8248 ( .IN0(\u_a23_core/u_execute/u_register_bank/r3[8] ), .IN1(n6090), 
        .SEL(n6206), .F(\u_a23_core/u_execute/u_register_bank/n4439 ) );
  MUX U8249 ( .IN0(\u_a23_core/u_execute/u_register_bank/r3[7] ), .IN1(n6091), 
        .SEL(n6206), .F(\u_a23_core/u_execute/u_register_bank/n4437 ) );
  MUX U8250 ( .IN0(\u_a23_core/u_execute/u_register_bank/r3[6] ), .IN1(n6092), 
        .SEL(n6206), .F(\u_a23_core/u_execute/u_register_bank/n4435 ) );
  MUX U8251 ( .IN0(\u_a23_core/u_execute/u_register_bank/r3[5] ), .IN1(n6093), 
        .SEL(n6206), .F(\u_a23_core/u_execute/u_register_bank/n4433 ) );
  MUX U8252 ( .IN0(\u_a23_core/u_execute/u_register_bank/r3[4] ), .IN1(n6094), 
        .SEL(n6206), .F(\u_a23_core/u_execute/u_register_bank/n4431 ) );
  MUX U8253 ( .IN0(\u_a23_core/u_execute/u_register_bank/r3[3] ), .IN1(n6095), 
        .SEL(n6206), .F(\u_a23_core/u_execute/u_register_bank/n4429 ) );
  MUX U8254 ( .IN0(\u_a23_core/u_execute/u_register_bank/r3[2] ), .IN1(n6096), 
        .SEL(n6206), .F(\u_a23_core/u_execute/u_register_bank/n4427 ) );
  MUX U8255 ( .IN0(\u_a23_core/u_execute/u_register_bank/r3[1] ), .IN1(n6097), 
        .SEL(n6206), .F(\u_a23_core/u_execute/u_register_bank/n4425 ) );
  MUX U8256 ( .IN0(\u_a23_core/u_execute/u_register_bank/r3[0] ), .IN1(n6098), 
        .SEL(n6206), .F(\u_a23_core/u_execute/u_register_bank/n4423 ) );
  ANDN U8257 ( .A(\u_a23_core/reg_bank_wen[3] ), .B(n6099), .Z(n6206) );
  MUX U8258 ( .IN0(\u_a23_core/u_execute/u_register_bank/r4[31] ), .IN1(n6066), 
        .SEL(n6207), .F(\u_a23_core/u_execute/u_register_bank/n4421 ) );
  MUX U8259 ( .IN0(\u_a23_core/u_execute/u_register_bank/r4[30] ), .IN1(n6068), 
        .SEL(n6207), .F(\u_a23_core/u_execute/u_register_bank/n4419 ) );
  MUX U8260 ( .IN0(\u_a23_core/u_execute/u_register_bank/r4[29] ), .IN1(n6069), 
        .SEL(n6207), .F(\u_a23_core/u_execute/u_register_bank/n4417 ) );
  MUX U8261 ( .IN0(\u_a23_core/u_execute/u_register_bank/r4[28] ), .IN1(n6070), 
        .SEL(n6207), .F(\u_a23_core/u_execute/u_register_bank/n4415 ) );
  MUX U8262 ( .IN0(\u_a23_core/u_execute/u_register_bank/r4[27] ), .IN1(n6071), 
        .SEL(n6207), .F(\u_a23_core/u_execute/u_register_bank/n4413 ) );
  MUX U8263 ( .IN0(\u_a23_core/u_execute/u_register_bank/r4[26] ), .IN1(n6072), 
        .SEL(n6207), .F(\u_a23_core/u_execute/u_register_bank/n4411 ) );
  MUX U8264 ( .IN0(\u_a23_core/u_execute/u_register_bank/r4[25] ), .IN1(n6073), 
        .SEL(n6207), .F(\u_a23_core/u_execute/u_register_bank/n4409 ) );
  MUX U8265 ( .IN0(\u_a23_core/u_execute/u_register_bank/r4[24] ), .IN1(n6074), 
        .SEL(n6207), .F(\u_a23_core/u_execute/u_register_bank/n4407 ) );
  MUX U8266 ( .IN0(\u_a23_core/u_execute/u_register_bank/r4[23] ), .IN1(n6075), 
        .SEL(n6207), .F(\u_a23_core/u_execute/u_register_bank/n4405 ) );
  MUX U8267 ( .IN0(\u_a23_core/u_execute/u_register_bank/r4[22] ), .IN1(n6076), 
        .SEL(n6207), .F(\u_a23_core/u_execute/u_register_bank/n4403 ) );
  MUX U8268 ( .IN0(\u_a23_core/u_execute/u_register_bank/r4[21] ), .IN1(n6077), 
        .SEL(n6207), .F(\u_a23_core/u_execute/u_register_bank/n4401 ) );
  MUX U8269 ( .IN0(\u_a23_core/u_execute/u_register_bank/r4[20] ), .IN1(n6078), 
        .SEL(n6207), .F(\u_a23_core/u_execute/u_register_bank/n4399 ) );
  MUX U8270 ( .IN0(\u_a23_core/u_execute/u_register_bank/r4[19] ), .IN1(n6079), 
        .SEL(n6207), .F(\u_a23_core/u_execute/u_register_bank/n4397 ) );
  MUX U8271 ( .IN0(\u_a23_core/u_execute/u_register_bank/r4[18] ), .IN1(n6080), 
        .SEL(n6207), .F(\u_a23_core/u_execute/u_register_bank/n4395 ) );
  MUX U8272 ( .IN0(\u_a23_core/u_execute/u_register_bank/r4[17] ), .IN1(n6081), 
        .SEL(n6207), .F(\u_a23_core/u_execute/u_register_bank/n4393 ) );
  MUX U8273 ( .IN0(\u_a23_core/u_execute/u_register_bank/r4[16] ), .IN1(n6082), 
        .SEL(n6207), .F(\u_a23_core/u_execute/u_register_bank/n4391 ) );
  MUX U8274 ( .IN0(\u_a23_core/u_execute/u_register_bank/r4[15] ), .IN1(n6083), 
        .SEL(n6207), .F(\u_a23_core/u_execute/u_register_bank/n4389 ) );
  MUX U8275 ( .IN0(\u_a23_core/u_execute/u_register_bank/r4[14] ), .IN1(n6084), 
        .SEL(n6207), .F(\u_a23_core/u_execute/u_register_bank/n4387 ) );
  MUX U8276 ( .IN0(\u_a23_core/u_execute/u_register_bank/r4[13] ), .IN1(n6085), 
        .SEL(n6207), .F(\u_a23_core/u_execute/u_register_bank/n4385 ) );
  MUX U8277 ( .IN0(\u_a23_core/u_execute/u_register_bank/r4[12] ), .IN1(n6086), 
        .SEL(n6207), .F(\u_a23_core/u_execute/u_register_bank/n4383 ) );
  MUX U8278 ( .IN0(\u_a23_core/u_execute/u_register_bank/r4[11] ), .IN1(n6087), 
        .SEL(n6207), .F(\u_a23_core/u_execute/u_register_bank/n4381 ) );
  MUX U8279 ( .IN0(\u_a23_core/u_execute/u_register_bank/r4[10] ), .IN1(n6088), 
        .SEL(n6207), .F(\u_a23_core/u_execute/u_register_bank/n4379 ) );
  MUX U8280 ( .IN0(\u_a23_core/u_execute/u_register_bank/r4[9] ), .IN1(n6089), 
        .SEL(n6207), .F(\u_a23_core/u_execute/u_register_bank/n4377 ) );
  MUX U8281 ( .IN0(\u_a23_core/u_execute/u_register_bank/r4[8] ), .IN1(n6090), 
        .SEL(n6207), .F(\u_a23_core/u_execute/u_register_bank/n4375 ) );
  MUX U8282 ( .IN0(\u_a23_core/u_execute/u_register_bank/r4[7] ), .IN1(n6091), 
        .SEL(n6207), .F(\u_a23_core/u_execute/u_register_bank/n4373 ) );
  MUX U8283 ( .IN0(\u_a23_core/u_execute/u_register_bank/r4[6] ), .IN1(n6092), 
        .SEL(n6207), .F(\u_a23_core/u_execute/u_register_bank/n4371 ) );
  MUX U8284 ( .IN0(\u_a23_core/u_execute/u_register_bank/r4[5] ), .IN1(n6093), 
        .SEL(n6207), .F(\u_a23_core/u_execute/u_register_bank/n4369 ) );
  MUX U8285 ( .IN0(\u_a23_core/u_execute/u_register_bank/r4[4] ), .IN1(n6094), 
        .SEL(n6207), .F(\u_a23_core/u_execute/u_register_bank/n4367 ) );
  MUX U8286 ( .IN0(\u_a23_core/u_execute/u_register_bank/r4[3] ), .IN1(n6095), 
        .SEL(n6207), .F(\u_a23_core/u_execute/u_register_bank/n4365 ) );
  MUX U8287 ( .IN0(\u_a23_core/u_execute/u_register_bank/r4[2] ), .IN1(n6096), 
        .SEL(n6207), .F(\u_a23_core/u_execute/u_register_bank/n4363 ) );
  MUX U8288 ( .IN0(\u_a23_core/u_execute/u_register_bank/r4[1] ), .IN1(n6097), 
        .SEL(n6207), .F(\u_a23_core/u_execute/u_register_bank/n4361 ) );
  MUX U8289 ( .IN0(\u_a23_core/u_execute/u_register_bank/r4[0] ), .IN1(n6098), 
        .SEL(n6207), .F(\u_a23_core/u_execute/u_register_bank/n4359 ) );
  ANDN U8290 ( .A(\u_a23_core/reg_bank_wen[4] ), .B(n6099), .Z(n6207) );
  MUX U8291 ( .IN0(\u_a23_core/u_execute/u_register_bank/r5[31] ), .IN1(n6066), 
        .SEL(n6208), .F(\u_a23_core/u_execute/u_register_bank/n4357 ) );
  MUX U8292 ( .IN0(\u_a23_core/u_execute/u_register_bank/r5[30] ), .IN1(n6068), 
        .SEL(n6208), .F(\u_a23_core/u_execute/u_register_bank/n4355 ) );
  MUX U8293 ( .IN0(\u_a23_core/u_execute/u_register_bank/r5[29] ), .IN1(n6069), 
        .SEL(n6208), .F(\u_a23_core/u_execute/u_register_bank/n4353 ) );
  MUX U8294 ( .IN0(\u_a23_core/u_execute/u_register_bank/r5[28] ), .IN1(n6070), 
        .SEL(n6208), .F(\u_a23_core/u_execute/u_register_bank/n4351 ) );
  MUX U8295 ( .IN0(\u_a23_core/u_execute/u_register_bank/r5[27] ), .IN1(n6071), 
        .SEL(n6208), .F(\u_a23_core/u_execute/u_register_bank/n4349 ) );
  MUX U8296 ( .IN0(\u_a23_core/u_execute/u_register_bank/r5[26] ), .IN1(n6072), 
        .SEL(n6208), .F(\u_a23_core/u_execute/u_register_bank/n4347 ) );
  MUX U8297 ( .IN0(\u_a23_core/u_execute/u_register_bank/r5[25] ), .IN1(n6073), 
        .SEL(n6208), .F(\u_a23_core/u_execute/u_register_bank/n4345 ) );
  MUX U8298 ( .IN0(\u_a23_core/u_execute/u_register_bank/r5[24] ), .IN1(n6074), 
        .SEL(n6208), .F(\u_a23_core/u_execute/u_register_bank/n4343 ) );
  MUX U8299 ( .IN0(\u_a23_core/u_execute/u_register_bank/r5[23] ), .IN1(n6075), 
        .SEL(n6208), .F(\u_a23_core/u_execute/u_register_bank/n4341 ) );
  MUX U8300 ( .IN0(\u_a23_core/u_execute/u_register_bank/r5[22] ), .IN1(n6076), 
        .SEL(n6208), .F(\u_a23_core/u_execute/u_register_bank/n4339 ) );
  MUX U8301 ( .IN0(\u_a23_core/u_execute/u_register_bank/r5[21] ), .IN1(n6077), 
        .SEL(n6208), .F(\u_a23_core/u_execute/u_register_bank/n4337 ) );
  MUX U8302 ( .IN0(\u_a23_core/u_execute/u_register_bank/r5[20] ), .IN1(n6078), 
        .SEL(n6208), .F(\u_a23_core/u_execute/u_register_bank/n4335 ) );
  MUX U8303 ( .IN0(\u_a23_core/u_execute/u_register_bank/r5[19] ), .IN1(n6079), 
        .SEL(n6208), .F(\u_a23_core/u_execute/u_register_bank/n4333 ) );
  MUX U8304 ( .IN0(\u_a23_core/u_execute/u_register_bank/r5[18] ), .IN1(n6080), 
        .SEL(n6208), .F(\u_a23_core/u_execute/u_register_bank/n4331 ) );
  MUX U8305 ( .IN0(\u_a23_core/u_execute/u_register_bank/r5[17] ), .IN1(n6081), 
        .SEL(n6208), .F(\u_a23_core/u_execute/u_register_bank/n4329 ) );
  MUX U8306 ( .IN0(\u_a23_core/u_execute/u_register_bank/r5[16] ), .IN1(n6082), 
        .SEL(n6208), .F(\u_a23_core/u_execute/u_register_bank/n4327 ) );
  MUX U8307 ( .IN0(\u_a23_core/u_execute/u_register_bank/r5[15] ), .IN1(n6083), 
        .SEL(n6208), .F(\u_a23_core/u_execute/u_register_bank/n4325 ) );
  MUX U8308 ( .IN0(\u_a23_core/u_execute/u_register_bank/r5[14] ), .IN1(n6084), 
        .SEL(n6208), .F(\u_a23_core/u_execute/u_register_bank/n4323 ) );
  MUX U8309 ( .IN0(\u_a23_core/u_execute/u_register_bank/r5[13] ), .IN1(n6085), 
        .SEL(n6208), .F(\u_a23_core/u_execute/u_register_bank/n4321 ) );
  MUX U8310 ( .IN0(\u_a23_core/u_execute/u_register_bank/r5[12] ), .IN1(n6086), 
        .SEL(n6208), .F(\u_a23_core/u_execute/u_register_bank/n4319 ) );
  MUX U8311 ( .IN0(\u_a23_core/u_execute/u_register_bank/r5[11] ), .IN1(n6087), 
        .SEL(n6208), .F(\u_a23_core/u_execute/u_register_bank/n4317 ) );
  MUX U8312 ( .IN0(\u_a23_core/u_execute/u_register_bank/r5[10] ), .IN1(n6088), 
        .SEL(n6208), .F(\u_a23_core/u_execute/u_register_bank/n4315 ) );
  MUX U8313 ( .IN0(\u_a23_core/u_execute/u_register_bank/r5[9] ), .IN1(n6089), 
        .SEL(n6208), .F(\u_a23_core/u_execute/u_register_bank/n4313 ) );
  MUX U8314 ( .IN0(\u_a23_core/u_execute/u_register_bank/r5[8] ), .IN1(n6090), 
        .SEL(n6208), .F(\u_a23_core/u_execute/u_register_bank/n4311 ) );
  MUX U8315 ( .IN0(\u_a23_core/u_execute/u_register_bank/r5[7] ), .IN1(n6091), 
        .SEL(n6208), .F(\u_a23_core/u_execute/u_register_bank/n4309 ) );
  MUX U8316 ( .IN0(\u_a23_core/u_execute/u_register_bank/r5[6] ), .IN1(n6092), 
        .SEL(n6208), .F(\u_a23_core/u_execute/u_register_bank/n4307 ) );
  MUX U8317 ( .IN0(\u_a23_core/u_execute/u_register_bank/r5[5] ), .IN1(n6093), 
        .SEL(n6208), .F(\u_a23_core/u_execute/u_register_bank/n4305 ) );
  MUX U8318 ( .IN0(\u_a23_core/u_execute/u_register_bank/r5[4] ), .IN1(n6094), 
        .SEL(n6208), .F(\u_a23_core/u_execute/u_register_bank/n4303 ) );
  MUX U8319 ( .IN0(\u_a23_core/u_execute/u_register_bank/r5[3] ), .IN1(n6095), 
        .SEL(n6208), .F(\u_a23_core/u_execute/u_register_bank/n4301 ) );
  MUX U8320 ( .IN0(\u_a23_core/u_execute/u_register_bank/r5[2] ), .IN1(n6096), 
        .SEL(n6208), .F(\u_a23_core/u_execute/u_register_bank/n4299 ) );
  MUX U8321 ( .IN0(\u_a23_core/u_execute/u_register_bank/r5[1] ), .IN1(n6097), 
        .SEL(n6208), .F(\u_a23_core/u_execute/u_register_bank/n4297 ) );
  MUX U8322 ( .IN0(\u_a23_core/u_execute/u_register_bank/r5[0] ), .IN1(n6098), 
        .SEL(n6208), .F(\u_a23_core/u_execute/u_register_bank/n4295 ) );
  ANDN U8323 ( .A(\u_a23_core/reg_bank_wen[5] ), .B(n6099), .Z(n6208) );
  MUX U8324 ( .IN0(\u_a23_core/u_execute/u_register_bank/r6[31] ), .IN1(n6066), 
        .SEL(n6209), .F(\u_a23_core/u_execute/u_register_bank/n4293 ) );
  MUX U8325 ( .IN0(\u_a23_core/u_execute/u_register_bank/r6[30] ), .IN1(n6068), 
        .SEL(n6209), .F(\u_a23_core/u_execute/u_register_bank/n4291 ) );
  MUX U8326 ( .IN0(\u_a23_core/u_execute/u_register_bank/r6[29] ), .IN1(n6069), 
        .SEL(n6209), .F(\u_a23_core/u_execute/u_register_bank/n4289 ) );
  MUX U8327 ( .IN0(\u_a23_core/u_execute/u_register_bank/r6[28] ), .IN1(n6070), 
        .SEL(n6209), .F(\u_a23_core/u_execute/u_register_bank/n4287 ) );
  MUX U8328 ( .IN0(\u_a23_core/u_execute/u_register_bank/r6[27] ), .IN1(n6071), 
        .SEL(n6209), .F(\u_a23_core/u_execute/u_register_bank/n4285 ) );
  MUX U8329 ( .IN0(\u_a23_core/u_execute/u_register_bank/r6[26] ), .IN1(n6072), 
        .SEL(n6209), .F(\u_a23_core/u_execute/u_register_bank/n4283 ) );
  MUX U8330 ( .IN0(\u_a23_core/u_execute/u_register_bank/r6[25] ), .IN1(n6073), 
        .SEL(n6209), .F(\u_a23_core/u_execute/u_register_bank/n4281 ) );
  MUX U8331 ( .IN0(\u_a23_core/u_execute/u_register_bank/r6[24] ), .IN1(n6074), 
        .SEL(n6209), .F(\u_a23_core/u_execute/u_register_bank/n4279 ) );
  MUX U8332 ( .IN0(\u_a23_core/u_execute/u_register_bank/r6[23] ), .IN1(n6075), 
        .SEL(n6209), .F(\u_a23_core/u_execute/u_register_bank/n4277 ) );
  MUX U8333 ( .IN0(\u_a23_core/u_execute/u_register_bank/r6[22] ), .IN1(n6076), 
        .SEL(n6209), .F(\u_a23_core/u_execute/u_register_bank/n4275 ) );
  MUX U8334 ( .IN0(\u_a23_core/u_execute/u_register_bank/r6[21] ), .IN1(n6077), 
        .SEL(n6209), .F(\u_a23_core/u_execute/u_register_bank/n4273 ) );
  MUX U8335 ( .IN0(\u_a23_core/u_execute/u_register_bank/r6[20] ), .IN1(n6078), 
        .SEL(n6209), .F(\u_a23_core/u_execute/u_register_bank/n4271 ) );
  MUX U8336 ( .IN0(\u_a23_core/u_execute/u_register_bank/r6[19] ), .IN1(n6079), 
        .SEL(n6209), .F(\u_a23_core/u_execute/u_register_bank/n4269 ) );
  MUX U8337 ( .IN0(\u_a23_core/u_execute/u_register_bank/r6[18] ), .IN1(n6080), 
        .SEL(n6209), .F(\u_a23_core/u_execute/u_register_bank/n4267 ) );
  MUX U8338 ( .IN0(\u_a23_core/u_execute/u_register_bank/r6[17] ), .IN1(n6081), 
        .SEL(n6209), .F(\u_a23_core/u_execute/u_register_bank/n4265 ) );
  MUX U8339 ( .IN0(\u_a23_core/u_execute/u_register_bank/r6[16] ), .IN1(n6082), 
        .SEL(n6209), .F(\u_a23_core/u_execute/u_register_bank/n4263 ) );
  MUX U8340 ( .IN0(\u_a23_core/u_execute/u_register_bank/r6[15] ), .IN1(n6083), 
        .SEL(n6209), .F(\u_a23_core/u_execute/u_register_bank/n4261 ) );
  MUX U8341 ( .IN0(\u_a23_core/u_execute/u_register_bank/r6[14] ), .IN1(n6084), 
        .SEL(n6209), .F(\u_a23_core/u_execute/u_register_bank/n4259 ) );
  MUX U8342 ( .IN0(\u_a23_core/u_execute/u_register_bank/r6[13] ), .IN1(n6085), 
        .SEL(n6209), .F(\u_a23_core/u_execute/u_register_bank/n4257 ) );
  MUX U8343 ( .IN0(\u_a23_core/u_execute/u_register_bank/r6[12] ), .IN1(n6086), 
        .SEL(n6209), .F(\u_a23_core/u_execute/u_register_bank/n4255 ) );
  MUX U8344 ( .IN0(\u_a23_core/u_execute/u_register_bank/r6[11] ), .IN1(n6087), 
        .SEL(n6209), .F(\u_a23_core/u_execute/u_register_bank/n4253 ) );
  MUX U8345 ( .IN0(\u_a23_core/u_execute/u_register_bank/r6[10] ), .IN1(n6088), 
        .SEL(n6209), .F(\u_a23_core/u_execute/u_register_bank/n4251 ) );
  MUX U8346 ( .IN0(\u_a23_core/u_execute/u_register_bank/r6[9] ), .IN1(n6089), 
        .SEL(n6209), .F(\u_a23_core/u_execute/u_register_bank/n4249 ) );
  MUX U8347 ( .IN0(\u_a23_core/u_execute/u_register_bank/r6[8] ), .IN1(n6090), 
        .SEL(n6209), .F(\u_a23_core/u_execute/u_register_bank/n4247 ) );
  MUX U8348 ( .IN0(\u_a23_core/u_execute/u_register_bank/r6[7] ), .IN1(n6091), 
        .SEL(n6209), .F(\u_a23_core/u_execute/u_register_bank/n4245 ) );
  MUX U8349 ( .IN0(\u_a23_core/u_execute/u_register_bank/r6[6] ), .IN1(n6092), 
        .SEL(n6209), .F(\u_a23_core/u_execute/u_register_bank/n4243 ) );
  MUX U8350 ( .IN0(\u_a23_core/u_execute/u_register_bank/r6[5] ), .IN1(n6093), 
        .SEL(n6209), .F(\u_a23_core/u_execute/u_register_bank/n4241 ) );
  MUX U8351 ( .IN0(\u_a23_core/u_execute/u_register_bank/r6[4] ), .IN1(n6094), 
        .SEL(n6209), .F(\u_a23_core/u_execute/u_register_bank/n4239 ) );
  MUX U8352 ( .IN0(\u_a23_core/u_execute/u_register_bank/r6[3] ), .IN1(n6095), 
        .SEL(n6209), .F(\u_a23_core/u_execute/u_register_bank/n4237 ) );
  MUX U8353 ( .IN0(\u_a23_core/u_execute/u_register_bank/r6[2] ), .IN1(n6096), 
        .SEL(n6209), .F(\u_a23_core/u_execute/u_register_bank/n4235 ) );
  MUX U8354 ( .IN0(\u_a23_core/u_execute/u_register_bank/r6[1] ), .IN1(n6097), 
        .SEL(n6209), .F(\u_a23_core/u_execute/u_register_bank/n4233 ) );
  MUX U8355 ( .IN0(\u_a23_core/u_execute/u_register_bank/r6[0] ), .IN1(n6098), 
        .SEL(n6209), .F(\u_a23_core/u_execute/u_register_bank/n4231 ) );
  ANDN U8356 ( .A(\u_a23_core/reg_bank_wen[6] ), .B(n6099), .Z(n6209) );
  MUX U8357 ( .IN0(\u_a23_core/u_execute/u_register_bank/r7[31] ), .IN1(n6066), 
        .SEL(n6210), .F(\u_a23_core/u_execute/u_register_bank/n4229 ) );
  MUX U8358 ( .IN0(\u_a23_core/u_execute/u_register_bank/r7[30] ), .IN1(n6068), 
        .SEL(n6210), .F(\u_a23_core/u_execute/u_register_bank/n4227 ) );
  MUX U8359 ( .IN0(\u_a23_core/u_execute/u_register_bank/r7[29] ), .IN1(n6069), 
        .SEL(n6210), .F(\u_a23_core/u_execute/u_register_bank/n4225 ) );
  MUX U8360 ( .IN0(\u_a23_core/u_execute/u_register_bank/r7[28] ), .IN1(n6070), 
        .SEL(n6210), .F(\u_a23_core/u_execute/u_register_bank/n4223 ) );
  MUX U8361 ( .IN0(\u_a23_core/u_execute/u_register_bank/r7[27] ), .IN1(n6071), 
        .SEL(n6210), .F(\u_a23_core/u_execute/u_register_bank/n4221 ) );
  MUX U8362 ( .IN0(\u_a23_core/u_execute/u_register_bank/r7[26] ), .IN1(n6072), 
        .SEL(n6210), .F(\u_a23_core/u_execute/u_register_bank/n4219 ) );
  MUX U8363 ( .IN0(\u_a23_core/u_execute/u_register_bank/r7[25] ), .IN1(n6073), 
        .SEL(n6210), .F(\u_a23_core/u_execute/u_register_bank/n4217 ) );
  MUX U8364 ( .IN0(\u_a23_core/u_execute/u_register_bank/r7[24] ), .IN1(n6074), 
        .SEL(n6210), .F(\u_a23_core/u_execute/u_register_bank/n4215 ) );
  MUX U8365 ( .IN0(\u_a23_core/u_execute/u_register_bank/r7[23] ), .IN1(n6075), 
        .SEL(n6210), .F(\u_a23_core/u_execute/u_register_bank/n4213 ) );
  MUX U8366 ( .IN0(\u_a23_core/u_execute/u_register_bank/r7[22] ), .IN1(n6076), 
        .SEL(n6210), .F(\u_a23_core/u_execute/u_register_bank/n4211 ) );
  MUX U8367 ( .IN0(\u_a23_core/u_execute/u_register_bank/r7[21] ), .IN1(n6077), 
        .SEL(n6210), .F(\u_a23_core/u_execute/u_register_bank/n4209 ) );
  MUX U8368 ( .IN0(\u_a23_core/u_execute/u_register_bank/r7[20] ), .IN1(n6078), 
        .SEL(n6210), .F(\u_a23_core/u_execute/u_register_bank/n4207 ) );
  MUX U8369 ( .IN0(\u_a23_core/u_execute/u_register_bank/r7[19] ), .IN1(n6079), 
        .SEL(n6210), .F(\u_a23_core/u_execute/u_register_bank/n4205 ) );
  MUX U8370 ( .IN0(\u_a23_core/u_execute/u_register_bank/r7[18] ), .IN1(n6080), 
        .SEL(n6210), .F(\u_a23_core/u_execute/u_register_bank/n4203 ) );
  MUX U8371 ( .IN0(\u_a23_core/u_execute/u_register_bank/r7[17] ), .IN1(n6081), 
        .SEL(n6210), .F(\u_a23_core/u_execute/u_register_bank/n4201 ) );
  MUX U8372 ( .IN0(\u_a23_core/u_execute/u_register_bank/r7[16] ), .IN1(n6082), 
        .SEL(n6210), .F(\u_a23_core/u_execute/u_register_bank/n4199 ) );
  MUX U8373 ( .IN0(\u_a23_core/u_execute/u_register_bank/r7[15] ), .IN1(n6083), 
        .SEL(n6210), .F(\u_a23_core/u_execute/u_register_bank/n4197 ) );
  MUX U8374 ( .IN0(\u_a23_core/u_execute/u_register_bank/r7[14] ), .IN1(n6084), 
        .SEL(n6210), .F(\u_a23_core/u_execute/u_register_bank/n4195 ) );
  MUX U8375 ( .IN0(\u_a23_core/u_execute/u_register_bank/r7[13] ), .IN1(n6085), 
        .SEL(n6210), .F(\u_a23_core/u_execute/u_register_bank/n4193 ) );
  MUX U8376 ( .IN0(\u_a23_core/u_execute/u_register_bank/r7[12] ), .IN1(n6086), 
        .SEL(n6210), .F(\u_a23_core/u_execute/u_register_bank/n4191 ) );
  MUX U8377 ( .IN0(\u_a23_core/u_execute/u_register_bank/r7[11] ), .IN1(n6087), 
        .SEL(n6210), .F(\u_a23_core/u_execute/u_register_bank/n4189 ) );
  MUX U8378 ( .IN0(\u_a23_core/u_execute/u_register_bank/r7[10] ), .IN1(n6088), 
        .SEL(n6210), .F(\u_a23_core/u_execute/u_register_bank/n4187 ) );
  MUX U8379 ( .IN0(\u_a23_core/u_execute/u_register_bank/r7[9] ), .IN1(n6089), 
        .SEL(n6210), .F(\u_a23_core/u_execute/u_register_bank/n4185 ) );
  MUX U8380 ( .IN0(\u_a23_core/u_execute/u_register_bank/r7[8] ), .IN1(n6090), 
        .SEL(n6210), .F(\u_a23_core/u_execute/u_register_bank/n4183 ) );
  MUX U8381 ( .IN0(\u_a23_core/u_execute/u_register_bank/r7[7] ), .IN1(n6091), 
        .SEL(n6210), .F(\u_a23_core/u_execute/u_register_bank/n4181 ) );
  MUX U8382 ( .IN0(\u_a23_core/u_execute/u_register_bank/r7[6] ), .IN1(n6092), 
        .SEL(n6210), .F(\u_a23_core/u_execute/u_register_bank/n4179 ) );
  MUX U8383 ( .IN0(\u_a23_core/u_execute/u_register_bank/r7[5] ), .IN1(n6093), 
        .SEL(n6210), .F(\u_a23_core/u_execute/u_register_bank/n4177 ) );
  MUX U8384 ( .IN0(\u_a23_core/u_execute/u_register_bank/r7[4] ), .IN1(n6094), 
        .SEL(n6210), .F(\u_a23_core/u_execute/u_register_bank/n4175 ) );
  MUX U8385 ( .IN0(\u_a23_core/u_execute/u_register_bank/r7[3] ), .IN1(n6095), 
        .SEL(n6210), .F(\u_a23_core/u_execute/u_register_bank/n4173 ) );
  MUX U8386 ( .IN0(\u_a23_core/u_execute/u_register_bank/r7[2] ), .IN1(n6096), 
        .SEL(n6210), .F(\u_a23_core/u_execute/u_register_bank/n4171 ) );
  MUX U8387 ( .IN0(\u_a23_core/u_execute/u_register_bank/r7[1] ), .IN1(n6097), 
        .SEL(n6210), .F(\u_a23_core/u_execute/u_register_bank/n4169 ) );
  MUX U8388 ( .IN0(\u_a23_core/u_execute/u_register_bank/r7[0] ), .IN1(n6098), 
        .SEL(n6210), .F(\u_a23_core/u_execute/u_register_bank/n4167 ) );
  ANDN U8389 ( .A(\u_a23_core/reg_bank_wen[7] ), .B(n6099), .Z(n6210) );
  MUX U8390 ( .IN0(\u_a23_core/u_execute/u_register_bank/r8[31] ), .IN1(n6066), 
        .SEL(n6211), .F(\u_a23_core/u_execute/u_register_bank/n4165 ) );
  MUX U8391 ( .IN0(\u_a23_core/u_execute/u_register_bank/r8[30] ), .IN1(n6068), 
        .SEL(n6211), .F(\u_a23_core/u_execute/u_register_bank/n4163 ) );
  MUX U8392 ( .IN0(\u_a23_core/u_execute/u_register_bank/r8[29] ), .IN1(n6069), 
        .SEL(n6211), .F(\u_a23_core/u_execute/u_register_bank/n4161 ) );
  MUX U8393 ( .IN0(\u_a23_core/u_execute/u_register_bank/r8[28] ), .IN1(n6070), 
        .SEL(n6211), .F(\u_a23_core/u_execute/u_register_bank/n4159 ) );
  MUX U8394 ( .IN0(\u_a23_core/u_execute/u_register_bank/r8[27] ), .IN1(n6071), 
        .SEL(n6211), .F(\u_a23_core/u_execute/u_register_bank/n4157 ) );
  MUX U8395 ( .IN0(\u_a23_core/u_execute/u_register_bank/r8[26] ), .IN1(n6072), 
        .SEL(n6211), .F(\u_a23_core/u_execute/u_register_bank/n4155 ) );
  MUX U8396 ( .IN0(\u_a23_core/u_execute/u_register_bank/r8[25] ), .IN1(n6073), 
        .SEL(n6211), .F(\u_a23_core/u_execute/u_register_bank/n4153 ) );
  MUX U8397 ( .IN0(\u_a23_core/u_execute/u_register_bank/r8[24] ), .IN1(n6074), 
        .SEL(n6211), .F(\u_a23_core/u_execute/u_register_bank/n4151 ) );
  MUX U8398 ( .IN0(\u_a23_core/u_execute/u_register_bank/r8[23] ), .IN1(n6075), 
        .SEL(n6211), .F(\u_a23_core/u_execute/u_register_bank/n4149 ) );
  MUX U8399 ( .IN0(\u_a23_core/u_execute/u_register_bank/r8[22] ), .IN1(n6076), 
        .SEL(n6211), .F(\u_a23_core/u_execute/u_register_bank/n4147 ) );
  MUX U8400 ( .IN0(\u_a23_core/u_execute/u_register_bank/r8[21] ), .IN1(n6077), 
        .SEL(n6211), .F(\u_a23_core/u_execute/u_register_bank/n4145 ) );
  MUX U8401 ( .IN0(\u_a23_core/u_execute/u_register_bank/r8[20] ), .IN1(n6078), 
        .SEL(n6211), .F(\u_a23_core/u_execute/u_register_bank/n4143 ) );
  MUX U8402 ( .IN0(\u_a23_core/u_execute/u_register_bank/r8[19] ), .IN1(n6079), 
        .SEL(n6211), .F(\u_a23_core/u_execute/u_register_bank/n4141 ) );
  MUX U8403 ( .IN0(\u_a23_core/u_execute/u_register_bank/r8[18] ), .IN1(n6080), 
        .SEL(n6211), .F(\u_a23_core/u_execute/u_register_bank/n4139 ) );
  MUX U8404 ( .IN0(\u_a23_core/u_execute/u_register_bank/r8[17] ), .IN1(n6081), 
        .SEL(n6211), .F(\u_a23_core/u_execute/u_register_bank/n4137 ) );
  MUX U8405 ( .IN0(\u_a23_core/u_execute/u_register_bank/r8[16] ), .IN1(n6082), 
        .SEL(n6211), .F(\u_a23_core/u_execute/u_register_bank/n4135 ) );
  MUX U8406 ( .IN0(\u_a23_core/u_execute/u_register_bank/r8[15] ), .IN1(n6083), 
        .SEL(n6211), .F(\u_a23_core/u_execute/u_register_bank/n4133 ) );
  MUX U8407 ( .IN0(\u_a23_core/u_execute/u_register_bank/r8[14] ), .IN1(n6084), 
        .SEL(n6211), .F(\u_a23_core/u_execute/u_register_bank/n4131 ) );
  MUX U8408 ( .IN0(\u_a23_core/u_execute/u_register_bank/r8[13] ), .IN1(n6085), 
        .SEL(n6211), .F(\u_a23_core/u_execute/u_register_bank/n4129 ) );
  MUX U8409 ( .IN0(\u_a23_core/u_execute/u_register_bank/r8[12] ), .IN1(n6086), 
        .SEL(n6211), .F(\u_a23_core/u_execute/u_register_bank/n4127 ) );
  MUX U8410 ( .IN0(\u_a23_core/u_execute/u_register_bank/r8[11] ), .IN1(n6087), 
        .SEL(n6211), .F(\u_a23_core/u_execute/u_register_bank/n4125 ) );
  MUX U8411 ( .IN0(\u_a23_core/u_execute/u_register_bank/r8[10] ), .IN1(n6088), 
        .SEL(n6211), .F(\u_a23_core/u_execute/u_register_bank/n4123 ) );
  MUX U8412 ( .IN0(\u_a23_core/u_execute/u_register_bank/r8[9] ), .IN1(n6089), 
        .SEL(n6211), .F(\u_a23_core/u_execute/u_register_bank/n4121 ) );
  MUX U8413 ( .IN0(\u_a23_core/u_execute/u_register_bank/r8[8] ), .IN1(n6090), 
        .SEL(n6211), .F(\u_a23_core/u_execute/u_register_bank/n4119 ) );
  MUX U8414 ( .IN0(\u_a23_core/u_execute/u_register_bank/r8[7] ), .IN1(n6091), 
        .SEL(n6211), .F(\u_a23_core/u_execute/u_register_bank/n4117 ) );
  MUX U8415 ( .IN0(\u_a23_core/u_execute/u_register_bank/r8[6] ), .IN1(n6092), 
        .SEL(n6211), .F(\u_a23_core/u_execute/u_register_bank/n4115 ) );
  MUX U8416 ( .IN0(\u_a23_core/u_execute/u_register_bank/r8[5] ), .IN1(n6093), 
        .SEL(n6211), .F(\u_a23_core/u_execute/u_register_bank/n4113 ) );
  MUX U8417 ( .IN0(\u_a23_core/u_execute/u_register_bank/r8[4] ), .IN1(n6094), 
        .SEL(n6211), .F(\u_a23_core/u_execute/u_register_bank/n4111 ) );
  MUX U8418 ( .IN0(\u_a23_core/u_execute/u_register_bank/r8[3] ), .IN1(n6095), 
        .SEL(n6211), .F(\u_a23_core/u_execute/u_register_bank/n4109 ) );
  MUX U8419 ( .IN0(\u_a23_core/u_execute/u_register_bank/r8[2] ), .IN1(n6096), 
        .SEL(n6211), .F(\u_a23_core/u_execute/u_register_bank/n4107 ) );
  MUX U8420 ( .IN0(\u_a23_core/u_execute/u_register_bank/r8[1] ), .IN1(n6097), 
        .SEL(n6211), .F(\u_a23_core/u_execute/u_register_bank/n4105 ) );
  MUX U8421 ( .IN0(\u_a23_core/u_execute/u_register_bank/r8[0] ), .IN1(n6098), 
        .SEL(n6211), .F(\u_a23_core/u_execute/u_register_bank/n4103 ) );
  ANDN U8422 ( .A(\u_a23_core/reg_bank_wen[8] ), .B(n6099), .Z(n6211) );
  MUX U8423 ( .IN0(\u_a23_core/u_execute/u_register_bank/r9[31] ), .IN1(n6066), 
        .SEL(n6212), .F(\u_a23_core/u_execute/u_register_bank/n4101 ) );
  MUX U8424 ( .IN0(\u_a23_core/u_execute/u_register_bank/r9[30] ), .IN1(n6068), 
        .SEL(n6212), .F(\u_a23_core/u_execute/u_register_bank/n4099 ) );
  MUX U8425 ( .IN0(\u_a23_core/u_execute/u_register_bank/r9[29] ), .IN1(n6069), 
        .SEL(n6212), .F(\u_a23_core/u_execute/u_register_bank/n4097 ) );
  MUX U8426 ( .IN0(\u_a23_core/u_execute/u_register_bank/r9[28] ), .IN1(n6070), 
        .SEL(n6212), .F(\u_a23_core/u_execute/u_register_bank/n4095 ) );
  MUX U8427 ( .IN0(\u_a23_core/u_execute/u_register_bank/r9[27] ), .IN1(n6071), 
        .SEL(n6212), .F(\u_a23_core/u_execute/u_register_bank/n4093 ) );
  MUX U8428 ( .IN0(\u_a23_core/u_execute/u_register_bank/r9[26] ), .IN1(n6072), 
        .SEL(n6212), .F(\u_a23_core/u_execute/u_register_bank/n4091 ) );
  MUX U8429 ( .IN0(\u_a23_core/u_execute/u_register_bank/r9[25] ), .IN1(n6073), 
        .SEL(n6212), .F(\u_a23_core/u_execute/u_register_bank/n4089 ) );
  MUX U8430 ( .IN0(\u_a23_core/u_execute/u_register_bank/r9[24] ), .IN1(n6074), 
        .SEL(n6212), .F(\u_a23_core/u_execute/u_register_bank/n4087 ) );
  MUX U8431 ( .IN0(\u_a23_core/u_execute/u_register_bank/r9[23] ), .IN1(n6075), 
        .SEL(n6212), .F(\u_a23_core/u_execute/u_register_bank/n4085 ) );
  MUX U8432 ( .IN0(\u_a23_core/u_execute/u_register_bank/r9[22] ), .IN1(n6076), 
        .SEL(n6212), .F(\u_a23_core/u_execute/u_register_bank/n4083 ) );
  MUX U8433 ( .IN0(\u_a23_core/u_execute/u_register_bank/r9[21] ), .IN1(n6077), 
        .SEL(n6212), .F(\u_a23_core/u_execute/u_register_bank/n4081 ) );
  MUX U8434 ( .IN0(\u_a23_core/u_execute/u_register_bank/r9[20] ), .IN1(n6078), 
        .SEL(n6212), .F(\u_a23_core/u_execute/u_register_bank/n4079 ) );
  MUX U8435 ( .IN0(\u_a23_core/u_execute/u_register_bank/r9[19] ), .IN1(n6079), 
        .SEL(n6212), .F(\u_a23_core/u_execute/u_register_bank/n4077 ) );
  MUX U8436 ( .IN0(\u_a23_core/u_execute/u_register_bank/r9[18] ), .IN1(n6080), 
        .SEL(n6212), .F(\u_a23_core/u_execute/u_register_bank/n4075 ) );
  MUX U8437 ( .IN0(\u_a23_core/u_execute/u_register_bank/r9[17] ), .IN1(n6081), 
        .SEL(n6212), .F(\u_a23_core/u_execute/u_register_bank/n4073 ) );
  MUX U8438 ( .IN0(\u_a23_core/u_execute/u_register_bank/r9[16] ), .IN1(n6082), 
        .SEL(n6212), .F(\u_a23_core/u_execute/u_register_bank/n4071 ) );
  MUX U8439 ( .IN0(\u_a23_core/u_execute/u_register_bank/r9[15] ), .IN1(n6083), 
        .SEL(n6212), .F(\u_a23_core/u_execute/u_register_bank/n4069 ) );
  MUX U8440 ( .IN0(\u_a23_core/u_execute/u_register_bank/r9[14] ), .IN1(n6084), 
        .SEL(n6212), .F(\u_a23_core/u_execute/u_register_bank/n4067 ) );
  MUX U8441 ( .IN0(\u_a23_core/u_execute/u_register_bank/r9[13] ), .IN1(n6085), 
        .SEL(n6212), .F(\u_a23_core/u_execute/u_register_bank/n4065 ) );
  MUX U8442 ( .IN0(\u_a23_core/u_execute/u_register_bank/r9[12] ), .IN1(n6086), 
        .SEL(n6212), .F(\u_a23_core/u_execute/u_register_bank/n4063 ) );
  MUX U8443 ( .IN0(\u_a23_core/u_execute/u_register_bank/r9[11] ), .IN1(n6087), 
        .SEL(n6212), .F(\u_a23_core/u_execute/u_register_bank/n4061 ) );
  MUX U8444 ( .IN0(\u_a23_core/u_execute/u_register_bank/r9[10] ), .IN1(n6088), 
        .SEL(n6212), .F(\u_a23_core/u_execute/u_register_bank/n4059 ) );
  MUX U8445 ( .IN0(\u_a23_core/u_execute/u_register_bank/r9[9] ), .IN1(n6089), 
        .SEL(n6212), .F(\u_a23_core/u_execute/u_register_bank/n4057 ) );
  MUX U8446 ( .IN0(\u_a23_core/u_execute/u_register_bank/r9[8] ), .IN1(n6090), 
        .SEL(n6212), .F(\u_a23_core/u_execute/u_register_bank/n4055 ) );
  MUX U8447 ( .IN0(\u_a23_core/u_execute/u_register_bank/r9[7] ), .IN1(n6091), 
        .SEL(n6212), .F(\u_a23_core/u_execute/u_register_bank/n4053 ) );
  MUX U8448 ( .IN0(\u_a23_core/u_execute/u_register_bank/r9[6] ), .IN1(n6092), 
        .SEL(n6212), .F(\u_a23_core/u_execute/u_register_bank/n4051 ) );
  MUX U8449 ( .IN0(\u_a23_core/u_execute/u_register_bank/r9[5] ), .IN1(n6093), 
        .SEL(n6212), .F(\u_a23_core/u_execute/u_register_bank/n4049 ) );
  MUX U8450 ( .IN0(\u_a23_core/u_execute/u_register_bank/r9[4] ), .IN1(n6094), 
        .SEL(n6212), .F(\u_a23_core/u_execute/u_register_bank/n4047 ) );
  MUX U8451 ( .IN0(\u_a23_core/u_execute/u_register_bank/r9[3] ), .IN1(n6095), 
        .SEL(n6212), .F(\u_a23_core/u_execute/u_register_bank/n4045 ) );
  MUX U8452 ( .IN0(\u_a23_core/u_execute/u_register_bank/r9[2] ), .IN1(n6096), 
        .SEL(n6212), .F(\u_a23_core/u_execute/u_register_bank/n4043 ) );
  MUX U8453 ( .IN0(\u_a23_core/u_execute/u_register_bank/r9[1] ), .IN1(n6097), 
        .SEL(n6212), .F(\u_a23_core/u_execute/u_register_bank/n4041 ) );
  MUX U8454 ( .IN0(\u_a23_core/u_execute/u_register_bank/r9[0] ), .IN1(n6098), 
        .SEL(n6212), .F(\u_a23_core/u_execute/u_register_bank/n4039 ) );
  ANDN U8455 ( .A(\u_a23_core/reg_bank_wen[9] ), .B(n6099), .Z(n6212) );
  MUX U8456 ( .IN0(\u_a23_core/u_execute/u_register_bank/r10[31] ), .IN1(n6066), .SEL(n6213), .F(\u_a23_core/u_execute/u_register_bank/n4037 ) );
  NAND U8457 ( .A(n6214), .B(n6215), .Z(n6066) );
  NAND U8458 ( .A(\u_a23_core/u_execute/multiply_out[31] ), .B(
        \u_a23_core/reg_write_sel[1] ), .Z(n6215) );
  AND U8459 ( .A(n6216), .B(n6217), .Z(n6214) );
  NAND U8460 ( .A(\u_a23_core/u_execute/save_int_pc_m4[31] ), .B(n6218), .Z(
        n6217) );
  NANDN U8461 ( .B(n6219), .A(\u_a23_core/u_execute/alu_out[31] ), .Z(n6216)
         );
  MUX U8462 ( .IN0(\u_a23_core/u_execute/u_register_bank/r10[30] ), .IN1(n6068), .SEL(n6213), .F(\u_a23_core/u_execute/u_register_bank/n4035 ) );
  NAND U8463 ( .A(n6220), .B(n6221), .Z(n6068) );
  NAND U8464 ( .A(\u_a23_core/reg_write_sel[1] ), .B(
        \u_a23_core/u_execute/multiply_out[30] ), .Z(n6221) );
  AND U8465 ( .A(n6222), .B(n6223), .Z(n6220) );
  NAND U8466 ( .A(\u_a23_core/u_execute/save_int_pc_m4[30] ), .B(n6218), .Z(
        n6223) );
  NANDN U8467 ( .B(n6219), .A(\u_a23_core/u_execute/alu_out[30] ), .Z(n6222)
         );
  MUX U8468 ( .IN0(\u_a23_core/u_execute/u_register_bank/r10[29] ), .IN1(n6069), .SEL(n6213), .F(\u_a23_core/u_execute/u_register_bank/n4033 ) );
  NAND U8469 ( .A(n6224), .B(n6225), .Z(n6069) );
  NAND U8470 ( .A(\u_a23_core/reg_write_sel[1] ), .B(
        \u_a23_core/u_execute/multiply_out[29] ), .Z(n6225) );
  AND U8471 ( .A(n6226), .B(n6227), .Z(n6224) );
  NAND U8472 ( .A(\u_a23_core/u_execute/save_int_pc_m4[29] ), .B(n6218), .Z(
        n6227) );
  NANDN U8473 ( .B(n6219), .A(\u_a23_core/u_execute/alu_out[29] ), .Z(n6226)
         );
  MUX U8474 ( .IN0(\u_a23_core/u_execute/u_register_bank/r10[28] ), .IN1(n6070), .SEL(n6213), .F(\u_a23_core/u_execute/u_register_bank/n4031 ) );
  NAND U8475 ( .A(n6228), .B(n6229), .Z(n6070) );
  NAND U8476 ( .A(\u_a23_core/reg_write_sel[1] ), .B(
        \u_a23_core/u_execute/multiply_out[28] ), .Z(n6229) );
  AND U8477 ( .A(n6230), .B(n6231), .Z(n6228) );
  NAND U8478 ( .A(\u_a23_core/u_execute/save_int_pc_m4[28] ), .B(n6218), .Z(
        n6231) );
  NANDN U8479 ( .B(n6219), .A(\u_a23_core/u_execute/alu_out[28] ), .Z(n6230)
         );
  MUX U8480 ( .IN0(\u_a23_core/u_execute/u_register_bank/r10[27] ), .IN1(n6071), .SEL(n6213), .F(\u_a23_core/u_execute/u_register_bank/n4029 ) );
  NAND U8481 ( .A(n6232), .B(n6233), .Z(n6071) );
  NAND U8482 ( .A(\u_a23_core/reg_write_sel[1] ), .B(
        \u_a23_core/u_execute/multiply_out[27] ), .Z(n6233) );
  AND U8483 ( .A(n6234), .B(n6235), .Z(n6232) );
  NANDN U8484 ( .B(n6219), .A(\u_a23_core/u_execute/alu_out[27] ), .Z(n6234)
         );
  MUX U8485 ( .IN0(\u_a23_core/u_execute/u_register_bank/r10[26] ), .IN1(n6072), .SEL(n6213), .F(\u_a23_core/u_execute/u_register_bank/n4027 ) );
  NAND U8486 ( .A(n6236), .B(n6237), .Z(n6072) );
  NAND U8487 ( .A(\u_a23_core/reg_write_sel[1] ), .B(
        \u_a23_core/u_execute/multiply_out[26] ), .Z(n6237) );
  AND U8488 ( .A(n6238), .B(n6235), .Z(n6236) );
  IV U8489 ( .A(n6218), .Z(n6235) );
  NANDN U8490 ( .B(n6219), .A(\u_a23_core/u_execute/alu_out[26] ), .Z(n6238)
         );
  MUX U8491 ( .IN0(\u_a23_core/u_execute/u_register_bank/r10[25] ), .IN1(n6073), .SEL(n6213), .F(\u_a23_core/u_execute/u_register_bank/n4025 ) );
  NAND U8492 ( .A(n6239), .B(n6240), .Z(n6073) );
  NAND U8493 ( .A(\u_a23_core/reg_write_sel[1] ), .B(
        \u_a23_core/u_execute/multiply_out[25] ), .Z(n6240) );
  AND U8494 ( .A(n6241), .B(n6242), .Z(n6239) );
  NAND U8495 ( .A(n6218), .B(\u_a23_core/u_execute/pc_minus4[25] ), .Z(n6242)
         );
  NANDN U8496 ( .B(n6219), .A(\u_a23_core/u_execute/alu_out_pc_filtered[25] ), 
        .Z(n6241) );
  MUX U8497 ( .IN0(\u_a23_core/u_execute/u_register_bank/r10[24] ), .IN1(n6074), .SEL(n6213), .F(\u_a23_core/u_execute/u_register_bank/n4023 ) );
  NAND U8498 ( .A(n6243), .B(n6244), .Z(n6074) );
  NAND U8499 ( .A(\u_a23_core/reg_write_sel[1] ), .B(
        \u_a23_core/u_execute/multiply_out[24] ), .Z(n6244) );
  AND U8500 ( .A(n6245), .B(n6246), .Z(n6243) );
  NAND U8501 ( .A(n6218), .B(\u_a23_core/u_execute/pc_minus4[24] ), .Z(n6246)
         );
  NANDN U8502 ( .B(n6219), .A(\u_a23_core/u_execute/alu_out_pc_filtered[24] ), 
        .Z(n6245) );
  MUX U8503 ( .IN0(\u_a23_core/u_execute/u_register_bank/r10[23] ), .IN1(n6075), .SEL(n6213), .F(\u_a23_core/u_execute/u_register_bank/n4021 ) );
  NAND U8504 ( .A(n6247), .B(n6248), .Z(n6075) );
  NAND U8505 ( .A(\u_a23_core/reg_write_sel[1] ), .B(
        \u_a23_core/u_execute/multiply_out[23] ), .Z(n6248) );
  AND U8506 ( .A(n6249), .B(n6250), .Z(n6247) );
  NAND U8507 ( .A(n6218), .B(\u_a23_core/u_execute/pc_minus4[23] ), .Z(n6250)
         );
  NANDN U8508 ( .B(n6219), .A(\u_a23_core/u_execute/alu_out_pc_filtered[23] ), 
        .Z(n6249) );
  MUX U8509 ( .IN0(\u_a23_core/u_execute/u_register_bank/r10[22] ), .IN1(n6076), .SEL(n6213), .F(\u_a23_core/u_execute/u_register_bank/n4019 ) );
  NAND U8510 ( .A(n6251), .B(n6252), .Z(n6076) );
  NAND U8511 ( .A(\u_a23_core/reg_write_sel[1] ), .B(
        \u_a23_core/u_execute/multiply_out[22] ), .Z(n6252) );
  AND U8512 ( .A(n6253), .B(n6254), .Z(n6251) );
  NAND U8513 ( .A(n6218), .B(\u_a23_core/u_execute/pc_minus4[22] ), .Z(n6254)
         );
  NANDN U8514 ( .B(n6219), .A(\u_a23_core/u_execute/alu_out_pc_filtered[22] ), 
        .Z(n6253) );
  MUX U8515 ( .IN0(\u_a23_core/u_execute/u_register_bank/r10[21] ), .IN1(n6077), .SEL(n6213), .F(\u_a23_core/u_execute/u_register_bank/n4017 ) );
  NAND U8516 ( .A(n6255), .B(n6256), .Z(n6077) );
  NAND U8517 ( .A(\u_a23_core/reg_write_sel[1] ), .B(
        \u_a23_core/u_execute/multiply_out[21] ), .Z(n6256) );
  AND U8518 ( .A(n6257), .B(n6258), .Z(n6255) );
  NAND U8519 ( .A(n6218), .B(\u_a23_core/u_execute/pc_minus4[21] ), .Z(n6258)
         );
  NANDN U8520 ( .B(n6219), .A(\u_a23_core/u_execute/alu_out_pc_filtered[21] ), 
        .Z(n6257) );
  MUX U8521 ( .IN0(\u_a23_core/u_execute/u_register_bank/r10[20] ), .IN1(n6078), .SEL(n6213), .F(\u_a23_core/u_execute/u_register_bank/n4015 ) );
  NAND U8522 ( .A(n6259), .B(n6260), .Z(n6078) );
  NAND U8523 ( .A(\u_a23_core/reg_write_sel[1] ), .B(
        \u_a23_core/u_execute/multiply_out[20] ), .Z(n6260) );
  AND U8524 ( .A(n6261), .B(n6262), .Z(n6259) );
  NAND U8525 ( .A(n6218), .B(\u_a23_core/u_execute/pc_minus4[20] ), .Z(n6262)
         );
  NANDN U8526 ( .B(n6219), .A(\u_a23_core/u_execute/alu_out_pc_filtered[20] ), 
        .Z(n6261) );
  MUX U8527 ( .IN0(\u_a23_core/u_execute/u_register_bank/r10[19] ), .IN1(n6079), .SEL(n6213), .F(\u_a23_core/u_execute/u_register_bank/n4013 ) );
  NAND U8528 ( .A(n6263), .B(n6264), .Z(n6079) );
  NAND U8529 ( .A(\u_a23_core/reg_write_sel[1] ), .B(
        \u_a23_core/u_execute/multiply_out[19] ), .Z(n6264) );
  AND U8530 ( .A(n6265), .B(n6266), .Z(n6263) );
  NAND U8531 ( .A(n6218), .B(\u_a23_core/u_execute/pc_minus4[19] ), .Z(n6266)
         );
  NANDN U8532 ( .B(n6219), .A(\u_a23_core/u_execute/alu_out_pc_filtered[19] ), 
        .Z(n6265) );
  MUX U8533 ( .IN0(\u_a23_core/u_execute/u_register_bank/r10[18] ), .IN1(n6080), .SEL(n6213), .F(\u_a23_core/u_execute/u_register_bank/n4011 ) );
  NAND U8534 ( .A(n6267), .B(n6268), .Z(n6080) );
  NAND U8535 ( .A(\u_a23_core/reg_write_sel[1] ), .B(
        \u_a23_core/u_execute/multiply_out[18] ), .Z(n6268) );
  AND U8536 ( .A(n6269), .B(n6270), .Z(n6267) );
  NAND U8537 ( .A(n6218), .B(\u_a23_core/u_execute/pc_minus4[18] ), .Z(n6270)
         );
  NANDN U8538 ( .B(n6219), .A(\u_a23_core/u_execute/alu_out_pc_filtered[18] ), 
        .Z(n6269) );
  MUX U8539 ( .IN0(\u_a23_core/u_execute/u_register_bank/r10[17] ), .IN1(n6081), .SEL(n6213), .F(\u_a23_core/u_execute/u_register_bank/n4009 ) );
  NAND U8540 ( .A(n6271), .B(n6272), .Z(n6081) );
  NAND U8541 ( .A(\u_a23_core/reg_write_sel[1] ), .B(
        \u_a23_core/u_execute/multiply_out[17] ), .Z(n6272) );
  AND U8542 ( .A(n6273), .B(n6274), .Z(n6271) );
  NAND U8543 ( .A(n6218), .B(\u_a23_core/u_execute/pc_minus4[17] ), .Z(n6274)
         );
  NANDN U8544 ( .B(n6219), .A(\u_a23_core/u_execute/alu_out_pc_filtered[17] ), 
        .Z(n6273) );
  MUX U8545 ( .IN0(\u_a23_core/u_execute/u_register_bank/r10[16] ), .IN1(n6082), .SEL(n6213), .F(\u_a23_core/u_execute/u_register_bank/n4007 ) );
  NAND U8546 ( .A(n6275), .B(n6276), .Z(n6082) );
  NAND U8547 ( .A(\u_a23_core/reg_write_sel[1] ), .B(
        \u_a23_core/u_execute/multiply_out[16] ), .Z(n6276) );
  AND U8548 ( .A(n6277), .B(n6278), .Z(n6275) );
  NAND U8549 ( .A(n6218), .B(\u_a23_core/u_execute/pc_minus4[16] ), .Z(n6278)
         );
  NANDN U8550 ( .B(n6219), .A(\u_a23_core/u_execute/alu_out_pc_filtered[16] ), 
        .Z(n6277) );
  MUX U8551 ( .IN0(\u_a23_core/u_execute/u_register_bank/r10[15] ), .IN1(n6083), .SEL(n6213), .F(\u_a23_core/u_execute/u_register_bank/n4005 ) );
  NAND U8552 ( .A(n6279), .B(n6280), .Z(n6083) );
  NAND U8553 ( .A(\u_a23_core/reg_write_sel[1] ), .B(
        \u_a23_core/u_execute/multiply_out[15] ), .Z(n6280) );
  AND U8554 ( .A(n6281), .B(n6282), .Z(n6279) );
  NAND U8555 ( .A(n6218), .B(\u_a23_core/u_execute/pc_minus4[15] ), .Z(n6282)
         );
  NANDN U8556 ( .B(n6219), .A(\u_a23_core/u_execute/alu_out_pc_filtered[15] ), 
        .Z(n6281) );
  MUX U8557 ( .IN0(\u_a23_core/u_execute/u_register_bank/r10[14] ), .IN1(n6084), .SEL(n6213), .F(\u_a23_core/u_execute/u_register_bank/n4003 ) );
  NAND U8558 ( .A(n6283), .B(n6284), .Z(n6084) );
  NAND U8559 ( .A(\u_a23_core/reg_write_sel[1] ), .B(
        \u_a23_core/u_execute/multiply_out[14] ), .Z(n6284) );
  AND U8560 ( .A(n6285), .B(n6286), .Z(n6283) );
  NAND U8561 ( .A(n6218), .B(\u_a23_core/u_execute/pc_minus4[14] ), .Z(n6286)
         );
  NANDN U8562 ( .B(n6219), .A(\u_a23_core/u_execute/alu_out_pc_filtered[14] ), 
        .Z(n6285) );
  MUX U8563 ( .IN0(\u_a23_core/u_execute/u_register_bank/r10[13] ), .IN1(n6085), .SEL(n6213), .F(\u_a23_core/u_execute/u_register_bank/n4001 ) );
  NAND U8564 ( .A(n6287), .B(n6288), .Z(n6085) );
  NAND U8565 ( .A(\u_a23_core/reg_write_sel[1] ), .B(
        \u_a23_core/u_execute/multiply_out[13] ), .Z(n6288) );
  AND U8566 ( .A(n6289), .B(n6290), .Z(n6287) );
  NAND U8567 ( .A(n6218), .B(\u_a23_core/u_execute/pc_minus4[13] ), .Z(n6290)
         );
  NANDN U8568 ( .B(n6219), .A(\u_a23_core/u_execute/alu_out_pc_filtered[13] ), 
        .Z(n6289) );
  MUX U8569 ( .IN0(\u_a23_core/u_execute/u_register_bank/r10[12] ), .IN1(n6086), .SEL(n6213), .F(\u_a23_core/u_execute/u_register_bank/n3999 ) );
  NAND U8570 ( .A(n6291), .B(n6292), .Z(n6086) );
  NAND U8571 ( .A(\u_a23_core/reg_write_sel[1] ), .B(
        \u_a23_core/u_execute/multiply_out[12] ), .Z(n6292) );
  AND U8572 ( .A(n6293), .B(n6294), .Z(n6291) );
  NAND U8573 ( .A(n6218), .B(\u_a23_core/u_execute/pc_minus4[12] ), .Z(n6294)
         );
  NANDN U8574 ( .B(n6219), .A(\u_a23_core/u_execute/alu_out_pc_filtered[12] ), 
        .Z(n6293) );
  MUX U8575 ( .IN0(\u_a23_core/u_execute/u_register_bank/r10[11] ), .IN1(n6087), .SEL(n6213), .F(\u_a23_core/u_execute/u_register_bank/n3997 ) );
  NAND U8576 ( .A(n6295), .B(n6296), .Z(n6087) );
  NAND U8577 ( .A(\u_a23_core/reg_write_sel[1] ), .B(
        \u_a23_core/u_execute/multiply_out[11] ), .Z(n6296) );
  AND U8578 ( .A(n6297), .B(n6298), .Z(n6295) );
  NAND U8579 ( .A(n6218), .B(\u_a23_core/u_execute/pc_minus4[11] ), .Z(n6298)
         );
  NANDN U8580 ( .B(n6219), .A(\u_a23_core/u_execute/alu_out_pc_filtered[11] ), 
        .Z(n6297) );
  MUX U8581 ( .IN0(\u_a23_core/u_execute/u_register_bank/r10[10] ), .IN1(n6088), .SEL(n6213), .F(\u_a23_core/u_execute/u_register_bank/n3995 ) );
  NAND U8582 ( .A(n6299), .B(n6300), .Z(n6088) );
  NAND U8583 ( .A(\u_a23_core/reg_write_sel[1] ), .B(
        \u_a23_core/u_execute/multiply_out[10] ), .Z(n6300) );
  AND U8584 ( .A(n6301), .B(n6302), .Z(n6299) );
  NAND U8585 ( .A(n6218), .B(\u_a23_core/u_execute/pc_minus4[10] ), .Z(n6302)
         );
  NANDN U8586 ( .B(n6219), .A(\u_a23_core/u_execute/alu_out_pc_filtered[10] ), 
        .Z(n6301) );
  MUX U8587 ( .IN0(\u_a23_core/u_execute/u_register_bank/r10[9] ), .IN1(n6089), 
        .SEL(n6213), .F(\u_a23_core/u_execute/u_register_bank/n3993 ) );
  NAND U8588 ( .A(n6303), .B(n6304), .Z(n6089) );
  NAND U8589 ( .A(\u_a23_core/reg_write_sel[1] ), .B(
        \u_a23_core/u_execute/multiply_out[9] ), .Z(n6304) );
  AND U8590 ( .A(n6305), .B(n6306), .Z(n6303) );
  NAND U8591 ( .A(n6218), .B(\u_a23_core/u_execute/pc_minus4[9] ), .Z(n6306)
         );
  NANDN U8592 ( .B(n6219), .A(\u_a23_core/u_execute/alu_out_pc_filtered[9] ), 
        .Z(n6305) );
  MUX U8593 ( .IN0(\u_a23_core/u_execute/u_register_bank/r10[8] ), .IN1(n6090), 
        .SEL(n6213), .F(\u_a23_core/u_execute/u_register_bank/n3991 ) );
  NAND U8594 ( .A(n6307), .B(n6308), .Z(n6090) );
  NAND U8595 ( .A(\u_a23_core/reg_write_sel[1] ), .B(
        \u_a23_core/u_execute/multiply_out[8] ), .Z(n6308) );
  AND U8596 ( .A(n6309), .B(n6310), .Z(n6307) );
  NAND U8597 ( .A(n6218), .B(\u_a23_core/u_execute/pc_minus4[8] ), .Z(n6310)
         );
  NANDN U8598 ( .B(n6219), .A(\u_a23_core/u_execute/alu_out_pc_filtered[8] ), 
        .Z(n6309) );
  MUX U8599 ( .IN0(\u_a23_core/u_execute/u_register_bank/r10[7] ), .IN1(n6091), 
        .SEL(n6213), .F(\u_a23_core/u_execute/u_register_bank/n3989 ) );
  NAND U8600 ( .A(n6311), .B(n6312), .Z(n6091) );
  NAND U8601 ( .A(\u_a23_core/reg_write_sel[1] ), .B(
        \u_a23_core/u_execute/multiply_out[7] ), .Z(n6312) );
  AND U8602 ( .A(n6313), .B(n6314), .Z(n6311) );
  NAND U8603 ( .A(n6218), .B(\u_a23_core/u_execute/pc_minus4[7] ), .Z(n6314)
         );
  NANDN U8604 ( .B(n6219), .A(\u_a23_core/u_execute/alu_out_pc_filtered[7] ), 
        .Z(n6313) );
  MUX U8605 ( .IN0(\u_a23_core/u_execute/u_register_bank/r10[6] ), .IN1(n6092), 
        .SEL(n6213), .F(\u_a23_core/u_execute/u_register_bank/n3987 ) );
  NAND U8606 ( .A(n6315), .B(n6316), .Z(n6092) );
  NAND U8607 ( .A(\u_a23_core/reg_write_sel[1] ), .B(
        \u_a23_core/u_execute/multiply_out[6] ), .Z(n6316) );
  AND U8608 ( .A(n6317), .B(n6318), .Z(n6315) );
  NAND U8609 ( .A(n6218), .B(\u_a23_core/u_execute/pc_minus4[6] ), .Z(n6318)
         );
  NANDN U8610 ( .B(n6219), .A(\u_a23_core/u_execute/alu_out_pc_filtered[6] ), 
        .Z(n6317) );
  MUX U8611 ( .IN0(\u_a23_core/u_execute/u_register_bank/r10[5] ), .IN1(n6093), 
        .SEL(n6213), .F(\u_a23_core/u_execute/u_register_bank/n3985 ) );
  NAND U8612 ( .A(n6319), .B(n6320), .Z(n6093) );
  NAND U8613 ( .A(\u_a23_core/reg_write_sel[1] ), .B(
        \u_a23_core/u_execute/multiply_out[5] ), .Z(n6320) );
  AND U8614 ( .A(n6321), .B(n6322), .Z(n6319) );
  NAND U8615 ( .A(n6218), .B(\u_a23_core/u_execute/pc_minus4[5] ), .Z(n6322)
         );
  NANDN U8616 ( .B(n6219), .A(\u_a23_core/u_execute/alu_out_pc_filtered[5] ), 
        .Z(n6321) );
  MUX U8617 ( .IN0(\u_a23_core/u_execute/u_register_bank/r10[4] ), .IN1(n6094), 
        .SEL(n6213), .F(\u_a23_core/u_execute/u_register_bank/n3983 ) );
  NAND U8618 ( .A(n6323), .B(n6324), .Z(n6094) );
  NAND U8619 ( .A(\u_a23_core/reg_write_sel[1] ), .B(
        \u_a23_core/u_execute/multiply_out[4] ), .Z(n6324) );
  AND U8620 ( .A(n6325), .B(n6326), .Z(n6323) );
  NAND U8621 ( .A(n6218), .B(\u_a23_core/u_execute/pc_minus4[4] ), .Z(n6326)
         );
  NANDN U8622 ( .B(n6219), .A(\u_a23_core/u_execute/alu_out_pc_filtered[4] ), 
        .Z(n6325) );
  MUX U8623 ( .IN0(\u_a23_core/u_execute/u_register_bank/r10[3] ), .IN1(n6095), 
        .SEL(n6213), .F(\u_a23_core/u_execute/u_register_bank/n3981 ) );
  NAND U8624 ( .A(n6327), .B(n6328), .Z(n6095) );
  NAND U8625 ( .A(\u_a23_core/reg_write_sel[1] ), .B(
        \u_a23_core/u_execute/multiply_out[3] ), .Z(n6328) );
  AND U8626 ( .A(n6329), .B(n6330), .Z(n6327) );
  NAND U8627 ( .A(n6218), .B(\u_a23_core/u_execute/pc_minus4[3] ), .Z(n6330)
         );
  NANDN U8628 ( .B(n6219), .A(\u_a23_core/u_execute/alu_out_pc_filtered[3] ), 
        .Z(n6329) );
  MUX U8629 ( .IN0(\u_a23_core/u_execute/u_register_bank/r10[2] ), .IN1(n6096), 
        .SEL(n6213), .F(\u_a23_core/u_execute/u_register_bank/n3979 ) );
  NAND U8630 ( .A(n6331), .B(n6332), .Z(n6096) );
  NAND U8631 ( .A(\u_a23_core/reg_write_sel[1] ), .B(
        \u_a23_core/u_execute/multiply_out[2] ), .Z(n6332) );
  AND U8632 ( .A(n6333), .B(n6334), .Z(n6331) );
  NAND U8633 ( .A(n6201), .B(n6218), .Z(n6334) );
  ANDN U8634 ( .A(\u_a23_core/reg_write_sel[0] ), .B(
        \u_a23_core/reg_write_sel[1] ), .Z(n6218) );
  IV U8635 ( .A(\u_a23_core/u_execute/pc[2] ), .Z(n6201) );
  NANDN U8636 ( .B(n6219), .A(\u_a23_core/u_execute/alu_out_pc_filtered[2] ), 
        .Z(n6333) );
  MUX U8637 ( .IN0(\u_a23_core/u_execute/u_register_bank/r10[1] ), .IN1(n6097), 
        .SEL(n6213), .F(\u_a23_core/u_execute/u_register_bank/n3977 ) );
  NAND U8638 ( .A(n6335), .B(n6336), .Z(n6097) );
  NANDN U8639 ( .B(n6219), .A(n6337), .Z(n6336) );
  NAND U8640 ( .A(\u_a23_core/reg_write_sel[1] ), .B(
        \u_a23_core/u_execute/multiply_out[1] ), .Z(n6335) );
  MUX U8641 ( .IN0(\u_a23_core/u_execute/u_register_bank/r10[0] ), .IN1(n6098), 
        .SEL(n6213), .F(\u_a23_core/u_execute/u_register_bank/n3975 ) );
  ANDN U8642 ( .A(\u_a23_core/reg_bank_wen[10] ), .B(n6099), .Z(n6213) );
  NAND U8643 ( .A(n6338), .B(n6339), .Z(n6098) );
  OR U8644 ( .A(n6219), .B(n6340), .Z(n6339) );
  OR U8645 ( .A(\u_a23_core/reg_write_sel[0] ), .B(
        \u_a23_core/reg_write_sel[1] ), .Z(n6219) );
  NAND U8646 ( .A(\u_a23_core/u_execute/multiply_out[0] ), .B(
        \u_a23_core/reg_write_sel[1] ), .Z(n6338) );
  NAND U8647 ( .A(n6341), .B(n6342), .Z(
        \u_a23_core/u_execute/u_multiply/sum34_b[9] ) );
  NAND U8648 ( .A(n6343), .B(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[9] ), .Z(n6342) );
  NAND U8649 ( .A(\u_a23_core/u_execute/rs[9] ), .B(n6344), .Z(n6341) );
  NAND U8650 ( .A(n6345), .B(n6346), .Z(
        \u_a23_core/u_execute/u_multiply/sum34_b[8] ) );
  NAND U8651 ( .A(n6343), .B(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[8] ), .Z(n6346) );
  NAND U8652 ( .A(\u_a23_core/u_execute/rs[8] ), .B(n6344), .Z(n6345) );
  NAND U8653 ( .A(n6347), .B(n6348), .Z(
        \u_a23_core/u_execute/u_multiply/sum34_b[7] ) );
  NAND U8654 ( .A(n6343), .B(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[7] ), .Z(n6348) );
  NAND U8655 ( .A(\u_a23_core/u_execute/rs[7] ), .B(n6344), .Z(n6347) );
  NAND U8656 ( .A(n6349), .B(n6350), .Z(
        \u_a23_core/u_execute/u_multiply/sum34_b[6] ) );
  NAND U8657 ( .A(n6343), .B(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[6] ), .Z(n6350) );
  NAND U8658 ( .A(\u_a23_core/u_execute/rs[6] ), .B(n6344), .Z(n6349) );
  NAND U8659 ( .A(n6351), .B(n6352), .Z(
        \u_a23_core/u_execute/u_multiply/sum34_b[5] ) );
  NAND U8660 ( .A(n6343), .B(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[5] ), .Z(n6352) );
  NAND U8661 ( .A(\u_a23_core/u_execute/rs[5] ), .B(n6344), .Z(n6351) );
  NAND U8662 ( .A(n6353), .B(n6354), .Z(
        \u_a23_core/u_execute/u_multiply/sum34_b[4] ) );
  NAND U8663 ( .A(n6343), .B(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[4] ), .Z(n6354) );
  NAND U8664 ( .A(\u_a23_core/u_execute/rs[4] ), .B(n6344), .Z(n6353) );
  NAND U8665 ( .A(n6355), .B(n6356), .Z(
        \u_a23_core/u_execute/u_multiply/sum34_b[3] ) );
  NAND U8666 ( .A(n6343), .B(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[3] ), .Z(n6356) );
  NAND U8667 ( .A(\u_a23_core/u_execute/rs[3] ), .B(n6344), .Z(n6355) );
  ANDN U8668 ( .A(n6343), .B(
        \u_a23_core/u_execute/u_multiply/add_90/carry[32] ), .Z(
        \u_a23_core/u_execute/u_multiply/sum34_b[33] ) );
  NAND U8669 ( .A(n6357), .B(n6358), .Z(
        \u_a23_core/u_execute/u_multiply/sum34_b[31] ) );
  NAND U8670 ( .A(n6343), .B(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[31] ), .Z(n6358) );
  NAND U8671 ( .A(\u_a23_core/u_execute/rs[31] ), .B(n6344), .Z(n6357) );
  NAND U8672 ( .A(n6359), .B(n6360), .Z(
        \u_a23_core/u_execute/u_multiply/sum34_b[30] ) );
  NAND U8673 ( .A(n6343), .B(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[30] ), .Z(n6360) );
  NAND U8674 ( .A(\u_a23_core/u_execute/rs[30] ), .B(n6344), .Z(n6359) );
  NAND U8675 ( .A(n6361), .B(n6362), .Z(
        \u_a23_core/u_execute/u_multiply/sum34_b[2] ) );
  NAND U8676 ( .A(n6343), .B(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[2] ), .Z(n6362) );
  NAND U8677 ( .A(\u_a23_core/u_execute/rs[2] ), .B(n6344), .Z(n6361) );
  NAND U8678 ( .A(n6363), .B(n6364), .Z(
        \u_a23_core/u_execute/u_multiply/sum34_b[29] ) );
  NAND U8679 ( .A(n6343), .B(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[29] ), .Z(n6364) );
  NAND U8680 ( .A(\u_a23_core/u_execute/rs[29] ), .B(n6344), .Z(n6363) );
  NAND U8681 ( .A(n6365), .B(n6366), .Z(
        \u_a23_core/u_execute/u_multiply/sum34_b[28] ) );
  NAND U8682 ( .A(n6343), .B(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[28] ), .Z(n6366) );
  NAND U8683 ( .A(\u_a23_core/u_execute/rs[28] ), .B(n6344), .Z(n6365) );
  NAND U8684 ( .A(n6367), .B(n6368), .Z(
        \u_a23_core/u_execute/u_multiply/sum34_b[27] ) );
  NAND U8685 ( .A(n6343), .B(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[27] ), .Z(n6368) );
  NAND U8686 ( .A(\u_a23_core/u_execute/rs[27] ), .B(n6344), .Z(n6367) );
  NAND U8687 ( .A(n6369), .B(n6370), .Z(
        \u_a23_core/u_execute/u_multiply/sum34_b[26] ) );
  NAND U8688 ( .A(n6343), .B(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[26] ), .Z(n6370) );
  NAND U8689 ( .A(\u_a23_core/u_execute/rs[26] ), .B(n6344), .Z(n6369) );
  NAND U8690 ( .A(n6371), .B(n6372), .Z(
        \u_a23_core/u_execute/u_multiply/sum34_b[25] ) );
  NAND U8691 ( .A(n6343), .B(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[25] ), .Z(n6372) );
  NAND U8692 ( .A(\u_a23_core/u_execute/rs[25] ), .B(n6344), .Z(n6371) );
  NAND U8693 ( .A(n6373), .B(n6374), .Z(
        \u_a23_core/u_execute/u_multiply/sum34_b[24] ) );
  NAND U8694 ( .A(n6343), .B(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[24] ), .Z(n6374) );
  NAND U8695 ( .A(\u_a23_core/u_execute/rs[24] ), .B(n6344), .Z(n6373) );
  NAND U8696 ( .A(n6375), .B(n6376), .Z(
        \u_a23_core/u_execute/u_multiply/sum34_b[23] ) );
  NAND U8697 ( .A(n6343), .B(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[23] ), .Z(n6376) );
  NAND U8698 ( .A(\u_a23_core/u_execute/rs[23] ), .B(n6344), .Z(n6375) );
  NAND U8699 ( .A(n6377), .B(n6378), .Z(
        \u_a23_core/u_execute/u_multiply/sum34_b[22] ) );
  NAND U8700 ( .A(n6343), .B(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[22] ), .Z(n6378) );
  NAND U8701 ( .A(\u_a23_core/u_execute/rs[22] ), .B(n6344), .Z(n6377) );
  NAND U8702 ( .A(n6379), .B(n6380), .Z(
        \u_a23_core/u_execute/u_multiply/sum34_b[21] ) );
  NAND U8703 ( .A(n6343), .B(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[21] ), .Z(n6380) );
  NAND U8704 ( .A(\u_a23_core/u_execute/rs[21] ), .B(n6344), .Z(n6379) );
  NAND U8705 ( .A(n6381), .B(n6382), .Z(
        \u_a23_core/u_execute/u_multiply/sum34_b[20] ) );
  NAND U8706 ( .A(n6343), .B(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[20] ), .Z(n6382) );
  NAND U8707 ( .A(\u_a23_core/u_execute/rs[20] ), .B(n6344), .Z(n6381) );
  NAND U8708 ( .A(n6383), .B(n6384), .Z(
        \u_a23_core/u_execute/u_multiply/sum34_b[1] ) );
  NAND U8709 ( .A(n6343), .B(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[1] ), .Z(n6384) );
  NAND U8710 ( .A(\u_a23_core/u_execute/rs[1] ), .B(n6344), .Z(n6383) );
  NAND U8711 ( .A(n6385), .B(n6386), .Z(
        \u_a23_core/u_execute/u_multiply/sum34_b[19] ) );
  NAND U8712 ( .A(n6343), .B(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[19] ), .Z(n6386) );
  NAND U8713 ( .A(\u_a23_core/u_execute/rs[19] ), .B(n6344), .Z(n6385) );
  NAND U8714 ( .A(n6387), .B(n6388), .Z(
        \u_a23_core/u_execute/u_multiply/sum34_b[18] ) );
  NAND U8715 ( .A(n6343), .B(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[18] ), .Z(n6388) );
  NAND U8716 ( .A(\u_a23_core/u_execute/rs[18] ), .B(n6344), .Z(n6387) );
  NAND U8717 ( .A(n6389), .B(n6390), .Z(
        \u_a23_core/u_execute/u_multiply/sum34_b[17] ) );
  NAND U8718 ( .A(n6343), .B(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[17] ), .Z(n6390) );
  NAND U8719 ( .A(\u_a23_core/u_execute/rs[17] ), .B(n6344), .Z(n6389) );
  NAND U8720 ( .A(n6391), .B(n6392), .Z(
        \u_a23_core/u_execute/u_multiply/sum34_b[16] ) );
  NAND U8721 ( .A(n6343), .B(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[16] ), .Z(n6392) );
  NAND U8722 ( .A(\u_a23_core/u_execute/rs[16] ), .B(n6344), .Z(n6391) );
  NAND U8723 ( .A(n6393), .B(n6394), .Z(
        \u_a23_core/u_execute/u_multiply/sum34_b[15] ) );
  NAND U8724 ( .A(n6343), .B(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[15] ), .Z(n6394) );
  NAND U8725 ( .A(\u_a23_core/u_execute/rs[15] ), .B(n6344), .Z(n6393) );
  NAND U8726 ( .A(n6395), .B(n6396), .Z(
        \u_a23_core/u_execute/u_multiply/sum34_b[14] ) );
  NAND U8727 ( .A(n6343), .B(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[14] ), .Z(n6396) );
  NAND U8728 ( .A(\u_a23_core/u_execute/rs[14] ), .B(n6344), .Z(n6395) );
  NAND U8729 ( .A(n6397), .B(n6398), .Z(
        \u_a23_core/u_execute/u_multiply/sum34_b[13] ) );
  NAND U8730 ( .A(n6343), .B(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[13] ), .Z(n6398) );
  NAND U8731 ( .A(\u_a23_core/u_execute/rs[13] ), .B(n6344), .Z(n6397) );
  NAND U8732 ( .A(n6399), .B(n6400), .Z(
        \u_a23_core/u_execute/u_multiply/sum34_b[12] ) );
  NAND U8733 ( .A(n6343), .B(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[12] ), .Z(n6400) );
  NAND U8734 ( .A(\u_a23_core/u_execute/rs[12] ), .B(n6344), .Z(n6399) );
  NAND U8735 ( .A(n6401), .B(n6402), .Z(
        \u_a23_core/u_execute/u_multiply/sum34_b[11] ) );
  NAND U8736 ( .A(n6343), .B(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[11] ), .Z(n6402) );
  NAND U8737 ( .A(\u_a23_core/u_execute/rs[11] ), .B(n6344), .Z(n6401) );
  NAND U8738 ( .A(n6403), .B(n6404), .Z(
        \u_a23_core/u_execute/u_multiply/sum34_b[10] ) );
  NAND U8739 ( .A(n6343), .B(
        \u_a23_core/u_execute/u_multiply/multiplier_bar[10] ), .Z(n6404) );
  NAND U8740 ( .A(\u_a23_core/u_execute/rs[10] ), .B(n6344), .Z(n6403) );
  AND U8741 ( .A(n6405), .B(\u_a23_core/u_execute/rs[0] ), .Z(
        \u_a23_core/u_execute/u_multiply/sum34_b[0] ) );
  OR U8742 ( .A(n6343), .B(n6344), .Z(n6405) );
  ANDN U8743 ( .A(\u_a23_core/u_execute/u_multiply/product_0 ), .B(
        \u_a23_core/u_execute/multiply_out[0] ), .Z(n6344) );
  NOR U8744 ( .A(n6406), .B(\u_a23_core/u_execute/u_multiply/product_0 ), .Z(
        n6343) );
  IV U8745 ( .A(n6407), .Z(\u_a23_core/u_execute/u_multiply/n611 ) );
  MUX U8746 ( .IN0(n6408), .IN1(n6409), .SEL(\u_a23_core/multiply_function[0] ), .F(n6407) );
  NAND U8747 ( .A(n6408), .B(n6410), .Z(n6409) );
  NAND U8748 ( .A(n6411), .B(n6412), .Z(\u_a23_core/u_execute/u_multiply/n610 ) );
  NANDN U8749 ( .B(n6413), .A(\u_a23_core/u_execute/multiply_out[0] ), .Z(
        n6412) );
  NAND U8750 ( .A(n6414), .B(\u_a23_core/u_execute/u_multiply/product_0 ), .Z(
        n6411) );
  NAND U8751 ( .A(n6415), .B(n6416), .Z(\u_a23_core/u_execute/u_multiply/n609 ) );
  NAND U8752 ( .A(n6417), .B(\u_a23_core/u_execute/u_multiply/sum[0] ), .Z(
        n6416) );
  NAND U8753 ( .A(n6418), .B(\u_a23_core/u_execute/u_multiply/product[33] ), 
        .Z(n6415) );
  NAND U8754 ( .A(n6419), .B(n6420), .Z(\u_a23_core/u_execute/u_multiply/n608 ) );
  AND U8755 ( .A(n6421), .B(n6422), .Z(n6420) );
  NAND U8756 ( .A(n6423), .B(\u_a23_core/u_execute/u_multiply/sum_acc1[0] ), 
        .Z(n6422) );
  NANDN U8757 ( .B(n6424), .A(n6425), .Z(n6421) );
  AND U8758 ( .A(n6426), .B(n6427), .Z(n6419) );
  NANDN U8759 ( .B(n6413), .A(\u_a23_core/u_execute/multiply_out[1] ), .Z(
        n6427) );
  NAND U8760 ( .A(\u_a23_core/u_execute/multiply_out[0] ), .B(n6414), .Z(n6426) );
  NAND U8761 ( .A(n6428), .B(n6429), .Z(\u_a23_core/u_execute/u_multiply/n607 ) );
  AND U8762 ( .A(n6430), .B(n6431), .Z(n6429) );
  NAND U8763 ( .A(n6423), .B(\u_a23_core/u_execute/u_multiply/sum_acc1[1] ), 
        .Z(n6431) );
  NANDN U8764 ( .B(n6432), .A(n6425), .Z(n6430) );
  AND U8765 ( .A(n6433), .B(n6434), .Z(n6428) );
  NANDN U8766 ( .B(n6413), .A(\u_a23_core/u_execute/multiply_out[2] ), .Z(
        n6434) );
  NAND U8767 ( .A(n6414), .B(\u_a23_core/u_execute/multiply_out[1] ), .Z(n6433) );
  NAND U8768 ( .A(n6435), .B(n6436), .Z(\u_a23_core/u_execute/u_multiply/n606 ) );
  AND U8769 ( .A(n6437), .B(n6438), .Z(n6436) );
  NAND U8770 ( .A(n6423), .B(\u_a23_core/u_execute/u_multiply/sum_acc1[2] ), 
        .Z(n6438) );
  NANDN U8771 ( .B(n6439), .A(n6425), .Z(n6437) );
  AND U8772 ( .A(n6440), .B(n6441), .Z(n6435) );
  NANDN U8773 ( .B(n6413), .A(\u_a23_core/u_execute/multiply_out[3] ), .Z(
        n6441) );
  NAND U8774 ( .A(n6414), .B(\u_a23_core/u_execute/multiply_out[2] ), .Z(n6440) );
  NAND U8775 ( .A(n6442), .B(n6443), .Z(\u_a23_core/u_execute/u_multiply/n605 ) );
  AND U8776 ( .A(n6444), .B(n6445), .Z(n6443) );
  NAND U8777 ( .A(n6423), .B(\u_a23_core/u_execute/u_multiply/sum_acc1[3] ), 
        .Z(n6445) );
  NANDN U8778 ( .B(n6446), .A(n6425), .Z(n6444) );
  AND U8779 ( .A(n6447), .B(n6448), .Z(n6442) );
  NANDN U8780 ( .B(n6413), .A(\u_a23_core/u_execute/multiply_out[4] ), .Z(
        n6448) );
  NAND U8781 ( .A(n6414), .B(\u_a23_core/u_execute/multiply_out[3] ), .Z(n6447) );
  NAND U8782 ( .A(n6449), .B(n6450), .Z(\u_a23_core/u_execute/u_multiply/n604 ) );
  AND U8783 ( .A(n6451), .B(n6452), .Z(n6450) );
  NAND U8784 ( .A(n6423), .B(\u_a23_core/u_execute/u_multiply/sum_acc1[4] ), 
        .Z(n6452) );
  NANDN U8785 ( .B(n6453), .A(n6425), .Z(n6451) );
  AND U8786 ( .A(n6454), .B(n6455), .Z(n6449) );
  NANDN U8787 ( .B(n6413), .A(\u_a23_core/u_execute/multiply_out[5] ), .Z(
        n6455) );
  NAND U8788 ( .A(n6414), .B(\u_a23_core/u_execute/multiply_out[4] ), .Z(n6454) );
  NAND U8789 ( .A(n6456), .B(n6457), .Z(\u_a23_core/u_execute/u_multiply/n603 ) );
  AND U8790 ( .A(n6458), .B(n6459), .Z(n6457) );
  NAND U8791 ( .A(n6423), .B(\u_a23_core/u_execute/u_multiply/sum_acc1[5] ), 
        .Z(n6459) );
  NANDN U8792 ( .B(n6460), .A(n6425), .Z(n6458) );
  AND U8793 ( .A(n6461), .B(n6462), .Z(n6456) );
  NANDN U8794 ( .B(n6413), .A(\u_a23_core/u_execute/multiply_out[6] ), .Z(
        n6462) );
  NAND U8795 ( .A(n6414), .B(\u_a23_core/u_execute/multiply_out[5] ), .Z(n6461) );
  NAND U8796 ( .A(n6463), .B(n6464), .Z(\u_a23_core/u_execute/u_multiply/n602 ) );
  AND U8797 ( .A(n6465), .B(n6466), .Z(n6464) );
  NAND U8798 ( .A(n6423), .B(\u_a23_core/u_execute/u_multiply/sum_acc1[6] ), 
        .Z(n6466) );
  NANDN U8799 ( .B(n6467), .A(n6425), .Z(n6465) );
  AND U8800 ( .A(n6468), .B(n6469), .Z(n6463) );
  NANDN U8801 ( .B(n6413), .A(\u_a23_core/u_execute/multiply_out[7] ), .Z(
        n6469) );
  NAND U8802 ( .A(n6414), .B(\u_a23_core/u_execute/multiply_out[6] ), .Z(n6468) );
  NAND U8803 ( .A(n6470), .B(n6471), .Z(\u_a23_core/u_execute/u_multiply/n601 ) );
  AND U8804 ( .A(n6472), .B(n6473), .Z(n6471) );
  NAND U8805 ( .A(n6423), .B(\u_a23_core/u_execute/u_multiply/sum_acc1[7] ), 
        .Z(n6473) );
  NANDN U8806 ( .B(n6474), .A(n6425), .Z(n6472) );
  AND U8807 ( .A(n6475), .B(n6476), .Z(n6470) );
  NANDN U8808 ( .B(n6413), .A(\u_a23_core/u_execute/multiply_out[8] ), .Z(
        n6476) );
  NAND U8809 ( .A(n6414), .B(\u_a23_core/u_execute/multiply_out[7] ), .Z(n6475) );
  NAND U8810 ( .A(n6477), .B(n6478), .Z(\u_a23_core/u_execute/u_multiply/n600 ) );
  AND U8811 ( .A(n6479), .B(n6480), .Z(n6478) );
  NAND U8812 ( .A(n6423), .B(\u_a23_core/u_execute/u_multiply/sum_acc1[8] ), 
        .Z(n6480) );
  NANDN U8813 ( .B(n6481), .A(n6425), .Z(n6479) );
  AND U8814 ( .A(n6482), .B(n6483), .Z(n6477) );
  NANDN U8815 ( .B(n6413), .A(\u_a23_core/u_execute/multiply_out[9] ), .Z(
        n6483) );
  NAND U8816 ( .A(n6414), .B(\u_a23_core/u_execute/multiply_out[8] ), .Z(n6482) );
  NAND U8817 ( .A(n6484), .B(n6485), .Z(\u_a23_core/u_execute/u_multiply/n599 ) );
  AND U8818 ( .A(n6486), .B(n6487), .Z(n6485) );
  NAND U8819 ( .A(n6423), .B(\u_a23_core/u_execute/u_multiply/sum_acc1[9] ), 
        .Z(n6487) );
  NANDN U8820 ( .B(n6488), .A(n6425), .Z(n6486) );
  AND U8821 ( .A(n6489), .B(n6490), .Z(n6484) );
  NANDN U8822 ( .B(n6413), .A(\u_a23_core/u_execute/multiply_out[10] ), .Z(
        n6490) );
  NAND U8823 ( .A(n6414), .B(\u_a23_core/u_execute/multiply_out[9] ), .Z(n6489) );
  NAND U8824 ( .A(n6491), .B(n6492), .Z(\u_a23_core/u_execute/u_multiply/n598 ) );
  AND U8825 ( .A(n6493), .B(n6494), .Z(n6492) );
  NAND U8826 ( .A(n6423), .B(\u_a23_core/u_execute/u_multiply/sum_acc1[10] ), 
        .Z(n6494) );
  NANDN U8827 ( .B(n6495), .A(n6425), .Z(n6493) );
  AND U8828 ( .A(n6496), .B(n6497), .Z(n6491) );
  NANDN U8829 ( .B(n6413), .A(\u_a23_core/u_execute/multiply_out[11] ), .Z(
        n6497) );
  NAND U8830 ( .A(n6414), .B(\u_a23_core/u_execute/multiply_out[10] ), .Z(
        n6496) );
  NAND U8831 ( .A(n6498), .B(n6499), .Z(\u_a23_core/u_execute/u_multiply/n597 ) );
  AND U8832 ( .A(n6500), .B(n6501), .Z(n6499) );
  NAND U8833 ( .A(n6423), .B(\u_a23_core/u_execute/u_multiply/sum_acc1[11] ), 
        .Z(n6501) );
  NANDN U8834 ( .B(n6502), .A(n6425), .Z(n6500) );
  AND U8835 ( .A(n6503), .B(n6504), .Z(n6498) );
  NANDN U8836 ( .B(n6413), .A(\u_a23_core/u_execute/multiply_out[12] ), .Z(
        n6504) );
  NAND U8837 ( .A(n6414), .B(\u_a23_core/u_execute/multiply_out[11] ), .Z(
        n6503) );
  NAND U8838 ( .A(n6505), .B(n6506), .Z(\u_a23_core/u_execute/u_multiply/n596 ) );
  AND U8839 ( .A(n6507), .B(n6508), .Z(n6506) );
  NAND U8840 ( .A(n6423), .B(\u_a23_core/u_execute/u_multiply/sum_acc1[12] ), 
        .Z(n6508) );
  NANDN U8841 ( .B(n6509), .A(n6425), .Z(n6507) );
  AND U8842 ( .A(n6510), .B(n6511), .Z(n6505) );
  NANDN U8843 ( .B(n6413), .A(\u_a23_core/u_execute/multiply_out[13] ), .Z(
        n6511) );
  NAND U8844 ( .A(n6414), .B(\u_a23_core/u_execute/multiply_out[12] ), .Z(
        n6510) );
  NAND U8845 ( .A(n6512), .B(n6513), .Z(\u_a23_core/u_execute/u_multiply/n595 ) );
  AND U8846 ( .A(n6514), .B(n6515), .Z(n6513) );
  NAND U8847 ( .A(n6423), .B(\u_a23_core/u_execute/u_multiply/sum_acc1[13] ), 
        .Z(n6515) );
  NANDN U8848 ( .B(n6516), .A(n6425), .Z(n6514) );
  AND U8849 ( .A(n6517), .B(n6518), .Z(n6512) );
  NANDN U8850 ( .B(n6413), .A(\u_a23_core/u_execute/multiply_out[14] ), .Z(
        n6518) );
  NAND U8851 ( .A(n6414), .B(\u_a23_core/u_execute/multiply_out[13] ), .Z(
        n6517) );
  NAND U8852 ( .A(n6519), .B(n6520), .Z(\u_a23_core/u_execute/u_multiply/n594 ) );
  AND U8853 ( .A(n6521), .B(n6522), .Z(n6520) );
  NAND U8854 ( .A(n6423), .B(\u_a23_core/u_execute/u_multiply/sum_acc1[14] ), 
        .Z(n6522) );
  NANDN U8855 ( .B(n6523), .A(n6425), .Z(n6521) );
  AND U8856 ( .A(n6524), .B(n6525), .Z(n6519) );
  NANDN U8857 ( .B(n6413), .A(\u_a23_core/u_execute/multiply_out[15] ), .Z(
        n6525) );
  NAND U8858 ( .A(n6414), .B(\u_a23_core/u_execute/multiply_out[14] ), .Z(
        n6524) );
  NAND U8859 ( .A(n6526), .B(n6527), .Z(\u_a23_core/u_execute/u_multiply/n593 ) );
  AND U8860 ( .A(n6528), .B(n6529), .Z(n6527) );
  NAND U8861 ( .A(n6423), .B(\u_a23_core/u_execute/u_multiply/sum_acc1[15] ), 
        .Z(n6529) );
  NANDN U8862 ( .B(n6530), .A(n6425), .Z(n6528) );
  AND U8863 ( .A(n6531), .B(n6532), .Z(n6526) );
  NANDN U8864 ( .B(n6413), .A(\u_a23_core/u_execute/multiply_out[16] ), .Z(
        n6532) );
  NAND U8865 ( .A(n6414), .B(\u_a23_core/u_execute/multiply_out[15] ), .Z(
        n6531) );
  NAND U8866 ( .A(n6533), .B(n6534), .Z(\u_a23_core/u_execute/u_multiply/n592 ) );
  AND U8867 ( .A(n6535), .B(n6536), .Z(n6534) );
  NAND U8868 ( .A(n6423), .B(\u_a23_core/u_execute/u_multiply/sum_acc1[16] ), 
        .Z(n6536) );
  NANDN U8869 ( .B(n6537), .A(n6425), .Z(n6535) );
  AND U8870 ( .A(n6538), .B(n6539), .Z(n6533) );
  NANDN U8871 ( .B(n6413), .A(\u_a23_core/u_execute/multiply_out[17] ), .Z(
        n6539) );
  NAND U8872 ( .A(n6414), .B(\u_a23_core/u_execute/multiply_out[16] ), .Z(
        n6538) );
  NAND U8873 ( .A(n6540), .B(n6541), .Z(\u_a23_core/u_execute/u_multiply/n591 ) );
  AND U8874 ( .A(n6542), .B(n6543), .Z(n6541) );
  NAND U8875 ( .A(n6423), .B(\u_a23_core/u_execute/u_multiply/sum_acc1[17] ), 
        .Z(n6543) );
  NANDN U8876 ( .B(n6544), .A(n6425), .Z(n6542) );
  AND U8877 ( .A(n6545), .B(n6546), .Z(n6540) );
  NANDN U8878 ( .B(n6413), .A(\u_a23_core/u_execute/multiply_out[18] ), .Z(
        n6546) );
  NAND U8879 ( .A(n6414), .B(\u_a23_core/u_execute/multiply_out[17] ), .Z(
        n6545) );
  NAND U8880 ( .A(n6547), .B(n6548), .Z(\u_a23_core/u_execute/u_multiply/n590 ) );
  AND U8881 ( .A(n6549), .B(n6550), .Z(n6548) );
  NAND U8882 ( .A(n6423), .B(\u_a23_core/u_execute/u_multiply/sum_acc1[18] ), 
        .Z(n6550) );
  NANDN U8883 ( .B(n6551), .A(n6425), .Z(n6549) );
  AND U8884 ( .A(n6552), .B(n6553), .Z(n6547) );
  NANDN U8885 ( .B(n6413), .A(\u_a23_core/u_execute/multiply_out[19] ), .Z(
        n6553) );
  NAND U8886 ( .A(n6414), .B(\u_a23_core/u_execute/multiply_out[18] ), .Z(
        n6552) );
  NAND U8887 ( .A(n6554), .B(n6555), .Z(\u_a23_core/u_execute/u_multiply/n589 ) );
  AND U8888 ( .A(n6556), .B(n6557), .Z(n6555) );
  NAND U8889 ( .A(n6423), .B(\u_a23_core/u_execute/u_multiply/sum_acc1[19] ), 
        .Z(n6557) );
  NANDN U8890 ( .B(n6558), .A(n6425), .Z(n6556) );
  AND U8891 ( .A(n6559), .B(n6560), .Z(n6554) );
  NANDN U8892 ( .B(n6413), .A(\u_a23_core/u_execute/multiply_out[20] ), .Z(
        n6560) );
  NAND U8893 ( .A(n6414), .B(\u_a23_core/u_execute/multiply_out[19] ), .Z(
        n6559) );
  NAND U8894 ( .A(n6561), .B(n6562), .Z(\u_a23_core/u_execute/u_multiply/n588 ) );
  AND U8895 ( .A(n6563), .B(n6564), .Z(n6562) );
  NAND U8896 ( .A(n6423), .B(\u_a23_core/u_execute/u_multiply/sum_acc1[20] ), 
        .Z(n6564) );
  NANDN U8897 ( .B(n6565), .A(n6425), .Z(n6563) );
  AND U8898 ( .A(n6566), .B(n6567), .Z(n6561) );
  NANDN U8899 ( .B(n6413), .A(\u_a23_core/u_execute/multiply_out[21] ), .Z(
        n6567) );
  NAND U8900 ( .A(n6414), .B(\u_a23_core/u_execute/multiply_out[20] ), .Z(
        n6566) );
  NAND U8901 ( .A(n6568), .B(n6569), .Z(\u_a23_core/u_execute/u_multiply/n587 ) );
  AND U8902 ( .A(n6570), .B(n6571), .Z(n6569) );
  NAND U8903 ( .A(n6423), .B(\u_a23_core/u_execute/u_multiply/sum_acc1[21] ), 
        .Z(n6571) );
  NANDN U8904 ( .B(n6572), .A(n6425), .Z(n6570) );
  AND U8905 ( .A(n6573), .B(n6574), .Z(n6568) );
  NANDN U8906 ( .B(n6413), .A(\u_a23_core/u_execute/multiply_out[22] ), .Z(
        n6574) );
  NAND U8907 ( .A(n6414), .B(\u_a23_core/u_execute/multiply_out[21] ), .Z(
        n6573) );
  NAND U8908 ( .A(n6575), .B(n6576), .Z(\u_a23_core/u_execute/u_multiply/n586 ) );
  AND U8909 ( .A(n6577), .B(n6578), .Z(n6576) );
  NAND U8910 ( .A(n6423), .B(\u_a23_core/u_execute/u_multiply/sum_acc1[22] ), 
        .Z(n6578) );
  NANDN U8911 ( .B(n6579), .A(n6425), .Z(n6577) );
  AND U8912 ( .A(n6580), .B(n6581), .Z(n6575) );
  NANDN U8913 ( .B(n6413), .A(\u_a23_core/u_execute/multiply_out[23] ), .Z(
        n6581) );
  NAND U8914 ( .A(n6414), .B(\u_a23_core/u_execute/multiply_out[22] ), .Z(
        n6580) );
  NAND U8915 ( .A(n6582), .B(n6583), .Z(\u_a23_core/u_execute/u_multiply/n585 ) );
  AND U8916 ( .A(n6584), .B(n6585), .Z(n6583) );
  NAND U8917 ( .A(n6423), .B(\u_a23_core/u_execute/u_multiply/sum_acc1[23] ), 
        .Z(n6585) );
  NANDN U8918 ( .B(n6586), .A(n6425), .Z(n6584) );
  AND U8919 ( .A(n6587), .B(n6588), .Z(n6582) );
  NANDN U8920 ( .B(n6413), .A(\u_a23_core/u_execute/multiply_out[24] ), .Z(
        n6588) );
  NAND U8921 ( .A(n6414), .B(\u_a23_core/u_execute/multiply_out[23] ), .Z(
        n6587) );
  NAND U8922 ( .A(n6589), .B(n6590), .Z(\u_a23_core/u_execute/u_multiply/n584 ) );
  AND U8923 ( .A(n6591), .B(n6592), .Z(n6590) );
  NAND U8924 ( .A(n6423), .B(\u_a23_core/u_execute/u_multiply/sum_acc1[24] ), 
        .Z(n6592) );
  NANDN U8925 ( .B(n6593), .A(n6425), .Z(n6591) );
  AND U8926 ( .A(n6594), .B(n6595), .Z(n6589) );
  NANDN U8927 ( .B(n6413), .A(\u_a23_core/u_execute/multiply_out[25] ), .Z(
        n6595) );
  NAND U8928 ( .A(n6414), .B(\u_a23_core/u_execute/multiply_out[24] ), .Z(
        n6594) );
  NAND U8929 ( .A(n6596), .B(n6597), .Z(\u_a23_core/u_execute/u_multiply/n583 ) );
  AND U8930 ( .A(n6598), .B(n6599), .Z(n6597) );
  NAND U8931 ( .A(n6423), .B(\u_a23_core/u_execute/u_multiply/sum_acc1[25] ), 
        .Z(n6599) );
  NANDN U8932 ( .B(n6600), .A(n6425), .Z(n6598) );
  AND U8933 ( .A(n6601), .B(n6602), .Z(n6596) );
  NANDN U8934 ( .B(n6413), .A(\u_a23_core/u_execute/multiply_out[26] ), .Z(
        n6602) );
  NAND U8935 ( .A(n6414), .B(\u_a23_core/u_execute/multiply_out[25] ), .Z(
        n6601) );
  NAND U8936 ( .A(n6603), .B(n6604), .Z(\u_a23_core/u_execute/u_multiply/n582 ) );
  AND U8937 ( .A(n6605), .B(n6606), .Z(n6604) );
  NAND U8938 ( .A(n6423), .B(\u_a23_core/u_execute/u_multiply/sum_acc1[26] ), 
        .Z(n6606) );
  NANDN U8939 ( .B(n6607), .A(n6425), .Z(n6605) );
  AND U8940 ( .A(n6608), .B(n6609), .Z(n6603) );
  NANDN U8941 ( .B(n6413), .A(\u_a23_core/u_execute/multiply_out[27] ), .Z(
        n6609) );
  NAND U8942 ( .A(n6414), .B(\u_a23_core/u_execute/multiply_out[26] ), .Z(
        n6608) );
  NAND U8943 ( .A(n6610), .B(n6611), .Z(\u_a23_core/u_execute/u_multiply/n581 ) );
  AND U8944 ( .A(n6612), .B(n6613), .Z(n6611) );
  NAND U8945 ( .A(n6423), .B(\u_a23_core/u_execute/u_multiply/sum_acc1[27] ), 
        .Z(n6613) );
  NANDN U8946 ( .B(n6614), .A(n6425), .Z(n6612) );
  AND U8947 ( .A(n6615), .B(n6616), .Z(n6610) );
  NANDN U8948 ( .B(n6413), .A(\u_a23_core/u_execute/multiply_out[28] ), .Z(
        n6616) );
  NAND U8949 ( .A(n6414), .B(\u_a23_core/u_execute/multiply_out[27] ), .Z(
        n6615) );
  NAND U8950 ( .A(n6617), .B(n6618), .Z(\u_a23_core/u_execute/u_multiply/n580 ) );
  AND U8951 ( .A(n6619), .B(n6620), .Z(n6618) );
  NAND U8952 ( .A(n6423), .B(\u_a23_core/u_execute/u_multiply/sum_acc1[28] ), 
        .Z(n6620) );
  NANDN U8953 ( .B(n6621), .A(n6425), .Z(n6619) );
  AND U8954 ( .A(n6622), .B(n6623), .Z(n6617) );
  NANDN U8955 ( .B(n6413), .A(\u_a23_core/u_execute/multiply_out[29] ), .Z(
        n6623) );
  NAND U8956 ( .A(n6414), .B(\u_a23_core/u_execute/multiply_out[28] ), .Z(
        n6622) );
  NAND U8957 ( .A(n6624), .B(n6625), .Z(\u_a23_core/u_execute/u_multiply/n579 ) );
  AND U8958 ( .A(n6626), .B(n6627), .Z(n6625) );
  NAND U8959 ( .A(n6423), .B(\u_a23_core/u_execute/u_multiply/sum_acc1[29] ), 
        .Z(n6627) );
  NANDN U8960 ( .B(n6628), .A(n6425), .Z(n6626) );
  AND U8961 ( .A(n6629), .B(n6630), .Z(n6624) );
  NANDN U8962 ( .B(n6413), .A(\u_a23_core/u_execute/multiply_out[30] ), .Z(
        n6630) );
  NAND U8963 ( .A(n6414), .B(\u_a23_core/u_execute/multiply_out[29] ), .Z(
        n6629) );
  NAND U8964 ( .A(n6631), .B(n6632), .Z(\u_a23_core/u_execute/u_multiply/n578 ) );
  AND U8965 ( .A(n6633), .B(n6634), .Z(n6632) );
  NAND U8966 ( .A(n6423), .B(\u_a23_core/u_execute/u_multiply/sum_acc1[30] ), 
        .Z(n6634) );
  NANDN U8967 ( .B(n6635), .A(n6425), .Z(n6633) );
  AND U8968 ( .A(n6636), .B(n6637), .Z(n6631) );
  NANDN U8969 ( .B(n6413), .A(\u_a23_core/u_execute/multiply_out[31] ), .Z(
        n6637) );
  NAND U8970 ( .A(n6414), .B(\u_a23_core/u_execute/multiply_out[30] ), .Z(
        n6636) );
  NAND U8971 ( .A(n6638), .B(n6639), .Z(\u_a23_core/u_execute/u_multiply/n577 ) );
  AND U8972 ( .A(n6640), .B(n6641), .Z(n6639) );
  NAND U8973 ( .A(n6423), .B(\u_a23_core/u_execute/u_multiply/sum_acc1[31] ), 
        .Z(n6641) );
  NOR U8974 ( .A(n6414), .B(n6642), .Z(n6423) );
  NANDN U8975 ( .B(n6643), .A(n6425), .Z(n6640) );
  ANDN U8976 ( .A(n6644), .B(n6645), .Z(n6425) );
  AND U8977 ( .A(n6646), .B(n6647), .Z(n6638) );
  NANDN U8978 ( .B(n6413), .A(\u_a23_core/u_execute/u_multiply/product[33] ), 
        .Z(n6647) );
  NAND U8979 ( .A(\u_a23_core/u_execute/multiply_out[31] ), .B(n6414), .Z(
        n6646) );
  NAND U8980 ( .A(n6648), .B(n6649), .Z(\u_a23_core/u_execute/u_multiply/n576 ) );
  NAND U8981 ( .A(n6417), .B(\u_a23_core/u_execute/u_multiply/sum[1] ), .Z(
        n6649) );
  NAND U8982 ( .A(n6418), .B(\u_a23_core/u_execute/u_multiply/product[34] ), 
        .Z(n6648) );
  NAND U8983 ( .A(n6650), .B(n6651), .Z(\u_a23_core/u_execute/u_multiply/n575 ) );
  NAND U8984 ( .A(n6417), .B(\u_a23_core/u_execute/u_multiply/sum[2] ), .Z(
        n6651) );
  NAND U8985 ( .A(n6418), .B(\u_a23_core/u_execute/u_multiply/product[35] ), 
        .Z(n6650) );
  NAND U8986 ( .A(n6652), .B(n6653), .Z(\u_a23_core/u_execute/u_multiply/n574 ) );
  NAND U8987 ( .A(n6417), .B(\u_a23_core/u_execute/u_multiply/sum[3] ), .Z(
        n6653) );
  NAND U8988 ( .A(n6418), .B(\u_a23_core/u_execute/u_multiply/product[36] ), 
        .Z(n6652) );
  NAND U8989 ( .A(n6654), .B(n6655), .Z(\u_a23_core/u_execute/u_multiply/n573 ) );
  NAND U8990 ( .A(n6417), .B(\u_a23_core/u_execute/u_multiply/sum[4] ), .Z(
        n6655) );
  NAND U8991 ( .A(n6418), .B(\u_a23_core/u_execute/u_multiply/product[37] ), 
        .Z(n6654) );
  NAND U8992 ( .A(n6656), .B(n6657), .Z(\u_a23_core/u_execute/u_multiply/n572 ) );
  NAND U8993 ( .A(n6417), .B(\u_a23_core/u_execute/u_multiply/sum[5] ), .Z(
        n6657) );
  NAND U8994 ( .A(n6418), .B(\u_a23_core/u_execute/u_multiply/product[38] ), 
        .Z(n6656) );
  NAND U8995 ( .A(n6658), .B(n6659), .Z(\u_a23_core/u_execute/u_multiply/n571 ) );
  NAND U8996 ( .A(n6417), .B(\u_a23_core/u_execute/u_multiply/sum[6] ), .Z(
        n6659) );
  NAND U8997 ( .A(n6418), .B(\u_a23_core/u_execute/u_multiply/product[39] ), 
        .Z(n6658) );
  NAND U8998 ( .A(n6660), .B(n6661), .Z(\u_a23_core/u_execute/u_multiply/n570 ) );
  NAND U8999 ( .A(n6417), .B(\u_a23_core/u_execute/u_multiply/sum[7] ), .Z(
        n6661) );
  NAND U9000 ( .A(n6418), .B(\u_a23_core/u_execute/u_multiply/product[40] ), 
        .Z(n6660) );
  NAND U9001 ( .A(n6662), .B(n6663), .Z(\u_a23_core/u_execute/u_multiply/n569 ) );
  NAND U9002 ( .A(n6417), .B(\u_a23_core/u_execute/u_multiply/sum[8] ), .Z(
        n6663) );
  NAND U9003 ( .A(n6418), .B(\u_a23_core/u_execute/u_multiply/product[41] ), 
        .Z(n6662) );
  NAND U9004 ( .A(n6664), .B(n6665), .Z(\u_a23_core/u_execute/u_multiply/n568 ) );
  NAND U9005 ( .A(n6417), .B(\u_a23_core/u_execute/u_multiply/sum[9] ), .Z(
        n6665) );
  NAND U9006 ( .A(n6418), .B(\u_a23_core/u_execute/u_multiply/product[42] ), 
        .Z(n6664) );
  NAND U9007 ( .A(n6666), .B(n6667), .Z(\u_a23_core/u_execute/u_multiply/n567 ) );
  NAND U9008 ( .A(n6417), .B(\u_a23_core/u_execute/u_multiply/sum[10] ), .Z(
        n6667) );
  NAND U9009 ( .A(n6418), .B(\u_a23_core/u_execute/u_multiply/product[43] ), 
        .Z(n6666) );
  NAND U9010 ( .A(n6668), .B(n6669), .Z(\u_a23_core/u_execute/u_multiply/n566 ) );
  NAND U9011 ( .A(n6417), .B(\u_a23_core/u_execute/u_multiply/sum[11] ), .Z(
        n6669) );
  NAND U9012 ( .A(n6418), .B(\u_a23_core/u_execute/u_multiply/product[44] ), 
        .Z(n6668) );
  NAND U9013 ( .A(n6670), .B(n6671), .Z(\u_a23_core/u_execute/u_multiply/n565 ) );
  NAND U9014 ( .A(n6417), .B(\u_a23_core/u_execute/u_multiply/sum[12] ), .Z(
        n6671) );
  NAND U9015 ( .A(n6418), .B(\u_a23_core/u_execute/u_multiply/product[45] ), 
        .Z(n6670) );
  NAND U9016 ( .A(n6672), .B(n6673), .Z(\u_a23_core/u_execute/u_multiply/n564 ) );
  NAND U9017 ( .A(n6417), .B(\u_a23_core/u_execute/u_multiply/sum[13] ), .Z(
        n6673) );
  NAND U9018 ( .A(n6418), .B(\u_a23_core/u_execute/u_multiply/product[46] ), 
        .Z(n6672) );
  NAND U9019 ( .A(n6674), .B(n6675), .Z(\u_a23_core/u_execute/u_multiply/n563 ) );
  NAND U9020 ( .A(n6417), .B(\u_a23_core/u_execute/u_multiply/sum[14] ), .Z(
        n6675) );
  NAND U9021 ( .A(n6418), .B(\u_a23_core/u_execute/u_multiply/product[47] ), 
        .Z(n6674) );
  NAND U9022 ( .A(n6676), .B(n6677), .Z(\u_a23_core/u_execute/u_multiply/n562 ) );
  NAND U9023 ( .A(n6417), .B(\u_a23_core/u_execute/u_multiply/sum[15] ), .Z(
        n6677) );
  NAND U9024 ( .A(n6418), .B(\u_a23_core/u_execute/u_multiply/product[48] ), 
        .Z(n6676) );
  NAND U9025 ( .A(n6678), .B(n6679), .Z(\u_a23_core/u_execute/u_multiply/n561 ) );
  NAND U9026 ( .A(n6417), .B(\u_a23_core/u_execute/u_multiply/sum[16] ), .Z(
        n6679) );
  NAND U9027 ( .A(n6418), .B(\u_a23_core/u_execute/u_multiply/product[49] ), 
        .Z(n6678) );
  NAND U9028 ( .A(n6680), .B(n6681), .Z(\u_a23_core/u_execute/u_multiply/n560 ) );
  NAND U9029 ( .A(n6417), .B(\u_a23_core/u_execute/u_multiply/sum[17] ), .Z(
        n6681) );
  NAND U9030 ( .A(n6418), .B(\u_a23_core/u_execute/u_multiply/product[50] ), 
        .Z(n6680) );
  NAND U9031 ( .A(n6682), .B(n6683), .Z(\u_a23_core/u_execute/u_multiply/n559 ) );
  NAND U9032 ( .A(n6417), .B(\u_a23_core/u_execute/u_multiply/sum[18] ), .Z(
        n6683) );
  NAND U9033 ( .A(n6418), .B(\u_a23_core/u_execute/u_multiply/product[51] ), 
        .Z(n6682) );
  NAND U9034 ( .A(n6684), .B(n6685), .Z(\u_a23_core/u_execute/u_multiply/n558 ) );
  NAND U9035 ( .A(n6417), .B(\u_a23_core/u_execute/u_multiply/sum[19] ), .Z(
        n6685) );
  NAND U9036 ( .A(n6418), .B(\u_a23_core/u_execute/u_multiply/product[52] ), 
        .Z(n6684) );
  NAND U9037 ( .A(n6686), .B(n6687), .Z(\u_a23_core/u_execute/u_multiply/n557 ) );
  NAND U9038 ( .A(n6417), .B(\u_a23_core/u_execute/u_multiply/sum[20] ), .Z(
        n6687) );
  NAND U9039 ( .A(n6418), .B(\u_a23_core/u_execute/u_multiply/product[53] ), 
        .Z(n6686) );
  NAND U9040 ( .A(n6688), .B(n6689), .Z(\u_a23_core/u_execute/u_multiply/n556 ) );
  NAND U9041 ( .A(n6417), .B(\u_a23_core/u_execute/u_multiply/sum[21] ), .Z(
        n6689) );
  NAND U9042 ( .A(n6418), .B(\u_a23_core/u_execute/u_multiply/product[54] ), 
        .Z(n6688) );
  NAND U9043 ( .A(n6690), .B(n6691), .Z(\u_a23_core/u_execute/u_multiply/n555 ) );
  NAND U9044 ( .A(n6417), .B(\u_a23_core/u_execute/u_multiply/sum[22] ), .Z(
        n6691) );
  NAND U9045 ( .A(n6418), .B(\u_a23_core/u_execute/u_multiply/product[55] ), 
        .Z(n6690) );
  NAND U9046 ( .A(n6692), .B(n6693), .Z(\u_a23_core/u_execute/u_multiply/n554 ) );
  NAND U9047 ( .A(n6417), .B(\u_a23_core/u_execute/u_multiply/sum[23] ), .Z(
        n6693) );
  NAND U9048 ( .A(n6418), .B(\u_a23_core/u_execute/u_multiply/product[56] ), 
        .Z(n6692) );
  NAND U9049 ( .A(n6694), .B(n6695), .Z(\u_a23_core/u_execute/u_multiply/n553 ) );
  NAND U9050 ( .A(n6417), .B(\u_a23_core/u_execute/u_multiply/sum[24] ), .Z(
        n6695) );
  NAND U9051 ( .A(n6418), .B(\u_a23_core/u_execute/u_multiply/product[57] ), 
        .Z(n6694) );
  NAND U9052 ( .A(n6696), .B(n6697), .Z(\u_a23_core/u_execute/u_multiply/n552 ) );
  NAND U9053 ( .A(n6417), .B(\u_a23_core/u_execute/u_multiply/sum[25] ), .Z(
        n6697) );
  NAND U9054 ( .A(n6418), .B(\u_a23_core/u_execute/u_multiply/product[58] ), 
        .Z(n6696) );
  NAND U9055 ( .A(n6698), .B(n6699), .Z(\u_a23_core/u_execute/u_multiply/n551 ) );
  NAND U9056 ( .A(n6417), .B(\u_a23_core/u_execute/u_multiply/sum[26] ), .Z(
        n6699) );
  NAND U9057 ( .A(n6418), .B(\u_a23_core/u_execute/u_multiply/product[59] ), 
        .Z(n6698) );
  NAND U9058 ( .A(n6700), .B(n6701), .Z(\u_a23_core/u_execute/u_multiply/n550 ) );
  NAND U9059 ( .A(n6417), .B(\u_a23_core/u_execute/u_multiply/sum[27] ), .Z(
        n6701) );
  NAND U9060 ( .A(n6418), .B(\u_a23_core/u_execute/u_multiply/product[60] ), 
        .Z(n6700) );
  NAND U9061 ( .A(n6702), .B(n6703), .Z(\u_a23_core/u_execute/u_multiply/n549 ) );
  NAND U9062 ( .A(n6417), .B(\u_a23_core/u_execute/u_multiply/sum[28] ), .Z(
        n6703) );
  NAND U9063 ( .A(n6418), .B(\u_a23_core/u_execute/u_multiply/product[61] ), 
        .Z(n6702) );
  NAND U9064 ( .A(n6704), .B(n6705), .Z(\u_a23_core/u_execute/u_multiply/n548 ) );
  NAND U9065 ( .A(n6417), .B(\u_a23_core/u_execute/u_multiply/sum[29] ), .Z(
        n6705) );
  NAND U9066 ( .A(n6418), .B(\u_a23_core/u_execute/u_multiply/product[62] ), 
        .Z(n6704) );
  NAND U9067 ( .A(n6706), .B(n6707), .Z(\u_a23_core/u_execute/u_multiply/n547 ) );
  NAND U9068 ( .A(n6417), .B(\u_a23_core/u_execute/u_multiply/sum[30] ), .Z(
        n6707) );
  NAND U9069 ( .A(n6418), .B(\u_a23_core/u_execute/u_multiply/product[63] ), 
        .Z(n6706) );
  NAND U9070 ( .A(n6708), .B(n6709), .Z(\u_a23_core/u_execute/u_multiply/n546 ) );
  NAND U9071 ( .A(n6417), .B(\u_a23_core/u_execute/u_multiply/sum[31] ), .Z(
        n6709) );
  NOR U9072 ( .A(n6710), .B(n6418), .Z(n6417) );
  NAND U9073 ( .A(n6418), .B(\u_a23_core/u_execute/u_multiply/product[64] ), 
        .Z(n6708) );
  NAND U9074 ( .A(n6711), .B(n6712), .Z(\u_a23_core/u_execute/u_multiply/n545 ) );
  NANDN U9075 ( .B(n6413), .A(\u_a23_core/u_execute/u_multiply/sum[32] ), .Z(
        n6712) );
  NAND U9076 ( .A(n6414), .B(\u_a23_core/u_execute/u_multiply/product[65] ), 
        .Z(n6711) );
  NAND U9077 ( .A(n6713), .B(n6714), .Z(\u_a23_core/u_execute/u_multiply/n544 ) );
  NAND U9078 ( .A(n6414), .B(\u_a23_core/u_execute/u_multiply/product[66] ), 
        .Z(n6713) );
  NAND U9079 ( .A(n6715), .B(n6714), .Z(\u_a23_core/u_execute/u_multiply/n543 ) );
  NANDN U9080 ( .B(n6413), .A(\u_a23_core/u_execute/u_multiply/sum[33] ), .Z(
        n6714) );
  NAND U9081 ( .A(n6716), .B(n6642), .Z(n6413) );
  AND U9082 ( .A(n6644), .B(n6645), .Z(n6716) );
  IV U9083 ( .A(n6710), .Z(n6645) );
  IV U9084 ( .A(n6414), .Z(n6644) );
  NAND U9085 ( .A(n6414), .B(\u_a23_core/u_execute/u_multiply/product[67] ), 
        .Z(n6715) );
  AND U9086 ( .A(n6717), .B(n6418), .Z(n6414) );
  NANDN U9087 ( .B(n6718), .A(n6719), .Z(n6418) );
  AND U9088 ( .A(n6642), .B(n5930), .Z(n6719) );
  NAND U9089 ( .A(n6720), .B(\u_a23_core/u_execute/u_multiply/count[5] ), .Z(
        n6642) );
  NAND U9090 ( .A(n6721), .B(n6722), .Z(n6720) );
  NAND U9091 ( .A(n6723), .B(n6724), .Z(n6717) );
  AND U9092 ( .A(n6725), .B(\u_a23_core/multiply_function[1] ), .Z(n6724) );
  AND U9093 ( .A(n6408), .B(n5930), .Z(n6725) );
  AND U9094 ( .A(n6722), .B(\u_a23_core/multiply_function[0] ), .Z(n6723) );
  IV U9095 ( .A(n6726), .Z(\u_a23_core/u_execute/u_multiply/n509 ) );
  MUX U9096 ( .IN0(n6721), .IN1(n6727), .SEL(\u_a23_core/multiply_function[0] ), .F(n6726) );
  NAND U9097 ( .A(n6728), .B(\u_a23_core/u_execute/u_multiply/N55 ), .Z(n6727)
         );
  AND U9098 ( .A(n6728), .B(n6729), .Z(\u_a23_core/u_execute/u_multiply/n507 )
         );
  MUX U9099 ( .IN0(\u_a23_core/u_execute/u_multiply/N56 ), .IN1(
        \u_a23_core/u_execute/u_multiply/count[2] ), .SEL(n6718), .F(n6729) );
  AND U9100 ( .A(n6728), .B(n6730), .Z(\u_a23_core/u_execute/u_multiply/n505 )
         );
  MUX U9101 ( .IN0(\u_a23_core/u_execute/u_multiply/N57 ), .IN1(
        \u_a23_core/u_execute/u_multiply/count[3] ), .SEL(n6718), .F(n6730) );
  AND U9102 ( .A(n6728), .B(n6731), .Z(\u_a23_core/u_execute/u_multiply/n503 )
         );
  MUX U9103 ( .IN0(\u_a23_core/u_execute/u_multiply/N58 ), .IN1(
        \u_a23_core/u_execute/u_multiply/count[4] ), .SEL(n6718), .F(n6731) );
  IV U9104 ( .A(\u_a23_core/multiply_function[0] ), .Z(n6718) );
  ANDN U9105 ( .A(n6410), .B(n6710), .Z(n6728) );
  ANDN U9106 ( .A(n6732), .B(\u_a23_core/u_execute/u_multiply/count[5] ), .Z(
        n6710) );
  NAND U9107 ( .A(n6733), .B(n6734), .Z(n6410) );
  ANDN U9108 ( .A(n6722), .B(n6735), .Z(n6734) );
  AND U9109 ( .A(\u_a23_core/u_execute/u_multiply/count[5] ), .B(
        \u_a23_core/u_execute/u_multiply/count[1] ), .Z(n6733) );
  MUX U9110 ( .IN0(n6736), .IN1(n6737), .SEL(
        \u_a23_core/u_execute/u_multiply/count[5] ), .F(
        \u_a23_core/u_execute/u_multiply/n501 ) );
  NAND U9111 ( .A(\u_a23_core/multiply_function[0] ), .B(n6738), .Z(n6737) );
  AND U9112 ( .A(n6739), .B(n6740), .Z(n6738) );
  NANDN U9113 ( .B(\u_a23_core/u_execute/u_multiply/add_139/carry[5] ), .A(
        n6741), .Z(n6740) );
  NANDN U9114 ( .B(n6735), .A(\u_a23_core/u_execute/u_multiply/count[1] ), .Z(
        n6741) );
  XOR U9115 ( .A(n6742), .B(n6408), .Z(n6735) );
  OR U9116 ( .A(n6722), .B(\u_a23_core/u_execute/u_multiply/add_139/carry[5] ), 
        .Z(n6739) );
  AND U9117 ( .A(n6743), .B(\u_a23_core/multiply_function[0] ), .Z(n6736) );
  ANDN U9118 ( .A(\u_a23_core/u_execute/u_multiply/add_139/carry[5] ), .B(
        n6732), .Z(n6743) );
  AND U9119 ( .A(n6744), .B(n6722), .Z(n6732) );
  ANDN U9120 ( .A(n6745), .B(\u_a23_core/u_execute/u_multiply/count[2] ), .Z(
        n6722) );
  NOR U9121 ( .A(\u_a23_core/u_execute/u_multiply/count[3] ), .B(
        \u_a23_core/u_execute/u_multiply/count[4] ), .Z(n6745) );
  AND U9122 ( .A(n6408), .B(n6721), .Z(n6744) );
  IV U9123 ( .A(\u_a23_core/u_execute/u_multiply/count[1] ), .Z(n6721) );
  IV U9124 ( .A(\u_a23_core/u_execute/u_multiply/count[0] ), .Z(n6408) );
  IV U9125 ( .A(n6746), .Z(\u_a23_core/u_execute/u_multiply/n499 ) );
  MUX U9126 ( .IN0(n6747), .IN1(n6748), .SEL(\u_a23_core/multiply_function[0] ), .F(n6746) );
  NAND U9127 ( .A(n6749), .B(n6750), .Z(n6748) );
  AND U9128 ( .A(n6751), .B(\u_a23_core/u_execute/u_multiply/count[1] ), .Z(
        n6750) );
  ANDN U9129 ( .A(\u_a23_core/u_execute/u_multiply/count[0] ), .B(
        \u_a23_core/u_execute/u_multiply/count[5] ), .Z(n6751) );
  AND U9130 ( .A(\u_a23_core/u_execute/u_multiply/count[4] ), .B(n6752), .Z(
        n6749) );
  AND U9131 ( .A(\u_a23_core/u_execute/u_multiply/count[2] ), .B(
        \u_a23_core/u_execute/u_multiply/count[3] ), .Z(n6752) );
  MUX U9132 ( .IN0(\u_a23_core/alu_function[5] ), .IN1(
        \u_a23_core/u_execute/save_int_pc_m4[29] ), .SEL(
        \u_a23_core/alu_function[6] ), .F(
        \u_a23_core/u_execute/u_alu/carry_in ) );
  IV U9133 ( .A(n16632), .Z(\u_a23_core/u_execute/rs[7] ) );
  IV U9134 ( .A(n16631), .Z(\u_a23_core/u_execute/rs[6] ) );
  IV U9135 ( .A(n16630), .Z(\u_a23_core/u_execute/rs[5] ) );
  NAND U9136 ( .A(n6753), .B(n6754), .Z(\u_a23_core/u_execute/n1076 ) );
  NAND U9137 ( .A(n6755), .B(n6756), .Z(n6754) );
  NAND U9138 ( .A(n6757), .B(n6758), .Z(n6755) );
  NAND U9139 ( .A(n6759), .B(n6760), .Z(n6758) );
  MUX U9140 ( .IN0(n6761), .IN1(n6762), .SEL(
        \u_a23_core/u_execute/u_alu/fadder_out[31] ), .F(n6760) );
  AND U9141 ( .A(n6763), .B(n6764), .Z(n6762) );
  AND U9142 ( .A(\u_a23_core/u_execute/u_alu/b_not[31] ), .B(
        \u_a23_core/u_execute/u_alu/a[31] ), .Z(n6761) );
  ANDN U9143 ( .A(n6765), .B(\u_a23_core/status_bits_sel[0] ), .Z(n6759) );
  NAND U9144 ( .A(\u_a23_core/u_execute/alu_out[28] ), .B(n6766), .Z(n6757) );
  NAND U9145 ( .A(\u_a23_core/u_execute/save_int_pc_m4[28] ), .B(n6767), .Z(
        n6753) );
  NANDN U9146 ( .B(\u_a23_core/status_bits_sel[2] ), .A(n6756), .Z(n6767) );
  MUX U9147 ( .IN0(\u_a23_core/u_execute/save_int_pc_m4[29] ), .IN1(n6768), 
        .SEL(n6756), .F(\u_a23_core/u_execute/n1075 ) );
  NOR U9148 ( .A(n6769), .B(n6770), .Z(n6756) );
  NAND U9149 ( .A(n6771), .B(n6772), .Z(n6768) );
  NAND U9150 ( .A(n6773), .B(n6774), .Z(n6772) );
  MUX U9151 ( .IN0(\u_a23_core/u_execute/u_alu/fadder_out[32] ), .IN1(n6775), 
        .SEL(\u_a23_core/alu_function[4] ), .F(n6773) );
  MUX U9152 ( .IN0(n6776), .IN1(n6777), .SEL(n6778), .F(n6775) );
  MUX U9153 ( .IN0(\u_a23_core/imm32[31] ), .IN1(
        \u_a23_core/u_execute/save_int_pc_m4[29] ), .SEL(n6779), .F(n6777) );
  AND U9154 ( .A(n6780), .B(n6781), .Z(n6779) );
  NOR U9155 ( .A(\u_a23_core/imm_shift_amount[3] ), .B(
        \u_a23_core/imm_shift_amount[4] ), .Z(n6781) );
  NOR U9156 ( .A(\u_a23_core/imm_shift_amount[1] ), .B(
        \u_a23_core/imm_shift_amount[2] ), .Z(n6780) );
  NAND U9157 ( .A(n6782), .B(n6783), .Z(n6776) );
  AND U9158 ( .A(n6784), .B(n6785), .Z(n6783) );
  NAND U9159 ( .A(n6786), .B(n6787), .Z(n6785) );
  NAND U9160 ( .A(n6788), .B(n6789), .Z(n6787) );
  AND U9161 ( .A(n6790), .B(n6791), .Z(n6789) );
  AND U9162 ( .A(n6792), .B(n6793), .Z(n6791) );
  AND U9163 ( .A(n6794), .B(n6795), .Z(n6793) );
  AND U9164 ( .A(n6796), .B(n6797), .Z(n6795) );
  NAND U9165 ( .A(n6798), .B(n6799), .Z(n6797) );
  AND U9166 ( .A(n6800), .B(n6801), .Z(n6796) );
  NAND U9167 ( .A(n6802), .B(n6803), .Z(n6801) );
  AND U9168 ( .A(n6804), .B(n6805), .Z(n6794) );
  NAND U9169 ( .A(n6806), .B(n6807), .Z(n6805) );
  NAND U9170 ( .A(n6808), .B(n6809), .Z(n6804) );
  AND U9171 ( .A(n6810), .B(n6811), .Z(n6792) );
  AND U9172 ( .A(n6812), .B(n6813), .Z(n6811) );
  AND U9173 ( .A(n6814), .B(n6815), .Z(n6810) );
  AND U9174 ( .A(n6816), .B(n6817), .Z(n6790) );
  AND U9175 ( .A(n6818), .B(n6819), .Z(n6817) );
  AND U9176 ( .A(n6820), .B(n6821), .Z(n6819) );
  NAND U9177 ( .A(n6822), .B(n6823), .Z(n6821) );
  AND U9178 ( .A(n6824), .B(n6825), .Z(n6818) );
  NAND U9179 ( .A(n6826), .B(n6827), .Z(n6824) );
  AND U9180 ( .A(n6828), .B(n6829), .Z(n6816) );
  AND U9181 ( .A(n6830), .B(n6831), .Z(n6829) );
  NAND U9182 ( .A(n6832), .B(n6833), .Z(n6831) );
  NAND U9183 ( .A(n6834), .B(n6835), .Z(n6830) );
  AND U9184 ( .A(n6836), .B(n6837), .Z(n6828) );
  NAND U9185 ( .A(n6838), .B(n6839), .Z(n6837) );
  NAND U9186 ( .A(n6840), .B(n6841), .Z(n6836) );
  AND U9187 ( .A(n6842), .B(n6843), .Z(n6788) );
  AND U9188 ( .A(n6844), .B(n6845), .Z(n6843) );
  AND U9189 ( .A(n6846), .B(n6847), .Z(n6845) );
  AND U9190 ( .A(n6848), .B(n6849), .Z(n6847) );
  NAND U9191 ( .A(n6850), .B(n6851), .Z(n6849) );
  NAND U9192 ( .A(n6852), .B(n6853), .Z(n6848) );
  AND U9193 ( .A(n6854), .B(n6855), .Z(n6846) );
  NAND U9194 ( .A(n6856), .B(n6857), .Z(n6855) );
  NAND U9195 ( .A(n6858), .B(n6859), .Z(n6854) );
  AND U9196 ( .A(n6860), .B(n6861), .Z(n6844) );
  AND U9197 ( .A(n6862), .B(n6863), .Z(n6861) );
  NAND U9198 ( .A(n6864), .B(n6865), .Z(n6863) );
  AND U9199 ( .A(n6866), .B(n6867), .Z(n6860) );
  AND U9200 ( .A(n6868), .B(n6869), .Z(n6842) );
  AND U9201 ( .A(n6870), .B(n6871), .Z(n6869) );
  AND U9202 ( .A(n6872), .B(n6873), .Z(n6871) );
  AND U9203 ( .A(n6874), .B(n6875), .Z(n6870) );
  AND U9204 ( .A(n6876), .B(n6877), .Z(n6868) );
  AND U9205 ( .A(n6878), .B(n6879), .Z(n6877) );
  AND U9206 ( .A(n6880), .B(n6881), .Z(n6876) );
  NAND U9207 ( .A(\u_a23_core/shift_imm_zero ), .B(n6882), .Z(n6880) );
  AND U9208 ( .A(n6883), .B(n6884), .Z(n6784) );
  NAND U9209 ( .A(n6885), .B(n6886), .Z(n6884) );
  NAND U9210 ( .A(n6887), .B(n6888), .Z(n6883) );
  NAND U9211 ( .A(n6889), .B(n6890), .Z(n6887) );
  AND U9212 ( .A(n6800), .B(n6891), .Z(n6890) );
  NANDN U9213 ( .B(n6892), .A(n6882), .Z(n6891) );
  NAND U9214 ( .A(n6893), .B(n6894), .Z(n6800) );
  ANDN U9215 ( .A(n6895), .B(n6896), .Z(n6889) );
  NAND U9216 ( .A(n6897), .B(n6898), .Z(n6895) );
  AND U9217 ( .A(n6899), .B(n6900), .Z(n6782) );
  NAND U9218 ( .A(n6901), .B(n6902), .Z(n6900) );
  NAND U9219 ( .A(n6903), .B(n6904), .Z(n6901) );
  AND U9220 ( .A(n6905), .B(n6906), .Z(n6904) );
  AND U9221 ( .A(n6907), .B(n6908), .Z(n6906) );
  AND U9222 ( .A(n6909), .B(n6910), .Z(n6908) );
  AND U9223 ( .A(n6911), .B(n6912), .Z(n6910) );
  NANDN U9224 ( .B(n6913), .A(n6898), .Z(n6912) );
  ANDN U9225 ( .A(n6914), .B(n6915), .Z(n6911) );
  NAND U9226 ( .A(n6894), .B(n6916), .Z(n6914) );
  AND U9227 ( .A(n6917), .B(n6918), .Z(n6909) );
  NAND U9228 ( .A(n6802), .B(n6919), .Z(n6918) );
  NAND U9229 ( .A(n6920), .B(n6798), .Z(n6917) );
  AND U9230 ( .A(n6921), .B(n6922), .Z(n6907) );
  AND U9231 ( .A(n6923), .B(n6924), .Z(n6922) );
  NAND U9232 ( .A(n6806), .B(n6925), .Z(n6924) );
  NAND U9233 ( .A(n6808), .B(n6926), .Z(n6923) );
  AND U9234 ( .A(n6927), .B(n6928), .Z(n6921) );
  AND U9235 ( .A(n6929), .B(n6930), .Z(n6905) );
  AND U9236 ( .A(n6931), .B(n6932), .Z(n6930) );
  AND U9237 ( .A(n6933), .B(n6934), .Z(n6932) );
  AND U9238 ( .A(n6935), .B(n6936), .Z(n6931) );
  NAND U9239 ( .A(n6937), .B(n6822), .Z(n6936) );
  AND U9240 ( .A(n6938), .B(n6939), .Z(n6929) );
  AND U9241 ( .A(n6940), .B(n6941), .Z(n6939) );
  NAND U9242 ( .A(n6942), .B(n6826), .Z(n6941) );
  NAND U9243 ( .A(n6832), .B(n6943), .Z(n6940) );
  AND U9244 ( .A(n6944), .B(n6945), .Z(n6938) );
  NAND U9245 ( .A(n6834), .B(n6946), .Z(n6945) );
  NAND U9246 ( .A(n6838), .B(n6947), .Z(n6944) );
  AND U9247 ( .A(n6948), .B(n6949), .Z(n6903) );
  AND U9248 ( .A(n6950), .B(n6951), .Z(n6949) );
  AND U9249 ( .A(n6952), .B(n6953), .Z(n6951) );
  AND U9250 ( .A(n6954), .B(n6955), .Z(n6953) );
  NAND U9251 ( .A(n6956), .B(n6840), .Z(n6955) );
  NAND U9252 ( .A(n6957), .B(n6851), .Z(n6954) );
  AND U9253 ( .A(n6958), .B(n6959), .Z(n6952) );
  NAND U9254 ( .A(n6852), .B(n6960), .Z(n6959) );
  NAND U9255 ( .A(n6961), .B(n6856), .Z(n6958) );
  AND U9256 ( .A(n6962), .B(n6963), .Z(n6950) );
  AND U9257 ( .A(n6964), .B(n6965), .Z(n6963) );
  NAND U9258 ( .A(n6966), .B(n6858), .Z(n6965) );
  NAND U9259 ( .A(n6967), .B(n6864), .Z(n6964) );
  AND U9260 ( .A(n6968), .B(n6969), .Z(n6962) );
  AND U9261 ( .A(n6970), .B(n6971), .Z(n6948) );
  AND U9262 ( .A(n6972), .B(n6973), .Z(n6971) );
  AND U9263 ( .A(n6974), .B(n6975), .Z(n6973) );
  AND U9264 ( .A(n6976), .B(n6977), .Z(n6972) );
  AND U9265 ( .A(n6978), .B(n6979), .Z(n6970) );
  AND U9266 ( .A(n6980), .B(n6981), .Z(n6979) );
  AND U9267 ( .A(n6982), .B(n6983), .Z(n6978) );
  NAND U9268 ( .A(n6882), .B(n6984), .Z(n6982) );
  NANDN U9269 ( .B(n6913), .A(n6985), .Z(n6899) );
  NAND U9270 ( .A(n6986), .B(n6987), .Z(n6913) );
  ANDN U9271 ( .A(n6988), .B(n6989), .Z(n6987) );
  ANDN U9272 ( .A(n6990), .B(n6991), .Z(n6986) );
  NAND U9273 ( .A(\u_a23_core/u_execute/alu_out[29] ), .B(n6766), .Z(n6771) );
  IV U9274 ( .A(n6992), .Z(\u_a23_core/u_execute/n1074 ) );
  MUX U9275 ( .IN0(n6993), .IN1(n6994), .SEL(n6995), .F(n6992) );
  ANDN U9276 ( .A(n6996), .B(n6997), .Z(n6994) );
  MUX U9277 ( .IN0(n6766), .IN1(n6998), .SEL(n6999), .F(n6997) );
  AND U9278 ( .A(n7000), .B(n7001), .Z(n6998) );
  AND U9279 ( .A(n7002), .B(n7003), .Z(n7001) );
  AND U9280 ( .A(n7004), .B(n7005), .Z(n7003) );
  AND U9281 ( .A(n7006), .B(n7007), .Z(n7005) );
  AND U9282 ( .A(n7008), .B(n7009), .Z(n7007) );
  AND U9283 ( .A(n7010), .B(n7011), .Z(n7006) );
  AND U9284 ( .A(n7012), .B(n7013), .Z(n7004) );
  AND U9285 ( .A(n7014), .B(n7015), .Z(n7013) );
  AND U9286 ( .A(n7016), .B(n7017), .Z(n7012) );
  AND U9287 ( .A(n7018), .B(n7019), .Z(n7002) );
  AND U9288 ( .A(n7020), .B(n7021), .Z(n7019) );
  AND U9289 ( .A(n7022), .B(n7023), .Z(n7021) );
  AND U9290 ( .A(n7024), .B(n7025), .Z(n7020) );
  AND U9291 ( .A(n7026), .B(n7027), .Z(n7018) );
  AND U9292 ( .A(n7028), .B(n7029), .Z(n7027) );
  AND U9293 ( .A(n7030), .B(n7031), .Z(n7026) );
  AND U9294 ( .A(n7032), .B(n7033), .Z(n7000) );
  AND U9295 ( .A(n7034), .B(n7035), .Z(n7033) );
  AND U9296 ( .A(n7036), .B(n7037), .Z(n7035) );
  AND U9297 ( .A(n7038), .B(n7039), .Z(n7037) );
  AND U9298 ( .A(n7040), .B(n7041), .Z(n7036) );
  AND U9299 ( .A(n7042), .B(n7043), .Z(n7034) );
  AND U9300 ( .A(n7044), .B(n7045), .Z(n7043) );
  AND U9301 ( .A(n7046), .B(n7047), .Z(n7042) );
  AND U9302 ( .A(n7048), .B(n7049), .Z(n7032) );
  AND U9303 ( .A(n7050), .B(n7051), .Z(n7049) );
  AND U9304 ( .A(n7052), .B(n7053), .Z(n7051) );
  AND U9305 ( .A(n7054), .B(n7055), .Z(n7050) );
  AND U9306 ( .A(n7056), .B(n7057), .Z(n7048) );
  AND U9307 ( .A(n6774), .B(n7058), .Z(n7057) );
  AND U9308 ( .A(n6340), .B(n7059), .Z(n7056) );
  NAND U9309 ( .A(n7060), .B(n7061), .Z(n6996) );
  AND U9310 ( .A(n7062), .B(n7063), .Z(n7061) );
  AND U9311 ( .A(n7064), .B(n7065), .Z(n7063) );
  AND U9312 ( .A(n7066), .B(n7067), .Z(n7065) );
  ANDN U9313 ( .A(n7068), .B(\u_a23_core/u_execute/multiply_out[7] ), .Z(n7067) );
  NOR U9314 ( .A(\u_a23_core/u_execute/multiply_out[8] ), .B(
        \u_a23_core/u_execute/multiply_out[9] ), .Z(n7068) );
  NOR U9315 ( .A(\u_a23_core/u_execute/multiply_out[5] ), .B(
        \u_a23_core/u_execute/multiply_out[6] ), .Z(n7066) );
  AND U9316 ( .A(n7069), .B(n7070), .Z(n7064) );
  NOR U9317 ( .A(\u_a23_core/u_execute/multiply_out[3] ), .B(
        \u_a23_core/u_execute/multiply_out[4] ), .Z(n7070) );
  ANDN U9318 ( .A(n7071), .B(\u_a23_core/u_execute/multiply_out[30] ), .Z(
        n7069) );
  IV U9319 ( .A(\u_a23_core/u_execute/multiply_out[31] ), .Z(n7071) );
  AND U9320 ( .A(n7072), .B(n7073), .Z(n7062) );
  AND U9321 ( .A(n7074), .B(n7075), .Z(n7073) );
  NOR U9322 ( .A(\u_a23_core/u_execute/multiply_out[29] ), .B(
        \u_a23_core/u_execute/multiply_out[2] ), .Z(n7075) );
  NOR U9323 ( .A(\u_a23_core/u_execute/multiply_out[27] ), .B(
        \u_a23_core/u_execute/multiply_out[28] ), .Z(n7074) );
  AND U9324 ( .A(n7076), .B(n7077), .Z(n7072) );
  NOR U9325 ( .A(\u_a23_core/u_execute/multiply_out[25] ), .B(
        \u_a23_core/u_execute/multiply_out[26] ), .Z(n7077) );
  NOR U9326 ( .A(\u_a23_core/u_execute/multiply_out[23] ), .B(
        \u_a23_core/u_execute/multiply_out[24] ), .Z(n7076) );
  AND U9327 ( .A(n7078), .B(n7079), .Z(n7060) );
  AND U9328 ( .A(n7080), .B(n7081), .Z(n7079) );
  AND U9329 ( .A(n7082), .B(n7083), .Z(n7081) );
  NOR U9330 ( .A(\u_a23_core/u_execute/multiply_out[21] ), .B(
        \u_a23_core/u_execute/multiply_out[22] ), .Z(n7083) );
  NOR U9331 ( .A(\u_a23_core/u_execute/multiply_out[1] ), .B(
        \u_a23_core/u_execute/multiply_out[20] ), .Z(n7082) );
  AND U9332 ( .A(n7084), .B(n7085), .Z(n7080) );
  NOR U9333 ( .A(\u_a23_core/u_execute/multiply_out[18] ), .B(
        \u_a23_core/u_execute/multiply_out[19] ), .Z(n7085) );
  NOR U9334 ( .A(\u_a23_core/u_execute/multiply_out[16] ), .B(
        \u_a23_core/u_execute/multiply_out[17] ), .Z(n7084) );
  AND U9335 ( .A(n7086), .B(n7087), .Z(n7078) );
  AND U9336 ( .A(n7088), .B(n7089), .Z(n7087) );
  NOR U9337 ( .A(\u_a23_core/u_execute/multiply_out[14] ), .B(
        \u_a23_core/u_execute/multiply_out[15] ), .Z(n7089) );
  NOR U9338 ( .A(\u_a23_core/u_execute/multiply_out[12] ), .B(
        \u_a23_core/u_execute/multiply_out[13] ), .Z(n7088) );
  AND U9339 ( .A(n7090), .B(n7091), .Z(n7086) );
  NOR U9340 ( .A(\u_a23_core/u_execute/multiply_out[10] ), .B(
        \u_a23_core/u_execute/multiply_out[11] ), .Z(n7091) );
  AND U9341 ( .A(n6770), .B(n6406), .Z(n7090) );
  IV U9342 ( .A(\u_a23_core/u_execute/multiply_out[0] ), .Z(n6406) );
  IV U9343 ( .A(n7092), .Z(\u_a23_core/u_execute/n1073 ) );
  MUX U9344 ( .IN0(n7093), .IN1(n7094), .SEL(n6769), .F(n7092) );
  IV U9345 ( .A(n6995), .Z(n6769) );
  ANDN U9346 ( .A(\u_a23_core/status_bits_flags_wen ), .B(n6099), .Z(n6995) );
  AND U9347 ( .A(n7095), .B(n7096), .Z(n7093) );
  NAND U9348 ( .A(\u_a23_core/u_execute/alu_out[31] ), .B(n7097), .Z(n7096) );
  OR U9349 ( .A(n6766), .B(n6774), .Z(n7097) );
  NOR U9350 ( .A(n6766), .B(n6770), .Z(n6774) );
  ANDN U9351 ( .A(\u_a23_core/status_bits_sel[0] ), .B(
        \u_a23_core/status_bits_sel[2] ), .Z(n6766) );
  NAND U9352 ( .A(\u_a23_core/u_execute/multiply_out[31] ), .B(n6770), .Z(
        n7095) );
  ANDN U9353 ( .A(\u_a23_core/status_bits_sel[2] ), .B(
        \u_a23_core/status_bits_sel[0] ), .Z(n6770) );
  NAND U9354 ( .A(\u_a23_core/byte_enable_sel[0] ), .B(n7098), .Z(
        \u_a23_core/u_execute/byte_enable_nxt[3] ) );
  NAND U9355 ( .A(\u_a23_core/execute_address_nxt[1] ), .B(
        \u_a23_core/execute_address_nxt[0] ), .Z(n7098) );
  NAND U9356 ( .A(\u_a23_core/byte_enable_sel[0] ), .B(n7099), .Z(
        \u_a23_core/u_execute/byte_enable_nxt[2] ) );
  NAND U9357 ( .A(n7100), .B(\u_a23_core/execute_address_nxt[1] ), .Z(n7099)
         );
  NAND U9358 ( .A(\u_a23_core/byte_enable_sel[0] ), .B(n7101), .Z(
        \u_a23_core/u_execute/byte_enable_nxt[1] ) );
  NAND U9359 ( .A(n7102), .B(\u_a23_core/execute_address_nxt[0] ), .Z(n7101)
         );
  NAND U9360 ( .A(\u_a23_core/byte_enable_sel[0] ), .B(n7103), .Z(
        \u_a23_core/u_execute/byte_enable_nxt[0] ) );
  NAND U9361 ( .A(n7102), .B(n7100), .Z(n7103) );
  IV U9362 ( .A(\u_a23_core/execute_address_nxt[1] ), .Z(n7102) );
  AND U9363 ( .A(n7104), .B(n7105), .Z(
        \u_a23_core/u_decode/write_data_wen_nxt ) );
  NANDN U9364 ( .B(n7106), .A(n7107), .Z(n7104) );
  NANDN U9365 ( .B(\u_a23_core/u_decode/alu_function_nxt[2] ), .A(n7108), .Z(
        \u_a23_core/u_decode/use_carry_in_nxt ) );
  NAND U9366 ( .A(n7109), .B(n7110), .Z(n7108) );
  NAND U9367 ( .A(n7111), .B(n7112), .Z(n7110) );
  NANDN U9368 ( .B(n7113), .A(n7114), .Z(n7112) );
  AND U9369 ( .A(n7115), .B(n7116), .Z(n7111) );
  NAND U9370 ( .A(n7117), .B(n7118), .Z(n7115) );
  AND U9371 ( .A(n7119), .B(\u_a23_core/u_decode/instruction[5] ), .Z(n7118)
         );
  AND U9372 ( .A(\u_a23_core/u_decode/instruction[6] ), .B(n7120), .Z(n7119)
         );
  AND U9373 ( .A(n7121), .B(n7122), .Z(n7117) );
  AND U9374 ( .A(n7123), .B(n7124), .Z(n7121) );
  NAND U9375 ( .A(n7125), .B(n7126), .Z(
        \u_a23_core/u_decode/status_bits_sel_nxt_0 ) );
  ANDN U9376 ( .A(n7127), .B(\u_a23_core/u_decode/alu_function_nxt[4] ), .Z(
        n7125) );
  NANDN U9377 ( .B(n7128), .A(n7129), .Z(n7127) );
  NAND U9378 ( .A(n7130), .B(n7131), .Z(
        \u_a23_core/u_decode/status_bits_sel_nxt[2] ) );
  NAND U9379 ( .A(n7128), .B(\u_a23_core/u_decode/alu_function_nxt[4] ), .Z(
        n7131) );
  NAND U9380 ( .A(n7132), .B(n7133), .Z(n7128) );
  AND U9381 ( .A(n7134), .B(n7135), .Z(n7132) );
  NAND U9382 ( .A(n7135), .B(n16637), .Z(n7130) );
  NAND U9383 ( .A(n7126), .B(n7136), .Z(
        \u_a23_core/u_decode/status_bits_flags_wen_nxt ) );
  NAND U9384 ( .A(n7135), .B(n7137), .Z(n7136) );
  NAND U9385 ( .A(n7138), .B(n7139), .Z(n7137) );
  NANDN U9386 ( .B(n7140), .A(n7114), .Z(n7126) );
  AND U9387 ( .A(n7141), .B(n7122), .Z(
        \u_a23_core/u_decode/shift_imm_zero_nxt ) );
  ANDN U9388 ( .A(\u_a23_core/u_decode/barrel_shift_amount_sel_nxt[1] ), .B(
        \u_a23_core/u_decode/barrel_shift_amount_sel_nxt[0] ), .Z(n7141) );
  AND U9389 ( .A(\u_a23_core/u_decode/pc_sel_nxt[1] ), .B(n7142), .Z(
        \u_a23_core/u_decode/reg_write_sel_nxt[0] ) );
  NOR U9390 ( .A(n7143), .B(n7144), .Z(\u_a23_core/u_decode/n1511 ) );
  NOR U9391 ( .A(n7144), .B(n7145), .Z(\u_a23_core/u_decode/n1510 ) );
  NOR U9392 ( .A(n7144), .B(n7146), .Z(\u_a23_core/u_decode/n1509 ) );
  ANDN U9393 ( .A(n7147), .B(n7144), .Z(\u_a23_core/u_decode/n1508 ) );
  NAND U9394 ( .A(n7148), .B(n7149), .Z(n7144) );
  ANDN U9395 ( .A(n7150), .B(n7143), .Z(\u_a23_core/u_decode/n1507 ) );
  ANDN U9396 ( .A(n7150), .B(n7145), .Z(\u_a23_core/u_decode/n1506 ) );
  ANDN U9397 ( .A(n7150), .B(n7146), .Z(\u_a23_core/u_decode/n1505 ) );
  ANDN U9398 ( .A(n7151), .B(n7145), .Z(\u_a23_core/u_decode/n1504 ) );
  ANDN U9399 ( .A(n7151), .B(n7146), .Z(\u_a23_core/u_decode/n1503 ) );
  AND U9400 ( .A(n7151), .B(n7147), .Z(\u_a23_core/u_decode/n1502 ) );
  AND U9401 ( .A(n7149), .B(n7152), .Z(n7151) );
  ANDN U9402 ( .A(n7153), .B(n7143), .Z(\u_a23_core/u_decode/n1501 ) );
  NAND U9403 ( .A(n7154), .B(n7155), .Z(n7143) );
  ANDN U9404 ( .A(n7153), .B(n7145), .Z(\u_a23_core/u_decode/n1500 ) );
  NAND U9405 ( .A(n7156), .B(n7155), .Z(n7145) );
  IV U9406 ( .A(n7154), .Z(n7156) );
  ANDN U9407 ( .A(n7153), .B(n7146), .Z(\u_a23_core/u_decode/n1499 ) );
  NANDN U9408 ( .B(n7155), .A(n7154), .Z(n7146) );
  AND U9409 ( .A(n7153), .B(n7147), .Z(\u_a23_core/u_decode/n1498 ) );
  NOR U9410 ( .A(n7148), .B(n7149), .Z(n7153) );
  IV U9411 ( .A(n7152), .Z(n7148) );
  MUX U9412 ( .IN0(\u_a23_core/u_decode/pre_fetch_instruction[0] ), .IN1(
        \u_a23_core/read_data_s2[0] ), .SEL(n7157), .F(
        \u_a23_core/u_decode/n1495 ) );
  NANDN U9413 ( .B(n7158), .A(n7159), .Z(\u_a23_core/u_decode/n1494 ) );
  NANDN U9414 ( .B(n7160), .A(\u_a23_core/multiply_function[0] ), .Z(n7159) );
  NAND U9415 ( .A(n7161), .B(n7162), .Z(\u_a23_core/u_decode/n1493 ) );
  NAND U9416 ( .A(n7163), .B(n7158), .Z(n7162) );
  NANDN U9417 ( .B(n7160), .A(\u_a23_core/multiply_function[1] ), .Z(n7161) );
  AND U9418 ( .A(n7164), .B(n7165), .Z(n7160) );
  MUX U9419 ( .IN0(\u_a23_core/u_decode/saved_current_instruction[16] ), .IN1(
        n7166), .SEL(n7167), .F(\u_a23_core/u_decode/n1492 ) );
  MUX U9420 ( .IN0(\u_a23_core/u_decode/saved_current_instruction[17] ), .IN1(
        n7168), .SEL(n7167), .F(\u_a23_core/u_decode/n1491 ) );
  MUX U9421 ( .IN0(\u_a23_core/u_decode/saved_current_instruction[18] ), .IN1(
        n7169), .SEL(n7167), .F(\u_a23_core/u_decode/n1490 ) );
  MUX U9422 ( .IN0(\u_a23_core/u_decode/saved_current_instruction[19] ), .IN1(
        n7170), .SEL(n7167), .F(\u_a23_core/u_decode/n1489 ) );
  MUX U9423 ( .IN0(\u_a23_core/u_decode/saved_current_instruction[20] ), .IN1(
        n7135), .SEL(n7167), .F(\u_a23_core/u_decode/n1488 ) );
  MUX U9424 ( .IN0(\u_a23_core/u_decode/saved_current_instruction[21] ), .IN1(
        n7163), .SEL(n7167), .F(\u_a23_core/u_decode/n1487 ) );
  MUX U9425 ( .IN0(\u_a23_core/u_decode/saved_current_instruction[22] ), .IN1(
        n7114), .SEL(n7167), .F(\u_a23_core/u_decode/n1486 ) );
  MUX U9426 ( .IN0(\u_a23_core/u_decode/saved_current_instruction[23] ), .IN1(
        n7171), .SEL(n7167), .F(\u_a23_core/u_decode/n1485 ) );
  MUX U9427 ( .IN0(\u_a23_core/u_decode/saved_current_instruction[24] ), .IN1(
        n7142), .SEL(n7167), .F(\u_a23_core/u_decode/n1484 ) );
  MUX U9428 ( .IN0(\u_a23_core/u_decode/saved_current_instruction[25] ), .IN1(
        n7172), .SEL(n7167), .F(\u_a23_core/u_decode/n1483 ) );
  MUX U9429 ( .IN0(\u_a23_core/u_decode/saved_current_instruction[26] ), .IN1(
        n7173), .SEL(n7167), .F(\u_a23_core/u_decode/n1482 ) );
  MUX U9430 ( .IN0(\u_a23_core/u_decode/saved_current_instruction[27] ), .IN1(
        n7174), .SEL(n7167), .F(\u_a23_core/u_decode/n1481 ) );
  NAND U9431 ( .A(n7175), .B(n7176), .Z(\u_a23_core/u_decode/n1480 ) );
  NAND U9432 ( .A(n7177), .B(
        \u_a23_core/u_decode/saved_current_instruction[0] ), .Z(n7176) );
  NAND U9433 ( .A(\u_a23_core/rm_sel_nxt[0] ), .B(n7178), .Z(n7175) );
  NAND U9434 ( .A(n7179), .B(n7180), .Z(\u_a23_core/u_decode/n1479 ) );
  NAND U9435 ( .A(n7181), .B(n7182), .Z(n7180) );
  AND U9436 ( .A(n7183), .B(n7184), .Z(n7179) );
  NAND U9437 ( .A(n7177), .B(
        \u_a23_core/u_decode/saved_current_instruction[1] ), .Z(n7184) );
  NAND U9438 ( .A(n7178), .B(\u_a23_core/rm_sel_nxt[1] ), .Z(n7183) );
  NAND U9439 ( .A(n7185), .B(n7186), .Z(\u_a23_core/u_decode/n1478 ) );
  NAND U9440 ( .A(\u_a23_core/rm_sel_nxt[2] ), .B(n7178), .Z(n7186) );
  AND U9441 ( .A(n7187), .B(n7188), .Z(n7185) );
  NAND U9442 ( .A(n7181), .B(n7189), .Z(n7188) );
  NAND U9443 ( .A(n7177), .B(
        \u_a23_core/u_decode/saved_current_instruction[2] ), .Z(n7187) );
  NAND U9444 ( .A(n7190), .B(n7191), .Z(\u_a23_core/u_decode/n1477 ) );
  NAND U9445 ( .A(\u_a23_core/rm_sel_nxt[3] ), .B(n7192), .Z(n7191) );
  NANDN U9446 ( .B(n7178), .A(n7193), .Z(n7192) );
  NAND U9447 ( .A(n7181), .B(n7194), .Z(n7193) );
  NAND U9448 ( .A(n7177), .B(
        \u_a23_core/u_decode/saved_current_instruction[3] ), .Z(n7190) );
  NAND U9449 ( .A(n7195), .B(n7196), .Z(\u_a23_core/u_decode/n1476 ) );
  NAND U9450 ( .A(n7181), .B(n7197), .Z(n7196) );
  AND U9451 ( .A(n7198), .B(n7199), .Z(n7195) );
  NAND U9452 ( .A(n7177), .B(
        \u_a23_core/u_decode/saved_current_instruction[4] ), .Z(n7199) );
  NAND U9453 ( .A(\u_a23_core/u_decode/instruction[4] ), .B(n7178), .Z(n7198)
         );
  NAND U9454 ( .A(n7200), .B(n7201), .Z(\u_a23_core/u_decode/n1475 ) );
  OR U9455 ( .A(n7202), .B(n7203), .Z(n7201) );
  NAND U9456 ( .A(n7177), .B(
        \u_a23_core/u_decode/saved_current_instruction[5] ), .Z(n7200) );
  NAND U9457 ( .A(n7204), .B(n7205), .Z(\u_a23_core/u_decode/n1474 ) );
  NANDN U9458 ( .B(n7206), .A(\u_a23_core/u_decode/instruction[6] ), .Z(n7205)
         );
  NAND U9459 ( .A(n7177), .B(
        \u_a23_core/u_decode/saved_current_instruction[6] ), .Z(n7204) );
  NAND U9460 ( .A(n7207), .B(n7208), .Z(\u_a23_core/u_decode/n1473 ) );
  NAND U9461 ( .A(\u_a23_core/u_decode/instruction[7] ), .B(n7209), .Z(n7208)
         );
  NAND U9462 ( .A(n7210), .B(n7206), .Z(n7209) );
  AND U9463 ( .A(n7202), .B(n7211), .Z(n7206) );
  NAND U9464 ( .A(\u_a23_core/u_decode/instruction[5] ), .B(n7181), .Z(n7211)
         );
  ANDN U9465 ( .A(n7212), .B(n7178), .Z(n7202) );
  OR U9466 ( .A(n7213), .B(n7214), .Z(n7212) );
  NAND U9467 ( .A(n7181), .B(\u_a23_core/u_decode/instruction[6] ), .Z(n7210)
         );
  NAND U9468 ( .A(n7177), .B(
        \u_a23_core/u_decode/saved_current_instruction[7] ), .Z(n7207) );
  NAND U9469 ( .A(n7215), .B(n7216), .Z(\u_a23_core/u_decode/n1472 ) );
  NAND U9470 ( .A(n7181), .B(n7217), .Z(n7216) );
  AND U9471 ( .A(n7218), .B(n7219), .Z(n7215) );
  NAND U9472 ( .A(n7177), .B(
        \u_a23_core/u_decode/saved_current_instruction[8] ), .Z(n7219) );
  NAND U9473 ( .A(\u_a23_core/u_decode/instruction[8] ), .B(n7178), .Z(n7218)
         );
  NAND U9474 ( .A(n7220), .B(n7221), .Z(\u_a23_core/u_decode/n1471 ) );
  NAND U9475 ( .A(\u_a23_core/u_decode/instruction[9] ), .B(n7222), .Z(n7221)
         );
  NANDN U9476 ( .B(n7178), .A(n7223), .Z(n7222) );
  OR U9477 ( .A(n7224), .B(n7214), .Z(n7223) );
  NAND U9478 ( .A(n7177), .B(
        \u_a23_core/u_decode/saved_current_instruction[9] ), .Z(n7220) );
  NAND U9479 ( .A(n7225), .B(n7226), .Z(\u_a23_core/u_decode/n1470 ) );
  NAND U9480 ( .A(\u_a23_core/u_decode/instruction[10] ), .B(n7178), .Z(n7226)
         );
  AND U9481 ( .A(n7227), .B(n7228), .Z(n7225) );
  NAND U9482 ( .A(n7181), .B(n7229), .Z(n7228) );
  NAND U9483 ( .A(n7177), .B(
        \u_a23_core/u_decode/saved_current_instruction[10] ), .Z(n7227) );
  NAND U9484 ( .A(n7230), .B(n7231), .Z(\u_a23_core/u_decode/n1469 ) );
  NAND U9485 ( .A(n7181), .B(n7232), .Z(n7231) );
  AND U9486 ( .A(n7233), .B(n7234), .Z(n7230) );
  NAND U9487 ( .A(n7177), .B(
        \u_a23_core/u_decode/saved_current_instruction[11] ), .Z(n7234) );
  NAND U9488 ( .A(\u_a23_core/u_decode/instruction[11] ), .B(n7178), .Z(n7233)
         );
  NAND U9489 ( .A(n7235), .B(n7236), .Z(\u_a23_core/u_decode/n1468 ) );
  NAND U9490 ( .A(n7237), .B(n7178), .Z(n7236) );
  AND U9491 ( .A(n7238), .B(n7239), .Z(n7235) );
  NAND U9492 ( .A(n7181), .B(n7240), .Z(n7239) );
  NAND U9493 ( .A(n7177), .B(
        \u_a23_core/u_decode/saved_current_instruction[12] ), .Z(n7238) );
  NAND U9494 ( .A(n7241), .B(n7242), .Z(\u_a23_core/u_decode/n1467 ) );
  NAND U9495 ( .A(n7181), .B(n7243), .Z(n7242) );
  AND U9496 ( .A(n7244), .B(n7245), .Z(n7241) );
  NAND U9497 ( .A(n7177), .B(
        \u_a23_core/u_decode/saved_current_instruction[13] ), .Z(n7245) );
  NAND U9498 ( .A(n7246), .B(n7178), .Z(n7244) );
  NAND U9499 ( .A(n7247), .B(n7248), .Z(\u_a23_core/u_decode/n1466 ) );
  NAND U9500 ( .A(n7249), .B(n7250), .Z(n7248) );
  NANDN U9501 ( .B(n7178), .A(n7251), .Z(n7250) );
  OR U9502 ( .A(n7252), .B(n7214), .Z(n7251) );
  NAND U9503 ( .A(n7177), .B(
        \u_a23_core/u_decode/saved_current_instruction[14] ), .Z(n7247) );
  NAND U9504 ( .A(n7253), .B(n7254), .Z(\u_a23_core/u_decode/n1465 ) );
  NAND U9505 ( .A(n7181), .B(n7255), .Z(n7254) );
  AND U9506 ( .A(n7256), .B(n7257), .Z(n7253) );
  NAND U9507 ( .A(n7177), .B(
        \u_a23_core/u_decode/saved_current_instruction[15] ), .Z(n7257) );
  NAND U9508 ( .A(n7258), .B(n7178), .Z(n7256) );
  MUX U9509 ( .IN0(\u_a23_core/u_decode/pre_fetch_instruction[1] ), .IN1(
        \u_a23_core/read_data_s2[1] ), .SEL(n7157), .F(
        \u_a23_core/u_decode/n1464 ) );
  MUX U9510 ( .IN0(\u_a23_core/u_decode/pre_fetch_instruction[2] ), .IN1(
        \u_a23_core/read_data_s2[2] ), .SEL(n7157), .F(
        \u_a23_core/u_decode/n1463 ) );
  MUX U9511 ( .IN0(\u_a23_core/u_decode/pre_fetch_instruction[3] ), .IN1(
        \u_a23_core/read_data_s2[3] ), .SEL(n7157), .F(
        \u_a23_core/u_decode/n1462 ) );
  MUX U9512 ( .IN0(\u_a23_core/u_decode/pre_fetch_instruction[4] ), .IN1(
        \u_a23_core/read_data_s2[4] ), .SEL(n7157), .F(
        \u_a23_core/u_decode/n1461 ) );
  MUX U9513 ( .IN0(\u_a23_core/u_decode/pre_fetch_instruction[5] ), .IN1(
        \u_a23_core/read_data_s2[5] ), .SEL(n7157), .F(
        \u_a23_core/u_decode/n1460 ) );
  MUX U9514 ( .IN0(\u_a23_core/u_decode/pre_fetch_instruction[6] ), .IN1(
        \u_a23_core/read_data_s2[6] ), .SEL(n7157), .F(
        \u_a23_core/u_decode/n1459 ) );
  MUX U9515 ( .IN0(\u_a23_core/u_decode/pre_fetch_instruction[7] ), .IN1(
        \u_a23_core/read_data_s2[7] ), .SEL(n7157), .F(
        \u_a23_core/u_decode/n1458 ) );
  MUX U9516 ( .IN0(\u_a23_core/u_decode/pre_fetch_instruction[8] ), .IN1(
        \u_a23_core/read_data_s2[8] ), .SEL(n7157), .F(
        \u_a23_core/u_decode/n1457 ) );
  MUX U9517 ( .IN0(\u_a23_core/u_decode/pre_fetch_instruction[9] ), .IN1(
        \u_a23_core/read_data_s2[9] ), .SEL(n7157), .F(
        \u_a23_core/u_decode/n1456 ) );
  MUX U9518 ( .IN0(\u_a23_core/u_decode/pre_fetch_instruction[10] ), .IN1(
        \u_a23_core/read_data_s2[10] ), .SEL(n7157), .F(
        \u_a23_core/u_decode/n1455 ) );
  MUX U9519 ( .IN0(\u_a23_core/u_decode/pre_fetch_instruction[11] ), .IN1(
        \u_a23_core/read_data_s2[11] ), .SEL(n7157), .F(
        \u_a23_core/u_decode/n1454 ) );
  MUX U9520 ( .IN0(\u_a23_core/u_decode/pre_fetch_instruction[12] ), .IN1(
        \u_a23_core/read_data_s2[12] ), .SEL(n7157), .F(
        \u_a23_core/u_decode/n1453 ) );
  MUX U9521 ( .IN0(\u_a23_core/u_decode/pre_fetch_instruction[13] ), .IN1(
        \u_a23_core/read_data_s2[13] ), .SEL(n7157), .F(
        \u_a23_core/u_decode/n1452 ) );
  MUX U9522 ( .IN0(\u_a23_core/u_decode/pre_fetch_instruction[14] ), .IN1(
        \u_a23_core/read_data_s2[14] ), .SEL(n7157), .F(
        \u_a23_core/u_decode/n1451 ) );
  MUX U9523 ( .IN0(\u_a23_core/u_decode/pre_fetch_instruction[15] ), .IN1(
        \u_a23_core/read_data_s2[15] ), .SEL(n7157), .F(
        \u_a23_core/u_decode/n1450 ) );
  MUX U9524 ( .IN0(\u_a23_core/u_decode/pre_fetch_instruction[16] ), .IN1(
        \u_a23_core/read_data_s2[16] ), .SEL(n7157), .F(
        \u_a23_core/u_decode/n1449 ) );
  MUX U9525 ( .IN0(\u_a23_core/u_decode/pre_fetch_instruction[17] ), .IN1(
        \u_a23_core/read_data_s2[17] ), .SEL(n7157), .F(
        \u_a23_core/u_decode/n1448 ) );
  MUX U9526 ( .IN0(\u_a23_core/u_decode/pre_fetch_instruction[18] ), .IN1(
        \u_a23_core/read_data_s2[18] ), .SEL(n7157), .F(
        \u_a23_core/u_decode/n1447 ) );
  MUX U9527 ( .IN0(\u_a23_core/u_decode/pre_fetch_instruction[19] ), .IN1(
        \u_a23_core/read_data_s2[19] ), .SEL(n7157), .F(
        \u_a23_core/u_decode/n1446 ) );
  MUX U9528 ( .IN0(\u_a23_core/u_decode/pre_fetch_instruction[20] ), .IN1(
        \u_a23_core/read_data_s2[20] ), .SEL(n7157), .F(
        \u_a23_core/u_decode/n1445 ) );
  MUX U9529 ( .IN0(\u_a23_core/u_decode/pre_fetch_instruction[21] ), .IN1(
        \u_a23_core/read_data_s2[21] ), .SEL(n7157), .F(
        \u_a23_core/u_decode/n1444 ) );
  MUX U9530 ( .IN0(\u_a23_core/u_decode/pre_fetch_instruction[22] ), .IN1(
        \u_a23_core/read_data_s2[22] ), .SEL(n7157), .F(
        \u_a23_core/u_decode/n1443 ) );
  MUX U9531 ( .IN0(\u_a23_core/u_decode/pre_fetch_instruction[23] ), .IN1(
        \u_a23_core/read_data_s2[23] ), .SEL(n7157), .F(
        \u_a23_core/u_decode/n1442 ) );
  MUX U9532 ( .IN0(\u_a23_core/u_decode/pre_fetch_instruction[24] ), .IN1(
        \u_a23_core/read_data_s2[24] ), .SEL(n7157), .F(
        \u_a23_core/u_decode/n1441 ) );
  MUX U9533 ( .IN0(\u_a23_core/u_decode/pre_fetch_instruction[25] ), .IN1(
        \u_a23_core/read_data_s2[25] ), .SEL(n7157), .F(
        \u_a23_core/u_decode/n1440 ) );
  MUX U9534 ( .IN0(\u_a23_core/u_decode/pre_fetch_instruction[26] ), .IN1(
        \u_a23_core/read_data_s2[26] ), .SEL(n7157), .F(
        \u_a23_core/u_decode/n1439 ) );
  MUX U9535 ( .IN0(\u_a23_core/u_decode/pre_fetch_instruction[27] ), .IN1(
        \u_a23_core/read_data_s2[27] ), .SEL(n7157), .F(
        \u_a23_core/u_decode/n1438 ) );
  MUX U9536 ( .IN0(\u_a23_core/u_decode/pre_fetch_instruction[28] ), .IN1(
        \u_a23_core/read_data_s2[28] ), .SEL(n7157), .F(
        \u_a23_core/u_decode/n1437 ) );
  IV U9537 ( .A(n7259), .Z(n7157) );
  MUX U9538 ( .IN0(\u_a23_core/read_data_s2[29] ), .IN1(
        \u_a23_core/u_decode/pre_fetch_instruction[29] ), .SEL(n7259), .F(
        \u_a23_core/u_decode/n1436 ) );
  MUX U9539 ( .IN0(\u_a23_core/read_data_s2[30] ), .IN1(
        \u_a23_core/u_decode/pre_fetch_instruction[30] ), .SEL(n7259), .F(
        \u_a23_core/u_decode/n1435 ) );
  MUX U9540 ( .IN0(\u_a23_core/read_data_s2[31] ), .IN1(
        \u_a23_core/u_decode/pre_fetch_instruction[31] ), .SEL(n7259), .F(
        \u_a23_core/u_decode/n1434 ) );
  AND U9541 ( .A(n7260), .B(n7261), .Z(n7259) );
  AND U9542 ( .A(n7262), .B(n7263), .Z(n7261) );
  IV U9543 ( .A(n7264), .Z(\u_a23_core/u_decode/n1433 ) );
  MUX U9544 ( .IN0(n7265), .IN1(n7266), .SEL(n7129), .F(n7264) );
  AND U9545 ( .A(n7267), .B(n7268), .Z(n7266) );
  NANDN U9546 ( .B(n7269), .A(\u_a23_core/read_data_s2[28] ), .Z(n7268) );
  NANDN U9547 ( .B(n7270), .A(\u_a23_core/u_decode/pre_fetch_instruction[28] ), 
        .Z(n7267) );
  IV U9548 ( .A(n7271), .Z(\u_a23_core/u_decode/n1431 ) );
  MUX U9549 ( .IN0(n7272), .IN1(n7273), .SEL(n7129), .F(n7271) );
  AND U9550 ( .A(n7274), .B(n7275), .Z(n7273) );
  NANDN U9551 ( .B(n7269), .A(\u_a23_core/read_data_s2[29] ), .Z(n7275) );
  NANDN U9552 ( .B(n7270), .A(\u_a23_core/u_decode/pre_fetch_instruction[29] ), 
        .Z(n7274) );
  MUX U9553 ( .IN0(n7276), .IN1(\u_a23_core/condition[2] ), .SEL(n7277), .F(
        \u_a23_core/u_decode/n1429 ) );
  NAND U9554 ( .A(n7278), .B(n7279), .Z(n7276) );
  NANDN U9555 ( .B(n7269), .A(\u_a23_core/read_data_s2[30] ), .Z(n7279) );
  NANDN U9556 ( .B(n7270), .A(\u_a23_core/u_decode/pre_fetch_instruction[30] ), 
        .Z(n7278) );
  MUX U9557 ( .IN0(n7280), .IN1(\u_a23_core/condition[3] ), .SEL(n7277), .F(
        \u_a23_core/u_decode/n1427 ) );
  NAND U9558 ( .A(n7281), .B(n7282), .Z(n7280) );
  NANDN U9559 ( .B(n7269), .A(\u_a23_core/read_data_s2[31] ), .Z(n7282) );
  NANDN U9560 ( .B(n7270), .A(\u_a23_core/u_decode/pre_fetch_instruction[31] ), 
        .Z(n7281) );
  IV U9561 ( .A(n7177), .Z(n7167) );
  ANDN U9562 ( .A(n7214), .B(n7178), .Z(n7177) );
  AND U9563 ( .A(n7284), .B(n7129), .Z(n7178) );
  NAND U9564 ( .A(n7285), .B(n7286), .Z(n7284) );
  IV U9565 ( .A(n7287), .Z(n7286) );
  NAND U9566 ( .A(n7288), .B(n7289), .Z(\u_a23_core/u_decode/imm32_nxt[9] ) );
  AND U9567 ( .A(n7290), .B(n7291), .Z(n7289) );
  NANDN U9568 ( .B(n7292), .A(\u_a23_core/u_decode/instruction[5] ), .Z(n7291)
         );
  AND U9569 ( .A(n7293), .B(n7294), .Z(n7290) );
  NAND U9570 ( .A(\u_a23_core/u_decode/instruction[7] ), .B(n7295), .Z(n7294)
         );
  NANDN U9571 ( .B(n7296), .A(\u_a23_core/rm_sel_nxt[3] ), .Z(n7293) );
  AND U9572 ( .A(n7297), .B(n7298), .Z(n7288) );
  NANDN U9573 ( .B(n7299), .A(\u_a23_core/rm_sel_nxt[1] ), .Z(n7298) );
  NAND U9574 ( .A(\u_a23_core/u_decode/instruction[9] ), .B(n7287), .Z(n7297)
         );
  NAND U9575 ( .A(n7300), .B(n7301), .Z(\u_a23_core/u_decode/imm32_nxt[8] ) );
  AND U9576 ( .A(n7302), .B(n7303), .Z(n7301) );
  NANDN U9577 ( .B(n7292), .A(\u_a23_core/u_decode/instruction[4] ), .Z(n7303)
         );
  AND U9578 ( .A(n7304), .B(n7305), .Z(n7302) );
  NAND U9579 ( .A(\u_a23_core/u_decode/instruction[6] ), .B(n7295), .Z(n7305)
         );
  NANDN U9580 ( .B(n7296), .A(\u_a23_core/rm_sel_nxt[2] ), .Z(n7304) );
  AND U9581 ( .A(n7306), .B(n7307), .Z(n7300) );
  NANDN U9582 ( .B(n7299), .A(\u_a23_core/rm_sel_nxt[0] ), .Z(n7307) );
  NAND U9583 ( .A(\u_a23_core/u_decode/instruction[8] ), .B(n7287), .Z(n7306)
         );
  NAND U9584 ( .A(n7308), .B(n7309), .Z(\u_a23_core/u_decode/imm32_nxt[7] ) );
  AND U9585 ( .A(n7310), .B(n7311), .Z(n7309) );
  NAND U9586 ( .A(\u_a23_core/u_decode/instruction[5] ), .B(n7295), .Z(n7311)
         );
  NANDN U9587 ( .B(n7296), .A(\u_a23_core/rm_sel_nxt[1] ), .Z(n7310) );
  AND U9588 ( .A(n7312), .B(n7313), .Z(n7308) );
  NANDN U9589 ( .B(n7292), .A(\u_a23_core/rm_sel_nxt[3] ), .Z(n7313) );
  NAND U9590 ( .A(\u_a23_core/u_decode/instruction[7] ), .B(n7314), .Z(n7312)
         );
  NAND U9591 ( .A(n7315), .B(n7316), .Z(\u_a23_core/u_decode/imm32_nxt[6] ) );
  AND U9592 ( .A(n7317), .B(n7318), .Z(n7316) );
  NANDN U9593 ( .B(n7292), .A(\u_a23_core/rm_sel_nxt[2] ), .Z(n7318) );
  AND U9594 ( .A(n7319), .B(n7320), .Z(n7317) );
  NAND U9595 ( .A(\u_a23_core/u_decode/instruction[4] ), .B(n7295), .Z(n7320)
         );
  NANDN U9596 ( .B(n7296), .A(\u_a23_core/rm_sel_nxt[0] ), .Z(n7319) );
  AND U9597 ( .A(n7321), .B(n7322), .Z(n7315) );
  NAND U9598 ( .A(\u_a23_core/u_decode/instruction[6] ), .B(n7314), .Z(n7322)
         );
  NAND U9599 ( .A(n7181), .B(\u_a23_core/u_decode/mtrans_num_registers[4] ), 
        .Z(n7321) );
  NAND U9600 ( .A(n7323), .B(n7324), .Z(\u_a23_core/u_decode/imm32_nxt[5] ) );
  AND U9601 ( .A(n7325), .B(n7326), .Z(n7324) );
  NANDN U9602 ( .B(n7327), .A(\u_a23_core/u_decode/instruction[7] ), .Z(n7326)
         );
  AND U9603 ( .A(n7328), .B(n7329), .Z(n7325) );
  NAND U9604 ( .A(\u_a23_core/rm_sel_nxt[3] ), .B(n7295), .Z(n7329) );
  NANDN U9605 ( .B(n7292), .A(\u_a23_core/rm_sel_nxt[1] ), .Z(n7328) );
  AND U9606 ( .A(n7330), .B(n7331), .Z(n7323) );
  NAND U9607 ( .A(\u_a23_core/u_decode/instruction[5] ), .B(n7314), .Z(n7331)
         );
  NAND U9608 ( .A(n7181), .B(\u_a23_core/u_decode/mtrans_num_registers[3] ), 
        .Z(n7330) );
  NAND U9609 ( .A(n7332), .B(n7333), .Z(\u_a23_core/u_decode/imm32_nxt[4] ) );
  AND U9610 ( .A(n7334), .B(n7335), .Z(n7333) );
  NANDN U9611 ( .B(n7327), .A(\u_a23_core/u_decode/instruction[6] ), .Z(n7335)
         );
  AND U9612 ( .A(n7336), .B(n7337), .Z(n7334) );
  NAND U9613 ( .A(\u_a23_core/rm_sel_nxt[2] ), .B(n7295), .Z(n7337) );
  NANDN U9614 ( .B(n7292), .A(\u_a23_core/rm_sel_nxt[0] ), .Z(n7336) );
  AND U9615 ( .A(n7338), .B(n7339), .Z(n7332) );
  NAND U9616 ( .A(\u_a23_core/u_decode/instruction[4] ), .B(n7314), .Z(n7339)
         );
  NAND U9617 ( .A(n7181), .B(\u_a23_core/u_decode/mtrans_num_registers[2] ), 
        .Z(n7338) );
  NAND U9618 ( .A(n7340), .B(n7341), .Z(\u_a23_core/u_decode/imm32_nxt[3] ) );
  AND U9619 ( .A(n7342), .B(n7343), .Z(n7341) );
  NANDN U9620 ( .B(n7327), .A(\u_a23_core/u_decode/instruction[5] ), .Z(n7343)
         );
  AND U9621 ( .A(n7344), .B(n7345), .Z(n7342) );
  NAND U9622 ( .A(\u_a23_core/rm_sel_nxt[1] ), .B(n7295), .Z(n7345) );
  NANDN U9623 ( .B(n7346), .A(\u_a23_core/u_decode/instruction[7] ), .Z(n7344)
         );
  AND U9624 ( .A(n7347), .B(n7348), .Z(n7340) );
  NAND U9625 ( .A(\u_a23_core/rm_sel_nxt[3] ), .B(n7314), .Z(n7348) );
  NAND U9626 ( .A(n7181), .B(\u_a23_core/u_decode/mtrans_num_registers[1] ), 
        .Z(n7347) );
  NAND U9627 ( .A(n7349), .B(n7350), .Z(\u_a23_core/u_decode/imm32_nxt[31] )
         );
  AND U9628 ( .A(n7351), .B(n7352), .Z(n7350) );
  NANDN U9629 ( .B(n7353), .A(\u_a23_core/u_decode/instruction[5] ), .Z(n7352)
         );
  AND U9630 ( .A(n7354), .B(n7355), .Z(n7351) );
  NANDN U9631 ( .B(n7356), .A(\u_a23_core/u_decode/instruction[7] ), .Z(n7355)
         );
  AND U9632 ( .A(n7357), .B(n7358), .Z(n7349) );
  NANDN U9633 ( .B(n7346), .A(\u_a23_core/rm_sel_nxt[3] ), .Z(n7358) );
  NANDN U9634 ( .B(n7327), .A(\u_a23_core/rm_sel_nxt[1] ), .Z(n7357) );
  NAND U9635 ( .A(n7359), .B(n7360), .Z(\u_a23_core/u_decode/imm32_nxt[30] )
         );
  AND U9636 ( .A(n7361), .B(n7362), .Z(n7360) );
  NANDN U9637 ( .B(n7353), .A(\u_a23_core/u_decode/instruction[4] ), .Z(n7362)
         );
  AND U9638 ( .A(n7354), .B(n7363), .Z(n7361) );
  NANDN U9639 ( .B(n7356), .A(\u_a23_core/u_decode/instruction[6] ), .Z(n7363)
         );
  AND U9640 ( .A(n7364), .B(n7365), .Z(n7359) );
  NANDN U9641 ( .B(n7346), .A(\u_a23_core/rm_sel_nxt[2] ), .Z(n7365) );
  NANDN U9642 ( .B(n7327), .A(\u_a23_core/rm_sel_nxt[0] ), .Z(n7364) );
  NAND U9643 ( .A(n7366), .B(n7367), .Z(\u_a23_core/u_decode/imm32_nxt[2] ) );
  AND U9644 ( .A(n7368), .B(n7369), .Z(n7367) );
  NANDN U9645 ( .B(n7327), .A(\u_a23_core/u_decode/instruction[4] ), .Z(n7369)
         );
  AND U9646 ( .A(n7370), .B(n7371), .Z(n7368) );
  NAND U9647 ( .A(\u_a23_core/rm_sel_nxt[0] ), .B(n7295), .Z(n7371) );
  NANDN U9648 ( .B(n7372), .A(n7373), .Z(n7295) );
  NAND U9649 ( .A(n7374), .B(n7375), .Z(n7373) );
  AND U9650 ( .A(n7376), .B(n7377), .Z(n7375) );
  IV U9651 ( .A(n7378), .Z(n7377) );
  AND U9652 ( .A(n7379), .B(n7380), .Z(n7374) );
  IV U9653 ( .A(n7381), .Z(n7380) );
  NANDN U9654 ( .B(n7346), .A(\u_a23_core/u_decode/instruction[6] ), .Z(n7370)
         );
  AND U9655 ( .A(n7382), .B(n7383), .Z(n7366) );
  NAND U9656 ( .A(\u_a23_core/rm_sel_nxt[2] ), .B(n7314), .Z(n7383) );
  NAND U9657 ( .A(n7181), .B(\u_a23_core/u_decode/mtrans_num_registers[0] ), 
        .Z(n7382) );
  NAND U9658 ( .A(n7384), .B(n7385), .Z(\u_a23_core/u_decode/imm32_nxt[29] )
         );
  AND U9659 ( .A(n7386), .B(n7387), .Z(n7385) );
  NANDN U9660 ( .B(n7388), .A(\u_a23_core/u_decode/instruction[7] ), .Z(n7387)
         );
  AND U9661 ( .A(n7354), .B(n7389), .Z(n7386) );
  NANDN U9662 ( .B(n7356), .A(\u_a23_core/u_decode/instruction[5] ), .Z(n7389)
         );
  AND U9663 ( .A(n7390), .B(n7391), .Z(n7384) );
  NANDN U9664 ( .B(n7353), .A(\u_a23_core/rm_sel_nxt[3] ), .Z(n7391) );
  NANDN U9665 ( .B(n7346), .A(\u_a23_core/rm_sel_nxt[1] ), .Z(n7390) );
  NAND U9666 ( .A(n7392), .B(n7393), .Z(\u_a23_core/u_decode/imm32_nxt[28] )
         );
  AND U9667 ( .A(n7394), .B(n7395), .Z(n7393) );
  NANDN U9668 ( .B(n7388), .A(\u_a23_core/u_decode/instruction[6] ), .Z(n7395)
         );
  AND U9669 ( .A(n7354), .B(n7396), .Z(n7394) );
  NANDN U9670 ( .B(n7356), .A(\u_a23_core/u_decode/instruction[4] ), .Z(n7396)
         );
  AND U9671 ( .A(n7397), .B(n7398), .Z(n7392) );
  NANDN U9672 ( .B(n7353), .A(\u_a23_core/rm_sel_nxt[2] ), .Z(n7398) );
  NANDN U9673 ( .B(n7346), .A(\u_a23_core/rm_sel_nxt[0] ), .Z(n7397) );
  NAND U9674 ( .A(n7399), .B(n7400), .Z(\u_a23_core/u_decode/imm32_nxt[27] )
         );
  AND U9675 ( .A(n7401), .B(n7402), .Z(n7400) );
  NANDN U9676 ( .B(n7388), .A(\u_a23_core/u_decode/instruction[5] ), .Z(n7402)
         );
  AND U9677 ( .A(n7354), .B(n7403), .Z(n7401) );
  NANDN U9678 ( .B(n7356), .A(\u_a23_core/rm_sel_nxt[3] ), .Z(n7403) );
  AND U9679 ( .A(n7404), .B(n7405), .Z(n7399) );
  NANDN U9680 ( .B(n7406), .A(\u_a23_core/u_decode/instruction[7] ), .Z(n7405)
         );
  NANDN U9681 ( .B(n7353), .A(\u_a23_core/rm_sel_nxt[1] ), .Z(n7404) );
  NAND U9682 ( .A(n7407), .B(n7408), .Z(\u_a23_core/u_decode/imm32_nxt[26] )
         );
  AND U9683 ( .A(n7409), .B(n7410), .Z(n7408) );
  NANDN U9684 ( .B(n7388), .A(\u_a23_core/u_decode/instruction[4] ), .Z(n7410)
         );
  AND U9685 ( .A(n7354), .B(n7411), .Z(n7409) );
  NANDN U9686 ( .B(n7356), .A(\u_a23_core/rm_sel_nxt[2] ), .Z(n7411) );
  AND U9687 ( .A(n7412), .B(n7413), .Z(n7407) );
  NANDN U9688 ( .B(n7406), .A(\u_a23_core/u_decode/instruction[6] ), .Z(n7413)
         );
  NANDN U9689 ( .B(n7353), .A(\u_a23_core/rm_sel_nxt[0] ), .Z(n7412) );
  NAND U9690 ( .A(n7414), .B(n7415), .Z(\u_a23_core/u_decode/imm32_nxt[25] )
         );
  AND U9691 ( .A(n7416), .B(n7417), .Z(n7415) );
  NANDN U9692 ( .B(n7388), .A(\u_a23_core/rm_sel_nxt[3] ), .Z(n7417) );
  AND U9693 ( .A(n7354), .B(n7418), .Z(n7416) );
  NANDN U9694 ( .B(n7356), .A(\u_a23_core/rm_sel_nxt[1] ), .Z(n7418) );
  NANDN U9695 ( .B(n7419), .A(n7171), .Z(n7354) );
  AND U9696 ( .A(n7420), .B(n7421), .Z(n7414) );
  NANDN U9697 ( .B(n7406), .A(\u_a23_core/u_decode/instruction[5] ), .Z(n7421)
         );
  NANDN U9698 ( .B(n7422), .A(\u_a23_core/u_decode/instruction[7] ), .Z(n7420)
         );
  NAND U9699 ( .A(n7423), .B(n7424), .Z(\u_a23_core/u_decode/imm32_nxt[24] )
         );
  AND U9700 ( .A(n7425), .B(n7426), .Z(n7424) );
  NANDN U9701 ( .B(n7406), .A(\u_a23_core/u_decode/instruction[4] ), .Z(n7426)
         );
  AND U9702 ( .A(n7427), .B(n7428), .Z(n7425) );
  NANDN U9703 ( .B(n7356), .A(\u_a23_core/rm_sel_nxt[0] ), .Z(n7428) );
  NAND U9704 ( .A(n7429), .B(n7430), .Z(n7356) );
  AND U9705 ( .A(n7431), .B(n7378), .Z(n7429) );
  NANDN U9706 ( .B(n7388), .A(\u_a23_core/rm_sel_nxt[2] ), .Z(n7427) );
  AND U9707 ( .A(n7432), .B(n7433), .Z(n7423) );
  NANDN U9708 ( .B(n7422), .A(\u_a23_core/u_decode/instruction[6] ), .Z(n7433)
         );
  NAND U9709 ( .A(n7114), .B(n7372), .Z(n7432) );
  NAND U9710 ( .A(n7434), .B(n7435), .Z(\u_a23_core/u_decode/imm32_nxt[23] )
         );
  AND U9711 ( .A(n7436), .B(n7437), .Z(n7435) );
  NANDN U9712 ( .B(n7422), .A(\u_a23_core/u_decode/instruction[5] ), .Z(n7437)
         );
  AND U9713 ( .A(n7438), .B(n7439), .Z(n7436) );
  NANDN U9714 ( .B(n7388), .A(\u_a23_core/rm_sel_nxt[1] ), .Z(n7439) );
  NANDN U9715 ( .B(n7406), .A(\u_a23_core/rm_sel_nxt[3] ), .Z(n7438) );
  AND U9716 ( .A(n7440), .B(n7441), .Z(n7434) );
  NANDN U9717 ( .B(n7442), .A(\u_a23_core/u_decode/instruction[7] ), .Z(n7441)
         );
  NAND U9718 ( .A(n7163), .B(n7372), .Z(n7440) );
  NAND U9719 ( .A(n7443), .B(n7444), .Z(\u_a23_core/u_decode/imm32_nxt[22] )
         );
  AND U9720 ( .A(n7445), .B(n7446), .Z(n7444) );
  NANDN U9721 ( .B(n7422), .A(\u_a23_core/u_decode/instruction[4] ), .Z(n7446)
         );
  AND U9722 ( .A(n7447), .B(n7448), .Z(n7445) );
  NANDN U9723 ( .B(n7388), .A(\u_a23_core/rm_sel_nxt[0] ), .Z(n7448) );
  NAND U9724 ( .A(n7381), .B(n7449), .Z(n7388) );
  AND U9725 ( .A(n7430), .B(n7450), .Z(n7449) );
  NANDN U9726 ( .B(n7406), .A(\u_a23_core/rm_sel_nxt[2] ), .Z(n7447) );
  AND U9727 ( .A(n7451), .B(n7452), .Z(n7443) );
  NANDN U9728 ( .B(n7442), .A(\u_a23_core/u_decode/instruction[6] ), .Z(n7452)
         );
  NAND U9729 ( .A(n7135), .B(n7372), .Z(n7451) );
  NAND U9730 ( .A(n7453), .B(n7454), .Z(\u_a23_core/u_decode/imm32_nxt[21] )
         );
  AND U9731 ( .A(n7455), .B(n7456), .Z(n7454) );
  NANDN U9732 ( .B(n7442), .A(\u_a23_core/u_decode/instruction[5] ), .Z(n7456)
         );
  AND U9733 ( .A(n7457), .B(n7458), .Z(n7455) );
  NANDN U9734 ( .B(n7406), .A(\u_a23_core/rm_sel_nxt[1] ), .Z(n7458) );
  NANDN U9735 ( .B(n7422), .A(\u_a23_core/rm_sel_nxt[3] ), .Z(n7457) );
  AND U9736 ( .A(n7459), .B(n7460), .Z(n7453) );
  NANDN U9737 ( .B(n7461), .A(\u_a23_core/u_decode/instruction[7] ), .Z(n7460)
         );
  NAND U9738 ( .A(n7372), .B(n7170), .Z(n7459) );
  NAND U9739 ( .A(n7462), .B(n7463), .Z(\u_a23_core/u_decode/imm32_nxt[20] )
         );
  AND U9740 ( .A(n7464), .B(n7465), .Z(n7463) );
  NANDN U9741 ( .B(n7442), .A(\u_a23_core/u_decode/instruction[4] ), .Z(n7465)
         );
  AND U9742 ( .A(n7466), .B(n7467), .Z(n7464) );
  NANDN U9743 ( .B(n7406), .A(\u_a23_core/rm_sel_nxt[0] ), .Z(n7467) );
  NAND U9744 ( .A(n7468), .B(n7469), .Z(n7406) );
  NANDN U9745 ( .B(n7422), .A(\u_a23_core/rm_sel_nxt[2] ), .Z(n7466) );
  AND U9746 ( .A(n7470), .B(n7471), .Z(n7462) );
  NANDN U9747 ( .B(n7461), .A(\u_a23_core/u_decode/instruction[6] ), .Z(n7471)
         );
  NAND U9748 ( .A(n7372), .B(n7169), .Z(n7470) );
  NAND U9749 ( .A(n7472), .B(n7473), .Z(\u_a23_core/u_decode/imm32_nxt[1] ) );
  AND U9750 ( .A(n7474), .B(n7475), .Z(n7473) );
  NANDN U9751 ( .B(n7353), .A(\u_a23_core/u_decode/instruction[7] ), .Z(n7475)
         );
  NANDN U9752 ( .B(n7346), .A(\u_a23_core/u_decode/instruction[5] ), .Z(n7474)
         );
  AND U9753 ( .A(n7476), .B(n7477), .Z(n7472) );
  NANDN U9754 ( .B(n7327), .A(\u_a23_core/rm_sel_nxt[3] ), .Z(n7477) );
  NAND U9755 ( .A(\u_a23_core/rm_sel_nxt[1] ), .B(n7314), .Z(n7476) );
  NAND U9756 ( .A(n7478), .B(n7479), .Z(\u_a23_core/u_decode/imm32_nxt[19] )
         );
  AND U9757 ( .A(n7480), .B(n7481), .Z(n7479) );
  NANDN U9758 ( .B(n7461), .A(\u_a23_core/u_decode/instruction[5] ), .Z(n7481)
         );
  AND U9759 ( .A(n7482), .B(n7483), .Z(n7480) );
  NANDN U9760 ( .B(n7422), .A(\u_a23_core/rm_sel_nxt[1] ), .Z(n7483) );
  NANDN U9761 ( .B(n7442), .A(\u_a23_core/rm_sel_nxt[3] ), .Z(n7482) );
  AND U9762 ( .A(n7484), .B(n7485), .Z(n7478) );
  NANDN U9763 ( .B(n7486), .A(\u_a23_core/u_decode/instruction[7] ), .Z(n7485)
         );
  NAND U9764 ( .A(n7372), .B(n7168), .Z(n7484) );
  NAND U9765 ( .A(n7487), .B(n7488), .Z(\u_a23_core/u_decode/imm32_nxt[18] )
         );
  AND U9766 ( .A(n7489), .B(n7490), .Z(n7488) );
  NANDN U9767 ( .B(n7461), .A(\u_a23_core/u_decode/instruction[4] ), .Z(n7490)
         );
  AND U9768 ( .A(n7491), .B(n7492), .Z(n7489) );
  NANDN U9769 ( .B(n7422), .A(\u_a23_core/rm_sel_nxt[0] ), .Z(n7492) );
  NAND U9770 ( .A(n7469), .B(n7493), .Z(n7422) );
  ANDN U9771 ( .A(n7430), .B(n7494), .Z(n7469) );
  NANDN U9772 ( .B(n7442), .A(\u_a23_core/rm_sel_nxt[2] ), .Z(n7491) );
  AND U9773 ( .A(n7495), .B(n7496), .Z(n7487) );
  NANDN U9774 ( .B(n7486), .A(\u_a23_core/u_decode/instruction[6] ), .Z(n7496)
         );
  NAND U9775 ( .A(n7372), .B(n7166), .Z(n7495) );
  NAND U9776 ( .A(n7497), .B(n7498), .Z(\u_a23_core/u_decode/imm32_nxt[17] )
         );
  AND U9777 ( .A(n7499), .B(n7500), .Z(n7498) );
  NANDN U9778 ( .B(n7486), .A(\u_a23_core/u_decode/instruction[5] ), .Z(n7500)
         );
  AND U9779 ( .A(n7501), .B(n7502), .Z(n7499) );
  NANDN U9780 ( .B(n7442), .A(\u_a23_core/rm_sel_nxt[1] ), .Z(n7502) );
  NANDN U9781 ( .B(n7461), .A(\u_a23_core/rm_sel_nxt[3] ), .Z(n7501) );
  AND U9782 ( .A(n7503), .B(n7504), .Z(n7497) );
  NANDN U9783 ( .B(n7505), .A(\u_a23_core/u_decode/instruction[7] ), .Z(n7504)
         );
  NAND U9784 ( .A(n7258), .B(n7372), .Z(n7503) );
  NAND U9785 ( .A(n7506), .B(n7507), .Z(\u_a23_core/u_decode/imm32_nxt[16] )
         );
  AND U9786 ( .A(n7508), .B(n7509), .Z(n7507) );
  NANDN U9787 ( .B(n7486), .A(\u_a23_core/u_decode/instruction[4] ), .Z(n7509)
         );
  AND U9788 ( .A(n7510), .B(n7511), .Z(n7508) );
  NANDN U9789 ( .B(n7442), .A(\u_a23_core/rm_sel_nxt[0] ), .Z(n7511) );
  NANDN U9790 ( .B(n7512), .A(n7513), .Z(n7442) );
  NANDN U9791 ( .B(n7461), .A(\u_a23_core/rm_sel_nxt[2] ), .Z(n7510) );
  AND U9792 ( .A(n7514), .B(n7515), .Z(n7506) );
  NANDN U9793 ( .B(n7505), .A(\u_a23_core/u_decode/instruction[6] ), .Z(n7515)
         );
  NAND U9794 ( .A(n7249), .B(n7372), .Z(n7514) );
  NAND U9795 ( .A(n7516), .B(n7517), .Z(\u_a23_core/u_decode/imm32_nxt[15] )
         );
  AND U9796 ( .A(n7518), .B(n7519), .Z(n7517) );
  NANDN U9797 ( .B(n7299), .A(\u_a23_core/u_decode/instruction[7] ), .Z(n7519)
         );
  AND U9798 ( .A(n7520), .B(n7521), .Z(n7518) );
  NANDN U9799 ( .B(n7461), .A(\u_a23_core/rm_sel_nxt[1] ), .Z(n7521) );
  NANDN U9800 ( .B(n7486), .A(\u_a23_core/rm_sel_nxt[3] ), .Z(n7520) );
  AND U9801 ( .A(n7522), .B(n7523), .Z(n7516) );
  NANDN U9802 ( .B(n7505), .A(\u_a23_core/u_decode/instruction[5] ), .Z(n7523)
         );
  NAND U9803 ( .A(n7246), .B(n7372), .Z(n7522) );
  NAND U9804 ( .A(n7524), .B(n7525), .Z(\u_a23_core/u_decode/imm32_nxt[14] )
         );
  AND U9805 ( .A(n7526), .B(n7527), .Z(n7525) );
  NANDN U9806 ( .B(n7299), .A(\u_a23_core/u_decode/instruction[6] ), .Z(n7527)
         );
  AND U9807 ( .A(n7528), .B(n7529), .Z(n7526) );
  NANDN U9808 ( .B(n7461), .A(\u_a23_core/rm_sel_nxt[0] ), .Z(n7529) );
  NAND U9809 ( .A(n7513), .B(n7530), .Z(n7461) );
  NANDN U9810 ( .B(n7486), .A(\u_a23_core/rm_sel_nxt[2] ), .Z(n7528) );
  AND U9811 ( .A(n7531), .B(n7532), .Z(n7524) );
  NANDN U9812 ( .B(n7505), .A(\u_a23_core/u_decode/instruction[4] ), .Z(n7532)
         );
  NAND U9813 ( .A(n7237), .B(n7372), .Z(n7531) );
  NAND U9814 ( .A(n7533), .B(n7534), .Z(\u_a23_core/u_decode/imm32_nxt[13] )
         );
  AND U9815 ( .A(n7535), .B(n7536), .Z(n7534) );
  NANDN U9816 ( .B(n7299), .A(\u_a23_core/u_decode/instruction[5] ), .Z(n7536)
         );
  AND U9817 ( .A(n7537), .B(n7538), .Z(n7535) );
  NANDN U9818 ( .B(n7486), .A(\u_a23_core/rm_sel_nxt[1] ), .Z(n7538) );
  NANDN U9819 ( .B(n7296), .A(\u_a23_core/u_decode/instruction[7] ), .Z(n7537)
         );
  AND U9820 ( .A(n7539), .B(n7540), .Z(n7533) );
  NANDN U9821 ( .B(n7505), .A(\u_a23_core/rm_sel_nxt[3] ), .Z(n7540) );
  NAND U9822 ( .A(\u_a23_core/u_decode/instruction[11] ), .B(n7372), .Z(n7539)
         );
  NAND U9823 ( .A(n7541), .B(n7542), .Z(\u_a23_core/u_decode/imm32_nxt[12] )
         );
  AND U9824 ( .A(n7543), .B(n7544), .Z(n7542) );
  NANDN U9825 ( .B(n7299), .A(\u_a23_core/u_decode/instruction[4] ), .Z(n7544)
         );
  AND U9826 ( .A(n7545), .B(n7546), .Z(n7543) );
  NANDN U9827 ( .B(n7486), .A(\u_a23_core/rm_sel_nxt[0] ), .Z(n7546) );
  NANDN U9828 ( .B(n7547), .A(n7548), .Z(n7486) );
  ANDN U9829 ( .A(n7468), .B(n7549), .Z(n7548) );
  NANDN U9830 ( .B(n7296), .A(\u_a23_core/u_decode/instruction[6] ), .Z(n7545)
         );
  AND U9831 ( .A(n7550), .B(n7551), .Z(n7541) );
  NANDN U9832 ( .B(n7505), .A(\u_a23_core/rm_sel_nxt[2] ), .Z(n7551) );
  NAND U9833 ( .A(\u_a23_core/u_decode/instruction[10] ), .B(n7372), .Z(n7550)
         );
  NAND U9834 ( .A(n7552), .B(n7553), .Z(\u_a23_core/u_decode/imm32_nxt[11] )
         );
  AND U9835 ( .A(n7554), .B(n7555), .Z(n7553) );
  NANDN U9836 ( .B(n7299), .A(\u_a23_core/rm_sel_nxt[3] ), .Z(n7555) );
  AND U9837 ( .A(n7556), .B(n7557), .Z(n7554) );
  NANDN U9838 ( .B(n7296), .A(\u_a23_core/u_decode/instruction[5] ), .Z(n7557)
         );
  NANDN U9839 ( .B(n7292), .A(\u_a23_core/u_decode/instruction[7] ), .Z(n7556)
         );
  AND U9840 ( .A(n7558), .B(n7559), .Z(n7552) );
  NAND U9841 ( .A(\u_a23_core/u_decode/instruction[9] ), .B(n7372), .Z(n7559)
         );
  AND U9842 ( .A(n7560), .B(n7561), .Z(n7558) );
  NANDN U9843 ( .B(n7505), .A(\u_a23_core/rm_sel_nxt[1] ), .Z(n7561) );
  NAND U9844 ( .A(\u_a23_core/u_decode/instruction[11] ), .B(n7287), .Z(n7560)
         );
  NAND U9845 ( .A(n7562), .B(n7563), .Z(\u_a23_core/u_decode/imm32_nxt[10] )
         );
  AND U9846 ( .A(n7564), .B(n7565), .Z(n7563) );
  NANDN U9847 ( .B(n7299), .A(\u_a23_core/rm_sel_nxt[2] ), .Z(n7565) );
  NAND U9848 ( .A(n7378), .B(n7379), .Z(n7299) );
  AND U9849 ( .A(n7566), .B(n7567), .Z(n7564) );
  NANDN U9850 ( .B(n7296), .A(\u_a23_core/u_decode/instruction[4] ), .Z(n7567)
         );
  NAND U9851 ( .A(n7381), .B(n7379), .Z(n7296) );
  NANDN U9852 ( .B(n7292), .A(\u_a23_core/u_decode/instruction[6] ), .Z(n7566)
         );
  NAND U9853 ( .A(n7468), .B(n7379), .Z(n7292) );
  ANDN U9854 ( .A(n7513), .B(n7568), .Z(n7379) );
  AND U9855 ( .A(n7569), .B(n7570), .Z(n7562) );
  NAND U9856 ( .A(\u_a23_core/u_decode/instruction[8] ), .B(n7372), .Z(n7570)
         );
  AND U9857 ( .A(n7571), .B(n7572), .Z(n7569) );
  NANDN U9858 ( .B(n7505), .A(\u_a23_core/rm_sel_nxt[0] ), .Z(n7572) );
  NANDN U9859 ( .B(n7547), .A(n7573), .Z(n7505) );
  ANDN U9860 ( .A(\u_a23_core/u_decode/instruction[8] ), .B(n7549), .Z(n7573)
         );
  NANDN U9861 ( .B(n7530), .A(n7513), .Z(n7547) );
  NOR U9862 ( .A(n7494), .B(n7430), .Z(n7513) );
  ANDN U9863 ( .A(\u_a23_core/u_decode/instruction[10] ), .B(
        \u_a23_core/u_decode/instruction[11] ), .Z(n7430) );
  IV U9864 ( .A(n7450), .Z(n7494) );
  AND U9865 ( .A(n7431), .B(n7574), .Z(n7450) );
  ANDN U9866 ( .A(n7381), .B(\u_a23_core/u_decode/instruction[10] ), .Z(n7530)
         );
  NAND U9867 ( .A(\u_a23_core/u_decode/instruction[10] ), .B(n7287), .Z(n7571)
         );
  NAND U9868 ( .A(n7575), .B(n7576), .Z(\u_a23_core/u_decode/imm32_nxt[0] ) );
  AND U9869 ( .A(n7577), .B(n7578), .Z(n7576) );
  NANDN U9870 ( .B(n7353), .A(\u_a23_core/u_decode/instruction[6] ), .Z(n7578)
         );
  NAND U9871 ( .A(n7579), .B(n7493), .Z(n7353) );
  ANDN U9872 ( .A(\u_a23_core/u_decode/instruction[9] ), .B(n7580), .Z(n7493)
         );
  NANDN U9873 ( .B(n7346), .A(\u_a23_core/u_decode/instruction[4] ), .Z(n7577)
         );
  NAND U9874 ( .A(n7581), .B(n7431), .Z(n7346) );
  AND U9875 ( .A(n7582), .B(n7468), .Z(n7581) );
  AND U9876 ( .A(n7583), .B(n7584), .Z(n7575) );
  NANDN U9877 ( .B(n7327), .A(\u_a23_core/rm_sel_nxt[2] ), .Z(n7584) );
  NAND U9878 ( .A(n7381), .B(n7579), .Z(n7327) );
  AND U9879 ( .A(n7431), .B(n7582), .Z(n7579) );
  AND U9880 ( .A(n7585), .B(n7586), .Z(n7431) );
  AND U9881 ( .A(n7285), .B(n7419), .Z(n7585) );
  ANDN U9882 ( .A(\u_a23_core/u_decode/instruction[8] ), .B(
        \u_a23_core/u_decode/instruction[9] ), .Z(n7381) );
  NAND U9883 ( .A(\u_a23_core/rm_sel_nxt[0] ), .B(n7314), .Z(n7583) );
  NANDN U9884 ( .B(n7287), .A(n7587), .Z(n7314) );
  NAND U9885 ( .A(n7588), .B(n7589), .Z(n7587) );
  AND U9886 ( .A(n7214), .B(n7285), .Z(n7589) );
  AND U9887 ( .A(n7590), .B(n7419), .Z(n7588) );
  NAND U9888 ( .A(n7591), .B(n7165), .Z(
        \u_a23_core/u_decode/control_state_nxt[4] ) );
  ANDN U9889 ( .A(n7592), .B(n7158), .Z(n7591) );
  NAND U9890 ( .A(\u_a23_core/u_decode/control_state[4] ), .B(n7593), .Z(n7592) );
  NAND U9891 ( .A(n7594), .B(n7595), .Z(n7593) );
  NAND U9892 ( .A(n7596), .B(n7597), .Z(
        \u_a23_core/u_decode/control_state_nxt[3] ) );
  AND U9893 ( .A(n7598), .B(n7263), .Z(n7597) );
  NOR U9894 ( .A(n7599), .B(n7600), .Z(n7598) );
  AND U9895 ( .A(n7601), .B(n7602), .Z(n7596) );
  NAND U9896 ( .A(\u_a23_core/u_decode/control_state[3] ), .B(n7603), .Z(n7602) );
  NAND U9897 ( .A(n7604), .B(n7605), .Z(
        \u_a23_core/u_decode/control_state_nxt[2] ) );
  AND U9898 ( .A(n7606), .B(n7607), .Z(n7605) );
  NOR U9899 ( .A(n7608), .B(n7609), .Z(n7607) );
  AND U9900 ( .A(n7610), .B(n7611), .Z(n7606) );
  NAND U9901 ( .A(n7612), .B(n7613), .Z(n7611) );
  AND U9902 ( .A(\u_a23_core/multiply_function[1] ), .B(
        \u_a23_core/multiply_done ), .Z(n7613) );
  NAND U9903 ( .A(n7614), .B(n7615), .Z(n7610) );
  ANDN U9904 ( .A(n7285), .B(n7600), .Z(n7615) );
  AND U9905 ( .A(n7616), .B(n7129), .Z(n7614) );
  NANDN U9906 ( .B(n7617), .A(n7181), .Z(n7616) );
  AND U9907 ( .A(n7618), .B(n7619), .Z(n7604) );
  AND U9908 ( .A(n7620), .B(n7621), .Z(n7619) );
  NAND U9909 ( .A(\u_a23_core/u_decode/control_state[2] ), .B(n7603), .Z(n7621) );
  NAND U9910 ( .A(n7622), .B(n7623), .Z(n7620) );
  IV U9911 ( .A(n7263), .Z(n7622) );
  AND U9912 ( .A(n7601), .B(n7624), .Z(n7618) );
  NOR U9913 ( .A(n7625), .B(n7626), .Z(n7601) );
  NAND U9914 ( .A(n7627), .B(n7628), .Z(
        \u_a23_core/u_decode/control_state_nxt[1] ) );
  AND U9915 ( .A(n7629), .B(n7630), .Z(n7628) );
  NAND U9916 ( .A(\u_a23_core/u_decode/control_state[1] ), .B(n7603), .Z(n7630) );
  AND U9917 ( .A(n7631), .B(n7632), .Z(n7629) );
  IV U9918 ( .A(n7633), .Z(n7632) );
  NANDN U9919 ( .B(n7617), .A(n7599), .Z(n7631) );
  AND U9920 ( .A(n7634), .B(n7635), .Z(n7617) );
  NOR U9921 ( .A(\u_a23_core/u_decode/mtrans_num_registers[1] ), .B(
        \u_a23_core/u_decode/mtrans_num_registers[2] ), .Z(n7634) );
  ANDN U9922 ( .A(n7636), .B(n7637), .Z(n7627) );
  NAND U9923 ( .A(n7638), .B(n7639), .Z(
        \u_a23_core/u_decode/control_state_nxt[0] ) );
  AND U9924 ( .A(n7165), .B(n7640), .Z(n7639) );
  AND U9925 ( .A(n7641), .B(n7642), .Z(n7640) );
  NANDN U9926 ( .B(n7643), .A(n7599), .Z(n7642) );
  AND U9927 ( .A(n7262), .B(n7644), .Z(n7165) );
  ANDN U9928 ( .A(n7645), .B(n7646), .Z(n7638) );
  MUX U9929 ( .IN0(n7647), .IN1(n7603), .SEL(
        \u_a23_core/u_decode/control_state[0] ), .F(n7646) );
  NAND U9930 ( .A(n7648), .B(n7595), .Z(n7603) );
  NAND U9931 ( .A(n7649), .B(n7650), .Z(n7595) );
  AND U9932 ( .A(n7651), .B(n7652), .Z(n7650) );
  AND U9933 ( .A(n7653), .B(n7654), .Z(n7652) );
  ANDN U9934 ( .A(n7277), .B(n7655), .Z(n7653) );
  AND U9935 ( .A(n7656), .B(n7263), .Z(n7651) );
  ANDN U9936 ( .A(n7644), .B(n7608), .Z(n7656) );
  NOR U9937 ( .A(\u_a23_core/u_decode/control_state[1] ), .B(n7657), .Z(n7608)
         );
  AND U9938 ( .A(n7658), .B(n7659), .Z(n7649) );
  ANDN U9939 ( .A(n7164), .B(n7625), .Z(n7659) );
  AND U9940 ( .A(n7139), .B(n7594), .Z(n7164) );
  NOR U9941 ( .A(n7609), .B(n7626), .Z(n7658) );
  ANDN U9942 ( .A(n7660), .B(n7643), .Z(n7626) );
  NAND U9943 ( .A(n7661), .B(n7662), .Z(n7643) );
  ANDN U9944 ( .A(n7635), .B(\u_a23_core/u_decode/mtrans_num_registers[2] ), 
        .Z(n7662) );
  NOR U9945 ( .A(\u_a23_core/u_decode/mtrans_num_registers[3] ), .B(
        \u_a23_core/u_decode/mtrans_num_registers[4] ), .Z(n7635) );
  ANDN U9946 ( .A(\u_a23_core/u_decode/mtrans_num_registers[0] ), .B(
        \u_a23_core/u_decode/mtrans_num_registers[1] ), .Z(n7661) );
  ANDN U9947 ( .A(n7663), .B(n7657), .Z(n7609) );
  NAND U9948 ( .A(n6747), .B(n7612), .Z(n7648) );
  IV U9949 ( .A(\u_a23_core/multiply_done ), .Z(n6747) );
  AND U9950 ( .A(n7664), .B(n7665), .Z(n7647) );
  ANDN U9951 ( .A(n7624), .B(n7637), .Z(n7645) );
  NAND U9952 ( .A(n7666), .B(n7667), .Z(n7637) );
  NAND U9953 ( .A(n7612), .B(n7668), .Z(n7667) );
  AND U9954 ( .A(n6742), .B(\u_a23_core/multiply_done ), .Z(n7668) );
  IV U9955 ( .A(\u_a23_core/multiply_function[1] ), .Z(n6742) );
  IV U9956 ( .A(n7594), .Z(n7612) );
  OR U9957 ( .A(n7623), .B(n7263), .Z(n7666) );
  AND U9958 ( .A(n7669), .B(n7670), .Z(n7623) );
  AND U9959 ( .A(n7671), .B(n7672), .Z(n7670) );
  AND U9960 ( .A(n7673), .B(n7674), .Z(n7672) );
  NOR U9961 ( .A(n7182), .B(n7189), .Z(n7674) );
  NOR U9962 ( .A(n7675), .B(n7676), .Z(n7189) );
  ANDN U9963 ( .A(\u_a23_core/rm_sel_nxt[1] ), .B(n7677), .Z(n7182) );
  NOR U9964 ( .A(n7197), .B(n7217), .Z(n7673) );
  NOR U9965 ( .A(n7580), .B(\u_a23_core/u_decode/N298 ), .Z(n7217) );
  NOR U9966 ( .A(n7120), .B(n7678), .Z(n7197) );
  ANDN U9967 ( .A(n7679), .B(n7240), .Z(n7671) );
  NOR U9968 ( .A(n7680), .B(n7681), .Z(n7240) );
  NOR U9969 ( .A(n7229), .B(n7232), .Z(n7679) );
  AND U9970 ( .A(n7682), .B(\u_a23_core/u_decode/instruction[11] ), .Z(n7232)
         );
  NAND U9971 ( .A(n7568), .B(n7683), .Z(n7682) );
  NOR U9972 ( .A(n7568), .B(n7683), .Z(n7229) );
  AND U9973 ( .A(n7684), .B(n7685), .Z(n7669) );
  AND U9974 ( .A(n7686), .B(n7687), .Z(n7685) );
  NOR U9975 ( .A(n7243), .B(n7255), .Z(n7687) );
  AND U9976 ( .A(n7688), .B(n7258), .Z(n7255) );
  NAND U9977 ( .A(n7689), .B(n7252), .Z(n7688) );
  AND U9978 ( .A(n7690), .B(n7246), .Z(n7243) );
  NAND U9979 ( .A(n7680), .B(n7681), .Z(n7690) );
  AND U9980 ( .A(n7691), .B(n7692), .Z(n7686) );
  NAND U9981 ( .A(\u_a23_core/u_decode/instruction[7] ), .B(n7693), .Z(n7692)
         );
  NAND U9982 ( .A(n7694), .B(n7213), .Z(n7693) );
  NAND U9983 ( .A(n7695), .B(n7696), .Z(n7691) );
  NAND U9984 ( .A(n7697), .B(n7213), .Z(n7696) );
  NAND U9985 ( .A(\u_a23_core/u_decode/instruction[5] ), .B(
        \u_a23_core/u_decode/instruction[6] ), .Z(n7697) );
  IV U9986 ( .A(n7694), .Z(n7695) );
  AND U9987 ( .A(n7698), .B(n7699), .Z(n7684) );
  NAND U9988 ( .A(\u_a23_core/rm_sel_nxt[3] ), .B(n7194), .Z(n7699) );
  NAND U9989 ( .A(n7675), .B(n7676), .Z(n7194) );
  AND U9990 ( .A(n7700), .B(n7701), .Z(n7698) );
  OR U9991 ( .A(n7252), .B(n7689), .Z(n7701) );
  AND U9992 ( .A(n7702), .B(n7681), .Z(n7252) );
  ANDN U9993 ( .A(n7683), .B(n7549), .Z(n7681) );
  NAND U9994 ( .A(n7568), .B(n7512), .Z(n7549) );
  NAND U9995 ( .A(n7378), .B(n7703), .Z(n7512) );
  AND U9996 ( .A(n7568), .B(\u_a23_core/u_decode/instruction[11] ), .Z(n7703)
         );
  ANDN U9997 ( .A(n7224), .B(n7468), .Z(n7683) );
  AND U9998 ( .A(n7704), .B(n7680), .Z(n7702) );
  OR U9999 ( .A(n7224), .B(n7705), .Z(n7700) );
  IV U10000 ( .A(\u_a23_core/u_decode/instruction[9] ), .Z(n7705) );
  ANDN U10001 ( .A(\u_a23_core/u_decode/N298 ), .B(
        \u_a23_core/u_decode/instruction[8] ), .Z(n7224) );
  ANDN U10002 ( .A(n7706), .B(n16637), .Z(n7624) );
  NANDN U10003 ( .B(n7600), .A(n7707), .Z(n7706) );
  NANDN U10004 ( .B(n7655), .A(n7654), .Z(n7707) );
  AND U10005 ( .A(\u_a23_core/u_decode/pc_wen_nxt ), .B(
        \u_a23_core/u_decode/pc_sel_nxt[0] ), .Z(n7600) );
  NAND U10006 ( .A(n7708), .B(n7709), .Z(\u_a23_core/u_decode/pc_sel_nxt[0] )
         );
  ANDN U10007 ( .A(n7710), .B(\u_a23_core/u_decode/pc_sel_nxt[1] ), .Z(n7708)
         );
  NAND U10008 ( .A(n7711), .B(n7712), .Z(n7710) );
  AND U10009 ( .A(n7713), .B(n7169), .Z(n7712) );
  AND U10010 ( .A(n7168), .B(\u_a23_core/rn_sel_nxt[0] ), .Z(n7713) );
  ANDN U10011 ( .A(n7170), .B(n7714), .Z(n7711) );
  AND U10012 ( .A(n7715), .B(n7716), .Z(\u_a23_core/u_decode/pc_wen_nxt ) );
  AND U10013 ( .A(n7717), .B(n7718), .Z(n7716) );
  NAND U10014 ( .A(n7129), .B(n7719), .Z(n7718) );
  NAND U10015 ( .A(n7285), .B(n7586), .Z(n7719) );
  AND U10016 ( .A(n7262), .B(n7594), .Z(n7717) );
  NANDN U10017 ( .B(n7720), .A(n7721), .Z(n7262) );
  AND U10018 ( .A(n7722), .B(n7723), .Z(n7721) );
  AND U10019 ( .A(n7107), .B(n7636), .Z(n7715) );
  AND U10020 ( .A(n7724), .B(n7633), .Z(
        \u_a23_core/u_decode/byte_enable_sel_nxt[0] ) );
  AND U10021 ( .A(n7114), .B(n7105), .Z(n7724) );
  NAND U10022 ( .A(n7725), .B(n7726), .Z(
        \u_a23_core/u_decode/barrel_shift_function_nxt[1] ) );
  NAND U10023 ( .A(\u_a23_core/u_decode/instruction[6] ), .B(n7727), .Z(n7725)
         );
  NAND U10024 ( .A(n7728), .B(n7726), .Z(
        \u_a23_core/u_decode/barrel_shift_function_nxt[0] ) );
  NAND U10025 ( .A(n7729), .B(n7730), .Z(n7726) );
  OR U10026 ( .A(\u_a23_core/u_execute/address_plus4[0] ), .B(
        \u_a23_core/execute_address[1] ), .Z(n7730) );
  NAND U10027 ( .A(\u_a23_core/u_decode/instruction[5] ), .B(n7727), .Z(n7728)
         );
  OR U10028 ( .A(n7731), .B(n7732), .Z(n7727) );
  NANDN U10029 ( .B(n7731), .A(n7733), .Z(
        \u_a23_core/u_decode/barrel_shift_data_sel_nxt[1] ) );
  NAND U10030 ( .A(n7172), .B(n7633), .Z(n7733) );
  NAND U10031 ( .A(n7734), .B(n7735), .Z(
        \u_a23_core/u_decode/barrel_shift_data_sel_nxt[0] ) );
  ANDN U10032 ( .A(n7736), .B(n7655), .Z(n7735) );
  NOR U10033 ( .A(n7729), .B(n7737), .Z(n7734) );
  NAND U10034 ( .A(n7738), .B(n7739), .Z(
        \u_a23_core/u_decode/barrel_shift_amount_sel_nxt[1] ) );
  NAND U10035 ( .A(n7120), .B(n7731), .Z(n7739) );
  ANDN U10036 ( .A(n7740), .B(n7732), .Z(n7738) );
  AND U10037 ( .A(n7741), .B(n7633), .Z(n7732) );
  AND U10038 ( .A(n7172), .B(n7742), .Z(n7741) );
  IV U10039 ( .A(n7122), .Z(n7742) );
  ANDN U10040 ( .A(n7590), .B(\u_a23_core/u_decode/instruction[7] ), .Z(n7122)
         );
  NAND U10041 ( .A(n7740), .B(n7743), .Z(
        \u_a23_core/u_decode/barrel_shift_amount_sel_nxt[0] ) );
  NAND U10042 ( .A(\u_a23_core/u_decode/instruction[4] ), .B(n7731), .Z(n7743)
         );
  ANDN U10043 ( .A(n7109), .B(n7172), .Z(n7731) );
  AND U10044 ( .A(n7744), .B(n7745), .Z(
        \u_a23_core/u_decode/alu_function_nxt[8] ) );
  AND U10045 ( .A(n7163), .B(n7746), .Z(n7745) );
  NAND U10046 ( .A(n7747), .B(n7748), .Z(
        \u_a23_core/u_decode/alu_function_nxt[7] ) );
  NAND U10047 ( .A(n7109), .B(n7749), .Z(n7748) );
  AND U10048 ( .A(n7750), .B(n7751), .Z(n7747) );
  NAND U10049 ( .A(n7752), .B(n7744), .Z(n7751) );
  NAND U10050 ( .A(n7753), .B(n7106), .Z(n7750) );
  AND U10051 ( .A(n7754), .B(n7109), .Z(
        \u_a23_core/u_decode/alu_function_nxt[6] ) );
  NOR U10052 ( .A(n7755), .B(n7113), .Z(n7754) );
  AND U10053 ( .A(n7756), .B(n7753), .Z(
        \u_a23_core/u_decode/alu_function_nxt[5] ) );
  NANDN U10054 ( .B(n7106), .A(n7757), .Z(n7756) );
  NAND U10055 ( .A(n7758), .B(n7744), .Z(n7757) );
  NAND U10056 ( .A(n7163), .B(n7142), .Z(n7758) );
  AND U10057 ( .A(n7759), .B(n7109), .Z(
        \u_a23_core/u_decode/alu_function_nxt[4] ) );
  NAND U10058 ( .A(n7116), .B(n7760), .Z(n7759) );
  NAND U10059 ( .A(n7753), .B(n7761), .Z(n7760) );
  MUX U10060 ( .IN0(n7762), .IN1(n7763), .SEL(n7753), .F(
        \u_a23_core/u_decode/alu_function_nxt[3] ) );
  AND U10061 ( .A(n7755), .B(n7109), .Z(n7763) );
  AND U10062 ( .A(n7744), .B(n7764), .Z(n7762) );
  ANDN U10063 ( .A(n7114), .B(n7138), .Z(n7744) );
  NANDN U10064 ( .B(\u_a23_core/u_decode/alu_function_nxt[2] ), .A(n7765), .Z(
        \u_a23_core/u_decode/alu_function_nxt[1] ) );
  AND U10065 ( .A(n7766), .B(n7109), .Z(
        \u_a23_core/u_decode/alu_function_nxt[2] ) );
  NAND U10066 ( .A(n7767), .B(n7768), .Z(n7766) );
  NAND U10067 ( .A(n7761), .B(n7769), .Z(n7768) );
  AND U10068 ( .A(n7163), .B(n7753), .Z(n7769) );
  NAND U10069 ( .A(n7770), .B(n7764), .Z(n7767) );
  AND U10070 ( .A(n7171), .B(n7761), .Z(n7770) );
  NAND U10071 ( .A(n7771), .B(n7772), .Z(
        \u_a23_core/u_decode/alu_function_nxt[0] ) );
  NOR U10072 ( .A(n7106), .B(\u_a23_core/u_decode/pc_sel_nxt[1] ), .Z(n7772)
         );
  ANDN U10073 ( .A(n7372), .B(n7277), .Z(\u_a23_core/u_decode/pc_sel_nxt[1] )
         );
  AND U10074 ( .A(n7765), .B(n7773), .Z(n7771) );
  NAND U10075 ( .A(n7109), .B(n7774), .Z(n7773) );
  OR U10076 ( .A(n7749), .B(n7123), .Z(n7774) );
  NAND U10077 ( .A(n7775), .B(n7776), .Z(n7123) );
  NAND U10078 ( .A(n7163), .B(n7777), .Z(n7776) );
  NAND U10079 ( .A(n7778), .B(n7113), .Z(n7777) );
  NAND U10080 ( .A(n7171), .B(n7746), .Z(n7113) );
  NAND U10081 ( .A(n7114), .B(n7779), .Z(n7778) );
  NAND U10082 ( .A(n7171), .B(n7755), .Z(n7775) );
  AND U10083 ( .A(n7780), .B(n7761), .Z(n7755) );
  AND U10084 ( .A(n7781), .B(n7114), .Z(n7749) );
  NAND U10085 ( .A(n7142), .B(n7782), .Z(n7781) );
  NAND U10086 ( .A(n7753), .B(n7780), .Z(n7782) );
  NAND U10087 ( .A(n7114), .B(n7729), .Z(n7765) );
  NAND U10088 ( .A(n7783), .B(n7107), .Z(
        \u_a23_core/u_decode/address_sel_nxt[2] ) );
  AND U10089 ( .A(n7784), .B(n7785), .Z(n7783) );
  NAND U10090 ( .A(n7746), .B(n7633), .Z(n7785) );
  ANDN U10091 ( .A(n7287), .B(n7277), .Z(n7633) );
  NANDN U10092 ( .B(n7779), .A(n7599), .Z(n7784) );
  NAND U10093 ( .A(n7786), .B(n7636), .Z(
        \u_a23_core/u_decode/address_sel_nxt[1] ) );
  AND U10094 ( .A(n7787), .B(n7594), .Z(n7786) );
  NAND U10095 ( .A(n7788), .B(n7599), .Z(n7787) );
  AND U10096 ( .A(n7181), .B(n7129), .Z(n7599) );
  NAND U10097 ( .A(n7116), .B(n7789), .Z(n7788) );
  NAND U10098 ( .A(n7753), .B(n7746), .Z(n7789) );
  IV U10099 ( .A(n7752), .Z(n7116) );
  ANDN U10100 ( .A(n7171), .B(n7746), .Z(n7752) );
  NAND U10101 ( .A(n7790), .B(n7791), .Z(
        \u_a23_core/u_decode/address_sel_nxt[0] ) );
  AND U10102 ( .A(n7107), .B(n7792), .Z(n7791) );
  AND U10103 ( .A(n7793), .B(n7594), .Z(n7792) );
  NANDN U10104 ( .B(n7720), .A(n7794), .Z(n7594) );
  AND U10105 ( .A(n7723), .B(\u_a23_core/u_decode/control_state[0] ), .Z(n7794) );
  NAND U10106 ( .A(n7142), .B(n7106), .Z(n7793) );
  NOR U10107 ( .A(n7277), .B(n7586), .Z(n7106) );
  ANDN U10108 ( .A(n7214), .B(n7287), .Z(n7586) );
  ANDN U10109 ( .A(n7263), .B(n7660), .Z(n7107) );
  NAND U10110 ( .A(n7795), .B(n7665), .Z(n7263) );
  ANDN U10111 ( .A(n7722), .B(n7664), .Z(n7795) );
  AND U10112 ( .A(n7636), .B(n7709), .Z(n7790) );
  AND U10113 ( .A(n7796), .B(n7140), .Z(n7709) );
  NAND U10114 ( .A(n7797), .B(n7798), .Z(n7140) );
  AND U10115 ( .A(\u_a23_core/u_decode/mtrans_reg_d2[0] ), .B(n7799), .Z(n7798) );
  AND U10116 ( .A(n7655), .B(n7135), .Z(n7799) );
  AND U10117 ( .A(\u_a23_core/u_decode/mtrans_reg_d2[3] ), .B(n7800), .Z(n7797) );
  AND U10118 ( .A(\u_a23_core/u_decode/mtrans_reg_d2[1] ), .B(
        \u_a23_core/u_decode/mtrans_reg_d2[2] ), .Z(n7800) );
  NAND U10119 ( .A(n7801), .B(n7133), .Z(n7796) );
  AND U10120 ( .A(n7802), .B(n7803), .Z(n7133) );
  AND U10121 ( .A(n7237), .B(n7249), .Z(n7803) );
  AND U10122 ( .A(n7246), .B(n7258), .Z(n7802) );
  NAND U10123 ( .A(n7740), .B(n7804), .Z(n7801) );
  AND U10124 ( .A(n7260), .B(n7805), .Z(n7636) );
  ANDN U10125 ( .A(n7644), .B(n7737), .Z(n7805) );
  NANDN U10126 ( .B(n7806), .A(n7807), .Z(n7644) );
  ANDN U10127 ( .A(n7722), .B(n7808), .Z(n7807) );
  ANDN U10128 ( .A(n7641), .B(n7625), .Z(n7260) );
  ANDN U10129 ( .A(\u_a23_core/u_decode/control_state[0] ), .B(n7809), .Z(
        n7625) );
  NANDN U10130 ( .B(n7810), .A(n7811), .Z(n7641) );
  AND U10131 ( .A(n7722), .B(n7663), .Z(n7811) );
  NAND U10132 ( .A(n7812), .B(n7813), .Z(\u_a23_core/u_decode/N524 ) );
  NAND U10133 ( .A(\u_a23_core/u_decode/instruction[9] ), .B(n7814), .Z(n7813)
         );
  NAND U10134 ( .A(\u_a23_core/u_decode/instruction[7] ), .B(
        \u_a23_core/u_decode/instruction[8] ), .Z(n7812) );
  XOR U10135 ( .A(n7814), .B(\u_a23_core/u_decode/instruction[9] ), .Z(
        \u_a23_core/u_decode/N523 ) );
  XNOR U10136 ( .A(\u_a23_core/u_decode/instruction[8] ), .B(n7815), .Z(n7814)
         );
  NANDN U10137 ( .B(n7816), .A(n7817), .Z(\u_a23_core/u_decode/N521 ) );
  NAND U10138 ( .A(n7574), .B(n7237), .Z(n7817) );
  XNOR U10139 ( .A(n7818), .B(n7237), .Z(\u_a23_core/u_decode/N520 ) );
  NANDN U10140 ( .B(n7816), .A(n7574), .Z(n7818) );
  ANDN U10141 ( .A(\u_a23_core/u_decode/instruction[10] ), .B(n7819), .Z(n7816) );
  NAND U10142 ( .A(n7820), .B(n7821), .Z(\u_a23_core/u_decode/N519 ) );
  NAND U10143 ( .A(n7258), .B(n7822), .Z(n7821) );
  NAND U10144 ( .A(n7249), .B(n7246), .Z(n7820) );
  XOR U10145 ( .A(n7822), .B(n7258), .Z(\u_a23_core/u_decode/N518 ) );
  XNOR U10146 ( .A(n7246), .B(n7689), .Z(n7822) );
  AND U10147 ( .A(n7147), .B(n7150), .Z(\u_a23_core/u_decode/N1089 ) );
  NOR U10148 ( .A(n7152), .B(n7149), .Z(n7150) );
  NAND U10149 ( .A(n7823), .B(n7824), .Z(n7149) );
  AND U10150 ( .A(n7825), .B(n7826), .Z(n7824) );
  NAND U10151 ( .A(n7827), .B(n7828), .Z(n7826) );
  AND U10152 ( .A(n7829), .B(n7740), .Z(n7827) );
  NAND U10153 ( .A(n7830), .B(n7831), .Z(n7829) );
  NANDN U10154 ( .B(n7832), .A(\u_a23_core/rn_sel_nxt[2] ), .Z(n7831) );
  NAND U10155 ( .A(n7833), .B(n7834), .Z(n7830) );
  NANDN U10156 ( .B(n7714), .A(n7835), .Z(n7834) );
  AND U10157 ( .A(n7836), .B(n7837), .Z(n7833) );
  NANDN U10158 ( .B(n7804), .A(n7689), .Z(n7837) );
  IV U10159 ( .A(n7249), .Z(n7689) );
  NAND U10160 ( .A(n7838), .B(n7839), .Z(n7825) );
  AND U10161 ( .A(n7169), .B(n16637), .Z(n7839) );
  AND U10162 ( .A(n7840), .B(n7841), .Z(n7823) );
  NAND U10163 ( .A(\u_a23_core/u_decode/mtrans_reg_d2[2] ), .B(n7842), .Z(
        n7841) );
  NANDN U10164 ( .B(n7843), .A(n7249), .Z(n7840) );
  NAND U10165 ( .A(n7844), .B(n7845), .Z(n7152) );
  AND U10166 ( .A(n7846), .B(n7847), .Z(n7845) );
  NAND U10167 ( .A(n7848), .B(n7828), .Z(n7847) );
  AND U10168 ( .A(n7849), .B(n7850), .Z(n7828) );
  ANDN U10169 ( .A(n7851), .B(n7852), .Z(n7849) );
  AND U10170 ( .A(n7853), .B(n7740), .Z(n7848) );
  IV U10171 ( .A(n7729), .Z(n7740) );
  NAND U10172 ( .A(n7854), .B(n7855), .Z(n7853) );
  NANDN U10173 ( .B(n7832), .A(\u_a23_core/rn_sel_nxt[3] ), .Z(n7855) );
  NAND U10174 ( .A(n7856), .B(n7857), .Z(n7854) );
  NANDN U10175 ( .B(n7714), .A(n7858), .Z(n7857) );
  AND U10176 ( .A(n7836), .B(n7859), .Z(n7856) );
  NANDN U10177 ( .B(n7804), .A(n7860), .Z(n7859) );
  IV U10178 ( .A(n7258), .Z(n7860) );
  NAND U10179 ( .A(n7838), .B(n7861), .Z(n7846) );
  AND U10180 ( .A(n7170), .B(n16637), .Z(n7861) );
  AND U10181 ( .A(n7862), .B(n7863), .Z(n7844) );
  NAND U10182 ( .A(n7842), .B(\u_a23_core/u_decode/mtrans_reg_d2[3] ), .Z(
        n7863) );
  NANDN U10183 ( .B(n7852), .A(n7864), .Z(n7842) );
  NANDN U10184 ( .B(n7843), .A(n7258), .Z(n7862) );
  NOR U10185 ( .A(n7729), .B(n7865), .Z(n7843) );
  NOR U10186 ( .A(n7154), .B(n7155), .Z(n7147) );
  NAND U10187 ( .A(n7866), .B(n7867), .Z(n7155) );
  AND U10188 ( .A(n7868), .B(n7869), .Z(n7867) );
  NAND U10189 ( .A(n7838), .B(n7870), .Z(n7869) );
  AND U10190 ( .A(n7168), .B(n16637), .Z(n7870) );
  NAND U10191 ( .A(n7871), .B(n7872), .Z(n7868) );
  AND U10192 ( .A(n7873), .B(n7874), .Z(n7872) );
  NAND U10193 ( .A(n7875), .B(n7876), .Z(n7874) );
  NAND U10194 ( .A(n7877), .B(n7878), .Z(n7876) );
  NANDN U10195 ( .B(n7714), .A(n7879), .Z(n7878) );
  NANDN U10196 ( .B(n7880), .A(n7129), .Z(n7714) );
  AND U10197 ( .A(n7836), .B(n7881), .Z(n7877) );
  NANDN U10198 ( .B(n7804), .A(n7704), .Z(n7881) );
  OR U10199 ( .A(n7779), .B(n7138), .Z(n7804) );
  IV U10200 ( .A(n7109), .Z(n7138) );
  ANDN U10201 ( .A(n7134), .B(n7277), .Z(n7109) );
  OR U10202 ( .A(n7832), .B(n7277), .Z(n7836) );
  IV U10203 ( .A(n7129), .Z(n7277) );
  NANDN U10204 ( .B(n7832), .A(\u_a23_core/rn_sel_nxt[1] ), .Z(n7875) );
  AND U10205 ( .A(n7851), .B(n7882), .Z(n7873) );
  NAND U10206 ( .A(n7729), .B(n7704), .Z(n7882) );
  AND U10207 ( .A(n7850), .B(n7883), .Z(n7871) );
  NANDN U10208 ( .B(\u_a23_core/u_decode/mtrans_reg_d2[1] ), .A(n7852), .Z(
        n7883) );
  AND U10209 ( .A(n7884), .B(n7885), .Z(n7866) );
  NAND U10210 ( .A(n7246), .B(n7865), .Z(n7885) );
  NANDN U10211 ( .B(n7864), .A(\u_a23_core/u_decode/mtrans_reg_d2[1] ), .Z(
        n7884) );
  NAND U10212 ( .A(n7886), .B(n7887), .Z(n7154) );
  AND U10213 ( .A(n7888), .B(n7889), .Z(n7887) );
  NAND U10214 ( .A(n7838), .B(n7890), .Z(n7889) );
  AND U10215 ( .A(n7166), .B(n16637), .Z(n7890) );
  NAND U10216 ( .A(n7891), .B(n7892), .Z(n7888) );
  AND U10217 ( .A(n7893), .B(n7894), .Z(n7892) );
  NAND U10218 ( .A(n7129), .B(n7895), .Z(n7894) );
  MUX U10219 ( .IN0(n7896), .IN1(n7897), .SEL(n7832), .F(n7895) );
  NAND U10220 ( .A(n7163), .B(n7181), .Z(n7832) );
  NAND U10221 ( .A(n7898), .B(n7899), .Z(n7897) );
  NAND U10222 ( .A(n7680), .B(n7900), .Z(n7899) );
  ANDN U10223 ( .A(n7134), .B(n7779), .Z(n7900) );
  AND U10224 ( .A(n7753), .B(n7142), .Z(n7779) );
  AND U10225 ( .A(n7901), .B(n7902), .Z(n7898) );
  NAND U10226 ( .A(n7142), .B(n7372), .Z(n7902) );
  IV U10227 ( .A(n7419), .Z(n7372) );
  NANDN U10228 ( .B(n7880), .A(n7896), .Z(n7901) );
  NANDN U10229 ( .B(n7764), .A(n7287), .Z(n7880) );
  AND U10230 ( .A(n7851), .B(n7903), .Z(n7893) );
  NAND U10231 ( .A(n7729), .B(n7680), .Z(n7903) );
  AND U10232 ( .A(n7904), .B(n7905), .Z(n7729) );
  IV U10233 ( .A(n7654), .Z(n7905) );
  NANDN U10234 ( .B(n7810), .A(n7906), .Z(n7654) );
  AND U10235 ( .A(n7663), .B(\u_a23_core/u_decode/control_state[0] ), .Z(n7906) );
  AND U10236 ( .A(n7135), .B(n7287), .Z(n7904) );
  AND U10237 ( .A(n7907), .B(n7908), .Z(n7287) );
  AND U10238 ( .A(n7909), .B(n7910), .Z(n7907) );
  AND U10239 ( .A(n7850), .B(n7911), .Z(n7891) );
  NANDN U10240 ( .B(\u_a23_core/u_decode/mtrans_reg_d2[0] ), .A(n7852), .Z(
        n7911) );
  ANDN U10241 ( .A(n7660), .B(n7105), .Z(n7852) );
  IV U10242 ( .A(n7736), .Z(n7660) );
  OR U10243 ( .A(n7664), .B(n7657), .Z(n7736) );
  NAND U10244 ( .A(\u_a23_core/u_decode/control_state[0] ), .B(n7665), .Z(
        n7657) );
  AND U10245 ( .A(n7912), .B(n7806), .Z(n7665) );
  NAND U10246 ( .A(\u_a23_core/u_decode/control_state[1] ), .B(
        \u_a23_core/u_decode/control_state[3] ), .Z(n7664) );
  ANDN U10247 ( .A(n7913), .B(n16637), .Z(n7850) );
  NAND U10248 ( .A(n7135), .B(n7655), .Z(n7913) );
  AND U10249 ( .A(n7914), .B(n7915), .Z(n7886) );
  NAND U10250 ( .A(n7237), .B(n7865), .Z(n7915) );
  ANDN U10251 ( .A(n16637), .B(n7838), .Z(n7865) );
  NANDN U10252 ( .B(n7864), .A(\u_a23_core/u_decode/mtrans_reg_d2[0] ), .Z(
        n7914) );
  ANDN U10253 ( .A(n7851), .B(n7655), .Z(n7864) );
  AND U10254 ( .A(n7916), .B(\u_a23_core/u_decode/control_state[3] ), .Z(n7655) );
  ANDN U10255 ( .A(n7722), .B(n7810), .Z(n7916) );
  NANDN U10256 ( .B(n7105), .A(n7737), .Z(n7851) );
  NOR U10257 ( .A(\u_a23_core/u_decode/control_state[0] ), .B(n7809), .Z(n7737) );
  NAND U10258 ( .A(n7917), .B(n7918), .Z(n7809) );
  AND U10259 ( .A(n7723), .B(n7806), .Z(n7918) );
  AND U10260 ( .A(\u_a23_core/u_decode/control_state[2] ), .B(
        \u_a23_core/u_decode/control_state[3] ), .Z(n7917) );
  IV U10261 ( .A(n7858), .Z(\u_a23_core/rn_sel_nxt[3] ) );
  ANDN U10262 ( .A(n7419), .B(n7170), .Z(n7858) );
  NAND U10263 ( .A(n7919), .B(n7920), .Z(n7170) );
  NANDN U10264 ( .B(n7270), .A(\u_a23_core/u_decode/pre_fetch_instruction[19] ), .Z(n7920) );
  AND U10265 ( .A(n7921), .B(n7922), .Z(n7919) );
  NANDN U10266 ( .B(n7269), .A(\u_a23_core/read_data_s2[19] ), .Z(n7922) );
  NAND U10267 ( .A(n7283), .B(
        \u_a23_core/u_decode/saved_current_instruction[19] ), .Z(n7921) );
  IV U10268 ( .A(n7835), .Z(\u_a23_core/rn_sel_nxt[2] ) );
  ANDN U10269 ( .A(n7419), .B(n7169), .Z(n7835) );
  NAND U10270 ( .A(n7923), .B(n7924), .Z(n7169) );
  NANDN U10271 ( .B(n7270), .A(\u_a23_core/u_decode/pre_fetch_instruction[18] ), .Z(n7924) );
  AND U10272 ( .A(n7925), .B(n7926), .Z(n7923) );
  NANDN U10273 ( .B(n7269), .A(\u_a23_core/read_data_s2[18] ), .Z(n7926) );
  NAND U10274 ( .A(n7283), .B(
        \u_a23_core/u_decode/saved_current_instruction[18] ), .Z(n7925) );
  IV U10275 ( .A(n7879), .Z(\u_a23_core/rn_sel_nxt[1] ) );
  ANDN U10276 ( .A(n7419), .B(n7168), .Z(n7879) );
  NAND U10277 ( .A(n7927), .B(n7928), .Z(n7168) );
  NANDN U10278 ( .B(n7270), .A(\u_a23_core/u_decode/pre_fetch_instruction[17] ), .Z(n7928) );
  AND U10279 ( .A(n7929), .B(n7930), .Z(n7927) );
  NANDN U10280 ( .B(n7269), .A(\u_a23_core/read_data_s2[17] ), .Z(n7930) );
  NAND U10281 ( .A(n7283), .B(
        \u_a23_core/u_decode/saved_current_instruction[17] ), .Z(n7929) );
  IV U10282 ( .A(n7896), .Z(\u_a23_core/rn_sel_nxt[0] ) );
  ANDN U10283 ( .A(n7419), .B(n7166), .Z(n7896) );
  NAND U10284 ( .A(n7931), .B(n7932), .Z(n7166) );
  NANDN U10285 ( .B(n7270), .A(\u_a23_core/u_decode/pre_fetch_instruction[16] ), .Z(n7932) );
  AND U10286 ( .A(n7933), .B(n7934), .Z(n7931) );
  NANDN U10287 ( .B(n7269), .A(\u_a23_core/read_data_s2[16] ), .Z(n7934) );
  NAND U10288 ( .A(n7283), .B(
        \u_a23_core/u_decode/saved_current_instruction[16] ), .Z(n7933) );
  NAND U10289 ( .A(n7935), .B(n7936), .Z(\u_a23_core/read_data[9] ) );
  AND U10290 ( .A(n7937), .B(n7938), .Z(n7936) );
  NAND U10291 ( .A(n7939), .B(\u_a23_mem/n21557 ), .Z(n7938) );
  AND U10292 ( .A(n7940), .B(n7941), .Z(n7937) );
  NANDN U10293 ( .B(n4962), .A(\u_a23_mem/n19901 ), .Z(n7941) );
  NAND U10294 ( .A(n7942), .B(\u_a23_mem/n21301 ), .Z(n7940) );
  AND U10295 ( .A(n7943), .B(n7944), .Z(n7935) );
  NAND U10296 ( .A(n5929), .B(\u_a23_mem/n21045 ), .Z(n7944) );
  NAND U10297 ( .A(n1007), .B(\u_a23_mem/n20789 ), .Z(n7943) );
  NAND U10298 ( .A(n7945), .B(n7946), .Z(\u_a23_core/read_data[8] ) );
  AND U10299 ( .A(n7947), .B(n7948), .Z(n7946) );
  NAND U10300 ( .A(n7939), .B(\u_a23_mem/n21528 ), .Z(n7948) );
  AND U10301 ( .A(n7949), .B(n7950), .Z(n7947) );
  NANDN U10302 ( .B(n4962), .A(\u_a23_mem/n19776 ), .Z(n7950) );
  NAND U10303 ( .A(n7942), .B(\u_a23_mem/n21272 ), .Z(n7949) );
  AND U10304 ( .A(n7951), .B(n7952), .Z(n7945) );
  NAND U10305 ( .A(n5929), .B(\u_a23_mem/n21016 ), .Z(n7952) );
  NAND U10306 ( .A(n1007), .B(\u_a23_mem/n20760 ), .Z(n7951) );
  NAND U10307 ( .A(n7953), .B(n7954), .Z(\u_a23_core/read_data[7] ) );
  AND U10308 ( .A(n7955), .B(n7956), .Z(n7954) );
  NAND U10309 ( .A(n7939), .B(\u_a23_mem/N1871 ), .Z(n7956) );
  AND U10310 ( .A(n7957), .B(n7958), .Z(n7955) );
  NANDN U10311 ( .B(n4962), .A(\u_a23_mem/N1839 ), .Z(n7958) );
  NAND U10312 ( .A(n7942), .B(\u_a23_mem/N1903 ), .Z(n7957) );
  AND U10313 ( .A(n7959), .B(n7960), .Z(n7953) );
  NAND U10314 ( .A(n5929), .B(\u_a23_mem/N1935 ), .Z(n7960) );
  NAND U10315 ( .A(n1007), .B(\u_a23_mem/N1967 ), .Z(n7959) );
  NAND U10316 ( .A(n7961), .B(n7962), .Z(\u_a23_core/read_data[6] ) );
  AND U10317 ( .A(n7963), .B(n7964), .Z(n7962) );
  NAND U10318 ( .A(n7939), .B(\u_a23_mem/N1872 ), .Z(n7964) );
  AND U10319 ( .A(n7965), .B(n7966), .Z(n7963) );
  NANDN U10320 ( .B(n4962), .A(\u_a23_mem/N1840 ), .Z(n7966) );
  NAND U10321 ( .A(n7942), .B(\u_a23_mem/N1904 ), .Z(n7965) );
  AND U10322 ( .A(n7967), .B(n7968), .Z(n7961) );
  NAND U10323 ( .A(n5929), .B(\u_a23_mem/N1936 ), .Z(n7968) );
  NAND U10324 ( .A(n1007), .B(\u_a23_mem/N1968 ), .Z(n7967) );
  NAND U10325 ( .A(n7969), .B(n7970), .Z(\u_a23_core/read_data[5] ) );
  AND U10326 ( .A(n7971), .B(n7972), .Z(n7970) );
  NAND U10327 ( .A(n7939), .B(\u_a23_mem/N1873 ), .Z(n7972) );
  AND U10328 ( .A(n7973), .B(n7974), .Z(n7971) );
  NANDN U10329 ( .B(n4962), .A(\u_a23_mem/N1841 ), .Z(n7974) );
  NAND U10330 ( .A(n7942), .B(\u_a23_mem/N1905 ), .Z(n7973) );
  AND U10331 ( .A(n7975), .B(n7976), .Z(n7969) );
  NAND U10332 ( .A(n5929), .B(\u_a23_mem/N1937 ), .Z(n7976) );
  NAND U10333 ( .A(n1007), .B(\u_a23_mem/N1969 ), .Z(n7975) );
  NAND U10334 ( .A(n7977), .B(n7978), .Z(\u_a23_core/read_data[4] ) );
  AND U10335 ( .A(n7979), .B(n7980), .Z(n7978) );
  NAND U10336 ( .A(n7939), .B(\u_a23_mem/N1874 ), .Z(n7980) );
  AND U10337 ( .A(n7981), .B(n7982), .Z(n7979) );
  NANDN U10338 ( .B(n4962), .A(\u_a23_mem/N1842 ), .Z(n7982) );
  NAND U10339 ( .A(n7942), .B(\u_a23_mem/N1906 ), .Z(n7981) );
  AND U10340 ( .A(n7983), .B(n7984), .Z(n7977) );
  NAND U10341 ( .A(n5929), .B(\u_a23_mem/N1938 ), .Z(n7984) );
  NAND U10342 ( .A(n1007), .B(\u_a23_mem/N1970 ), .Z(n7983) );
  NAND U10343 ( .A(n7985), .B(n7986), .Z(\u_a23_core/read_data[3] ) );
  AND U10344 ( .A(n7987), .B(n7988), .Z(n7986) );
  NAND U10345 ( .A(n7939), .B(\u_a23_mem/N1875 ), .Z(n7988) );
  AND U10346 ( .A(n7989), .B(n7990), .Z(n7987) );
  NANDN U10347 ( .B(n4962), .A(\u_a23_mem/N1843 ), .Z(n7990) );
  NAND U10348 ( .A(n7942), .B(\u_a23_mem/N1907 ), .Z(n7989) );
  AND U10349 ( .A(n7991), .B(n7992), .Z(n7985) );
  NAND U10350 ( .A(n5929), .B(\u_a23_mem/N1939 ), .Z(n7992) );
  NAND U10351 ( .A(n1007), .B(\u_a23_mem/N1971 ), .Z(n7991) );
  NAND U10352 ( .A(n7993), .B(n7994), .Z(\u_a23_core/read_data[31] ) );
  AND U10353 ( .A(n7995), .B(n7996), .Z(n7994) );
  NAND U10354 ( .A(n7939), .B(\u_a23_mem/n21724 ), .Z(n7996) );
  AND U10355 ( .A(n7997), .B(n7998), .Z(n7995) );
  NANDN U10356 ( .B(n4962), .A(\u_a23_mem/n20620 ), .Z(n7998) );
  NAND U10357 ( .A(n7942), .B(\u_a23_mem/n21468 ), .Z(n7997) );
  AND U10358 ( .A(n7999), .B(n8000), .Z(n7993) );
  NAND U10359 ( .A(n5929), .B(\u_a23_mem/n21212 ), .Z(n8000) );
  NAND U10360 ( .A(n1007), .B(\u_a23_mem/n20956 ), .Z(n7999) );
  NAND U10361 ( .A(n8001), .B(n8002), .Z(\u_a23_core/read_data[30] ) );
  AND U10362 ( .A(n8003), .B(n8004), .Z(n8002) );
  NAND U10363 ( .A(n7939), .B(\u_a23_mem/n21695 ), .Z(n8004) );
  AND U10364 ( .A(n8005), .B(n8006), .Z(n8003) );
  NANDN U10365 ( .B(n4962), .A(\u_a23_mem/n20495 ), .Z(n8006) );
  NAND U10366 ( .A(n7942), .B(\u_a23_mem/n21439 ), .Z(n8005) );
  AND U10367 ( .A(n8007), .B(n8008), .Z(n8001) );
  NAND U10368 ( .A(n5929), .B(\u_a23_mem/n21183 ), .Z(n8008) );
  NAND U10369 ( .A(n1007), .B(\u_a23_mem/n20927 ), .Z(n8007) );
  NAND U10370 ( .A(n8009), .B(n8010), .Z(\u_a23_core/read_data[2] ) );
  AND U10371 ( .A(n8011), .B(n8012), .Z(n8010) );
  NAND U10372 ( .A(n7939), .B(\u_a23_mem/N1876 ), .Z(n8012) );
  AND U10373 ( .A(n8013), .B(n8014), .Z(n8011) );
  NANDN U10374 ( .B(n4962), .A(\u_a23_mem/N1844 ), .Z(n8014) );
  NAND U10375 ( .A(n7942), .B(\u_a23_mem/N1908 ), .Z(n8013) );
  AND U10376 ( .A(n8015), .B(n8016), .Z(n8009) );
  NAND U10377 ( .A(n5929), .B(\u_a23_mem/N1940 ), .Z(n8016) );
  NAND U10378 ( .A(n1007), .B(\u_a23_mem/N1972 ), .Z(n8015) );
  NAND U10379 ( .A(n8017), .B(n8018), .Z(\u_a23_core/read_data[29] ) );
  AND U10380 ( .A(n8019), .B(n8020), .Z(n8018) );
  NAND U10381 ( .A(n7939), .B(\u_a23_mem/n21666 ), .Z(n8020) );
  AND U10382 ( .A(n8021), .B(n8022), .Z(n8019) );
  NANDN U10383 ( .B(n4962), .A(\u_a23_mem/n20370 ), .Z(n8022) );
  NAND U10384 ( .A(n7942), .B(\u_a23_mem/n21410 ), .Z(n8021) );
  AND U10385 ( .A(n8023), .B(n8024), .Z(n8017) );
  NAND U10386 ( .A(n5929), .B(\u_a23_mem/n21154 ), .Z(n8024) );
  NAND U10387 ( .A(n1007), .B(\u_a23_mem/n20898 ), .Z(n8023) );
  NAND U10388 ( .A(n8025), .B(n8026), .Z(\u_a23_core/read_data[28] ) );
  AND U10389 ( .A(n8027), .B(n8028), .Z(n8026) );
  NAND U10390 ( .A(n7939), .B(\u_a23_mem/n21637 ), .Z(n8028) );
  AND U10391 ( .A(n8029), .B(n8030), .Z(n8027) );
  NANDN U10392 ( .B(n4962), .A(\u_a23_mem/n20245 ), .Z(n8030) );
  NAND U10393 ( .A(n7942), .B(\u_a23_mem/n21381 ), .Z(n8029) );
  AND U10394 ( .A(n8031), .B(n8032), .Z(n8025) );
  NAND U10395 ( .A(n5929), .B(\u_a23_mem/n21125 ), .Z(n8032) );
  NAND U10396 ( .A(n1007), .B(\u_a23_mem/n20869 ), .Z(n8031) );
  NAND U10397 ( .A(n8033), .B(n8034), .Z(\u_a23_core/read_data[27] ) );
  AND U10398 ( .A(n8035), .B(n8036), .Z(n8034) );
  NAND U10399 ( .A(n7939), .B(\u_a23_mem/n21608 ), .Z(n8036) );
  AND U10400 ( .A(n8037), .B(n8038), .Z(n8035) );
  NANDN U10401 ( .B(n4962), .A(\u_a23_mem/n20120 ), .Z(n8038) );
  NAND U10402 ( .A(n7942), .B(\u_a23_mem/n21352 ), .Z(n8037) );
  AND U10403 ( .A(n8039), .B(n8040), .Z(n8033) );
  NAND U10404 ( .A(n5929), .B(\u_a23_mem/n21096 ), .Z(n8040) );
  NAND U10405 ( .A(n1007), .B(\u_a23_mem/n20840 ), .Z(n8039) );
  NAND U10406 ( .A(n8041), .B(n8042), .Z(\u_a23_core/read_data[26] ) );
  AND U10407 ( .A(n8043), .B(n8044), .Z(n8042) );
  NAND U10408 ( .A(n7939), .B(\u_a23_mem/n21579 ), .Z(n8044) );
  AND U10409 ( .A(n8045), .B(n8046), .Z(n8043) );
  NANDN U10410 ( .B(n4962), .A(\u_a23_mem/n19995 ), .Z(n8046) );
  NAND U10411 ( .A(n7942), .B(\u_a23_mem/n21323 ), .Z(n8045) );
  AND U10412 ( .A(n8047), .B(n8048), .Z(n8041) );
  NAND U10413 ( .A(n5929), .B(\u_a23_mem/n21067 ), .Z(n8048) );
  NAND U10414 ( .A(n1007), .B(\u_a23_mem/n20811 ), .Z(n8047) );
  NAND U10415 ( .A(n8049), .B(n8050), .Z(\u_a23_core/read_data[25] ) );
  AND U10416 ( .A(n8051), .B(n8052), .Z(n8050) );
  NAND U10417 ( .A(n7939), .B(\u_a23_mem/n21550 ), .Z(n8052) );
  AND U10418 ( .A(n8053), .B(n8054), .Z(n8051) );
  NANDN U10419 ( .B(n4962), .A(\u_a23_mem/n19870 ), .Z(n8054) );
  NAND U10420 ( .A(n7942), .B(\u_a23_mem/n21294 ), .Z(n8053) );
  AND U10421 ( .A(n8055), .B(n8056), .Z(n8049) );
  NAND U10422 ( .A(n5929), .B(\u_a23_mem/n21038 ), .Z(n8056) );
  NAND U10423 ( .A(n1007), .B(\u_a23_mem/n20782 ), .Z(n8055) );
  NAND U10424 ( .A(n8057), .B(n8058), .Z(\u_a23_core/read_data[24] ) );
  AND U10425 ( .A(n8059), .B(n8060), .Z(n8058) );
  NAND U10426 ( .A(n7939), .B(\u_a23_mem/n21521 ), .Z(n8060) );
  AND U10427 ( .A(n8061), .B(n8062), .Z(n8059) );
  NANDN U10428 ( .B(n4962), .A(\u_a23_mem/n19745 ), .Z(n8062) );
  NAND U10429 ( .A(n7942), .B(\u_a23_mem/n21265 ), .Z(n8061) );
  AND U10430 ( .A(n8063), .B(n8064), .Z(n8057) );
  NAND U10431 ( .A(n5929), .B(\u_a23_mem/n21009 ), .Z(n8064) );
  NAND U10432 ( .A(n1007), .B(\u_a23_mem/n20753 ), .Z(n8063) );
  NAND U10433 ( .A(n8065), .B(n8066), .Z(\u_a23_core/read_data[23] ) );
  AND U10434 ( .A(n8067), .B(n8068), .Z(n8066) );
  NAND U10435 ( .A(n7939), .B(\u_a23_mem/n21716 ), .Z(n8068) );
  AND U10436 ( .A(n8069), .B(n8070), .Z(n8067) );
  NANDN U10437 ( .B(n4962), .A(\u_a23_mem/n20588 ), .Z(n8070) );
  NAND U10438 ( .A(n7942), .B(\u_a23_mem/n21460 ), .Z(n8069) );
  AND U10439 ( .A(n8071), .B(n8072), .Z(n8065) );
  NAND U10440 ( .A(n5929), .B(\u_a23_mem/n21204 ), .Z(n8072) );
  NAND U10441 ( .A(n1007), .B(\u_a23_mem/n20948 ), .Z(n8071) );
  NAND U10442 ( .A(n8073), .B(n8074), .Z(\u_a23_core/read_data[22] ) );
  AND U10443 ( .A(n8075), .B(n8076), .Z(n8074) );
  NAND U10444 ( .A(n7939), .B(\u_a23_mem/n21687 ), .Z(n8076) );
  AND U10445 ( .A(n8077), .B(n8078), .Z(n8075) );
  NANDN U10446 ( .B(n4962), .A(\u_a23_mem/n20463 ), .Z(n8078) );
  NAND U10447 ( .A(n7942), .B(\u_a23_mem/n21431 ), .Z(n8077) );
  AND U10448 ( .A(n8079), .B(n8080), .Z(n8073) );
  NAND U10449 ( .A(n5929), .B(\u_a23_mem/n21175 ), .Z(n8080) );
  NAND U10450 ( .A(n1007), .B(\u_a23_mem/n20919 ), .Z(n8079) );
  NAND U10451 ( .A(n8081), .B(n8082), .Z(\u_a23_core/read_data[21] ) );
  AND U10452 ( .A(n8083), .B(n8084), .Z(n8082) );
  NAND U10453 ( .A(n7939), .B(\u_a23_mem/n21658 ), .Z(n8084) );
  AND U10454 ( .A(n8085), .B(n8086), .Z(n8083) );
  NANDN U10455 ( .B(n4962), .A(\u_a23_mem/n20338 ), .Z(n8086) );
  NAND U10456 ( .A(n7942), .B(\u_a23_mem/n21402 ), .Z(n8085) );
  AND U10457 ( .A(n8087), .B(n8088), .Z(n8081) );
  NAND U10458 ( .A(n5929), .B(\u_a23_mem/n21146 ), .Z(n8088) );
  NAND U10459 ( .A(n1007), .B(\u_a23_mem/n20890 ), .Z(n8087) );
  NAND U10460 ( .A(n8089), .B(n8090), .Z(\u_a23_core/read_data[20] ) );
  AND U10461 ( .A(n8091), .B(n8092), .Z(n8090) );
  NAND U10462 ( .A(n7939), .B(\u_a23_mem/n21629 ), .Z(n8092) );
  AND U10463 ( .A(n8093), .B(n8094), .Z(n8091) );
  NANDN U10464 ( .B(n4962), .A(\u_a23_mem/n20213 ), .Z(n8094) );
  NAND U10465 ( .A(n7942), .B(\u_a23_mem/n21373 ), .Z(n8093) );
  AND U10466 ( .A(n8095), .B(n8096), .Z(n8089) );
  NAND U10467 ( .A(n5929), .B(\u_a23_mem/n21117 ), .Z(n8096) );
  NAND U10468 ( .A(n1007), .B(\u_a23_mem/n20861 ), .Z(n8095) );
  NAND U10469 ( .A(n8097), .B(n8098), .Z(\u_a23_core/read_data[1] ) );
  AND U10470 ( .A(n8099), .B(n8100), .Z(n8098) );
  NAND U10471 ( .A(n7939), .B(\u_a23_mem/N1877 ), .Z(n8100) );
  AND U10472 ( .A(n8101), .B(n8102), .Z(n8099) );
  NANDN U10473 ( .B(n4962), .A(\u_a23_mem/N1845 ), .Z(n8102) );
  NAND U10474 ( .A(n7942), .B(\u_a23_mem/N1909 ), .Z(n8101) );
  AND U10475 ( .A(n8103), .B(n8104), .Z(n8097) );
  NAND U10476 ( .A(n5929), .B(\u_a23_mem/N1941 ), .Z(n8104) );
  NAND U10477 ( .A(n1007), .B(\u_a23_mem/N1973 ), .Z(n8103) );
  NAND U10478 ( .A(n8105), .B(n8106), .Z(\u_a23_core/read_data[19] ) );
  AND U10479 ( .A(n8107), .B(n8108), .Z(n8106) );
  NAND U10480 ( .A(n7939), .B(\u_a23_mem/n21600 ), .Z(n8108) );
  AND U10481 ( .A(n8109), .B(n8110), .Z(n8107) );
  NANDN U10482 ( .B(n4962), .A(\u_a23_mem/n20088 ), .Z(n8110) );
  NAND U10483 ( .A(n7942), .B(\u_a23_mem/n21344 ), .Z(n8109) );
  AND U10484 ( .A(n8111), .B(n8112), .Z(n8105) );
  NAND U10485 ( .A(n5929), .B(\u_a23_mem/n21088 ), .Z(n8112) );
  NAND U10486 ( .A(n1007), .B(\u_a23_mem/n20832 ), .Z(n8111) );
  NAND U10487 ( .A(n8113), .B(n8114), .Z(\u_a23_core/read_data[18] ) );
  AND U10488 ( .A(n8115), .B(n8116), .Z(n8114) );
  NAND U10489 ( .A(n7939), .B(\u_a23_mem/n21571 ), .Z(n8116) );
  AND U10490 ( .A(n8117), .B(n8118), .Z(n8115) );
  NANDN U10491 ( .B(n4962), .A(\u_a23_mem/n19963 ), .Z(n8118) );
  NAND U10492 ( .A(n7942), .B(\u_a23_mem/n21315 ), .Z(n8117) );
  AND U10493 ( .A(n8119), .B(n8120), .Z(n8113) );
  NAND U10494 ( .A(n5929), .B(\u_a23_mem/n21059 ), .Z(n8120) );
  NAND U10495 ( .A(n1007), .B(\u_a23_mem/n20803 ), .Z(n8119) );
  NAND U10496 ( .A(n8121), .B(n8122), .Z(\u_a23_core/read_data[17] ) );
  AND U10497 ( .A(n8123), .B(n8124), .Z(n8122) );
  NAND U10498 ( .A(n7939), .B(\u_a23_mem/n21542 ), .Z(n8124) );
  AND U10499 ( .A(n8125), .B(n8126), .Z(n8123) );
  NANDN U10500 ( .B(n4962), .A(\u_a23_mem/n19838 ), .Z(n8126) );
  NAND U10501 ( .A(n7942), .B(\u_a23_mem/n21286 ), .Z(n8125) );
  AND U10502 ( .A(n8127), .B(n8128), .Z(n8121) );
  NAND U10503 ( .A(n5929), .B(\u_a23_mem/n21030 ), .Z(n8128) );
  NAND U10504 ( .A(n1007), .B(\u_a23_mem/n20774 ), .Z(n8127) );
  NAND U10505 ( .A(n8129), .B(n8130), .Z(\u_a23_core/read_data[16] ) );
  AND U10506 ( .A(n8131), .B(n8132), .Z(n8130) );
  NAND U10507 ( .A(n7939), .B(\u_a23_mem/n21513 ), .Z(n8132) );
  AND U10508 ( .A(n8133), .B(n8134), .Z(n8131) );
  NANDN U10509 ( .B(n4962), .A(\u_a23_mem/n19713 ), .Z(n8134) );
  NAND U10510 ( .A(n7942), .B(\u_a23_mem/n21257 ), .Z(n8133) );
  AND U10511 ( .A(n8135), .B(n8136), .Z(n8129) );
  NAND U10512 ( .A(n5929), .B(\u_a23_mem/n21001 ), .Z(n8136) );
  NAND U10513 ( .A(n1007), .B(\u_a23_mem/n20745 ), .Z(n8135) );
  NAND U10514 ( .A(n8137), .B(n8138), .Z(\u_a23_core/read_data[15] ) );
  AND U10515 ( .A(n8139), .B(n8140), .Z(n8138) );
  NAND U10516 ( .A(n7939), .B(\u_a23_mem/n21731 ), .Z(n8140) );
  AND U10517 ( .A(n8141), .B(n8142), .Z(n8139) );
  NANDN U10518 ( .B(n4962), .A(\u_a23_mem/n20651 ), .Z(n8142) );
  NAND U10519 ( .A(n7942), .B(\u_a23_mem/n21475 ), .Z(n8141) );
  AND U10520 ( .A(n8143), .B(n8144), .Z(n8137) );
  NAND U10521 ( .A(n5929), .B(\u_a23_mem/n21219 ), .Z(n8144) );
  NAND U10522 ( .A(n1007), .B(\u_a23_mem/n20963 ), .Z(n8143) );
  NAND U10523 ( .A(n8145), .B(n8146), .Z(\u_a23_core/read_data[14] ) );
  AND U10524 ( .A(n8147), .B(n8148), .Z(n8146) );
  NAND U10525 ( .A(n7939), .B(\u_a23_mem/n21702 ), .Z(n8148) );
  AND U10526 ( .A(n8149), .B(n8150), .Z(n8147) );
  NANDN U10527 ( .B(n4962), .A(\u_a23_mem/n20526 ), .Z(n8150) );
  NAND U10528 ( .A(n7942), .B(\u_a23_mem/n21446 ), .Z(n8149) );
  AND U10529 ( .A(n8151), .B(n8152), .Z(n8145) );
  NAND U10530 ( .A(n5929), .B(\u_a23_mem/n21190 ), .Z(n8152) );
  NAND U10531 ( .A(n1007), .B(\u_a23_mem/n20934 ), .Z(n8151) );
  NAND U10532 ( .A(n8153), .B(n8154), .Z(\u_a23_core/read_data[13] ) );
  AND U10533 ( .A(n8155), .B(n8156), .Z(n8154) );
  NAND U10534 ( .A(n7939), .B(\u_a23_mem/n21673 ), .Z(n8156) );
  AND U10535 ( .A(n8157), .B(n8158), .Z(n8155) );
  NANDN U10536 ( .B(n4962), .A(\u_a23_mem/n20401 ), .Z(n8158) );
  NAND U10537 ( .A(n7942), .B(\u_a23_mem/n21417 ), .Z(n8157) );
  AND U10538 ( .A(n8159), .B(n8160), .Z(n8153) );
  NAND U10539 ( .A(n5929), .B(\u_a23_mem/n21161 ), .Z(n8160) );
  NAND U10540 ( .A(n1007), .B(\u_a23_mem/n20905 ), .Z(n8159) );
  NAND U10541 ( .A(n8161), .B(n8162), .Z(\u_a23_core/read_data[12] ) );
  AND U10542 ( .A(n8163), .B(n8164), .Z(n8162) );
  NAND U10543 ( .A(n7939), .B(\u_a23_mem/n21644 ), .Z(n8164) );
  AND U10544 ( .A(n8165), .B(n8166), .Z(n8163) );
  NANDN U10545 ( .B(n4962), .A(\u_a23_mem/n20276 ), .Z(n8166) );
  NAND U10546 ( .A(n7942), .B(\u_a23_mem/n21388 ), .Z(n8165) );
  AND U10547 ( .A(n8167), .B(n8168), .Z(n8161) );
  NAND U10548 ( .A(n5929), .B(\u_a23_mem/n21132 ), .Z(n8168) );
  NAND U10549 ( .A(n1007), .B(\u_a23_mem/n20876 ), .Z(n8167) );
  NAND U10550 ( .A(n8169), .B(n8170), .Z(\u_a23_core/read_data[11] ) );
  AND U10551 ( .A(n8171), .B(n8172), .Z(n8170) );
  NAND U10552 ( .A(n7939), .B(\u_a23_mem/n21615 ), .Z(n8172) );
  AND U10553 ( .A(n8173), .B(n8174), .Z(n8171) );
  NANDN U10554 ( .B(n4962), .A(\u_a23_mem/n20151 ), .Z(n8174) );
  NAND U10555 ( .A(n7942), .B(\u_a23_mem/n21359 ), .Z(n8173) );
  AND U10556 ( .A(n8175), .B(n8176), .Z(n8169) );
  NAND U10557 ( .A(n5929), .B(\u_a23_mem/n21103 ), .Z(n8176) );
  NAND U10558 ( .A(n1007), .B(\u_a23_mem/n20847 ), .Z(n8175) );
  NAND U10559 ( .A(n8177), .B(n8178), .Z(\u_a23_core/read_data[10] ) );
  AND U10560 ( .A(n8179), .B(n8180), .Z(n8178) );
  NAND U10561 ( .A(n7939), .B(\u_a23_mem/n21586 ), .Z(n8180) );
  AND U10562 ( .A(n8181), .B(n8182), .Z(n8179) );
  NANDN U10563 ( .B(n4962), .A(\u_a23_mem/n20026 ), .Z(n8182) );
  NAND U10564 ( .A(n7942), .B(\u_a23_mem/n21330 ), .Z(n8181) );
  AND U10565 ( .A(n8183), .B(n8184), .Z(n8177) );
  NAND U10566 ( .A(n5929), .B(\u_a23_mem/n21074 ), .Z(n8184) );
  NAND U10567 ( .A(n1007), .B(\u_a23_mem/n20818 ), .Z(n8183) );
  NAND U10568 ( .A(n8185), .B(n8186), .Z(\u_a23_core/read_data[0] ) );
  AND U10569 ( .A(n8187), .B(n8188), .Z(n8186) );
  NAND U10570 ( .A(n7939), .B(\u_a23_mem/N1878 ), .Z(n8188) );
  AND U10571 ( .A(n8189), .B(n8190), .Z(n7939) );
  AND U10572 ( .A(n8191), .B(n8192), .Z(n8190) );
  AND U10573 ( .A(n8193), .B(m_address[24]), .Z(n8189) );
  AND U10574 ( .A(n8194), .B(n8195), .Z(n8187) );
  NANDN U10575 ( .B(n4962), .A(\u_a23_mem/N1846 ), .Z(n8195) );
  NAND U10576 ( .A(n7942), .B(\u_a23_mem/N1910 ), .Z(n8194) );
  AND U10577 ( .A(n8196), .B(n8197), .Z(n7942) );
  AND U10578 ( .A(n8198), .B(n8192), .Z(n8197) );
  AND U10579 ( .A(m_address[25]), .B(n8193), .Z(n8196) );
  AND U10580 ( .A(n8199), .B(n8200), .Z(n8185) );
  NAND U10581 ( .A(n5929), .B(\u_a23_mem/N1942 ), .Z(n8200) );
  AND U10582 ( .A(n8201), .B(n8202), .Z(n5929) );
  AND U10583 ( .A(n8192), .B(n8193), .Z(n8202) );
  AND U10584 ( .A(m_address[24]), .B(m_address[25]), .Z(n8201) );
  NAND U10585 ( .A(n1007), .B(\u_a23_mem/N1974 ), .Z(n8199) );
  AND U10586 ( .A(n8203), .B(m_address[26]), .Z(n1007) );
  NAND U10587 ( .A(n8204), .B(n8205), .Z(\u_a23_core/rds_sel_nxt[3] ) );
  AND U10588 ( .A(n8206), .B(n7419), .Z(n8205) );
  NANDN U10589 ( .B(n8207), .A(n7258), .Z(n8206) );
  NAND U10590 ( .A(n8208), .B(n8209), .Z(n7258) );
  NANDN U10591 ( .B(n7270), .A(\u_a23_core/u_decode/pre_fetch_instruction[15] ), .Z(n8209) );
  AND U10592 ( .A(n8210), .B(n8211), .Z(n8208) );
  NANDN U10593 ( .B(n7269), .A(\u_a23_core/read_data_s2[15] ), .Z(n8211) );
  NAND U10594 ( .A(n7283), .B(
        \u_a23_core/u_decode/saved_current_instruction[15] ), .Z(n8210) );
  AND U10595 ( .A(n8212), .B(n8213), .Z(n8204) );
  NAND U10596 ( .A(\u_a23_core/u_decode/instruction[11] ), .B(n8214), .Z(n8213) );
  NAND U10597 ( .A(n7181), .B(\u_a23_core/u_decode/N298 ), .Z(n8212) );
  AND U10598 ( .A(n8215), .B(n7213), .Z(\u_a23_core/u_decode/N298 ) );
  ANDN U10599 ( .A(n7678), .B(\u_a23_core/u_decode/instruction[4] ), .Z(n7213)
         );
  AND U10600 ( .A(n7815), .B(n7694), .Z(n8215) );
  NAND U10601 ( .A(n8216), .B(n8217), .Z(\u_a23_core/rds_sel_nxt[2] ) );
  AND U10602 ( .A(n8218), .B(n7419), .Z(n8217) );
  NANDN U10603 ( .B(n8207), .A(n7249), .Z(n8218) );
  AND U10604 ( .A(n8219), .B(n8220), .Z(n8216) );
  NAND U10605 ( .A(\u_a23_core/u_decode/instruction[10] ), .B(n8214), .Z(n8220) );
  NAND U10606 ( .A(n7181), .B(\u_a23_core/u_decode/N319 ), .Z(n8219) );
  AND U10607 ( .A(n8221), .B(n7678), .Z(\u_a23_core/u_decode/N319 ) );
  AND U10608 ( .A(n8222), .B(n7676), .Z(n7678) );
  NAND U10609 ( .A(n8223), .B(n8224), .Z(n8221) );
  AND U10610 ( .A(n7815), .B(n7120), .Z(n8224) );
  ANDN U10611 ( .A(n7694), .B(n7590), .Z(n8223) );
  ANDN U10612 ( .A(n7378), .B(n7574), .Z(n7590) );
  IV U10613 ( .A(n7582), .Z(n7574) );
  NAND U10614 ( .A(n8225), .B(n8226), .Z(\u_a23_core/rds_sel_nxt[1] ) );
  AND U10615 ( .A(n8227), .B(n7419), .Z(n8226) );
  NANDN U10616 ( .B(n8207), .A(n7246), .Z(n8227) );
  AND U10617 ( .A(n8228), .B(n8229), .Z(n8225) );
  NAND U10618 ( .A(\u_a23_core/u_decode/instruction[9] ), .B(n8214), .Z(n8229)
         );
  NAND U10619 ( .A(n7181), .B(\u_a23_core/u_decode/N348 ), .Z(n8228) );
  AND U10620 ( .A(n8230), .B(n7676), .Z(\u_a23_core/u_decode/N348 ) );
  ANDN U10621 ( .A(n7677), .B(\u_a23_core/rm_sel_nxt[1] ), .Z(n7676) );
  IV U10622 ( .A(\u_a23_core/rm_sel_nxt[0] ), .Z(n7677) );
  NAND U10623 ( .A(n8222), .B(n8231), .Z(n8230) );
  NAND U10624 ( .A(n8232), .B(n8233), .Z(n8231) );
  NAND U10625 ( .A(n8234), .B(n8235), .Z(n8233) );
  NAND U10626 ( .A(n7378), .B(n8236), .Z(n8235) );
  NAND U10627 ( .A(n7582), .B(n8237), .Z(n8236) );
  NAND U10628 ( .A(n7704), .B(n7680), .Z(n8237) );
  ANDN U10629 ( .A(n7568), .B(\u_a23_core/u_decode/instruction[11] ), .Z(n7582) );
  ANDN U10630 ( .A(n7580), .B(\u_a23_core/u_decode/instruction[9] ), .Z(n7378)
         );
  ANDN U10631 ( .A(n7815), .B(\u_a23_core/u_decode/instruction[6] ), .Z(n8234)
         );
  AND U10632 ( .A(n7203), .B(n7120), .Z(n8232) );
  AND U10633 ( .A(n8238), .B(n7675), .Z(n8222) );
  NAND U10634 ( .A(n8239), .B(n8240), .Z(\u_a23_core/rds_sel_nxt[0] ) );
  AND U10635 ( .A(n8241), .B(n7419), .Z(n8240) );
  NANDN U10636 ( .B(n7909), .A(n8242), .Z(n7419) );
  AND U10637 ( .A(n7174), .B(n7910), .Z(n8242) );
  NANDN U10638 ( .B(n8207), .A(n7237), .Z(n8241) );
  NANDN U10639 ( .B(n8214), .A(n7214), .Z(n8207) );
  IV U10640 ( .A(n7181), .Z(n7214) );
  AND U10641 ( .A(n8243), .B(n8244), .Z(n8239) );
  NAND U10642 ( .A(\u_a23_core/u_decode/instruction[8] ), .B(n8214), .Z(n8244)
         );
  NAND U10643 ( .A(n8245), .B(n8246), .Z(n8214) );
  NAND U10644 ( .A(n8247), .B(n7134), .Z(n8246) );
  ANDN U10645 ( .A(n8248), .B(n7909), .Z(n7134) );
  AND U10646 ( .A(n7908), .B(n8249), .Z(n8248) );
  AND U10647 ( .A(\u_a23_core/u_decode/instruction[4] ), .B(n7124), .Z(n8247)
         );
  ANDN U10648 ( .A(n8250), .B(n7158), .Z(n8245) );
  AND U10649 ( .A(n7838), .B(n7129), .Z(n7158) );
  NAND U10650 ( .A(n7838), .B(n8251), .Z(n8250) );
  ANDN U10651 ( .A(n7723), .B(n7720), .Z(n8251) );
  IV U10652 ( .A(n7285), .Z(n7838) );
  NANDN U10653 ( .B(n7909), .A(n8252), .Z(n7285) );
  AND U10654 ( .A(n7910), .B(n7908), .Z(n8252) );
  NANDN U10655 ( .B(n7173), .A(n8253), .Z(n7909) );
  NAND U10656 ( .A(n8254), .B(n7764), .Z(n8253) );
  ANDN U10657 ( .A(n7780), .B(n7746), .Z(n7764) );
  IV U10658 ( .A(n7163), .Z(n7780) );
  NAND U10659 ( .A(n8255), .B(n8256), .Z(n7163) );
  NANDN U10660 ( .B(n7270), .A(\u_a23_core/u_decode/pre_fetch_instruction[21] ), .Z(n8256) );
  AND U10661 ( .A(n8257), .B(n8258), .Z(n8255) );
  NANDN U10662 ( .B(n7269), .A(\u_a23_core/read_data_s2[21] ), .Z(n8258) );
  NAND U10663 ( .A(n7283), .B(
        \u_a23_core/u_decode/saved_current_instruction[21] ), .Z(n8257) );
  AND U10664 ( .A(n8259), .B(n7105), .Z(n8254) );
  IV U10665 ( .A(n7135), .Z(n7105) );
  NAND U10666 ( .A(n8260), .B(n8261), .Z(n7135) );
  NANDN U10667 ( .B(n7270), .A(\u_a23_core/u_decode/pre_fetch_instruction[20] ), .Z(n8261) );
  AND U10668 ( .A(n8262), .B(n8263), .Z(n8260) );
  NANDN U10669 ( .B(n7269), .A(\u_a23_core/read_data_s2[20] ), .Z(n8263) );
  NAND U10670 ( .A(n7283), .B(
        \u_a23_core/u_decode/saved_current_instruction[20] ), .Z(n8262) );
  NAND U10671 ( .A(n7181), .B(\u_a23_core/u_decode/N384 ), .Z(n8243) );
  ANDN U10672 ( .A(n8264), .B(\u_a23_core/rm_sel_nxt[0] ), .Z(
        \u_a23_core/u_decode/N384 ) );
  NAND U10673 ( .A(n8265), .B(n8266), .Z(\u_a23_core/rm_sel_nxt[0] ) );
  NANDN U10674 ( .B(n7270), .A(\u_a23_core/u_decode/pre_fetch_instruction[0] ), 
        .Z(n8266) );
  AND U10675 ( .A(n8267), .B(n8268), .Z(n8265) );
  NANDN U10676 ( .B(n7269), .A(\u_a23_core/read_data_s2[0] ), .Z(n8268) );
  NAND U10677 ( .A(n7283), .B(
        \u_a23_core/u_decode/saved_current_instruction[0] ), .Z(n8267) );
  NANDN U10678 ( .B(\u_a23_core/rm_sel_nxt[1] ), .A(n8269), .Z(n8264) );
  NAND U10679 ( .A(n7675), .B(n8270), .Z(n8269) );
  NAND U10680 ( .A(n8238), .B(n8271), .Z(n8270) );
  NAND U10681 ( .A(n7120), .B(n8272), .Z(n8271) );
  NAND U10682 ( .A(n7203), .B(n8273), .Z(n8272) );
  NANDN U10683 ( .B(\u_a23_core/u_decode/instruction[6] ), .A(n8274), .Z(n8273) );
  NAND U10684 ( .A(n8275), .B(n8276), .Z(n8274) );
  NAND U10685 ( .A(n8277), .B(n8278), .Z(n8276) );
  NAND U10686 ( .A(n7819), .B(n8279), .Z(n8278) );
  NAND U10687 ( .A(n7680), .B(n8280), .Z(n8279) );
  NAND U10688 ( .A(n7249), .B(n7704), .Z(n8280) );
  IV U10689 ( .A(n7246), .Z(n7704) );
  NAND U10690 ( .A(n8281), .B(n8282), .Z(n7246) );
  NANDN U10691 ( .B(n7270), .A(\u_a23_core/u_decode/pre_fetch_instruction[13] ), .Z(n8282) );
  AND U10692 ( .A(n8283), .B(n8284), .Z(n8281) );
  NANDN U10693 ( .B(n7269), .A(\u_a23_core/read_data_s2[13] ), .Z(n8284) );
  NAND U10694 ( .A(n7283), .B(
        \u_a23_core/u_decode/saved_current_instruction[13] ), .Z(n8283) );
  NAND U10695 ( .A(n8285), .B(n8286), .Z(n7249) );
  NANDN U10696 ( .B(n7270), .A(\u_a23_core/u_decode/pre_fetch_instruction[14] ), .Z(n8286) );
  AND U10697 ( .A(n8287), .B(n8288), .Z(n8285) );
  NANDN U10698 ( .B(n7269), .A(\u_a23_core/read_data_s2[14] ), .Z(n8288) );
  NAND U10699 ( .A(n7283), .B(
        \u_a23_core/u_decode/saved_current_instruction[14] ), .Z(n8287) );
  IV U10700 ( .A(n7237), .Z(n7680) );
  NAND U10701 ( .A(n8289), .B(n8290), .Z(n7237) );
  NANDN U10702 ( .B(n7270), .A(\u_a23_core/u_decode/pre_fetch_instruction[12] ), .Z(n8290) );
  AND U10703 ( .A(n8291), .B(n8292), .Z(n8289) );
  NANDN U10704 ( .B(n7269), .A(\u_a23_core/read_data_s2[12] ), .Z(n8292) );
  NAND U10705 ( .A(n7283), .B(
        \u_a23_core/u_decode/saved_current_instruction[12] ), .Z(n8291) );
  IV U10706 ( .A(\u_a23_core/u_decode/instruction[11] ), .Z(n7819) );
  NAND U10707 ( .A(n8293), .B(n8294), .Z(\u_a23_core/u_decode/instruction[11] ) );
  NANDN U10708 ( .B(n7270), .A(\u_a23_core/u_decode/pre_fetch_instruction[11] ), .Z(n8294) );
  AND U10709 ( .A(n8295), .B(n8296), .Z(n8293) );
  NANDN U10710 ( .B(n7269), .A(\u_a23_core/read_data_s2[11] ), .Z(n8296) );
  NAND U10711 ( .A(n7283), .B(
        \u_a23_core/u_decode/saved_current_instruction[11] ), .Z(n8295) );
  AND U10712 ( .A(n7580), .B(n7568), .Z(n8277) );
  IV U10713 ( .A(\u_a23_core/u_decode/instruction[10] ), .Z(n7568) );
  NAND U10714 ( .A(n8297), .B(n8298), .Z(\u_a23_core/u_decode/instruction[10] ) );
  NANDN U10715 ( .B(n7270), .A(\u_a23_core/u_decode/pre_fetch_instruction[10] ), .Z(n8298) );
  AND U10716 ( .A(n8299), .B(n8300), .Z(n8297) );
  NANDN U10717 ( .B(n7269), .A(\u_a23_core/read_data_s2[10] ), .Z(n8300) );
  NAND U10718 ( .A(n7283), .B(
        \u_a23_core/u_decode/saved_current_instruction[10] ), .Z(n8299) );
  IV U10719 ( .A(\u_a23_core/u_decode/instruction[8] ), .Z(n7580) );
  AND U10720 ( .A(n7815), .B(n7376), .Z(n8275) );
  IV U10721 ( .A(n7468), .Z(n7376) );
  ANDN U10722 ( .A(\u_a23_core/u_decode/instruction[9] ), .B(
        \u_a23_core/u_decode/instruction[8] ), .Z(n7468) );
  NAND U10723 ( .A(n8301), .B(n8302), .Z(\u_a23_core/u_decode/instruction[8] )
         );
  NANDN U10724 ( .B(n7270), .A(\u_a23_core/u_decode/pre_fetch_instruction[8] ), 
        .Z(n8302) );
  AND U10725 ( .A(n8303), .B(n8304), .Z(n8301) );
  NANDN U10726 ( .B(n7269), .A(\u_a23_core/read_data_s2[8] ), .Z(n8304) );
  NAND U10727 ( .A(n7283), .B(
        \u_a23_core/u_decode/saved_current_instruction[8] ), .Z(n8303) );
  NAND U10728 ( .A(n8305), .B(n8306), .Z(\u_a23_core/u_decode/instruction[9] )
         );
  NANDN U10729 ( .B(n7270), .A(\u_a23_core/u_decode/pre_fetch_instruction[9] ), 
        .Z(n8306) );
  AND U10730 ( .A(n8307), .B(n8308), .Z(n8305) );
  NANDN U10731 ( .B(n7269), .A(\u_a23_core/read_data_s2[9] ), .Z(n8308) );
  NAND U10732 ( .A(n7283), .B(
        \u_a23_core/u_decode/saved_current_instruction[9] ), .Z(n8307) );
  IV U10733 ( .A(\u_a23_core/u_decode/instruction[7] ), .Z(n7815) );
  IV U10734 ( .A(\u_a23_core/u_decode/instruction[4] ), .Z(n7120) );
  IV U10735 ( .A(\u_a23_core/rm_sel_nxt[3] ), .Z(n8238) );
  NAND U10736 ( .A(n8309), .B(n8310), .Z(\u_a23_core/rm_sel_nxt[3] ) );
  NANDN U10737 ( .B(n7270), .A(\u_a23_core/u_decode/pre_fetch_instruction[3] ), 
        .Z(n8310) );
  AND U10738 ( .A(n8311), .B(n8312), .Z(n8309) );
  NANDN U10739 ( .B(n7269), .A(\u_a23_core/read_data_s2[3] ), .Z(n8312) );
  NAND U10740 ( .A(n7283), .B(
        \u_a23_core/u_decode/saved_current_instruction[3] ), .Z(n8311) );
  IV U10741 ( .A(\u_a23_core/rm_sel_nxt[2] ), .Z(n7675) );
  NAND U10742 ( .A(n8313), .B(n8314), .Z(\u_a23_core/rm_sel_nxt[2] ) );
  NANDN U10743 ( .B(n7270), .A(\u_a23_core/u_decode/pre_fetch_instruction[2] ), 
        .Z(n8314) );
  AND U10744 ( .A(n8315), .B(n8316), .Z(n8313) );
  NANDN U10745 ( .B(n7269), .A(\u_a23_core/read_data_s2[2] ), .Z(n8316) );
  NAND U10746 ( .A(n7283), .B(
        \u_a23_core/u_decode/saved_current_instruction[2] ), .Z(n8315) );
  NAND U10747 ( .A(n8317), .B(n8318), .Z(\u_a23_core/rm_sel_nxt[1] ) );
  NANDN U10748 ( .B(n7270), .A(\u_a23_core/u_decode/pre_fetch_instruction[1] ), 
        .Z(n8318) );
  AND U10749 ( .A(n8319), .B(n8320), .Z(n8317) );
  NANDN U10750 ( .B(n7269), .A(\u_a23_core/read_data_s2[1] ), .Z(n8320) );
  NAND U10751 ( .A(n7283), .B(
        \u_a23_core/u_decode/saved_current_instruction[1] ), .Z(n8319) );
  ANDN U10752 ( .A(n8249), .B(n7908), .Z(n7181) );
  IV U10753 ( .A(n7910), .Z(n8249) );
  OR U10754 ( .A(n7173), .B(n8321), .Z(n7910) );
  MUX U10755 ( .IN0(n7172), .IN1(n8322), .SEL(n7908), .F(n8321) );
  IV U10756 ( .A(n7174), .Z(n7908) );
  NAND U10757 ( .A(n8323), .B(n8324), .Z(n7174) );
  NANDN U10758 ( .B(n7270), .A(\u_a23_core/u_decode/pre_fetch_instruction[27] ), .Z(n8324) );
  AND U10759 ( .A(n8325), .B(n8326), .Z(n8323) );
  NANDN U10760 ( .B(n7269), .A(\u_a23_core/read_data_s2[27] ), .Z(n8326) );
  NAND U10761 ( .A(n7283), .B(
        \u_a23_core/u_decode/saved_current_instruction[27] ), .Z(n8325) );
  AND U10762 ( .A(n8259), .B(n8327), .Z(n8322) );
  AND U10763 ( .A(n7746), .B(n7761), .Z(n8327) );
  IV U10764 ( .A(n7114), .Z(n7761) );
  NAND U10765 ( .A(n8328), .B(n8329), .Z(n7114) );
  NANDN U10766 ( .B(n7270), .A(\u_a23_core/u_decode/pre_fetch_instruction[22] ), .Z(n8329) );
  AND U10767 ( .A(n8330), .B(n8331), .Z(n8328) );
  NANDN U10768 ( .B(n7269), .A(\u_a23_core/read_data_s2[22] ), .Z(n8331) );
  NAND U10769 ( .A(n7283), .B(
        \u_a23_core/u_decode/saved_current_instruction[22] ), .Z(n8330) );
  IV U10770 ( .A(n7142), .Z(n7746) );
  NAND U10771 ( .A(n8332), .B(n8333), .Z(n7142) );
  NANDN U10772 ( .B(n7270), .A(\u_a23_core/u_decode/pre_fetch_instruction[24] ), .Z(n8333) );
  AND U10773 ( .A(n8334), .B(n8335), .Z(n8332) );
  NANDN U10774 ( .B(n7269), .A(\u_a23_core/read_data_s2[24] ), .Z(n8335) );
  NAND U10775 ( .A(n7283), .B(
        \u_a23_core/u_decode/saved_current_instruction[24] ), .Z(n8334) );
  AND U10776 ( .A(n8336), .B(n8337), .Z(n8259) );
  AND U10777 ( .A(n8338), .B(n7753), .Z(n8337) );
  IV U10778 ( .A(n7171), .Z(n7753) );
  NAND U10779 ( .A(n8339), .B(n8340), .Z(n7171) );
  NANDN U10780 ( .B(n7270), .A(\u_a23_core/u_decode/pre_fetch_instruction[23] ), .Z(n8340) );
  AND U10781 ( .A(n8341), .B(n8342), .Z(n8339) );
  NANDN U10782 ( .B(n7269), .A(\u_a23_core/read_data_s2[23] ), .Z(n8342) );
  NAND U10783 ( .A(n7283), .B(
        \u_a23_core/u_decode/saved_current_instruction[23] ), .Z(n8341) );
  AND U10784 ( .A(\u_a23_core/u_decode/instruction[7] ), .B(
        \u_a23_core/u_decode/instruction[4] ), .Z(n8338) );
  NAND U10785 ( .A(n8343), .B(n8344), .Z(\u_a23_core/u_decode/instruction[4] )
         );
  NANDN U10786 ( .B(n7270), .A(\u_a23_core/u_decode/pre_fetch_instruction[4] ), 
        .Z(n8344) );
  AND U10787 ( .A(n8345), .B(n8346), .Z(n8343) );
  NANDN U10788 ( .B(n7269), .A(\u_a23_core/read_data_s2[4] ), .Z(n8346) );
  NAND U10789 ( .A(n7283), .B(
        \u_a23_core/u_decode/saved_current_instruction[4] ), .Z(n8345) );
  NAND U10790 ( .A(n8347), .B(n8348), .Z(\u_a23_core/u_decode/instruction[7] )
         );
  NANDN U10791 ( .B(n7270), .A(\u_a23_core/u_decode/pre_fetch_instruction[7] ), 
        .Z(n8348) );
  AND U10792 ( .A(n8349), .B(n8350), .Z(n8347) );
  NANDN U10793 ( .B(n7269), .A(\u_a23_core/read_data_s2[7] ), .Z(n8350) );
  NAND U10794 ( .A(n7283), .B(
        \u_a23_core/u_decode/saved_current_instruction[7] ), .Z(n8349) );
  AND U10795 ( .A(n7124), .B(n7694), .Z(n8336) );
  ANDN U10796 ( .A(n7203), .B(\u_a23_core/u_decode/instruction[6] ), .Z(n7694)
         );
  NAND U10797 ( .A(n8351), .B(n8352), .Z(\u_a23_core/u_decode/instruction[6] )
         );
  NANDN U10798 ( .B(n7270), .A(\u_a23_core/u_decode/pre_fetch_instruction[6] ), 
        .Z(n8352) );
  AND U10799 ( .A(n8353), .B(n8354), .Z(n8351) );
  NANDN U10800 ( .B(n7269), .A(\u_a23_core/read_data_s2[6] ), .Z(n8354) );
  NAND U10801 ( .A(n7283), .B(
        \u_a23_core/u_decode/saved_current_instruction[6] ), .Z(n8353) );
  IV U10802 ( .A(\u_a23_core/u_decode/instruction[5] ), .Z(n7203) );
  NAND U10803 ( .A(n8355), .B(n8356), .Z(\u_a23_core/u_decode/instruction[5] )
         );
  NANDN U10804 ( .B(n7270), .A(\u_a23_core/u_decode/pre_fetch_instruction[5] ), 
        .Z(n8356) );
  AND U10805 ( .A(n8357), .B(n8358), .Z(n8355) );
  NANDN U10806 ( .B(n7269), .A(\u_a23_core/read_data_s2[5] ), .Z(n8358) );
  NAND U10807 ( .A(n7283), .B(
        \u_a23_core/u_decode/saved_current_instruction[5] ), .Z(n8357) );
  IV U10808 ( .A(n7172), .Z(n7124) );
  NAND U10809 ( .A(n8359), .B(n8360), .Z(n7172) );
  NANDN U10810 ( .B(n7270), .A(\u_a23_core/u_decode/pre_fetch_instruction[25] ), .Z(n8360) );
  AND U10811 ( .A(n8361), .B(n8362), .Z(n8359) );
  NANDN U10812 ( .B(n7269), .A(\u_a23_core/read_data_s2[25] ), .Z(n8362) );
  NAND U10813 ( .A(n7283), .B(
        \u_a23_core/u_decode/saved_current_instruction[25] ), .Z(n8361) );
  NAND U10814 ( .A(n8363), .B(n8364), .Z(n7173) );
  NANDN U10815 ( .B(n7270), .A(\u_a23_core/u_decode/pre_fetch_instruction[26] ), .Z(n8364) );
  AND U10816 ( .A(n8365), .B(n8366), .Z(n8363) );
  NANDN U10817 ( .B(n7269), .A(\u_a23_core/read_data_s2[26] ), .Z(n8366) );
  NAND U10818 ( .A(n8367), .B(n7270), .Z(n7269) );
  NAND U10819 ( .A(n7129), .B(\u_a23_core/u_decode/control_state[0] ), .Z(
        n7270) );
  ANDN U10820 ( .A(n7806), .B(n7808), .Z(n7129) );
  NAND U10821 ( .A(\u_a23_core/u_decode/control_state[2] ), .B(n8368), .Z(
        n7808) );
  AND U10822 ( .A(n7723), .B(n7663), .Z(n8368) );
  NAND U10823 ( .A(n7283), .B(
        \u_a23_core/u_decode/saved_current_instruction[26] ), .Z(n8365) );
  IV U10824 ( .A(n8367), .Z(n7283) );
  AND U10825 ( .A(n8369), .B(n8370), .Z(n8367) );
  MUX U10826 ( .IN0(n8371), .IN1(n8372), .SEL(
        \u_a23_core/u_decode/control_state[3] ), .F(n8370) );
  NAND U10827 ( .A(n7806), .B(n8373), .Z(n8372) );
  XOR U10828 ( .A(n7912), .B(n7723), .Z(n8373) );
  IV U10829 ( .A(\u_a23_core/u_decode/control_state[1] ), .Z(n7723) );
  AND U10830 ( .A(n7810), .B(n8374), .Z(n8371) );
  NANDN U10831 ( .B(n8375), .A(\u_a23_core/u_decode/control_state[4] ), .Z(
        n8374) );
  MUX U10832 ( .IN0(\u_a23_core/u_decode/control_state[2] ), .IN1(
        \u_a23_core/u_decode/control_state[1] ), .SEL(n7722), .F(n8375) );
  NANDN U10833 ( .B(n7810), .A(n7722), .Z(n8369) );
  IV U10834 ( .A(\u_a23_core/u_decode/control_state[0] ), .Z(n7722) );
  NAND U10835 ( .A(\u_a23_core/u_decode/control_state[1] ), .B(n8376), .Z(
        n7810) );
  AND U10836 ( .A(n7806), .B(\u_a23_core/u_decode/control_state[2] ), .Z(n8376) );
  IV U10837 ( .A(\u_a23_core/u_decode/control_state[4] ), .Z(n7806) );
  AND U10838 ( .A(n8377), .B(n8378), .Z(terminate) );
  AND U10839 ( .A(n8379), .B(n8380), .Z(n8378) );
  AND U10840 ( .A(n8381), .B(n8382), .Z(n8380) );
  AND U10841 ( .A(n8383), .B(n8384), .Z(n8382) );
  ANDN U10842 ( .A(n8385), .B(\u_a23_core/execute_address_nxt[7] ), .Z(n8384)
         );
  NAND U10843 ( .A(n8386), .B(n8387), .Z(\u_a23_core/execute_address_nxt[7] )
         );
  AND U10844 ( .A(n8388), .B(n8389), .Z(n8387) );
  AND U10845 ( .A(n8390), .B(n8391), .Z(n8389) );
  NANDN U10846 ( .B(n8392), .A(\u_a23_core/u_execute/pc_minus4[7] ), .Z(n8391)
         );
  NAND U10847 ( .A(n8393), .B(\u_a23_core/u_execute/alu_out_pc_filtered[7] ), 
        .Z(n8390) );
  IV U10848 ( .A(n7010), .Z(\u_a23_core/u_execute/alu_out_pc_filtered[7] ) );
  AND U10849 ( .A(n8394), .B(n8395), .Z(n7010) );
  MUX U10850 ( .IN0(n8396), .IN1(n8397), .SEL(
        \u_a23_core/u_execute/u_alu/b_not[7] ), .F(n8395) );
  ANDN U10851 ( .A(n8398), .B(n8399), .Z(n8397) );
  MUX U10852 ( .IN0(n8400), .IN1(\u_a23_core/alu_function[3] ), .SEL(
        \u_a23_core/u_execute/u_alu/a[7] ), .F(n8399) );
  NAND U10853 ( .A(\u_a23_core/u_execute/u_alu/a[7] ), .B(n8400), .Z(n8396) );
  IV U10854 ( .A(n8401), .Z(\u_a23_core/u_execute/u_alu/a[7] ) );
  MUX U10855 ( .IN0(n8402), .IN1(n8403), .SEL(\u_a23_core/alu_function[8] ), 
        .F(n8401) );
  IV U10856 ( .A(\u_a23_core/u_execute/rn[7] ), .Z(n8402) );
  NAND U10857 ( .A(n6765), .B(\u_a23_core/u_execute/u_alu/fadder_out[7] ), .Z(
        n8394) );
  AND U10858 ( .A(n8404), .B(n8405), .Z(n8388) );
  NANDN U10859 ( .B(n8406), .A(\u_a23_core/u_execute/rn_plus4[7] ), .Z(n8405)
         );
  NANDN U10860 ( .B(n8407), .A(\u_a23_core/u_execute/alu_plus4[7] ), .Z(n8404)
         );
  AND U10861 ( .A(n8408), .B(n8409), .Z(n8386) );
  AND U10862 ( .A(n8410), .B(n8411), .Z(n8409) );
  NAND U10863 ( .A(n8412), .B(\u_a23_core/u_execute/address_plus4[7] ), .Z(
        n8411) );
  NAND U10864 ( .A(\u_a23_core/u_execute/rn[7] ), .B(n8413), .Z(n8410) );
  AND U10865 ( .A(n8414), .B(n8415), .Z(n8408) );
  NAND U10866 ( .A(\u_a23_core/u_execute/pc[7] ), .B(n8416), .Z(n8415) );
  NAND U10867 ( .A(n8417), .B(\u_a23_core/u_execute/pc_plus4[7] ), .Z(n8414)
         );
  NOR U10868 ( .A(\u_a23_core/execute_address_nxt[8] ), .B(
        \u_a23_core/execute_address_nxt[9] ), .Z(n8385) );
  NAND U10869 ( .A(n8418), .B(n8419), .Z(\u_a23_core/execute_address_nxt[9] )
         );
  AND U10870 ( .A(n8420), .B(n8421), .Z(n8419) );
  AND U10871 ( .A(n8422), .B(n8423), .Z(n8421) );
  NANDN U10872 ( .B(n8392), .A(\u_a23_core/u_execute/pc_minus4[9] ), .Z(n8423)
         );
  NAND U10873 ( .A(n8393), .B(\u_a23_core/u_execute/alu_out_pc_filtered[9] ), 
        .Z(n8422) );
  IV U10874 ( .A(n7008), .Z(\u_a23_core/u_execute/alu_out_pc_filtered[9] ) );
  AND U10875 ( .A(n8424), .B(n8425), .Z(n7008) );
  MUX U10876 ( .IN0(n8426), .IN1(n8427), .SEL(
        \u_a23_core/u_execute/u_alu/b_not[9] ), .F(n8425) );
  NAND U10877 ( .A(n8428), .B(n8429), .Z(\u_a23_core/u_execute/u_alu/b_not[9] ) );
  MUX U10878 ( .IN0(n8430), .IN1(n8431), .SEL(n8432), .F(n8429) );
  MUX U10879 ( .IN0(n8433), .IN1(n8434), .SEL(\u_a23_core/u_execute/rn[9] ), 
        .F(n8428) );
  ANDN U10880 ( .A(n8435), .B(n8436), .Z(n8427) );
  MUX U10881 ( .IN0(n8400), .IN1(\u_a23_core/alu_function[3] ), .SEL(
        \u_a23_core/u_execute/u_alu/a[9] ), .F(n8436) );
  NAND U10882 ( .A(\u_a23_core/u_execute/u_alu/a[9] ), .B(n8400), .Z(n8426) );
  IV U10883 ( .A(n8437), .Z(\u_a23_core/u_execute/u_alu/a[9] ) );
  MUX U10884 ( .IN0(n8438), .IN1(n8432), .SEL(\u_a23_core/alu_function[8] ), 
        .F(n8437) );
  AND U10885 ( .A(n8439), .B(n8440), .Z(n8432) );
  AND U10886 ( .A(n8441), .B(n8442), .Z(n8440) );
  NAND U10887 ( .A(n8443), .B(n8444), .Z(n8442) );
  NAND U10888 ( .A(n8445), .B(n8446), .Z(n8444) );
  NAND U10889 ( .A(n6882), .B(n8447), .Z(n8445) );
  NAND U10890 ( .A(n8448), .B(n8449), .Z(n8447) );
  AND U10891 ( .A(n8450), .B(n8451), .Z(n8441) );
  NANDN U10892 ( .B(n8446), .A(n8452), .Z(n8451) );
  AND U10893 ( .A(n8453), .B(n8454), .Z(n8446) );
  AND U10894 ( .A(n8455), .B(n8456), .Z(n8454) );
  AND U10895 ( .A(n8457), .B(n8458), .Z(n8456) );
  AND U10896 ( .A(n8459), .B(n8460), .Z(n8458) );
  NAND U10897 ( .A(n8461), .B(n6839), .Z(n8460) );
  AND U10898 ( .A(n8462), .B(n8463), .Z(n8459) );
  NAND U10899 ( .A(n8464), .B(n6833), .Z(n8463) );
  NAND U10900 ( .A(n8465), .B(n6835), .Z(n8462) );
  AND U10901 ( .A(n8466), .B(n8467), .Z(n8457) );
  AND U10902 ( .A(n8468), .B(n8469), .Z(n8466) );
  NAND U10903 ( .A(n6850), .B(n8470), .Z(n8469) );
  AND U10904 ( .A(n8471), .B(n8472), .Z(n8455) );
  AND U10905 ( .A(n8473), .B(n8474), .Z(n8472) );
  NAND U10906 ( .A(n6856), .B(n6799), .Z(n8474) );
  AND U10907 ( .A(n8475), .B(n8476), .Z(n8473) );
  NAND U10908 ( .A(n6840), .B(n6807), .Z(n8476) );
  NAND U10909 ( .A(n6852), .B(n6809), .Z(n8475) );
  AND U10910 ( .A(n8477), .B(n8478), .Z(n8471) );
  NAND U10911 ( .A(n6858), .B(n6803), .Z(n8478) );
  NAND U10912 ( .A(n6864), .B(n6823), .Z(n8477) );
  AND U10913 ( .A(n8479), .B(n8480), .Z(n8453) );
  AND U10914 ( .A(n8481), .B(n8482), .Z(n8480) );
  AND U10915 ( .A(n8483), .B(n8484), .Z(n8482) );
  AND U10916 ( .A(n8485), .B(n8486), .Z(n8483) );
  NAND U10917 ( .A(n6827), .B(n8487), .Z(n8486) );
  AND U10918 ( .A(n8488), .B(n8489), .Z(n8481) );
  AND U10919 ( .A(n8490), .B(n8491), .Z(n8488) );
  AND U10920 ( .A(n8492), .B(n8493), .Z(n8479) );
  AND U10921 ( .A(n8494), .B(n8495), .Z(n8493) );
  AND U10922 ( .A(n8496), .B(n8497), .Z(n8494) );
  AND U10923 ( .A(n8498), .B(n8499), .Z(n8492) );
  NAND U10924 ( .A(n6893), .B(n6947), .Z(n8498) );
  NAND U10925 ( .A(n8500), .B(n6888), .Z(n8450) );
  NAND U10926 ( .A(n8501), .B(n8502), .Z(n8500) );
  AND U10927 ( .A(n8503), .B(n8504), .Z(n8502) );
  AND U10928 ( .A(n8505), .B(n8506), .Z(n8504) );
  AND U10929 ( .A(n8507), .B(n8508), .Z(n8506) );
  AND U10930 ( .A(n8509), .B(n8510), .Z(n8508) );
  NANDN U10931 ( .B(n8511), .A(n6919), .Z(n8510) );
  NAND U10932 ( .A(n6947), .B(n8512), .Z(n8509) );
  AND U10933 ( .A(n8513), .B(n8514), .Z(n8507) );
  NANDN U10934 ( .B(n8515), .A(n6920), .Z(n8514) );
  NANDN U10935 ( .B(n8516), .A(n6946), .Z(n8513) );
  AND U10936 ( .A(n8517), .B(n8518), .Z(n8505) );
  AND U10937 ( .A(n8519), .B(n8520), .Z(n8518) );
  NANDN U10938 ( .B(n8521), .A(n6925), .Z(n8520) );
  NANDN U10939 ( .B(n8522), .A(n6943), .Z(n8519) );
  AND U10940 ( .A(n8523), .B(n8524), .Z(n8517) );
  NANDN U10941 ( .B(n8525), .A(n6926), .Z(n8524) );
  NANDN U10942 ( .B(n8526), .A(n6942), .Z(n8523) );
  AND U10943 ( .A(n8527), .B(n8528), .Z(n8503) );
  AND U10944 ( .A(n8529), .B(n8530), .Z(n8528) );
  AND U10945 ( .A(n8531), .B(n8532), .Z(n8530) );
  NANDN U10946 ( .B(n8533), .A(n6898), .Z(n8532) );
  NANDN U10947 ( .B(n8534), .A(n6937), .Z(n8531) );
  AND U10948 ( .A(n8535), .B(n8536), .Z(n8529) );
  NANDN U10949 ( .B(n8537), .A(n6882), .Z(n8536) );
  NANDN U10950 ( .B(n8538), .A(n6809), .Z(n8535) );
  AND U10951 ( .A(n8539), .B(n8540), .Z(n8527) );
  AND U10952 ( .A(n8541), .B(n8542), .Z(n8540) );
  NANDN U10953 ( .B(n8543), .A(n6807), .Z(n8542) );
  NANDN U10954 ( .B(n8544), .A(n6799), .Z(n8541) );
  AND U10955 ( .A(n8545), .B(n8546), .Z(n8539) );
  NANDN U10956 ( .B(n8547), .A(n6803), .Z(n8546) );
  NANDN U10957 ( .B(n8548), .A(n6823), .Z(n8545) );
  AND U10958 ( .A(n8549), .B(n8550), .Z(n8501) );
  AND U10959 ( .A(n8551), .B(n8552), .Z(n8550) );
  AND U10960 ( .A(n8553), .B(n8554), .Z(n8552) );
  AND U10961 ( .A(n8555), .B(n8556), .Z(n8554) );
  NANDN U10962 ( .B(n8557), .A(n6827), .Z(n8556) );
  NANDN U10963 ( .B(n8558), .A(n6833), .Z(n8555) );
  AND U10964 ( .A(n8559), .B(n8560), .Z(n8553) );
  NANDN U10965 ( .B(n8561), .A(n6835), .Z(n8560) );
  NANDN U10966 ( .B(n8562), .A(n6839), .Z(n8559) );
  AND U10967 ( .A(n8563), .B(n8564), .Z(n8551) );
  AND U10968 ( .A(n8565), .B(n8566), .Z(n8564) );
  NANDN U10969 ( .B(n8567), .A(n6850), .Z(n8566) );
  NANDN U10970 ( .B(n8568), .A(n6853), .Z(n8565) );
  AND U10971 ( .A(n8569), .B(n8570), .Z(n8563) );
  NANDN U10972 ( .B(n8571), .A(n6841), .Z(n8570) );
  NANDN U10973 ( .B(n8572), .A(n6857), .Z(n8569) );
  AND U10974 ( .A(n8573), .B(n8574), .Z(n8549) );
  AND U10975 ( .A(n8575), .B(n8576), .Z(n8574) );
  AND U10976 ( .A(n8577), .B(n8578), .Z(n8576) );
  NANDN U10977 ( .B(n8579), .A(n6859), .Z(n8578) );
  NANDN U10978 ( .B(n8580), .A(n6865), .Z(n8577) );
  AND U10979 ( .A(n8581), .B(n8582), .Z(n8575) );
  NANDN U10980 ( .B(n8583), .A(n6967), .Z(n8582) );
  NANDN U10981 ( .B(n8584), .A(n6966), .Z(n8581) );
  AND U10982 ( .A(n8585), .B(n8586), .Z(n8573) );
  AND U10983 ( .A(n8587), .B(n8588), .Z(n8586) );
  NANDN U10984 ( .B(n8589), .A(n6961), .Z(n8588) );
  NANDN U10985 ( .B(n8590), .A(n6956), .Z(n8587) );
  AND U10986 ( .A(n8591), .B(n8592), .Z(n8585) );
  NANDN U10987 ( .B(n8593), .A(n6960), .Z(n8592) );
  NAND U10988 ( .A(n6957), .B(n6897), .Z(n8591) );
  AND U10989 ( .A(n8594), .B(n8595), .Z(n8439) );
  NAND U10990 ( .A(n8596), .B(n6902), .Z(n8595) );
  NAND U10991 ( .A(n8597), .B(n8598), .Z(n8596) );
  AND U10992 ( .A(n8599), .B(n8600), .Z(n8598) );
  AND U10993 ( .A(n8601), .B(n8602), .Z(n8600) );
  NAND U10994 ( .A(n8603), .B(n6898), .Z(n8602) );
  AND U10995 ( .A(n8604), .B(n8605), .Z(n8601) );
  NAND U10996 ( .A(n6947), .B(n6916), .Z(n8605) );
  NAND U10997 ( .A(n8606), .B(n6925), .Z(n8604) );
  AND U10998 ( .A(n8607), .B(n8608), .Z(n8599) );
  NAND U10999 ( .A(n8609), .B(n6926), .Z(n8608) );
  NAND U11000 ( .A(n8610), .B(n6920), .Z(n8607) );
  AND U11001 ( .A(n8611), .B(n8612), .Z(n8597) );
  AND U11002 ( .A(n8613), .B(n8614), .Z(n8612) );
  AND U11003 ( .A(n8615), .B(n6875), .Z(n8613) );
  NAND U11004 ( .A(n8616), .B(n6919), .Z(n6875) );
  AND U11005 ( .A(n8617), .B(n8618), .Z(n8611) );
  NAND U11006 ( .A(n6985), .B(n6851), .Z(n8594) );
  IV U11007 ( .A(\u_a23_core/u_execute/rn[9] ), .Z(n8438) );
  AND U11008 ( .A(n8619), .B(n8620), .Z(n8424) );
  NAND U11009 ( .A(n6765), .B(\u_a23_core/u_execute/u_alu/fadder_out[9] ), .Z(
        n8619) );
  AND U11010 ( .A(n8621), .B(n8622), .Z(n8420) );
  NANDN U11011 ( .B(n8406), .A(\u_a23_core/u_execute/rn_plus4[9] ), .Z(n8622)
         );
  NANDN U11012 ( .B(n8407), .A(\u_a23_core/u_execute/alu_plus4[9] ), .Z(n8621)
         );
  AND U11013 ( .A(n8623), .B(n8624), .Z(n8418) );
  AND U11014 ( .A(n8625), .B(n8626), .Z(n8624) );
  NAND U11015 ( .A(n8412), .B(\u_a23_core/u_execute/address_plus4[9] ), .Z(
        n8626) );
  NAND U11016 ( .A(\u_a23_core/u_execute/rn[9] ), .B(n8413), .Z(n8625) );
  NAND U11017 ( .A(n8627), .B(n8628), .Z(\u_a23_core/u_execute/rn[9] ) );
  AND U11018 ( .A(n8629), .B(n8630), .Z(n8628) );
  AND U11019 ( .A(n8631), .B(n8632), .Z(n8630) );
  AND U11020 ( .A(n8633), .B(n8634), .Z(n8632) );
  NANDN U11021 ( .B(n8635), .A(\u_a23_core/u_execute/pc[9] ), .Z(n8634) );
  NANDN U11022 ( .B(n8636), .A(\u_a23_core/u_execute/u_register_bank/r14[9] ), 
        .Z(n8633) );
  AND U11023 ( .A(n8637), .B(n8638), .Z(n8631) );
  NANDN U11024 ( .B(n8639), .A(\u_a23_core/u_execute/u_register_bank/r13[9] ), 
        .Z(n8638) );
  NANDN U11025 ( .B(n8640), .A(\u_a23_core/u_execute/u_register_bank/r12[9] ), 
        .Z(n8637) );
  AND U11026 ( .A(n8641), .B(n8642), .Z(n8629) );
  AND U11027 ( .A(n8643), .B(n8644), .Z(n8642) );
  NANDN U11028 ( .B(n8645), .A(\u_a23_core/u_execute/u_register_bank/r11[9] ), 
        .Z(n8644) );
  NANDN U11029 ( .B(n8646), .A(\u_a23_core/u_execute/u_register_bank/r10[9] ), 
        .Z(n8643) );
  AND U11030 ( .A(n8647), .B(n8648), .Z(n8641) );
  NANDN U11031 ( .B(n8649), .A(\u_a23_core/u_execute/u_register_bank/r9[9] ), 
        .Z(n8648) );
  NANDN U11032 ( .B(n8650), .A(\u_a23_core/u_execute/u_register_bank/r8[9] ), 
        .Z(n8647) );
  AND U11033 ( .A(n8651), .B(n8652), .Z(n8627) );
  AND U11034 ( .A(n8653), .B(n8654), .Z(n8652) );
  AND U11035 ( .A(n8655), .B(n8656), .Z(n8654) );
  NANDN U11036 ( .B(n8657), .A(\u_a23_core/u_execute/u_register_bank/r7[9] ), 
        .Z(n8656) );
  NANDN U11037 ( .B(n8658), .A(\u_a23_core/u_execute/u_register_bank/r6[9] ), 
        .Z(n8655) );
  AND U11038 ( .A(n8659), .B(n8660), .Z(n8653) );
  NANDN U11039 ( .B(n8661), .A(\u_a23_core/u_execute/u_register_bank/r5[9] ), 
        .Z(n8660) );
  NANDN U11040 ( .B(n8662), .A(\u_a23_core/u_execute/u_register_bank/r4[9] ), 
        .Z(n8659) );
  AND U11041 ( .A(n8663), .B(n8664), .Z(n8651) );
  AND U11042 ( .A(n8665), .B(n8666), .Z(n8664) );
  NANDN U11043 ( .B(n8667), .A(\u_a23_core/u_execute/u_register_bank/r3[9] ), 
        .Z(n8666) );
  NANDN U11044 ( .B(n8668), .A(\u_a23_core/u_execute/u_register_bank/r0[9] ), 
        .Z(n8665) );
  AND U11045 ( .A(n8669), .B(n8670), .Z(n8663) );
  NANDN U11046 ( .B(n8671), .A(\u_a23_core/u_execute/u_register_bank/r2[9] ), 
        .Z(n8670) );
  NANDN U11047 ( .B(n8672), .A(\u_a23_core/u_execute/u_register_bank/r1[9] ), 
        .Z(n8669) );
  AND U11048 ( .A(n8673), .B(n8674), .Z(n8623) );
  NAND U11049 ( .A(\u_a23_core/u_execute/pc[9] ), .B(n8416), .Z(n8674) );
  NAND U11050 ( .A(n8417), .B(\u_a23_core/u_execute/pc_plus4[9] ), .Z(n8673)
         );
  NAND U11051 ( .A(n8675), .B(n8676), .Z(\u_a23_core/execute_address_nxt[8] )
         );
  AND U11052 ( .A(n8677), .B(n8678), .Z(n8676) );
  AND U11053 ( .A(n8679), .B(n8680), .Z(n8678) );
  NANDN U11054 ( .B(n8392), .A(\u_a23_core/u_execute/pc_minus4[8] ), .Z(n8680)
         );
  NAND U11055 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[8] ), .B(n8393), 
        .Z(n8679) );
  IV U11056 ( .A(n7009), .Z(\u_a23_core/u_execute/alu_out_pc_filtered[8] ) );
  AND U11057 ( .A(n8681), .B(n8682), .Z(n7009) );
  MUX U11058 ( .IN0(n8683), .IN1(n8684), .SEL(
        \u_a23_core/u_execute/u_alu/b_not[8] ), .F(n8682) );
  NAND U11059 ( .A(n8685), .B(n8686), .Z(\u_a23_core/u_execute/u_alu/b_not[8] ) );
  MUX U11060 ( .IN0(n8430), .IN1(n8431), .SEL(n8687), .F(n8686) );
  MUX U11061 ( .IN0(n8433), .IN1(n8434), .SEL(\u_a23_core/u_execute/rn[8] ), 
        .F(n8685) );
  ANDN U11062 ( .A(n8435), .B(n8688), .Z(n8684) );
  MUX U11063 ( .IN0(n8400), .IN1(\u_a23_core/alu_function[3] ), .SEL(
        \u_a23_core/u_execute/u_alu/a[8] ), .F(n8688) );
  NAND U11064 ( .A(\u_a23_core/u_execute/u_alu/a[8] ), .B(n8400), .Z(n8683) );
  IV U11065 ( .A(n8689), .Z(\u_a23_core/u_execute/u_alu/a[8] ) );
  MUX U11066 ( .IN0(n8690), .IN1(n8687), .SEL(\u_a23_core/alu_function[8] ), 
        .F(n8689) );
  AND U11067 ( .A(n8691), .B(n8692), .Z(n8687) );
  AND U11068 ( .A(n8693), .B(n8694), .Z(n8692) );
  NAND U11069 ( .A(n6886), .B(n8695), .Z(n8694) );
  NAND U11070 ( .A(n8696), .B(n8448), .Z(n8695) );
  NAND U11071 ( .A(n6786), .B(n8697), .Z(n8693) );
  NAND U11072 ( .A(n8698), .B(n8699), .Z(n8697) );
  AND U11073 ( .A(n8700), .B(n8701), .Z(n8699) );
  AND U11074 ( .A(n8702), .B(n8703), .Z(n8701) );
  AND U11075 ( .A(n8704), .B(n8705), .Z(n8703) );
  NOR U11076 ( .A(n8706), .B(n8707), .Z(n8705) );
  AND U11077 ( .A(n8708), .B(n8709), .Z(n8702) );
  NAND U11078 ( .A(n8465), .B(n6839), .Z(n8709) );
  ANDN U11079 ( .A(n8710), .B(n8711), .Z(n8708) );
  NAND U11080 ( .A(n8464), .B(n6835), .Z(n8710) );
  AND U11081 ( .A(n8712), .B(n8713), .Z(n8700) );
  AND U11082 ( .A(n8714), .B(n8715), .Z(n8713) );
  AND U11083 ( .A(n6933), .B(n8716), .Z(n8714) );
  NAND U11084 ( .A(n6850), .B(n8461), .Z(n8716) );
  NAND U11085 ( .A(n8470), .B(n6853), .Z(n6933) );
  AND U11086 ( .A(n8717), .B(n8718), .Z(n8712) );
  NAND U11087 ( .A(n6840), .B(n6799), .Z(n8718) );
  AND U11088 ( .A(n8719), .B(n8720), .Z(n8717) );
  NAND U11089 ( .A(n6882), .B(n6838), .Z(n8719) );
  AND U11090 ( .A(n8721), .B(n8722), .Z(n8698) );
  AND U11091 ( .A(n8723), .B(n8724), .Z(n8722) );
  AND U11092 ( .A(n8725), .B(n8726), .Z(n8724) );
  NAND U11093 ( .A(n6856), .B(n6803), .Z(n8726) );
  AND U11094 ( .A(n8727), .B(n8728), .Z(n8725) );
  NAND U11095 ( .A(n6809), .B(n6851), .Z(n8728) );
  NAND U11096 ( .A(n6852), .B(n6807), .Z(n8727) );
  AND U11097 ( .A(n8729), .B(n8730), .Z(n8723) );
  NAND U11098 ( .A(n6833), .B(n8487), .Z(n8730) );
  AND U11099 ( .A(n8731), .B(n8732), .Z(n8729) );
  NAND U11100 ( .A(n6858), .B(n6823), .Z(n8732) );
  NAND U11101 ( .A(n6864), .B(n6827), .Z(n8731) );
  AND U11102 ( .A(n8733), .B(n8734), .Z(n8721) );
  AND U11103 ( .A(n8735), .B(n8736), .Z(n8734) );
  AND U11104 ( .A(n8737), .B(n8738), .Z(n8735) );
  AND U11105 ( .A(n8739), .B(n8740), .Z(n8733) );
  NAND U11106 ( .A(n6893), .B(n6946), .Z(n8740) );
  AND U11107 ( .A(n8741), .B(n8742), .Z(n8739) );
  AND U11108 ( .A(n8743), .B(n8744), .Z(n8691) );
  NAND U11109 ( .A(n8745), .B(n6888), .Z(n8744) );
  NAND U11110 ( .A(n8746), .B(n8747), .Z(n8745) );
  AND U11111 ( .A(n8748), .B(n8749), .Z(n8747) );
  AND U11112 ( .A(n8750), .B(n8751), .Z(n8749) );
  AND U11113 ( .A(n8752), .B(n8753), .Z(n8751) );
  AND U11114 ( .A(n8754), .B(n8755), .Z(n8753) );
  NANDN U11115 ( .B(n8534), .A(n6919), .Z(n8755) );
  NAND U11116 ( .A(n6946), .B(n8512), .Z(n8754) );
  AND U11117 ( .A(n8756), .B(n8757), .Z(n8752) );
  NANDN U11118 ( .B(n8511), .A(n6920), .Z(n8757) );
  NANDN U11119 ( .B(n8516), .A(n6943), .Z(n8756) );
  AND U11120 ( .A(n8758), .B(n8759), .Z(n8750) );
  AND U11121 ( .A(n8760), .B(n8761), .Z(n8759) );
  NANDN U11122 ( .B(n8515), .A(n6925), .Z(n8761) );
  NANDN U11123 ( .B(n8522), .A(n6942), .Z(n8760) );
  AND U11124 ( .A(n8762), .B(n8763), .Z(n8758) );
  NANDN U11125 ( .B(n8521), .A(n6926), .Z(n8763) );
  NANDN U11126 ( .B(n8526), .A(n6937), .Z(n8762) );
  AND U11127 ( .A(n8764), .B(n8765), .Z(n8748) );
  AND U11128 ( .A(n8766), .B(n8767), .Z(n8765) );
  AND U11129 ( .A(n8768), .B(n8769), .Z(n8767) );
  NANDN U11130 ( .B(n8525), .A(n6898), .Z(n8769) );
  NANDN U11131 ( .B(n8533), .A(n6882), .Z(n8768) );
  AND U11132 ( .A(n8770), .B(n8771), .Z(n8766) );
  NANDN U11133 ( .B(n8537), .A(n6809), .Z(n8771) );
  NANDN U11134 ( .B(n8538), .A(n6807), .Z(n8770) );
  AND U11135 ( .A(n8772), .B(n8773), .Z(n8764) );
  AND U11136 ( .A(n8774), .B(n8775), .Z(n8773) );
  NANDN U11137 ( .B(n8543), .A(n6799), .Z(n8775) );
  NANDN U11138 ( .B(n8544), .A(n6803), .Z(n8774) );
  AND U11139 ( .A(n8776), .B(n8777), .Z(n8772) );
  NANDN U11140 ( .B(n8547), .A(n6823), .Z(n8777) );
  NANDN U11141 ( .B(n8548), .A(n6827), .Z(n8776) );
  AND U11142 ( .A(n8778), .B(n8779), .Z(n8746) );
  AND U11143 ( .A(n8780), .B(n8781), .Z(n8779) );
  AND U11144 ( .A(n8782), .B(n8783), .Z(n8781) );
  AND U11145 ( .A(n8784), .B(n8785), .Z(n8783) );
  NANDN U11146 ( .B(n8557), .A(n6833), .Z(n8785) );
  NANDN U11147 ( .B(n8558), .A(n6835), .Z(n8784) );
  AND U11148 ( .A(n8786), .B(n8787), .Z(n8782) );
  NANDN U11149 ( .B(n8561), .A(n6839), .Z(n8787) );
  NANDN U11150 ( .B(n8562), .A(n6850), .Z(n8786) );
  AND U11151 ( .A(n8788), .B(n8789), .Z(n8780) );
  AND U11152 ( .A(n8790), .B(n8791), .Z(n8789) );
  NANDN U11153 ( .B(n8567), .A(n6853), .Z(n8791) );
  NANDN U11154 ( .B(n8568), .A(n6841), .Z(n8790) );
  AND U11155 ( .A(n8792), .B(n8793), .Z(n8788) );
  NANDN U11156 ( .B(n8571), .A(n6857), .Z(n8793) );
  NANDN U11157 ( .B(n8572), .A(n6859), .Z(n8792) );
  AND U11158 ( .A(n8794), .B(n8795), .Z(n8778) );
  AND U11159 ( .A(n8796), .B(n8797), .Z(n8795) );
  AND U11160 ( .A(n8798), .B(n8799), .Z(n8797) );
  NANDN U11161 ( .B(n8579), .A(n6865), .Z(n8799) );
  NANDN U11162 ( .B(n8580), .A(n6967), .Z(n8798) );
  AND U11163 ( .A(n8800), .B(n8801), .Z(n8796) );
  NANDN U11164 ( .B(n8583), .A(n6966), .Z(n8801) );
  NANDN U11165 ( .B(n8584), .A(n6961), .Z(n8800) );
  AND U11166 ( .A(n8802), .B(n8803), .Z(n8794) );
  AND U11167 ( .A(n8804), .B(n8805), .Z(n8803) );
  NANDN U11168 ( .B(n8589), .A(n6956), .Z(n8805) );
  NANDN U11169 ( .B(n8590), .A(n6960), .Z(n8804) );
  AND U11170 ( .A(n8806), .B(n8807), .Z(n8802) );
  NANDN U11171 ( .B(n8593), .A(n6957), .Z(n8807) );
  NAND U11172 ( .A(n6947), .B(n6897), .Z(n8806) );
  NAND U11173 ( .A(n8808), .B(n6902), .Z(n8743) );
  NAND U11174 ( .A(n8809), .B(n8810), .Z(n8808) );
  AND U11175 ( .A(n8811), .B(n8812), .Z(n8810) );
  AND U11176 ( .A(n8813), .B(n8814), .Z(n8812) );
  NAND U11177 ( .A(n8609), .B(n6898), .Z(n8814) );
  AND U11178 ( .A(n8815), .B(n8816), .Z(n8813) );
  NAND U11179 ( .A(n6946), .B(n6916), .Z(n8816) );
  NAND U11180 ( .A(n8606), .B(n6926), .Z(n8815) );
  AND U11181 ( .A(n8817), .B(n8818), .Z(n8811) );
  NAND U11182 ( .A(n8610), .B(n6925), .Z(n8818) );
  NAND U11183 ( .A(n8616), .B(n6920), .Z(n8817) );
  AND U11184 ( .A(n8819), .B(n8820), .Z(n8809) );
  AND U11185 ( .A(n8821), .B(n8822), .Z(n8820) );
  AND U11186 ( .A(n8823), .B(n8824), .Z(n8819) );
  IV U11187 ( .A(\u_a23_core/u_execute/rn[8] ), .Z(n8690) );
  AND U11188 ( .A(n8825), .B(n8620), .Z(n8681) );
  NAND U11189 ( .A(n6765), .B(\u_a23_core/u_execute/u_alu/fadder_out[8] ), .Z(
        n8825) );
  AND U11190 ( .A(n8826), .B(n8827), .Z(n8677) );
  NANDN U11191 ( .B(n8406), .A(\u_a23_core/u_execute/rn_plus4[8] ), .Z(n8827)
         );
  NANDN U11192 ( .B(n8407), .A(\u_a23_core/u_execute/alu_plus4[8] ), .Z(n8826)
         );
  AND U11193 ( .A(n8828), .B(n8829), .Z(n8675) );
  AND U11194 ( .A(n8830), .B(n8831), .Z(n8829) );
  NAND U11195 ( .A(n8412), .B(\u_a23_core/u_execute/address_plus4[8] ), .Z(
        n8831) );
  NAND U11196 ( .A(\u_a23_core/u_execute/rn[8] ), .B(n8413), .Z(n8830) );
  NAND U11197 ( .A(n8832), .B(n8833), .Z(\u_a23_core/u_execute/rn[8] ) );
  AND U11198 ( .A(n8834), .B(n8835), .Z(n8833) );
  AND U11199 ( .A(n8836), .B(n8837), .Z(n8835) );
  AND U11200 ( .A(n8838), .B(n8839), .Z(n8837) );
  NANDN U11201 ( .B(n8635), .A(\u_a23_core/u_execute/pc[8] ), .Z(n8839) );
  NANDN U11202 ( .B(n8636), .A(\u_a23_core/u_execute/u_register_bank/r14[8] ), 
        .Z(n8838) );
  AND U11203 ( .A(n8840), .B(n8841), .Z(n8836) );
  NANDN U11204 ( .B(n8639), .A(\u_a23_core/u_execute/u_register_bank/r13[8] ), 
        .Z(n8841) );
  NANDN U11205 ( .B(n8640), .A(\u_a23_core/u_execute/u_register_bank/r12[8] ), 
        .Z(n8840) );
  AND U11206 ( .A(n8842), .B(n8843), .Z(n8834) );
  AND U11207 ( .A(n8844), .B(n8845), .Z(n8843) );
  NANDN U11208 ( .B(n8645), .A(\u_a23_core/u_execute/u_register_bank/r11[8] ), 
        .Z(n8845) );
  NANDN U11209 ( .B(n8646), .A(\u_a23_core/u_execute/u_register_bank/r10[8] ), 
        .Z(n8844) );
  AND U11210 ( .A(n8846), .B(n8847), .Z(n8842) );
  NANDN U11211 ( .B(n8649), .A(\u_a23_core/u_execute/u_register_bank/r9[8] ), 
        .Z(n8847) );
  NANDN U11212 ( .B(n8650), .A(\u_a23_core/u_execute/u_register_bank/r8[8] ), 
        .Z(n8846) );
  AND U11213 ( .A(n8848), .B(n8849), .Z(n8832) );
  AND U11214 ( .A(n8850), .B(n8851), .Z(n8849) );
  AND U11215 ( .A(n8852), .B(n8853), .Z(n8851) );
  NANDN U11216 ( .B(n8657), .A(\u_a23_core/u_execute/u_register_bank/r7[8] ), 
        .Z(n8853) );
  NANDN U11217 ( .B(n8658), .A(\u_a23_core/u_execute/u_register_bank/r6[8] ), 
        .Z(n8852) );
  AND U11218 ( .A(n8854), .B(n8855), .Z(n8850) );
  NANDN U11219 ( .B(n8661), .A(\u_a23_core/u_execute/u_register_bank/r5[8] ), 
        .Z(n8855) );
  NANDN U11220 ( .B(n8662), .A(\u_a23_core/u_execute/u_register_bank/r4[8] ), 
        .Z(n8854) );
  AND U11221 ( .A(n8856), .B(n8857), .Z(n8848) );
  AND U11222 ( .A(n8858), .B(n8859), .Z(n8857) );
  NANDN U11223 ( .B(n8667), .A(\u_a23_core/u_execute/u_register_bank/r3[8] ), 
        .Z(n8859) );
  NANDN U11224 ( .B(n8668), .A(\u_a23_core/u_execute/u_register_bank/r0[8] ), 
        .Z(n8858) );
  AND U11225 ( .A(n8860), .B(n8861), .Z(n8856) );
  NANDN U11226 ( .B(n8671), .A(\u_a23_core/u_execute/u_register_bank/r2[8] ), 
        .Z(n8861) );
  NANDN U11227 ( .B(n8672), .A(\u_a23_core/u_execute/u_register_bank/r1[8] ), 
        .Z(n8860) );
  AND U11228 ( .A(n8862), .B(n8863), .Z(n8828) );
  NAND U11229 ( .A(\u_a23_core/u_execute/pc[8] ), .B(n8416), .Z(n8863) );
  NAND U11230 ( .A(n8417), .B(\u_a23_core/u_execute/pc_plus4[8] ), .Z(n8862)
         );
  NOR U11231 ( .A(\u_a23_core/execute_address_nxt[5] ), .B(
        \u_a23_core/execute_address_nxt[6] ), .Z(n8383) );
  NAND U11232 ( .A(n8864), .B(n8865), .Z(\u_a23_core/execute_address_nxt[6] )
         );
  AND U11233 ( .A(n8866), .B(n8867), .Z(n8865) );
  AND U11234 ( .A(n8868), .B(n8869), .Z(n8867) );
  NANDN U11235 ( .B(n8392), .A(\u_a23_core/u_execute/pc_minus4[6] ), .Z(n8869)
         );
  NAND U11236 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[6] ), .B(n8393), 
        .Z(n8868) );
  IV U11237 ( .A(n7011), .Z(\u_a23_core/u_execute/alu_out_pc_filtered[6] ) );
  AND U11238 ( .A(n8870), .B(n8871), .Z(n7011) );
  MUX U11239 ( .IN0(n8872), .IN1(n8873), .SEL(
        \u_a23_core/u_execute/u_alu/b_not[6] ), .F(n8871) );
  NAND U11240 ( .A(n8874), .B(n8875), .Z(\u_a23_core/u_execute/u_alu/b_not[6] ) );
  MUX U11241 ( .IN0(n8430), .IN1(n8431), .SEL(n8876), .F(n8875) );
  MUX U11242 ( .IN0(n8433), .IN1(n8434), .SEL(\u_a23_core/u_execute/rn[6] ), 
        .F(n8874) );
  ANDN U11243 ( .A(n8398), .B(n8877), .Z(n8873) );
  MUX U11244 ( .IN0(n8400), .IN1(\u_a23_core/alu_function[3] ), .SEL(
        \u_a23_core/u_execute/u_alu/a[6] ), .F(n8877) );
  NAND U11245 ( .A(\u_a23_core/u_execute/u_alu/a[6] ), .B(n8400), .Z(n8872) );
  IV U11246 ( .A(n8878), .Z(\u_a23_core/u_execute/u_alu/a[6] ) );
  MUX U11247 ( .IN0(n8879), .IN1(n8876), .SEL(\u_a23_core/alu_function[8] ), 
        .F(n8878) );
  AND U11248 ( .A(n8880), .B(n8881), .Z(n8876) );
  AND U11249 ( .A(n8882), .B(n8883), .Z(n8881) );
  NAND U11250 ( .A(n8884), .B(n6888), .Z(n8883) );
  NAND U11251 ( .A(n8885), .B(n8886), .Z(n8884) );
  AND U11252 ( .A(n8887), .B(n8888), .Z(n8886) );
  AND U11253 ( .A(n8889), .B(n8890), .Z(n8888) );
  AND U11254 ( .A(n8891), .B(n8892), .Z(n8890) );
  AND U11255 ( .A(n8893), .B(n8894), .Z(n8892) );
  NANDN U11256 ( .B(n8522), .A(n6919), .Z(n8894) );
  NAND U11257 ( .A(n6942), .B(n8512), .Z(n8893) );
  AND U11258 ( .A(n8895), .B(n8896), .Z(n8891) );
  NANDN U11259 ( .B(n8526), .A(n6920), .Z(n8896) );
  NANDN U11260 ( .B(n8516), .A(n6937), .Z(n8895) );
  AND U11261 ( .A(n8897), .B(n8898), .Z(n8889) );
  AND U11262 ( .A(n8899), .B(n8900), .Z(n8898) );
  NANDN U11263 ( .B(n8534), .A(n6925), .Z(n8900) );
  NANDN U11264 ( .B(n8511), .A(n6926), .Z(n8899) );
  AND U11265 ( .A(n8901), .B(n8902), .Z(n8897) );
  NANDN U11266 ( .B(n8515), .A(n6898), .Z(n8902) );
  NANDN U11267 ( .B(n8521), .A(n6882), .Z(n8901) );
  AND U11268 ( .A(n8903), .B(n8904), .Z(n8887) );
  AND U11269 ( .A(n8905), .B(n8906), .Z(n8904) );
  AND U11270 ( .A(n8907), .B(n8908), .Z(n8906) );
  NANDN U11271 ( .B(n8525), .A(n6809), .Z(n8908) );
  NANDN U11272 ( .B(n8533), .A(n6807), .Z(n8907) );
  AND U11273 ( .A(n8909), .B(n8910), .Z(n8905) );
  NANDN U11274 ( .B(n8537), .A(n6799), .Z(n8910) );
  NANDN U11275 ( .B(n8538), .A(n6803), .Z(n8909) );
  AND U11276 ( .A(n8911), .B(n8912), .Z(n8903) );
  AND U11277 ( .A(n8913), .B(n8914), .Z(n8912) );
  NANDN U11278 ( .B(n8543), .A(n6823), .Z(n8914) );
  NANDN U11279 ( .B(n8544), .A(n6827), .Z(n8913) );
  AND U11280 ( .A(n8915), .B(n8916), .Z(n8911) );
  NANDN U11281 ( .B(n8547), .A(n6833), .Z(n8916) );
  NANDN U11282 ( .B(n8548), .A(n6835), .Z(n8915) );
  AND U11283 ( .A(n8917), .B(n8918), .Z(n8885) );
  AND U11284 ( .A(n8919), .B(n8920), .Z(n8918) );
  AND U11285 ( .A(n8921), .B(n8922), .Z(n8920) );
  AND U11286 ( .A(n8923), .B(n8924), .Z(n8922) );
  NANDN U11287 ( .B(n8557), .A(n6839), .Z(n8924) );
  NANDN U11288 ( .B(n8558), .A(n6850), .Z(n8923) );
  AND U11289 ( .A(n8925), .B(n8926), .Z(n8921) );
  NANDN U11290 ( .B(n8561), .A(n6853), .Z(n8926) );
  NANDN U11291 ( .B(n8562), .A(n6841), .Z(n8925) );
  AND U11292 ( .A(n8927), .B(n8928), .Z(n8919) );
  AND U11293 ( .A(n8929), .B(n8930), .Z(n8928) );
  NANDN U11294 ( .B(n8567), .A(n6857), .Z(n8930) );
  NANDN U11295 ( .B(n8568), .A(n6859), .Z(n8929) );
  AND U11296 ( .A(n8931), .B(n8932), .Z(n8927) );
  NANDN U11297 ( .B(n8571), .A(n6865), .Z(n8932) );
  NANDN U11298 ( .B(n8572), .A(n6967), .Z(n8931) );
  AND U11299 ( .A(n8933), .B(n8934), .Z(n8917) );
  AND U11300 ( .A(n8935), .B(n8936), .Z(n8934) );
  AND U11301 ( .A(n8937), .B(n8938), .Z(n8936) );
  NANDN U11302 ( .B(n8579), .A(n6966), .Z(n8938) );
  NANDN U11303 ( .B(n8580), .A(n6961), .Z(n8937) );
  AND U11304 ( .A(n8939), .B(n8940), .Z(n8935) );
  NANDN U11305 ( .B(n8583), .A(n6956), .Z(n8940) );
  NANDN U11306 ( .B(n8584), .A(n6960), .Z(n8939) );
  AND U11307 ( .A(n8941), .B(n8942), .Z(n8933) );
  AND U11308 ( .A(n8943), .B(n8944), .Z(n8942) );
  NANDN U11309 ( .B(n8589), .A(n6957), .Z(n8944) );
  NANDN U11310 ( .B(n8590), .A(n6947), .Z(n8943) );
  AND U11311 ( .A(n8945), .B(n8946), .Z(n8941) );
  NANDN U11312 ( .B(n8593), .A(n6946), .Z(n8946) );
  NAND U11313 ( .A(n6943), .B(n6897), .Z(n8945) );
  AND U11314 ( .A(n8947), .B(n8948), .Z(n8882) );
  NAND U11315 ( .A(n8949), .B(n6902), .Z(n8948) );
  NAND U11316 ( .A(n8950), .B(n8951), .Z(n8949) );
  AND U11317 ( .A(n8952), .B(n8953), .Z(n8951) );
  AND U11318 ( .A(n8954), .B(n8955), .Z(n8953) );
  NAND U11319 ( .A(n6942), .B(n6916), .Z(n8955) );
  NAND U11320 ( .A(n8610), .B(n6898), .Z(n8954) );
  AND U11321 ( .A(n8956), .B(n8957), .Z(n8952) );
  NAND U11322 ( .A(n8616), .B(n6926), .Z(n8957) );
  NAND U11323 ( .A(n8958), .B(n6925), .Z(n8956) );
  AND U11324 ( .A(n8959), .B(n8960), .Z(n8950) );
  AND U11325 ( .A(n8961), .B(n8962), .Z(n8959) );
  NAND U11326 ( .A(n6786), .B(n8963), .Z(n8947) );
  NAND U11327 ( .A(n8964), .B(n8965), .Z(n8963) );
  AND U11328 ( .A(n8966), .B(n8967), .Z(n8965) );
  AND U11329 ( .A(n8968), .B(n8969), .Z(n8967) );
  AND U11330 ( .A(n8970), .B(n8971), .Z(n8969) );
  ANDN U11331 ( .A(n8972), .B(n8973), .Z(n8971) );
  NOR U11332 ( .A(n8974), .B(n8975), .Z(n8970) );
  AND U11333 ( .A(n8976), .B(n6934), .Z(n8968) );
  NAND U11334 ( .A(n8461), .B(n6841), .Z(n6934) );
  AND U11335 ( .A(n8977), .B(n8978), .Z(n8976) );
  NAND U11336 ( .A(n6850), .B(n8464), .Z(n8978) );
  NAND U11337 ( .A(n8465), .B(n6853), .Z(n8977) );
  AND U11338 ( .A(n8979), .B(n8980), .Z(n8966) );
  AND U11339 ( .A(n8981), .B(n8982), .Z(n8980) );
  AND U11340 ( .A(n8983), .B(n8984), .Z(n8981) );
  AND U11341 ( .A(n8985), .B(n8986), .Z(n8979) );
  NAND U11342 ( .A(n6838), .B(n6807), .Z(n8986) );
  AND U11343 ( .A(n8987), .B(n8988), .Z(n8985) );
  NAND U11344 ( .A(n6882), .B(n6832), .Z(n8988) );
  NAND U11345 ( .A(n6834), .B(n6809), .Z(n8987) );
  AND U11346 ( .A(n8989), .B(n8990), .Z(n8964) );
  AND U11347 ( .A(n8991), .B(n8992), .Z(n8990) );
  AND U11348 ( .A(n8993), .B(n8994), .Z(n8992) );
  AND U11349 ( .A(n8995), .B(n8996), .Z(n8994) );
  NAND U11350 ( .A(n6840), .B(n6823), .Z(n8996) );
  NAND U11351 ( .A(n6799), .B(n6851), .Z(n8995) );
  AND U11352 ( .A(n8997), .B(n8998), .Z(n8993) );
  NAND U11353 ( .A(n6852), .B(n6803), .Z(n8998) );
  NAND U11354 ( .A(n6856), .B(n6827), .Z(n8997) );
  AND U11355 ( .A(n8999), .B(n9000), .Z(n8991) );
  NAND U11356 ( .A(n6839), .B(n8487), .Z(n9000) );
  AND U11357 ( .A(n9001), .B(n9002), .Z(n8999) );
  NAND U11358 ( .A(n6858), .B(n6833), .Z(n9002) );
  NAND U11359 ( .A(n6864), .B(n6835), .Z(n9001) );
  AND U11360 ( .A(n9003), .B(n9004), .Z(n8989) );
  AND U11361 ( .A(n9005), .B(n9006), .Z(n9004) );
  AND U11362 ( .A(n9007), .B(n9008), .Z(n9005) );
  AND U11363 ( .A(n9009), .B(n9010), .Z(n9003) );
  NAND U11364 ( .A(n6893), .B(n6942), .Z(n9010) );
  AND U11365 ( .A(n8823), .B(n9011), .Z(n9009) );
  NAND U11366 ( .A(n6984), .B(n6943), .Z(n8823) );
  AND U11367 ( .A(n9012), .B(n9013), .Z(n8880) );
  NAND U11368 ( .A(n6886), .B(n6826), .Z(n9013) );
  IV U11369 ( .A(\u_a23_core/u_execute/rn[6] ), .Z(n8879) );
  NAND U11370 ( .A(n6765), .B(\u_a23_core/u_execute/u_alu/fadder_out[6] ), .Z(
        n8870) );
  AND U11371 ( .A(n9014), .B(n9015), .Z(n8866) );
  NANDN U11372 ( .B(n8406), .A(\u_a23_core/u_execute/rn_plus4[6] ), .Z(n9015)
         );
  NANDN U11373 ( .B(n8407), .A(\u_a23_core/u_execute/alu_plus4[6] ), .Z(n9014)
         );
  AND U11374 ( .A(n9016), .B(n9017), .Z(n8864) );
  AND U11375 ( .A(n9018), .B(n9019), .Z(n9017) );
  NAND U11376 ( .A(n8412), .B(\u_a23_core/u_execute/address_plus4[6] ), .Z(
        n9019) );
  NAND U11377 ( .A(\u_a23_core/u_execute/rn[6] ), .B(n8413), .Z(n9018) );
  NAND U11378 ( .A(n9020), .B(n9021), .Z(\u_a23_core/u_execute/rn[6] ) );
  AND U11379 ( .A(n9022), .B(n9023), .Z(n9021) );
  AND U11380 ( .A(n9024), .B(n9025), .Z(n9023) );
  AND U11381 ( .A(n9026), .B(n9027), .Z(n9025) );
  NANDN U11382 ( .B(n8635), .A(\u_a23_core/u_execute/pc[6] ), .Z(n9027) );
  NANDN U11383 ( .B(n8636), .A(\u_a23_core/u_execute/u_register_bank/r14[6] ), 
        .Z(n9026) );
  AND U11384 ( .A(n9028), .B(n9029), .Z(n9024) );
  NANDN U11385 ( .B(n8639), .A(\u_a23_core/u_execute/u_register_bank/r13[6] ), 
        .Z(n9029) );
  NANDN U11386 ( .B(n8640), .A(\u_a23_core/u_execute/u_register_bank/r12[6] ), 
        .Z(n9028) );
  AND U11387 ( .A(n9030), .B(n9031), .Z(n9022) );
  AND U11388 ( .A(n9032), .B(n9033), .Z(n9031) );
  NANDN U11389 ( .B(n8645), .A(\u_a23_core/u_execute/u_register_bank/r11[6] ), 
        .Z(n9033) );
  NANDN U11390 ( .B(n8646), .A(\u_a23_core/u_execute/u_register_bank/r10[6] ), 
        .Z(n9032) );
  AND U11391 ( .A(n9034), .B(n9035), .Z(n9030) );
  NANDN U11392 ( .B(n8649), .A(\u_a23_core/u_execute/u_register_bank/r9[6] ), 
        .Z(n9035) );
  NANDN U11393 ( .B(n8650), .A(\u_a23_core/u_execute/u_register_bank/r8[6] ), 
        .Z(n9034) );
  AND U11394 ( .A(n9036), .B(n9037), .Z(n9020) );
  AND U11395 ( .A(n9038), .B(n9039), .Z(n9037) );
  AND U11396 ( .A(n9040), .B(n9041), .Z(n9039) );
  NANDN U11397 ( .B(n8657), .A(\u_a23_core/u_execute/u_register_bank/r7[6] ), 
        .Z(n9041) );
  NANDN U11398 ( .B(n8658), .A(\u_a23_core/u_execute/u_register_bank/r6[6] ), 
        .Z(n9040) );
  AND U11399 ( .A(n9042), .B(n9043), .Z(n9038) );
  NANDN U11400 ( .B(n8661), .A(\u_a23_core/u_execute/u_register_bank/r5[6] ), 
        .Z(n9043) );
  NANDN U11401 ( .B(n8662), .A(\u_a23_core/u_execute/u_register_bank/r4[6] ), 
        .Z(n9042) );
  AND U11402 ( .A(n9044), .B(n9045), .Z(n9036) );
  AND U11403 ( .A(n9046), .B(n9047), .Z(n9045) );
  NANDN U11404 ( .B(n8667), .A(\u_a23_core/u_execute/u_register_bank/r3[6] ), 
        .Z(n9047) );
  NANDN U11405 ( .B(n8668), .A(\u_a23_core/u_execute/u_register_bank/r0[6] ), 
        .Z(n9046) );
  AND U11406 ( .A(n9048), .B(n9049), .Z(n9044) );
  NANDN U11407 ( .B(n8671), .A(\u_a23_core/u_execute/u_register_bank/r2[6] ), 
        .Z(n9049) );
  NANDN U11408 ( .B(n8672), .A(\u_a23_core/u_execute/u_register_bank/r1[6] ), 
        .Z(n9048) );
  AND U11409 ( .A(n9050), .B(n9051), .Z(n9016) );
  NAND U11410 ( .A(\u_a23_core/u_execute/pc[6] ), .B(n8416), .Z(n9051) );
  NAND U11411 ( .A(n8417), .B(\u_a23_core/u_execute/pc_plus4[6] ), .Z(n9050)
         );
  NAND U11412 ( .A(n9052), .B(n9053), .Z(\u_a23_core/execute_address_nxt[5] )
         );
  AND U11413 ( .A(n9054), .B(n9055), .Z(n9053) );
  AND U11414 ( .A(n9056), .B(n9057), .Z(n9055) );
  NANDN U11415 ( .B(n8392), .A(\u_a23_core/u_execute/pc_minus4[5] ), .Z(n9057)
         );
  NAND U11416 ( .A(n8393), .B(\u_a23_core/u_execute/alu_out_pc_filtered[5] ), 
        .Z(n9056) );
  IV U11417 ( .A(n7014), .Z(\u_a23_core/u_execute/alu_out_pc_filtered[5] ) );
  AND U11418 ( .A(n9058), .B(n9059), .Z(n7014) );
  MUX U11419 ( .IN0(n9060), .IN1(n9061), .SEL(
        \u_a23_core/u_execute/u_alu/b_not[5] ), .F(n9059) );
  NAND U11420 ( .A(n9062), .B(n9063), .Z(\u_a23_core/u_execute/u_alu/b_not[5] ) );
  MUX U11421 ( .IN0(n8430), .IN1(n8431), .SEL(n9064), .F(n9063) );
  MUX U11422 ( .IN0(n8433), .IN1(n8434), .SEL(\u_a23_core/u_execute/rn[5] ), 
        .F(n9062) );
  ANDN U11423 ( .A(n8398), .B(n9065), .Z(n9061) );
  MUX U11424 ( .IN0(n8400), .IN1(\u_a23_core/alu_function[3] ), .SEL(
        \u_a23_core/u_execute/u_alu/a[5] ), .F(n9065) );
  NAND U11425 ( .A(\u_a23_core/u_execute/u_alu/a[5] ), .B(n8400), .Z(n9060) );
  IV U11426 ( .A(n9066), .Z(\u_a23_core/u_execute/u_alu/a[5] ) );
  MUX U11427 ( .IN0(n9067), .IN1(n9064), .SEL(\u_a23_core/alu_function[8] ), 
        .F(n9066) );
  AND U11428 ( .A(n9068), .B(n9069), .Z(n9064) );
  AND U11429 ( .A(n9070), .B(n9071), .Z(n9069) );
  NAND U11430 ( .A(n9072), .B(n6902), .Z(n9071) );
  NAND U11431 ( .A(n9073), .B(n9074), .Z(n9072) );
  AND U11432 ( .A(n9075), .B(n9076), .Z(n9074) );
  NAND U11433 ( .A(n8958), .B(n6926), .Z(n9076) );
  AND U11434 ( .A(n9077), .B(n9078), .Z(n9075) );
  NAND U11435 ( .A(n6937), .B(n6916), .Z(n9078) );
  NAND U11436 ( .A(n8616), .B(n6898), .Z(n9077) );
  AND U11437 ( .A(n9079), .B(n9080), .Z(n9073) );
  AND U11438 ( .A(n9081), .B(n6879), .Z(n9079) );
  NAND U11439 ( .A(n9082), .B(n6925), .Z(n6879) );
  NAND U11440 ( .A(n6786), .B(n9083), .Z(n9070) );
  NAND U11441 ( .A(n9084), .B(n9085), .Z(n9083) );
  AND U11442 ( .A(n9086), .B(n9087), .Z(n9085) );
  AND U11443 ( .A(n9088), .B(n9089), .Z(n9087) );
  AND U11444 ( .A(n9090), .B(n9091), .Z(n9089) );
  AND U11445 ( .A(n9092), .B(n9093), .Z(n9091) );
  NAND U11446 ( .A(n8464), .B(n6853), .Z(n9093) );
  NAND U11447 ( .A(n8465), .B(n6841), .Z(n9092) );
  AND U11448 ( .A(n9094), .B(n9095), .Z(n9090) );
  AND U11449 ( .A(n9096), .B(n9097), .Z(n9088) );
  NAND U11450 ( .A(n6882), .B(n6826), .Z(n9097) );
  AND U11451 ( .A(n9098), .B(n9099), .Z(n9096) );
  AND U11452 ( .A(n9100), .B(n9101), .Z(n9086) );
  AND U11453 ( .A(n9102), .B(n9103), .Z(n9101) );
  AND U11454 ( .A(n9104), .B(n9105), .Z(n9103) );
  NAND U11455 ( .A(n6832), .B(n6809), .Z(n9105) );
  NAND U11456 ( .A(n6834), .B(n6807), .Z(n9104) );
  AND U11457 ( .A(n9106), .B(n9107), .Z(n9102) );
  NAND U11458 ( .A(n6838), .B(n6799), .Z(n9107) );
  NAND U11459 ( .A(n6840), .B(n6827), .Z(n9106) );
  AND U11460 ( .A(n9108), .B(n9109), .Z(n9100) );
  NAND U11461 ( .A(n6856), .B(n6833), .Z(n9109) );
  AND U11462 ( .A(n9110), .B(n9111), .Z(n9108) );
  NAND U11463 ( .A(n6803), .B(n6851), .Z(n9111) );
  NAND U11464 ( .A(n6852), .B(n6823), .Z(n9110) );
  AND U11465 ( .A(n9112), .B(n9113), .Z(n9084) );
  AND U11466 ( .A(n9114), .B(n9115), .Z(n9113) );
  AND U11467 ( .A(n9116), .B(n9117), .Z(n9115) );
  AND U11468 ( .A(n9118), .B(n9119), .Z(n9117) );
  NAND U11469 ( .A(n6858), .B(n6835), .Z(n9119) );
  NAND U11470 ( .A(n6864), .B(n6839), .Z(n9118) );
  AND U11471 ( .A(n9120), .B(n9121), .Z(n9116) );
  NAND U11472 ( .A(n6850), .B(n8487), .Z(n9121) );
  AND U11473 ( .A(n9122), .B(n9123), .Z(n9114) );
  AND U11474 ( .A(n9124), .B(n9125), .Z(n9122) );
  AND U11475 ( .A(n9126), .B(n9127), .Z(n9112) );
  AND U11476 ( .A(n9128), .B(n9129), .Z(n9127) );
  AND U11477 ( .A(n9130), .B(n9131), .Z(n9128) );
  AND U11478 ( .A(n9132), .B(n9133), .Z(n9126) );
  NAND U11479 ( .A(n6893), .B(n6937), .Z(n9133) );
  AND U11480 ( .A(n9134), .B(n8618), .Z(n9132) );
  NAND U11481 ( .A(n9135), .B(n6943), .Z(n8618) );
  AND U11482 ( .A(n9012), .B(n9136), .Z(n9068) );
  NAND U11483 ( .A(n9137), .B(n6888), .Z(n9136) );
  NAND U11484 ( .A(n9138), .B(n9139), .Z(n9137) );
  AND U11485 ( .A(n9140), .B(n9141), .Z(n9139) );
  AND U11486 ( .A(n9142), .B(n9143), .Z(n9141) );
  AND U11487 ( .A(n9144), .B(n9145), .Z(n9143) );
  AND U11488 ( .A(n9146), .B(n9147), .Z(n9145) );
  NANDN U11489 ( .B(n8516), .A(n6919), .Z(n9147) );
  NAND U11490 ( .A(n6937), .B(n8512), .Z(n9146) );
  AND U11491 ( .A(n9148), .B(n9149), .Z(n9144) );
  NANDN U11492 ( .B(n8522), .A(n6920), .Z(n9149) );
  NANDN U11493 ( .B(n8526), .A(n6925), .Z(n9148) );
  AND U11494 ( .A(n9150), .B(n9151), .Z(n9142) );
  AND U11495 ( .A(n9152), .B(n9153), .Z(n9151) );
  NANDN U11496 ( .B(n8534), .A(n6926), .Z(n9153) );
  NANDN U11497 ( .B(n8511), .A(n6898), .Z(n9152) );
  AND U11498 ( .A(n9154), .B(n9155), .Z(n9150) );
  NANDN U11499 ( .B(n8515), .A(n6882), .Z(n9155) );
  NANDN U11500 ( .B(n8521), .A(n6809), .Z(n9154) );
  AND U11501 ( .A(n9156), .B(n9157), .Z(n9140) );
  AND U11502 ( .A(n9158), .B(n9159), .Z(n9157) );
  AND U11503 ( .A(n9160), .B(n9161), .Z(n9159) );
  NANDN U11504 ( .B(n8525), .A(n6807), .Z(n9161) );
  NANDN U11505 ( .B(n8533), .A(n6799), .Z(n9160) );
  AND U11506 ( .A(n9162), .B(n9163), .Z(n9158) );
  NANDN U11507 ( .B(n8537), .A(n6803), .Z(n9163) );
  NANDN U11508 ( .B(n8538), .A(n6823), .Z(n9162) );
  AND U11509 ( .A(n9164), .B(n9165), .Z(n9156) );
  AND U11510 ( .A(n9166), .B(n9167), .Z(n9165) );
  NANDN U11511 ( .B(n8543), .A(n6827), .Z(n9167) );
  NANDN U11512 ( .B(n8544), .A(n6833), .Z(n9166) );
  AND U11513 ( .A(n9168), .B(n9169), .Z(n9164) );
  NANDN U11514 ( .B(n8547), .A(n6835), .Z(n9169) );
  NANDN U11515 ( .B(n8548), .A(n6839), .Z(n9168) );
  AND U11516 ( .A(n9170), .B(n9171), .Z(n9138) );
  AND U11517 ( .A(n9172), .B(n9173), .Z(n9171) );
  AND U11518 ( .A(n9174), .B(n9175), .Z(n9173) );
  AND U11519 ( .A(n9176), .B(n9177), .Z(n9175) );
  NANDN U11520 ( .B(n8557), .A(n6850), .Z(n9177) );
  NANDN U11521 ( .B(n8558), .A(n6853), .Z(n9176) );
  AND U11522 ( .A(n9178), .B(n9179), .Z(n9174) );
  NANDN U11523 ( .B(n8561), .A(n6841), .Z(n9179) );
  NANDN U11524 ( .B(n8562), .A(n6857), .Z(n9178) );
  AND U11525 ( .A(n9180), .B(n9181), .Z(n9172) );
  AND U11526 ( .A(n9182), .B(n9183), .Z(n9181) );
  NANDN U11527 ( .B(n8567), .A(n6859), .Z(n9183) );
  NANDN U11528 ( .B(n8568), .A(n6865), .Z(n9182) );
  AND U11529 ( .A(n9184), .B(n9185), .Z(n9180) );
  NANDN U11530 ( .B(n8571), .A(n6967), .Z(n9185) );
  NANDN U11531 ( .B(n8572), .A(n6966), .Z(n9184) );
  AND U11532 ( .A(n9186), .B(n9187), .Z(n9170) );
  AND U11533 ( .A(n9188), .B(n9189), .Z(n9187) );
  AND U11534 ( .A(n9190), .B(n9191), .Z(n9189) );
  NANDN U11535 ( .B(n8579), .A(n6961), .Z(n9191) );
  NANDN U11536 ( .B(n8580), .A(n6956), .Z(n9190) );
  AND U11537 ( .A(n9192), .B(n9193), .Z(n9188) );
  NANDN U11538 ( .B(n8583), .A(n6960), .Z(n9193) );
  NANDN U11539 ( .B(n8584), .A(n6957), .Z(n9192) );
  AND U11540 ( .A(n9194), .B(n9195), .Z(n9186) );
  AND U11541 ( .A(n9196), .B(n9197), .Z(n9195) );
  NANDN U11542 ( .B(n8589), .A(n6947), .Z(n9197) );
  NANDN U11543 ( .B(n8590), .A(n6946), .Z(n9196) );
  AND U11544 ( .A(n9198), .B(n9199), .Z(n9194) );
  NANDN U11545 ( .B(n8593), .A(n6943), .Z(n9199) );
  NAND U11546 ( .A(n6942), .B(n6897), .Z(n9198) );
  ANDN U11547 ( .A(n9200), .B(n9201), .Z(n9012) );
  NAND U11548 ( .A(n6886), .B(n6822), .Z(n9200) );
  IV U11549 ( .A(\u_a23_core/u_execute/rn[5] ), .Z(n9067) );
  NAND U11550 ( .A(n6765), .B(\u_a23_core/u_execute/u_alu/fadder_out[5] ), .Z(
        n9058) );
  AND U11551 ( .A(n9202), .B(n9203), .Z(n9054) );
  NANDN U11552 ( .B(n8406), .A(\u_a23_core/u_execute/rn_plus4[5] ), .Z(n9203)
         );
  NANDN U11553 ( .B(n8407), .A(\u_a23_core/u_execute/alu_plus4[5] ), .Z(n9202)
         );
  AND U11554 ( .A(n9204), .B(n9205), .Z(n9052) );
  AND U11555 ( .A(n9206), .B(n9207), .Z(n9205) );
  NAND U11556 ( .A(n8412), .B(\u_a23_core/u_execute/address_plus4[5] ), .Z(
        n9207) );
  NAND U11557 ( .A(\u_a23_core/u_execute/rn[5] ), .B(n8413), .Z(n9206) );
  NAND U11558 ( .A(n9208), .B(n9209), .Z(\u_a23_core/u_execute/rn[5] ) );
  AND U11559 ( .A(n9210), .B(n9211), .Z(n9209) );
  AND U11560 ( .A(n9212), .B(n9213), .Z(n9211) );
  AND U11561 ( .A(n9214), .B(n9215), .Z(n9213) );
  NANDN U11562 ( .B(n8635), .A(\u_a23_core/u_execute/pc[5] ), .Z(n9215) );
  NANDN U11563 ( .B(n8636), .A(\u_a23_core/u_execute/u_register_bank/r14[5] ), 
        .Z(n9214) );
  AND U11564 ( .A(n9216), .B(n9217), .Z(n9212) );
  NANDN U11565 ( .B(n8639), .A(\u_a23_core/u_execute/u_register_bank/r13[5] ), 
        .Z(n9217) );
  NANDN U11566 ( .B(n8640), .A(\u_a23_core/u_execute/u_register_bank/r12[5] ), 
        .Z(n9216) );
  AND U11567 ( .A(n9218), .B(n9219), .Z(n9210) );
  AND U11568 ( .A(n9220), .B(n9221), .Z(n9219) );
  NANDN U11569 ( .B(n8645), .A(\u_a23_core/u_execute/u_register_bank/r11[5] ), 
        .Z(n9221) );
  NANDN U11570 ( .B(n8646), .A(\u_a23_core/u_execute/u_register_bank/r10[5] ), 
        .Z(n9220) );
  AND U11571 ( .A(n9222), .B(n9223), .Z(n9218) );
  NANDN U11572 ( .B(n8649), .A(\u_a23_core/u_execute/u_register_bank/r9[5] ), 
        .Z(n9223) );
  NANDN U11573 ( .B(n8650), .A(\u_a23_core/u_execute/u_register_bank/r8[5] ), 
        .Z(n9222) );
  AND U11574 ( .A(n9224), .B(n9225), .Z(n9208) );
  AND U11575 ( .A(n9226), .B(n9227), .Z(n9225) );
  AND U11576 ( .A(n9228), .B(n9229), .Z(n9227) );
  NANDN U11577 ( .B(n8657), .A(\u_a23_core/u_execute/u_register_bank/r7[5] ), 
        .Z(n9229) );
  NANDN U11578 ( .B(n8658), .A(\u_a23_core/u_execute/u_register_bank/r6[5] ), 
        .Z(n9228) );
  AND U11579 ( .A(n9230), .B(n9231), .Z(n9226) );
  NANDN U11580 ( .B(n8661), .A(\u_a23_core/u_execute/u_register_bank/r5[5] ), 
        .Z(n9231) );
  NANDN U11581 ( .B(n8662), .A(\u_a23_core/u_execute/u_register_bank/r4[5] ), 
        .Z(n9230) );
  AND U11582 ( .A(n9232), .B(n9233), .Z(n9224) );
  AND U11583 ( .A(n9234), .B(n9235), .Z(n9233) );
  NANDN U11584 ( .B(n8667), .A(\u_a23_core/u_execute/u_register_bank/r3[5] ), 
        .Z(n9235) );
  NANDN U11585 ( .B(n8668), .A(\u_a23_core/u_execute/u_register_bank/r0[5] ), 
        .Z(n9234) );
  AND U11586 ( .A(n9236), .B(n9237), .Z(n9232) );
  NANDN U11587 ( .B(n8671), .A(\u_a23_core/u_execute/u_register_bank/r2[5] ), 
        .Z(n9237) );
  NANDN U11588 ( .B(n8672), .A(\u_a23_core/u_execute/u_register_bank/r1[5] ), 
        .Z(n9236) );
  AND U11589 ( .A(n9238), .B(n9239), .Z(n9204) );
  NAND U11590 ( .A(\u_a23_core/u_execute/pc[5] ), .B(n8416), .Z(n9239) );
  NAND U11591 ( .A(n8417), .B(\u_a23_core/u_execute/pc_plus4[5] ), .Z(n9238)
         );
  AND U11592 ( .A(n9240), .B(n9241), .Z(n8381) );
  NOR U11593 ( .A(\u_a23_core/execute_address_nxt[30] ), .B(
        \u_a23_core/execute_address_nxt[31] ), .Z(n9241) );
  NAND U11594 ( .A(n9242), .B(n9243), .Z(\u_a23_core/execute_address_nxt[31] )
         );
  AND U11595 ( .A(n9244), .B(n9245), .Z(n9243) );
  NANDN U11596 ( .B(n8406), .A(\u_a23_core/u_execute/rn_plus4[31] ), .Z(n9245)
         );
  AND U11597 ( .A(n9246), .B(n9247), .Z(n9244) );
  NAND U11598 ( .A(\u_a23_core/u_execute/alu_out[31] ), .B(n9248), .Z(n9247)
         );
  IV U11599 ( .A(n7052), .Z(\u_a23_core/u_execute/alu_out[31] ) );
  AND U11600 ( .A(n9249), .B(n9250), .Z(n7052) );
  MUX U11601 ( .IN0(n9251), .IN1(n9252), .SEL(n6763), .F(n9250) );
  IV U11602 ( .A(\u_a23_core/u_execute/u_alu/b_not[31] ), .Z(n6763) );
  NAND U11603 ( .A(n9253), .B(n9254), .Z(
        \u_a23_core/u_execute/u_alu/b_not[31] ) );
  MUX U11604 ( .IN0(n8430), .IN1(n8431), .SEL(n9255), .F(n9254) );
  MUX U11605 ( .IN0(n8433), .IN1(n8434), .SEL(\u_a23_core/u_execute/rn[31] ), 
        .F(n9253) );
  NAND U11606 ( .A(\u_a23_core/u_execute/u_alu/a[31] ), .B(n8400), .Z(n9252)
         );
  ANDN U11607 ( .A(n9256), .B(n9257), .Z(n9251) );
  MUX U11608 ( .IN0(n8400), .IN1(\u_a23_core/alu_function[3] ), .SEL(
        \u_a23_core/u_execute/u_alu/a[31] ), .F(n9257) );
  IV U11609 ( .A(n6764), .Z(\u_a23_core/u_execute/u_alu/a[31] ) );
  MUX U11610 ( .IN0(n9258), .IN1(n9255), .SEL(\u_a23_core/alu_function[8] ), 
        .F(n6764) );
  AND U11611 ( .A(n9259), .B(n9260), .Z(n9255) );
  AND U11612 ( .A(n9261), .B(n9262), .Z(n9260) );
  NAND U11613 ( .A(n9263), .B(n6888), .Z(n9261) );
  NAND U11614 ( .A(n9264), .B(n9265), .Z(n9263) );
  AND U11615 ( .A(n9266), .B(n9267), .Z(n9265) );
  NAND U11616 ( .A(n9268), .B(n9269), .Z(n9267) );
  AND U11617 ( .A(n6898), .B(n6988), .Z(n9269) );
  AND U11618 ( .A(n9270), .B(n9271), .Z(n9268) );
  NAND U11619 ( .A(\u_a23_core/shift_imm_zero ), .B(n6894), .Z(n9266) );
  ANDN U11620 ( .A(\u_a23_core/use_carry_in ), .B(n9272), .Z(n6894) );
  ANDN U11621 ( .A(n9273), .B(n6896), .Z(n9264) );
  NAND U11622 ( .A(n9274), .B(n9275), .Z(n6896) );
  AND U11623 ( .A(n9276), .B(n9277), .Z(n9275) );
  AND U11624 ( .A(n9278), .B(n9279), .Z(n9277) );
  AND U11625 ( .A(n9280), .B(n9281), .Z(n9279) );
  AND U11626 ( .A(n9282), .B(n9283), .Z(n9281) );
  NANDN U11627 ( .B(n8584), .A(n6919), .Z(n9283) );
  NANDN U11628 ( .B(n8589), .A(n6920), .Z(n9282) );
  AND U11629 ( .A(n9284), .B(n9285), .Z(n9280) );
  NANDN U11630 ( .B(n8516), .A(n6809), .Z(n9285) );
  NANDN U11631 ( .B(n8590), .A(n6925), .Z(n9284) );
  AND U11632 ( .A(n9286), .B(n9287), .Z(n9278) );
  AND U11633 ( .A(n9288), .B(n9289), .Z(n9287) );
  NANDN U11634 ( .B(n8522), .A(n6807), .Z(n9289) );
  NANDN U11635 ( .B(n8593), .A(n6926), .Z(n9288) );
  AND U11636 ( .A(n9290), .B(n9291), .Z(n9286) );
  NANDN U11637 ( .B(n8526), .A(n6799), .Z(n9291) );
  NANDN U11638 ( .B(n8534), .A(n6803), .Z(n9290) );
  AND U11639 ( .A(n9292), .B(n9293), .Z(n9276) );
  AND U11640 ( .A(n9294), .B(n9295), .Z(n9293) );
  AND U11641 ( .A(n9296), .B(n9297), .Z(n9295) );
  NANDN U11642 ( .B(n8511), .A(n6823), .Z(n9297) );
  NANDN U11643 ( .B(n8515), .A(n6827), .Z(n9296) );
  AND U11644 ( .A(n9298), .B(n9299), .Z(n9294) );
  NANDN U11645 ( .B(n8521), .A(n6833), .Z(n9299) );
  NANDN U11646 ( .B(n8525), .A(n6835), .Z(n9298) );
  AND U11647 ( .A(n9300), .B(n9301), .Z(n9292) );
  NANDN U11648 ( .B(n8538), .A(n6853), .Z(n9301) );
  AND U11649 ( .A(n9302), .B(n9303), .Z(n9300) );
  NANDN U11650 ( .B(n8533), .A(n6839), .Z(n9303) );
  NANDN U11651 ( .B(n8537), .A(n6850), .Z(n9302) );
  AND U11652 ( .A(n9304), .B(n9305), .Z(n9274) );
  AND U11653 ( .A(n9306), .B(n9307), .Z(n9305) );
  AND U11654 ( .A(n9308), .B(n9309), .Z(n9307) );
  AND U11655 ( .A(n9310), .B(n9311), .Z(n9309) );
  NANDN U11656 ( .B(n8543), .A(n6841), .Z(n9311) );
  NANDN U11657 ( .B(n8544), .A(n6857), .Z(n9310) );
  AND U11658 ( .A(n9312), .B(n9313), .Z(n9308) );
  NANDN U11659 ( .B(n8547), .A(n6859), .Z(n9313) );
  NANDN U11660 ( .B(n8548), .A(n6865), .Z(n9312) );
  AND U11661 ( .A(n9314), .B(n9315), .Z(n9306) );
  AND U11662 ( .A(n9316), .B(n9317), .Z(n9315) );
  NANDN U11663 ( .B(n8557), .A(n6967), .Z(n9317) );
  NANDN U11664 ( .B(n8558), .A(n6966), .Z(n9316) );
  AND U11665 ( .A(n9318), .B(n9319), .Z(n9314) );
  NANDN U11666 ( .B(n8561), .A(n6961), .Z(n9319) );
  NANDN U11667 ( .B(n8562), .A(n6956), .Z(n9318) );
  AND U11668 ( .A(n9320), .B(n9321), .Z(n9304) );
  AND U11669 ( .A(n9322), .B(n9323), .Z(n9321) );
  AND U11670 ( .A(n9324), .B(n9325), .Z(n9323) );
  NANDN U11671 ( .B(n8567), .A(n6960), .Z(n9325) );
  NANDN U11672 ( .B(n8568), .A(n6957), .Z(n9324) );
  AND U11673 ( .A(n9326), .B(n9327), .Z(n9322) );
  NANDN U11674 ( .B(n8571), .A(n6947), .Z(n9327) );
  NANDN U11675 ( .B(n8572), .A(n6946), .Z(n9326) );
  AND U11676 ( .A(n9328), .B(n9329), .Z(n9320) );
  NANDN U11677 ( .B(n8583), .A(n6937), .Z(n9329) );
  AND U11678 ( .A(n9330), .B(n9331), .Z(n9328) );
  NANDN U11679 ( .B(n8579), .A(n6943), .Z(n9331) );
  NANDN U11680 ( .B(n8580), .A(n6942), .Z(n9330) );
  NAND U11681 ( .A(n6882), .B(n8512), .Z(n9273) );
  AND U11682 ( .A(n9332), .B(n9333), .Z(n9259) );
  NAND U11683 ( .A(n9334), .B(n6902), .Z(n9333) );
  NAND U11684 ( .A(n9335), .B(n9336), .Z(n9334) );
  AND U11685 ( .A(n9337), .B(n9338), .Z(n9336) );
  AND U11686 ( .A(n9339), .B(n9340), .Z(n9338) );
  AND U11687 ( .A(n9341), .B(n9342), .Z(n9340) );
  AND U11688 ( .A(n9343), .B(n9344), .Z(n9342) );
  NAND U11689 ( .A(n6802), .B(n6920), .Z(n9344) );
  AND U11690 ( .A(n9345), .B(n9346), .Z(n9341) );
  NAND U11691 ( .A(n6925), .B(n6798), .Z(n9346) );
  NAND U11692 ( .A(n6806), .B(n6926), .Z(n9345) );
  AND U11693 ( .A(n9347), .B(n9348), .Z(n9339) );
  AND U11694 ( .A(n9349), .B(n9350), .Z(n9348) );
  NAND U11695 ( .A(n6898), .B(n6808), .Z(n9350) );
  NAND U11696 ( .A(n6882), .B(n6916), .Z(n9349) );
  AND U11697 ( .A(n9351), .B(n9352), .Z(n9347) );
  AND U11698 ( .A(n9353), .B(n9354), .Z(n9337) );
  AND U11699 ( .A(n9355), .B(n9356), .Z(n9354) );
  AND U11700 ( .A(n9357), .B(n9095), .Z(n9356) );
  NAND U11701 ( .A(n8461), .B(n6857), .Z(n9095) );
  AND U11702 ( .A(n8468), .B(n9358), .Z(n9355) );
  NAND U11703 ( .A(n6919), .B(n6822), .Z(n9358) );
  NAND U11704 ( .A(n9359), .B(n6853), .Z(n8468) );
  AND U11705 ( .A(n9360), .B(n9361), .Z(n9353) );
  AND U11706 ( .A(n9362), .B(n9363), .Z(n9361) );
  NAND U11707 ( .A(n6937), .B(n6826), .Z(n9362) );
  AND U11708 ( .A(n9364), .B(n9365), .Z(n9360) );
  NAND U11709 ( .A(n6832), .B(n6942), .Z(n9365) );
  NAND U11710 ( .A(n6834), .B(n6943), .Z(n9364) );
  AND U11711 ( .A(n9366), .B(n9367), .Z(n9335) );
  AND U11712 ( .A(n9368), .B(n9369), .Z(n9367) );
  AND U11713 ( .A(n9370), .B(n9371), .Z(n9369) );
  AND U11714 ( .A(n9372), .B(n9373), .Z(n9371) );
  NAND U11715 ( .A(n6838), .B(n6946), .Z(n9373) );
  NAND U11716 ( .A(n6840), .B(n6960), .Z(n9372) );
  AND U11717 ( .A(n9374), .B(n9375), .Z(n9370) );
  NAND U11718 ( .A(n6947), .B(n6851), .Z(n9375) );
  NAND U11719 ( .A(n6852), .B(n6957), .Z(n9374) );
  AND U11720 ( .A(n9376), .B(n9377), .Z(n9368) );
  AND U11721 ( .A(n9378), .B(n9379), .Z(n9377) );
  NAND U11722 ( .A(n6956), .B(n6856), .Z(n9379) );
  NAND U11723 ( .A(n6961), .B(n6858), .Z(n9378) );
  AND U11724 ( .A(n6862), .B(n9380), .Z(n9376) );
  NAND U11725 ( .A(n6966), .B(n6864), .Z(n9380) );
  NAND U11726 ( .A(n6967), .B(n8487), .Z(n6862) );
  AND U11727 ( .A(n9381), .B(n9382), .Z(n9366) );
  AND U11728 ( .A(n9383), .B(n9384), .Z(n9382) );
  AND U11729 ( .A(n9385), .B(n9386), .Z(n9384) );
  AND U11730 ( .A(n9387), .B(n9388), .Z(n9383) );
  AND U11731 ( .A(n9389), .B(n9390), .Z(n9381) );
  AND U11732 ( .A(n9391), .B(n9392), .Z(n9390) );
  AND U11733 ( .A(n9393), .B(n9394), .Z(n9389) );
  NAND U11734 ( .A(n6985), .B(n6893), .Z(n9332) );
  IV U11735 ( .A(\u_a23_core/u_execute/rn[31] ), .Z(n9258) );
  AND U11736 ( .A(n9395), .B(n9396), .Z(n9249) );
  NAND U11737 ( .A(n6765), .B(\u_a23_core/u_execute/u_alu/fadder_out[31] ), 
        .Z(n9396) );
  AND U11738 ( .A(n9397), .B(n9398), .Z(n9242) );
  NAND U11739 ( .A(\u_a23_core/u_execute/rn[31] ), .B(n8413), .Z(n9398) );
  NAND U11740 ( .A(n9399), .B(n9400), .Z(\u_a23_core/u_execute/rn[31] ) );
  AND U11741 ( .A(n9401), .B(n9402), .Z(n9400) );
  AND U11742 ( .A(n9403), .B(n9404), .Z(n9402) );
  AND U11743 ( .A(n9405), .B(n9406), .Z(n9404) );
  NANDN U11744 ( .B(n8636), .A(\u_a23_core/u_execute/u_register_bank/r14[31] ), 
        .Z(n9406) );
  NANDN U11745 ( .B(n8639), .A(\u_a23_core/u_execute/u_register_bank/r13[31] ), 
        .Z(n9405) );
  AND U11746 ( .A(n9407), .B(n9408), .Z(n9403) );
  NANDN U11747 ( .B(n8640), .A(\u_a23_core/u_execute/u_register_bank/r12[31] ), 
        .Z(n9408) );
  NANDN U11748 ( .B(n8645), .A(\u_a23_core/u_execute/u_register_bank/r11[31] ), 
        .Z(n9407) );
  AND U11749 ( .A(n9409), .B(n9410), .Z(n9401) );
  AND U11750 ( .A(n9411), .B(n9412), .Z(n9410) );
  NANDN U11751 ( .B(n8646), .A(\u_a23_core/u_execute/u_register_bank/r10[31] ), 
        .Z(n9412) );
  NANDN U11752 ( .B(n8649), .A(\u_a23_core/u_execute/u_register_bank/r9[31] ), 
        .Z(n9411) );
  AND U11753 ( .A(n9413), .B(n9414), .Z(n9409) );
  NANDN U11754 ( .B(n8650), .A(\u_a23_core/u_execute/u_register_bank/r8[31] ), 
        .Z(n9414) );
  NANDN U11755 ( .B(n8657), .A(\u_a23_core/u_execute/u_register_bank/r7[31] ), 
        .Z(n9413) );
  AND U11756 ( .A(n9415), .B(n9416), .Z(n9399) );
  AND U11757 ( .A(n9417), .B(n9418), .Z(n9416) );
  AND U11758 ( .A(n9419), .B(n9420), .Z(n9418) );
  NANDN U11759 ( .B(n8658), .A(\u_a23_core/u_execute/u_register_bank/r6[31] ), 
        .Z(n9420) );
  NANDN U11760 ( .B(n8661), .A(\u_a23_core/u_execute/u_register_bank/r5[31] ), 
        .Z(n9419) );
  AND U11761 ( .A(n9421), .B(n9422), .Z(n9417) );
  NANDN U11762 ( .B(n8662), .A(\u_a23_core/u_execute/u_register_bank/r4[31] ), 
        .Z(n9422) );
  NANDN U11763 ( .B(n8667), .A(\u_a23_core/u_execute/u_register_bank/r3[31] ), 
        .Z(n9421) );
  AND U11764 ( .A(n9423), .B(n9424), .Z(n9415) );
  NANDN U11765 ( .B(n8672), .A(\u_a23_core/u_execute/u_register_bank/r1[31] ), 
        .Z(n9424) );
  AND U11766 ( .A(n9425), .B(n9426), .Z(n9423) );
  NANDN U11767 ( .B(n8668), .A(\u_a23_core/u_execute/u_register_bank/r0[31] ), 
        .Z(n9426) );
  NANDN U11768 ( .B(n8671), .A(\u_a23_core/u_execute/u_register_bank/r2[31] ), 
        .Z(n9425) );
  AND U11769 ( .A(n9427), .B(n9428), .Z(n9397) );
  NANDN U11770 ( .B(n8407), .A(\u_a23_core/u_execute/alu_plus4[31] ), .Z(n9428) );
  NAND U11771 ( .A(n8412), .B(\u_a23_core/u_execute/address_plus4[31] ), .Z(
        n9427) );
  NAND U11772 ( .A(n9429), .B(n9430), .Z(\u_a23_core/execute_address_nxt[30] )
         );
  AND U11773 ( .A(n9431), .B(n9432), .Z(n9430) );
  NANDN U11774 ( .B(n8406), .A(\u_a23_core/u_execute/rn_plus4[30] ), .Z(n9432)
         );
  AND U11775 ( .A(n9246), .B(n9433), .Z(n9431) );
  NAND U11776 ( .A(\u_a23_core/u_execute/alu_out[30] ), .B(n9248), .Z(n9433)
         );
  IV U11777 ( .A(n6999), .Z(\u_a23_core/u_execute/alu_out[30] ) );
  AND U11778 ( .A(n9434), .B(n9435), .Z(n6999) );
  MUX U11779 ( .IN0(n9436), .IN1(n9437), .SEL(
        \u_a23_core/u_execute/u_alu/b_not[30] ), .F(n9435) );
  NAND U11780 ( .A(n9438), .B(n9439), .Z(
        \u_a23_core/u_execute/u_alu/b_not[30] ) );
  MUX U11781 ( .IN0(n8430), .IN1(n8431), .SEL(n9440), .F(n9439) );
  MUX U11782 ( .IN0(n8433), .IN1(n8434), .SEL(\u_a23_core/u_execute/rn[30] ), 
        .F(n9438) );
  ANDN U11783 ( .A(n9256), .B(n9441), .Z(n9437) );
  MUX U11784 ( .IN0(n8400), .IN1(\u_a23_core/alu_function[3] ), .SEL(
        \u_a23_core/u_execute/u_alu/a[30] ), .F(n9441) );
  NAND U11785 ( .A(\u_a23_core/u_execute/u_alu/a[30] ), .B(n8400), .Z(n9436)
         );
  IV U11786 ( .A(n9442), .Z(\u_a23_core/u_execute/u_alu/a[30] ) );
  MUX U11787 ( .IN0(n9443), .IN1(n9440), .SEL(\u_a23_core/alu_function[8] ), 
        .F(n9442) );
  AND U11788 ( .A(n9444), .B(n9445), .Z(n9440) );
  AND U11789 ( .A(n9446), .B(n9447), .Z(n9445) );
  NAND U11790 ( .A(n9448), .B(n6902), .Z(n9447) );
  NAND U11791 ( .A(n9449), .B(n9450), .Z(n9448) );
  AND U11792 ( .A(n9451), .B(n9452), .Z(n9450) );
  AND U11793 ( .A(n9453), .B(n9454), .Z(n9452) );
  AND U11794 ( .A(n9455), .B(n9456), .Z(n9454) );
  AND U11795 ( .A(n9457), .B(n9458), .Z(n9456) );
  NAND U11796 ( .A(n6802), .B(n6925), .Z(n9458) );
  AND U11797 ( .A(n9459), .B(n9460), .Z(n9455) );
  NAND U11798 ( .A(n6926), .B(n6798), .Z(n9460) );
  NAND U11799 ( .A(n6806), .B(n6898), .Z(n9459) );
  AND U11800 ( .A(n9461), .B(n9462), .Z(n9453) );
  AND U11801 ( .A(n9463), .B(n9464), .Z(n9462) );
  NAND U11802 ( .A(n6916), .B(n6809), .Z(n9464) );
  AND U11803 ( .A(n9465), .B(n9466), .Z(n9461) );
  AND U11804 ( .A(n9467), .B(n9468), .Z(n9451) );
  AND U11805 ( .A(n9469), .B(n9470), .Z(n9468) );
  AND U11806 ( .A(n9471), .B(n8984), .Z(n9470) );
  NAND U11807 ( .A(n8470), .B(n6857), .Z(n8984) );
  NAND U11808 ( .A(n6920), .B(n6822), .Z(n9471) );
  AND U11809 ( .A(n9472), .B(n8715), .Z(n9469) );
  NAND U11810 ( .A(n9359), .B(n6841), .Z(n8715) );
  NAND U11811 ( .A(n6919), .B(n6826), .Z(n9472) );
  AND U11812 ( .A(n9473), .B(n9474), .Z(n9467) );
  AND U11813 ( .A(n9475), .B(n9476), .Z(n9474) );
  NAND U11814 ( .A(n6832), .B(n6937), .Z(n9476) );
  NAND U11815 ( .A(n6834), .B(n6942), .Z(n9475) );
  AND U11816 ( .A(n9477), .B(n9478), .Z(n9473) );
  NAND U11817 ( .A(n6838), .B(n6943), .Z(n9478) );
  NAND U11818 ( .A(n6840), .B(n6957), .Z(n9477) );
  AND U11819 ( .A(n9479), .B(n9480), .Z(n9449) );
  AND U11820 ( .A(n9481), .B(n9482), .Z(n9480) );
  AND U11821 ( .A(n9483), .B(n9484), .Z(n9482) );
  AND U11822 ( .A(n9485), .B(n9486), .Z(n9484) );
  NAND U11823 ( .A(n6946), .B(n6851), .Z(n9486) );
  NAND U11824 ( .A(n6852), .B(n6947), .Z(n9485) );
  AND U11825 ( .A(n9487), .B(n9488), .Z(n9483) );
  NAND U11826 ( .A(n6856), .B(n6960), .Z(n9488) );
  NAND U11827 ( .A(n6956), .B(n6858), .Z(n9487) );
  AND U11828 ( .A(n9489), .B(n9490), .Z(n9481) );
  AND U11829 ( .A(n9491), .B(n9492), .Z(n9490) );
  NAND U11830 ( .A(n6961), .B(n6864), .Z(n9492) );
  NAND U11831 ( .A(n6966), .B(n8487), .Z(n9491) );
  AND U11832 ( .A(n9493), .B(n9494), .Z(n9489) );
  AND U11833 ( .A(n9495), .B(n9496), .Z(n9479) );
  AND U11834 ( .A(n9497), .B(n9498), .Z(n9496) );
  AND U11835 ( .A(n9499), .B(n9500), .Z(n9498) );
  AND U11836 ( .A(n9501), .B(n9502), .Z(n9497) );
  AND U11837 ( .A(n9503), .B(n9504), .Z(n9495) );
  AND U11838 ( .A(n9505), .B(n9506), .Z(n9503) );
  AND U11839 ( .A(n9507), .B(n9508), .Z(n9446) );
  NAND U11840 ( .A(n6886), .B(n9509), .Z(n9508) );
  NAND U11841 ( .A(n9510), .B(n9511), .Z(n9509) );
  AND U11842 ( .A(n9512), .B(n9513), .Z(n9511) );
  IV U11843 ( .A(n9135), .Z(n9513) );
  IV U11844 ( .A(n6984), .Z(n9512) );
  AND U11845 ( .A(n9514), .B(n9515), .Z(n9510) );
  NAND U11846 ( .A(n9516), .B(n6888), .Z(n9507) );
  NAND U11847 ( .A(n9517), .B(n9518), .Z(n9516) );
  AND U11848 ( .A(n9519), .B(n9520), .Z(n9518) );
  AND U11849 ( .A(n9521), .B(n9522), .Z(n9520) );
  AND U11850 ( .A(n9523), .B(n9524), .Z(n9522) );
  AND U11851 ( .A(n9525), .B(n9526), .Z(n9524) );
  NANDN U11852 ( .B(n8583), .A(n6919), .Z(n9526) );
  NAND U11853 ( .A(n6809), .B(n8512), .Z(n9525) );
  AND U11854 ( .A(n9527), .B(n9528), .Z(n9523) );
  NANDN U11855 ( .B(n8584), .A(n6920), .Z(n9528) );
  NANDN U11856 ( .B(n8516), .A(n6807), .Z(n9527) );
  AND U11857 ( .A(n9529), .B(n9530), .Z(n9521) );
  AND U11858 ( .A(n9531), .B(n9532), .Z(n9530) );
  NANDN U11859 ( .B(n8589), .A(n6925), .Z(n9532) );
  NANDN U11860 ( .B(n8522), .A(n6799), .Z(n9531) );
  AND U11861 ( .A(n9533), .B(n9534), .Z(n9529) );
  NANDN U11862 ( .B(n8590), .A(n6926), .Z(n9534) );
  NANDN U11863 ( .B(n8526), .A(n6803), .Z(n9533) );
  AND U11864 ( .A(n9535), .B(n9536), .Z(n9519) );
  AND U11865 ( .A(n9537), .B(n9538), .Z(n9536) );
  AND U11866 ( .A(n9539), .B(n9540), .Z(n9538) );
  NANDN U11867 ( .B(n8593), .A(n6898), .Z(n9540) );
  NANDN U11868 ( .B(n8534), .A(n6823), .Z(n9539) );
  AND U11869 ( .A(n9541), .B(n9542), .Z(n9537) );
  NANDN U11870 ( .B(n8511), .A(n6827), .Z(n9542) );
  NAND U11871 ( .A(n6882), .B(n6897), .Z(n9541) );
  AND U11872 ( .A(n9543), .B(n9544), .Z(n9535) );
  AND U11873 ( .A(n9545), .B(n9546), .Z(n9544) );
  NANDN U11874 ( .B(n8515), .A(n6833), .Z(n9546) );
  NANDN U11875 ( .B(n8521), .A(n6835), .Z(n9545) );
  AND U11876 ( .A(n9547), .B(n9548), .Z(n9543) );
  NANDN U11877 ( .B(n8525), .A(n6839), .Z(n9548) );
  NANDN U11878 ( .B(n8533), .A(n6850), .Z(n9547) );
  AND U11879 ( .A(n9549), .B(n9550), .Z(n9517) );
  AND U11880 ( .A(n9551), .B(n9552), .Z(n9550) );
  AND U11881 ( .A(n9553), .B(n9554), .Z(n9552) );
  AND U11882 ( .A(n9555), .B(n9556), .Z(n9554) );
  NANDN U11883 ( .B(n8537), .A(n6853), .Z(n9556) );
  NANDN U11884 ( .B(n8538), .A(n6841), .Z(n9555) );
  AND U11885 ( .A(n9557), .B(n9558), .Z(n9553) );
  NANDN U11886 ( .B(n8543), .A(n6857), .Z(n9558) );
  NANDN U11887 ( .B(n8544), .A(n6859), .Z(n9557) );
  AND U11888 ( .A(n9559), .B(n9560), .Z(n9551) );
  AND U11889 ( .A(n9561), .B(n9562), .Z(n9560) );
  NANDN U11890 ( .B(n8547), .A(n6865), .Z(n9562) );
  NANDN U11891 ( .B(n8548), .A(n6967), .Z(n9561) );
  AND U11892 ( .A(n9563), .B(n9564), .Z(n9559) );
  NANDN U11893 ( .B(n8557), .A(n6966), .Z(n9564) );
  NANDN U11894 ( .B(n8558), .A(n6961), .Z(n9563) );
  AND U11895 ( .A(n9565), .B(n9566), .Z(n9549) );
  AND U11896 ( .A(n9567), .B(n9568), .Z(n9566) );
  AND U11897 ( .A(n9569), .B(n9570), .Z(n9568) );
  NANDN U11898 ( .B(n8561), .A(n6956), .Z(n9570) );
  NANDN U11899 ( .B(n8562), .A(n6960), .Z(n9569) );
  AND U11900 ( .A(n9571), .B(n9572), .Z(n9567) );
  NANDN U11901 ( .B(n8567), .A(n6957), .Z(n9572) );
  NANDN U11902 ( .B(n8568), .A(n6947), .Z(n9571) );
  AND U11903 ( .A(n9573), .B(n9574), .Z(n9565) );
  AND U11904 ( .A(n9575), .B(n9576), .Z(n9574) );
  NANDN U11905 ( .B(n8571), .A(n6946), .Z(n9576) );
  NANDN U11906 ( .B(n8572), .A(n6943), .Z(n9575) );
  AND U11907 ( .A(n9577), .B(n9578), .Z(n9573) );
  NANDN U11908 ( .B(n8579), .A(n6942), .Z(n9578) );
  NANDN U11909 ( .B(n8580), .A(n6937), .Z(n9577) );
  AND U11910 ( .A(n9579), .B(n9580), .Z(n9444) );
  NAND U11911 ( .A(n6984), .B(n6985), .Z(n9580) );
  NAND U11912 ( .A(n6893), .B(n6809), .Z(n9579) );
  IV U11913 ( .A(\u_a23_core/u_execute/rn[30] ), .Z(n9443) );
  AND U11914 ( .A(n9395), .B(n9581), .Z(n9434) );
  NAND U11915 ( .A(n6765), .B(\u_a23_core/u_execute/u_alu/fadder_out[30] ), 
        .Z(n9581) );
  AND U11916 ( .A(n9582), .B(n9583), .Z(n9429) );
  NAND U11917 ( .A(\u_a23_core/u_execute/rn[30] ), .B(n8413), .Z(n9583) );
  NAND U11918 ( .A(n9584), .B(n9585), .Z(\u_a23_core/u_execute/rn[30] ) );
  AND U11919 ( .A(n9586), .B(n9587), .Z(n9585) );
  AND U11920 ( .A(n9588), .B(n9589), .Z(n9587) );
  AND U11921 ( .A(n9590), .B(n9591), .Z(n9589) );
  NANDN U11922 ( .B(n8636), .A(\u_a23_core/u_execute/u_register_bank/r14[30] ), 
        .Z(n9591) );
  NANDN U11923 ( .B(n8639), .A(\u_a23_core/u_execute/u_register_bank/r13[30] ), 
        .Z(n9590) );
  AND U11924 ( .A(n9592), .B(n9593), .Z(n9588) );
  NANDN U11925 ( .B(n8640), .A(\u_a23_core/u_execute/u_register_bank/r12[30] ), 
        .Z(n9593) );
  NANDN U11926 ( .B(n8645), .A(\u_a23_core/u_execute/u_register_bank/r11[30] ), 
        .Z(n9592) );
  AND U11927 ( .A(n9594), .B(n9595), .Z(n9586) );
  AND U11928 ( .A(n9596), .B(n9597), .Z(n9595) );
  NANDN U11929 ( .B(n8646), .A(\u_a23_core/u_execute/u_register_bank/r10[30] ), 
        .Z(n9597) );
  NANDN U11930 ( .B(n8649), .A(\u_a23_core/u_execute/u_register_bank/r9[30] ), 
        .Z(n9596) );
  AND U11931 ( .A(n9598), .B(n9599), .Z(n9594) );
  NANDN U11932 ( .B(n8650), .A(\u_a23_core/u_execute/u_register_bank/r8[30] ), 
        .Z(n9599) );
  NANDN U11933 ( .B(n8657), .A(\u_a23_core/u_execute/u_register_bank/r7[30] ), 
        .Z(n9598) );
  AND U11934 ( .A(n9600), .B(n9601), .Z(n9584) );
  AND U11935 ( .A(n9602), .B(n9603), .Z(n9601) );
  AND U11936 ( .A(n9604), .B(n9605), .Z(n9603) );
  NANDN U11937 ( .B(n8658), .A(\u_a23_core/u_execute/u_register_bank/r6[30] ), 
        .Z(n9605) );
  NANDN U11938 ( .B(n8661), .A(\u_a23_core/u_execute/u_register_bank/r5[30] ), 
        .Z(n9604) );
  AND U11939 ( .A(n9606), .B(n9607), .Z(n9602) );
  NANDN U11940 ( .B(n8662), .A(\u_a23_core/u_execute/u_register_bank/r4[30] ), 
        .Z(n9607) );
  NANDN U11941 ( .B(n8667), .A(\u_a23_core/u_execute/u_register_bank/r3[30] ), 
        .Z(n9606) );
  AND U11942 ( .A(n9608), .B(n9609), .Z(n9600) );
  NANDN U11943 ( .B(n8672), .A(\u_a23_core/u_execute/u_register_bank/r1[30] ), 
        .Z(n9609) );
  AND U11944 ( .A(n9610), .B(n9611), .Z(n9608) );
  NANDN U11945 ( .B(n8668), .A(\u_a23_core/u_execute/u_register_bank/r0[30] ), 
        .Z(n9611) );
  NANDN U11946 ( .B(n8671), .A(\u_a23_core/u_execute/u_register_bank/r2[30] ), 
        .Z(n9610) );
  AND U11947 ( .A(n9612), .B(n9613), .Z(n9582) );
  NANDN U11948 ( .B(n8407), .A(\u_a23_core/u_execute/alu_plus4[30] ), .Z(n9613) );
  NAND U11949 ( .A(n8412), .B(\u_a23_core/u_execute/address_plus4[30] ), .Z(
        n9612) );
  NOR U11950 ( .A(\u_a23_core/execute_address_nxt[28] ), .B(
        \u_a23_core/execute_address_nxt[29] ), .Z(n9240) );
  NAND U11951 ( .A(n9614), .B(n9615), .Z(\u_a23_core/execute_address_nxt[29] )
         );
  AND U11952 ( .A(n9616), .B(n9617), .Z(n9615) );
  NANDN U11953 ( .B(n8406), .A(\u_a23_core/u_execute/rn_plus4[29] ), .Z(n9617)
         );
  AND U11954 ( .A(n9246), .B(n9618), .Z(n9616) );
  NAND U11955 ( .A(\u_a23_core/u_execute/alu_out[29] ), .B(n9248), .Z(n9618)
         );
  IV U11956 ( .A(n7053), .Z(\u_a23_core/u_execute/alu_out[29] ) );
  AND U11957 ( .A(n9619), .B(n9620), .Z(n7053) );
  MUX U11958 ( .IN0(n9621), .IN1(n9622), .SEL(
        \u_a23_core/u_execute/u_alu/b_not[29] ), .F(n9620) );
  NAND U11959 ( .A(n9623), .B(n9624), .Z(
        \u_a23_core/u_execute/u_alu/b_not[29] ) );
  MUX U11960 ( .IN0(n8430), .IN1(n8431), .SEL(n9625), .F(n9624) );
  MUX U11961 ( .IN0(n8433), .IN1(n8434), .SEL(\u_a23_core/u_execute/rn[29] ), 
        .F(n9623) );
  ANDN U11962 ( .A(n9256), .B(n9626), .Z(n9622) );
  MUX U11963 ( .IN0(n8400), .IN1(\u_a23_core/alu_function[3] ), .SEL(
        \u_a23_core/u_execute/u_alu/a[29] ), .F(n9626) );
  NAND U11964 ( .A(\u_a23_core/u_execute/u_alu/a[29] ), .B(n8400), .Z(n9621)
         );
  IV U11965 ( .A(n9627), .Z(\u_a23_core/u_execute/u_alu/a[29] ) );
  MUX U11966 ( .IN0(n9628), .IN1(n9625), .SEL(\u_a23_core/alu_function[8] ), 
        .F(n9627) );
  AND U11967 ( .A(n9629), .B(n9630), .Z(n9625) );
  AND U11968 ( .A(n9631), .B(n9632), .Z(n9630) );
  AND U11969 ( .A(n9633), .B(n9634), .Z(n9631) );
  NAND U11970 ( .A(n6786), .B(n9635), .Z(n9634) );
  NAND U11971 ( .A(n9636), .B(n9343), .Z(n9635) );
  NAND U11972 ( .A(n6984), .B(n6809), .Z(n9343) );
  NAND U11973 ( .A(n6893), .B(n6807), .Z(n9636) );
  NAND U11974 ( .A(n9135), .B(n9637), .Z(n9633) );
  NAND U11975 ( .A(n9262), .B(n9638), .Z(n9637) );
  IV U11976 ( .A(n6985), .Z(n9638) );
  AND U11977 ( .A(n9639), .B(n9640), .Z(n9629) );
  NAND U11978 ( .A(n9641), .B(n6888), .Z(n9640) );
  NAND U11979 ( .A(n9642), .B(n9643), .Z(n9641) );
  AND U11980 ( .A(n9644), .B(n9645), .Z(n9643) );
  AND U11981 ( .A(n9646), .B(n9647), .Z(n9645) );
  AND U11982 ( .A(n9648), .B(n9649), .Z(n9647) );
  AND U11983 ( .A(n9650), .B(n9651), .Z(n9649) );
  NANDN U11984 ( .B(n8580), .A(n6919), .Z(n9651) );
  NAND U11985 ( .A(n6807), .B(n8512), .Z(n9650) );
  AND U11986 ( .A(n9652), .B(n9653), .Z(n9648) );
  NANDN U11987 ( .B(n8583), .A(n6920), .Z(n9653) );
  NANDN U11988 ( .B(n8516), .A(n6799), .Z(n9652) );
  AND U11989 ( .A(n9654), .B(n9655), .Z(n9646) );
  AND U11990 ( .A(n9656), .B(n9657), .Z(n9655) );
  NANDN U11991 ( .B(n8584), .A(n6925), .Z(n9657) );
  NANDN U11992 ( .B(n8522), .A(n6803), .Z(n9656) );
  AND U11993 ( .A(n9658), .B(n9659), .Z(n9654) );
  NANDN U11994 ( .B(n8589), .A(n6926), .Z(n9659) );
  NANDN U11995 ( .B(n8526), .A(n6823), .Z(n9658) );
  AND U11996 ( .A(n9660), .B(n9661), .Z(n9644) );
  AND U11997 ( .A(n9662), .B(n9663), .Z(n9661) );
  AND U11998 ( .A(n9664), .B(n9665), .Z(n9663) );
  NANDN U11999 ( .B(n8590), .A(n6898), .Z(n9665) );
  NANDN U12000 ( .B(n8534), .A(n6827), .Z(n9664) );
  AND U12001 ( .A(n9666), .B(n9667), .Z(n9662) );
  NANDN U12002 ( .B(n8511), .A(n6833), .Z(n9667) );
  NANDN U12003 ( .B(n8593), .A(n6882), .Z(n9666) );
  AND U12004 ( .A(n9668), .B(n9669), .Z(n9660) );
  AND U12005 ( .A(n9670), .B(n9671), .Z(n9669) );
  NANDN U12006 ( .B(n8515), .A(n6835), .Z(n9671) );
  NAND U12007 ( .A(n6809), .B(n6897), .Z(n9670) );
  AND U12008 ( .A(n9672), .B(n9673), .Z(n9668) );
  NANDN U12009 ( .B(n8521), .A(n6839), .Z(n9673) );
  NANDN U12010 ( .B(n8525), .A(n6850), .Z(n9672) );
  AND U12011 ( .A(n9674), .B(n9675), .Z(n9642) );
  AND U12012 ( .A(n9676), .B(n9677), .Z(n9675) );
  AND U12013 ( .A(n9678), .B(n9679), .Z(n9677) );
  AND U12014 ( .A(n9680), .B(n9681), .Z(n9679) );
  NANDN U12015 ( .B(n8533), .A(n6853), .Z(n9681) );
  NANDN U12016 ( .B(n8537), .A(n6841), .Z(n9680) );
  AND U12017 ( .A(n9682), .B(n9683), .Z(n9678) );
  NANDN U12018 ( .B(n8538), .A(n6857), .Z(n9683) );
  NANDN U12019 ( .B(n8543), .A(n6859), .Z(n9682) );
  AND U12020 ( .A(n9684), .B(n9685), .Z(n9676) );
  AND U12021 ( .A(n9686), .B(n9687), .Z(n9685) );
  NANDN U12022 ( .B(n8544), .A(n6865), .Z(n9687) );
  NANDN U12023 ( .B(n8547), .A(n6967), .Z(n9686) );
  AND U12024 ( .A(n9688), .B(n9689), .Z(n9684) );
  NANDN U12025 ( .B(n8548), .A(n6966), .Z(n9689) );
  NANDN U12026 ( .B(n8557), .A(n6961), .Z(n9688) );
  AND U12027 ( .A(n9690), .B(n9691), .Z(n9674) );
  AND U12028 ( .A(n9692), .B(n9693), .Z(n9691) );
  AND U12029 ( .A(n9694), .B(n9695), .Z(n9693) );
  NANDN U12030 ( .B(n8558), .A(n6956), .Z(n9695) );
  NANDN U12031 ( .B(n8561), .A(n6960), .Z(n9694) );
  AND U12032 ( .A(n9696), .B(n9697), .Z(n9692) );
  NANDN U12033 ( .B(n8562), .A(n6957), .Z(n9697) );
  NANDN U12034 ( .B(n8567), .A(n6947), .Z(n9696) );
  AND U12035 ( .A(n9698), .B(n9699), .Z(n9690) );
  AND U12036 ( .A(n9700), .B(n9701), .Z(n9699) );
  NANDN U12037 ( .B(n8568), .A(n6946), .Z(n9701) );
  NANDN U12038 ( .B(n8571), .A(n6943), .Z(n9700) );
  AND U12039 ( .A(n9702), .B(n9703), .Z(n9698) );
  NANDN U12040 ( .B(n8572), .A(n6942), .Z(n9703) );
  NANDN U12041 ( .B(n8579), .A(n6937), .Z(n9702) );
  NAND U12042 ( .A(n9704), .B(n6902), .Z(n9639) );
  NAND U12043 ( .A(n9705), .B(n9706), .Z(n9704) );
  AND U12044 ( .A(n9707), .B(n9708), .Z(n9706) );
  AND U12045 ( .A(n9709), .B(n9710), .Z(n9708) );
  AND U12046 ( .A(n9711), .B(n9712), .Z(n9710) );
  AND U12047 ( .A(n9713), .B(n9714), .Z(n9712) );
  NAND U12048 ( .A(n6802), .B(n6926), .Z(n9714) );
  NAND U12049 ( .A(n6898), .B(n6798), .Z(n9713) );
  AND U12050 ( .A(n6813), .B(n9715), .Z(n9711) );
  NAND U12051 ( .A(n6916), .B(n6807), .Z(n9715) );
  NAND U12052 ( .A(n8464), .B(n6966), .Z(n6813) );
  AND U12053 ( .A(n9716), .B(n9717), .Z(n9709) );
  AND U12054 ( .A(n9718), .B(n9719), .Z(n9717) );
  AND U12055 ( .A(n9720), .B(n9094), .Z(n9716) );
  NAND U12056 ( .A(n8470), .B(n6859), .Z(n9094) );
  NAND U12057 ( .A(n6925), .B(n6822), .Z(n9720) );
  AND U12058 ( .A(n9721), .B(n9722), .Z(n9707) );
  AND U12059 ( .A(n9723), .B(n9724), .Z(n9722) );
  AND U12060 ( .A(n8467), .B(n9725), .Z(n9724) );
  NAND U12061 ( .A(n9726), .B(n6841), .Z(n8467) );
  AND U12062 ( .A(n9727), .B(n9728), .Z(n9723) );
  NAND U12063 ( .A(n6920), .B(n6826), .Z(n9728) );
  NAND U12064 ( .A(n6832), .B(n6919), .Z(n9727) );
  AND U12065 ( .A(n9729), .B(n9730), .Z(n9721) );
  NAND U12066 ( .A(n6840), .B(n6947), .Z(n9730) );
  AND U12067 ( .A(n9731), .B(n9732), .Z(n9729) );
  NAND U12068 ( .A(n6834), .B(n6937), .Z(n9732) );
  NAND U12069 ( .A(n6838), .B(n6942), .Z(n9731) );
  AND U12070 ( .A(n9733), .B(n9734), .Z(n9705) );
  AND U12071 ( .A(n9735), .B(n9736), .Z(n9734) );
  AND U12072 ( .A(n9737), .B(n9738), .Z(n9736) );
  AND U12073 ( .A(n9739), .B(n9740), .Z(n9738) );
  NAND U12074 ( .A(n6943), .B(n6851), .Z(n9740) );
  NAND U12075 ( .A(n6852), .B(n6946), .Z(n9739) );
  AND U12076 ( .A(n9741), .B(n9742), .Z(n9737) );
  NAND U12077 ( .A(n6856), .B(n6957), .Z(n9742) );
  NAND U12078 ( .A(n6858), .B(n6960), .Z(n9741) );
  AND U12079 ( .A(n9743), .B(n9744), .Z(n9735) );
  AND U12080 ( .A(n9745), .B(n9746), .Z(n9744) );
  NAND U12081 ( .A(n6956), .B(n6864), .Z(n9746) );
  NAND U12082 ( .A(n6961), .B(n8487), .Z(n9745) );
  AND U12083 ( .A(n9747), .B(n9748), .Z(n9743) );
  AND U12084 ( .A(n9749), .B(n9750), .Z(n9733) );
  AND U12085 ( .A(n9751), .B(n9752), .Z(n9750) );
  AND U12086 ( .A(n9753), .B(n9754), .Z(n9752) );
  AND U12087 ( .A(n9755), .B(n9756), .Z(n9751) );
  AND U12088 ( .A(n9757), .B(n9758), .Z(n9749) );
  AND U12089 ( .A(n9759), .B(n9760), .Z(n9757) );
  IV U12090 ( .A(\u_a23_core/u_execute/rn[29] ), .Z(n9628) );
  AND U12091 ( .A(n9395), .B(n9761), .Z(n9619) );
  NAND U12092 ( .A(n6765), .B(\u_a23_core/u_execute/u_alu/fadder_out[29] ), 
        .Z(n9761) );
  AND U12093 ( .A(n9762), .B(n9763), .Z(n9614) );
  NAND U12094 ( .A(\u_a23_core/u_execute/rn[29] ), .B(n8413), .Z(n9763) );
  NAND U12095 ( .A(n9764), .B(n9765), .Z(\u_a23_core/u_execute/rn[29] ) );
  AND U12096 ( .A(n9766), .B(n9767), .Z(n9765) );
  AND U12097 ( .A(n9768), .B(n9769), .Z(n9767) );
  AND U12098 ( .A(n9770), .B(n9771), .Z(n9769) );
  NANDN U12099 ( .B(n8636), .A(\u_a23_core/u_execute/u_register_bank/r14[29] ), 
        .Z(n9771) );
  NANDN U12100 ( .B(n8639), .A(\u_a23_core/u_execute/u_register_bank/r13[29] ), 
        .Z(n9770) );
  AND U12101 ( .A(n9772), .B(n9773), .Z(n9768) );
  NANDN U12102 ( .B(n8640), .A(\u_a23_core/u_execute/u_register_bank/r12[29] ), 
        .Z(n9773) );
  NANDN U12103 ( .B(n8645), .A(\u_a23_core/u_execute/u_register_bank/r11[29] ), 
        .Z(n9772) );
  AND U12104 ( .A(n9774), .B(n9775), .Z(n9766) );
  AND U12105 ( .A(n9776), .B(n9777), .Z(n9775) );
  NANDN U12106 ( .B(n8646), .A(\u_a23_core/u_execute/u_register_bank/r10[29] ), 
        .Z(n9777) );
  NANDN U12107 ( .B(n8649), .A(\u_a23_core/u_execute/u_register_bank/r9[29] ), 
        .Z(n9776) );
  AND U12108 ( .A(n9778), .B(n9779), .Z(n9774) );
  NANDN U12109 ( .B(n8650), .A(\u_a23_core/u_execute/u_register_bank/r8[29] ), 
        .Z(n9779) );
  NANDN U12110 ( .B(n8657), .A(\u_a23_core/u_execute/u_register_bank/r7[29] ), 
        .Z(n9778) );
  AND U12111 ( .A(n9780), .B(n9781), .Z(n9764) );
  AND U12112 ( .A(n9782), .B(n9783), .Z(n9781) );
  AND U12113 ( .A(n9784), .B(n9785), .Z(n9783) );
  NANDN U12114 ( .B(n8658), .A(\u_a23_core/u_execute/u_register_bank/r6[29] ), 
        .Z(n9785) );
  NANDN U12115 ( .B(n8661), .A(\u_a23_core/u_execute/u_register_bank/r5[29] ), 
        .Z(n9784) );
  AND U12116 ( .A(n9786), .B(n9787), .Z(n9782) );
  NANDN U12117 ( .B(n8662), .A(\u_a23_core/u_execute/u_register_bank/r4[29] ), 
        .Z(n9787) );
  NANDN U12118 ( .B(n8667), .A(\u_a23_core/u_execute/u_register_bank/r3[29] ), 
        .Z(n9786) );
  AND U12119 ( .A(n9788), .B(n9789), .Z(n9780) );
  NANDN U12120 ( .B(n8672), .A(\u_a23_core/u_execute/u_register_bank/r1[29] ), 
        .Z(n9789) );
  AND U12121 ( .A(n9790), .B(n9791), .Z(n9788) );
  NANDN U12122 ( .B(n8668), .A(\u_a23_core/u_execute/u_register_bank/r0[29] ), 
        .Z(n9791) );
  NANDN U12123 ( .B(n8671), .A(\u_a23_core/u_execute/u_register_bank/r2[29] ), 
        .Z(n9790) );
  AND U12124 ( .A(n9792), .B(n9793), .Z(n9762) );
  NANDN U12125 ( .B(n8407), .A(\u_a23_core/u_execute/alu_plus4[29] ), .Z(n9793) );
  NAND U12126 ( .A(n8412), .B(\u_a23_core/u_execute/address_plus4[29] ), .Z(
        n9792) );
  NAND U12127 ( .A(n9794), .B(n9795), .Z(\u_a23_core/execute_address_nxt[28] )
         );
  AND U12128 ( .A(n9796), .B(n9797), .Z(n9795) );
  NANDN U12129 ( .B(n8406), .A(\u_a23_core/u_execute/rn_plus4[28] ), .Z(n9797)
         );
  AND U12130 ( .A(n9246), .B(n9798), .Z(n9796) );
  NAND U12131 ( .A(\u_a23_core/u_execute/alu_out[28] ), .B(n9248), .Z(n9798)
         );
  IV U12132 ( .A(n7054), .Z(\u_a23_core/u_execute/alu_out[28] ) );
  AND U12133 ( .A(n9799), .B(n9800), .Z(n7054) );
  MUX U12134 ( .IN0(n9801), .IN1(n9802), .SEL(
        \u_a23_core/u_execute/u_alu/b_not[28] ), .F(n9800) );
  NAND U12135 ( .A(n9803), .B(n9804), .Z(
        \u_a23_core/u_execute/u_alu/b_not[28] ) );
  MUX U12136 ( .IN0(n8430), .IN1(n8431), .SEL(n9805), .F(n9804) );
  MUX U12137 ( .IN0(n8433), .IN1(n8434), .SEL(\u_a23_core/u_execute/rn[28] ), 
        .F(n9803) );
  ANDN U12138 ( .A(n9256), .B(n9806), .Z(n9802) );
  MUX U12139 ( .IN0(n8400), .IN1(\u_a23_core/alu_function[3] ), .SEL(
        \u_a23_core/u_execute/u_alu/a[28] ), .F(n9806) );
  NAND U12140 ( .A(\u_a23_core/u_execute/u_alu/a[28] ), .B(n8400), .Z(n9801)
         );
  IV U12141 ( .A(n9807), .Z(\u_a23_core/u_execute/u_alu/a[28] ) );
  MUX U12142 ( .IN0(n9808), .IN1(n9805), .SEL(\u_a23_core/alu_function[8] ), 
        .F(n9807) );
  AND U12143 ( .A(n9809), .B(n9810), .Z(n9805) );
  AND U12144 ( .A(n9811), .B(n9812), .Z(n9810) );
  NAND U12145 ( .A(n9813), .B(n6888), .Z(n9812) );
  NAND U12146 ( .A(n9814), .B(n9815), .Z(n9813) );
  AND U12147 ( .A(n9816), .B(n9817), .Z(n9815) );
  AND U12148 ( .A(n9818), .B(n9819), .Z(n9817) );
  AND U12149 ( .A(n9820), .B(n9821), .Z(n9819) );
  AND U12150 ( .A(n9822), .B(n9823), .Z(n9821) );
  NANDN U12151 ( .B(n8579), .A(n6919), .Z(n9823) );
  NAND U12152 ( .A(n6799), .B(n8512), .Z(n9822) );
  AND U12153 ( .A(n9824), .B(n9825), .Z(n9820) );
  NANDN U12154 ( .B(n8580), .A(n6920), .Z(n9825) );
  NANDN U12155 ( .B(n8516), .A(n6803), .Z(n9824) );
  AND U12156 ( .A(n9826), .B(n9827), .Z(n9818) );
  AND U12157 ( .A(n9828), .B(n9829), .Z(n9827) );
  NANDN U12158 ( .B(n8583), .A(n6925), .Z(n9829) );
  NANDN U12159 ( .B(n8522), .A(n6823), .Z(n9828) );
  AND U12160 ( .A(n9830), .B(n9831), .Z(n9826) );
  NANDN U12161 ( .B(n8584), .A(n6926), .Z(n9831) );
  NANDN U12162 ( .B(n8526), .A(n6827), .Z(n9830) );
  AND U12163 ( .A(n9832), .B(n9833), .Z(n9816) );
  AND U12164 ( .A(n9834), .B(n9835), .Z(n9833) );
  AND U12165 ( .A(n9836), .B(n9837), .Z(n9835) );
  NANDN U12166 ( .B(n8589), .A(n6898), .Z(n9837) );
  NANDN U12167 ( .B(n8534), .A(n6833), .Z(n9836) );
  AND U12168 ( .A(n9838), .B(n9839), .Z(n9834) );
  NANDN U12169 ( .B(n8511), .A(n6835), .Z(n9839) );
  NANDN U12170 ( .B(n8590), .A(n6882), .Z(n9838) );
  AND U12171 ( .A(n9840), .B(n9841), .Z(n9832) );
  AND U12172 ( .A(n9842), .B(n9843), .Z(n9841) );
  NANDN U12173 ( .B(n8515), .A(n6839), .Z(n9843) );
  NANDN U12174 ( .B(n8593), .A(n6809), .Z(n9842) );
  AND U12175 ( .A(n9844), .B(n9845), .Z(n9840) );
  NANDN U12176 ( .B(n8521), .A(n6850), .Z(n9845) );
  NAND U12177 ( .A(n6807), .B(n6897), .Z(n9844) );
  AND U12178 ( .A(n9846), .B(n9847), .Z(n9814) );
  AND U12179 ( .A(n9848), .B(n9849), .Z(n9847) );
  AND U12180 ( .A(n9850), .B(n9851), .Z(n9849) );
  AND U12181 ( .A(n9852), .B(n9853), .Z(n9851) );
  NANDN U12182 ( .B(n8525), .A(n6853), .Z(n9853) );
  NANDN U12183 ( .B(n8533), .A(n6841), .Z(n9852) );
  AND U12184 ( .A(n9854), .B(n9855), .Z(n9850) );
  NANDN U12185 ( .B(n8537), .A(n6857), .Z(n9855) );
  NANDN U12186 ( .B(n8538), .A(n6859), .Z(n9854) );
  AND U12187 ( .A(n9856), .B(n9857), .Z(n9848) );
  AND U12188 ( .A(n9858), .B(n9859), .Z(n9857) );
  NANDN U12189 ( .B(n8543), .A(n6865), .Z(n9859) );
  NANDN U12190 ( .B(n8544), .A(n6967), .Z(n9858) );
  AND U12191 ( .A(n9860), .B(n9861), .Z(n9856) );
  NANDN U12192 ( .B(n8547), .A(n6966), .Z(n9861) );
  NANDN U12193 ( .B(n8548), .A(n6961), .Z(n9860) );
  AND U12194 ( .A(n9862), .B(n9863), .Z(n9846) );
  AND U12195 ( .A(n9864), .B(n9865), .Z(n9863) );
  AND U12196 ( .A(n9866), .B(n9867), .Z(n9865) );
  NANDN U12197 ( .B(n8557), .A(n6956), .Z(n9867) );
  NANDN U12198 ( .B(n8558), .A(n6960), .Z(n9866) );
  AND U12199 ( .A(n9868), .B(n9869), .Z(n9864) );
  NANDN U12200 ( .B(n8561), .A(n6957), .Z(n9869) );
  NANDN U12201 ( .B(n8562), .A(n6947), .Z(n9868) );
  AND U12202 ( .A(n9870), .B(n9871), .Z(n9862) );
  AND U12203 ( .A(n9872), .B(n9873), .Z(n9871) );
  NANDN U12204 ( .B(n8567), .A(n6946), .Z(n9873) );
  NANDN U12205 ( .B(n8568), .A(n6943), .Z(n9872) );
  AND U12206 ( .A(n9874), .B(n9875), .Z(n9870) );
  NANDN U12207 ( .B(n8571), .A(n6942), .Z(n9875) );
  NANDN U12208 ( .B(n8572), .A(n6937), .Z(n9874) );
  AND U12209 ( .A(n9876), .B(n9632), .Z(n9811) );
  NAND U12210 ( .A(n6886), .B(n9877), .Z(n9632) );
  NAND U12211 ( .A(n9878), .B(n9514), .Z(n9877) );
  ANDN U12212 ( .A(n9879), .B(n9880), .Z(n9514) );
  IV U12213 ( .A(n9881), .Z(n9880) );
  AND U12214 ( .A(n9882), .B(n9883), .Z(n9879) );
  IV U12215 ( .A(n9082), .Z(n9883) );
  AND U12216 ( .A(n9884), .B(n9885), .Z(n9878) );
  NAND U12217 ( .A(n6786), .B(n9886), .Z(n9876) );
  NAND U12218 ( .A(n9887), .B(n9888), .Z(n9886) );
  NAND U12219 ( .A(n6893), .B(n6799), .Z(n9888) );
  AND U12220 ( .A(n9504), .B(n6983), .Z(n9887) );
  NAND U12221 ( .A(n9135), .B(n6809), .Z(n6983) );
  NAND U12222 ( .A(n6984), .B(n6807), .Z(n9504) );
  AND U12223 ( .A(n9889), .B(n9890), .Z(n9809) );
  NAND U12224 ( .A(n9891), .B(n6902), .Z(n9890) );
  NAND U12225 ( .A(n9892), .B(n9893), .Z(n9891) );
  AND U12226 ( .A(n9894), .B(n9895), .Z(n9893) );
  AND U12227 ( .A(n9896), .B(n9897), .Z(n9895) );
  AND U12228 ( .A(n9898), .B(n9899), .Z(n9897) );
  AND U12229 ( .A(n9900), .B(n9901), .Z(n9899) );
  NAND U12230 ( .A(n6802), .B(n6898), .Z(n9901) );
  NAND U12231 ( .A(n6916), .B(n6799), .Z(n9900) );
  AND U12232 ( .A(n9902), .B(n9903), .Z(n9898) );
  NAND U12233 ( .A(n6961), .B(n8464), .Z(n9903) );
  AND U12234 ( .A(n9904), .B(n9905), .Z(n9896) );
  AND U12235 ( .A(n9906), .B(n9907), .Z(n9905) );
  AND U12236 ( .A(n8983), .B(n9908), .Z(n9904) );
  NAND U12237 ( .A(n6926), .B(n6822), .Z(n9908) );
  NAND U12238 ( .A(n9359), .B(n6859), .Z(n8983) );
  AND U12239 ( .A(n9909), .B(n9910), .Z(n9894) );
  AND U12240 ( .A(n9911), .B(n9912), .Z(n9910) );
  AND U12241 ( .A(n9913), .B(n8720), .Z(n9912) );
  NAND U12242 ( .A(n9726), .B(n6857), .Z(n8720) );
  NAND U12243 ( .A(n6925), .B(n6826), .Z(n9913) );
  AND U12244 ( .A(n9914), .B(n9915), .Z(n9911) );
  NAND U12245 ( .A(n6832), .B(n6920), .Z(n9915) );
  NAND U12246 ( .A(n6834), .B(n6919), .Z(n9914) );
  AND U12247 ( .A(n9916), .B(n9917), .Z(n9909) );
  NAND U12248 ( .A(n6942), .B(n6851), .Z(n9917) );
  AND U12249 ( .A(n9918), .B(n9919), .Z(n9916) );
  NAND U12250 ( .A(n6838), .B(n6937), .Z(n9919) );
  NAND U12251 ( .A(n6840), .B(n6946), .Z(n9918) );
  AND U12252 ( .A(n9920), .B(n9921), .Z(n9892) );
  AND U12253 ( .A(n9922), .B(n9923), .Z(n9921) );
  AND U12254 ( .A(n9924), .B(n9925), .Z(n9923) );
  AND U12255 ( .A(n9926), .B(n9927), .Z(n9925) );
  NAND U12256 ( .A(n6852), .B(n6943), .Z(n9927) );
  NAND U12257 ( .A(n6856), .B(n6947), .Z(n9926) );
  AND U12258 ( .A(n9928), .B(n9929), .Z(n9924) );
  NAND U12259 ( .A(n6858), .B(n6957), .Z(n9929) );
  NAND U12260 ( .A(n6864), .B(n6960), .Z(n9928) );
  AND U12261 ( .A(n9930), .B(n9931), .Z(n9922) );
  AND U12262 ( .A(n9932), .B(n9933), .Z(n9930) );
  NAND U12263 ( .A(n6956), .B(n8487), .Z(n9933) );
  AND U12264 ( .A(n9934), .B(n9935), .Z(n9920) );
  AND U12265 ( .A(n9936), .B(n9937), .Z(n9935) );
  AND U12266 ( .A(n9938), .B(n9939), .Z(n9937) );
  AND U12267 ( .A(n9940), .B(n9941), .Z(n9936) );
  AND U12268 ( .A(n9942), .B(n9943), .Z(n9934) );
  AND U12269 ( .A(n9944), .B(n9945), .Z(n9942) );
  NAND U12270 ( .A(n9082), .B(n6985), .Z(n9889) );
  IV U12271 ( .A(\u_a23_core/u_execute/rn[28] ), .Z(n9808) );
  AND U12272 ( .A(n9395), .B(n9946), .Z(n9799) );
  NAND U12273 ( .A(n6765), .B(\u_a23_core/u_execute/u_alu/fadder_out[28] ), 
        .Z(n9946) );
  AND U12274 ( .A(n9947), .B(n9948), .Z(n9794) );
  NAND U12275 ( .A(\u_a23_core/u_execute/rn[28] ), .B(n8413), .Z(n9948) );
  NAND U12276 ( .A(n9949), .B(n9950), .Z(\u_a23_core/u_execute/rn[28] ) );
  AND U12277 ( .A(n9951), .B(n9952), .Z(n9950) );
  AND U12278 ( .A(n9953), .B(n9954), .Z(n9952) );
  AND U12279 ( .A(n9955), .B(n9956), .Z(n9954) );
  NANDN U12280 ( .B(n8636), .A(\u_a23_core/u_execute/u_register_bank/r14[28] ), 
        .Z(n9956) );
  NANDN U12281 ( .B(n8639), .A(\u_a23_core/u_execute/u_register_bank/r13[28] ), 
        .Z(n9955) );
  AND U12282 ( .A(n9957), .B(n9958), .Z(n9953) );
  NANDN U12283 ( .B(n8640), .A(\u_a23_core/u_execute/u_register_bank/r12[28] ), 
        .Z(n9958) );
  NANDN U12284 ( .B(n8645), .A(\u_a23_core/u_execute/u_register_bank/r11[28] ), 
        .Z(n9957) );
  AND U12285 ( .A(n9959), .B(n9960), .Z(n9951) );
  AND U12286 ( .A(n9961), .B(n9962), .Z(n9960) );
  NANDN U12287 ( .B(n8646), .A(\u_a23_core/u_execute/u_register_bank/r10[28] ), 
        .Z(n9962) );
  NANDN U12288 ( .B(n8649), .A(\u_a23_core/u_execute/u_register_bank/r9[28] ), 
        .Z(n9961) );
  AND U12289 ( .A(n9963), .B(n9964), .Z(n9959) );
  NANDN U12290 ( .B(n8650), .A(\u_a23_core/u_execute/u_register_bank/r8[28] ), 
        .Z(n9964) );
  NANDN U12291 ( .B(n8657), .A(\u_a23_core/u_execute/u_register_bank/r7[28] ), 
        .Z(n9963) );
  AND U12292 ( .A(n9965), .B(n9966), .Z(n9949) );
  AND U12293 ( .A(n9967), .B(n9968), .Z(n9966) );
  AND U12294 ( .A(n9969), .B(n9970), .Z(n9968) );
  NANDN U12295 ( .B(n8658), .A(\u_a23_core/u_execute/u_register_bank/r6[28] ), 
        .Z(n9970) );
  NANDN U12296 ( .B(n8661), .A(\u_a23_core/u_execute/u_register_bank/r5[28] ), 
        .Z(n9969) );
  AND U12297 ( .A(n9971), .B(n9972), .Z(n9967) );
  NANDN U12298 ( .B(n8662), .A(\u_a23_core/u_execute/u_register_bank/r4[28] ), 
        .Z(n9972) );
  NANDN U12299 ( .B(n8667), .A(\u_a23_core/u_execute/u_register_bank/r3[28] ), 
        .Z(n9971) );
  AND U12300 ( .A(n9973), .B(n9974), .Z(n9965) );
  NANDN U12301 ( .B(n8672), .A(\u_a23_core/u_execute/u_register_bank/r1[28] ), 
        .Z(n9974) );
  AND U12302 ( .A(n9975), .B(n9976), .Z(n9973) );
  NANDN U12303 ( .B(n8668), .A(\u_a23_core/u_execute/u_register_bank/r0[28] ), 
        .Z(n9976) );
  NANDN U12304 ( .B(n8671), .A(\u_a23_core/u_execute/u_register_bank/r2[28] ), 
        .Z(n9975) );
  AND U12305 ( .A(n9977), .B(n9978), .Z(n9947) );
  NANDN U12306 ( .B(n8407), .A(\u_a23_core/u_execute/alu_plus4[28] ), .Z(n9978) );
  NAND U12307 ( .A(n8412), .B(\u_a23_core/u_execute/address_plus4[28] ), .Z(
        n9977) );
  AND U12308 ( .A(n9979), .B(n9980), .Z(n8379) );
  AND U12309 ( .A(n9981), .B(n9982), .Z(n9980) );
  NOR U12310 ( .A(\u_a23_core/execute_address_nxt[26] ), .B(
        \u_a23_core/execute_address_nxt[27] ), .Z(n9982) );
  NAND U12311 ( .A(n9983), .B(n9984), .Z(\u_a23_core/execute_address_nxt[27] )
         );
  AND U12312 ( .A(n9985), .B(n9986), .Z(n9984) );
  NANDN U12313 ( .B(n8406), .A(\u_a23_core/u_execute/rn_plus4[27] ), .Z(n9986)
         );
  AND U12314 ( .A(n9246), .B(n9987), .Z(n9985) );
  NAND U12315 ( .A(\u_a23_core/u_execute/alu_out[27] ), .B(n9248), .Z(n9987)
         );
  IV U12316 ( .A(n7055), .Z(\u_a23_core/u_execute/alu_out[27] ) );
  AND U12317 ( .A(n9988), .B(n9989), .Z(n7055) );
  MUX U12318 ( .IN0(n9990), .IN1(n9991), .SEL(
        \u_a23_core/u_execute/u_alu/b_not[27] ), .F(n9989) );
  NAND U12319 ( .A(n9992), .B(n9993), .Z(
        \u_a23_core/u_execute/u_alu/b_not[27] ) );
  MUX U12320 ( .IN0(n8430), .IN1(n8431), .SEL(n9994), .F(n9993) );
  MUX U12321 ( .IN0(n8433), .IN1(n8434), .SEL(\u_a23_core/u_execute/rn[27] ), 
        .F(n9992) );
  ANDN U12322 ( .A(n9256), .B(n9995), .Z(n9991) );
  MUX U12323 ( .IN0(n8400), .IN1(\u_a23_core/alu_function[3] ), .SEL(
        \u_a23_core/u_execute/u_alu/a[27] ), .F(n9995) );
  NAND U12324 ( .A(\u_a23_core/u_execute/u_alu/a[27] ), .B(n8400), .Z(n9990)
         );
  IV U12325 ( .A(n9996), .Z(\u_a23_core/u_execute/u_alu/a[27] ) );
  MUX U12326 ( .IN0(n9997), .IN1(n9994), .SEL(\u_a23_core/alu_function[8] ), 
        .F(n9996) );
  AND U12327 ( .A(n9998), .B(n9999), .Z(n9994) );
  AND U12328 ( .A(n10000), .B(n10001), .Z(n9999) );
  NAND U12329 ( .A(n10002), .B(n6888), .Z(n10001) );
  NAND U12330 ( .A(n10003), .B(n10004), .Z(n10002) );
  AND U12331 ( .A(n10005), .B(n10006), .Z(n10004) );
  AND U12332 ( .A(n10007), .B(n10008), .Z(n10006) );
  AND U12333 ( .A(n10009), .B(n10010), .Z(n10008) );
  AND U12334 ( .A(n10011), .B(n10012), .Z(n10010) );
  NANDN U12335 ( .B(n8572), .A(n6919), .Z(n10012) );
  NAND U12336 ( .A(n6803), .B(n8512), .Z(n10011) );
  AND U12337 ( .A(n10013), .B(n10014), .Z(n10009) );
  NANDN U12338 ( .B(n8579), .A(n6920), .Z(n10014) );
  NANDN U12339 ( .B(n8516), .A(n6823), .Z(n10013) );
  AND U12340 ( .A(n10015), .B(n10016), .Z(n10007) );
  AND U12341 ( .A(n10017), .B(n10018), .Z(n10016) );
  NANDN U12342 ( .B(n8580), .A(n6925), .Z(n10018) );
  NANDN U12343 ( .B(n8522), .A(n6827), .Z(n10017) );
  AND U12344 ( .A(n10019), .B(n10020), .Z(n10015) );
  NANDN U12345 ( .B(n8583), .A(n6926), .Z(n10020) );
  NANDN U12346 ( .B(n8526), .A(n6833), .Z(n10019) );
  AND U12347 ( .A(n10021), .B(n10022), .Z(n10005) );
  AND U12348 ( .A(n10023), .B(n10024), .Z(n10022) );
  AND U12349 ( .A(n10025), .B(n10026), .Z(n10024) );
  NANDN U12350 ( .B(n8584), .A(n6898), .Z(n10026) );
  NANDN U12351 ( .B(n8534), .A(n6835), .Z(n10025) );
  AND U12352 ( .A(n10027), .B(n10028), .Z(n10023) );
  NANDN U12353 ( .B(n8511), .A(n6839), .Z(n10028) );
  NANDN U12354 ( .B(n8589), .A(n6882), .Z(n10027) );
  AND U12355 ( .A(n10029), .B(n10030), .Z(n10021) );
  AND U12356 ( .A(n10031), .B(n10032), .Z(n10030) );
  NANDN U12357 ( .B(n8515), .A(n6850), .Z(n10032) );
  NANDN U12358 ( .B(n8590), .A(n6809), .Z(n10031) );
  AND U12359 ( .A(n10033), .B(n10034), .Z(n10029) );
  NANDN U12360 ( .B(n8521), .A(n6853), .Z(n10034) );
  NANDN U12361 ( .B(n8593), .A(n6807), .Z(n10033) );
  AND U12362 ( .A(n10035), .B(n10036), .Z(n10003) );
  AND U12363 ( .A(n10037), .B(n10038), .Z(n10036) );
  AND U12364 ( .A(n10039), .B(n10040), .Z(n10038) );
  AND U12365 ( .A(n10041), .B(n10042), .Z(n10040) );
  NANDN U12366 ( .B(n8525), .A(n6841), .Z(n10042) );
  NAND U12367 ( .A(n6799), .B(n6897), .Z(n10041) );
  AND U12368 ( .A(n10043), .B(n10044), .Z(n10039) );
  NANDN U12369 ( .B(n8533), .A(n6857), .Z(n10044) );
  NANDN U12370 ( .B(n8537), .A(n6859), .Z(n10043) );
  AND U12371 ( .A(n10045), .B(n10046), .Z(n10037) );
  AND U12372 ( .A(n10047), .B(n10048), .Z(n10046) );
  NANDN U12373 ( .B(n8538), .A(n6865), .Z(n10048) );
  NANDN U12374 ( .B(n8543), .A(n6967), .Z(n10047) );
  AND U12375 ( .A(n10049), .B(n10050), .Z(n10045) );
  NANDN U12376 ( .B(n8544), .A(n6966), .Z(n10050) );
  NANDN U12377 ( .B(n8547), .A(n6961), .Z(n10049) );
  AND U12378 ( .A(n10051), .B(n10052), .Z(n10035) );
  AND U12379 ( .A(n10053), .B(n10054), .Z(n10052) );
  AND U12380 ( .A(n10055), .B(n10056), .Z(n10054) );
  NANDN U12381 ( .B(n8548), .A(n6956), .Z(n10056) );
  NANDN U12382 ( .B(n8557), .A(n6960), .Z(n10055) );
  AND U12383 ( .A(n10057), .B(n10058), .Z(n10053) );
  NANDN U12384 ( .B(n8558), .A(n6957), .Z(n10058) );
  NANDN U12385 ( .B(n8561), .A(n6947), .Z(n10057) );
  AND U12386 ( .A(n10059), .B(n10060), .Z(n10051) );
  AND U12387 ( .A(n10061), .B(n10062), .Z(n10060) );
  NANDN U12388 ( .B(n8562), .A(n6946), .Z(n10062) );
  NANDN U12389 ( .B(n8567), .A(n6943), .Z(n10061) );
  AND U12390 ( .A(n10063), .B(n10064), .Z(n10059) );
  NANDN U12391 ( .B(n8568), .A(n6942), .Z(n10064) );
  NANDN U12392 ( .B(n8571), .A(n6937), .Z(n10063) );
  AND U12393 ( .A(n10065), .B(n10066), .Z(n10000) );
  NAND U12394 ( .A(n6886), .B(n10067), .Z(n10066) );
  NAND U12395 ( .A(n9881), .B(n10068), .Z(n10067) );
  AND U12396 ( .A(n9882), .B(n9515), .Z(n10068) );
  IV U12397 ( .A(n8958), .Z(n9882) );
  NAND U12398 ( .A(n6786), .B(n10069), .Z(n10065) );
  NAND U12399 ( .A(n10070), .B(n10071), .Z(n10069) );
  AND U12400 ( .A(n9393), .B(n10072), .Z(n10071) );
  NAND U12401 ( .A(n9082), .B(n6809), .Z(n10072) );
  NAND U12402 ( .A(n9135), .B(n6807), .Z(n9393) );
  AND U12403 ( .A(n10073), .B(n9758), .Z(n10070) );
  NAND U12404 ( .A(n6984), .B(n6799), .Z(n9758) );
  NAND U12405 ( .A(n6893), .B(n6803), .Z(n10073) );
  AND U12406 ( .A(n10074), .B(n10075), .Z(n9998) );
  NAND U12407 ( .A(n10076), .B(n6902), .Z(n10075) );
  NAND U12408 ( .A(n10077), .B(n10078), .Z(n10076) );
  AND U12409 ( .A(n10079), .B(n10080), .Z(n10078) );
  AND U12410 ( .A(n10081), .B(n10082), .Z(n10080) );
  AND U12411 ( .A(n10083), .B(n10084), .Z(n10082) );
  AND U12412 ( .A(n10085), .B(n10086), .Z(n10084) );
  NAND U12413 ( .A(n6916), .B(n6803), .Z(n10086) );
  NAND U12414 ( .A(n6956), .B(n8464), .Z(n10085) );
  AND U12415 ( .A(n10087), .B(n6812), .Z(n10083) );
  NAND U12416 ( .A(n8465), .B(n6961), .Z(n6812) );
  AND U12417 ( .A(n10088), .B(n9099), .Z(n10081) );
  NAND U12418 ( .A(n6865), .B(n9359), .Z(n9099) );
  AND U12419 ( .A(n10089), .B(n10090), .Z(n10088) );
  NAND U12420 ( .A(n6898), .B(n6822), .Z(n10089) );
  AND U12421 ( .A(n10091), .B(n10092), .Z(n10079) );
  AND U12422 ( .A(n10093), .B(n10094), .Z(n10092) );
  AND U12423 ( .A(n10095), .B(n10096), .Z(n10094) );
  NAND U12424 ( .A(n6926), .B(n6826), .Z(n10095) );
  AND U12425 ( .A(n10097), .B(n10098), .Z(n10093) );
  NAND U12426 ( .A(n6832), .B(n6925), .Z(n10098) );
  NAND U12427 ( .A(n6834), .B(n6920), .Z(n10097) );
  AND U12428 ( .A(n10099), .B(n10100), .Z(n10091) );
  NAND U12429 ( .A(n6937), .B(n6851), .Z(n10100) );
  AND U12430 ( .A(n10101), .B(n10102), .Z(n10099) );
  NAND U12431 ( .A(n6838), .B(n6919), .Z(n10102) );
  NAND U12432 ( .A(n6840), .B(n6943), .Z(n10101) );
  AND U12433 ( .A(n10103), .B(n10104), .Z(n10077) );
  AND U12434 ( .A(n10105), .B(n10106), .Z(n10104) );
  AND U12435 ( .A(n10107), .B(n10108), .Z(n10106) );
  AND U12436 ( .A(n10109), .B(n10110), .Z(n10108) );
  NAND U12437 ( .A(n6852), .B(n6942), .Z(n10110) );
  NAND U12438 ( .A(n6856), .B(n6946), .Z(n10109) );
  AND U12439 ( .A(n10111), .B(n10112), .Z(n10107) );
  NAND U12440 ( .A(n6858), .B(n6947), .Z(n10112) );
  NAND U12441 ( .A(n6864), .B(n6957), .Z(n10111) );
  AND U12442 ( .A(n10113), .B(n8484), .Z(n10105) );
  NAND U12443 ( .A(n8603), .B(n6857), .Z(n8484) );
  AND U12444 ( .A(n10114), .B(n10115), .Z(n10113) );
  NAND U12445 ( .A(n6960), .B(n8487), .Z(n10115) );
  AND U12446 ( .A(n10116), .B(n10117), .Z(n10103) );
  AND U12447 ( .A(n10118), .B(n10119), .Z(n10117) );
  AND U12448 ( .A(n10120), .B(n10121), .Z(n10119) );
  AND U12449 ( .A(n10122), .B(n10123), .Z(n10118) );
  AND U12450 ( .A(n10124), .B(n10125), .Z(n10116) );
  AND U12451 ( .A(n10126), .B(n10127), .Z(n10124) );
  NAND U12452 ( .A(n8958), .B(n6985), .Z(n10074) );
  IV U12453 ( .A(\u_a23_core/u_execute/rn[27] ), .Z(n9997) );
  AND U12454 ( .A(n9395), .B(n10128), .Z(n9988) );
  NAND U12455 ( .A(n6765), .B(\u_a23_core/u_execute/u_alu/fadder_out[27] ), 
        .Z(n10128) );
  AND U12456 ( .A(n10129), .B(n10130), .Z(n9983) );
  NAND U12457 ( .A(\u_a23_core/u_execute/rn[27] ), .B(n8413), .Z(n10130) );
  NAND U12458 ( .A(n10131), .B(n10132), .Z(\u_a23_core/u_execute/rn[27] ) );
  AND U12459 ( .A(n10133), .B(n10134), .Z(n10132) );
  AND U12460 ( .A(n10135), .B(n10136), .Z(n10134) );
  AND U12461 ( .A(n10137), .B(n10138), .Z(n10136) );
  NANDN U12462 ( .B(n8636), .A(\u_a23_core/u_execute/u_register_bank/r14[27] ), 
        .Z(n10138) );
  NANDN U12463 ( .B(n8639), .A(\u_a23_core/u_execute/u_register_bank/r13[27] ), 
        .Z(n10137) );
  AND U12464 ( .A(n10139), .B(n10140), .Z(n10135) );
  NANDN U12465 ( .B(n8640), .A(\u_a23_core/u_execute/u_register_bank/r12[27] ), 
        .Z(n10140) );
  NANDN U12466 ( .B(n8645), .A(\u_a23_core/u_execute/u_register_bank/r11[27] ), 
        .Z(n10139) );
  AND U12467 ( .A(n10141), .B(n10142), .Z(n10133) );
  AND U12468 ( .A(n10143), .B(n10144), .Z(n10142) );
  NANDN U12469 ( .B(n8646), .A(\u_a23_core/u_execute/u_register_bank/r10[27] ), 
        .Z(n10144) );
  NANDN U12470 ( .B(n8649), .A(\u_a23_core/u_execute/u_register_bank/r9[27] ), 
        .Z(n10143) );
  AND U12471 ( .A(n10145), .B(n10146), .Z(n10141) );
  NANDN U12472 ( .B(n8650), .A(\u_a23_core/u_execute/u_register_bank/r8[27] ), 
        .Z(n10146) );
  NANDN U12473 ( .B(n8657), .A(\u_a23_core/u_execute/u_register_bank/r7[27] ), 
        .Z(n10145) );
  AND U12474 ( .A(n10147), .B(n10148), .Z(n10131) );
  AND U12475 ( .A(n10149), .B(n10150), .Z(n10148) );
  AND U12476 ( .A(n10151), .B(n10152), .Z(n10150) );
  NANDN U12477 ( .B(n8658), .A(\u_a23_core/u_execute/u_register_bank/r6[27] ), 
        .Z(n10152) );
  NANDN U12478 ( .B(n8661), .A(\u_a23_core/u_execute/u_register_bank/r5[27] ), 
        .Z(n10151) );
  AND U12479 ( .A(n10153), .B(n10154), .Z(n10149) );
  NANDN U12480 ( .B(n8662), .A(\u_a23_core/u_execute/u_register_bank/r4[27] ), 
        .Z(n10154) );
  NANDN U12481 ( .B(n8667), .A(\u_a23_core/u_execute/u_register_bank/r3[27] ), 
        .Z(n10153) );
  AND U12482 ( .A(n10155), .B(n10156), .Z(n10147) );
  NANDN U12483 ( .B(n8672), .A(\u_a23_core/u_execute/u_register_bank/r1[27] ), 
        .Z(n10156) );
  AND U12484 ( .A(n10157), .B(n10158), .Z(n10155) );
  NANDN U12485 ( .B(n8668), .A(\u_a23_core/u_execute/u_register_bank/r0[27] ), 
        .Z(n10158) );
  NANDN U12486 ( .B(n8671), .A(\u_a23_core/u_execute/u_register_bank/r2[27] ), 
        .Z(n10157) );
  AND U12487 ( .A(n10159), .B(n10160), .Z(n10129) );
  NANDN U12488 ( .B(n8407), .A(\u_a23_core/u_execute/alu_plus4[27] ), .Z(
        n10160) );
  NAND U12489 ( .A(n8412), .B(\u_a23_core/u_execute/address_plus4[27] ), .Z(
        n10159) );
  NAND U12490 ( .A(n10161), .B(n10162), .Z(
        \u_a23_core/execute_address_nxt[26] ) );
  AND U12491 ( .A(n10163), .B(n10164), .Z(n10162) );
  AND U12492 ( .A(n9246), .B(n10165), .Z(n10164) );
  NAND U12493 ( .A(\u_a23_core/u_execute/alu_out[26] ), .B(n9248), .Z(n10165)
         );
  IV U12494 ( .A(n7058), .Z(\u_a23_core/u_execute/alu_out[26] ) );
  AND U12495 ( .A(n10166), .B(n10167), .Z(n7058) );
  MUX U12496 ( .IN0(n10168), .IN1(n10169), .SEL(
        \u_a23_core/u_execute/u_alu/b_not[26] ), .F(n10167) );
  NAND U12497 ( .A(n10170), .B(n10171), .Z(
        \u_a23_core/u_execute/u_alu/b_not[26] ) );
  MUX U12498 ( .IN0(n8430), .IN1(n8431), .SEL(n10172), .F(n10171) );
  MUX U12499 ( .IN0(n8433), .IN1(n8434), .SEL(\u_a23_core/u_execute/rn[26] ), 
        .F(n10170) );
  ANDN U12500 ( .A(n9256), .B(n10173), .Z(n10169) );
  MUX U12501 ( .IN0(n8400), .IN1(\u_a23_core/alu_function[3] ), .SEL(
        \u_a23_core/u_execute/u_alu/a[26] ), .F(n10173) );
  NAND U12502 ( .A(\u_a23_core/u_execute/u_alu/a[26] ), .B(n8400), .Z(n10168)
         );
  IV U12503 ( .A(n10174), .Z(\u_a23_core/u_execute/u_alu/a[26] ) );
  MUX U12504 ( .IN0(n10175), .IN1(n10172), .SEL(\u_a23_core/alu_function[8] ), 
        .F(n10174) );
  AND U12505 ( .A(n10176), .B(n10177), .Z(n10172) );
  AND U12506 ( .A(n10178), .B(n10179), .Z(n10177) );
  NAND U12507 ( .A(n8616), .B(n6985), .Z(n10179) );
  AND U12508 ( .A(n10180), .B(n10181), .Z(n10178) );
  NAND U12509 ( .A(n6886), .B(n10182), .Z(n10181) );
  NAND U12510 ( .A(n9515), .B(n9881), .Z(n10182) );
  AND U12511 ( .A(n10183), .B(n10184), .Z(n9881) );
  AND U12512 ( .A(n10185), .B(n10186), .Z(n10184) );
  IV U12513 ( .A(n8616), .Z(n10185) );
  ANDN U12514 ( .A(n10187), .B(n10188), .Z(n10183) );
  NAND U12515 ( .A(n6786), .B(n10189), .Z(n10180) );
  NAND U12516 ( .A(n10190), .B(n10191), .Z(n10189) );
  AND U12517 ( .A(n10192), .B(n9505), .Z(n10191) );
  NAND U12518 ( .A(n9135), .B(n6799), .Z(n9505) );
  AND U12519 ( .A(n6980), .B(n10193), .Z(n10192) );
  NAND U12520 ( .A(n8958), .B(n6809), .Z(n10193) );
  NAND U12521 ( .A(n9082), .B(n6807), .Z(n6980) );
  AND U12522 ( .A(n10194), .B(n9943), .Z(n10190) );
  NAND U12523 ( .A(n6984), .B(n6803), .Z(n9943) );
  NAND U12524 ( .A(n6893), .B(n6823), .Z(n10194) );
  AND U12525 ( .A(n10195), .B(n10196), .Z(n10176) );
  NAND U12526 ( .A(n10197), .B(n6888), .Z(n10196) );
  NAND U12527 ( .A(n10198), .B(n10199), .Z(n10197) );
  AND U12528 ( .A(n10200), .B(n10201), .Z(n10199) );
  AND U12529 ( .A(n10202), .B(n10203), .Z(n10201) );
  AND U12530 ( .A(n10204), .B(n10205), .Z(n10203) );
  AND U12531 ( .A(n10206), .B(n10207), .Z(n10205) );
  NANDN U12532 ( .B(n8571), .A(n6919), .Z(n10207) );
  NAND U12533 ( .A(n6823), .B(n8512), .Z(n10206) );
  AND U12534 ( .A(n10208), .B(n10209), .Z(n10204) );
  NANDN U12535 ( .B(n8572), .A(n6920), .Z(n10209) );
  NANDN U12536 ( .B(n8516), .A(n6827), .Z(n10208) );
  AND U12537 ( .A(n10210), .B(n10211), .Z(n10202) );
  AND U12538 ( .A(n10212), .B(n10213), .Z(n10211) );
  NANDN U12539 ( .B(n8579), .A(n6925), .Z(n10213) );
  NANDN U12540 ( .B(n8522), .A(n6833), .Z(n10212) );
  AND U12541 ( .A(n10214), .B(n10215), .Z(n10210) );
  NANDN U12542 ( .B(n8580), .A(n6926), .Z(n10215) );
  NANDN U12543 ( .B(n8526), .A(n6835), .Z(n10214) );
  AND U12544 ( .A(n10216), .B(n10217), .Z(n10200) );
  AND U12545 ( .A(n10218), .B(n10219), .Z(n10217) );
  AND U12546 ( .A(n10220), .B(n10221), .Z(n10219) );
  NANDN U12547 ( .B(n8583), .A(n6898), .Z(n10221) );
  NANDN U12548 ( .B(n8534), .A(n6839), .Z(n10220) );
  AND U12549 ( .A(n10222), .B(n10223), .Z(n10218) );
  NANDN U12550 ( .B(n8511), .A(n6850), .Z(n10223) );
  NANDN U12551 ( .B(n8584), .A(n6882), .Z(n10222) );
  AND U12552 ( .A(n10224), .B(n10225), .Z(n10216) );
  AND U12553 ( .A(n10226), .B(n10227), .Z(n10225) );
  NANDN U12554 ( .B(n8515), .A(n6853), .Z(n10227) );
  NANDN U12555 ( .B(n8589), .A(n6809), .Z(n10226) );
  AND U12556 ( .A(n10228), .B(n10229), .Z(n10224) );
  NANDN U12557 ( .B(n8521), .A(n6841), .Z(n10229) );
  NANDN U12558 ( .B(n8590), .A(n6807), .Z(n10228) );
  AND U12559 ( .A(n10230), .B(n10231), .Z(n10198) );
  AND U12560 ( .A(n10232), .B(n10233), .Z(n10231) );
  AND U12561 ( .A(n10234), .B(n10235), .Z(n10233) );
  AND U12562 ( .A(n10236), .B(n10237), .Z(n10235) );
  NANDN U12563 ( .B(n8525), .A(n6857), .Z(n10237) );
  NANDN U12564 ( .B(n8593), .A(n6799), .Z(n10236) );
  AND U12565 ( .A(n10238), .B(n10239), .Z(n10234) );
  NAND U12566 ( .A(n6803), .B(n6897), .Z(n10239) );
  NANDN U12567 ( .B(n8533), .A(n6859), .Z(n10238) );
  AND U12568 ( .A(n10240), .B(n10241), .Z(n10232) );
  AND U12569 ( .A(n10242), .B(n10243), .Z(n10241) );
  NANDN U12570 ( .B(n8537), .A(n6865), .Z(n10243) );
  NANDN U12571 ( .B(n8538), .A(n6967), .Z(n10242) );
  AND U12572 ( .A(n10244), .B(n10245), .Z(n10240) );
  NANDN U12573 ( .B(n8543), .A(n6966), .Z(n10245) );
  NANDN U12574 ( .B(n8544), .A(n6961), .Z(n10244) );
  AND U12575 ( .A(n10246), .B(n10247), .Z(n10230) );
  AND U12576 ( .A(n10248), .B(n10249), .Z(n10247) );
  AND U12577 ( .A(n10250), .B(n10251), .Z(n10249) );
  NANDN U12578 ( .B(n8547), .A(n6956), .Z(n10251) );
  NANDN U12579 ( .B(n8548), .A(n6960), .Z(n10250) );
  AND U12580 ( .A(n10252), .B(n10253), .Z(n10248) );
  NANDN U12581 ( .B(n8557), .A(n6957), .Z(n10253) );
  NANDN U12582 ( .B(n8558), .A(n6947), .Z(n10252) );
  AND U12583 ( .A(n10254), .B(n10255), .Z(n10246) );
  AND U12584 ( .A(n10256), .B(n10257), .Z(n10255) );
  NANDN U12585 ( .B(n8561), .A(n6946), .Z(n10257) );
  NANDN U12586 ( .B(n8562), .A(n6943), .Z(n10256) );
  AND U12587 ( .A(n10258), .B(n10259), .Z(n10254) );
  NANDN U12588 ( .B(n8567), .A(n6942), .Z(n10259) );
  NANDN U12589 ( .B(n8568), .A(n6937), .Z(n10258) );
  NAND U12590 ( .A(n10260), .B(n6902), .Z(n10195) );
  NAND U12591 ( .A(n10261), .B(n10262), .Z(n10260) );
  AND U12592 ( .A(n10263), .B(n10264), .Z(n10262) );
  AND U12593 ( .A(n10265), .B(n10266), .Z(n10264) );
  AND U12594 ( .A(n10267), .B(n10268), .Z(n10266) );
  AND U12595 ( .A(n8704), .B(n10269), .Z(n10268) );
  NAND U12596 ( .A(n6916), .B(n6823), .Z(n10269) );
  NAND U12597 ( .A(n8603), .B(n6859), .Z(n8704) );
  AND U12598 ( .A(n10270), .B(n10271), .Z(n10267) );
  NAND U12599 ( .A(n8464), .B(n6960), .Z(n10271) );
  NAND U12600 ( .A(n6956), .B(n8465), .Z(n10270) );
  AND U12601 ( .A(n10272), .B(n10273), .Z(n10265) );
  AND U12602 ( .A(n10274), .B(n10275), .Z(n10272) );
  AND U12603 ( .A(n10276), .B(n10277), .Z(n10263) );
  AND U12604 ( .A(n10278), .B(n10279), .Z(n10277) );
  AND U12605 ( .A(n10280), .B(n8982), .Z(n10279) );
  NAND U12606 ( .A(n6865), .B(n9726), .Z(n8982) );
  NAND U12607 ( .A(n6898), .B(n6826), .Z(n10280) );
  AND U12608 ( .A(n10281), .B(n10282), .Z(n10278) );
  NAND U12609 ( .A(n6832), .B(n6926), .Z(n10282) );
  NAND U12610 ( .A(n6834), .B(n6925), .Z(n10281) );
  AND U12611 ( .A(n10283), .B(n10284), .Z(n10276) );
  NAND U12612 ( .A(n6919), .B(n6851), .Z(n10284) );
  AND U12613 ( .A(n10285), .B(n10286), .Z(n10283) );
  NAND U12614 ( .A(n6838), .B(n6920), .Z(n10286) );
  NAND U12615 ( .A(n6840), .B(n6942), .Z(n10285) );
  AND U12616 ( .A(n10287), .B(n10288), .Z(n10261) );
  AND U12617 ( .A(n10289), .B(n10290), .Z(n10288) );
  AND U12618 ( .A(n10291), .B(n10292), .Z(n10290) );
  AND U12619 ( .A(n10293), .B(n10294), .Z(n10292) );
  NAND U12620 ( .A(n6852), .B(n6937), .Z(n10294) );
  NAND U12621 ( .A(n6856), .B(n6943), .Z(n10293) );
  AND U12622 ( .A(n10295), .B(n10296), .Z(n10291) );
  NAND U12623 ( .A(n6858), .B(n6946), .Z(n10296) );
  NAND U12624 ( .A(n6864), .B(n6947), .Z(n10295) );
  AND U12625 ( .A(n10297), .B(n10298), .Z(n10289) );
  AND U12626 ( .A(n10299), .B(n10300), .Z(n10297) );
  NAND U12627 ( .A(n6957), .B(n8487), .Z(n10300) );
  AND U12628 ( .A(n10301), .B(n10302), .Z(n10287) );
  AND U12629 ( .A(n10303), .B(n10304), .Z(n10302) );
  AND U12630 ( .A(n10305), .B(n10306), .Z(n10303) );
  AND U12631 ( .A(n10307), .B(n10308), .Z(n10301) );
  AND U12632 ( .A(n10309), .B(n10310), .Z(n10307) );
  IV U12633 ( .A(\u_a23_core/u_execute/rn[26] ), .Z(n10175) );
  AND U12634 ( .A(n9395), .B(n10311), .Z(n10166) );
  NAND U12635 ( .A(n6765), .B(\u_a23_core/u_execute/u_alu/fadder_out[26] ), 
        .Z(n10311) );
  OR U12636 ( .A(\u_a23_core/u_execute/sub_166/carry[26] ), .B(n8392), .Z(
        n9246) );
  AND U12637 ( .A(n10312), .B(n10313), .Z(n10163) );
  NANDN U12638 ( .B(n8406), .A(\u_a23_core/u_execute/rn_plus4[26] ), .Z(n10313) );
  NANDN U12639 ( .B(n8407), .A(\u_a23_core/u_execute/alu_plus4[26] ), .Z(
        n10312) );
  AND U12640 ( .A(n10314), .B(n10315), .Z(n10161) );
  NAND U12641 ( .A(n8417), .B(\u_a23_core/u_execute/pc_plus4[26] ), .Z(n10315)
         );
  AND U12642 ( .A(n10316), .B(n10317), .Z(n10314) );
  NAND U12643 ( .A(n8412), .B(\u_a23_core/u_execute/address_plus4[26] ), .Z(
        n10317) );
  NAND U12644 ( .A(\u_a23_core/u_execute/rn[26] ), .B(n8413), .Z(n10316) );
  NAND U12645 ( .A(n10318), .B(n10319), .Z(\u_a23_core/u_execute/rn[26] ) );
  AND U12646 ( .A(n10320), .B(n10321), .Z(n10319) );
  AND U12647 ( .A(n10322), .B(n10323), .Z(n10321) );
  AND U12648 ( .A(n10324), .B(n10325), .Z(n10323) );
  NANDN U12649 ( .B(n8636), .A(\u_a23_core/u_execute/u_register_bank/r14[26] ), 
        .Z(n10325) );
  NANDN U12650 ( .B(n8639), .A(\u_a23_core/u_execute/u_register_bank/r13[26] ), 
        .Z(n10324) );
  AND U12651 ( .A(n10326), .B(n10327), .Z(n10322) );
  NANDN U12652 ( .B(n8640), .A(\u_a23_core/u_execute/u_register_bank/r12[26] ), 
        .Z(n10327) );
  NANDN U12653 ( .B(n8645), .A(\u_a23_core/u_execute/u_register_bank/r11[26] ), 
        .Z(n10326) );
  AND U12654 ( .A(n10328), .B(n10329), .Z(n10320) );
  AND U12655 ( .A(n10330), .B(n10331), .Z(n10329) );
  NANDN U12656 ( .B(n8646), .A(\u_a23_core/u_execute/u_register_bank/r10[26] ), 
        .Z(n10331) );
  NANDN U12657 ( .B(n8649), .A(\u_a23_core/u_execute/u_register_bank/r9[26] ), 
        .Z(n10330) );
  AND U12658 ( .A(n10332), .B(n10333), .Z(n10328) );
  NANDN U12659 ( .B(n8650), .A(\u_a23_core/u_execute/u_register_bank/r8[26] ), 
        .Z(n10333) );
  NANDN U12660 ( .B(n8657), .A(\u_a23_core/u_execute/u_register_bank/r7[26] ), 
        .Z(n10332) );
  AND U12661 ( .A(n10334), .B(n10335), .Z(n10318) );
  AND U12662 ( .A(n10336), .B(n10337), .Z(n10335) );
  AND U12663 ( .A(n10338), .B(n10339), .Z(n10337) );
  NANDN U12664 ( .B(n8658), .A(\u_a23_core/u_execute/u_register_bank/r6[26] ), 
        .Z(n10339) );
  NANDN U12665 ( .B(n8661), .A(\u_a23_core/u_execute/u_register_bank/r5[26] ), 
        .Z(n10338) );
  AND U12666 ( .A(n10340), .B(n10341), .Z(n10336) );
  NANDN U12667 ( .B(n8662), .A(\u_a23_core/u_execute/u_register_bank/r4[26] ), 
        .Z(n10341) );
  NANDN U12668 ( .B(n8667), .A(\u_a23_core/u_execute/u_register_bank/r3[26] ), 
        .Z(n10340) );
  AND U12669 ( .A(n10342), .B(n10343), .Z(n10334) );
  NANDN U12670 ( .B(n8672), .A(\u_a23_core/u_execute/u_register_bank/r1[26] ), 
        .Z(n10343) );
  AND U12671 ( .A(n10344), .B(n10345), .Z(n10342) );
  NANDN U12672 ( .B(n8668), .A(\u_a23_core/u_execute/u_register_bank/r0[26] ), 
        .Z(n10345) );
  NANDN U12673 ( .B(n8671), .A(\u_a23_core/u_execute/u_register_bank/r2[26] ), 
        .Z(n10344) );
  NOR U12674 ( .A(\u_a23_core/execute_address_nxt[24] ), .B(
        \u_a23_core/execute_address_nxt[25] ), .Z(n9981) );
  NAND U12675 ( .A(n10346), .B(n10347), .Z(
        \u_a23_core/execute_address_nxt[25] ) );
  AND U12676 ( .A(n10348), .B(n10349), .Z(n10347) );
  AND U12677 ( .A(n10350), .B(n10351), .Z(n10349) );
  NANDN U12678 ( .B(n8392), .A(\u_a23_core/u_execute/pc_minus4[25] ), .Z(
        n10351) );
  NAND U12679 ( .A(n8393), .B(\u_a23_core/u_execute/alu_out_pc_filtered[25] ), 
        .Z(n10350) );
  IV U12680 ( .A(n7022), .Z(\u_a23_core/u_execute/alu_out_pc_filtered[25] ) );
  AND U12681 ( .A(n10352), .B(n10353), .Z(n7022) );
  MUX U12682 ( .IN0(n10354), .IN1(n10355), .SEL(
        \u_a23_core/u_execute/u_alu/b_not[25] ), .F(n10353) );
  NAND U12683 ( .A(n10356), .B(n10357), .Z(
        \u_a23_core/u_execute/u_alu/b_not[25] ) );
  MUX U12684 ( .IN0(n8430), .IN1(n8431), .SEL(n10358), .F(n10357) );
  MUX U12685 ( .IN0(n8433), .IN1(n8434), .SEL(\u_a23_core/u_execute/rn[25] ), 
        .F(n10356) );
  ANDN U12686 ( .A(n9256), .B(n10359), .Z(n10355) );
  MUX U12687 ( .IN0(n8400), .IN1(\u_a23_core/alu_function[3] ), .SEL(
        \u_a23_core/u_execute/u_alu/a[25] ), .F(n10359) );
  NAND U12688 ( .A(\u_a23_core/u_execute/u_alu/a[25] ), .B(n8400), .Z(n10354)
         );
  IV U12689 ( .A(n10360), .Z(\u_a23_core/u_execute/u_alu/a[25] ) );
  MUX U12690 ( .IN0(n10361), .IN1(n10358), .SEL(\u_a23_core/alu_function[8] ), 
        .F(n10360) );
  AND U12691 ( .A(n10362), .B(n10363), .Z(n10358) );
  AND U12692 ( .A(n10364), .B(n10365), .Z(n10363) );
  NAND U12693 ( .A(n10366), .B(n6888), .Z(n10365) );
  NAND U12694 ( .A(n10367), .B(n10368), .Z(n10366) );
  AND U12695 ( .A(n10369), .B(n10370), .Z(n10368) );
  AND U12696 ( .A(n10371), .B(n10372), .Z(n10370) );
  AND U12697 ( .A(n10373), .B(n10374), .Z(n10372) );
  AND U12698 ( .A(n10375), .B(n10376), .Z(n10374) );
  NANDN U12699 ( .B(n8568), .A(n6919), .Z(n10376) );
  NAND U12700 ( .A(n6827), .B(n8512), .Z(n10375) );
  AND U12701 ( .A(n10377), .B(n10378), .Z(n10373) );
  NANDN U12702 ( .B(n8571), .A(n6920), .Z(n10378) );
  NANDN U12703 ( .B(n8516), .A(n6833), .Z(n10377) );
  AND U12704 ( .A(n10379), .B(n10380), .Z(n10371) );
  AND U12705 ( .A(n10381), .B(n10382), .Z(n10380) );
  NANDN U12706 ( .B(n8572), .A(n6925), .Z(n10382) );
  NANDN U12707 ( .B(n8522), .A(n6835), .Z(n10381) );
  AND U12708 ( .A(n10383), .B(n10384), .Z(n10379) );
  NANDN U12709 ( .B(n8579), .A(n6926), .Z(n10384) );
  NANDN U12710 ( .B(n8526), .A(n6839), .Z(n10383) );
  AND U12711 ( .A(n10385), .B(n10386), .Z(n10369) );
  AND U12712 ( .A(n10387), .B(n10388), .Z(n10386) );
  AND U12713 ( .A(n10389), .B(n10390), .Z(n10388) );
  NANDN U12714 ( .B(n8580), .A(n6898), .Z(n10390) );
  NANDN U12715 ( .B(n8534), .A(n6850), .Z(n10389) );
  AND U12716 ( .A(n10391), .B(n10392), .Z(n10387) );
  NANDN U12717 ( .B(n8511), .A(n6853), .Z(n10392) );
  NANDN U12718 ( .B(n8583), .A(n6882), .Z(n10391) );
  AND U12719 ( .A(n10393), .B(n10394), .Z(n10385) );
  AND U12720 ( .A(n10395), .B(n10396), .Z(n10394) );
  NANDN U12721 ( .B(n8515), .A(n6841), .Z(n10396) );
  NANDN U12722 ( .B(n8584), .A(n6809), .Z(n10395) );
  AND U12723 ( .A(n10397), .B(n10398), .Z(n10393) );
  NANDN U12724 ( .B(n8521), .A(n6857), .Z(n10398) );
  NANDN U12725 ( .B(n8589), .A(n6807), .Z(n10397) );
  AND U12726 ( .A(n10399), .B(n10400), .Z(n10367) );
  AND U12727 ( .A(n10401), .B(n10402), .Z(n10400) );
  AND U12728 ( .A(n10403), .B(n10404), .Z(n10402) );
  AND U12729 ( .A(n10405), .B(n10406), .Z(n10404) );
  NANDN U12730 ( .B(n8525), .A(n6859), .Z(n10406) );
  NANDN U12731 ( .B(n8590), .A(n6799), .Z(n10405) );
  AND U12732 ( .A(n10407), .B(n10408), .Z(n10403) );
  NANDN U12733 ( .B(n8593), .A(n6803), .Z(n10408) );
  NANDN U12734 ( .B(n8533), .A(n6865), .Z(n10407) );
  AND U12735 ( .A(n10409), .B(n10410), .Z(n10401) );
  AND U12736 ( .A(n10411), .B(n10412), .Z(n10410) );
  NAND U12737 ( .A(n6823), .B(n6897), .Z(n10412) );
  NANDN U12738 ( .B(n8537), .A(n6967), .Z(n10411) );
  AND U12739 ( .A(n10413), .B(n10414), .Z(n10409) );
  NANDN U12740 ( .B(n8538), .A(n6966), .Z(n10414) );
  NANDN U12741 ( .B(n8543), .A(n6961), .Z(n10413) );
  AND U12742 ( .A(n10415), .B(n10416), .Z(n10399) );
  AND U12743 ( .A(n10417), .B(n10418), .Z(n10416) );
  AND U12744 ( .A(n10419), .B(n10420), .Z(n10418) );
  NANDN U12745 ( .B(n8544), .A(n6956), .Z(n10420) );
  NANDN U12746 ( .B(n8547), .A(n6960), .Z(n10419) );
  AND U12747 ( .A(n10421), .B(n10422), .Z(n10417) );
  NANDN U12748 ( .B(n8548), .A(n6957), .Z(n10422) );
  NANDN U12749 ( .B(n8557), .A(n6947), .Z(n10421) );
  AND U12750 ( .A(n10423), .B(n10424), .Z(n10415) );
  AND U12751 ( .A(n10425), .B(n10426), .Z(n10424) );
  NANDN U12752 ( .B(n8558), .A(n6946), .Z(n10426) );
  NANDN U12753 ( .B(n8561), .A(n6943), .Z(n10425) );
  AND U12754 ( .A(n10427), .B(n10428), .Z(n10423) );
  NANDN U12755 ( .B(n8562), .A(n6942), .Z(n10428) );
  NANDN U12756 ( .B(n8567), .A(n6937), .Z(n10427) );
  AND U12757 ( .A(n10429), .B(n10430), .Z(n10364) );
  NAND U12758 ( .A(n6886), .B(n10431), .Z(n10430) );
  NAND U12759 ( .A(n10432), .B(n10433), .Z(n10431) );
  AND U12760 ( .A(n10186), .B(n10187), .Z(n10433) );
  IV U12761 ( .A(n8610), .Z(n10186) );
  ANDN U12762 ( .A(n9515), .B(n10188), .Z(n10432) );
  NAND U12763 ( .A(n6786), .B(n10434), .Z(n10429) );
  NAND U12764 ( .A(n10435), .B(n10436), .Z(n10434) );
  AND U12765 ( .A(n10437), .B(n9394), .Z(n10436) );
  NAND U12766 ( .A(n9082), .B(n6799), .Z(n9394) );
  AND U12767 ( .A(n10438), .B(n10439), .Z(n10437) );
  NAND U12768 ( .A(n8616), .B(n6809), .Z(n10439) );
  NAND U12769 ( .A(n8958), .B(n6807), .Z(n10438) );
  AND U12770 ( .A(n10440), .B(n10441), .Z(n10435) );
  NAND U12771 ( .A(n6893), .B(n6827), .Z(n10441) );
  AND U12772 ( .A(n10125), .B(n9759), .Z(n10440) );
  NAND U12773 ( .A(n9135), .B(n6803), .Z(n9759) );
  NAND U12774 ( .A(n6984), .B(n6823), .Z(n10125) );
  AND U12775 ( .A(n10442), .B(n10443), .Z(n10362) );
  NAND U12776 ( .A(n10444), .B(n6902), .Z(n10443) );
  NAND U12777 ( .A(n10445), .B(n10446), .Z(n10444) );
  AND U12778 ( .A(n10447), .B(n10448), .Z(n10446) );
  AND U12779 ( .A(n10449), .B(n10450), .Z(n10448) );
  AND U12780 ( .A(n10451), .B(n10452), .Z(n10450) );
  ANDN U12781 ( .A(n10453), .B(n10454), .Z(n10452) );
  NAND U12782 ( .A(n6916), .B(n6827), .Z(n10453) );
  AND U12783 ( .A(n10455), .B(n10456), .Z(n10451) );
  NAND U12784 ( .A(n8464), .B(n6957), .Z(n10456) );
  NAND U12785 ( .A(n8465), .B(n6960), .Z(n10455) );
  AND U12786 ( .A(n10457), .B(n10458), .Z(n10449) );
  AND U12787 ( .A(n10459), .B(n6815), .Z(n10457) );
  NAND U12788 ( .A(n8461), .B(n6956), .Z(n6815) );
  AND U12789 ( .A(n10460), .B(n10461), .Z(n10447) );
  AND U12790 ( .A(n10462), .B(n10463), .Z(n10461) );
  NAND U12791 ( .A(n6834), .B(n6926), .Z(n10463) );
  AND U12792 ( .A(n10464), .B(n9098), .Z(n10462) );
  NAND U12793 ( .A(n6967), .B(n9726), .Z(n9098) );
  NAND U12794 ( .A(n6832), .B(n6898), .Z(n10464) );
  AND U12795 ( .A(n10465), .B(n10466), .Z(n10460) );
  NAND U12796 ( .A(n6920), .B(n6851), .Z(n10466) );
  AND U12797 ( .A(n10467), .B(n10468), .Z(n10465) );
  NAND U12798 ( .A(n6838), .B(n6925), .Z(n10468) );
  NAND U12799 ( .A(n6840), .B(n6937), .Z(n10467) );
  AND U12800 ( .A(n10469), .B(n10470), .Z(n10445) );
  AND U12801 ( .A(n10471), .B(n10472), .Z(n10470) );
  AND U12802 ( .A(n10473), .B(n10474), .Z(n10472) );
  AND U12803 ( .A(n10475), .B(n10476), .Z(n10474) );
  NAND U12804 ( .A(n6852), .B(n6919), .Z(n10476) );
  NAND U12805 ( .A(n6856), .B(n6942), .Z(n10475) );
  AND U12806 ( .A(n10477), .B(n10478), .Z(n10473) );
  NAND U12807 ( .A(n6858), .B(n6943), .Z(n10478) );
  NAND U12808 ( .A(n6864), .B(n6946), .Z(n10477) );
  AND U12809 ( .A(n10479), .B(n8491), .Z(n10471) );
  NAND U12810 ( .A(n8609), .B(n6859), .Z(n8491) );
  AND U12811 ( .A(n10480), .B(n10481), .Z(n10479) );
  NAND U12812 ( .A(n6947), .B(n8487), .Z(n10481) );
  AND U12813 ( .A(n10482), .B(n10483), .Z(n10469) );
  AND U12814 ( .A(n10484), .B(n10485), .Z(n10483) );
  AND U12815 ( .A(n10486), .B(n10487), .Z(n10484) );
  AND U12816 ( .A(n10488), .B(n10489), .Z(n10482) );
  AND U12817 ( .A(n10490), .B(n10491), .Z(n10488) );
  NAND U12818 ( .A(n8610), .B(n6985), .Z(n10442) );
  IV U12819 ( .A(\u_a23_core/u_execute/rn[25] ), .Z(n10361) );
  AND U12820 ( .A(n9395), .B(n10492), .Z(n10352) );
  NAND U12821 ( .A(n6765), .B(\u_a23_core/u_execute/u_alu/fadder_out[25] ), 
        .Z(n10492) );
  AND U12822 ( .A(n10493), .B(n10494), .Z(n10348) );
  NANDN U12823 ( .B(n8406), .A(\u_a23_core/u_execute/rn_plus4[25] ), .Z(n10494) );
  NANDN U12824 ( .B(n8407), .A(\u_a23_core/u_execute/alu_plus4[25] ), .Z(
        n10493) );
  AND U12825 ( .A(n10495), .B(n10496), .Z(n10346) );
  AND U12826 ( .A(n10497), .B(n10498), .Z(n10496) );
  NAND U12827 ( .A(n8412), .B(\u_a23_core/u_execute/address_plus4[25] ), .Z(
        n10498) );
  NAND U12828 ( .A(\u_a23_core/u_execute/rn[25] ), .B(n8413), .Z(n10497) );
  NAND U12829 ( .A(n10499), .B(n10500), .Z(\u_a23_core/u_execute/rn[25] ) );
  AND U12830 ( .A(n10501), .B(n10502), .Z(n10500) );
  AND U12831 ( .A(n10503), .B(n10504), .Z(n10502) );
  AND U12832 ( .A(n10505), .B(n10506), .Z(n10504) );
  NANDN U12833 ( .B(n8635), .A(\u_a23_core/u_execute/pc[25] ), .Z(n10506) );
  NANDN U12834 ( .B(n8636), .A(\u_a23_core/u_execute/u_register_bank/r14[25] ), 
        .Z(n10505) );
  AND U12835 ( .A(n10507), .B(n10508), .Z(n10503) );
  NANDN U12836 ( .B(n8639), .A(\u_a23_core/u_execute/u_register_bank/r13[25] ), 
        .Z(n10508) );
  NANDN U12837 ( .B(n8640), .A(\u_a23_core/u_execute/u_register_bank/r12[25] ), 
        .Z(n10507) );
  AND U12838 ( .A(n10509), .B(n10510), .Z(n10501) );
  AND U12839 ( .A(n10511), .B(n10512), .Z(n10510) );
  NANDN U12840 ( .B(n8645), .A(\u_a23_core/u_execute/u_register_bank/r11[25] ), 
        .Z(n10512) );
  NANDN U12841 ( .B(n8646), .A(\u_a23_core/u_execute/u_register_bank/r10[25] ), 
        .Z(n10511) );
  AND U12842 ( .A(n10513), .B(n10514), .Z(n10509) );
  NANDN U12843 ( .B(n8649), .A(\u_a23_core/u_execute/u_register_bank/r9[25] ), 
        .Z(n10514) );
  NANDN U12844 ( .B(n8650), .A(\u_a23_core/u_execute/u_register_bank/r8[25] ), 
        .Z(n10513) );
  AND U12845 ( .A(n10515), .B(n10516), .Z(n10499) );
  AND U12846 ( .A(n10517), .B(n10518), .Z(n10516) );
  AND U12847 ( .A(n10519), .B(n10520), .Z(n10518) );
  NANDN U12848 ( .B(n8657), .A(\u_a23_core/u_execute/u_register_bank/r7[25] ), 
        .Z(n10520) );
  NANDN U12849 ( .B(n8658), .A(\u_a23_core/u_execute/u_register_bank/r6[25] ), 
        .Z(n10519) );
  AND U12850 ( .A(n10521), .B(n10522), .Z(n10517) );
  NANDN U12851 ( .B(n8661), .A(\u_a23_core/u_execute/u_register_bank/r5[25] ), 
        .Z(n10522) );
  NANDN U12852 ( .B(n8662), .A(\u_a23_core/u_execute/u_register_bank/r4[25] ), 
        .Z(n10521) );
  AND U12853 ( .A(n10523), .B(n10524), .Z(n10515) );
  AND U12854 ( .A(n10525), .B(n10526), .Z(n10524) );
  NANDN U12855 ( .B(n8667), .A(\u_a23_core/u_execute/u_register_bank/r3[25] ), 
        .Z(n10526) );
  NANDN U12856 ( .B(n8668), .A(\u_a23_core/u_execute/u_register_bank/r0[25] ), 
        .Z(n10525) );
  AND U12857 ( .A(n10527), .B(n10528), .Z(n10523) );
  NANDN U12858 ( .B(n8671), .A(\u_a23_core/u_execute/u_register_bank/r2[25] ), 
        .Z(n10528) );
  NANDN U12859 ( .B(n8672), .A(\u_a23_core/u_execute/u_register_bank/r1[25] ), 
        .Z(n10527) );
  AND U12860 ( .A(n10529), .B(n10530), .Z(n10495) );
  NAND U12861 ( .A(\u_a23_core/u_execute/pc[25] ), .B(n8416), .Z(n10530) );
  NAND U12862 ( .A(n8417), .B(\u_a23_core/u_execute/pc_plus4[25] ), .Z(n10529)
         );
  NAND U12863 ( .A(n10531), .B(n10532), .Z(
        \u_a23_core/execute_address_nxt[24] ) );
  AND U12864 ( .A(n10533), .B(n10534), .Z(n10532) );
  AND U12865 ( .A(n10535), .B(n10536), .Z(n10534) );
  NANDN U12866 ( .B(n8392), .A(\u_a23_core/u_execute/pc_minus4[24] ), .Z(
        n10536) );
  NAND U12867 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[24] ), .B(n8393), 
        .Z(n10535) );
  IV U12868 ( .A(n7023), .Z(\u_a23_core/u_execute/alu_out_pc_filtered[24] ) );
  AND U12869 ( .A(n10537), .B(n10538), .Z(n7023) );
  MUX U12870 ( .IN0(n10539), .IN1(n10540), .SEL(
        \u_a23_core/u_execute/u_alu/b_not[24] ), .F(n10538) );
  NAND U12871 ( .A(n10541), .B(n10542), .Z(
        \u_a23_core/u_execute/u_alu/b_not[24] ) );
  MUX U12872 ( .IN0(n8430), .IN1(n8431), .SEL(n10543), .F(n10542) );
  MUX U12873 ( .IN0(n8433), .IN1(n8434), .SEL(\u_a23_core/u_execute/rn[24] ), 
        .F(n10541) );
  ANDN U12874 ( .A(n9256), .B(n10544), .Z(n10540) );
  MUX U12875 ( .IN0(n8400), .IN1(\u_a23_core/alu_function[3] ), .SEL(
        \u_a23_core/u_execute/u_alu/a[24] ), .F(n10544) );
  NAND U12876 ( .A(\u_a23_core/u_execute/u_alu/a[24] ), .B(n8400), .Z(n10539)
         );
  IV U12877 ( .A(n10545), .Z(\u_a23_core/u_execute/u_alu/a[24] ) );
  MUX U12878 ( .IN0(n10546), .IN1(n10543), .SEL(\u_a23_core/alu_function[8] ), 
        .F(n10545) );
  AND U12879 ( .A(n10547), .B(n10548), .Z(n10543) );
  AND U12880 ( .A(n10549), .B(n10550), .Z(n10548) );
  NAND U12881 ( .A(n10551), .B(n10552), .Z(n10550) );
  NAND U12882 ( .A(n10187), .B(n10553), .Z(n10551) );
  NAND U12883 ( .A(n8443), .B(n10554), .Z(n10553) );
  IV U12884 ( .A(n8606), .Z(n10187) );
  NAND U12885 ( .A(n6786), .B(n10555), .Z(n10549) );
  NAND U12886 ( .A(n10556), .B(n10557), .Z(n10555) );
  AND U12887 ( .A(n10558), .B(n10559), .Z(n10557) );
  AND U12888 ( .A(n10560), .B(n10561), .Z(n10559) );
  NAND U12889 ( .A(n8610), .B(n6809), .Z(n10561) );
  NAND U12890 ( .A(n8616), .B(n6807), .Z(n10560) );
  AND U12891 ( .A(n9506), .B(n6981), .Z(n10558) );
  NAND U12892 ( .A(n8958), .B(n6799), .Z(n6981) );
  NAND U12893 ( .A(n9082), .B(n6803), .Z(n9506) );
  AND U12894 ( .A(n10562), .B(n10563), .Z(n10556) );
  NAND U12895 ( .A(n6893), .B(n6833), .Z(n10563) );
  AND U12896 ( .A(n10308), .B(n9944), .Z(n10562) );
  NAND U12897 ( .A(n9135), .B(n6823), .Z(n9944) );
  NAND U12898 ( .A(n6984), .B(n6827), .Z(n10308) );
  AND U12899 ( .A(n10564), .B(n10565), .Z(n10547) );
  NAND U12900 ( .A(n10566), .B(n6888), .Z(n10565) );
  NAND U12901 ( .A(n10567), .B(n10568), .Z(n10566) );
  AND U12902 ( .A(n10569), .B(n10570), .Z(n10568) );
  AND U12903 ( .A(n10571), .B(n10572), .Z(n10570) );
  AND U12904 ( .A(n10573), .B(n10574), .Z(n10572) );
  AND U12905 ( .A(n10575), .B(n10576), .Z(n10574) );
  NANDN U12906 ( .B(n8567), .A(n6919), .Z(n10576) );
  NAND U12907 ( .A(n6833), .B(n8512), .Z(n10575) );
  AND U12908 ( .A(n10577), .B(n10578), .Z(n10573) );
  NANDN U12909 ( .B(n8568), .A(n6920), .Z(n10578) );
  NANDN U12910 ( .B(n8516), .A(n6835), .Z(n10577) );
  AND U12911 ( .A(n10579), .B(n10580), .Z(n10571) );
  AND U12912 ( .A(n10581), .B(n10582), .Z(n10580) );
  NANDN U12913 ( .B(n8571), .A(n6925), .Z(n10582) );
  NANDN U12914 ( .B(n8522), .A(n6839), .Z(n10581) );
  AND U12915 ( .A(n10583), .B(n10584), .Z(n10579) );
  NANDN U12916 ( .B(n8572), .A(n6926), .Z(n10584) );
  NANDN U12917 ( .B(n8526), .A(n6850), .Z(n10583) );
  AND U12918 ( .A(n10585), .B(n10586), .Z(n10569) );
  AND U12919 ( .A(n10587), .B(n10588), .Z(n10586) );
  AND U12920 ( .A(n10589), .B(n10590), .Z(n10588) );
  NANDN U12921 ( .B(n8579), .A(n6898), .Z(n10590) );
  NANDN U12922 ( .B(n8534), .A(n6853), .Z(n10589) );
  AND U12923 ( .A(n10591), .B(n10592), .Z(n10587) );
  NANDN U12924 ( .B(n8511), .A(n6841), .Z(n10592) );
  NANDN U12925 ( .B(n8580), .A(n6882), .Z(n10591) );
  AND U12926 ( .A(n10593), .B(n10594), .Z(n10585) );
  AND U12927 ( .A(n10595), .B(n10596), .Z(n10594) );
  NANDN U12928 ( .B(n8515), .A(n6857), .Z(n10596) );
  NANDN U12929 ( .B(n8583), .A(n6809), .Z(n10595) );
  AND U12930 ( .A(n10597), .B(n10598), .Z(n10593) );
  NANDN U12931 ( .B(n8521), .A(n6859), .Z(n10598) );
  NANDN U12932 ( .B(n8584), .A(n6807), .Z(n10597) );
  AND U12933 ( .A(n10599), .B(n10600), .Z(n10567) );
  AND U12934 ( .A(n10601), .B(n10602), .Z(n10600) );
  AND U12935 ( .A(n10603), .B(n10604), .Z(n10602) );
  AND U12936 ( .A(n10605), .B(n10606), .Z(n10604) );
  NANDN U12937 ( .B(n8525), .A(n6865), .Z(n10606) );
  NANDN U12938 ( .B(n8589), .A(n6799), .Z(n10605) );
  AND U12939 ( .A(n10607), .B(n10608), .Z(n10603) );
  NANDN U12940 ( .B(n8590), .A(n6803), .Z(n10608) );
  NANDN U12941 ( .B(n8533), .A(n6967), .Z(n10607) );
  AND U12942 ( .A(n10609), .B(n10610), .Z(n10601) );
  AND U12943 ( .A(n10611), .B(n10612), .Z(n10610) );
  NANDN U12944 ( .B(n8593), .A(n6823), .Z(n10612) );
  NANDN U12945 ( .B(n8537), .A(n6966), .Z(n10611) );
  AND U12946 ( .A(n10613), .B(n10614), .Z(n10609) );
  NAND U12947 ( .A(n6827), .B(n6897), .Z(n10614) );
  NANDN U12948 ( .B(n8538), .A(n6961), .Z(n10613) );
  AND U12949 ( .A(n10615), .B(n10616), .Z(n10599) );
  AND U12950 ( .A(n10617), .B(n10618), .Z(n10616) );
  AND U12951 ( .A(n10619), .B(n10620), .Z(n10618) );
  NANDN U12952 ( .B(n8543), .A(n6956), .Z(n10620) );
  NANDN U12953 ( .B(n8544), .A(n6960), .Z(n10619) );
  AND U12954 ( .A(n10621), .B(n10622), .Z(n10617) );
  NANDN U12955 ( .B(n8547), .A(n6957), .Z(n10622) );
  NANDN U12956 ( .B(n8548), .A(n6947), .Z(n10621) );
  AND U12957 ( .A(n10623), .B(n10624), .Z(n10615) );
  AND U12958 ( .A(n10625), .B(n10626), .Z(n10624) );
  NANDN U12959 ( .B(n8557), .A(n6946), .Z(n10626) );
  NANDN U12960 ( .B(n8558), .A(n6943), .Z(n10625) );
  AND U12961 ( .A(n10627), .B(n10628), .Z(n10623) );
  NANDN U12962 ( .B(n8561), .A(n6942), .Z(n10628) );
  NANDN U12963 ( .B(n8562), .A(n6937), .Z(n10627) );
  NAND U12964 ( .A(n10629), .B(n6902), .Z(n10564) );
  NAND U12965 ( .A(n10630), .B(n10631), .Z(n10629) );
  AND U12966 ( .A(n10632), .B(n10633), .Z(n10631) );
  AND U12967 ( .A(n10634), .B(n10635), .Z(n10633) );
  AND U12968 ( .A(n10636), .B(n10637), .Z(n10635) );
  NOR U12969 ( .A(n8707), .B(n8974), .Z(n10637) );
  ANDN U12970 ( .A(n8603), .B(n10638), .Z(n8974) );
  ANDN U12971 ( .A(n8609), .B(n10639), .Z(n8707) );
  AND U12972 ( .A(n10640), .B(n10641), .Z(n10636) );
  NAND U12973 ( .A(n6916), .B(n6833), .Z(n10641) );
  NAND U12974 ( .A(n8464), .B(n6947), .Z(n10640) );
  AND U12975 ( .A(n10642), .B(n10643), .Z(n10634) );
  AND U12976 ( .A(n10644), .B(n10645), .Z(n10642) );
  NAND U12977 ( .A(n8465), .B(n6957), .Z(n10645) );
  NAND U12978 ( .A(n8461), .B(n6960), .Z(n10644) );
  AND U12979 ( .A(n10646), .B(n10647), .Z(n10632) );
  AND U12980 ( .A(n10648), .B(n10649), .Z(n10647) );
  NAND U12981 ( .A(n6834), .B(n6898), .Z(n10649) );
  AND U12982 ( .A(n10650), .B(n10651), .Z(n10648) );
  AND U12983 ( .A(n10652), .B(n10653), .Z(n10646) );
  NAND U12984 ( .A(n6925), .B(n6851), .Z(n10653) );
  AND U12985 ( .A(n10654), .B(n10655), .Z(n10652) );
  NAND U12986 ( .A(n6838), .B(n6926), .Z(n10655) );
  NAND U12987 ( .A(n6840), .B(n6919), .Z(n10654) );
  AND U12988 ( .A(n10656), .B(n10657), .Z(n10630) );
  AND U12989 ( .A(n10658), .B(n10659), .Z(n10657) );
  AND U12990 ( .A(n10660), .B(n10661), .Z(n10659) );
  NAND U12991 ( .A(n6858), .B(n6942), .Z(n10661) );
  AND U12992 ( .A(n10662), .B(n10663), .Z(n10660) );
  NAND U12993 ( .A(n6852), .B(n6920), .Z(n10663) );
  NAND U12994 ( .A(n6856), .B(n6937), .Z(n10662) );
  AND U12995 ( .A(n10664), .B(n10665), .Z(n10658) );
  AND U12996 ( .A(n10666), .B(n10667), .Z(n10664) );
  NAND U12997 ( .A(n6864), .B(n6943), .Z(n10667) );
  NAND U12998 ( .A(n6946), .B(n8487), .Z(n10666) );
  AND U12999 ( .A(n10668), .B(n10669), .Z(n10656) );
  AND U13000 ( .A(n10670), .B(n10671), .Z(n10669) );
  AND U13001 ( .A(n10672), .B(n10673), .Z(n10670) );
  AND U13002 ( .A(n10674), .B(n10675), .Z(n10668) );
  AND U13003 ( .A(n10676), .B(n10677), .Z(n10674) );
  IV U13004 ( .A(\u_a23_core/u_execute/rn[24] ), .Z(n10546) );
  AND U13005 ( .A(n9395), .B(n10678), .Z(n10537) );
  NAND U13006 ( .A(n6765), .B(\u_a23_core/u_execute/u_alu/fadder_out[24] ), 
        .Z(n10678) );
  AND U13007 ( .A(n10679), .B(n10680), .Z(n10533) );
  NANDN U13008 ( .B(n8406), .A(\u_a23_core/u_execute/rn_plus4[24] ), .Z(n10680) );
  NANDN U13009 ( .B(n8407), .A(\u_a23_core/u_execute/alu_plus4[24] ), .Z(
        n10679) );
  AND U13010 ( .A(n10681), .B(n10682), .Z(n10531) );
  AND U13011 ( .A(n10683), .B(n10684), .Z(n10682) );
  NAND U13012 ( .A(n8412), .B(\u_a23_core/u_execute/address_plus4[24] ), .Z(
        n10684) );
  NAND U13013 ( .A(\u_a23_core/u_execute/rn[24] ), .B(n8413), .Z(n10683) );
  NAND U13014 ( .A(n10685), .B(n10686), .Z(\u_a23_core/u_execute/rn[24] ) );
  AND U13015 ( .A(n10687), .B(n10688), .Z(n10686) );
  AND U13016 ( .A(n10689), .B(n10690), .Z(n10688) );
  AND U13017 ( .A(n10691), .B(n10692), .Z(n10690) );
  NANDN U13018 ( .B(n8635), .A(\u_a23_core/u_execute/pc[24] ), .Z(n10692) );
  NANDN U13019 ( .B(n8636), .A(\u_a23_core/u_execute/u_register_bank/r14[24] ), 
        .Z(n10691) );
  AND U13020 ( .A(n10693), .B(n10694), .Z(n10689) );
  NANDN U13021 ( .B(n8639), .A(\u_a23_core/u_execute/u_register_bank/r13[24] ), 
        .Z(n10694) );
  NANDN U13022 ( .B(n8640), .A(\u_a23_core/u_execute/u_register_bank/r12[24] ), 
        .Z(n10693) );
  AND U13023 ( .A(n10695), .B(n10696), .Z(n10687) );
  AND U13024 ( .A(n10697), .B(n10698), .Z(n10696) );
  NANDN U13025 ( .B(n8645), .A(\u_a23_core/u_execute/u_register_bank/r11[24] ), 
        .Z(n10698) );
  NANDN U13026 ( .B(n8646), .A(\u_a23_core/u_execute/u_register_bank/r10[24] ), 
        .Z(n10697) );
  AND U13027 ( .A(n10699), .B(n10700), .Z(n10695) );
  NANDN U13028 ( .B(n8649), .A(\u_a23_core/u_execute/u_register_bank/r9[24] ), 
        .Z(n10700) );
  NANDN U13029 ( .B(n8650), .A(\u_a23_core/u_execute/u_register_bank/r8[24] ), 
        .Z(n10699) );
  AND U13030 ( .A(n10701), .B(n10702), .Z(n10685) );
  AND U13031 ( .A(n10703), .B(n10704), .Z(n10702) );
  AND U13032 ( .A(n10705), .B(n10706), .Z(n10704) );
  NANDN U13033 ( .B(n8657), .A(\u_a23_core/u_execute/u_register_bank/r7[24] ), 
        .Z(n10706) );
  NANDN U13034 ( .B(n8658), .A(\u_a23_core/u_execute/u_register_bank/r6[24] ), 
        .Z(n10705) );
  AND U13035 ( .A(n10707), .B(n10708), .Z(n10703) );
  NANDN U13036 ( .B(n8661), .A(\u_a23_core/u_execute/u_register_bank/r5[24] ), 
        .Z(n10708) );
  NANDN U13037 ( .B(n8662), .A(\u_a23_core/u_execute/u_register_bank/r4[24] ), 
        .Z(n10707) );
  AND U13038 ( .A(n10709), .B(n10710), .Z(n10701) );
  AND U13039 ( .A(n10711), .B(n10712), .Z(n10710) );
  NANDN U13040 ( .B(n8667), .A(\u_a23_core/u_execute/u_register_bank/r3[24] ), 
        .Z(n10712) );
  NANDN U13041 ( .B(n8668), .A(\u_a23_core/u_execute/u_register_bank/r0[24] ), 
        .Z(n10711) );
  AND U13042 ( .A(n10713), .B(n10714), .Z(n10709) );
  NANDN U13043 ( .B(n8671), .A(\u_a23_core/u_execute/u_register_bank/r2[24] ), 
        .Z(n10714) );
  NANDN U13044 ( .B(n8672), .A(\u_a23_core/u_execute/u_register_bank/r1[24] ), 
        .Z(n10713) );
  AND U13045 ( .A(n10715), .B(n10716), .Z(n10681) );
  NAND U13046 ( .A(\u_a23_core/u_execute/pc[24] ), .B(n8416), .Z(n10716) );
  NAND U13047 ( .A(n8417), .B(\u_a23_core/u_execute/pc_plus4[24] ), .Z(n10715)
         );
  AND U13048 ( .A(n10717), .B(n10718), .Z(n9979) );
  NOR U13049 ( .A(\u_a23_core/execute_address_nxt[22] ), .B(
        \u_a23_core/execute_address_nxt[23] ), .Z(n10718) );
  NAND U13050 ( .A(n10719), .B(n10720), .Z(
        \u_a23_core/execute_address_nxt[23] ) );
  AND U13051 ( .A(n10721), .B(n10722), .Z(n10720) );
  AND U13052 ( .A(n10723), .B(n10724), .Z(n10722) );
  NANDN U13053 ( .B(n8392), .A(\u_a23_core/u_execute/pc_minus4[23] ), .Z(
        n10724) );
  NAND U13054 ( .A(n8393), .B(\u_a23_core/u_execute/alu_out_pc_filtered[23] ), 
        .Z(n10723) );
  IV U13055 ( .A(n7024), .Z(\u_a23_core/u_execute/alu_out_pc_filtered[23] ) );
  AND U13056 ( .A(n10725), .B(n10726), .Z(n7024) );
  MUX U13057 ( .IN0(n10727), .IN1(n10728), .SEL(
        \u_a23_core/u_execute/u_alu/b_not[23] ), .F(n10726) );
  NAND U13058 ( .A(n10729), .B(n10730), .Z(
        \u_a23_core/u_execute/u_alu/b_not[23] ) );
  MUX U13059 ( .IN0(n8430), .IN1(n8431), .SEL(n10731), .F(n10730) );
  MUX U13060 ( .IN0(n8433), .IN1(n8434), .SEL(\u_a23_core/u_execute/rn[23] ), 
        .F(n10729) );
  ANDN U13061 ( .A(n9256), .B(n10732), .Z(n10728) );
  MUX U13062 ( .IN0(n8400), .IN1(\u_a23_core/alu_function[3] ), .SEL(
        \u_a23_core/u_execute/u_alu/a[23] ), .F(n10732) );
  NAND U13063 ( .A(\u_a23_core/u_execute/u_alu/a[23] ), .B(n8400), .Z(n10727)
         );
  IV U13064 ( .A(n10733), .Z(\u_a23_core/u_execute/u_alu/a[23] ) );
  MUX U13065 ( .IN0(n10734), .IN1(n10731), .SEL(\u_a23_core/alu_function[8] ), 
        .F(n10733) );
  AND U13066 ( .A(n10735), .B(n10736), .Z(n10731) );
  AND U13067 ( .A(n10737), .B(n10738), .Z(n10736) );
  NAND U13068 ( .A(n10739), .B(n10552), .Z(n10738) );
  AND U13069 ( .A(n10554), .B(n10740), .Z(n10739) );
  NAND U13070 ( .A(n10741), .B(n10742), .Z(n10740) );
  IV U13071 ( .A(n8443), .Z(n10742) );
  NAND U13072 ( .A(n9885), .B(n10743), .Z(n10554) );
  ANDN U13073 ( .A(n9884), .B(n10188), .Z(n10743) );
  NAND U13074 ( .A(n10744), .B(n10745), .Z(n10188) );
  AND U13075 ( .A(n10741), .B(n10746), .Z(n10745) );
  IV U13076 ( .A(n8609), .Z(n10741) );
  NAND U13077 ( .A(n6786), .B(n10747), .Z(n10737) );
  NAND U13078 ( .A(n10748), .B(n10749), .Z(n10747) );
  AND U13079 ( .A(n10750), .B(n10751), .Z(n10749) );
  AND U13080 ( .A(n10752), .B(n10753), .Z(n10751) );
  NAND U13081 ( .A(n8606), .B(n6809), .Z(n10753) );
  NAND U13082 ( .A(n8610), .B(n6807), .Z(n10752) );
  AND U13083 ( .A(n9391), .B(n10754), .Z(n10750) );
  NAND U13084 ( .A(n8616), .B(n6799), .Z(n10754) );
  NAND U13085 ( .A(n8958), .B(n6803), .Z(n9391) );
  AND U13086 ( .A(n10755), .B(n10756), .Z(n10748) );
  AND U13087 ( .A(n10126), .B(n9760), .Z(n10756) );
  NAND U13088 ( .A(n9082), .B(n6823), .Z(n9760) );
  NAND U13089 ( .A(n9135), .B(n6827), .Z(n10126) );
  AND U13090 ( .A(n10757), .B(n10489), .Z(n10755) );
  NAND U13091 ( .A(n6984), .B(n6833), .Z(n10489) );
  NAND U13092 ( .A(n6893), .B(n6835), .Z(n10757) );
  AND U13093 ( .A(n10758), .B(n10759), .Z(n10735) );
  NAND U13094 ( .A(n10760), .B(n6888), .Z(n10759) );
  NAND U13095 ( .A(n10761), .B(n10762), .Z(n10760) );
  AND U13096 ( .A(n10763), .B(n10764), .Z(n10762) );
  AND U13097 ( .A(n10765), .B(n10766), .Z(n10764) );
  AND U13098 ( .A(n10767), .B(n10768), .Z(n10766) );
  AND U13099 ( .A(n10769), .B(n10770), .Z(n10768) );
  NANDN U13100 ( .B(n8562), .A(n6919), .Z(n10770) );
  NAND U13101 ( .A(n6835), .B(n8512), .Z(n10769) );
  AND U13102 ( .A(n10771), .B(n10772), .Z(n10767) );
  NANDN U13103 ( .B(n8567), .A(n6920), .Z(n10772) );
  NANDN U13104 ( .B(n8516), .A(n6839), .Z(n10771) );
  AND U13105 ( .A(n10773), .B(n10774), .Z(n10765) );
  AND U13106 ( .A(n10775), .B(n10776), .Z(n10774) );
  NANDN U13107 ( .B(n8568), .A(n6925), .Z(n10776) );
  NANDN U13108 ( .B(n8522), .A(n6850), .Z(n10775) );
  AND U13109 ( .A(n10777), .B(n10778), .Z(n10773) );
  NANDN U13110 ( .B(n8571), .A(n6926), .Z(n10778) );
  NANDN U13111 ( .B(n8526), .A(n6853), .Z(n10777) );
  AND U13112 ( .A(n10779), .B(n10780), .Z(n10763) );
  AND U13113 ( .A(n10781), .B(n10782), .Z(n10780) );
  AND U13114 ( .A(n10783), .B(n10784), .Z(n10782) );
  NANDN U13115 ( .B(n8572), .A(n6898), .Z(n10784) );
  NANDN U13116 ( .B(n8534), .A(n6841), .Z(n10783) );
  AND U13117 ( .A(n10785), .B(n10786), .Z(n10781) );
  NANDN U13118 ( .B(n8511), .A(n6857), .Z(n10786) );
  NANDN U13119 ( .B(n8579), .A(n6882), .Z(n10785) );
  AND U13120 ( .A(n10787), .B(n10788), .Z(n10779) );
  AND U13121 ( .A(n10789), .B(n10790), .Z(n10788) );
  NANDN U13122 ( .B(n8515), .A(n6859), .Z(n10790) );
  NANDN U13123 ( .B(n8580), .A(n6809), .Z(n10789) );
  AND U13124 ( .A(n10791), .B(n10792), .Z(n10787) );
  NANDN U13125 ( .B(n8521), .A(n6865), .Z(n10792) );
  NANDN U13126 ( .B(n8583), .A(n6807), .Z(n10791) );
  AND U13127 ( .A(n10793), .B(n10794), .Z(n10761) );
  AND U13128 ( .A(n10795), .B(n10796), .Z(n10794) );
  AND U13129 ( .A(n10797), .B(n10798), .Z(n10796) );
  AND U13130 ( .A(n10799), .B(n10800), .Z(n10798) );
  NANDN U13131 ( .B(n8525), .A(n6967), .Z(n10800) );
  NANDN U13132 ( .B(n8584), .A(n6799), .Z(n10799) );
  AND U13133 ( .A(n10801), .B(n10802), .Z(n10797) );
  NANDN U13134 ( .B(n8589), .A(n6803), .Z(n10802) );
  NANDN U13135 ( .B(n8533), .A(n6966), .Z(n10801) );
  AND U13136 ( .A(n10803), .B(n10804), .Z(n10795) );
  AND U13137 ( .A(n10805), .B(n10806), .Z(n10804) );
  NANDN U13138 ( .B(n8590), .A(n6823), .Z(n10806) );
  NANDN U13139 ( .B(n8537), .A(n6961), .Z(n10805) );
  AND U13140 ( .A(n10807), .B(n10808), .Z(n10803) );
  NANDN U13141 ( .B(n8593), .A(n6827), .Z(n10808) );
  NANDN U13142 ( .B(n8538), .A(n6956), .Z(n10807) );
  AND U13143 ( .A(n10809), .B(n10810), .Z(n10793) );
  AND U13144 ( .A(n10811), .B(n10812), .Z(n10810) );
  AND U13145 ( .A(n10813), .B(n10814), .Z(n10812) );
  NAND U13146 ( .A(n6833), .B(n6897), .Z(n10814) );
  NANDN U13147 ( .B(n8543), .A(n6960), .Z(n10813) );
  AND U13148 ( .A(n10815), .B(n10816), .Z(n10811) );
  NANDN U13149 ( .B(n8544), .A(n6957), .Z(n10816) );
  NANDN U13150 ( .B(n8547), .A(n6947), .Z(n10815) );
  AND U13151 ( .A(n10817), .B(n10818), .Z(n10809) );
  AND U13152 ( .A(n10819), .B(n10820), .Z(n10818) );
  NANDN U13153 ( .B(n8548), .A(n6946), .Z(n10820) );
  NANDN U13154 ( .B(n8557), .A(n6943), .Z(n10819) );
  AND U13155 ( .A(n10821), .B(n10822), .Z(n10817) );
  NANDN U13156 ( .B(n8558), .A(n6942), .Z(n10822) );
  NANDN U13157 ( .B(n8561), .A(n6937), .Z(n10821) );
  NAND U13158 ( .A(n10823), .B(n6902), .Z(n10758) );
  NAND U13159 ( .A(n10824), .B(n10825), .Z(n10823) );
  AND U13160 ( .A(n10826), .B(n10827), .Z(n10825) );
  AND U13161 ( .A(n10828), .B(n10829), .Z(n10827) );
  AND U13162 ( .A(n10830), .B(n10831), .Z(n10829) );
  NAND U13163 ( .A(n8464), .B(n6946), .Z(n10831) );
  AND U13164 ( .A(n10832), .B(n10833), .Z(n10830) );
  NAND U13165 ( .A(n6916), .B(n6835), .Z(n10833) );
  AND U13166 ( .A(n10834), .B(n6814), .Z(n10828) );
  NAND U13167 ( .A(n8470), .B(n6960), .Z(n6814) );
  AND U13168 ( .A(n10835), .B(n10836), .Z(n10834) );
  NAND U13169 ( .A(n8465), .B(n6947), .Z(n10836) );
  NAND U13170 ( .A(n8461), .B(n6957), .Z(n10835) );
  AND U13171 ( .A(n10837), .B(n10838), .Z(n10826) );
  AND U13172 ( .A(n10839), .B(n10840), .Z(n10838) );
  NAND U13173 ( .A(n6838), .B(n6898), .Z(n10840) );
  AND U13174 ( .A(n10841), .B(n10842), .Z(n10839) );
  AND U13175 ( .A(n10843), .B(n10844), .Z(n10837) );
  NAND U13176 ( .A(n6852), .B(n6925), .Z(n10844) );
  AND U13177 ( .A(n10845), .B(n10846), .Z(n10843) );
  NAND U13178 ( .A(n6840), .B(n6920), .Z(n10846) );
  NAND U13179 ( .A(n6926), .B(n6851), .Z(n10845) );
  AND U13180 ( .A(n10847), .B(n10848), .Z(n10824) );
  AND U13181 ( .A(n10849), .B(n10850), .Z(n10848) );
  AND U13182 ( .A(n10851), .B(n10852), .Z(n10850) );
  NAND U13183 ( .A(n6864), .B(n6942), .Z(n10852) );
  AND U13184 ( .A(n10853), .B(n10854), .Z(n10851) );
  NAND U13185 ( .A(n6856), .B(n6919), .Z(n10854) );
  NAND U13186 ( .A(n6858), .B(n6937), .Z(n10853) );
  AND U13187 ( .A(n10855), .B(n9125), .Z(n10849) );
  NAND U13188 ( .A(n6966), .B(n8603), .Z(n9125) );
  AND U13189 ( .A(n8485), .B(n10856), .Z(n10855) );
  NAND U13190 ( .A(n6943), .B(n8487), .Z(n10856) );
  NAND U13191 ( .A(n6865), .B(n8606), .Z(n8485) );
  AND U13192 ( .A(n10857), .B(n10858), .Z(n10847) );
  AND U13193 ( .A(n10859), .B(n10860), .Z(n10858) );
  AND U13194 ( .A(n10861), .B(n10862), .Z(n10859) );
  AND U13195 ( .A(n10863), .B(n10864), .Z(n10857) );
  AND U13196 ( .A(n10865), .B(n10866), .Z(n10863) );
  IV U13197 ( .A(\u_a23_core/u_execute/rn[23] ), .Z(n10734) );
  AND U13198 ( .A(n9395), .B(n10867), .Z(n10725) );
  NAND U13199 ( .A(n6765), .B(\u_a23_core/u_execute/u_alu/fadder_out[23] ), 
        .Z(n10867) );
  AND U13200 ( .A(n10868), .B(n10869), .Z(n10721) );
  NANDN U13201 ( .B(n8406), .A(\u_a23_core/u_execute/rn_plus4[23] ), .Z(n10869) );
  NANDN U13202 ( .B(n8407), .A(\u_a23_core/u_execute/alu_plus4[23] ), .Z(
        n10868) );
  AND U13203 ( .A(n10870), .B(n10871), .Z(n10719) );
  AND U13204 ( .A(n10872), .B(n10873), .Z(n10871) );
  NAND U13205 ( .A(n8412), .B(\u_a23_core/u_execute/address_plus4[23] ), .Z(
        n10873) );
  NAND U13206 ( .A(\u_a23_core/u_execute/rn[23] ), .B(n8413), .Z(n10872) );
  NAND U13207 ( .A(n10874), .B(n10875), .Z(\u_a23_core/u_execute/rn[23] ) );
  AND U13208 ( .A(n10876), .B(n10877), .Z(n10875) );
  AND U13209 ( .A(n10878), .B(n10879), .Z(n10877) );
  AND U13210 ( .A(n10880), .B(n10881), .Z(n10879) );
  NANDN U13211 ( .B(n8635), .A(\u_a23_core/u_execute/pc[23] ), .Z(n10881) );
  NANDN U13212 ( .B(n8636), .A(\u_a23_core/u_execute/u_register_bank/r14[23] ), 
        .Z(n10880) );
  AND U13213 ( .A(n10882), .B(n10883), .Z(n10878) );
  NANDN U13214 ( .B(n8639), .A(\u_a23_core/u_execute/u_register_bank/r13[23] ), 
        .Z(n10883) );
  NANDN U13215 ( .B(n8640), .A(\u_a23_core/u_execute/u_register_bank/r12[23] ), 
        .Z(n10882) );
  AND U13216 ( .A(n10884), .B(n10885), .Z(n10876) );
  AND U13217 ( .A(n10886), .B(n10887), .Z(n10885) );
  NANDN U13218 ( .B(n8645), .A(\u_a23_core/u_execute/u_register_bank/r11[23] ), 
        .Z(n10887) );
  NANDN U13219 ( .B(n8646), .A(\u_a23_core/u_execute/u_register_bank/r10[23] ), 
        .Z(n10886) );
  AND U13220 ( .A(n10888), .B(n10889), .Z(n10884) );
  NANDN U13221 ( .B(n8649), .A(\u_a23_core/u_execute/u_register_bank/r9[23] ), 
        .Z(n10889) );
  NANDN U13222 ( .B(n8650), .A(\u_a23_core/u_execute/u_register_bank/r8[23] ), 
        .Z(n10888) );
  AND U13223 ( .A(n10890), .B(n10891), .Z(n10874) );
  AND U13224 ( .A(n10892), .B(n10893), .Z(n10891) );
  AND U13225 ( .A(n10894), .B(n10895), .Z(n10893) );
  NANDN U13226 ( .B(n8657), .A(\u_a23_core/u_execute/u_register_bank/r7[23] ), 
        .Z(n10895) );
  NANDN U13227 ( .B(n8658), .A(\u_a23_core/u_execute/u_register_bank/r6[23] ), 
        .Z(n10894) );
  AND U13228 ( .A(n10896), .B(n10897), .Z(n10892) );
  NANDN U13229 ( .B(n8661), .A(\u_a23_core/u_execute/u_register_bank/r5[23] ), 
        .Z(n10897) );
  NANDN U13230 ( .B(n8662), .A(\u_a23_core/u_execute/u_register_bank/r4[23] ), 
        .Z(n10896) );
  AND U13231 ( .A(n10898), .B(n10899), .Z(n10890) );
  AND U13232 ( .A(n10900), .B(n10901), .Z(n10899) );
  NANDN U13233 ( .B(n8667), .A(\u_a23_core/u_execute/u_register_bank/r3[23] ), 
        .Z(n10901) );
  NANDN U13234 ( .B(n8668), .A(\u_a23_core/u_execute/u_register_bank/r0[23] ), 
        .Z(n10900) );
  AND U13235 ( .A(n10902), .B(n10903), .Z(n10898) );
  NANDN U13236 ( .B(n8671), .A(\u_a23_core/u_execute/u_register_bank/r2[23] ), 
        .Z(n10903) );
  NANDN U13237 ( .B(n8672), .A(\u_a23_core/u_execute/u_register_bank/r1[23] ), 
        .Z(n10902) );
  AND U13238 ( .A(n10904), .B(n10905), .Z(n10870) );
  NAND U13239 ( .A(\u_a23_core/u_execute/pc[23] ), .B(n8416), .Z(n10905) );
  NAND U13240 ( .A(n8417), .B(\u_a23_core/u_execute/pc_plus4[23] ), .Z(n10904)
         );
  NAND U13241 ( .A(n10906), .B(n10907), .Z(
        \u_a23_core/execute_address_nxt[22] ) );
  AND U13242 ( .A(n10908), .B(n10909), .Z(n10907) );
  AND U13243 ( .A(n10910), .B(n10911), .Z(n10909) );
  NANDN U13244 ( .B(n8392), .A(\u_a23_core/u_execute/pc_minus4[22] ), .Z(
        n10911) );
  NAND U13245 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[22] ), .B(n8393), 
        .Z(n10910) );
  IV U13246 ( .A(n7025), .Z(\u_a23_core/u_execute/alu_out_pc_filtered[22] ) );
  AND U13247 ( .A(n10912), .B(n10913), .Z(n7025) );
  MUX U13248 ( .IN0(n10914), .IN1(n10915), .SEL(
        \u_a23_core/u_execute/u_alu/b_not[22] ), .F(n10913) );
  NAND U13249 ( .A(n10916), .B(n10917), .Z(
        \u_a23_core/u_execute/u_alu/b_not[22] ) );
  MUX U13250 ( .IN0(n8430), .IN1(n8431), .SEL(n10918), .F(n10917) );
  MUX U13251 ( .IN0(n8433), .IN1(n8434), .SEL(\u_a23_core/u_execute/rn[22] ), 
        .F(n10916) );
  ANDN U13252 ( .A(n9256), .B(n10919), .Z(n10915) );
  MUX U13253 ( .IN0(n8400), .IN1(\u_a23_core/alu_function[3] ), .SEL(
        \u_a23_core/u_execute/u_alu/a[22] ), .F(n10919) );
  NAND U13254 ( .A(\u_a23_core/u_execute/u_alu/a[22] ), .B(n8400), .Z(n10914)
         );
  IV U13255 ( .A(n10920), .Z(\u_a23_core/u_execute/u_alu/a[22] ) );
  MUX U13256 ( .IN0(n10921), .IN1(n10918), .SEL(\u_a23_core/alu_function[8] ), 
        .F(n10920) );
  AND U13257 ( .A(n10922), .B(n10923), .Z(n10918) );
  AND U13258 ( .A(n10924), .B(n10925), .Z(n10923) );
  NAND U13259 ( .A(n10926), .B(n10552), .Z(n10925) );
  NAND U13260 ( .A(n10746), .B(n10927), .Z(n10926) );
  NAND U13261 ( .A(n8443), .B(n10928), .Z(n10927) );
  NAND U13262 ( .A(n10744), .B(n9515), .Z(n10928) );
  IV U13263 ( .A(n10929), .Z(n9515) );
  IV U13264 ( .A(n8603), .Z(n10746) );
  NAND U13265 ( .A(n6786), .B(n10930), .Z(n10924) );
  NAND U13266 ( .A(n10931), .B(n10932), .Z(n10930) );
  AND U13267 ( .A(n10933), .B(n10934), .Z(n10932) );
  AND U13268 ( .A(n10935), .B(n10936), .Z(n10934) );
  NAND U13269 ( .A(n8610), .B(n6799), .Z(n10936) );
  AND U13270 ( .A(n10937), .B(n10938), .Z(n10935) );
  NAND U13271 ( .A(n8606), .B(n6807), .Z(n10938) );
  NAND U13272 ( .A(n8609), .B(n6809), .Z(n10937) );
  AND U13273 ( .A(n9501), .B(n6976), .Z(n10933) );
  NAND U13274 ( .A(n8616), .B(n6803), .Z(n6976) );
  NAND U13275 ( .A(n8958), .B(n6823), .Z(n9501) );
  AND U13276 ( .A(n10939), .B(n10940), .Z(n10931) );
  AND U13277 ( .A(n10309), .B(n9945), .Z(n10940) );
  NAND U13278 ( .A(n9082), .B(n6827), .Z(n9945) );
  NAND U13279 ( .A(n9135), .B(n6833), .Z(n10309) );
  AND U13280 ( .A(n10941), .B(n10675), .Z(n10939) );
  NAND U13281 ( .A(n6984), .B(n6835), .Z(n10675) );
  NAND U13282 ( .A(n6893), .B(n6839), .Z(n10941) );
  AND U13283 ( .A(n10942), .B(n10943), .Z(n10922) );
  NAND U13284 ( .A(n10944), .B(n6888), .Z(n10943) );
  NAND U13285 ( .A(n10945), .B(n10946), .Z(n10944) );
  AND U13286 ( .A(n10947), .B(n10948), .Z(n10946) );
  AND U13287 ( .A(n10949), .B(n10950), .Z(n10948) );
  AND U13288 ( .A(n10951), .B(n10952), .Z(n10950) );
  AND U13289 ( .A(n10953), .B(n10954), .Z(n10952) );
  NANDN U13290 ( .B(n8561), .A(n6919), .Z(n10954) );
  NAND U13291 ( .A(n6839), .B(n8512), .Z(n10953) );
  AND U13292 ( .A(n10955), .B(n10956), .Z(n10951) );
  NANDN U13293 ( .B(n8562), .A(n6920), .Z(n10956) );
  NANDN U13294 ( .B(n8516), .A(n6850), .Z(n10955) );
  AND U13295 ( .A(n10957), .B(n10958), .Z(n10949) );
  AND U13296 ( .A(n10959), .B(n10960), .Z(n10958) );
  NANDN U13297 ( .B(n8567), .A(n6925), .Z(n10960) );
  NANDN U13298 ( .B(n8522), .A(n6853), .Z(n10959) );
  AND U13299 ( .A(n10961), .B(n10962), .Z(n10957) );
  NANDN U13300 ( .B(n8568), .A(n6926), .Z(n10962) );
  NANDN U13301 ( .B(n8526), .A(n6841), .Z(n10961) );
  AND U13302 ( .A(n10963), .B(n10964), .Z(n10947) );
  AND U13303 ( .A(n10965), .B(n10966), .Z(n10964) );
  AND U13304 ( .A(n10967), .B(n10968), .Z(n10966) );
  NANDN U13305 ( .B(n8571), .A(n6898), .Z(n10968) );
  NANDN U13306 ( .B(n8534), .A(n6857), .Z(n10967) );
  AND U13307 ( .A(n10969), .B(n10970), .Z(n10965) );
  NANDN U13308 ( .B(n8511), .A(n6859), .Z(n10970) );
  NANDN U13309 ( .B(n8572), .A(n6882), .Z(n10969) );
  AND U13310 ( .A(n10971), .B(n10972), .Z(n10963) );
  AND U13311 ( .A(n10973), .B(n10974), .Z(n10972) );
  NANDN U13312 ( .B(n8515), .A(n6865), .Z(n10974) );
  NANDN U13313 ( .B(n8579), .A(n6809), .Z(n10973) );
  AND U13314 ( .A(n10975), .B(n10976), .Z(n10971) );
  NANDN U13315 ( .B(n8521), .A(n6967), .Z(n10976) );
  NANDN U13316 ( .B(n8580), .A(n6807), .Z(n10975) );
  AND U13317 ( .A(n10977), .B(n10978), .Z(n10945) );
  AND U13318 ( .A(n10979), .B(n10980), .Z(n10978) );
  AND U13319 ( .A(n10981), .B(n10982), .Z(n10980) );
  AND U13320 ( .A(n10983), .B(n10984), .Z(n10982) );
  NANDN U13321 ( .B(n8525), .A(n6966), .Z(n10984) );
  NANDN U13322 ( .B(n8583), .A(n6799), .Z(n10983) );
  AND U13323 ( .A(n10985), .B(n10986), .Z(n10981) );
  NANDN U13324 ( .B(n8584), .A(n6803), .Z(n10986) );
  NANDN U13325 ( .B(n8533), .A(n6961), .Z(n10985) );
  AND U13326 ( .A(n10987), .B(n10988), .Z(n10979) );
  AND U13327 ( .A(n10989), .B(n10990), .Z(n10988) );
  NANDN U13328 ( .B(n8589), .A(n6823), .Z(n10990) );
  NANDN U13329 ( .B(n8537), .A(n6956), .Z(n10989) );
  AND U13330 ( .A(n10991), .B(n10992), .Z(n10987) );
  NANDN U13331 ( .B(n8590), .A(n6827), .Z(n10992) );
  NANDN U13332 ( .B(n8538), .A(n6960), .Z(n10991) );
  AND U13333 ( .A(n10993), .B(n10994), .Z(n10977) );
  AND U13334 ( .A(n10995), .B(n10996), .Z(n10994) );
  AND U13335 ( .A(n10997), .B(n10998), .Z(n10996) );
  NANDN U13336 ( .B(n8593), .A(n6833), .Z(n10998) );
  NANDN U13337 ( .B(n8543), .A(n6957), .Z(n10997) );
  AND U13338 ( .A(n10999), .B(n11000), .Z(n10995) );
  NAND U13339 ( .A(n6835), .B(n6897), .Z(n11000) );
  NANDN U13340 ( .B(n8544), .A(n6947), .Z(n10999) );
  AND U13341 ( .A(n11001), .B(n11002), .Z(n10993) );
  AND U13342 ( .A(n11003), .B(n11004), .Z(n11002) );
  NANDN U13343 ( .B(n8547), .A(n6946), .Z(n11004) );
  NANDN U13344 ( .B(n8548), .A(n6943), .Z(n11003) );
  AND U13345 ( .A(n11005), .B(n11006), .Z(n11001) );
  NANDN U13346 ( .B(n8557), .A(n6942), .Z(n11006) );
  NANDN U13347 ( .B(n8558), .A(n6937), .Z(n11005) );
  NAND U13348 ( .A(n11007), .B(n6902), .Z(n10942) );
  NAND U13349 ( .A(n11008), .B(n11009), .Z(n11007) );
  AND U13350 ( .A(n11010), .B(n11011), .Z(n11009) );
  AND U13351 ( .A(n11012), .B(n11013), .Z(n11011) );
  AND U13352 ( .A(n11014), .B(n11015), .Z(n11013) );
  NAND U13353 ( .A(n6916), .B(n6839), .Z(n11015) );
  ANDN U13354 ( .A(n8972), .B(n8711), .Z(n11014) );
  ANDN U13355 ( .A(n8606), .B(n10638), .Z(n8711) );
  IV U13356 ( .A(n6967), .Z(n10638) );
  NAND U13357 ( .A(n6966), .B(n8609), .Z(n8972) );
  AND U13358 ( .A(n11016), .B(n11017), .Z(n11012) );
  NAND U13359 ( .A(n8461), .B(n6947), .Z(n11017) );
  AND U13360 ( .A(n11018), .B(n11019), .Z(n11016) );
  NAND U13361 ( .A(n8464), .B(n6943), .Z(n11019) );
  NAND U13362 ( .A(n8465), .B(n6946), .Z(n11018) );
  AND U13363 ( .A(n11020), .B(n11021), .Z(n11010) );
  AND U13364 ( .A(n11022), .B(n11023), .Z(n11021) );
  AND U13365 ( .A(n11024), .B(n11025), .Z(n11022) );
  NAND U13366 ( .A(n8470), .B(n6957), .Z(n11025) );
  AND U13367 ( .A(n11026), .B(n11027), .Z(n11020) );
  NAND U13368 ( .A(n6852), .B(n6926), .Z(n11027) );
  AND U13369 ( .A(n11028), .B(n11029), .Z(n11026) );
  NAND U13370 ( .A(n6840), .B(n6925), .Z(n11029) );
  NAND U13371 ( .A(n6898), .B(n6851), .Z(n11028) );
  AND U13372 ( .A(n11030), .B(n11031), .Z(n11008) );
  AND U13373 ( .A(n11032), .B(n11033), .Z(n11031) );
  AND U13374 ( .A(n11034), .B(n11035), .Z(n11033) );
  NAND U13375 ( .A(n6864), .B(n6937), .Z(n11035) );
  AND U13376 ( .A(n11036), .B(n11037), .Z(n11034) );
  NAND U13377 ( .A(n6856), .B(n6920), .Z(n11037) );
  NAND U13378 ( .A(n6858), .B(n6919), .Z(n11036) );
  AND U13379 ( .A(n11038), .B(n11039), .Z(n11032) );
  AND U13380 ( .A(n11040), .B(n11041), .Z(n11038) );
  NAND U13381 ( .A(n6942), .B(n8487), .Z(n11041) );
  AND U13382 ( .A(n11042), .B(n11043), .Z(n11030) );
  AND U13383 ( .A(n11044), .B(n11045), .Z(n11043) );
  AND U13384 ( .A(n11046), .B(n11047), .Z(n11044) );
  AND U13385 ( .A(n11048), .B(n11049), .Z(n11042) );
  IV U13386 ( .A(\u_a23_core/u_execute/rn[22] ), .Z(n10921) );
  AND U13387 ( .A(n9395), .B(n11050), .Z(n10912) );
  NAND U13388 ( .A(n6765), .B(\u_a23_core/u_execute/u_alu/fadder_out[22] ), 
        .Z(n11050) );
  AND U13389 ( .A(n11051), .B(n11052), .Z(n10908) );
  NANDN U13390 ( .B(n8406), .A(\u_a23_core/u_execute/rn_plus4[22] ), .Z(n11052) );
  NANDN U13391 ( .B(n8407), .A(\u_a23_core/u_execute/alu_plus4[22] ), .Z(
        n11051) );
  AND U13392 ( .A(n11053), .B(n11054), .Z(n10906) );
  AND U13393 ( .A(n11055), .B(n11056), .Z(n11054) );
  NAND U13394 ( .A(n8412), .B(\u_a23_core/u_execute/address_plus4[22] ), .Z(
        n11056) );
  NAND U13395 ( .A(\u_a23_core/u_execute/rn[22] ), .B(n8413), .Z(n11055) );
  NAND U13396 ( .A(n11057), .B(n11058), .Z(\u_a23_core/u_execute/rn[22] ) );
  AND U13397 ( .A(n11059), .B(n11060), .Z(n11058) );
  AND U13398 ( .A(n11061), .B(n11062), .Z(n11060) );
  AND U13399 ( .A(n11063), .B(n11064), .Z(n11062) );
  NANDN U13400 ( .B(n8635), .A(\u_a23_core/u_execute/pc[22] ), .Z(n11064) );
  NANDN U13401 ( .B(n8636), .A(\u_a23_core/u_execute/u_register_bank/r14[22] ), 
        .Z(n11063) );
  AND U13402 ( .A(n11065), .B(n11066), .Z(n11061) );
  NANDN U13403 ( .B(n8639), .A(\u_a23_core/u_execute/u_register_bank/r13[22] ), 
        .Z(n11066) );
  NANDN U13404 ( .B(n8640), .A(\u_a23_core/u_execute/u_register_bank/r12[22] ), 
        .Z(n11065) );
  AND U13405 ( .A(n11067), .B(n11068), .Z(n11059) );
  AND U13406 ( .A(n11069), .B(n11070), .Z(n11068) );
  NANDN U13407 ( .B(n8645), .A(\u_a23_core/u_execute/u_register_bank/r11[22] ), 
        .Z(n11070) );
  NANDN U13408 ( .B(n8646), .A(\u_a23_core/u_execute/u_register_bank/r10[22] ), 
        .Z(n11069) );
  AND U13409 ( .A(n11071), .B(n11072), .Z(n11067) );
  NANDN U13410 ( .B(n8649), .A(\u_a23_core/u_execute/u_register_bank/r9[22] ), 
        .Z(n11072) );
  NANDN U13411 ( .B(n8650), .A(\u_a23_core/u_execute/u_register_bank/r8[22] ), 
        .Z(n11071) );
  AND U13412 ( .A(n11073), .B(n11074), .Z(n11057) );
  AND U13413 ( .A(n11075), .B(n11076), .Z(n11074) );
  AND U13414 ( .A(n11077), .B(n11078), .Z(n11076) );
  NANDN U13415 ( .B(n8657), .A(\u_a23_core/u_execute/u_register_bank/r7[22] ), 
        .Z(n11078) );
  NANDN U13416 ( .B(n8658), .A(\u_a23_core/u_execute/u_register_bank/r6[22] ), 
        .Z(n11077) );
  AND U13417 ( .A(n11079), .B(n11080), .Z(n11075) );
  NANDN U13418 ( .B(n8661), .A(\u_a23_core/u_execute/u_register_bank/r5[22] ), 
        .Z(n11080) );
  NANDN U13419 ( .B(n8662), .A(\u_a23_core/u_execute/u_register_bank/r4[22] ), 
        .Z(n11079) );
  AND U13420 ( .A(n11081), .B(n11082), .Z(n11073) );
  AND U13421 ( .A(n11083), .B(n11084), .Z(n11082) );
  NANDN U13422 ( .B(n8667), .A(\u_a23_core/u_execute/u_register_bank/r3[22] ), 
        .Z(n11084) );
  NANDN U13423 ( .B(n8668), .A(\u_a23_core/u_execute/u_register_bank/r0[22] ), 
        .Z(n11083) );
  AND U13424 ( .A(n11085), .B(n11086), .Z(n11081) );
  NANDN U13425 ( .B(n8671), .A(\u_a23_core/u_execute/u_register_bank/r2[22] ), 
        .Z(n11086) );
  NANDN U13426 ( .B(n8672), .A(\u_a23_core/u_execute/u_register_bank/r1[22] ), 
        .Z(n11085) );
  AND U13427 ( .A(n11087), .B(n11088), .Z(n11053) );
  NAND U13428 ( .A(\u_a23_core/u_execute/pc[22] ), .B(n8416), .Z(n11088) );
  NAND U13429 ( .A(n8417), .B(\u_a23_core/u_execute/pc_plus4[22] ), .Z(n11087)
         );
  NOR U13430 ( .A(\u_a23_core/execute_address_nxt[20] ), .B(
        \u_a23_core/execute_address_nxt[21] ), .Z(n10717) );
  NAND U13431 ( .A(n11089), .B(n11090), .Z(
        \u_a23_core/execute_address_nxt[21] ) );
  AND U13432 ( .A(n11091), .B(n11092), .Z(n11090) );
  AND U13433 ( .A(n11093), .B(n11094), .Z(n11092) );
  NANDN U13434 ( .B(n8392), .A(\u_a23_core/u_execute/pc_minus4[21] ), .Z(
        n11094) );
  NAND U13435 ( .A(n8393), .B(\u_a23_core/u_execute/alu_out_pc_filtered[21] ), 
        .Z(n11093) );
  IV U13436 ( .A(n7028), .Z(\u_a23_core/u_execute/alu_out_pc_filtered[21] ) );
  AND U13437 ( .A(n11095), .B(n11096), .Z(n7028) );
  MUX U13438 ( .IN0(n11097), .IN1(n11098), .SEL(
        \u_a23_core/u_execute/u_alu/b_not[21] ), .F(n11096) );
  NAND U13439 ( .A(n11099), .B(n11100), .Z(
        \u_a23_core/u_execute/u_alu/b_not[21] ) );
  MUX U13440 ( .IN0(n8430), .IN1(n8431), .SEL(n11101), .F(n11100) );
  MUX U13441 ( .IN0(n8433), .IN1(n8434), .SEL(\u_a23_core/u_execute/rn[21] ), 
        .F(n11099) );
  ANDN U13442 ( .A(n9256), .B(n11102), .Z(n11098) );
  MUX U13443 ( .IN0(n8400), .IN1(\u_a23_core/alu_function[3] ), .SEL(
        \u_a23_core/u_execute/u_alu/a[21] ), .F(n11102) );
  NAND U13444 ( .A(\u_a23_core/u_execute/u_alu/a[21] ), .B(n8400), .Z(n11097)
         );
  IV U13445 ( .A(n11103), .Z(\u_a23_core/u_execute/u_alu/a[21] ) );
  MUX U13446 ( .IN0(n11104), .IN1(n11101), .SEL(\u_a23_core/alu_function[8] ), 
        .F(n11103) );
  AND U13447 ( .A(n11105), .B(n11106), .Z(n11101) );
  AND U13448 ( .A(n11107), .B(n11108), .Z(n11106) );
  NAND U13449 ( .A(n11109), .B(n10552), .Z(n11108) );
  ANDN U13450 ( .A(n6786), .B(n11110), .Z(n10552) );
  NAND U13451 ( .A(n10744), .B(n11111), .Z(n11109) );
  NAND U13452 ( .A(n10929), .B(n8443), .Z(n11111) );
  IV U13453 ( .A(n9726), .Z(n10744) );
  NAND U13454 ( .A(n6786), .B(n11112), .Z(n11107) );
  NAND U13455 ( .A(n11113), .B(n11114), .Z(n11112) );
  AND U13456 ( .A(n11115), .B(n11116), .Z(n11114) );
  AND U13457 ( .A(n11117), .B(n11118), .Z(n11116) );
  NAND U13458 ( .A(n8609), .B(n6807), .Z(n11118) );
  AND U13459 ( .A(n11119), .B(n11120), .Z(n11117) );
  NAND U13460 ( .A(n8606), .B(n6799), .Z(n11120) );
  NAND U13461 ( .A(n8603), .B(n6809), .Z(n11119) );
  AND U13462 ( .A(n9392), .B(n11121), .Z(n11115) );
  NAND U13463 ( .A(n8610), .B(n6803), .Z(n11121) );
  NAND U13464 ( .A(n8616), .B(n6823), .Z(n9392) );
  AND U13465 ( .A(n11122), .B(n11123), .Z(n11113) );
  AND U13466 ( .A(n11124), .B(n10490), .Z(n11123) );
  NAND U13467 ( .A(n9135), .B(n6835), .Z(n10490) );
  AND U13468 ( .A(n10127), .B(n9755), .Z(n11124) );
  NAND U13469 ( .A(n8958), .B(n6827), .Z(n9755) );
  NAND U13470 ( .A(n9082), .B(n6833), .Z(n10127) );
  AND U13471 ( .A(n11125), .B(n10864), .Z(n11122) );
  NAND U13472 ( .A(n6984), .B(n6839), .Z(n10864) );
  NAND U13473 ( .A(n6850), .B(n6893), .Z(n11125) );
  AND U13474 ( .A(n11126), .B(n11127), .Z(n11105) );
  NAND U13475 ( .A(n11128), .B(n6888), .Z(n11127) );
  NAND U13476 ( .A(n11129), .B(n11130), .Z(n11128) );
  AND U13477 ( .A(n11131), .B(n11132), .Z(n11130) );
  AND U13478 ( .A(n11133), .B(n11134), .Z(n11132) );
  AND U13479 ( .A(n11135), .B(n11136), .Z(n11134) );
  AND U13480 ( .A(n11137), .B(n11138), .Z(n11136) );
  NANDN U13481 ( .B(n8558), .A(n6919), .Z(n11138) );
  NAND U13482 ( .A(n6850), .B(n8512), .Z(n11137) );
  AND U13483 ( .A(n11139), .B(n11140), .Z(n11135) );
  NANDN U13484 ( .B(n8561), .A(n6920), .Z(n11140) );
  NANDN U13485 ( .B(n8516), .A(n6853), .Z(n11139) );
  AND U13486 ( .A(n11141), .B(n11142), .Z(n11133) );
  AND U13487 ( .A(n11143), .B(n11144), .Z(n11142) );
  NANDN U13488 ( .B(n8562), .A(n6925), .Z(n11144) );
  NANDN U13489 ( .B(n8522), .A(n6841), .Z(n11143) );
  AND U13490 ( .A(n11145), .B(n11146), .Z(n11141) );
  NANDN U13491 ( .B(n8567), .A(n6926), .Z(n11146) );
  NANDN U13492 ( .B(n8526), .A(n6857), .Z(n11145) );
  AND U13493 ( .A(n11147), .B(n11148), .Z(n11131) );
  AND U13494 ( .A(n11149), .B(n11150), .Z(n11148) );
  AND U13495 ( .A(n11151), .B(n11152), .Z(n11150) );
  NANDN U13496 ( .B(n8568), .A(n6898), .Z(n11152) );
  NANDN U13497 ( .B(n8534), .A(n6859), .Z(n11151) );
  AND U13498 ( .A(n11153), .B(n11154), .Z(n11149) );
  NANDN U13499 ( .B(n8511), .A(n6865), .Z(n11154) );
  NANDN U13500 ( .B(n8571), .A(n6882), .Z(n11153) );
  AND U13501 ( .A(n11155), .B(n11156), .Z(n11147) );
  AND U13502 ( .A(n11157), .B(n11158), .Z(n11156) );
  NANDN U13503 ( .B(n8515), .A(n6967), .Z(n11158) );
  NANDN U13504 ( .B(n8572), .A(n6809), .Z(n11157) );
  AND U13505 ( .A(n11159), .B(n11160), .Z(n11155) );
  NANDN U13506 ( .B(n8521), .A(n6966), .Z(n11160) );
  NANDN U13507 ( .B(n8579), .A(n6807), .Z(n11159) );
  AND U13508 ( .A(n11161), .B(n11162), .Z(n11129) );
  AND U13509 ( .A(n11163), .B(n11164), .Z(n11162) );
  AND U13510 ( .A(n11165), .B(n11166), .Z(n11164) );
  AND U13511 ( .A(n11167), .B(n11168), .Z(n11166) );
  NANDN U13512 ( .B(n8525), .A(n6961), .Z(n11168) );
  NANDN U13513 ( .B(n8580), .A(n6799), .Z(n11167) );
  AND U13514 ( .A(n11169), .B(n11170), .Z(n11165) );
  NANDN U13515 ( .B(n8583), .A(n6803), .Z(n11170) );
  NANDN U13516 ( .B(n8533), .A(n6956), .Z(n11169) );
  AND U13517 ( .A(n11171), .B(n11172), .Z(n11163) );
  AND U13518 ( .A(n11173), .B(n11174), .Z(n11172) );
  NANDN U13519 ( .B(n8584), .A(n6823), .Z(n11174) );
  NANDN U13520 ( .B(n8537), .A(n6960), .Z(n11173) );
  AND U13521 ( .A(n11175), .B(n11176), .Z(n11171) );
  NANDN U13522 ( .B(n8589), .A(n6827), .Z(n11176) );
  NANDN U13523 ( .B(n8538), .A(n6957), .Z(n11175) );
  AND U13524 ( .A(n11177), .B(n11178), .Z(n11161) );
  AND U13525 ( .A(n11179), .B(n11180), .Z(n11178) );
  AND U13526 ( .A(n11181), .B(n11182), .Z(n11180) );
  NANDN U13527 ( .B(n8590), .A(n6833), .Z(n11182) );
  NANDN U13528 ( .B(n8543), .A(n6947), .Z(n11181) );
  AND U13529 ( .A(n11183), .B(n11184), .Z(n11179) );
  NANDN U13530 ( .B(n8593), .A(n6835), .Z(n11184) );
  NANDN U13531 ( .B(n8544), .A(n6946), .Z(n11183) );
  AND U13532 ( .A(n11185), .B(n11186), .Z(n11177) );
  AND U13533 ( .A(n11187), .B(n11188), .Z(n11186) );
  NAND U13534 ( .A(n6839), .B(n6897), .Z(n11188) );
  NANDN U13535 ( .B(n8547), .A(n6943), .Z(n11187) );
  AND U13536 ( .A(n11189), .B(n11190), .Z(n11185) );
  NANDN U13537 ( .B(n8548), .A(n6942), .Z(n11190) );
  NANDN U13538 ( .B(n8557), .A(n6937), .Z(n11189) );
  NAND U13539 ( .A(n11191), .B(n6902), .Z(n11126) );
  NAND U13540 ( .A(n11192), .B(n11193), .Z(n11191) );
  AND U13541 ( .A(n11194), .B(n11195), .Z(n11193) );
  AND U13542 ( .A(n11196), .B(n11197), .Z(n11195) );
  AND U13543 ( .A(n11198), .B(n11199), .Z(n11197) );
  NAND U13544 ( .A(n8464), .B(n6942), .Z(n11199) );
  ANDN U13545 ( .A(n11200), .B(n11201), .Z(n11198) );
  NAND U13546 ( .A(n6850), .B(n6916), .Z(n11200) );
  AND U13547 ( .A(n11202), .B(n11203), .Z(n11196) );
  NAND U13548 ( .A(n8470), .B(n6947), .Z(n11203) );
  AND U13549 ( .A(n11204), .B(n11205), .Z(n11202) );
  NAND U13550 ( .A(n8465), .B(n6943), .Z(n11205) );
  NAND U13551 ( .A(n8461), .B(n6946), .Z(n11204) );
  AND U13552 ( .A(n11206), .B(n11207), .Z(n11194) );
  AND U13553 ( .A(n11208), .B(n11209), .Z(n11207) );
  NAND U13554 ( .A(n6840), .B(n6926), .Z(n11209) );
  AND U13555 ( .A(n11210), .B(n6820), .Z(n11208) );
  NAND U13556 ( .A(n9359), .B(n6957), .Z(n6820) );
  AND U13557 ( .A(n11211), .B(n11212), .Z(n11206) );
  NAND U13558 ( .A(n6852), .B(n6898), .Z(n11212) );
  NAND U13559 ( .A(n6856), .B(n6925), .Z(n11211) );
  AND U13560 ( .A(n11213), .B(n11214), .Z(n11192) );
  AND U13561 ( .A(n11215), .B(n11216), .Z(n11214) );
  AND U13562 ( .A(n11217), .B(n11218), .Z(n11216) );
  NAND U13563 ( .A(n6937), .B(n8487), .Z(n11218) );
  AND U13564 ( .A(n11219), .B(n11220), .Z(n11217) );
  NAND U13565 ( .A(n6858), .B(n6920), .Z(n11220) );
  NAND U13566 ( .A(n6864), .B(n6919), .Z(n11219) );
  AND U13567 ( .A(n11221), .B(n8490), .Z(n11215) );
  NAND U13568 ( .A(n6967), .B(n8610), .Z(n8490) );
  AND U13569 ( .A(n9124), .B(n11222), .Z(n11221) );
  NAND U13570 ( .A(n6961), .B(n8609), .Z(n9124) );
  AND U13571 ( .A(n11223), .B(n11224), .Z(n11213) );
  AND U13572 ( .A(n11225), .B(n11226), .Z(n11224) );
  AND U13573 ( .A(n11227), .B(n11228), .Z(n11225) );
  AND U13574 ( .A(n11229), .B(n11230), .Z(n11223) );
  IV U13575 ( .A(\u_a23_core/u_execute/rn[21] ), .Z(n11104) );
  AND U13576 ( .A(n9395), .B(n11231), .Z(n11095) );
  NAND U13577 ( .A(n6765), .B(\u_a23_core/u_execute/u_alu/fadder_out[21] ), 
        .Z(n11231) );
  AND U13578 ( .A(n11232), .B(n11233), .Z(n11091) );
  NANDN U13579 ( .B(n8406), .A(\u_a23_core/u_execute/rn_plus4[21] ), .Z(n11233) );
  NANDN U13580 ( .B(n8407), .A(\u_a23_core/u_execute/alu_plus4[21] ), .Z(
        n11232) );
  AND U13581 ( .A(n11234), .B(n11235), .Z(n11089) );
  AND U13582 ( .A(n11236), .B(n11237), .Z(n11235) );
  NAND U13583 ( .A(n8412), .B(\u_a23_core/u_execute/address_plus4[21] ), .Z(
        n11237) );
  NAND U13584 ( .A(\u_a23_core/u_execute/rn[21] ), .B(n8413), .Z(n11236) );
  NAND U13585 ( .A(n11238), .B(n11239), .Z(\u_a23_core/u_execute/rn[21] ) );
  AND U13586 ( .A(n11240), .B(n11241), .Z(n11239) );
  AND U13587 ( .A(n11242), .B(n11243), .Z(n11241) );
  AND U13588 ( .A(n11244), .B(n11245), .Z(n11243) );
  NANDN U13589 ( .B(n8635), .A(\u_a23_core/u_execute/pc[21] ), .Z(n11245) );
  NANDN U13590 ( .B(n8636), .A(\u_a23_core/u_execute/u_register_bank/r14[21] ), 
        .Z(n11244) );
  AND U13591 ( .A(n11246), .B(n11247), .Z(n11242) );
  NANDN U13592 ( .B(n8639), .A(\u_a23_core/u_execute/u_register_bank/r13[21] ), 
        .Z(n11247) );
  NANDN U13593 ( .B(n8640), .A(\u_a23_core/u_execute/u_register_bank/r12[21] ), 
        .Z(n11246) );
  AND U13594 ( .A(n11248), .B(n11249), .Z(n11240) );
  AND U13595 ( .A(n11250), .B(n11251), .Z(n11249) );
  NANDN U13596 ( .B(n8645), .A(\u_a23_core/u_execute/u_register_bank/r11[21] ), 
        .Z(n11251) );
  NANDN U13597 ( .B(n8646), .A(\u_a23_core/u_execute/u_register_bank/r10[21] ), 
        .Z(n11250) );
  AND U13598 ( .A(n11252), .B(n11253), .Z(n11248) );
  NANDN U13599 ( .B(n8649), .A(\u_a23_core/u_execute/u_register_bank/r9[21] ), 
        .Z(n11253) );
  NANDN U13600 ( .B(n8650), .A(\u_a23_core/u_execute/u_register_bank/r8[21] ), 
        .Z(n11252) );
  AND U13601 ( .A(n11254), .B(n11255), .Z(n11238) );
  AND U13602 ( .A(n11256), .B(n11257), .Z(n11255) );
  AND U13603 ( .A(n11258), .B(n11259), .Z(n11257) );
  NANDN U13604 ( .B(n8657), .A(\u_a23_core/u_execute/u_register_bank/r7[21] ), 
        .Z(n11259) );
  NANDN U13605 ( .B(n8658), .A(\u_a23_core/u_execute/u_register_bank/r6[21] ), 
        .Z(n11258) );
  AND U13606 ( .A(n11260), .B(n11261), .Z(n11256) );
  NANDN U13607 ( .B(n8661), .A(\u_a23_core/u_execute/u_register_bank/r5[21] ), 
        .Z(n11261) );
  NANDN U13608 ( .B(n8662), .A(\u_a23_core/u_execute/u_register_bank/r4[21] ), 
        .Z(n11260) );
  AND U13609 ( .A(n11262), .B(n11263), .Z(n11254) );
  AND U13610 ( .A(n11264), .B(n11265), .Z(n11263) );
  NANDN U13611 ( .B(n8667), .A(\u_a23_core/u_execute/u_register_bank/r3[21] ), 
        .Z(n11265) );
  NANDN U13612 ( .B(n8668), .A(\u_a23_core/u_execute/u_register_bank/r0[21] ), 
        .Z(n11264) );
  AND U13613 ( .A(n11266), .B(n11267), .Z(n11262) );
  NANDN U13614 ( .B(n8671), .A(\u_a23_core/u_execute/u_register_bank/r2[21] ), 
        .Z(n11267) );
  NANDN U13615 ( .B(n8672), .A(\u_a23_core/u_execute/u_register_bank/r1[21] ), 
        .Z(n11266) );
  AND U13616 ( .A(n11268), .B(n11269), .Z(n11234) );
  NAND U13617 ( .A(\u_a23_core/u_execute/pc[21] ), .B(n8416), .Z(n11269) );
  NAND U13618 ( .A(n8417), .B(\u_a23_core/u_execute/pc_plus4[21] ), .Z(n11268)
         );
  NAND U13619 ( .A(n11270), .B(n11271), .Z(
        \u_a23_core/execute_address_nxt[20] ) );
  AND U13620 ( .A(n11272), .B(n11273), .Z(n11271) );
  AND U13621 ( .A(n11274), .B(n11275), .Z(n11273) );
  NANDN U13622 ( .B(n8392), .A(\u_a23_core/u_execute/pc_minus4[20] ), .Z(
        n11275) );
  NAND U13623 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[20] ), .B(n8393), 
        .Z(n11274) );
  IV U13624 ( .A(n7029), .Z(\u_a23_core/u_execute/alu_out_pc_filtered[20] ) );
  AND U13625 ( .A(n11276), .B(n11277), .Z(n7029) );
  MUX U13626 ( .IN0(n11278), .IN1(n11279), .SEL(
        \u_a23_core/u_execute/u_alu/b_not[20] ), .F(n11277) );
  NAND U13627 ( .A(n11280), .B(n11281), .Z(
        \u_a23_core/u_execute/u_alu/b_not[20] ) );
  MUX U13628 ( .IN0(n8430), .IN1(n8431), .SEL(n11282), .F(n11281) );
  MUX U13629 ( .IN0(n8433), .IN1(n8434), .SEL(\u_a23_core/u_execute/rn[20] ), 
        .F(n11280) );
  ANDN U13630 ( .A(n9256), .B(n11283), .Z(n11279) );
  MUX U13631 ( .IN0(n8400), .IN1(\u_a23_core/alu_function[3] ), .SEL(
        \u_a23_core/u_execute/u_alu/a[20] ), .F(n11283) );
  NAND U13632 ( .A(\u_a23_core/u_execute/u_alu/a[20] ), .B(n8400), .Z(n11278)
         );
  IV U13633 ( .A(n11284), .Z(\u_a23_core/u_execute/u_alu/a[20] ) );
  MUX U13634 ( .IN0(n11285), .IN1(n11282), .SEL(\u_a23_core/alu_function[8] ), 
        .F(n11284) );
  AND U13635 ( .A(n11286), .B(n11287), .Z(n11282) );
  AND U13636 ( .A(n11288), .B(n11289), .Z(n11287) );
  NAND U13637 ( .A(n6786), .B(n11290), .Z(n11289) );
  NAND U13638 ( .A(n11291), .B(n11292), .Z(n11290) );
  AND U13639 ( .A(n11293), .B(n11294), .Z(n11292) );
  AND U13640 ( .A(n11295), .B(n11296), .Z(n11294) );
  NAND U13641 ( .A(n8603), .B(n6807), .Z(n11296) );
  AND U13642 ( .A(n11297), .B(n11298), .Z(n11295) );
  NAND U13643 ( .A(n9726), .B(n6809), .Z(n11298) );
  NAND U13644 ( .A(n8606), .B(n6803), .Z(n11297) );
  AND U13645 ( .A(n11299), .B(n9502), .Z(n11293) );
  NAND U13646 ( .A(n8616), .B(n6827), .Z(n9502) );
  AND U13647 ( .A(n6977), .B(n11300), .Z(n11299) );
  NAND U13648 ( .A(n8609), .B(n6799), .Z(n11300) );
  NAND U13649 ( .A(n8610), .B(n6823), .Z(n6977) );
  AND U13650 ( .A(n11301), .B(n11302), .Z(n11291) );
  AND U13651 ( .A(n11303), .B(n10676), .Z(n11302) );
  NAND U13652 ( .A(n9135), .B(n6839), .Z(n10676) );
  AND U13653 ( .A(n10310), .B(n9940), .Z(n11303) );
  NAND U13654 ( .A(n8958), .B(n6833), .Z(n9940) );
  NAND U13655 ( .A(n9082), .B(n6835), .Z(n10310) );
  AND U13656 ( .A(n11304), .B(n11048), .Z(n11301) );
  NAND U13657 ( .A(n6850), .B(n6984), .Z(n11048) );
  NAND U13658 ( .A(n6893), .B(n6853), .Z(n11304) );
  AND U13659 ( .A(n11305), .B(n11306), .Z(n11288) );
  NAND U13660 ( .A(n10929), .B(n6886), .Z(n11306) );
  NAND U13661 ( .A(n11307), .B(n11308), .Z(n10929) );
  AND U13662 ( .A(n9884), .B(n11309), .Z(n11308) );
  IV U13663 ( .A(n9359), .Z(n9884) );
  AND U13664 ( .A(n11310), .B(n11311), .Z(n11307) );
  NAND U13665 ( .A(n9359), .B(n6985), .Z(n11305) );
  AND U13666 ( .A(n11312), .B(n11313), .Z(n11286) );
  NAND U13667 ( .A(n11314), .B(n6888), .Z(n11313) );
  NAND U13668 ( .A(n11315), .B(n11316), .Z(n11314) );
  AND U13669 ( .A(n11317), .B(n11318), .Z(n11316) );
  AND U13670 ( .A(n11319), .B(n11320), .Z(n11318) );
  AND U13671 ( .A(n11321), .B(n11322), .Z(n11320) );
  AND U13672 ( .A(n11323), .B(n11324), .Z(n11322) );
  NANDN U13673 ( .B(n8557), .A(n6919), .Z(n11324) );
  NAND U13674 ( .A(n6853), .B(n8512), .Z(n11323) );
  AND U13675 ( .A(n11325), .B(n11326), .Z(n11321) );
  NANDN U13676 ( .B(n8558), .A(n6920), .Z(n11326) );
  NANDN U13677 ( .B(n8516), .A(n6841), .Z(n11325) );
  AND U13678 ( .A(n11327), .B(n11328), .Z(n11319) );
  AND U13679 ( .A(n11329), .B(n11330), .Z(n11328) );
  NANDN U13680 ( .B(n8561), .A(n6925), .Z(n11330) );
  NANDN U13681 ( .B(n8522), .A(n6857), .Z(n11329) );
  AND U13682 ( .A(n11331), .B(n11332), .Z(n11327) );
  NANDN U13683 ( .B(n8562), .A(n6926), .Z(n11332) );
  NANDN U13684 ( .B(n8526), .A(n6859), .Z(n11331) );
  AND U13685 ( .A(n11333), .B(n11334), .Z(n11317) );
  AND U13686 ( .A(n11335), .B(n11336), .Z(n11334) );
  AND U13687 ( .A(n11337), .B(n11338), .Z(n11336) );
  NANDN U13688 ( .B(n8567), .A(n6898), .Z(n11338) );
  NANDN U13689 ( .B(n8534), .A(n6865), .Z(n11337) );
  AND U13690 ( .A(n11339), .B(n11340), .Z(n11335) );
  NANDN U13691 ( .B(n8511), .A(n6967), .Z(n11340) );
  NANDN U13692 ( .B(n8568), .A(n6882), .Z(n11339) );
  AND U13693 ( .A(n11341), .B(n11342), .Z(n11333) );
  AND U13694 ( .A(n11343), .B(n11344), .Z(n11342) );
  NANDN U13695 ( .B(n8515), .A(n6966), .Z(n11344) );
  NANDN U13696 ( .B(n8571), .A(n6809), .Z(n11343) );
  AND U13697 ( .A(n11345), .B(n11346), .Z(n11341) );
  NANDN U13698 ( .B(n8521), .A(n6961), .Z(n11346) );
  NANDN U13699 ( .B(n8572), .A(n6807), .Z(n11345) );
  AND U13700 ( .A(n11347), .B(n11348), .Z(n11315) );
  AND U13701 ( .A(n11349), .B(n11350), .Z(n11348) );
  AND U13702 ( .A(n11351), .B(n11352), .Z(n11350) );
  AND U13703 ( .A(n11353), .B(n11354), .Z(n11352) );
  NANDN U13704 ( .B(n8525), .A(n6956), .Z(n11354) );
  NANDN U13705 ( .B(n8579), .A(n6799), .Z(n11353) );
  AND U13706 ( .A(n11355), .B(n11356), .Z(n11351) );
  NANDN U13707 ( .B(n8580), .A(n6803), .Z(n11356) );
  NANDN U13708 ( .B(n8533), .A(n6960), .Z(n11355) );
  AND U13709 ( .A(n11357), .B(n11358), .Z(n11349) );
  AND U13710 ( .A(n11359), .B(n11360), .Z(n11358) );
  NANDN U13711 ( .B(n8583), .A(n6823), .Z(n11360) );
  NANDN U13712 ( .B(n8537), .A(n6957), .Z(n11359) );
  AND U13713 ( .A(n11361), .B(n11362), .Z(n11357) );
  NANDN U13714 ( .B(n8584), .A(n6827), .Z(n11362) );
  NANDN U13715 ( .B(n8538), .A(n6947), .Z(n11361) );
  AND U13716 ( .A(n11363), .B(n11364), .Z(n11347) );
  AND U13717 ( .A(n11365), .B(n11366), .Z(n11364) );
  AND U13718 ( .A(n11367), .B(n11368), .Z(n11366) );
  NANDN U13719 ( .B(n8589), .A(n6833), .Z(n11368) );
  NANDN U13720 ( .B(n8543), .A(n6946), .Z(n11367) );
  AND U13721 ( .A(n11369), .B(n11370), .Z(n11365) );
  NANDN U13722 ( .B(n8590), .A(n6835), .Z(n11370) );
  NANDN U13723 ( .B(n8544), .A(n6943), .Z(n11369) );
  AND U13724 ( .A(n11371), .B(n11372), .Z(n11363) );
  AND U13725 ( .A(n11373), .B(n11374), .Z(n11372) );
  NANDN U13726 ( .B(n8593), .A(n6839), .Z(n11374) );
  NANDN U13727 ( .B(n8547), .A(n6942), .Z(n11373) );
  AND U13728 ( .A(n11375), .B(n11376), .Z(n11371) );
  NAND U13729 ( .A(n6850), .B(n6897), .Z(n11376) );
  NANDN U13730 ( .B(n8548), .A(n6937), .Z(n11375) );
  NAND U13731 ( .A(n11377), .B(n6902), .Z(n11312) );
  NAND U13732 ( .A(n11378), .B(n11379), .Z(n11377) );
  AND U13733 ( .A(n11380), .B(n11381), .Z(n11379) );
  AND U13734 ( .A(n11382), .B(n11383), .Z(n11381) );
  AND U13735 ( .A(n11384), .B(n11385), .Z(n11383) );
  NAND U13736 ( .A(n6916), .B(n6853), .Z(n11385) );
  NOR U13737 ( .A(n8975), .B(n8706), .Z(n11384) );
  ANDN U13738 ( .A(n8610), .B(n11386), .Z(n8706) );
  ANDN U13739 ( .A(n8606), .B(n11387), .Z(n8975) );
  IV U13740 ( .A(n6961), .Z(n11387) );
  AND U13741 ( .A(n11388), .B(n11389), .Z(n11382) );
  NAND U13742 ( .A(n8461), .B(n6943), .Z(n11389) );
  AND U13743 ( .A(n11390), .B(n11391), .Z(n11388) );
  NAND U13744 ( .A(n8464), .B(n6937), .Z(n11391) );
  NAND U13745 ( .A(n8465), .B(n6942), .Z(n11390) );
  AND U13746 ( .A(n11392), .B(n11393), .Z(n11380) );
  AND U13747 ( .A(n11394), .B(n11395), .Z(n11393) );
  AND U13748 ( .A(n11396), .B(n11397), .Z(n11394) );
  NAND U13749 ( .A(n8470), .B(n6946), .Z(n11397) );
  NAND U13750 ( .A(n9359), .B(n6947), .Z(n11396) );
  AND U13751 ( .A(n11398), .B(n11399), .Z(n11392) );
  NAND U13752 ( .A(n6840), .B(n6898), .Z(n11399) );
  NAND U13753 ( .A(n6856), .B(n6926), .Z(n11398) );
  AND U13754 ( .A(n11400), .B(n11401), .Z(n11378) );
  AND U13755 ( .A(n11402), .B(n11403), .Z(n11401) );
  AND U13756 ( .A(n11404), .B(n11405), .Z(n11403) );
  NAND U13757 ( .A(n6919), .B(n8487), .Z(n11405) );
  AND U13758 ( .A(n11406), .B(n11407), .Z(n11404) );
  NAND U13759 ( .A(n6858), .B(n6925), .Z(n11407) );
  NAND U13760 ( .A(n6864), .B(n6920), .Z(n11406) );
  AND U13761 ( .A(n11408), .B(n11409), .Z(n11402) );
  AND U13762 ( .A(n11410), .B(n11411), .Z(n11400) );
  AND U13763 ( .A(n11412), .B(n11413), .Z(n11411) );
  AND U13764 ( .A(n11414), .B(n11415), .Z(n11412) );
  AND U13765 ( .A(n11416), .B(n11417), .Z(n11410) );
  IV U13766 ( .A(\u_a23_core/u_execute/rn[20] ), .Z(n11285) );
  AND U13767 ( .A(n9395), .B(n11418), .Z(n11276) );
  NAND U13768 ( .A(n6765), .B(\u_a23_core/u_execute/u_alu/fadder_out[20] ), 
        .Z(n11418) );
  AND U13769 ( .A(n11419), .B(n11420), .Z(n11272) );
  NANDN U13770 ( .B(n8406), .A(\u_a23_core/u_execute/rn_plus4[20] ), .Z(n11420) );
  NANDN U13771 ( .B(n8407), .A(\u_a23_core/u_execute/alu_plus4[20] ), .Z(
        n11419) );
  AND U13772 ( .A(n11421), .B(n11422), .Z(n11270) );
  AND U13773 ( .A(n11423), .B(n11424), .Z(n11422) );
  NAND U13774 ( .A(n8412), .B(\u_a23_core/u_execute/address_plus4[20] ), .Z(
        n11424) );
  NAND U13775 ( .A(\u_a23_core/u_execute/rn[20] ), .B(n8413), .Z(n11423) );
  NAND U13776 ( .A(n11425), .B(n11426), .Z(\u_a23_core/u_execute/rn[20] ) );
  AND U13777 ( .A(n11427), .B(n11428), .Z(n11426) );
  AND U13778 ( .A(n11429), .B(n11430), .Z(n11428) );
  AND U13779 ( .A(n11431), .B(n11432), .Z(n11430) );
  NANDN U13780 ( .B(n8635), .A(\u_a23_core/u_execute/pc[20] ), .Z(n11432) );
  NANDN U13781 ( .B(n8636), .A(\u_a23_core/u_execute/u_register_bank/r14[20] ), 
        .Z(n11431) );
  AND U13782 ( .A(n11433), .B(n11434), .Z(n11429) );
  NANDN U13783 ( .B(n8639), .A(\u_a23_core/u_execute/u_register_bank/r13[20] ), 
        .Z(n11434) );
  NANDN U13784 ( .B(n8640), .A(\u_a23_core/u_execute/u_register_bank/r12[20] ), 
        .Z(n11433) );
  AND U13785 ( .A(n11435), .B(n11436), .Z(n11427) );
  AND U13786 ( .A(n11437), .B(n11438), .Z(n11436) );
  NANDN U13787 ( .B(n8645), .A(\u_a23_core/u_execute/u_register_bank/r11[20] ), 
        .Z(n11438) );
  NANDN U13788 ( .B(n8646), .A(\u_a23_core/u_execute/u_register_bank/r10[20] ), 
        .Z(n11437) );
  AND U13789 ( .A(n11439), .B(n11440), .Z(n11435) );
  NANDN U13790 ( .B(n8649), .A(\u_a23_core/u_execute/u_register_bank/r9[20] ), 
        .Z(n11440) );
  NANDN U13791 ( .B(n8650), .A(\u_a23_core/u_execute/u_register_bank/r8[20] ), 
        .Z(n11439) );
  AND U13792 ( .A(n11441), .B(n11442), .Z(n11425) );
  AND U13793 ( .A(n11443), .B(n11444), .Z(n11442) );
  AND U13794 ( .A(n11445), .B(n11446), .Z(n11444) );
  NANDN U13795 ( .B(n8657), .A(\u_a23_core/u_execute/u_register_bank/r7[20] ), 
        .Z(n11446) );
  NANDN U13796 ( .B(n8658), .A(\u_a23_core/u_execute/u_register_bank/r6[20] ), 
        .Z(n11445) );
  AND U13797 ( .A(n11447), .B(n11448), .Z(n11443) );
  NANDN U13798 ( .B(n8661), .A(\u_a23_core/u_execute/u_register_bank/r5[20] ), 
        .Z(n11448) );
  NANDN U13799 ( .B(n8662), .A(\u_a23_core/u_execute/u_register_bank/r4[20] ), 
        .Z(n11447) );
  AND U13800 ( .A(n11449), .B(n11450), .Z(n11441) );
  AND U13801 ( .A(n11451), .B(n11452), .Z(n11450) );
  NANDN U13802 ( .B(n8667), .A(\u_a23_core/u_execute/u_register_bank/r3[20] ), 
        .Z(n11452) );
  NANDN U13803 ( .B(n8668), .A(\u_a23_core/u_execute/u_register_bank/r0[20] ), 
        .Z(n11451) );
  AND U13804 ( .A(n11453), .B(n11454), .Z(n11449) );
  NANDN U13805 ( .B(n8671), .A(\u_a23_core/u_execute/u_register_bank/r2[20] ), 
        .Z(n11454) );
  NANDN U13806 ( .B(n8672), .A(\u_a23_core/u_execute/u_register_bank/r1[20] ), 
        .Z(n11453) );
  AND U13807 ( .A(n11455), .B(n11456), .Z(n11421) );
  NAND U13808 ( .A(\u_a23_core/u_execute/pc[20] ), .B(n8416), .Z(n11456) );
  NAND U13809 ( .A(n8417), .B(\u_a23_core/u_execute/pc_plus4[20] ), .Z(n11455)
         );
  AND U13810 ( .A(n11457), .B(n11458), .Z(n8377) );
  AND U13811 ( .A(n11459), .B(n11460), .Z(n11458) );
  AND U13812 ( .A(n11461), .B(n11462), .Z(n11460) );
  ANDN U13813 ( .A(n11463), .B(\u_a23_core/execute_address_nxt[18] ), .Z(
        n11462) );
  NAND U13814 ( .A(n11464), .B(n11465), .Z(
        \u_a23_core/execute_address_nxt[18] ) );
  AND U13815 ( .A(n11466), .B(n11467), .Z(n11465) );
  AND U13816 ( .A(n11468), .B(n11469), .Z(n11467) );
  NANDN U13817 ( .B(n8392), .A(\u_a23_core/u_execute/pc_minus4[18] ), .Z(
        n11469) );
  NAND U13818 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[18] ), .B(n8393), 
        .Z(n11468) );
  IV U13819 ( .A(n7031), .Z(\u_a23_core/u_execute/alu_out_pc_filtered[18] ) );
  AND U13820 ( .A(n11470), .B(n11471), .Z(n7031) );
  MUX U13821 ( .IN0(n11472), .IN1(n11473), .SEL(
        \u_a23_core/u_execute/u_alu/b_not[18] ), .F(n11471) );
  NAND U13822 ( .A(n11474), .B(n11475), .Z(
        \u_a23_core/u_execute/u_alu/b_not[18] ) );
  MUX U13823 ( .IN0(n8430), .IN1(n8431), .SEL(n11476), .F(n11475) );
  MUX U13824 ( .IN0(n8433), .IN1(n8434), .SEL(\u_a23_core/u_execute/rn[18] ), 
        .F(n11474) );
  ANDN U13825 ( .A(n9256), .B(n11477), .Z(n11473) );
  MUX U13826 ( .IN0(n8400), .IN1(\u_a23_core/alu_function[3] ), .SEL(
        \u_a23_core/u_execute/u_alu/a[18] ), .F(n11477) );
  NAND U13827 ( .A(\u_a23_core/u_execute/u_alu/a[18] ), .B(n8400), .Z(n11472)
         );
  IV U13828 ( .A(n11478), .Z(\u_a23_core/u_execute/u_alu/a[18] ) );
  MUX U13829 ( .IN0(n11479), .IN1(n11476), .SEL(\u_a23_core/alu_function[8] ), 
        .F(n11478) );
  AND U13830 ( .A(n11480), .B(n11481), .Z(n11476) );
  AND U13831 ( .A(n11482), .B(n11483), .Z(n11481) );
  NAND U13832 ( .A(n6786), .B(n11484), .Z(n11483) );
  NAND U13833 ( .A(n11485), .B(n11486), .Z(n11484) );
  AND U13834 ( .A(n11487), .B(n11488), .Z(n11486) );
  AND U13835 ( .A(n11489), .B(n11490), .Z(n11488) );
  AND U13836 ( .A(n11491), .B(n11492), .Z(n11490) );
  NAND U13837 ( .A(n8470), .B(n6809), .Z(n11492) );
  NAND U13838 ( .A(n9359), .B(n6807), .Z(n11491) );
  AND U13839 ( .A(n6968), .B(n11493), .Z(n11489) );
  NAND U13840 ( .A(n9726), .B(n6799), .Z(n11493) );
  NAND U13841 ( .A(n8606), .B(n6827), .Z(n6968) );
  AND U13842 ( .A(n11494), .B(n9499), .Z(n11487) );
  NAND U13843 ( .A(n8610), .B(n6833), .Z(n9499) );
  AND U13844 ( .A(n11495), .B(n11496), .Z(n11494) );
  NAND U13845 ( .A(n8603), .B(n6803), .Z(n11496) );
  NAND U13846 ( .A(n8609), .B(n6823), .Z(n11495) );
  AND U13847 ( .A(n11497), .B(n11498), .Z(n11485) );
  AND U13848 ( .A(n11499), .B(n10677), .Z(n11498) );
  NAND U13849 ( .A(n6850), .B(n9082), .Z(n10677) );
  AND U13850 ( .A(n10304), .B(n9941), .Z(n11499) );
  NAND U13851 ( .A(n8616), .B(n6835), .Z(n9941) );
  NAND U13852 ( .A(n8958), .B(n6839), .Z(n10304) );
  AND U13853 ( .A(n11500), .B(n11501), .Z(n11497) );
  NAND U13854 ( .A(n6893), .B(n6857), .Z(n11501) );
  AND U13855 ( .A(n11416), .B(n11049), .Z(n11500) );
  NAND U13856 ( .A(n9135), .B(n6853), .Z(n11049) );
  NAND U13857 ( .A(n6984), .B(n6841), .Z(n11416) );
  AND U13858 ( .A(n11502), .B(n11503), .Z(n11482) );
  NAND U13859 ( .A(n6886), .B(n11504), .Z(n11503) );
  NAND U13860 ( .A(n8461), .B(n6985), .Z(n11502) );
  AND U13861 ( .A(n11505), .B(n11506), .Z(n11480) );
  NAND U13862 ( .A(n11507), .B(n6888), .Z(n11506) );
  NAND U13863 ( .A(n11508), .B(n11509), .Z(n11507) );
  AND U13864 ( .A(n11510), .B(n11511), .Z(n11509) );
  AND U13865 ( .A(n11512), .B(n11513), .Z(n11511) );
  AND U13866 ( .A(n11514), .B(n11515), .Z(n11513) );
  AND U13867 ( .A(n11516), .B(n11517), .Z(n11515) );
  NANDN U13868 ( .B(n8547), .A(n6919), .Z(n11517) );
  NAND U13869 ( .A(n6857), .B(n8512), .Z(n11516) );
  AND U13870 ( .A(n11518), .B(n11519), .Z(n11514) );
  NANDN U13871 ( .B(n8548), .A(n6920), .Z(n11519) );
  NANDN U13872 ( .B(n8516), .A(n6859), .Z(n11518) );
  AND U13873 ( .A(n11520), .B(n11521), .Z(n11512) );
  AND U13874 ( .A(n11522), .B(n11523), .Z(n11521) );
  NANDN U13875 ( .B(n8557), .A(n6925), .Z(n11523) );
  NANDN U13876 ( .B(n8522), .A(n6865), .Z(n11522) );
  AND U13877 ( .A(n11524), .B(n11525), .Z(n11520) );
  NANDN U13878 ( .B(n8558), .A(n6926), .Z(n11525) );
  NANDN U13879 ( .B(n8526), .A(n6967), .Z(n11524) );
  AND U13880 ( .A(n11526), .B(n11527), .Z(n11510) );
  AND U13881 ( .A(n11528), .B(n11529), .Z(n11527) );
  AND U13882 ( .A(n11530), .B(n11531), .Z(n11529) );
  NANDN U13883 ( .B(n8561), .A(n6898), .Z(n11531) );
  NANDN U13884 ( .B(n8534), .A(n6966), .Z(n11530) );
  AND U13885 ( .A(n11532), .B(n11533), .Z(n11528) );
  NANDN U13886 ( .B(n8511), .A(n6961), .Z(n11533) );
  NANDN U13887 ( .B(n8562), .A(n6882), .Z(n11532) );
  AND U13888 ( .A(n11534), .B(n11535), .Z(n11526) );
  AND U13889 ( .A(n11536), .B(n11537), .Z(n11535) );
  NANDN U13890 ( .B(n8515), .A(n6956), .Z(n11537) );
  NANDN U13891 ( .B(n8567), .A(n6809), .Z(n11536) );
  AND U13892 ( .A(n11538), .B(n11539), .Z(n11534) );
  NANDN U13893 ( .B(n8521), .A(n6960), .Z(n11539) );
  NANDN U13894 ( .B(n8568), .A(n6807), .Z(n11538) );
  AND U13895 ( .A(n11540), .B(n11541), .Z(n11508) );
  AND U13896 ( .A(n11542), .B(n11543), .Z(n11541) );
  AND U13897 ( .A(n11544), .B(n11545), .Z(n11543) );
  AND U13898 ( .A(n11546), .B(n11547), .Z(n11545) );
  NANDN U13899 ( .B(n8525), .A(n6957), .Z(n11547) );
  NANDN U13900 ( .B(n8571), .A(n6799), .Z(n11546) );
  AND U13901 ( .A(n11548), .B(n11549), .Z(n11544) );
  NANDN U13902 ( .B(n8572), .A(n6803), .Z(n11549) );
  NANDN U13903 ( .B(n8533), .A(n6947), .Z(n11548) );
  AND U13904 ( .A(n11550), .B(n11551), .Z(n11542) );
  AND U13905 ( .A(n11552), .B(n11553), .Z(n11551) );
  NANDN U13906 ( .B(n8579), .A(n6823), .Z(n11553) );
  NANDN U13907 ( .B(n8537), .A(n6946), .Z(n11552) );
  AND U13908 ( .A(n11554), .B(n11555), .Z(n11550) );
  NANDN U13909 ( .B(n8580), .A(n6827), .Z(n11555) );
  NANDN U13910 ( .B(n8538), .A(n6943), .Z(n11554) );
  AND U13911 ( .A(n11556), .B(n11557), .Z(n11540) );
  AND U13912 ( .A(n11558), .B(n11559), .Z(n11557) );
  AND U13913 ( .A(n11560), .B(n11561), .Z(n11559) );
  NANDN U13914 ( .B(n8583), .A(n6833), .Z(n11561) );
  NANDN U13915 ( .B(n8543), .A(n6942), .Z(n11560) );
  AND U13916 ( .A(n11562), .B(n11563), .Z(n11558) );
  NANDN U13917 ( .B(n8584), .A(n6835), .Z(n11563) );
  NANDN U13918 ( .B(n8544), .A(n6937), .Z(n11562) );
  AND U13919 ( .A(n11564), .B(n11565), .Z(n11556) );
  AND U13920 ( .A(n11566), .B(n11567), .Z(n11565) );
  NANDN U13921 ( .B(n8589), .A(n6839), .Z(n11567) );
  NANDN U13922 ( .B(n8590), .A(n6850), .Z(n11566) );
  AND U13923 ( .A(n11568), .B(n11569), .Z(n11564) );
  NANDN U13924 ( .B(n8593), .A(n6853), .Z(n11569) );
  NAND U13925 ( .A(n6841), .B(n6897), .Z(n11568) );
  NAND U13926 ( .A(n11570), .B(n6902), .Z(n11505) );
  NAND U13927 ( .A(n11571), .B(n11572), .Z(n11570) );
  AND U13928 ( .A(n11573), .B(n11574), .Z(n11572) );
  AND U13929 ( .A(n11575), .B(n11576), .Z(n11574) );
  AND U13930 ( .A(n11577), .B(n11578), .Z(n11576) );
  NAND U13931 ( .A(n8464), .B(n6920), .Z(n11578) );
  ANDN U13932 ( .A(n11579), .B(n8973), .Z(n11577) );
  ANDN U13933 ( .A(n8610), .B(n11580), .Z(n8973) );
  IV U13934 ( .A(n6956), .Z(n11580) );
  NAND U13935 ( .A(n6916), .B(n6857), .Z(n11579) );
  AND U13936 ( .A(n11581), .B(n11582), .Z(n11575) );
  NAND U13937 ( .A(n8465), .B(n6919), .Z(n11582) );
  NAND U13938 ( .A(n8461), .B(n6937), .Z(n11581) );
  AND U13939 ( .A(n11583), .B(n11584), .Z(n11573) );
  AND U13940 ( .A(n11585), .B(n11586), .Z(n11584) );
  NAND U13941 ( .A(n9726), .B(n6946), .Z(n11586) );
  AND U13942 ( .A(n11587), .B(n11588), .Z(n11585) );
  NAND U13943 ( .A(n8470), .B(n6942), .Z(n11588) );
  NAND U13944 ( .A(n9359), .B(n6943), .Z(n11587) );
  AND U13945 ( .A(n11589), .B(n11590), .Z(n11583) );
  NAND U13946 ( .A(n6858), .B(n6898), .Z(n11590) );
  NAND U13947 ( .A(n6864), .B(n6926), .Z(n11589) );
  AND U13948 ( .A(n11591), .B(n11592), .Z(n11571) );
  AND U13949 ( .A(n11593), .B(n11594), .Z(n11592) );
  AND U13950 ( .A(n11595), .B(n11596), .Z(n11594) );
  AND U13951 ( .A(n11597), .B(n11598), .Z(n11595) );
  NAND U13952 ( .A(n6925), .B(n8487), .Z(n11598) );
  AND U13953 ( .A(n8738), .B(n11599), .Z(n11593) );
  NAND U13954 ( .A(n6961), .B(n8616), .Z(n8738) );
  AND U13955 ( .A(n11600), .B(n11601), .Z(n11591) );
  AND U13956 ( .A(n11602), .B(n11603), .Z(n11601) );
  AND U13957 ( .A(n11604), .B(n11605), .Z(n11600) );
  IV U13958 ( .A(\u_a23_core/u_execute/rn[18] ), .Z(n11479) );
  AND U13959 ( .A(n9395), .B(n11606), .Z(n11470) );
  NAND U13960 ( .A(n6765), .B(\u_a23_core/u_execute/u_alu/fadder_out[18] ), 
        .Z(n11606) );
  AND U13961 ( .A(n11607), .B(n11608), .Z(n11466) );
  NANDN U13962 ( .B(n8406), .A(\u_a23_core/u_execute/rn_plus4[18] ), .Z(n11608) );
  NANDN U13963 ( .B(n8407), .A(\u_a23_core/u_execute/alu_plus4[18] ), .Z(
        n11607) );
  AND U13964 ( .A(n11609), .B(n11610), .Z(n11464) );
  AND U13965 ( .A(n11611), .B(n11612), .Z(n11610) );
  NAND U13966 ( .A(n8412), .B(\u_a23_core/u_execute/address_plus4[18] ), .Z(
        n11612) );
  NAND U13967 ( .A(\u_a23_core/u_execute/rn[18] ), .B(n8413), .Z(n11611) );
  NAND U13968 ( .A(n11613), .B(n11614), .Z(\u_a23_core/u_execute/rn[18] ) );
  AND U13969 ( .A(n11615), .B(n11616), .Z(n11614) );
  AND U13970 ( .A(n11617), .B(n11618), .Z(n11616) );
  AND U13971 ( .A(n11619), .B(n11620), .Z(n11618) );
  NANDN U13972 ( .B(n8635), .A(\u_a23_core/u_execute/pc[18] ), .Z(n11620) );
  NANDN U13973 ( .B(n8636), .A(\u_a23_core/u_execute/u_register_bank/r14[18] ), 
        .Z(n11619) );
  AND U13974 ( .A(n11621), .B(n11622), .Z(n11617) );
  NANDN U13975 ( .B(n8639), .A(\u_a23_core/u_execute/u_register_bank/r13[18] ), 
        .Z(n11622) );
  NANDN U13976 ( .B(n8640), .A(\u_a23_core/u_execute/u_register_bank/r12[18] ), 
        .Z(n11621) );
  AND U13977 ( .A(n11623), .B(n11624), .Z(n11615) );
  AND U13978 ( .A(n11625), .B(n11626), .Z(n11624) );
  NANDN U13979 ( .B(n8645), .A(\u_a23_core/u_execute/u_register_bank/r11[18] ), 
        .Z(n11626) );
  NANDN U13980 ( .B(n8646), .A(\u_a23_core/u_execute/u_register_bank/r10[18] ), 
        .Z(n11625) );
  AND U13981 ( .A(n11627), .B(n11628), .Z(n11623) );
  NANDN U13982 ( .B(n8649), .A(\u_a23_core/u_execute/u_register_bank/r9[18] ), 
        .Z(n11628) );
  NANDN U13983 ( .B(n8650), .A(\u_a23_core/u_execute/u_register_bank/r8[18] ), 
        .Z(n11627) );
  AND U13984 ( .A(n11629), .B(n11630), .Z(n11613) );
  AND U13985 ( .A(n11631), .B(n11632), .Z(n11630) );
  AND U13986 ( .A(n11633), .B(n11634), .Z(n11632) );
  NANDN U13987 ( .B(n8657), .A(\u_a23_core/u_execute/u_register_bank/r7[18] ), 
        .Z(n11634) );
  NANDN U13988 ( .B(n8658), .A(\u_a23_core/u_execute/u_register_bank/r6[18] ), 
        .Z(n11633) );
  AND U13989 ( .A(n11635), .B(n11636), .Z(n11631) );
  NANDN U13990 ( .B(n8661), .A(\u_a23_core/u_execute/u_register_bank/r5[18] ), 
        .Z(n11636) );
  NANDN U13991 ( .B(n8662), .A(\u_a23_core/u_execute/u_register_bank/r4[18] ), 
        .Z(n11635) );
  AND U13992 ( .A(n11637), .B(n11638), .Z(n11629) );
  AND U13993 ( .A(n11639), .B(n11640), .Z(n11638) );
  NANDN U13994 ( .B(n8667), .A(\u_a23_core/u_execute/u_register_bank/r3[18] ), 
        .Z(n11640) );
  NANDN U13995 ( .B(n8668), .A(\u_a23_core/u_execute/u_register_bank/r0[18] ), 
        .Z(n11639) );
  AND U13996 ( .A(n11641), .B(n11642), .Z(n11637) );
  NANDN U13997 ( .B(n8671), .A(\u_a23_core/u_execute/u_register_bank/r2[18] ), 
        .Z(n11642) );
  NANDN U13998 ( .B(n8672), .A(\u_a23_core/u_execute/u_register_bank/r1[18] ), 
        .Z(n11641) );
  AND U13999 ( .A(n11643), .B(n11644), .Z(n11609) );
  NAND U14000 ( .A(\u_a23_core/u_execute/pc[18] ), .B(n8416), .Z(n11644) );
  NAND U14001 ( .A(n8417), .B(\u_a23_core/u_execute/pc_plus4[18] ), .Z(n11643)
         );
  NOR U14002 ( .A(\u_a23_core/execute_address_nxt[1] ), .B(
        \u_a23_core/execute_address_nxt[19] ), .Z(n11463) );
  NAND U14003 ( .A(n11645), .B(n11646), .Z(
        \u_a23_core/execute_address_nxt[19] ) );
  AND U14004 ( .A(n11647), .B(n11648), .Z(n11646) );
  AND U14005 ( .A(n11649), .B(n11650), .Z(n11648) );
  NANDN U14006 ( .B(n8392), .A(\u_a23_core/u_execute/pc_minus4[19] ), .Z(
        n11650) );
  NAND U14007 ( .A(n8393), .B(\u_a23_core/u_execute/alu_out_pc_filtered[19] ), 
        .Z(n11649) );
  IV U14008 ( .A(n7030), .Z(\u_a23_core/u_execute/alu_out_pc_filtered[19] ) );
  AND U14009 ( .A(n11651), .B(n11652), .Z(n7030) );
  MUX U14010 ( .IN0(n11653), .IN1(n11654), .SEL(
        \u_a23_core/u_execute/u_alu/b_not[19] ), .F(n11652) );
  NAND U14011 ( .A(n11655), .B(n11656), .Z(
        \u_a23_core/u_execute/u_alu/b_not[19] ) );
  MUX U14012 ( .IN0(n8430), .IN1(n8431), .SEL(n11657), .F(n11656) );
  MUX U14013 ( .IN0(n8433), .IN1(n8434), .SEL(\u_a23_core/u_execute/rn[19] ), 
        .F(n11655) );
  ANDN U14014 ( .A(n9256), .B(n11658), .Z(n11654) );
  MUX U14015 ( .IN0(n8400), .IN1(\u_a23_core/alu_function[3] ), .SEL(
        \u_a23_core/u_execute/u_alu/a[19] ), .F(n11658) );
  NAND U14016 ( .A(\u_a23_core/u_execute/u_alu/a[19] ), .B(n8400), .Z(n11653)
         );
  IV U14017 ( .A(n11659), .Z(\u_a23_core/u_execute/u_alu/a[19] ) );
  MUX U14018 ( .IN0(n11660), .IN1(n11657), .SEL(\u_a23_core/alu_function[8] ), 
        .F(n11659) );
  AND U14019 ( .A(n11661), .B(n11662), .Z(n11657) );
  AND U14020 ( .A(n11663), .B(n11664), .Z(n11662) );
  NAND U14021 ( .A(n6786), .B(n11665), .Z(n11664) );
  NAND U14022 ( .A(n11666), .B(n11667), .Z(n11665) );
  AND U14023 ( .A(n11668), .B(n11669), .Z(n11667) );
  AND U14024 ( .A(n11670), .B(n11671), .Z(n11669) );
  NAND U14025 ( .A(n8606), .B(n6823), .Z(n11671) );
  AND U14026 ( .A(n11672), .B(n11673), .Z(n11670) );
  NAND U14027 ( .A(n9359), .B(n6809), .Z(n11673) );
  NAND U14028 ( .A(n9726), .B(n6807), .Z(n11672) );
  AND U14029 ( .A(n11674), .B(n9387), .Z(n11668) );
  NAND U14030 ( .A(n8610), .B(n6827), .Z(n9387) );
  AND U14031 ( .A(n11675), .B(n11676), .Z(n11674) );
  NAND U14032 ( .A(n8603), .B(n6799), .Z(n11676) );
  NAND U14033 ( .A(n8609), .B(n6803), .Z(n11675) );
  AND U14034 ( .A(n11677), .B(n11678), .Z(n11666) );
  AND U14035 ( .A(n11679), .B(n10491), .Z(n11678) );
  NAND U14036 ( .A(n9082), .B(n6839), .Z(n10491) );
  AND U14037 ( .A(n10122), .B(n9756), .Z(n11679) );
  NAND U14038 ( .A(n8616), .B(n6833), .Z(n9756) );
  NAND U14039 ( .A(n8958), .B(n6835), .Z(n10122) );
  AND U14040 ( .A(n11680), .B(n11681), .Z(n11677) );
  NAND U14041 ( .A(n6893), .B(n6841), .Z(n11681) );
  AND U14042 ( .A(n11229), .B(n10865), .Z(n11680) );
  NAND U14043 ( .A(n6850), .B(n9135), .Z(n10865) );
  NAND U14044 ( .A(n6984), .B(n6853), .Z(n11229) );
  AND U14045 ( .A(n11682), .B(n11683), .Z(n11663) );
  NAND U14046 ( .A(n11684), .B(n6886), .Z(n11683) );
  IV U14047 ( .A(n9885), .Z(n11684) );
  ANDN U14048 ( .A(n11309), .B(n11504), .Z(n9885) );
  NAND U14049 ( .A(n11685), .B(n11686), .Z(n11504) );
  AND U14050 ( .A(n11687), .B(n11311), .Z(n11686) );
  AND U14051 ( .A(n11688), .B(n11689), .Z(n11687) );
  IV U14052 ( .A(n8465), .Z(n11688) );
  AND U14053 ( .A(n11690), .B(n8448), .Z(n11685) );
  IV U14054 ( .A(n8470), .Z(n11309) );
  NAND U14055 ( .A(n8470), .B(n6985), .Z(n11682) );
  AND U14056 ( .A(n11691), .B(n11692), .Z(n11661) );
  NAND U14057 ( .A(n11693), .B(n6888), .Z(n11692) );
  NAND U14058 ( .A(n11694), .B(n11695), .Z(n11693) );
  AND U14059 ( .A(n11696), .B(n11697), .Z(n11695) );
  AND U14060 ( .A(n11698), .B(n11699), .Z(n11697) );
  AND U14061 ( .A(n11700), .B(n11701), .Z(n11699) );
  AND U14062 ( .A(n11702), .B(n11703), .Z(n11701) );
  NANDN U14063 ( .B(n8548), .A(n6919), .Z(n11703) );
  NAND U14064 ( .A(n6841), .B(n8512), .Z(n11702) );
  AND U14065 ( .A(n11704), .B(n11705), .Z(n11700) );
  NANDN U14066 ( .B(n8557), .A(n6920), .Z(n11705) );
  NANDN U14067 ( .B(n8516), .A(n6857), .Z(n11704) );
  AND U14068 ( .A(n11706), .B(n11707), .Z(n11698) );
  AND U14069 ( .A(n11708), .B(n11709), .Z(n11707) );
  NANDN U14070 ( .B(n8558), .A(n6925), .Z(n11709) );
  NANDN U14071 ( .B(n8522), .A(n6859), .Z(n11708) );
  AND U14072 ( .A(n11710), .B(n11711), .Z(n11706) );
  NANDN U14073 ( .B(n8561), .A(n6926), .Z(n11711) );
  NANDN U14074 ( .B(n8526), .A(n6865), .Z(n11710) );
  AND U14075 ( .A(n11712), .B(n11713), .Z(n11696) );
  AND U14076 ( .A(n11714), .B(n11715), .Z(n11713) );
  AND U14077 ( .A(n11716), .B(n11717), .Z(n11715) );
  NANDN U14078 ( .B(n8562), .A(n6898), .Z(n11717) );
  NANDN U14079 ( .B(n8534), .A(n6967), .Z(n11716) );
  AND U14080 ( .A(n11718), .B(n11719), .Z(n11714) );
  NANDN U14081 ( .B(n8511), .A(n6966), .Z(n11719) );
  NANDN U14082 ( .B(n8567), .A(n6882), .Z(n11718) );
  AND U14083 ( .A(n11720), .B(n11721), .Z(n11712) );
  AND U14084 ( .A(n11722), .B(n11723), .Z(n11721) );
  NANDN U14085 ( .B(n8515), .A(n6961), .Z(n11723) );
  NANDN U14086 ( .B(n8568), .A(n6809), .Z(n11722) );
  AND U14087 ( .A(n11724), .B(n11725), .Z(n11720) );
  NANDN U14088 ( .B(n8521), .A(n6956), .Z(n11725) );
  NANDN U14089 ( .B(n8571), .A(n6807), .Z(n11724) );
  AND U14090 ( .A(n11726), .B(n11727), .Z(n11694) );
  AND U14091 ( .A(n11728), .B(n11729), .Z(n11727) );
  AND U14092 ( .A(n11730), .B(n11731), .Z(n11729) );
  AND U14093 ( .A(n11732), .B(n11733), .Z(n11731) );
  NANDN U14094 ( .B(n8525), .A(n6960), .Z(n11733) );
  NANDN U14095 ( .B(n8572), .A(n6799), .Z(n11732) );
  AND U14096 ( .A(n11734), .B(n11735), .Z(n11730) );
  NANDN U14097 ( .B(n8579), .A(n6803), .Z(n11735) );
  NANDN U14098 ( .B(n8533), .A(n6957), .Z(n11734) );
  AND U14099 ( .A(n11736), .B(n11737), .Z(n11728) );
  AND U14100 ( .A(n11738), .B(n11739), .Z(n11737) );
  NANDN U14101 ( .B(n8580), .A(n6823), .Z(n11739) );
  NANDN U14102 ( .B(n8537), .A(n6947), .Z(n11738) );
  AND U14103 ( .A(n11740), .B(n11741), .Z(n11736) );
  NANDN U14104 ( .B(n8583), .A(n6827), .Z(n11741) );
  NANDN U14105 ( .B(n8538), .A(n6946), .Z(n11740) );
  AND U14106 ( .A(n11742), .B(n11743), .Z(n11726) );
  AND U14107 ( .A(n11744), .B(n11745), .Z(n11743) );
  AND U14108 ( .A(n11746), .B(n11747), .Z(n11745) );
  NANDN U14109 ( .B(n8584), .A(n6833), .Z(n11747) );
  NANDN U14110 ( .B(n8543), .A(n6943), .Z(n11746) );
  AND U14111 ( .A(n11748), .B(n11749), .Z(n11744) );
  NANDN U14112 ( .B(n8589), .A(n6835), .Z(n11749) );
  NANDN U14113 ( .B(n8544), .A(n6942), .Z(n11748) );
  AND U14114 ( .A(n11750), .B(n11751), .Z(n11742) );
  AND U14115 ( .A(n11752), .B(n11753), .Z(n11751) );
  NANDN U14116 ( .B(n8590), .A(n6839), .Z(n11753) );
  NANDN U14117 ( .B(n8547), .A(n6937), .Z(n11752) );
  AND U14118 ( .A(n11754), .B(n11755), .Z(n11750) );
  NANDN U14119 ( .B(n8593), .A(n6850), .Z(n11755) );
  NAND U14120 ( .A(n6853), .B(n6897), .Z(n11754) );
  NAND U14121 ( .A(n11756), .B(n6902), .Z(n11691) );
  NAND U14122 ( .A(n11757), .B(n11758), .Z(n11756) );
  AND U14123 ( .A(n11759), .B(n11760), .Z(n11758) );
  AND U14124 ( .A(n11761), .B(n11762), .Z(n11760) );
  AND U14125 ( .A(n11763), .B(n11764), .Z(n11762) );
  NAND U14126 ( .A(n8464), .B(n6919), .Z(n11764) );
  AND U14127 ( .A(n11765), .B(n11766), .Z(n11763) );
  NAND U14128 ( .A(n6916), .B(n6841), .Z(n11766) );
  AND U14129 ( .A(n11767), .B(n11768), .Z(n11761) );
  NAND U14130 ( .A(n8465), .B(n6937), .Z(n11768) );
  NAND U14131 ( .A(n8461), .B(n6942), .Z(n11767) );
  AND U14132 ( .A(n11769), .B(n11770), .Z(n11759) );
  AND U14133 ( .A(n11771), .B(n6825), .Z(n11770) );
  NAND U14134 ( .A(n9726), .B(n6947), .Z(n6825) );
  AND U14135 ( .A(n11772), .B(n11773), .Z(n11771) );
  NAND U14136 ( .A(n8470), .B(n6943), .Z(n11773) );
  NAND U14137 ( .A(n9359), .B(n6946), .Z(n11772) );
  AND U14138 ( .A(n11774), .B(n11775), .Z(n11769) );
  NAND U14139 ( .A(n6856), .B(n6898), .Z(n11775) );
  NAND U14140 ( .A(n6858), .B(n6926), .Z(n11774) );
  AND U14141 ( .A(n11776), .B(n11777), .Z(n11757) );
  AND U14142 ( .A(n11778), .B(n11779), .Z(n11777) );
  AND U14143 ( .A(n11780), .B(n9120), .Z(n11779) );
  NAND U14144 ( .A(n6956), .B(n8606), .Z(n9120) );
  AND U14145 ( .A(n11781), .B(n11782), .Z(n11780) );
  NAND U14146 ( .A(n6864), .B(n6925), .Z(n11782) );
  NAND U14147 ( .A(n6920), .B(n8487), .Z(n11781) );
  AND U14148 ( .A(n11783), .B(n11784), .Z(n11778) );
  AND U14149 ( .A(n11785), .B(n11786), .Z(n11776) );
  AND U14150 ( .A(n11787), .B(n11788), .Z(n11786) );
  AND U14151 ( .A(n11789), .B(n8489), .Z(n11787) );
  NAND U14152 ( .A(n6966), .B(n8616), .Z(n8489) );
  AND U14153 ( .A(n11790), .B(n11791), .Z(n11785) );
  IV U14154 ( .A(\u_a23_core/u_execute/rn[19] ), .Z(n11660) );
  AND U14155 ( .A(n9395), .B(n11792), .Z(n11651) );
  NAND U14156 ( .A(n6765), .B(\u_a23_core/u_execute/u_alu/fadder_out[19] ), 
        .Z(n11792) );
  AND U14157 ( .A(n11793), .B(n11794), .Z(n11647) );
  NANDN U14158 ( .B(n8406), .A(\u_a23_core/u_execute/rn_plus4[19] ), .Z(n11794) );
  NANDN U14159 ( .B(n8407), .A(\u_a23_core/u_execute/alu_plus4[19] ), .Z(
        n11793) );
  AND U14160 ( .A(n11795), .B(n11796), .Z(n11645) );
  AND U14161 ( .A(n11797), .B(n11798), .Z(n11796) );
  NAND U14162 ( .A(n8412), .B(\u_a23_core/u_execute/address_plus4[19] ), .Z(
        n11798) );
  NAND U14163 ( .A(\u_a23_core/u_execute/rn[19] ), .B(n8413), .Z(n11797) );
  NAND U14164 ( .A(n11799), .B(n11800), .Z(\u_a23_core/u_execute/rn[19] ) );
  AND U14165 ( .A(n11801), .B(n11802), .Z(n11800) );
  AND U14166 ( .A(n11803), .B(n11804), .Z(n11802) );
  AND U14167 ( .A(n11805), .B(n11806), .Z(n11804) );
  NANDN U14168 ( .B(n8635), .A(\u_a23_core/u_execute/pc[19] ), .Z(n11806) );
  NANDN U14169 ( .B(n8636), .A(\u_a23_core/u_execute/u_register_bank/r14[19] ), 
        .Z(n11805) );
  AND U14170 ( .A(n11807), .B(n11808), .Z(n11803) );
  NANDN U14171 ( .B(n8639), .A(\u_a23_core/u_execute/u_register_bank/r13[19] ), 
        .Z(n11808) );
  NANDN U14172 ( .B(n8640), .A(\u_a23_core/u_execute/u_register_bank/r12[19] ), 
        .Z(n11807) );
  AND U14173 ( .A(n11809), .B(n11810), .Z(n11801) );
  AND U14174 ( .A(n11811), .B(n11812), .Z(n11810) );
  NANDN U14175 ( .B(n8645), .A(\u_a23_core/u_execute/u_register_bank/r11[19] ), 
        .Z(n11812) );
  NANDN U14176 ( .B(n8646), .A(\u_a23_core/u_execute/u_register_bank/r10[19] ), 
        .Z(n11811) );
  AND U14177 ( .A(n11813), .B(n11814), .Z(n11809) );
  NANDN U14178 ( .B(n8649), .A(\u_a23_core/u_execute/u_register_bank/r9[19] ), 
        .Z(n11814) );
  NANDN U14179 ( .B(n8650), .A(\u_a23_core/u_execute/u_register_bank/r8[19] ), 
        .Z(n11813) );
  AND U14180 ( .A(n11815), .B(n11816), .Z(n11799) );
  AND U14181 ( .A(n11817), .B(n11818), .Z(n11816) );
  AND U14182 ( .A(n11819), .B(n11820), .Z(n11818) );
  NANDN U14183 ( .B(n8657), .A(\u_a23_core/u_execute/u_register_bank/r7[19] ), 
        .Z(n11820) );
  NANDN U14184 ( .B(n8658), .A(\u_a23_core/u_execute/u_register_bank/r6[19] ), 
        .Z(n11819) );
  AND U14185 ( .A(n11821), .B(n11822), .Z(n11817) );
  NANDN U14186 ( .B(n8661), .A(\u_a23_core/u_execute/u_register_bank/r5[19] ), 
        .Z(n11822) );
  NANDN U14187 ( .B(n8662), .A(\u_a23_core/u_execute/u_register_bank/r4[19] ), 
        .Z(n11821) );
  AND U14188 ( .A(n11823), .B(n11824), .Z(n11815) );
  AND U14189 ( .A(n11825), .B(n11826), .Z(n11824) );
  NANDN U14190 ( .B(n8667), .A(\u_a23_core/u_execute/u_register_bank/r3[19] ), 
        .Z(n11826) );
  NANDN U14191 ( .B(n8668), .A(\u_a23_core/u_execute/u_register_bank/r0[19] ), 
        .Z(n11825) );
  AND U14192 ( .A(n11827), .B(n11828), .Z(n11823) );
  NANDN U14193 ( .B(n8671), .A(\u_a23_core/u_execute/u_register_bank/r2[19] ), 
        .Z(n11828) );
  NANDN U14194 ( .B(n8672), .A(\u_a23_core/u_execute/u_register_bank/r1[19] ), 
        .Z(n11827) );
  AND U14195 ( .A(n11829), .B(n11830), .Z(n11795) );
  NAND U14196 ( .A(\u_a23_core/u_execute/pc[19] ), .B(n8416), .Z(n11830) );
  NAND U14197 ( .A(n8417), .B(\u_a23_core/u_execute/pc_plus4[19] ), .Z(n11829)
         );
  NAND U14198 ( .A(n11831), .B(n11832), .Z(\u_a23_core/execute_address_nxt[1] ) );
  NAND U14199 ( .A(n8412), .B(\u_a23_core/execute_address[1] ), .Z(n11832) );
  AND U14200 ( .A(n11833), .B(n11834), .Z(n11831) );
  NANDN U14201 ( .B(n11835), .A(n6337), .Z(n11834) );
  IV U14202 ( .A(n7059), .Z(n6337) );
  AND U14203 ( .A(n11836), .B(n11837), .Z(n7059) );
  MUX U14204 ( .IN0(n11838), .IN1(n11839), .SEL(
        \u_a23_core/u_execute/u_alu/b_not[1] ), .F(n11837) );
  NAND U14205 ( .A(n11840), .B(n11841), .Z(
        \u_a23_core/u_execute/u_alu/b_not[1] ) );
  MUX U14206 ( .IN0(n8430), .IN1(n8431), .SEL(n11842), .F(n11841) );
  MUX U14207 ( .IN0(n8434), .IN1(n8433), .SEL(n11843), .F(n11840) );
  ANDN U14208 ( .A(n8398), .B(n11844), .Z(n11839) );
  MUX U14209 ( .IN0(n8400), .IN1(\u_a23_core/alu_function[3] ), .SEL(
        \u_a23_core/u_execute/u_alu/a[1] ), .F(n11844) );
  NAND U14210 ( .A(\u_a23_core/u_execute/u_alu/a[1] ), .B(n8400), .Z(n11838)
         );
  IV U14211 ( .A(n11845), .Z(\u_a23_core/u_execute/u_alu/a[1] ) );
  MUX U14212 ( .IN0(n11843), .IN1(n11842), .SEL(\u_a23_core/alu_function[8] ), 
        .F(n11845) );
  AND U14213 ( .A(n11846), .B(n11847), .Z(n11842) );
  AND U14214 ( .A(n11848), .B(n11849), .Z(n11847) );
  NAND U14215 ( .A(n11850), .B(n6902), .Z(n11849) );
  NAND U14216 ( .A(n6881), .B(n11851), .Z(n11850) );
  NAND U14217 ( .A(n6926), .B(n6916), .Z(n11851) );
  NAND U14218 ( .A(n6984), .B(n6898), .Z(n6881) );
  AND U14219 ( .A(n11852), .B(n11853), .Z(n11846) );
  NAND U14220 ( .A(n6786), .B(n11854), .Z(n11853) );
  NAND U14221 ( .A(n11855), .B(n11856), .Z(n11854) );
  AND U14222 ( .A(n11857), .B(n11858), .Z(n11856) );
  AND U14223 ( .A(n11859), .B(n11860), .Z(n11858) );
  AND U14224 ( .A(n11861), .B(n11862), .Z(n11860) );
  AND U14225 ( .A(n11863), .B(n11864), .Z(n11862) );
  NAND U14226 ( .A(n6802), .B(n6807), .Z(n11864) );
  NAND U14227 ( .A(n6809), .B(n6798), .Z(n11863) );
  AND U14228 ( .A(n9352), .B(n11865), .Z(n11861) );
  NAND U14229 ( .A(n6882), .B(n6806), .Z(n11865) );
  NAND U14230 ( .A(n6865), .B(n8464), .Z(n9352) );
  AND U14231 ( .A(n11866), .B(n11867), .Z(n11859) );
  AND U14232 ( .A(n10087), .B(n9719), .Z(n11867) );
  NAND U14233 ( .A(n6967), .B(n8465), .Z(n9719) );
  NAND U14234 ( .A(n6966), .B(n8461), .Z(n10087) );
  AND U14235 ( .A(n11868), .B(n10459), .Z(n11866) );
  NAND U14236 ( .A(n6961), .B(n8470), .Z(n10459) );
  NAND U14237 ( .A(n6799), .B(n6822), .Z(n11868) );
  AND U14238 ( .A(n11869), .B(n11870), .Z(n11857) );
  AND U14239 ( .A(n11871), .B(n11872), .Z(n11870) );
  AND U14240 ( .A(n11210), .B(n10842), .Z(n11872) );
  NAND U14241 ( .A(n6956), .B(n9359), .Z(n10842) );
  NAND U14242 ( .A(n9726), .B(n6960), .Z(n11210) );
  AND U14243 ( .A(n11873), .B(n11874), .Z(n11871) );
  NAND U14244 ( .A(n6803), .B(n6826), .Z(n11874) );
  NAND U14245 ( .A(n6832), .B(n6823), .Z(n11873) );
  AND U14246 ( .A(n11875), .B(n11876), .Z(n11869) );
  AND U14247 ( .A(n11877), .B(n11878), .Z(n11876) );
  NAND U14248 ( .A(n6834), .B(n6827), .Z(n11878) );
  NAND U14249 ( .A(n6838), .B(n6833), .Z(n11877) );
  AND U14250 ( .A(n11879), .B(n11880), .Z(n11875) );
  NAND U14251 ( .A(n6850), .B(n6840), .Z(n11880) );
  NAND U14252 ( .A(n6835), .B(n6851), .Z(n11879) );
  AND U14253 ( .A(n11881), .B(n11882), .Z(n11855) );
  AND U14254 ( .A(n11883), .B(n11884), .Z(n11882) );
  AND U14255 ( .A(n11885), .B(n11886), .Z(n11884) );
  AND U14256 ( .A(n11887), .B(n11888), .Z(n11886) );
  NAND U14257 ( .A(n6852), .B(n6839), .Z(n11888) );
  NAND U14258 ( .A(n6856), .B(n6853), .Z(n11887) );
  AND U14259 ( .A(n11889), .B(n11890), .Z(n11885) );
  NAND U14260 ( .A(n6858), .B(n6841), .Z(n11890) );
  NAND U14261 ( .A(n6864), .B(n6857), .Z(n11889) );
  AND U14262 ( .A(n11891), .B(n11892), .Z(n11883) );
  AND U14263 ( .A(n11893), .B(n11894), .Z(n11892) );
  NAND U14264 ( .A(n6859), .B(n8487), .Z(n11894) );
  AND U14265 ( .A(n11895), .B(n11784), .Z(n11891) );
  NAND U14266 ( .A(n8603), .B(n6957), .Z(n11784) );
  AND U14267 ( .A(n11896), .B(n11897), .Z(n11881) );
  AND U14268 ( .A(n11898), .B(n11899), .Z(n11897) );
  AND U14269 ( .A(n11900), .B(n11901), .Z(n11899) );
  AND U14270 ( .A(n11902), .B(n8615), .Z(n11898) );
  NAND U14271 ( .A(n8958), .B(n6937), .Z(n8615) );
  AND U14272 ( .A(n11903), .B(n11904), .Z(n11896) );
  NAND U14273 ( .A(n6893), .B(n6926), .Z(n11904) );
  AND U14274 ( .A(n11905), .B(n9081), .Z(n11903) );
  NAND U14275 ( .A(n9135), .B(n6920), .Z(n9081) );
  NAND U14276 ( .A(n11906), .B(n6888), .Z(n11852) );
  NAND U14277 ( .A(n11907), .B(n11908), .Z(n11906) );
  AND U14278 ( .A(n11909), .B(n11910), .Z(n11908) );
  AND U14279 ( .A(n11911), .B(n11912), .Z(n11910) );
  AND U14280 ( .A(n11913), .B(n11914), .Z(n11912) );
  AND U14281 ( .A(n11915), .B(n11916), .Z(n11914) );
  NANDN U14282 ( .B(n8590), .A(n6919), .Z(n11916) );
  NAND U14283 ( .A(n6926), .B(n8512), .Z(n11915) );
  AND U14284 ( .A(n11917), .B(n11918), .Z(n11913) );
  NANDN U14285 ( .B(n8593), .A(n6920), .Z(n11918) );
  NANDN U14286 ( .B(n8516), .A(n6898), .Z(n11917) );
  AND U14287 ( .A(n11919), .B(n11920), .Z(n11911) );
  AND U14288 ( .A(n11921), .B(n11922), .Z(n11920) );
  NAND U14289 ( .A(n6925), .B(n6897), .Z(n11922) );
  NANDN U14290 ( .B(n8522), .A(n6882), .Z(n11921) );
  AND U14291 ( .A(n11923), .B(n11924), .Z(n11919) );
  NANDN U14292 ( .B(n8526), .A(n6809), .Z(n11924) );
  NANDN U14293 ( .B(n8534), .A(n6807), .Z(n11923) );
  AND U14294 ( .A(n11925), .B(n11926), .Z(n11909) );
  AND U14295 ( .A(n11927), .B(n11928), .Z(n11926) );
  AND U14296 ( .A(n11929), .B(n11930), .Z(n11928) );
  NANDN U14297 ( .B(n8511), .A(n6799), .Z(n11930) );
  NANDN U14298 ( .B(n8515), .A(n6803), .Z(n11929) );
  AND U14299 ( .A(n11931), .B(n11932), .Z(n11927) );
  NANDN U14300 ( .B(n8521), .A(n6823), .Z(n11932) );
  NANDN U14301 ( .B(n8525), .A(n6827), .Z(n11931) );
  AND U14302 ( .A(n11933), .B(n11934), .Z(n11925) );
  AND U14303 ( .A(n11935), .B(n11936), .Z(n11934) );
  NANDN U14304 ( .B(n8533), .A(n6833), .Z(n11936) );
  NANDN U14305 ( .B(n8537), .A(n6835), .Z(n11935) );
  AND U14306 ( .A(n11937), .B(n11938), .Z(n11933) );
  NANDN U14307 ( .B(n8538), .A(n6839), .Z(n11938) );
  NANDN U14308 ( .B(n8543), .A(n6850), .Z(n11937) );
  AND U14309 ( .A(n11939), .B(n11940), .Z(n11907) );
  AND U14310 ( .A(n11941), .B(n11942), .Z(n11940) );
  AND U14311 ( .A(n11943), .B(n11944), .Z(n11942) );
  AND U14312 ( .A(n11945), .B(n11946), .Z(n11944) );
  NANDN U14313 ( .B(n8544), .A(n6853), .Z(n11946) );
  NANDN U14314 ( .B(n8547), .A(n6841), .Z(n11945) );
  AND U14315 ( .A(n11947), .B(n11948), .Z(n11943) );
  NANDN U14316 ( .B(n8548), .A(n6857), .Z(n11948) );
  NANDN U14317 ( .B(n8557), .A(n6859), .Z(n11947) );
  AND U14318 ( .A(n11949), .B(n11950), .Z(n11941) );
  AND U14319 ( .A(n11951), .B(n11952), .Z(n11950) );
  NANDN U14320 ( .B(n8558), .A(n6865), .Z(n11952) );
  NANDN U14321 ( .B(n8561), .A(n6967), .Z(n11951) );
  AND U14322 ( .A(n11953), .B(n11954), .Z(n11949) );
  NANDN U14323 ( .B(n8562), .A(n6966), .Z(n11954) );
  NANDN U14324 ( .B(n8567), .A(n6961), .Z(n11953) );
  AND U14325 ( .A(n11955), .B(n11956), .Z(n11939) );
  AND U14326 ( .A(n11957), .B(n11958), .Z(n11956) );
  AND U14327 ( .A(n11959), .B(n11960), .Z(n11958) );
  NANDN U14328 ( .B(n8568), .A(n6956), .Z(n11960) );
  NANDN U14329 ( .B(n8571), .A(n6960), .Z(n11959) );
  AND U14330 ( .A(n11961), .B(n11962), .Z(n11957) );
  NANDN U14331 ( .B(n8572), .A(n6957), .Z(n11962) );
  NANDN U14332 ( .B(n8579), .A(n6947), .Z(n11961) );
  AND U14333 ( .A(n11963), .B(n11964), .Z(n11955) );
  AND U14334 ( .A(n11965), .B(n11966), .Z(n11964) );
  NANDN U14335 ( .B(n8580), .A(n6946), .Z(n11966) );
  NANDN U14336 ( .B(n8583), .A(n6943), .Z(n11965) );
  AND U14337 ( .A(n11967), .B(n11968), .Z(n11963) );
  NANDN U14338 ( .B(n8584), .A(n6942), .Z(n11968) );
  NANDN U14339 ( .B(n8589), .A(n6937), .Z(n11967) );
  NAND U14340 ( .A(n6765), .B(\u_a23_core/u_execute/u_alu/fadder_out[1] ), .Z(
        n11836) );
  OR U14341 ( .A(n11969), .B(n11843), .Z(n11833) );
  AND U14342 ( .A(n11970), .B(n11971), .Z(n11843) );
  AND U14343 ( .A(n11972), .B(n11973), .Z(n11971) );
  AND U14344 ( .A(n11974), .B(n11975), .Z(n11973) );
  AND U14345 ( .A(n11976), .B(n11977), .Z(n11975) );
  NANDN U14346 ( .B(n8636), .A(\u_a23_core/u_execute/u_register_bank/r14[1] ), 
        .Z(n11977) );
  NANDN U14347 ( .B(n8639), .A(\u_a23_core/u_execute/u_register_bank/r13[1] ), 
        .Z(n11976) );
  AND U14348 ( .A(n11978), .B(n11979), .Z(n11974) );
  NANDN U14349 ( .B(n8640), .A(\u_a23_core/u_execute/u_register_bank/r12[1] ), 
        .Z(n11979) );
  NANDN U14350 ( .B(n8645), .A(\u_a23_core/u_execute/u_register_bank/r11[1] ), 
        .Z(n11978) );
  AND U14351 ( .A(n11980), .B(n11981), .Z(n11972) );
  AND U14352 ( .A(n11982), .B(n11983), .Z(n11981) );
  NANDN U14353 ( .B(n8646), .A(\u_a23_core/u_execute/u_register_bank/r10[1] ), 
        .Z(n11983) );
  NANDN U14354 ( .B(n8649), .A(\u_a23_core/u_execute/u_register_bank/r9[1] ), 
        .Z(n11982) );
  AND U14355 ( .A(n11984), .B(n11985), .Z(n11980) );
  NANDN U14356 ( .B(n8650), .A(\u_a23_core/u_execute/u_register_bank/r8[1] ), 
        .Z(n11985) );
  NANDN U14357 ( .B(n8657), .A(\u_a23_core/u_execute/u_register_bank/r7[1] ), 
        .Z(n11984) );
  AND U14358 ( .A(n11986), .B(n11987), .Z(n11970) );
  AND U14359 ( .A(n11988), .B(n11989), .Z(n11987) );
  AND U14360 ( .A(n11990), .B(n11991), .Z(n11989) );
  NANDN U14361 ( .B(n8658), .A(\u_a23_core/u_execute/u_register_bank/r6[1] ), 
        .Z(n11991) );
  NANDN U14362 ( .B(n8661), .A(\u_a23_core/u_execute/u_register_bank/r5[1] ), 
        .Z(n11990) );
  AND U14363 ( .A(n11992), .B(n11993), .Z(n11988) );
  NANDN U14364 ( .B(n8662), .A(\u_a23_core/u_execute/u_register_bank/r4[1] ), 
        .Z(n11993) );
  NANDN U14365 ( .B(n8667), .A(\u_a23_core/u_execute/u_register_bank/r3[1] ), 
        .Z(n11992) );
  AND U14366 ( .A(n11994), .B(n11995), .Z(n11986) );
  NANDN U14367 ( .B(n8672), .A(\u_a23_core/u_execute/u_register_bank/r1[1] ), 
        .Z(n11995) );
  AND U14368 ( .A(n11996), .B(n11997), .Z(n11994) );
  NANDN U14369 ( .B(n8668), .A(\u_a23_core/u_execute/u_register_bank/r0[1] ), 
        .Z(n11997) );
  NANDN U14370 ( .B(n8671), .A(\u_a23_core/u_execute/u_register_bank/r2[1] ), 
        .Z(n11996) );
  NOR U14371 ( .A(\u_a23_core/execute_address_nxt[16] ), .B(
        \u_a23_core/execute_address_nxt[17] ), .Z(n11461) );
  NAND U14372 ( .A(n11998), .B(n11999), .Z(
        \u_a23_core/execute_address_nxt[17] ) );
  AND U14373 ( .A(n12000), .B(n12001), .Z(n11999) );
  AND U14374 ( .A(n12002), .B(n12003), .Z(n12001) );
  NANDN U14375 ( .B(n8392), .A(\u_a23_core/u_execute/pc_minus4[17] ), .Z(
        n12003) );
  NAND U14376 ( .A(n8393), .B(\u_a23_core/u_execute/alu_out_pc_filtered[17] ), 
        .Z(n12002) );
  IV U14377 ( .A(n7038), .Z(\u_a23_core/u_execute/alu_out_pc_filtered[17] ) );
  AND U14378 ( .A(n12004), .B(n12005), .Z(n7038) );
  MUX U14379 ( .IN0(n12006), .IN1(n12007), .SEL(
        \u_a23_core/u_execute/u_alu/b_not[17] ), .F(n12005) );
  NAND U14380 ( .A(n12008), .B(n12009), .Z(
        \u_a23_core/u_execute/u_alu/b_not[17] ) );
  MUX U14381 ( .IN0(n8430), .IN1(n8431), .SEL(n12010), .F(n12009) );
  MUX U14382 ( .IN0(n8433), .IN1(n8434), .SEL(\u_a23_core/u_execute/rn[17] ), 
        .F(n12008) );
  ANDN U14383 ( .A(n9256), .B(n12011), .Z(n12007) );
  MUX U14384 ( .IN0(n8400), .IN1(\u_a23_core/alu_function[3] ), .SEL(
        \u_a23_core/u_execute/u_alu/a[17] ), .F(n12011) );
  NAND U14385 ( .A(\u_a23_core/u_execute/u_alu/a[17] ), .B(n8400), .Z(n12006)
         );
  IV U14386 ( .A(n12012), .Z(\u_a23_core/u_execute/u_alu/a[17] ) );
  MUX U14387 ( .IN0(n12013), .IN1(n12010), .SEL(\u_a23_core/alu_function[8] ), 
        .F(n12012) );
  AND U14388 ( .A(n12014), .B(n12015), .Z(n12010) );
  AND U14389 ( .A(n12016), .B(n12017), .Z(n12015) );
  NAND U14390 ( .A(n6786), .B(n12018), .Z(n12017) );
  NAND U14391 ( .A(n12019), .B(n12020), .Z(n12018) );
  AND U14392 ( .A(n12021), .B(n12022), .Z(n12020) );
  AND U14393 ( .A(n12023), .B(n12024), .Z(n12022) );
  AND U14394 ( .A(n12025), .B(n12026), .Z(n12024) );
  NAND U14395 ( .A(n8461), .B(n6809), .Z(n12026) );
  NAND U14396 ( .A(n8470), .B(n6807), .Z(n12025) );
  AND U14397 ( .A(n12027), .B(n12028), .Z(n12023) );
  NAND U14398 ( .A(n9359), .B(n6799), .Z(n12028) );
  NAND U14399 ( .A(n9726), .B(n6803), .Z(n12027) );
  AND U14400 ( .A(n12029), .B(n12030), .Z(n12021) );
  NAND U14401 ( .A(n8609), .B(n6827), .Z(n12030) );
  AND U14402 ( .A(n12031), .B(n9386), .Z(n12029) );
  NAND U14403 ( .A(n8606), .B(n6833), .Z(n9386) );
  NAND U14404 ( .A(n8603), .B(n6823), .Z(n12031) );
  AND U14405 ( .A(n12032), .B(n12033), .Z(n12019) );
  AND U14406 ( .A(n12034), .B(n12035), .Z(n12033) );
  AND U14407 ( .A(n10123), .B(n9753), .Z(n12035) );
  NAND U14408 ( .A(n8610), .B(n6835), .Z(n9753) );
  NAND U14409 ( .A(n8616), .B(n6839), .Z(n10123) );
  AND U14410 ( .A(n10866), .B(n10485), .Z(n12034) );
  NAND U14411 ( .A(n6850), .B(n8958), .Z(n10485) );
  NAND U14412 ( .A(n9082), .B(n6853), .Z(n10866) );
  AND U14413 ( .A(n12036), .B(n12037), .Z(n12032) );
  NAND U14414 ( .A(n6893), .B(n6859), .Z(n12037) );
  AND U14415 ( .A(n11790), .B(n11230), .Z(n12036) );
  NAND U14416 ( .A(n9135), .B(n6841), .Z(n11230) );
  NAND U14417 ( .A(n6984), .B(n6857), .Z(n11790) );
  AND U14418 ( .A(n12038), .B(n12039), .Z(n12016) );
  NANDN U14419 ( .B(n11310), .A(n6886), .Z(n12039) );
  ANDN U14420 ( .A(n12040), .B(n8465), .Z(n11310) );
  NAND U14421 ( .A(n8465), .B(n6985), .Z(n12038) );
  AND U14422 ( .A(n12041), .B(n12042), .Z(n12014) );
  NAND U14423 ( .A(n12043), .B(n6888), .Z(n12042) );
  NAND U14424 ( .A(n12044), .B(n12045), .Z(n12043) );
  AND U14425 ( .A(n12046), .B(n12047), .Z(n12045) );
  AND U14426 ( .A(n12048), .B(n12049), .Z(n12047) );
  AND U14427 ( .A(n12050), .B(n12051), .Z(n12049) );
  AND U14428 ( .A(n12052), .B(n12053), .Z(n12051) );
  NANDN U14429 ( .B(n8544), .A(n6919), .Z(n12053) );
  NAND U14430 ( .A(n6859), .B(n8512), .Z(n12052) );
  AND U14431 ( .A(n12054), .B(n12055), .Z(n12050) );
  NANDN U14432 ( .B(n8547), .A(n6920), .Z(n12055) );
  NANDN U14433 ( .B(n8516), .A(n6865), .Z(n12054) );
  AND U14434 ( .A(n12056), .B(n12057), .Z(n12048) );
  AND U14435 ( .A(n12058), .B(n12059), .Z(n12057) );
  NANDN U14436 ( .B(n8548), .A(n6925), .Z(n12059) );
  NANDN U14437 ( .B(n8522), .A(n6967), .Z(n12058) );
  AND U14438 ( .A(n12060), .B(n12061), .Z(n12056) );
  NANDN U14439 ( .B(n8557), .A(n6926), .Z(n12061) );
  NANDN U14440 ( .B(n8526), .A(n6966), .Z(n12060) );
  AND U14441 ( .A(n12062), .B(n12063), .Z(n12046) );
  AND U14442 ( .A(n12064), .B(n12065), .Z(n12063) );
  AND U14443 ( .A(n12066), .B(n12067), .Z(n12065) );
  NANDN U14444 ( .B(n8558), .A(n6898), .Z(n12067) );
  NANDN U14445 ( .B(n8534), .A(n6961), .Z(n12066) );
  AND U14446 ( .A(n12068), .B(n12069), .Z(n12064) );
  NANDN U14447 ( .B(n8511), .A(n6956), .Z(n12069) );
  NANDN U14448 ( .B(n8561), .A(n6882), .Z(n12068) );
  AND U14449 ( .A(n12070), .B(n12071), .Z(n12062) );
  AND U14450 ( .A(n12072), .B(n12073), .Z(n12071) );
  NANDN U14451 ( .B(n8515), .A(n6960), .Z(n12073) );
  NANDN U14452 ( .B(n8562), .A(n6809), .Z(n12072) );
  AND U14453 ( .A(n12074), .B(n12075), .Z(n12070) );
  NANDN U14454 ( .B(n8521), .A(n6957), .Z(n12075) );
  NANDN U14455 ( .B(n8567), .A(n6807), .Z(n12074) );
  AND U14456 ( .A(n12076), .B(n12077), .Z(n12044) );
  AND U14457 ( .A(n12078), .B(n12079), .Z(n12077) );
  AND U14458 ( .A(n12080), .B(n12081), .Z(n12079) );
  AND U14459 ( .A(n12082), .B(n12083), .Z(n12081) );
  NANDN U14460 ( .B(n8525), .A(n6947), .Z(n12083) );
  NANDN U14461 ( .B(n8568), .A(n6799), .Z(n12082) );
  AND U14462 ( .A(n12084), .B(n12085), .Z(n12080) );
  NANDN U14463 ( .B(n8571), .A(n6803), .Z(n12085) );
  NANDN U14464 ( .B(n8533), .A(n6946), .Z(n12084) );
  AND U14465 ( .A(n12086), .B(n12087), .Z(n12078) );
  AND U14466 ( .A(n12088), .B(n12089), .Z(n12087) );
  NANDN U14467 ( .B(n8572), .A(n6823), .Z(n12089) );
  NANDN U14468 ( .B(n8537), .A(n6943), .Z(n12088) );
  AND U14469 ( .A(n12090), .B(n12091), .Z(n12086) );
  NANDN U14470 ( .B(n8579), .A(n6827), .Z(n12091) );
  NANDN U14471 ( .B(n8538), .A(n6942), .Z(n12090) );
  AND U14472 ( .A(n12092), .B(n12093), .Z(n12076) );
  AND U14473 ( .A(n12094), .B(n12095), .Z(n12093) );
  AND U14474 ( .A(n12096), .B(n12097), .Z(n12095) );
  NANDN U14475 ( .B(n8580), .A(n6833), .Z(n12097) );
  NANDN U14476 ( .B(n8543), .A(n6937), .Z(n12096) );
  AND U14477 ( .A(n12098), .B(n12099), .Z(n12094) );
  NANDN U14478 ( .B(n8583), .A(n6835), .Z(n12099) );
  NANDN U14479 ( .B(n8584), .A(n6839), .Z(n12098) );
  AND U14480 ( .A(n12100), .B(n12101), .Z(n12092) );
  AND U14481 ( .A(n12102), .B(n12103), .Z(n12101) );
  NANDN U14482 ( .B(n8589), .A(n6850), .Z(n12103) );
  NANDN U14483 ( .B(n8590), .A(n6853), .Z(n12102) );
  AND U14484 ( .A(n12104), .B(n12105), .Z(n12100) );
  NANDN U14485 ( .B(n8593), .A(n6841), .Z(n12105) );
  NAND U14486 ( .A(n6857), .B(n6897), .Z(n12104) );
  NAND U14487 ( .A(n12106), .B(n6902), .Z(n12041) );
  NAND U14488 ( .A(n12107), .B(n12108), .Z(n12106) );
  AND U14489 ( .A(n12109), .B(n12110), .Z(n12108) );
  AND U14490 ( .A(n12111), .B(n12112), .Z(n12110) );
  AND U14491 ( .A(n12113), .B(n12114), .Z(n12112) );
  NAND U14492 ( .A(n8465), .B(n6920), .Z(n12114) );
  AND U14493 ( .A(n12115), .B(n12116), .Z(n12113) );
  NAND U14494 ( .A(n6916), .B(n6859), .Z(n12116) );
  NAND U14495 ( .A(n8464), .B(n6925), .Z(n12115) );
  AND U14496 ( .A(n12117), .B(n12118), .Z(n12111) );
  NAND U14497 ( .A(n8461), .B(n6919), .Z(n12118) );
  NAND U14498 ( .A(n8470), .B(n6937), .Z(n12117) );
  AND U14499 ( .A(n12119), .B(n12120), .Z(n12109) );
  AND U14500 ( .A(n12121), .B(n12122), .Z(n12120) );
  NAND U14501 ( .A(n9359), .B(n6942), .Z(n12122) );
  NAND U14502 ( .A(n9726), .B(n6943), .Z(n12121) );
  AND U14503 ( .A(n12123), .B(n12124), .Z(n12119) );
  NAND U14504 ( .A(n6864), .B(n6898), .Z(n12124) );
  NAND U14505 ( .A(n6926), .B(n8487), .Z(n12123) );
  AND U14506 ( .A(n12125), .B(n12126), .Z(n12107) );
  AND U14507 ( .A(n12127), .B(n12128), .Z(n12126) );
  AND U14508 ( .A(n12129), .B(n11895), .Z(n12128) );
  NAND U14509 ( .A(n8609), .B(n6947), .Z(n11895) );
  AND U14510 ( .A(n6866), .B(n12130), .Z(n12129) );
  NAND U14511 ( .A(n8603), .B(n6946), .Z(n6866) );
  AND U14512 ( .A(n12131), .B(n9123), .Z(n12127) );
  NAND U14513 ( .A(n8610), .B(n6960), .Z(n9123) );
  AND U14514 ( .A(n12132), .B(n12133), .Z(n12125) );
  AND U14515 ( .A(n12134), .B(n8497), .Z(n12133) );
  NAND U14516 ( .A(n6961), .B(n8958), .Z(n8497) );
  AND U14517 ( .A(n12135), .B(n12136), .Z(n12132) );
  IV U14518 ( .A(\u_a23_core/u_execute/rn[17] ), .Z(n12013) );
  AND U14519 ( .A(n9395), .B(n12137), .Z(n12004) );
  NAND U14520 ( .A(n6765), .B(\u_a23_core/u_execute/u_alu/fadder_out[17] ), 
        .Z(n12137) );
  AND U14521 ( .A(n12138), .B(n12139), .Z(n12000) );
  NANDN U14522 ( .B(n8406), .A(\u_a23_core/u_execute/rn_plus4[17] ), .Z(n12139) );
  NANDN U14523 ( .B(n8407), .A(\u_a23_core/u_execute/alu_plus4[17] ), .Z(
        n12138) );
  AND U14524 ( .A(n12140), .B(n12141), .Z(n11998) );
  AND U14525 ( .A(n12142), .B(n12143), .Z(n12141) );
  NAND U14526 ( .A(n8412), .B(\u_a23_core/u_execute/address_plus4[17] ), .Z(
        n12143) );
  NAND U14527 ( .A(\u_a23_core/u_execute/rn[17] ), .B(n8413), .Z(n12142) );
  NAND U14528 ( .A(n12144), .B(n12145), .Z(\u_a23_core/u_execute/rn[17] ) );
  AND U14529 ( .A(n12146), .B(n12147), .Z(n12145) );
  AND U14530 ( .A(n12148), .B(n12149), .Z(n12147) );
  AND U14531 ( .A(n12150), .B(n12151), .Z(n12149) );
  NANDN U14532 ( .B(n8635), .A(\u_a23_core/u_execute/pc[17] ), .Z(n12151) );
  NANDN U14533 ( .B(n8636), .A(\u_a23_core/u_execute/u_register_bank/r14[17] ), 
        .Z(n12150) );
  AND U14534 ( .A(n12152), .B(n12153), .Z(n12148) );
  NANDN U14535 ( .B(n8639), .A(\u_a23_core/u_execute/u_register_bank/r13[17] ), 
        .Z(n12153) );
  NANDN U14536 ( .B(n8640), .A(\u_a23_core/u_execute/u_register_bank/r12[17] ), 
        .Z(n12152) );
  AND U14537 ( .A(n12154), .B(n12155), .Z(n12146) );
  AND U14538 ( .A(n12156), .B(n12157), .Z(n12155) );
  NANDN U14539 ( .B(n8645), .A(\u_a23_core/u_execute/u_register_bank/r11[17] ), 
        .Z(n12157) );
  NANDN U14540 ( .B(n8646), .A(\u_a23_core/u_execute/u_register_bank/r10[17] ), 
        .Z(n12156) );
  AND U14541 ( .A(n12158), .B(n12159), .Z(n12154) );
  NANDN U14542 ( .B(n8649), .A(\u_a23_core/u_execute/u_register_bank/r9[17] ), 
        .Z(n12159) );
  NANDN U14543 ( .B(n8650), .A(\u_a23_core/u_execute/u_register_bank/r8[17] ), 
        .Z(n12158) );
  AND U14544 ( .A(n12160), .B(n12161), .Z(n12144) );
  AND U14545 ( .A(n12162), .B(n12163), .Z(n12161) );
  AND U14546 ( .A(n12164), .B(n12165), .Z(n12163) );
  NANDN U14547 ( .B(n8657), .A(\u_a23_core/u_execute/u_register_bank/r7[17] ), 
        .Z(n12165) );
  NANDN U14548 ( .B(n8658), .A(\u_a23_core/u_execute/u_register_bank/r6[17] ), 
        .Z(n12164) );
  AND U14549 ( .A(n12166), .B(n12167), .Z(n12162) );
  NANDN U14550 ( .B(n8661), .A(\u_a23_core/u_execute/u_register_bank/r5[17] ), 
        .Z(n12167) );
  NANDN U14551 ( .B(n8662), .A(\u_a23_core/u_execute/u_register_bank/r4[17] ), 
        .Z(n12166) );
  AND U14552 ( .A(n12168), .B(n12169), .Z(n12160) );
  AND U14553 ( .A(n12170), .B(n12171), .Z(n12169) );
  NANDN U14554 ( .B(n8667), .A(\u_a23_core/u_execute/u_register_bank/r3[17] ), 
        .Z(n12171) );
  NANDN U14555 ( .B(n8668), .A(\u_a23_core/u_execute/u_register_bank/r0[17] ), 
        .Z(n12170) );
  AND U14556 ( .A(n12172), .B(n12173), .Z(n12168) );
  NANDN U14557 ( .B(n8671), .A(\u_a23_core/u_execute/u_register_bank/r2[17] ), 
        .Z(n12173) );
  NANDN U14558 ( .B(n8672), .A(\u_a23_core/u_execute/u_register_bank/r1[17] ), 
        .Z(n12172) );
  AND U14559 ( .A(n12174), .B(n12175), .Z(n12140) );
  NAND U14560 ( .A(\u_a23_core/u_execute/pc[17] ), .B(n8416), .Z(n12175) );
  NAND U14561 ( .A(n8417), .B(\u_a23_core/u_execute/pc_plus4[17] ), .Z(n12174)
         );
  NAND U14562 ( .A(n12176), .B(n12177), .Z(
        \u_a23_core/execute_address_nxt[16] ) );
  AND U14563 ( .A(n12178), .B(n12179), .Z(n12177) );
  AND U14564 ( .A(n12180), .B(n12181), .Z(n12179) );
  NANDN U14565 ( .B(n8392), .A(\u_a23_core/u_execute/pc_minus4[16] ), .Z(
        n12181) );
  NAND U14566 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[16] ), .B(n8393), 
        .Z(n12180) );
  IV U14567 ( .A(n7039), .Z(\u_a23_core/u_execute/alu_out_pc_filtered[16] ) );
  AND U14568 ( .A(n12182), .B(n12183), .Z(n7039) );
  MUX U14569 ( .IN0(n12184), .IN1(n12185), .SEL(
        \u_a23_core/u_execute/u_alu/b_not[16] ), .F(n12183) );
  NAND U14570 ( .A(n12186), .B(n12187), .Z(
        \u_a23_core/u_execute/u_alu/b_not[16] ) );
  MUX U14571 ( .IN0(n8430), .IN1(n8431), .SEL(n12188), .F(n12187) );
  MUX U14572 ( .IN0(n8433), .IN1(n8434), .SEL(\u_a23_core/u_execute/rn[16] ), 
        .F(n12186) );
  ANDN U14573 ( .A(n9256), .B(n12189), .Z(n12185) );
  MUX U14574 ( .IN0(n8400), .IN1(\u_a23_core/alu_function[3] ), .SEL(
        \u_a23_core/u_execute/u_alu/a[16] ), .F(n12189) );
  NAND U14575 ( .A(\u_a23_core/u_execute/u_alu/a[16] ), .B(n8400), .Z(n12184)
         );
  IV U14576 ( .A(n12190), .Z(\u_a23_core/u_execute/u_alu/a[16] ) );
  MUX U14577 ( .IN0(n12191), .IN1(n12188), .SEL(\u_a23_core/alu_function[8] ), 
        .F(n12190) );
  AND U14578 ( .A(n12192), .B(n12193), .Z(n12188) );
  AND U14579 ( .A(n12194), .B(n12195), .Z(n12193) );
  NAND U14580 ( .A(n6786), .B(n12196), .Z(n12195) );
  NAND U14581 ( .A(n12197), .B(n12198), .Z(n12196) );
  AND U14582 ( .A(n12199), .B(n12200), .Z(n12198) );
  AND U14583 ( .A(n12201), .B(n12202), .Z(n12200) );
  AND U14584 ( .A(n12203), .B(n12204), .Z(n12202) );
  NAND U14585 ( .A(n8465), .B(n6809), .Z(n12204) );
  NAND U14586 ( .A(n8461), .B(n6807), .Z(n12203) );
  AND U14587 ( .A(n12205), .B(n12206), .Z(n12201) );
  NAND U14588 ( .A(n8470), .B(n6799), .Z(n12206) );
  NAND U14589 ( .A(n9359), .B(n6803), .Z(n12205) );
  AND U14590 ( .A(n12207), .B(n12208), .Z(n12199) );
  AND U14591 ( .A(n9494), .B(n12209), .Z(n12208) );
  NAND U14592 ( .A(n9726), .B(n6823), .Z(n12209) );
  NAND U14593 ( .A(n8606), .B(n6835), .Z(n9494) );
  AND U14594 ( .A(n6974), .B(n12210), .Z(n12207) );
  NAND U14595 ( .A(n8603), .B(n6827), .Z(n12210) );
  NAND U14596 ( .A(n8609), .B(n6833), .Z(n6974) );
  AND U14597 ( .A(n12211), .B(n12212), .Z(n12197) );
  AND U14598 ( .A(n12213), .B(n12214), .Z(n12212) );
  AND U14599 ( .A(n10305), .B(n9938), .Z(n12214) );
  NAND U14600 ( .A(n8610), .B(n6839), .Z(n9938) );
  NAND U14601 ( .A(n6850), .B(n8616), .Z(n10305) );
  AND U14602 ( .A(n11045), .B(n10671), .Z(n12213) );
  NAND U14603 ( .A(n8958), .B(n6853), .Z(n10671) );
  NAND U14604 ( .A(n9082), .B(n6841), .Z(n11045) );
  AND U14605 ( .A(n12215), .B(n12216), .Z(n12211) );
  NAND U14606 ( .A(n6865), .B(n6893), .Z(n12216) );
  AND U14607 ( .A(n11604), .B(n11417), .Z(n12215) );
  NAND U14608 ( .A(n9135), .B(n6857), .Z(n11417) );
  NAND U14609 ( .A(n6984), .B(n6859), .Z(n11604) );
  AND U14610 ( .A(n12217), .B(n12218), .Z(n12194) );
  NANDN U14611 ( .B(n12040), .A(n6886), .Z(n12218) );
  AND U14612 ( .A(n12219), .B(n11690), .Z(n12040) );
  AND U14613 ( .A(n12220), .B(n11689), .Z(n12219) );
  IV U14614 ( .A(n8464), .Z(n11689) );
  NAND U14615 ( .A(n8464), .B(n6985), .Z(n12217) );
  AND U14616 ( .A(n12221), .B(n12222), .Z(n12192) );
  NAND U14617 ( .A(n12223), .B(n6888), .Z(n12222) );
  NAND U14618 ( .A(n12224), .B(n12225), .Z(n12223) );
  AND U14619 ( .A(n12226), .B(n12227), .Z(n12225) );
  AND U14620 ( .A(n12228), .B(n12229), .Z(n12227) );
  AND U14621 ( .A(n12230), .B(n12231), .Z(n12229) );
  AND U14622 ( .A(n12232), .B(n12233), .Z(n12231) );
  NANDN U14623 ( .B(n8543), .A(n6919), .Z(n12233) );
  NAND U14624 ( .A(n6865), .B(n8512), .Z(n12232) );
  AND U14625 ( .A(n12234), .B(n12235), .Z(n12230) );
  NANDN U14626 ( .B(n8544), .A(n6920), .Z(n12235) );
  NANDN U14627 ( .B(n8516), .A(n6967), .Z(n12234) );
  AND U14628 ( .A(n12236), .B(n12237), .Z(n12228) );
  AND U14629 ( .A(n12238), .B(n12239), .Z(n12237) );
  NANDN U14630 ( .B(n8547), .A(n6925), .Z(n12239) );
  NANDN U14631 ( .B(n8522), .A(n6966), .Z(n12238) );
  AND U14632 ( .A(n12240), .B(n12241), .Z(n12236) );
  NANDN U14633 ( .B(n8548), .A(n6926), .Z(n12241) );
  NANDN U14634 ( .B(n8526), .A(n6961), .Z(n12240) );
  AND U14635 ( .A(n12242), .B(n12243), .Z(n12226) );
  AND U14636 ( .A(n12244), .B(n12245), .Z(n12243) );
  AND U14637 ( .A(n12246), .B(n12247), .Z(n12245) );
  NANDN U14638 ( .B(n8557), .A(n6898), .Z(n12247) );
  NANDN U14639 ( .B(n8534), .A(n6956), .Z(n12246) );
  AND U14640 ( .A(n12248), .B(n12249), .Z(n12244) );
  NANDN U14641 ( .B(n8511), .A(n6960), .Z(n12249) );
  NANDN U14642 ( .B(n8558), .A(n6882), .Z(n12248) );
  AND U14643 ( .A(n12250), .B(n12251), .Z(n12242) );
  AND U14644 ( .A(n12252), .B(n12253), .Z(n12251) );
  NANDN U14645 ( .B(n8515), .A(n6957), .Z(n12253) );
  NANDN U14646 ( .B(n8561), .A(n6809), .Z(n12252) );
  AND U14647 ( .A(n12254), .B(n12255), .Z(n12250) );
  NANDN U14648 ( .B(n8521), .A(n6947), .Z(n12255) );
  NANDN U14649 ( .B(n8562), .A(n6807), .Z(n12254) );
  AND U14650 ( .A(n12256), .B(n12257), .Z(n12224) );
  AND U14651 ( .A(n12258), .B(n12259), .Z(n12257) );
  AND U14652 ( .A(n12260), .B(n12261), .Z(n12259) );
  AND U14653 ( .A(n12262), .B(n12263), .Z(n12261) );
  NANDN U14654 ( .B(n8525), .A(n6946), .Z(n12263) );
  NANDN U14655 ( .B(n8567), .A(n6799), .Z(n12262) );
  AND U14656 ( .A(n12264), .B(n12265), .Z(n12260) );
  NANDN U14657 ( .B(n8568), .A(n6803), .Z(n12265) );
  NANDN U14658 ( .B(n8533), .A(n6943), .Z(n12264) );
  AND U14659 ( .A(n12266), .B(n12267), .Z(n12258) );
  AND U14660 ( .A(n12268), .B(n12269), .Z(n12267) );
  NANDN U14661 ( .B(n8571), .A(n6823), .Z(n12269) );
  NANDN U14662 ( .B(n8537), .A(n6942), .Z(n12268) );
  AND U14663 ( .A(n12270), .B(n12271), .Z(n12266) );
  NANDN U14664 ( .B(n8572), .A(n6827), .Z(n12271) );
  NANDN U14665 ( .B(n8538), .A(n6937), .Z(n12270) );
  AND U14666 ( .A(n12272), .B(n12273), .Z(n12256) );
  AND U14667 ( .A(n12274), .B(n12275), .Z(n12273) );
  AND U14668 ( .A(n12276), .B(n12277), .Z(n12275) );
  NANDN U14669 ( .B(n8579), .A(n6833), .Z(n12277) );
  NANDN U14670 ( .B(n8580), .A(n6835), .Z(n12276) );
  AND U14671 ( .A(n12278), .B(n12279), .Z(n12274) );
  NANDN U14672 ( .B(n8583), .A(n6839), .Z(n12279) );
  NANDN U14673 ( .B(n8584), .A(n6850), .Z(n12278) );
  AND U14674 ( .A(n12280), .B(n12281), .Z(n12272) );
  AND U14675 ( .A(n12282), .B(n12283), .Z(n12281) );
  NANDN U14676 ( .B(n8589), .A(n6853), .Z(n12283) );
  NANDN U14677 ( .B(n8590), .A(n6841), .Z(n12282) );
  AND U14678 ( .A(n12284), .B(n12285), .Z(n12280) );
  NANDN U14679 ( .B(n8593), .A(n6857), .Z(n12285) );
  NAND U14680 ( .A(n6859), .B(n6897), .Z(n12284) );
  NAND U14681 ( .A(n12286), .B(n6902), .Z(n12221) );
  NAND U14682 ( .A(n12287), .B(n12288), .Z(n12286) );
  AND U14683 ( .A(n12289), .B(n12290), .Z(n12288) );
  AND U14684 ( .A(n12291), .B(n12292), .Z(n12290) );
  AND U14685 ( .A(n12293), .B(n12294), .Z(n12292) );
  NAND U14686 ( .A(n8465), .B(n6925), .Z(n12294) );
  AND U14687 ( .A(n12295), .B(n12296), .Z(n12293) );
  NAND U14688 ( .A(n6865), .B(n6916), .Z(n12296) );
  NAND U14689 ( .A(n8464), .B(n6926), .Z(n12295) );
  AND U14690 ( .A(n12297), .B(n12298), .Z(n12291) );
  NAND U14691 ( .A(n8461), .B(n6920), .Z(n12298) );
  NAND U14692 ( .A(n8470), .B(n6919), .Z(n12297) );
  AND U14693 ( .A(n12299), .B(n12300), .Z(n12289) );
  AND U14694 ( .A(n12301), .B(n12302), .Z(n12300) );
  NAND U14695 ( .A(n9359), .B(n6937), .Z(n12302) );
  NAND U14696 ( .A(n9726), .B(n6942), .Z(n12301) );
  AND U14697 ( .A(n12303), .B(n12304), .Z(n12299) );
  NAND U14698 ( .A(n6898), .B(n8487), .Z(n12304) );
  AND U14699 ( .A(n12305), .B(n12306), .Z(n12287) );
  AND U14700 ( .A(n12307), .B(n12308), .Z(n12306) );
  AND U14701 ( .A(n12309), .B(n12310), .Z(n12308) );
  NAND U14702 ( .A(n8603), .B(n6943), .Z(n12310) );
  AND U14703 ( .A(n9008), .B(n12311), .Z(n12307) );
  NAND U14704 ( .A(n8616), .B(n6960), .Z(n9008) );
  AND U14705 ( .A(n12312), .B(n12313), .Z(n12305) );
  AND U14706 ( .A(n12314), .B(n8737), .Z(n12313) );
  NAND U14707 ( .A(n6956), .B(n8958), .Z(n8737) );
  AND U14708 ( .A(n12315), .B(n12316), .Z(n12312) );
  IV U14709 ( .A(\u_a23_core/u_execute/rn[16] ), .Z(n12191) );
  AND U14710 ( .A(n9395), .B(n12317), .Z(n12182) );
  NAND U14711 ( .A(n6765), .B(\u_a23_core/u_execute/u_alu/fadder_out[16] ), 
        .Z(n12317) );
  ANDN U14712 ( .A(n12318), .B(n12319), .Z(n9395) );
  NAND U14713 ( .A(n12320), .B(\u_a23_core/u_execute/u_alu/b_not[15] ), .Z(
        n12318) );
  AND U14714 ( .A(n12321), .B(n12322), .Z(n12178) );
  NANDN U14715 ( .B(n8406), .A(\u_a23_core/u_execute/rn_plus4[16] ), .Z(n12322) );
  NANDN U14716 ( .B(n8407), .A(\u_a23_core/u_execute/alu_plus4[16] ), .Z(
        n12321) );
  AND U14717 ( .A(n12323), .B(n12324), .Z(n12176) );
  AND U14718 ( .A(n12325), .B(n12326), .Z(n12324) );
  NAND U14719 ( .A(n8412), .B(\u_a23_core/u_execute/address_plus4[16] ), .Z(
        n12326) );
  NAND U14720 ( .A(\u_a23_core/u_execute/rn[16] ), .B(n8413), .Z(n12325) );
  NAND U14721 ( .A(n12327), .B(n12328), .Z(\u_a23_core/u_execute/rn[16] ) );
  AND U14722 ( .A(n12329), .B(n12330), .Z(n12328) );
  AND U14723 ( .A(n12331), .B(n12332), .Z(n12330) );
  AND U14724 ( .A(n12333), .B(n12334), .Z(n12332) );
  NANDN U14725 ( .B(n8635), .A(\u_a23_core/u_execute/pc[16] ), .Z(n12334) );
  NANDN U14726 ( .B(n8636), .A(\u_a23_core/u_execute/u_register_bank/r14[16] ), 
        .Z(n12333) );
  AND U14727 ( .A(n12335), .B(n12336), .Z(n12331) );
  NANDN U14728 ( .B(n8639), .A(\u_a23_core/u_execute/u_register_bank/r13[16] ), 
        .Z(n12336) );
  NANDN U14729 ( .B(n8640), .A(\u_a23_core/u_execute/u_register_bank/r12[16] ), 
        .Z(n12335) );
  AND U14730 ( .A(n12337), .B(n12338), .Z(n12329) );
  AND U14731 ( .A(n12339), .B(n12340), .Z(n12338) );
  NANDN U14732 ( .B(n8645), .A(\u_a23_core/u_execute/u_register_bank/r11[16] ), 
        .Z(n12340) );
  NANDN U14733 ( .B(n8646), .A(\u_a23_core/u_execute/u_register_bank/r10[16] ), 
        .Z(n12339) );
  AND U14734 ( .A(n12341), .B(n12342), .Z(n12337) );
  NANDN U14735 ( .B(n8649), .A(\u_a23_core/u_execute/u_register_bank/r9[16] ), 
        .Z(n12342) );
  NANDN U14736 ( .B(n8650), .A(\u_a23_core/u_execute/u_register_bank/r8[16] ), 
        .Z(n12341) );
  AND U14737 ( .A(n12343), .B(n12344), .Z(n12327) );
  AND U14738 ( .A(n12345), .B(n12346), .Z(n12344) );
  AND U14739 ( .A(n12347), .B(n12348), .Z(n12346) );
  NANDN U14740 ( .B(n8657), .A(\u_a23_core/u_execute/u_register_bank/r7[16] ), 
        .Z(n12348) );
  NANDN U14741 ( .B(n8658), .A(\u_a23_core/u_execute/u_register_bank/r6[16] ), 
        .Z(n12347) );
  AND U14742 ( .A(n12349), .B(n12350), .Z(n12345) );
  NANDN U14743 ( .B(n8661), .A(\u_a23_core/u_execute/u_register_bank/r5[16] ), 
        .Z(n12350) );
  NANDN U14744 ( .B(n8662), .A(\u_a23_core/u_execute/u_register_bank/r4[16] ), 
        .Z(n12349) );
  AND U14745 ( .A(n12351), .B(n12352), .Z(n12343) );
  AND U14746 ( .A(n12353), .B(n12354), .Z(n12352) );
  NANDN U14747 ( .B(n8667), .A(\u_a23_core/u_execute/u_register_bank/r3[16] ), 
        .Z(n12354) );
  NANDN U14748 ( .B(n8668), .A(\u_a23_core/u_execute/u_register_bank/r0[16] ), 
        .Z(n12353) );
  AND U14749 ( .A(n12355), .B(n12356), .Z(n12351) );
  NANDN U14750 ( .B(n8671), .A(\u_a23_core/u_execute/u_register_bank/r2[16] ), 
        .Z(n12356) );
  NANDN U14751 ( .B(n8672), .A(\u_a23_core/u_execute/u_register_bank/r1[16] ), 
        .Z(n12355) );
  AND U14752 ( .A(n12357), .B(n12358), .Z(n12323) );
  NAND U14753 ( .A(\u_a23_core/u_execute/pc[16] ), .B(n8416), .Z(n12358) );
  NAND U14754 ( .A(n8417), .B(\u_a23_core/u_execute/pc_plus4[16] ), .Z(n12357)
         );
  AND U14755 ( .A(n12359), .B(n12360), .Z(n11459) );
  NOR U14756 ( .A(\u_a23_core/execute_address_nxt[14] ), .B(
        \u_a23_core/execute_address_nxt[15] ), .Z(n12360) );
  NAND U14757 ( .A(n12361), .B(n12362), .Z(
        \u_a23_core/execute_address_nxt[15] ) );
  AND U14758 ( .A(n12363), .B(n12364), .Z(n12362) );
  AND U14759 ( .A(n12365), .B(n12366), .Z(n12364) );
  NANDN U14760 ( .B(n8392), .A(\u_a23_core/u_execute/pc_minus4[15] ), .Z(
        n12366) );
  NAND U14761 ( .A(n8393), .B(\u_a23_core/u_execute/alu_out_pc_filtered[15] ), 
        .Z(n12365) );
  IV U14762 ( .A(n7040), .Z(\u_a23_core/u_execute/alu_out_pc_filtered[15] ) );
  AND U14763 ( .A(n12367), .B(n12368), .Z(n7040) );
  MUX U14764 ( .IN0(n12369), .IN1(n12370), .SEL(
        \u_a23_core/u_execute/u_alu/b_not[15] ), .F(n12368) );
  NAND U14765 ( .A(n12371), .B(n12372), .Z(
        \u_a23_core/u_execute/u_alu/b_not[15] ) );
  MUX U14766 ( .IN0(n8430), .IN1(n8431), .SEL(n12373), .F(n12372) );
  MUX U14767 ( .IN0(n8433), .IN1(n8434), .SEL(\u_a23_core/u_execute/rn[15] ), 
        .F(n12371) );
  ANDN U14768 ( .A(n8435), .B(n12374), .Z(n12370) );
  MUX U14769 ( .IN0(n8400), .IN1(\u_a23_core/alu_function[3] ), .SEL(
        \u_a23_core/u_execute/u_alu/a[15] ), .F(n12374) );
  NAND U14770 ( .A(\u_a23_core/u_execute/u_alu/a[15] ), .B(n8400), .Z(n12369)
         );
  IV U14771 ( .A(n12375), .Z(\u_a23_core/u_execute/u_alu/a[15] ) );
  MUX U14772 ( .IN0(n12376), .IN1(n12373), .SEL(\u_a23_core/alu_function[8] ), 
        .F(n12375) );
  AND U14773 ( .A(n12377), .B(n12378), .Z(n12373) );
  AND U14774 ( .A(n12379), .B(n12380), .Z(n12378) );
  NAND U14775 ( .A(n8443), .B(n12381), .Z(n12380) );
  AND U14776 ( .A(n12382), .B(n6882), .Z(n12381) );
  NAND U14777 ( .A(n12220), .B(n11690), .Z(n12382) );
  NOR U14778 ( .A(n8487), .B(n12383), .Z(n11690) );
  AND U14779 ( .A(n12384), .B(n12385), .Z(n12379) );
  NAND U14780 ( .A(n6985), .B(n8487), .Z(n12385) );
  NAND U14781 ( .A(n6786), .B(n12386), .Z(n12384) );
  NAND U14782 ( .A(n12387), .B(n12388), .Z(n12386) );
  AND U14783 ( .A(n12389), .B(n12390), .Z(n12388) );
  AND U14784 ( .A(n12391), .B(n12392), .Z(n12390) );
  AND U14785 ( .A(n12393), .B(n12394), .Z(n12392) );
  NAND U14786 ( .A(n8464), .B(n6809), .Z(n12394) );
  NAND U14787 ( .A(n8465), .B(n6807), .Z(n12393) );
  AND U14788 ( .A(n12395), .B(n12396), .Z(n12391) );
  NAND U14789 ( .A(n8461), .B(n6799), .Z(n12396) );
  NAND U14790 ( .A(n8470), .B(n6803), .Z(n12395) );
  AND U14791 ( .A(n12397), .B(n12398), .Z(n12389) );
  AND U14792 ( .A(n12399), .B(n12400), .Z(n12398) );
  NAND U14793 ( .A(n9359), .B(n6823), .Z(n12400) );
  NAND U14794 ( .A(n9726), .B(n6827), .Z(n12399) );
  AND U14795 ( .A(n12401), .B(n9748), .Z(n12397) );
  NAND U14796 ( .A(n8606), .B(n6839), .Z(n9748) );
  NAND U14797 ( .A(n8603), .B(n6833), .Z(n12401) );
  AND U14798 ( .A(n12402), .B(n12403), .Z(n12387) );
  AND U14799 ( .A(n12404), .B(n12405), .Z(n12403) );
  AND U14800 ( .A(n10120), .B(n9388), .Z(n12405) );
  NAND U14801 ( .A(n8609), .B(n6835), .Z(n9388) );
  NAND U14802 ( .A(n6850), .B(n8610), .Z(n10120) );
  AND U14803 ( .A(n10860), .B(n10486), .Z(n12404) );
  NAND U14804 ( .A(n8616), .B(n6853), .Z(n10486) );
  NAND U14805 ( .A(n8958), .B(n6841), .Z(n10860) );
  AND U14806 ( .A(n12406), .B(n12407), .Z(n12402) );
  AND U14807 ( .A(n11791), .B(n11226), .Z(n12407) );
  NAND U14808 ( .A(n9082), .B(n6857), .Z(n11226) );
  NAND U14809 ( .A(n9135), .B(n6859), .Z(n11791) );
  AND U14810 ( .A(n12408), .B(n12135), .Z(n12406) );
  NAND U14811 ( .A(n6865), .B(n6984), .Z(n12135) );
  NAND U14812 ( .A(n6967), .B(n6893), .Z(n12408) );
  AND U14813 ( .A(n12409), .B(n12410), .Z(n12377) );
  NAND U14814 ( .A(n12411), .B(n6888), .Z(n12410) );
  NAND U14815 ( .A(n12412), .B(n12413), .Z(n12411) );
  AND U14816 ( .A(n12414), .B(n12415), .Z(n12413) );
  AND U14817 ( .A(n12416), .B(n12417), .Z(n12415) );
  AND U14818 ( .A(n12418), .B(n12419), .Z(n12417) );
  AND U14819 ( .A(n12420), .B(n12421), .Z(n12419) );
  NANDN U14820 ( .B(n8538), .A(n6919), .Z(n12421) );
  NAND U14821 ( .A(n6967), .B(n8512), .Z(n12420) );
  AND U14822 ( .A(n12422), .B(n12423), .Z(n12418) );
  NANDN U14823 ( .B(n8543), .A(n6920), .Z(n12423) );
  NANDN U14824 ( .B(n8516), .A(n6966), .Z(n12422) );
  AND U14825 ( .A(n12424), .B(n12425), .Z(n12416) );
  AND U14826 ( .A(n12426), .B(n12427), .Z(n12425) );
  NANDN U14827 ( .B(n8544), .A(n6925), .Z(n12427) );
  NANDN U14828 ( .B(n8522), .A(n6961), .Z(n12426) );
  AND U14829 ( .A(n12428), .B(n12429), .Z(n12424) );
  NANDN U14830 ( .B(n8547), .A(n6926), .Z(n12429) );
  NANDN U14831 ( .B(n8526), .A(n6956), .Z(n12428) );
  AND U14832 ( .A(n12430), .B(n12431), .Z(n12414) );
  AND U14833 ( .A(n12432), .B(n12433), .Z(n12431) );
  AND U14834 ( .A(n12434), .B(n12435), .Z(n12433) );
  NANDN U14835 ( .B(n8548), .A(n6898), .Z(n12435) );
  NANDN U14836 ( .B(n8534), .A(n6960), .Z(n12434) );
  AND U14837 ( .A(n12436), .B(n12437), .Z(n12432) );
  NANDN U14838 ( .B(n8511), .A(n6957), .Z(n12437) );
  NANDN U14839 ( .B(n8557), .A(n6882), .Z(n12436) );
  AND U14840 ( .A(n12438), .B(n12439), .Z(n12430) );
  AND U14841 ( .A(n12440), .B(n12441), .Z(n12439) );
  NANDN U14842 ( .B(n8515), .A(n6947), .Z(n12441) );
  NANDN U14843 ( .B(n8558), .A(n6809), .Z(n12440) );
  AND U14844 ( .A(n12442), .B(n12443), .Z(n12438) );
  NANDN U14845 ( .B(n8521), .A(n6946), .Z(n12443) );
  NANDN U14846 ( .B(n8561), .A(n6807), .Z(n12442) );
  AND U14847 ( .A(n12444), .B(n12445), .Z(n12412) );
  AND U14848 ( .A(n12446), .B(n12447), .Z(n12445) );
  AND U14849 ( .A(n12448), .B(n12449), .Z(n12447) );
  AND U14850 ( .A(n12450), .B(n12451), .Z(n12449) );
  NANDN U14851 ( .B(n8525), .A(n6943), .Z(n12451) );
  NANDN U14852 ( .B(n8562), .A(n6799), .Z(n12450) );
  AND U14853 ( .A(n12452), .B(n12453), .Z(n12448) );
  NANDN U14854 ( .B(n8567), .A(n6803), .Z(n12453) );
  NANDN U14855 ( .B(n8533), .A(n6942), .Z(n12452) );
  AND U14856 ( .A(n12454), .B(n12455), .Z(n12446) );
  AND U14857 ( .A(n12456), .B(n12457), .Z(n12455) );
  NANDN U14858 ( .B(n8568), .A(n6823), .Z(n12457) );
  NANDN U14859 ( .B(n8537), .A(n6937), .Z(n12456) );
  AND U14860 ( .A(n12458), .B(n12459), .Z(n12454) );
  NANDN U14861 ( .B(n8571), .A(n6827), .Z(n12459) );
  NANDN U14862 ( .B(n8572), .A(n6833), .Z(n12458) );
  AND U14863 ( .A(n12460), .B(n12461), .Z(n12444) );
  AND U14864 ( .A(n12462), .B(n12463), .Z(n12461) );
  AND U14865 ( .A(n12464), .B(n12465), .Z(n12463) );
  NANDN U14866 ( .B(n8579), .A(n6835), .Z(n12465) );
  NANDN U14867 ( .B(n8580), .A(n6839), .Z(n12464) );
  AND U14868 ( .A(n12466), .B(n12467), .Z(n12462) );
  NANDN U14869 ( .B(n8583), .A(n6850), .Z(n12467) );
  NANDN U14870 ( .B(n8584), .A(n6853), .Z(n12466) );
  AND U14871 ( .A(n12468), .B(n12469), .Z(n12460) );
  AND U14872 ( .A(n12470), .B(n12471), .Z(n12469) );
  NANDN U14873 ( .B(n8589), .A(n6841), .Z(n12471) );
  NANDN U14874 ( .B(n8590), .A(n6857), .Z(n12470) );
  AND U14875 ( .A(n12472), .B(n12473), .Z(n12468) );
  NANDN U14876 ( .B(n8593), .A(n6859), .Z(n12473) );
  NAND U14877 ( .A(n6865), .B(n6897), .Z(n12472) );
  NAND U14878 ( .A(n12474), .B(n6902), .Z(n12409) );
  NAND U14879 ( .A(n12475), .B(n12476), .Z(n12474) );
  AND U14880 ( .A(n12477), .B(n12478), .Z(n12476) );
  AND U14881 ( .A(n12479), .B(n12480), .Z(n12478) );
  AND U14882 ( .A(n12481), .B(n12482), .Z(n12480) );
  NAND U14883 ( .A(n6967), .B(n6916), .Z(n12482) );
  NAND U14884 ( .A(n8464), .B(n6898), .Z(n12481) );
  AND U14885 ( .A(n12483), .B(n12484), .Z(n12479) );
  NAND U14886 ( .A(n8465), .B(n6926), .Z(n12484) );
  NAND U14887 ( .A(n8461), .B(n6925), .Z(n12483) );
  AND U14888 ( .A(n12485), .B(n12486), .Z(n12477) );
  AND U14889 ( .A(n12487), .B(n12488), .Z(n12486) );
  NAND U14890 ( .A(n8470), .B(n6920), .Z(n12488) );
  NAND U14891 ( .A(n9359), .B(n6919), .Z(n12487) );
  AND U14892 ( .A(n11893), .B(n12489), .Z(n12485) );
  NAND U14893 ( .A(n9726), .B(n6937), .Z(n12489) );
  NAND U14894 ( .A(n8606), .B(n6946), .Z(n11893) );
  AND U14895 ( .A(n12490), .B(n12491), .Z(n12475) );
  AND U14896 ( .A(n12492), .B(n12493), .Z(n12491) );
  AND U14897 ( .A(n6873), .B(n12494), .Z(n12493) );
  NAND U14898 ( .A(n8603), .B(n6942), .Z(n12494) );
  NAND U14899 ( .A(n8609), .B(n6943), .Z(n6873) );
  AND U14900 ( .A(n9131), .B(n12495), .Z(n12492) );
  NAND U14901 ( .A(n8616), .B(n6957), .Z(n9131) );
  AND U14902 ( .A(n12496), .B(n12497), .Z(n12490) );
  AND U14903 ( .A(n8496), .B(n12498), .Z(n12497) );
  NAND U14904 ( .A(n6956), .B(n9082), .Z(n8496) );
  AND U14905 ( .A(n12499), .B(n12500), .Z(n12496) );
  IV U14906 ( .A(\u_a23_core/u_execute/rn[15] ), .Z(n12376) );
  AND U14907 ( .A(n12501), .B(n8620), .Z(n12367) );
  NAND U14908 ( .A(n6765), .B(\u_a23_core/u_execute/u_alu/fadder_out[15] ), 
        .Z(n12501) );
  AND U14909 ( .A(n12502), .B(n12503), .Z(n12363) );
  NANDN U14910 ( .B(n8406), .A(\u_a23_core/u_execute/rn_plus4[15] ), .Z(n12503) );
  NANDN U14911 ( .B(n8407), .A(\u_a23_core/u_execute/alu_plus4[15] ), .Z(
        n12502) );
  AND U14912 ( .A(n12504), .B(n12505), .Z(n12361) );
  AND U14913 ( .A(n12506), .B(n12507), .Z(n12505) );
  NAND U14914 ( .A(n8412), .B(\u_a23_core/u_execute/address_plus4[15] ), .Z(
        n12507) );
  NAND U14915 ( .A(\u_a23_core/u_execute/rn[15] ), .B(n8413), .Z(n12506) );
  NAND U14916 ( .A(n12508), .B(n12509), .Z(\u_a23_core/u_execute/rn[15] ) );
  AND U14917 ( .A(n12510), .B(n12511), .Z(n12509) );
  AND U14918 ( .A(n12512), .B(n12513), .Z(n12511) );
  AND U14919 ( .A(n12514), .B(n12515), .Z(n12513) );
  NANDN U14920 ( .B(n8635), .A(\u_a23_core/u_execute/pc[15] ), .Z(n12515) );
  NANDN U14921 ( .B(n8636), .A(\u_a23_core/u_execute/u_register_bank/r14[15] ), 
        .Z(n12514) );
  AND U14922 ( .A(n12516), .B(n12517), .Z(n12512) );
  NANDN U14923 ( .B(n8639), .A(\u_a23_core/u_execute/u_register_bank/r13[15] ), 
        .Z(n12517) );
  NANDN U14924 ( .B(n8640), .A(\u_a23_core/u_execute/u_register_bank/r12[15] ), 
        .Z(n12516) );
  AND U14925 ( .A(n12518), .B(n12519), .Z(n12510) );
  AND U14926 ( .A(n12520), .B(n12521), .Z(n12519) );
  NANDN U14927 ( .B(n8645), .A(\u_a23_core/u_execute/u_register_bank/r11[15] ), 
        .Z(n12521) );
  NANDN U14928 ( .B(n8646), .A(\u_a23_core/u_execute/u_register_bank/r10[15] ), 
        .Z(n12520) );
  AND U14929 ( .A(n12522), .B(n12523), .Z(n12518) );
  NANDN U14930 ( .B(n8649), .A(\u_a23_core/u_execute/u_register_bank/r9[15] ), 
        .Z(n12523) );
  NANDN U14931 ( .B(n8650), .A(\u_a23_core/u_execute/u_register_bank/r8[15] ), 
        .Z(n12522) );
  AND U14932 ( .A(n12524), .B(n12525), .Z(n12508) );
  AND U14933 ( .A(n12526), .B(n12527), .Z(n12525) );
  AND U14934 ( .A(n12528), .B(n12529), .Z(n12527) );
  NANDN U14935 ( .B(n8657), .A(\u_a23_core/u_execute/u_register_bank/r7[15] ), 
        .Z(n12529) );
  NANDN U14936 ( .B(n8658), .A(\u_a23_core/u_execute/u_register_bank/r6[15] ), 
        .Z(n12528) );
  AND U14937 ( .A(n12530), .B(n12531), .Z(n12526) );
  NANDN U14938 ( .B(n8661), .A(\u_a23_core/u_execute/u_register_bank/r5[15] ), 
        .Z(n12531) );
  NANDN U14939 ( .B(n8662), .A(\u_a23_core/u_execute/u_register_bank/r4[15] ), 
        .Z(n12530) );
  AND U14940 ( .A(n12532), .B(n12533), .Z(n12524) );
  AND U14941 ( .A(n12534), .B(n12535), .Z(n12533) );
  NANDN U14942 ( .B(n8667), .A(\u_a23_core/u_execute/u_register_bank/r3[15] ), 
        .Z(n12535) );
  NANDN U14943 ( .B(n8668), .A(\u_a23_core/u_execute/u_register_bank/r0[15] ), 
        .Z(n12534) );
  AND U14944 ( .A(n12536), .B(n12537), .Z(n12532) );
  NANDN U14945 ( .B(n8671), .A(\u_a23_core/u_execute/u_register_bank/r2[15] ), 
        .Z(n12537) );
  NANDN U14946 ( .B(n8672), .A(\u_a23_core/u_execute/u_register_bank/r1[15] ), 
        .Z(n12536) );
  AND U14947 ( .A(n12538), .B(n12539), .Z(n12504) );
  NAND U14948 ( .A(\u_a23_core/u_execute/pc[15] ), .B(n8416), .Z(n12539) );
  NAND U14949 ( .A(n8417), .B(\u_a23_core/u_execute/pc_plus4[15] ), .Z(n12538)
         );
  NAND U14950 ( .A(n12540), .B(n12541), .Z(
        \u_a23_core/execute_address_nxt[14] ) );
  AND U14951 ( .A(n12542), .B(n12543), .Z(n12541) );
  AND U14952 ( .A(n12544), .B(n12545), .Z(n12543) );
  NANDN U14953 ( .B(n8392), .A(\u_a23_core/u_execute/pc_minus4[14] ), .Z(
        n12545) );
  NAND U14954 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[14] ), .B(n8393), 
        .Z(n12544) );
  IV U14955 ( .A(n7041), .Z(\u_a23_core/u_execute/alu_out_pc_filtered[14] ) );
  AND U14956 ( .A(n12546), .B(n12547), .Z(n7041) );
  MUX U14957 ( .IN0(n12548), .IN1(n12549), .SEL(
        \u_a23_core/u_execute/u_alu/b_not[14] ), .F(n12547) );
  NAND U14958 ( .A(n12550), .B(n12551), .Z(
        \u_a23_core/u_execute/u_alu/b_not[14] ) );
  MUX U14959 ( .IN0(n8430), .IN1(n8431), .SEL(n12552), .F(n12551) );
  MUX U14960 ( .IN0(n8433), .IN1(n8434), .SEL(\u_a23_core/u_execute/rn[14] ), 
        .F(n12550) );
  ANDN U14961 ( .A(n8435), .B(n12553), .Z(n12549) );
  MUX U14962 ( .IN0(n8400), .IN1(\u_a23_core/alu_function[3] ), .SEL(
        \u_a23_core/u_execute/u_alu/a[14] ), .F(n12553) );
  NAND U14963 ( .A(\u_a23_core/u_execute/u_alu/a[14] ), .B(n8400), .Z(n12548)
         );
  IV U14964 ( .A(n12554), .Z(\u_a23_core/u_execute/u_alu/a[14] ) );
  MUX U14965 ( .IN0(n12555), .IN1(n12552), .SEL(\u_a23_core/alu_function[8] ), 
        .F(n12554) );
  AND U14966 ( .A(n12556), .B(n12557), .Z(n12552) );
  AND U14967 ( .A(n12558), .B(n12559), .Z(n12557) );
  NAND U14968 ( .A(n6786), .B(n12560), .Z(n12559) );
  NAND U14969 ( .A(n12561), .B(n12562), .Z(n12560) );
  AND U14970 ( .A(n12563), .B(n12564), .Z(n12562) );
  AND U14971 ( .A(n12565), .B(n12566), .Z(n12564) );
  AND U14972 ( .A(n12567), .B(n12568), .Z(n12566) );
  NAND U14973 ( .A(n8461), .B(n6803), .Z(n12568) );
  AND U14974 ( .A(n12569), .B(n12570), .Z(n12567) );
  NAND U14975 ( .A(n8464), .B(n6807), .Z(n12570) );
  NAND U14976 ( .A(n8465), .B(n6799), .Z(n12569) );
  AND U14977 ( .A(n12571), .B(n12572), .Z(n12565) );
  NAND U14978 ( .A(n8470), .B(n6823), .Z(n12572) );
  NAND U14979 ( .A(n9359), .B(n6827), .Z(n12571) );
  AND U14980 ( .A(n12573), .B(n12574), .Z(n12563) );
  AND U14981 ( .A(n12575), .B(n12576), .Z(n12574) );
  NAND U14982 ( .A(n9726), .B(n6833), .Z(n12576) );
  NAND U14983 ( .A(n6809), .B(n8487), .Z(n12575) );
  AND U14984 ( .A(n6975), .B(n9932), .Z(n12573) );
  NAND U14985 ( .A(n6850), .B(n8606), .Z(n9932) );
  NAND U14986 ( .A(n8603), .B(n6835), .Z(n6975) );
  AND U14987 ( .A(n12577), .B(n12578), .Z(n12561) );
  AND U14988 ( .A(n12579), .B(n12580), .Z(n12578) );
  AND U14989 ( .A(n10306), .B(n9500), .Z(n12580) );
  NAND U14990 ( .A(n8609), .B(n6839), .Z(n9500) );
  NAND U14991 ( .A(n8610), .B(n6853), .Z(n10306) );
  AND U14992 ( .A(n11046), .B(n10672), .Z(n12579) );
  NAND U14993 ( .A(n8616), .B(n6841), .Z(n10672) );
  NAND U14994 ( .A(n8958), .B(n6857), .Z(n11046) );
  AND U14995 ( .A(n12581), .B(n12582), .Z(n12577) );
  AND U14996 ( .A(n11605), .B(n11413), .Z(n12582) );
  NAND U14997 ( .A(n9082), .B(n6859), .Z(n11413) );
  NAND U14998 ( .A(n6865), .B(n9135), .Z(n11605) );
  AND U14999 ( .A(n12583), .B(n12315), .Z(n12581) );
  NAND U15000 ( .A(n6967), .B(n6984), .Z(n12315) );
  NAND U15001 ( .A(n6966), .B(n6893), .Z(n12583) );
  AND U15002 ( .A(n12584), .B(n12585), .Z(n12558) );
  NAND U15003 ( .A(n6886), .B(n12586), .Z(n12585) );
  NANDN U15004 ( .B(n12383), .A(n8448), .Z(n12586) );
  NAND U15005 ( .A(n12587), .B(n12588), .Z(n12383) );
  AND U15006 ( .A(n12589), .B(n12590), .Z(n12588) );
  AND U15007 ( .A(n12591), .B(n12592), .Z(n12589) );
  IV U15008 ( .A(n6864), .Z(n12591) );
  AND U15009 ( .A(n8449), .B(n12593), .Z(n12587) );
  AND U15010 ( .A(n12594), .B(n12595), .Z(n12593) );
  NAND U15011 ( .A(n6864), .B(n6985), .Z(n12584) );
  AND U15012 ( .A(n12596), .B(n12597), .Z(n12556) );
  NAND U15013 ( .A(n12598), .B(n6888), .Z(n12597) );
  NAND U15014 ( .A(n12599), .B(n12600), .Z(n12598) );
  AND U15015 ( .A(n12601), .B(n12602), .Z(n12600) );
  AND U15016 ( .A(n12603), .B(n12604), .Z(n12602) );
  AND U15017 ( .A(n12605), .B(n12606), .Z(n12604) );
  AND U15018 ( .A(n12607), .B(n12608), .Z(n12606) );
  NANDN U15019 ( .B(n8537), .A(n6919), .Z(n12608) );
  NAND U15020 ( .A(n6966), .B(n8512), .Z(n12607) );
  AND U15021 ( .A(n12609), .B(n12610), .Z(n12605) );
  NANDN U15022 ( .B(n8538), .A(n6920), .Z(n12610) );
  NANDN U15023 ( .B(n8516), .A(n6961), .Z(n12609) );
  AND U15024 ( .A(n12611), .B(n12612), .Z(n12603) );
  AND U15025 ( .A(n12613), .B(n12614), .Z(n12612) );
  NANDN U15026 ( .B(n8543), .A(n6925), .Z(n12614) );
  NANDN U15027 ( .B(n8522), .A(n6956), .Z(n12613) );
  AND U15028 ( .A(n12615), .B(n12616), .Z(n12611) );
  NANDN U15029 ( .B(n8544), .A(n6926), .Z(n12616) );
  NANDN U15030 ( .B(n8526), .A(n6960), .Z(n12615) );
  AND U15031 ( .A(n12617), .B(n12618), .Z(n12601) );
  AND U15032 ( .A(n12619), .B(n12620), .Z(n12618) );
  AND U15033 ( .A(n12621), .B(n12622), .Z(n12620) );
  NANDN U15034 ( .B(n8547), .A(n6898), .Z(n12622) );
  NANDN U15035 ( .B(n8534), .A(n6957), .Z(n12621) );
  AND U15036 ( .A(n12623), .B(n12624), .Z(n12619) );
  NANDN U15037 ( .B(n8511), .A(n6947), .Z(n12624) );
  NANDN U15038 ( .B(n8548), .A(n6882), .Z(n12623) );
  AND U15039 ( .A(n12625), .B(n12626), .Z(n12617) );
  AND U15040 ( .A(n12627), .B(n12628), .Z(n12626) );
  NANDN U15041 ( .B(n8515), .A(n6946), .Z(n12628) );
  NANDN U15042 ( .B(n8557), .A(n6809), .Z(n12627) );
  AND U15043 ( .A(n12629), .B(n12630), .Z(n12625) );
  NANDN U15044 ( .B(n8521), .A(n6943), .Z(n12630) );
  NANDN U15045 ( .B(n8558), .A(n6807), .Z(n12629) );
  AND U15046 ( .A(n12631), .B(n12632), .Z(n12599) );
  AND U15047 ( .A(n12633), .B(n12634), .Z(n12632) );
  AND U15048 ( .A(n12635), .B(n12636), .Z(n12634) );
  AND U15049 ( .A(n12637), .B(n12638), .Z(n12636) );
  NANDN U15050 ( .B(n8525), .A(n6942), .Z(n12638) );
  NANDN U15051 ( .B(n8561), .A(n6799), .Z(n12637) );
  AND U15052 ( .A(n12639), .B(n12640), .Z(n12635) );
  NANDN U15053 ( .B(n8562), .A(n6803), .Z(n12640) );
  NANDN U15054 ( .B(n8533), .A(n6937), .Z(n12639) );
  AND U15055 ( .A(n12641), .B(n12642), .Z(n12633) );
  AND U15056 ( .A(n12643), .B(n12644), .Z(n12642) );
  NANDN U15057 ( .B(n8567), .A(n6823), .Z(n12644) );
  NANDN U15058 ( .B(n8568), .A(n6827), .Z(n12643) );
  AND U15059 ( .A(n12645), .B(n12646), .Z(n12641) );
  NANDN U15060 ( .B(n8571), .A(n6833), .Z(n12646) );
  NANDN U15061 ( .B(n8572), .A(n6835), .Z(n12645) );
  AND U15062 ( .A(n12647), .B(n12648), .Z(n12631) );
  AND U15063 ( .A(n12649), .B(n12650), .Z(n12648) );
  AND U15064 ( .A(n12651), .B(n12652), .Z(n12650) );
  NANDN U15065 ( .B(n8579), .A(n6839), .Z(n12652) );
  NANDN U15066 ( .B(n8580), .A(n6850), .Z(n12651) );
  AND U15067 ( .A(n12653), .B(n12654), .Z(n12649) );
  NANDN U15068 ( .B(n8583), .A(n6853), .Z(n12654) );
  NANDN U15069 ( .B(n8584), .A(n6841), .Z(n12653) );
  AND U15070 ( .A(n12655), .B(n12656), .Z(n12647) );
  AND U15071 ( .A(n12657), .B(n12658), .Z(n12656) );
  NANDN U15072 ( .B(n8589), .A(n6857), .Z(n12658) );
  NANDN U15073 ( .B(n8590), .A(n6859), .Z(n12657) );
  AND U15074 ( .A(n12659), .B(n12660), .Z(n12655) );
  NANDN U15075 ( .B(n8593), .A(n6865), .Z(n12660) );
  NAND U15076 ( .A(n6967), .B(n6897), .Z(n12659) );
  NAND U15077 ( .A(n12661), .B(n6902), .Z(n12596) );
  NAND U15078 ( .A(n12662), .B(n12663), .Z(n12661) );
  AND U15079 ( .A(n12664), .B(n12665), .Z(n12663) );
  AND U15080 ( .A(n12666), .B(n12667), .Z(n12665) );
  AND U15081 ( .A(n12668), .B(n12669), .Z(n12667) );
  NAND U15082 ( .A(n6966), .B(n6916), .Z(n12669) );
  NAND U15083 ( .A(n8465), .B(n6898), .Z(n12668) );
  AND U15084 ( .A(n12670), .B(n12671), .Z(n12666) );
  NAND U15085 ( .A(n8461), .B(n6926), .Z(n12671) );
  NAND U15086 ( .A(n8470), .B(n6925), .Z(n12670) );
  AND U15087 ( .A(n12672), .B(n12673), .Z(n12664) );
  AND U15088 ( .A(n12674), .B(n12675), .Z(n12673) );
  NAND U15089 ( .A(n9359), .B(n6920), .Z(n12675) );
  NAND U15090 ( .A(n9726), .B(n6919), .Z(n12674) );
  AND U15091 ( .A(n12676), .B(n12677), .Z(n12672) );
  NAND U15092 ( .A(n8603), .B(n6937), .Z(n12676) );
  AND U15093 ( .A(n12678), .B(n12679), .Z(n12662) );
  AND U15094 ( .A(n12680), .B(n12681), .Z(n12679) );
  AND U15095 ( .A(n12682), .B(n12683), .Z(n12681) );
  NAND U15096 ( .A(n8609), .B(n6942), .Z(n12683) );
  AND U15097 ( .A(n9007), .B(n12684), .Z(n12680) );
  NAND U15098 ( .A(n8958), .B(n6957), .Z(n9007) );
  AND U15099 ( .A(n12685), .B(n12686), .Z(n12678) );
  AND U15100 ( .A(n12687), .B(n8736), .Z(n12685) );
  NAND U15101 ( .A(n9082), .B(n6960), .Z(n8736) );
  IV U15102 ( .A(\u_a23_core/u_execute/rn[14] ), .Z(n12555) );
  AND U15103 ( .A(n12688), .B(n8620), .Z(n12546) );
  NAND U15104 ( .A(n6765), .B(\u_a23_core/u_execute/u_alu/fadder_out[14] ), 
        .Z(n12688) );
  AND U15105 ( .A(n12689), .B(n12690), .Z(n12542) );
  NANDN U15106 ( .B(n8406), .A(\u_a23_core/u_execute/rn_plus4[14] ), .Z(n12690) );
  NANDN U15107 ( .B(n8407), .A(\u_a23_core/u_execute/alu_plus4[14] ), .Z(
        n12689) );
  AND U15108 ( .A(n12691), .B(n12692), .Z(n12540) );
  AND U15109 ( .A(n12693), .B(n12694), .Z(n12692) );
  NAND U15110 ( .A(n8412), .B(\u_a23_core/u_execute/address_plus4[14] ), .Z(
        n12694) );
  NAND U15111 ( .A(\u_a23_core/u_execute/rn[14] ), .B(n8413), .Z(n12693) );
  NAND U15112 ( .A(n12695), .B(n12696), .Z(\u_a23_core/u_execute/rn[14] ) );
  AND U15113 ( .A(n12697), .B(n12698), .Z(n12696) );
  AND U15114 ( .A(n12699), .B(n12700), .Z(n12698) );
  AND U15115 ( .A(n12701), .B(n12702), .Z(n12700) );
  NANDN U15116 ( .B(n8635), .A(\u_a23_core/u_execute/pc[14] ), .Z(n12702) );
  NANDN U15117 ( .B(n8636), .A(\u_a23_core/u_execute/u_register_bank/r14[14] ), 
        .Z(n12701) );
  AND U15118 ( .A(n12703), .B(n12704), .Z(n12699) );
  NANDN U15119 ( .B(n8639), .A(\u_a23_core/u_execute/u_register_bank/r13[14] ), 
        .Z(n12704) );
  NANDN U15120 ( .B(n8640), .A(\u_a23_core/u_execute/u_register_bank/r12[14] ), 
        .Z(n12703) );
  AND U15121 ( .A(n12705), .B(n12706), .Z(n12697) );
  AND U15122 ( .A(n12707), .B(n12708), .Z(n12706) );
  NANDN U15123 ( .B(n8645), .A(\u_a23_core/u_execute/u_register_bank/r11[14] ), 
        .Z(n12708) );
  NANDN U15124 ( .B(n8646), .A(\u_a23_core/u_execute/u_register_bank/r10[14] ), 
        .Z(n12707) );
  AND U15125 ( .A(n12709), .B(n12710), .Z(n12705) );
  NANDN U15126 ( .B(n8649), .A(\u_a23_core/u_execute/u_register_bank/r9[14] ), 
        .Z(n12710) );
  NANDN U15127 ( .B(n8650), .A(\u_a23_core/u_execute/u_register_bank/r8[14] ), 
        .Z(n12709) );
  AND U15128 ( .A(n12711), .B(n12712), .Z(n12695) );
  AND U15129 ( .A(n12713), .B(n12714), .Z(n12712) );
  AND U15130 ( .A(n12715), .B(n12716), .Z(n12714) );
  NANDN U15131 ( .B(n8657), .A(\u_a23_core/u_execute/u_register_bank/r7[14] ), 
        .Z(n12716) );
  NANDN U15132 ( .B(n8658), .A(\u_a23_core/u_execute/u_register_bank/r6[14] ), 
        .Z(n12715) );
  AND U15133 ( .A(n12717), .B(n12718), .Z(n12713) );
  NANDN U15134 ( .B(n8661), .A(\u_a23_core/u_execute/u_register_bank/r5[14] ), 
        .Z(n12718) );
  NANDN U15135 ( .B(n8662), .A(\u_a23_core/u_execute/u_register_bank/r4[14] ), 
        .Z(n12717) );
  AND U15136 ( .A(n12719), .B(n12720), .Z(n12711) );
  AND U15137 ( .A(n12721), .B(n12722), .Z(n12720) );
  NANDN U15138 ( .B(n8667), .A(\u_a23_core/u_execute/u_register_bank/r3[14] ), 
        .Z(n12722) );
  NANDN U15139 ( .B(n8668), .A(\u_a23_core/u_execute/u_register_bank/r0[14] ), 
        .Z(n12721) );
  AND U15140 ( .A(n12723), .B(n12724), .Z(n12719) );
  NANDN U15141 ( .B(n8671), .A(\u_a23_core/u_execute/u_register_bank/r2[14] ), 
        .Z(n12724) );
  NANDN U15142 ( .B(n8672), .A(\u_a23_core/u_execute/u_register_bank/r1[14] ), 
        .Z(n12723) );
  AND U15143 ( .A(n12725), .B(n12726), .Z(n12691) );
  NAND U15144 ( .A(\u_a23_core/u_execute/pc[14] ), .B(n8416), .Z(n12726) );
  NAND U15145 ( .A(n8417), .B(\u_a23_core/u_execute/pc_plus4[14] ), .Z(n12725)
         );
  NOR U15146 ( .A(\u_a23_core/execute_address_nxt[12] ), .B(
        \u_a23_core/execute_address_nxt[13] ), .Z(n12359) );
  NAND U15147 ( .A(n12727), .B(n12728), .Z(
        \u_a23_core/execute_address_nxt[13] ) );
  AND U15148 ( .A(n12729), .B(n12730), .Z(n12728) );
  AND U15149 ( .A(n12731), .B(n12732), .Z(n12730) );
  NANDN U15150 ( .B(n8392), .A(\u_a23_core/u_execute/pc_minus4[13] ), .Z(
        n12732) );
  NAND U15151 ( .A(n8393), .B(\u_a23_core/u_execute/alu_out_pc_filtered[13] ), 
        .Z(n12731) );
  IV U15152 ( .A(n7044), .Z(\u_a23_core/u_execute/alu_out_pc_filtered[13] ) );
  AND U15153 ( .A(n12733), .B(n12734), .Z(n7044) );
  MUX U15154 ( .IN0(n12735), .IN1(n12736), .SEL(
        \u_a23_core/u_execute/u_alu/b_not[13] ), .F(n12734) );
  NAND U15155 ( .A(n12737), .B(n12738), .Z(
        \u_a23_core/u_execute/u_alu/b_not[13] ) );
  MUX U15156 ( .IN0(n8430), .IN1(n8431), .SEL(n12739), .F(n12738) );
  MUX U15157 ( .IN0(n8433), .IN1(n8434), .SEL(\u_a23_core/u_execute/rn[13] ), 
        .F(n12737) );
  ANDN U15158 ( .A(n8435), .B(n12740), .Z(n12736) );
  MUX U15159 ( .IN0(n8400), .IN1(\u_a23_core/alu_function[3] ), .SEL(
        \u_a23_core/u_execute/u_alu/a[13] ), .F(n12740) );
  NAND U15160 ( .A(\u_a23_core/u_execute/u_alu/a[13] ), .B(n8400), .Z(n12735)
         );
  IV U15161 ( .A(n12741), .Z(\u_a23_core/u_execute/u_alu/a[13] ) );
  MUX U15162 ( .IN0(n12742), .IN1(n12739), .SEL(\u_a23_core/alu_function[8] ), 
        .F(n12741) );
  AND U15163 ( .A(n12743), .B(n12744), .Z(n12739) );
  AND U15164 ( .A(n12745), .B(n12746), .Z(n12744) );
  NAND U15165 ( .A(n8443), .B(n12747), .Z(n12746) );
  AND U15166 ( .A(n12748), .B(n6882), .Z(n12747) );
  NAND U15167 ( .A(n12749), .B(n12750), .Z(n12748) );
  AND U15168 ( .A(n12751), .B(n12594), .Z(n12750) );
  AND U15169 ( .A(n12592), .B(n12590), .Z(n12751) );
  IV U15170 ( .A(n6858), .Z(n12592) );
  AND U15171 ( .A(n8449), .B(n12752), .Z(n12749) );
  AND U15172 ( .A(n8448), .B(n12595), .Z(n12752) );
  AND U15173 ( .A(n12753), .B(n12754), .Z(n8448) );
  AND U15174 ( .A(n12755), .B(n12756), .Z(n12754) );
  NOR U15175 ( .A(n6806), .B(n6798), .Z(n12755) );
  AND U15176 ( .A(n12757), .B(n12758), .Z(n12753) );
  NOR U15177 ( .A(n6802), .B(n6826), .Z(n12757) );
  AND U15178 ( .A(n12759), .B(n12760), .Z(n12745) );
  NAND U15179 ( .A(n6858), .B(n6985), .Z(n12760) );
  NAND U15180 ( .A(n6786), .B(n12761), .Z(n12759) );
  NAND U15181 ( .A(n12762), .B(n12763), .Z(n12761) );
  AND U15182 ( .A(n12764), .B(n12765), .Z(n12763) );
  AND U15183 ( .A(n12766), .B(n12767), .Z(n12765) );
  AND U15184 ( .A(n12768), .B(n12769), .Z(n12767) );
  NAND U15185 ( .A(n8461), .B(n6823), .Z(n12769) );
  AND U15186 ( .A(n12770), .B(n12771), .Z(n12768) );
  NAND U15187 ( .A(n8464), .B(n6799), .Z(n12771) );
  NAND U15188 ( .A(n8465), .B(n6803), .Z(n12770) );
  AND U15189 ( .A(n12772), .B(n12773), .Z(n12766) );
  NAND U15190 ( .A(n8470), .B(n6827), .Z(n12773) );
  NAND U15191 ( .A(n9359), .B(n6833), .Z(n12772) );
  AND U15192 ( .A(n12774), .B(n12775), .Z(n12764) );
  AND U15193 ( .A(n12776), .B(n12777), .Z(n12775) );
  NAND U15194 ( .A(n9726), .B(n6835), .Z(n12777) );
  NAND U15195 ( .A(n6864), .B(n6809), .Z(n12776) );
  AND U15196 ( .A(n10114), .B(n12778), .Z(n12774) );
  NAND U15197 ( .A(n6807), .B(n8487), .Z(n12778) );
  NAND U15198 ( .A(n8606), .B(n6853), .Z(n10114) );
  AND U15199 ( .A(n12779), .B(n12780), .Z(n12762) );
  AND U15200 ( .A(n12781), .B(n12782), .Z(n12780) );
  AND U15201 ( .A(n12783), .B(n10487), .Z(n12782) );
  NAND U15202 ( .A(n8610), .B(n6841), .Z(n10487) );
  AND U15203 ( .A(n9754), .B(n9385), .Z(n12783) );
  NAND U15204 ( .A(n8603), .B(n6839), .Z(n9385) );
  NAND U15205 ( .A(n6850), .B(n8609), .Z(n9754) );
  AND U15206 ( .A(n11227), .B(n10861), .Z(n12781) );
  NAND U15207 ( .A(n8616), .B(n6857), .Z(n10861) );
  NAND U15208 ( .A(n8958), .B(n6859), .Z(n11227) );
  AND U15209 ( .A(n12784), .B(n12785), .Z(n12779) );
  AND U15210 ( .A(n12136), .B(n11788), .Z(n12785) );
  NAND U15211 ( .A(n6865), .B(n9082), .Z(n11788) );
  NAND U15212 ( .A(n6967), .B(n9135), .Z(n12136) );
  AND U15213 ( .A(n12786), .B(n12499), .Z(n12784) );
  NAND U15214 ( .A(n6966), .B(n6984), .Z(n12499) );
  NAND U15215 ( .A(n6961), .B(n6893), .Z(n12786) );
  AND U15216 ( .A(n12787), .B(n12788), .Z(n12743) );
  NAND U15217 ( .A(n12789), .B(n6888), .Z(n12788) );
  NAND U15218 ( .A(n12790), .B(n12791), .Z(n12789) );
  AND U15219 ( .A(n12792), .B(n12793), .Z(n12791) );
  AND U15220 ( .A(n12794), .B(n12795), .Z(n12793) );
  AND U15221 ( .A(n12796), .B(n12797), .Z(n12795) );
  AND U15222 ( .A(n12798), .B(n12799), .Z(n12797) );
  NANDN U15223 ( .B(n8533), .A(n6919), .Z(n12799) );
  NAND U15224 ( .A(n6961), .B(n8512), .Z(n12798) );
  AND U15225 ( .A(n12800), .B(n12801), .Z(n12796) );
  NANDN U15226 ( .B(n8537), .A(n6920), .Z(n12801) );
  NANDN U15227 ( .B(n8516), .A(n6956), .Z(n12800) );
  AND U15228 ( .A(n12802), .B(n12803), .Z(n12794) );
  AND U15229 ( .A(n12804), .B(n12805), .Z(n12803) );
  NANDN U15230 ( .B(n8538), .A(n6925), .Z(n12805) );
  NANDN U15231 ( .B(n8522), .A(n6960), .Z(n12804) );
  AND U15232 ( .A(n12806), .B(n12807), .Z(n12802) );
  NANDN U15233 ( .B(n8543), .A(n6926), .Z(n12807) );
  NANDN U15234 ( .B(n8526), .A(n6957), .Z(n12806) );
  AND U15235 ( .A(n12808), .B(n12809), .Z(n12792) );
  AND U15236 ( .A(n12810), .B(n12811), .Z(n12809) );
  AND U15237 ( .A(n12812), .B(n12813), .Z(n12811) );
  NANDN U15238 ( .B(n8544), .A(n6898), .Z(n12813) );
  NANDN U15239 ( .B(n8534), .A(n6947), .Z(n12812) );
  AND U15240 ( .A(n12814), .B(n12815), .Z(n12810) );
  NANDN U15241 ( .B(n8511), .A(n6946), .Z(n12815) );
  NANDN U15242 ( .B(n8547), .A(n6882), .Z(n12814) );
  AND U15243 ( .A(n12816), .B(n12817), .Z(n12808) );
  AND U15244 ( .A(n12818), .B(n12819), .Z(n12817) );
  NANDN U15245 ( .B(n8515), .A(n6943), .Z(n12819) );
  NANDN U15246 ( .B(n8548), .A(n6809), .Z(n12818) );
  AND U15247 ( .A(n12820), .B(n12821), .Z(n12816) );
  NANDN U15248 ( .B(n8521), .A(n6942), .Z(n12821) );
  NANDN U15249 ( .B(n8557), .A(n6807), .Z(n12820) );
  AND U15250 ( .A(n12822), .B(n12823), .Z(n12790) );
  AND U15251 ( .A(n12824), .B(n12825), .Z(n12823) );
  AND U15252 ( .A(n12826), .B(n12827), .Z(n12825) );
  AND U15253 ( .A(n12828), .B(n12829), .Z(n12827) );
  NANDN U15254 ( .B(n8525), .A(n6937), .Z(n12829) );
  NANDN U15255 ( .B(n8558), .A(n6799), .Z(n12828) );
  AND U15256 ( .A(n12830), .B(n12831), .Z(n12826) );
  NANDN U15257 ( .B(n8561), .A(n6803), .Z(n12831) );
  NANDN U15258 ( .B(n8562), .A(n6823), .Z(n12830) );
  AND U15259 ( .A(n12832), .B(n12833), .Z(n12824) );
  AND U15260 ( .A(n12834), .B(n12835), .Z(n12833) );
  NANDN U15261 ( .B(n8567), .A(n6827), .Z(n12835) );
  NANDN U15262 ( .B(n8568), .A(n6833), .Z(n12834) );
  AND U15263 ( .A(n12836), .B(n12837), .Z(n12832) );
  NANDN U15264 ( .B(n8571), .A(n6835), .Z(n12837) );
  NANDN U15265 ( .B(n8572), .A(n6839), .Z(n12836) );
  AND U15266 ( .A(n12838), .B(n12839), .Z(n12822) );
  AND U15267 ( .A(n12840), .B(n12841), .Z(n12839) );
  AND U15268 ( .A(n12842), .B(n12843), .Z(n12841) );
  NANDN U15269 ( .B(n8579), .A(n6850), .Z(n12843) );
  NANDN U15270 ( .B(n8580), .A(n6853), .Z(n12842) );
  AND U15271 ( .A(n12844), .B(n12845), .Z(n12840) );
  NANDN U15272 ( .B(n8583), .A(n6841), .Z(n12845) );
  NANDN U15273 ( .B(n8584), .A(n6857), .Z(n12844) );
  AND U15274 ( .A(n12846), .B(n12847), .Z(n12838) );
  AND U15275 ( .A(n12848), .B(n12849), .Z(n12847) );
  NANDN U15276 ( .B(n8589), .A(n6859), .Z(n12849) );
  NANDN U15277 ( .B(n8590), .A(n6865), .Z(n12848) );
  AND U15278 ( .A(n12850), .B(n12851), .Z(n12846) );
  NANDN U15279 ( .B(n8593), .A(n6967), .Z(n12851) );
  NAND U15280 ( .A(n6966), .B(n6897), .Z(n12850) );
  NAND U15281 ( .A(n12852), .B(n6902), .Z(n12787) );
  NAND U15282 ( .A(n12853), .B(n12854), .Z(n12852) );
  AND U15283 ( .A(n12855), .B(n12856), .Z(n12854) );
  AND U15284 ( .A(n12857), .B(n12858), .Z(n12856) );
  AND U15285 ( .A(n12859), .B(n12860), .Z(n12858) );
  NAND U15286 ( .A(n6961), .B(n6916), .Z(n12860) );
  NAND U15287 ( .A(n8461), .B(n6898), .Z(n12859) );
  AND U15288 ( .A(n12861), .B(n12862), .Z(n12857) );
  NAND U15289 ( .A(n8470), .B(n6926), .Z(n12862) );
  NAND U15290 ( .A(n9359), .B(n6925), .Z(n12861) );
  AND U15291 ( .A(n12863), .B(n12864), .Z(n12855) );
  NAND U15292 ( .A(n8603), .B(n6919), .Z(n12864) );
  AND U15293 ( .A(n6867), .B(n12865), .Z(n12863) );
  NAND U15294 ( .A(n9726), .B(n6920), .Z(n12865) );
  NAND U15295 ( .A(n8606), .B(n6942), .Z(n6867) );
  AND U15296 ( .A(n12866), .B(n12867), .Z(n12853) );
  AND U15297 ( .A(n12868), .B(n12869), .Z(n12867) );
  AND U15298 ( .A(n11901), .B(n12870), .Z(n12869) );
  NAND U15299 ( .A(n8609), .B(n6937), .Z(n12870) );
  NAND U15300 ( .A(n8610), .B(n6943), .Z(n11901) );
  AND U15301 ( .A(n9130), .B(n12871), .Z(n12868) );
  NAND U15302 ( .A(n8958), .B(n6947), .Z(n9130) );
  AND U15303 ( .A(n12872), .B(n12873), .Z(n12866) );
  AND U15304 ( .A(n8495), .B(n12874), .Z(n12872) );
  NAND U15305 ( .A(n9135), .B(n6960), .Z(n8495) );
  IV U15306 ( .A(\u_a23_core/u_execute/rn[13] ), .Z(n12742) );
  AND U15307 ( .A(n12875), .B(n8620), .Z(n12733) );
  NAND U15308 ( .A(n6765), .B(\u_a23_core/u_execute/u_alu/fadder_out[13] ), 
        .Z(n12875) );
  AND U15309 ( .A(n12876), .B(n12877), .Z(n12729) );
  NANDN U15310 ( .B(n8406), .A(\u_a23_core/u_execute/rn_plus4[13] ), .Z(n12877) );
  NANDN U15311 ( .B(n8407), .A(\u_a23_core/u_execute/alu_plus4[13] ), .Z(
        n12876) );
  AND U15312 ( .A(n12878), .B(n12879), .Z(n12727) );
  AND U15313 ( .A(n12880), .B(n12881), .Z(n12879) );
  NAND U15314 ( .A(n8412), .B(\u_a23_core/u_execute/address_plus4[13] ), .Z(
        n12881) );
  NAND U15315 ( .A(\u_a23_core/u_execute/rn[13] ), .B(n8413), .Z(n12880) );
  NAND U15316 ( .A(n12882), .B(n12883), .Z(\u_a23_core/u_execute/rn[13] ) );
  AND U15317 ( .A(n12884), .B(n12885), .Z(n12883) );
  AND U15318 ( .A(n12886), .B(n12887), .Z(n12885) );
  AND U15319 ( .A(n12888), .B(n12889), .Z(n12887) );
  NANDN U15320 ( .B(n8635), .A(\u_a23_core/u_execute/pc[13] ), .Z(n12889) );
  NANDN U15321 ( .B(n8636), .A(\u_a23_core/u_execute/u_register_bank/r14[13] ), 
        .Z(n12888) );
  AND U15322 ( .A(n12890), .B(n12891), .Z(n12886) );
  NANDN U15323 ( .B(n8639), .A(\u_a23_core/u_execute/u_register_bank/r13[13] ), 
        .Z(n12891) );
  NANDN U15324 ( .B(n8640), .A(\u_a23_core/u_execute/u_register_bank/r12[13] ), 
        .Z(n12890) );
  AND U15325 ( .A(n12892), .B(n12893), .Z(n12884) );
  AND U15326 ( .A(n12894), .B(n12895), .Z(n12893) );
  NANDN U15327 ( .B(n8645), .A(\u_a23_core/u_execute/u_register_bank/r11[13] ), 
        .Z(n12895) );
  NANDN U15328 ( .B(n8646), .A(\u_a23_core/u_execute/u_register_bank/r10[13] ), 
        .Z(n12894) );
  AND U15329 ( .A(n12896), .B(n12897), .Z(n12892) );
  NANDN U15330 ( .B(n8649), .A(\u_a23_core/u_execute/u_register_bank/r9[13] ), 
        .Z(n12897) );
  NANDN U15331 ( .B(n8650), .A(\u_a23_core/u_execute/u_register_bank/r8[13] ), 
        .Z(n12896) );
  AND U15332 ( .A(n12898), .B(n12899), .Z(n12882) );
  AND U15333 ( .A(n12900), .B(n12901), .Z(n12899) );
  AND U15334 ( .A(n12902), .B(n12903), .Z(n12901) );
  NANDN U15335 ( .B(n8657), .A(\u_a23_core/u_execute/u_register_bank/r7[13] ), 
        .Z(n12903) );
  NANDN U15336 ( .B(n8658), .A(\u_a23_core/u_execute/u_register_bank/r6[13] ), 
        .Z(n12902) );
  AND U15337 ( .A(n12904), .B(n12905), .Z(n12900) );
  NANDN U15338 ( .B(n8661), .A(\u_a23_core/u_execute/u_register_bank/r5[13] ), 
        .Z(n12905) );
  NANDN U15339 ( .B(n8662), .A(\u_a23_core/u_execute/u_register_bank/r4[13] ), 
        .Z(n12904) );
  AND U15340 ( .A(n12906), .B(n12907), .Z(n12898) );
  AND U15341 ( .A(n12908), .B(n12909), .Z(n12907) );
  NANDN U15342 ( .B(n8667), .A(\u_a23_core/u_execute/u_register_bank/r3[13] ), 
        .Z(n12909) );
  NANDN U15343 ( .B(n8668), .A(\u_a23_core/u_execute/u_register_bank/r0[13] ), 
        .Z(n12908) );
  AND U15344 ( .A(n12910), .B(n12911), .Z(n12906) );
  NANDN U15345 ( .B(n8671), .A(\u_a23_core/u_execute/u_register_bank/r2[13] ), 
        .Z(n12911) );
  NANDN U15346 ( .B(n8672), .A(\u_a23_core/u_execute/u_register_bank/r1[13] ), 
        .Z(n12910) );
  AND U15347 ( .A(n12912), .B(n12913), .Z(n12878) );
  NAND U15348 ( .A(\u_a23_core/u_execute/pc[13] ), .B(n8416), .Z(n12913) );
  NAND U15349 ( .A(n8417), .B(\u_a23_core/u_execute/pc_plus4[13] ), .Z(n12912)
         );
  NAND U15350 ( .A(n12914), .B(n12915), .Z(
        \u_a23_core/execute_address_nxt[12] ) );
  AND U15351 ( .A(n12916), .B(n12917), .Z(n12915) );
  AND U15352 ( .A(n12918), .B(n12919), .Z(n12917) );
  NANDN U15353 ( .B(n8392), .A(\u_a23_core/u_execute/pc_minus4[12] ), .Z(
        n12919) );
  NAND U15354 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[12] ), .B(n8393), 
        .Z(n12918) );
  IV U15355 ( .A(n7045), .Z(\u_a23_core/u_execute/alu_out_pc_filtered[12] ) );
  AND U15356 ( .A(n12920), .B(n12921), .Z(n7045) );
  MUX U15357 ( .IN0(n12922), .IN1(n12923), .SEL(
        \u_a23_core/u_execute/u_alu/b_not[12] ), .F(n12921) );
  NAND U15358 ( .A(n12924), .B(n12925), .Z(
        \u_a23_core/u_execute/u_alu/b_not[12] ) );
  MUX U15359 ( .IN0(n8430), .IN1(n8431), .SEL(n12926), .F(n12925) );
  MUX U15360 ( .IN0(n8433), .IN1(n8434), .SEL(\u_a23_core/u_execute/rn[12] ), 
        .F(n12924) );
  ANDN U15361 ( .A(n8435), .B(n12927), .Z(n12923) );
  MUX U15362 ( .IN0(n8400), .IN1(\u_a23_core/alu_function[3] ), .SEL(
        \u_a23_core/u_execute/u_alu/a[12] ), .F(n12927) );
  NAND U15363 ( .A(\u_a23_core/u_execute/u_alu/a[12] ), .B(n8400), .Z(n12922)
         );
  IV U15364 ( .A(n12928), .Z(\u_a23_core/u_execute/u_alu/a[12] ) );
  MUX U15365 ( .IN0(n12929), .IN1(n12926), .SEL(\u_a23_core/alu_function[8] ), 
        .F(n12928) );
  AND U15366 ( .A(n12930), .B(n12931), .Z(n12926) );
  AND U15367 ( .A(n12932), .B(n12933), .Z(n12931) );
  NAND U15368 ( .A(n12934), .B(n6888), .Z(n12933) );
  NAND U15369 ( .A(n12935), .B(n12936), .Z(n12934) );
  AND U15370 ( .A(n12937), .B(n12938), .Z(n12936) );
  AND U15371 ( .A(n12939), .B(n12940), .Z(n12938) );
  AND U15372 ( .A(n12941), .B(n12942), .Z(n12940) );
  AND U15373 ( .A(n12943), .B(n12944), .Z(n12942) );
  NANDN U15374 ( .B(n8525), .A(n6919), .Z(n12944) );
  NAND U15375 ( .A(n6956), .B(n8512), .Z(n12943) );
  AND U15376 ( .A(n12945), .B(n12946), .Z(n12941) );
  NANDN U15377 ( .B(n8533), .A(n6920), .Z(n12946) );
  NANDN U15378 ( .B(n8516), .A(n6960), .Z(n12945) );
  AND U15379 ( .A(n12947), .B(n12948), .Z(n12939) );
  AND U15380 ( .A(n12949), .B(n12950), .Z(n12948) );
  NANDN U15381 ( .B(n8537), .A(n6925), .Z(n12950) );
  NANDN U15382 ( .B(n8522), .A(n6957), .Z(n12949) );
  AND U15383 ( .A(n12951), .B(n12952), .Z(n12947) );
  NANDN U15384 ( .B(n8538), .A(n6926), .Z(n12952) );
  NANDN U15385 ( .B(n8526), .A(n6947), .Z(n12951) );
  AND U15386 ( .A(n12953), .B(n12954), .Z(n12937) );
  AND U15387 ( .A(n12955), .B(n12956), .Z(n12954) );
  AND U15388 ( .A(n12957), .B(n12958), .Z(n12956) );
  NANDN U15389 ( .B(n8543), .A(n6898), .Z(n12958) );
  NANDN U15390 ( .B(n8534), .A(n6946), .Z(n12957) );
  AND U15391 ( .A(n12959), .B(n12960), .Z(n12955) );
  NANDN U15392 ( .B(n8511), .A(n6943), .Z(n12960) );
  NANDN U15393 ( .B(n8544), .A(n6882), .Z(n12959) );
  AND U15394 ( .A(n12961), .B(n12962), .Z(n12953) );
  AND U15395 ( .A(n12963), .B(n12964), .Z(n12962) );
  NANDN U15396 ( .B(n8515), .A(n6942), .Z(n12964) );
  NANDN U15397 ( .B(n8547), .A(n6809), .Z(n12963) );
  AND U15398 ( .A(n12965), .B(n12966), .Z(n12961) );
  NANDN U15399 ( .B(n8521), .A(n6937), .Z(n12966) );
  NANDN U15400 ( .B(n8548), .A(n6807), .Z(n12965) );
  AND U15401 ( .A(n12967), .B(n12968), .Z(n12935) );
  AND U15402 ( .A(n12969), .B(n12970), .Z(n12968) );
  AND U15403 ( .A(n12971), .B(n12972), .Z(n12970) );
  AND U15404 ( .A(n12973), .B(n12974), .Z(n12972) );
  NANDN U15405 ( .B(n8557), .A(n6799), .Z(n12974) );
  NANDN U15406 ( .B(n8558), .A(n6803), .Z(n12973) );
  AND U15407 ( .A(n12975), .B(n12976), .Z(n12971) );
  NANDN U15408 ( .B(n8561), .A(n6823), .Z(n12976) );
  NANDN U15409 ( .B(n8562), .A(n6827), .Z(n12975) );
  AND U15410 ( .A(n12977), .B(n12978), .Z(n12969) );
  AND U15411 ( .A(n12979), .B(n12980), .Z(n12978) );
  NANDN U15412 ( .B(n8567), .A(n6833), .Z(n12980) );
  NANDN U15413 ( .B(n8568), .A(n6835), .Z(n12979) );
  AND U15414 ( .A(n12981), .B(n12982), .Z(n12977) );
  NANDN U15415 ( .B(n8571), .A(n6839), .Z(n12982) );
  NANDN U15416 ( .B(n8572), .A(n6850), .Z(n12981) );
  AND U15417 ( .A(n12983), .B(n12984), .Z(n12967) );
  AND U15418 ( .A(n12985), .B(n12986), .Z(n12984) );
  AND U15419 ( .A(n12987), .B(n12988), .Z(n12986) );
  NANDN U15420 ( .B(n8579), .A(n6853), .Z(n12988) );
  NANDN U15421 ( .B(n8580), .A(n6841), .Z(n12987) );
  AND U15422 ( .A(n12989), .B(n12990), .Z(n12985) );
  NANDN U15423 ( .B(n8583), .A(n6857), .Z(n12990) );
  NANDN U15424 ( .B(n8584), .A(n6859), .Z(n12989) );
  AND U15425 ( .A(n12991), .B(n12992), .Z(n12983) );
  AND U15426 ( .A(n12993), .B(n12994), .Z(n12992) );
  NANDN U15427 ( .B(n8589), .A(n6865), .Z(n12994) );
  NANDN U15428 ( .B(n8590), .A(n6967), .Z(n12993) );
  AND U15429 ( .A(n12995), .B(n12996), .Z(n12991) );
  NANDN U15430 ( .B(n8593), .A(n6966), .Z(n12996) );
  NAND U15431 ( .A(n6961), .B(n6897), .Z(n12995) );
  AND U15432 ( .A(n12997), .B(n12998), .Z(n12932) );
  NAND U15433 ( .A(n12999), .B(n8452), .Z(n12998) );
  NAND U15434 ( .A(n6856), .B(n6985), .Z(n12997) );
  AND U15435 ( .A(n13000), .B(n13001), .Z(n12930) );
  NAND U15436 ( .A(n8443), .B(n13002), .Z(n13001) );
  NAND U15437 ( .A(n13003), .B(n13004), .Z(n13002) );
  ANDN U15438 ( .A(n13005), .B(n13006), .Z(n13004) );
  NAND U15439 ( .A(n6882), .B(n6856), .Z(n13005) );
  IV U15440 ( .A(n12999), .Z(n13003) );
  NAND U15441 ( .A(n13007), .B(n13008), .Z(n12999) );
  AND U15442 ( .A(n13009), .B(n13010), .Z(n13008) );
  AND U15443 ( .A(n13011), .B(n13012), .Z(n13010) );
  AND U15444 ( .A(n13013), .B(n13014), .Z(n13012) );
  NAND U15445 ( .A(n8461), .B(n6827), .Z(n13014) );
  AND U15446 ( .A(n13015), .B(n13016), .Z(n13013) );
  NAND U15447 ( .A(n8464), .B(n6803), .Z(n13016) );
  NAND U15448 ( .A(n8465), .B(n6823), .Z(n13015) );
  AND U15449 ( .A(n13017), .B(n13018), .Z(n13011) );
  NAND U15450 ( .A(n8470), .B(n6833), .Z(n13018) );
  NAND U15451 ( .A(n9359), .B(n6835), .Z(n13017) );
  AND U15452 ( .A(n13019), .B(n13020), .Z(n13009) );
  AND U15453 ( .A(n13021), .B(n13022), .Z(n13020) );
  NAND U15454 ( .A(n6864), .B(n6807), .Z(n13022) );
  AND U15455 ( .A(n13023), .B(n6935), .Z(n13021) );
  NAND U15456 ( .A(n9726), .B(n6839), .Z(n6935) );
  NAND U15457 ( .A(n6858), .B(n6809), .Z(n13023) );
  AND U15458 ( .A(n10299), .B(n13024), .Z(n13019) );
  NAND U15459 ( .A(n6799), .B(n8487), .Z(n13024) );
  NAND U15460 ( .A(n8606), .B(n6841), .Z(n10299) );
  AND U15461 ( .A(n13025), .B(n13026), .Z(n13007) );
  AND U15462 ( .A(n13027), .B(n13028), .Z(n13026) );
  AND U15463 ( .A(n13029), .B(n10673), .Z(n13028) );
  NAND U15464 ( .A(n8610), .B(n6857), .Z(n10673) );
  AND U15465 ( .A(n9939), .B(n9493), .Z(n13029) );
  NAND U15466 ( .A(n6850), .B(n8603), .Z(n9493) );
  NAND U15467 ( .A(n8609), .B(n6853), .Z(n9939) );
  AND U15468 ( .A(n11414), .B(n11047), .Z(n13027) );
  NAND U15469 ( .A(n8616), .B(n6859), .Z(n11047) );
  NAND U15470 ( .A(n6865), .B(n8958), .Z(n11414) );
  AND U15471 ( .A(n13030), .B(n13031), .Z(n13025) );
  AND U15472 ( .A(n12316), .B(n11602), .Z(n13031) );
  NAND U15473 ( .A(n6967), .B(n9082), .Z(n11602) );
  NAND U15474 ( .A(n6966), .B(n9135), .Z(n12316) );
  AND U15475 ( .A(n13032), .B(n12686), .Z(n13030) );
  NAND U15476 ( .A(n6961), .B(n6984), .Z(n12686) );
  NAND U15477 ( .A(n6956), .B(n6893), .Z(n13032) );
  NAND U15478 ( .A(n13033), .B(n6902), .Z(n13000) );
  NAND U15479 ( .A(n13034), .B(n13035), .Z(n13033) );
  AND U15480 ( .A(n13036), .B(n13037), .Z(n13035) );
  AND U15481 ( .A(n13038), .B(n13039), .Z(n13037) );
  AND U15482 ( .A(n13040), .B(n13041), .Z(n13039) );
  NAND U15483 ( .A(n6956), .B(n6916), .Z(n13041) );
  NAND U15484 ( .A(n8470), .B(n6898), .Z(n13040) );
  AND U15485 ( .A(n13042), .B(n13043), .Z(n13038) );
  NAND U15486 ( .A(n9359), .B(n6926), .Z(n13043) );
  NAND U15487 ( .A(n9726), .B(n6925), .Z(n13042) );
  AND U15488 ( .A(n13044), .B(n13045), .Z(n13036) );
  NAND U15489 ( .A(n8609), .B(n6919), .Z(n13045) );
  AND U15490 ( .A(n13046), .B(n13047), .Z(n13044) );
  NAND U15491 ( .A(n8606), .B(n6937), .Z(n13047) );
  NAND U15492 ( .A(n8603), .B(n6920), .Z(n13046) );
  AND U15493 ( .A(n13048), .B(n13049), .Z(n13034) );
  AND U15494 ( .A(n13050), .B(n13051), .Z(n13049) );
  AND U15495 ( .A(n13052), .B(n13053), .Z(n13050) );
  AND U15496 ( .A(n13054), .B(n13055), .Z(n13048) );
  AND U15497 ( .A(n8742), .B(n9006), .Z(n13054) );
  NAND U15498 ( .A(n9082), .B(n6947), .Z(n9006) );
  NAND U15499 ( .A(n9135), .B(n6957), .Z(n8742) );
  IV U15500 ( .A(\u_a23_core/u_execute/rn[12] ), .Z(n12929) );
  AND U15501 ( .A(n13056), .B(n8620), .Z(n12920) );
  NAND U15502 ( .A(n6765), .B(\u_a23_core/u_execute/u_alu/fadder_out[12] ), 
        .Z(n13056) );
  AND U15503 ( .A(n13057), .B(n13058), .Z(n12916) );
  NANDN U15504 ( .B(n8406), .A(\u_a23_core/u_execute/rn_plus4[12] ), .Z(n13058) );
  NANDN U15505 ( .B(n8407), .A(\u_a23_core/u_execute/alu_plus4[12] ), .Z(
        n13057) );
  AND U15506 ( .A(n13059), .B(n13060), .Z(n12914) );
  AND U15507 ( .A(n13061), .B(n13062), .Z(n13060) );
  NAND U15508 ( .A(n8412), .B(\u_a23_core/u_execute/address_plus4[12] ), .Z(
        n13062) );
  NAND U15509 ( .A(\u_a23_core/u_execute/rn[12] ), .B(n8413), .Z(n13061) );
  NAND U15510 ( .A(n13063), .B(n13064), .Z(\u_a23_core/u_execute/rn[12] ) );
  AND U15511 ( .A(n13065), .B(n13066), .Z(n13064) );
  AND U15512 ( .A(n13067), .B(n13068), .Z(n13066) );
  AND U15513 ( .A(n13069), .B(n13070), .Z(n13068) );
  NANDN U15514 ( .B(n8635), .A(\u_a23_core/u_execute/pc[12] ), .Z(n13070) );
  NANDN U15515 ( .B(n8636), .A(\u_a23_core/u_execute/u_register_bank/r14[12] ), 
        .Z(n13069) );
  AND U15516 ( .A(n13071), .B(n13072), .Z(n13067) );
  NANDN U15517 ( .B(n8639), .A(\u_a23_core/u_execute/u_register_bank/r13[12] ), 
        .Z(n13072) );
  NANDN U15518 ( .B(n8640), .A(\u_a23_core/u_execute/u_register_bank/r12[12] ), 
        .Z(n13071) );
  AND U15519 ( .A(n13073), .B(n13074), .Z(n13065) );
  AND U15520 ( .A(n13075), .B(n13076), .Z(n13074) );
  NANDN U15521 ( .B(n8645), .A(\u_a23_core/u_execute/u_register_bank/r11[12] ), 
        .Z(n13076) );
  NANDN U15522 ( .B(n8646), .A(\u_a23_core/u_execute/u_register_bank/r10[12] ), 
        .Z(n13075) );
  AND U15523 ( .A(n13077), .B(n13078), .Z(n13073) );
  NANDN U15524 ( .B(n8649), .A(\u_a23_core/u_execute/u_register_bank/r9[12] ), 
        .Z(n13078) );
  NANDN U15525 ( .B(n8650), .A(\u_a23_core/u_execute/u_register_bank/r8[12] ), 
        .Z(n13077) );
  AND U15526 ( .A(n13079), .B(n13080), .Z(n13063) );
  AND U15527 ( .A(n13081), .B(n13082), .Z(n13080) );
  AND U15528 ( .A(n13083), .B(n13084), .Z(n13082) );
  NANDN U15529 ( .B(n8657), .A(\u_a23_core/u_execute/u_register_bank/r7[12] ), 
        .Z(n13084) );
  NANDN U15530 ( .B(n8658), .A(\u_a23_core/u_execute/u_register_bank/r6[12] ), 
        .Z(n13083) );
  AND U15531 ( .A(n13085), .B(n13086), .Z(n13081) );
  NANDN U15532 ( .B(n8661), .A(\u_a23_core/u_execute/u_register_bank/r5[12] ), 
        .Z(n13086) );
  NANDN U15533 ( .B(n8662), .A(\u_a23_core/u_execute/u_register_bank/r4[12] ), 
        .Z(n13085) );
  AND U15534 ( .A(n13087), .B(n13088), .Z(n13079) );
  AND U15535 ( .A(n13089), .B(n13090), .Z(n13088) );
  NANDN U15536 ( .B(n8667), .A(\u_a23_core/u_execute/u_register_bank/r3[12] ), 
        .Z(n13090) );
  NANDN U15537 ( .B(n8668), .A(\u_a23_core/u_execute/u_register_bank/r0[12] ), 
        .Z(n13089) );
  AND U15538 ( .A(n13091), .B(n13092), .Z(n13087) );
  NANDN U15539 ( .B(n8671), .A(\u_a23_core/u_execute/u_register_bank/r2[12] ), 
        .Z(n13092) );
  NANDN U15540 ( .B(n8672), .A(\u_a23_core/u_execute/u_register_bank/r1[12] ), 
        .Z(n13091) );
  AND U15541 ( .A(n13093), .B(n13094), .Z(n13059) );
  NAND U15542 ( .A(\u_a23_core/u_execute/pc[12] ), .B(n8416), .Z(n13094) );
  NAND U15543 ( .A(n8417), .B(\u_a23_core/u_execute/pc_plus4[12] ), .Z(n13093)
         );
  AND U15544 ( .A(n13095), .B(n13096), .Z(n11457) );
  AND U15545 ( .A(n13097), .B(n13098), .Z(n13096) );
  NOR U15546 ( .A(\u_a23_core/execute_address_nxt[10] ), .B(
        \u_a23_core/execute_address_nxt[11] ), .Z(n13098) );
  NAND U15547 ( .A(n13099), .B(n13100), .Z(
        \u_a23_core/execute_address_nxt[11] ) );
  AND U15548 ( .A(n13101), .B(n13102), .Z(n13100) );
  AND U15549 ( .A(n13103), .B(n13104), .Z(n13102) );
  NANDN U15550 ( .B(n8392), .A(\u_a23_core/u_execute/pc_minus4[11] ), .Z(
        n13104) );
  NAND U15551 ( .A(n8393), .B(\u_a23_core/u_execute/alu_out_pc_filtered[11] ), 
        .Z(n13103) );
  IV U15552 ( .A(n7046), .Z(\u_a23_core/u_execute/alu_out_pc_filtered[11] ) );
  AND U15553 ( .A(n13105), .B(n13106), .Z(n7046) );
  MUX U15554 ( .IN0(n13107), .IN1(n13108), .SEL(
        \u_a23_core/u_execute/u_alu/b_not[11] ), .F(n13106) );
  NAND U15555 ( .A(n13109), .B(n13110), .Z(
        \u_a23_core/u_execute/u_alu/b_not[11] ) );
  MUX U15556 ( .IN0(n8430), .IN1(n8431), .SEL(n13111), .F(n13110) );
  MUX U15557 ( .IN0(n8433), .IN1(n8434), .SEL(\u_a23_core/u_execute/rn[11] ), 
        .F(n13109) );
  ANDN U15558 ( .A(n8435), .B(n13112), .Z(n13108) );
  MUX U15559 ( .IN0(n8400), .IN1(\u_a23_core/alu_function[3] ), .SEL(
        \u_a23_core/u_execute/u_alu/a[11] ), .F(n13112) );
  NAND U15560 ( .A(\u_a23_core/u_execute/u_alu/a[11] ), .B(n8400), .Z(n13107)
         );
  IV U15561 ( .A(n13113), .Z(\u_a23_core/u_execute/u_alu/a[11] ) );
  MUX U15562 ( .IN0(n13114), .IN1(n13111), .SEL(\u_a23_core/alu_function[8] ), 
        .F(n13113) );
  AND U15563 ( .A(n13115), .B(n13116), .Z(n13111) );
  AND U15564 ( .A(n13117), .B(n13118), .Z(n13116) );
  NAND U15565 ( .A(n6840), .B(n6985), .Z(n13118) );
  AND U15566 ( .A(n13119), .B(n13120), .Z(n13117) );
  NAND U15567 ( .A(n8443), .B(n13121), .Z(n13120) );
  NANDN U15568 ( .B(n13006), .A(n13122), .Z(n13121) );
  NAND U15569 ( .A(n13123), .B(n13124), .Z(n13006) );
  NAND U15570 ( .A(n6882), .B(n13125), .Z(n13123) );
  NAND U15571 ( .A(n13126), .B(n13127), .Z(n13125) );
  AND U15572 ( .A(n12590), .B(n12594), .Z(n13127) );
  IV U15573 ( .A(n6840), .Z(n12594) );
  ANDN U15574 ( .A(n8449), .B(n13128), .Z(n13126) );
  NANDN U15575 ( .B(n13122), .A(n8452), .Z(n13119) );
  AND U15576 ( .A(n13129), .B(n13130), .Z(n13122) );
  AND U15577 ( .A(n13131), .B(n13132), .Z(n13130) );
  AND U15578 ( .A(n13133), .B(n13134), .Z(n13132) );
  AND U15579 ( .A(n13135), .B(n13136), .Z(n13134) );
  NAND U15580 ( .A(n8461), .B(n6833), .Z(n13136) );
  AND U15581 ( .A(n13137), .B(n13138), .Z(n13135) );
  NAND U15582 ( .A(n8464), .B(n6823), .Z(n13138) );
  NAND U15583 ( .A(n8465), .B(n6827), .Z(n13137) );
  AND U15584 ( .A(n13139), .B(n13140), .Z(n13133) );
  NAND U15585 ( .A(n8470), .B(n6835), .Z(n13140) );
  NAND U15586 ( .A(n9359), .B(n6839), .Z(n13139) );
  AND U15587 ( .A(n13141), .B(n13142), .Z(n13131) );
  AND U15588 ( .A(n13143), .B(n13144), .Z(n13142) );
  NAND U15589 ( .A(n6858), .B(n6807), .Z(n13144) );
  AND U15590 ( .A(n13145), .B(n9363), .Z(n13143) );
  NAND U15591 ( .A(n6850), .B(n9726), .Z(n9363) );
  NAND U15592 ( .A(n6856), .B(n6809), .Z(n13145) );
  AND U15593 ( .A(n13146), .B(n13147), .Z(n13141) );
  NAND U15594 ( .A(n6864), .B(n6799), .Z(n13147) );
  NAND U15595 ( .A(n6803), .B(n8487), .Z(n13146) );
  AND U15596 ( .A(n13148), .B(n13149), .Z(n13129) );
  AND U15597 ( .A(n13150), .B(n13151), .Z(n13149) );
  AND U15598 ( .A(n13152), .B(n10121), .Z(n13151) );
  NAND U15599 ( .A(n8609), .B(n6841), .Z(n10121) );
  AND U15600 ( .A(n9747), .B(n10480), .Z(n13152) );
  NAND U15601 ( .A(n8606), .B(n6857), .Z(n10480) );
  NAND U15602 ( .A(n8603), .B(n6853), .Z(n9747) );
  AND U15603 ( .A(n11228), .B(n10862), .Z(n13150) );
  NAND U15604 ( .A(n8610), .B(n6859), .Z(n10862) );
  NAND U15605 ( .A(n6865), .B(n8616), .Z(n11228) );
  AND U15606 ( .A(n13153), .B(n13154), .Z(n13148) );
  AND U15607 ( .A(n13155), .B(n12500), .Z(n13154) );
  NAND U15608 ( .A(n6961), .B(n9135), .Z(n12500) );
  AND U15609 ( .A(n12134), .B(n11789), .Z(n13155) );
  NAND U15610 ( .A(n6967), .B(n8958), .Z(n11789) );
  NAND U15611 ( .A(n6966), .B(n9082), .Z(n12134) );
  AND U15612 ( .A(n13156), .B(n12873), .Z(n13153) );
  NAND U15613 ( .A(n6956), .B(n6984), .Z(n12873) );
  NAND U15614 ( .A(n6893), .B(n6960), .Z(n13156) );
  AND U15615 ( .A(n13157), .B(n13158), .Z(n13115) );
  NAND U15616 ( .A(n13159), .B(n6888), .Z(n13158) );
  NAND U15617 ( .A(n13160), .B(n13161), .Z(n13159) );
  AND U15618 ( .A(n13162), .B(n13163), .Z(n13161) );
  AND U15619 ( .A(n13164), .B(n13165), .Z(n13163) );
  AND U15620 ( .A(n13166), .B(n13167), .Z(n13165) );
  AND U15621 ( .A(n13168), .B(n13169), .Z(n13167) );
  NANDN U15622 ( .B(n8521), .A(n6919), .Z(n13169) );
  NAND U15623 ( .A(n6960), .B(n8512), .Z(n13168) );
  AND U15624 ( .A(n13170), .B(n13171), .Z(n13166) );
  NANDN U15625 ( .B(n8525), .A(n6920), .Z(n13171) );
  NANDN U15626 ( .B(n8516), .A(n6957), .Z(n13170) );
  AND U15627 ( .A(n13172), .B(n13173), .Z(n13164) );
  AND U15628 ( .A(n13174), .B(n13175), .Z(n13173) );
  NANDN U15629 ( .B(n8533), .A(n6925), .Z(n13175) );
  NANDN U15630 ( .B(n8522), .A(n6947), .Z(n13174) );
  AND U15631 ( .A(n13176), .B(n13177), .Z(n13172) );
  NANDN U15632 ( .B(n8537), .A(n6926), .Z(n13177) );
  NANDN U15633 ( .B(n8526), .A(n6946), .Z(n13176) );
  AND U15634 ( .A(n13178), .B(n13179), .Z(n13162) );
  AND U15635 ( .A(n13180), .B(n13181), .Z(n13179) );
  AND U15636 ( .A(n13182), .B(n13183), .Z(n13181) );
  NANDN U15637 ( .B(n8538), .A(n6898), .Z(n13183) );
  NANDN U15638 ( .B(n8534), .A(n6943), .Z(n13182) );
  AND U15639 ( .A(n13184), .B(n13185), .Z(n13180) );
  NANDN U15640 ( .B(n8511), .A(n6942), .Z(n13185) );
  NANDN U15641 ( .B(n8543), .A(n6882), .Z(n13184) );
  AND U15642 ( .A(n13186), .B(n13187), .Z(n13178) );
  AND U15643 ( .A(n13188), .B(n13189), .Z(n13187) );
  NANDN U15644 ( .B(n8515), .A(n6937), .Z(n13189) );
  NANDN U15645 ( .B(n8544), .A(n6809), .Z(n13188) );
  AND U15646 ( .A(n13190), .B(n13191), .Z(n13186) );
  NANDN U15647 ( .B(n8547), .A(n6807), .Z(n13191) );
  NANDN U15648 ( .B(n8548), .A(n6799), .Z(n13190) );
  AND U15649 ( .A(n13192), .B(n13193), .Z(n13160) );
  AND U15650 ( .A(n13194), .B(n13195), .Z(n13193) );
  AND U15651 ( .A(n13196), .B(n13197), .Z(n13195) );
  AND U15652 ( .A(n13198), .B(n13199), .Z(n13197) );
  NANDN U15653 ( .B(n8557), .A(n6803), .Z(n13199) );
  NANDN U15654 ( .B(n8558), .A(n6823), .Z(n13198) );
  AND U15655 ( .A(n13200), .B(n13201), .Z(n13196) );
  NANDN U15656 ( .B(n8561), .A(n6827), .Z(n13201) );
  NANDN U15657 ( .B(n8562), .A(n6833), .Z(n13200) );
  AND U15658 ( .A(n13202), .B(n13203), .Z(n13194) );
  AND U15659 ( .A(n13204), .B(n13205), .Z(n13203) );
  NANDN U15660 ( .B(n8567), .A(n6835), .Z(n13205) );
  NANDN U15661 ( .B(n8568), .A(n6839), .Z(n13204) );
  AND U15662 ( .A(n13206), .B(n13207), .Z(n13202) );
  NANDN U15663 ( .B(n8571), .A(n6850), .Z(n13207) );
  NANDN U15664 ( .B(n8572), .A(n6853), .Z(n13206) );
  AND U15665 ( .A(n13208), .B(n13209), .Z(n13192) );
  AND U15666 ( .A(n13210), .B(n13211), .Z(n13209) );
  AND U15667 ( .A(n13212), .B(n13213), .Z(n13211) );
  NANDN U15668 ( .B(n8579), .A(n6841), .Z(n13213) );
  NANDN U15669 ( .B(n8580), .A(n6857), .Z(n13212) );
  AND U15670 ( .A(n13214), .B(n13215), .Z(n13210) );
  NANDN U15671 ( .B(n8583), .A(n6859), .Z(n13215) );
  NANDN U15672 ( .B(n8584), .A(n6865), .Z(n13214) );
  AND U15673 ( .A(n13216), .B(n13217), .Z(n13208) );
  AND U15674 ( .A(n13218), .B(n13219), .Z(n13217) );
  NANDN U15675 ( .B(n8589), .A(n6967), .Z(n13219) );
  NANDN U15676 ( .B(n8590), .A(n6966), .Z(n13218) );
  AND U15677 ( .A(n13220), .B(n13221), .Z(n13216) );
  NANDN U15678 ( .B(n8593), .A(n6961), .Z(n13221) );
  NAND U15679 ( .A(n6956), .B(n6897), .Z(n13220) );
  NAND U15680 ( .A(n13222), .B(n6902), .Z(n13157) );
  NAND U15681 ( .A(n13223), .B(n13224), .Z(n13222) );
  AND U15682 ( .A(n13225), .B(n13226), .Z(n13224) );
  AND U15683 ( .A(n13227), .B(n13228), .Z(n13226) );
  NAND U15684 ( .A(n9726), .B(n6926), .Z(n13228) );
  AND U15685 ( .A(n13229), .B(n13230), .Z(n13227) );
  NAND U15686 ( .A(n6916), .B(n6960), .Z(n13230) );
  NAND U15687 ( .A(n9359), .B(n6898), .Z(n13229) );
  AND U15688 ( .A(n13231), .B(n13232), .Z(n13225) );
  NAND U15689 ( .A(n8609), .B(n6920), .Z(n13232) );
  AND U15690 ( .A(n13233), .B(n13234), .Z(n13231) );
  NAND U15691 ( .A(n8606), .B(n6919), .Z(n13234) );
  NAND U15692 ( .A(n8603), .B(n6925), .Z(n13233) );
  AND U15693 ( .A(n13235), .B(n13236), .Z(n13223) );
  AND U15694 ( .A(n13237), .B(n13238), .Z(n13236) );
  AND U15695 ( .A(n11900), .B(n6872), .Z(n13237) );
  NAND U15696 ( .A(n8610), .B(n6937), .Z(n6872) );
  NAND U15697 ( .A(n8616), .B(n6942), .Z(n11900) );
  AND U15698 ( .A(n13239), .B(n8499), .Z(n13235) );
  NAND U15699 ( .A(n6984), .B(n6957), .Z(n8499) );
  AND U15700 ( .A(n13240), .B(n9129), .Z(n13239) );
  NAND U15701 ( .A(n9082), .B(n6946), .Z(n9129) );
  IV U15702 ( .A(\u_a23_core/u_execute/rn[11] ), .Z(n13114) );
  AND U15703 ( .A(n13241), .B(n8620), .Z(n13105) );
  NAND U15704 ( .A(n6765), .B(\u_a23_core/u_execute/u_alu/fadder_out[11] ), 
        .Z(n13241) );
  AND U15705 ( .A(n13242), .B(n13243), .Z(n13101) );
  NANDN U15706 ( .B(n8406), .A(\u_a23_core/u_execute/rn_plus4[11] ), .Z(n13243) );
  NANDN U15707 ( .B(n8407), .A(\u_a23_core/u_execute/alu_plus4[11] ), .Z(
        n13242) );
  AND U15708 ( .A(n13244), .B(n13245), .Z(n13099) );
  AND U15709 ( .A(n13246), .B(n13247), .Z(n13245) );
  NAND U15710 ( .A(n8412), .B(\u_a23_core/u_execute/address_plus4[11] ), .Z(
        n13247) );
  NAND U15711 ( .A(\u_a23_core/u_execute/rn[11] ), .B(n8413), .Z(n13246) );
  NAND U15712 ( .A(n13248), .B(n13249), .Z(\u_a23_core/u_execute/rn[11] ) );
  AND U15713 ( .A(n13250), .B(n13251), .Z(n13249) );
  AND U15714 ( .A(n13252), .B(n13253), .Z(n13251) );
  AND U15715 ( .A(n13254), .B(n13255), .Z(n13253) );
  NANDN U15716 ( .B(n8635), .A(\u_a23_core/u_execute/pc[11] ), .Z(n13255) );
  NANDN U15717 ( .B(n8636), .A(\u_a23_core/u_execute/u_register_bank/r14[11] ), 
        .Z(n13254) );
  AND U15718 ( .A(n13256), .B(n13257), .Z(n13252) );
  NANDN U15719 ( .B(n8639), .A(\u_a23_core/u_execute/u_register_bank/r13[11] ), 
        .Z(n13257) );
  NANDN U15720 ( .B(n8640), .A(\u_a23_core/u_execute/u_register_bank/r12[11] ), 
        .Z(n13256) );
  AND U15721 ( .A(n13258), .B(n13259), .Z(n13250) );
  AND U15722 ( .A(n13260), .B(n13261), .Z(n13259) );
  NANDN U15723 ( .B(n8645), .A(\u_a23_core/u_execute/u_register_bank/r11[11] ), 
        .Z(n13261) );
  NANDN U15724 ( .B(n8646), .A(\u_a23_core/u_execute/u_register_bank/r10[11] ), 
        .Z(n13260) );
  AND U15725 ( .A(n13262), .B(n13263), .Z(n13258) );
  NANDN U15726 ( .B(n8649), .A(\u_a23_core/u_execute/u_register_bank/r9[11] ), 
        .Z(n13263) );
  NANDN U15727 ( .B(n8650), .A(\u_a23_core/u_execute/u_register_bank/r8[11] ), 
        .Z(n13262) );
  AND U15728 ( .A(n13264), .B(n13265), .Z(n13248) );
  AND U15729 ( .A(n13266), .B(n13267), .Z(n13265) );
  AND U15730 ( .A(n13268), .B(n13269), .Z(n13267) );
  NANDN U15731 ( .B(n8657), .A(\u_a23_core/u_execute/u_register_bank/r7[11] ), 
        .Z(n13269) );
  NANDN U15732 ( .B(n8658), .A(\u_a23_core/u_execute/u_register_bank/r6[11] ), 
        .Z(n13268) );
  AND U15733 ( .A(n13270), .B(n13271), .Z(n13266) );
  NANDN U15734 ( .B(n8661), .A(\u_a23_core/u_execute/u_register_bank/r5[11] ), 
        .Z(n13271) );
  NANDN U15735 ( .B(n8662), .A(\u_a23_core/u_execute/u_register_bank/r4[11] ), 
        .Z(n13270) );
  AND U15736 ( .A(n13272), .B(n13273), .Z(n13264) );
  AND U15737 ( .A(n13274), .B(n13275), .Z(n13273) );
  NANDN U15738 ( .B(n8667), .A(\u_a23_core/u_execute/u_register_bank/r3[11] ), 
        .Z(n13275) );
  NANDN U15739 ( .B(n8668), .A(\u_a23_core/u_execute/u_register_bank/r0[11] ), 
        .Z(n13274) );
  AND U15740 ( .A(n13276), .B(n13277), .Z(n13272) );
  NANDN U15741 ( .B(n8671), .A(\u_a23_core/u_execute/u_register_bank/r2[11] ), 
        .Z(n13277) );
  NANDN U15742 ( .B(n8672), .A(\u_a23_core/u_execute/u_register_bank/r1[11] ), 
        .Z(n13276) );
  AND U15743 ( .A(n13278), .B(n13279), .Z(n13244) );
  NAND U15744 ( .A(\u_a23_core/u_execute/pc[11] ), .B(n8416), .Z(n13279) );
  NAND U15745 ( .A(n8417), .B(\u_a23_core/u_execute/pc_plus4[11] ), .Z(n13278)
         );
  NAND U15746 ( .A(n13280), .B(n13281), .Z(
        \u_a23_core/execute_address_nxt[10] ) );
  AND U15747 ( .A(n13282), .B(n13283), .Z(n13281) );
  AND U15748 ( .A(n13284), .B(n13285), .Z(n13283) );
  NANDN U15749 ( .B(n8392), .A(\u_a23_core/u_execute/pc_minus4[10] ), .Z(
        n13285) );
  NAND U15750 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[10] ), .B(n8393), 
        .Z(n13284) );
  IV U15751 ( .A(n7047), .Z(\u_a23_core/u_execute/alu_out_pc_filtered[10] ) );
  AND U15752 ( .A(n13286), .B(n13287), .Z(n7047) );
  MUX U15753 ( .IN0(n13288), .IN1(n13289), .SEL(
        \u_a23_core/u_execute/u_alu/b_not[10] ), .F(n13287) );
  NAND U15754 ( .A(n13290), .B(n13291), .Z(
        \u_a23_core/u_execute/u_alu/b_not[10] ) );
  MUX U15755 ( .IN0(n8430), .IN1(n8431), .SEL(n13292), .F(n13291) );
  MUX U15756 ( .IN0(n8433), .IN1(n8434), .SEL(\u_a23_core/u_execute/rn[10] ), 
        .F(n13290) );
  ANDN U15757 ( .A(n8435), .B(n13293), .Z(n13289) );
  MUX U15758 ( .IN0(n8400), .IN1(\u_a23_core/alu_function[3] ), .SEL(
        \u_a23_core/u_execute/u_alu/a[10] ), .F(n13293) );
  AND U15759 ( .A(n13294), .B(n13295), .Z(n8435) );
  AND U15760 ( .A(n13296), .B(n13297), .Z(n13294) );
  NAND U15761 ( .A(\u_a23_core/u_execute/u_alu/a[10] ), .B(n8400), .Z(n13288)
         );
  IV U15762 ( .A(n13298), .Z(\u_a23_core/u_execute/u_alu/a[10] ) );
  MUX U15763 ( .IN0(n13299), .IN1(n13292), .SEL(\u_a23_core/alu_function[8] ), 
        .F(n13298) );
  AND U15764 ( .A(n13300), .B(n13301), .Z(n13292) );
  AND U15765 ( .A(n13302), .B(n13303), .Z(n13301) );
  NAND U15766 ( .A(n6886), .B(n13304), .Z(n13303) );
  NAND U15767 ( .A(n8449), .B(n12220), .Z(n13304) );
  ANDN U15768 ( .A(n13305), .B(n13128), .Z(n12220) );
  AND U15769 ( .A(n13306), .B(n13307), .Z(n13305) );
  ANDN U15770 ( .A(n13308), .B(n6851), .Z(n8449) );
  AND U15771 ( .A(n13309), .B(n8696), .Z(n13308) );
  IV U15772 ( .A(n6834), .Z(n8696) );
  IV U15773 ( .A(n6838), .Z(n13309) );
  NAND U15774 ( .A(n6786), .B(n13310), .Z(n13302) );
  NAND U15775 ( .A(n13311), .B(n13312), .Z(n13310) );
  AND U15776 ( .A(n13313), .B(n13314), .Z(n13312) );
  AND U15777 ( .A(n13315), .B(n13316), .Z(n13314) );
  AND U15778 ( .A(n13317), .B(n13318), .Z(n13316) );
  NAND U15779 ( .A(n8464), .B(n6827), .Z(n13318) );
  ANDN U15780 ( .A(n9457), .B(n6915), .Z(n13317) );
  ANDN U15781 ( .A(n9359), .B(n13319), .Z(n6915) );
  IV U15782 ( .A(n6850), .Z(n13319) );
  NAND U15783 ( .A(n9726), .B(n6853), .Z(n9457) );
  AND U15784 ( .A(n13320), .B(n13321), .Z(n13315) );
  NAND U15785 ( .A(n8470), .B(n6839), .Z(n13321) );
  AND U15786 ( .A(n13322), .B(n13323), .Z(n13320) );
  NAND U15787 ( .A(n8465), .B(n6833), .Z(n13323) );
  NAND U15788 ( .A(n8461), .B(n6835), .Z(n13322) );
  AND U15789 ( .A(n13324), .B(n13325), .Z(n13313) );
  AND U15790 ( .A(n13326), .B(n13327), .Z(n13325) );
  NAND U15791 ( .A(n6856), .B(n6807), .Z(n13327) );
  AND U15792 ( .A(n13328), .B(n13329), .Z(n13326) );
  NAND U15793 ( .A(n6840), .B(n6809), .Z(n13329) );
  NAND U15794 ( .A(n6882), .B(n6852), .Z(n13328) );
  AND U15795 ( .A(n13330), .B(n13331), .Z(n13324) );
  NAND U15796 ( .A(n6858), .B(n6799), .Z(n13331) );
  NAND U15797 ( .A(n6864), .B(n6803), .Z(n13330) );
  AND U15798 ( .A(n13332), .B(n13333), .Z(n13311) );
  AND U15799 ( .A(n13334), .B(n13335), .Z(n13333) );
  AND U15800 ( .A(n13336), .B(n9931), .Z(n13335) );
  NAND U15801 ( .A(n8603), .B(n6841), .Z(n9931) );
  AND U15802 ( .A(n10665), .B(n13337), .Z(n13336) );
  NAND U15803 ( .A(n6823), .B(n8487), .Z(n13337) );
  NAND U15804 ( .A(n8606), .B(n6859), .Z(n10665) );
  AND U15805 ( .A(n13338), .B(n11415), .Z(n13334) );
  NAND U15806 ( .A(n6967), .B(n8616), .Z(n11415) );
  AND U15807 ( .A(n11039), .B(n10298), .Z(n13338) );
  NAND U15808 ( .A(n8609), .B(n6857), .Z(n10298) );
  NAND U15809 ( .A(n6865), .B(n8610), .Z(n11039) );
  AND U15810 ( .A(n13339), .B(n13340), .Z(n13332) );
  AND U15811 ( .A(n13341), .B(n12687), .Z(n13340) );
  NAND U15812 ( .A(n6956), .B(n9135), .Z(n12687) );
  AND U15813 ( .A(n12314), .B(n11603), .Z(n13341) );
  NAND U15814 ( .A(n6966), .B(n8958), .Z(n11603) );
  NAND U15815 ( .A(n6961), .B(n9082), .Z(n12314) );
  AND U15816 ( .A(n13342), .B(n13055), .Z(n13339) );
  NAND U15817 ( .A(n6984), .B(n6960), .Z(n13055) );
  NAND U15818 ( .A(n6893), .B(n6957), .Z(n13342) );
  AND U15819 ( .A(n13343), .B(n13344), .Z(n13300) );
  NAND U15820 ( .A(n13345), .B(n6888), .Z(n13344) );
  NAND U15821 ( .A(n13346), .B(n13347), .Z(n13345) );
  AND U15822 ( .A(n13348), .B(n13349), .Z(n13347) );
  AND U15823 ( .A(n13350), .B(n13351), .Z(n13349) );
  AND U15824 ( .A(n13352), .B(n13353), .Z(n13351) );
  AND U15825 ( .A(n13354), .B(n13355), .Z(n13353) );
  NANDN U15826 ( .B(n8515), .A(n6919), .Z(n13355) );
  NAND U15827 ( .A(n6957), .B(n8512), .Z(n13354) );
  AND U15828 ( .A(n13356), .B(n13357), .Z(n13352) );
  NANDN U15829 ( .B(n8521), .A(n6920), .Z(n13357) );
  NANDN U15830 ( .B(n8516), .A(n6947), .Z(n13356) );
  AND U15831 ( .A(n13358), .B(n13359), .Z(n13350) );
  AND U15832 ( .A(n13360), .B(n13361), .Z(n13359) );
  NANDN U15833 ( .B(n8525), .A(n6925), .Z(n13361) );
  NANDN U15834 ( .B(n8522), .A(n6946), .Z(n13360) );
  AND U15835 ( .A(n13362), .B(n13363), .Z(n13358) );
  NANDN U15836 ( .B(n8533), .A(n6926), .Z(n13363) );
  NANDN U15837 ( .B(n8526), .A(n6943), .Z(n13362) );
  AND U15838 ( .A(n13364), .B(n13365), .Z(n13348) );
  AND U15839 ( .A(n13366), .B(n13367), .Z(n13365) );
  AND U15840 ( .A(n13368), .B(n13369), .Z(n13367) );
  NANDN U15841 ( .B(n8537), .A(n6898), .Z(n13369) );
  NANDN U15842 ( .B(n8534), .A(n6942), .Z(n13368) );
  AND U15843 ( .A(n13370), .B(n13371), .Z(n13366) );
  NANDN U15844 ( .B(n8511), .A(n6937), .Z(n13371) );
  NANDN U15845 ( .B(n8538), .A(n6882), .Z(n13370) );
  AND U15846 ( .A(n13372), .B(n13373), .Z(n13364) );
  AND U15847 ( .A(n13374), .B(n13375), .Z(n13373) );
  NANDN U15848 ( .B(n8543), .A(n6809), .Z(n13375) );
  NANDN U15849 ( .B(n8544), .A(n6807), .Z(n13374) );
  AND U15850 ( .A(n13376), .B(n13377), .Z(n13372) );
  NANDN U15851 ( .B(n8547), .A(n6799), .Z(n13377) );
  NANDN U15852 ( .B(n8548), .A(n6803), .Z(n13376) );
  AND U15853 ( .A(n13378), .B(n13379), .Z(n13346) );
  AND U15854 ( .A(n13380), .B(n13381), .Z(n13379) );
  AND U15855 ( .A(n13382), .B(n13383), .Z(n13381) );
  AND U15856 ( .A(n13384), .B(n13385), .Z(n13383) );
  NANDN U15857 ( .B(n8557), .A(n6823), .Z(n13385) );
  NANDN U15858 ( .B(n8558), .A(n6827), .Z(n13384) );
  AND U15859 ( .A(n13386), .B(n13387), .Z(n13382) );
  NANDN U15860 ( .B(n8561), .A(n6833), .Z(n13387) );
  NANDN U15861 ( .B(n8562), .A(n6835), .Z(n13386) );
  AND U15862 ( .A(n13388), .B(n13389), .Z(n13380) );
  AND U15863 ( .A(n13390), .B(n13391), .Z(n13389) );
  NANDN U15864 ( .B(n8567), .A(n6839), .Z(n13391) );
  NANDN U15865 ( .B(n8568), .A(n6850), .Z(n13390) );
  AND U15866 ( .A(n13392), .B(n13393), .Z(n13388) );
  NANDN U15867 ( .B(n8571), .A(n6853), .Z(n13393) );
  NANDN U15868 ( .B(n8572), .A(n6841), .Z(n13392) );
  AND U15869 ( .A(n13394), .B(n13395), .Z(n13378) );
  AND U15870 ( .A(n13396), .B(n13397), .Z(n13395) );
  AND U15871 ( .A(n13398), .B(n13399), .Z(n13397) );
  NANDN U15872 ( .B(n8579), .A(n6857), .Z(n13399) );
  NANDN U15873 ( .B(n8580), .A(n6859), .Z(n13398) );
  AND U15874 ( .A(n13400), .B(n13401), .Z(n13396) );
  NANDN U15875 ( .B(n8583), .A(n6865), .Z(n13401) );
  NANDN U15876 ( .B(n8584), .A(n6967), .Z(n13400) );
  AND U15877 ( .A(n13402), .B(n13403), .Z(n13394) );
  AND U15878 ( .A(n13404), .B(n13405), .Z(n13403) );
  NANDN U15879 ( .B(n8589), .A(n6966), .Z(n13405) );
  NANDN U15880 ( .B(n8590), .A(n6961), .Z(n13404) );
  AND U15881 ( .A(n13406), .B(n13407), .Z(n13402) );
  NANDN U15882 ( .B(n8593), .A(n6956), .Z(n13407) );
  NAND U15883 ( .A(n6960), .B(n6897), .Z(n13406) );
  NAND U15884 ( .A(n13408), .B(n6902), .Z(n13343) );
  NAND U15885 ( .A(n13409), .B(n13410), .Z(n13408) );
  AND U15886 ( .A(n13411), .B(n13412), .Z(n13410) );
  AND U15887 ( .A(n13413), .B(n13414), .Z(n13412) );
  NAND U15888 ( .A(n8606), .B(n6920), .Z(n13414) );
  AND U15889 ( .A(n13415), .B(n13416), .Z(n13413) );
  NAND U15890 ( .A(n6916), .B(n6957), .Z(n13416) );
  NAND U15891 ( .A(n9726), .B(n6898), .Z(n13415) );
  AND U15892 ( .A(n13417), .B(n13418), .Z(n13411) );
  NAND U15893 ( .A(n8610), .B(n6919), .Z(n13418) );
  AND U15894 ( .A(n13419), .B(n13420), .Z(n13417) );
  NAND U15895 ( .A(n8603), .B(n6926), .Z(n13420) );
  NAND U15896 ( .A(n8609), .B(n6925), .Z(n13419) );
  AND U15897 ( .A(n13421), .B(n13422), .Z(n13409) );
  AND U15898 ( .A(n13423), .B(n13424), .Z(n13422) );
  AND U15899 ( .A(n13425), .B(n13426), .Z(n13423) );
  AND U15900 ( .A(n8741), .B(n9011), .Z(n13421) );
  NAND U15901 ( .A(n9135), .B(n6946), .Z(n9011) );
  NAND U15902 ( .A(n6984), .B(n6947), .Z(n8741) );
  IV U15903 ( .A(\u_a23_core/u_execute/rn[10] ), .Z(n13299) );
  AND U15904 ( .A(n13427), .B(n8620), .Z(n13286) );
  IV U15905 ( .A(n12319), .Z(n8620) );
  ANDN U15906 ( .A(\u_a23_core/u_execute/u_alu/b_not[7] ), .B(n13428), .Z(
        n12319) );
  NAND U15907 ( .A(n13429), .B(n13430), .Z(
        \u_a23_core/u_execute/u_alu/b_not[7] ) );
  MUX U15908 ( .IN0(n8430), .IN1(n8431), .SEL(n8403), .F(n13430) );
  AND U15909 ( .A(n13431), .B(n13432), .Z(n8403) );
  AND U15910 ( .A(n13433), .B(n13434), .Z(n13432) );
  NAND U15911 ( .A(n6886), .B(n13128), .Z(n13434) );
  NANDN U15912 ( .B(n6826), .A(n12756), .Z(n13128) );
  NOR U15913 ( .A(n6832), .B(n6822), .Z(n12756) );
  AND U15914 ( .A(n13435), .B(n13436), .Z(n13433) );
  NAND U15915 ( .A(n6786), .B(n13437), .Z(n13435) );
  NAND U15916 ( .A(n13438), .B(n13439), .Z(n13437) );
  AND U15917 ( .A(n13440), .B(n13441), .Z(n13439) );
  AND U15918 ( .A(n13442), .B(n13443), .Z(n13441) );
  AND U15919 ( .A(n13444), .B(n13445), .Z(n13443) );
  ANDN U15920 ( .A(n11765), .B(n11201), .Z(n13445) );
  ANDN U15921 ( .A(n8606), .B(n11386), .Z(n11201) );
  IV U15922 ( .A(n6966), .Z(n11386) );
  NAND U15923 ( .A(n6961), .B(n8610), .Z(n11765) );
  ANDN U15924 ( .A(n10832), .B(n10454), .Z(n13444) );
  ANDN U15925 ( .A(n8603), .B(n10639), .Z(n10454) );
  IV U15926 ( .A(n6865), .Z(n10639) );
  NAND U15927 ( .A(n6967), .B(n8609), .Z(n10832) );
  AND U15928 ( .A(n13446), .B(n13447), .Z(n13442) );
  NAND U15929 ( .A(n8461), .B(n6853), .Z(n13447) );
  AND U15930 ( .A(n13448), .B(n13449), .Z(n13446) );
  NAND U15931 ( .A(n8464), .B(n6839), .Z(n13449) );
  NAND U15932 ( .A(n6850), .B(n8465), .Z(n13448) );
  AND U15933 ( .A(n13450), .B(n13451), .Z(n13440) );
  AND U15934 ( .A(n13452), .B(n10096), .Z(n13451) );
  NAND U15935 ( .A(n9726), .B(n6859), .Z(n10096) );
  AND U15936 ( .A(n9725), .B(n9357), .Z(n13452) );
  NAND U15937 ( .A(n8470), .B(n6841), .Z(n9357) );
  NAND U15938 ( .A(n9359), .B(n6857), .Z(n9725) );
  AND U15939 ( .A(n13453), .B(n13454), .Z(n13450) );
  NAND U15940 ( .A(n6840), .B(n6803), .Z(n13454) );
  AND U15941 ( .A(n13455), .B(n13456), .Z(n13453) );
  NAND U15942 ( .A(n6882), .B(n6834), .Z(n13456) );
  NAND U15943 ( .A(n6838), .B(n6809), .Z(n13455) );
  AND U15944 ( .A(n13457), .B(n13458), .Z(n13438) );
  AND U15945 ( .A(n13459), .B(n13460), .Z(n13458) );
  AND U15946 ( .A(n13461), .B(n13462), .Z(n13460) );
  NAND U15947 ( .A(n6856), .B(n6823), .Z(n13462) );
  AND U15948 ( .A(n13463), .B(n13464), .Z(n13461) );
  NAND U15949 ( .A(n6807), .B(n6851), .Z(n13464) );
  NAND U15950 ( .A(n6852), .B(n6799), .Z(n13463) );
  AND U15951 ( .A(n13465), .B(n13466), .Z(n13459) );
  NAND U15952 ( .A(n6835), .B(n8487), .Z(n13466) );
  AND U15953 ( .A(n13467), .B(n13468), .Z(n13465) );
  NAND U15954 ( .A(n6858), .B(n6827), .Z(n13468) );
  NAND U15955 ( .A(n6864), .B(n6833), .Z(n13467) );
  AND U15956 ( .A(n13469), .B(n13470), .Z(n13457) );
  AND U15957 ( .A(n13471), .B(n12874), .Z(n13470) );
  NAND U15958 ( .A(n9082), .B(n6957), .Z(n12874) );
  AND U15959 ( .A(n12498), .B(n12131), .Z(n13471) );
  NAND U15960 ( .A(n6956), .B(n8616), .Z(n12131) );
  NAND U15961 ( .A(n8958), .B(n6960), .Z(n12498) );
  AND U15962 ( .A(n13472), .B(n13473), .Z(n13469) );
  NAND U15963 ( .A(n6893), .B(n6943), .Z(n13473) );
  AND U15964 ( .A(n8617), .B(n13240), .Z(n13472) );
  NAND U15965 ( .A(n9135), .B(n6947), .Z(n13240) );
  NAND U15966 ( .A(n6984), .B(n6946), .Z(n8617) );
  AND U15967 ( .A(n13474), .B(n13475), .Z(n13431) );
  NAND U15968 ( .A(n13476), .B(n6888), .Z(n13475) );
  NAND U15969 ( .A(n13477), .B(n13478), .Z(n13476) );
  AND U15970 ( .A(n13479), .B(n13480), .Z(n13478) );
  AND U15971 ( .A(n13481), .B(n13482), .Z(n13480) );
  AND U15972 ( .A(n13483), .B(n13484), .Z(n13482) );
  AND U15973 ( .A(n13485), .B(n13486), .Z(n13484) );
  NANDN U15974 ( .B(n8526), .A(n6919), .Z(n13486) );
  NAND U15975 ( .A(n6943), .B(n8512), .Z(n13485) );
  AND U15976 ( .A(n13487), .B(n13488), .Z(n13483) );
  NANDN U15977 ( .B(n8534), .A(n6920), .Z(n13488) );
  NANDN U15978 ( .B(n8516), .A(n6942), .Z(n13487) );
  AND U15979 ( .A(n13489), .B(n13490), .Z(n13481) );
  AND U15980 ( .A(n13491), .B(n13492), .Z(n13490) );
  NANDN U15981 ( .B(n8511), .A(n6925), .Z(n13492) );
  NANDN U15982 ( .B(n8522), .A(n6937), .Z(n13491) );
  AND U15983 ( .A(n13493), .B(n13494), .Z(n13489) );
  NANDN U15984 ( .B(n8515), .A(n6926), .Z(n13494) );
  NANDN U15985 ( .B(n8521), .A(n6898), .Z(n13493) );
  AND U15986 ( .A(n13495), .B(n13496), .Z(n13479) );
  AND U15987 ( .A(n13497), .B(n13498), .Z(n13496) );
  AND U15988 ( .A(n13499), .B(n13500), .Z(n13498) );
  NANDN U15989 ( .B(n8525), .A(n6882), .Z(n13500) );
  NANDN U15990 ( .B(n8533), .A(n6809), .Z(n13499) );
  AND U15991 ( .A(n13501), .B(n13502), .Z(n13497) );
  NANDN U15992 ( .B(n8537), .A(n6807), .Z(n13502) );
  NANDN U15993 ( .B(n8538), .A(n6799), .Z(n13501) );
  AND U15994 ( .A(n13503), .B(n13504), .Z(n13495) );
  AND U15995 ( .A(n13505), .B(n13506), .Z(n13504) );
  NANDN U15996 ( .B(n8543), .A(n6803), .Z(n13506) );
  NANDN U15997 ( .B(n8544), .A(n6823), .Z(n13505) );
  AND U15998 ( .A(n13507), .B(n13508), .Z(n13503) );
  NANDN U15999 ( .B(n8547), .A(n6827), .Z(n13508) );
  NANDN U16000 ( .B(n8548), .A(n6833), .Z(n13507) );
  AND U16001 ( .A(n13509), .B(n13510), .Z(n13477) );
  AND U16002 ( .A(n13511), .B(n13512), .Z(n13510) );
  AND U16003 ( .A(n13513), .B(n13514), .Z(n13512) );
  AND U16004 ( .A(n13515), .B(n13516), .Z(n13514) );
  NANDN U16005 ( .B(n8557), .A(n6835), .Z(n13516) );
  NANDN U16006 ( .B(n8558), .A(n6839), .Z(n13515) );
  AND U16007 ( .A(n13517), .B(n13518), .Z(n13513) );
  NANDN U16008 ( .B(n8561), .A(n6850), .Z(n13518) );
  NANDN U16009 ( .B(n8562), .A(n6853), .Z(n13517) );
  AND U16010 ( .A(n13519), .B(n13520), .Z(n13511) );
  AND U16011 ( .A(n13521), .B(n13522), .Z(n13520) );
  NANDN U16012 ( .B(n8567), .A(n6841), .Z(n13522) );
  NANDN U16013 ( .B(n8568), .A(n6857), .Z(n13521) );
  AND U16014 ( .A(n13523), .B(n13524), .Z(n13519) );
  NANDN U16015 ( .B(n8571), .A(n6859), .Z(n13524) );
  NANDN U16016 ( .B(n8572), .A(n6865), .Z(n13523) );
  AND U16017 ( .A(n13525), .B(n13526), .Z(n13509) );
  AND U16018 ( .A(n13527), .B(n13528), .Z(n13526) );
  AND U16019 ( .A(n13529), .B(n13530), .Z(n13528) );
  NANDN U16020 ( .B(n8579), .A(n6967), .Z(n13530) );
  NANDN U16021 ( .B(n8580), .A(n6966), .Z(n13529) );
  AND U16022 ( .A(n13531), .B(n13532), .Z(n13527) );
  NANDN U16023 ( .B(n8583), .A(n6961), .Z(n13532) );
  NANDN U16024 ( .B(n8584), .A(n6956), .Z(n13531) );
  AND U16025 ( .A(n13533), .B(n13534), .Z(n13525) );
  AND U16026 ( .A(n13535), .B(n13536), .Z(n13534) );
  NANDN U16027 ( .B(n8589), .A(n6960), .Z(n13536) );
  NANDN U16028 ( .B(n8590), .A(n6957), .Z(n13535) );
  AND U16029 ( .A(n13537), .B(n13538), .Z(n13533) );
  NANDN U16030 ( .B(n8593), .A(n6947), .Z(n13538) );
  NAND U16031 ( .A(n6946), .B(n6897), .Z(n13537) );
  NAND U16032 ( .A(n13539), .B(n6902), .Z(n13474) );
  NAND U16033 ( .A(n13540), .B(n13541), .Z(n13539) );
  AND U16034 ( .A(n13542), .B(n13543), .Z(n13541) );
  AND U16035 ( .A(n13544), .B(n13545), .Z(n13543) );
  NAND U16036 ( .A(n6943), .B(n6916), .Z(n13545) );
  NAND U16037 ( .A(n8606), .B(n6898), .Z(n13544) );
  AND U16038 ( .A(n13546), .B(n13547), .Z(n13542) );
  NAND U16039 ( .A(n8610), .B(n6926), .Z(n13547) );
  NAND U16040 ( .A(n8616), .B(n6925), .Z(n13546) );
  AND U16041 ( .A(n13548), .B(n13549), .Z(n13540) );
  AND U16042 ( .A(n11902), .B(n6874), .Z(n13549) );
  NAND U16043 ( .A(n8958), .B(n6920), .Z(n6874) );
  NAND U16044 ( .A(n9082), .B(n6919), .Z(n11902) );
  AND U16045 ( .A(n9134), .B(n13550), .Z(n13548) );
  NAND U16046 ( .A(n6984), .B(n6942), .Z(n9134) );
  MUX U16047 ( .IN0(n8433), .IN1(n8434), .SEL(\u_a23_core/u_execute/rn[7] ), 
        .F(n13429) );
  NAND U16048 ( .A(n13551), .B(n13552), .Z(\u_a23_core/u_execute/rn[7] ) );
  AND U16049 ( .A(n13553), .B(n13554), .Z(n13552) );
  AND U16050 ( .A(n13555), .B(n13556), .Z(n13554) );
  AND U16051 ( .A(n13557), .B(n13558), .Z(n13556) );
  NANDN U16052 ( .B(n8635), .A(\u_a23_core/u_execute/pc[7] ), .Z(n13558) );
  NANDN U16053 ( .B(n8636), .A(\u_a23_core/u_execute/u_register_bank/r14[7] ), 
        .Z(n13557) );
  AND U16054 ( .A(n13559), .B(n13560), .Z(n13555) );
  NANDN U16055 ( .B(n8639), .A(\u_a23_core/u_execute/u_register_bank/r13[7] ), 
        .Z(n13560) );
  NANDN U16056 ( .B(n8640), .A(\u_a23_core/u_execute/u_register_bank/r12[7] ), 
        .Z(n13559) );
  AND U16057 ( .A(n13561), .B(n13562), .Z(n13553) );
  AND U16058 ( .A(n13563), .B(n13564), .Z(n13562) );
  NANDN U16059 ( .B(n8645), .A(\u_a23_core/u_execute/u_register_bank/r11[7] ), 
        .Z(n13564) );
  NANDN U16060 ( .B(n8646), .A(\u_a23_core/u_execute/u_register_bank/r10[7] ), 
        .Z(n13563) );
  AND U16061 ( .A(n13565), .B(n13566), .Z(n13561) );
  NANDN U16062 ( .B(n8649), .A(\u_a23_core/u_execute/u_register_bank/r9[7] ), 
        .Z(n13566) );
  NANDN U16063 ( .B(n8650), .A(\u_a23_core/u_execute/u_register_bank/r8[7] ), 
        .Z(n13565) );
  AND U16064 ( .A(n13567), .B(n13568), .Z(n13551) );
  AND U16065 ( .A(n13569), .B(n13570), .Z(n13568) );
  AND U16066 ( .A(n13571), .B(n13572), .Z(n13570) );
  NANDN U16067 ( .B(n8657), .A(\u_a23_core/u_execute/u_register_bank/r7[7] ), 
        .Z(n13572) );
  NANDN U16068 ( .B(n8658), .A(\u_a23_core/u_execute/u_register_bank/r6[7] ), 
        .Z(n13571) );
  AND U16069 ( .A(n13573), .B(n13574), .Z(n13569) );
  NANDN U16070 ( .B(n8661), .A(\u_a23_core/u_execute/u_register_bank/r5[7] ), 
        .Z(n13574) );
  NANDN U16071 ( .B(n8662), .A(\u_a23_core/u_execute/u_register_bank/r4[7] ), 
        .Z(n13573) );
  AND U16072 ( .A(n13575), .B(n13576), .Z(n13567) );
  AND U16073 ( .A(n13577), .B(n13578), .Z(n13576) );
  NANDN U16074 ( .B(n8667), .A(\u_a23_core/u_execute/u_register_bank/r3[7] ), 
        .Z(n13578) );
  NANDN U16075 ( .B(n8668), .A(\u_a23_core/u_execute/u_register_bank/r0[7] ), 
        .Z(n13577) );
  AND U16076 ( .A(n13579), .B(n13580), .Z(n13575) );
  NANDN U16077 ( .B(n8671), .A(\u_a23_core/u_execute/u_register_bank/r2[7] ), 
        .Z(n13580) );
  NANDN U16078 ( .B(n8672), .A(\u_a23_core/u_execute/u_register_bank/r1[7] ), 
        .Z(n13579) );
  NAND U16079 ( .A(n6765), .B(\u_a23_core/u_execute/u_alu/fadder_out[10] ), 
        .Z(n13427) );
  AND U16080 ( .A(n13581), .B(n13582), .Z(n13282) );
  NANDN U16081 ( .B(n8406), .A(\u_a23_core/u_execute/rn_plus4[10] ), .Z(n13582) );
  NANDN U16082 ( .B(n8407), .A(\u_a23_core/u_execute/alu_plus4[10] ), .Z(
        n13581) );
  AND U16083 ( .A(n13583), .B(n13584), .Z(n13280) );
  AND U16084 ( .A(n13585), .B(n13586), .Z(n13584) );
  NAND U16085 ( .A(n8412), .B(\u_a23_core/u_execute/address_plus4[10] ), .Z(
        n13586) );
  NAND U16086 ( .A(\u_a23_core/u_execute/rn[10] ), .B(n8413), .Z(n13585) );
  NAND U16087 ( .A(n13587), .B(n13588), .Z(\u_a23_core/u_execute/rn[10] ) );
  AND U16088 ( .A(n13589), .B(n13590), .Z(n13588) );
  AND U16089 ( .A(n13591), .B(n13592), .Z(n13590) );
  AND U16090 ( .A(n13593), .B(n13594), .Z(n13592) );
  NANDN U16091 ( .B(n8635), .A(\u_a23_core/u_execute/pc[10] ), .Z(n13594) );
  NANDN U16092 ( .B(n8636), .A(\u_a23_core/u_execute/u_register_bank/r14[10] ), 
        .Z(n13593) );
  AND U16093 ( .A(n13595), .B(n13596), .Z(n13591) );
  NANDN U16094 ( .B(n8639), .A(\u_a23_core/u_execute/u_register_bank/r13[10] ), 
        .Z(n13596) );
  NANDN U16095 ( .B(n8640), .A(\u_a23_core/u_execute/u_register_bank/r12[10] ), 
        .Z(n13595) );
  AND U16096 ( .A(n13597), .B(n13598), .Z(n13589) );
  AND U16097 ( .A(n13599), .B(n13600), .Z(n13598) );
  NANDN U16098 ( .B(n8645), .A(\u_a23_core/u_execute/u_register_bank/r11[10] ), 
        .Z(n13600) );
  NANDN U16099 ( .B(n8646), .A(\u_a23_core/u_execute/u_register_bank/r10[10] ), 
        .Z(n13599) );
  AND U16100 ( .A(n13601), .B(n13602), .Z(n13597) );
  NANDN U16101 ( .B(n8649), .A(\u_a23_core/u_execute/u_register_bank/r9[10] ), 
        .Z(n13602) );
  NANDN U16102 ( .B(n8650), .A(\u_a23_core/u_execute/u_register_bank/r8[10] ), 
        .Z(n13601) );
  AND U16103 ( .A(n13603), .B(n13604), .Z(n13587) );
  AND U16104 ( .A(n13605), .B(n13606), .Z(n13604) );
  AND U16105 ( .A(n13607), .B(n13608), .Z(n13606) );
  NANDN U16106 ( .B(n8657), .A(\u_a23_core/u_execute/u_register_bank/r7[10] ), 
        .Z(n13608) );
  NANDN U16107 ( .B(n8658), .A(\u_a23_core/u_execute/u_register_bank/r6[10] ), 
        .Z(n13607) );
  AND U16108 ( .A(n13609), .B(n13610), .Z(n13605) );
  NANDN U16109 ( .B(n8661), .A(\u_a23_core/u_execute/u_register_bank/r5[10] ), 
        .Z(n13610) );
  NANDN U16110 ( .B(n8662), .A(\u_a23_core/u_execute/u_register_bank/r4[10] ), 
        .Z(n13609) );
  AND U16111 ( .A(n13611), .B(n13612), .Z(n13603) );
  AND U16112 ( .A(n13613), .B(n13614), .Z(n13612) );
  NANDN U16113 ( .B(n8667), .A(\u_a23_core/u_execute/u_register_bank/r3[10] ), 
        .Z(n13614) );
  NANDN U16114 ( .B(n8668), .A(\u_a23_core/u_execute/u_register_bank/r0[10] ), 
        .Z(n13613) );
  AND U16115 ( .A(n13615), .B(n13616), .Z(n13611) );
  NANDN U16116 ( .B(n8671), .A(\u_a23_core/u_execute/u_register_bank/r2[10] ), 
        .Z(n13616) );
  NANDN U16117 ( .B(n8672), .A(\u_a23_core/u_execute/u_register_bank/r1[10] ), 
        .Z(n13615) );
  AND U16118 ( .A(n13617), .B(n13618), .Z(n13583) );
  NAND U16119 ( .A(\u_a23_core/u_execute/pc[10] ), .B(n8416), .Z(n13618) );
  NAND U16120 ( .A(n8417), .B(\u_a23_core/u_execute/pc_plus4[10] ), .Z(n13617)
         );
  AND U16121 ( .A(n879), .B(n7100), .Z(n13097) );
  IV U16122 ( .A(\u_a23_core/execute_address_nxt[0] ), .Z(n7100) );
  NAND U16123 ( .A(n13619), .B(n13620), .Z(\u_a23_core/execute_address_nxt[0] ) );
  NAND U16124 ( .A(n8412), .B(\u_a23_core/u_execute/address_plus4[0] ), .Z(
        n13620) );
  AND U16125 ( .A(n13621), .B(n13622), .Z(n13619) );
  OR U16126 ( .A(n11835), .B(n6340), .Z(n13622) );
  AND U16127 ( .A(n13623), .B(n13624), .Z(n6340) );
  MUX U16128 ( .IN0(n13625), .IN1(n13626), .SEL(
        \u_a23_core/u_execute/u_alu/b_not[0] ), .F(n13624) );
  OR U16129 ( .A(n13627), .B(n13628), .Z(\u_a23_core/u_execute/u_alu/b_not[0] ) );
  MUX U16130 ( .IN0(n13629), .IN1(n13630), .SEL(n13631), .F(n13628) );
  MUX U16131 ( .IN0(n13632), .IN1(n13633), .SEL(n13634), .F(n13627) );
  ANDN U16132 ( .A(n8398), .B(n13635), .Z(n13626) );
  MUX U16133 ( .IN0(n8400), .IN1(\u_a23_core/alu_function[3] ), .SEL(
        \u_a23_core/u_execute/u_alu/a[0] ), .F(n13635) );
  NAND U16134 ( .A(\u_a23_core/u_execute/u_alu/a[0] ), .B(n8400), .Z(n13625)
         );
  IV U16135 ( .A(n13636), .Z(\u_a23_core/u_execute/u_alu/a[0] ) );
  MUX U16136 ( .IN0(n13634), .IN1(n13631), .SEL(\u_a23_core/alu_function[8] ), 
        .F(n13636) );
  AND U16137 ( .A(n13637), .B(n13638), .Z(n13631) );
  AND U16138 ( .A(n13639), .B(n13640), .Z(n13638) );
  NAND U16139 ( .A(n6985), .B(n6808), .Z(n13640) );
  AND U16140 ( .A(n11848), .B(n13641), .Z(n13639) );
  NAND U16141 ( .A(n13642), .B(n6902), .Z(n13641) );
  AND U16142 ( .A(n6898), .B(n6916), .Z(n13642) );
  OR U16143 ( .A(n12758), .B(n9262), .Z(n11848) );
  ANDN U16144 ( .A(n13643), .B(\u_a23_core/shift_imm_zero ), .Z(n12758) );
  AND U16145 ( .A(n13644), .B(n13645), .Z(n13637) );
  NAND U16146 ( .A(n6786), .B(n13646), .Z(n13645) );
  NAND U16147 ( .A(n13647), .B(n13648), .Z(n13646) );
  AND U16148 ( .A(n13649), .B(n13650), .Z(n13648) );
  AND U16149 ( .A(n13651), .B(n13652), .Z(n13650) );
  AND U16150 ( .A(n13653), .B(n13654), .Z(n13652) );
  AND U16151 ( .A(n13655), .B(n13656), .Z(n13654) );
  NAND U16152 ( .A(n6802), .B(n6799), .Z(n13656) );
  NAND U16153 ( .A(n6807), .B(n6798), .Z(n13655) );
  AND U16154 ( .A(n9463), .B(n13657), .Z(n13653) );
  NAND U16155 ( .A(n6806), .B(n6809), .Z(n13657) );
  NAND U16156 ( .A(n6967), .B(n8464), .Z(n9463) );
  AND U16157 ( .A(n13658), .B(n13659), .Z(n13651) );
  AND U16158 ( .A(n10275), .B(n9902), .Z(n13659) );
  NAND U16159 ( .A(n6966), .B(n8465), .Z(n9902) );
  NAND U16160 ( .A(n6961), .B(n8461), .Z(n10275) );
  AND U16161 ( .A(n13660), .B(n10643), .Z(n13658) );
  NAND U16162 ( .A(n6956), .B(n8470), .Z(n10643) );
  NAND U16163 ( .A(n6803), .B(n6822), .Z(n13660) );
  AND U16164 ( .A(n13661), .B(n13662), .Z(n13649) );
  AND U16165 ( .A(n13663), .B(n13664), .Z(n13662) );
  AND U16166 ( .A(n11395), .B(n11024), .Z(n13664) );
  NAND U16167 ( .A(n9359), .B(n6960), .Z(n11024) );
  NAND U16168 ( .A(n9726), .B(n6957), .Z(n11395) );
  AND U16169 ( .A(n13665), .B(n13666), .Z(n13663) );
  NAND U16170 ( .A(n6823), .B(n6826), .Z(n13666) );
  NAND U16171 ( .A(n6832), .B(n6827), .Z(n13665) );
  AND U16172 ( .A(n13667), .B(n13668), .Z(n13661) );
  AND U16173 ( .A(n13669), .B(n13670), .Z(n13668) );
  NAND U16174 ( .A(n6834), .B(n6833), .Z(n13670) );
  NAND U16175 ( .A(n6838), .B(n6835), .Z(n13669) );
  AND U16176 ( .A(n13671), .B(n13672), .Z(n13667) );
  NAND U16177 ( .A(n6840), .B(n6853), .Z(n13672) );
  NAND U16178 ( .A(n6839), .B(n6851), .Z(n13671) );
  AND U16179 ( .A(n13673), .B(n13674), .Z(n13647) );
  AND U16180 ( .A(n13675), .B(n13676), .Z(n13674) );
  AND U16181 ( .A(n13677), .B(n13678), .Z(n13676) );
  AND U16182 ( .A(n13679), .B(n13680), .Z(n13678) );
  NAND U16183 ( .A(n6850), .B(n6852), .Z(n13680) );
  NAND U16184 ( .A(n6856), .B(n6841), .Z(n13679) );
  AND U16185 ( .A(n13681), .B(n13682), .Z(n13677) );
  NAND U16186 ( .A(n6858), .B(n6857), .Z(n13682) );
  NAND U16187 ( .A(n6864), .B(n6859), .Z(n13681) );
  AND U16188 ( .A(n13683), .B(n13684), .Z(n13675) );
  AND U16189 ( .A(n12677), .B(n6969), .Z(n13684) );
  NAND U16190 ( .A(n6865), .B(n8487), .Z(n6969) );
  NAND U16191 ( .A(n8606), .B(n6943), .Z(n12677) );
  AND U16192 ( .A(n12309), .B(n11596), .Z(n13683) );
  NAND U16193 ( .A(n8603), .B(n6947), .Z(n11596) );
  NAND U16194 ( .A(n8609), .B(n6946), .Z(n12309) );
  AND U16195 ( .A(n13685), .B(n13686), .Z(n13673) );
  AND U16196 ( .A(n13687), .B(n13688), .Z(n13686) );
  AND U16197 ( .A(n13426), .B(n13053), .Z(n13688) );
  NAND U16198 ( .A(n8610), .B(n6942), .Z(n13053) );
  NAND U16199 ( .A(n8616), .B(n6937), .Z(n13426) );
  AND U16200 ( .A(n8962), .B(n8822), .Z(n13687) );
  NAND U16201 ( .A(n8958), .B(n6919), .Z(n8822) );
  NAND U16202 ( .A(n9082), .B(n6920), .Z(n8962) );
  AND U16203 ( .A(n13689), .B(n13690), .Z(n13685) );
  NAND U16204 ( .A(n6893), .B(n6898), .Z(n13690) );
  AND U16205 ( .A(n13691), .B(n13692), .Z(n13689) );
  NAND U16206 ( .A(n13693), .B(n6888), .Z(n13644) );
  NAND U16207 ( .A(n13694), .B(n13695), .Z(n13693) );
  AND U16208 ( .A(n13696), .B(n13697), .Z(n13695) );
  AND U16209 ( .A(n13698), .B(n13699), .Z(n13697) );
  AND U16210 ( .A(n13700), .B(n13701), .Z(n13699) );
  AND U16211 ( .A(n13702), .B(n13703), .Z(n13701) );
  NANDN U16212 ( .B(n8589), .A(n6919), .Z(n13703) );
  NAND U16213 ( .A(n8512), .B(n6898), .Z(n13702) );
  AND U16214 ( .A(n13704), .B(n13705), .Z(n13700) );
  NANDN U16215 ( .B(n8590), .A(n6920), .Z(n13705) );
  NANDN U16216 ( .B(n8516), .A(n6882), .Z(n13704) );
  AND U16217 ( .A(n13706), .B(n13707), .Z(n13698) );
  AND U16218 ( .A(n13708), .B(n13709), .Z(n13707) );
  NANDN U16219 ( .B(n8593), .A(n6925), .Z(n13709) );
  NANDN U16220 ( .B(n8522), .A(n6809), .Z(n13708) );
  AND U16221 ( .A(n13710), .B(n13711), .Z(n13706) );
  NAND U16222 ( .A(n6926), .B(n6897), .Z(n13711) );
  NANDN U16223 ( .B(n8526), .A(n6807), .Z(n13710) );
  AND U16224 ( .A(n13712), .B(n13713), .Z(n13696) );
  AND U16225 ( .A(n13714), .B(n13715), .Z(n13713) );
  AND U16226 ( .A(n13716), .B(n13717), .Z(n13715) );
  NANDN U16227 ( .B(n8534), .A(n6799), .Z(n13717) );
  NANDN U16228 ( .B(n8511), .A(n6803), .Z(n13716) );
  AND U16229 ( .A(n13718), .B(n13719), .Z(n13714) );
  NANDN U16230 ( .B(n8515), .A(n6823), .Z(n13719) );
  NANDN U16231 ( .B(n8521), .A(n6827), .Z(n13718) );
  AND U16232 ( .A(n13720), .B(n13721), .Z(n13712) );
  AND U16233 ( .A(n13722), .B(n13723), .Z(n13721) );
  NANDN U16234 ( .B(n8525), .A(n6833), .Z(n13723) );
  NANDN U16235 ( .B(n8533), .A(n6835), .Z(n13722) );
  AND U16236 ( .A(n13724), .B(n13725), .Z(n13720) );
  NANDN U16237 ( .B(n8537), .A(n6839), .Z(n13725) );
  NANDN U16238 ( .B(n8538), .A(n6850), .Z(n13724) );
  AND U16239 ( .A(n13726), .B(n13727), .Z(n13694) );
  AND U16240 ( .A(n13728), .B(n13729), .Z(n13727) );
  AND U16241 ( .A(n13730), .B(n13731), .Z(n13729) );
  AND U16242 ( .A(n13732), .B(n13733), .Z(n13731) );
  NANDN U16243 ( .B(n8543), .A(n6853), .Z(n13733) );
  NANDN U16244 ( .B(n8544), .A(n6841), .Z(n13732) );
  AND U16245 ( .A(n13734), .B(n13735), .Z(n13730) );
  NANDN U16246 ( .B(n8547), .A(n6857), .Z(n13735) );
  NANDN U16247 ( .B(n8548), .A(n6859), .Z(n13734) );
  AND U16248 ( .A(n13736), .B(n13737), .Z(n13728) );
  AND U16249 ( .A(n13738), .B(n13739), .Z(n13737) );
  NANDN U16250 ( .B(n8557), .A(n6865), .Z(n13739) );
  NANDN U16251 ( .B(n8558), .A(n6967), .Z(n13738) );
  AND U16252 ( .A(n13740), .B(n13741), .Z(n13736) );
  NANDN U16253 ( .B(n8561), .A(n6966), .Z(n13741) );
  NANDN U16254 ( .B(n8562), .A(n6961), .Z(n13740) );
  AND U16255 ( .A(n13742), .B(n13743), .Z(n13726) );
  AND U16256 ( .A(n13744), .B(n13745), .Z(n13743) );
  AND U16257 ( .A(n13746), .B(n13747), .Z(n13745) );
  NANDN U16258 ( .B(n8567), .A(n6956), .Z(n13747) );
  NANDN U16259 ( .B(n8568), .A(n6960), .Z(n13746) );
  AND U16260 ( .A(n13748), .B(n13749), .Z(n13744) );
  NANDN U16261 ( .B(n8571), .A(n6957), .Z(n13749) );
  NANDN U16262 ( .B(n8572), .A(n6947), .Z(n13748) );
  AND U16263 ( .A(n13750), .B(n13751), .Z(n13742) );
  AND U16264 ( .A(n13752), .B(n13753), .Z(n13751) );
  NANDN U16265 ( .B(n8579), .A(n6946), .Z(n13753) );
  NANDN U16266 ( .B(n8580), .A(n6943), .Z(n13752) );
  AND U16267 ( .A(n13754), .B(n13755), .Z(n13750) );
  NANDN U16268 ( .B(n8583), .A(n6942), .Z(n13755) );
  NANDN U16269 ( .B(n8584), .A(n6937), .Z(n13754) );
  NAND U16270 ( .A(n6765), .B(\u_a23_core/u_execute/u_alu/fadder_out[0] ), .Z(
        n13623) );
  ANDN U16271 ( .A(n8407), .B(n9248), .Z(n11835) );
  AND U16272 ( .A(n13756), .B(n8393), .Z(n9248) );
  NAND U16273 ( .A(n13757), .B(\u_a23_core/pc_wen ), .Z(n13756) );
  ANDN U16274 ( .A(\u_a23_core/pc_sel[0] ), .B(\u_a23_core/pc_sel[1] ), .Z(
        n13757) );
  OR U16275 ( .A(n11969), .B(n13634), .Z(n13621) );
  AND U16276 ( .A(n13758), .B(n13759), .Z(n13634) );
  AND U16277 ( .A(n13760), .B(n13761), .Z(n13759) );
  AND U16278 ( .A(n13762), .B(n13763), .Z(n13761) );
  AND U16279 ( .A(n13764), .B(n13765), .Z(n13763) );
  NANDN U16280 ( .B(n8636), .A(\u_a23_core/u_execute/u_register_bank/r14[0] ), 
        .Z(n13765) );
  NANDN U16281 ( .B(n8639), .A(\u_a23_core/u_execute/u_register_bank/r13[0] ), 
        .Z(n13764) );
  AND U16282 ( .A(n13766), .B(n13767), .Z(n13762) );
  NANDN U16283 ( .B(n8640), .A(\u_a23_core/u_execute/u_register_bank/r12[0] ), 
        .Z(n13767) );
  NANDN U16284 ( .B(n8645), .A(\u_a23_core/u_execute/u_register_bank/r11[0] ), 
        .Z(n13766) );
  AND U16285 ( .A(n13768), .B(n13769), .Z(n13760) );
  AND U16286 ( .A(n13770), .B(n13771), .Z(n13769) );
  NANDN U16287 ( .B(n8646), .A(\u_a23_core/u_execute/u_register_bank/r10[0] ), 
        .Z(n13771) );
  NANDN U16288 ( .B(n8649), .A(\u_a23_core/u_execute/u_register_bank/r9[0] ), 
        .Z(n13770) );
  AND U16289 ( .A(n13772), .B(n13773), .Z(n13768) );
  NANDN U16290 ( .B(n8650), .A(\u_a23_core/u_execute/u_register_bank/r8[0] ), 
        .Z(n13773) );
  NANDN U16291 ( .B(n8657), .A(\u_a23_core/u_execute/u_register_bank/r7[0] ), 
        .Z(n13772) );
  AND U16292 ( .A(n13774), .B(n13775), .Z(n13758) );
  AND U16293 ( .A(n13776), .B(n13777), .Z(n13775) );
  AND U16294 ( .A(n13778), .B(n13779), .Z(n13777) );
  NANDN U16295 ( .B(n8658), .A(\u_a23_core/u_execute/u_register_bank/r6[0] ), 
        .Z(n13779) );
  NANDN U16296 ( .B(n8661), .A(\u_a23_core/u_execute/u_register_bank/r5[0] ), 
        .Z(n13778) );
  AND U16297 ( .A(n13780), .B(n13781), .Z(n13776) );
  NANDN U16298 ( .B(n8662), .A(\u_a23_core/u_execute/u_register_bank/r4[0] ), 
        .Z(n13781) );
  NANDN U16299 ( .B(n8667), .A(\u_a23_core/u_execute/u_register_bank/r3[0] ), 
        .Z(n13780) );
  AND U16300 ( .A(n13782), .B(n13783), .Z(n13774) );
  NANDN U16301 ( .B(n8672), .A(\u_a23_core/u_execute/u_register_bank/r1[0] ), 
        .Z(n13783) );
  AND U16302 ( .A(n13784), .B(n13785), .Z(n13782) );
  NANDN U16303 ( .B(n8668), .A(\u_a23_core/u_execute/u_register_bank/r0[0] ), 
        .Z(n13785) );
  NANDN U16304 ( .B(n8671), .A(\u_a23_core/u_execute/u_register_bank/r2[0] ), 
        .Z(n13784) );
  ANDN U16305 ( .A(n8406), .B(n8413), .Z(n11969) );
  ANDN U16306 ( .A(n13786), .B(n1939), .Z(n879) );
  IV U16307 ( .A(m_address[4]), .Z(n1939) );
  AND U16308 ( .A(n5081), .B(m_address[3]), .Z(n13786) );
  ANDN U16309 ( .A(n4963), .B(m_address[2]), .Z(n5081) );
  ANDN U16310 ( .A(n1940), .B(n4518), .Z(n4963) );
  IV U16311 ( .A(n4148), .Z(n4518) );
  AND U16312 ( .A(n13787), .B(n13788), .Z(n4148) );
  AND U16313 ( .A(n13789), .B(n13790), .Z(n13788) );
  AND U16314 ( .A(n13791), .B(n13792), .Z(n13790) );
  ANDN U16315 ( .A(n13793), .B(m_address[7]), .Z(n13792) );
  NOR U16316 ( .A(m_address[9]), .B(m_address[8]), .Z(n13793) );
  NOR U16317 ( .A(m_address[23]), .B(m_address[22]), .Z(n13791) );
  AND U16318 ( .A(n13794), .B(n13795), .Z(n13789) );
  NOR U16319 ( .A(m_address[21]), .B(m_address[20]), .Z(n13795) );
  NOR U16320 ( .A(m_address[19]), .B(m_address[18]), .Z(n13794) );
  AND U16321 ( .A(n13796), .B(n13797), .Z(n13787) );
  AND U16322 ( .A(n13798), .B(n13799), .Z(n13797) );
  NOR U16323 ( .A(m_address[17]), .B(m_address[16]), .Z(n13799) );
  NOR U16324 ( .A(m_address[15]), .B(m_address[14]), .Z(n13798) );
  AND U16325 ( .A(n13800), .B(n13801), .Z(n13796) );
  NOR U16326 ( .A(m_address[13]), .B(m_address[12]), .Z(n13801) );
  NOR U16327 ( .A(m_address[11]), .B(m_address[10]), .Z(n13800) );
  AND U16328 ( .A(n2428), .B(n2429), .Z(n1940) );
  IV U16329 ( .A(m_address[6]), .Z(n2429) );
  IV U16330 ( .A(m_address[5]), .Z(n2428) );
  AND U16331 ( .A(n13802), .B(n13803), .Z(n13095) );
  AND U16332 ( .A(\u_a23_core/execute_address_nxt[4] ), .B(
        \u_a23_core/execute_address_nxt[3] ), .Z(n13803) );
  NAND U16333 ( .A(n13804), .B(n13805), .Z(\u_a23_core/execute_address_nxt[3] ) );
  AND U16334 ( .A(n13806), .B(n13807), .Z(n13805) );
  AND U16335 ( .A(n13808), .B(n13809), .Z(n13807) );
  NANDN U16336 ( .B(n8392), .A(\u_a23_core/u_execute/pc_minus4[3] ), .Z(n13809) );
  NAND U16337 ( .A(n8393), .B(\u_a23_core/u_execute/alu_out_pc_filtered[3] ), 
        .Z(n13808) );
  IV U16338 ( .A(n7016), .Z(\u_a23_core/u_execute/alu_out_pc_filtered[3] ) );
  AND U16339 ( .A(n13810), .B(n13811), .Z(n7016) );
  MUX U16340 ( .IN0(n13812), .IN1(n13813), .SEL(
        \u_a23_core/u_execute/u_alu/b_not[3] ), .F(n13811) );
  NAND U16341 ( .A(n13814), .B(n13815), .Z(
        \u_a23_core/u_execute/u_alu/b_not[3] ) );
  MUX U16342 ( .IN0(n8430), .IN1(n8431), .SEL(n13816), .F(n13815) );
  MUX U16343 ( .IN0(n8433), .IN1(n8434), .SEL(\u_a23_core/u_execute/rn[3] ), 
        .F(n13814) );
  ANDN U16344 ( .A(n8398), .B(n13817), .Z(n13813) );
  MUX U16345 ( .IN0(n8400), .IN1(\u_a23_core/alu_function[3] ), .SEL(
        \u_a23_core/u_execute/u_alu/a[3] ), .F(n13817) );
  NAND U16346 ( .A(\u_a23_core/u_execute/u_alu/a[3] ), .B(n8400), .Z(n13812)
         );
  IV U16347 ( .A(n13818), .Z(\u_a23_core/u_execute/u_alu/a[3] ) );
  MUX U16348 ( .IN0(n13819), .IN1(n13816), .SEL(\u_a23_core/alu_function[8] ), 
        .F(n13818) );
  AND U16349 ( .A(n13820), .B(n13821), .Z(n13816) );
  AND U16350 ( .A(n13822), .B(n13823), .Z(n13821) );
  NAND U16351 ( .A(n6985), .B(n6802), .Z(n13823) );
  AND U16352 ( .A(n13824), .B(n13436), .Z(n13822) );
  NAND U16353 ( .A(n13825), .B(n6902), .Z(n13824) );
  NAND U16354 ( .A(n13826), .B(n13827), .Z(n13825) );
  AND U16355 ( .A(n13828), .B(n13829), .Z(n13827) );
  NAND U16356 ( .A(n6920), .B(n6916), .Z(n13829) );
  NAND U16357 ( .A(n9082), .B(n6898), .Z(n13828) );
  AND U16358 ( .A(n11905), .B(n6878), .Z(n13826) );
  NAND U16359 ( .A(n9135), .B(n6926), .Z(n6878) );
  NAND U16360 ( .A(n6984), .B(n6925), .Z(n11905) );
  AND U16361 ( .A(n13830), .B(n13831), .Z(n13820) );
  NAND U16362 ( .A(n6786), .B(n13832), .Z(n13831) );
  NAND U16363 ( .A(n13833), .B(n13834), .Z(n13832) );
  AND U16364 ( .A(n13835), .B(n13836), .Z(n13834) );
  AND U16365 ( .A(n13837), .B(n13838), .Z(n13836) );
  AND U16366 ( .A(n13839), .B(n13840), .Z(n13838) );
  AND U16367 ( .A(n9351), .B(n13841), .Z(n13840) );
  NAND U16368 ( .A(n8464), .B(n6857), .Z(n13841) );
  NAND U16369 ( .A(n8465), .B(n6859), .Z(n9351) );
  AND U16370 ( .A(n10090), .B(n9718), .Z(n13839) );
  NAND U16371 ( .A(n6865), .B(n8461), .Z(n9718) );
  NAND U16372 ( .A(n6967), .B(n8470), .Z(n10090) );
  AND U16373 ( .A(n13842), .B(n10841), .Z(n13837) );
  NAND U16374 ( .A(n6961), .B(n9726), .Z(n10841) );
  AND U16375 ( .A(n10458), .B(n13843), .Z(n13842) );
  NAND U16376 ( .A(n6809), .B(n6822), .Z(n13843) );
  NAND U16377 ( .A(n6966), .B(n9359), .Z(n10458) );
  AND U16378 ( .A(n13844), .B(n13845), .Z(n13835) );
  AND U16379 ( .A(n13846), .B(n13847), .Z(n13845) );
  AND U16380 ( .A(n13848), .B(n13849), .Z(n13847) );
  NAND U16381 ( .A(n6807), .B(n6826), .Z(n13849) );
  NAND U16382 ( .A(n6832), .B(n6799), .Z(n13848) );
  AND U16383 ( .A(n13850), .B(n13851), .Z(n13846) );
  NAND U16384 ( .A(n6834), .B(n6803), .Z(n13851) );
  NAND U16385 ( .A(n6838), .B(n6823), .Z(n13850) );
  AND U16386 ( .A(n13852), .B(n13853), .Z(n13844) );
  NAND U16387 ( .A(n6852), .B(n6833), .Z(n13853) );
  AND U16388 ( .A(n13854), .B(n13855), .Z(n13852) );
  NAND U16389 ( .A(n6840), .B(n6835), .Z(n13855) );
  NAND U16390 ( .A(n6827), .B(n6851), .Z(n13854) );
  AND U16391 ( .A(n13856), .B(n13857), .Z(n13833) );
  AND U16392 ( .A(n13858), .B(n13859), .Z(n13857) );
  AND U16393 ( .A(n13860), .B(n13861), .Z(n13859) );
  AND U16394 ( .A(n13862), .B(n13863), .Z(n13861) );
  NAND U16395 ( .A(n6856), .B(n6839), .Z(n13863) );
  NAND U16396 ( .A(n6850), .B(n6858), .Z(n13862) );
  AND U16397 ( .A(n13864), .B(n13865), .Z(n13860) );
  NAND U16398 ( .A(n6864), .B(n6853), .Z(n13865) );
  NAND U16399 ( .A(n6841), .B(n8487), .Z(n13864) );
  AND U16400 ( .A(n13866), .B(n11783), .Z(n13858) );
  NAND U16401 ( .A(n8609), .B(n6960), .Z(n11783) );
  AND U16402 ( .A(n11222), .B(n12130), .Z(n13866) );
  NAND U16403 ( .A(n8606), .B(n6957), .Z(n12130) );
  NAND U16404 ( .A(n6956), .B(n8603), .Z(n11222) );
  AND U16405 ( .A(n13867), .B(n13868), .Z(n13856) );
  AND U16406 ( .A(n13869), .B(n13870), .Z(n13868) );
  AND U16407 ( .A(n12871), .B(n12495), .Z(n13870) );
  NAND U16408 ( .A(n8610), .B(n6947), .Z(n12495) );
  NAND U16409 ( .A(n8616), .B(n6946), .Z(n12871) );
  AND U16410 ( .A(n8614), .B(n13238), .Z(n13869) );
  NAND U16411 ( .A(n8958), .B(n6943), .Z(n13238) );
  NAND U16412 ( .A(n9082), .B(n6942), .Z(n8614) );
  AND U16413 ( .A(n13871), .B(n13872), .Z(n13867) );
  NAND U16414 ( .A(n6893), .B(n6920), .Z(n13872) );
  AND U16415 ( .A(n9080), .B(n13550), .Z(n13871) );
  NAND U16416 ( .A(n9135), .B(n6937), .Z(n13550) );
  NAND U16417 ( .A(n6984), .B(n6919), .Z(n9080) );
  NAND U16418 ( .A(n13873), .B(n6888), .Z(n13830) );
  NAND U16419 ( .A(n13874), .B(n13875), .Z(n13873) );
  AND U16420 ( .A(n13876), .B(n13877), .Z(n13875) );
  AND U16421 ( .A(n13878), .B(n13879), .Z(n13877) );
  AND U16422 ( .A(n13880), .B(n13881), .Z(n13879) );
  AND U16423 ( .A(n13882), .B(n13883), .Z(n13881) );
  NAND U16424 ( .A(n6919), .B(n6897), .Z(n13883) );
  NAND U16425 ( .A(n6920), .B(n8512), .Z(n13882) );
  AND U16426 ( .A(n13884), .B(n13885), .Z(n13880) );
  NANDN U16427 ( .B(n8516), .A(n6925), .Z(n13885) );
  NANDN U16428 ( .B(n8522), .A(n6926), .Z(n13884) );
  AND U16429 ( .A(n13886), .B(n13887), .Z(n13878) );
  AND U16430 ( .A(n13888), .B(n13889), .Z(n13887) );
  NANDN U16431 ( .B(n8526), .A(n6898), .Z(n13889) );
  NANDN U16432 ( .B(n8534), .A(n6882), .Z(n13888) );
  AND U16433 ( .A(n13890), .B(n13891), .Z(n13886) );
  NANDN U16434 ( .B(n8511), .A(n6809), .Z(n13891) );
  NANDN U16435 ( .B(n8515), .A(n6807), .Z(n13890) );
  AND U16436 ( .A(n13892), .B(n13893), .Z(n13876) );
  AND U16437 ( .A(n13894), .B(n13895), .Z(n13893) );
  AND U16438 ( .A(n13896), .B(n13897), .Z(n13895) );
  NANDN U16439 ( .B(n8521), .A(n6799), .Z(n13897) );
  NANDN U16440 ( .B(n8525), .A(n6803), .Z(n13896) );
  AND U16441 ( .A(n13898), .B(n13899), .Z(n13894) );
  NANDN U16442 ( .B(n8533), .A(n6823), .Z(n13899) );
  NANDN U16443 ( .B(n8537), .A(n6827), .Z(n13898) );
  AND U16444 ( .A(n13900), .B(n13901), .Z(n13892) );
  AND U16445 ( .A(n13902), .B(n13903), .Z(n13901) );
  NANDN U16446 ( .B(n8538), .A(n6833), .Z(n13903) );
  NANDN U16447 ( .B(n8543), .A(n6835), .Z(n13902) );
  AND U16448 ( .A(n13904), .B(n13905), .Z(n13900) );
  NANDN U16449 ( .B(n8544), .A(n6839), .Z(n13905) );
  NANDN U16450 ( .B(n8547), .A(n6850), .Z(n13904) );
  AND U16451 ( .A(n13906), .B(n13907), .Z(n13874) );
  AND U16452 ( .A(n13908), .B(n13909), .Z(n13907) );
  AND U16453 ( .A(n13910), .B(n13911), .Z(n13909) );
  AND U16454 ( .A(n13912), .B(n13913), .Z(n13911) );
  NANDN U16455 ( .B(n8548), .A(n6853), .Z(n13913) );
  NANDN U16456 ( .B(n8557), .A(n6841), .Z(n13912) );
  AND U16457 ( .A(n13914), .B(n13915), .Z(n13910) );
  NANDN U16458 ( .B(n8558), .A(n6857), .Z(n13915) );
  NANDN U16459 ( .B(n8561), .A(n6859), .Z(n13914) );
  AND U16460 ( .A(n13916), .B(n13917), .Z(n13908) );
  AND U16461 ( .A(n13918), .B(n13919), .Z(n13917) );
  NANDN U16462 ( .B(n8562), .A(n6865), .Z(n13919) );
  NANDN U16463 ( .B(n8567), .A(n6967), .Z(n13918) );
  AND U16464 ( .A(n13920), .B(n13921), .Z(n13916) );
  NANDN U16465 ( .B(n8568), .A(n6966), .Z(n13921) );
  NANDN U16466 ( .B(n8571), .A(n6961), .Z(n13920) );
  AND U16467 ( .A(n13922), .B(n13923), .Z(n13906) );
  AND U16468 ( .A(n13924), .B(n13925), .Z(n13923) );
  AND U16469 ( .A(n13926), .B(n13927), .Z(n13925) );
  NANDN U16470 ( .B(n8572), .A(n6956), .Z(n13927) );
  NANDN U16471 ( .B(n8579), .A(n6960), .Z(n13926) );
  AND U16472 ( .A(n13928), .B(n13929), .Z(n13924) );
  NANDN U16473 ( .B(n8580), .A(n6957), .Z(n13929) );
  NANDN U16474 ( .B(n8583), .A(n6947), .Z(n13928) );
  AND U16475 ( .A(n13930), .B(n13931), .Z(n13922) );
  AND U16476 ( .A(n13932), .B(n13933), .Z(n13931) );
  NANDN U16477 ( .B(n8584), .A(n6946), .Z(n13933) );
  NANDN U16478 ( .B(n8589), .A(n6943), .Z(n13932) );
  AND U16479 ( .A(n13934), .B(n13935), .Z(n13930) );
  NANDN U16480 ( .B(n8590), .A(n6942), .Z(n13935) );
  NANDN U16481 ( .B(n8593), .A(n6937), .Z(n13934) );
  IV U16482 ( .A(\u_a23_core/u_execute/rn[3] ), .Z(n13819) );
  NAND U16483 ( .A(n6765), .B(\u_a23_core/u_execute/u_alu/fadder_out[3] ), .Z(
        n13810) );
  AND U16484 ( .A(n13936), .B(n13937), .Z(n13806) );
  NANDN U16485 ( .B(n8406), .A(\u_a23_core/u_execute/rn_plus4[3] ), .Z(n13937)
         );
  NANDN U16486 ( .B(n8407), .A(\u_a23_core/u_execute/alu_plus4[3] ), .Z(n13936) );
  AND U16487 ( .A(n13938), .B(n13939), .Z(n13804) );
  AND U16488 ( .A(n13940), .B(n13941), .Z(n13939) );
  NAND U16489 ( .A(n8412), .B(\u_a23_core/u_execute/address_plus4[3] ), .Z(
        n13941) );
  NAND U16490 ( .A(\u_a23_core/u_execute/rn[3] ), .B(n8413), .Z(n13940) );
  NAND U16491 ( .A(n13942), .B(n13943), .Z(\u_a23_core/u_execute/rn[3] ) );
  AND U16492 ( .A(n13944), .B(n13945), .Z(n13943) );
  AND U16493 ( .A(n13946), .B(n13947), .Z(n13945) );
  AND U16494 ( .A(n13948), .B(n13949), .Z(n13947) );
  NANDN U16495 ( .B(n8635), .A(\u_a23_core/u_execute/pc[3] ), .Z(n13949) );
  NANDN U16496 ( .B(n8636), .A(\u_a23_core/u_execute/u_register_bank/r14[3] ), 
        .Z(n13948) );
  AND U16497 ( .A(n13950), .B(n13951), .Z(n13946) );
  NANDN U16498 ( .B(n8639), .A(\u_a23_core/u_execute/u_register_bank/r13[3] ), 
        .Z(n13951) );
  NANDN U16499 ( .B(n8640), .A(\u_a23_core/u_execute/u_register_bank/r12[3] ), 
        .Z(n13950) );
  AND U16500 ( .A(n13952), .B(n13953), .Z(n13944) );
  AND U16501 ( .A(n13954), .B(n13955), .Z(n13953) );
  NANDN U16502 ( .B(n8645), .A(\u_a23_core/u_execute/u_register_bank/r11[3] ), 
        .Z(n13955) );
  NANDN U16503 ( .B(n8646), .A(\u_a23_core/u_execute/u_register_bank/r10[3] ), 
        .Z(n13954) );
  AND U16504 ( .A(n13956), .B(n13957), .Z(n13952) );
  NANDN U16505 ( .B(n8649), .A(\u_a23_core/u_execute/u_register_bank/r9[3] ), 
        .Z(n13957) );
  NANDN U16506 ( .B(n8650), .A(\u_a23_core/u_execute/u_register_bank/r8[3] ), 
        .Z(n13956) );
  AND U16507 ( .A(n13958), .B(n13959), .Z(n13942) );
  AND U16508 ( .A(n13960), .B(n13961), .Z(n13959) );
  AND U16509 ( .A(n13962), .B(n13963), .Z(n13961) );
  NANDN U16510 ( .B(n8657), .A(\u_a23_core/u_execute/u_register_bank/r7[3] ), 
        .Z(n13963) );
  NANDN U16511 ( .B(n8658), .A(\u_a23_core/u_execute/u_register_bank/r6[3] ), 
        .Z(n13962) );
  AND U16512 ( .A(n13964), .B(n13965), .Z(n13960) );
  NANDN U16513 ( .B(n8661), .A(\u_a23_core/u_execute/u_register_bank/r5[3] ), 
        .Z(n13965) );
  NANDN U16514 ( .B(n8662), .A(\u_a23_core/u_execute/u_register_bank/r4[3] ), 
        .Z(n13964) );
  AND U16515 ( .A(n13966), .B(n13967), .Z(n13958) );
  AND U16516 ( .A(n13968), .B(n13969), .Z(n13967) );
  NANDN U16517 ( .B(n8667), .A(\u_a23_core/u_execute/u_register_bank/r3[3] ), 
        .Z(n13969) );
  NANDN U16518 ( .B(n8668), .A(\u_a23_core/u_execute/u_register_bank/r0[3] ), 
        .Z(n13968) );
  AND U16519 ( .A(n13970), .B(n13971), .Z(n13966) );
  NANDN U16520 ( .B(n8671), .A(\u_a23_core/u_execute/u_register_bank/r2[3] ), 
        .Z(n13971) );
  NANDN U16521 ( .B(n8672), .A(\u_a23_core/u_execute/u_register_bank/r1[3] ), 
        .Z(n13970) );
  AND U16522 ( .A(n13972), .B(n13973), .Z(n13938) );
  NAND U16523 ( .A(\u_a23_core/u_execute/pc[3] ), .B(n8416), .Z(n13973) );
  NAND U16524 ( .A(n8417), .B(\u_a23_core/u_execute/pc_plus4[3] ), .Z(n13972)
         );
  NAND U16525 ( .A(n13974), .B(n13975), .Z(\u_a23_core/execute_address_nxt[4] ) );
  AND U16526 ( .A(n13976), .B(n13977), .Z(n13975) );
  AND U16527 ( .A(n13978), .B(n13979), .Z(n13977) );
  NANDN U16528 ( .B(n8392), .A(\u_a23_core/u_execute/pc_minus4[4] ), .Z(n13979) );
  NAND U16529 ( .A(\u_a23_core/u_execute/alu_out_pc_filtered[4] ), .B(n8393), 
        .Z(n13978) );
  IV U16530 ( .A(n7015), .Z(\u_a23_core/u_execute/alu_out_pc_filtered[4] ) );
  AND U16531 ( .A(n13980), .B(n13981), .Z(n7015) );
  MUX U16532 ( .IN0(n13982), .IN1(n13983), .SEL(
        \u_a23_core/u_execute/u_alu/b_not[4] ), .F(n13981) );
  NAND U16533 ( .A(n13984), .B(n13985), .Z(
        \u_a23_core/u_execute/u_alu/b_not[4] ) );
  MUX U16534 ( .IN0(n8430), .IN1(n8431), .SEL(n13986), .F(n13985) );
  MUX U16535 ( .IN0(n8433), .IN1(n8434), .SEL(\u_a23_core/u_execute/rn[4] ), 
        .F(n13984) );
  ANDN U16536 ( .A(n8398), .B(n13987), .Z(n13983) );
  MUX U16537 ( .IN0(n8400), .IN1(\u_a23_core/alu_function[3] ), .SEL(
        \u_a23_core/u_execute/u_alu/a[4] ), .F(n13987) );
  NAND U16538 ( .A(\u_a23_core/u_execute/u_alu/a[4] ), .B(n8400), .Z(n13982)
         );
  IV U16539 ( .A(n13988), .Z(\u_a23_core/u_execute/u_alu/a[4] ) );
  MUX U16540 ( .IN0(n13989), .IN1(n13986), .SEL(\u_a23_core/alu_function[8] ), 
        .F(n13988) );
  AND U16541 ( .A(n13990), .B(n13991), .Z(n13986) );
  AND U16542 ( .A(n13992), .B(n13436), .Z(n13991) );
  IV U16543 ( .A(n9201), .Z(n13436) );
  ANDN U16544 ( .A(n8443), .B(n13124), .Z(n9201) );
  NAND U16545 ( .A(n6882), .B(n13993), .Z(n13124) );
  NAND U16546 ( .A(n13307), .B(n13306), .Z(n13993) );
  NAND U16547 ( .A(n13994), .B(n6902), .Z(n13992) );
  NAND U16548 ( .A(n13995), .B(n13996), .Z(n13994) );
  AND U16549 ( .A(n13997), .B(n13998), .Z(n13996) );
  NAND U16550 ( .A(n9082), .B(n6926), .Z(n13998) );
  AND U16551 ( .A(n13999), .B(n14000), .Z(n13997) );
  NAND U16552 ( .A(n6919), .B(n6916), .Z(n14000) );
  NAND U16553 ( .A(n8958), .B(n6898), .Z(n13999) );
  AND U16554 ( .A(n14001), .B(n13692), .Z(n13995) );
  NAND U16555 ( .A(n9135), .B(n6925), .Z(n13692) );
  AND U16556 ( .A(n14002), .B(n14003), .Z(n13990) );
  NAND U16557 ( .A(n6786), .B(n14004), .Z(n14003) );
  NAND U16558 ( .A(n14005), .B(n14006), .Z(n14004) );
  AND U16559 ( .A(n14007), .B(n14008), .Z(n14006) );
  AND U16560 ( .A(n14009), .B(n14010), .Z(n14008) );
  AND U16561 ( .A(n14011), .B(n14012), .Z(n14010) );
  AND U16562 ( .A(n6927), .B(n14013), .Z(n14012) );
  NAND U16563 ( .A(n8464), .B(n6841), .Z(n14013) );
  NAND U16564 ( .A(n8465), .B(n6857), .Z(n6927) );
  AND U16565 ( .A(n9906), .B(n9465), .Z(n14011) );
  NAND U16566 ( .A(n8461), .B(n6859), .Z(n9465) );
  NAND U16567 ( .A(n6865), .B(n8470), .Z(n9906) );
  AND U16568 ( .A(n14014), .B(n10650), .Z(n14009) );
  NAND U16569 ( .A(n6966), .B(n9726), .Z(n10650) );
  AND U16570 ( .A(n10273), .B(n14015), .Z(n14014) );
  NAND U16571 ( .A(n6882), .B(n6822), .Z(n14015) );
  NAND U16572 ( .A(n6967), .B(n9359), .Z(n10273) );
  AND U16573 ( .A(n14016), .B(n14017), .Z(n14007) );
  AND U16574 ( .A(n14018), .B(n14019), .Z(n14017) );
  AND U16575 ( .A(n14020), .B(n14021), .Z(n14019) );
  NAND U16576 ( .A(n6809), .B(n6826), .Z(n14021) );
  NAND U16577 ( .A(n6832), .B(n6807), .Z(n14020) );
  AND U16578 ( .A(n14022), .B(n14023), .Z(n14018) );
  NAND U16579 ( .A(n6834), .B(n6799), .Z(n14023) );
  NAND U16580 ( .A(n6838), .B(n6803), .Z(n14022) );
  AND U16581 ( .A(n14024), .B(n14025), .Z(n14016) );
  NAND U16582 ( .A(n6852), .B(n6827), .Z(n14025) );
  AND U16583 ( .A(n14026), .B(n14027), .Z(n14024) );
  NAND U16584 ( .A(n6840), .B(n6833), .Z(n14027) );
  NAND U16585 ( .A(n6823), .B(n6851), .Z(n14026) );
  AND U16586 ( .A(n14028), .B(n14029), .Z(n14005) );
  AND U16587 ( .A(n14030), .B(n14031), .Z(n14029) );
  AND U16588 ( .A(n14032), .B(n14033), .Z(n14031) );
  AND U16589 ( .A(n14034), .B(n14035), .Z(n14033) );
  NAND U16590 ( .A(n6856), .B(n6835), .Z(n14035) );
  NAND U16591 ( .A(n6858), .B(n6839), .Z(n14034) );
  AND U16592 ( .A(n14036), .B(n14037), .Z(n14032) );
  NAND U16593 ( .A(n6850), .B(n6864), .Z(n14037) );
  NAND U16594 ( .A(n6853), .B(n8487), .Z(n14036) );
  AND U16595 ( .A(n14038), .B(n11408), .Z(n14030) );
  NAND U16596 ( .A(n6956), .B(n8609), .Z(n11408) );
  AND U16597 ( .A(n11040), .B(n11597), .Z(n14038) );
  NAND U16598 ( .A(n8606), .B(n6960), .Z(n11597) );
  NAND U16599 ( .A(n6961), .B(n8603), .Z(n11040) );
  AND U16600 ( .A(n14039), .B(n14040), .Z(n14028) );
  AND U16601 ( .A(n14041), .B(n14042), .Z(n14040) );
  AND U16602 ( .A(n12684), .B(n12311), .Z(n14042) );
  NAND U16603 ( .A(n8610), .B(n6957), .Z(n12311) );
  NAND U16604 ( .A(n8616), .B(n6947), .Z(n12684) );
  AND U16605 ( .A(n13424), .B(n13051), .Z(n14041) );
  NAND U16606 ( .A(n8958), .B(n6946), .Z(n13051) );
  NAND U16607 ( .A(n9082), .B(n6943), .Z(n13424) );
  AND U16608 ( .A(n14043), .B(n14044), .Z(n14039) );
  NAND U16609 ( .A(n6893), .B(n6919), .Z(n14044) );
  AND U16610 ( .A(n8960), .B(n8824), .Z(n14043) );
  NAND U16611 ( .A(n9135), .B(n6942), .Z(n8824) );
  NAND U16612 ( .A(n6984), .B(n6937), .Z(n8960) );
  NAND U16613 ( .A(n14045), .B(n6888), .Z(n14002) );
  NAND U16614 ( .A(n14046), .B(n14047), .Z(n14045) );
  AND U16615 ( .A(n14048), .B(n14049), .Z(n14047) );
  AND U16616 ( .A(n14050), .B(n14051), .Z(n14049) );
  AND U16617 ( .A(n14052), .B(n14053), .Z(n14051) );
  AND U16618 ( .A(n14054), .B(n14055), .Z(n14053) );
  NAND U16619 ( .A(n6919), .B(n8512), .Z(n14055) );
  NANDN U16620 ( .B(n8516), .A(n6920), .Z(n14054) );
  AND U16621 ( .A(n14056), .B(n14057), .Z(n14052) );
  NANDN U16622 ( .B(n8522), .A(n6925), .Z(n14057) );
  NANDN U16623 ( .B(n8526), .A(n6926), .Z(n14056) );
  AND U16624 ( .A(n14058), .B(n14059), .Z(n14050) );
  AND U16625 ( .A(n14060), .B(n14061), .Z(n14059) );
  NANDN U16626 ( .B(n8534), .A(n6898), .Z(n14061) );
  NANDN U16627 ( .B(n8511), .A(n6882), .Z(n14060) );
  AND U16628 ( .A(n14062), .B(n14063), .Z(n14058) );
  NANDN U16629 ( .B(n8515), .A(n6809), .Z(n14063) );
  NANDN U16630 ( .B(n8521), .A(n6807), .Z(n14062) );
  AND U16631 ( .A(n14064), .B(n14065), .Z(n14048) );
  AND U16632 ( .A(n14066), .B(n14067), .Z(n14065) );
  AND U16633 ( .A(n14068), .B(n14069), .Z(n14067) );
  NANDN U16634 ( .B(n8525), .A(n6799), .Z(n14069) );
  NANDN U16635 ( .B(n8533), .A(n6803), .Z(n14068) );
  AND U16636 ( .A(n14070), .B(n14071), .Z(n14066) );
  NANDN U16637 ( .B(n8537), .A(n6823), .Z(n14071) );
  NANDN U16638 ( .B(n8538), .A(n6827), .Z(n14070) );
  AND U16639 ( .A(n14072), .B(n14073), .Z(n14064) );
  AND U16640 ( .A(n14074), .B(n14075), .Z(n14073) );
  NANDN U16641 ( .B(n8543), .A(n6833), .Z(n14075) );
  NANDN U16642 ( .B(n8544), .A(n6835), .Z(n14074) );
  AND U16643 ( .A(n14076), .B(n14077), .Z(n14072) );
  NANDN U16644 ( .B(n8547), .A(n6839), .Z(n14077) );
  NANDN U16645 ( .B(n8548), .A(n6850), .Z(n14076) );
  AND U16646 ( .A(n14078), .B(n14079), .Z(n14046) );
  AND U16647 ( .A(n14080), .B(n14081), .Z(n14079) );
  AND U16648 ( .A(n14082), .B(n14083), .Z(n14081) );
  AND U16649 ( .A(n14084), .B(n14085), .Z(n14083) );
  NANDN U16650 ( .B(n8557), .A(n6853), .Z(n14085) );
  NANDN U16651 ( .B(n8558), .A(n6841), .Z(n14084) );
  AND U16652 ( .A(n14086), .B(n14087), .Z(n14082) );
  NANDN U16653 ( .B(n8561), .A(n6857), .Z(n14087) );
  NANDN U16654 ( .B(n8562), .A(n6859), .Z(n14086) );
  AND U16655 ( .A(n14088), .B(n14089), .Z(n14080) );
  AND U16656 ( .A(n14090), .B(n14091), .Z(n14089) );
  NANDN U16657 ( .B(n8567), .A(n6865), .Z(n14091) );
  NANDN U16658 ( .B(n8568), .A(n6967), .Z(n14090) );
  AND U16659 ( .A(n14092), .B(n14093), .Z(n14088) );
  NANDN U16660 ( .B(n8571), .A(n6966), .Z(n14093) );
  NANDN U16661 ( .B(n8572), .A(n6961), .Z(n14092) );
  AND U16662 ( .A(n14094), .B(n14095), .Z(n14078) );
  AND U16663 ( .A(n14096), .B(n14097), .Z(n14095) );
  AND U16664 ( .A(n14098), .B(n14099), .Z(n14097) );
  NANDN U16665 ( .B(n8579), .A(n6956), .Z(n14099) );
  NANDN U16666 ( .B(n8580), .A(n6960), .Z(n14098) );
  AND U16667 ( .A(n14100), .B(n14101), .Z(n14096) );
  NANDN U16668 ( .B(n8583), .A(n6957), .Z(n14101) );
  NANDN U16669 ( .B(n8584), .A(n6947), .Z(n14100) );
  AND U16670 ( .A(n14102), .B(n14103), .Z(n14094) );
  AND U16671 ( .A(n14104), .B(n14105), .Z(n14103) );
  NANDN U16672 ( .B(n8589), .A(n6946), .Z(n14105) );
  NANDN U16673 ( .B(n8590), .A(n6943), .Z(n14104) );
  AND U16674 ( .A(n14106), .B(n14107), .Z(n14102) );
  NANDN U16675 ( .B(n8593), .A(n6942), .Z(n14107) );
  NAND U16676 ( .A(n6937), .B(n6897), .Z(n14106) );
  IV U16677 ( .A(\u_a23_core/u_execute/rn[4] ), .Z(n13989) );
  NAND U16678 ( .A(n6765), .B(\u_a23_core/u_execute/u_alu/fadder_out[4] ), .Z(
        n13980) );
  AND U16679 ( .A(n14108), .B(n14109), .Z(n13976) );
  NANDN U16680 ( .B(n8406), .A(\u_a23_core/u_execute/rn_plus4[4] ), .Z(n14109)
         );
  NANDN U16681 ( .B(n8407), .A(\u_a23_core/u_execute/alu_plus4[4] ), .Z(n14108) );
  AND U16682 ( .A(n14110), .B(n14111), .Z(n13974) );
  AND U16683 ( .A(n14112), .B(n14113), .Z(n14111) );
  NAND U16684 ( .A(n8412), .B(\u_a23_core/u_execute/address_plus4[4] ), .Z(
        n14113) );
  NAND U16685 ( .A(\u_a23_core/u_execute/rn[4] ), .B(n8413), .Z(n14112) );
  NAND U16686 ( .A(n14114), .B(n14115), .Z(\u_a23_core/u_execute/rn[4] ) );
  AND U16687 ( .A(n14116), .B(n14117), .Z(n14115) );
  AND U16688 ( .A(n14118), .B(n14119), .Z(n14117) );
  AND U16689 ( .A(n14120), .B(n14121), .Z(n14119) );
  NANDN U16690 ( .B(n8635), .A(\u_a23_core/u_execute/pc[4] ), .Z(n14121) );
  NANDN U16691 ( .B(n8636), .A(\u_a23_core/u_execute/u_register_bank/r14[4] ), 
        .Z(n14120) );
  AND U16692 ( .A(n14122), .B(n14123), .Z(n14118) );
  NANDN U16693 ( .B(n8639), .A(\u_a23_core/u_execute/u_register_bank/r13[4] ), 
        .Z(n14123) );
  NANDN U16694 ( .B(n8640), .A(\u_a23_core/u_execute/u_register_bank/r12[4] ), 
        .Z(n14122) );
  AND U16695 ( .A(n14124), .B(n14125), .Z(n14116) );
  AND U16696 ( .A(n14126), .B(n14127), .Z(n14125) );
  NANDN U16697 ( .B(n8645), .A(\u_a23_core/u_execute/u_register_bank/r11[4] ), 
        .Z(n14127) );
  NANDN U16698 ( .B(n8646), .A(\u_a23_core/u_execute/u_register_bank/r10[4] ), 
        .Z(n14126) );
  AND U16699 ( .A(n14128), .B(n14129), .Z(n14124) );
  NANDN U16700 ( .B(n8649), .A(\u_a23_core/u_execute/u_register_bank/r9[4] ), 
        .Z(n14129) );
  NANDN U16701 ( .B(n8650), .A(\u_a23_core/u_execute/u_register_bank/r8[4] ), 
        .Z(n14128) );
  AND U16702 ( .A(n14130), .B(n14131), .Z(n14114) );
  AND U16703 ( .A(n14132), .B(n14133), .Z(n14131) );
  AND U16704 ( .A(n14134), .B(n14135), .Z(n14133) );
  NANDN U16705 ( .B(n8657), .A(\u_a23_core/u_execute/u_register_bank/r7[4] ), 
        .Z(n14135) );
  NANDN U16706 ( .B(n8658), .A(\u_a23_core/u_execute/u_register_bank/r6[4] ), 
        .Z(n14134) );
  AND U16707 ( .A(n14136), .B(n14137), .Z(n14132) );
  NANDN U16708 ( .B(n8661), .A(\u_a23_core/u_execute/u_register_bank/r5[4] ), 
        .Z(n14137) );
  NANDN U16709 ( .B(n8662), .A(\u_a23_core/u_execute/u_register_bank/r4[4] ), 
        .Z(n14136) );
  AND U16710 ( .A(n14138), .B(n14139), .Z(n14130) );
  AND U16711 ( .A(n14140), .B(n14141), .Z(n14139) );
  NANDN U16712 ( .B(n8667), .A(\u_a23_core/u_execute/u_register_bank/r3[4] ), 
        .Z(n14141) );
  NANDN U16713 ( .B(n8668), .A(\u_a23_core/u_execute/u_register_bank/r0[4] ), 
        .Z(n14140) );
  AND U16714 ( .A(n14142), .B(n14143), .Z(n14138) );
  NANDN U16715 ( .B(n8671), .A(\u_a23_core/u_execute/u_register_bank/r2[4] ), 
        .Z(n14143) );
  NANDN U16716 ( .B(n8672), .A(\u_a23_core/u_execute/u_register_bank/r1[4] ), 
        .Z(n14142) );
  AND U16717 ( .A(n14144), .B(n14145), .Z(n14110) );
  NAND U16718 ( .A(\u_a23_core/u_execute/pc[4] ), .B(n8416), .Z(n14145) );
  NAND U16719 ( .A(n8417), .B(\u_a23_core/u_execute/pc_plus4[4] ), .Z(n14144)
         );
  IV U16720 ( .A(n14146), .Z(n8417) );
  ANDN U16721 ( .A(\u_a23_core/execute_address_nxt[2] ), .B(n4962), .Z(n13802)
         );
  NAND U16722 ( .A(n8192), .B(n8203), .Z(n4962) );
  ANDN U16723 ( .A(n14147), .B(n14148), .Z(n8203) );
  IV U16724 ( .A(n8193), .Z(n14148) );
  AND U16725 ( .A(n14149), .B(n14150), .Z(n8193) );
  ANDN U16726 ( .A(n14151), .B(m_address[29]), .Z(n14150) );
  NOR U16727 ( .A(m_address[31]), .B(m_address[30]), .Z(n14151) );
  NOR U16728 ( .A(m_address[28]), .B(m_address[27]), .Z(n14149) );
  AND U16729 ( .A(n8198), .B(n8191), .Z(n14147) );
  IV U16730 ( .A(m_address[25]), .Z(n8191) );
  IV U16731 ( .A(m_address[24]), .Z(n8198) );
  IV U16732 ( .A(m_address[26]), .Z(n8192) );
  NAND U16733 ( .A(n14152), .B(n14153), .Z(\u_a23_core/execute_address_nxt[2] ) );
  ANDN U16734 ( .A(n14154), .B(n14155), .Z(n14153) );
  MUX U16735 ( .IN0(n14156), .IN1(n8416), .SEL(\u_a23_core/u_execute/pc[2] ), 
        .F(n14155) );
  NOR U16736 ( .A(\u_a23_core/address_sel[2] ), .B(n14157), .Z(n8416) );
  NAND U16737 ( .A(n14146), .B(n8392), .Z(n14156) );
  NANDN U16738 ( .B(n14158), .A(n6099), .Z(n8392) );
  NAND U16739 ( .A(n14159), .B(n14160), .Z(n14146) );
  NAND U16740 ( .A(n4146), .B(n8412), .Z(n14154) );
  ANDN U16741 ( .A(n14161), .B(n14162), .Z(n8412) );
  AND U16742 ( .A(n14160), .B(\u_a23_core/address_sel[0] ), .Z(n14161) );
  IV U16743 ( .A(m_address[2]), .Z(n4146) );
  AND U16744 ( .A(n14163), .B(n14164), .Z(n14152) );
  MUX U16745 ( .IN0(n8407), .IN1(n14165), .SEL(
        \u_a23_core/u_execute/alu_out_pc_filtered[2] ), .F(n14164) );
  IV U16746 ( .A(n7017), .Z(\u_a23_core/u_execute/alu_out_pc_filtered[2] ) );
  AND U16747 ( .A(n14166), .B(n14167), .Z(n7017) );
  MUX U16748 ( .IN0(n14168), .IN1(n14169), .SEL(
        \u_a23_core/u_execute/u_alu/b_not[2] ), .F(n14167) );
  NAND U16749 ( .A(n14170), .B(n14171), .Z(
        \u_a23_core/u_execute/u_alu/b_not[2] ) );
  MUX U16750 ( .IN0(n8430), .IN1(n8431), .SEL(n14172), .F(n14171) );
  IV U16751 ( .A(n13630), .Z(n8431) );
  ANDN U16752 ( .A(n14173), .B(n14174), .Z(n13630) );
  IV U16753 ( .A(n13629), .Z(n8430) );
  ANDN U16754 ( .A(n14173), .B(\u_a23_core/alu_function[7] ), .Z(n13629) );
  MUX U16755 ( .IN0(n8433), .IN1(n8434), .SEL(\u_a23_core/u_execute/rn[2] ), 
        .F(n14170) );
  IV U16756 ( .A(n13632), .Z(n8434) );
  NOR U16757 ( .A(n14173), .B(\u_a23_core/alu_function[7] ), .Z(n13632) );
  IV U16758 ( .A(\u_a23_core/alu_function[8] ), .Z(n14173) );
  IV U16759 ( .A(n13633), .Z(n8433) );
  ANDN U16760 ( .A(\u_a23_core/alu_function[8] ), .B(n14174), .Z(n13633) );
  IV U16761 ( .A(\u_a23_core/alu_function[7] ), .Z(n14174) );
  ANDN U16762 ( .A(n8398), .B(n14175), .Z(n14169) );
  MUX U16763 ( .IN0(n8400), .IN1(\u_a23_core/alu_function[3] ), .SEL(
        \u_a23_core/u_execute/u_alu/a[2] ), .F(n14175) );
  AND U16764 ( .A(n14176), .B(n14177), .Z(n8398) );
  AND U16765 ( .A(n13428), .B(n13297), .Z(n14177) );
  IV U16766 ( .A(n12320), .Z(n13297) );
  NOR U16767 ( .A(\u_a23_core/alu_function[0] ), .B(n14178), .Z(n12320) );
  NANDN U16768 ( .B(n14178), .A(\u_a23_core/alu_function[0] ), .Z(n13428) );
  NAND U16769 ( .A(\u_a23_core/alu_function[2] ), .B(n14179), .Z(n14178) );
  ANDN U16770 ( .A(n14180), .B(\u_a23_core/alu_function[3] ), .Z(n14179) );
  AND U16771 ( .A(n9256), .B(n14181), .Z(n14176) );
  NAND U16772 ( .A(\u_a23_core/alu_function[1] ), .B(n14182), .Z(n14181) );
  AND U16773 ( .A(n14183), .B(n13296), .Z(n9256) );
  NAND U16774 ( .A(n8400), .B(\u_a23_core/alu_function[0] ), .Z(n13296) );
  NANDN U16775 ( .B(n13295), .A(n14180), .Z(n14183) );
  NANDN U16776 ( .B(\u_a23_core/alu_function[0] ), .A(n14182), .Z(n13295) );
  NAND U16777 ( .A(\u_a23_core/u_execute/u_alu/a[2] ), .B(n8400), .Z(n14168)
         );
  AND U16778 ( .A(n14184), .B(\u_a23_core/alu_function[1] ), .Z(n8400) );
  ANDN U16779 ( .A(\u_a23_core/alu_function[2] ), .B(
        \u_a23_core/alu_function[3] ), .Z(n14184) );
  IV U16780 ( .A(n14185), .Z(\u_a23_core/u_execute/u_alu/a[2] ) );
  MUX U16781 ( .IN0(n14186), .IN1(n14172), .SEL(\u_a23_core/alu_function[8] ), 
        .F(n14185) );
  AND U16782 ( .A(n14187), .B(n14188), .Z(n14172) );
  AND U16783 ( .A(n14189), .B(n14190), .Z(n14188) );
  NAND U16784 ( .A(n6985), .B(n6798), .Z(n14190) );
  ANDN U16785 ( .A(n8452), .B(n11110), .Z(n6985) );
  AND U16786 ( .A(n14191), .B(n14192), .Z(n14189) );
  NAND U16787 ( .A(n14193), .B(n6902), .Z(n14192) );
  NOR U16788 ( .A(\u_a23_core/barrel_shift_function[1] ), .B(
        \u_a23_core/barrel_shift_function[0] ), .Z(n6902) );
  NAND U16789 ( .A(n14194), .B(n13691), .Z(n14193) );
  NAND U16790 ( .A(n6984), .B(n6926), .Z(n13691) );
  AND U16791 ( .A(n14195), .B(n14196), .Z(n14194) );
  NAND U16792 ( .A(n6925), .B(n6916), .Z(n14196) );
  OR U16793 ( .A(n6893), .B(\u_a23_core/shift_imm_zero ), .Z(n6916) );
  NAND U16794 ( .A(n9135), .B(n6898), .Z(n14195) );
  OR U16795 ( .A(n13306), .B(n9262), .Z(n14191) );
  IV U16796 ( .A(n6886), .Z(n9262) );
  ANDN U16797 ( .A(n8443), .B(n11110), .Z(n6886) );
  IV U16798 ( .A(n6882), .Z(n11110) );
  AND U16799 ( .A(n14197), .B(n14198), .Z(n13306) );
  NOR U16800 ( .A(\u_a23_core/shift_imm_zero ), .B(n6806), .Z(n14198) );
  ANDN U16801 ( .A(n14199), .B(n6991), .Z(n6806) );
  ANDN U16802 ( .A(n13643), .B(n6798), .Z(n14197) );
  AND U16803 ( .A(n14200), .B(n14201), .Z(n6798) );
  NOR U16804 ( .A(n6885), .B(n6808), .Z(n13643) );
  ANDN U16805 ( .A(n14201), .B(n6991), .Z(n6808) );
  NAND U16806 ( .A(n14202), .B(n14203), .Z(n6991) );
  NAND U16807 ( .A(n14204), .B(n14205), .Z(n14202) );
  AND U16808 ( .A(n14206), .B(n14207), .Z(n14187) );
  NAND U16809 ( .A(n6786), .B(n14208), .Z(n14207) );
  NAND U16810 ( .A(n14209), .B(n14210), .Z(n14208) );
  AND U16811 ( .A(n14211), .B(n14212), .Z(n14210) );
  AND U16812 ( .A(n14213), .B(n14214), .Z(n14212) );
  AND U16813 ( .A(n14215), .B(n14216), .Z(n14214) );
  AND U16814 ( .A(n6928), .B(n14217), .Z(n14216) );
  NAND U16815 ( .A(n6802), .B(n6809), .Z(n14217) );
  IV U16816 ( .A(n13307), .Z(n6802) );
  NAND U16817 ( .A(n14200), .B(n14199), .Z(n13307) );
  AND U16818 ( .A(n14204), .B(n14218), .Z(n14199) );
  AND U16819 ( .A(n14203), .B(n14205), .Z(n14200) );
  ANDN U16820 ( .A(n14219), .B(n14220), .Z(n14203) );
  AND U16821 ( .A(n14221), .B(n14222), .Z(n14219) );
  NAND U16822 ( .A(n8464), .B(n6859), .Z(n6928) );
  ANDN U16823 ( .A(n14223), .B(n14224), .Z(n8464) );
  ANDN U16824 ( .A(n14225), .B(n14226), .Z(n14223) );
  AND U16825 ( .A(n9907), .B(n9466), .Z(n14215) );
  NAND U16826 ( .A(n6865), .B(n8465), .Z(n9466) );
  AND U16827 ( .A(n14227), .B(n14228), .Z(n8465) );
  ANDN U16828 ( .A(n14218), .B(n14226), .Z(n14227) );
  NAND U16829 ( .A(n6967), .B(n8461), .Z(n9907) );
  IV U16830 ( .A(n11311), .Z(n8461) );
  NANDN U16831 ( .B(n14229), .A(n14230), .Z(n11311) );
  AND U16832 ( .A(n14231), .B(n14232), .Z(n14213) );
  AND U16833 ( .A(n14233), .B(n10274), .Z(n14232) );
  NAND U16834 ( .A(n6966), .B(n8470), .Z(n10274) );
  AND U16835 ( .A(n14234), .B(n14230), .Z(n8470) );
  AND U16836 ( .A(n14235), .B(n14218), .Z(n14234) );
  NAND U16837 ( .A(n6807), .B(n6822), .Z(n14233) );
  ANDN U16838 ( .A(n14236), .B(n14222), .Z(n6822) );
  NAND U16839 ( .A(n14237), .B(n14201), .Z(n14222) );
  AND U16840 ( .A(n14204), .B(n14225), .Z(n14201) );
  AND U16841 ( .A(n11023), .B(n10651), .Z(n14231) );
  NAND U16842 ( .A(n6961), .B(n9359), .Z(n10651) );
  AND U16843 ( .A(n14238), .B(n14235), .Z(n9359) );
  ANDN U16844 ( .A(n14237), .B(n14226), .Z(n14238) );
  NAND U16845 ( .A(n6956), .B(n9726), .Z(n11023) );
  AND U16846 ( .A(n14239), .B(n14240), .Z(n9726) );
  ANDN U16847 ( .A(n14241), .B(n14226), .Z(n14239) );
  AND U16848 ( .A(n14242), .B(n14243), .Z(n14211) );
  AND U16849 ( .A(n14244), .B(n14245), .Z(n14243) );
  AND U16850 ( .A(n14246), .B(n14247), .Z(n14245) );
  NAND U16851 ( .A(n6799), .B(n6826), .Z(n14247) );
  NOR U16852 ( .A(n14220), .B(n14221), .Z(n6826) );
  NANDN U16853 ( .B(n6885), .A(n14240), .Z(n14221) );
  IV U16854 ( .A(n14236), .Z(n14220) );
  ANDN U16855 ( .A(n14248), .B(n14249), .Z(n14236) );
  NAND U16856 ( .A(n14204), .B(n6988), .Z(n14248) );
  NAND U16857 ( .A(n6832), .B(n6803), .Z(n14246) );
  ANDN U16858 ( .A(n14250), .B(n14249), .Z(n6832) );
  NAND U16859 ( .A(n14251), .B(n14252), .Z(n14249) );
  AND U16860 ( .A(n14253), .B(n14254), .Z(n14251) );
  NAND U16861 ( .A(n14204), .B(n14255), .Z(n14253) );
  AND U16862 ( .A(n14204), .B(n6988), .Z(n14250) );
  AND U16863 ( .A(n14256), .B(n14257), .Z(n14244) );
  NAND U16864 ( .A(n6834), .B(n6823), .Z(n14257) );
  AND U16865 ( .A(n14258), .B(n14252), .Z(n6834) );
  AND U16866 ( .A(n14204), .B(n14255), .Z(n14258) );
  NAND U16867 ( .A(n6838), .B(n6827), .Z(n14256) );
  ANDN U16868 ( .A(n14252), .B(n14254), .Z(n6838) );
  ANDN U16869 ( .A(n14259), .B(n14260), .Z(n14252) );
  AND U16870 ( .A(n14261), .B(n14262), .Z(n14242) );
  NAND U16871 ( .A(n6852), .B(n6835), .Z(n14262) );
  IV U16872 ( .A(n12590), .Z(n6852) );
  NAND U16873 ( .A(n14263), .B(n14264), .Z(n12590) );
  AND U16874 ( .A(n14225), .B(n14265), .Z(n14264) );
  AND U16875 ( .A(n14205), .B(n14266), .Z(n14263) );
  AND U16876 ( .A(n14267), .B(n14268), .Z(n14261) );
  NAND U16877 ( .A(n6840), .B(n6839), .Z(n14268) );
  ANDN U16878 ( .A(n14269), .B(n14270), .Z(n6840) );
  AND U16879 ( .A(n14260), .B(n14205), .Z(n14269) );
  NAND U16880 ( .A(n6833), .B(n6851), .Z(n14267) );
  AND U16881 ( .A(n14259), .B(n14260), .Z(n6851) );
  ANDN U16882 ( .A(n14271), .B(n14270), .Z(n14259) );
  IV U16883 ( .A(n14266), .Z(n14270) );
  NOR U16884 ( .A(n14272), .B(n14273), .Z(n14266) );
  NAND U16885 ( .A(n14265), .B(n14205), .Z(n14271) );
  AND U16886 ( .A(n14274), .B(n14275), .Z(n14209) );
  AND U16887 ( .A(n14276), .B(n14277), .Z(n14275) );
  AND U16888 ( .A(n14278), .B(n14279), .Z(n14277) );
  AND U16889 ( .A(n14280), .B(n14281), .Z(n14279) );
  NAND U16890 ( .A(n6850), .B(n6856), .Z(n14281) );
  IV U16891 ( .A(n12595), .Z(n6856) );
  NANDN U16892 ( .B(n14273), .A(n14272), .Z(n12595) );
  NAND U16893 ( .A(n14282), .B(n14283), .Z(n14273) );
  NANDN U16894 ( .B(n14284), .A(n14265), .Z(n14282) );
  NAND U16895 ( .A(n6858), .B(n6853), .Z(n14280) );
  AND U16896 ( .A(n14285), .B(n14272), .Z(n6858) );
  ANDN U16897 ( .A(n14237), .B(n14254), .Z(n14272) );
  IV U16898 ( .A(n14265), .Z(n14254) );
  AND U16899 ( .A(n14283), .B(n14218), .Z(n14285) );
  AND U16900 ( .A(n14286), .B(n14287), .Z(n14278) );
  NAND U16901 ( .A(n6864), .B(n6841), .Z(n14287) );
  AND U16902 ( .A(n14288), .B(n14283), .Z(n6864) );
  ANDN U16903 ( .A(n14289), .B(n14224), .Z(n14283) );
  ANDN U16904 ( .A(n14226), .B(n14290), .Z(n14289) );
  AND U16905 ( .A(n14265), .B(n6988), .Z(n14288) );
  NAND U16906 ( .A(n6857), .B(n8487), .Z(n14286) );
  ANDN U16907 ( .A(n14290), .B(n14224), .Z(n8487) );
  IV U16908 ( .A(n14228), .Z(n14224) );
  NOR U16909 ( .A(n14230), .B(n14229), .Z(n14228) );
  NAND U16910 ( .A(n14291), .B(n14235), .Z(n14229) );
  ANDN U16911 ( .A(n14292), .B(n14293), .Z(n14235) );
  OR U16912 ( .A(n14284), .B(n14226), .Z(n14292) );
  OR U16913 ( .A(n14294), .B(n14226), .Z(n14291) );
  ANDN U16914 ( .A(n14205), .B(n14226), .Z(n14230) );
  AND U16915 ( .A(n14260), .B(n6988), .Z(n14290) );
  AND U16916 ( .A(n14218), .B(n14265), .Z(n14260) );
  NOR U16917 ( .A(n6885), .B(n14295), .Z(n14265) );
  IV U16918 ( .A(n14204), .Z(n6885) );
  AND U16919 ( .A(n14296), .B(n11599), .Z(n14276) );
  NAND U16920 ( .A(n8609), .B(n6957), .Z(n11599) );
  ANDN U16921 ( .A(n14297), .B(n14298), .Z(n8609) );
  ANDN U16922 ( .A(n14255), .B(n14226), .Z(n14297) );
  AND U16923 ( .A(n11409), .B(n12303), .Z(n14296) );
  NAND U16924 ( .A(n8606), .B(n6947), .Z(n12303) );
  ANDN U16925 ( .A(n14299), .B(n14298), .Z(n8606) );
  NAND U16926 ( .A(n8603), .B(n6960), .Z(n11409) );
  ANDN U16927 ( .A(n14300), .B(n14293), .Z(n8603) );
  IV U16928 ( .A(n14241), .Z(n14293) );
  ANDN U16929 ( .A(n14301), .B(n14298), .Z(n14241) );
  NAND U16930 ( .A(n14302), .B(n14303), .Z(n14298) );
  NAND U16931 ( .A(n14299), .B(n14304), .Z(n14302) );
  NAND U16932 ( .A(n14305), .B(n14225), .Z(n14304) );
  ANDN U16933 ( .A(n14306), .B(n14299), .Z(n14301) );
  NANDN U16934 ( .B(n14226), .A(n14255), .Z(n14306) );
  ANDN U16935 ( .A(n6988), .B(n14226), .Z(n14300) );
  AND U16936 ( .A(n14307), .B(n14308), .Z(n14274) );
  AND U16937 ( .A(n14309), .B(n14310), .Z(n14308) );
  AND U16938 ( .A(n13052), .B(n12682), .Z(n14310) );
  NAND U16939 ( .A(n8610), .B(n6946), .Z(n12682) );
  AND U16940 ( .A(n14311), .B(n14303), .Z(n8610) );
  AND U16941 ( .A(n14299), .B(n14218), .Z(n14311) );
  NAND U16942 ( .A(n8616), .B(n6943), .Z(n13052) );
  AND U16943 ( .A(n14312), .B(n14303), .Z(n8616) );
  ANDN U16944 ( .A(n14313), .B(n14314), .Z(n14303) );
  NOR U16945 ( .A(n14315), .B(n14316), .Z(n14313) );
  AND U16946 ( .A(n14299), .B(n14205), .Z(n14312) );
  AND U16947 ( .A(n8821), .B(n13425), .Z(n14309) );
  NAND U16948 ( .A(n8958), .B(n6942), .Z(n13425) );
  ANDN U16949 ( .A(n14316), .B(n14314), .Z(n8958) );
  AND U16950 ( .A(n14317), .B(n14299), .Z(n14316) );
  NAND U16951 ( .A(n9082), .B(n6937), .Z(n8821) );
  ANDN U16952 ( .A(n14315), .B(n14314), .Z(n9082) );
  NANDN U16953 ( .B(n14318), .A(n14319), .Z(n14314) );
  ANDN U16954 ( .A(n14320), .B(n14321), .Z(n14319) );
  AND U16955 ( .A(n14322), .B(n14323), .Z(n14307) );
  NAND U16956 ( .A(n6893), .B(n6925), .Z(n14323) );
  AND U16957 ( .A(n14001), .B(n8961), .Z(n14322) );
  NAND U16958 ( .A(n9135), .B(n6919), .Z(n8961) );
  ANDN U16959 ( .A(n14321), .B(n14318), .Z(n9135) );
  ANDN U16960 ( .A(n14315), .B(n14225), .Z(n14321) );
  ANDN U16961 ( .A(n14299), .B(n14324), .Z(n14315) );
  NAND U16962 ( .A(n6984), .B(n6920), .Z(n14001) );
  ANDN U16963 ( .A(n9270), .B(n14320), .Z(n6984) );
  IV U16964 ( .A(n14325), .Z(n14320) );
  OR U16965 ( .A(n8452), .B(n8443), .Z(n6786) );
  ANDN U16966 ( .A(\u_a23_core/barrel_shift_function[1] ), .B(
        \u_a23_core/barrel_shift_function[0] ), .Z(n8443) );
  ANDN U16967 ( .A(\u_a23_core/barrel_shift_function[0] ), .B(
        \u_a23_core/barrel_shift_function[1] ), .Z(n8452) );
  NAND U16968 ( .A(n14326), .B(n6888), .Z(n14206) );
  AND U16969 ( .A(\u_a23_core/barrel_shift_function[0] ), .B(
        \u_a23_core/barrel_shift_function[1] ), .Z(n6888) );
  NAND U16970 ( .A(n14327), .B(n14328), .Z(n14326) );
  AND U16971 ( .A(n14329), .B(n14330), .Z(n14328) );
  AND U16972 ( .A(n14331), .B(n14332), .Z(n14330) );
  AND U16973 ( .A(n14333), .B(n14334), .Z(n14332) );
  AND U16974 ( .A(n14335), .B(n14336), .Z(n14334) );
  NANDN U16975 ( .B(n8593), .A(n6919), .Z(n14336) );
  NAND U16976 ( .A(n14337), .B(n14338), .Z(n6919) );
  NAND U16977 ( .A(n6778), .B(\u_a23_core/imm32[4] ), .Z(n14338) );
  AND U16978 ( .A(n14339), .B(n14340), .Z(n14337) );
  NANDN U16979 ( .B(n6453), .A(\u_a23_core/barrel_shift_data_sel[1] ), .Z(
        n14340) );
  AND U16980 ( .A(n14341), .B(n14342), .Z(n6453) );
  AND U16981 ( .A(n14343), .B(n14344), .Z(n14342) );
  AND U16982 ( .A(n14345), .B(n14346), .Z(n14344) );
  AND U16983 ( .A(n14347), .B(n14348), .Z(n14346) );
  NAND U16984 ( .A(n14349), .B(\u_a23_core/u_execute/pc[4] ), .Z(n14348) );
  NANDN U16985 ( .B(n14350), .A(\u_a23_core/u_execute/u_register_bank/r14[4] ), 
        .Z(n14347) );
  AND U16986 ( .A(n14351), .B(n14352), .Z(n14345) );
  NANDN U16987 ( .B(n14353), .A(\u_a23_core/u_execute/u_register_bank/r13[4] ), 
        .Z(n14352) );
  NANDN U16988 ( .B(n14354), .A(\u_a23_core/u_execute/u_register_bank/r12[4] ), 
        .Z(n14351) );
  AND U16989 ( .A(n14355), .B(n14356), .Z(n14343) );
  AND U16990 ( .A(n14357), .B(n14358), .Z(n14356) );
  NANDN U16991 ( .B(n14359), .A(\u_a23_core/u_execute/u_register_bank/r11[4] ), 
        .Z(n14358) );
  NANDN U16992 ( .B(n14360), .A(\u_a23_core/u_execute/u_register_bank/r10[4] ), 
        .Z(n14357) );
  AND U16993 ( .A(n14361), .B(n14362), .Z(n14355) );
  NANDN U16994 ( .B(n14363), .A(\u_a23_core/u_execute/u_register_bank/r9[4] ), 
        .Z(n14362) );
  NANDN U16995 ( .B(n14364), .A(\u_a23_core/u_execute/u_register_bank/r8[4] ), 
        .Z(n14361) );
  AND U16996 ( .A(n14365), .B(n14366), .Z(n14341) );
  AND U16997 ( .A(n14367), .B(n14368), .Z(n14366) );
  AND U16998 ( .A(n14369), .B(n14370), .Z(n14368) );
  NANDN U16999 ( .B(n14371), .A(\u_a23_core/u_execute/u_register_bank/r7[4] ), 
        .Z(n14370) );
  NANDN U17000 ( .B(n14372), .A(\u_a23_core/u_execute/u_register_bank/r6[4] ), 
        .Z(n14369) );
  AND U17001 ( .A(n14373), .B(n14374), .Z(n14367) );
  NANDN U17002 ( .B(n14375), .A(\u_a23_core/u_execute/u_register_bank/r5[4] ), 
        .Z(n14374) );
  NANDN U17003 ( .B(n14376), .A(\u_a23_core/u_execute/u_register_bank/r4[4] ), 
        .Z(n14373) );
  AND U17004 ( .A(n14377), .B(n14378), .Z(n14365) );
  AND U17005 ( .A(n14379), .B(n14380), .Z(n14378) );
  NANDN U17006 ( .B(n14381), .A(\u_a23_core/u_execute/u_register_bank/r3[4] ), 
        .Z(n14380) );
  NANDN U17007 ( .B(n14382), .A(\u_a23_core/u_execute/u_register_bank/r0[4] ), 
        .Z(n14379) );
  AND U17008 ( .A(n14383), .B(n14384), .Z(n14377) );
  NANDN U17009 ( .B(n14385), .A(\u_a23_core/u_execute/u_register_bank/r2[4] ), 
        .Z(n14384) );
  NANDN U17010 ( .B(n14386), .A(\u_a23_core/u_execute/u_register_bank/r1[4] ), 
        .Z(n14383) );
  NANDN U17011 ( .B(n14387), .A(\u_a23_core/read_data_s2[4] ), .Z(n14339) );
  NAND U17012 ( .A(n14388), .B(n14389), .Z(n8593) );
  AND U17013 ( .A(n14390), .B(n14237), .Z(n14389) );
  AND U17014 ( .A(n6990), .B(n9270), .Z(n14388) );
  NAND U17015 ( .A(n6925), .B(n8512), .Z(n14335) );
  NANDN U17016 ( .B(n6893), .A(n6892), .Z(n8512) );
  NAND U17017 ( .A(n14391), .B(n6990), .Z(n6892) );
  AND U17018 ( .A(n6988), .B(n9270), .Z(n14391) );
  AND U17019 ( .A(n14392), .B(n14325), .Z(n6893) );
  AND U17020 ( .A(n14393), .B(n14218), .Z(n14392) );
  IV U17021 ( .A(\u_a23_core/shift_imm_zero ), .Z(n14393) );
  NAND U17022 ( .A(n14394), .B(n14395), .Z(n6925) );
  NAND U17023 ( .A(n6778), .B(\u_a23_core/imm32[2] ), .Z(n14395) );
  AND U17024 ( .A(n14396), .B(n14397), .Z(n14394) );
  NANDN U17025 ( .B(n6439), .A(\u_a23_core/barrel_shift_data_sel[1] ), .Z(
        n14397) );
  AND U17026 ( .A(n14398), .B(n14399), .Z(n6439) );
  AND U17027 ( .A(n14400), .B(n14401), .Z(n14399) );
  AND U17028 ( .A(n14402), .B(n14403), .Z(n14401) );
  AND U17029 ( .A(n14404), .B(n14405), .Z(n14403) );
  NAND U17030 ( .A(\u_a23_core/u_execute/pc[2] ), .B(n14349), .Z(n14405) );
  NANDN U17031 ( .B(n14350), .A(\u_a23_core/u_execute/u_register_bank/r14[2] ), 
        .Z(n14404) );
  AND U17032 ( .A(n14406), .B(n14407), .Z(n14402) );
  NANDN U17033 ( .B(n14353), .A(\u_a23_core/u_execute/u_register_bank/r13[2] ), 
        .Z(n14407) );
  NANDN U17034 ( .B(n14354), .A(\u_a23_core/u_execute/u_register_bank/r12[2] ), 
        .Z(n14406) );
  AND U17035 ( .A(n14408), .B(n14409), .Z(n14400) );
  AND U17036 ( .A(n14410), .B(n14411), .Z(n14409) );
  NANDN U17037 ( .B(n14359), .A(\u_a23_core/u_execute/u_register_bank/r11[2] ), 
        .Z(n14411) );
  NANDN U17038 ( .B(n14360), .A(\u_a23_core/u_execute/u_register_bank/r10[2] ), 
        .Z(n14410) );
  AND U17039 ( .A(n14412), .B(n14413), .Z(n14408) );
  NANDN U17040 ( .B(n14363), .A(\u_a23_core/u_execute/u_register_bank/r9[2] ), 
        .Z(n14413) );
  NANDN U17041 ( .B(n14364), .A(\u_a23_core/u_execute/u_register_bank/r8[2] ), 
        .Z(n14412) );
  AND U17042 ( .A(n14414), .B(n14415), .Z(n14398) );
  AND U17043 ( .A(n14416), .B(n14417), .Z(n14415) );
  AND U17044 ( .A(n14418), .B(n14419), .Z(n14417) );
  NANDN U17045 ( .B(n14371), .A(\u_a23_core/u_execute/u_register_bank/r7[2] ), 
        .Z(n14419) );
  NANDN U17046 ( .B(n14372), .A(\u_a23_core/u_execute/u_register_bank/r6[2] ), 
        .Z(n14418) );
  AND U17047 ( .A(n14420), .B(n14421), .Z(n14416) );
  NANDN U17048 ( .B(n14375), .A(\u_a23_core/u_execute/u_register_bank/r5[2] ), 
        .Z(n14421) );
  NANDN U17049 ( .B(n14376), .A(\u_a23_core/u_execute/u_register_bank/r4[2] ), 
        .Z(n14420) );
  AND U17050 ( .A(n14422), .B(n14423), .Z(n14414) );
  AND U17051 ( .A(n14424), .B(n14425), .Z(n14423) );
  NANDN U17052 ( .B(n14381), .A(\u_a23_core/u_execute/u_register_bank/r3[2] ), 
        .Z(n14425) );
  NANDN U17053 ( .B(n14382), .A(\u_a23_core/u_execute/u_register_bank/r0[2] ), 
        .Z(n14424) );
  AND U17054 ( .A(n14426), .B(n14427), .Z(n14422) );
  NANDN U17055 ( .B(n14385), .A(\u_a23_core/u_execute/u_register_bank/r2[2] ), 
        .Z(n14427) );
  NANDN U17056 ( .B(n14386), .A(\u_a23_core/u_execute/u_register_bank/r1[2] ), 
        .Z(n14426) );
  NANDN U17057 ( .B(n14387), .A(\u_a23_core/read_data_s2[2] ), .Z(n14396) );
  AND U17058 ( .A(n14428), .B(n14429), .Z(n14333) );
  NAND U17059 ( .A(n6920), .B(n6897), .Z(n14429) );
  NANDN U17060 ( .B(\u_a23_core/shift_imm_zero ), .A(n14430), .Z(n6897) );
  NAND U17061 ( .A(n6988), .B(n9271), .Z(n14430) );
  NAND U17062 ( .A(n14431), .B(n14432), .Z(n6920) );
  NAND U17063 ( .A(n6778), .B(\u_a23_core/imm32[3] ), .Z(n14432) );
  AND U17064 ( .A(n14433), .B(n14434), .Z(n14431) );
  NANDN U17065 ( .B(n6446), .A(\u_a23_core/barrel_shift_data_sel[1] ), .Z(
        n14434) );
  AND U17066 ( .A(n14435), .B(n14436), .Z(n6446) );
  AND U17067 ( .A(n14437), .B(n14438), .Z(n14436) );
  AND U17068 ( .A(n14439), .B(n14440), .Z(n14438) );
  AND U17069 ( .A(n14441), .B(n14442), .Z(n14440) );
  NAND U17070 ( .A(n14349), .B(\u_a23_core/u_execute/pc[3] ), .Z(n14442) );
  NANDN U17071 ( .B(n14350), .A(\u_a23_core/u_execute/u_register_bank/r14[3] ), 
        .Z(n14441) );
  AND U17072 ( .A(n14443), .B(n14444), .Z(n14439) );
  NANDN U17073 ( .B(n14353), .A(\u_a23_core/u_execute/u_register_bank/r13[3] ), 
        .Z(n14444) );
  NANDN U17074 ( .B(n14354), .A(\u_a23_core/u_execute/u_register_bank/r12[3] ), 
        .Z(n14443) );
  AND U17075 ( .A(n14445), .B(n14446), .Z(n14437) );
  AND U17076 ( .A(n14447), .B(n14448), .Z(n14446) );
  NANDN U17077 ( .B(n14359), .A(\u_a23_core/u_execute/u_register_bank/r11[3] ), 
        .Z(n14448) );
  NANDN U17078 ( .B(n14360), .A(\u_a23_core/u_execute/u_register_bank/r10[3] ), 
        .Z(n14447) );
  AND U17079 ( .A(n14449), .B(n14450), .Z(n14445) );
  NANDN U17080 ( .B(n14363), .A(\u_a23_core/u_execute/u_register_bank/r9[3] ), 
        .Z(n14450) );
  NANDN U17081 ( .B(n14364), .A(\u_a23_core/u_execute/u_register_bank/r8[3] ), 
        .Z(n14449) );
  AND U17082 ( .A(n14451), .B(n14452), .Z(n14435) );
  AND U17083 ( .A(n14453), .B(n14454), .Z(n14452) );
  AND U17084 ( .A(n14455), .B(n14456), .Z(n14454) );
  NANDN U17085 ( .B(n14371), .A(\u_a23_core/u_execute/u_register_bank/r7[3] ), 
        .Z(n14456) );
  NANDN U17086 ( .B(n14372), .A(\u_a23_core/u_execute/u_register_bank/r6[3] ), 
        .Z(n14455) );
  AND U17087 ( .A(n14457), .B(n14458), .Z(n14453) );
  NANDN U17088 ( .B(n14375), .A(\u_a23_core/u_execute/u_register_bank/r5[3] ), 
        .Z(n14458) );
  NANDN U17089 ( .B(n14376), .A(\u_a23_core/u_execute/u_register_bank/r4[3] ), 
        .Z(n14457) );
  AND U17090 ( .A(n14459), .B(n14460), .Z(n14451) );
  AND U17091 ( .A(n14461), .B(n14462), .Z(n14460) );
  NANDN U17092 ( .B(n14381), .A(\u_a23_core/u_execute/u_register_bank/r3[3] ), 
        .Z(n14462) );
  NANDN U17093 ( .B(n14382), .A(\u_a23_core/u_execute/u_register_bank/r0[3] ), 
        .Z(n14461) );
  AND U17094 ( .A(n14463), .B(n14464), .Z(n14459) );
  NANDN U17095 ( .B(n14385), .A(\u_a23_core/u_execute/u_register_bank/r2[3] ), 
        .Z(n14464) );
  NANDN U17096 ( .B(n14386), .A(\u_a23_core/u_execute/u_register_bank/r1[3] ), 
        .Z(n14463) );
  NANDN U17097 ( .B(n14387), .A(\u_a23_core/read_data_s2[3] ), .Z(n14433) );
  NANDN U17098 ( .B(n8516), .A(n6926), .Z(n14428) );
  NAND U17099 ( .A(n14465), .B(n14466), .Z(n6926) );
  NAND U17100 ( .A(n6778), .B(\u_a23_core/imm32[1] ), .Z(n14466) );
  AND U17101 ( .A(n14467), .B(n14468), .Z(n14465) );
  NANDN U17102 ( .B(n6432), .A(\u_a23_core/barrel_shift_data_sel[1] ), .Z(
        n14468) );
  AND U17103 ( .A(n14469), .B(n14470), .Z(n6432) );
  AND U17104 ( .A(n14471), .B(n14472), .Z(n14470) );
  AND U17105 ( .A(n14473), .B(n14474), .Z(n14472) );
  AND U17106 ( .A(n14475), .B(n14476), .Z(n14474) );
  NANDN U17107 ( .B(n14350), .A(\u_a23_core/u_execute/u_register_bank/r14[1] ), 
        .Z(n14476) );
  NANDN U17108 ( .B(n14353), .A(\u_a23_core/u_execute/u_register_bank/r13[1] ), 
        .Z(n14475) );
  AND U17109 ( .A(n14477), .B(n14478), .Z(n14473) );
  NANDN U17110 ( .B(n14354), .A(\u_a23_core/u_execute/u_register_bank/r12[1] ), 
        .Z(n14478) );
  NANDN U17111 ( .B(n14359), .A(\u_a23_core/u_execute/u_register_bank/r11[1] ), 
        .Z(n14477) );
  AND U17112 ( .A(n14479), .B(n14480), .Z(n14471) );
  AND U17113 ( .A(n14481), .B(n14482), .Z(n14480) );
  NANDN U17114 ( .B(n14360), .A(\u_a23_core/u_execute/u_register_bank/r10[1] ), 
        .Z(n14482) );
  NANDN U17115 ( .B(n14363), .A(\u_a23_core/u_execute/u_register_bank/r9[1] ), 
        .Z(n14481) );
  AND U17116 ( .A(n14483), .B(n14484), .Z(n14479) );
  NANDN U17117 ( .B(n14364), .A(\u_a23_core/u_execute/u_register_bank/r8[1] ), 
        .Z(n14484) );
  NANDN U17118 ( .B(n14371), .A(\u_a23_core/u_execute/u_register_bank/r7[1] ), 
        .Z(n14483) );
  AND U17119 ( .A(n14485), .B(n14486), .Z(n14469) );
  AND U17120 ( .A(n14487), .B(n14488), .Z(n14486) );
  AND U17121 ( .A(n14489), .B(n14490), .Z(n14488) );
  NANDN U17122 ( .B(n14372), .A(\u_a23_core/u_execute/u_register_bank/r6[1] ), 
        .Z(n14490) );
  NANDN U17123 ( .B(n14375), .A(\u_a23_core/u_execute/u_register_bank/r5[1] ), 
        .Z(n14489) );
  AND U17124 ( .A(n14491), .B(n14492), .Z(n14487) );
  NANDN U17125 ( .B(n14376), .A(\u_a23_core/u_execute/u_register_bank/r4[1] ), 
        .Z(n14492) );
  NANDN U17126 ( .B(n14381), .A(\u_a23_core/u_execute/u_register_bank/r3[1] ), 
        .Z(n14491) );
  AND U17127 ( .A(n14493), .B(n14494), .Z(n14485) );
  NANDN U17128 ( .B(n14386), .A(\u_a23_core/u_execute/u_register_bank/r1[1] ), 
        .Z(n14494) );
  AND U17129 ( .A(n14495), .B(n14496), .Z(n14493) );
  NANDN U17130 ( .B(n14382), .A(\u_a23_core/u_execute/u_register_bank/r0[1] ), 
        .Z(n14496) );
  NANDN U17131 ( .B(n14385), .A(\u_a23_core/u_execute/u_register_bank/r2[1] ), 
        .Z(n14495) );
  NANDN U17132 ( .B(n14387), .A(\u_a23_core/read_data_s2[1] ), .Z(n14467) );
  NAND U17133 ( .A(n14497), .B(n14498), .Z(n8516) );
  AND U17134 ( .A(n14305), .B(n14225), .Z(n14497) );
  AND U17135 ( .A(n14499), .B(n14500), .Z(n14331) );
  AND U17136 ( .A(n14501), .B(n14502), .Z(n14500) );
  NANDN U17137 ( .B(n8522), .A(n6898), .Z(n14502) );
  NAND U17138 ( .A(n14503), .B(n14504), .Z(n6898) );
  NAND U17139 ( .A(n6778), .B(\u_a23_core/imm32[0] ), .Z(n14504) );
  AND U17140 ( .A(n14505), .B(n14506), .Z(n14503) );
  NANDN U17141 ( .B(n6424), .A(\u_a23_core/barrel_shift_data_sel[1] ), .Z(
        n14506) );
  AND U17142 ( .A(n14507), .B(n14508), .Z(n6424) );
  AND U17143 ( .A(n14509), .B(n14510), .Z(n14508) );
  AND U17144 ( .A(n14511), .B(n14512), .Z(n14510) );
  AND U17145 ( .A(n14513), .B(n14514), .Z(n14512) );
  NANDN U17146 ( .B(n14350), .A(\u_a23_core/u_execute/u_register_bank/r14[0] ), 
        .Z(n14514) );
  NANDN U17147 ( .B(n14353), .A(\u_a23_core/u_execute/u_register_bank/r13[0] ), 
        .Z(n14513) );
  AND U17148 ( .A(n14515), .B(n14516), .Z(n14511) );
  NANDN U17149 ( .B(n14354), .A(\u_a23_core/u_execute/u_register_bank/r12[0] ), 
        .Z(n14516) );
  NANDN U17150 ( .B(n14359), .A(\u_a23_core/u_execute/u_register_bank/r11[0] ), 
        .Z(n14515) );
  AND U17151 ( .A(n14517), .B(n14518), .Z(n14509) );
  AND U17152 ( .A(n14519), .B(n14520), .Z(n14518) );
  NANDN U17153 ( .B(n14360), .A(\u_a23_core/u_execute/u_register_bank/r10[0] ), 
        .Z(n14520) );
  NANDN U17154 ( .B(n14363), .A(\u_a23_core/u_execute/u_register_bank/r9[0] ), 
        .Z(n14519) );
  AND U17155 ( .A(n14521), .B(n14522), .Z(n14517) );
  NANDN U17156 ( .B(n14364), .A(\u_a23_core/u_execute/u_register_bank/r8[0] ), 
        .Z(n14522) );
  NANDN U17157 ( .B(n14371), .A(\u_a23_core/u_execute/u_register_bank/r7[0] ), 
        .Z(n14521) );
  AND U17158 ( .A(n14523), .B(n14524), .Z(n14507) );
  AND U17159 ( .A(n14525), .B(n14526), .Z(n14524) );
  AND U17160 ( .A(n14527), .B(n14528), .Z(n14526) );
  NANDN U17161 ( .B(n14372), .A(\u_a23_core/u_execute/u_register_bank/r6[0] ), 
        .Z(n14528) );
  NANDN U17162 ( .B(n14375), .A(\u_a23_core/u_execute/u_register_bank/r5[0] ), 
        .Z(n14527) );
  AND U17163 ( .A(n14529), .B(n14530), .Z(n14525) );
  NANDN U17164 ( .B(n14376), .A(\u_a23_core/u_execute/u_register_bank/r4[0] ), 
        .Z(n14530) );
  NANDN U17165 ( .B(n14381), .A(\u_a23_core/u_execute/u_register_bank/r3[0] ), 
        .Z(n14529) );
  AND U17166 ( .A(n14531), .B(n14532), .Z(n14523) );
  NANDN U17167 ( .B(n14386), .A(\u_a23_core/u_execute/u_register_bank/r1[0] ), 
        .Z(n14532) );
  AND U17168 ( .A(n14533), .B(n14534), .Z(n14531) );
  NANDN U17169 ( .B(n14382), .A(\u_a23_core/u_execute/u_register_bank/r0[0] ), 
        .Z(n14534) );
  NANDN U17170 ( .B(n14385), .A(\u_a23_core/u_execute/u_register_bank/r2[0] ), 
        .Z(n14533) );
  NANDN U17171 ( .B(n14387), .A(\u_a23_core/read_data_s2[0] ), .Z(n14505) );
  NAND U17172 ( .A(n14218), .B(n14498), .Z(n8522) );
  NANDN U17173 ( .B(n8526), .A(n6882), .Z(n14501) );
  NAND U17174 ( .A(n14535), .B(n14536), .Z(n6882) );
  NAND U17175 ( .A(\u_a23_core/imm32[31] ), .B(n6778), .Z(n14536) );
  AND U17176 ( .A(n14537), .B(n14538), .Z(n14535) );
  NANDN U17177 ( .B(n6643), .A(\u_a23_core/barrel_shift_data_sel[1] ), .Z(
        n14538) );
  AND U17178 ( .A(n14539), .B(n14540), .Z(n6643) );
  AND U17179 ( .A(n14541), .B(n14542), .Z(n14540) );
  AND U17180 ( .A(n14543), .B(n14544), .Z(n14542) );
  AND U17181 ( .A(n14545), .B(n14546), .Z(n14544) );
  NAND U17182 ( .A(\u_a23_core/u_execute/save_int_pc_m4[31] ), .B(n14349), .Z(
        n14546) );
  NANDN U17183 ( .B(n14350), .A(\u_a23_core/u_execute/u_register_bank/r14[31] ), .Z(n14545) );
  AND U17184 ( .A(n14547), .B(n14548), .Z(n14543) );
  NANDN U17185 ( .B(n14353), .A(\u_a23_core/u_execute/u_register_bank/r13[31] ), .Z(n14548) );
  NANDN U17186 ( .B(n14354), .A(\u_a23_core/u_execute/u_register_bank/r12[31] ), .Z(n14547) );
  AND U17187 ( .A(n14549), .B(n14550), .Z(n14541) );
  AND U17188 ( .A(n14551), .B(n14552), .Z(n14550) );
  NANDN U17189 ( .B(n14359), .A(\u_a23_core/u_execute/u_register_bank/r11[31] ), .Z(n14552) );
  NANDN U17190 ( .B(n14360), .A(\u_a23_core/u_execute/u_register_bank/r10[31] ), .Z(n14551) );
  AND U17191 ( .A(n14553), .B(n14554), .Z(n14549) );
  NANDN U17192 ( .B(n14363), .A(\u_a23_core/u_execute/u_register_bank/r9[31] ), 
        .Z(n14554) );
  NANDN U17193 ( .B(n14364), .A(\u_a23_core/u_execute/u_register_bank/r8[31] ), 
        .Z(n14553) );
  AND U17194 ( .A(n14555), .B(n14556), .Z(n14539) );
  AND U17195 ( .A(n14557), .B(n14558), .Z(n14556) );
  AND U17196 ( .A(n14559), .B(n14560), .Z(n14558) );
  NANDN U17197 ( .B(n14371), .A(\u_a23_core/u_execute/u_register_bank/r7[31] ), 
        .Z(n14560) );
  NANDN U17198 ( .B(n14372), .A(\u_a23_core/u_execute/u_register_bank/r6[31] ), 
        .Z(n14559) );
  AND U17199 ( .A(n14561), .B(n14562), .Z(n14557) );
  NANDN U17200 ( .B(n14375), .A(\u_a23_core/u_execute/u_register_bank/r5[31] ), 
        .Z(n14562) );
  NANDN U17201 ( .B(n14376), .A(\u_a23_core/u_execute/u_register_bank/r4[31] ), 
        .Z(n14561) );
  AND U17202 ( .A(n14563), .B(n14564), .Z(n14555) );
  AND U17203 ( .A(n14565), .B(n14566), .Z(n14564) );
  NANDN U17204 ( .B(n14381), .A(\u_a23_core/u_execute/u_register_bank/r3[31] ), 
        .Z(n14566) );
  NANDN U17205 ( .B(n14382), .A(\u_a23_core/u_execute/u_register_bank/r0[31] ), 
        .Z(n14565) );
  AND U17206 ( .A(n14567), .B(n14568), .Z(n14563) );
  NANDN U17207 ( .B(n14385), .A(\u_a23_core/u_execute/u_register_bank/r2[31] ), 
        .Z(n14568) );
  NANDN U17208 ( .B(n14386), .A(\u_a23_core/u_execute/u_register_bank/r1[31] ), 
        .Z(n14567) );
  NANDN U17209 ( .B(n14387), .A(\u_a23_core/read_data_s2[31] ), .Z(n14537) );
  NAND U17210 ( .A(n14205), .B(n14498), .Z(n8526) );
  ANDN U17211 ( .A(n14294), .B(n14569), .Z(n14498) );
  IV U17212 ( .A(n14570), .Z(n14569) );
  AND U17213 ( .A(n14571), .B(n14324), .Z(n14294) );
  NAND U17214 ( .A(n14218), .B(n14205), .Z(n14571) );
  AND U17215 ( .A(n14572), .B(n14573), .Z(n14499) );
  NANDN U17216 ( .B(n8534), .A(n6809), .Z(n14573) );
  NAND U17217 ( .A(n14574), .B(n14575), .Z(n6809) );
  NAND U17218 ( .A(n6778), .B(\u_a23_core/imm32[30] ), .Z(n14575) );
  AND U17219 ( .A(n14576), .B(n14577), .Z(n14574) );
  NANDN U17220 ( .B(n6635), .A(\u_a23_core/barrel_shift_data_sel[1] ), .Z(
        n14577) );
  AND U17221 ( .A(n14578), .B(n14579), .Z(n6635) );
  AND U17222 ( .A(n14580), .B(n14581), .Z(n14579) );
  AND U17223 ( .A(n14582), .B(n14583), .Z(n14581) );
  AND U17224 ( .A(n14584), .B(n14585), .Z(n14583) );
  NAND U17225 ( .A(\u_a23_core/u_execute/save_int_pc_m4[30] ), .B(n14349), .Z(
        n14585) );
  NANDN U17226 ( .B(n14350), .A(\u_a23_core/u_execute/u_register_bank/r14[30] ), .Z(n14584) );
  AND U17227 ( .A(n14586), .B(n14587), .Z(n14582) );
  NANDN U17228 ( .B(n14353), .A(\u_a23_core/u_execute/u_register_bank/r13[30] ), .Z(n14587) );
  NANDN U17229 ( .B(n14354), .A(\u_a23_core/u_execute/u_register_bank/r12[30] ), .Z(n14586) );
  AND U17230 ( .A(n14588), .B(n14589), .Z(n14580) );
  AND U17231 ( .A(n14590), .B(n14591), .Z(n14589) );
  NANDN U17232 ( .B(n14359), .A(\u_a23_core/u_execute/u_register_bank/r11[30] ), .Z(n14591) );
  NANDN U17233 ( .B(n14360), .A(\u_a23_core/u_execute/u_register_bank/r10[30] ), .Z(n14590) );
  AND U17234 ( .A(n14592), .B(n14593), .Z(n14588) );
  NANDN U17235 ( .B(n14363), .A(\u_a23_core/u_execute/u_register_bank/r9[30] ), 
        .Z(n14593) );
  NANDN U17236 ( .B(n14364), .A(\u_a23_core/u_execute/u_register_bank/r8[30] ), 
        .Z(n14592) );
  AND U17237 ( .A(n14594), .B(n14595), .Z(n14578) );
  AND U17238 ( .A(n14596), .B(n14597), .Z(n14595) );
  AND U17239 ( .A(n14598), .B(n14599), .Z(n14597) );
  NANDN U17240 ( .B(n14371), .A(\u_a23_core/u_execute/u_register_bank/r7[30] ), 
        .Z(n14599) );
  NANDN U17241 ( .B(n14372), .A(\u_a23_core/u_execute/u_register_bank/r6[30] ), 
        .Z(n14598) );
  AND U17242 ( .A(n14600), .B(n14601), .Z(n14596) );
  NANDN U17243 ( .B(n14375), .A(\u_a23_core/u_execute/u_register_bank/r5[30] ), 
        .Z(n14601) );
  NANDN U17244 ( .B(n14376), .A(\u_a23_core/u_execute/u_register_bank/r4[30] ), 
        .Z(n14600) );
  AND U17245 ( .A(n14602), .B(n14603), .Z(n14594) );
  AND U17246 ( .A(n14604), .B(n14605), .Z(n14603) );
  NANDN U17247 ( .B(n14381), .A(\u_a23_core/u_execute/u_register_bank/r3[30] ), 
        .Z(n14605) );
  NANDN U17248 ( .B(n14382), .A(\u_a23_core/u_execute/u_register_bank/r0[30] ), 
        .Z(n14604) );
  AND U17249 ( .A(n14606), .B(n14607), .Z(n14602) );
  NANDN U17250 ( .B(n14385), .A(\u_a23_core/u_execute/u_register_bank/r2[30] ), 
        .Z(n14607) );
  NANDN U17251 ( .B(n14386), .A(\u_a23_core/u_execute/u_register_bank/r1[30] ), 
        .Z(n14606) );
  NANDN U17252 ( .B(n14387), .A(\u_a23_core/read_data_s2[30] ), .Z(n14576) );
  NAND U17253 ( .A(n14570), .B(n14317), .Z(n8534) );
  AND U17254 ( .A(n14218), .B(n14205), .Z(n14317) );
  NANDN U17255 ( .B(n8511), .A(n6807), .Z(n14572) );
  NAND U17256 ( .A(n14608), .B(n14609), .Z(n6807) );
  NAND U17257 ( .A(n6778), .B(\u_a23_core/imm32[29] ), .Z(n14609) );
  AND U17258 ( .A(n14610), .B(n14611), .Z(n14608) );
  NANDN U17259 ( .B(n6628), .A(\u_a23_core/barrel_shift_data_sel[1] ), .Z(
        n14611) );
  AND U17260 ( .A(n14612), .B(n14613), .Z(n6628) );
  AND U17261 ( .A(n14614), .B(n14615), .Z(n14613) );
  AND U17262 ( .A(n14616), .B(n14617), .Z(n14615) );
  AND U17263 ( .A(n14618), .B(n14619), .Z(n14617) );
  NAND U17264 ( .A(\u_a23_core/u_execute/save_int_pc_m4[29] ), .B(n14349), .Z(
        n14619) );
  NANDN U17265 ( .B(n14350), .A(\u_a23_core/u_execute/u_register_bank/r14[29] ), .Z(n14618) );
  AND U17266 ( .A(n14620), .B(n14621), .Z(n14616) );
  NANDN U17267 ( .B(n14353), .A(\u_a23_core/u_execute/u_register_bank/r13[29] ), .Z(n14621) );
  NANDN U17268 ( .B(n14354), .A(\u_a23_core/u_execute/u_register_bank/r12[29] ), .Z(n14620) );
  AND U17269 ( .A(n14622), .B(n14623), .Z(n14614) );
  AND U17270 ( .A(n14624), .B(n14625), .Z(n14623) );
  NANDN U17271 ( .B(n14359), .A(\u_a23_core/u_execute/u_register_bank/r11[29] ), .Z(n14625) );
  NANDN U17272 ( .B(n14360), .A(\u_a23_core/u_execute/u_register_bank/r10[29] ), .Z(n14624) );
  AND U17273 ( .A(n14626), .B(n14627), .Z(n14622) );
  NANDN U17274 ( .B(n14363), .A(\u_a23_core/u_execute/u_register_bank/r9[29] ), 
        .Z(n14627) );
  NANDN U17275 ( .B(n14364), .A(\u_a23_core/u_execute/u_register_bank/r8[29] ), 
        .Z(n14626) );
  AND U17276 ( .A(n14628), .B(n14629), .Z(n14612) );
  AND U17277 ( .A(n14630), .B(n14631), .Z(n14629) );
  AND U17278 ( .A(n14632), .B(n14633), .Z(n14631) );
  NANDN U17279 ( .B(n14371), .A(\u_a23_core/u_execute/u_register_bank/r7[29] ), 
        .Z(n14633) );
  NANDN U17280 ( .B(n14372), .A(\u_a23_core/u_execute/u_register_bank/r6[29] ), 
        .Z(n14632) );
  AND U17281 ( .A(n14634), .B(n14635), .Z(n14630) );
  NANDN U17282 ( .B(n14375), .A(\u_a23_core/u_execute/u_register_bank/r5[29] ), 
        .Z(n14635) );
  NANDN U17283 ( .B(n14376), .A(\u_a23_core/u_execute/u_register_bank/r4[29] ), 
        .Z(n14634) );
  AND U17284 ( .A(n14636), .B(n14637), .Z(n14628) );
  AND U17285 ( .A(n14638), .B(n14639), .Z(n14637) );
  NANDN U17286 ( .B(n14381), .A(\u_a23_core/u_execute/u_register_bank/r3[29] ), 
        .Z(n14639) );
  NANDN U17287 ( .B(n14382), .A(\u_a23_core/u_execute/u_register_bank/r0[29] ), 
        .Z(n14638) );
  AND U17288 ( .A(n14640), .B(n14641), .Z(n14636) );
  NANDN U17289 ( .B(n14385), .A(\u_a23_core/u_execute/u_register_bank/r2[29] ), 
        .Z(n14641) );
  NANDN U17290 ( .B(n14386), .A(\u_a23_core/u_execute/u_register_bank/r1[29] ), 
        .Z(n14640) );
  NANDN U17291 ( .B(n14387), .A(\u_a23_core/read_data_s2[29] ), .Z(n14610) );
  NAND U17292 ( .A(n14237), .B(n14570), .Z(n8511) );
  AND U17293 ( .A(n14642), .B(n14284), .Z(n14570) );
  ANDN U17294 ( .A(n14390), .B(n14240), .Z(n14284) );
  AND U17295 ( .A(n14643), .B(n14644), .Z(n14329) );
  AND U17296 ( .A(n14645), .B(n14646), .Z(n14644) );
  AND U17297 ( .A(n14647), .B(n14648), .Z(n14646) );
  NANDN U17298 ( .B(n8515), .A(n6799), .Z(n14648) );
  NAND U17299 ( .A(n14649), .B(n14650), .Z(n6799) );
  NAND U17300 ( .A(n6778), .B(\u_a23_core/imm32[28] ), .Z(n14650) );
  AND U17301 ( .A(n14651), .B(n14652), .Z(n14649) );
  NANDN U17302 ( .B(n6621), .A(\u_a23_core/barrel_shift_data_sel[1] ), .Z(
        n14652) );
  AND U17303 ( .A(n14653), .B(n14654), .Z(n6621) );
  AND U17304 ( .A(n14655), .B(n14656), .Z(n14654) );
  AND U17305 ( .A(n14657), .B(n14658), .Z(n14656) );
  AND U17306 ( .A(n14659), .B(n14660), .Z(n14658) );
  NAND U17307 ( .A(\u_a23_core/u_execute/save_int_pc_m4[28] ), .B(n14349), .Z(
        n14660) );
  NANDN U17308 ( .B(n14350), .A(\u_a23_core/u_execute/u_register_bank/r14[28] ), .Z(n14659) );
  AND U17309 ( .A(n14661), .B(n14662), .Z(n14657) );
  NANDN U17310 ( .B(n14353), .A(\u_a23_core/u_execute/u_register_bank/r13[28] ), .Z(n14662) );
  NANDN U17311 ( .B(n14354), .A(\u_a23_core/u_execute/u_register_bank/r12[28] ), .Z(n14661) );
  AND U17312 ( .A(n14663), .B(n14664), .Z(n14655) );
  AND U17313 ( .A(n14665), .B(n14666), .Z(n14664) );
  NANDN U17314 ( .B(n14359), .A(\u_a23_core/u_execute/u_register_bank/r11[28] ), .Z(n14666) );
  NANDN U17315 ( .B(n14360), .A(\u_a23_core/u_execute/u_register_bank/r10[28] ), .Z(n14665) );
  AND U17316 ( .A(n14667), .B(n14668), .Z(n14663) );
  NANDN U17317 ( .B(n14363), .A(\u_a23_core/u_execute/u_register_bank/r9[28] ), 
        .Z(n14668) );
  NANDN U17318 ( .B(n14364), .A(\u_a23_core/u_execute/u_register_bank/r8[28] ), 
        .Z(n14667) );
  AND U17319 ( .A(n14669), .B(n14670), .Z(n14653) );
  AND U17320 ( .A(n14671), .B(n14672), .Z(n14670) );
  AND U17321 ( .A(n14673), .B(n14674), .Z(n14672) );
  NANDN U17322 ( .B(n14371), .A(\u_a23_core/u_execute/u_register_bank/r7[28] ), 
        .Z(n14674) );
  NANDN U17323 ( .B(n14372), .A(\u_a23_core/u_execute/u_register_bank/r6[28] ), 
        .Z(n14673) );
  AND U17324 ( .A(n14675), .B(n14676), .Z(n14671) );
  NANDN U17325 ( .B(n14375), .A(\u_a23_core/u_execute/u_register_bank/r5[28] ), 
        .Z(n14676) );
  NANDN U17326 ( .B(n14376), .A(\u_a23_core/u_execute/u_register_bank/r4[28] ), 
        .Z(n14675) );
  AND U17327 ( .A(n14677), .B(n14678), .Z(n14669) );
  AND U17328 ( .A(n14679), .B(n14680), .Z(n14678) );
  NANDN U17329 ( .B(n14381), .A(\u_a23_core/u_execute/u_register_bank/r3[28] ), 
        .Z(n14680) );
  NANDN U17330 ( .B(n14382), .A(\u_a23_core/u_execute/u_register_bank/r0[28] ), 
        .Z(n14679) );
  AND U17331 ( .A(n14681), .B(n14682), .Z(n14677) );
  NANDN U17332 ( .B(n14385), .A(\u_a23_core/u_execute/u_register_bank/r2[28] ), 
        .Z(n14682) );
  NANDN U17333 ( .B(n14386), .A(\u_a23_core/u_execute/u_register_bank/r1[28] ), 
        .Z(n14681) );
  NANDN U17334 ( .B(n14387), .A(\u_a23_core/read_data_s2[28] ), .Z(n14651) );
  NAND U17335 ( .A(n14240), .B(n14642), .Z(n8515) );
  ANDN U17336 ( .A(n14237), .B(n14225), .Z(n14240) );
  NANDN U17337 ( .B(n8521), .A(n6803), .Z(n14647) );
  NAND U17338 ( .A(n14683), .B(n14684), .Z(n6803) );
  NAND U17339 ( .A(n6778), .B(\u_a23_core/imm32[27] ), .Z(n14684) );
  AND U17340 ( .A(n14685), .B(n14686), .Z(n14683) );
  NANDN U17341 ( .B(n6614), .A(\u_a23_core/barrel_shift_data_sel[1] ), .Z(
        n14686) );
  AND U17342 ( .A(n14687), .B(n14688), .Z(n6614) );
  AND U17343 ( .A(n14689), .B(n14690), .Z(n14688) );
  AND U17344 ( .A(n14691), .B(n14692), .Z(n14690) );
  ANDN U17345 ( .A(n14693), .B(n14349), .Z(n14692) );
  NANDN U17346 ( .B(n14350), .A(\u_a23_core/u_execute/u_register_bank/r14[27] ), .Z(n14693) );
  AND U17347 ( .A(n14694), .B(n14695), .Z(n14691) );
  NANDN U17348 ( .B(n14353), .A(\u_a23_core/u_execute/u_register_bank/r13[27] ), .Z(n14695) );
  NANDN U17349 ( .B(n14354), .A(\u_a23_core/u_execute/u_register_bank/r12[27] ), .Z(n14694) );
  AND U17350 ( .A(n14696), .B(n14697), .Z(n14689) );
  AND U17351 ( .A(n14698), .B(n14699), .Z(n14697) );
  NANDN U17352 ( .B(n14359), .A(\u_a23_core/u_execute/u_register_bank/r11[27] ), .Z(n14699) );
  NANDN U17353 ( .B(n14360), .A(\u_a23_core/u_execute/u_register_bank/r10[27] ), .Z(n14698) );
  AND U17354 ( .A(n14700), .B(n14701), .Z(n14696) );
  NANDN U17355 ( .B(n14363), .A(\u_a23_core/u_execute/u_register_bank/r9[27] ), 
        .Z(n14701) );
  NANDN U17356 ( .B(n14364), .A(\u_a23_core/u_execute/u_register_bank/r8[27] ), 
        .Z(n14700) );
  AND U17357 ( .A(n14702), .B(n14703), .Z(n14687) );
  AND U17358 ( .A(n14704), .B(n14705), .Z(n14703) );
  AND U17359 ( .A(n14706), .B(n14707), .Z(n14705) );
  NANDN U17360 ( .B(n14371), .A(\u_a23_core/u_execute/u_register_bank/r7[27] ), 
        .Z(n14707) );
  NANDN U17361 ( .B(n14372), .A(\u_a23_core/u_execute/u_register_bank/r6[27] ), 
        .Z(n14706) );
  AND U17362 ( .A(n14708), .B(n14709), .Z(n14704) );
  NANDN U17363 ( .B(n14375), .A(\u_a23_core/u_execute/u_register_bank/r5[27] ), 
        .Z(n14709) );
  NANDN U17364 ( .B(n14376), .A(\u_a23_core/u_execute/u_register_bank/r4[27] ), 
        .Z(n14708) );
  AND U17365 ( .A(n14710), .B(n14711), .Z(n14702) );
  AND U17366 ( .A(n14712), .B(n14713), .Z(n14711) );
  NANDN U17367 ( .B(n14381), .A(\u_a23_core/u_execute/u_register_bank/r3[27] ), 
        .Z(n14713) );
  NANDN U17368 ( .B(n14382), .A(\u_a23_core/u_execute/u_register_bank/r0[27] ), 
        .Z(n14712) );
  AND U17369 ( .A(n14714), .B(n14715), .Z(n14710) );
  NANDN U17370 ( .B(n14385), .A(\u_a23_core/u_execute/u_register_bank/r2[27] ), 
        .Z(n14715) );
  NANDN U17371 ( .B(n14386), .A(\u_a23_core/u_execute/u_register_bank/r1[27] ), 
        .Z(n14714) );
  NANDN U17372 ( .B(n14387), .A(\u_a23_core/read_data_s2[27] ), .Z(n14685) );
  NAND U17373 ( .A(n6988), .B(n14642), .Z(n8521) );
  AND U17374 ( .A(n14716), .B(n14717), .Z(n14642) );
  AND U17375 ( .A(n14718), .B(n14719), .Z(n14716) );
  IV U17376 ( .A(n14255), .Z(n14719) );
  AND U17377 ( .A(n14720), .B(n14721), .Z(n14645) );
  NANDN U17378 ( .B(n8525), .A(n6823), .Z(n14721) );
  NAND U17379 ( .A(n14722), .B(n14723), .Z(n6823) );
  NAND U17380 ( .A(n6778), .B(\u_a23_core/imm32[26] ), .Z(n14723) );
  AND U17381 ( .A(n14724), .B(n14725), .Z(n14722) );
  NANDN U17382 ( .B(n6607), .A(\u_a23_core/barrel_shift_data_sel[1] ), .Z(
        n14725) );
  AND U17383 ( .A(n14726), .B(n14727), .Z(n6607) );
  AND U17384 ( .A(n14728), .B(n14729), .Z(n14727) );
  AND U17385 ( .A(n14730), .B(n14731), .Z(n14729) );
  ANDN U17386 ( .A(n14732), .B(n14349), .Z(n14731) );
  NANDN U17387 ( .B(n14350), .A(\u_a23_core/u_execute/u_register_bank/r14[26] ), .Z(n14732) );
  AND U17388 ( .A(n14733), .B(n14734), .Z(n14730) );
  NANDN U17389 ( .B(n14353), .A(\u_a23_core/u_execute/u_register_bank/r13[26] ), .Z(n14734) );
  NANDN U17390 ( .B(n14354), .A(\u_a23_core/u_execute/u_register_bank/r12[26] ), .Z(n14733) );
  AND U17391 ( .A(n14735), .B(n14736), .Z(n14728) );
  AND U17392 ( .A(n14737), .B(n14738), .Z(n14736) );
  NANDN U17393 ( .B(n14359), .A(\u_a23_core/u_execute/u_register_bank/r11[26] ), .Z(n14738) );
  NANDN U17394 ( .B(n14360), .A(\u_a23_core/u_execute/u_register_bank/r10[26] ), .Z(n14737) );
  AND U17395 ( .A(n14739), .B(n14740), .Z(n14735) );
  NANDN U17396 ( .B(n14363), .A(\u_a23_core/u_execute/u_register_bank/r9[26] ), 
        .Z(n14740) );
  NANDN U17397 ( .B(n14364), .A(\u_a23_core/u_execute/u_register_bank/r8[26] ), 
        .Z(n14739) );
  AND U17398 ( .A(n14741), .B(n14742), .Z(n14726) );
  AND U17399 ( .A(n14743), .B(n14744), .Z(n14742) );
  AND U17400 ( .A(n14745), .B(n14746), .Z(n14744) );
  NANDN U17401 ( .B(n14371), .A(\u_a23_core/u_execute/u_register_bank/r7[26] ), 
        .Z(n14746) );
  NANDN U17402 ( .B(n14372), .A(\u_a23_core/u_execute/u_register_bank/r6[26] ), 
        .Z(n14745) );
  AND U17403 ( .A(n14747), .B(n14748), .Z(n14743) );
  NANDN U17404 ( .B(n14375), .A(\u_a23_core/u_execute/u_register_bank/r5[26] ), 
        .Z(n14748) );
  NANDN U17405 ( .B(n14376), .A(\u_a23_core/u_execute/u_register_bank/r4[26] ), 
        .Z(n14747) );
  AND U17406 ( .A(n14749), .B(n14750), .Z(n14741) );
  AND U17407 ( .A(n14751), .B(n14752), .Z(n14750) );
  NANDN U17408 ( .B(n14381), .A(\u_a23_core/u_execute/u_register_bank/r3[26] ), 
        .Z(n14752) );
  NANDN U17409 ( .B(n14382), .A(\u_a23_core/u_execute/u_register_bank/r0[26] ), 
        .Z(n14751) );
  AND U17410 ( .A(n14753), .B(n14754), .Z(n14749) );
  NANDN U17411 ( .B(n14385), .A(\u_a23_core/u_execute/u_register_bank/r2[26] ), 
        .Z(n14754) );
  NANDN U17412 ( .B(n14386), .A(\u_a23_core/u_execute/u_register_bank/r1[26] ), 
        .Z(n14753) );
  NANDN U17413 ( .B(n14387), .A(\u_a23_core/read_data_s2[26] ), .Z(n14724) );
  NAND U17414 ( .A(n14255), .B(n14718), .Z(n8525) );
  ANDN U17415 ( .A(n6988), .B(n14225), .Z(n14255) );
  NANDN U17416 ( .B(n8533), .A(n6827), .Z(n14720) );
  NAND U17417 ( .A(n14755), .B(n14756), .Z(n6827) );
  NAND U17418 ( .A(n6778), .B(\u_a23_core/imm32[25] ), .Z(n14756) );
  AND U17419 ( .A(n14757), .B(n14758), .Z(n14755) );
  NANDN U17420 ( .B(n6600), .A(\u_a23_core/barrel_shift_data_sel[1] ), .Z(
        n14758) );
  AND U17421 ( .A(n14759), .B(n14760), .Z(n6600) );
  AND U17422 ( .A(n14761), .B(n14762), .Z(n14760) );
  AND U17423 ( .A(n14763), .B(n14764), .Z(n14762) );
  AND U17424 ( .A(n14765), .B(n14766), .Z(n14764) );
  NAND U17425 ( .A(n14349), .B(\u_a23_core/u_execute/pc[25] ), .Z(n14766) );
  NANDN U17426 ( .B(n14350), .A(\u_a23_core/u_execute/u_register_bank/r14[25] ), .Z(n14765) );
  AND U17427 ( .A(n14767), .B(n14768), .Z(n14763) );
  NANDN U17428 ( .B(n14353), .A(\u_a23_core/u_execute/u_register_bank/r13[25] ), .Z(n14768) );
  NANDN U17429 ( .B(n14354), .A(\u_a23_core/u_execute/u_register_bank/r12[25] ), .Z(n14767) );
  AND U17430 ( .A(n14769), .B(n14770), .Z(n14761) );
  AND U17431 ( .A(n14771), .B(n14772), .Z(n14770) );
  NANDN U17432 ( .B(n14359), .A(\u_a23_core/u_execute/u_register_bank/r11[25] ), .Z(n14772) );
  NANDN U17433 ( .B(n14360), .A(\u_a23_core/u_execute/u_register_bank/r10[25] ), .Z(n14771) );
  AND U17434 ( .A(n14773), .B(n14774), .Z(n14769) );
  NANDN U17435 ( .B(n14363), .A(\u_a23_core/u_execute/u_register_bank/r9[25] ), 
        .Z(n14774) );
  NANDN U17436 ( .B(n14364), .A(\u_a23_core/u_execute/u_register_bank/r8[25] ), 
        .Z(n14773) );
  AND U17437 ( .A(n14775), .B(n14776), .Z(n14759) );
  AND U17438 ( .A(n14777), .B(n14778), .Z(n14776) );
  AND U17439 ( .A(n14779), .B(n14780), .Z(n14778) );
  NANDN U17440 ( .B(n14371), .A(\u_a23_core/u_execute/u_register_bank/r7[25] ), 
        .Z(n14780) );
  NANDN U17441 ( .B(n14372), .A(\u_a23_core/u_execute/u_register_bank/r6[25] ), 
        .Z(n14779) );
  AND U17442 ( .A(n14781), .B(n14782), .Z(n14777) );
  NANDN U17443 ( .B(n14375), .A(\u_a23_core/u_execute/u_register_bank/r5[25] ), 
        .Z(n14782) );
  NANDN U17444 ( .B(n14376), .A(\u_a23_core/u_execute/u_register_bank/r4[25] ), 
        .Z(n14781) );
  AND U17445 ( .A(n14783), .B(n14784), .Z(n14775) );
  AND U17446 ( .A(n14785), .B(n14786), .Z(n14784) );
  NANDN U17447 ( .B(n14381), .A(\u_a23_core/u_execute/u_register_bank/r3[25] ), 
        .Z(n14786) );
  NANDN U17448 ( .B(n14382), .A(\u_a23_core/u_execute/u_register_bank/r0[25] ), 
        .Z(n14785) );
  AND U17449 ( .A(n14787), .B(n14788), .Z(n14783) );
  NANDN U17450 ( .B(n14385), .A(\u_a23_core/u_execute/u_register_bank/r2[25] ), 
        .Z(n14788) );
  NANDN U17451 ( .B(n14386), .A(\u_a23_core/u_execute/u_register_bank/r1[25] ), 
        .Z(n14787) );
  NANDN U17452 ( .B(n14387), .A(\u_a23_core/read_data_s2[25] ), .Z(n14757) );
  NAND U17453 ( .A(n14718), .B(n14789), .Z(n8533) );
  AND U17454 ( .A(n14790), .B(n14791), .Z(n14643) );
  AND U17455 ( .A(n14792), .B(n14793), .Z(n14791) );
  NANDN U17456 ( .B(n8537), .A(n6833), .Z(n14793) );
  NAND U17457 ( .A(n14794), .B(n14795), .Z(n6833) );
  NAND U17458 ( .A(n6778), .B(\u_a23_core/imm32[24] ), .Z(n14795) );
  AND U17459 ( .A(n14796), .B(n14797), .Z(n14794) );
  NANDN U17460 ( .B(n6593), .A(\u_a23_core/barrel_shift_data_sel[1] ), .Z(
        n14797) );
  AND U17461 ( .A(n14798), .B(n14799), .Z(n6593) );
  AND U17462 ( .A(n14800), .B(n14801), .Z(n14799) );
  AND U17463 ( .A(n14802), .B(n14803), .Z(n14801) );
  AND U17464 ( .A(n14804), .B(n14805), .Z(n14803) );
  NAND U17465 ( .A(n14349), .B(\u_a23_core/u_execute/pc[24] ), .Z(n14805) );
  NANDN U17466 ( .B(n14350), .A(\u_a23_core/u_execute/u_register_bank/r14[24] ), .Z(n14804) );
  AND U17467 ( .A(n14806), .B(n14807), .Z(n14802) );
  NANDN U17468 ( .B(n14353), .A(\u_a23_core/u_execute/u_register_bank/r13[24] ), .Z(n14807) );
  NANDN U17469 ( .B(n14354), .A(\u_a23_core/u_execute/u_register_bank/r12[24] ), .Z(n14806) );
  AND U17470 ( .A(n14808), .B(n14809), .Z(n14800) );
  AND U17471 ( .A(n14810), .B(n14811), .Z(n14809) );
  NANDN U17472 ( .B(n14359), .A(\u_a23_core/u_execute/u_register_bank/r11[24] ), .Z(n14811) );
  NANDN U17473 ( .B(n14360), .A(\u_a23_core/u_execute/u_register_bank/r10[24] ), .Z(n14810) );
  AND U17474 ( .A(n14812), .B(n14813), .Z(n14808) );
  NANDN U17475 ( .B(n14363), .A(\u_a23_core/u_execute/u_register_bank/r9[24] ), 
        .Z(n14813) );
  NANDN U17476 ( .B(n14364), .A(\u_a23_core/u_execute/u_register_bank/r8[24] ), 
        .Z(n14812) );
  AND U17477 ( .A(n14814), .B(n14815), .Z(n14798) );
  AND U17478 ( .A(n14816), .B(n14817), .Z(n14815) );
  AND U17479 ( .A(n14818), .B(n14819), .Z(n14817) );
  NANDN U17480 ( .B(n14371), .A(\u_a23_core/u_execute/u_register_bank/r7[24] ), 
        .Z(n14819) );
  NANDN U17481 ( .B(n14372), .A(\u_a23_core/u_execute/u_register_bank/r6[24] ), 
        .Z(n14818) );
  AND U17482 ( .A(n14820), .B(n14821), .Z(n14816) );
  NANDN U17483 ( .B(n14375), .A(\u_a23_core/u_execute/u_register_bank/r5[24] ), 
        .Z(n14821) );
  NANDN U17484 ( .B(n14376), .A(\u_a23_core/u_execute/u_register_bank/r4[24] ), 
        .Z(n14820) );
  AND U17485 ( .A(n14822), .B(n14823), .Z(n14814) );
  AND U17486 ( .A(n14824), .B(n14825), .Z(n14823) );
  NANDN U17487 ( .B(n14381), .A(\u_a23_core/u_execute/u_register_bank/r3[24] ), 
        .Z(n14825) );
  NANDN U17488 ( .B(n14382), .A(\u_a23_core/u_execute/u_register_bank/r0[24] ), 
        .Z(n14824) );
  AND U17489 ( .A(n14826), .B(n14827), .Z(n14822) );
  NANDN U17490 ( .B(n14385), .A(\u_a23_core/u_execute/u_register_bank/r2[24] ), 
        .Z(n14827) );
  NANDN U17491 ( .B(n14386), .A(\u_a23_core/u_execute/u_register_bank/r1[24] ), 
        .Z(n14826) );
  NANDN U17492 ( .B(n14387), .A(\u_a23_core/read_data_s2[24] ), .Z(n14796) );
  NAND U17493 ( .A(n14828), .B(n14718), .Z(n8537) );
  ANDN U17494 ( .A(n14829), .B(n14830), .Z(n14718) );
  OR U17495 ( .A(n14717), .B(n14305), .Z(n14829) );
  NANDN U17496 ( .B(n8538), .A(n6835), .Z(n14792) );
  NAND U17497 ( .A(n14831), .B(n14832), .Z(n6835) );
  NAND U17498 ( .A(n6778), .B(\u_a23_core/imm32[23] ), .Z(n14832) );
  AND U17499 ( .A(n14833), .B(n14834), .Z(n14831) );
  NANDN U17500 ( .B(n6586), .A(\u_a23_core/barrel_shift_data_sel[1] ), .Z(
        n14834) );
  AND U17501 ( .A(n14835), .B(n14836), .Z(n6586) );
  AND U17502 ( .A(n14837), .B(n14838), .Z(n14836) );
  AND U17503 ( .A(n14839), .B(n14840), .Z(n14838) );
  AND U17504 ( .A(n14841), .B(n14842), .Z(n14840) );
  NAND U17505 ( .A(n14349), .B(\u_a23_core/u_execute/pc[23] ), .Z(n14842) );
  NANDN U17506 ( .B(n14350), .A(\u_a23_core/u_execute/u_register_bank/r14[23] ), .Z(n14841) );
  AND U17507 ( .A(n14843), .B(n14844), .Z(n14839) );
  NANDN U17508 ( .B(n14353), .A(\u_a23_core/u_execute/u_register_bank/r13[23] ), .Z(n14844) );
  NANDN U17509 ( .B(n14354), .A(\u_a23_core/u_execute/u_register_bank/r12[23] ), .Z(n14843) );
  AND U17510 ( .A(n14845), .B(n14846), .Z(n14837) );
  AND U17511 ( .A(n14847), .B(n14848), .Z(n14846) );
  NANDN U17512 ( .B(n14359), .A(\u_a23_core/u_execute/u_register_bank/r11[23] ), .Z(n14848) );
  NANDN U17513 ( .B(n14360), .A(\u_a23_core/u_execute/u_register_bank/r10[23] ), .Z(n14847) );
  AND U17514 ( .A(n14849), .B(n14850), .Z(n14845) );
  NANDN U17515 ( .B(n14363), .A(\u_a23_core/u_execute/u_register_bank/r9[23] ), 
        .Z(n14850) );
  NANDN U17516 ( .B(n14364), .A(\u_a23_core/u_execute/u_register_bank/r8[23] ), 
        .Z(n14849) );
  AND U17517 ( .A(n14851), .B(n14852), .Z(n14835) );
  AND U17518 ( .A(n14853), .B(n14854), .Z(n14852) );
  AND U17519 ( .A(n14855), .B(n14856), .Z(n14854) );
  NANDN U17520 ( .B(n14371), .A(\u_a23_core/u_execute/u_register_bank/r7[23] ), 
        .Z(n14856) );
  NANDN U17521 ( .B(n14372), .A(\u_a23_core/u_execute/u_register_bank/r6[23] ), 
        .Z(n14855) );
  AND U17522 ( .A(n14857), .B(n14858), .Z(n14853) );
  NANDN U17523 ( .B(n14375), .A(\u_a23_core/u_execute/u_register_bank/r5[23] ), 
        .Z(n14858) );
  NANDN U17524 ( .B(n14376), .A(\u_a23_core/u_execute/u_register_bank/r4[23] ), 
        .Z(n14857) );
  AND U17525 ( .A(n14859), .B(n14860), .Z(n14851) );
  AND U17526 ( .A(n14861), .B(n14862), .Z(n14860) );
  NANDN U17527 ( .B(n14381), .A(\u_a23_core/u_execute/u_register_bank/r3[23] ), 
        .Z(n14862) );
  NANDN U17528 ( .B(n14382), .A(\u_a23_core/u_execute/u_register_bank/r0[23] ), 
        .Z(n14861) );
  AND U17529 ( .A(n14863), .B(n14864), .Z(n14859) );
  NANDN U17530 ( .B(n14385), .A(\u_a23_core/u_execute/u_register_bank/r2[23] ), 
        .Z(n14864) );
  NANDN U17531 ( .B(n14386), .A(\u_a23_core/u_execute/u_register_bank/r1[23] ), 
        .Z(n14863) );
  NANDN U17532 ( .B(n14387), .A(\u_a23_core/read_data_s2[23] ), .Z(n14833) );
  NAND U17533 ( .A(n14865), .B(n14789), .Z(n8538) );
  AND U17534 ( .A(n14866), .B(n14867), .Z(n14790) );
  NANDN U17535 ( .B(n8543), .A(n6839), .Z(n14867) );
  NAND U17536 ( .A(n14868), .B(n14869), .Z(n6839) );
  NAND U17537 ( .A(n6778), .B(\u_a23_core/imm32[22] ), .Z(n14869) );
  AND U17538 ( .A(n14870), .B(n14871), .Z(n14868) );
  NANDN U17539 ( .B(n6579), .A(\u_a23_core/barrel_shift_data_sel[1] ), .Z(
        n14871) );
  AND U17540 ( .A(n14872), .B(n14873), .Z(n6579) );
  AND U17541 ( .A(n14874), .B(n14875), .Z(n14873) );
  AND U17542 ( .A(n14876), .B(n14877), .Z(n14875) );
  AND U17543 ( .A(n14878), .B(n14879), .Z(n14877) );
  NAND U17544 ( .A(n14349), .B(\u_a23_core/u_execute/pc[22] ), .Z(n14879) );
  NANDN U17545 ( .B(n14350), .A(\u_a23_core/u_execute/u_register_bank/r14[22] ), .Z(n14878) );
  AND U17546 ( .A(n14880), .B(n14881), .Z(n14876) );
  NANDN U17547 ( .B(n14353), .A(\u_a23_core/u_execute/u_register_bank/r13[22] ), .Z(n14881) );
  NANDN U17548 ( .B(n14354), .A(\u_a23_core/u_execute/u_register_bank/r12[22] ), .Z(n14880) );
  AND U17549 ( .A(n14882), .B(n14883), .Z(n14874) );
  AND U17550 ( .A(n14884), .B(n14885), .Z(n14883) );
  NANDN U17551 ( .B(n14359), .A(\u_a23_core/u_execute/u_register_bank/r11[22] ), .Z(n14885) );
  NANDN U17552 ( .B(n14360), .A(\u_a23_core/u_execute/u_register_bank/r10[22] ), .Z(n14884) );
  AND U17553 ( .A(n14886), .B(n14887), .Z(n14882) );
  NANDN U17554 ( .B(n14363), .A(\u_a23_core/u_execute/u_register_bank/r9[22] ), 
        .Z(n14887) );
  NANDN U17555 ( .B(n14364), .A(\u_a23_core/u_execute/u_register_bank/r8[22] ), 
        .Z(n14886) );
  AND U17556 ( .A(n14888), .B(n14889), .Z(n14872) );
  AND U17557 ( .A(n14890), .B(n14891), .Z(n14889) );
  AND U17558 ( .A(n14892), .B(n14893), .Z(n14891) );
  NANDN U17559 ( .B(n14371), .A(\u_a23_core/u_execute/u_register_bank/r7[22] ), 
        .Z(n14893) );
  NANDN U17560 ( .B(n14372), .A(\u_a23_core/u_execute/u_register_bank/r6[22] ), 
        .Z(n14892) );
  AND U17561 ( .A(n14894), .B(n14895), .Z(n14890) );
  NANDN U17562 ( .B(n14375), .A(\u_a23_core/u_execute/u_register_bank/r5[22] ), 
        .Z(n14895) );
  NANDN U17563 ( .B(n14376), .A(\u_a23_core/u_execute/u_register_bank/r4[22] ), 
        .Z(n14894) );
  AND U17564 ( .A(n14896), .B(n14897), .Z(n14888) );
  AND U17565 ( .A(n14898), .B(n14899), .Z(n14897) );
  NANDN U17566 ( .B(n14381), .A(\u_a23_core/u_execute/u_register_bank/r3[22] ), 
        .Z(n14899) );
  NANDN U17567 ( .B(n14382), .A(\u_a23_core/u_execute/u_register_bank/r0[22] ), 
        .Z(n14898) );
  AND U17568 ( .A(n14900), .B(n14901), .Z(n14896) );
  NANDN U17569 ( .B(n14385), .A(\u_a23_core/u_execute/u_register_bank/r2[22] ), 
        .Z(n14901) );
  NANDN U17570 ( .B(n14386), .A(\u_a23_core/u_execute/u_register_bank/r1[22] ), 
        .Z(n14900) );
  NANDN U17571 ( .B(n14387), .A(\u_a23_core/read_data_s2[22] ), .Z(n14870) );
  NAND U17572 ( .A(n14828), .B(n14865), .Z(n8543) );
  AND U17573 ( .A(n14902), .B(n14205), .Z(n14865) );
  IV U17574 ( .A(n14830), .Z(n14902) );
  NAND U17575 ( .A(n14903), .B(n14904), .Z(n14830) );
  OR U17576 ( .A(n14717), .B(n14324), .Z(n14903) );
  NANDN U17577 ( .B(n8544), .A(n6850), .Z(n14866) );
  NAND U17578 ( .A(n14905), .B(n14906), .Z(n6850) );
  NAND U17579 ( .A(n6778), .B(\u_a23_core/imm32[21] ), .Z(n14906) );
  AND U17580 ( .A(n14907), .B(n14908), .Z(n14905) );
  NANDN U17581 ( .B(n6572), .A(\u_a23_core/barrel_shift_data_sel[1] ), .Z(
        n14908) );
  AND U17582 ( .A(n14909), .B(n14910), .Z(n6572) );
  AND U17583 ( .A(n14911), .B(n14912), .Z(n14910) );
  AND U17584 ( .A(n14913), .B(n14914), .Z(n14912) );
  AND U17585 ( .A(n14915), .B(n14916), .Z(n14914) );
  NAND U17586 ( .A(n14349), .B(\u_a23_core/u_execute/pc[21] ), .Z(n14916) );
  NANDN U17587 ( .B(n14350), .A(\u_a23_core/u_execute/u_register_bank/r14[21] ), .Z(n14915) );
  AND U17588 ( .A(n14917), .B(n14918), .Z(n14913) );
  NANDN U17589 ( .B(n14353), .A(\u_a23_core/u_execute/u_register_bank/r13[21] ), .Z(n14918) );
  NANDN U17590 ( .B(n14354), .A(\u_a23_core/u_execute/u_register_bank/r12[21] ), .Z(n14917) );
  AND U17591 ( .A(n14919), .B(n14920), .Z(n14911) );
  AND U17592 ( .A(n14921), .B(n14922), .Z(n14920) );
  NANDN U17593 ( .B(n14359), .A(\u_a23_core/u_execute/u_register_bank/r11[21] ), .Z(n14922) );
  NANDN U17594 ( .B(n14360), .A(\u_a23_core/u_execute/u_register_bank/r10[21] ), .Z(n14921) );
  AND U17595 ( .A(n14923), .B(n14924), .Z(n14919) );
  NANDN U17596 ( .B(n14363), .A(\u_a23_core/u_execute/u_register_bank/r9[21] ), 
        .Z(n14924) );
  NANDN U17597 ( .B(n14364), .A(\u_a23_core/u_execute/u_register_bank/r8[21] ), 
        .Z(n14923) );
  AND U17598 ( .A(n14925), .B(n14926), .Z(n14909) );
  AND U17599 ( .A(n14927), .B(n14928), .Z(n14926) );
  AND U17600 ( .A(n14929), .B(n14930), .Z(n14928) );
  NANDN U17601 ( .B(n14371), .A(\u_a23_core/u_execute/u_register_bank/r7[21] ), 
        .Z(n14930) );
  NANDN U17602 ( .B(n14372), .A(\u_a23_core/u_execute/u_register_bank/r6[21] ), 
        .Z(n14929) );
  AND U17603 ( .A(n14931), .B(n14932), .Z(n14927) );
  NANDN U17604 ( .B(n14375), .A(\u_a23_core/u_execute/u_register_bank/r5[21] ), 
        .Z(n14932) );
  NANDN U17605 ( .B(n14376), .A(\u_a23_core/u_execute/u_register_bank/r4[21] ), 
        .Z(n14931) );
  AND U17606 ( .A(n14933), .B(n14934), .Z(n14925) );
  AND U17607 ( .A(n14935), .B(n14936), .Z(n14934) );
  NANDN U17608 ( .B(n14381), .A(\u_a23_core/u_execute/u_register_bank/r3[21] ), 
        .Z(n14936) );
  NANDN U17609 ( .B(n14382), .A(\u_a23_core/u_execute/u_register_bank/r0[21] ), 
        .Z(n14935) );
  AND U17610 ( .A(n14937), .B(n14938), .Z(n14933) );
  NANDN U17611 ( .B(n14385), .A(\u_a23_core/u_execute/u_register_bank/r2[21] ), 
        .Z(n14938) );
  NANDN U17612 ( .B(n14386), .A(\u_a23_core/u_execute/u_register_bank/r1[21] ), 
        .Z(n14937) );
  NANDN U17613 ( .B(n14387), .A(\u_a23_core/read_data_s2[21] ), .Z(n14907) );
  NAND U17614 ( .A(n14939), .B(n14789), .Z(n8544) );
  AND U17615 ( .A(n14940), .B(n14941), .Z(n14327) );
  AND U17616 ( .A(n14942), .B(n14943), .Z(n14941) );
  AND U17617 ( .A(n14944), .B(n14945), .Z(n14943) );
  AND U17618 ( .A(n14946), .B(n14947), .Z(n14945) );
  NANDN U17619 ( .B(n8547), .A(n6853), .Z(n14947) );
  NAND U17620 ( .A(n14948), .B(n14949), .Z(n6853) );
  NAND U17621 ( .A(n6778), .B(\u_a23_core/imm32[20] ), .Z(n14949) );
  AND U17622 ( .A(n14950), .B(n14951), .Z(n14948) );
  NANDN U17623 ( .B(n6565), .A(\u_a23_core/barrel_shift_data_sel[1] ), .Z(
        n14951) );
  AND U17624 ( .A(n14952), .B(n14953), .Z(n6565) );
  AND U17625 ( .A(n14954), .B(n14955), .Z(n14953) );
  AND U17626 ( .A(n14956), .B(n14957), .Z(n14955) );
  AND U17627 ( .A(n14958), .B(n14959), .Z(n14957) );
  NAND U17628 ( .A(n14349), .B(\u_a23_core/u_execute/pc[20] ), .Z(n14959) );
  NANDN U17629 ( .B(n14350), .A(\u_a23_core/u_execute/u_register_bank/r14[20] ), .Z(n14958) );
  AND U17630 ( .A(n14960), .B(n14961), .Z(n14956) );
  NANDN U17631 ( .B(n14353), .A(\u_a23_core/u_execute/u_register_bank/r13[20] ), .Z(n14961) );
  NANDN U17632 ( .B(n14354), .A(\u_a23_core/u_execute/u_register_bank/r12[20] ), .Z(n14960) );
  AND U17633 ( .A(n14962), .B(n14963), .Z(n14954) );
  AND U17634 ( .A(n14964), .B(n14965), .Z(n14963) );
  NANDN U17635 ( .B(n14359), .A(\u_a23_core/u_execute/u_register_bank/r11[20] ), .Z(n14965) );
  NANDN U17636 ( .B(n14360), .A(\u_a23_core/u_execute/u_register_bank/r10[20] ), .Z(n14964) );
  AND U17637 ( .A(n14966), .B(n14967), .Z(n14962) );
  NANDN U17638 ( .B(n14363), .A(\u_a23_core/u_execute/u_register_bank/r9[20] ), 
        .Z(n14967) );
  NANDN U17639 ( .B(n14364), .A(\u_a23_core/u_execute/u_register_bank/r8[20] ), 
        .Z(n14966) );
  AND U17640 ( .A(n14968), .B(n14969), .Z(n14952) );
  AND U17641 ( .A(n14970), .B(n14971), .Z(n14969) );
  AND U17642 ( .A(n14972), .B(n14973), .Z(n14971) );
  NANDN U17643 ( .B(n14371), .A(\u_a23_core/u_execute/u_register_bank/r7[20] ), 
        .Z(n14973) );
  NANDN U17644 ( .B(n14372), .A(\u_a23_core/u_execute/u_register_bank/r6[20] ), 
        .Z(n14972) );
  AND U17645 ( .A(n14974), .B(n14975), .Z(n14970) );
  NANDN U17646 ( .B(n14375), .A(\u_a23_core/u_execute/u_register_bank/r5[20] ), 
        .Z(n14975) );
  NANDN U17647 ( .B(n14376), .A(\u_a23_core/u_execute/u_register_bank/r4[20] ), 
        .Z(n14974) );
  AND U17648 ( .A(n14976), .B(n14977), .Z(n14968) );
  AND U17649 ( .A(n14978), .B(n14979), .Z(n14977) );
  NANDN U17650 ( .B(n14381), .A(\u_a23_core/u_execute/u_register_bank/r3[20] ), 
        .Z(n14979) );
  NANDN U17651 ( .B(n14382), .A(\u_a23_core/u_execute/u_register_bank/r0[20] ), 
        .Z(n14978) );
  AND U17652 ( .A(n14980), .B(n14981), .Z(n14976) );
  NANDN U17653 ( .B(n14385), .A(\u_a23_core/u_execute/u_register_bank/r2[20] ), 
        .Z(n14981) );
  NANDN U17654 ( .B(n14386), .A(\u_a23_core/u_execute/u_register_bank/r1[20] ), 
        .Z(n14980) );
  NANDN U17655 ( .B(n14387), .A(\u_a23_core/read_data_s2[20] ), .Z(n14950) );
  NAND U17656 ( .A(n14828), .B(n14939), .Z(n8547) );
  AND U17657 ( .A(n14904), .B(n14237), .Z(n14939) );
  ANDN U17658 ( .A(n14982), .B(n14983), .Z(n14904) );
  AND U17659 ( .A(n14984), .B(n14985), .Z(n14982) );
  OR U17660 ( .A(n14717), .B(n14390), .Z(n14985) );
  ANDN U17661 ( .A(n14986), .B(n14789), .Z(n14717) );
  IV U17662 ( .A(n14828), .Z(n14986) );
  NANDN U17663 ( .B(n8548), .A(n6841), .Z(n14946) );
  NAND U17664 ( .A(n14987), .B(n14988), .Z(n6841) );
  NAND U17665 ( .A(n6778), .B(\u_a23_core/imm32[19] ), .Z(n14988) );
  AND U17666 ( .A(n14989), .B(n14990), .Z(n14987) );
  NANDN U17667 ( .B(n6558), .A(\u_a23_core/barrel_shift_data_sel[1] ), .Z(
        n14990) );
  AND U17668 ( .A(n14991), .B(n14992), .Z(n6558) );
  AND U17669 ( .A(n14993), .B(n14994), .Z(n14992) );
  AND U17670 ( .A(n14995), .B(n14996), .Z(n14994) );
  AND U17671 ( .A(n14997), .B(n14998), .Z(n14996) );
  NAND U17672 ( .A(n14349), .B(\u_a23_core/u_execute/pc[19] ), .Z(n14998) );
  NANDN U17673 ( .B(n14350), .A(\u_a23_core/u_execute/u_register_bank/r14[19] ), .Z(n14997) );
  AND U17674 ( .A(n14999), .B(n15000), .Z(n14995) );
  NANDN U17675 ( .B(n14353), .A(\u_a23_core/u_execute/u_register_bank/r13[19] ), .Z(n15000) );
  NANDN U17676 ( .B(n14354), .A(\u_a23_core/u_execute/u_register_bank/r12[19] ), .Z(n14999) );
  AND U17677 ( .A(n15001), .B(n15002), .Z(n14993) );
  AND U17678 ( .A(n15003), .B(n15004), .Z(n15002) );
  NANDN U17679 ( .B(n14359), .A(\u_a23_core/u_execute/u_register_bank/r11[19] ), .Z(n15004) );
  NANDN U17680 ( .B(n14360), .A(\u_a23_core/u_execute/u_register_bank/r10[19] ), .Z(n15003) );
  AND U17681 ( .A(n15005), .B(n15006), .Z(n15001) );
  NANDN U17682 ( .B(n14363), .A(\u_a23_core/u_execute/u_register_bank/r9[19] ), 
        .Z(n15006) );
  NANDN U17683 ( .B(n14364), .A(\u_a23_core/u_execute/u_register_bank/r8[19] ), 
        .Z(n15005) );
  AND U17684 ( .A(n15007), .B(n15008), .Z(n14991) );
  AND U17685 ( .A(n15009), .B(n15010), .Z(n15008) );
  AND U17686 ( .A(n15011), .B(n15012), .Z(n15010) );
  NANDN U17687 ( .B(n14371), .A(\u_a23_core/u_execute/u_register_bank/r7[19] ), 
        .Z(n15012) );
  NANDN U17688 ( .B(n14372), .A(\u_a23_core/u_execute/u_register_bank/r6[19] ), 
        .Z(n15011) );
  AND U17689 ( .A(n15013), .B(n15014), .Z(n15009) );
  NANDN U17690 ( .B(n14375), .A(\u_a23_core/u_execute/u_register_bank/r5[19] ), 
        .Z(n15014) );
  NANDN U17691 ( .B(n14376), .A(\u_a23_core/u_execute/u_register_bank/r4[19] ), 
        .Z(n15013) );
  AND U17692 ( .A(n15015), .B(n15016), .Z(n15007) );
  AND U17693 ( .A(n15017), .B(n15018), .Z(n15016) );
  NANDN U17694 ( .B(n14381), .A(\u_a23_core/u_execute/u_register_bank/r3[19] ), 
        .Z(n15018) );
  NANDN U17695 ( .B(n14382), .A(\u_a23_core/u_execute/u_register_bank/r0[19] ), 
        .Z(n15017) );
  AND U17696 ( .A(n15019), .B(n15020), .Z(n15015) );
  NANDN U17697 ( .B(n14385), .A(\u_a23_core/u_execute/u_register_bank/r2[19] ), 
        .Z(n15020) );
  NANDN U17698 ( .B(n14386), .A(\u_a23_core/u_execute/u_register_bank/r1[19] ), 
        .Z(n15019) );
  NANDN U17699 ( .B(n14387), .A(\u_a23_core/read_data_s2[19] ), .Z(n14989) );
  NAND U17700 ( .A(n15021), .B(n14789), .Z(n8548) );
  ANDN U17701 ( .A(n15022), .B(n14218), .Z(n14789) );
  AND U17702 ( .A(n15023), .B(n15024), .Z(n14944) );
  NANDN U17703 ( .B(n8557), .A(n6857), .Z(n15024) );
  NAND U17704 ( .A(n15025), .B(n15026), .Z(n6857) );
  NAND U17705 ( .A(n6778), .B(\u_a23_core/imm32[18] ), .Z(n15026) );
  AND U17706 ( .A(n15027), .B(n15028), .Z(n15025) );
  NANDN U17707 ( .B(n6551), .A(\u_a23_core/barrel_shift_data_sel[1] ), .Z(
        n15028) );
  AND U17708 ( .A(n15029), .B(n15030), .Z(n6551) );
  AND U17709 ( .A(n15031), .B(n15032), .Z(n15030) );
  AND U17710 ( .A(n15033), .B(n15034), .Z(n15032) );
  AND U17711 ( .A(n15035), .B(n15036), .Z(n15034) );
  NAND U17712 ( .A(n14349), .B(\u_a23_core/u_execute/pc[18] ), .Z(n15036) );
  NANDN U17713 ( .B(n14350), .A(\u_a23_core/u_execute/u_register_bank/r14[18] ), .Z(n15035) );
  AND U17714 ( .A(n15037), .B(n15038), .Z(n15033) );
  NANDN U17715 ( .B(n14353), .A(\u_a23_core/u_execute/u_register_bank/r13[18] ), .Z(n15038) );
  NANDN U17716 ( .B(n14354), .A(\u_a23_core/u_execute/u_register_bank/r12[18] ), .Z(n15037) );
  AND U17717 ( .A(n15039), .B(n15040), .Z(n15031) );
  AND U17718 ( .A(n15041), .B(n15042), .Z(n15040) );
  NANDN U17719 ( .B(n14359), .A(\u_a23_core/u_execute/u_register_bank/r11[18] ), .Z(n15042) );
  NANDN U17720 ( .B(n14360), .A(\u_a23_core/u_execute/u_register_bank/r10[18] ), .Z(n15041) );
  AND U17721 ( .A(n15043), .B(n15044), .Z(n15039) );
  NANDN U17722 ( .B(n14363), .A(\u_a23_core/u_execute/u_register_bank/r9[18] ), 
        .Z(n15044) );
  NANDN U17723 ( .B(n14364), .A(\u_a23_core/u_execute/u_register_bank/r8[18] ), 
        .Z(n15043) );
  AND U17724 ( .A(n15045), .B(n15046), .Z(n15029) );
  AND U17725 ( .A(n15047), .B(n15048), .Z(n15046) );
  AND U17726 ( .A(n15049), .B(n15050), .Z(n15048) );
  NANDN U17727 ( .B(n14371), .A(\u_a23_core/u_execute/u_register_bank/r7[18] ), 
        .Z(n15050) );
  NANDN U17728 ( .B(n14372), .A(\u_a23_core/u_execute/u_register_bank/r6[18] ), 
        .Z(n15049) );
  AND U17729 ( .A(n15051), .B(n15052), .Z(n15047) );
  NANDN U17730 ( .B(n14375), .A(\u_a23_core/u_execute/u_register_bank/r5[18] ), 
        .Z(n15052) );
  NANDN U17731 ( .B(n14376), .A(\u_a23_core/u_execute/u_register_bank/r4[18] ), 
        .Z(n15051) );
  AND U17732 ( .A(n15053), .B(n15054), .Z(n15045) );
  AND U17733 ( .A(n15055), .B(n15056), .Z(n15054) );
  NANDN U17734 ( .B(n14381), .A(\u_a23_core/u_execute/u_register_bank/r3[18] ), 
        .Z(n15056) );
  NANDN U17735 ( .B(n14382), .A(\u_a23_core/u_execute/u_register_bank/r0[18] ), 
        .Z(n15055) );
  AND U17736 ( .A(n15057), .B(n15058), .Z(n15053) );
  NANDN U17737 ( .B(n14385), .A(\u_a23_core/u_execute/u_register_bank/r2[18] ), 
        .Z(n15058) );
  NANDN U17738 ( .B(n14386), .A(\u_a23_core/u_execute/u_register_bank/r1[18] ), 
        .Z(n15057) );
  NANDN U17739 ( .B(n14387), .A(\u_a23_core/read_data_s2[18] ), .Z(n15027) );
  NAND U17740 ( .A(n14828), .B(n15021), .Z(n8557) );
  ANDN U17741 ( .A(n14984), .B(n14390), .Z(n15021) );
  NOR U17742 ( .A(n14295), .B(n14225), .Z(n14828) );
  NANDN U17743 ( .B(n8558), .A(n6859), .Z(n15023) );
  NAND U17744 ( .A(n15059), .B(n15060), .Z(n6859) );
  NAND U17745 ( .A(n6778), .B(\u_a23_core/imm32[17] ), .Z(n15060) );
  AND U17746 ( .A(n15061), .B(n15062), .Z(n15059) );
  NANDN U17747 ( .B(n6544), .A(\u_a23_core/barrel_shift_data_sel[1] ), .Z(
        n15062) );
  AND U17748 ( .A(n15063), .B(n15064), .Z(n6544) );
  AND U17749 ( .A(n15065), .B(n15066), .Z(n15064) );
  AND U17750 ( .A(n15067), .B(n15068), .Z(n15066) );
  AND U17751 ( .A(n15069), .B(n15070), .Z(n15068) );
  NAND U17752 ( .A(n14349), .B(\u_a23_core/u_execute/pc[17] ), .Z(n15070) );
  NANDN U17753 ( .B(n14350), .A(\u_a23_core/u_execute/u_register_bank/r14[17] ), .Z(n15069) );
  AND U17754 ( .A(n15071), .B(n15072), .Z(n15067) );
  NANDN U17755 ( .B(n14353), .A(\u_a23_core/u_execute/u_register_bank/r13[17] ), .Z(n15072) );
  NANDN U17756 ( .B(n14354), .A(\u_a23_core/u_execute/u_register_bank/r12[17] ), .Z(n15071) );
  AND U17757 ( .A(n15073), .B(n15074), .Z(n15065) );
  AND U17758 ( .A(n15075), .B(n15076), .Z(n15074) );
  NANDN U17759 ( .B(n14359), .A(\u_a23_core/u_execute/u_register_bank/r11[17] ), .Z(n15076) );
  NANDN U17760 ( .B(n14360), .A(\u_a23_core/u_execute/u_register_bank/r10[17] ), .Z(n15075) );
  AND U17761 ( .A(n15077), .B(n15078), .Z(n15073) );
  NANDN U17762 ( .B(n14363), .A(\u_a23_core/u_execute/u_register_bank/r9[17] ), 
        .Z(n15078) );
  NANDN U17763 ( .B(n14364), .A(\u_a23_core/u_execute/u_register_bank/r8[17] ), 
        .Z(n15077) );
  AND U17764 ( .A(n15079), .B(n15080), .Z(n15063) );
  AND U17765 ( .A(n15081), .B(n15082), .Z(n15080) );
  AND U17766 ( .A(n15083), .B(n15084), .Z(n15082) );
  NANDN U17767 ( .B(n14371), .A(\u_a23_core/u_execute/u_register_bank/r7[17] ), 
        .Z(n15084) );
  NANDN U17768 ( .B(n14372), .A(\u_a23_core/u_execute/u_register_bank/r6[17] ), 
        .Z(n15083) );
  AND U17769 ( .A(n15085), .B(n15086), .Z(n15081) );
  NANDN U17770 ( .B(n14375), .A(\u_a23_core/u_execute/u_register_bank/r5[17] ), 
        .Z(n15086) );
  NANDN U17771 ( .B(n14376), .A(\u_a23_core/u_execute/u_register_bank/r4[17] ), 
        .Z(n15085) );
  AND U17772 ( .A(n15087), .B(n15088), .Z(n15079) );
  AND U17773 ( .A(n15089), .B(n15090), .Z(n15088) );
  NANDN U17774 ( .B(n14381), .A(\u_a23_core/u_execute/u_register_bank/r3[17] ), 
        .Z(n15090) );
  NANDN U17775 ( .B(n14382), .A(\u_a23_core/u_execute/u_register_bank/r0[17] ), 
        .Z(n15089) );
  AND U17776 ( .A(n15091), .B(n15092), .Z(n15087) );
  NANDN U17777 ( .B(n14385), .A(\u_a23_core/u_execute/u_register_bank/r2[17] ), 
        .Z(n15092) );
  NANDN U17778 ( .B(n14386), .A(\u_a23_core/u_execute/u_register_bank/r1[17] ), 
        .Z(n15091) );
  NANDN U17779 ( .B(n14387), .A(\u_a23_core/read_data_s2[17] ), .Z(n15061) );
  NAND U17780 ( .A(n15093), .B(n14984), .Z(n8558) );
  AND U17781 ( .A(n15094), .B(n15095), .Z(n14942) );
  AND U17782 ( .A(n15096), .B(n15097), .Z(n15095) );
  NANDN U17783 ( .B(n8561), .A(n6865), .Z(n15097) );
  NAND U17784 ( .A(n15098), .B(n15099), .Z(n6865) );
  NAND U17785 ( .A(n6778), .B(\u_a23_core/imm32[16] ), .Z(n15099) );
  AND U17786 ( .A(n15100), .B(n15101), .Z(n15098) );
  NANDN U17787 ( .B(n6537), .A(\u_a23_core/barrel_shift_data_sel[1] ), .Z(
        n15101) );
  AND U17788 ( .A(n15102), .B(n15103), .Z(n6537) );
  AND U17789 ( .A(n15104), .B(n15105), .Z(n15103) );
  AND U17790 ( .A(n15106), .B(n15107), .Z(n15105) );
  AND U17791 ( .A(n15108), .B(n15109), .Z(n15107) );
  NAND U17792 ( .A(n14349), .B(\u_a23_core/u_execute/pc[16] ), .Z(n15109) );
  NANDN U17793 ( .B(n14350), .A(\u_a23_core/u_execute/u_register_bank/r14[16] ), .Z(n15108) );
  AND U17794 ( .A(n15110), .B(n15111), .Z(n15106) );
  NANDN U17795 ( .B(n14353), .A(\u_a23_core/u_execute/u_register_bank/r13[16] ), .Z(n15111) );
  NANDN U17796 ( .B(n14354), .A(\u_a23_core/u_execute/u_register_bank/r12[16] ), .Z(n15110) );
  AND U17797 ( .A(n15112), .B(n15113), .Z(n15104) );
  AND U17798 ( .A(n15114), .B(n15115), .Z(n15113) );
  NANDN U17799 ( .B(n14359), .A(\u_a23_core/u_execute/u_register_bank/r11[16] ), .Z(n15115) );
  NANDN U17800 ( .B(n14360), .A(\u_a23_core/u_execute/u_register_bank/r10[16] ), .Z(n15114) );
  AND U17801 ( .A(n15116), .B(n15117), .Z(n15112) );
  NANDN U17802 ( .B(n14363), .A(\u_a23_core/u_execute/u_register_bank/r9[16] ), 
        .Z(n15117) );
  NANDN U17803 ( .B(n14364), .A(\u_a23_core/u_execute/u_register_bank/r8[16] ), 
        .Z(n15116) );
  AND U17804 ( .A(n15118), .B(n15119), .Z(n15102) );
  AND U17805 ( .A(n15120), .B(n15121), .Z(n15119) );
  AND U17806 ( .A(n15122), .B(n15123), .Z(n15121) );
  NANDN U17807 ( .B(n14371), .A(\u_a23_core/u_execute/u_register_bank/r7[16] ), 
        .Z(n15123) );
  NANDN U17808 ( .B(n14372), .A(\u_a23_core/u_execute/u_register_bank/r6[16] ), 
        .Z(n15122) );
  AND U17809 ( .A(n15124), .B(n15125), .Z(n15120) );
  NANDN U17810 ( .B(n14375), .A(\u_a23_core/u_execute/u_register_bank/r5[16] ), 
        .Z(n15125) );
  NANDN U17811 ( .B(n14376), .A(\u_a23_core/u_execute/u_register_bank/r4[16] ), 
        .Z(n15124) );
  AND U17812 ( .A(n15126), .B(n15127), .Z(n15118) );
  AND U17813 ( .A(n15128), .B(n15129), .Z(n15127) );
  NANDN U17814 ( .B(n14381), .A(\u_a23_core/u_execute/u_register_bank/r3[16] ), 
        .Z(n15129) );
  NANDN U17815 ( .B(n14382), .A(\u_a23_core/u_execute/u_register_bank/r0[16] ), 
        .Z(n15128) );
  AND U17816 ( .A(n15130), .B(n15131), .Z(n15126) );
  NANDN U17817 ( .B(n14385), .A(\u_a23_core/u_execute/u_register_bank/r2[16] ), 
        .Z(n15131) );
  NANDN U17818 ( .B(n14386), .A(\u_a23_core/u_execute/u_register_bank/r1[16] ), 
        .Z(n15130) );
  NANDN U17819 ( .B(n14387), .A(\u_a23_core/read_data_s2[16] ), .Z(n15100) );
  NAND U17820 ( .A(n15132), .B(n14984), .Z(n8561) );
  AND U17821 ( .A(n15133), .B(n15134), .Z(n14984) );
  NAND U17822 ( .A(n14205), .B(n14983), .Z(n15133) );
  NANDN U17823 ( .B(n8562), .A(n6967), .Z(n15096) );
  NAND U17824 ( .A(n15135), .B(n15136), .Z(n6967) );
  NAND U17825 ( .A(n6778), .B(\u_a23_core/imm32[15] ), .Z(n15136) );
  AND U17826 ( .A(n15137), .B(n15138), .Z(n15135) );
  NANDN U17827 ( .B(n6530), .A(\u_a23_core/barrel_shift_data_sel[1] ), .Z(
        n15138) );
  AND U17828 ( .A(n15139), .B(n15140), .Z(n6530) );
  AND U17829 ( .A(n15141), .B(n15142), .Z(n15140) );
  AND U17830 ( .A(n15143), .B(n15144), .Z(n15142) );
  AND U17831 ( .A(n15145), .B(n15146), .Z(n15144) );
  NAND U17832 ( .A(n14349), .B(\u_a23_core/u_execute/pc[15] ), .Z(n15146) );
  NANDN U17833 ( .B(n14350), .A(\u_a23_core/u_execute/u_register_bank/r14[15] ), .Z(n15145) );
  AND U17834 ( .A(n15147), .B(n15148), .Z(n15143) );
  NANDN U17835 ( .B(n14353), .A(\u_a23_core/u_execute/u_register_bank/r13[15] ), .Z(n15148) );
  NANDN U17836 ( .B(n14354), .A(\u_a23_core/u_execute/u_register_bank/r12[15] ), .Z(n15147) );
  AND U17837 ( .A(n15149), .B(n15150), .Z(n15141) );
  AND U17838 ( .A(n15151), .B(n15152), .Z(n15150) );
  NANDN U17839 ( .B(n14359), .A(\u_a23_core/u_execute/u_register_bank/r11[15] ), .Z(n15152) );
  NANDN U17840 ( .B(n14360), .A(\u_a23_core/u_execute/u_register_bank/r10[15] ), .Z(n15151) );
  AND U17841 ( .A(n15153), .B(n15154), .Z(n15149) );
  NANDN U17842 ( .B(n14363), .A(\u_a23_core/u_execute/u_register_bank/r9[15] ), 
        .Z(n15154) );
  NANDN U17843 ( .B(n14364), .A(\u_a23_core/u_execute/u_register_bank/r8[15] ), 
        .Z(n15153) );
  AND U17844 ( .A(n15155), .B(n15156), .Z(n15139) );
  AND U17845 ( .A(n15157), .B(n15158), .Z(n15156) );
  AND U17846 ( .A(n15159), .B(n15160), .Z(n15158) );
  NANDN U17847 ( .B(n14371), .A(\u_a23_core/u_execute/u_register_bank/r7[15] ), 
        .Z(n15160) );
  NANDN U17848 ( .B(n14372), .A(\u_a23_core/u_execute/u_register_bank/r6[15] ), 
        .Z(n15159) );
  AND U17849 ( .A(n15161), .B(n15162), .Z(n15157) );
  NANDN U17850 ( .B(n14375), .A(\u_a23_core/u_execute/u_register_bank/r5[15] ), 
        .Z(n15162) );
  NANDN U17851 ( .B(n14376), .A(\u_a23_core/u_execute/u_register_bank/r4[15] ), 
        .Z(n15161) );
  AND U17852 ( .A(n15163), .B(n15164), .Z(n15155) );
  AND U17853 ( .A(n15165), .B(n15166), .Z(n15164) );
  NANDN U17854 ( .B(n14381), .A(\u_a23_core/u_execute/u_register_bank/r3[15] ), 
        .Z(n15166) );
  NANDN U17855 ( .B(n14382), .A(\u_a23_core/u_execute/u_register_bank/r0[15] ), 
        .Z(n15165) );
  AND U17856 ( .A(n15167), .B(n15168), .Z(n15163) );
  NANDN U17857 ( .B(n14385), .A(\u_a23_core/u_execute/u_register_bank/r2[15] ), 
        .Z(n15168) );
  NANDN U17858 ( .B(n14386), .A(\u_a23_core/u_execute/u_register_bank/r1[15] ), 
        .Z(n15167) );
  NANDN U17859 ( .B(n14387), .A(\u_a23_core/read_data_s2[15] ), .Z(n15137) );
  NAND U17860 ( .A(n15169), .B(n15134), .Z(n8562) );
  AND U17861 ( .A(n15093), .B(n14205), .Z(n15169) );
  AND U17862 ( .A(n15170), .B(n15171), .Z(n15094) );
  NANDN U17863 ( .B(n8567), .A(n6966), .Z(n15171) );
  NAND U17864 ( .A(n15172), .B(n15173), .Z(n6966) );
  NAND U17865 ( .A(n6778), .B(\u_a23_core/imm32[14] ), .Z(n15173) );
  AND U17866 ( .A(n15174), .B(n15175), .Z(n15172) );
  NANDN U17867 ( .B(n6523), .A(\u_a23_core/barrel_shift_data_sel[1] ), .Z(
        n15175) );
  AND U17868 ( .A(n15176), .B(n15177), .Z(n6523) );
  AND U17869 ( .A(n15178), .B(n15179), .Z(n15177) );
  AND U17870 ( .A(n15180), .B(n15181), .Z(n15179) );
  AND U17871 ( .A(n15182), .B(n15183), .Z(n15181) );
  NAND U17872 ( .A(n14349), .B(\u_a23_core/u_execute/pc[14] ), .Z(n15183) );
  NANDN U17873 ( .B(n14350), .A(\u_a23_core/u_execute/u_register_bank/r14[14] ), .Z(n15182) );
  AND U17874 ( .A(n15184), .B(n15185), .Z(n15180) );
  NANDN U17875 ( .B(n14353), .A(\u_a23_core/u_execute/u_register_bank/r13[14] ), .Z(n15185) );
  NANDN U17876 ( .B(n14354), .A(\u_a23_core/u_execute/u_register_bank/r12[14] ), .Z(n15184) );
  AND U17877 ( .A(n15186), .B(n15187), .Z(n15178) );
  AND U17878 ( .A(n15188), .B(n15189), .Z(n15187) );
  NANDN U17879 ( .B(n14359), .A(\u_a23_core/u_execute/u_register_bank/r11[14] ), .Z(n15189) );
  NANDN U17880 ( .B(n14360), .A(\u_a23_core/u_execute/u_register_bank/r10[14] ), .Z(n15188) );
  AND U17881 ( .A(n15190), .B(n15191), .Z(n15186) );
  NANDN U17882 ( .B(n14363), .A(\u_a23_core/u_execute/u_register_bank/r9[14] ), 
        .Z(n15191) );
  NANDN U17883 ( .B(n14364), .A(\u_a23_core/u_execute/u_register_bank/r8[14] ), 
        .Z(n15190) );
  AND U17884 ( .A(n15192), .B(n15193), .Z(n15176) );
  AND U17885 ( .A(n15194), .B(n15195), .Z(n15193) );
  AND U17886 ( .A(n15196), .B(n15197), .Z(n15195) );
  NANDN U17887 ( .B(n14371), .A(\u_a23_core/u_execute/u_register_bank/r7[14] ), 
        .Z(n15197) );
  NANDN U17888 ( .B(n14372), .A(\u_a23_core/u_execute/u_register_bank/r6[14] ), 
        .Z(n15196) );
  AND U17889 ( .A(n15198), .B(n15199), .Z(n15194) );
  NANDN U17890 ( .B(n14375), .A(\u_a23_core/u_execute/u_register_bank/r5[14] ), 
        .Z(n15199) );
  NANDN U17891 ( .B(n14376), .A(\u_a23_core/u_execute/u_register_bank/r4[14] ), 
        .Z(n15198) );
  AND U17892 ( .A(n15200), .B(n15201), .Z(n15192) );
  AND U17893 ( .A(n15202), .B(n15203), .Z(n15201) );
  NANDN U17894 ( .B(n14381), .A(\u_a23_core/u_execute/u_register_bank/r3[14] ), 
        .Z(n15203) );
  NANDN U17895 ( .B(n14382), .A(\u_a23_core/u_execute/u_register_bank/r0[14] ), 
        .Z(n15202) );
  AND U17896 ( .A(n15204), .B(n15205), .Z(n15200) );
  NANDN U17897 ( .B(n14385), .A(\u_a23_core/u_execute/u_register_bank/r2[14] ), 
        .Z(n15205) );
  NANDN U17898 ( .B(n14386), .A(\u_a23_core/u_execute/u_register_bank/r1[14] ), 
        .Z(n15204) );
  NANDN U17899 ( .B(n14387), .A(\u_a23_core/read_data_s2[14] ), .Z(n15174) );
  NAND U17900 ( .A(n15206), .B(n15134), .Z(n8567) );
  AND U17901 ( .A(n15207), .B(n15208), .Z(n15134) );
  NAND U17902 ( .A(n14237), .B(n14983), .Z(n15207) );
  AND U17903 ( .A(n15132), .B(n14205), .Z(n15206) );
  NANDN U17904 ( .B(n8568), .A(n6961), .Z(n15170) );
  NAND U17905 ( .A(n15209), .B(n15210), .Z(n6961) );
  NAND U17906 ( .A(n6778), .B(\u_a23_core/imm32[13] ), .Z(n15210) );
  AND U17907 ( .A(n15211), .B(n15212), .Z(n15209) );
  NANDN U17908 ( .B(n6516), .A(\u_a23_core/barrel_shift_data_sel[1] ), .Z(
        n15212) );
  AND U17909 ( .A(n15213), .B(n15214), .Z(n6516) );
  AND U17910 ( .A(n15215), .B(n15216), .Z(n15214) );
  AND U17911 ( .A(n15217), .B(n15218), .Z(n15216) );
  AND U17912 ( .A(n15219), .B(n15220), .Z(n15218) );
  NAND U17913 ( .A(n14349), .B(\u_a23_core/u_execute/pc[13] ), .Z(n15220) );
  NANDN U17914 ( .B(n14350), .A(\u_a23_core/u_execute/u_register_bank/r14[13] ), .Z(n15219) );
  AND U17915 ( .A(n15221), .B(n15222), .Z(n15217) );
  NANDN U17916 ( .B(n14353), .A(\u_a23_core/u_execute/u_register_bank/r13[13] ), .Z(n15222) );
  NANDN U17917 ( .B(n14354), .A(\u_a23_core/u_execute/u_register_bank/r12[13] ), .Z(n15221) );
  AND U17918 ( .A(n15223), .B(n15224), .Z(n15215) );
  AND U17919 ( .A(n15225), .B(n15226), .Z(n15224) );
  NANDN U17920 ( .B(n14359), .A(\u_a23_core/u_execute/u_register_bank/r11[13] ), .Z(n15226) );
  NANDN U17921 ( .B(n14360), .A(\u_a23_core/u_execute/u_register_bank/r10[13] ), .Z(n15225) );
  AND U17922 ( .A(n15227), .B(n15228), .Z(n15223) );
  NANDN U17923 ( .B(n14363), .A(\u_a23_core/u_execute/u_register_bank/r9[13] ), 
        .Z(n15228) );
  NANDN U17924 ( .B(n14364), .A(\u_a23_core/u_execute/u_register_bank/r8[13] ), 
        .Z(n15227) );
  AND U17925 ( .A(n15229), .B(n15230), .Z(n15213) );
  AND U17926 ( .A(n15231), .B(n15232), .Z(n15230) );
  AND U17927 ( .A(n15233), .B(n15234), .Z(n15232) );
  NANDN U17928 ( .B(n14371), .A(\u_a23_core/u_execute/u_register_bank/r7[13] ), 
        .Z(n15234) );
  NANDN U17929 ( .B(n14372), .A(\u_a23_core/u_execute/u_register_bank/r6[13] ), 
        .Z(n15233) );
  AND U17930 ( .A(n15235), .B(n15236), .Z(n15231) );
  NANDN U17931 ( .B(n14375), .A(\u_a23_core/u_execute/u_register_bank/r5[13] ), 
        .Z(n15236) );
  NANDN U17932 ( .B(n14376), .A(\u_a23_core/u_execute/u_register_bank/r4[13] ), 
        .Z(n15235) );
  AND U17933 ( .A(n15237), .B(n15238), .Z(n15229) );
  AND U17934 ( .A(n15239), .B(n15240), .Z(n15238) );
  NANDN U17935 ( .B(n14381), .A(\u_a23_core/u_execute/u_register_bank/r3[13] ), 
        .Z(n15240) );
  NANDN U17936 ( .B(n14382), .A(\u_a23_core/u_execute/u_register_bank/r0[13] ), 
        .Z(n15239) );
  AND U17937 ( .A(n15241), .B(n15242), .Z(n15237) );
  NANDN U17938 ( .B(n14385), .A(\u_a23_core/u_execute/u_register_bank/r2[13] ), 
        .Z(n15242) );
  NANDN U17939 ( .B(n14386), .A(\u_a23_core/u_execute/u_register_bank/r1[13] ), 
        .Z(n15241) );
  NANDN U17940 ( .B(n14387), .A(\u_a23_core/read_data_s2[13] ), .Z(n15211) );
  NAND U17941 ( .A(n15243), .B(n15208), .Z(n8568) );
  AND U17942 ( .A(n15093), .B(n14237), .Z(n15243) );
  AND U17943 ( .A(n15244), .B(n15245), .Z(n14940) );
  AND U17944 ( .A(n15246), .B(n15247), .Z(n15245) );
  AND U17945 ( .A(n15248), .B(n15249), .Z(n15247) );
  NANDN U17946 ( .B(n8571), .A(n6956), .Z(n15249) );
  NAND U17947 ( .A(n15250), .B(n15251), .Z(n6956) );
  NAND U17948 ( .A(n6778), .B(\u_a23_core/imm32[12] ), .Z(n15251) );
  AND U17949 ( .A(n15252), .B(n15253), .Z(n15250) );
  NANDN U17950 ( .B(n6509), .A(\u_a23_core/barrel_shift_data_sel[1] ), .Z(
        n15253) );
  AND U17951 ( .A(n15254), .B(n15255), .Z(n6509) );
  AND U17952 ( .A(n15256), .B(n15257), .Z(n15255) );
  AND U17953 ( .A(n15258), .B(n15259), .Z(n15257) );
  AND U17954 ( .A(n15260), .B(n15261), .Z(n15259) );
  NAND U17955 ( .A(n14349), .B(\u_a23_core/u_execute/pc[12] ), .Z(n15261) );
  NANDN U17956 ( .B(n14350), .A(\u_a23_core/u_execute/u_register_bank/r14[12] ), .Z(n15260) );
  AND U17957 ( .A(n15262), .B(n15263), .Z(n15258) );
  NANDN U17958 ( .B(n14353), .A(\u_a23_core/u_execute/u_register_bank/r13[12] ), .Z(n15263) );
  NANDN U17959 ( .B(n14354), .A(\u_a23_core/u_execute/u_register_bank/r12[12] ), .Z(n15262) );
  AND U17960 ( .A(n15264), .B(n15265), .Z(n15256) );
  AND U17961 ( .A(n15266), .B(n15267), .Z(n15265) );
  NANDN U17962 ( .B(n14359), .A(\u_a23_core/u_execute/u_register_bank/r11[12] ), .Z(n15267) );
  NANDN U17963 ( .B(n14360), .A(\u_a23_core/u_execute/u_register_bank/r10[12] ), .Z(n15266) );
  AND U17964 ( .A(n15268), .B(n15269), .Z(n15264) );
  NANDN U17965 ( .B(n14363), .A(\u_a23_core/u_execute/u_register_bank/r9[12] ), 
        .Z(n15269) );
  NANDN U17966 ( .B(n14364), .A(\u_a23_core/u_execute/u_register_bank/r8[12] ), 
        .Z(n15268) );
  AND U17967 ( .A(n15270), .B(n15271), .Z(n15254) );
  AND U17968 ( .A(n15272), .B(n15273), .Z(n15271) );
  AND U17969 ( .A(n15274), .B(n15275), .Z(n15273) );
  NANDN U17970 ( .B(n14371), .A(\u_a23_core/u_execute/u_register_bank/r7[12] ), 
        .Z(n15275) );
  NANDN U17971 ( .B(n14372), .A(\u_a23_core/u_execute/u_register_bank/r6[12] ), 
        .Z(n15274) );
  AND U17972 ( .A(n15276), .B(n15277), .Z(n15272) );
  NANDN U17973 ( .B(n14375), .A(\u_a23_core/u_execute/u_register_bank/r5[12] ), 
        .Z(n15277) );
  NANDN U17974 ( .B(n14376), .A(\u_a23_core/u_execute/u_register_bank/r4[12] ), 
        .Z(n15276) );
  AND U17975 ( .A(n15278), .B(n15279), .Z(n15270) );
  AND U17976 ( .A(n15280), .B(n15281), .Z(n15279) );
  NANDN U17977 ( .B(n14381), .A(\u_a23_core/u_execute/u_register_bank/r3[12] ), 
        .Z(n15281) );
  NANDN U17978 ( .B(n14382), .A(\u_a23_core/u_execute/u_register_bank/r0[12] ), 
        .Z(n15280) );
  AND U17979 ( .A(n15282), .B(n15283), .Z(n15278) );
  NANDN U17980 ( .B(n14385), .A(\u_a23_core/u_execute/u_register_bank/r2[12] ), 
        .Z(n15283) );
  NANDN U17981 ( .B(n14386), .A(\u_a23_core/u_execute/u_register_bank/r1[12] ), 
        .Z(n15282) );
  NANDN U17982 ( .B(n14387), .A(\u_a23_core/read_data_s2[12] ), .Z(n15252) );
  NAND U17983 ( .A(n15284), .B(n15208), .Z(n8571) );
  AND U17984 ( .A(n15285), .B(n15286), .Z(n15208) );
  AND U17985 ( .A(n15287), .B(n15288), .Z(n15285) );
  NAND U17986 ( .A(n6988), .B(n14983), .Z(n15288) );
  OR U17987 ( .A(n15093), .B(n15132), .Z(n14983) );
  AND U17988 ( .A(n15132), .B(n14237), .Z(n15284) );
  NANDN U17989 ( .B(n8572), .A(n6960), .Z(n15248) );
  NAND U17990 ( .A(n15289), .B(n15290), .Z(n6960) );
  NAND U17991 ( .A(n6778), .B(\u_a23_core/imm32[11] ), .Z(n15290) );
  AND U17992 ( .A(n15291), .B(n15292), .Z(n15289) );
  NANDN U17993 ( .B(n6502), .A(\u_a23_core/barrel_shift_data_sel[1] ), .Z(
        n15292) );
  AND U17994 ( .A(n15293), .B(n15294), .Z(n6502) );
  AND U17995 ( .A(n15295), .B(n15296), .Z(n15294) );
  AND U17996 ( .A(n15297), .B(n15298), .Z(n15296) );
  AND U17997 ( .A(n15299), .B(n15300), .Z(n15298) );
  NAND U17998 ( .A(n14349), .B(\u_a23_core/u_execute/pc[11] ), .Z(n15300) );
  NANDN U17999 ( .B(n14350), .A(\u_a23_core/u_execute/u_register_bank/r14[11] ), .Z(n15299) );
  AND U18000 ( .A(n15301), .B(n15302), .Z(n15297) );
  NANDN U18001 ( .B(n14353), .A(\u_a23_core/u_execute/u_register_bank/r13[11] ), .Z(n15302) );
  NANDN U18002 ( .B(n14354), .A(\u_a23_core/u_execute/u_register_bank/r12[11] ), .Z(n15301) );
  AND U18003 ( .A(n15303), .B(n15304), .Z(n15295) );
  AND U18004 ( .A(n15305), .B(n15306), .Z(n15304) );
  NANDN U18005 ( .B(n14359), .A(\u_a23_core/u_execute/u_register_bank/r11[11] ), .Z(n15306) );
  NANDN U18006 ( .B(n14360), .A(\u_a23_core/u_execute/u_register_bank/r10[11] ), .Z(n15305) );
  AND U18007 ( .A(n15307), .B(n15308), .Z(n15303) );
  NANDN U18008 ( .B(n14363), .A(\u_a23_core/u_execute/u_register_bank/r9[11] ), 
        .Z(n15308) );
  NANDN U18009 ( .B(n14364), .A(\u_a23_core/u_execute/u_register_bank/r8[11] ), 
        .Z(n15307) );
  AND U18010 ( .A(n15309), .B(n15310), .Z(n15293) );
  AND U18011 ( .A(n15311), .B(n15312), .Z(n15310) );
  AND U18012 ( .A(n15313), .B(n15314), .Z(n15312) );
  NANDN U18013 ( .B(n14371), .A(\u_a23_core/u_execute/u_register_bank/r7[11] ), 
        .Z(n15314) );
  NANDN U18014 ( .B(n14372), .A(\u_a23_core/u_execute/u_register_bank/r6[11] ), 
        .Z(n15313) );
  AND U18015 ( .A(n15315), .B(n15316), .Z(n15311) );
  NANDN U18016 ( .B(n14375), .A(\u_a23_core/u_execute/u_register_bank/r5[11] ), 
        .Z(n15316) );
  NANDN U18017 ( .B(n14376), .A(\u_a23_core/u_execute/u_register_bank/r4[11] ), 
        .Z(n15315) );
  AND U18018 ( .A(n15317), .B(n15318), .Z(n15309) );
  AND U18019 ( .A(n15319), .B(n15320), .Z(n15318) );
  NANDN U18020 ( .B(n14381), .A(\u_a23_core/u_execute/u_register_bank/r3[11] ), 
        .Z(n15320) );
  NANDN U18021 ( .B(n14382), .A(\u_a23_core/u_execute/u_register_bank/r0[11] ), 
        .Z(n15319) );
  AND U18022 ( .A(n15321), .B(n15322), .Z(n15317) );
  NANDN U18023 ( .B(n14385), .A(\u_a23_core/u_execute/u_register_bank/r2[11] ), 
        .Z(n15322) );
  NANDN U18024 ( .B(n14386), .A(\u_a23_core/u_execute/u_register_bank/r1[11] ), 
        .Z(n15321) );
  NANDN U18025 ( .B(n14387), .A(\u_a23_core/read_data_s2[11] ), .Z(n15291) );
  NAND U18026 ( .A(n15323), .B(n15093), .Z(n8572) );
  AND U18027 ( .A(n15324), .B(n15325), .Z(n15246) );
  NANDN U18028 ( .B(n8579), .A(n6957), .Z(n15325) );
  NAND U18029 ( .A(n15326), .B(n15327), .Z(n6957) );
  NAND U18030 ( .A(n6778), .B(\u_a23_core/imm32[10] ), .Z(n15327) );
  AND U18031 ( .A(n15328), .B(n15329), .Z(n15326) );
  NANDN U18032 ( .B(n6495), .A(\u_a23_core/barrel_shift_data_sel[1] ), .Z(
        n15329) );
  AND U18033 ( .A(n15330), .B(n15331), .Z(n6495) );
  AND U18034 ( .A(n15332), .B(n15333), .Z(n15331) );
  AND U18035 ( .A(n15334), .B(n15335), .Z(n15333) );
  AND U18036 ( .A(n15336), .B(n15337), .Z(n15335) );
  NAND U18037 ( .A(n14349), .B(\u_a23_core/u_execute/pc[10] ), .Z(n15337) );
  NANDN U18038 ( .B(n14350), .A(\u_a23_core/u_execute/u_register_bank/r14[10] ), .Z(n15336) );
  AND U18039 ( .A(n15338), .B(n15339), .Z(n15334) );
  NANDN U18040 ( .B(n14353), .A(\u_a23_core/u_execute/u_register_bank/r13[10] ), .Z(n15339) );
  NANDN U18041 ( .B(n14354), .A(\u_a23_core/u_execute/u_register_bank/r12[10] ), .Z(n15338) );
  AND U18042 ( .A(n15340), .B(n15341), .Z(n15332) );
  AND U18043 ( .A(n15342), .B(n15343), .Z(n15341) );
  NANDN U18044 ( .B(n14359), .A(\u_a23_core/u_execute/u_register_bank/r11[10] ), .Z(n15343) );
  NANDN U18045 ( .B(n14360), .A(\u_a23_core/u_execute/u_register_bank/r10[10] ), .Z(n15342) );
  AND U18046 ( .A(n15344), .B(n15345), .Z(n15340) );
  NANDN U18047 ( .B(n14363), .A(\u_a23_core/u_execute/u_register_bank/r9[10] ), 
        .Z(n15345) );
  NANDN U18048 ( .B(n14364), .A(\u_a23_core/u_execute/u_register_bank/r8[10] ), 
        .Z(n15344) );
  AND U18049 ( .A(n15346), .B(n15347), .Z(n15330) );
  AND U18050 ( .A(n15348), .B(n15349), .Z(n15347) );
  AND U18051 ( .A(n15350), .B(n15351), .Z(n15349) );
  NANDN U18052 ( .B(n14371), .A(\u_a23_core/u_execute/u_register_bank/r7[10] ), 
        .Z(n15351) );
  NANDN U18053 ( .B(n14372), .A(\u_a23_core/u_execute/u_register_bank/r6[10] ), 
        .Z(n15350) );
  AND U18054 ( .A(n15352), .B(n15353), .Z(n15348) );
  NANDN U18055 ( .B(n14375), .A(\u_a23_core/u_execute/u_register_bank/r5[10] ), 
        .Z(n15353) );
  NANDN U18056 ( .B(n14376), .A(\u_a23_core/u_execute/u_register_bank/r4[10] ), 
        .Z(n15352) );
  AND U18057 ( .A(n15354), .B(n15355), .Z(n15346) );
  AND U18058 ( .A(n15356), .B(n15357), .Z(n15355) );
  NANDN U18059 ( .B(n14381), .A(\u_a23_core/u_execute/u_register_bank/r3[10] ), 
        .Z(n15357) );
  NANDN U18060 ( .B(n14382), .A(\u_a23_core/u_execute/u_register_bank/r0[10] ), 
        .Z(n15356) );
  AND U18061 ( .A(n15358), .B(n15359), .Z(n15354) );
  NANDN U18062 ( .B(n14385), .A(\u_a23_core/u_execute/u_register_bank/r2[10] ), 
        .Z(n15359) );
  NANDN U18063 ( .B(n14386), .A(\u_a23_core/u_execute/u_register_bank/r1[10] ), 
        .Z(n15358) );
  NANDN U18064 ( .B(n14387), .A(\u_a23_core/read_data_s2[10] ), .Z(n15328) );
  NAND U18065 ( .A(n15132), .B(n15323), .Z(n8579) );
  ANDN U18066 ( .A(n15287), .B(n14390), .Z(n15323) );
  NANDN U18067 ( .B(n8580), .A(n6947), .Z(n15324) );
  NAND U18068 ( .A(n15360), .B(n15361), .Z(n6947) );
  NAND U18069 ( .A(n6778), .B(\u_a23_core/imm32[9] ), .Z(n15361) );
  AND U18070 ( .A(n15362), .B(n15363), .Z(n15360) );
  NANDN U18071 ( .B(n6488), .A(\u_a23_core/barrel_shift_data_sel[1] ), .Z(
        n15363) );
  AND U18072 ( .A(n15364), .B(n15365), .Z(n6488) );
  AND U18073 ( .A(n15366), .B(n15367), .Z(n15365) );
  AND U18074 ( .A(n15368), .B(n15369), .Z(n15367) );
  AND U18075 ( .A(n15370), .B(n15371), .Z(n15369) );
  NAND U18076 ( .A(n14349), .B(\u_a23_core/u_execute/pc[9] ), .Z(n15371) );
  NANDN U18077 ( .B(n14350), .A(\u_a23_core/u_execute/u_register_bank/r14[9] ), 
        .Z(n15370) );
  AND U18078 ( .A(n15372), .B(n15373), .Z(n15368) );
  NANDN U18079 ( .B(n14353), .A(\u_a23_core/u_execute/u_register_bank/r13[9] ), 
        .Z(n15373) );
  NANDN U18080 ( .B(n14354), .A(\u_a23_core/u_execute/u_register_bank/r12[9] ), 
        .Z(n15372) );
  AND U18081 ( .A(n15374), .B(n15375), .Z(n15366) );
  AND U18082 ( .A(n15376), .B(n15377), .Z(n15375) );
  NANDN U18083 ( .B(n14359), .A(\u_a23_core/u_execute/u_register_bank/r11[9] ), 
        .Z(n15377) );
  NANDN U18084 ( .B(n14360), .A(\u_a23_core/u_execute/u_register_bank/r10[9] ), 
        .Z(n15376) );
  AND U18085 ( .A(n15378), .B(n15379), .Z(n15374) );
  NANDN U18086 ( .B(n14363), .A(\u_a23_core/u_execute/u_register_bank/r9[9] ), 
        .Z(n15379) );
  NANDN U18087 ( .B(n14364), .A(\u_a23_core/u_execute/u_register_bank/r8[9] ), 
        .Z(n15378) );
  AND U18088 ( .A(n15380), .B(n15381), .Z(n15364) );
  AND U18089 ( .A(n15382), .B(n15383), .Z(n15381) );
  AND U18090 ( .A(n15384), .B(n15385), .Z(n15383) );
  NANDN U18091 ( .B(n14371), .A(\u_a23_core/u_execute/u_register_bank/r7[9] ), 
        .Z(n15385) );
  NANDN U18092 ( .B(n14372), .A(\u_a23_core/u_execute/u_register_bank/r6[9] ), 
        .Z(n15384) );
  AND U18093 ( .A(n15386), .B(n15387), .Z(n15382) );
  NANDN U18094 ( .B(n14375), .A(\u_a23_core/u_execute/u_register_bank/r5[9] ), 
        .Z(n15387) );
  NANDN U18095 ( .B(n14376), .A(\u_a23_core/u_execute/u_register_bank/r4[9] ), 
        .Z(n15386) );
  AND U18096 ( .A(n15388), .B(n15389), .Z(n15380) );
  AND U18097 ( .A(n15390), .B(n15391), .Z(n15389) );
  NANDN U18098 ( .B(n14381), .A(\u_a23_core/u_execute/u_register_bank/r3[9] ), 
        .Z(n15391) );
  NANDN U18099 ( .B(n14382), .A(\u_a23_core/u_execute/u_register_bank/r0[9] ), 
        .Z(n15390) );
  AND U18100 ( .A(n15392), .B(n15393), .Z(n15388) );
  NANDN U18101 ( .B(n14385), .A(\u_a23_core/u_execute/u_register_bank/r2[9] ), 
        .Z(n15393) );
  NANDN U18102 ( .B(n14386), .A(\u_a23_core/u_execute/u_register_bank/r1[9] ), 
        .Z(n15392) );
  NANDN U18103 ( .B(n14387), .A(\u_a23_core/read_data_s2[9] ), .Z(n15362) );
  NAND U18104 ( .A(n9271), .B(n15287), .Z(n8580) );
  AND U18105 ( .A(n15394), .B(n15395), .Z(n15244) );
  AND U18106 ( .A(n15396), .B(n15397), .Z(n15395) );
  NANDN U18107 ( .B(n8583), .A(n6946), .Z(n15397) );
  NAND U18108 ( .A(n15398), .B(n15399), .Z(n6946) );
  NAND U18109 ( .A(n6778), .B(\u_a23_core/imm32[8] ), .Z(n15399) );
  AND U18110 ( .A(n15400), .B(n15401), .Z(n15398) );
  NANDN U18111 ( .B(n6481), .A(\u_a23_core/barrel_shift_data_sel[1] ), .Z(
        n15401) );
  AND U18112 ( .A(n15402), .B(n15403), .Z(n6481) );
  AND U18113 ( .A(n15404), .B(n15405), .Z(n15403) );
  AND U18114 ( .A(n15406), .B(n15407), .Z(n15405) );
  AND U18115 ( .A(n15408), .B(n15409), .Z(n15407) );
  NAND U18116 ( .A(n14349), .B(\u_a23_core/u_execute/pc[8] ), .Z(n15409) );
  NANDN U18117 ( .B(n14350), .A(\u_a23_core/u_execute/u_register_bank/r14[8] ), 
        .Z(n15408) );
  AND U18118 ( .A(n15410), .B(n15411), .Z(n15406) );
  NANDN U18119 ( .B(n14353), .A(\u_a23_core/u_execute/u_register_bank/r13[8] ), 
        .Z(n15411) );
  NANDN U18120 ( .B(n14354), .A(\u_a23_core/u_execute/u_register_bank/r12[8] ), 
        .Z(n15410) );
  AND U18121 ( .A(n15412), .B(n15413), .Z(n15404) );
  AND U18122 ( .A(n15414), .B(n15415), .Z(n15413) );
  NANDN U18123 ( .B(n14359), .A(\u_a23_core/u_execute/u_register_bank/r11[8] ), 
        .Z(n15415) );
  NANDN U18124 ( .B(n14360), .A(\u_a23_core/u_execute/u_register_bank/r10[8] ), 
        .Z(n15414) );
  AND U18125 ( .A(n15416), .B(n15417), .Z(n15412) );
  NANDN U18126 ( .B(n14363), .A(\u_a23_core/u_execute/u_register_bank/r9[8] ), 
        .Z(n15417) );
  NANDN U18127 ( .B(n14364), .A(\u_a23_core/u_execute/u_register_bank/r8[8] ), 
        .Z(n15416) );
  AND U18128 ( .A(n15418), .B(n15419), .Z(n15402) );
  AND U18129 ( .A(n15420), .B(n15421), .Z(n15419) );
  AND U18130 ( .A(n15422), .B(n15423), .Z(n15421) );
  NANDN U18131 ( .B(n14371), .A(\u_a23_core/u_execute/u_register_bank/r7[8] ), 
        .Z(n15423) );
  NANDN U18132 ( .B(n14372), .A(\u_a23_core/u_execute/u_register_bank/r6[8] ), 
        .Z(n15422) );
  AND U18133 ( .A(n15424), .B(n15425), .Z(n15420) );
  NANDN U18134 ( .B(n14375), .A(\u_a23_core/u_execute/u_register_bank/r5[8] ), 
        .Z(n15425) );
  NANDN U18135 ( .B(n14376), .A(\u_a23_core/u_execute/u_register_bank/r4[8] ), 
        .Z(n15424) );
  AND U18136 ( .A(n15426), .B(n15427), .Z(n15418) );
  AND U18137 ( .A(n15428), .B(n15429), .Z(n15427) );
  NANDN U18138 ( .B(n14381), .A(\u_a23_core/u_execute/u_register_bank/r3[8] ), 
        .Z(n15429) );
  NANDN U18139 ( .B(n14382), .A(\u_a23_core/u_execute/u_register_bank/r0[8] ), 
        .Z(n15428) );
  AND U18140 ( .A(n15430), .B(n15431), .Z(n15426) );
  NANDN U18141 ( .B(n14385), .A(\u_a23_core/u_execute/u_register_bank/r2[8] ), 
        .Z(n15431) );
  NANDN U18142 ( .B(n14386), .A(\u_a23_core/u_execute/u_register_bank/r1[8] ), 
        .Z(n15430) );
  NANDN U18143 ( .B(n14387), .A(\u_a23_core/read_data_s2[8] ), .Z(n15400) );
  NAND U18144 ( .A(n6990), .B(n15287), .Z(n8583) );
  AND U18145 ( .A(n15432), .B(n15433), .Z(n15287) );
  AND U18146 ( .A(n15434), .B(n15435), .Z(n15432) );
  OR U18147 ( .A(n15286), .B(n14305), .Z(n15435) );
  NAND U18148 ( .A(n14237), .B(n9271), .Z(n15434) );
  NANDN U18149 ( .B(n8584), .A(n6943), .Z(n15396) );
  NAND U18150 ( .A(n15436), .B(n15437), .Z(n6943) );
  NAND U18151 ( .A(n6778), .B(\u_a23_core/imm32[7] ), .Z(n15437) );
  AND U18152 ( .A(n15438), .B(n15439), .Z(n15436) );
  NANDN U18153 ( .B(n6474), .A(\u_a23_core/barrel_shift_data_sel[1] ), .Z(
        n15439) );
  AND U18154 ( .A(n15440), .B(n15441), .Z(n6474) );
  AND U18155 ( .A(n15442), .B(n15443), .Z(n15441) );
  AND U18156 ( .A(n15444), .B(n15445), .Z(n15443) );
  AND U18157 ( .A(n15446), .B(n15447), .Z(n15445) );
  NAND U18158 ( .A(n14349), .B(\u_a23_core/u_execute/pc[7] ), .Z(n15447) );
  NANDN U18159 ( .B(n14350), .A(\u_a23_core/u_execute/u_register_bank/r14[7] ), 
        .Z(n15446) );
  AND U18160 ( .A(n15448), .B(n15449), .Z(n15444) );
  NANDN U18161 ( .B(n14353), .A(\u_a23_core/u_execute/u_register_bank/r13[7] ), 
        .Z(n15449) );
  NANDN U18162 ( .B(n14354), .A(\u_a23_core/u_execute/u_register_bank/r12[7] ), 
        .Z(n15448) );
  AND U18163 ( .A(n15450), .B(n15451), .Z(n15442) );
  AND U18164 ( .A(n15452), .B(n15453), .Z(n15451) );
  NANDN U18165 ( .B(n14359), .A(\u_a23_core/u_execute/u_register_bank/r11[7] ), 
        .Z(n15453) );
  NANDN U18166 ( .B(n14360), .A(\u_a23_core/u_execute/u_register_bank/r10[7] ), 
        .Z(n15452) );
  AND U18167 ( .A(n15454), .B(n15455), .Z(n15450) );
  NANDN U18168 ( .B(n14363), .A(\u_a23_core/u_execute/u_register_bank/r9[7] ), 
        .Z(n15455) );
  NANDN U18169 ( .B(n14364), .A(\u_a23_core/u_execute/u_register_bank/r8[7] ), 
        .Z(n15454) );
  AND U18170 ( .A(n15456), .B(n15457), .Z(n15440) );
  AND U18171 ( .A(n15458), .B(n15459), .Z(n15457) );
  AND U18172 ( .A(n15460), .B(n15461), .Z(n15459) );
  NANDN U18173 ( .B(n14371), .A(\u_a23_core/u_execute/u_register_bank/r7[7] ), 
        .Z(n15461) );
  NANDN U18174 ( .B(n14372), .A(\u_a23_core/u_execute/u_register_bank/r6[7] ), 
        .Z(n15460) );
  AND U18175 ( .A(n15462), .B(n15463), .Z(n15458) );
  NANDN U18176 ( .B(n14375), .A(\u_a23_core/u_execute/u_register_bank/r5[7] ), 
        .Z(n15463) );
  NANDN U18177 ( .B(n14376), .A(\u_a23_core/u_execute/u_register_bank/r4[7] ), 
        .Z(n15462) );
  AND U18178 ( .A(n15464), .B(n15465), .Z(n15456) );
  AND U18179 ( .A(n15466), .B(n15467), .Z(n15465) );
  NANDN U18180 ( .B(n14381), .A(\u_a23_core/u_execute/u_register_bank/r3[7] ), 
        .Z(n15467) );
  NANDN U18181 ( .B(n14382), .A(\u_a23_core/u_execute/u_register_bank/r0[7] ), 
        .Z(n15466) );
  AND U18182 ( .A(n15468), .B(n15469), .Z(n15464) );
  NANDN U18183 ( .B(n14385), .A(\u_a23_core/u_execute/u_register_bank/r2[7] ), 
        .Z(n15469) );
  NANDN U18184 ( .B(n14386), .A(\u_a23_core/u_execute/u_register_bank/r1[7] ), 
        .Z(n15468) );
  NANDN U18185 ( .B(n14387), .A(\u_a23_core/read_data_s2[7] ), .Z(n15438) );
  NAND U18186 ( .A(n15470), .B(n15433), .Z(n8584) );
  AND U18187 ( .A(n14205), .B(n9271), .Z(n15470) );
  AND U18188 ( .A(n15471), .B(n15472), .Z(n15394) );
  NANDN U18189 ( .B(n8589), .A(n6942), .Z(n15472) );
  NAND U18190 ( .A(n15473), .B(n15474), .Z(n6942) );
  NAND U18191 ( .A(n6778), .B(\u_a23_core/imm32[6] ), .Z(n15474) );
  AND U18192 ( .A(n15475), .B(n15476), .Z(n15473) );
  NANDN U18193 ( .B(n6467), .A(\u_a23_core/barrel_shift_data_sel[1] ), .Z(
        n15476) );
  AND U18194 ( .A(n15477), .B(n15478), .Z(n6467) );
  AND U18195 ( .A(n15479), .B(n15480), .Z(n15478) );
  AND U18196 ( .A(n15481), .B(n15482), .Z(n15480) );
  AND U18197 ( .A(n15483), .B(n15484), .Z(n15482) );
  NAND U18198 ( .A(n14349), .B(\u_a23_core/u_execute/pc[6] ), .Z(n15484) );
  NANDN U18199 ( .B(n14350), .A(\u_a23_core/u_execute/u_register_bank/r14[6] ), 
        .Z(n15483) );
  AND U18200 ( .A(n15485), .B(n15486), .Z(n15481) );
  NANDN U18201 ( .B(n14353), .A(\u_a23_core/u_execute/u_register_bank/r13[6] ), 
        .Z(n15486) );
  NANDN U18202 ( .B(n14354), .A(\u_a23_core/u_execute/u_register_bank/r12[6] ), 
        .Z(n15485) );
  AND U18203 ( .A(n15487), .B(n15488), .Z(n15479) );
  AND U18204 ( .A(n15489), .B(n15490), .Z(n15488) );
  NANDN U18205 ( .B(n14359), .A(\u_a23_core/u_execute/u_register_bank/r11[6] ), 
        .Z(n15490) );
  NANDN U18206 ( .B(n14360), .A(\u_a23_core/u_execute/u_register_bank/r10[6] ), 
        .Z(n15489) );
  AND U18207 ( .A(n15491), .B(n15492), .Z(n15487) );
  NANDN U18208 ( .B(n14363), .A(\u_a23_core/u_execute/u_register_bank/r9[6] ), 
        .Z(n15492) );
  NANDN U18209 ( .B(n14364), .A(\u_a23_core/u_execute/u_register_bank/r8[6] ), 
        .Z(n15491) );
  AND U18210 ( .A(n15493), .B(n15494), .Z(n15477) );
  AND U18211 ( .A(n15495), .B(n15496), .Z(n15494) );
  AND U18212 ( .A(n15497), .B(n15498), .Z(n15496) );
  NANDN U18213 ( .B(n14371), .A(\u_a23_core/u_execute/u_register_bank/r7[6] ), 
        .Z(n15498) );
  NANDN U18214 ( .B(n14372), .A(\u_a23_core/u_execute/u_register_bank/r6[6] ), 
        .Z(n15497) );
  AND U18215 ( .A(n15499), .B(n15500), .Z(n15495) );
  NANDN U18216 ( .B(n14375), .A(\u_a23_core/u_execute/u_register_bank/r5[6] ), 
        .Z(n15500) );
  NANDN U18217 ( .B(n14376), .A(\u_a23_core/u_execute/u_register_bank/r4[6] ), 
        .Z(n15499) );
  AND U18218 ( .A(n15501), .B(n15502), .Z(n15493) );
  AND U18219 ( .A(n15503), .B(n15504), .Z(n15502) );
  NANDN U18220 ( .B(n14381), .A(\u_a23_core/u_execute/u_register_bank/r3[6] ), 
        .Z(n15504) );
  NANDN U18221 ( .B(n14382), .A(\u_a23_core/u_execute/u_register_bank/r0[6] ), 
        .Z(n15503) );
  AND U18222 ( .A(n15505), .B(n15506), .Z(n15501) );
  NANDN U18223 ( .B(n14385), .A(\u_a23_core/u_execute/u_register_bank/r2[6] ), 
        .Z(n15506) );
  NANDN U18224 ( .B(n14386), .A(\u_a23_core/u_execute/u_register_bank/r1[6] ), 
        .Z(n15505) );
  NANDN U18225 ( .B(n14387), .A(\u_a23_core/read_data_s2[6] ), .Z(n15475) );
  NAND U18226 ( .A(n15507), .B(n15433), .Z(n8589) );
  AND U18227 ( .A(n6990), .B(n14205), .Z(n15507) );
  NANDN U18228 ( .B(n8590), .A(n6937), .Z(n15471) );
  NAND U18229 ( .A(n15508), .B(n15509), .Z(n6937) );
  NAND U18230 ( .A(n6778), .B(\u_a23_core/imm32[5] ), .Z(n15509) );
  NOR U18231 ( .A(\u_a23_core/barrel_shift_data_sel[1] ), .B(
        \u_a23_core/barrel_shift_data_sel[0] ), .Z(n6778) );
  AND U18232 ( .A(n15510), .B(n15511), .Z(n15508) );
  NANDN U18233 ( .B(n6460), .A(\u_a23_core/barrel_shift_data_sel[1] ), .Z(
        n15511) );
  AND U18234 ( .A(n15512), .B(n15513), .Z(n6460) );
  AND U18235 ( .A(n15514), .B(n15515), .Z(n15513) );
  AND U18236 ( .A(n15516), .B(n15517), .Z(n15515) );
  AND U18237 ( .A(n15518), .B(n15519), .Z(n15517) );
  NAND U18238 ( .A(n14349), .B(\u_a23_core/u_execute/pc[5] ), .Z(n15519) );
  AND U18239 ( .A(n15520), .B(n15521), .Z(n14349) );
  NANDN U18240 ( .B(n14350), .A(\u_a23_core/u_execute/u_register_bank/r14[5] ), 
        .Z(n15518) );
  NAND U18241 ( .A(n15521), .B(n15522), .Z(n14350) );
  AND U18242 ( .A(n15523), .B(n15524), .Z(n15516) );
  NANDN U18243 ( .B(n14353), .A(\u_a23_core/u_execute/u_register_bank/r13[5] ), 
        .Z(n15524) );
  NAND U18244 ( .A(n15521), .B(n15525), .Z(n14353) );
  NANDN U18245 ( .B(n14354), .A(\u_a23_core/u_execute/u_register_bank/r12[5] ), 
        .Z(n15523) );
  NAND U18246 ( .A(n15521), .B(n15526), .Z(n14354) );
  AND U18247 ( .A(\u_a23_core/rm_sel[3] ), .B(\u_a23_core/rm_sel[2] ), .Z(
        n15521) );
  AND U18248 ( .A(n15527), .B(n15528), .Z(n15514) );
  AND U18249 ( .A(n15529), .B(n15530), .Z(n15528) );
  NANDN U18250 ( .B(n14359), .A(\u_a23_core/u_execute/u_register_bank/r11[5] ), 
        .Z(n15530) );
  NAND U18251 ( .A(n15531), .B(n15520), .Z(n14359) );
  NANDN U18252 ( .B(n14360), .A(\u_a23_core/u_execute/u_register_bank/r10[5] ), 
        .Z(n15529) );
  NAND U18253 ( .A(n15522), .B(n15531), .Z(n14360) );
  AND U18254 ( .A(n15532), .B(n15533), .Z(n15527) );
  NANDN U18255 ( .B(n14363), .A(\u_a23_core/u_execute/u_register_bank/r9[5] ), 
        .Z(n15533) );
  NAND U18256 ( .A(n15525), .B(n15531), .Z(n14363) );
  NANDN U18257 ( .B(n14364), .A(\u_a23_core/u_execute/u_register_bank/r8[5] ), 
        .Z(n15532) );
  NAND U18258 ( .A(n15526), .B(n15531), .Z(n14364) );
  AND U18259 ( .A(\u_a23_core/rm_sel[3] ), .B(n15534), .Z(n15531) );
  AND U18260 ( .A(n15535), .B(n15536), .Z(n15512) );
  AND U18261 ( .A(n15537), .B(n15538), .Z(n15536) );
  AND U18262 ( .A(n15539), .B(n15540), .Z(n15538) );
  NANDN U18263 ( .B(n14371), .A(\u_a23_core/u_execute/u_register_bank/r7[5] ), 
        .Z(n15540) );
  NAND U18264 ( .A(n15541), .B(n15520), .Z(n14371) );
  NANDN U18265 ( .B(n14372), .A(\u_a23_core/u_execute/u_register_bank/r6[5] ), 
        .Z(n15539) );
  NAND U18266 ( .A(n15522), .B(n15541), .Z(n14372) );
  AND U18267 ( .A(n15542), .B(n15543), .Z(n15537) );
  NANDN U18268 ( .B(n14375), .A(\u_a23_core/u_execute/u_register_bank/r5[5] ), 
        .Z(n15543) );
  NAND U18269 ( .A(n15525), .B(n15541), .Z(n14375) );
  NANDN U18270 ( .B(n14376), .A(\u_a23_core/u_execute/u_register_bank/r4[5] ), 
        .Z(n15542) );
  NAND U18271 ( .A(n15526), .B(n15541), .Z(n14376) );
  NOR U18272 ( .A(n15534), .B(\u_a23_core/rm_sel[3] ), .Z(n15541) );
  IV U18273 ( .A(\u_a23_core/rm_sel[2] ), .Z(n15534) );
  AND U18274 ( .A(n15544), .B(n15545), .Z(n15535) );
  AND U18275 ( .A(n15546), .B(n15547), .Z(n15545) );
  NANDN U18276 ( .B(n14381), .A(\u_a23_core/u_execute/u_register_bank/r3[5] ), 
        .Z(n15547) );
  NAND U18277 ( .A(n15548), .B(n15520), .Z(n14381) );
  ANDN U18278 ( .A(\u_a23_core/rm_sel[0] ), .B(n15549), .Z(n15520) );
  NANDN U18279 ( .B(n14382), .A(\u_a23_core/u_execute/u_register_bank/r0[5] ), 
        .Z(n15546) );
  NAND U18280 ( .A(n15526), .B(n15548), .Z(n14382) );
  ANDN U18281 ( .A(n15550), .B(\u_a23_core/rm_sel[1] ), .Z(n15526) );
  AND U18282 ( .A(n15551), .B(n15552), .Z(n15544) );
  NANDN U18283 ( .B(n14385), .A(\u_a23_core/u_execute/u_register_bank/r2[5] ), 
        .Z(n15552) );
  NAND U18284 ( .A(n15522), .B(n15548), .Z(n14385) );
  ANDN U18285 ( .A(\u_a23_core/rm_sel[1] ), .B(\u_a23_core/rm_sel[0] ), .Z(
        n15522) );
  NANDN U18286 ( .B(n14386), .A(\u_a23_core/u_execute/u_register_bank/r1[5] ), 
        .Z(n15551) );
  NAND U18287 ( .A(n15525), .B(n15548), .Z(n14386) );
  NOR U18288 ( .A(\u_a23_core/rm_sel[2] ), .B(\u_a23_core/rm_sel[3] ), .Z(
        n15548) );
  ANDN U18289 ( .A(n15549), .B(n15550), .Z(n15525) );
  IV U18290 ( .A(\u_a23_core/rm_sel[0] ), .Z(n15550) );
  IV U18291 ( .A(\u_a23_core/rm_sel[1] ), .Z(n15549) );
  NANDN U18292 ( .B(n14387), .A(\u_a23_core/read_data_s2[5] ), .Z(n15510) );
  NANDN U18293 ( .B(\u_a23_core/barrel_shift_data_sel[1] ), .A(
        \u_a23_core/barrel_shift_data_sel[0] ), .Z(n14387) );
  NAND U18294 ( .A(n15553), .B(n15433), .Z(n8590) );
  ANDN U18295 ( .A(n15554), .B(n14318), .Z(n15433) );
  IV U18296 ( .A(n9270), .Z(n14318) );
  ANDN U18297 ( .A(n15555), .B(\u_a23_core/shift_imm_zero ), .Z(n9270) );
  NAND U18298 ( .A(n14218), .B(n14325), .Z(n15555) );
  ANDN U18299 ( .A(n14299), .B(n14390), .Z(n14325) );
  ANDN U18300 ( .A(n15022), .B(n14226), .Z(n14299) );
  NANDN U18301 ( .B(n15556), .A(n14204), .Z(n14226) );
  NANDN U18302 ( .B(n15557), .A(n15558), .Z(n14204) );
  NANDN U18303 ( .B(n6989), .A(n16630), .Z(n15558) );
  NAND U18304 ( .A(n16632), .B(n16631), .Z(n6989) );
  IV U18305 ( .A(n14225), .Z(n14218) );
  AND U18306 ( .A(n15559), .B(n15560), .Z(n15554) );
  OR U18307 ( .A(n15286), .B(n14390), .Z(n15560) );
  IV U18308 ( .A(n6988), .Z(n14390) );
  ANDN U18309 ( .A(n14205), .B(n14324), .Z(n6988) );
  IV U18310 ( .A(n14305), .Z(n14205) );
  NAND U18311 ( .A(n15561), .B(n15562), .Z(n14305) );
  NANDN U18312 ( .B(n15557), .A(\u_a23_core/u_execute/rs[1] ), .Z(n15562) );
  NAND U18313 ( .A(n15563), .B(\u_a23_core/imm_shift_amount[1] ), .Z(n15561)
         );
  ANDN U18314 ( .A(n15564), .B(n6990), .Z(n15286) );
  IV U18315 ( .A(n9271), .Z(n15564) );
  NAND U18316 ( .A(n14237), .B(n6990), .Z(n15559) );
  ANDN U18317 ( .A(n15132), .B(n14295), .Z(n6990) );
  NOR U18318 ( .A(n14225), .B(n15556), .Z(n15132) );
  AND U18319 ( .A(n14237), .B(n9271), .Z(n15553) );
  ANDN U18320 ( .A(n15093), .B(n14295), .Z(n9271) );
  IV U18321 ( .A(n15022), .Z(n14295) );
  AND U18322 ( .A(n15565), .B(n15566), .Z(n15022) );
  NAND U18323 ( .A(n15563), .B(\u_a23_core/imm_shift_amount[3] ), .Z(n15566)
         );
  AND U18324 ( .A(n15567), .B(n15568), .Z(n15565) );
  NAND U18325 ( .A(n15569), .B(\u_a23_core/read_data_alignment[3] ), .Z(n15568) );
  NANDN U18326 ( .B(n15557), .A(\u_a23_core/u_execute/rs[3] ), .Z(n15567) );
  IV U18327 ( .A(n16628), .Z(\u_a23_core/u_execute/rs[3] ) );
  ANDN U18328 ( .A(n14225), .B(n15556), .Z(n15093) );
  NAND U18329 ( .A(n15570), .B(n15571), .Z(n15556) );
  NAND U18330 ( .A(n15563), .B(\u_a23_core/imm_shift_amount[4] ), .Z(n15571)
         );
  AND U18331 ( .A(n15572), .B(n15573), .Z(n15570) );
  NAND U18332 ( .A(n15569), .B(\u_a23_core/read_data_alignment[4] ), .Z(n15573) );
  AND U18333 ( .A(\u_a23_core/barrel_shift_amount_sel[0] ), .B(
        \u_a23_core/barrel_shift_amount_sel[1] ), .Z(n15569) );
  NANDN U18334 ( .B(n15557), .A(\u_a23_core/u_execute/rs[4] ), .Z(n15572) );
  IV U18335 ( .A(n16629), .Z(\u_a23_core/u_execute/rs[4] ) );
  NAND U18336 ( .A(n15574), .B(n15575), .Z(n14225) );
  NANDN U18337 ( .B(n15557), .A(\u_a23_core/u_execute/rs[0] ), .Z(n15575) );
  NAND U18338 ( .A(n15563), .B(\u_a23_core/imm_shift_amount[0] ), .Z(n15574)
         );
  IV U18339 ( .A(n14324), .Z(n14237) );
  NAND U18340 ( .A(n15576), .B(n15577), .Z(n14324) );
  NANDN U18341 ( .B(n15557), .A(\u_a23_core/u_execute/rs[2] ), .Z(n15577) );
  IV U18342 ( .A(n16625), .Z(\u_a23_core/u_execute/rs[2] ) );
  NAND U18343 ( .A(n15578), .B(\u_a23_core/barrel_shift_amount_sel[0] ), .Z(
        n15557) );
  NAND U18344 ( .A(n15563), .B(\u_a23_core/imm_shift_amount[2] ), .Z(n15576)
         );
  NOR U18345 ( .A(n15578), .B(\u_a23_core/barrel_shift_amount_sel[0] ), .Z(
        n15563) );
  IV U18346 ( .A(\u_a23_core/barrel_shift_amount_sel[1] ), .Z(n15578) );
  IV U18347 ( .A(\u_a23_core/u_execute/rn[2] ), .Z(n14186) );
  NAND U18348 ( .A(n6765), .B(\u_a23_core/u_execute/u_alu/fadder_out[2] ), .Z(
        n14166) );
  AND U18349 ( .A(n15579), .B(n14182), .Z(n6765) );
  ANDN U18350 ( .A(n15580), .B(\u_a23_core/alu_function[3] ), .Z(n14182) );
  IV U18351 ( .A(\u_a23_core/alu_function[2] ), .Z(n15580) );
  AND U18352 ( .A(\u_a23_core/alu_function[0] ), .B(n14180), .Z(n15579) );
  IV U18353 ( .A(\u_a23_core/alu_function[1] ), .Z(n14180) );
  IV U18354 ( .A(n8393), .Z(n14165) );
  NAND U18355 ( .A(n15581), .B(n15582), .Z(n8393) );
  NAND U18356 ( .A(\u_a23_core/address_sel[0] ), .B(n15583), .Z(n15582) );
  AND U18357 ( .A(n14160), .B(n14162), .Z(n15583) );
  NANDN U18358 ( .B(n14158), .A(n5930), .Z(n15581) );
  IV U18359 ( .A(n6099), .Z(n5930) );
  MUX U18360 ( .IN0(n15584), .IN1(n15585), .SEL(\u_a23_core/condition[3] ), 
        .F(n6099) );
  NAND U18361 ( .A(n15586), .B(n15587), .Z(n15585) );
  NAND U18362 ( .A(n15588), .B(n15589), .Z(n15587) );
  NAND U18363 ( .A(n6993), .B(n15590), .Z(n15588) );
  MUX U18364 ( .IN0(\u_a23_core/u_execute/save_int_pc_m4[29] ), .IN1(n15591), 
        .SEL(\u_a23_core/condition[2] ), .F(n15590) );
  XNOR U18365 ( .A(n7094), .B(n15592), .Z(n15591) );
  AND U18366 ( .A(n15593), .B(n15594), .Z(n15586) );
  NANDN U18367 ( .B(n15595), .A(n15596), .Z(n15594) );
  MUX U18368 ( .IN0(n15597), .IN1(n15598), .SEL(\u_a23_core/condition[2] ), 
        .F(n15595) );
  XOR U18369 ( .A(n7094), .B(n15592), .Z(n15598) );
  IV U18370 ( .A(\u_a23_core/u_execute/save_int_pc_m4[28] ), .Z(n15592) );
  NAND U18371 ( .A(\u_a23_core/u_execute/save_int_pc_m4[29] ), .B(n7272), .Z(
        n15597) );
  NANDN U18372 ( .B(n15599), .A(\u_a23_core/condition[1] ), .Z(n15593) );
  MUX U18373 ( .IN0(n15600), .IN1(n7265), .SEL(\u_a23_core/condition[2] ), .F(
        n15599) );
  XOR U18374 ( .A(n7094), .B(n15601), .Z(n15600) );
  IV U18375 ( .A(\u_a23_core/u_execute/save_int_pc_m4[31] ), .Z(n7094) );
  MUX U18376 ( .IN0(n15602), .IN1(n15603), .SEL(\u_a23_core/condition[2] ), 
        .F(n15584) );
  ANDN U18377 ( .A(n15604), .B(n15605), .Z(n15603) );
  MUX U18378 ( .IN0(n15606), .IN1(n15589), .SEL(
        \u_a23_core/u_execute/save_int_pc_m4[31] ), .F(n15605) );
  AND U18379 ( .A(\u_a23_core/condition[0] ), .B(n7272), .Z(n15606) );
  IV U18380 ( .A(\u_a23_core/condition[1] ), .Z(n7272) );
  NAND U18381 ( .A(\u_a23_core/condition[1] ), .B(n15601), .Z(n15604) );
  XNOR U18382 ( .A(n7265), .B(\u_a23_core/u_execute/save_int_pc_m4[28] ), .Z(
        n15601) );
  ANDN U18383 ( .A(n15607), .B(n15608), .Z(n15602) );
  MUX U18384 ( .IN0(n15596), .IN1(n15609), .SEL(\u_a23_core/condition[1] ), 
        .F(n15608) );
  XOR U18385 ( .A(n9272), .B(n7265), .Z(n15609) );
  IV U18386 ( .A(\u_a23_core/u_execute/save_int_pc_m4[29] ), .Z(n9272) );
  AND U18387 ( .A(n6993), .B(\u_a23_core/condition[0] ), .Z(n15596) );
  IV U18388 ( .A(\u_a23_core/u_execute/save_int_pc_m4[30] ), .Z(n6993) );
  NAND U18389 ( .A(\u_a23_core/u_execute/save_int_pc_m4[30] ), .B(n15589), .Z(
        n15607) );
  ANDN U18390 ( .A(n7265), .B(\u_a23_core/condition[1] ), .Z(n15589) );
  IV U18391 ( .A(\u_a23_core/condition[0] ), .Z(n7265) );
  ANDN U18392 ( .A(n15610), .B(\u_a23_core/address_sel[3] ), .Z(n14158) );
  NAND U18393 ( .A(n14159), .B(\u_a23_core/address_sel[1] ), .Z(n15610) );
  AND U18394 ( .A(n15611), .B(n14162), .Z(n14159) );
  IV U18395 ( .A(\u_a23_core/address_sel[2] ), .Z(n14162) );
  NAND U18396 ( .A(n15612), .B(n15613), .Z(n8407) );
  AND U18397 ( .A(n15611), .B(n15614), .Z(n15613) );
  AND U18398 ( .A(\u_a23_core/address_sel[1] ), .B(\u_a23_core/address_sel[2] ), .Z(n15612) );
  MUX U18399 ( .IN0(n8406), .IN1(n15615), .SEL(\u_a23_core/u_execute/rn[2] ), 
        .F(n14163) );
  NAND U18400 ( .A(n15616), .B(n15617), .Z(\u_a23_core/u_execute/rn[2] ) );
  AND U18401 ( .A(n15618), .B(n15619), .Z(n15617) );
  AND U18402 ( .A(n15620), .B(n15621), .Z(n15619) );
  AND U18403 ( .A(n15622), .B(n15623), .Z(n15621) );
  NANDN U18404 ( .B(n8635), .A(\u_a23_core/u_execute/pc[2] ), .Z(n15623) );
  NAND U18405 ( .A(n15624), .B(n15625), .Z(n8635) );
  NANDN U18406 ( .B(n8636), .A(\u_a23_core/u_execute/u_register_bank/r14[2] ), 
        .Z(n15622) );
  NAND U18407 ( .A(n15625), .B(n15626), .Z(n8636) );
  AND U18408 ( .A(n15627), .B(n15628), .Z(n15620) );
  NANDN U18409 ( .B(n8639), .A(\u_a23_core/u_execute/u_register_bank/r13[2] ), 
        .Z(n15628) );
  NAND U18410 ( .A(n15625), .B(n15629), .Z(n8639) );
  NANDN U18411 ( .B(n8640), .A(\u_a23_core/u_execute/u_register_bank/r12[2] ), 
        .Z(n15627) );
  NAND U18412 ( .A(n15625), .B(n15630), .Z(n8640) );
  AND U18413 ( .A(\u_a23_core/rn_sel[3] ), .B(\u_a23_core/rn_sel[2] ), .Z(
        n15625) );
  AND U18414 ( .A(n15631), .B(n15632), .Z(n15618) );
  AND U18415 ( .A(n15633), .B(n15634), .Z(n15632) );
  NANDN U18416 ( .B(n8645), .A(\u_a23_core/u_execute/u_register_bank/r11[2] ), 
        .Z(n15634) );
  NAND U18417 ( .A(n15635), .B(n15624), .Z(n8645) );
  NANDN U18418 ( .B(n8646), .A(\u_a23_core/u_execute/u_register_bank/r10[2] ), 
        .Z(n15633) );
  NAND U18419 ( .A(n15626), .B(n15635), .Z(n8646) );
  AND U18420 ( .A(n15636), .B(n15637), .Z(n15631) );
  NANDN U18421 ( .B(n8649), .A(\u_a23_core/u_execute/u_register_bank/r9[2] ), 
        .Z(n15637) );
  NAND U18422 ( .A(n15629), .B(n15635), .Z(n8649) );
  NANDN U18423 ( .B(n8650), .A(\u_a23_core/u_execute/u_register_bank/r8[2] ), 
        .Z(n15636) );
  NAND U18424 ( .A(n15630), .B(n15635), .Z(n8650) );
  AND U18425 ( .A(\u_a23_core/rn_sel[3] ), .B(n15638), .Z(n15635) );
  AND U18426 ( .A(n15639), .B(n15640), .Z(n15616) );
  AND U18427 ( .A(n15641), .B(n15642), .Z(n15640) );
  AND U18428 ( .A(n15643), .B(n15644), .Z(n15642) );
  NANDN U18429 ( .B(n8657), .A(\u_a23_core/u_execute/u_register_bank/r7[2] ), 
        .Z(n15644) );
  NAND U18430 ( .A(n15645), .B(n15624), .Z(n8657) );
  NANDN U18431 ( .B(n8658), .A(\u_a23_core/u_execute/u_register_bank/r6[2] ), 
        .Z(n15643) );
  NAND U18432 ( .A(n15626), .B(n15645), .Z(n8658) );
  AND U18433 ( .A(n15646), .B(n15647), .Z(n15641) );
  NANDN U18434 ( .B(n8661), .A(\u_a23_core/u_execute/u_register_bank/r5[2] ), 
        .Z(n15647) );
  NAND U18435 ( .A(n15629), .B(n15645), .Z(n8661) );
  NANDN U18436 ( .B(n8662), .A(\u_a23_core/u_execute/u_register_bank/r4[2] ), 
        .Z(n15646) );
  NAND U18437 ( .A(n15630), .B(n15645), .Z(n8662) );
  NOR U18438 ( .A(n15638), .B(\u_a23_core/rn_sel[3] ), .Z(n15645) );
  IV U18439 ( .A(\u_a23_core/rn_sel[2] ), .Z(n15638) );
  AND U18440 ( .A(n15648), .B(n15649), .Z(n15639) );
  AND U18441 ( .A(n15650), .B(n15651), .Z(n15649) );
  NANDN U18442 ( .B(n8667), .A(\u_a23_core/u_execute/u_register_bank/r3[2] ), 
        .Z(n15651) );
  NAND U18443 ( .A(n15652), .B(n15624), .Z(n8667) );
  ANDN U18444 ( .A(\u_a23_core/rn_sel[0] ), .B(n15653), .Z(n15624) );
  NANDN U18445 ( .B(n8668), .A(\u_a23_core/u_execute/u_register_bank/r0[2] ), 
        .Z(n15650) );
  NAND U18446 ( .A(n15630), .B(n15652), .Z(n8668) );
  ANDN U18447 ( .A(n15654), .B(\u_a23_core/rn_sel[1] ), .Z(n15630) );
  AND U18448 ( .A(n15655), .B(n15656), .Z(n15648) );
  NANDN U18449 ( .B(n8671), .A(\u_a23_core/u_execute/u_register_bank/r2[2] ), 
        .Z(n15656) );
  NAND U18450 ( .A(n15626), .B(n15652), .Z(n8671) );
  ANDN U18451 ( .A(\u_a23_core/rn_sel[1] ), .B(\u_a23_core/rn_sel[0] ), .Z(
        n15626) );
  NANDN U18452 ( .B(n8672), .A(\u_a23_core/u_execute/u_register_bank/r1[2] ), 
        .Z(n15655) );
  NAND U18453 ( .A(n15629), .B(n15652), .Z(n8672) );
  NOR U18454 ( .A(\u_a23_core/rn_sel[2] ), .B(\u_a23_core/rn_sel[3] ), .Z(
        n15652) );
  ANDN U18455 ( .A(n15653), .B(n15654), .Z(n15629) );
  IV U18456 ( .A(\u_a23_core/rn_sel[0] ), .Z(n15654) );
  IV U18457 ( .A(\u_a23_core/rn_sel[1] ), .Z(n15653) );
  IV U18458 ( .A(n8413), .Z(n15615) );
  AND U18459 ( .A(n15657), .B(\u_a23_core/address_sel[2] ), .Z(n8413) );
  AND U18460 ( .A(n14160), .B(n15611), .Z(n15657) );
  IV U18461 ( .A(\u_a23_core/address_sel[0] ), .Z(n15611) );
  NOR U18462 ( .A(\u_a23_core/address_sel[3] ), .B(\u_a23_core/address_sel[1] ), .Z(n14160) );
  NANDN U18463 ( .B(n14157), .A(\u_a23_core/address_sel[2] ), .Z(n8406) );
  NAND U18464 ( .A(n15658), .B(\u_a23_core/address_sel[1] ), .Z(n14157) );
  AND U18465 ( .A(n15614), .B(\u_a23_core/address_sel[0] ), .Z(n15658) );
  IV U18466 ( .A(\u_a23_core/address_sel[3] ), .Z(n15614) );
  IV U18467 ( .A(\u_a23_core/u_execute/rs[10] ), .Z(n16605) );
  NANDN U18468 ( .B(n6060), .A(n15659), .Z(\u_a23_core/u_execute/rs[10] ) );
  NAND U18469 ( .A(\u_a23_core/u_execute/pc[10] ), .B(n6025), .Z(n15659) );
  NAND U18470 ( .A(n15660), .B(n15661), .Z(n6060) );
  AND U18471 ( .A(n15662), .B(n15663), .Z(n15661) );
  AND U18472 ( .A(n15664), .B(n15665), .Z(n15663) );
  AND U18473 ( .A(n15666), .B(n15667), .Z(n15665) );
  NAND U18474 ( .A(\u_a23_core/u_execute/u_register_bank/r14[10] ), .B(n15668), 
        .Z(n15667) );
  NANDN U18475 ( .B(n15669), .A(\u_a23_core/u_execute/u_register_bank/r13[10] ), .Z(n15666) );
  AND U18476 ( .A(n15670), .B(n15671), .Z(n15664) );
  NANDN U18477 ( .B(n15672), .A(\u_a23_core/u_execute/u_register_bank/r12[10] ), .Z(n15671) );
  NANDN U18478 ( .B(n15673), .A(\u_a23_core/u_execute/u_register_bank/r11[10] ), .Z(n15670) );
  AND U18479 ( .A(n15674), .B(n15675), .Z(n15662) );
  AND U18480 ( .A(n15676), .B(n15677), .Z(n15675) );
  NANDN U18481 ( .B(n15678), .A(\u_a23_core/u_execute/u_register_bank/r10[10] ), .Z(n15677) );
  NANDN U18482 ( .B(n15679), .A(\u_a23_core/u_execute/u_register_bank/r9[10] ), 
        .Z(n15676) );
  AND U18483 ( .A(n15680), .B(n15681), .Z(n15674) );
  NANDN U18484 ( .B(n15682), .A(\u_a23_core/u_execute/u_register_bank/r8[10] ), 
        .Z(n15681) );
  NANDN U18485 ( .B(n15683), .A(\u_a23_core/u_execute/u_register_bank/r7[10] ), 
        .Z(n15680) );
  AND U18486 ( .A(n15684), .B(n15685), .Z(n15660) );
  AND U18487 ( .A(n15686), .B(n15687), .Z(n15685) );
  AND U18488 ( .A(n15688), .B(n15689), .Z(n15687) );
  NANDN U18489 ( .B(n15690), .A(\u_a23_core/u_execute/u_register_bank/r6[10] ), 
        .Z(n15689) );
  NANDN U18490 ( .B(n15691), .A(\u_a23_core/u_execute/u_register_bank/r5[10] ), 
        .Z(n15688) );
  AND U18491 ( .A(n15692), .B(n15693), .Z(n15686) );
  NANDN U18492 ( .B(n15694), .A(\u_a23_core/u_execute/u_register_bank/r4[10] ), 
        .Z(n15693) );
  NANDN U18493 ( .B(n15695), .A(\u_a23_core/u_execute/u_register_bank/r3[10] ), 
        .Z(n15692) );
  AND U18494 ( .A(n15696), .B(n15697), .Z(n15684) );
  NANDN U18495 ( .B(n15698), .A(\u_a23_core/u_execute/u_register_bank/r2[10] ), 
        .Z(n15697) );
  AND U18496 ( .A(n15699), .B(n15700), .Z(n15696) );
  NANDN U18497 ( .B(n15701), .A(\u_a23_core/u_execute/u_register_bank/r1[10] ), 
        .Z(n15700) );
  NANDN U18498 ( .B(n15702), .A(\u_a23_core/u_execute/u_register_bank/r0[10] ), 
        .Z(n15699) );
  IV U18499 ( .A(\u_a23_core/u_execute/rs[11] ), .Z(n16606) );
  NANDN U18500 ( .B(n6052), .A(n15703), .Z(\u_a23_core/u_execute/rs[11] ) );
  NAND U18501 ( .A(n6025), .B(\u_a23_core/u_execute/pc[11] ), .Z(n15703) );
  NAND U18502 ( .A(n15704), .B(n15705), .Z(n6052) );
  AND U18503 ( .A(n15706), .B(n15707), .Z(n15705) );
  AND U18504 ( .A(n15708), .B(n15709), .Z(n15707) );
  AND U18505 ( .A(n15710), .B(n15711), .Z(n15709) );
  NAND U18506 ( .A(\u_a23_core/u_execute/u_register_bank/r14[11] ), .B(n15668), 
        .Z(n15711) );
  NANDN U18507 ( .B(n15669), .A(\u_a23_core/u_execute/u_register_bank/r13[11] ), .Z(n15710) );
  AND U18508 ( .A(n15712), .B(n15713), .Z(n15708) );
  NANDN U18509 ( .B(n15672), .A(\u_a23_core/u_execute/u_register_bank/r12[11] ), .Z(n15713) );
  NANDN U18510 ( .B(n15673), .A(\u_a23_core/u_execute/u_register_bank/r11[11] ), .Z(n15712) );
  AND U18511 ( .A(n15714), .B(n15715), .Z(n15706) );
  AND U18512 ( .A(n15716), .B(n15717), .Z(n15715) );
  NANDN U18513 ( .B(n15678), .A(\u_a23_core/u_execute/u_register_bank/r10[11] ), .Z(n15717) );
  NANDN U18514 ( .B(n15679), .A(\u_a23_core/u_execute/u_register_bank/r9[11] ), 
        .Z(n15716) );
  AND U18515 ( .A(n15718), .B(n15719), .Z(n15714) );
  NANDN U18516 ( .B(n15682), .A(\u_a23_core/u_execute/u_register_bank/r8[11] ), 
        .Z(n15719) );
  NANDN U18517 ( .B(n15683), .A(\u_a23_core/u_execute/u_register_bank/r7[11] ), 
        .Z(n15718) );
  AND U18518 ( .A(n15720), .B(n15721), .Z(n15704) );
  AND U18519 ( .A(n15722), .B(n15723), .Z(n15721) );
  AND U18520 ( .A(n15724), .B(n15725), .Z(n15723) );
  NANDN U18521 ( .B(n15690), .A(\u_a23_core/u_execute/u_register_bank/r6[11] ), 
        .Z(n15725) );
  NANDN U18522 ( .B(n15691), .A(\u_a23_core/u_execute/u_register_bank/r5[11] ), 
        .Z(n15724) );
  AND U18523 ( .A(n15726), .B(n15727), .Z(n15722) );
  NANDN U18524 ( .B(n15694), .A(\u_a23_core/u_execute/u_register_bank/r4[11] ), 
        .Z(n15727) );
  NANDN U18525 ( .B(n15695), .A(\u_a23_core/u_execute/u_register_bank/r3[11] ), 
        .Z(n15726) );
  AND U18526 ( .A(n15728), .B(n15729), .Z(n15720) );
  NANDN U18527 ( .B(n15698), .A(\u_a23_core/u_execute/u_register_bank/r2[11] ), 
        .Z(n15729) );
  AND U18528 ( .A(n15730), .B(n15731), .Z(n15728) );
  NANDN U18529 ( .B(n15701), .A(\u_a23_core/u_execute/u_register_bank/r1[11] ), 
        .Z(n15731) );
  NANDN U18530 ( .B(n15702), .A(\u_a23_core/u_execute/u_register_bank/r0[11] ), 
        .Z(n15730) );
  IV U18531 ( .A(\u_a23_core/u_execute/rs[12] ), .Z(n16607) );
  NANDN U18532 ( .B(n6044), .A(n15732), .Z(\u_a23_core/u_execute/rs[12] ) );
  NAND U18533 ( .A(n6025), .B(\u_a23_core/u_execute/pc[12] ), .Z(n15732) );
  NAND U18534 ( .A(n15733), .B(n15734), .Z(n6044) );
  AND U18535 ( .A(n15735), .B(n15736), .Z(n15734) );
  AND U18536 ( .A(n15737), .B(n15738), .Z(n15736) );
  AND U18537 ( .A(n15739), .B(n15740), .Z(n15738) );
  NAND U18538 ( .A(n15668), .B(\u_a23_core/u_execute/u_register_bank/r14[12] ), 
        .Z(n15740) );
  NANDN U18539 ( .B(n15669), .A(\u_a23_core/u_execute/u_register_bank/r13[12] ), .Z(n15739) );
  AND U18540 ( .A(n15741), .B(n15742), .Z(n15737) );
  NANDN U18541 ( .B(n15672), .A(\u_a23_core/u_execute/u_register_bank/r12[12] ), .Z(n15742) );
  NANDN U18542 ( .B(n15673), .A(\u_a23_core/u_execute/u_register_bank/r11[12] ), .Z(n15741) );
  AND U18543 ( .A(n15743), .B(n15744), .Z(n15735) );
  AND U18544 ( .A(n15745), .B(n15746), .Z(n15744) );
  NANDN U18545 ( .B(n15678), .A(\u_a23_core/u_execute/u_register_bank/r10[12] ), .Z(n15746) );
  NANDN U18546 ( .B(n15679), .A(\u_a23_core/u_execute/u_register_bank/r9[12] ), 
        .Z(n15745) );
  AND U18547 ( .A(n15747), .B(n15748), .Z(n15743) );
  NANDN U18548 ( .B(n15682), .A(\u_a23_core/u_execute/u_register_bank/r8[12] ), 
        .Z(n15748) );
  NANDN U18549 ( .B(n15683), .A(\u_a23_core/u_execute/u_register_bank/r7[12] ), 
        .Z(n15747) );
  AND U18550 ( .A(n15749), .B(n15750), .Z(n15733) );
  AND U18551 ( .A(n15751), .B(n15752), .Z(n15750) );
  AND U18552 ( .A(n15753), .B(n15754), .Z(n15752) );
  NANDN U18553 ( .B(n15690), .A(\u_a23_core/u_execute/u_register_bank/r6[12] ), 
        .Z(n15754) );
  NANDN U18554 ( .B(n15691), .A(\u_a23_core/u_execute/u_register_bank/r5[12] ), 
        .Z(n15753) );
  AND U18555 ( .A(n15755), .B(n15756), .Z(n15751) );
  NANDN U18556 ( .B(n15694), .A(\u_a23_core/u_execute/u_register_bank/r4[12] ), 
        .Z(n15756) );
  NANDN U18557 ( .B(n15695), .A(\u_a23_core/u_execute/u_register_bank/r3[12] ), 
        .Z(n15755) );
  AND U18558 ( .A(n15757), .B(n15758), .Z(n15749) );
  NANDN U18559 ( .B(n15698), .A(\u_a23_core/u_execute/u_register_bank/r2[12] ), 
        .Z(n15758) );
  AND U18560 ( .A(n15759), .B(n15760), .Z(n15757) );
  NANDN U18561 ( .B(n15701), .A(\u_a23_core/u_execute/u_register_bank/r1[12] ), 
        .Z(n15760) );
  NANDN U18562 ( .B(n15702), .A(\u_a23_core/u_execute/u_register_bank/r0[12] ), 
        .Z(n15759) );
  IV U18563 ( .A(\u_a23_core/u_execute/rs[13] ), .Z(n16608) );
  NANDN U18564 ( .B(n6036), .A(n15761), .Z(\u_a23_core/u_execute/rs[13] ) );
  NAND U18565 ( .A(n6025), .B(\u_a23_core/u_execute/pc[13] ), .Z(n15761) );
  NAND U18566 ( .A(n15762), .B(n15763), .Z(n6036) );
  AND U18567 ( .A(n15764), .B(n15765), .Z(n15763) );
  AND U18568 ( .A(n15766), .B(n15767), .Z(n15765) );
  AND U18569 ( .A(n15768), .B(n15769), .Z(n15767) );
  NAND U18570 ( .A(n15668), .B(\u_a23_core/u_execute/u_register_bank/r14[13] ), 
        .Z(n15769) );
  NANDN U18571 ( .B(n15669), .A(\u_a23_core/u_execute/u_register_bank/r13[13] ), .Z(n15768) );
  AND U18572 ( .A(n15770), .B(n15771), .Z(n15766) );
  NANDN U18573 ( .B(n15672), .A(\u_a23_core/u_execute/u_register_bank/r12[13] ), .Z(n15771) );
  NANDN U18574 ( .B(n15673), .A(\u_a23_core/u_execute/u_register_bank/r11[13] ), .Z(n15770) );
  AND U18575 ( .A(n15772), .B(n15773), .Z(n15764) );
  AND U18576 ( .A(n15774), .B(n15775), .Z(n15773) );
  NANDN U18577 ( .B(n15678), .A(\u_a23_core/u_execute/u_register_bank/r10[13] ), .Z(n15775) );
  NANDN U18578 ( .B(n15679), .A(\u_a23_core/u_execute/u_register_bank/r9[13] ), 
        .Z(n15774) );
  AND U18579 ( .A(n15776), .B(n15777), .Z(n15772) );
  NANDN U18580 ( .B(n15682), .A(\u_a23_core/u_execute/u_register_bank/r8[13] ), 
        .Z(n15777) );
  NANDN U18581 ( .B(n15683), .A(\u_a23_core/u_execute/u_register_bank/r7[13] ), 
        .Z(n15776) );
  AND U18582 ( .A(n15778), .B(n15779), .Z(n15762) );
  AND U18583 ( .A(n15780), .B(n15781), .Z(n15779) );
  AND U18584 ( .A(n15782), .B(n15783), .Z(n15781) );
  NANDN U18585 ( .B(n15690), .A(\u_a23_core/u_execute/u_register_bank/r6[13] ), 
        .Z(n15783) );
  NANDN U18586 ( .B(n15691), .A(\u_a23_core/u_execute/u_register_bank/r5[13] ), 
        .Z(n15782) );
  AND U18587 ( .A(n15784), .B(n15785), .Z(n15780) );
  NANDN U18588 ( .B(n15694), .A(\u_a23_core/u_execute/u_register_bank/r4[13] ), 
        .Z(n15785) );
  NANDN U18589 ( .B(n15695), .A(\u_a23_core/u_execute/u_register_bank/r3[13] ), 
        .Z(n15784) );
  AND U18590 ( .A(n15786), .B(n15787), .Z(n15778) );
  NANDN U18591 ( .B(n15698), .A(\u_a23_core/u_execute/u_register_bank/r2[13] ), 
        .Z(n15787) );
  AND U18592 ( .A(n15788), .B(n15789), .Z(n15786) );
  NANDN U18593 ( .B(n15701), .A(\u_a23_core/u_execute/u_register_bank/r1[13] ), 
        .Z(n15789) );
  NANDN U18594 ( .B(n15702), .A(\u_a23_core/u_execute/u_register_bank/r0[13] ), 
        .Z(n15788) );
  IV U18595 ( .A(\u_a23_core/u_execute/rs[14] ), .Z(n16609) );
  NANDN U18596 ( .B(n6028), .A(n15790), .Z(\u_a23_core/u_execute/rs[14] ) );
  NAND U18597 ( .A(n6025), .B(\u_a23_core/u_execute/pc[14] ), .Z(n15790) );
  NAND U18598 ( .A(n15791), .B(n15792), .Z(n6028) );
  AND U18599 ( .A(n15793), .B(n15794), .Z(n15792) );
  AND U18600 ( .A(n15795), .B(n15796), .Z(n15794) );
  AND U18601 ( .A(n15797), .B(n15798), .Z(n15796) );
  NAND U18602 ( .A(n15668), .B(\u_a23_core/u_execute/u_register_bank/r14[14] ), 
        .Z(n15798) );
  NANDN U18603 ( .B(n15669), .A(\u_a23_core/u_execute/u_register_bank/r13[14] ), .Z(n15797) );
  AND U18604 ( .A(n15799), .B(n15800), .Z(n15795) );
  NANDN U18605 ( .B(n15672), .A(\u_a23_core/u_execute/u_register_bank/r12[14] ), .Z(n15800) );
  NANDN U18606 ( .B(n15673), .A(\u_a23_core/u_execute/u_register_bank/r11[14] ), .Z(n15799) );
  AND U18607 ( .A(n15801), .B(n15802), .Z(n15793) );
  AND U18608 ( .A(n15803), .B(n15804), .Z(n15802) );
  NANDN U18609 ( .B(n15678), .A(\u_a23_core/u_execute/u_register_bank/r10[14] ), .Z(n15804) );
  NANDN U18610 ( .B(n15679), .A(\u_a23_core/u_execute/u_register_bank/r9[14] ), 
        .Z(n15803) );
  AND U18611 ( .A(n15805), .B(n15806), .Z(n15801) );
  NANDN U18612 ( .B(n15682), .A(\u_a23_core/u_execute/u_register_bank/r8[14] ), 
        .Z(n15806) );
  NANDN U18613 ( .B(n15683), .A(\u_a23_core/u_execute/u_register_bank/r7[14] ), 
        .Z(n15805) );
  AND U18614 ( .A(n15807), .B(n15808), .Z(n15791) );
  AND U18615 ( .A(n15809), .B(n15810), .Z(n15808) );
  AND U18616 ( .A(n15811), .B(n15812), .Z(n15810) );
  NANDN U18617 ( .B(n15690), .A(\u_a23_core/u_execute/u_register_bank/r6[14] ), 
        .Z(n15812) );
  NANDN U18618 ( .B(n15691), .A(\u_a23_core/u_execute/u_register_bank/r5[14] ), 
        .Z(n15811) );
  AND U18619 ( .A(n15813), .B(n15814), .Z(n15809) );
  NANDN U18620 ( .B(n15694), .A(\u_a23_core/u_execute/u_register_bank/r4[14] ), 
        .Z(n15814) );
  NANDN U18621 ( .B(n15695), .A(\u_a23_core/u_execute/u_register_bank/r3[14] ), 
        .Z(n15813) );
  AND U18622 ( .A(n15815), .B(n15816), .Z(n15807) );
  NANDN U18623 ( .B(n15698), .A(\u_a23_core/u_execute/u_register_bank/r2[14] ), 
        .Z(n15816) );
  AND U18624 ( .A(n15817), .B(n15818), .Z(n15815) );
  NANDN U18625 ( .B(n15701), .A(\u_a23_core/u_execute/u_register_bank/r1[14] ), 
        .Z(n15818) );
  NANDN U18626 ( .B(n15702), .A(\u_a23_core/u_execute/u_register_bank/r0[14] ), 
        .Z(n15817) );
  IV U18627 ( .A(\u_a23_core/u_execute/rs[15] ), .Z(n16610) );
  NANDN U18628 ( .B(n6019), .A(n15819), .Z(\u_a23_core/u_execute/rs[15] ) );
  NAND U18629 ( .A(n6025), .B(\u_a23_core/u_execute/pc[15] ), .Z(n15819) );
  NAND U18630 ( .A(n15820), .B(n15821), .Z(n6019) );
  AND U18631 ( .A(n15822), .B(n15823), .Z(n15821) );
  AND U18632 ( .A(n15824), .B(n15825), .Z(n15823) );
  AND U18633 ( .A(n15826), .B(n15827), .Z(n15825) );
  NAND U18634 ( .A(n15668), .B(\u_a23_core/u_execute/u_register_bank/r14[15] ), 
        .Z(n15827) );
  NANDN U18635 ( .B(n15669), .A(\u_a23_core/u_execute/u_register_bank/r13[15] ), .Z(n15826) );
  AND U18636 ( .A(n15828), .B(n15829), .Z(n15824) );
  NANDN U18637 ( .B(n15672), .A(\u_a23_core/u_execute/u_register_bank/r12[15] ), .Z(n15829) );
  NANDN U18638 ( .B(n15673), .A(\u_a23_core/u_execute/u_register_bank/r11[15] ), .Z(n15828) );
  AND U18639 ( .A(n15830), .B(n15831), .Z(n15822) );
  AND U18640 ( .A(n15832), .B(n15833), .Z(n15831) );
  NANDN U18641 ( .B(n15678), .A(\u_a23_core/u_execute/u_register_bank/r10[15] ), .Z(n15833) );
  NANDN U18642 ( .B(n15679), .A(\u_a23_core/u_execute/u_register_bank/r9[15] ), 
        .Z(n15832) );
  AND U18643 ( .A(n15834), .B(n15835), .Z(n15830) );
  NANDN U18644 ( .B(n15682), .A(\u_a23_core/u_execute/u_register_bank/r8[15] ), 
        .Z(n15835) );
  NANDN U18645 ( .B(n15683), .A(\u_a23_core/u_execute/u_register_bank/r7[15] ), 
        .Z(n15834) );
  AND U18646 ( .A(n15836), .B(n15837), .Z(n15820) );
  AND U18647 ( .A(n15838), .B(n15839), .Z(n15837) );
  AND U18648 ( .A(n15840), .B(n15841), .Z(n15839) );
  NANDN U18649 ( .B(n15690), .A(\u_a23_core/u_execute/u_register_bank/r6[15] ), 
        .Z(n15841) );
  NANDN U18650 ( .B(n15691), .A(\u_a23_core/u_execute/u_register_bank/r5[15] ), 
        .Z(n15840) );
  AND U18651 ( .A(n15842), .B(n15843), .Z(n15838) );
  NANDN U18652 ( .B(n15694), .A(\u_a23_core/u_execute/u_register_bank/r4[15] ), 
        .Z(n15843) );
  NANDN U18653 ( .B(n15695), .A(\u_a23_core/u_execute/u_register_bank/r3[15] ), 
        .Z(n15842) );
  AND U18654 ( .A(n15844), .B(n15845), .Z(n15836) );
  NANDN U18655 ( .B(n15698), .A(\u_a23_core/u_execute/u_register_bank/r2[15] ), 
        .Z(n15845) );
  AND U18656 ( .A(n15846), .B(n15847), .Z(n15844) );
  NANDN U18657 ( .B(n15701), .A(\u_a23_core/u_execute/u_register_bank/r1[15] ), 
        .Z(n15847) );
  NANDN U18658 ( .B(n15702), .A(\u_a23_core/u_execute/u_register_bank/r0[15] ), 
        .Z(n15846) );
  IV U18659 ( .A(\u_a23_core/u_execute/rs[16] ), .Z(n16611) );
  NANDN U18660 ( .B(n6014), .A(n15848), .Z(\u_a23_core/u_execute/rs[16] ) );
  NAND U18661 ( .A(n6025), .B(\u_a23_core/u_execute/pc[16] ), .Z(n15848) );
  NAND U18662 ( .A(n15849), .B(n15850), .Z(n6014) );
  AND U18663 ( .A(n15851), .B(n15852), .Z(n15850) );
  AND U18664 ( .A(n15853), .B(n15854), .Z(n15852) );
  AND U18665 ( .A(n15855), .B(n15856), .Z(n15854) );
  NAND U18666 ( .A(n15668), .B(\u_a23_core/u_execute/u_register_bank/r14[16] ), 
        .Z(n15856) );
  NANDN U18667 ( .B(n15669), .A(\u_a23_core/u_execute/u_register_bank/r13[16] ), .Z(n15855) );
  AND U18668 ( .A(n15857), .B(n15858), .Z(n15853) );
  NANDN U18669 ( .B(n15672), .A(\u_a23_core/u_execute/u_register_bank/r12[16] ), .Z(n15858) );
  NANDN U18670 ( .B(n15673), .A(\u_a23_core/u_execute/u_register_bank/r11[16] ), .Z(n15857) );
  AND U18671 ( .A(n15859), .B(n15860), .Z(n15851) );
  AND U18672 ( .A(n15861), .B(n15862), .Z(n15860) );
  NANDN U18673 ( .B(n15678), .A(\u_a23_core/u_execute/u_register_bank/r10[16] ), .Z(n15862) );
  NANDN U18674 ( .B(n15679), .A(\u_a23_core/u_execute/u_register_bank/r9[16] ), 
        .Z(n15861) );
  AND U18675 ( .A(n15863), .B(n15864), .Z(n15859) );
  NANDN U18676 ( .B(n15682), .A(\u_a23_core/u_execute/u_register_bank/r8[16] ), 
        .Z(n15864) );
  NANDN U18677 ( .B(n15683), .A(\u_a23_core/u_execute/u_register_bank/r7[16] ), 
        .Z(n15863) );
  AND U18678 ( .A(n15865), .B(n15866), .Z(n15849) );
  AND U18679 ( .A(n15867), .B(n15868), .Z(n15866) );
  AND U18680 ( .A(n15869), .B(n15870), .Z(n15868) );
  NANDN U18681 ( .B(n15690), .A(\u_a23_core/u_execute/u_register_bank/r6[16] ), 
        .Z(n15870) );
  NANDN U18682 ( .B(n15691), .A(\u_a23_core/u_execute/u_register_bank/r5[16] ), 
        .Z(n15869) );
  AND U18683 ( .A(n15871), .B(n15872), .Z(n15867) );
  NANDN U18684 ( .B(n15694), .A(\u_a23_core/u_execute/u_register_bank/r4[16] ), 
        .Z(n15872) );
  NANDN U18685 ( .B(n15695), .A(\u_a23_core/u_execute/u_register_bank/r3[16] ), 
        .Z(n15871) );
  AND U18686 ( .A(n15873), .B(n15874), .Z(n15865) );
  NANDN U18687 ( .B(n15698), .A(\u_a23_core/u_execute/u_register_bank/r2[16] ), 
        .Z(n15874) );
  AND U18688 ( .A(n15875), .B(n15876), .Z(n15873) );
  NANDN U18689 ( .B(n15701), .A(\u_a23_core/u_execute/u_register_bank/r1[16] ), 
        .Z(n15876) );
  NANDN U18690 ( .B(n15702), .A(\u_a23_core/u_execute/u_register_bank/r0[16] ), 
        .Z(n15875) );
  IV U18691 ( .A(\u_a23_core/u_execute/rs[17] ), .Z(n16612) );
  NANDN U18692 ( .B(n6009), .A(n15877), .Z(\u_a23_core/u_execute/rs[17] ) );
  NAND U18693 ( .A(n6025), .B(\u_a23_core/u_execute/pc[17] ), .Z(n15877) );
  NAND U18694 ( .A(n15878), .B(n15879), .Z(n6009) );
  AND U18695 ( .A(n15880), .B(n15881), .Z(n15879) );
  AND U18696 ( .A(n15882), .B(n15883), .Z(n15881) );
  AND U18697 ( .A(n15884), .B(n15885), .Z(n15883) );
  NAND U18698 ( .A(n15668), .B(\u_a23_core/u_execute/u_register_bank/r14[17] ), 
        .Z(n15885) );
  NANDN U18699 ( .B(n15669), .A(\u_a23_core/u_execute/u_register_bank/r13[17] ), .Z(n15884) );
  AND U18700 ( .A(n15886), .B(n15887), .Z(n15882) );
  NANDN U18701 ( .B(n15672), .A(\u_a23_core/u_execute/u_register_bank/r12[17] ), .Z(n15887) );
  NANDN U18702 ( .B(n15673), .A(\u_a23_core/u_execute/u_register_bank/r11[17] ), .Z(n15886) );
  AND U18703 ( .A(n15888), .B(n15889), .Z(n15880) );
  AND U18704 ( .A(n15890), .B(n15891), .Z(n15889) );
  NANDN U18705 ( .B(n15678), .A(\u_a23_core/u_execute/u_register_bank/r10[17] ), .Z(n15891) );
  NANDN U18706 ( .B(n15679), .A(\u_a23_core/u_execute/u_register_bank/r9[17] ), 
        .Z(n15890) );
  AND U18707 ( .A(n15892), .B(n15893), .Z(n15888) );
  NANDN U18708 ( .B(n15682), .A(\u_a23_core/u_execute/u_register_bank/r8[17] ), 
        .Z(n15893) );
  NANDN U18709 ( .B(n15683), .A(\u_a23_core/u_execute/u_register_bank/r7[17] ), 
        .Z(n15892) );
  AND U18710 ( .A(n15894), .B(n15895), .Z(n15878) );
  AND U18711 ( .A(n15896), .B(n15897), .Z(n15895) );
  AND U18712 ( .A(n15898), .B(n15899), .Z(n15897) );
  NANDN U18713 ( .B(n15690), .A(\u_a23_core/u_execute/u_register_bank/r6[17] ), 
        .Z(n15899) );
  NANDN U18714 ( .B(n15691), .A(\u_a23_core/u_execute/u_register_bank/r5[17] ), 
        .Z(n15898) );
  AND U18715 ( .A(n15900), .B(n15901), .Z(n15896) );
  NANDN U18716 ( .B(n15694), .A(\u_a23_core/u_execute/u_register_bank/r4[17] ), 
        .Z(n15901) );
  NANDN U18717 ( .B(n15695), .A(\u_a23_core/u_execute/u_register_bank/r3[17] ), 
        .Z(n15900) );
  AND U18718 ( .A(n15902), .B(n15903), .Z(n15894) );
  NANDN U18719 ( .B(n15698), .A(\u_a23_core/u_execute/u_register_bank/r2[17] ), 
        .Z(n15903) );
  AND U18720 ( .A(n15904), .B(n15905), .Z(n15902) );
  NANDN U18721 ( .B(n15701), .A(\u_a23_core/u_execute/u_register_bank/r1[17] ), 
        .Z(n15905) );
  NANDN U18722 ( .B(n15702), .A(\u_a23_core/u_execute/u_register_bank/r0[17] ), 
        .Z(n15904) );
  IV U18723 ( .A(\u_a23_core/u_execute/rs[18] ), .Z(n16613) );
  NANDN U18724 ( .B(n6004), .A(n15906), .Z(\u_a23_core/u_execute/rs[18] ) );
  NAND U18725 ( .A(n6025), .B(\u_a23_core/u_execute/pc[18] ), .Z(n15906) );
  NAND U18726 ( .A(n15907), .B(n15908), .Z(n6004) );
  AND U18727 ( .A(n15909), .B(n15910), .Z(n15908) );
  AND U18728 ( .A(n15911), .B(n15912), .Z(n15910) );
  AND U18729 ( .A(n15913), .B(n15914), .Z(n15912) );
  NAND U18730 ( .A(n15668), .B(\u_a23_core/u_execute/u_register_bank/r14[18] ), 
        .Z(n15914) );
  NANDN U18731 ( .B(n15669), .A(\u_a23_core/u_execute/u_register_bank/r13[18] ), .Z(n15913) );
  AND U18732 ( .A(n15915), .B(n15916), .Z(n15911) );
  NANDN U18733 ( .B(n15672), .A(\u_a23_core/u_execute/u_register_bank/r12[18] ), .Z(n15916) );
  NANDN U18734 ( .B(n15673), .A(\u_a23_core/u_execute/u_register_bank/r11[18] ), .Z(n15915) );
  AND U18735 ( .A(n15917), .B(n15918), .Z(n15909) );
  AND U18736 ( .A(n15919), .B(n15920), .Z(n15918) );
  NANDN U18737 ( .B(n15678), .A(\u_a23_core/u_execute/u_register_bank/r10[18] ), .Z(n15920) );
  NANDN U18738 ( .B(n15679), .A(\u_a23_core/u_execute/u_register_bank/r9[18] ), 
        .Z(n15919) );
  AND U18739 ( .A(n15921), .B(n15922), .Z(n15917) );
  NANDN U18740 ( .B(n15682), .A(\u_a23_core/u_execute/u_register_bank/r8[18] ), 
        .Z(n15922) );
  NANDN U18741 ( .B(n15683), .A(\u_a23_core/u_execute/u_register_bank/r7[18] ), 
        .Z(n15921) );
  AND U18742 ( .A(n15923), .B(n15924), .Z(n15907) );
  AND U18743 ( .A(n15925), .B(n15926), .Z(n15924) );
  AND U18744 ( .A(n15927), .B(n15928), .Z(n15926) );
  NANDN U18745 ( .B(n15690), .A(\u_a23_core/u_execute/u_register_bank/r6[18] ), 
        .Z(n15928) );
  NANDN U18746 ( .B(n15691), .A(\u_a23_core/u_execute/u_register_bank/r5[18] ), 
        .Z(n15927) );
  AND U18747 ( .A(n15929), .B(n15930), .Z(n15925) );
  NANDN U18748 ( .B(n15694), .A(\u_a23_core/u_execute/u_register_bank/r4[18] ), 
        .Z(n15930) );
  NANDN U18749 ( .B(n15695), .A(\u_a23_core/u_execute/u_register_bank/r3[18] ), 
        .Z(n15929) );
  AND U18750 ( .A(n15931), .B(n15932), .Z(n15923) );
  NANDN U18751 ( .B(n15698), .A(\u_a23_core/u_execute/u_register_bank/r2[18] ), 
        .Z(n15932) );
  AND U18752 ( .A(n15933), .B(n15934), .Z(n15931) );
  NANDN U18753 ( .B(n15701), .A(\u_a23_core/u_execute/u_register_bank/r1[18] ), 
        .Z(n15934) );
  NANDN U18754 ( .B(n15702), .A(\u_a23_core/u_execute/u_register_bank/r0[18] ), 
        .Z(n15933) );
  IV U18755 ( .A(\u_a23_core/u_execute/rs[19] ), .Z(n16614) );
  NANDN U18756 ( .B(n5999), .A(n15935), .Z(\u_a23_core/u_execute/rs[19] ) );
  NAND U18757 ( .A(n6025), .B(\u_a23_core/u_execute/pc[19] ), .Z(n15935) );
  NAND U18758 ( .A(n15936), .B(n15937), .Z(n5999) );
  AND U18759 ( .A(n15938), .B(n15939), .Z(n15937) );
  AND U18760 ( .A(n15940), .B(n15941), .Z(n15939) );
  AND U18761 ( .A(n15942), .B(n15943), .Z(n15941) );
  NAND U18762 ( .A(n15668), .B(\u_a23_core/u_execute/u_register_bank/r14[19] ), 
        .Z(n15943) );
  NANDN U18763 ( .B(n15669), .A(\u_a23_core/u_execute/u_register_bank/r13[19] ), .Z(n15942) );
  AND U18764 ( .A(n15944), .B(n15945), .Z(n15940) );
  NANDN U18765 ( .B(n15672), .A(\u_a23_core/u_execute/u_register_bank/r12[19] ), .Z(n15945) );
  NANDN U18766 ( .B(n15673), .A(\u_a23_core/u_execute/u_register_bank/r11[19] ), .Z(n15944) );
  AND U18767 ( .A(n15946), .B(n15947), .Z(n15938) );
  AND U18768 ( .A(n15948), .B(n15949), .Z(n15947) );
  NANDN U18769 ( .B(n15678), .A(\u_a23_core/u_execute/u_register_bank/r10[19] ), .Z(n15949) );
  NANDN U18770 ( .B(n15679), .A(\u_a23_core/u_execute/u_register_bank/r9[19] ), 
        .Z(n15948) );
  AND U18771 ( .A(n15950), .B(n15951), .Z(n15946) );
  NANDN U18772 ( .B(n15682), .A(\u_a23_core/u_execute/u_register_bank/r8[19] ), 
        .Z(n15951) );
  NANDN U18773 ( .B(n15683), .A(\u_a23_core/u_execute/u_register_bank/r7[19] ), 
        .Z(n15950) );
  AND U18774 ( .A(n15952), .B(n15953), .Z(n15936) );
  AND U18775 ( .A(n15954), .B(n15955), .Z(n15953) );
  AND U18776 ( .A(n15956), .B(n15957), .Z(n15955) );
  NANDN U18777 ( .B(n15690), .A(\u_a23_core/u_execute/u_register_bank/r6[19] ), 
        .Z(n15957) );
  NANDN U18778 ( .B(n15691), .A(\u_a23_core/u_execute/u_register_bank/r5[19] ), 
        .Z(n15956) );
  AND U18779 ( .A(n15958), .B(n15959), .Z(n15954) );
  NANDN U18780 ( .B(n15694), .A(\u_a23_core/u_execute/u_register_bank/r4[19] ), 
        .Z(n15959) );
  NANDN U18781 ( .B(n15695), .A(\u_a23_core/u_execute/u_register_bank/r3[19] ), 
        .Z(n15958) );
  AND U18782 ( .A(n15960), .B(n15961), .Z(n15952) );
  NANDN U18783 ( .B(n15698), .A(\u_a23_core/u_execute/u_register_bank/r2[19] ), 
        .Z(n15961) );
  AND U18784 ( .A(n15962), .B(n15963), .Z(n15960) );
  NANDN U18785 ( .B(n15701), .A(\u_a23_core/u_execute/u_register_bank/r1[19] ), 
        .Z(n15963) );
  NANDN U18786 ( .B(n15702), .A(\u_a23_core/u_execute/u_register_bank/r0[19] ), 
        .Z(n15962) );
  IV U18787 ( .A(\u_a23_core/u_execute/rs[20] ), .Z(n16615) );
  NANDN U18788 ( .B(n5994), .A(n15964), .Z(\u_a23_core/u_execute/rs[20] ) );
  NAND U18789 ( .A(n6025), .B(\u_a23_core/u_execute/pc[20] ), .Z(n15964) );
  NAND U18790 ( .A(n15965), .B(n15966), .Z(n5994) );
  AND U18791 ( .A(n15967), .B(n15968), .Z(n15966) );
  AND U18792 ( .A(n15969), .B(n15970), .Z(n15968) );
  AND U18793 ( .A(n15971), .B(n15972), .Z(n15970) );
  NAND U18794 ( .A(n15668), .B(\u_a23_core/u_execute/u_register_bank/r14[20] ), 
        .Z(n15972) );
  NANDN U18795 ( .B(n15669), .A(\u_a23_core/u_execute/u_register_bank/r13[20] ), .Z(n15971) );
  AND U18796 ( .A(n15973), .B(n15974), .Z(n15969) );
  NANDN U18797 ( .B(n15672), .A(\u_a23_core/u_execute/u_register_bank/r12[20] ), .Z(n15974) );
  NANDN U18798 ( .B(n15673), .A(\u_a23_core/u_execute/u_register_bank/r11[20] ), .Z(n15973) );
  AND U18799 ( .A(n15975), .B(n15976), .Z(n15967) );
  AND U18800 ( .A(n15977), .B(n15978), .Z(n15976) );
  NANDN U18801 ( .B(n15678), .A(\u_a23_core/u_execute/u_register_bank/r10[20] ), .Z(n15978) );
  NANDN U18802 ( .B(n15679), .A(\u_a23_core/u_execute/u_register_bank/r9[20] ), 
        .Z(n15977) );
  AND U18803 ( .A(n15979), .B(n15980), .Z(n15975) );
  NANDN U18804 ( .B(n15682), .A(\u_a23_core/u_execute/u_register_bank/r8[20] ), 
        .Z(n15980) );
  NANDN U18805 ( .B(n15683), .A(\u_a23_core/u_execute/u_register_bank/r7[20] ), 
        .Z(n15979) );
  AND U18806 ( .A(n15981), .B(n15982), .Z(n15965) );
  AND U18807 ( .A(n15983), .B(n15984), .Z(n15982) );
  AND U18808 ( .A(n15985), .B(n15986), .Z(n15984) );
  NANDN U18809 ( .B(n15690), .A(\u_a23_core/u_execute/u_register_bank/r6[20] ), 
        .Z(n15986) );
  NANDN U18810 ( .B(n15691), .A(\u_a23_core/u_execute/u_register_bank/r5[20] ), 
        .Z(n15985) );
  AND U18811 ( .A(n15987), .B(n15988), .Z(n15983) );
  NANDN U18812 ( .B(n15694), .A(\u_a23_core/u_execute/u_register_bank/r4[20] ), 
        .Z(n15988) );
  NANDN U18813 ( .B(n15695), .A(\u_a23_core/u_execute/u_register_bank/r3[20] ), 
        .Z(n15987) );
  AND U18814 ( .A(n15989), .B(n15990), .Z(n15981) );
  NANDN U18815 ( .B(n15698), .A(\u_a23_core/u_execute/u_register_bank/r2[20] ), 
        .Z(n15990) );
  AND U18816 ( .A(n15991), .B(n15992), .Z(n15989) );
  NANDN U18817 ( .B(n15701), .A(\u_a23_core/u_execute/u_register_bank/r1[20] ), 
        .Z(n15992) );
  NANDN U18818 ( .B(n15702), .A(\u_a23_core/u_execute/u_register_bank/r0[20] ), 
        .Z(n15991) );
  IV U18819 ( .A(\u_a23_core/u_execute/rs[21] ), .Z(n16616) );
  NANDN U18820 ( .B(n5989), .A(n15993), .Z(\u_a23_core/u_execute/rs[21] ) );
  NAND U18821 ( .A(n6025), .B(\u_a23_core/u_execute/pc[21] ), .Z(n15993) );
  NAND U18822 ( .A(n15994), .B(n15995), .Z(n5989) );
  AND U18823 ( .A(n15996), .B(n15997), .Z(n15995) );
  AND U18824 ( .A(n15998), .B(n15999), .Z(n15997) );
  AND U18825 ( .A(n16000), .B(n16001), .Z(n15999) );
  NAND U18826 ( .A(n15668), .B(\u_a23_core/u_execute/u_register_bank/r14[21] ), 
        .Z(n16001) );
  NANDN U18827 ( .B(n15669), .A(\u_a23_core/u_execute/u_register_bank/r13[21] ), .Z(n16000) );
  AND U18828 ( .A(n16002), .B(n16003), .Z(n15998) );
  NANDN U18829 ( .B(n15672), .A(\u_a23_core/u_execute/u_register_bank/r12[21] ), .Z(n16003) );
  NANDN U18830 ( .B(n15673), .A(\u_a23_core/u_execute/u_register_bank/r11[21] ), .Z(n16002) );
  AND U18831 ( .A(n16004), .B(n16005), .Z(n15996) );
  AND U18832 ( .A(n16006), .B(n16007), .Z(n16005) );
  NANDN U18833 ( .B(n15678), .A(\u_a23_core/u_execute/u_register_bank/r10[21] ), .Z(n16007) );
  NANDN U18834 ( .B(n15679), .A(\u_a23_core/u_execute/u_register_bank/r9[21] ), 
        .Z(n16006) );
  AND U18835 ( .A(n16008), .B(n16009), .Z(n16004) );
  NANDN U18836 ( .B(n15682), .A(\u_a23_core/u_execute/u_register_bank/r8[21] ), 
        .Z(n16009) );
  NANDN U18837 ( .B(n15683), .A(\u_a23_core/u_execute/u_register_bank/r7[21] ), 
        .Z(n16008) );
  AND U18838 ( .A(n16010), .B(n16011), .Z(n15994) );
  AND U18839 ( .A(n16012), .B(n16013), .Z(n16011) );
  AND U18840 ( .A(n16014), .B(n16015), .Z(n16013) );
  NANDN U18841 ( .B(n15690), .A(\u_a23_core/u_execute/u_register_bank/r6[21] ), 
        .Z(n16015) );
  NANDN U18842 ( .B(n15691), .A(\u_a23_core/u_execute/u_register_bank/r5[21] ), 
        .Z(n16014) );
  AND U18843 ( .A(n16016), .B(n16017), .Z(n16012) );
  NANDN U18844 ( .B(n15694), .A(\u_a23_core/u_execute/u_register_bank/r4[21] ), 
        .Z(n16017) );
  NANDN U18845 ( .B(n15695), .A(\u_a23_core/u_execute/u_register_bank/r3[21] ), 
        .Z(n16016) );
  AND U18846 ( .A(n16018), .B(n16019), .Z(n16010) );
  NANDN U18847 ( .B(n15698), .A(\u_a23_core/u_execute/u_register_bank/r2[21] ), 
        .Z(n16019) );
  AND U18848 ( .A(n16020), .B(n16021), .Z(n16018) );
  NANDN U18849 ( .B(n15701), .A(\u_a23_core/u_execute/u_register_bank/r1[21] ), 
        .Z(n16021) );
  NANDN U18850 ( .B(n15702), .A(\u_a23_core/u_execute/u_register_bank/r0[21] ), 
        .Z(n16020) );
  IV U18851 ( .A(\u_a23_core/u_execute/rs[22] ), .Z(n16617) );
  NANDN U18852 ( .B(n5984), .A(n16022), .Z(\u_a23_core/u_execute/rs[22] ) );
  NAND U18853 ( .A(n6025), .B(\u_a23_core/u_execute/pc[22] ), .Z(n16022) );
  NAND U18854 ( .A(n16023), .B(n16024), .Z(n5984) );
  AND U18855 ( .A(n16025), .B(n16026), .Z(n16024) );
  AND U18856 ( .A(n16027), .B(n16028), .Z(n16026) );
  AND U18857 ( .A(n16029), .B(n16030), .Z(n16028) );
  NAND U18858 ( .A(n15668), .B(\u_a23_core/u_execute/u_register_bank/r14[22] ), 
        .Z(n16030) );
  NANDN U18859 ( .B(n15669), .A(\u_a23_core/u_execute/u_register_bank/r13[22] ), .Z(n16029) );
  AND U18860 ( .A(n16031), .B(n16032), .Z(n16027) );
  NANDN U18861 ( .B(n15672), .A(\u_a23_core/u_execute/u_register_bank/r12[22] ), .Z(n16032) );
  NANDN U18862 ( .B(n15673), .A(\u_a23_core/u_execute/u_register_bank/r11[22] ), .Z(n16031) );
  AND U18863 ( .A(n16033), .B(n16034), .Z(n16025) );
  AND U18864 ( .A(n16035), .B(n16036), .Z(n16034) );
  NANDN U18865 ( .B(n15678), .A(\u_a23_core/u_execute/u_register_bank/r10[22] ), .Z(n16036) );
  NANDN U18866 ( .B(n15679), .A(\u_a23_core/u_execute/u_register_bank/r9[22] ), 
        .Z(n16035) );
  AND U18867 ( .A(n16037), .B(n16038), .Z(n16033) );
  NANDN U18868 ( .B(n15682), .A(\u_a23_core/u_execute/u_register_bank/r8[22] ), 
        .Z(n16038) );
  NANDN U18869 ( .B(n15683), .A(\u_a23_core/u_execute/u_register_bank/r7[22] ), 
        .Z(n16037) );
  AND U18870 ( .A(n16039), .B(n16040), .Z(n16023) );
  AND U18871 ( .A(n16041), .B(n16042), .Z(n16040) );
  AND U18872 ( .A(n16043), .B(n16044), .Z(n16042) );
  NANDN U18873 ( .B(n15690), .A(\u_a23_core/u_execute/u_register_bank/r6[22] ), 
        .Z(n16044) );
  NANDN U18874 ( .B(n15691), .A(\u_a23_core/u_execute/u_register_bank/r5[22] ), 
        .Z(n16043) );
  AND U18875 ( .A(n16045), .B(n16046), .Z(n16041) );
  NANDN U18876 ( .B(n15694), .A(\u_a23_core/u_execute/u_register_bank/r4[22] ), 
        .Z(n16046) );
  NANDN U18877 ( .B(n15695), .A(\u_a23_core/u_execute/u_register_bank/r3[22] ), 
        .Z(n16045) );
  AND U18878 ( .A(n16047), .B(n16048), .Z(n16039) );
  NANDN U18879 ( .B(n15698), .A(\u_a23_core/u_execute/u_register_bank/r2[22] ), 
        .Z(n16048) );
  AND U18880 ( .A(n16049), .B(n16050), .Z(n16047) );
  NANDN U18881 ( .B(n15701), .A(\u_a23_core/u_execute/u_register_bank/r1[22] ), 
        .Z(n16050) );
  NANDN U18882 ( .B(n15702), .A(\u_a23_core/u_execute/u_register_bank/r0[22] ), 
        .Z(n16049) );
  IV U18883 ( .A(\u_a23_core/u_execute/rs[23] ), .Z(n16618) );
  NANDN U18884 ( .B(n5979), .A(n16051), .Z(\u_a23_core/u_execute/rs[23] ) );
  NAND U18885 ( .A(n6025), .B(\u_a23_core/u_execute/pc[23] ), .Z(n16051) );
  NAND U18886 ( .A(n16052), .B(n16053), .Z(n5979) );
  AND U18887 ( .A(n16054), .B(n16055), .Z(n16053) );
  AND U18888 ( .A(n16056), .B(n16057), .Z(n16055) );
  AND U18889 ( .A(n16058), .B(n16059), .Z(n16057) );
  NAND U18890 ( .A(n15668), .B(\u_a23_core/u_execute/u_register_bank/r14[23] ), 
        .Z(n16059) );
  NANDN U18891 ( .B(n15669), .A(\u_a23_core/u_execute/u_register_bank/r13[23] ), .Z(n16058) );
  AND U18892 ( .A(n16060), .B(n16061), .Z(n16056) );
  NANDN U18893 ( .B(n15672), .A(\u_a23_core/u_execute/u_register_bank/r12[23] ), .Z(n16061) );
  NANDN U18894 ( .B(n15673), .A(\u_a23_core/u_execute/u_register_bank/r11[23] ), .Z(n16060) );
  AND U18895 ( .A(n16062), .B(n16063), .Z(n16054) );
  AND U18896 ( .A(n16064), .B(n16065), .Z(n16063) );
  NANDN U18897 ( .B(n15678), .A(\u_a23_core/u_execute/u_register_bank/r10[23] ), .Z(n16065) );
  NANDN U18898 ( .B(n15679), .A(\u_a23_core/u_execute/u_register_bank/r9[23] ), 
        .Z(n16064) );
  AND U18899 ( .A(n16066), .B(n16067), .Z(n16062) );
  NANDN U18900 ( .B(n15682), .A(\u_a23_core/u_execute/u_register_bank/r8[23] ), 
        .Z(n16067) );
  NANDN U18901 ( .B(n15683), .A(\u_a23_core/u_execute/u_register_bank/r7[23] ), 
        .Z(n16066) );
  AND U18902 ( .A(n16068), .B(n16069), .Z(n16052) );
  AND U18903 ( .A(n16070), .B(n16071), .Z(n16069) );
  AND U18904 ( .A(n16072), .B(n16073), .Z(n16071) );
  NANDN U18905 ( .B(n15690), .A(\u_a23_core/u_execute/u_register_bank/r6[23] ), 
        .Z(n16073) );
  NANDN U18906 ( .B(n15691), .A(\u_a23_core/u_execute/u_register_bank/r5[23] ), 
        .Z(n16072) );
  AND U18907 ( .A(n16074), .B(n16075), .Z(n16070) );
  NANDN U18908 ( .B(n15694), .A(\u_a23_core/u_execute/u_register_bank/r4[23] ), 
        .Z(n16075) );
  NANDN U18909 ( .B(n15695), .A(\u_a23_core/u_execute/u_register_bank/r3[23] ), 
        .Z(n16074) );
  AND U18910 ( .A(n16076), .B(n16077), .Z(n16068) );
  NANDN U18911 ( .B(n15698), .A(\u_a23_core/u_execute/u_register_bank/r2[23] ), 
        .Z(n16077) );
  AND U18912 ( .A(n16078), .B(n16079), .Z(n16076) );
  NANDN U18913 ( .B(n15701), .A(\u_a23_core/u_execute/u_register_bank/r1[23] ), 
        .Z(n16079) );
  NANDN U18914 ( .B(n15702), .A(\u_a23_core/u_execute/u_register_bank/r0[23] ), 
        .Z(n16078) );
  IV U18915 ( .A(\u_a23_core/u_execute/rs[24] ), .Z(n16619) );
  NANDN U18916 ( .B(n5974), .A(n16080), .Z(\u_a23_core/u_execute/rs[24] ) );
  NAND U18917 ( .A(n6025), .B(\u_a23_core/u_execute/pc[24] ), .Z(n16080) );
  NAND U18918 ( .A(n16081), .B(n16082), .Z(n5974) );
  AND U18919 ( .A(n16083), .B(n16084), .Z(n16082) );
  AND U18920 ( .A(n16085), .B(n16086), .Z(n16084) );
  AND U18921 ( .A(n16087), .B(n16088), .Z(n16086) );
  NAND U18922 ( .A(n15668), .B(\u_a23_core/u_execute/u_register_bank/r14[24] ), 
        .Z(n16088) );
  NANDN U18923 ( .B(n15669), .A(\u_a23_core/u_execute/u_register_bank/r13[24] ), .Z(n16087) );
  AND U18924 ( .A(n16089), .B(n16090), .Z(n16085) );
  NANDN U18925 ( .B(n15672), .A(\u_a23_core/u_execute/u_register_bank/r12[24] ), .Z(n16090) );
  NANDN U18926 ( .B(n15673), .A(\u_a23_core/u_execute/u_register_bank/r11[24] ), .Z(n16089) );
  AND U18927 ( .A(n16091), .B(n16092), .Z(n16083) );
  AND U18928 ( .A(n16093), .B(n16094), .Z(n16092) );
  NANDN U18929 ( .B(n15678), .A(\u_a23_core/u_execute/u_register_bank/r10[24] ), .Z(n16094) );
  NANDN U18930 ( .B(n15679), .A(\u_a23_core/u_execute/u_register_bank/r9[24] ), 
        .Z(n16093) );
  AND U18931 ( .A(n16095), .B(n16096), .Z(n16091) );
  NANDN U18932 ( .B(n15682), .A(\u_a23_core/u_execute/u_register_bank/r8[24] ), 
        .Z(n16096) );
  NANDN U18933 ( .B(n15683), .A(\u_a23_core/u_execute/u_register_bank/r7[24] ), 
        .Z(n16095) );
  AND U18934 ( .A(n16097), .B(n16098), .Z(n16081) );
  AND U18935 ( .A(n16099), .B(n16100), .Z(n16098) );
  AND U18936 ( .A(n16101), .B(n16102), .Z(n16100) );
  NANDN U18937 ( .B(n15690), .A(\u_a23_core/u_execute/u_register_bank/r6[24] ), 
        .Z(n16102) );
  NANDN U18938 ( .B(n15691), .A(\u_a23_core/u_execute/u_register_bank/r5[24] ), 
        .Z(n16101) );
  AND U18939 ( .A(n16103), .B(n16104), .Z(n16099) );
  NANDN U18940 ( .B(n15694), .A(\u_a23_core/u_execute/u_register_bank/r4[24] ), 
        .Z(n16104) );
  NANDN U18941 ( .B(n15695), .A(\u_a23_core/u_execute/u_register_bank/r3[24] ), 
        .Z(n16103) );
  AND U18942 ( .A(n16105), .B(n16106), .Z(n16097) );
  NANDN U18943 ( .B(n15698), .A(\u_a23_core/u_execute/u_register_bank/r2[24] ), 
        .Z(n16106) );
  AND U18944 ( .A(n16107), .B(n16108), .Z(n16105) );
  NANDN U18945 ( .B(n15701), .A(\u_a23_core/u_execute/u_register_bank/r1[24] ), 
        .Z(n16108) );
  NANDN U18946 ( .B(n15702), .A(\u_a23_core/u_execute/u_register_bank/r0[24] ), 
        .Z(n16107) );
  IV U18947 ( .A(\u_a23_core/u_execute/rs[25] ), .Z(n16620) );
  NANDN U18948 ( .B(n5969), .A(n16109), .Z(\u_a23_core/u_execute/rs[25] ) );
  NAND U18949 ( .A(n6025), .B(\u_a23_core/u_execute/pc[25] ), .Z(n16109) );
  NAND U18950 ( .A(n16110), .B(n16111), .Z(n5969) );
  AND U18951 ( .A(n16112), .B(n16113), .Z(n16111) );
  AND U18952 ( .A(n16114), .B(n16115), .Z(n16113) );
  AND U18953 ( .A(n16116), .B(n16117), .Z(n16115) );
  NAND U18954 ( .A(n15668), .B(\u_a23_core/u_execute/u_register_bank/r14[25] ), 
        .Z(n16117) );
  NANDN U18955 ( .B(n15669), .A(\u_a23_core/u_execute/u_register_bank/r13[25] ), .Z(n16116) );
  AND U18956 ( .A(n16118), .B(n16119), .Z(n16114) );
  NANDN U18957 ( .B(n15672), .A(\u_a23_core/u_execute/u_register_bank/r12[25] ), .Z(n16119) );
  NANDN U18958 ( .B(n15673), .A(\u_a23_core/u_execute/u_register_bank/r11[25] ), .Z(n16118) );
  AND U18959 ( .A(n16120), .B(n16121), .Z(n16112) );
  AND U18960 ( .A(n16122), .B(n16123), .Z(n16121) );
  NANDN U18961 ( .B(n15678), .A(\u_a23_core/u_execute/u_register_bank/r10[25] ), .Z(n16123) );
  NANDN U18962 ( .B(n15679), .A(\u_a23_core/u_execute/u_register_bank/r9[25] ), 
        .Z(n16122) );
  AND U18963 ( .A(n16124), .B(n16125), .Z(n16120) );
  NANDN U18964 ( .B(n15682), .A(\u_a23_core/u_execute/u_register_bank/r8[25] ), 
        .Z(n16125) );
  NANDN U18965 ( .B(n15683), .A(\u_a23_core/u_execute/u_register_bank/r7[25] ), 
        .Z(n16124) );
  AND U18966 ( .A(n16126), .B(n16127), .Z(n16110) );
  AND U18967 ( .A(n16128), .B(n16129), .Z(n16127) );
  AND U18968 ( .A(n16130), .B(n16131), .Z(n16129) );
  NANDN U18969 ( .B(n15690), .A(\u_a23_core/u_execute/u_register_bank/r6[25] ), 
        .Z(n16131) );
  NANDN U18970 ( .B(n15691), .A(\u_a23_core/u_execute/u_register_bank/r5[25] ), 
        .Z(n16130) );
  AND U18971 ( .A(n16132), .B(n16133), .Z(n16128) );
  NANDN U18972 ( .B(n15694), .A(\u_a23_core/u_execute/u_register_bank/r4[25] ), 
        .Z(n16133) );
  NANDN U18973 ( .B(n15695), .A(\u_a23_core/u_execute/u_register_bank/r3[25] ), 
        .Z(n16132) );
  AND U18974 ( .A(n16134), .B(n16135), .Z(n16126) );
  NANDN U18975 ( .B(n15698), .A(\u_a23_core/u_execute/u_register_bank/r2[25] ), 
        .Z(n16135) );
  AND U18976 ( .A(n16136), .B(n16137), .Z(n16134) );
  NANDN U18977 ( .B(n15701), .A(\u_a23_core/u_execute/u_register_bank/r1[25] ), 
        .Z(n16137) );
  NANDN U18978 ( .B(n15702), .A(\u_a23_core/u_execute/u_register_bank/r0[25] ), 
        .Z(n16136) );
  IV U18979 ( .A(\u_a23_core/u_execute/rs[26] ), .Z(n16621) );
  NAND U18980 ( .A(n16138), .B(n16139), .Z(\u_a23_core/u_execute/rs[26] ) );
  AND U18981 ( .A(n16140), .B(n16141), .Z(n16139) );
  AND U18982 ( .A(n16142), .B(n16143), .Z(n16141) );
  AND U18983 ( .A(n16144), .B(n16145), .Z(n16143) );
  NAND U18984 ( .A(n15668), .B(\u_a23_core/u_execute/u_register_bank/r14[26] ), 
        .Z(n16145) );
  NANDN U18985 ( .B(n15669), .A(\u_a23_core/u_execute/u_register_bank/r13[26] ), .Z(n16144) );
  AND U18986 ( .A(n16146), .B(n16147), .Z(n16142) );
  NANDN U18987 ( .B(n15672), .A(\u_a23_core/u_execute/u_register_bank/r12[26] ), .Z(n16147) );
  NANDN U18988 ( .B(n15673), .A(\u_a23_core/u_execute/u_register_bank/r11[26] ), .Z(n16146) );
  AND U18989 ( .A(n16148), .B(n16149), .Z(n16140) );
  AND U18990 ( .A(n16150), .B(n16151), .Z(n16149) );
  NANDN U18991 ( .B(n15678), .A(\u_a23_core/u_execute/u_register_bank/r10[26] ), .Z(n16151) );
  NANDN U18992 ( .B(n15679), .A(\u_a23_core/u_execute/u_register_bank/r9[26] ), 
        .Z(n16150) );
  AND U18993 ( .A(n16152), .B(n16153), .Z(n16148) );
  NANDN U18994 ( .B(n15682), .A(\u_a23_core/u_execute/u_register_bank/r8[26] ), 
        .Z(n16153) );
  NANDN U18995 ( .B(n15683), .A(\u_a23_core/u_execute/u_register_bank/r7[26] ), 
        .Z(n16152) );
  AND U18996 ( .A(n16154), .B(n16155), .Z(n16138) );
  AND U18997 ( .A(n16156), .B(n16157), .Z(n16155) );
  AND U18998 ( .A(n16158), .B(n16159), .Z(n16157) );
  NANDN U18999 ( .B(n15690), .A(\u_a23_core/u_execute/u_register_bank/r6[26] ), 
        .Z(n16159) );
  NANDN U19000 ( .B(n15691), .A(\u_a23_core/u_execute/u_register_bank/r5[26] ), 
        .Z(n16158) );
  AND U19001 ( .A(n16160), .B(n16161), .Z(n16156) );
  NANDN U19002 ( .B(n15694), .A(\u_a23_core/u_execute/u_register_bank/r4[26] ), 
        .Z(n16161) );
  NANDN U19003 ( .B(n15695), .A(\u_a23_core/u_execute/u_register_bank/r3[26] ), 
        .Z(n16160) );
  AND U19004 ( .A(n16162), .B(n16163), .Z(n16154) );
  NANDN U19005 ( .B(n15698), .A(\u_a23_core/u_execute/u_register_bank/r2[26] ), 
        .Z(n16163) );
  AND U19006 ( .A(n16164), .B(n16165), .Z(n16162) );
  NANDN U19007 ( .B(n15701), .A(\u_a23_core/u_execute/u_register_bank/r1[26] ), 
        .Z(n16165) );
  NANDN U19008 ( .B(n15702), .A(\u_a23_core/u_execute/u_register_bank/r0[26] ), 
        .Z(n16164) );
  IV U19009 ( .A(\u_a23_core/u_execute/rs[27] ), .Z(n16622) );
  NAND U19010 ( .A(n16166), .B(n16167), .Z(\u_a23_core/u_execute/rs[27] ) );
  AND U19011 ( .A(n16168), .B(n16169), .Z(n16167) );
  AND U19012 ( .A(n16170), .B(n16171), .Z(n16169) );
  AND U19013 ( .A(n16172), .B(n16173), .Z(n16171) );
  NAND U19014 ( .A(n15668), .B(\u_a23_core/u_execute/u_register_bank/r14[27] ), 
        .Z(n16173) );
  NANDN U19015 ( .B(n15669), .A(\u_a23_core/u_execute/u_register_bank/r13[27] ), .Z(n16172) );
  AND U19016 ( .A(n16174), .B(n16175), .Z(n16170) );
  NANDN U19017 ( .B(n15672), .A(\u_a23_core/u_execute/u_register_bank/r12[27] ), .Z(n16175) );
  NANDN U19018 ( .B(n15673), .A(\u_a23_core/u_execute/u_register_bank/r11[27] ), .Z(n16174) );
  AND U19019 ( .A(n16176), .B(n16177), .Z(n16168) );
  AND U19020 ( .A(n16178), .B(n16179), .Z(n16177) );
  NANDN U19021 ( .B(n15678), .A(\u_a23_core/u_execute/u_register_bank/r10[27] ), .Z(n16179) );
  NANDN U19022 ( .B(n15679), .A(\u_a23_core/u_execute/u_register_bank/r9[27] ), 
        .Z(n16178) );
  AND U19023 ( .A(n16180), .B(n16181), .Z(n16176) );
  NANDN U19024 ( .B(n15682), .A(\u_a23_core/u_execute/u_register_bank/r8[27] ), 
        .Z(n16181) );
  NANDN U19025 ( .B(n15683), .A(\u_a23_core/u_execute/u_register_bank/r7[27] ), 
        .Z(n16180) );
  AND U19026 ( .A(n16182), .B(n16183), .Z(n16166) );
  AND U19027 ( .A(n16184), .B(n16185), .Z(n16183) );
  AND U19028 ( .A(n16186), .B(n16187), .Z(n16185) );
  NANDN U19029 ( .B(n15690), .A(\u_a23_core/u_execute/u_register_bank/r6[27] ), 
        .Z(n16187) );
  NANDN U19030 ( .B(n15691), .A(\u_a23_core/u_execute/u_register_bank/r5[27] ), 
        .Z(n16186) );
  AND U19031 ( .A(n16188), .B(n16189), .Z(n16184) );
  NANDN U19032 ( .B(n15694), .A(\u_a23_core/u_execute/u_register_bank/r4[27] ), 
        .Z(n16189) );
  NANDN U19033 ( .B(n15695), .A(\u_a23_core/u_execute/u_register_bank/r3[27] ), 
        .Z(n16188) );
  AND U19034 ( .A(n16190), .B(n16191), .Z(n16182) );
  NANDN U19035 ( .B(n15698), .A(\u_a23_core/u_execute/u_register_bank/r2[27] ), 
        .Z(n16191) );
  AND U19036 ( .A(n16192), .B(n16193), .Z(n16190) );
  NANDN U19037 ( .B(n15701), .A(\u_a23_core/u_execute/u_register_bank/r1[27] ), 
        .Z(n16193) );
  NANDN U19038 ( .B(n15702), .A(\u_a23_core/u_execute/u_register_bank/r0[27] ), 
        .Z(n16192) );
  IV U19039 ( .A(\u_a23_core/u_execute/rs[28] ), .Z(n16623) );
  NAND U19040 ( .A(n16194), .B(n16195), .Z(\u_a23_core/u_execute/rs[28] ) );
  AND U19041 ( .A(n16196), .B(n16197), .Z(n16195) );
  AND U19042 ( .A(n16198), .B(n16199), .Z(n16197) );
  AND U19043 ( .A(n16200), .B(n16201), .Z(n16199) );
  NAND U19044 ( .A(n15668), .B(\u_a23_core/u_execute/u_register_bank/r14[28] ), 
        .Z(n16201) );
  NANDN U19045 ( .B(n15669), .A(\u_a23_core/u_execute/u_register_bank/r13[28] ), .Z(n16200) );
  AND U19046 ( .A(n16202), .B(n16203), .Z(n16198) );
  NANDN U19047 ( .B(n15672), .A(\u_a23_core/u_execute/u_register_bank/r12[28] ), .Z(n16203) );
  NANDN U19048 ( .B(n15673), .A(\u_a23_core/u_execute/u_register_bank/r11[28] ), .Z(n16202) );
  AND U19049 ( .A(n16204), .B(n16205), .Z(n16196) );
  AND U19050 ( .A(n16206), .B(n16207), .Z(n16205) );
  NANDN U19051 ( .B(n15678), .A(\u_a23_core/u_execute/u_register_bank/r10[28] ), .Z(n16207) );
  NANDN U19052 ( .B(n15679), .A(\u_a23_core/u_execute/u_register_bank/r9[28] ), 
        .Z(n16206) );
  AND U19053 ( .A(n16208), .B(n16209), .Z(n16204) );
  NANDN U19054 ( .B(n15682), .A(\u_a23_core/u_execute/u_register_bank/r8[28] ), 
        .Z(n16209) );
  NANDN U19055 ( .B(n15683), .A(\u_a23_core/u_execute/u_register_bank/r7[28] ), 
        .Z(n16208) );
  AND U19056 ( .A(n16210), .B(n16211), .Z(n16194) );
  AND U19057 ( .A(n16212), .B(n16213), .Z(n16211) );
  AND U19058 ( .A(n16214), .B(n16215), .Z(n16213) );
  NANDN U19059 ( .B(n15690), .A(\u_a23_core/u_execute/u_register_bank/r6[28] ), 
        .Z(n16215) );
  NANDN U19060 ( .B(n15691), .A(\u_a23_core/u_execute/u_register_bank/r5[28] ), 
        .Z(n16214) );
  AND U19061 ( .A(n16216), .B(n16217), .Z(n16212) );
  NANDN U19062 ( .B(n15694), .A(\u_a23_core/u_execute/u_register_bank/r4[28] ), 
        .Z(n16217) );
  NANDN U19063 ( .B(n15695), .A(\u_a23_core/u_execute/u_register_bank/r3[28] ), 
        .Z(n16216) );
  AND U19064 ( .A(n16218), .B(n16219), .Z(n16210) );
  NANDN U19065 ( .B(n15698), .A(\u_a23_core/u_execute/u_register_bank/r2[28] ), 
        .Z(n16219) );
  AND U19066 ( .A(n16220), .B(n16221), .Z(n16218) );
  NANDN U19067 ( .B(n15701), .A(\u_a23_core/u_execute/u_register_bank/r1[28] ), 
        .Z(n16221) );
  NANDN U19068 ( .B(n15702), .A(\u_a23_core/u_execute/u_register_bank/r0[28] ), 
        .Z(n16220) );
  IV U19069 ( .A(\u_a23_core/u_execute/rs[29] ), .Z(n16624) );
  NAND U19070 ( .A(n16222), .B(n16223), .Z(\u_a23_core/u_execute/rs[29] ) );
  AND U19071 ( .A(n16224), .B(n16225), .Z(n16223) );
  AND U19072 ( .A(n16226), .B(n16227), .Z(n16225) );
  AND U19073 ( .A(n16228), .B(n16229), .Z(n16227) );
  NAND U19074 ( .A(n15668), .B(\u_a23_core/u_execute/u_register_bank/r14[29] ), 
        .Z(n16229) );
  NANDN U19075 ( .B(n15669), .A(\u_a23_core/u_execute/u_register_bank/r13[29] ), .Z(n16228) );
  AND U19076 ( .A(n16230), .B(n16231), .Z(n16226) );
  NANDN U19077 ( .B(n15672), .A(\u_a23_core/u_execute/u_register_bank/r12[29] ), .Z(n16231) );
  NANDN U19078 ( .B(n15673), .A(\u_a23_core/u_execute/u_register_bank/r11[29] ), .Z(n16230) );
  AND U19079 ( .A(n16232), .B(n16233), .Z(n16224) );
  AND U19080 ( .A(n16234), .B(n16235), .Z(n16233) );
  NANDN U19081 ( .B(n15678), .A(\u_a23_core/u_execute/u_register_bank/r10[29] ), .Z(n16235) );
  NANDN U19082 ( .B(n15679), .A(\u_a23_core/u_execute/u_register_bank/r9[29] ), 
        .Z(n16234) );
  AND U19083 ( .A(n16236), .B(n16237), .Z(n16232) );
  NANDN U19084 ( .B(n15682), .A(\u_a23_core/u_execute/u_register_bank/r8[29] ), 
        .Z(n16237) );
  NANDN U19085 ( .B(n15683), .A(\u_a23_core/u_execute/u_register_bank/r7[29] ), 
        .Z(n16236) );
  AND U19086 ( .A(n16238), .B(n16239), .Z(n16222) );
  AND U19087 ( .A(n16240), .B(n16241), .Z(n16239) );
  AND U19088 ( .A(n16242), .B(n16243), .Z(n16241) );
  NANDN U19089 ( .B(n15690), .A(\u_a23_core/u_execute/u_register_bank/r6[29] ), 
        .Z(n16243) );
  NANDN U19090 ( .B(n15691), .A(\u_a23_core/u_execute/u_register_bank/r5[29] ), 
        .Z(n16242) );
  AND U19091 ( .A(n16244), .B(n16245), .Z(n16240) );
  NANDN U19092 ( .B(n15694), .A(\u_a23_core/u_execute/u_register_bank/r4[29] ), 
        .Z(n16245) );
  NANDN U19093 ( .B(n15695), .A(\u_a23_core/u_execute/u_register_bank/r3[29] ), 
        .Z(n16244) );
  AND U19094 ( .A(n16246), .B(n16247), .Z(n16238) );
  NANDN U19095 ( .B(n15698), .A(\u_a23_core/u_execute/u_register_bank/r2[29] ), 
        .Z(n16247) );
  AND U19096 ( .A(n16248), .B(n16249), .Z(n16246) );
  NANDN U19097 ( .B(n15701), .A(\u_a23_core/u_execute/u_register_bank/r1[29] ), 
        .Z(n16249) );
  NANDN U19098 ( .B(n15702), .A(\u_a23_core/u_execute/u_register_bank/r0[29] ), 
        .Z(n16248) );
  AND U19099 ( .A(n16250), .B(n6064), .Z(n16625) );
  AND U19100 ( .A(n16251), .B(n16252), .Z(n6064) );
  AND U19101 ( .A(n16253), .B(n16254), .Z(n16252) );
  AND U19102 ( .A(n16255), .B(n16256), .Z(n16254) );
  AND U19103 ( .A(n16257), .B(n16258), .Z(n16256) );
  NAND U19104 ( .A(n15668), .B(\u_a23_core/u_execute/u_register_bank/r14[2] ), 
        .Z(n16258) );
  NANDN U19105 ( .B(n15669), .A(\u_a23_core/u_execute/u_register_bank/r13[2] ), 
        .Z(n16257) );
  AND U19106 ( .A(n16259), .B(n16260), .Z(n16255) );
  NANDN U19107 ( .B(n15672), .A(\u_a23_core/u_execute/u_register_bank/r12[2] ), 
        .Z(n16260) );
  NANDN U19108 ( .B(n15673), .A(\u_a23_core/u_execute/u_register_bank/r11[2] ), 
        .Z(n16259) );
  AND U19109 ( .A(n16261), .B(n16262), .Z(n16253) );
  AND U19110 ( .A(n16263), .B(n16264), .Z(n16262) );
  NANDN U19111 ( .B(n15678), .A(\u_a23_core/u_execute/u_register_bank/r10[2] ), 
        .Z(n16264) );
  NANDN U19112 ( .B(n15679), .A(\u_a23_core/u_execute/u_register_bank/r9[2] ), 
        .Z(n16263) );
  AND U19113 ( .A(n16265), .B(n16266), .Z(n16261) );
  NANDN U19114 ( .B(n15682), .A(\u_a23_core/u_execute/u_register_bank/r8[2] ), 
        .Z(n16266) );
  NANDN U19115 ( .B(n15683), .A(\u_a23_core/u_execute/u_register_bank/r7[2] ), 
        .Z(n16265) );
  AND U19116 ( .A(n16267), .B(n16268), .Z(n16251) );
  AND U19117 ( .A(n16269), .B(n16270), .Z(n16268) );
  AND U19118 ( .A(n16271), .B(n16272), .Z(n16270) );
  NANDN U19119 ( .B(n15690), .A(\u_a23_core/u_execute/u_register_bank/r6[2] ), 
        .Z(n16272) );
  NANDN U19120 ( .B(n15691), .A(\u_a23_core/u_execute/u_register_bank/r5[2] ), 
        .Z(n16271) );
  AND U19121 ( .A(n16273), .B(n16274), .Z(n16269) );
  NANDN U19122 ( .B(n15694), .A(\u_a23_core/u_execute/u_register_bank/r4[2] ), 
        .Z(n16274) );
  NANDN U19123 ( .B(n15695), .A(\u_a23_core/u_execute/u_register_bank/r3[2] ), 
        .Z(n16273) );
  AND U19124 ( .A(n16275), .B(n16276), .Z(n16267) );
  NANDN U19125 ( .B(n15698), .A(\u_a23_core/u_execute/u_register_bank/r2[2] ), 
        .Z(n16276) );
  AND U19126 ( .A(n16277), .B(n16278), .Z(n16275) );
  NANDN U19127 ( .B(n15701), .A(\u_a23_core/u_execute/u_register_bank/r1[2] ), 
        .Z(n16278) );
  NANDN U19128 ( .B(n15702), .A(\u_a23_core/u_execute/u_register_bank/r0[2] ), 
        .Z(n16277) );
  NAND U19129 ( .A(\u_a23_core/u_execute/pc[2] ), .B(n6025), .Z(n16250) );
  IV U19130 ( .A(\u_a23_core/u_execute/rs[30] ), .Z(n16626) );
  NAND U19131 ( .A(n16279), .B(n16280), .Z(\u_a23_core/u_execute/rs[30] ) );
  AND U19132 ( .A(n16281), .B(n16282), .Z(n16280) );
  AND U19133 ( .A(n16283), .B(n16284), .Z(n16282) );
  AND U19134 ( .A(n16285), .B(n16286), .Z(n16284) );
  NAND U19135 ( .A(n15668), .B(\u_a23_core/u_execute/u_register_bank/r14[30] ), 
        .Z(n16286) );
  NANDN U19136 ( .B(n15669), .A(\u_a23_core/u_execute/u_register_bank/r13[30] ), .Z(n16285) );
  AND U19137 ( .A(n16287), .B(n16288), .Z(n16283) );
  NANDN U19138 ( .B(n15672), .A(\u_a23_core/u_execute/u_register_bank/r12[30] ), .Z(n16288) );
  NANDN U19139 ( .B(n15673), .A(\u_a23_core/u_execute/u_register_bank/r11[30] ), .Z(n16287) );
  AND U19140 ( .A(n16289), .B(n16290), .Z(n16281) );
  AND U19141 ( .A(n16291), .B(n16292), .Z(n16290) );
  NANDN U19142 ( .B(n15678), .A(\u_a23_core/u_execute/u_register_bank/r10[30] ), .Z(n16292) );
  NANDN U19143 ( .B(n15679), .A(\u_a23_core/u_execute/u_register_bank/r9[30] ), 
        .Z(n16291) );
  AND U19144 ( .A(n16293), .B(n16294), .Z(n16289) );
  NANDN U19145 ( .B(n15682), .A(\u_a23_core/u_execute/u_register_bank/r8[30] ), 
        .Z(n16294) );
  NANDN U19146 ( .B(n15683), .A(\u_a23_core/u_execute/u_register_bank/r7[30] ), 
        .Z(n16293) );
  AND U19147 ( .A(n16295), .B(n16296), .Z(n16279) );
  AND U19148 ( .A(n16297), .B(n16298), .Z(n16296) );
  AND U19149 ( .A(n16299), .B(n16300), .Z(n16298) );
  NANDN U19150 ( .B(n15690), .A(\u_a23_core/u_execute/u_register_bank/r6[30] ), 
        .Z(n16300) );
  NANDN U19151 ( .B(n15691), .A(\u_a23_core/u_execute/u_register_bank/r5[30] ), 
        .Z(n16299) );
  AND U19152 ( .A(n16301), .B(n16302), .Z(n16297) );
  NANDN U19153 ( .B(n15694), .A(\u_a23_core/u_execute/u_register_bank/r4[30] ), 
        .Z(n16302) );
  NANDN U19154 ( .B(n15695), .A(\u_a23_core/u_execute/u_register_bank/r3[30] ), 
        .Z(n16301) );
  AND U19155 ( .A(n16303), .B(n16304), .Z(n16295) );
  NANDN U19156 ( .B(n15698), .A(\u_a23_core/u_execute/u_register_bank/r2[30] ), 
        .Z(n16304) );
  AND U19157 ( .A(n16305), .B(n16306), .Z(n16303) );
  NANDN U19158 ( .B(n15701), .A(\u_a23_core/u_execute/u_register_bank/r1[30] ), 
        .Z(n16306) );
  NANDN U19159 ( .B(n15702), .A(\u_a23_core/u_execute/u_register_bank/r0[30] ), 
        .Z(n16305) );
  IV U19160 ( .A(\u_a23_core/u_execute/rs[31] ), .Z(n16627) );
  NAND U19161 ( .A(n16307), .B(n16308), .Z(\u_a23_core/u_execute/rs[31] ) );
  AND U19162 ( .A(n16309), .B(n16310), .Z(n16308) );
  AND U19163 ( .A(n16311), .B(n16312), .Z(n16310) );
  AND U19164 ( .A(n16313), .B(n16314), .Z(n16312) );
  NAND U19165 ( .A(n15668), .B(\u_a23_core/u_execute/u_register_bank/r14[31] ), 
        .Z(n16314) );
  NANDN U19166 ( .B(n15669), .A(\u_a23_core/u_execute/u_register_bank/r13[31] ), .Z(n16313) );
  AND U19167 ( .A(n16315), .B(n16316), .Z(n16311) );
  NANDN U19168 ( .B(n15672), .A(\u_a23_core/u_execute/u_register_bank/r12[31] ), .Z(n16316) );
  NANDN U19169 ( .B(n15673), .A(\u_a23_core/u_execute/u_register_bank/r11[31] ), .Z(n16315) );
  AND U19170 ( .A(n16317), .B(n16318), .Z(n16309) );
  AND U19171 ( .A(n16319), .B(n16320), .Z(n16318) );
  NANDN U19172 ( .B(n15678), .A(\u_a23_core/u_execute/u_register_bank/r10[31] ), .Z(n16320) );
  NANDN U19173 ( .B(n15679), .A(\u_a23_core/u_execute/u_register_bank/r9[31] ), 
        .Z(n16319) );
  AND U19174 ( .A(n16321), .B(n16322), .Z(n16317) );
  NANDN U19175 ( .B(n15682), .A(\u_a23_core/u_execute/u_register_bank/r8[31] ), 
        .Z(n16322) );
  NANDN U19176 ( .B(n15683), .A(\u_a23_core/u_execute/u_register_bank/r7[31] ), 
        .Z(n16321) );
  AND U19177 ( .A(n16323), .B(n16324), .Z(n16307) );
  AND U19178 ( .A(n16325), .B(n16326), .Z(n16324) );
  AND U19179 ( .A(n16327), .B(n16328), .Z(n16326) );
  NANDN U19180 ( .B(n15690), .A(\u_a23_core/u_execute/u_register_bank/r6[31] ), 
        .Z(n16328) );
  NANDN U19181 ( .B(n15691), .A(\u_a23_core/u_execute/u_register_bank/r5[31] ), 
        .Z(n16327) );
  AND U19182 ( .A(n16329), .B(n16330), .Z(n16325) );
  NANDN U19183 ( .B(n15694), .A(\u_a23_core/u_execute/u_register_bank/r4[31] ), 
        .Z(n16330) );
  NANDN U19184 ( .B(n15695), .A(\u_a23_core/u_execute/u_register_bank/r3[31] ), 
        .Z(n16329) );
  AND U19185 ( .A(n16331), .B(n16332), .Z(n16323) );
  NANDN U19186 ( .B(n15698), .A(\u_a23_core/u_execute/u_register_bank/r2[31] ), 
        .Z(n16332) );
  AND U19187 ( .A(n16333), .B(n16334), .Z(n16331) );
  NANDN U19188 ( .B(n15701), .A(\u_a23_core/u_execute/u_register_bank/r1[31] ), 
        .Z(n16334) );
  NANDN U19189 ( .B(n15702), .A(\u_a23_core/u_execute/u_register_bank/r0[31] ), 
        .Z(n16333) );
  AND U19190 ( .A(n16335), .B(n6056), .Z(n16628) );
  AND U19191 ( .A(n16336), .B(n16337), .Z(n6056) );
  AND U19192 ( .A(n16338), .B(n16339), .Z(n16337) );
  AND U19193 ( .A(n16340), .B(n16341), .Z(n16339) );
  AND U19194 ( .A(n16342), .B(n16343), .Z(n16341) );
  NAND U19195 ( .A(n15668), .B(\u_a23_core/u_execute/u_register_bank/r14[3] ), 
        .Z(n16343) );
  NANDN U19196 ( .B(n15669), .A(\u_a23_core/u_execute/u_register_bank/r13[3] ), 
        .Z(n16342) );
  AND U19197 ( .A(n16344), .B(n16345), .Z(n16340) );
  NANDN U19198 ( .B(n15672), .A(\u_a23_core/u_execute/u_register_bank/r12[3] ), 
        .Z(n16345) );
  NANDN U19199 ( .B(n15673), .A(\u_a23_core/u_execute/u_register_bank/r11[3] ), 
        .Z(n16344) );
  AND U19200 ( .A(n16346), .B(n16347), .Z(n16338) );
  AND U19201 ( .A(n16348), .B(n16349), .Z(n16347) );
  NANDN U19202 ( .B(n15678), .A(\u_a23_core/u_execute/u_register_bank/r10[3] ), 
        .Z(n16349) );
  NANDN U19203 ( .B(n15679), .A(\u_a23_core/u_execute/u_register_bank/r9[3] ), 
        .Z(n16348) );
  AND U19204 ( .A(n16350), .B(n16351), .Z(n16346) );
  NANDN U19205 ( .B(n15682), .A(\u_a23_core/u_execute/u_register_bank/r8[3] ), 
        .Z(n16351) );
  NANDN U19206 ( .B(n15683), .A(\u_a23_core/u_execute/u_register_bank/r7[3] ), 
        .Z(n16350) );
  AND U19207 ( .A(n16352), .B(n16353), .Z(n16336) );
  AND U19208 ( .A(n16354), .B(n16355), .Z(n16353) );
  AND U19209 ( .A(n16356), .B(n16357), .Z(n16355) );
  NANDN U19210 ( .B(n15690), .A(\u_a23_core/u_execute/u_register_bank/r6[3] ), 
        .Z(n16357) );
  NANDN U19211 ( .B(n15691), .A(\u_a23_core/u_execute/u_register_bank/r5[3] ), 
        .Z(n16356) );
  AND U19212 ( .A(n16358), .B(n16359), .Z(n16354) );
  NANDN U19213 ( .B(n15694), .A(\u_a23_core/u_execute/u_register_bank/r4[3] ), 
        .Z(n16359) );
  NANDN U19214 ( .B(n15695), .A(\u_a23_core/u_execute/u_register_bank/r3[3] ), 
        .Z(n16358) );
  AND U19215 ( .A(n16360), .B(n16361), .Z(n16352) );
  NANDN U19216 ( .B(n15698), .A(\u_a23_core/u_execute/u_register_bank/r2[3] ), 
        .Z(n16361) );
  AND U19217 ( .A(n16362), .B(n16363), .Z(n16360) );
  NANDN U19218 ( .B(n15701), .A(\u_a23_core/u_execute/u_register_bank/r1[3] ), 
        .Z(n16363) );
  NANDN U19219 ( .B(n15702), .A(\u_a23_core/u_execute/u_register_bank/r0[3] ), 
        .Z(n16362) );
  NAND U19220 ( .A(n6025), .B(\u_a23_core/u_execute/pc[3] ), .Z(n16335) );
  AND U19221 ( .A(n16364), .B(n6048), .Z(n16629) );
  AND U19222 ( .A(n16365), .B(n16366), .Z(n6048) );
  AND U19223 ( .A(n16367), .B(n16368), .Z(n16366) );
  AND U19224 ( .A(n16369), .B(n16370), .Z(n16368) );
  AND U19225 ( .A(n16371), .B(n16372), .Z(n16370) );
  NAND U19226 ( .A(n15668), .B(\u_a23_core/u_execute/u_register_bank/r14[4] ), 
        .Z(n16372) );
  NANDN U19227 ( .B(n15669), .A(\u_a23_core/u_execute/u_register_bank/r13[4] ), 
        .Z(n16371) );
  AND U19228 ( .A(n16373), .B(n16374), .Z(n16369) );
  NANDN U19229 ( .B(n15672), .A(\u_a23_core/u_execute/u_register_bank/r12[4] ), 
        .Z(n16374) );
  NANDN U19230 ( .B(n15673), .A(\u_a23_core/u_execute/u_register_bank/r11[4] ), 
        .Z(n16373) );
  AND U19231 ( .A(n16375), .B(n16376), .Z(n16367) );
  AND U19232 ( .A(n16377), .B(n16378), .Z(n16376) );
  NANDN U19233 ( .B(n15678), .A(\u_a23_core/u_execute/u_register_bank/r10[4] ), 
        .Z(n16378) );
  NANDN U19234 ( .B(n15679), .A(\u_a23_core/u_execute/u_register_bank/r9[4] ), 
        .Z(n16377) );
  AND U19235 ( .A(n16379), .B(n16380), .Z(n16375) );
  NANDN U19236 ( .B(n15682), .A(\u_a23_core/u_execute/u_register_bank/r8[4] ), 
        .Z(n16380) );
  NANDN U19237 ( .B(n15683), .A(\u_a23_core/u_execute/u_register_bank/r7[4] ), 
        .Z(n16379) );
  AND U19238 ( .A(n16381), .B(n16382), .Z(n16365) );
  AND U19239 ( .A(n16383), .B(n16384), .Z(n16382) );
  AND U19240 ( .A(n16385), .B(n16386), .Z(n16384) );
  NANDN U19241 ( .B(n15690), .A(\u_a23_core/u_execute/u_register_bank/r6[4] ), 
        .Z(n16386) );
  NANDN U19242 ( .B(n15691), .A(\u_a23_core/u_execute/u_register_bank/r5[4] ), 
        .Z(n16385) );
  AND U19243 ( .A(n16387), .B(n16388), .Z(n16383) );
  NANDN U19244 ( .B(n15694), .A(\u_a23_core/u_execute/u_register_bank/r4[4] ), 
        .Z(n16388) );
  NANDN U19245 ( .B(n15695), .A(\u_a23_core/u_execute/u_register_bank/r3[4] ), 
        .Z(n16387) );
  AND U19246 ( .A(n16389), .B(n16390), .Z(n16381) );
  NANDN U19247 ( .B(n15698), .A(\u_a23_core/u_execute/u_register_bank/r2[4] ), 
        .Z(n16390) );
  AND U19248 ( .A(n16391), .B(n16392), .Z(n16389) );
  NANDN U19249 ( .B(n15701), .A(\u_a23_core/u_execute/u_register_bank/r1[4] ), 
        .Z(n16392) );
  NANDN U19250 ( .B(n15702), .A(\u_a23_core/u_execute/u_register_bank/r0[4] ), 
        .Z(n16391) );
  NAND U19251 ( .A(n6025), .B(\u_a23_core/u_execute/pc[4] ), .Z(n16364) );
  AND U19252 ( .A(n16393), .B(n6040), .Z(n16630) );
  AND U19253 ( .A(n16394), .B(n16395), .Z(n6040) );
  AND U19254 ( .A(n16396), .B(n16397), .Z(n16395) );
  AND U19255 ( .A(n16398), .B(n16399), .Z(n16397) );
  AND U19256 ( .A(n16400), .B(n16401), .Z(n16399) );
  NAND U19257 ( .A(n15668), .B(\u_a23_core/u_execute/u_register_bank/r14[5] ), 
        .Z(n16401) );
  NANDN U19258 ( .B(n15669), .A(\u_a23_core/u_execute/u_register_bank/r13[5] ), 
        .Z(n16400) );
  AND U19259 ( .A(n16402), .B(n16403), .Z(n16398) );
  NANDN U19260 ( .B(n15672), .A(\u_a23_core/u_execute/u_register_bank/r12[5] ), 
        .Z(n16403) );
  NANDN U19261 ( .B(n15673), .A(\u_a23_core/u_execute/u_register_bank/r11[5] ), 
        .Z(n16402) );
  AND U19262 ( .A(n16404), .B(n16405), .Z(n16396) );
  AND U19263 ( .A(n16406), .B(n16407), .Z(n16405) );
  NANDN U19264 ( .B(n15678), .A(\u_a23_core/u_execute/u_register_bank/r10[5] ), 
        .Z(n16407) );
  NANDN U19265 ( .B(n15679), .A(\u_a23_core/u_execute/u_register_bank/r9[5] ), 
        .Z(n16406) );
  AND U19266 ( .A(n16408), .B(n16409), .Z(n16404) );
  NANDN U19267 ( .B(n15682), .A(\u_a23_core/u_execute/u_register_bank/r8[5] ), 
        .Z(n16409) );
  NANDN U19268 ( .B(n15683), .A(\u_a23_core/u_execute/u_register_bank/r7[5] ), 
        .Z(n16408) );
  AND U19269 ( .A(n16410), .B(n16411), .Z(n16394) );
  AND U19270 ( .A(n16412), .B(n16413), .Z(n16411) );
  AND U19271 ( .A(n16414), .B(n16415), .Z(n16413) );
  NANDN U19272 ( .B(n15690), .A(\u_a23_core/u_execute/u_register_bank/r6[5] ), 
        .Z(n16415) );
  NANDN U19273 ( .B(n15691), .A(\u_a23_core/u_execute/u_register_bank/r5[5] ), 
        .Z(n16414) );
  AND U19274 ( .A(n16416), .B(n16417), .Z(n16412) );
  NANDN U19275 ( .B(n15694), .A(\u_a23_core/u_execute/u_register_bank/r4[5] ), 
        .Z(n16417) );
  NANDN U19276 ( .B(n15695), .A(\u_a23_core/u_execute/u_register_bank/r3[5] ), 
        .Z(n16416) );
  AND U19277 ( .A(n16418), .B(n16419), .Z(n16410) );
  NANDN U19278 ( .B(n15698), .A(\u_a23_core/u_execute/u_register_bank/r2[5] ), 
        .Z(n16419) );
  AND U19279 ( .A(n16420), .B(n16421), .Z(n16418) );
  NANDN U19280 ( .B(n15701), .A(\u_a23_core/u_execute/u_register_bank/r1[5] ), 
        .Z(n16421) );
  NANDN U19281 ( .B(n15702), .A(\u_a23_core/u_execute/u_register_bank/r0[5] ), 
        .Z(n16420) );
  NAND U19282 ( .A(n6025), .B(\u_a23_core/u_execute/pc[5] ), .Z(n16393) );
  AND U19283 ( .A(n16422), .B(n6032), .Z(n16631) );
  AND U19284 ( .A(n16423), .B(n16424), .Z(n6032) );
  AND U19285 ( .A(n16425), .B(n16426), .Z(n16424) );
  AND U19286 ( .A(n16427), .B(n16428), .Z(n16426) );
  AND U19287 ( .A(n16429), .B(n16430), .Z(n16428) );
  NAND U19288 ( .A(n15668), .B(\u_a23_core/u_execute/u_register_bank/r14[6] ), 
        .Z(n16430) );
  NANDN U19289 ( .B(n15669), .A(\u_a23_core/u_execute/u_register_bank/r13[6] ), 
        .Z(n16429) );
  AND U19290 ( .A(n16431), .B(n16432), .Z(n16427) );
  NANDN U19291 ( .B(n15672), .A(\u_a23_core/u_execute/u_register_bank/r12[6] ), 
        .Z(n16432) );
  NANDN U19292 ( .B(n15673), .A(\u_a23_core/u_execute/u_register_bank/r11[6] ), 
        .Z(n16431) );
  AND U19293 ( .A(n16433), .B(n16434), .Z(n16425) );
  AND U19294 ( .A(n16435), .B(n16436), .Z(n16434) );
  NANDN U19295 ( .B(n15678), .A(\u_a23_core/u_execute/u_register_bank/r10[6] ), 
        .Z(n16436) );
  NANDN U19296 ( .B(n15679), .A(\u_a23_core/u_execute/u_register_bank/r9[6] ), 
        .Z(n16435) );
  AND U19297 ( .A(n16437), .B(n16438), .Z(n16433) );
  NANDN U19298 ( .B(n15682), .A(\u_a23_core/u_execute/u_register_bank/r8[6] ), 
        .Z(n16438) );
  NANDN U19299 ( .B(n15683), .A(\u_a23_core/u_execute/u_register_bank/r7[6] ), 
        .Z(n16437) );
  AND U19300 ( .A(n16439), .B(n16440), .Z(n16423) );
  AND U19301 ( .A(n16441), .B(n16442), .Z(n16440) );
  AND U19302 ( .A(n16443), .B(n16444), .Z(n16442) );
  NANDN U19303 ( .B(n15690), .A(\u_a23_core/u_execute/u_register_bank/r6[6] ), 
        .Z(n16444) );
  NANDN U19304 ( .B(n15691), .A(\u_a23_core/u_execute/u_register_bank/r5[6] ), 
        .Z(n16443) );
  AND U19305 ( .A(n16445), .B(n16446), .Z(n16441) );
  NANDN U19306 ( .B(n15694), .A(\u_a23_core/u_execute/u_register_bank/r4[6] ), 
        .Z(n16446) );
  NANDN U19307 ( .B(n15695), .A(\u_a23_core/u_execute/u_register_bank/r3[6] ), 
        .Z(n16445) );
  AND U19308 ( .A(n16447), .B(n16448), .Z(n16439) );
  NANDN U19309 ( .B(n15698), .A(\u_a23_core/u_execute/u_register_bank/r2[6] ), 
        .Z(n16448) );
  AND U19310 ( .A(n16449), .B(n16450), .Z(n16447) );
  NANDN U19311 ( .B(n15701), .A(\u_a23_core/u_execute/u_register_bank/r1[6] ), 
        .Z(n16450) );
  NANDN U19312 ( .B(n15702), .A(\u_a23_core/u_execute/u_register_bank/r0[6] ), 
        .Z(n16449) );
  NAND U19313 ( .A(n6025), .B(\u_a23_core/u_execute/pc[6] ), .Z(n16422) );
  AND U19314 ( .A(n16451), .B(n6023), .Z(n16632) );
  AND U19315 ( .A(n16452), .B(n16453), .Z(n6023) );
  AND U19316 ( .A(n16454), .B(n16455), .Z(n16453) );
  AND U19317 ( .A(n16456), .B(n16457), .Z(n16455) );
  AND U19318 ( .A(n16458), .B(n16459), .Z(n16457) );
  NAND U19319 ( .A(n15668), .B(\u_a23_core/u_execute/u_register_bank/r14[7] ), 
        .Z(n16459) );
  NANDN U19320 ( .B(n15669), .A(\u_a23_core/u_execute/u_register_bank/r13[7] ), 
        .Z(n16458) );
  AND U19321 ( .A(n16460), .B(n16461), .Z(n16456) );
  NANDN U19322 ( .B(n15672), .A(\u_a23_core/u_execute/u_register_bank/r12[7] ), 
        .Z(n16461) );
  NANDN U19323 ( .B(n15673), .A(\u_a23_core/u_execute/u_register_bank/r11[7] ), 
        .Z(n16460) );
  AND U19324 ( .A(n16462), .B(n16463), .Z(n16454) );
  AND U19325 ( .A(n16464), .B(n16465), .Z(n16463) );
  NANDN U19326 ( .B(n15678), .A(\u_a23_core/u_execute/u_register_bank/r10[7] ), 
        .Z(n16465) );
  NANDN U19327 ( .B(n15679), .A(\u_a23_core/u_execute/u_register_bank/r9[7] ), 
        .Z(n16464) );
  AND U19328 ( .A(n16466), .B(n16467), .Z(n16462) );
  NANDN U19329 ( .B(n15682), .A(\u_a23_core/u_execute/u_register_bank/r8[7] ), 
        .Z(n16467) );
  NANDN U19330 ( .B(n15683), .A(\u_a23_core/u_execute/u_register_bank/r7[7] ), 
        .Z(n16466) );
  AND U19331 ( .A(n16468), .B(n16469), .Z(n16452) );
  AND U19332 ( .A(n16470), .B(n16471), .Z(n16469) );
  AND U19333 ( .A(n16472), .B(n16473), .Z(n16471) );
  NANDN U19334 ( .B(n15690), .A(\u_a23_core/u_execute/u_register_bank/r6[7] ), 
        .Z(n16473) );
  NANDN U19335 ( .B(n15691), .A(\u_a23_core/u_execute/u_register_bank/r5[7] ), 
        .Z(n16472) );
  AND U19336 ( .A(n16474), .B(n16475), .Z(n16470) );
  NANDN U19337 ( .B(n15694), .A(\u_a23_core/u_execute/u_register_bank/r4[7] ), 
        .Z(n16475) );
  NANDN U19338 ( .B(n15695), .A(\u_a23_core/u_execute/u_register_bank/r3[7] ), 
        .Z(n16474) );
  AND U19339 ( .A(n16476), .B(n16477), .Z(n16468) );
  NANDN U19340 ( .B(n15698), .A(\u_a23_core/u_execute/u_register_bank/r2[7] ), 
        .Z(n16477) );
  AND U19341 ( .A(n16478), .B(n16479), .Z(n16476) );
  NANDN U19342 ( .B(n15701), .A(\u_a23_core/u_execute/u_register_bank/r1[7] ), 
        .Z(n16479) );
  NANDN U19343 ( .B(n15702), .A(\u_a23_core/u_execute/u_register_bank/r0[7] ), 
        .Z(n16478) );
  NAND U19344 ( .A(n6025), .B(\u_a23_core/u_execute/pc[7] ), .Z(n16451) );
  IV U19345 ( .A(\u_a23_core/u_execute/rs[8] ), .Z(n16633) );
  NANDN U19346 ( .B(n5941), .A(n16480), .Z(\u_a23_core/u_execute/rs[8] ) );
  NAND U19347 ( .A(n6025), .B(\u_a23_core/u_execute/pc[8] ), .Z(n16480) );
  NAND U19348 ( .A(n16481), .B(n16482), .Z(n5941) );
  AND U19349 ( .A(n16483), .B(n16484), .Z(n16482) );
  AND U19350 ( .A(n16485), .B(n16486), .Z(n16484) );
  AND U19351 ( .A(n16487), .B(n16488), .Z(n16486) );
  NAND U19352 ( .A(n15668), .B(\u_a23_core/u_execute/u_register_bank/r14[8] ), 
        .Z(n16488) );
  NANDN U19353 ( .B(n15669), .A(\u_a23_core/u_execute/u_register_bank/r13[8] ), 
        .Z(n16487) );
  AND U19354 ( .A(n16489), .B(n16490), .Z(n16485) );
  NANDN U19355 ( .B(n15672), .A(\u_a23_core/u_execute/u_register_bank/r12[8] ), 
        .Z(n16490) );
  NANDN U19356 ( .B(n15673), .A(\u_a23_core/u_execute/u_register_bank/r11[8] ), 
        .Z(n16489) );
  AND U19357 ( .A(n16491), .B(n16492), .Z(n16483) );
  AND U19358 ( .A(n16493), .B(n16494), .Z(n16492) );
  NANDN U19359 ( .B(n15678), .A(\u_a23_core/u_execute/u_register_bank/r10[8] ), 
        .Z(n16494) );
  NANDN U19360 ( .B(n15679), .A(\u_a23_core/u_execute/u_register_bank/r9[8] ), 
        .Z(n16493) );
  AND U19361 ( .A(n16495), .B(n16496), .Z(n16491) );
  NANDN U19362 ( .B(n15682), .A(\u_a23_core/u_execute/u_register_bank/r8[8] ), 
        .Z(n16496) );
  NANDN U19363 ( .B(n15683), .A(\u_a23_core/u_execute/u_register_bank/r7[8] ), 
        .Z(n16495) );
  AND U19364 ( .A(n16497), .B(n16498), .Z(n16481) );
  AND U19365 ( .A(n16499), .B(n16500), .Z(n16498) );
  AND U19366 ( .A(n16501), .B(n16502), .Z(n16500) );
  NANDN U19367 ( .B(n15690), .A(\u_a23_core/u_execute/u_register_bank/r6[8] ), 
        .Z(n16502) );
  NANDN U19368 ( .B(n15691), .A(\u_a23_core/u_execute/u_register_bank/r5[8] ), 
        .Z(n16501) );
  AND U19369 ( .A(n16503), .B(n16504), .Z(n16499) );
  NANDN U19370 ( .B(n15694), .A(\u_a23_core/u_execute/u_register_bank/r4[8] ), 
        .Z(n16504) );
  NANDN U19371 ( .B(n15695), .A(\u_a23_core/u_execute/u_register_bank/r3[8] ), 
        .Z(n16503) );
  AND U19372 ( .A(n16505), .B(n16506), .Z(n16497) );
  NANDN U19373 ( .B(n15698), .A(\u_a23_core/u_execute/u_register_bank/r2[8] ), 
        .Z(n16506) );
  AND U19374 ( .A(n16507), .B(n16508), .Z(n16505) );
  NANDN U19375 ( .B(n15701), .A(\u_a23_core/u_execute/u_register_bank/r1[8] ), 
        .Z(n16508) );
  NANDN U19376 ( .B(n15702), .A(\u_a23_core/u_execute/u_register_bank/r0[8] ), 
        .Z(n16507) );
  IV U19377 ( .A(\u_a23_core/u_execute/rs[9] ), .Z(n16634) );
  NANDN U19378 ( .B(n5934), .A(n16509), .Z(\u_a23_core/u_execute/rs[9] ) );
  NAND U19379 ( .A(n6025), .B(\u_a23_core/u_execute/pc[9] ), .Z(n16509) );
  AND U19380 ( .A(n16510), .B(n16511), .Z(n6025) );
  NAND U19381 ( .A(n16512), .B(n16513), .Z(n5934) );
  AND U19382 ( .A(n16514), .B(n16515), .Z(n16513) );
  AND U19383 ( .A(n16516), .B(n16517), .Z(n16515) );
  AND U19384 ( .A(n16518), .B(n16519), .Z(n16517) );
  NAND U19385 ( .A(n15668), .B(\u_a23_core/u_execute/u_register_bank/r14[9] ), 
        .Z(n16519) );
  NANDN U19386 ( .B(n15669), .A(\u_a23_core/u_execute/u_register_bank/r13[9] ), 
        .Z(n16518) );
  AND U19387 ( .A(n16520), .B(n16521), .Z(n16516) );
  NANDN U19388 ( .B(n15672), .A(\u_a23_core/u_execute/u_register_bank/r12[9] ), 
        .Z(n16521) );
  NANDN U19389 ( .B(n15673), .A(\u_a23_core/u_execute/u_register_bank/r11[9] ), 
        .Z(n16520) );
  AND U19390 ( .A(n16522), .B(n16523), .Z(n16514) );
  AND U19391 ( .A(n16524), .B(n16525), .Z(n16523) );
  NANDN U19392 ( .B(n15678), .A(\u_a23_core/u_execute/u_register_bank/r10[9] ), 
        .Z(n16525) );
  NANDN U19393 ( .B(n15679), .A(\u_a23_core/u_execute/u_register_bank/r9[9] ), 
        .Z(n16524) );
  AND U19394 ( .A(n16526), .B(n16527), .Z(n16522) );
  NANDN U19395 ( .B(n15682), .A(\u_a23_core/u_execute/u_register_bank/r8[9] ), 
        .Z(n16527) );
  NANDN U19396 ( .B(n15683), .A(\u_a23_core/u_execute/u_register_bank/r7[9] ), 
        .Z(n16526) );
  AND U19397 ( .A(n16528), .B(n16529), .Z(n16512) );
  AND U19398 ( .A(n16530), .B(n16531), .Z(n16529) );
  AND U19399 ( .A(n16532), .B(n16533), .Z(n16531) );
  NANDN U19400 ( .B(n15690), .A(\u_a23_core/u_execute/u_register_bank/r6[9] ), 
        .Z(n16533) );
  NANDN U19401 ( .B(n15691), .A(\u_a23_core/u_execute/u_register_bank/r5[9] ), 
        .Z(n16532) );
  AND U19402 ( .A(n16534), .B(n16535), .Z(n16530) );
  NANDN U19403 ( .B(n15694), .A(\u_a23_core/u_execute/u_register_bank/r4[9] ), 
        .Z(n16535) );
  NANDN U19404 ( .B(n15695), .A(\u_a23_core/u_execute/u_register_bank/r3[9] ), 
        .Z(n16534) );
  AND U19405 ( .A(n16536), .B(n16537), .Z(n16528) );
  NANDN U19406 ( .B(n15698), .A(\u_a23_core/u_execute/u_register_bank/r2[9] ), 
        .Z(n16537) );
  AND U19407 ( .A(n16538), .B(n16539), .Z(n16536) );
  NANDN U19408 ( .B(n15701), .A(\u_a23_core/u_execute/u_register_bank/r1[9] ), 
        .Z(n16539) );
  NANDN U19409 ( .B(n15702), .A(\u_a23_core/u_execute/u_register_bank/r0[9] ), 
        .Z(n16538) );
  IV U19410 ( .A(\u_a23_core/u_execute/rs[0] ), .Z(n16635) );
  NAND U19411 ( .A(n16540), .B(n16541), .Z(\u_a23_core/u_execute/rs[0] ) );
  AND U19412 ( .A(n16542), .B(n16543), .Z(n16541) );
  AND U19413 ( .A(n16544), .B(n16545), .Z(n16543) );
  AND U19414 ( .A(n16546), .B(n16547), .Z(n16545) );
  NAND U19415 ( .A(n15668), .B(\u_a23_core/u_execute/u_register_bank/r14[0] ), 
        .Z(n16547) );
  NANDN U19416 ( .B(n15669), .A(\u_a23_core/u_execute/u_register_bank/r13[0] ), 
        .Z(n16546) );
  AND U19417 ( .A(n16548), .B(n16549), .Z(n16544) );
  NANDN U19418 ( .B(n15672), .A(\u_a23_core/u_execute/u_register_bank/r12[0] ), 
        .Z(n16549) );
  NANDN U19419 ( .B(n15673), .A(\u_a23_core/u_execute/u_register_bank/r11[0] ), 
        .Z(n16548) );
  AND U19420 ( .A(n16550), .B(n16551), .Z(n16542) );
  AND U19421 ( .A(n16552), .B(n16553), .Z(n16551) );
  NANDN U19422 ( .B(n15678), .A(\u_a23_core/u_execute/u_register_bank/r10[0] ), 
        .Z(n16553) );
  NANDN U19423 ( .B(n15679), .A(\u_a23_core/u_execute/u_register_bank/r9[0] ), 
        .Z(n16552) );
  AND U19424 ( .A(n16554), .B(n16555), .Z(n16550) );
  NANDN U19425 ( .B(n15682), .A(\u_a23_core/u_execute/u_register_bank/r8[0] ), 
        .Z(n16555) );
  NANDN U19426 ( .B(n15683), .A(\u_a23_core/u_execute/u_register_bank/r7[0] ), 
        .Z(n16554) );
  AND U19427 ( .A(n16556), .B(n16557), .Z(n16540) );
  AND U19428 ( .A(n16558), .B(n16559), .Z(n16557) );
  AND U19429 ( .A(n16560), .B(n16561), .Z(n16559) );
  NANDN U19430 ( .B(n15690), .A(\u_a23_core/u_execute/u_register_bank/r6[0] ), 
        .Z(n16561) );
  NANDN U19431 ( .B(n15691), .A(\u_a23_core/u_execute/u_register_bank/r5[0] ), 
        .Z(n16560) );
  AND U19432 ( .A(n16562), .B(n16563), .Z(n16558) );
  NANDN U19433 ( .B(n15694), .A(\u_a23_core/u_execute/u_register_bank/r4[0] ), 
        .Z(n16563) );
  NANDN U19434 ( .B(n15695), .A(\u_a23_core/u_execute/u_register_bank/r3[0] ), 
        .Z(n16562) );
  AND U19435 ( .A(n16564), .B(n16565), .Z(n16556) );
  NANDN U19436 ( .B(n15698), .A(\u_a23_core/u_execute/u_register_bank/r2[0] ), 
        .Z(n16565) );
  AND U19437 ( .A(n16566), .B(n16567), .Z(n16564) );
  NANDN U19438 ( .B(n15701), .A(\u_a23_core/u_execute/u_register_bank/r1[0] ), 
        .Z(n16567) );
  NANDN U19439 ( .B(n15702), .A(\u_a23_core/u_execute/u_register_bank/r0[0] ), 
        .Z(n16566) );
  IV U19440 ( .A(\u_a23_core/u_execute/rs[1] ), .Z(n16636) );
  NAND U19441 ( .A(n16568), .B(n16569), .Z(\u_a23_core/u_execute/rs[1] ) );
  AND U19442 ( .A(n16570), .B(n16571), .Z(n16569) );
  AND U19443 ( .A(n16572), .B(n16573), .Z(n16571) );
  AND U19444 ( .A(n16574), .B(n16575), .Z(n16573) );
  NAND U19445 ( .A(n15668), .B(\u_a23_core/u_execute/u_register_bank/r14[1] ), 
        .Z(n16575) );
  AND U19446 ( .A(n16576), .B(n16510), .Z(n15668) );
  NANDN U19447 ( .B(n15669), .A(\u_a23_core/u_execute/u_register_bank/r13[1] ), 
        .Z(n16574) );
  NAND U19448 ( .A(n16510), .B(n16577), .Z(n15669) );
  AND U19449 ( .A(n16578), .B(n16579), .Z(n16572) );
  NANDN U19450 ( .B(n15672), .A(\u_a23_core/u_execute/u_register_bank/r12[1] ), 
        .Z(n16579) );
  NAND U19451 ( .A(n16510), .B(n16580), .Z(n15672) );
  AND U19452 ( .A(\u_a23_core/rds_sel[2] ), .B(\u_a23_core/rds_sel[3] ), .Z(
        n16510) );
  NANDN U19453 ( .B(n15673), .A(\u_a23_core/u_execute/u_register_bank/r11[1] ), 
        .Z(n16578) );
  NANDN U19454 ( .B(n16581), .A(n16511), .Z(n15673) );
  AND U19455 ( .A(n16582), .B(n16583), .Z(n16570) );
  AND U19456 ( .A(n16584), .B(n16585), .Z(n16583) );
  NANDN U19457 ( .B(n15678), .A(\u_a23_core/u_execute/u_register_bank/r10[1] ), 
        .Z(n16585) );
  NANDN U19458 ( .B(n16581), .A(n16576), .Z(n15678) );
  NANDN U19459 ( .B(n15679), .A(\u_a23_core/u_execute/u_register_bank/r9[1] ), 
        .Z(n16584) );
  NANDN U19460 ( .B(n16581), .A(n16577), .Z(n15679) );
  AND U19461 ( .A(n16586), .B(n16587), .Z(n16582) );
  NANDN U19462 ( .B(n15682), .A(\u_a23_core/u_execute/u_register_bank/r8[1] ), 
        .Z(n16587) );
  NANDN U19463 ( .B(n16581), .A(n16580), .Z(n15682) );
  NANDN U19464 ( .B(\u_a23_core/rds_sel[2] ), .A(\u_a23_core/rds_sel[3] ), .Z(
        n16581) );
  NANDN U19465 ( .B(n15683), .A(\u_a23_core/u_execute/u_register_bank/r7[1] ), 
        .Z(n16586) );
  NAND U19466 ( .A(n16588), .B(n16511), .Z(n15683) );
  AND U19467 ( .A(n16589), .B(n16590), .Z(n16568) );
  AND U19468 ( .A(n16591), .B(n16592), .Z(n16590) );
  AND U19469 ( .A(n16593), .B(n16594), .Z(n16592) );
  NANDN U19470 ( .B(n15690), .A(\u_a23_core/u_execute/u_register_bank/r6[1] ), 
        .Z(n16594) );
  NAND U19471 ( .A(n16576), .B(n16588), .Z(n15690) );
  NANDN U19472 ( .B(n15691), .A(\u_a23_core/u_execute/u_register_bank/r5[1] ), 
        .Z(n16593) );
  NAND U19473 ( .A(n16577), .B(n16588), .Z(n15691) );
  AND U19474 ( .A(n16595), .B(n16596), .Z(n16591) );
  NANDN U19475 ( .B(n15694), .A(\u_a23_core/u_execute/u_register_bank/r4[1] ), 
        .Z(n16596) );
  NAND U19476 ( .A(n16580), .B(n16588), .Z(n15694) );
  ANDN U19477 ( .A(\u_a23_core/rds_sel[2] ), .B(\u_a23_core/rds_sel[3] ), .Z(
        n16588) );
  NANDN U19478 ( .B(n15695), .A(\u_a23_core/u_execute/u_register_bank/r3[1] ), 
        .Z(n16595) );
  NAND U19479 ( .A(n16597), .B(n16511), .Z(n15695) );
  AND U19480 ( .A(\u_a23_core/rds_sel[1] ), .B(\u_a23_core/rds_sel[0] ), .Z(
        n16511) );
  AND U19481 ( .A(n16598), .B(n16599), .Z(n16589) );
  NANDN U19482 ( .B(n15698), .A(\u_a23_core/u_execute/u_register_bank/r2[1] ), 
        .Z(n16599) );
  NAND U19483 ( .A(n16576), .B(n16597), .Z(n15698) );
  AND U19484 ( .A(\u_a23_core/rds_sel[1] ), .B(n16600), .Z(n16576) );
  AND U19485 ( .A(n16601), .B(n16602), .Z(n16598) );
  NANDN U19486 ( .B(n15701), .A(\u_a23_core/u_execute/u_register_bank/r1[1] ), 
        .Z(n16602) );
  NAND U19487 ( .A(n16577), .B(n16597), .Z(n15701) );
  NOR U19488 ( .A(n16600), .B(\u_a23_core/rds_sel[1] ), .Z(n16577) );
  IV U19489 ( .A(\u_a23_core/rds_sel[0] ), .Z(n16600) );
  NANDN U19490 ( .B(n15702), .A(\u_a23_core/u_execute/u_register_bank/r0[1] ), 
        .Z(n16601) );
  NAND U19491 ( .A(n16580), .B(n16597), .Z(n15702) );
  NOR U19492 ( .A(\u_a23_core/rds_sel[3] ), .B(\u_a23_core/rds_sel[2] ), .Z(
        n16597) );
  NOR U19493 ( .A(\u_a23_core/rds_sel[0] ), .B(\u_a23_core/rds_sel[1] ), .Z(
        n16580) );
  IV U19494 ( .A(n7139), .Z(n16637) );
  NANDN U19495 ( .B(n7720), .A(n16603), .Z(n7139) );
  AND U19496 ( .A(\u_a23_core/u_decode/control_state[0] ), .B(
        \u_a23_core/u_decode/control_state[1] ), .Z(n16603) );
  NAND U19497 ( .A(\u_a23_core/u_decode/control_state[4] ), .B(n16604), .Z(
        n7720) );
  AND U19498 ( .A(n7912), .B(n7663), .Z(n16604) );
  IV U19499 ( .A(\u_a23_core/u_decode/control_state[3] ), .Z(n7663) );
  IV U19500 ( .A(\u_a23_core/u_decode/control_state[2] ), .Z(n7912) );
endmodule

