
module sum_N256_CC4 ( clk, rst, a, b, c );
  input [63:0] a;
  input [63:0] b;
  output [63:0] c;
  input clk, rst;
  wire   carry_on, carry_on_d, \ADD_/c[63] , \ADD_/c[62] , \ADD_/c[61] ,
         \ADD_/c[60] , \ADD_/c[59] , \ADD_/c[58] , \ADD_/c[57] , \ADD_/c[56] ,
         \ADD_/c[55] , \ADD_/c[54] , \ADD_/c[53] , \ADD_/c[52] , \ADD_/c[51] ,
         \ADD_/c[50] , \ADD_/c[49] , \ADD_/c[48] , \ADD_/c[47] , \ADD_/c[46] ,
         \ADD_/c[45] , \ADD_/c[44] , \ADD_/c[43] , \ADD_/c[42] , \ADD_/c[41] ,
         \ADD_/c[40] , \ADD_/c[39] , \ADD_/c[38] , \ADD_/c[37] , \ADD_/c[36] ,
         \ADD_/c[35] , \ADD_/c[34] , \ADD_/c[33] , \ADD_/c[32] , \ADD_/c[31] ,
         \ADD_/c[30] , \ADD_/c[29] , \ADD_/c[28] , \ADD_/c[27] , \ADD_/c[26] ,
         \ADD_/c[25] , \ADD_/c[24] , \ADD_/c[23] , \ADD_/c[22] , \ADD_/c[21] ,
         \ADD_/c[20] , \ADD_/c[19] , \ADD_/c[18] , \ADD_/c[17] , \ADD_/c[16] ,
         \ADD_/c[15] , \ADD_/c[14] , \ADD_/c[13] , \ADD_/c[12] , \ADD_/c[11] ,
         \ADD_/c[10] , \ADD_/c[9] , \ADD_/c[8] , \ADD_/c[7] , \ADD_/c[6] ,
         \ADD_/c[5] , \ADD_/c[4] , \ADD_/c[3] , \ADD_/c[2] , \ADD_/c[1] ,
         \ADD_/FAINST[0].FA_/n3 , \ADD_/FAINST[0].FA_/n2 ,
         \ADD_/FAINST[0].FA_/n1 , \ADD_/FAINST[63].FA_/n3 ,
         \ADD_/FAINST[63].FA_/n2 , \ADD_/FAINST[63].FA_/n1 ,
         \ADD_/FAINST[62].FA_/n3 , \ADD_/FAINST[62].FA_/n2 ,
         \ADD_/FAINST[62].FA_/n1 , \ADD_/FAINST[61].FA_/n3 ,
         \ADD_/FAINST[61].FA_/n2 , \ADD_/FAINST[61].FA_/n1 ,
         \ADD_/FAINST[60].FA_/n3 , \ADD_/FAINST[60].FA_/n2 ,
         \ADD_/FAINST[60].FA_/n1 , \ADD_/FAINST[59].FA_/n3 ,
         \ADD_/FAINST[59].FA_/n2 , \ADD_/FAINST[59].FA_/n1 ,
         \ADD_/FAINST[58].FA_/n3 , \ADD_/FAINST[58].FA_/n2 ,
         \ADD_/FAINST[58].FA_/n1 , \ADD_/FAINST[57].FA_/n3 ,
         \ADD_/FAINST[57].FA_/n2 , \ADD_/FAINST[57].FA_/n1 ,
         \ADD_/FAINST[56].FA_/n3 , \ADD_/FAINST[56].FA_/n2 ,
         \ADD_/FAINST[56].FA_/n1 , \ADD_/FAINST[55].FA_/n3 ,
         \ADD_/FAINST[55].FA_/n2 , \ADD_/FAINST[55].FA_/n1 ,
         \ADD_/FAINST[54].FA_/n3 , \ADD_/FAINST[54].FA_/n2 ,
         \ADD_/FAINST[54].FA_/n1 , \ADD_/FAINST[53].FA_/n3 ,
         \ADD_/FAINST[53].FA_/n2 , \ADD_/FAINST[53].FA_/n1 ,
         \ADD_/FAINST[52].FA_/n3 , \ADD_/FAINST[52].FA_/n2 ,
         \ADD_/FAINST[52].FA_/n1 , \ADD_/FAINST[51].FA_/n3 ,
         \ADD_/FAINST[51].FA_/n2 , \ADD_/FAINST[51].FA_/n1 ,
         \ADD_/FAINST[50].FA_/n3 , \ADD_/FAINST[50].FA_/n2 ,
         \ADD_/FAINST[50].FA_/n1 , \ADD_/FAINST[49].FA_/n3 ,
         \ADD_/FAINST[49].FA_/n2 , \ADD_/FAINST[49].FA_/n1 ,
         \ADD_/FAINST[48].FA_/n3 , \ADD_/FAINST[48].FA_/n2 ,
         \ADD_/FAINST[48].FA_/n1 , \ADD_/FAINST[47].FA_/n3 ,
         \ADD_/FAINST[47].FA_/n2 , \ADD_/FAINST[47].FA_/n1 ,
         \ADD_/FAINST[46].FA_/n3 , \ADD_/FAINST[46].FA_/n2 ,
         \ADD_/FAINST[46].FA_/n1 , \ADD_/FAINST[45].FA_/n3 ,
         \ADD_/FAINST[45].FA_/n2 , \ADD_/FAINST[45].FA_/n1 ,
         \ADD_/FAINST[44].FA_/n3 , \ADD_/FAINST[44].FA_/n2 ,
         \ADD_/FAINST[44].FA_/n1 , \ADD_/FAINST[43].FA_/n3 ,
         \ADD_/FAINST[43].FA_/n2 , \ADD_/FAINST[43].FA_/n1 ,
         \ADD_/FAINST[42].FA_/n3 , \ADD_/FAINST[42].FA_/n2 ,
         \ADD_/FAINST[42].FA_/n1 , \ADD_/FAINST[41].FA_/n3 ,
         \ADD_/FAINST[41].FA_/n2 , \ADD_/FAINST[41].FA_/n1 ,
         \ADD_/FAINST[40].FA_/n3 , \ADD_/FAINST[40].FA_/n2 ,
         \ADD_/FAINST[40].FA_/n1 , \ADD_/FAINST[39].FA_/n3 ,
         \ADD_/FAINST[39].FA_/n2 , \ADD_/FAINST[39].FA_/n1 ,
         \ADD_/FAINST[38].FA_/n3 , \ADD_/FAINST[38].FA_/n2 ,
         \ADD_/FAINST[38].FA_/n1 , \ADD_/FAINST[37].FA_/n3 ,
         \ADD_/FAINST[37].FA_/n2 , \ADD_/FAINST[37].FA_/n1 ,
         \ADD_/FAINST[36].FA_/n3 , \ADD_/FAINST[36].FA_/n2 ,
         \ADD_/FAINST[36].FA_/n1 , \ADD_/FAINST[35].FA_/n3 ,
         \ADD_/FAINST[35].FA_/n2 , \ADD_/FAINST[35].FA_/n1 ,
         \ADD_/FAINST[34].FA_/n3 , \ADD_/FAINST[34].FA_/n2 ,
         \ADD_/FAINST[34].FA_/n1 , \ADD_/FAINST[33].FA_/n3 ,
         \ADD_/FAINST[33].FA_/n2 , \ADD_/FAINST[33].FA_/n1 ,
         \ADD_/FAINST[32].FA_/n3 , \ADD_/FAINST[32].FA_/n2 ,
         \ADD_/FAINST[32].FA_/n1 , \ADD_/FAINST[31].FA_/n3 ,
         \ADD_/FAINST[31].FA_/n2 , \ADD_/FAINST[31].FA_/n1 ,
         \ADD_/FAINST[30].FA_/n3 , \ADD_/FAINST[30].FA_/n2 ,
         \ADD_/FAINST[30].FA_/n1 , \ADD_/FAINST[29].FA_/n3 ,
         \ADD_/FAINST[29].FA_/n2 , \ADD_/FAINST[29].FA_/n1 ,
         \ADD_/FAINST[28].FA_/n3 , \ADD_/FAINST[28].FA_/n2 ,
         \ADD_/FAINST[28].FA_/n1 , \ADD_/FAINST[27].FA_/n3 ,
         \ADD_/FAINST[27].FA_/n2 , \ADD_/FAINST[27].FA_/n1 ,
         \ADD_/FAINST[26].FA_/n3 , \ADD_/FAINST[26].FA_/n2 ,
         \ADD_/FAINST[26].FA_/n1 , \ADD_/FAINST[25].FA_/n3 ,
         \ADD_/FAINST[25].FA_/n2 , \ADD_/FAINST[25].FA_/n1 ,
         \ADD_/FAINST[24].FA_/n3 , \ADD_/FAINST[24].FA_/n2 ,
         \ADD_/FAINST[24].FA_/n1 , \ADD_/FAINST[23].FA_/n3 ,
         \ADD_/FAINST[23].FA_/n2 , \ADD_/FAINST[23].FA_/n1 ,
         \ADD_/FAINST[22].FA_/n3 , \ADD_/FAINST[22].FA_/n2 ,
         \ADD_/FAINST[22].FA_/n1 , \ADD_/FAINST[21].FA_/n3 ,
         \ADD_/FAINST[21].FA_/n2 , \ADD_/FAINST[21].FA_/n1 ,
         \ADD_/FAINST[20].FA_/n3 , \ADD_/FAINST[20].FA_/n2 ,
         \ADD_/FAINST[20].FA_/n1 , \ADD_/FAINST[19].FA_/n3 ,
         \ADD_/FAINST[19].FA_/n2 , \ADD_/FAINST[19].FA_/n1 ,
         \ADD_/FAINST[18].FA_/n3 , \ADD_/FAINST[18].FA_/n2 ,
         \ADD_/FAINST[18].FA_/n1 , \ADD_/FAINST[17].FA_/n3 ,
         \ADD_/FAINST[17].FA_/n2 , \ADD_/FAINST[17].FA_/n1 ,
         \ADD_/FAINST[16].FA_/n3 , \ADD_/FAINST[16].FA_/n2 ,
         \ADD_/FAINST[16].FA_/n1 , \ADD_/FAINST[15].FA_/n3 ,
         \ADD_/FAINST[15].FA_/n2 , \ADD_/FAINST[15].FA_/n1 ,
         \ADD_/FAINST[14].FA_/n3 , \ADD_/FAINST[14].FA_/n2 ,
         \ADD_/FAINST[14].FA_/n1 , \ADD_/FAINST[13].FA_/n3 ,
         \ADD_/FAINST[13].FA_/n2 , \ADD_/FAINST[13].FA_/n1 ,
         \ADD_/FAINST[12].FA_/n3 , \ADD_/FAINST[12].FA_/n2 ,
         \ADD_/FAINST[12].FA_/n1 , \ADD_/FAINST[11].FA_/n3 ,
         \ADD_/FAINST[11].FA_/n2 , \ADD_/FAINST[11].FA_/n1 ,
         \ADD_/FAINST[10].FA_/n3 , \ADD_/FAINST[10].FA_/n2 ,
         \ADD_/FAINST[10].FA_/n1 , \ADD_/FAINST[9].FA_/n3 ,
         \ADD_/FAINST[9].FA_/n2 , \ADD_/FAINST[9].FA_/n1 ,
         \ADD_/FAINST[8].FA_/n3 , \ADD_/FAINST[8].FA_/n2 ,
         \ADD_/FAINST[8].FA_/n1 , \ADD_/FAINST[7].FA_/n3 ,
         \ADD_/FAINST[7].FA_/n2 , \ADD_/FAINST[7].FA_/n1 ,
         \ADD_/FAINST[6].FA_/n3 , \ADD_/FAINST[6].FA_/n2 ,
         \ADD_/FAINST[6].FA_/n1 , \ADD_/FAINST[5].FA_/n3 ,
         \ADD_/FAINST[5].FA_/n2 , \ADD_/FAINST[5].FA_/n1 ,
         \ADD_/FAINST[4].FA_/n3 , \ADD_/FAINST[4].FA_/n2 ,
         \ADD_/FAINST[4].FA_/n1 , \ADD_/FAINST[3].FA_/n3 ,
         \ADD_/FAINST[3].FA_/n2 , \ADD_/FAINST[3].FA_/n1 ,
         \ADD_/FAINST[2].FA_/n3 , \ADD_/FAINST[2].FA_/n2 ,
         \ADD_/FAINST[2].FA_/n1 , \ADD_/FAINST[1].FA_/n3 ,
         \ADD_/FAINST[1].FA_/n2 , \ADD_/FAINST[1].FA_/n1 ;

  DFF carry_on_reg ( .D(carry_on_d), .CLK(clk), .RST(rst), .Q(carry_on) );
  XOR \ADD_/FAINST[0].FA_/U5  ( .A(\ADD_/FAINST[0].FA_/n3 ), .B(carry_on), .Z(
        \ADD_/c[1] ) );
  XOR \ADD_/FAINST[0].FA_/U4  ( .A(\ADD_/FAINST[0].FA_/n1 ), .B(b[0]), .Z(c[0]) );
  AND \ADD_/FAINST[0].FA_/U3  ( .A(\ADD_/FAINST[0].FA_/n1 ), .B(
        \ADD_/FAINST[0].FA_/n2 ), .Z(\ADD_/FAINST[0].FA_/n3 ) );
  XOR \ADD_/FAINST[0].FA_/U2  ( .A(b[0]), .B(carry_on), .Z(
        \ADD_/FAINST[0].FA_/n2 ) );
  XOR \ADD_/FAINST[0].FA_/U1  ( .A(a[0]), .B(carry_on), .Z(
        \ADD_/FAINST[0].FA_/n1 ) );
  XOR \ADD_/FAINST[63].FA_/U5  ( .A(\ADD_/FAINST[63].FA_/n3 ), .B(\ADD_/c[63] ), .Z(carry_on_d) );
  XOR \ADD_/FAINST[63].FA_/U4  ( .A(\ADD_/FAINST[63].FA_/n1 ), .B(b[63]), .Z(
        c[63]) );
  AND \ADD_/FAINST[63].FA_/U3  ( .A(\ADD_/FAINST[63].FA_/n1 ), .B(
        \ADD_/FAINST[63].FA_/n2 ), .Z(\ADD_/FAINST[63].FA_/n3 ) );
  XOR \ADD_/FAINST[63].FA_/U2  ( .A(b[63]), .B(\ADD_/c[63] ), .Z(
        \ADD_/FAINST[63].FA_/n2 ) );
  XOR \ADD_/FAINST[63].FA_/U1  ( .A(a[63]), .B(\ADD_/c[63] ), .Z(
        \ADD_/FAINST[63].FA_/n1 ) );
  XOR \ADD_/FAINST[62].FA_/U5  ( .A(\ADD_/FAINST[62].FA_/n3 ), .B(\ADD_/c[62] ), .Z(\ADD_/c[63] ) );
  XOR \ADD_/FAINST[62].FA_/U4  ( .A(\ADD_/FAINST[62].FA_/n1 ), .B(b[62]), .Z(
        c[62]) );
  AND \ADD_/FAINST[62].FA_/U3  ( .A(\ADD_/FAINST[62].FA_/n1 ), .B(
        \ADD_/FAINST[62].FA_/n2 ), .Z(\ADD_/FAINST[62].FA_/n3 ) );
  XOR \ADD_/FAINST[62].FA_/U2  ( .A(b[62]), .B(\ADD_/c[62] ), .Z(
        \ADD_/FAINST[62].FA_/n2 ) );
  XOR \ADD_/FAINST[62].FA_/U1  ( .A(a[62]), .B(\ADD_/c[62] ), .Z(
        \ADD_/FAINST[62].FA_/n1 ) );
  XOR \ADD_/FAINST[61].FA_/U5  ( .A(\ADD_/FAINST[61].FA_/n3 ), .B(\ADD_/c[61] ), .Z(\ADD_/c[62] ) );
  XOR \ADD_/FAINST[61].FA_/U4  ( .A(\ADD_/FAINST[61].FA_/n1 ), .B(b[61]), .Z(
        c[61]) );
  AND \ADD_/FAINST[61].FA_/U3  ( .A(\ADD_/FAINST[61].FA_/n1 ), .B(
        \ADD_/FAINST[61].FA_/n2 ), .Z(\ADD_/FAINST[61].FA_/n3 ) );
  XOR \ADD_/FAINST[61].FA_/U2  ( .A(b[61]), .B(\ADD_/c[61] ), .Z(
        \ADD_/FAINST[61].FA_/n2 ) );
  XOR \ADD_/FAINST[61].FA_/U1  ( .A(a[61]), .B(\ADD_/c[61] ), .Z(
        \ADD_/FAINST[61].FA_/n1 ) );
  XOR \ADD_/FAINST[60].FA_/U5  ( .A(\ADD_/FAINST[60].FA_/n3 ), .B(\ADD_/c[60] ), .Z(\ADD_/c[61] ) );
  XOR \ADD_/FAINST[60].FA_/U4  ( .A(\ADD_/FAINST[60].FA_/n1 ), .B(b[60]), .Z(
        c[60]) );
  AND \ADD_/FAINST[60].FA_/U3  ( .A(\ADD_/FAINST[60].FA_/n1 ), .B(
        \ADD_/FAINST[60].FA_/n2 ), .Z(\ADD_/FAINST[60].FA_/n3 ) );
  XOR \ADD_/FAINST[60].FA_/U2  ( .A(b[60]), .B(\ADD_/c[60] ), .Z(
        \ADD_/FAINST[60].FA_/n2 ) );
  XOR \ADD_/FAINST[60].FA_/U1  ( .A(a[60]), .B(\ADD_/c[60] ), .Z(
        \ADD_/FAINST[60].FA_/n1 ) );
  XOR \ADD_/FAINST[59].FA_/U5  ( .A(\ADD_/FAINST[59].FA_/n3 ), .B(\ADD_/c[59] ), .Z(\ADD_/c[60] ) );
  XOR \ADD_/FAINST[59].FA_/U4  ( .A(\ADD_/FAINST[59].FA_/n1 ), .B(b[59]), .Z(
        c[59]) );
  AND \ADD_/FAINST[59].FA_/U3  ( .A(\ADD_/FAINST[59].FA_/n1 ), .B(
        \ADD_/FAINST[59].FA_/n2 ), .Z(\ADD_/FAINST[59].FA_/n3 ) );
  XOR \ADD_/FAINST[59].FA_/U2  ( .A(b[59]), .B(\ADD_/c[59] ), .Z(
        \ADD_/FAINST[59].FA_/n2 ) );
  XOR \ADD_/FAINST[59].FA_/U1  ( .A(a[59]), .B(\ADD_/c[59] ), .Z(
        \ADD_/FAINST[59].FA_/n1 ) );
  XOR \ADD_/FAINST[58].FA_/U5  ( .A(\ADD_/FAINST[58].FA_/n3 ), .B(\ADD_/c[58] ), .Z(\ADD_/c[59] ) );
  XOR \ADD_/FAINST[58].FA_/U4  ( .A(\ADD_/FAINST[58].FA_/n1 ), .B(b[58]), .Z(
        c[58]) );
  AND \ADD_/FAINST[58].FA_/U3  ( .A(\ADD_/FAINST[58].FA_/n1 ), .B(
        \ADD_/FAINST[58].FA_/n2 ), .Z(\ADD_/FAINST[58].FA_/n3 ) );
  XOR \ADD_/FAINST[58].FA_/U2  ( .A(b[58]), .B(\ADD_/c[58] ), .Z(
        \ADD_/FAINST[58].FA_/n2 ) );
  XOR \ADD_/FAINST[58].FA_/U1  ( .A(a[58]), .B(\ADD_/c[58] ), .Z(
        \ADD_/FAINST[58].FA_/n1 ) );
  XOR \ADD_/FAINST[57].FA_/U5  ( .A(\ADD_/FAINST[57].FA_/n3 ), .B(\ADD_/c[57] ), .Z(\ADD_/c[58] ) );
  XOR \ADD_/FAINST[57].FA_/U4  ( .A(\ADD_/FAINST[57].FA_/n1 ), .B(b[57]), .Z(
        c[57]) );
  AND \ADD_/FAINST[57].FA_/U3  ( .A(\ADD_/FAINST[57].FA_/n1 ), .B(
        \ADD_/FAINST[57].FA_/n2 ), .Z(\ADD_/FAINST[57].FA_/n3 ) );
  XOR \ADD_/FAINST[57].FA_/U2  ( .A(b[57]), .B(\ADD_/c[57] ), .Z(
        \ADD_/FAINST[57].FA_/n2 ) );
  XOR \ADD_/FAINST[57].FA_/U1  ( .A(a[57]), .B(\ADD_/c[57] ), .Z(
        \ADD_/FAINST[57].FA_/n1 ) );
  XOR \ADD_/FAINST[56].FA_/U5  ( .A(\ADD_/FAINST[56].FA_/n3 ), .B(\ADD_/c[56] ), .Z(\ADD_/c[57] ) );
  XOR \ADD_/FAINST[56].FA_/U4  ( .A(\ADD_/FAINST[56].FA_/n1 ), .B(b[56]), .Z(
        c[56]) );
  AND \ADD_/FAINST[56].FA_/U3  ( .A(\ADD_/FAINST[56].FA_/n1 ), .B(
        \ADD_/FAINST[56].FA_/n2 ), .Z(\ADD_/FAINST[56].FA_/n3 ) );
  XOR \ADD_/FAINST[56].FA_/U2  ( .A(b[56]), .B(\ADD_/c[56] ), .Z(
        \ADD_/FAINST[56].FA_/n2 ) );
  XOR \ADD_/FAINST[56].FA_/U1  ( .A(a[56]), .B(\ADD_/c[56] ), .Z(
        \ADD_/FAINST[56].FA_/n1 ) );
  XOR \ADD_/FAINST[55].FA_/U5  ( .A(\ADD_/FAINST[55].FA_/n3 ), .B(\ADD_/c[55] ), .Z(\ADD_/c[56] ) );
  XOR \ADD_/FAINST[55].FA_/U4  ( .A(\ADD_/FAINST[55].FA_/n1 ), .B(b[55]), .Z(
        c[55]) );
  AND \ADD_/FAINST[55].FA_/U3  ( .A(\ADD_/FAINST[55].FA_/n1 ), .B(
        \ADD_/FAINST[55].FA_/n2 ), .Z(\ADD_/FAINST[55].FA_/n3 ) );
  XOR \ADD_/FAINST[55].FA_/U2  ( .A(b[55]), .B(\ADD_/c[55] ), .Z(
        \ADD_/FAINST[55].FA_/n2 ) );
  XOR \ADD_/FAINST[55].FA_/U1  ( .A(a[55]), .B(\ADD_/c[55] ), .Z(
        \ADD_/FAINST[55].FA_/n1 ) );
  XOR \ADD_/FAINST[54].FA_/U5  ( .A(\ADD_/FAINST[54].FA_/n3 ), .B(\ADD_/c[54] ), .Z(\ADD_/c[55] ) );
  XOR \ADD_/FAINST[54].FA_/U4  ( .A(\ADD_/FAINST[54].FA_/n1 ), .B(b[54]), .Z(
        c[54]) );
  AND \ADD_/FAINST[54].FA_/U3  ( .A(\ADD_/FAINST[54].FA_/n1 ), .B(
        \ADD_/FAINST[54].FA_/n2 ), .Z(\ADD_/FAINST[54].FA_/n3 ) );
  XOR \ADD_/FAINST[54].FA_/U2  ( .A(b[54]), .B(\ADD_/c[54] ), .Z(
        \ADD_/FAINST[54].FA_/n2 ) );
  XOR \ADD_/FAINST[54].FA_/U1  ( .A(a[54]), .B(\ADD_/c[54] ), .Z(
        \ADD_/FAINST[54].FA_/n1 ) );
  XOR \ADD_/FAINST[53].FA_/U5  ( .A(\ADD_/FAINST[53].FA_/n3 ), .B(\ADD_/c[53] ), .Z(\ADD_/c[54] ) );
  XOR \ADD_/FAINST[53].FA_/U4  ( .A(\ADD_/FAINST[53].FA_/n1 ), .B(b[53]), .Z(
        c[53]) );
  AND \ADD_/FAINST[53].FA_/U3  ( .A(\ADD_/FAINST[53].FA_/n1 ), .B(
        \ADD_/FAINST[53].FA_/n2 ), .Z(\ADD_/FAINST[53].FA_/n3 ) );
  XOR \ADD_/FAINST[53].FA_/U2  ( .A(b[53]), .B(\ADD_/c[53] ), .Z(
        \ADD_/FAINST[53].FA_/n2 ) );
  XOR \ADD_/FAINST[53].FA_/U1  ( .A(a[53]), .B(\ADD_/c[53] ), .Z(
        \ADD_/FAINST[53].FA_/n1 ) );
  XOR \ADD_/FAINST[52].FA_/U5  ( .A(\ADD_/FAINST[52].FA_/n3 ), .B(\ADD_/c[52] ), .Z(\ADD_/c[53] ) );
  XOR \ADD_/FAINST[52].FA_/U4  ( .A(\ADD_/FAINST[52].FA_/n1 ), .B(b[52]), .Z(
        c[52]) );
  AND \ADD_/FAINST[52].FA_/U3  ( .A(\ADD_/FAINST[52].FA_/n1 ), .B(
        \ADD_/FAINST[52].FA_/n2 ), .Z(\ADD_/FAINST[52].FA_/n3 ) );
  XOR \ADD_/FAINST[52].FA_/U2  ( .A(b[52]), .B(\ADD_/c[52] ), .Z(
        \ADD_/FAINST[52].FA_/n2 ) );
  XOR \ADD_/FAINST[52].FA_/U1  ( .A(a[52]), .B(\ADD_/c[52] ), .Z(
        \ADD_/FAINST[52].FA_/n1 ) );
  XOR \ADD_/FAINST[51].FA_/U5  ( .A(\ADD_/FAINST[51].FA_/n3 ), .B(\ADD_/c[51] ), .Z(\ADD_/c[52] ) );
  XOR \ADD_/FAINST[51].FA_/U4  ( .A(\ADD_/FAINST[51].FA_/n1 ), .B(b[51]), .Z(
        c[51]) );
  AND \ADD_/FAINST[51].FA_/U3  ( .A(\ADD_/FAINST[51].FA_/n1 ), .B(
        \ADD_/FAINST[51].FA_/n2 ), .Z(\ADD_/FAINST[51].FA_/n3 ) );
  XOR \ADD_/FAINST[51].FA_/U2  ( .A(b[51]), .B(\ADD_/c[51] ), .Z(
        \ADD_/FAINST[51].FA_/n2 ) );
  XOR \ADD_/FAINST[51].FA_/U1  ( .A(a[51]), .B(\ADD_/c[51] ), .Z(
        \ADD_/FAINST[51].FA_/n1 ) );
  XOR \ADD_/FAINST[50].FA_/U5  ( .A(\ADD_/FAINST[50].FA_/n3 ), .B(\ADD_/c[50] ), .Z(\ADD_/c[51] ) );
  XOR \ADD_/FAINST[50].FA_/U4  ( .A(\ADD_/FAINST[50].FA_/n1 ), .B(b[50]), .Z(
        c[50]) );
  AND \ADD_/FAINST[50].FA_/U3  ( .A(\ADD_/FAINST[50].FA_/n1 ), .B(
        \ADD_/FAINST[50].FA_/n2 ), .Z(\ADD_/FAINST[50].FA_/n3 ) );
  XOR \ADD_/FAINST[50].FA_/U2  ( .A(b[50]), .B(\ADD_/c[50] ), .Z(
        \ADD_/FAINST[50].FA_/n2 ) );
  XOR \ADD_/FAINST[50].FA_/U1  ( .A(a[50]), .B(\ADD_/c[50] ), .Z(
        \ADD_/FAINST[50].FA_/n1 ) );
  XOR \ADD_/FAINST[49].FA_/U5  ( .A(\ADD_/FAINST[49].FA_/n3 ), .B(\ADD_/c[49] ), .Z(\ADD_/c[50] ) );
  XOR \ADD_/FAINST[49].FA_/U4  ( .A(\ADD_/FAINST[49].FA_/n1 ), .B(b[49]), .Z(
        c[49]) );
  AND \ADD_/FAINST[49].FA_/U3  ( .A(\ADD_/FAINST[49].FA_/n1 ), .B(
        \ADD_/FAINST[49].FA_/n2 ), .Z(\ADD_/FAINST[49].FA_/n3 ) );
  XOR \ADD_/FAINST[49].FA_/U2  ( .A(b[49]), .B(\ADD_/c[49] ), .Z(
        \ADD_/FAINST[49].FA_/n2 ) );
  XOR \ADD_/FAINST[49].FA_/U1  ( .A(a[49]), .B(\ADD_/c[49] ), .Z(
        \ADD_/FAINST[49].FA_/n1 ) );
  XOR \ADD_/FAINST[48].FA_/U5  ( .A(\ADD_/FAINST[48].FA_/n3 ), .B(\ADD_/c[48] ), .Z(\ADD_/c[49] ) );
  XOR \ADD_/FAINST[48].FA_/U4  ( .A(\ADD_/FAINST[48].FA_/n1 ), .B(b[48]), .Z(
        c[48]) );
  AND \ADD_/FAINST[48].FA_/U3  ( .A(\ADD_/FAINST[48].FA_/n1 ), .B(
        \ADD_/FAINST[48].FA_/n2 ), .Z(\ADD_/FAINST[48].FA_/n3 ) );
  XOR \ADD_/FAINST[48].FA_/U2  ( .A(b[48]), .B(\ADD_/c[48] ), .Z(
        \ADD_/FAINST[48].FA_/n2 ) );
  XOR \ADD_/FAINST[48].FA_/U1  ( .A(a[48]), .B(\ADD_/c[48] ), .Z(
        \ADD_/FAINST[48].FA_/n1 ) );
  XOR \ADD_/FAINST[47].FA_/U5  ( .A(\ADD_/FAINST[47].FA_/n3 ), .B(\ADD_/c[47] ), .Z(\ADD_/c[48] ) );
  XOR \ADD_/FAINST[47].FA_/U4  ( .A(\ADD_/FAINST[47].FA_/n1 ), .B(b[47]), .Z(
        c[47]) );
  AND \ADD_/FAINST[47].FA_/U3  ( .A(\ADD_/FAINST[47].FA_/n1 ), .B(
        \ADD_/FAINST[47].FA_/n2 ), .Z(\ADD_/FAINST[47].FA_/n3 ) );
  XOR \ADD_/FAINST[47].FA_/U2  ( .A(b[47]), .B(\ADD_/c[47] ), .Z(
        \ADD_/FAINST[47].FA_/n2 ) );
  XOR \ADD_/FAINST[47].FA_/U1  ( .A(a[47]), .B(\ADD_/c[47] ), .Z(
        \ADD_/FAINST[47].FA_/n1 ) );
  XOR \ADD_/FAINST[46].FA_/U5  ( .A(\ADD_/FAINST[46].FA_/n3 ), .B(\ADD_/c[46] ), .Z(\ADD_/c[47] ) );
  XOR \ADD_/FAINST[46].FA_/U4  ( .A(\ADD_/FAINST[46].FA_/n1 ), .B(b[46]), .Z(
        c[46]) );
  AND \ADD_/FAINST[46].FA_/U3  ( .A(\ADD_/FAINST[46].FA_/n1 ), .B(
        \ADD_/FAINST[46].FA_/n2 ), .Z(\ADD_/FAINST[46].FA_/n3 ) );
  XOR \ADD_/FAINST[46].FA_/U2  ( .A(b[46]), .B(\ADD_/c[46] ), .Z(
        \ADD_/FAINST[46].FA_/n2 ) );
  XOR \ADD_/FAINST[46].FA_/U1  ( .A(a[46]), .B(\ADD_/c[46] ), .Z(
        \ADD_/FAINST[46].FA_/n1 ) );
  XOR \ADD_/FAINST[45].FA_/U5  ( .A(\ADD_/FAINST[45].FA_/n3 ), .B(\ADD_/c[45] ), .Z(\ADD_/c[46] ) );
  XOR \ADD_/FAINST[45].FA_/U4  ( .A(\ADD_/FAINST[45].FA_/n1 ), .B(b[45]), .Z(
        c[45]) );
  AND \ADD_/FAINST[45].FA_/U3  ( .A(\ADD_/FAINST[45].FA_/n1 ), .B(
        \ADD_/FAINST[45].FA_/n2 ), .Z(\ADD_/FAINST[45].FA_/n3 ) );
  XOR \ADD_/FAINST[45].FA_/U2  ( .A(b[45]), .B(\ADD_/c[45] ), .Z(
        \ADD_/FAINST[45].FA_/n2 ) );
  XOR \ADD_/FAINST[45].FA_/U1  ( .A(a[45]), .B(\ADD_/c[45] ), .Z(
        \ADD_/FAINST[45].FA_/n1 ) );
  XOR \ADD_/FAINST[44].FA_/U5  ( .A(\ADD_/FAINST[44].FA_/n3 ), .B(\ADD_/c[44] ), .Z(\ADD_/c[45] ) );
  XOR \ADD_/FAINST[44].FA_/U4  ( .A(\ADD_/FAINST[44].FA_/n1 ), .B(b[44]), .Z(
        c[44]) );
  AND \ADD_/FAINST[44].FA_/U3  ( .A(\ADD_/FAINST[44].FA_/n1 ), .B(
        \ADD_/FAINST[44].FA_/n2 ), .Z(\ADD_/FAINST[44].FA_/n3 ) );
  XOR \ADD_/FAINST[44].FA_/U2  ( .A(b[44]), .B(\ADD_/c[44] ), .Z(
        \ADD_/FAINST[44].FA_/n2 ) );
  XOR \ADD_/FAINST[44].FA_/U1  ( .A(a[44]), .B(\ADD_/c[44] ), .Z(
        \ADD_/FAINST[44].FA_/n1 ) );
  XOR \ADD_/FAINST[43].FA_/U5  ( .A(\ADD_/FAINST[43].FA_/n3 ), .B(\ADD_/c[43] ), .Z(\ADD_/c[44] ) );
  XOR \ADD_/FAINST[43].FA_/U4  ( .A(\ADD_/FAINST[43].FA_/n1 ), .B(b[43]), .Z(
        c[43]) );
  AND \ADD_/FAINST[43].FA_/U3  ( .A(\ADD_/FAINST[43].FA_/n1 ), .B(
        \ADD_/FAINST[43].FA_/n2 ), .Z(\ADD_/FAINST[43].FA_/n3 ) );
  XOR \ADD_/FAINST[43].FA_/U2  ( .A(b[43]), .B(\ADD_/c[43] ), .Z(
        \ADD_/FAINST[43].FA_/n2 ) );
  XOR \ADD_/FAINST[43].FA_/U1  ( .A(a[43]), .B(\ADD_/c[43] ), .Z(
        \ADD_/FAINST[43].FA_/n1 ) );
  XOR \ADD_/FAINST[42].FA_/U5  ( .A(\ADD_/FAINST[42].FA_/n3 ), .B(\ADD_/c[42] ), .Z(\ADD_/c[43] ) );
  XOR \ADD_/FAINST[42].FA_/U4  ( .A(\ADD_/FAINST[42].FA_/n1 ), .B(b[42]), .Z(
        c[42]) );
  AND \ADD_/FAINST[42].FA_/U3  ( .A(\ADD_/FAINST[42].FA_/n1 ), .B(
        \ADD_/FAINST[42].FA_/n2 ), .Z(\ADD_/FAINST[42].FA_/n3 ) );
  XOR \ADD_/FAINST[42].FA_/U2  ( .A(b[42]), .B(\ADD_/c[42] ), .Z(
        \ADD_/FAINST[42].FA_/n2 ) );
  XOR \ADD_/FAINST[42].FA_/U1  ( .A(a[42]), .B(\ADD_/c[42] ), .Z(
        \ADD_/FAINST[42].FA_/n1 ) );
  XOR \ADD_/FAINST[41].FA_/U5  ( .A(\ADD_/FAINST[41].FA_/n3 ), .B(\ADD_/c[41] ), .Z(\ADD_/c[42] ) );
  XOR \ADD_/FAINST[41].FA_/U4  ( .A(\ADD_/FAINST[41].FA_/n1 ), .B(b[41]), .Z(
        c[41]) );
  AND \ADD_/FAINST[41].FA_/U3  ( .A(\ADD_/FAINST[41].FA_/n1 ), .B(
        \ADD_/FAINST[41].FA_/n2 ), .Z(\ADD_/FAINST[41].FA_/n3 ) );
  XOR \ADD_/FAINST[41].FA_/U2  ( .A(b[41]), .B(\ADD_/c[41] ), .Z(
        \ADD_/FAINST[41].FA_/n2 ) );
  XOR \ADD_/FAINST[41].FA_/U1  ( .A(a[41]), .B(\ADD_/c[41] ), .Z(
        \ADD_/FAINST[41].FA_/n1 ) );
  XOR \ADD_/FAINST[40].FA_/U5  ( .A(\ADD_/FAINST[40].FA_/n3 ), .B(\ADD_/c[40] ), .Z(\ADD_/c[41] ) );
  XOR \ADD_/FAINST[40].FA_/U4  ( .A(\ADD_/FAINST[40].FA_/n1 ), .B(b[40]), .Z(
        c[40]) );
  AND \ADD_/FAINST[40].FA_/U3  ( .A(\ADD_/FAINST[40].FA_/n1 ), .B(
        \ADD_/FAINST[40].FA_/n2 ), .Z(\ADD_/FAINST[40].FA_/n3 ) );
  XOR \ADD_/FAINST[40].FA_/U2  ( .A(b[40]), .B(\ADD_/c[40] ), .Z(
        \ADD_/FAINST[40].FA_/n2 ) );
  XOR \ADD_/FAINST[40].FA_/U1  ( .A(a[40]), .B(\ADD_/c[40] ), .Z(
        \ADD_/FAINST[40].FA_/n1 ) );
  XOR \ADD_/FAINST[39].FA_/U5  ( .A(\ADD_/FAINST[39].FA_/n3 ), .B(\ADD_/c[39] ), .Z(\ADD_/c[40] ) );
  XOR \ADD_/FAINST[39].FA_/U4  ( .A(\ADD_/FAINST[39].FA_/n1 ), .B(b[39]), .Z(
        c[39]) );
  AND \ADD_/FAINST[39].FA_/U3  ( .A(\ADD_/FAINST[39].FA_/n1 ), .B(
        \ADD_/FAINST[39].FA_/n2 ), .Z(\ADD_/FAINST[39].FA_/n3 ) );
  XOR \ADD_/FAINST[39].FA_/U2  ( .A(b[39]), .B(\ADD_/c[39] ), .Z(
        \ADD_/FAINST[39].FA_/n2 ) );
  XOR \ADD_/FAINST[39].FA_/U1  ( .A(a[39]), .B(\ADD_/c[39] ), .Z(
        \ADD_/FAINST[39].FA_/n1 ) );
  XOR \ADD_/FAINST[38].FA_/U5  ( .A(\ADD_/FAINST[38].FA_/n3 ), .B(\ADD_/c[38] ), .Z(\ADD_/c[39] ) );
  XOR \ADD_/FAINST[38].FA_/U4  ( .A(\ADD_/FAINST[38].FA_/n1 ), .B(b[38]), .Z(
        c[38]) );
  AND \ADD_/FAINST[38].FA_/U3  ( .A(\ADD_/FAINST[38].FA_/n1 ), .B(
        \ADD_/FAINST[38].FA_/n2 ), .Z(\ADD_/FAINST[38].FA_/n3 ) );
  XOR \ADD_/FAINST[38].FA_/U2  ( .A(b[38]), .B(\ADD_/c[38] ), .Z(
        \ADD_/FAINST[38].FA_/n2 ) );
  XOR \ADD_/FAINST[38].FA_/U1  ( .A(a[38]), .B(\ADD_/c[38] ), .Z(
        \ADD_/FAINST[38].FA_/n1 ) );
  XOR \ADD_/FAINST[37].FA_/U5  ( .A(\ADD_/FAINST[37].FA_/n3 ), .B(\ADD_/c[37] ), .Z(\ADD_/c[38] ) );
  XOR \ADD_/FAINST[37].FA_/U4  ( .A(\ADD_/FAINST[37].FA_/n1 ), .B(b[37]), .Z(
        c[37]) );
  AND \ADD_/FAINST[37].FA_/U3  ( .A(\ADD_/FAINST[37].FA_/n1 ), .B(
        \ADD_/FAINST[37].FA_/n2 ), .Z(\ADD_/FAINST[37].FA_/n3 ) );
  XOR \ADD_/FAINST[37].FA_/U2  ( .A(b[37]), .B(\ADD_/c[37] ), .Z(
        \ADD_/FAINST[37].FA_/n2 ) );
  XOR \ADD_/FAINST[37].FA_/U1  ( .A(a[37]), .B(\ADD_/c[37] ), .Z(
        \ADD_/FAINST[37].FA_/n1 ) );
  XOR \ADD_/FAINST[36].FA_/U5  ( .A(\ADD_/FAINST[36].FA_/n3 ), .B(\ADD_/c[36] ), .Z(\ADD_/c[37] ) );
  XOR \ADD_/FAINST[36].FA_/U4  ( .A(\ADD_/FAINST[36].FA_/n1 ), .B(b[36]), .Z(
        c[36]) );
  AND \ADD_/FAINST[36].FA_/U3  ( .A(\ADD_/FAINST[36].FA_/n1 ), .B(
        \ADD_/FAINST[36].FA_/n2 ), .Z(\ADD_/FAINST[36].FA_/n3 ) );
  XOR \ADD_/FAINST[36].FA_/U2  ( .A(b[36]), .B(\ADD_/c[36] ), .Z(
        \ADD_/FAINST[36].FA_/n2 ) );
  XOR \ADD_/FAINST[36].FA_/U1  ( .A(a[36]), .B(\ADD_/c[36] ), .Z(
        \ADD_/FAINST[36].FA_/n1 ) );
  XOR \ADD_/FAINST[35].FA_/U5  ( .A(\ADD_/FAINST[35].FA_/n3 ), .B(\ADD_/c[35] ), .Z(\ADD_/c[36] ) );
  XOR \ADD_/FAINST[35].FA_/U4  ( .A(\ADD_/FAINST[35].FA_/n1 ), .B(b[35]), .Z(
        c[35]) );
  AND \ADD_/FAINST[35].FA_/U3  ( .A(\ADD_/FAINST[35].FA_/n1 ), .B(
        \ADD_/FAINST[35].FA_/n2 ), .Z(\ADD_/FAINST[35].FA_/n3 ) );
  XOR \ADD_/FAINST[35].FA_/U2  ( .A(b[35]), .B(\ADD_/c[35] ), .Z(
        \ADD_/FAINST[35].FA_/n2 ) );
  XOR \ADD_/FAINST[35].FA_/U1  ( .A(a[35]), .B(\ADD_/c[35] ), .Z(
        \ADD_/FAINST[35].FA_/n1 ) );
  XOR \ADD_/FAINST[34].FA_/U5  ( .A(\ADD_/FAINST[34].FA_/n3 ), .B(\ADD_/c[34] ), .Z(\ADD_/c[35] ) );
  XOR \ADD_/FAINST[34].FA_/U4  ( .A(\ADD_/FAINST[34].FA_/n1 ), .B(b[34]), .Z(
        c[34]) );
  AND \ADD_/FAINST[34].FA_/U3  ( .A(\ADD_/FAINST[34].FA_/n1 ), .B(
        \ADD_/FAINST[34].FA_/n2 ), .Z(\ADD_/FAINST[34].FA_/n3 ) );
  XOR \ADD_/FAINST[34].FA_/U2  ( .A(b[34]), .B(\ADD_/c[34] ), .Z(
        \ADD_/FAINST[34].FA_/n2 ) );
  XOR \ADD_/FAINST[34].FA_/U1  ( .A(a[34]), .B(\ADD_/c[34] ), .Z(
        \ADD_/FAINST[34].FA_/n1 ) );
  XOR \ADD_/FAINST[33].FA_/U5  ( .A(\ADD_/FAINST[33].FA_/n3 ), .B(\ADD_/c[33] ), .Z(\ADD_/c[34] ) );
  XOR \ADD_/FAINST[33].FA_/U4  ( .A(\ADD_/FAINST[33].FA_/n1 ), .B(b[33]), .Z(
        c[33]) );
  AND \ADD_/FAINST[33].FA_/U3  ( .A(\ADD_/FAINST[33].FA_/n1 ), .B(
        \ADD_/FAINST[33].FA_/n2 ), .Z(\ADD_/FAINST[33].FA_/n3 ) );
  XOR \ADD_/FAINST[33].FA_/U2  ( .A(b[33]), .B(\ADD_/c[33] ), .Z(
        \ADD_/FAINST[33].FA_/n2 ) );
  XOR \ADD_/FAINST[33].FA_/U1  ( .A(a[33]), .B(\ADD_/c[33] ), .Z(
        \ADD_/FAINST[33].FA_/n1 ) );
  XOR \ADD_/FAINST[32].FA_/U5  ( .A(\ADD_/FAINST[32].FA_/n3 ), .B(\ADD_/c[32] ), .Z(\ADD_/c[33] ) );
  XOR \ADD_/FAINST[32].FA_/U4  ( .A(\ADD_/FAINST[32].FA_/n1 ), .B(b[32]), .Z(
        c[32]) );
  AND \ADD_/FAINST[32].FA_/U3  ( .A(\ADD_/FAINST[32].FA_/n1 ), .B(
        \ADD_/FAINST[32].FA_/n2 ), .Z(\ADD_/FAINST[32].FA_/n3 ) );
  XOR \ADD_/FAINST[32].FA_/U2  ( .A(b[32]), .B(\ADD_/c[32] ), .Z(
        \ADD_/FAINST[32].FA_/n2 ) );
  XOR \ADD_/FAINST[32].FA_/U1  ( .A(a[32]), .B(\ADD_/c[32] ), .Z(
        \ADD_/FAINST[32].FA_/n1 ) );
  XOR \ADD_/FAINST[31].FA_/U5  ( .A(\ADD_/FAINST[31].FA_/n3 ), .B(\ADD_/c[31] ), .Z(\ADD_/c[32] ) );
  XOR \ADD_/FAINST[31].FA_/U4  ( .A(\ADD_/FAINST[31].FA_/n1 ), .B(b[31]), .Z(
        c[31]) );
  AND \ADD_/FAINST[31].FA_/U3  ( .A(\ADD_/FAINST[31].FA_/n1 ), .B(
        \ADD_/FAINST[31].FA_/n2 ), .Z(\ADD_/FAINST[31].FA_/n3 ) );
  XOR \ADD_/FAINST[31].FA_/U2  ( .A(b[31]), .B(\ADD_/c[31] ), .Z(
        \ADD_/FAINST[31].FA_/n2 ) );
  XOR \ADD_/FAINST[31].FA_/U1  ( .A(a[31]), .B(\ADD_/c[31] ), .Z(
        \ADD_/FAINST[31].FA_/n1 ) );
  XOR \ADD_/FAINST[30].FA_/U5  ( .A(\ADD_/FAINST[30].FA_/n3 ), .B(\ADD_/c[30] ), .Z(\ADD_/c[31] ) );
  XOR \ADD_/FAINST[30].FA_/U4  ( .A(\ADD_/FAINST[30].FA_/n1 ), .B(b[30]), .Z(
        c[30]) );
  AND \ADD_/FAINST[30].FA_/U3  ( .A(\ADD_/FAINST[30].FA_/n1 ), .B(
        \ADD_/FAINST[30].FA_/n2 ), .Z(\ADD_/FAINST[30].FA_/n3 ) );
  XOR \ADD_/FAINST[30].FA_/U2  ( .A(b[30]), .B(\ADD_/c[30] ), .Z(
        \ADD_/FAINST[30].FA_/n2 ) );
  XOR \ADD_/FAINST[30].FA_/U1  ( .A(a[30]), .B(\ADD_/c[30] ), .Z(
        \ADD_/FAINST[30].FA_/n1 ) );
  XOR \ADD_/FAINST[29].FA_/U5  ( .A(\ADD_/FAINST[29].FA_/n3 ), .B(\ADD_/c[29] ), .Z(\ADD_/c[30] ) );
  XOR \ADD_/FAINST[29].FA_/U4  ( .A(\ADD_/FAINST[29].FA_/n1 ), .B(b[29]), .Z(
        c[29]) );
  AND \ADD_/FAINST[29].FA_/U3  ( .A(\ADD_/FAINST[29].FA_/n1 ), .B(
        \ADD_/FAINST[29].FA_/n2 ), .Z(\ADD_/FAINST[29].FA_/n3 ) );
  XOR \ADD_/FAINST[29].FA_/U2  ( .A(b[29]), .B(\ADD_/c[29] ), .Z(
        \ADD_/FAINST[29].FA_/n2 ) );
  XOR \ADD_/FAINST[29].FA_/U1  ( .A(a[29]), .B(\ADD_/c[29] ), .Z(
        \ADD_/FAINST[29].FA_/n1 ) );
  XOR \ADD_/FAINST[28].FA_/U5  ( .A(\ADD_/FAINST[28].FA_/n3 ), .B(\ADD_/c[28] ), .Z(\ADD_/c[29] ) );
  XOR \ADD_/FAINST[28].FA_/U4  ( .A(\ADD_/FAINST[28].FA_/n1 ), .B(b[28]), .Z(
        c[28]) );
  AND \ADD_/FAINST[28].FA_/U3  ( .A(\ADD_/FAINST[28].FA_/n1 ), .B(
        \ADD_/FAINST[28].FA_/n2 ), .Z(\ADD_/FAINST[28].FA_/n3 ) );
  XOR \ADD_/FAINST[28].FA_/U2  ( .A(b[28]), .B(\ADD_/c[28] ), .Z(
        \ADD_/FAINST[28].FA_/n2 ) );
  XOR \ADD_/FAINST[28].FA_/U1  ( .A(a[28]), .B(\ADD_/c[28] ), .Z(
        \ADD_/FAINST[28].FA_/n1 ) );
  XOR \ADD_/FAINST[27].FA_/U5  ( .A(\ADD_/FAINST[27].FA_/n3 ), .B(\ADD_/c[27] ), .Z(\ADD_/c[28] ) );
  XOR \ADD_/FAINST[27].FA_/U4  ( .A(\ADD_/FAINST[27].FA_/n1 ), .B(b[27]), .Z(
        c[27]) );
  AND \ADD_/FAINST[27].FA_/U3  ( .A(\ADD_/FAINST[27].FA_/n1 ), .B(
        \ADD_/FAINST[27].FA_/n2 ), .Z(\ADD_/FAINST[27].FA_/n3 ) );
  XOR \ADD_/FAINST[27].FA_/U2  ( .A(b[27]), .B(\ADD_/c[27] ), .Z(
        \ADD_/FAINST[27].FA_/n2 ) );
  XOR \ADD_/FAINST[27].FA_/U1  ( .A(a[27]), .B(\ADD_/c[27] ), .Z(
        \ADD_/FAINST[27].FA_/n1 ) );
  XOR \ADD_/FAINST[26].FA_/U5  ( .A(\ADD_/FAINST[26].FA_/n3 ), .B(\ADD_/c[26] ), .Z(\ADD_/c[27] ) );
  XOR \ADD_/FAINST[26].FA_/U4  ( .A(\ADD_/FAINST[26].FA_/n1 ), .B(b[26]), .Z(
        c[26]) );
  AND \ADD_/FAINST[26].FA_/U3  ( .A(\ADD_/FAINST[26].FA_/n1 ), .B(
        \ADD_/FAINST[26].FA_/n2 ), .Z(\ADD_/FAINST[26].FA_/n3 ) );
  XOR \ADD_/FAINST[26].FA_/U2  ( .A(b[26]), .B(\ADD_/c[26] ), .Z(
        \ADD_/FAINST[26].FA_/n2 ) );
  XOR \ADD_/FAINST[26].FA_/U1  ( .A(a[26]), .B(\ADD_/c[26] ), .Z(
        \ADD_/FAINST[26].FA_/n1 ) );
  XOR \ADD_/FAINST[25].FA_/U5  ( .A(\ADD_/FAINST[25].FA_/n3 ), .B(\ADD_/c[25] ), .Z(\ADD_/c[26] ) );
  XOR \ADD_/FAINST[25].FA_/U4  ( .A(\ADD_/FAINST[25].FA_/n1 ), .B(b[25]), .Z(
        c[25]) );
  AND \ADD_/FAINST[25].FA_/U3  ( .A(\ADD_/FAINST[25].FA_/n1 ), .B(
        \ADD_/FAINST[25].FA_/n2 ), .Z(\ADD_/FAINST[25].FA_/n3 ) );
  XOR \ADD_/FAINST[25].FA_/U2  ( .A(b[25]), .B(\ADD_/c[25] ), .Z(
        \ADD_/FAINST[25].FA_/n2 ) );
  XOR \ADD_/FAINST[25].FA_/U1  ( .A(a[25]), .B(\ADD_/c[25] ), .Z(
        \ADD_/FAINST[25].FA_/n1 ) );
  XOR \ADD_/FAINST[24].FA_/U5  ( .A(\ADD_/FAINST[24].FA_/n3 ), .B(\ADD_/c[24] ), .Z(\ADD_/c[25] ) );
  XOR \ADD_/FAINST[24].FA_/U4  ( .A(\ADD_/FAINST[24].FA_/n1 ), .B(b[24]), .Z(
        c[24]) );
  AND \ADD_/FAINST[24].FA_/U3  ( .A(\ADD_/FAINST[24].FA_/n1 ), .B(
        \ADD_/FAINST[24].FA_/n2 ), .Z(\ADD_/FAINST[24].FA_/n3 ) );
  XOR \ADD_/FAINST[24].FA_/U2  ( .A(b[24]), .B(\ADD_/c[24] ), .Z(
        \ADD_/FAINST[24].FA_/n2 ) );
  XOR \ADD_/FAINST[24].FA_/U1  ( .A(a[24]), .B(\ADD_/c[24] ), .Z(
        \ADD_/FAINST[24].FA_/n1 ) );
  XOR \ADD_/FAINST[23].FA_/U5  ( .A(\ADD_/FAINST[23].FA_/n3 ), .B(\ADD_/c[23] ), .Z(\ADD_/c[24] ) );
  XOR \ADD_/FAINST[23].FA_/U4  ( .A(\ADD_/FAINST[23].FA_/n1 ), .B(b[23]), .Z(
        c[23]) );
  AND \ADD_/FAINST[23].FA_/U3  ( .A(\ADD_/FAINST[23].FA_/n1 ), .B(
        \ADD_/FAINST[23].FA_/n2 ), .Z(\ADD_/FAINST[23].FA_/n3 ) );
  XOR \ADD_/FAINST[23].FA_/U2  ( .A(b[23]), .B(\ADD_/c[23] ), .Z(
        \ADD_/FAINST[23].FA_/n2 ) );
  XOR \ADD_/FAINST[23].FA_/U1  ( .A(a[23]), .B(\ADD_/c[23] ), .Z(
        \ADD_/FAINST[23].FA_/n1 ) );
  XOR \ADD_/FAINST[22].FA_/U5  ( .A(\ADD_/FAINST[22].FA_/n3 ), .B(\ADD_/c[22] ), .Z(\ADD_/c[23] ) );
  XOR \ADD_/FAINST[22].FA_/U4  ( .A(\ADD_/FAINST[22].FA_/n1 ), .B(b[22]), .Z(
        c[22]) );
  AND \ADD_/FAINST[22].FA_/U3  ( .A(\ADD_/FAINST[22].FA_/n1 ), .B(
        \ADD_/FAINST[22].FA_/n2 ), .Z(\ADD_/FAINST[22].FA_/n3 ) );
  XOR \ADD_/FAINST[22].FA_/U2  ( .A(b[22]), .B(\ADD_/c[22] ), .Z(
        \ADD_/FAINST[22].FA_/n2 ) );
  XOR \ADD_/FAINST[22].FA_/U1  ( .A(a[22]), .B(\ADD_/c[22] ), .Z(
        \ADD_/FAINST[22].FA_/n1 ) );
  XOR \ADD_/FAINST[21].FA_/U5  ( .A(\ADD_/FAINST[21].FA_/n3 ), .B(\ADD_/c[21] ), .Z(\ADD_/c[22] ) );
  XOR \ADD_/FAINST[21].FA_/U4  ( .A(\ADD_/FAINST[21].FA_/n1 ), .B(b[21]), .Z(
        c[21]) );
  AND \ADD_/FAINST[21].FA_/U3  ( .A(\ADD_/FAINST[21].FA_/n1 ), .B(
        \ADD_/FAINST[21].FA_/n2 ), .Z(\ADD_/FAINST[21].FA_/n3 ) );
  XOR \ADD_/FAINST[21].FA_/U2  ( .A(b[21]), .B(\ADD_/c[21] ), .Z(
        \ADD_/FAINST[21].FA_/n2 ) );
  XOR \ADD_/FAINST[21].FA_/U1  ( .A(a[21]), .B(\ADD_/c[21] ), .Z(
        \ADD_/FAINST[21].FA_/n1 ) );
  XOR \ADD_/FAINST[20].FA_/U5  ( .A(\ADD_/FAINST[20].FA_/n3 ), .B(\ADD_/c[20] ), .Z(\ADD_/c[21] ) );
  XOR \ADD_/FAINST[20].FA_/U4  ( .A(\ADD_/FAINST[20].FA_/n1 ), .B(b[20]), .Z(
        c[20]) );
  AND \ADD_/FAINST[20].FA_/U3  ( .A(\ADD_/FAINST[20].FA_/n1 ), .B(
        \ADD_/FAINST[20].FA_/n2 ), .Z(\ADD_/FAINST[20].FA_/n3 ) );
  XOR \ADD_/FAINST[20].FA_/U2  ( .A(b[20]), .B(\ADD_/c[20] ), .Z(
        \ADD_/FAINST[20].FA_/n2 ) );
  XOR \ADD_/FAINST[20].FA_/U1  ( .A(a[20]), .B(\ADD_/c[20] ), .Z(
        \ADD_/FAINST[20].FA_/n1 ) );
  XOR \ADD_/FAINST[19].FA_/U5  ( .A(\ADD_/FAINST[19].FA_/n3 ), .B(\ADD_/c[19] ), .Z(\ADD_/c[20] ) );
  XOR \ADD_/FAINST[19].FA_/U4  ( .A(\ADD_/FAINST[19].FA_/n1 ), .B(b[19]), .Z(
        c[19]) );
  AND \ADD_/FAINST[19].FA_/U3  ( .A(\ADD_/FAINST[19].FA_/n1 ), .B(
        \ADD_/FAINST[19].FA_/n2 ), .Z(\ADD_/FAINST[19].FA_/n3 ) );
  XOR \ADD_/FAINST[19].FA_/U2  ( .A(b[19]), .B(\ADD_/c[19] ), .Z(
        \ADD_/FAINST[19].FA_/n2 ) );
  XOR \ADD_/FAINST[19].FA_/U1  ( .A(a[19]), .B(\ADD_/c[19] ), .Z(
        \ADD_/FAINST[19].FA_/n1 ) );
  XOR \ADD_/FAINST[18].FA_/U5  ( .A(\ADD_/FAINST[18].FA_/n3 ), .B(\ADD_/c[18] ), .Z(\ADD_/c[19] ) );
  XOR \ADD_/FAINST[18].FA_/U4  ( .A(\ADD_/FAINST[18].FA_/n1 ), .B(b[18]), .Z(
        c[18]) );
  AND \ADD_/FAINST[18].FA_/U3  ( .A(\ADD_/FAINST[18].FA_/n1 ), .B(
        \ADD_/FAINST[18].FA_/n2 ), .Z(\ADD_/FAINST[18].FA_/n3 ) );
  XOR \ADD_/FAINST[18].FA_/U2  ( .A(b[18]), .B(\ADD_/c[18] ), .Z(
        \ADD_/FAINST[18].FA_/n2 ) );
  XOR \ADD_/FAINST[18].FA_/U1  ( .A(a[18]), .B(\ADD_/c[18] ), .Z(
        \ADD_/FAINST[18].FA_/n1 ) );
  XOR \ADD_/FAINST[17].FA_/U5  ( .A(\ADD_/FAINST[17].FA_/n3 ), .B(\ADD_/c[17] ), .Z(\ADD_/c[18] ) );
  XOR \ADD_/FAINST[17].FA_/U4  ( .A(\ADD_/FAINST[17].FA_/n1 ), .B(b[17]), .Z(
        c[17]) );
  AND \ADD_/FAINST[17].FA_/U3  ( .A(\ADD_/FAINST[17].FA_/n1 ), .B(
        \ADD_/FAINST[17].FA_/n2 ), .Z(\ADD_/FAINST[17].FA_/n3 ) );
  XOR \ADD_/FAINST[17].FA_/U2  ( .A(b[17]), .B(\ADD_/c[17] ), .Z(
        \ADD_/FAINST[17].FA_/n2 ) );
  XOR \ADD_/FAINST[17].FA_/U1  ( .A(a[17]), .B(\ADD_/c[17] ), .Z(
        \ADD_/FAINST[17].FA_/n1 ) );
  XOR \ADD_/FAINST[16].FA_/U5  ( .A(\ADD_/FAINST[16].FA_/n3 ), .B(\ADD_/c[16] ), .Z(\ADD_/c[17] ) );
  XOR \ADD_/FAINST[16].FA_/U4  ( .A(\ADD_/FAINST[16].FA_/n1 ), .B(b[16]), .Z(
        c[16]) );
  AND \ADD_/FAINST[16].FA_/U3  ( .A(\ADD_/FAINST[16].FA_/n1 ), .B(
        \ADD_/FAINST[16].FA_/n2 ), .Z(\ADD_/FAINST[16].FA_/n3 ) );
  XOR \ADD_/FAINST[16].FA_/U2  ( .A(b[16]), .B(\ADD_/c[16] ), .Z(
        \ADD_/FAINST[16].FA_/n2 ) );
  XOR \ADD_/FAINST[16].FA_/U1  ( .A(a[16]), .B(\ADD_/c[16] ), .Z(
        \ADD_/FAINST[16].FA_/n1 ) );
  XOR \ADD_/FAINST[15].FA_/U5  ( .A(\ADD_/FAINST[15].FA_/n3 ), .B(\ADD_/c[15] ), .Z(\ADD_/c[16] ) );
  XOR \ADD_/FAINST[15].FA_/U4  ( .A(\ADD_/FAINST[15].FA_/n1 ), .B(b[15]), .Z(
        c[15]) );
  AND \ADD_/FAINST[15].FA_/U3  ( .A(\ADD_/FAINST[15].FA_/n1 ), .B(
        \ADD_/FAINST[15].FA_/n2 ), .Z(\ADD_/FAINST[15].FA_/n3 ) );
  XOR \ADD_/FAINST[15].FA_/U2  ( .A(b[15]), .B(\ADD_/c[15] ), .Z(
        \ADD_/FAINST[15].FA_/n2 ) );
  XOR \ADD_/FAINST[15].FA_/U1  ( .A(a[15]), .B(\ADD_/c[15] ), .Z(
        \ADD_/FAINST[15].FA_/n1 ) );
  XOR \ADD_/FAINST[14].FA_/U5  ( .A(\ADD_/FAINST[14].FA_/n3 ), .B(\ADD_/c[14] ), .Z(\ADD_/c[15] ) );
  XOR \ADD_/FAINST[14].FA_/U4  ( .A(\ADD_/FAINST[14].FA_/n1 ), .B(b[14]), .Z(
        c[14]) );
  AND \ADD_/FAINST[14].FA_/U3  ( .A(\ADD_/FAINST[14].FA_/n1 ), .B(
        \ADD_/FAINST[14].FA_/n2 ), .Z(\ADD_/FAINST[14].FA_/n3 ) );
  XOR \ADD_/FAINST[14].FA_/U2  ( .A(b[14]), .B(\ADD_/c[14] ), .Z(
        \ADD_/FAINST[14].FA_/n2 ) );
  XOR \ADD_/FAINST[14].FA_/U1  ( .A(a[14]), .B(\ADD_/c[14] ), .Z(
        \ADD_/FAINST[14].FA_/n1 ) );
  XOR \ADD_/FAINST[13].FA_/U5  ( .A(\ADD_/FAINST[13].FA_/n3 ), .B(\ADD_/c[13] ), .Z(\ADD_/c[14] ) );
  XOR \ADD_/FAINST[13].FA_/U4  ( .A(\ADD_/FAINST[13].FA_/n1 ), .B(b[13]), .Z(
        c[13]) );
  AND \ADD_/FAINST[13].FA_/U3  ( .A(\ADD_/FAINST[13].FA_/n1 ), .B(
        \ADD_/FAINST[13].FA_/n2 ), .Z(\ADD_/FAINST[13].FA_/n3 ) );
  XOR \ADD_/FAINST[13].FA_/U2  ( .A(b[13]), .B(\ADD_/c[13] ), .Z(
        \ADD_/FAINST[13].FA_/n2 ) );
  XOR \ADD_/FAINST[13].FA_/U1  ( .A(a[13]), .B(\ADD_/c[13] ), .Z(
        \ADD_/FAINST[13].FA_/n1 ) );
  XOR \ADD_/FAINST[12].FA_/U5  ( .A(\ADD_/FAINST[12].FA_/n3 ), .B(\ADD_/c[12] ), .Z(\ADD_/c[13] ) );
  XOR \ADD_/FAINST[12].FA_/U4  ( .A(\ADD_/FAINST[12].FA_/n1 ), .B(b[12]), .Z(
        c[12]) );
  AND \ADD_/FAINST[12].FA_/U3  ( .A(\ADD_/FAINST[12].FA_/n1 ), .B(
        \ADD_/FAINST[12].FA_/n2 ), .Z(\ADD_/FAINST[12].FA_/n3 ) );
  XOR \ADD_/FAINST[12].FA_/U2  ( .A(b[12]), .B(\ADD_/c[12] ), .Z(
        \ADD_/FAINST[12].FA_/n2 ) );
  XOR \ADD_/FAINST[12].FA_/U1  ( .A(a[12]), .B(\ADD_/c[12] ), .Z(
        \ADD_/FAINST[12].FA_/n1 ) );
  XOR \ADD_/FAINST[11].FA_/U5  ( .A(\ADD_/FAINST[11].FA_/n3 ), .B(\ADD_/c[11] ), .Z(\ADD_/c[12] ) );
  XOR \ADD_/FAINST[11].FA_/U4  ( .A(\ADD_/FAINST[11].FA_/n1 ), .B(b[11]), .Z(
        c[11]) );
  AND \ADD_/FAINST[11].FA_/U3  ( .A(\ADD_/FAINST[11].FA_/n1 ), .B(
        \ADD_/FAINST[11].FA_/n2 ), .Z(\ADD_/FAINST[11].FA_/n3 ) );
  XOR \ADD_/FAINST[11].FA_/U2  ( .A(b[11]), .B(\ADD_/c[11] ), .Z(
        \ADD_/FAINST[11].FA_/n2 ) );
  XOR \ADD_/FAINST[11].FA_/U1  ( .A(a[11]), .B(\ADD_/c[11] ), .Z(
        \ADD_/FAINST[11].FA_/n1 ) );
  XOR \ADD_/FAINST[10].FA_/U5  ( .A(\ADD_/FAINST[10].FA_/n3 ), .B(\ADD_/c[10] ), .Z(\ADD_/c[11] ) );
  XOR \ADD_/FAINST[10].FA_/U4  ( .A(\ADD_/FAINST[10].FA_/n1 ), .B(b[10]), .Z(
        c[10]) );
  AND \ADD_/FAINST[10].FA_/U3  ( .A(\ADD_/FAINST[10].FA_/n1 ), .B(
        \ADD_/FAINST[10].FA_/n2 ), .Z(\ADD_/FAINST[10].FA_/n3 ) );
  XOR \ADD_/FAINST[10].FA_/U2  ( .A(b[10]), .B(\ADD_/c[10] ), .Z(
        \ADD_/FAINST[10].FA_/n2 ) );
  XOR \ADD_/FAINST[10].FA_/U1  ( .A(a[10]), .B(\ADD_/c[10] ), .Z(
        \ADD_/FAINST[10].FA_/n1 ) );
  XOR \ADD_/FAINST[9].FA_/U5  ( .A(\ADD_/FAINST[9].FA_/n3 ), .B(\ADD_/c[9] ), 
        .Z(\ADD_/c[10] ) );
  XOR \ADD_/FAINST[9].FA_/U4  ( .A(\ADD_/FAINST[9].FA_/n1 ), .B(b[9]), .Z(c[9]) );
  AND \ADD_/FAINST[9].FA_/U3  ( .A(\ADD_/FAINST[9].FA_/n1 ), .B(
        \ADD_/FAINST[9].FA_/n2 ), .Z(\ADD_/FAINST[9].FA_/n3 ) );
  XOR \ADD_/FAINST[9].FA_/U2  ( .A(b[9]), .B(\ADD_/c[9] ), .Z(
        \ADD_/FAINST[9].FA_/n2 ) );
  XOR \ADD_/FAINST[9].FA_/U1  ( .A(a[9]), .B(\ADD_/c[9] ), .Z(
        \ADD_/FAINST[9].FA_/n1 ) );
  XOR \ADD_/FAINST[8].FA_/U5  ( .A(\ADD_/FAINST[8].FA_/n3 ), .B(\ADD_/c[8] ), 
        .Z(\ADD_/c[9] ) );
  XOR \ADD_/FAINST[8].FA_/U4  ( .A(\ADD_/FAINST[8].FA_/n1 ), .B(b[8]), .Z(c[8]) );
  AND \ADD_/FAINST[8].FA_/U3  ( .A(\ADD_/FAINST[8].FA_/n1 ), .B(
        \ADD_/FAINST[8].FA_/n2 ), .Z(\ADD_/FAINST[8].FA_/n3 ) );
  XOR \ADD_/FAINST[8].FA_/U2  ( .A(b[8]), .B(\ADD_/c[8] ), .Z(
        \ADD_/FAINST[8].FA_/n2 ) );
  XOR \ADD_/FAINST[8].FA_/U1  ( .A(a[8]), .B(\ADD_/c[8] ), .Z(
        \ADD_/FAINST[8].FA_/n1 ) );
  XOR \ADD_/FAINST[7].FA_/U5  ( .A(\ADD_/FAINST[7].FA_/n3 ), .B(\ADD_/c[7] ), 
        .Z(\ADD_/c[8] ) );
  XOR \ADD_/FAINST[7].FA_/U4  ( .A(\ADD_/FAINST[7].FA_/n1 ), .B(b[7]), .Z(c[7]) );
  AND \ADD_/FAINST[7].FA_/U3  ( .A(\ADD_/FAINST[7].FA_/n1 ), .B(
        \ADD_/FAINST[7].FA_/n2 ), .Z(\ADD_/FAINST[7].FA_/n3 ) );
  XOR \ADD_/FAINST[7].FA_/U2  ( .A(b[7]), .B(\ADD_/c[7] ), .Z(
        \ADD_/FAINST[7].FA_/n2 ) );
  XOR \ADD_/FAINST[7].FA_/U1  ( .A(a[7]), .B(\ADD_/c[7] ), .Z(
        \ADD_/FAINST[7].FA_/n1 ) );
  XOR \ADD_/FAINST[6].FA_/U5  ( .A(\ADD_/FAINST[6].FA_/n3 ), .B(\ADD_/c[6] ), 
        .Z(\ADD_/c[7] ) );
  XOR \ADD_/FAINST[6].FA_/U4  ( .A(\ADD_/FAINST[6].FA_/n1 ), .B(b[6]), .Z(c[6]) );
  AND \ADD_/FAINST[6].FA_/U3  ( .A(\ADD_/FAINST[6].FA_/n1 ), .B(
        \ADD_/FAINST[6].FA_/n2 ), .Z(\ADD_/FAINST[6].FA_/n3 ) );
  XOR \ADD_/FAINST[6].FA_/U2  ( .A(b[6]), .B(\ADD_/c[6] ), .Z(
        \ADD_/FAINST[6].FA_/n2 ) );
  XOR \ADD_/FAINST[6].FA_/U1  ( .A(a[6]), .B(\ADD_/c[6] ), .Z(
        \ADD_/FAINST[6].FA_/n1 ) );
  XOR \ADD_/FAINST[5].FA_/U5  ( .A(\ADD_/FAINST[5].FA_/n3 ), .B(\ADD_/c[5] ), 
        .Z(\ADD_/c[6] ) );
  XOR \ADD_/FAINST[5].FA_/U4  ( .A(\ADD_/FAINST[5].FA_/n1 ), .B(b[5]), .Z(c[5]) );
  AND \ADD_/FAINST[5].FA_/U3  ( .A(\ADD_/FAINST[5].FA_/n1 ), .B(
        \ADD_/FAINST[5].FA_/n2 ), .Z(\ADD_/FAINST[5].FA_/n3 ) );
  XOR \ADD_/FAINST[5].FA_/U2  ( .A(b[5]), .B(\ADD_/c[5] ), .Z(
        \ADD_/FAINST[5].FA_/n2 ) );
  XOR \ADD_/FAINST[5].FA_/U1  ( .A(a[5]), .B(\ADD_/c[5] ), .Z(
        \ADD_/FAINST[5].FA_/n1 ) );
  XOR \ADD_/FAINST[4].FA_/U5  ( .A(\ADD_/FAINST[4].FA_/n3 ), .B(\ADD_/c[4] ), 
        .Z(\ADD_/c[5] ) );
  XOR \ADD_/FAINST[4].FA_/U4  ( .A(\ADD_/FAINST[4].FA_/n1 ), .B(b[4]), .Z(c[4]) );
  AND \ADD_/FAINST[4].FA_/U3  ( .A(\ADD_/FAINST[4].FA_/n1 ), .B(
        \ADD_/FAINST[4].FA_/n2 ), .Z(\ADD_/FAINST[4].FA_/n3 ) );
  XOR \ADD_/FAINST[4].FA_/U2  ( .A(b[4]), .B(\ADD_/c[4] ), .Z(
        \ADD_/FAINST[4].FA_/n2 ) );
  XOR \ADD_/FAINST[4].FA_/U1  ( .A(a[4]), .B(\ADD_/c[4] ), .Z(
        \ADD_/FAINST[4].FA_/n1 ) );
  XOR \ADD_/FAINST[3].FA_/U5  ( .A(\ADD_/FAINST[3].FA_/n3 ), .B(\ADD_/c[3] ), 
        .Z(\ADD_/c[4] ) );
  XOR \ADD_/FAINST[3].FA_/U4  ( .A(\ADD_/FAINST[3].FA_/n1 ), .B(b[3]), .Z(c[3]) );
  AND \ADD_/FAINST[3].FA_/U3  ( .A(\ADD_/FAINST[3].FA_/n1 ), .B(
        \ADD_/FAINST[3].FA_/n2 ), .Z(\ADD_/FAINST[3].FA_/n3 ) );
  XOR \ADD_/FAINST[3].FA_/U2  ( .A(b[3]), .B(\ADD_/c[3] ), .Z(
        \ADD_/FAINST[3].FA_/n2 ) );
  XOR \ADD_/FAINST[3].FA_/U1  ( .A(a[3]), .B(\ADD_/c[3] ), .Z(
        \ADD_/FAINST[3].FA_/n1 ) );
  XOR \ADD_/FAINST[2].FA_/U5  ( .A(\ADD_/FAINST[2].FA_/n3 ), .B(\ADD_/c[2] ), 
        .Z(\ADD_/c[3] ) );
  XOR \ADD_/FAINST[2].FA_/U4  ( .A(\ADD_/FAINST[2].FA_/n1 ), .B(b[2]), .Z(c[2]) );
  AND \ADD_/FAINST[2].FA_/U3  ( .A(\ADD_/FAINST[2].FA_/n1 ), .B(
        \ADD_/FAINST[2].FA_/n2 ), .Z(\ADD_/FAINST[2].FA_/n3 ) );
  XOR \ADD_/FAINST[2].FA_/U2  ( .A(b[2]), .B(\ADD_/c[2] ), .Z(
        \ADD_/FAINST[2].FA_/n2 ) );
  XOR \ADD_/FAINST[2].FA_/U1  ( .A(a[2]), .B(\ADD_/c[2] ), .Z(
        \ADD_/FAINST[2].FA_/n1 ) );
  XOR \ADD_/FAINST[1].FA_/U5  ( .A(\ADD_/FAINST[1].FA_/n3 ), .B(\ADD_/c[1] ), 
        .Z(\ADD_/c[2] ) );
  XOR \ADD_/FAINST[1].FA_/U4  ( .A(\ADD_/FAINST[1].FA_/n1 ), .B(b[1]), .Z(c[1]) );
  AND \ADD_/FAINST[1].FA_/U3  ( .A(\ADD_/FAINST[1].FA_/n1 ), .B(
        \ADD_/FAINST[1].FA_/n2 ), .Z(\ADD_/FAINST[1].FA_/n3 ) );
  XOR \ADD_/FAINST[1].FA_/U2  ( .A(b[1]), .B(\ADD_/c[1] ), .Z(
        \ADD_/FAINST[1].FA_/n2 ) );
  XOR \ADD_/FAINST[1].FA_/U1  ( .A(a[1]), .B(\ADD_/c[1] ), .Z(
        \ADD_/FAINST[1].FA_/n1 ) );
endmodule

